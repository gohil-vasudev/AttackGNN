module add_mul_mix_8_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, c_0_, c_1_, c_2_, c_3_, 
        c_4_, c_5_, c_6_, c_7_, d_0_, d_1_, d_2_, d_3_, d_4_, d_5_, d_6_, d_7_, 
        Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_, 
        Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_, 
        Result_12_, Result_13_, Result_14_, Result_15_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_,
         b_4_, b_5_, b_6_, b_7_, c_0_, c_1_, c_2_, c_3_, c_4_, c_5_, c_6_,
         c_7_, d_0_, d_1_, d_2_, d_3_, d_4_, d_5_, d_6_, d_7_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_;
  wire   n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957;

  XNOR2_X1 U492 ( .A(n477), .B(n478), .ZN(Result_9_) );
  XOR2_X1 U493 ( .A(n479), .B(n480), .Z(n478) );
  XNOR2_X1 U494 ( .A(n481), .B(n482), .ZN(Result_8_) );
  XOR2_X1 U495 ( .A(n483), .B(n484), .Z(n482) );
  XOR2_X1 U496 ( .A(n485), .B(n486), .Z(Result_7_) );
  AND2_X1 U497 ( .A1(n487), .A2(n488), .ZN(Result_6_) );
  INV_X1 U498 ( .A(n489), .ZN(n487) );
  AND2_X1 U499 ( .A1(n490), .A2(n491), .ZN(n489) );
  OR2_X1 U500 ( .A1(n485), .A2(n486), .ZN(n490) );
  XOR2_X1 U501 ( .A(n488), .B(n492), .Z(Result_5_) );
  OR2_X1 U502 ( .A1(n493), .A2(n494), .ZN(n492) );
  INV_X1 U503 ( .A(n495), .ZN(n494) );
  AND2_X1 U504 ( .A1(n496), .A2(n497), .ZN(n493) );
  OR2_X1 U505 ( .A1(n498), .A2(n499), .ZN(n496) );
  XNOR2_X1 U506 ( .A(n500), .B(n501), .ZN(Result_4_) );
  XOR2_X1 U507 ( .A(n502), .B(n503), .Z(Result_3_) );
  AND2_X1 U508 ( .A1(n504), .A2(n505), .ZN(n503) );
  OR2_X1 U509 ( .A1(n506), .A2(n507), .ZN(n505) );
  AND2_X1 U510 ( .A1(n508), .A2(n509), .ZN(n507) );
  INV_X1 U511 ( .A(n510), .ZN(n504) );
  XOR2_X1 U512 ( .A(n511), .B(n512), .Z(Result_2_) );
  XOR2_X1 U513 ( .A(n513), .B(n514), .Z(Result_1_) );
  AND2_X1 U514 ( .A1(n515), .A2(n516), .ZN(n514) );
  OR2_X1 U515 ( .A1(n517), .A2(n518), .ZN(n516) );
  AND2_X1 U516 ( .A1(n519), .A2(n520), .ZN(n517) );
  INV_X1 U517 ( .A(n521), .ZN(n515) );
  INV_X1 U518 ( .A(n522), .ZN(Result_15_) );
  XOR2_X1 U519 ( .A(n523), .B(n524), .Z(Result_14_) );
  OR2_X1 U520 ( .A1(n525), .A2(n526), .ZN(n524) );
  XNOR2_X1 U521 ( .A(n527), .B(n528), .ZN(Result_13_) );
  XOR2_X1 U522 ( .A(n529), .B(n530), .Z(n528) );
  XOR2_X1 U523 ( .A(n531), .B(n532), .Z(Result_12_) );
  XNOR2_X1 U524 ( .A(n533), .B(n534), .ZN(n532) );
  XNOR2_X1 U525 ( .A(n535), .B(n536), .ZN(Result_11_) );
  XOR2_X1 U526 ( .A(n537), .B(n538), .Z(n536) );
  XNOR2_X1 U527 ( .A(n539), .B(n540), .ZN(Result_10_) );
  XOR2_X1 U528 ( .A(n541), .B(n542), .Z(n540) );
  OR3_X1 U529 ( .A1(n521), .A2(n543), .A3(n544), .ZN(Result_0_) );
  INV_X1 U530 ( .A(n545), .ZN(n544) );
  OR2_X1 U531 ( .A1(n546), .A2(n547), .ZN(n545) );
  AND2_X1 U532 ( .A1(n513), .A2(n518), .ZN(n543) );
  AND2_X1 U533 ( .A1(n511), .A2(n512), .ZN(n513) );
  XNOR2_X1 U534 ( .A(n520), .B(n548), .ZN(n512) );
  OR2_X1 U535 ( .A1(n549), .A2(n550), .ZN(n511) );
  OR2_X1 U536 ( .A1(n551), .A2(n510), .ZN(n549) );
  AND3_X1 U537 ( .A1(n509), .A2(n508), .A3(n506), .ZN(n510) );
  INV_X1 U538 ( .A(n552), .ZN(n508) );
  AND2_X1 U539 ( .A1(n502), .A2(n506), .ZN(n551) );
  INV_X1 U540 ( .A(n553), .ZN(n506) );
  OR2_X1 U541 ( .A1(n554), .A2(n550), .ZN(n553) );
  INV_X1 U542 ( .A(n555), .ZN(n550) );
  OR2_X1 U543 ( .A1(n556), .A2(n557), .ZN(n555) );
  AND2_X1 U544 ( .A1(n556), .A2(n557), .ZN(n554) );
  OR2_X1 U545 ( .A1(n558), .A2(n559), .ZN(n557) );
  AND2_X1 U546 ( .A1(n560), .A2(n561), .ZN(n559) );
  AND2_X1 U547 ( .A1(n562), .A2(n563), .ZN(n558) );
  OR2_X1 U548 ( .A1(n561), .A2(n560), .ZN(n563) );
  XOR2_X1 U549 ( .A(n564), .B(n565), .Z(n556) );
  XOR2_X1 U550 ( .A(n566), .B(n567), .Z(n565) );
  AND2_X1 U551 ( .A1(n568), .A2(n501), .ZN(n502) );
  XNOR2_X1 U552 ( .A(n509), .B(n552), .ZN(n501) );
  OR2_X1 U553 ( .A1(n569), .A2(n570), .ZN(n552) );
  AND2_X1 U554 ( .A1(n571), .A2(n572), .ZN(n570) );
  AND2_X1 U555 ( .A1(n573), .A2(n574), .ZN(n569) );
  OR2_X1 U556 ( .A1(n572), .A2(n571), .ZN(n574) );
  XOR2_X1 U557 ( .A(n575), .B(n562), .Z(n509) );
  XOR2_X1 U558 ( .A(n576), .B(n577), .Z(n562) );
  XOR2_X1 U559 ( .A(n578), .B(n579), .Z(n577) );
  XNOR2_X1 U560 ( .A(n561), .B(n560), .ZN(n575) );
  OR2_X1 U561 ( .A1(n580), .A2(n581), .ZN(n560) );
  AND2_X1 U562 ( .A1(n582), .A2(n583), .ZN(n581) );
  AND2_X1 U563 ( .A1(n584), .A2(n585), .ZN(n580) );
  OR2_X1 U564 ( .A1(n583), .A2(n582), .ZN(n585) );
  OR2_X1 U565 ( .A1(n586), .A2(n547), .ZN(n561) );
  INV_X1 U566 ( .A(n500), .ZN(n568) );
  AND2_X1 U567 ( .A1(n587), .A2(n588), .ZN(n500) );
  AND2_X1 U568 ( .A1(n589), .A2(n495), .ZN(n587) );
  OR3_X1 U569 ( .A1(n499), .A2(n498), .A3(n497), .ZN(n495) );
  OR2_X1 U570 ( .A1(n488), .A2(n497), .ZN(n589) );
  OR2_X1 U571 ( .A1(n590), .A2(n591), .ZN(n497) );
  INV_X1 U572 ( .A(n588), .ZN(n591) );
  OR2_X1 U573 ( .A1(n592), .A2(n593), .ZN(n588) );
  AND2_X1 U574 ( .A1(n592), .A2(n593), .ZN(n590) );
  OR2_X1 U575 ( .A1(n594), .A2(n595), .ZN(n593) );
  AND2_X1 U576 ( .A1(n596), .A2(n597), .ZN(n595) );
  AND2_X1 U577 ( .A1(n598), .A2(n599), .ZN(n594) );
  OR2_X1 U578 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U579 ( .A(n573), .B(n600), .Z(n592) );
  XOR2_X1 U580 ( .A(n572), .B(n571), .Z(n600) );
  OR2_X1 U581 ( .A1(n601), .A2(n547), .ZN(n571) );
  OR2_X1 U582 ( .A1(n602), .A2(n603), .ZN(n572) );
  AND2_X1 U583 ( .A1(n604), .A2(n605), .ZN(n603) );
  AND2_X1 U584 ( .A1(n606), .A2(n607), .ZN(n602) );
  OR2_X1 U585 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U586 ( .A(n608), .B(n584), .ZN(n573) );
  XNOR2_X1 U587 ( .A(n609), .B(n610), .ZN(n584) );
  XNOR2_X1 U588 ( .A(n611), .B(n612), .ZN(n609) );
  XNOR2_X1 U589 ( .A(n583), .B(n582), .ZN(n608) );
  OR2_X1 U590 ( .A1(n613), .A2(n614), .ZN(n582) );
  AND2_X1 U591 ( .A1(n615), .A2(n616), .ZN(n614) );
  AND2_X1 U592 ( .A1(n617), .A2(n618), .ZN(n613) );
  OR2_X1 U593 ( .A1(n616), .A2(n615), .ZN(n618) );
  OR2_X1 U594 ( .A1(n586), .A2(n619), .ZN(n583) );
  OR3_X1 U595 ( .A1(n486), .A2(n485), .A3(n491), .ZN(n488) );
  XNOR2_X1 U596 ( .A(n498), .B(n499), .ZN(n491) );
  OR2_X1 U597 ( .A1(n620), .A2(n621), .ZN(n499) );
  AND2_X1 U598 ( .A1(n622), .A2(n623), .ZN(n621) );
  AND2_X1 U599 ( .A1(n624), .A2(n625), .ZN(n620) );
  OR2_X1 U600 ( .A1(n623), .A2(n622), .ZN(n625) );
  XNOR2_X1 U601 ( .A(n626), .B(n596), .ZN(n498) );
  XNOR2_X1 U602 ( .A(n627), .B(n604), .ZN(n596) );
  XNOR2_X1 U603 ( .A(n628), .B(n617), .ZN(n604) );
  XNOR2_X1 U604 ( .A(n629), .B(n630), .ZN(n617) );
  XNOR2_X1 U605 ( .A(n631), .B(n632), .ZN(n629) );
  XNOR2_X1 U606 ( .A(n616), .B(n615), .ZN(n628) );
  OR2_X1 U607 ( .A1(n633), .A2(n634), .ZN(n615) );
  AND2_X1 U608 ( .A1(n635), .A2(n636), .ZN(n634) );
  AND2_X1 U609 ( .A1(n637), .A2(n638), .ZN(n633) );
  OR2_X1 U610 ( .A1(n636), .A2(n635), .ZN(n638) );
  OR2_X1 U611 ( .A1(n586), .A2(n639), .ZN(n616) );
  XNOR2_X1 U612 ( .A(n607), .B(n605), .ZN(n627) );
  OR2_X1 U613 ( .A1(n601), .A2(n619), .ZN(n605) );
  OR2_X1 U614 ( .A1(n640), .A2(n641), .ZN(n607) );
  AND2_X1 U615 ( .A1(n642), .A2(n643), .ZN(n641) );
  AND2_X1 U616 ( .A1(n644), .A2(n645), .ZN(n640) );
  OR2_X1 U617 ( .A1(n643), .A2(n642), .ZN(n645) );
  XNOR2_X1 U618 ( .A(n599), .B(n597), .ZN(n626) );
  OR2_X1 U619 ( .A1(n646), .A2(n547), .ZN(n597) );
  OR2_X1 U620 ( .A1(n647), .A2(n648), .ZN(n599) );
  AND2_X1 U621 ( .A1(n649), .A2(n650), .ZN(n648) );
  AND2_X1 U622 ( .A1(n651), .A2(n652), .ZN(n647) );
  OR2_X1 U623 ( .A1(n650), .A2(n649), .ZN(n652) );
  OR2_X1 U624 ( .A1(n653), .A2(n654), .ZN(n485) );
  AND2_X1 U625 ( .A1(n484), .A2(n483), .ZN(n654) );
  AND2_X1 U626 ( .A1(n481), .A2(n655), .ZN(n653) );
  OR2_X1 U627 ( .A1(n483), .A2(n484), .ZN(n655) );
  OR2_X1 U628 ( .A1(n525), .A2(n547), .ZN(n484) );
  OR2_X1 U629 ( .A1(n656), .A2(n657), .ZN(n483) );
  AND2_X1 U630 ( .A1(n480), .A2(n479), .ZN(n657) );
  AND2_X1 U631 ( .A1(n477), .A2(n658), .ZN(n656) );
  OR2_X1 U632 ( .A1(n479), .A2(n480), .ZN(n658) );
  OR2_X1 U633 ( .A1(n619), .A2(n525), .ZN(n480) );
  OR2_X1 U634 ( .A1(n659), .A2(n660), .ZN(n479) );
  AND2_X1 U635 ( .A1(n542), .A2(n541), .ZN(n660) );
  AND2_X1 U636 ( .A1(n539), .A2(n661), .ZN(n659) );
  OR2_X1 U637 ( .A1(n542), .A2(n541), .ZN(n661) );
  OR2_X1 U638 ( .A1(n662), .A2(n663), .ZN(n541) );
  AND2_X1 U639 ( .A1(n538), .A2(n537), .ZN(n663) );
  AND2_X1 U640 ( .A1(n535), .A2(n664), .ZN(n662) );
  OR2_X1 U641 ( .A1(n538), .A2(n537), .ZN(n664) );
  OR2_X1 U642 ( .A1(n665), .A2(n666), .ZN(n537) );
  AND2_X1 U643 ( .A1(n533), .A2(n534), .ZN(n666) );
  AND2_X1 U644 ( .A1(n531), .A2(n667), .ZN(n665) );
  OR2_X1 U645 ( .A1(n533), .A2(n534), .ZN(n667) );
  OR2_X1 U646 ( .A1(n668), .A2(n669), .ZN(n534) );
  AND2_X1 U647 ( .A1(n530), .A2(n529), .ZN(n669) );
  AND2_X1 U648 ( .A1(n527), .A2(n670), .ZN(n668) );
  OR2_X1 U649 ( .A1(n530), .A2(n529), .ZN(n670) );
  OR2_X1 U650 ( .A1(n671), .A2(n525), .ZN(n529) );
  OR2_X1 U651 ( .A1(n672), .A2(n522), .ZN(n530) );
  OR2_X1 U652 ( .A1(n673), .A2(n525), .ZN(n522) );
  XNOR2_X1 U653 ( .A(n672), .B(n674), .ZN(n527) );
  OR2_X1 U654 ( .A1(n646), .A2(n673), .ZN(n674) );
  OR2_X1 U655 ( .A1(n526), .A2(n675), .ZN(n672) );
  OR2_X1 U656 ( .A1(n676), .A2(n525), .ZN(n533) );
  XNOR2_X1 U657 ( .A(n677), .B(n678), .ZN(n531) );
  XNOR2_X1 U658 ( .A(n679), .B(n680), .ZN(n677) );
  OR2_X1 U659 ( .A1(n681), .A2(n525), .ZN(n538) );
  XOR2_X1 U660 ( .A(n682), .B(n683), .Z(n535) );
  XOR2_X1 U661 ( .A(n684), .B(n685), .Z(n683) );
  OR2_X1 U662 ( .A1(n639), .A2(n525), .ZN(n542) );
  OR2_X1 U663 ( .A1(n686), .A2(n687), .ZN(n525) );
  INV_X1 U664 ( .A(n688), .ZN(n686) );
  OR2_X1 U665 ( .A1(c_7_), .A2(d_7_), .ZN(n688) );
  XOR2_X1 U666 ( .A(n689), .B(n690), .Z(n539) );
  XOR2_X1 U667 ( .A(n691), .B(n692), .Z(n690) );
  XOR2_X1 U668 ( .A(n693), .B(n694), .Z(n477) );
  XOR2_X1 U669 ( .A(n695), .B(n696), .Z(n694) );
  XOR2_X1 U670 ( .A(n697), .B(n698), .Z(n481) );
  XOR2_X1 U671 ( .A(n699), .B(n700), .Z(n698) );
  XOR2_X1 U672 ( .A(n624), .B(n701), .Z(n486) );
  XOR2_X1 U673 ( .A(n623), .B(n622), .Z(n701) );
  OR2_X1 U674 ( .A1(n675), .A2(n547), .ZN(n622) );
  OR2_X1 U675 ( .A1(n702), .A2(n703), .ZN(n623) );
  AND2_X1 U676 ( .A1(n700), .A2(n699), .ZN(n703) );
  AND2_X1 U677 ( .A1(n697), .A2(n704), .ZN(n702) );
  OR2_X1 U678 ( .A1(n699), .A2(n700), .ZN(n704) );
  OR2_X1 U679 ( .A1(n675), .A2(n619), .ZN(n700) );
  OR2_X1 U680 ( .A1(n705), .A2(n706), .ZN(n699) );
  AND2_X1 U681 ( .A1(n696), .A2(n695), .ZN(n706) );
  AND2_X1 U682 ( .A1(n693), .A2(n707), .ZN(n705) );
  OR2_X1 U683 ( .A1(n695), .A2(n696), .ZN(n707) );
  OR2_X1 U684 ( .A1(n675), .A2(n639), .ZN(n696) );
  OR2_X1 U685 ( .A1(n708), .A2(n709), .ZN(n695) );
  AND2_X1 U686 ( .A1(n692), .A2(n691), .ZN(n709) );
  AND2_X1 U687 ( .A1(n689), .A2(n710), .ZN(n708) );
  OR2_X1 U688 ( .A1(n692), .A2(n691), .ZN(n710) );
  OR2_X1 U689 ( .A1(n711), .A2(n712), .ZN(n691) );
  AND2_X1 U690 ( .A1(n685), .A2(n684), .ZN(n712) );
  AND2_X1 U691 ( .A1(n682), .A2(n713), .ZN(n711) );
  OR2_X1 U692 ( .A1(n685), .A2(n684), .ZN(n713) );
  OR2_X1 U693 ( .A1(n714), .A2(n715), .ZN(n684) );
  AND2_X1 U694 ( .A1(n678), .A2(n680), .ZN(n715) );
  AND2_X1 U695 ( .A1(n716), .A2(n679), .ZN(n714) );
  OR2_X1 U696 ( .A1(n717), .A2(n718), .ZN(n679) );
  INV_X1 U697 ( .A(n719), .ZN(n718) );
  AND2_X1 U698 ( .A1(n720), .A2(n721), .ZN(n717) );
  OR2_X1 U699 ( .A1(n678), .A2(n680), .ZN(n716) );
  OR2_X1 U700 ( .A1(n721), .A2(n523), .ZN(n680) );
  OR2_X1 U701 ( .A1(n675), .A2(n673), .ZN(n523) );
  OR2_X1 U702 ( .A1(n675), .A2(n671), .ZN(n678) );
  OR2_X1 U703 ( .A1(n676), .A2(n675), .ZN(n685) );
  XNOR2_X1 U704 ( .A(n722), .B(n723), .ZN(n682) );
  XNOR2_X1 U705 ( .A(n724), .B(n719), .ZN(n722) );
  OR2_X1 U706 ( .A1(n681), .A2(n675), .ZN(n692) );
  XNOR2_X1 U707 ( .A(n687), .B(n725), .ZN(n675) );
  XOR2_X1 U708 ( .A(d_6_), .B(c_6_), .Z(n725) );
  XOR2_X1 U709 ( .A(n726), .B(n727), .Z(n689) );
  XOR2_X1 U710 ( .A(n728), .B(n729), .Z(n727) );
  XOR2_X1 U711 ( .A(n730), .B(n731), .Z(n693) );
  XOR2_X1 U712 ( .A(n732), .B(n733), .Z(n731) );
  XOR2_X1 U713 ( .A(n734), .B(n735), .Z(n697) );
  XOR2_X1 U714 ( .A(n736), .B(n737), .Z(n735) );
  XOR2_X1 U715 ( .A(n651), .B(n738), .Z(n624) );
  XOR2_X1 U716 ( .A(n650), .B(n649), .Z(n738) );
  OR2_X1 U717 ( .A1(n619), .A2(n646), .ZN(n649) );
  OR2_X1 U718 ( .A1(n739), .A2(n740), .ZN(n650) );
  AND2_X1 U719 ( .A1(n737), .A2(n736), .ZN(n740) );
  AND2_X1 U720 ( .A1(n734), .A2(n741), .ZN(n739) );
  OR2_X1 U721 ( .A1(n736), .A2(n737), .ZN(n741) );
  OR2_X1 U722 ( .A1(n639), .A2(n646), .ZN(n737) );
  OR2_X1 U723 ( .A1(n742), .A2(n743), .ZN(n736) );
  AND2_X1 U724 ( .A1(n733), .A2(n732), .ZN(n743) );
  AND2_X1 U725 ( .A1(n730), .A2(n744), .ZN(n742) );
  OR2_X1 U726 ( .A1(n732), .A2(n733), .ZN(n744) );
  OR2_X1 U727 ( .A1(n681), .A2(n646), .ZN(n733) );
  OR2_X1 U728 ( .A1(n745), .A2(n746), .ZN(n732) );
  AND2_X1 U729 ( .A1(n729), .A2(n728), .ZN(n746) );
  AND2_X1 U730 ( .A1(n726), .A2(n747), .ZN(n745) );
  OR2_X1 U731 ( .A1(n729), .A2(n728), .ZN(n747) );
  OR2_X1 U732 ( .A1(n748), .A2(n749), .ZN(n728) );
  AND2_X1 U733 ( .A1(n723), .A2(n719), .ZN(n749) );
  AND2_X1 U734 ( .A1(n750), .A2(n724), .ZN(n748) );
  OR2_X1 U735 ( .A1(n751), .A2(n752), .ZN(n724) );
  INV_X1 U736 ( .A(n753), .ZN(n752) );
  AND2_X1 U737 ( .A1(n754), .A2(n755), .ZN(n751) );
  OR2_X1 U738 ( .A1(n723), .A2(n719), .ZN(n750) );
  OR2_X1 U739 ( .A1(n720), .A2(n721), .ZN(n719) );
  OR2_X1 U740 ( .A1(n526), .A2(n646), .ZN(n721) );
  OR2_X1 U741 ( .A1(n601), .A2(n673), .ZN(n720) );
  OR2_X1 U742 ( .A1(n671), .A2(n646), .ZN(n723) );
  OR2_X1 U743 ( .A1(n676), .A2(n646), .ZN(n729) );
  XOR2_X1 U744 ( .A(n756), .B(n757), .Z(n646) );
  XNOR2_X1 U745 ( .A(n758), .B(c_5_), .ZN(n757) );
  XNOR2_X1 U746 ( .A(n759), .B(n760), .ZN(n726) );
  XNOR2_X1 U747 ( .A(n761), .B(n753), .ZN(n759) );
  XOR2_X1 U748 ( .A(n762), .B(n763), .Z(n730) );
  XOR2_X1 U749 ( .A(n764), .B(n765), .Z(n763) );
  XOR2_X1 U750 ( .A(n766), .B(n767), .Z(n734) );
  XOR2_X1 U751 ( .A(n768), .B(n769), .Z(n767) );
  XOR2_X1 U752 ( .A(n644), .B(n770), .Z(n651) );
  XOR2_X1 U753 ( .A(n643), .B(n642), .Z(n770) );
  OR2_X1 U754 ( .A1(n601), .A2(n639), .ZN(n642) );
  OR2_X1 U755 ( .A1(n771), .A2(n772), .ZN(n643) );
  AND2_X1 U756 ( .A1(n769), .A2(n768), .ZN(n772) );
  AND2_X1 U757 ( .A1(n766), .A2(n773), .ZN(n771) );
  OR2_X1 U758 ( .A1(n768), .A2(n769), .ZN(n773) );
  OR2_X1 U759 ( .A1(n601), .A2(n681), .ZN(n769) );
  OR2_X1 U760 ( .A1(n774), .A2(n775), .ZN(n768) );
  AND2_X1 U761 ( .A1(n765), .A2(n764), .ZN(n775) );
  AND2_X1 U762 ( .A1(n762), .A2(n776), .ZN(n774) );
  OR2_X1 U763 ( .A1(n764), .A2(n765), .ZN(n776) );
  OR2_X1 U764 ( .A1(n601), .A2(n676), .ZN(n765) );
  OR2_X1 U765 ( .A1(n777), .A2(n778), .ZN(n764) );
  AND2_X1 U766 ( .A1(n760), .A2(n753), .ZN(n778) );
  AND2_X1 U767 ( .A1(n779), .A2(n761), .ZN(n777) );
  OR2_X1 U768 ( .A1(n780), .A2(n781), .ZN(n761) );
  INV_X1 U769 ( .A(n782), .ZN(n781) );
  AND2_X1 U770 ( .A1(n783), .A2(n784), .ZN(n780) );
  OR2_X1 U771 ( .A1(n760), .A2(n753), .ZN(n779) );
  OR2_X1 U772 ( .A1(n754), .A2(n755), .ZN(n753) );
  OR2_X1 U773 ( .A1(n586), .A2(n673), .ZN(n755) );
  OR2_X1 U774 ( .A1(n526), .A2(n601), .ZN(n754) );
  OR2_X1 U775 ( .A1(n601), .A2(n671), .ZN(n760) );
  XNOR2_X1 U776 ( .A(n785), .B(n786), .ZN(n601) );
  XNOR2_X1 U777 ( .A(c_4_), .B(d_4_), .ZN(n785) );
  XNOR2_X1 U778 ( .A(n787), .B(n782), .ZN(n762) );
  XNOR2_X1 U779 ( .A(n788), .B(n789), .ZN(n787) );
  XOR2_X1 U780 ( .A(n790), .B(n791), .Z(n766) );
  XOR2_X1 U781 ( .A(n792), .B(n793), .Z(n791) );
  XNOR2_X1 U782 ( .A(n794), .B(n637), .ZN(n644) );
  XNOR2_X1 U783 ( .A(n795), .B(n796), .ZN(n637) );
  XNOR2_X1 U784 ( .A(n797), .B(n798), .ZN(n795) );
  XNOR2_X1 U785 ( .A(n635), .B(n636), .ZN(n794) );
  OR2_X1 U786 ( .A1(n586), .A2(n681), .ZN(n636) );
  OR2_X1 U787 ( .A1(n799), .A2(n800), .ZN(n635) );
  AND2_X1 U788 ( .A1(n793), .A2(n792), .ZN(n800) );
  AND2_X1 U789 ( .A1(n790), .A2(n801), .ZN(n799) );
  OR2_X1 U790 ( .A1(n792), .A2(n793), .ZN(n801) );
  OR2_X1 U791 ( .A1(n802), .A2(n803), .ZN(n793) );
  AND2_X1 U792 ( .A1(n782), .A2(n789), .ZN(n803) );
  AND2_X1 U793 ( .A1(n804), .A2(n788), .ZN(n802) );
  OR2_X1 U794 ( .A1(n805), .A2(n806), .ZN(n788) );
  INV_X1 U795 ( .A(n807), .ZN(n806) );
  AND2_X1 U796 ( .A1(n808), .A2(n809), .ZN(n805) );
  OR2_X1 U797 ( .A1(n810), .A2(n673), .ZN(n809) );
  OR2_X1 U798 ( .A1(n811), .A2(n526), .ZN(n808) );
  OR2_X1 U799 ( .A1(n789), .A2(n782), .ZN(n804) );
  OR2_X1 U800 ( .A1(n783), .A2(n784), .ZN(n782) );
  OR2_X1 U801 ( .A1(n526), .A2(n586), .ZN(n783) );
  OR2_X1 U802 ( .A1(n586), .A2(n671), .ZN(n789) );
  OR2_X1 U803 ( .A1(n586), .A2(n676), .ZN(n792) );
  XNOR2_X1 U804 ( .A(n812), .B(n813), .ZN(n586) );
  XNOR2_X1 U805 ( .A(c_3_), .B(d_3_), .ZN(n812) );
  XNOR2_X1 U806 ( .A(n814), .B(n815), .ZN(n790) );
  XNOR2_X1 U807 ( .A(n816), .B(n807), .ZN(n814) );
  AND3_X1 U808 ( .A1(n520), .A2(n518), .A3(n519), .ZN(n521) );
  INV_X1 U809 ( .A(n548), .ZN(n519) );
  OR2_X1 U810 ( .A1(n817), .A2(n818), .ZN(n548) );
  AND2_X1 U811 ( .A1(n567), .A2(n566), .ZN(n818) );
  AND2_X1 U812 ( .A1(n564), .A2(n819), .ZN(n817) );
  OR2_X1 U813 ( .A1(n566), .A2(n567), .ZN(n819) );
  OR2_X1 U814 ( .A1(n811), .A2(n547), .ZN(n567) );
  OR2_X1 U815 ( .A1(n820), .A2(n821), .ZN(n566) );
  AND2_X1 U816 ( .A1(n579), .A2(n578), .ZN(n821) );
  AND2_X1 U817 ( .A1(n576), .A2(n822), .ZN(n820) );
  OR2_X1 U818 ( .A1(n578), .A2(n579), .ZN(n822) );
  OR2_X1 U819 ( .A1(n811), .A2(n619), .ZN(n579) );
  OR2_X1 U820 ( .A1(n823), .A2(n824), .ZN(n578) );
  AND2_X1 U821 ( .A1(n612), .A2(n611), .ZN(n824) );
  AND2_X1 U822 ( .A1(n610), .A2(n825), .ZN(n823) );
  OR2_X1 U823 ( .A1(n611), .A2(n612), .ZN(n825) );
  OR2_X1 U824 ( .A1(n826), .A2(n827), .ZN(n612) );
  AND2_X1 U825 ( .A1(n632), .A2(n631), .ZN(n827) );
  AND2_X1 U826 ( .A1(n630), .A2(n828), .ZN(n826) );
  OR2_X1 U827 ( .A1(n631), .A2(n632), .ZN(n828) );
  OR2_X1 U828 ( .A1(n829), .A2(n830), .ZN(n632) );
  AND2_X1 U829 ( .A1(n798), .A2(n797), .ZN(n830) );
  AND2_X1 U830 ( .A1(n796), .A2(n831), .ZN(n829) );
  OR2_X1 U831 ( .A1(n797), .A2(n798), .ZN(n831) );
  OR2_X1 U832 ( .A1(n811), .A2(n676), .ZN(n798) );
  OR2_X1 U833 ( .A1(n832), .A2(n833), .ZN(n797) );
  AND2_X1 U834 ( .A1(n815), .A2(n807), .ZN(n833) );
  AND2_X1 U835 ( .A1(n834), .A2(n816), .ZN(n832) );
  OR2_X1 U836 ( .A1(n835), .A2(n836), .ZN(n816) );
  AND2_X1 U837 ( .A1(n837), .A2(n838), .ZN(n835) );
  OR2_X1 U838 ( .A1(n807), .A2(n815), .ZN(n834) );
  OR2_X1 U839 ( .A1(n811), .A2(n671), .ZN(n815) );
  OR2_X1 U840 ( .A1(n784), .A2(n838), .ZN(n807) );
  OR2_X1 U841 ( .A1(n811), .A2(n673), .ZN(n784) );
  XNOR2_X1 U842 ( .A(n839), .B(n840), .ZN(n796) );
  OR2_X1 U843 ( .A1(n836), .A2(n841), .ZN(n839) );
  INV_X1 U844 ( .A(n842), .ZN(n836) );
  OR2_X1 U845 ( .A1(n811), .A2(n681), .ZN(n631) );
  XOR2_X1 U846 ( .A(n843), .B(n844), .Z(n630) );
  XOR2_X1 U847 ( .A(n845), .B(n846), .Z(n843) );
  OR2_X1 U848 ( .A1(n811), .A2(n639), .ZN(n611) );
  XNOR2_X1 U849 ( .A(n847), .B(n848), .ZN(n811) );
  XNOR2_X1 U850 ( .A(c_2_), .B(d_2_), .ZN(n847) );
  XOR2_X1 U851 ( .A(n849), .B(n850), .Z(n610) );
  XOR2_X1 U852 ( .A(n851), .B(n852), .Z(n850) );
  XOR2_X1 U853 ( .A(n853), .B(n854), .Z(n576) );
  XOR2_X1 U854 ( .A(n855), .B(n856), .Z(n854) );
  XOR2_X1 U855 ( .A(n857), .B(n858), .Z(n564) );
  XOR2_X1 U856 ( .A(n859), .B(n860), .Z(n858) );
  XOR2_X1 U857 ( .A(n861), .B(n546), .Z(n518) );
  OR2_X1 U858 ( .A1(n862), .A2(n863), .ZN(n546) );
  AND2_X1 U859 ( .A1(n864), .A2(n865), .ZN(n863) );
  AND2_X1 U860 ( .A1(n866), .A2(n867), .ZN(n862) );
  OR2_X1 U861 ( .A1(n865), .A2(n864), .ZN(n866) );
  OR2_X1 U862 ( .A1(n868), .A2(n547), .ZN(n861) );
  XNOR2_X1 U863 ( .A(n864), .B(n869), .ZN(n520) );
  XOR2_X1 U864 ( .A(n865), .B(n867), .Z(n869) );
  OR2_X1 U865 ( .A1(n810), .A2(n547), .ZN(n867) );
  XNOR2_X1 U866 ( .A(n870), .B(n871), .ZN(n547) );
  XOR2_X1 U867 ( .A(b_0_), .B(a_0_), .Z(n871) );
  OR2_X1 U868 ( .A1(n872), .A2(n873), .ZN(n870) );
  AND2_X1 U869 ( .A1(n874), .A2(a_1_), .ZN(n873) );
  AND2_X1 U870 ( .A1(b_1_), .A2(n875), .ZN(n872) );
  OR2_X1 U871 ( .A1(n874), .A2(a_1_), .ZN(n875) );
  INV_X1 U872 ( .A(n876), .ZN(n874) );
  OR2_X1 U873 ( .A1(n877), .A2(n878), .ZN(n865) );
  AND2_X1 U874 ( .A1(n857), .A2(n859), .ZN(n878) );
  AND2_X1 U875 ( .A1(n879), .A2(n860), .ZN(n877) );
  OR2_X1 U876 ( .A1(n810), .A2(n619), .ZN(n860) );
  OR2_X1 U877 ( .A1(n859), .A2(n857), .ZN(n879) );
  OR2_X1 U878 ( .A1(n639), .A2(n868), .ZN(n857) );
  OR2_X1 U879 ( .A1(n880), .A2(n881), .ZN(n859) );
  AND2_X1 U880 ( .A1(n853), .A2(n855), .ZN(n881) );
  AND2_X1 U881 ( .A1(n882), .A2(n856), .ZN(n880) );
  OR2_X1 U882 ( .A1(n681), .A2(n868), .ZN(n856) );
  OR2_X1 U883 ( .A1(n855), .A2(n853), .ZN(n882) );
  OR2_X1 U884 ( .A1(n810), .A2(n639), .ZN(n853) );
  XNOR2_X1 U885 ( .A(n883), .B(n884), .ZN(n639) );
  XNOR2_X1 U886 ( .A(a_2_), .B(b_2_), .ZN(n883) );
  OR2_X1 U887 ( .A1(n885), .A2(n886), .ZN(n855) );
  AND2_X1 U888 ( .A1(n849), .A2(n851), .ZN(n886) );
  AND2_X1 U889 ( .A1(n887), .A2(n852), .ZN(n885) );
  OR2_X1 U890 ( .A1(n810), .A2(n681), .ZN(n852) );
  XNOR2_X1 U891 ( .A(n888), .B(n889), .ZN(n681) );
  XNOR2_X1 U892 ( .A(a_3_), .B(b_3_), .ZN(n888) );
  OR2_X1 U893 ( .A1(n851), .A2(n849), .ZN(n887) );
  OR2_X1 U894 ( .A1(n676), .A2(n868), .ZN(n849) );
  OR2_X1 U895 ( .A1(n890), .A2(n891), .ZN(n851) );
  AND2_X1 U896 ( .A1(n844), .A2(n846), .ZN(n891) );
  AND2_X1 U897 ( .A1(n845), .A2(n892), .ZN(n890) );
  OR2_X1 U898 ( .A1(n846), .A2(n844), .ZN(n892) );
  OR2_X1 U899 ( .A1(n671), .A2(n868), .ZN(n844) );
  OR2_X1 U900 ( .A1(n810), .A2(n676), .ZN(n846) );
  XNOR2_X1 U901 ( .A(n893), .B(n894), .ZN(n676) );
  XNOR2_X1 U902 ( .A(a_4_), .B(b_4_), .ZN(n893) );
  AND2_X1 U903 ( .A1(n842), .A2(n895), .ZN(n845) );
  OR2_X1 U904 ( .A1(n840), .A2(n841), .ZN(n895) );
  OR2_X1 U905 ( .A1(n526), .A2(n868), .ZN(n841) );
  OR2_X1 U906 ( .A1(n810), .A2(n671), .ZN(n840) );
  XNOR2_X1 U907 ( .A(n896), .B(n897), .ZN(n671) );
  XNOR2_X1 U908 ( .A(n898), .B(a_5_), .ZN(n897) );
  OR2_X1 U909 ( .A1(n838), .A2(n837), .ZN(n842) );
  OR2_X1 U910 ( .A1(n673), .A2(n868), .ZN(n837) );
  OR2_X1 U911 ( .A1(n899), .A2(n900), .ZN(n673) );
  INV_X1 U912 ( .A(n901), .ZN(n899) );
  OR2_X1 U913 ( .A1(a_7_), .A2(b_7_), .ZN(n901) );
  OR2_X1 U914 ( .A1(n526), .A2(n810), .ZN(n838) );
  XNOR2_X1 U915 ( .A(n902), .B(n903), .ZN(n810) );
  XNOR2_X1 U916 ( .A(c_1_), .B(d_1_), .ZN(n902) );
  XNOR2_X1 U917 ( .A(n900), .B(n904), .ZN(n526) );
  XOR2_X1 U918 ( .A(b_6_), .B(a_6_), .Z(n904) );
  OR2_X1 U919 ( .A1(n619), .A2(n868), .ZN(n864) );
  XNOR2_X1 U920 ( .A(n905), .B(n906), .ZN(n868) );
  XOR2_X1 U921 ( .A(d_0_), .B(c_0_), .Z(n906) );
  OR2_X1 U922 ( .A1(n907), .A2(n908), .ZN(n905) );
  AND2_X1 U923 ( .A1(n909), .A2(c_1_), .ZN(n908) );
  AND2_X1 U924 ( .A1(d_1_), .A2(n910), .ZN(n907) );
  OR2_X1 U925 ( .A1(n909), .A2(c_1_), .ZN(n910) );
  INV_X1 U926 ( .A(n903), .ZN(n909) );
  OR2_X1 U927 ( .A1(n911), .A2(n912), .ZN(n903) );
  AND2_X1 U928 ( .A1(n848), .A2(n913), .ZN(n912) );
  AND2_X1 U929 ( .A1(n914), .A2(n915), .ZN(n911) );
  INV_X1 U930 ( .A(d_2_), .ZN(n915) );
  OR2_X1 U931 ( .A1(n913), .A2(n848), .ZN(n914) );
  OR2_X1 U932 ( .A1(n916), .A2(n917), .ZN(n848) );
  AND2_X1 U933 ( .A1(n813), .A2(n918), .ZN(n917) );
  AND2_X1 U934 ( .A1(n919), .A2(n920), .ZN(n916) );
  INV_X1 U935 ( .A(d_3_), .ZN(n920) );
  OR2_X1 U936 ( .A1(n813), .A2(n918), .ZN(n919) );
  INV_X1 U937 ( .A(c_3_), .ZN(n918) );
  OR2_X1 U938 ( .A1(n921), .A2(n922), .ZN(n813) );
  AND2_X1 U939 ( .A1(n786), .A2(n923), .ZN(n922) );
  AND2_X1 U940 ( .A1(n924), .A2(n925), .ZN(n921) );
  INV_X1 U941 ( .A(d_4_), .ZN(n925) );
  OR2_X1 U942 ( .A1(n786), .A2(n923), .ZN(n924) );
  INV_X1 U943 ( .A(c_4_), .ZN(n923) );
  OR2_X1 U944 ( .A1(n926), .A2(n927), .ZN(n786) );
  AND2_X1 U945 ( .A1(n756), .A2(n928), .ZN(n927) );
  AND2_X1 U946 ( .A1(n929), .A2(n758), .ZN(n926) );
  INV_X1 U947 ( .A(d_5_), .ZN(n758) );
  OR2_X1 U948 ( .A1(n756), .A2(n928), .ZN(n929) );
  INV_X1 U949 ( .A(c_5_), .ZN(n928) );
  INV_X1 U950 ( .A(n930), .ZN(n756) );
  OR2_X1 U951 ( .A1(n931), .A2(n932), .ZN(n930) );
  AND2_X1 U952 ( .A1(c_6_), .A2(n687), .ZN(n932) );
  AND2_X1 U953 ( .A1(d_6_), .A2(n933), .ZN(n931) );
  OR2_X1 U954 ( .A1(n687), .A2(c_6_), .ZN(n933) );
  AND2_X1 U955 ( .A1(c_7_), .A2(d_7_), .ZN(n687) );
  INV_X1 U956 ( .A(c_2_), .ZN(n913) );
  XNOR2_X1 U957 ( .A(n934), .B(n876), .ZN(n619) );
  OR2_X1 U958 ( .A1(n935), .A2(n936), .ZN(n876) );
  AND2_X1 U959 ( .A1(n884), .A2(n937), .ZN(n936) );
  AND2_X1 U960 ( .A1(n938), .A2(n939), .ZN(n935) );
  INV_X1 U961 ( .A(b_2_), .ZN(n939) );
  OR2_X1 U962 ( .A1(n937), .A2(n884), .ZN(n938) );
  OR2_X1 U963 ( .A1(n940), .A2(n941), .ZN(n884) );
  AND2_X1 U964 ( .A1(n889), .A2(n942), .ZN(n941) );
  AND2_X1 U965 ( .A1(n943), .A2(n944), .ZN(n940) );
  INV_X1 U966 ( .A(b_3_), .ZN(n944) );
  OR2_X1 U967 ( .A1(n942), .A2(n889), .ZN(n943) );
  OR2_X1 U968 ( .A1(n945), .A2(n946), .ZN(n889) );
  AND2_X1 U969 ( .A1(n894), .A2(n947), .ZN(n946) );
  AND2_X1 U970 ( .A1(n948), .A2(n949), .ZN(n945) );
  INV_X1 U971 ( .A(b_4_), .ZN(n949) );
  OR2_X1 U972 ( .A1(n947), .A2(n894), .ZN(n948) );
  OR2_X1 U973 ( .A1(n950), .A2(n951), .ZN(n894) );
  AND2_X1 U974 ( .A1(n952), .A2(n953), .ZN(n951) );
  AND2_X1 U975 ( .A1(n954), .A2(n898), .ZN(n950) );
  INV_X1 U976 ( .A(b_5_), .ZN(n898) );
  OR2_X1 U977 ( .A1(n952), .A2(n953), .ZN(n954) );
  INV_X1 U978 ( .A(a_5_), .ZN(n953) );
  INV_X1 U979 ( .A(n896), .ZN(n952) );
  OR2_X1 U980 ( .A1(n955), .A2(n956), .ZN(n896) );
  AND2_X1 U981 ( .A1(n900), .A2(a_6_), .ZN(n956) );
  AND2_X1 U982 ( .A1(b_6_), .A2(n957), .ZN(n955) );
  OR2_X1 U983 ( .A1(n900), .A2(a_6_), .ZN(n957) );
  AND2_X1 U984 ( .A1(a_7_), .A2(b_7_), .ZN(n900) );
  INV_X1 U985 ( .A(a_4_), .ZN(n947) );
  INV_X1 U986 ( .A(a_3_), .ZN(n942) );
  INV_X1 U987 ( .A(a_2_), .ZN(n937) );
  XNOR2_X1 U988 ( .A(a_1_), .B(b_1_), .ZN(n934) );
endmodule

