module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n614_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n421_, new_n620_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n636_, new_n456_, new_n246_, new_n682_, new_n679_, new_n266_, new_n667_, new_n367_, new_n542_, new_n548_, new_n669_, new_n220_, new_n419_, new_n624_, new_n534_, new_n637_, new_n451_, new_n489_, new_n424_, new_n602_, new_n695_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n626_, new_n152_, new_n701_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n655_, new_n630_, new_n167_, new_n385_, new_n478_, new_n694_, new_n461_, new_n297_, new_n361_, new_n683_, new_n183_, new_n511_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n530_, new_n318_, new_n622_, new_n629_, new_n702_, new_n321_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n650_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n506_, new_n680_, new_n256_, new_n452_, new_n381_, new_n656_, new_n388_, new_n508_, new_n194_, new_n483_, new_n394_, new_n299_, new_n657_, new_n652_, new_n314_, new_n582_, new_n363_, new_n165_, new_n441_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n187_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n438_, new_n696_, new_n208_, new_n632_, new_n671_, new_n528_, new_n572_, new_n436_, new_n397_, new_n399_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n628_, new_n162_, new_n409_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n688_, new_n155_, new_n384_, new_n410_, new_n543_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n232_, new_n258_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n654_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n310_, new_n275_, new_n352_, new_n575_, new_n562_, new_n525_, new_n578_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n379_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n520_, new_n253_, new_n403_, new_n475_, new_n237_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n605_, new_n182_, new_n407_, new_n666_, new_n480_, new_n625_, new_n151_, new_n513_, new_n592_, new_n558_, new_n231_, new_n219_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n522_, new_n588_, new_n428_, new_n199_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n191_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n515_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n662_, new_n440_, new_n531_, new_n593_, new_n252_, new_n585_, new_n312_, new_n535_, new_n372_, new_n242_, new_n527_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n651_, new_n433_, new_n435_, new_n265_, new_n687_, new_n370_, new_n689_, new_n584_, new_n278_, new_n304_, new_n523_, new_n638_, new_n550_, new_n217_, new_n269_, new_n512_, new_n644_, new_n599_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n594_, new_n561_, new_n495_, new_n431_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n490_, new_n560_, new_n358_, new_n348_, new_n610_, new_n322_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n226_, new_n697_, new_n185_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n618_, new_n521_, new_n406_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n573_, new_n405_;

not g000 ( new_n151_, N75 );
nand g001 ( new_n152_, N29, N42 );
nor g002 ( N388, new_n152_, new_n151_ );
not g003 ( new_n154_, N29 );
not g004 ( new_n155_, N36 );
nor g005 ( new_n156_, new_n154_, new_n155_ );
and g006 ( N389, new_n156_, N80 );
nand g007 ( new_n158_, new_n156_, N42 );
not g008 ( N390, new_n158_ );
and g009 ( N391, N85, N86 );
not g010 ( new_n161_, N17 );
not g011 ( new_n162_, N13 );
nand g012 ( new_n163_, N1, N8 );
nor g013 ( new_n164_, new_n163_, new_n162_ );
not g014 ( new_n165_, new_n164_ );
nor g015 ( N418, new_n165_, new_n161_ );
nand g016 ( new_n167_, N1, N26 );
nand g017 ( new_n168_, N13, N17 );
nor g018 ( new_n169_, new_n167_, new_n168_ );
nand g019 ( N419, new_n158_, new_n169_ );
not g020 ( new_n171_, N59 );
nor g021 ( new_n172_, new_n171_, new_n151_ );
nand g022 ( N420, new_n172_, N80 );
nor g023 ( new_n174_, new_n155_, new_n171_ );
nand g024 ( N421, new_n174_, N80 );
nand g025 ( N422, new_n174_, N42 );
not g026 ( new_n177_, N90 );
nor g027 ( new_n178_, N87, N88 );
nor g028 ( N423, new_n178_, new_n177_ );
nand g029 ( N446, N390, new_n169_ );
and g030 ( new_n181_, N1, N26 );
nand g031 ( new_n182_, new_n181_, N51 );
nand g032 ( new_n183_, new_n182_, keyIn_0_0 );
not g033 ( new_n184_, keyIn_0_0 );
not g034 ( new_n185_, N51 );
nor g035 ( new_n186_, new_n167_, new_n185_ );
nand g036 ( new_n187_, new_n186_, new_n184_ );
nand g037 ( N447, new_n183_, new_n187_ );
not g038 ( new_n189_, N55 );
nor g039 ( new_n190_, new_n165_, new_n189_ );
not g040 ( new_n191_, new_n190_ );
nand g041 ( new_n192_, N29, N68 );
nor g042 ( N448, new_n191_, new_n192_ );
nand g043 ( new_n194_, N59, N68 );
nor g044 ( new_n195_, new_n191_, new_n194_ );
and g045 ( N449, new_n195_, N74 );
not g046 ( new_n197_, N89 );
nor g047 ( N450, new_n178_, new_n197_ );
not g048 ( new_n199_, keyIn_0_21 );
not g049 ( new_n200_, N135 );
xnor g050 ( new_n201_, N111, N116 );
xnor g051 ( new_n202_, N121, N126 );
xnor g052 ( new_n203_, new_n201_, new_n202_ );
nand g053 ( new_n204_, new_n203_, new_n200_ );
nand g054 ( new_n205_, new_n204_, new_n199_ );
nor g055 ( new_n206_, new_n204_, new_n199_ );
nor g056 ( new_n207_, new_n203_, new_n200_ );
nor g057 ( new_n208_, new_n206_, new_n207_ );
nand g058 ( new_n209_, new_n208_, new_n205_ );
xor g059 ( new_n210_, N101, N106 );
xnor g060 ( new_n211_, N91, N96 );
xnor g061 ( new_n212_, new_n210_, new_n211_ );
xor g062 ( new_n213_, new_n212_, N130 );
xnor g063 ( N767, new_n209_, new_n213_ );
nand g064 ( new_n215_, N183, N189 );
xnor g065 ( new_n216_, new_n215_, keyIn_0_6 );
not g066 ( new_n217_, N183 );
not g067 ( new_n218_, N189 );
nand g068 ( new_n219_, new_n217_, new_n218_ );
nand g069 ( new_n220_, new_n216_, new_n219_ );
xnor g070 ( new_n221_, N195, N201 );
xnor g071 ( new_n222_, new_n220_, new_n221_ );
xnor g072 ( new_n223_, new_n222_, N207 );
xor g073 ( new_n224_, N159, N165 );
xnor g074 ( new_n225_, N171, N177 );
xnor g075 ( new_n226_, new_n224_, new_n225_ );
xnor g076 ( new_n227_, new_n226_, N130 );
xnor g077 ( N768, new_n223_, new_n227_ );
not g078 ( new_n229_, N201 );
not g079 ( new_n230_, keyIn_0_16 );
xnor g080 ( new_n231_, N447, keyIn_0_8 );
nand g081 ( new_n232_, new_n231_, keyIn_0_12 );
not g082 ( new_n233_, keyIn_0_12 );
not g083 ( new_n234_, keyIn_0_8 );
nand g084 ( new_n235_, N447, new_n234_ );
xnor g085 ( new_n236_, new_n186_, keyIn_0_0 );
nand g086 ( new_n237_, new_n236_, keyIn_0_8 );
nand g087 ( new_n238_, new_n237_, new_n235_ );
nand g088 ( new_n239_, new_n238_, new_n233_ );
nand g089 ( new_n240_, new_n232_, new_n239_ );
nand g090 ( new_n241_, N59, N156 );
xnor g091 ( new_n242_, new_n241_, keyIn_0_3 );
nor g092 ( new_n243_, new_n242_, new_n161_ );
nand g093 ( new_n244_, new_n240_, new_n243_ );
nand g094 ( new_n245_, new_n244_, new_n230_ );
not g095 ( new_n246_, N1 );
nor g096 ( new_n247_, new_n244_, new_n230_ );
nor g097 ( new_n248_, new_n247_, new_n246_ );
nand g098 ( new_n249_, new_n248_, new_n245_ );
xnor g099 ( new_n250_, new_n249_, keyIn_0_18 );
nand g100 ( new_n251_, new_n250_, N153 );
not g101 ( new_n252_, keyIn_0_17 );
not g102 ( new_n253_, keyIn_0_15 );
not g103 ( new_n254_, keyIn_0_11 );
nand g104 ( new_n255_, N17, N42 );
xor g105 ( new_n256_, new_n255_, keyIn_0_5 );
nor g106 ( new_n257_, N17, N42 );
xnor g107 ( new_n258_, new_n257_, keyIn_0_4 );
nor g108 ( new_n259_, new_n256_, new_n258_ );
nor g109 ( new_n260_, new_n259_, new_n254_ );
not g110 ( new_n261_, new_n241_ );
nand g111 ( new_n262_, new_n259_, new_n254_ );
nand g112 ( new_n263_, new_n262_, new_n261_ );
nor g113 ( new_n264_, new_n263_, new_n260_ );
nand g114 ( new_n265_, new_n240_, new_n264_ );
xnor g115 ( new_n266_, new_n265_, new_n253_ );
nand g116 ( new_n267_, N17, N51 );
nor g117 ( new_n268_, new_n163_, new_n267_ );
xor g118 ( new_n269_, new_n268_, keyIn_0_1 );
xnor g119 ( new_n270_, new_n269_, keyIn_0_9 );
nand g120 ( new_n271_, N42, N59 );
nor g121 ( new_n272_, new_n271_, new_n151_ );
xor g122 ( new_n273_, new_n272_, keyIn_0_2 );
xnor g123 ( new_n274_, new_n273_, keyIn_0_10 );
nand g124 ( new_n275_, new_n270_, new_n274_ );
xnor g125 ( new_n276_, new_n275_, keyIn_0_13 );
nor g126 ( new_n277_, new_n266_, new_n276_ );
nand g127 ( new_n278_, new_n277_, new_n252_ );
xnor g128 ( new_n279_, new_n265_, keyIn_0_15 );
not g129 ( new_n280_, new_n276_ );
nand g130 ( new_n281_, new_n279_, new_n280_ );
nand g131 ( new_n282_, new_n281_, keyIn_0_17 );
nand g132 ( new_n283_, new_n278_, new_n282_ );
nand g133 ( new_n284_, new_n283_, N126 );
nand g134 ( new_n285_, new_n251_, new_n284_ );
xnor g135 ( new_n286_, new_n285_, keyIn_0_27 );
not g136 ( new_n287_, keyIn_0_14 );
nor g137 ( new_n288_, new_n154_, new_n151_ );
and g138 ( new_n289_, new_n288_, N80 );
and g139 ( new_n290_, new_n240_, new_n289_ );
nand g140 ( new_n291_, new_n290_, N55 );
not g141 ( new_n292_, new_n291_ );
nor g142 ( new_n293_, new_n292_, new_n287_ );
not g143 ( new_n294_, N268 );
nand g144 ( new_n295_, new_n292_, new_n287_ );
nand g145 ( new_n296_, new_n295_, new_n294_ );
nor g146 ( new_n297_, new_n296_, new_n293_ );
not g147 ( new_n298_, new_n297_ );
nand g148 ( new_n299_, new_n286_, new_n298_ );
xor g149 ( new_n300_, new_n299_, keyIn_0_30 );
nand g150 ( new_n301_, new_n300_, new_n229_ );
xnor g151 ( new_n302_, new_n301_, keyIn_0_35 );
not g152 ( new_n303_, new_n302_ );
nor g153 ( new_n304_, new_n300_, new_n229_ );
nor g154 ( new_n305_, new_n303_, new_n304_ );
nand g155 ( new_n306_, new_n305_, N261 );
not g156 ( new_n307_, N219 );
nor g157 ( new_n308_, new_n305_, N261 );
nor g158 ( new_n309_, new_n308_, new_n307_ );
nand g159 ( new_n310_, new_n309_, new_n306_ );
and g160 ( new_n311_, new_n305_, N228 );
nand g161 ( new_n312_, new_n304_, N237 );
not g162 ( new_n313_, N246 );
nor g163 ( new_n314_, new_n300_, new_n313_ );
not g164 ( new_n315_, N73 );
nand g165 ( new_n316_, N42, N72 );
nor g166 ( new_n317_, new_n316_, new_n315_ );
nand g167 ( new_n318_, new_n195_, new_n317_ );
not g168 ( new_n319_, new_n318_ );
nand g169 ( new_n320_, new_n319_, N201 );
not g170 ( new_n321_, keyIn_0_7 );
nand g171 ( new_n322_, N121, N210 );
nor g172 ( new_n323_, new_n322_, new_n321_ );
nand g173 ( new_n324_, new_n322_, new_n321_ );
nand g174 ( new_n325_, N255, N267 );
nand g175 ( new_n326_, new_n324_, new_n325_ );
nor g176 ( new_n327_, new_n326_, new_n323_ );
nand g177 ( new_n328_, new_n320_, new_n327_ );
nor g178 ( new_n329_, new_n314_, new_n328_ );
nand g179 ( new_n330_, new_n329_, new_n312_ );
nor g180 ( new_n331_, new_n311_, new_n330_ );
nand g181 ( N850, new_n310_, new_n331_ );
not g182 ( new_n333_, keyIn_0_42 );
not g183 ( new_n334_, keyIn_0_39 );
not g184 ( new_n335_, keyIn_0_36 );
not g185 ( new_n336_, keyIn_0_31 );
not g186 ( new_n337_, keyIn_0_28 );
nand g187 ( new_n338_, new_n283_, N116 );
xnor g188 ( new_n339_, new_n338_, keyIn_0_23 );
nand g189 ( new_n340_, new_n250_, N146 );
xnor g190 ( new_n341_, new_n340_, keyIn_0_22 );
nand g191 ( new_n342_, new_n341_, new_n339_ );
xnor g192 ( new_n343_, new_n342_, keyIn_0_25 );
xor g193 ( new_n344_, new_n297_, keyIn_0_20 );
nor g194 ( new_n345_, new_n343_, new_n344_ );
nand g195 ( new_n346_, new_n345_, new_n337_ );
not g196 ( new_n347_, keyIn_0_25 );
xnor g197 ( new_n348_, new_n342_, new_n347_ );
not g198 ( new_n349_, new_n344_ );
nand g199 ( new_n350_, new_n348_, new_n349_ );
nand g200 ( new_n351_, new_n350_, keyIn_0_28 );
nand g201 ( new_n352_, new_n346_, new_n351_ );
nor g202 ( new_n353_, new_n352_, new_n218_ );
nand g203 ( new_n354_, new_n353_, new_n336_ );
xnor g204 ( new_n355_, new_n350_, new_n337_ );
nand g205 ( new_n356_, new_n355_, N189 );
nand g206 ( new_n357_, new_n356_, keyIn_0_31 );
nand g207 ( new_n358_, new_n357_, new_n354_ );
xnor g208 ( new_n359_, new_n358_, new_n335_ );
nand g209 ( new_n360_, new_n359_, new_n334_ );
not g210 ( new_n361_, N195 );
not g211 ( new_n362_, keyIn_0_24 );
nand g212 ( new_n363_, new_n283_, N121 );
nand g213 ( new_n364_, new_n363_, new_n362_ );
nor g214 ( new_n365_, new_n363_, new_n362_ );
not g215 ( new_n366_, N149 );
not g216 ( new_n367_, keyIn_0_18 );
xnor g217 ( new_n368_, new_n249_, new_n367_ );
nor g218 ( new_n369_, new_n368_, new_n366_ );
nor g219 ( new_n370_, new_n365_, new_n369_ );
nand g220 ( new_n371_, new_n370_, new_n364_ );
nor g221 ( new_n372_, new_n371_, keyIn_0_26 );
nand g222 ( new_n373_, new_n371_, keyIn_0_26 );
nand g223 ( new_n374_, new_n373_, new_n298_ );
nor g224 ( new_n375_, new_n374_, new_n372_ );
nand g225 ( new_n376_, new_n375_, keyIn_0_29 );
not g226 ( new_n377_, keyIn_0_29 );
not g227 ( new_n378_, new_n372_ );
and g228 ( new_n379_, new_n373_, new_n298_ );
nand g229 ( new_n380_, new_n379_, new_n378_ );
nand g230 ( new_n381_, new_n380_, new_n377_ );
nand g231 ( new_n382_, new_n381_, new_n376_ );
nand g232 ( new_n383_, new_n382_, new_n361_ );
xnor g233 ( new_n384_, new_n383_, keyIn_0_34 );
not g234 ( new_n385_, new_n384_ );
nand g235 ( new_n386_, new_n352_, new_n218_ );
xnor g236 ( new_n387_, new_n386_, keyIn_0_32 );
nand g237 ( new_n388_, new_n302_, N261 );
nor g238 ( new_n389_, new_n387_, new_n388_ );
nand g239 ( new_n390_, new_n389_, new_n385_ );
nand g240 ( new_n391_, new_n390_, keyIn_0_38 );
nand g241 ( new_n392_, new_n360_, new_n391_ );
not g242 ( new_n393_, new_n392_ );
xnor g243 ( new_n394_, new_n358_, keyIn_0_36 );
nand g244 ( new_n395_, new_n394_, keyIn_0_39 );
not g245 ( new_n396_, keyIn_0_38 );
not g246 ( new_n397_, keyIn_0_32 );
xnor g247 ( new_n398_, new_n386_, new_n397_ );
and g248 ( new_n399_, new_n302_, N261 );
nand g249 ( new_n400_, new_n398_, new_n399_ );
nor g250 ( new_n401_, new_n400_, new_n384_ );
nand g251 ( new_n402_, new_n401_, new_n396_ );
and g252 ( new_n403_, new_n395_, new_n402_ );
nand g253 ( new_n404_, new_n393_, new_n403_ );
not g254 ( new_n405_, keyIn_0_41 );
nand g255 ( new_n406_, new_n398_, new_n304_ );
nor g256 ( new_n407_, new_n406_, new_n384_ );
xnor g257 ( new_n408_, new_n407_, new_n405_ );
not g258 ( new_n409_, keyIn_0_37 );
nor g259 ( new_n410_, new_n382_, new_n361_ );
nand g260 ( new_n411_, new_n410_, keyIn_0_33 );
not g261 ( new_n412_, keyIn_0_33 );
xnor g262 ( new_n413_, new_n375_, new_n377_ );
nand g263 ( new_n414_, new_n413_, N195 );
nand g264 ( new_n415_, new_n414_, new_n412_ );
nand g265 ( new_n416_, new_n415_, new_n411_ );
xnor g266 ( new_n417_, new_n416_, new_n409_ );
nand g267 ( new_n418_, new_n417_, new_n398_ );
xnor g268 ( new_n419_, new_n418_, keyIn_0_40 );
nand g269 ( new_n420_, new_n419_, new_n408_ );
nor g270 ( new_n421_, new_n420_, new_n404_ );
nand g271 ( new_n422_, new_n421_, new_n333_ );
nand g272 ( new_n423_, new_n395_, new_n402_ );
nor g273 ( new_n424_, new_n423_, new_n392_ );
xnor g274 ( new_n425_, new_n407_, keyIn_0_41 );
xnor g275 ( new_n426_, new_n416_, keyIn_0_37 );
nor g276 ( new_n427_, new_n426_, new_n387_ );
nand g277 ( new_n428_, new_n427_, keyIn_0_40 );
not g278 ( new_n429_, keyIn_0_40 );
nand g279 ( new_n430_, new_n418_, new_n429_ );
nand g280 ( new_n431_, new_n428_, new_n430_ );
nor g281 ( new_n432_, new_n431_, new_n425_ );
nand g282 ( new_n433_, new_n432_, new_n424_ );
nand g283 ( new_n434_, new_n433_, keyIn_0_42 );
nand g284 ( new_n435_, new_n422_, new_n434_ );
nand g285 ( new_n436_, new_n283_, N111 );
not g286 ( new_n437_, N143 );
nor g287 ( new_n438_, new_n368_, new_n437_ );
xor g288 ( new_n439_, new_n297_, keyIn_0_19 );
nor g289 ( new_n440_, new_n439_, new_n438_ );
nand g290 ( new_n441_, new_n440_, new_n436_ );
nor g291 ( new_n442_, new_n441_, N183 );
not g292 ( new_n443_, new_n442_ );
nand g293 ( new_n444_, new_n435_, new_n443_ );
nand g294 ( new_n445_, new_n441_, N183 );
not g295 ( new_n446_, new_n445_ );
nor g296 ( new_n447_, new_n444_, new_n446_ );
not g297 ( new_n448_, new_n435_ );
nand g298 ( new_n449_, new_n443_, new_n445_ );
nand g299 ( new_n450_, new_n448_, new_n449_ );
nand g300 ( new_n451_, new_n450_, N219 );
or g301 ( new_n452_, new_n451_, new_n447_ );
not g302 ( new_n453_, N228 );
nor g303 ( new_n454_, new_n449_, new_n453_ );
nand g304 ( new_n455_, new_n446_, N237 );
nand g305 ( new_n456_, new_n441_, N246 );
nor g306 ( new_n457_, new_n318_, new_n217_ );
and g307 ( new_n458_, N106, N210 );
nor g308 ( new_n459_, new_n457_, new_n458_ );
and g309 ( new_n460_, new_n456_, new_n459_ );
nand g310 ( new_n461_, new_n455_, new_n460_ );
nor g311 ( new_n462_, new_n454_, new_n461_ );
nand g312 ( N863, new_n452_, new_n462_ );
or g313 ( new_n464_, new_n399_, new_n304_ );
nand g314 ( new_n465_, new_n464_, new_n385_ );
nand g315 ( new_n466_, new_n465_, new_n426_ );
nor g316 ( new_n467_, new_n387_, new_n358_ );
nor g317 ( new_n468_, new_n466_, new_n467_ );
nand g318 ( new_n469_, new_n466_, new_n467_ );
nand g319 ( new_n470_, new_n469_, N219 );
nor g320 ( new_n471_, new_n470_, new_n468_ );
and g321 ( new_n472_, N111, N210 );
nor g322 ( new_n473_, new_n471_, new_n472_ );
xnor g323 ( new_n474_, new_n473_, keyIn_0_50 );
not g324 ( new_n475_, N237 );
nor g325 ( new_n476_, new_n359_, new_n475_ );
nand g326 ( new_n477_, new_n467_, N228 );
nor g327 ( new_n478_, new_n352_, new_n313_ );
nand g328 ( new_n479_, new_n319_, N189 );
nand g329 ( new_n480_, N255, N259 );
nand g330 ( new_n481_, new_n479_, new_n480_ );
nor g331 ( new_n482_, new_n478_, new_n481_ );
nand g332 ( new_n483_, new_n477_, new_n482_ );
nor g333 ( new_n484_, new_n476_, new_n483_ );
nand g334 ( N864, new_n474_, new_n484_ );
not g335 ( new_n486_, new_n416_ );
nor g336 ( new_n487_, new_n486_, new_n384_ );
or g337 ( new_n488_, new_n464_, new_n487_ );
nor g338 ( new_n489_, new_n465_, new_n486_ );
nor g339 ( new_n490_, new_n489_, new_n307_ );
nand g340 ( new_n491_, new_n490_, new_n488_ );
nor g341 ( new_n492_, new_n426_, new_n475_ );
nand g342 ( new_n493_, new_n487_, N228 );
nor g343 ( new_n494_, new_n382_, new_n313_ );
nand g344 ( new_n495_, new_n319_, N195 );
nand g345 ( new_n496_, N255, N260 );
nand g346 ( new_n497_, N116, N210 );
and g347 ( new_n498_, new_n496_, new_n497_ );
nand g348 ( new_n499_, new_n495_, new_n498_ );
nor g349 ( new_n500_, new_n494_, new_n499_ );
nand g350 ( new_n501_, new_n493_, new_n500_ );
nor g351 ( new_n502_, new_n501_, new_n492_ );
nand g352 ( N865, new_n491_, new_n502_ );
not g353 ( new_n504_, keyIn_0_44 );
not g354 ( new_n505_, keyIn_0_43 );
xnor g355 ( new_n506_, new_n444_, new_n505_ );
nor g356 ( new_n507_, new_n506_, new_n446_ );
nand g357 ( new_n508_, new_n507_, new_n504_ );
xnor g358 ( new_n509_, new_n444_, keyIn_0_43 );
nand g359 ( new_n510_, new_n509_, new_n445_ );
nand g360 ( new_n511_, new_n510_, keyIn_0_44 );
nand g361 ( new_n512_, new_n508_, new_n511_ );
nand g362 ( new_n513_, new_n283_, N96 );
not g363 ( new_n514_, N146 );
nor g364 ( new_n515_, new_n242_, new_n189_ );
nand g365 ( new_n516_, new_n240_, new_n515_ );
nor g366 ( new_n517_, new_n516_, new_n514_ );
nor g367 ( new_n518_, new_n161_, N268 );
nand g368 ( new_n519_, new_n290_, new_n518_ );
nand g369 ( new_n520_, N51, N138 );
nand g370 ( new_n521_, new_n519_, new_n520_ );
nor g371 ( new_n522_, new_n521_, new_n517_ );
nand g372 ( new_n523_, new_n513_, new_n522_ );
nor g373 ( new_n524_, new_n523_, N165 );
nand g374 ( new_n525_, new_n283_, N101 );
nor g375 ( new_n526_, new_n516_, new_n366_ );
nand g376 ( new_n527_, N17, N138 );
nand g377 ( new_n528_, new_n519_, new_n527_ );
nor g378 ( new_n529_, new_n528_, new_n526_ );
nand g379 ( new_n530_, new_n525_, new_n529_ );
nor g380 ( new_n531_, new_n530_, N171 );
nor g381 ( new_n532_, new_n524_, new_n531_ );
nand g382 ( new_n533_, new_n283_, N106 );
not g383 ( new_n534_, N153 );
nor g384 ( new_n535_, new_n516_, new_n534_ );
nand g385 ( new_n536_, N138, N152 );
nand g386 ( new_n537_, new_n519_, new_n536_ );
nor g387 ( new_n538_, new_n537_, new_n535_ );
nand g388 ( new_n539_, new_n533_, new_n538_ );
nor g389 ( new_n540_, new_n539_, N177 );
not g390 ( new_n541_, new_n540_ );
nand g391 ( new_n542_, new_n532_, new_n541_ );
not g392 ( new_n543_, new_n542_ );
nand g393 ( new_n544_, new_n512_, new_n543_ );
nor g394 ( new_n545_, new_n544_, keyIn_0_47 );
nand g395 ( new_n546_, new_n544_, keyIn_0_47 );
nand g396 ( new_n547_, new_n539_, N177 );
nand g397 ( new_n548_, new_n530_, N171 );
nand g398 ( new_n549_, new_n547_, new_n548_ );
nand g399 ( new_n550_, new_n532_, new_n549_ );
nand g400 ( new_n551_, new_n523_, N165 );
and g401 ( new_n552_, new_n550_, new_n551_ );
nand g402 ( new_n553_, new_n546_, new_n552_ );
nor g403 ( new_n554_, new_n553_, new_n545_ );
xnor g404 ( new_n555_, new_n554_, keyIn_0_48 );
nand g405 ( new_n556_, new_n283_, N91 );
nor g406 ( new_n557_, new_n516_, new_n437_ );
nand g407 ( new_n558_, N8, N138 );
nand g408 ( new_n559_, new_n519_, new_n558_ );
nor g409 ( new_n560_, new_n559_, new_n557_ );
nand g410 ( new_n561_, new_n556_, new_n560_ );
or g411 ( new_n562_, new_n561_, N159 );
nand g412 ( new_n563_, new_n555_, new_n562_ );
nand g413 ( new_n564_, new_n561_, N159 );
nand g414 ( N866, new_n563_, new_n564_ );
not g415 ( new_n566_, keyIn_0_55 );
not g416 ( new_n567_, keyIn_0_49 );
not g417 ( new_n568_, new_n512_ );
nand g418 ( new_n569_, new_n541_, new_n547_ );
nor g419 ( new_n570_, new_n568_, new_n569_ );
xnor g420 ( new_n571_, new_n570_, keyIn_0_46 );
nand g421 ( new_n572_, new_n568_, new_n569_ );
xor g422 ( new_n573_, new_n572_, keyIn_0_45 );
nand g423 ( new_n574_, new_n573_, new_n571_ );
nor g424 ( new_n575_, new_n574_, new_n567_ );
nand g425 ( new_n576_, new_n574_, new_n567_ );
nand g426 ( new_n577_, new_n576_, N219 );
nor g427 ( new_n578_, new_n577_, new_n575_ );
xor g428 ( new_n579_, new_n578_, keyIn_0_53 );
nand g429 ( new_n580_, N101, N210 );
nand g430 ( new_n581_, new_n579_, new_n580_ );
nor g431 ( new_n582_, new_n581_, new_n566_ );
nand g432 ( new_n583_, new_n581_, new_n566_ );
nor g433 ( new_n584_, new_n569_, new_n453_ );
nor g434 ( new_n585_, new_n547_, new_n475_ );
nand g435 ( new_n586_, new_n539_, N246 );
nand g436 ( new_n587_, new_n319_, N177 );
nand g437 ( new_n588_, new_n586_, new_n587_ );
or g438 ( new_n589_, new_n585_, new_n588_ );
nor g439 ( new_n590_, new_n584_, new_n589_ );
nand g440 ( new_n591_, new_n583_, new_n590_ );
nor g441 ( new_n592_, new_n591_, new_n582_ );
xnor g442 ( new_n593_, new_n592_, keyIn_0_57 );
xor g443 ( new_n594_, new_n593_, keyIn_0_59 );
xnor g444 ( N874, new_n594_, keyIn_0_61 );
not g445 ( new_n596_, keyIn_0_63 );
not g446 ( new_n597_, keyIn_0_58 );
not g447 ( new_n598_, keyIn_0_56 );
not g448 ( new_n599_, keyIn_0_54 );
not g449 ( new_n600_, keyIn_0_48 );
nand g450 ( new_n601_, new_n554_, new_n600_ );
not g451 ( new_n602_, new_n545_ );
and g452 ( new_n603_, new_n546_, new_n552_ );
nand g453 ( new_n604_, new_n603_, new_n602_ );
nand g454 ( new_n605_, new_n604_, keyIn_0_48 );
nand g455 ( new_n606_, new_n605_, new_n601_ );
nand g456 ( new_n607_, new_n562_, new_n564_ );
nand g457 ( new_n608_, new_n606_, new_n607_ );
nand g458 ( new_n609_, new_n608_, keyIn_0_51 );
not g459 ( new_n610_, new_n607_ );
nand g460 ( new_n611_, new_n555_, new_n610_ );
nand g461 ( new_n612_, new_n611_, keyIn_0_52 );
and g462 ( new_n613_, new_n612_, new_n609_ );
nor g463 ( new_n614_, new_n611_, keyIn_0_52 );
nor g464 ( new_n615_, new_n608_, keyIn_0_51 );
nor g465 ( new_n616_, new_n614_, new_n615_ );
nand g466 ( new_n617_, new_n613_, new_n616_ );
nand g467 ( new_n618_, new_n617_, new_n599_ );
nand g468 ( new_n619_, new_n612_, new_n609_ );
not g469 ( new_n620_, keyIn_0_52 );
nor g470 ( new_n621_, new_n606_, new_n607_ );
nand g471 ( new_n622_, new_n621_, new_n620_ );
not g472 ( new_n623_, keyIn_0_51 );
nor g473 ( new_n624_, new_n555_, new_n610_ );
nand g474 ( new_n625_, new_n624_, new_n623_ );
nand g475 ( new_n626_, new_n625_, new_n622_ );
nor g476 ( new_n627_, new_n626_, new_n619_ );
nand g477 ( new_n628_, new_n627_, keyIn_0_54 );
nand g478 ( new_n629_, new_n618_, new_n628_ );
nand g479 ( new_n630_, new_n629_, N219 );
xnor g480 ( new_n631_, new_n630_, new_n598_ );
not g481 ( new_n632_, N210 );
nor g482 ( new_n633_, new_n632_, new_n294_ );
nor g483 ( new_n634_, new_n631_, new_n633_ );
nor g484 ( new_n635_, new_n634_, new_n597_ );
not g485 ( new_n636_, new_n635_ );
nand g486 ( new_n637_, new_n630_, keyIn_0_56 );
and g487 ( new_n638_, new_n629_, N219 );
nand g488 ( new_n639_, new_n638_, new_n598_ );
nand g489 ( new_n640_, new_n639_, new_n637_ );
not g490 ( new_n641_, new_n633_ );
nand g491 ( new_n642_, new_n640_, new_n641_ );
nor g492 ( new_n643_, new_n642_, keyIn_0_58 );
nor g493 ( new_n644_, new_n607_, new_n453_ );
nor g494 ( new_n645_, new_n564_, new_n475_ );
nand g495 ( new_n646_, new_n561_, N246 );
nand g496 ( new_n647_, new_n319_, N159 );
nand g497 ( new_n648_, new_n646_, new_n647_ );
nor g498 ( new_n649_, new_n645_, new_n648_ );
not g499 ( new_n650_, new_n649_ );
nor g500 ( new_n651_, new_n650_, new_n644_ );
not g501 ( new_n652_, new_n651_ );
nor g502 ( new_n653_, new_n643_, new_n652_ );
nand g503 ( new_n654_, new_n653_, new_n636_ );
nand g504 ( new_n655_, new_n654_, keyIn_0_60 );
not g505 ( new_n656_, keyIn_0_60 );
nand g506 ( new_n657_, new_n634_, new_n597_ );
nand g507 ( new_n658_, new_n657_, new_n651_ );
nor g508 ( new_n659_, new_n658_, new_n635_ );
nand g509 ( new_n660_, new_n659_, new_n656_ );
nand g510 ( new_n661_, new_n660_, new_n655_ );
xnor g511 ( new_n662_, new_n661_, keyIn_0_62 );
nand g512 ( new_n663_, new_n662_, new_n596_ );
not g513 ( new_n664_, keyIn_0_62 );
nand g514 ( new_n665_, new_n661_, new_n664_ );
xnor g515 ( new_n666_, new_n654_, new_n656_ );
nand g516 ( new_n667_, new_n666_, keyIn_0_62 );
nand g517 ( new_n668_, new_n667_, new_n665_ );
nand g518 ( new_n669_, new_n668_, keyIn_0_63 );
nand g519 ( N878, new_n663_, new_n669_ );
not g520 ( new_n671_, new_n531_ );
nand g521 ( new_n672_, new_n512_, new_n541_ );
nand g522 ( new_n673_, new_n672_, new_n547_ );
nand g523 ( new_n674_, new_n673_, new_n671_ );
nand g524 ( new_n675_, new_n674_, new_n548_ );
not g525 ( new_n676_, new_n551_ );
nor g526 ( new_n677_, new_n676_, new_n524_ );
nor g527 ( new_n678_, new_n675_, new_n677_ );
nand g528 ( new_n679_, new_n675_, new_n677_ );
nand g529 ( new_n680_, new_n679_, N219 );
or g530 ( new_n681_, new_n680_, new_n678_ );
and g531 ( new_n682_, new_n677_, N228 );
nand g532 ( new_n683_, new_n676_, N237 );
and g533 ( new_n684_, new_n523_, N246 );
nand g534 ( new_n685_, new_n319_, N165 );
nand g535 ( new_n686_, N91, N210 );
nand g536 ( new_n687_, new_n685_, new_n686_ );
nor g537 ( new_n688_, new_n684_, new_n687_ );
nand g538 ( new_n689_, new_n688_, new_n683_ );
nor g539 ( new_n690_, new_n682_, new_n689_ );
nand g540 ( N879, new_n681_, new_n690_ );
not g541 ( new_n692_, new_n548_ );
nor g542 ( new_n693_, new_n692_, new_n531_ );
nor g543 ( new_n694_, new_n673_, new_n693_ );
nand g544 ( new_n695_, new_n673_, new_n693_ );
nand g545 ( new_n696_, new_n695_, N219 );
or g546 ( new_n697_, new_n696_, new_n694_ );
and g547 ( new_n698_, new_n693_, N228 );
nand g548 ( new_n699_, new_n692_, N237 );
and g549 ( new_n700_, new_n530_, N246 );
nand g550 ( new_n701_, new_n319_, N171 );
nand g551 ( new_n702_, N96, N210 );
nand g552 ( new_n703_, new_n701_, new_n702_ );
nor g553 ( new_n704_, new_n700_, new_n703_ );
nand g554 ( new_n705_, new_n704_, new_n699_ );
nor g555 ( new_n706_, new_n698_, new_n705_ );
nand g556 ( N880, new_n697_, new_n706_ );
endmodule