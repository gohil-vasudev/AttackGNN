module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n155_, new_n384_, new_n410_, new_n445_, new_n236_, new_n238_, new_n479_, new_n92_, new_n79_, new_n543_, new_n250_, new_n113_, new_n501_, new_n288_, new_n371_, new_n509_, new_n97_, new_n454_, new_n421_, new_n202_, new_n296_, new_n308_, new_n368_, new_n232_, new_n258_, new_n76_, new_n439_, new_n176_, new_n283_, new_n223_, new_n390_, new_n156_, new_n306_, new_n366_, new_n494_, new_n291_, new_n241_, new_n261_, new_n309_, new_n186_, new_n365_, new_n339_, new_n197_, new_n529_, new_n386_, new_n82_, new_n401_, new_n389_, new_n323_, new_n259_, new_n362_, new_n556_, new_n227_, new_n416_, new_n222_, new_n456_, new_n170_, new_n246_, new_n400_, new_n328_, new_n460_, new_n266_, new_n367_, new_n542_, new_n548_, new_n173_, new_n220_, new_n130_, new_n505_, new_n419_, new_n471_, new_n268_, new_n374_, new_n534_, new_n376_, new_n380_, new_n214_, new_n451_, new_n489_, new_n424_, new_n138_, new_n310_, new_n144_, new_n275_, new_n114_, new_n188_, new_n240_, new_n413_, new_n526_, new_n352_, new_n442_, new_n485_, new_n525_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n126_, new_n462_, new_n177_, new_n493_, new_n264_, new_n379_, new_n500_, new_n273_, new_n224_, new_n270_, new_n317_, new_n102_, new_n344_, new_n143_, new_n520_, new_n287_, new_n125_, new_n145_, new_n253_, new_n504_, new_n403_, new_n475_, new_n90_, new_n237_, new_n427_, new_n234_, new_n532_, new_n149_, new_n472_, new_n557_, new_n393_, new_n260_, new_n418_, new_n251_, new_n189_, new_n300_, new_n292_, new_n106_, new_n411_, new_n215_, new_n507_, new_n152_, new_n157_, new_n107_, new_n93_, new_n182_, new_n153_, new_n407_, new_n81_, new_n480_, new_n133_, new_n257_, new_n481_, new_n212_, new_n151_, new_n513_, new_n364_, new_n449_, new_n558_, new_n484_, new_n219_, new_n231_, new_n313_, new_n78_, new_n239_, new_n272_, new_n282_, new_n382_, new_n522_, new_n201_, new_n428_, new_n192_, new_n414_, new_n199_, new_n146_, new_n88_, new_n487_, new_n360_, new_n98_, new_n546_, new_n110_, new_n315_, new_n302_, new_n191_, new_n124_, new_n326_, new_n554_, new_n95_, new_n225_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n87_, new_n387_, new_n544_, new_n103_, new_n476_, new_n112_, new_n248_, new_n350_, new_n117_, new_n121_, new_n415_, new_n167_, new_n537_, new_n221_, new_n385_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n478_, new_n461_, new_n459_, new_n555_, new_n174_, new_n297_, new_n361_, new_n468_, new_n150_, new_n354_, new_n392_, new_n444_, new_n518_, new_n108_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n105_, new_n340_, new_n147_, new_n510_, new_n285_, new_n502_, new_n80_, new_n351_, new_n209_, new_n337_, new_n446_, new_n203_, new_n316_, new_n517_, new_n325_, new_n417_, new_n180_, new_n515_, new_n530_, new_n332_, new_n318_, new_n453_, new_n516_, new_n163_, new_n519_, new_n148_, new_n321_, new_n440_, new_n443_, new_n324_, new_n122_, new_n531_, new_n111_, new_n252_, new_n486_, new_n491_, new_n549_, new_n466_, new_n262_, new_n160_, new_n312_, new_n271_, new_n535_, new_n274_, new_n372_, new_n100_, new_n242_, new_n503_, new_n527_, new_n218_, new_n497_, new_n115_, new_n307_, new_n190_, new_n305_, new_n420_, new_n470_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n213_, new_n134_, new_n433_, new_n435_, new_n206_, new_n109_, new_n254_, new_n429_, new_n355_, new_n353_, new_n85_, new_n432_, new_n265_, new_n506_, new_n370_, new_n256_, new_n452_, new_n278_, new_n304_, new_n381_, new_n523_, new_n388_, new_n550_, new_n217_, new_n101_, new_n269_, new_n508_, new_n512_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n129_, new_n142_, new_n139_, new_n314_, new_n118_, new_n363_, new_n412_, new_n165_, new_n441_, new_n477_, new_n327_, new_n216_, new_n495_, new_n431_, new_n77_, new_n196_, new_n280_, new_n426_, new_n319_, new_n235_, new_n398_, new_n301_, new_n169_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n338_, new_n207_, new_n267_, new_n473_, new_n140_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n187_, new_n311_, new_n86_, new_n465_, new_n84_, new_n195_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n357_, new_n320_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n245_, new_n402_, new_n474_, new_n89_, new_n467_, new_n286_, new_n404_, new_n335_, new_n347_, new_n193_, new_n490_, new_n560_, new_n91_, new_n346_, new_n396_, new_n198_, new_n438_, new_n128_, new_n358_, new_n208_, new_n348_, new_n159_, new_n83_, new_n322_, new_n228_, new_n545_, new_n289_, new_n528_, new_n179_, new_n425_, new_n436_, new_n175_, new_n226_, new_n397_, new_n104_, new_n185_, new_n399_, new_n373_, new_n171_, new_n559_, new_n540_, new_n434_, new_n200_, new_n422_, new_n99_, new_n329_, new_n249_, new_n233_, new_n136_, new_n469_, new_n119_, new_n293_, new_n391_, new_n96_, new_n178_, new_n437_, new_n551_, new_n168_, new_n279_, new_n455_, new_n295_, new_n359_, new_n132_, new_n120_, new_n521_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n553_, new_n406_, new_n356_, new_n333_, new_n229_, new_n536_, new_n290_, new_n464_, new_n94_, new_n204_, new_n369_, new_n181_, new_n135_, new_n448_, new_n276_, new_n405_;

not g000 ( new_n76_, keyIn_0_6 );
not g001 ( new_n77_, keyIn_0_4 );
not g002 ( new_n78_, N69 );
and g003 ( new_n79_, keyIn_0_1, N63 );
not g004 ( new_n80_, new_n79_ );
or g005 ( new_n81_, keyIn_0_1, N63 );
and g006 ( new_n82_, new_n80_, new_n81_ );
or g007 ( new_n83_, new_n82_, new_n78_ );
and g008 ( new_n84_, new_n83_, new_n77_ );
not g009 ( new_n85_, keyIn_0_1 );
not g010 ( new_n86_, N63 );
and g011 ( new_n87_, new_n85_, new_n86_ );
or g012 ( new_n88_, new_n87_, new_n79_ );
and g013 ( new_n89_, new_n88_, N69 );
and g014 ( new_n90_, new_n89_, keyIn_0_4 );
or g015 ( new_n91_, new_n84_, new_n90_ );
not g016 ( new_n92_, N24 );
and g017 ( new_n93_, new_n92_, N30 );
not g018 ( new_n94_, N102 );
and g019 ( new_n95_, new_n94_, N108 );
or g020 ( new_n96_, new_n93_, new_n95_ );
not g021 ( new_n97_, new_n96_ );
not g022 ( new_n98_, N82 );
or g023 ( new_n99_, new_n98_, N76 );
not g024 ( new_n100_, N43 );
or g025 ( new_n101_, new_n100_, N37 );
and g026 ( new_n102_, new_n99_, new_n101_ );
not g027 ( new_n103_, N4 );
or g028 ( new_n104_, new_n103_, N1 );
not g029 ( new_n105_, N56 );
or g030 ( new_n106_, new_n105_, N50 );
and g031 ( new_n107_, new_n104_, new_n106_ );
and g032 ( new_n108_, new_n102_, new_n107_ );
and g033 ( new_n109_, new_n108_, new_n97_ );
not g034 ( new_n110_, new_n109_ );
or g035 ( new_n111_, new_n91_, new_n110_ );
not g036 ( new_n112_, keyIn_0_5 );
not g037 ( new_n113_, keyIn_0_2 );
and g038 ( new_n114_, new_n113_, N89 );
not g039 ( new_n115_, N95 );
not g040 ( new_n116_, N89 );
and g041 ( new_n117_, new_n116_, keyIn_0_2 );
or g042 ( new_n118_, new_n117_, new_n115_ );
or g043 ( new_n119_, new_n118_, new_n114_ );
or g044 ( new_n120_, new_n119_, new_n112_ );
not g045 ( new_n121_, new_n114_ );
or g046 ( new_n122_, new_n113_, N89 );
and g047 ( new_n123_, new_n122_, N95 );
and g048 ( new_n124_, new_n123_, new_n121_ );
or g049 ( new_n125_, new_n124_, keyIn_0_5 );
and g050 ( new_n126_, new_n120_, new_n125_ );
not g051 ( new_n127_, keyIn_0_3 );
not g052 ( new_n128_, keyIn_0_0 );
not g053 ( new_n129_, N11 );
and g054 ( new_n130_, new_n128_, new_n129_ );
and g055 ( new_n131_, keyIn_0_0, N11 );
or g056 ( new_n132_, new_n130_, new_n131_ );
and g057 ( new_n133_, new_n132_, N17 );
or g058 ( new_n134_, new_n133_, new_n127_ );
not g059 ( new_n135_, N17 );
or g060 ( new_n136_, keyIn_0_0, N11 );
not g061 ( new_n137_, new_n131_ );
and g062 ( new_n138_, new_n137_, new_n136_ );
or g063 ( new_n139_, new_n138_, new_n135_ );
or g064 ( new_n140_, new_n139_, keyIn_0_3 );
and g065 ( new_n141_, new_n134_, new_n140_ );
or g066 ( new_n142_, new_n126_, new_n141_ );
or g067 ( new_n143_, new_n142_, new_n111_ );
and g068 ( new_n144_, new_n143_, new_n76_ );
or g069 ( new_n145_, new_n89_, keyIn_0_4 );
or g070 ( new_n146_, new_n83_, new_n77_ );
and g071 ( new_n147_, new_n145_, new_n146_ );
and g072 ( new_n148_, new_n147_, new_n109_ );
and g073 ( new_n149_, new_n124_, keyIn_0_5 );
and g074 ( new_n150_, new_n119_, new_n112_ );
or g075 ( new_n151_, new_n150_, new_n149_ );
and g076 ( new_n152_, new_n139_, keyIn_0_3 );
and g077 ( new_n153_, new_n133_, new_n127_ );
or g078 ( new_n154_, new_n152_, new_n153_ );
and g079 ( new_n155_, new_n154_, new_n151_ );
and g080 ( new_n156_, new_n155_, new_n148_ );
and g081 ( new_n157_, new_n156_, keyIn_0_6 );
or g082 ( N223, new_n144_, new_n157_ );
not g083 ( new_n159_, keyIn_0_13 );
not g084 ( new_n160_, keyIn_0_10 );
not g085 ( new_n161_, keyIn_0_7 );
and g086 ( new_n162_, N223, new_n161_ );
or g087 ( new_n163_, new_n156_, keyIn_0_6 );
or g088 ( new_n164_, new_n143_, new_n76_ );
and g089 ( new_n165_, new_n164_, new_n163_ );
and g090 ( new_n166_, new_n165_, keyIn_0_7 );
or g091 ( new_n167_, new_n162_, new_n166_ );
and g092 ( new_n168_, new_n167_, new_n151_ );
or g093 ( new_n169_, new_n165_, keyIn_0_7 );
or g094 ( new_n170_, N223, new_n161_ );
and g095 ( new_n171_, new_n169_, new_n170_ );
and g096 ( new_n172_, new_n171_, new_n126_ );
or g097 ( new_n173_, new_n168_, new_n172_ );
and g098 ( new_n174_, new_n173_, new_n160_ );
not g099 ( new_n175_, new_n174_ );
or g100 ( new_n176_, new_n173_, new_n160_ );
and g101 ( new_n177_, new_n175_, new_n176_ );
or g102 ( new_n178_, new_n177_, new_n115_ );
or g103 ( new_n179_, new_n178_, N99 );
not g104 ( new_n180_, new_n179_ );
and g105 ( new_n181_, new_n180_, keyIn_0_12 );
not g106 ( new_n182_, keyIn_0_12 );
and g107 ( new_n183_, new_n179_, new_n182_ );
or g108 ( new_n184_, new_n181_, new_n183_ );
not g109 ( new_n185_, keyIn_0_11 );
not g110 ( new_n186_, keyIn_0_8 );
and g111 ( new_n187_, new_n167_, new_n104_ );
not g112 ( new_n188_, new_n104_ );
and g113 ( new_n189_, new_n171_, new_n188_ );
or g114 ( new_n190_, new_n187_, new_n189_ );
or g115 ( new_n191_, new_n190_, new_n186_ );
or g116 ( new_n192_, new_n171_, new_n188_ );
or g117 ( new_n193_, new_n167_, new_n104_ );
and g118 ( new_n194_, new_n193_, new_n192_ );
or g119 ( new_n195_, new_n194_, keyIn_0_8 );
and g120 ( new_n196_, new_n191_, new_n195_ );
or g121 ( new_n197_, new_n196_, new_n103_ );
or g122 ( new_n198_, new_n197_, N8 );
or g123 ( new_n199_, new_n198_, new_n185_ );
not g124 ( new_n200_, N8 );
and g125 ( new_n201_, new_n194_, keyIn_0_8 );
and g126 ( new_n202_, new_n190_, new_n186_ );
or g127 ( new_n203_, new_n202_, new_n201_ );
and g128 ( new_n204_, new_n203_, N4 );
and g129 ( new_n205_, new_n204_, new_n200_ );
or g130 ( new_n206_, new_n205_, keyIn_0_11 );
and g131 ( new_n207_, new_n199_, new_n206_ );
not g132 ( new_n208_, N34 );
not g133 ( new_n209_, new_n93_ );
and g134 ( new_n210_, new_n167_, new_n209_ );
and g135 ( new_n211_, new_n171_, new_n93_ );
or g136 ( new_n212_, new_n210_, new_n211_ );
and g137 ( new_n213_, new_n212_, N30 );
and g138 ( new_n214_, new_n213_, new_n208_ );
not g139 ( new_n215_, N86 );
and g140 ( new_n216_, new_n167_, new_n99_ );
not g141 ( new_n217_, new_n216_ );
or g142 ( new_n218_, new_n167_, new_n99_ );
and g143 ( new_n219_, new_n217_, new_n218_ );
not g144 ( new_n220_, new_n219_ );
and g145 ( new_n221_, new_n220_, N82 );
and g146 ( new_n222_, new_n221_, new_n215_ );
or g147 ( new_n223_, new_n222_, new_n214_ );
not g148 ( new_n224_, N60 );
not g149 ( new_n225_, new_n106_ );
and g150 ( new_n226_, new_n171_, new_n225_ );
and g151 ( new_n227_, new_n167_, new_n106_ );
or g152 ( new_n228_, new_n227_, new_n226_ );
and g153 ( new_n229_, new_n228_, N56 );
and g154 ( new_n230_, new_n229_, new_n224_ );
not g155 ( new_n231_, N112 );
and g156 ( new_n232_, new_n171_, new_n95_ );
not g157 ( new_n233_, new_n232_ );
or g158 ( new_n234_, new_n171_, new_n95_ );
and g159 ( new_n235_, new_n233_, new_n234_ );
not g160 ( new_n236_, new_n235_ );
and g161 ( new_n237_, new_n236_, N108 );
and g162 ( new_n238_, new_n237_, new_n231_ );
or g163 ( new_n239_, new_n238_, new_n230_ );
or g164 ( new_n240_, new_n223_, new_n239_ );
not g165 ( new_n241_, keyIn_0_9 );
and g166 ( new_n242_, new_n167_, new_n154_ );
and g167 ( new_n243_, new_n171_, new_n141_ );
or g168 ( new_n244_, new_n242_, new_n243_ );
or g169 ( new_n245_, new_n244_, new_n241_ );
and g170 ( new_n246_, new_n245_, N17 );
and g171 ( new_n247_, new_n244_, new_n241_ );
or g172 ( new_n248_, new_n247_, N21 );
not g173 ( new_n249_, new_n248_ );
and g174 ( new_n250_, new_n249_, new_n246_ );
not g175 ( new_n251_, N73 );
and g176 ( new_n252_, new_n167_, new_n147_ );
and g177 ( new_n253_, new_n171_, new_n91_ );
or g178 ( new_n254_, new_n252_, new_n253_ );
and g179 ( new_n255_, new_n254_, N69 );
and g180 ( new_n256_, new_n255_, new_n251_ );
not g181 ( new_n257_, N47 );
and g182 ( new_n258_, new_n167_, new_n101_ );
or g183 ( new_n259_, new_n167_, new_n101_ );
not g184 ( new_n260_, new_n259_ );
or g185 ( new_n261_, new_n260_, new_n258_ );
and g186 ( new_n262_, new_n261_, N43 );
and g187 ( new_n263_, new_n262_, new_n257_ );
or g188 ( new_n264_, new_n263_, new_n256_ );
or g189 ( new_n265_, new_n264_, new_n250_ );
or g190 ( new_n266_, new_n240_, new_n265_ );
or g191 ( new_n267_, new_n207_, new_n266_ );
or g192 ( new_n268_, new_n267_, new_n184_ );
and g193 ( new_n269_, new_n268_, new_n159_ );
or g194 ( new_n270_, new_n179_, new_n182_ );
not g195 ( new_n271_, new_n183_ );
and g196 ( new_n272_, new_n271_, new_n270_ );
and g197 ( new_n273_, new_n205_, keyIn_0_11 );
and g198 ( new_n274_, new_n198_, new_n185_ );
or g199 ( new_n275_, new_n274_, new_n273_ );
not g200 ( new_n276_, new_n223_ );
not g201 ( new_n277_, new_n239_ );
and g202 ( new_n278_, new_n276_, new_n277_ );
not g203 ( new_n279_, new_n265_ );
and g204 ( new_n280_, new_n278_, new_n279_ );
and g205 ( new_n281_, new_n275_, new_n280_ );
and g206 ( new_n282_, new_n281_, new_n272_ );
and g207 ( new_n283_, new_n282_, keyIn_0_13 );
or g208 ( N329, new_n269_, new_n283_ );
not g209 ( new_n285_, keyIn_0_20 );
not g210 ( new_n286_, keyIn_0_16 );
and g211 ( new_n287_, N329, keyIn_0_15 );
not g212 ( new_n288_, keyIn_0_15 );
or g213 ( new_n289_, new_n282_, keyIn_0_13 );
or g214 ( new_n290_, new_n268_, new_n159_ );
and g215 ( new_n291_, new_n290_, new_n289_ );
and g216 ( new_n292_, new_n291_, new_n288_ );
or g217 ( new_n293_, new_n287_, new_n292_ );
and g218 ( new_n294_, new_n293_, new_n275_ );
or g219 ( new_n295_, new_n291_, new_n288_ );
or g220 ( new_n296_, N329, keyIn_0_15 );
and g221 ( new_n297_, new_n295_, new_n296_ );
and g222 ( new_n298_, new_n297_, new_n207_ );
or g223 ( new_n299_, new_n294_, new_n298_ );
not g224 ( new_n300_, new_n299_ );
and g225 ( new_n301_, new_n300_, new_n286_ );
not g226 ( new_n302_, new_n301_ );
and g227 ( new_n303_, new_n299_, keyIn_0_16 );
not g228 ( new_n304_, new_n303_ );
or g229 ( new_n305_, new_n197_, N14 );
and g230 ( new_n306_, new_n305_, keyIn_0_14 );
not g231 ( new_n307_, new_n306_ );
or g232 ( new_n308_, new_n305_, keyIn_0_14 );
and g233 ( new_n309_, new_n307_, new_n308_ );
and g234 ( new_n310_, new_n304_, new_n309_ );
and g235 ( new_n311_, new_n310_, new_n302_ );
and g236 ( new_n312_, new_n311_, keyIn_0_18 );
not g237 ( new_n313_, new_n312_ );
or g238 ( new_n314_, new_n311_, keyIn_0_18 );
and g239 ( new_n315_, new_n313_, new_n314_ );
not g240 ( new_n316_, keyIn_0_19 );
not g241 ( new_n317_, keyIn_0_17 );
not g242 ( new_n318_, new_n230_ );
and g243 ( new_n319_, new_n293_, new_n318_ );
and g244 ( new_n320_, new_n297_, new_n230_ );
or g245 ( new_n321_, new_n319_, new_n320_ );
or g246 ( new_n322_, new_n321_, new_n317_ );
or g247 ( new_n323_, new_n297_, new_n230_ );
or g248 ( new_n324_, new_n293_, new_n318_ );
and g249 ( new_n325_, new_n324_, new_n323_ );
or g250 ( new_n326_, new_n325_, keyIn_0_17 );
and g251 ( new_n327_, new_n322_, new_n326_ );
not g252 ( new_n328_, N66 );
and g253 ( new_n329_, new_n229_, new_n328_ );
not g254 ( new_n330_, new_n329_ );
or g255 ( new_n331_, new_n327_, new_n330_ );
or g256 ( new_n332_, new_n331_, new_n316_ );
and g257 ( new_n333_, new_n325_, keyIn_0_17 );
and g258 ( new_n334_, new_n321_, new_n317_ );
or g259 ( new_n335_, new_n334_, new_n333_ );
and g260 ( new_n336_, new_n335_, new_n329_ );
or g261 ( new_n337_, new_n336_, keyIn_0_19 );
and g262 ( new_n338_, new_n332_, new_n337_ );
and g263 ( new_n339_, new_n293_, new_n272_ );
and g264 ( new_n340_, new_n297_, new_n184_ );
or g265 ( new_n341_, new_n339_, new_n340_ );
not g266 ( new_n342_, N105 );
not g267 ( new_n343_, new_n178_ );
and g268 ( new_n344_, new_n343_, new_n342_ );
and g269 ( new_n345_, new_n341_, new_n344_ );
not g270 ( new_n346_, new_n250_ );
and g271 ( new_n347_, new_n293_, new_n346_ );
and g272 ( new_n348_, new_n297_, new_n250_ );
or g273 ( new_n349_, new_n347_, new_n348_ );
not g274 ( new_n350_, N27 );
not g275 ( new_n351_, new_n247_ );
and g276 ( new_n352_, new_n351_, new_n350_ );
and g277 ( new_n353_, new_n352_, new_n246_ );
and g278 ( new_n354_, new_n349_, new_n353_ );
not g279 ( new_n355_, new_n222_ );
and g280 ( new_n356_, new_n293_, new_n355_ );
and g281 ( new_n357_, new_n297_, new_n222_ );
or g282 ( new_n358_, new_n356_, new_n357_ );
not g283 ( new_n359_, N92 );
and g284 ( new_n360_, new_n221_, new_n359_ );
and g285 ( new_n361_, new_n358_, new_n360_ );
or g286 ( new_n362_, new_n354_, new_n361_ );
or g287 ( new_n363_, new_n362_, new_n345_ );
not g288 ( new_n364_, new_n256_ );
and g289 ( new_n365_, new_n293_, new_n364_ );
and g290 ( new_n366_, new_n297_, new_n256_ );
or g291 ( new_n367_, new_n365_, new_n366_ );
not g292 ( new_n368_, N79 );
and g293 ( new_n369_, new_n255_, new_n368_ );
and g294 ( new_n370_, new_n367_, new_n369_ );
not g295 ( new_n371_, new_n238_ );
and g296 ( new_n372_, new_n293_, new_n371_ );
and g297 ( new_n373_, new_n297_, new_n238_ );
or g298 ( new_n374_, new_n372_, new_n373_ );
not g299 ( new_n375_, N115 );
and g300 ( new_n376_, new_n237_, new_n375_ );
and g301 ( new_n377_, new_n374_, new_n376_ );
or g302 ( new_n378_, new_n370_, new_n377_ );
not g303 ( new_n379_, new_n263_ );
and g304 ( new_n380_, new_n293_, new_n379_ );
and g305 ( new_n381_, new_n297_, new_n263_ );
or g306 ( new_n382_, new_n380_, new_n381_ );
not g307 ( new_n383_, N53 );
and g308 ( new_n384_, new_n262_, new_n383_ );
and g309 ( new_n385_, new_n382_, new_n384_ );
not g310 ( new_n386_, new_n214_ );
and g311 ( new_n387_, new_n293_, new_n386_ );
and g312 ( new_n388_, new_n297_, new_n214_ );
or g313 ( new_n389_, new_n387_, new_n388_ );
not g314 ( new_n390_, N40 );
and g315 ( new_n391_, new_n213_, new_n390_ );
and g316 ( new_n392_, new_n389_, new_n391_ );
or g317 ( new_n393_, new_n385_, new_n392_ );
or g318 ( new_n394_, new_n378_, new_n393_ );
or g319 ( new_n395_, new_n394_, new_n363_ );
or g320 ( new_n396_, new_n338_, new_n395_ );
or g321 ( new_n397_, new_n396_, new_n315_ );
and g322 ( new_n398_, new_n397_, new_n285_ );
not g323 ( new_n399_, new_n314_ );
or g324 ( new_n400_, new_n399_, new_n312_ );
and g325 ( new_n401_, new_n336_, keyIn_0_19 );
and g326 ( new_n402_, new_n331_, new_n316_ );
or g327 ( new_n403_, new_n402_, new_n401_ );
not g328 ( new_n404_, new_n395_ );
and g329 ( new_n405_, new_n403_, new_n404_ );
and g330 ( new_n406_, new_n405_, new_n400_ );
and g331 ( new_n407_, new_n406_, keyIn_0_20 );
or g332 ( N370, new_n398_, new_n407_ );
or g333 ( new_n409_, new_n406_, keyIn_0_20 );
or g334 ( new_n410_, new_n397_, new_n285_ );
and g335 ( new_n411_, new_n410_, new_n409_ );
and g336 ( new_n412_, new_n411_, keyIn_0_21 );
not g337 ( new_n413_, keyIn_0_21 );
and g338 ( new_n414_, N370, new_n413_ );
or g339 ( new_n415_, new_n412_, new_n414_ );
and g340 ( new_n416_, new_n415_, N40 );
and g341 ( new_n417_, new_n416_, keyIn_0_22 );
not g342 ( new_n418_, keyIn_0_22 );
or g343 ( new_n419_, N370, new_n413_ );
or g344 ( new_n420_, new_n411_, keyIn_0_21 );
and g345 ( new_n421_, new_n419_, new_n420_ );
or g346 ( new_n422_, new_n421_, new_n390_ );
and g347 ( new_n423_, new_n422_, new_n418_ );
and g348 ( new_n424_, N329, N34 );
not g349 ( new_n425_, N30 );
and g350 ( new_n426_, N223, N24 );
or g351 ( new_n427_, new_n426_, new_n425_ );
or g352 ( new_n428_, new_n424_, new_n427_ );
or g353 ( new_n429_, new_n423_, new_n428_ );
or g354 ( new_n430_, new_n429_, new_n417_ );
and g355 ( new_n431_, new_n430_, keyIn_0_24 );
not g356 ( new_n432_, keyIn_0_24 );
not g357 ( new_n433_, new_n417_ );
or g358 ( new_n434_, new_n416_, keyIn_0_22 );
not g359 ( new_n435_, new_n428_ );
and g360 ( new_n436_, new_n434_, new_n435_ );
and g361 ( new_n437_, new_n436_, new_n433_ );
and g362 ( new_n438_, new_n437_, new_n432_ );
or g363 ( new_n439_, new_n431_, new_n438_ );
and g364 ( new_n440_, new_n415_, N27 );
and g365 ( new_n441_, N329, N21 );
and g366 ( new_n442_, N223, N11 );
or g367 ( new_n443_, new_n442_, new_n135_ );
or g368 ( new_n444_, new_n441_, new_n443_ );
or g369 ( new_n445_, new_n440_, new_n444_ );
and g370 ( new_n446_, new_n439_, new_n445_ );
and g371 ( new_n447_, new_n415_, N66 );
and g372 ( new_n448_, N329, N60 );
and g373 ( new_n449_, N223, N50 );
or g374 ( new_n450_, new_n449_, new_n105_ );
or g375 ( new_n451_, new_n448_, new_n450_ );
or g376 ( new_n452_, new_n447_, new_n451_ );
and g377 ( new_n453_, new_n446_, new_n452_ );
not g378 ( new_n454_, new_n453_ );
not g379 ( new_n455_, keyIn_0_25 );
and g380 ( new_n456_, new_n415_, N53 );
and g381 ( new_n457_, new_n456_, keyIn_0_23 );
not g382 ( new_n458_, keyIn_0_23 );
or g383 ( new_n459_, new_n421_, new_n383_ );
and g384 ( new_n460_, new_n459_, new_n458_ );
and g385 ( new_n461_, N329, N47 );
and g386 ( new_n462_, N223, N37 );
or g387 ( new_n463_, new_n462_, new_n100_ );
or g388 ( new_n464_, new_n461_, new_n463_ );
or g389 ( new_n465_, new_n460_, new_n464_ );
or g390 ( new_n466_, new_n465_, new_n457_ );
and g391 ( new_n467_, new_n466_, new_n455_ );
not g392 ( new_n468_, new_n457_ );
or g393 ( new_n469_, new_n456_, keyIn_0_23 );
not g394 ( new_n470_, new_n464_ );
and g395 ( new_n471_, new_n469_, new_n470_ );
and g396 ( new_n472_, new_n471_, new_n468_ );
and g397 ( new_n473_, new_n472_, keyIn_0_25 );
or g398 ( new_n474_, new_n467_, new_n473_ );
not g399 ( new_n475_, new_n474_ );
and g400 ( new_n476_, new_n415_, N92 );
and g401 ( new_n477_, N329, N86 );
and g402 ( new_n478_, N223, N76 );
or g403 ( new_n479_, new_n478_, new_n98_ );
or g404 ( new_n480_, new_n477_, new_n479_ );
or g405 ( new_n481_, new_n476_, new_n480_ );
not g406 ( new_n482_, new_n481_ );
and g407 ( new_n483_, new_n415_, N79 );
and g408 ( new_n484_, N329, N73 );
and g409 ( new_n485_, N223, N63 );
or g410 ( new_n486_, new_n485_, new_n78_ );
or g411 ( new_n487_, new_n484_, new_n486_ );
or g412 ( new_n488_, new_n483_, new_n487_ );
not g413 ( new_n489_, new_n488_ );
or g414 ( new_n490_, new_n482_, new_n489_ );
and g415 ( new_n491_, new_n415_, N105 );
and g416 ( new_n492_, N329, N99 );
and g417 ( new_n493_, N223, N89 );
or g418 ( new_n494_, new_n493_, new_n115_ );
or g419 ( new_n495_, new_n492_, new_n494_ );
or g420 ( new_n496_, new_n491_, new_n495_ );
not g421 ( new_n497_, new_n496_ );
or g422 ( new_n498_, new_n421_, new_n375_ );
or g423 ( new_n499_, new_n291_, new_n231_ );
or g424 ( new_n500_, new_n165_, new_n94_ );
and g425 ( new_n501_, new_n500_, N108 );
and g426 ( new_n502_, new_n499_, new_n501_ );
and g427 ( new_n503_, new_n498_, new_n502_ );
or g428 ( new_n504_, new_n497_, new_n503_ );
or g429 ( new_n505_, new_n490_, new_n504_ );
or g430 ( new_n506_, new_n475_, new_n505_ );
or g431 ( new_n507_, new_n454_, new_n506_ );
and g432 ( new_n508_, new_n415_, N14 );
and g433 ( new_n509_, N329, N8 );
and g434 ( new_n510_, N223, N1 );
or g435 ( new_n511_, new_n510_, new_n103_ );
or g436 ( new_n512_, new_n509_, new_n511_ );
or g437 ( new_n513_, new_n508_, new_n512_ );
and g438 ( N421, new_n507_, new_n513_ );
not g439 ( new_n515_, keyIn_0_30 );
not g440 ( new_n516_, keyIn_0_27 );
or g441 ( new_n517_, new_n474_, keyIn_0_26 );
not g442 ( new_n518_, new_n517_ );
and g443 ( new_n519_, new_n474_, keyIn_0_26 );
or g444 ( new_n520_, new_n518_, new_n519_ );
and g445 ( new_n521_, new_n520_, new_n439_ );
or g446 ( new_n522_, new_n521_, new_n516_ );
not g447 ( new_n523_, new_n439_ );
not g448 ( new_n524_, new_n519_ );
and g449 ( new_n525_, new_n524_, new_n517_ );
or g450 ( new_n526_, new_n525_, new_n523_ );
or g451 ( new_n527_, new_n526_, keyIn_0_27 );
and g452 ( new_n528_, new_n522_, new_n527_ );
and g453 ( new_n529_, new_n528_, new_n453_ );
not g454 ( new_n530_, new_n529_ );
and g455 ( new_n531_, new_n530_, new_n515_ );
and g456 ( new_n532_, new_n529_, keyIn_0_30 );
or g457 ( N430, new_n531_, new_n532_ );
and g458 ( new_n534_, new_n439_, new_n474_ );
and g459 ( new_n535_, new_n489_, new_n452_ );
and g460 ( new_n536_, new_n534_, new_n535_ );
not g461 ( new_n537_, new_n536_ );
or g462 ( new_n538_, new_n537_, keyIn_0_28 );
not g463 ( new_n539_, keyIn_0_28 );
or g464 ( new_n540_, new_n536_, new_n539_ );
and g465 ( new_n541_, new_n538_, new_n540_ );
not g466 ( new_n542_, new_n541_ );
not g467 ( new_n543_, new_n446_ );
and g468 ( new_n544_, new_n482_, new_n452_ );
and g469 ( new_n545_, new_n474_, new_n544_ );
or g470 ( new_n546_, new_n543_, new_n545_ );
or g471 ( N431, new_n542_, new_n546_ );
and g472 ( new_n548_, new_n497_, new_n481_ );
and g473 ( new_n549_, new_n534_, new_n548_ );
not g474 ( new_n550_, new_n549_ );
or g475 ( new_n551_, new_n550_, keyIn_0_29 );
not g476 ( new_n552_, keyIn_0_29 );
or g477 ( new_n553_, new_n549_, new_n552_ );
and g478 ( new_n554_, new_n553_, new_n445_ );
and g479 ( new_n555_, new_n554_, new_n551_ );
and g480 ( new_n556_, new_n555_, new_n541_ );
and g481 ( new_n557_, new_n556_, new_n528_ );
and g482 ( new_n558_, new_n557_, keyIn_0_31 );
not g483 ( new_n559_, new_n558_ );
or g484 ( new_n560_, new_n557_, keyIn_0_31 );
and g485 ( N432, new_n559_, new_n560_ );
endmodule