module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n595_, new_n614_, new_n445_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n421_, new_n620_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n456_, new_n246_, new_n170_, new_n266_, new_n367_, new_n542_, new_n548_, new_n173_, new_n220_, new_n419_, new_n624_, new_n534_, new_n214_, new_n451_, new_n489_, new_n424_, new_n602_, new_n188_, new_n240_, new_n413_, new_n526_, new_n442_, new_n211_, new_n552_, new_n342_, new_n462_, new_n603_, new_n564_, new_n500_, new_n317_, new_n287_, new_n504_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n626_, new_n152_, new_n153_, new_n257_, new_n481_, new_n212_, new_n449_, new_n364_, new_n580_, new_n484_, new_n272_, new_n282_, new_n201_, new_n192_, new_n414_, new_n315_, new_n326_, new_n554_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n630_, new_n167_, new_n385_, new_n478_, new_n461_, new_n297_, new_n361_, new_n565_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n622_, new_n629_, new_n321_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n549_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n506_, new_n256_, new_n452_, new_n381_, new_n388_, new_n508_, new_n483_, new_n394_, new_n299_, new_n314_, new_n582_, new_n363_, new_n165_, new_n441_, new_n477_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n488_, new_n524_, new_n277_, new_n402_, new_n579_, new_n286_, new_n335_, new_n347_, new_n346_, new_n396_, new_n198_, new_n438_, new_n208_, new_n528_, new_n572_, new_n436_, new_n397_, new_n399_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n628_, new_n162_, new_n409_, new_n457_, new_n553_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n155_, new_n384_, new_n410_, new_n543_, new_n371_, new_n509_, new_n202_, new_n296_, new_n308_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n604_, new_n227_, new_n416_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n310_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n562_, new_n578_, new_n493_, new_n264_, new_n379_, new_n273_, new_n270_, new_n598_, new_n570_, new_n520_, new_n253_, new_n403_, new_n475_, new_n237_, new_n557_, new_n260_, new_n189_, new_n300_, new_n411_, new_n507_, new_n605_, new_n407_, new_n480_, new_n625_, new_n151_, new_n513_, new_n592_, new_n558_, new_n219_, new_n583_, new_n231_, new_n313_, new_n382_, new_n239_, new_n617_, new_n522_, new_n588_, new_n199_, new_n487_, new_n360_, new_n546_, new_n612_, new_n302_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n285_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n591_, new_n515_, new_n332_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n440_, new_n531_, new_n593_, new_n252_, new_n585_, new_n312_, new_n535_, new_n372_, new_n242_, new_n503_, new_n527_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n433_, new_n435_, new_n265_, new_n370_, new_n584_, new_n278_, new_n304_, new_n523_, new_n550_, new_n217_, new_n269_, new_n512_, new_n599_, new_n412_, new_n607_, new_n327_, new_n594_, new_n561_, new_n495_, new_n431_, new_n196_, new_n574_, new_n319_, new_n338_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n627_, new_n195_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n358_, new_n348_, new_n610_, new_n159_, new_n322_, new_n228_, new_n545_, new_n289_, new_n425_, new_n226_, new_n185_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n551_, new_n168_, new_n279_, new_n455_, new_n618_, new_n521_, new_n406_, new_n356_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n573_, new_n405_;

not g000 ( new_n151_, N75 );
nand g001 ( new_n152_, N29, N42 );
nor g002 ( new_n153_, new_n152_, new_n151_ );
xnor g003 ( N388, new_n153_, keyIn_0_3 );
not g004 ( new_n155_, N80 );
nand g005 ( new_n156_, N29, N36 );
nor g006 ( N389, new_n156_, new_n155_ );
not g007 ( new_n158_, N42 );
nor g008 ( new_n159_, new_n156_, new_n158_ );
xor g009 ( N390, new_n159_, keyIn_0_4 );
and g010 ( N391, N85, N86 );
not g011 ( new_n162_, N13 );
nand g012 ( new_n163_, N1, N8 );
nor g013 ( new_n164_, new_n163_, new_n162_ );
nand g014 ( new_n165_, new_n164_, N17 );
xnor g015 ( N418, new_n165_, keyIn_0_0 );
xnor g016 ( new_n167_, new_n159_, keyIn_0_1 );
not g017 ( new_n168_, new_n167_ );
nand g018 ( new_n169_, N1, N26 );
nand g019 ( new_n170_, N13, N17 );
nor g020 ( new_n171_, new_n169_, new_n170_ );
nand g021 ( N419, new_n168_, new_n171_ );
not g022 ( new_n173_, N59 );
nor g023 ( new_n174_, new_n173_, new_n151_ );
nand g024 ( N420, new_n174_, N80 );
nand g025 ( new_n176_, N36, N59 );
or g026 ( N421, new_n176_, new_n155_ );
nor g027 ( new_n178_, new_n176_, new_n158_ );
xnor g028 ( N422, new_n178_, keyIn_0_5 );
not g029 ( new_n180_, N90 );
nor g030 ( new_n181_, N87, N88 );
nor g031 ( N423, new_n181_, new_n180_ );
nand g032 ( N446, new_n167_, new_n171_ );
not g033 ( new_n184_, keyIn_0_2 );
not g034 ( new_n185_, N51 );
nor g035 ( new_n186_, new_n169_, new_n185_ );
xnor g036 ( N447, new_n186_, new_n184_ );
not g037 ( new_n188_, N29 );
and g038 ( new_n189_, N55, N68 );
nand g039 ( new_n190_, new_n164_, new_n189_ );
nor g040 ( N448, new_n190_, new_n188_ );
nand g041 ( new_n192_, N59, N74 );
nor g042 ( new_n193_, new_n190_, new_n192_ );
xnor g043 ( N449, new_n193_, keyIn_0_12 );
not g044 ( new_n195_, N89 );
nor g045 ( new_n196_, new_n181_, new_n195_ );
xnor g046 ( N450, new_n196_, keyIn_0_9 );
not g047 ( new_n198_, keyIn_0_32 );
not g048 ( new_n199_, N135 );
not g049 ( new_n200_, keyIn_0_6 );
nor g050 ( new_n201_, N111, N116 );
nand g051 ( new_n202_, new_n201_, new_n200_ );
and g052 ( new_n203_, N111, N116 );
nor g053 ( new_n204_, new_n201_, new_n200_ );
nor g054 ( new_n205_, new_n204_, new_n203_ );
nand g055 ( new_n206_, new_n205_, new_n202_ );
xnor g056 ( new_n207_, N121, N126 );
xnor g057 ( new_n208_, new_n206_, new_n207_ );
nand g058 ( new_n209_, new_n208_, new_n199_ );
nor g059 ( new_n210_, new_n209_, keyIn_0_19 );
or g060 ( new_n211_, new_n208_, new_n199_ );
nand g061 ( new_n212_, new_n209_, keyIn_0_19 );
nand g062 ( new_n213_, new_n212_, new_n211_ );
nor g063 ( new_n214_, new_n213_, new_n210_ );
xnor g064 ( new_n215_, N91, N96 );
xnor g065 ( new_n216_, N101, N106 );
xnor g066 ( new_n217_, new_n215_, new_n216_ );
xnor g067 ( new_n218_, new_n217_, N130 );
and g068 ( new_n219_, new_n214_, new_n218_ );
nor g069 ( new_n220_, new_n219_, new_n198_ );
or g070 ( new_n221_, new_n214_, new_n218_ );
nand g071 ( new_n222_, new_n219_, new_n198_ );
nand g072 ( new_n223_, new_n222_, new_n221_ );
nor g073 ( N767, new_n223_, new_n220_ );
not g074 ( new_n225_, keyIn_0_25 );
xor g075 ( new_n226_, N171, N177 );
not g076 ( new_n227_, N159 );
not g077 ( new_n228_, N165 );
nand g078 ( new_n229_, new_n227_, new_n228_ );
nor g079 ( new_n230_, new_n227_, new_n228_ );
nor g080 ( new_n231_, new_n230_, keyIn_0_13 );
nand g081 ( new_n232_, new_n231_, new_n229_ );
xnor g082 ( new_n233_, new_n232_, new_n226_ );
nor g083 ( new_n234_, new_n233_, N130 );
nor g084 ( new_n235_, new_n234_, new_n225_ );
nand g085 ( new_n236_, new_n234_, new_n225_ );
nand g086 ( new_n237_, new_n233_, N130 );
and g087 ( new_n238_, new_n237_, keyIn_0_31 );
nand g088 ( new_n239_, new_n238_, new_n236_ );
nor g089 ( new_n240_, new_n239_, new_n235_ );
not g090 ( new_n241_, N207 );
xnor g091 ( new_n242_, N183, N189 );
xnor g092 ( new_n243_, N195, N201 );
xnor g093 ( new_n244_, new_n242_, new_n243_ );
nand g094 ( new_n245_, new_n244_, new_n241_ );
nand g095 ( new_n246_, new_n245_, keyIn_0_26 );
nor g096 ( new_n247_, new_n245_, keyIn_0_26 );
nor g097 ( new_n248_, new_n244_, new_n241_ );
nor g098 ( new_n249_, new_n247_, new_n248_ );
nand g099 ( new_n250_, new_n249_, new_n246_ );
xnor g100 ( N768, new_n240_, new_n250_ );
not g101 ( new_n252_, keyIn_0_56 );
not g102 ( new_n253_, N201 );
not g103 ( new_n254_, keyIn_0_15 );
nor g104 ( new_n255_, new_n188_, new_n151_ );
nand g105 ( new_n256_, new_n255_, N80 );
nand g106 ( new_n257_, N447, N55 );
nor g107 ( new_n258_, new_n257_, new_n256_ );
nor g108 ( new_n259_, new_n258_, new_n254_ );
xor g109 ( new_n260_, keyIn_0_10, N268 );
nand g110 ( new_n261_, new_n258_, new_n254_ );
nand g111 ( new_n262_, new_n261_, new_n260_ );
nor g112 ( new_n263_, new_n262_, new_n259_ );
and g113 ( new_n264_, N59, N156 );
not g114 ( new_n265_, new_n264_ );
not g115 ( new_n266_, N17 );
and g116 ( new_n267_, N1, N26 );
nand g117 ( new_n268_, new_n267_, N51 );
nand g118 ( new_n269_, new_n268_, new_n184_ );
nand g119 ( new_n270_, new_n186_, keyIn_0_2 );
nand g120 ( new_n271_, new_n269_, new_n270_ );
nor g121 ( new_n272_, new_n271_, new_n266_ );
nand g122 ( new_n273_, new_n272_, new_n265_ );
nand g123 ( new_n274_, new_n273_, N1 );
nand g124 ( new_n275_, new_n274_, N153 );
not g125 ( new_n276_, keyIn_0_24 );
not g126 ( new_n277_, N126 );
nor g127 ( new_n278_, N17, N42 );
nand g128 ( new_n279_, N17, N42 );
nand g129 ( new_n280_, new_n264_, new_n279_ );
or g130 ( new_n281_, new_n280_, new_n278_ );
nor g131 ( new_n282_, new_n271_, new_n281_ );
nor g132 ( new_n283_, new_n158_, new_n173_ );
and g133 ( new_n284_, new_n283_, N75 );
nand g134 ( new_n285_, N17, N51 );
or g135 ( new_n286_, new_n163_, new_n285_ );
nor g136 ( new_n287_, new_n284_, new_n286_ );
nor g137 ( new_n288_, new_n282_, new_n287_ );
nor g138 ( new_n289_, new_n288_, new_n277_ );
nand g139 ( new_n290_, new_n289_, new_n276_ );
nor g140 ( new_n291_, new_n280_, new_n278_ );
nand g141 ( new_n292_, N447, new_n291_ );
not g142 ( new_n293_, new_n287_ );
nand g143 ( new_n294_, new_n292_, new_n293_ );
nand g144 ( new_n295_, new_n294_, N126 );
nand g145 ( new_n296_, new_n295_, keyIn_0_24 );
nand g146 ( new_n297_, new_n290_, new_n296_ );
nand g147 ( new_n298_, new_n297_, new_n275_ );
nor g148 ( new_n299_, new_n298_, new_n263_ );
or g149 ( new_n300_, new_n299_, new_n253_ );
xnor g150 ( new_n301_, new_n300_, keyIn_0_37 );
not g151 ( new_n302_, new_n301_ );
nand g152 ( new_n303_, new_n299_, new_n253_ );
xnor g153 ( new_n304_, new_n303_, keyIn_0_38 );
nor g154 ( new_n305_, new_n302_, new_n304_ );
xnor g155 ( new_n306_, new_n305_, N261 );
nand g156 ( new_n307_, new_n306_, keyIn_0_52 );
not g157 ( new_n308_, N219 );
nor g158 ( new_n309_, new_n306_, keyIn_0_52 );
nor g159 ( new_n310_, new_n309_, new_n308_ );
nand g160 ( new_n311_, new_n310_, new_n307_ );
nand g161 ( new_n312_, N121, N210 );
nand g162 ( new_n313_, new_n311_, new_n312_ );
nand g163 ( new_n314_, new_n313_, new_n252_ );
nor g164 ( new_n315_, new_n313_, new_n252_ );
not g165 ( new_n316_, keyIn_0_28 );
nand g166 ( new_n317_, new_n283_, N72 );
nor g167 ( new_n318_, new_n190_, new_n317_ );
nand g168 ( new_n319_, new_n318_, keyIn_0_8 );
or g169 ( new_n320_, new_n318_, keyIn_0_8 );
and g170 ( new_n321_, new_n320_, N73 );
nand g171 ( new_n322_, new_n321_, new_n319_ );
xnor g172 ( new_n323_, new_n322_, keyIn_0_11 );
xnor g173 ( new_n324_, new_n323_, keyIn_0_14 );
xor g174 ( new_n325_, new_n324_, keyIn_0_16 );
not g175 ( new_n326_, new_n325_ );
nand g176 ( new_n327_, new_n326_, N201 );
nor g177 ( new_n328_, new_n327_, new_n316_ );
nand g178 ( new_n329_, new_n327_, new_n316_ );
not g179 ( new_n330_, N246 );
nor g180 ( new_n331_, new_n299_, new_n330_ );
and g181 ( new_n332_, N255, N267 );
nor g182 ( new_n333_, new_n331_, new_n332_ );
nand g183 ( new_n334_, new_n329_, new_n333_ );
nor g184 ( new_n335_, new_n334_, new_n328_ );
nand g185 ( new_n336_, new_n302_, N237 );
nor g186 ( new_n337_, new_n336_, keyIn_0_50 );
nand g187 ( new_n338_, new_n305_, N228 );
nand g188 ( new_n339_, new_n336_, keyIn_0_50 );
nand g189 ( new_n340_, new_n338_, new_n339_ );
nor g190 ( new_n341_, new_n340_, new_n337_ );
nand g191 ( new_n342_, new_n335_, new_n341_ );
nor g192 ( new_n343_, new_n315_, new_n342_ );
nand g193 ( N850, new_n343_, new_n314_ );
not g194 ( new_n345_, keyIn_0_53 );
not g195 ( new_n346_, keyIn_0_51 );
not g196 ( new_n347_, keyIn_0_23 );
nand g197 ( new_n348_, new_n294_, N116 );
nor g198 ( new_n349_, new_n348_, new_n347_ );
not g199 ( new_n350_, new_n349_ );
nand g200 ( new_n351_, new_n348_, new_n347_ );
nand g201 ( new_n352_, new_n274_, N146 );
and g202 ( new_n353_, new_n351_, new_n352_ );
nand g203 ( new_n354_, new_n353_, new_n350_ );
nor g204 ( new_n355_, new_n354_, new_n263_ );
nand g205 ( new_n356_, new_n355_, keyIn_0_30 );
not g206 ( new_n357_, keyIn_0_30 );
not g207 ( new_n358_, new_n263_ );
nand g208 ( new_n359_, new_n351_, new_n352_ );
nor g209 ( new_n360_, new_n359_, new_n349_ );
nand g210 ( new_n361_, new_n360_, new_n358_ );
nand g211 ( new_n362_, new_n361_, new_n357_ );
nand g212 ( new_n363_, new_n356_, new_n362_ );
nor g213 ( new_n364_, new_n363_, N189 );
nand g214 ( new_n365_, new_n294_, N121 );
nand g215 ( new_n366_, new_n274_, N149 );
nand g216 ( new_n367_, new_n366_, new_n365_ );
or g217 ( new_n368_, new_n263_, new_n367_ );
nor g218 ( new_n369_, new_n368_, N195 );
nor g219 ( new_n370_, new_n364_, new_n369_ );
nand g220 ( new_n371_, new_n302_, new_n370_ );
xnor g221 ( new_n372_, new_n371_, new_n346_ );
not g222 ( new_n373_, N261 );
nor g223 ( new_n374_, new_n304_, new_n373_ );
nand g224 ( new_n375_, new_n374_, new_n370_ );
nor g225 ( new_n376_, new_n375_, keyIn_0_42 );
nand g226 ( new_n377_, new_n375_, keyIn_0_42 );
nand g227 ( new_n378_, new_n368_, N195 );
nor g228 ( new_n379_, new_n364_, new_n378_ );
nand g229 ( new_n380_, new_n363_, N189 );
not g230 ( new_n381_, new_n380_ );
nor g231 ( new_n382_, new_n379_, new_n381_ );
nand g232 ( new_n383_, new_n377_, new_n382_ );
nor g233 ( new_n384_, new_n383_, new_n376_ );
nand g234 ( new_n385_, new_n384_, new_n372_ );
not g235 ( new_n386_, new_n385_ );
not g236 ( new_n387_, keyIn_0_36 );
not g237 ( new_n388_, keyIn_0_29 );
nand g238 ( new_n389_, new_n294_, N111 );
nor g239 ( new_n390_, new_n389_, keyIn_0_22 );
nand g240 ( new_n391_, new_n274_, N143 );
nand g241 ( new_n392_, new_n389_, keyIn_0_22 );
nand g242 ( new_n393_, new_n392_, new_n391_ );
nor g243 ( new_n394_, new_n393_, new_n390_ );
nand g244 ( new_n395_, new_n394_, new_n358_ );
xnor g245 ( new_n396_, new_n395_, new_n388_ );
nand g246 ( new_n397_, new_n396_, N183 );
xnor g247 ( new_n398_, new_n397_, new_n387_ );
or g248 ( new_n399_, new_n396_, N183 );
nand g249 ( new_n400_, new_n398_, new_n399_ );
or g250 ( new_n401_, new_n386_, new_n400_ );
nor g251 ( new_n402_, new_n401_, new_n345_ );
nand g252 ( new_n403_, new_n386_, new_n400_ );
nand g253 ( new_n404_, new_n401_, new_n345_ );
nand g254 ( new_n405_, new_n404_, new_n403_ );
nor g255 ( new_n406_, new_n405_, new_n402_ );
nor g256 ( new_n407_, new_n406_, keyIn_0_55 );
nand g257 ( new_n408_, new_n406_, keyIn_0_55 );
nand g258 ( new_n409_, new_n408_, N219 );
or g259 ( new_n410_, new_n409_, new_n407_ );
not g260 ( new_n411_, keyIn_0_40 );
xnor g261 ( new_n412_, new_n398_, new_n411_ );
nand g262 ( new_n413_, new_n412_, N237 );
not g263 ( new_n414_, keyIn_0_27 );
nand g264 ( new_n415_, new_n326_, N183 );
nor g265 ( new_n416_, new_n415_, new_n414_ );
nand g266 ( new_n417_, new_n415_, new_n414_ );
nand g267 ( new_n418_, new_n396_, N246 );
nand g268 ( new_n419_, N106, N210 );
and g269 ( new_n420_, new_n418_, new_n419_ );
nand g270 ( new_n421_, new_n417_, new_n420_ );
nor g271 ( new_n422_, new_n421_, new_n416_ );
nand g272 ( new_n423_, new_n422_, new_n413_ );
not g273 ( new_n424_, N228 );
nor g274 ( new_n425_, new_n400_, new_n424_ );
xnor g275 ( new_n426_, new_n425_, keyIn_0_47 );
nor g276 ( new_n427_, new_n426_, new_n423_ );
nand g277 ( N863, new_n410_, new_n427_ );
nor g278 ( new_n429_, new_n381_, new_n364_ );
not g279 ( new_n430_, new_n369_ );
or g280 ( new_n431_, new_n302_, new_n374_ );
nand g281 ( new_n432_, new_n431_, new_n430_ );
xnor g282 ( new_n433_, new_n378_, keyIn_0_49 );
nand g283 ( new_n434_, new_n432_, new_n433_ );
nand g284 ( new_n435_, new_n434_, new_n429_ );
nor g285 ( new_n436_, new_n434_, new_n429_ );
nor g286 ( new_n437_, new_n436_, new_n308_ );
nand g287 ( new_n438_, new_n437_, new_n435_ );
nand g288 ( new_n439_, new_n363_, N246 );
nand g289 ( new_n440_, N255, N259 );
and g290 ( new_n441_, new_n439_, new_n440_ );
nand g291 ( new_n442_, new_n441_, keyIn_0_41 );
nor g292 ( new_n443_, new_n441_, keyIn_0_41 );
nand g293 ( new_n444_, new_n381_, N237 );
nand g294 ( new_n445_, new_n326_, N189 );
nand g295 ( new_n446_, N111, N210 );
and g296 ( new_n447_, new_n445_, new_n446_ );
nand g297 ( new_n448_, new_n447_, new_n444_ );
nor g298 ( new_n449_, new_n448_, new_n443_ );
nand g299 ( new_n450_, new_n449_, new_n442_ );
nand g300 ( new_n451_, new_n429_, N228 );
xor g301 ( new_n452_, new_n451_, keyIn_0_48 );
nor g302 ( new_n453_, new_n450_, new_n452_ );
nand g303 ( N864, new_n453_, new_n438_ );
not g304 ( new_n455_, new_n378_ );
or g305 ( new_n456_, new_n432_, new_n455_ );
nor g306 ( new_n457_, new_n455_, new_n369_ );
nor g307 ( new_n458_, new_n431_, new_n457_ );
nor g308 ( new_n459_, new_n458_, new_n308_ );
nand g309 ( new_n460_, new_n456_, new_n459_ );
and g310 ( new_n461_, new_n326_, N195 );
nand g311 ( new_n462_, new_n457_, N228 );
not g312 ( new_n463_, N237 );
nor g313 ( new_n464_, new_n378_, new_n463_ );
nand g314 ( new_n465_, new_n368_, N246 );
nand g315 ( new_n466_, N255, N260 );
nand g316 ( new_n467_, N116, N210 );
and g317 ( new_n468_, new_n466_, new_n467_ );
nand g318 ( new_n469_, new_n465_, new_n468_ );
nor g319 ( new_n470_, new_n464_, new_n469_ );
nand g320 ( new_n471_, new_n462_, new_n470_ );
nor g321 ( new_n472_, new_n461_, new_n471_ );
nand g322 ( N865, new_n460_, new_n472_ );
nor g323 ( new_n474_, new_n256_, N268 );
nand g324 ( new_n475_, new_n272_, new_n474_ );
nor g325 ( new_n476_, new_n475_, keyIn_0_18 );
and g326 ( new_n477_, N138, N152 );
nor g327 ( new_n478_, new_n476_, new_n477_ );
nor g328 ( new_n479_, new_n257_, new_n264_ );
and g329 ( new_n480_, new_n479_, N153 );
nand g330 ( new_n481_, new_n475_, keyIn_0_18 );
nand g331 ( new_n482_, new_n294_, N106 );
nand g332 ( new_n483_, new_n482_, new_n481_ );
nor g333 ( new_n484_, new_n483_, new_n480_ );
nand g334 ( new_n485_, new_n484_, new_n478_ );
nand g335 ( new_n486_, new_n485_, N177 );
or g336 ( new_n487_, new_n485_, N177 );
xnor g337 ( new_n488_, new_n398_, keyIn_0_40 );
nand g338 ( new_n489_, new_n488_, keyIn_0_46 );
not g339 ( new_n490_, keyIn_0_46 );
nand g340 ( new_n491_, new_n412_, new_n490_ );
nand g341 ( new_n492_, new_n489_, new_n491_ );
nand g342 ( new_n493_, new_n385_, new_n399_ );
nand g343 ( new_n494_, new_n493_, new_n492_ );
xnor g344 ( new_n495_, new_n494_, keyIn_0_54 );
nand g345 ( new_n496_, new_n495_, new_n487_ );
nand g346 ( new_n497_, new_n496_, new_n486_ );
nand g347 ( new_n498_, new_n479_, N149 );
nor g348 ( new_n499_, new_n498_, keyIn_0_17 );
nand g349 ( new_n500_, new_n498_, keyIn_0_17 );
nand g350 ( new_n501_, new_n294_, N101 );
not g351 ( new_n502_, new_n501_ );
nand g352 ( new_n503_, N17, N138 );
nand g353 ( new_n504_, new_n475_, new_n503_ );
nor g354 ( new_n505_, new_n502_, new_n504_ );
nand g355 ( new_n506_, new_n505_, new_n500_ );
nor g356 ( new_n507_, new_n506_, new_n499_ );
not g357 ( new_n508_, new_n507_ );
nor g358 ( new_n509_, new_n508_, N171 );
not g359 ( new_n510_, new_n509_ );
nand g360 ( new_n511_, new_n497_, new_n510_ );
nand g361 ( new_n512_, new_n508_, N171 );
xnor g362 ( new_n513_, new_n512_, keyIn_0_35 );
nand g363 ( new_n514_, new_n511_, new_n513_ );
not g364 ( new_n515_, keyIn_0_21 );
nand g365 ( new_n516_, new_n479_, N146 );
nand g366 ( new_n517_, new_n516_, new_n475_ );
nand g367 ( new_n518_, new_n517_, new_n515_ );
nor g368 ( new_n519_, new_n517_, new_n515_ );
nand g369 ( new_n520_, new_n294_, N96 );
nand g370 ( new_n521_, N51, N138 );
nand g371 ( new_n522_, new_n520_, new_n521_ );
nor g372 ( new_n523_, new_n519_, new_n522_ );
nand g373 ( new_n524_, new_n523_, new_n518_ );
not g374 ( new_n525_, new_n524_ );
nand g375 ( new_n526_, new_n525_, new_n228_ );
nand g376 ( new_n527_, new_n514_, new_n526_ );
nand g377 ( new_n528_, new_n524_, N165 );
nand g378 ( new_n529_, new_n527_, new_n528_ );
nand g379 ( new_n530_, new_n479_, N143 );
nand g380 ( new_n531_, new_n530_, new_n475_ );
nand g381 ( new_n532_, new_n531_, keyIn_0_20 );
nor g382 ( new_n533_, new_n531_, keyIn_0_20 );
nand g383 ( new_n534_, N8, N138 );
nand g384 ( new_n535_, new_n294_, N91 );
nand g385 ( new_n536_, new_n535_, new_n534_ );
nor g386 ( new_n537_, new_n533_, new_n536_ );
nand g387 ( new_n538_, new_n537_, new_n532_ );
not g388 ( new_n539_, new_n538_ );
nand g389 ( new_n540_, new_n539_, new_n227_ );
xor g390 ( new_n541_, new_n540_, keyIn_0_33 );
not g391 ( new_n542_, new_n541_ );
nand g392 ( new_n543_, new_n529_, new_n542_ );
nor g393 ( new_n544_, new_n539_, new_n227_ );
xor g394 ( new_n545_, new_n544_, keyIn_0_43 );
nand g395 ( new_n546_, new_n543_, new_n545_ );
xnor g396 ( N866, new_n546_, keyIn_0_59 );
not g397 ( new_n548_, keyIn_0_57 );
not g398 ( new_n549_, new_n495_ );
nand g399 ( new_n550_, new_n487_, new_n486_ );
nand g400 ( new_n551_, new_n549_, new_n550_ );
nor g401 ( new_n552_, new_n551_, new_n548_ );
nand g402 ( new_n553_, new_n551_, new_n548_ );
nor g403 ( new_n554_, new_n549_, new_n550_ );
nor g404 ( new_n555_, new_n554_, new_n308_ );
nand g405 ( new_n556_, new_n555_, new_n553_ );
nor g406 ( new_n557_, new_n556_, new_n552_ );
nand g407 ( new_n558_, new_n326_, N177 );
nor g408 ( new_n559_, new_n550_, new_n424_ );
nor g409 ( new_n560_, new_n486_, new_n463_ );
nand g410 ( new_n561_, new_n485_, N246 );
nand g411 ( new_n562_, N101, N210 );
nand g412 ( new_n563_, new_n561_, new_n562_ );
or g413 ( new_n564_, new_n560_, new_n563_ );
nor g414 ( new_n565_, new_n559_, new_n564_ );
nand g415 ( new_n566_, new_n558_, new_n565_ );
nor g416 ( new_n567_, new_n557_, new_n566_ );
xnor g417 ( N874, new_n567_, keyIn_0_62 );
or g418 ( new_n569_, new_n543_, new_n544_ );
nor g419 ( new_n570_, new_n541_, new_n544_ );
nor g420 ( new_n571_, new_n529_, new_n570_ );
nor g421 ( new_n572_, new_n571_, new_n308_ );
nand g422 ( new_n573_, new_n569_, new_n572_ );
nand g423 ( new_n574_, new_n570_, N228 );
and g424 ( new_n575_, new_n544_, N237 );
not g425 ( new_n576_, N210 );
nor g426 ( new_n577_, new_n260_, new_n576_ );
nor g427 ( new_n578_, new_n575_, new_n577_ );
nand g428 ( new_n579_, new_n574_, new_n578_ );
nand g429 ( new_n580_, new_n326_, N159 );
nand g430 ( new_n581_, new_n538_, N246 );
xor g431 ( new_n582_, new_n581_, keyIn_0_34 );
nand g432 ( new_n583_, new_n580_, new_n582_ );
xnor g433 ( new_n584_, new_n583_, keyIn_0_39 );
nor g434 ( new_n585_, new_n584_, new_n579_ );
nand g435 ( N878, new_n573_, new_n585_ );
nand g436 ( new_n587_, new_n526_, new_n528_ );
not g437 ( new_n588_, new_n587_ );
xnor g438 ( new_n589_, new_n513_, keyIn_0_44 );
nand g439 ( new_n590_, new_n511_, new_n589_ );
nor g440 ( new_n591_, new_n590_, new_n588_ );
nand g441 ( new_n592_, new_n591_, keyIn_0_58 );
nor g442 ( new_n593_, new_n591_, keyIn_0_58 );
nand g443 ( new_n594_, new_n590_, new_n588_ );
nand g444 ( new_n595_, new_n594_, N219 );
nor g445 ( new_n596_, new_n593_, new_n595_ );
nand g446 ( new_n597_, new_n596_, new_n592_ );
nand g447 ( new_n598_, N91, N210 );
xor g448 ( new_n599_, new_n598_, keyIn_0_7 );
nand g449 ( new_n600_, new_n597_, new_n599_ );
or g450 ( new_n601_, new_n600_, keyIn_0_60 );
nand g451 ( new_n602_, new_n600_, keyIn_0_60 );
nor g452 ( new_n603_, new_n587_, new_n424_ );
nand g453 ( new_n604_, new_n326_, N165 );
nor g454 ( new_n605_, new_n528_, new_n463_ );
nor g455 ( new_n606_, new_n525_, new_n330_ );
nor g456 ( new_n607_, new_n605_, new_n606_ );
nand g457 ( new_n608_, new_n604_, new_n607_ );
nor g458 ( new_n609_, new_n608_, new_n603_ );
and g459 ( new_n610_, new_n602_, new_n609_ );
nand g460 ( N879, new_n610_, new_n601_ );
not g461 ( new_n612_, keyIn_0_63 );
not g462 ( new_n613_, new_n513_ );
nor g463 ( new_n614_, new_n613_, new_n509_ );
nand g464 ( new_n615_, new_n497_, new_n614_ );
nor g465 ( new_n616_, new_n497_, new_n614_ );
nor g466 ( new_n617_, new_n616_, new_n308_ );
nand g467 ( new_n618_, new_n617_, new_n615_ );
nand g468 ( new_n619_, N96, N210 );
nand g469 ( new_n620_, new_n618_, new_n619_ );
xnor g470 ( new_n621_, new_n620_, keyIn_0_61 );
nand g471 ( new_n622_, new_n613_, N237 );
xnor g472 ( new_n623_, new_n622_, keyIn_0_45 );
and g473 ( new_n624_, new_n614_, N228 );
nand g474 ( new_n625_, new_n508_, N246 );
nand g475 ( new_n626_, new_n326_, N171 );
nand g476 ( new_n627_, new_n626_, new_n625_ );
nor g477 ( new_n628_, new_n624_, new_n627_ );
nand g478 ( new_n629_, new_n628_, new_n623_ );
nor g479 ( new_n630_, new_n621_, new_n629_ );
xnor g480 ( N880, new_n630_, new_n612_ );
endmodule