module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n445_, new_n699_, new_n236_, new_n1009_, new_n238_, new_n479_, new_n1105_, new_n955_, new_n608_, new_n847_, new_n250_, new_n888_, new_n501_, new_n288_, new_n1157_, new_n798_, new_n1180_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1048_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n1025_, new_n566_, new_n641_, new_n339_, new_n365_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n1176_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n1057_, new_n670_, new_n456_, new_n691_, new_n1024_, new_n1125_, new_n246_, new_n682_, new_n1075_, new_n812_, new_n911_, new_n679_, new_n937_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n1071_, new_n1131_, new_n1120_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n695_, new_n240_, new_n660_, new_n413_, new_n1060_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n1119_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n1045_, new_n1132_, new_n500_, new_n898_, new_n1163_, new_n786_, new_n799_, new_n946_, new_n317_, new_n1188_, new_n344_, new_n287_, new_n721_, new_n504_, new_n1108_, new_n862_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n1167_, new_n215_, new_n626_, new_n959_, new_n990_, new_n774_, new_n716_, new_n701_, new_n792_, new_n1058_, new_n953_, new_n257_, new_n1162_, new_n481_, new_n212_, new_n1073_, new_n1110_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n1059_, new_n634_, new_n414_, new_n1101_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n1050_, new_n903_, new_n230_, new_n983_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n1151_, new_n1082_, new_n849_, new_n1018_, new_n855_, new_n606_, new_n1037_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n1054_, new_n1083_, new_n385_, new_n1049_, new_n829_, new_n988_, new_n478_, new_n694_, new_n461_, new_n710_, new_n971_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n683_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n1184_, new_n517_, new_n325_, new_n609_, new_n1031_, new_n961_, new_n530_, new_n890_, new_n318_, new_n1006_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n1005_, new_n999_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n1086_, new_n956_, new_n763_, new_n960_, new_n1138_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n970_, new_n995_, new_n1035_, new_n271_, new_n674_, new_n274_, new_n991_, new_n1044_, new_n218_, new_n497_, new_n816_, new_n1170_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n1051_, new_n1053_, new_n423_, new_n205_, new_n492_, new_n498_, new_n496_, new_n1046_, new_n650_, new_n708_, new_n750_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n734_, new_n925_, new_n1062_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n256_, new_n778_, new_n452_, new_n381_, new_n656_, new_n1121_, new_n820_, new_n1127_, new_n771_, new_n388_, new_n979_, new_n1028_, new_n508_, new_n714_, new_n483_, new_n1004_, new_n1152_, new_n394_, new_n299_, new_n1007_, new_n882_, new_n657_, new_n1150_, new_n929_, new_n652_, new_n314_, new_n582_, new_n986_, new_n1020_, new_n363_, new_n1159_, new_n1113_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n917_, new_n1041_, new_n426_, new_n1036_, new_n235_, new_n1133_, new_n398_, new_n301_, new_n1177_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n1026_, new_n207_, new_n267_, new_n473_, new_n1147_, new_n790_, new_n1081_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n969_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n996_, new_n621_, new_n846_, new_n915_, new_n349_, new_n244_, new_n488_, new_n524_, new_n705_, new_n277_, new_n848_, new_n874_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n438_, new_n1003_, new_n696_, new_n208_, new_n632_, new_n1039_, new_n671_, new_n965_, new_n528_, new_n952_, new_n1158_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n397_, new_n729_, new_n1111_, new_n975_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n1115_, new_n559_, new_n948_, new_n762_, new_n1055_, new_n1193_, new_n838_, new_n923_, new_n233_, new_n1187_, new_n469_, new_n391_, new_n1154_, new_n437_, new_n1085_, new_n295_, new_n359_, new_n794_, new_n628_, new_n409_, new_n1090_, new_n745_, new_n457_, new_n553_, new_n1084_, new_n1061_, new_n668_, new_n333_, new_n1128_, new_n1002_, new_n290_, new_n834_, new_n1169_, new_n369_, new_n448_, new_n867_, new_n1032_, new_n901_, new_n1171_, new_n276_, new_n688_, new_n384_, new_n900_, new_n1161_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n1096_, new_n454_, new_n202_, new_n1034_, new_n296_, new_n661_, new_n1124_, new_n308_, new_n1000_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n1070_, new_n1109_, new_n860_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n938_, new_n1166_, new_n809_, new_n1142_, new_n654_, new_n713_, new_n880_, new_n1102_, new_n604_, new_n227_, new_n1104_, new_n690_, new_n416_, new_n222_, new_n1043_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n1136_, new_n693_, new_n1175_, new_n505_, new_n619_, new_n471_, new_n967_, new_n268_, new_n374_, new_n577_, new_n1135_, new_n376_, new_n380_, new_n1079_, new_n747_, new_n749_, new_n861_, new_n1091_, new_n310_, new_n1095_, new_n275_, new_n998_, new_n1056_, new_n352_, new_n1094_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n1064_, new_n1065_, new_n1118_, new_n493_, new_n547_, new_n907_, new_n264_, new_n665_, new_n800_, new_n379_, new_n897_, new_n1012_, new_n719_, new_n869_, new_n273_, new_n1178_, new_n224_, new_n586_, new_n963_, new_n270_, new_n570_, new_n598_, new_n893_, new_n993_, new_n1063_, new_n1191_, new_n824_, new_n520_, new_n1001_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n557_, new_n260_, new_n936_, new_n251_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1016_, new_n1074_, new_n748_, new_n1144_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n807_, new_n736_, new_n879_, new_n513_, new_n592_, new_n726_, new_n1123_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n1080_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n487_, new_n360_, new_n675_, new_n1126_, new_n1155_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n302_, new_n755_, new_n225_, new_n1040_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n1179_, new_n298_, new_n499_, new_n255_, new_n533_, new_n1088_, new_n1130_, new_n1148_, new_n795_, new_n1146_, new_n459_, new_n569_, new_n555_, new_n468_, new_n977_, new_n1139_, new_n782_, new_n1185_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n1174_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n972_, new_n1067_, new_n891_, new_n631_, new_n453_, new_n516_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n1076_, new_n252_, new_n585_, new_n751_, new_n312_, new_n535_, new_n1038_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n1181_, new_n597_, new_n978_, new_n1093_, new_n1092_, new_n408_, new_n1143_, new_n470_, new_n213_, new_n1072_, new_n769_, new_n1097_, new_n1069_, new_n651_, new_n433_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n265_, new_n732_, new_n687_, new_n370_, new_n1029_, new_n689_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n1052_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n989_, new_n1117_, new_n1112_, new_n711_, new_n1156_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n1116_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n327_, new_n681_, new_n1087_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n319_, new_n1008_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n957_, new_n754_, new_n1047_, new_n787_, new_n653_, new_n1134_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n330_, new_n727_, new_n375_, new_n294_, new_n760_, new_n627_, new_n1173_, new_n704_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n1189_, new_n1153_, new_n357_, new_n320_, new_n780_, new_n1183_, new_n245_, new_n643_, new_n474_, new_n1129_, new_n467_, new_n1013_, new_n404_, new_n1077_, new_n490_, new_n560_, new_n1100_, new_n865_, new_n1027_, new_n358_, new_n877_, new_n348_, new_n610_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n1011_, new_n1165_, new_n425_, new_n896_, new_n226_, new_n802_, new_n697_, new_n1099_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n866_, new_n540_, new_n1066_, new_n434_, new_n947_, new_n994_, new_n982_, new_n422_, new_n964_, new_n1078_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n551_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n1140_, new_n521_, new_n1042_, new_n793_, new_n863_, new_n406_, new_n828_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n1089_, new_n1192_, new_n573_, new_n765_, new_n405_, new_n1103_;

not g000 ( new_n202_, N1 );
not g001 ( new_n203_, keyIn_0_64 );
not g002 ( new_n204_, keyIn_0_60 );
not g003 ( new_n205_, N81 );
not g004 ( new_n206_, N85 );
nand g005 ( new_n207_, new_n205_, new_n206_ );
nand g006 ( new_n208_, N81, N85 );
nand g007 ( new_n209_, new_n207_, new_n208_ );
nand g008 ( new_n210_, new_n209_, keyIn_0_10 );
not g009 ( new_n211_, keyIn_0_10 );
nand g010 ( new_n212_, new_n207_, new_n211_, new_n208_ );
not g011 ( new_n213_, N89 );
not g012 ( new_n214_, N93 );
nand g013 ( new_n215_, new_n213_, new_n214_ );
nand g014 ( new_n216_, N89, N93 );
nand g015 ( new_n217_, new_n215_, new_n216_ );
nand g016 ( new_n218_, new_n217_, keyIn_0_11 );
not g017 ( new_n219_, keyIn_0_11 );
nand g018 ( new_n220_, new_n215_, new_n219_, new_n216_ );
nand g019 ( new_n221_, new_n210_, new_n218_, new_n212_, new_n220_ );
nand g020 ( new_n222_, new_n210_, new_n212_ );
nand g021 ( new_n223_, new_n218_, new_n220_ );
nand g022 ( new_n224_, new_n222_, new_n223_ );
nand g023 ( new_n225_, new_n224_, new_n221_ );
nand g024 ( new_n226_, new_n225_, keyIn_0_45 );
not g025 ( new_n227_, keyIn_0_45 );
nand g026 ( new_n228_, new_n224_, new_n227_, new_n221_ );
not g027 ( new_n229_, keyIn_0_44 );
not g028 ( new_n230_, N65 );
not g029 ( new_n231_, N69 );
nand g030 ( new_n232_, new_n230_, new_n231_ );
nand g031 ( new_n233_, N65, N69 );
nand g032 ( new_n234_, new_n232_, new_n233_ );
nand g033 ( new_n235_, new_n234_, keyIn_0_8 );
not g034 ( new_n236_, keyIn_0_8 );
nand g035 ( new_n237_, new_n232_, new_n236_, new_n233_ );
not g036 ( new_n238_, N73 );
not g037 ( new_n239_, N77 );
nand g038 ( new_n240_, new_n238_, new_n239_ );
nand g039 ( new_n241_, N73, N77 );
nand g040 ( new_n242_, new_n240_, new_n241_ );
nand g041 ( new_n243_, new_n242_, keyIn_0_9 );
not g042 ( new_n244_, keyIn_0_9 );
nand g043 ( new_n245_, new_n240_, new_n244_, new_n241_ );
nand g044 ( new_n246_, new_n235_, new_n243_, new_n237_, new_n245_ );
nand g045 ( new_n247_, new_n235_, new_n237_ );
nand g046 ( new_n248_, new_n243_, new_n245_ );
nand g047 ( new_n249_, new_n247_, new_n248_ );
nand g048 ( new_n250_, new_n249_, new_n246_ );
nand g049 ( new_n251_, new_n250_, new_n229_ );
nand g050 ( new_n252_, new_n249_, keyIn_0_44, new_n246_ );
nand g051 ( new_n253_, new_n226_, new_n251_, new_n228_, new_n252_ );
nand g052 ( new_n254_, new_n226_, new_n228_ );
nand g053 ( new_n255_, new_n251_, new_n252_ );
nand g054 ( new_n256_, new_n254_, new_n255_ );
nand g055 ( new_n257_, new_n256_, new_n204_, new_n253_ );
nand g056 ( new_n258_, new_n256_, new_n253_ );
nand g057 ( new_n259_, new_n258_, keyIn_0_60 );
nand g058 ( new_n260_, N129, N137 );
nand g059 ( new_n261_, new_n260_, keyIn_0_16 );
not g060 ( new_n262_, keyIn_0_16 );
nand g061 ( new_n263_, new_n262_, N129, N137 );
nand g062 ( new_n264_, new_n259_, new_n257_, new_n261_, new_n263_ );
nand g063 ( new_n265_, new_n259_, new_n257_ );
nand g064 ( new_n266_, new_n261_, new_n263_ );
nand g065 ( new_n267_, new_n265_, new_n266_ );
nand g066 ( new_n268_, new_n267_, new_n264_ );
nand g067 ( new_n269_, new_n268_, new_n203_ );
nand g068 ( new_n270_, new_n267_, keyIn_0_64, new_n264_ );
nand g069 ( new_n271_, new_n269_, new_n270_ );
nor g070 ( new_n272_, N1, N17 );
not g071 ( new_n273_, new_n272_ );
nand g072 ( new_n274_, N1, N17 );
nand g073 ( new_n275_, new_n273_, new_n274_ );
nand g074 ( new_n276_, new_n275_, keyIn_0_24 );
not g075 ( new_n277_, new_n276_ );
nor g076 ( new_n278_, new_n275_, keyIn_0_24 );
nor g077 ( new_n279_, new_n277_, new_n278_ );
not g078 ( new_n280_, new_n279_ );
nor g079 ( new_n281_, N33, N49 );
not g080 ( new_n282_, new_n281_ );
nand g081 ( new_n283_, N33, N49 );
nand g082 ( new_n284_, new_n282_, new_n283_ );
nand g083 ( new_n285_, new_n284_, keyIn_0_25 );
not g084 ( new_n286_, new_n285_ );
nor g085 ( new_n287_, new_n284_, keyIn_0_25 );
nor g086 ( new_n288_, new_n286_, new_n287_ );
not g087 ( new_n289_, new_n288_ );
nand g088 ( new_n290_, new_n280_, new_n289_ );
nand g089 ( new_n291_, new_n279_, new_n288_ );
nand g090 ( new_n292_, new_n290_, new_n291_ );
nand g091 ( new_n293_, new_n292_, keyIn_0_48 );
not g092 ( new_n294_, keyIn_0_48 );
nand g093 ( new_n295_, new_n290_, new_n294_, new_n291_ );
nand g094 ( new_n296_, new_n293_, new_n295_ );
not g095 ( new_n297_, new_n296_ );
nand g096 ( new_n298_, new_n271_, new_n297_ );
nand g097 ( new_n299_, new_n269_, new_n270_, new_n296_ );
nand g098 ( new_n300_, new_n298_, keyIn_0_72, new_n299_ );
not g099 ( new_n301_, keyIn_0_72 );
nand g100 ( new_n302_, new_n298_, new_n299_ );
nand g101 ( new_n303_, new_n302_, new_n301_ );
nand g102 ( new_n304_, new_n303_, new_n300_ );
not g103 ( new_n305_, new_n304_ );
not g104 ( new_n306_, keyIn_0_82 );
not g105 ( new_n307_, keyIn_0_74 );
not g106 ( new_n308_, keyIn_0_66 );
not g107 ( new_n309_, keyIn_0_62 );
not g108 ( new_n310_, N97 );
not g109 ( new_n311_, N101 );
nand g110 ( new_n312_, new_n310_, new_n311_ );
nand g111 ( new_n313_, N97, N101 );
nand g112 ( new_n314_, new_n312_, new_n313_ );
nand g113 ( new_n315_, new_n314_, keyIn_0_12 );
not g114 ( new_n316_, keyIn_0_12 );
nand g115 ( new_n317_, new_n312_, new_n316_, new_n313_ );
not g116 ( new_n318_, N105 );
not g117 ( new_n319_, N109 );
nand g118 ( new_n320_, new_n318_, new_n319_ );
nand g119 ( new_n321_, N105, N109 );
nand g120 ( new_n322_, new_n320_, new_n321_ );
nand g121 ( new_n323_, new_n322_, keyIn_0_13 );
not g122 ( new_n324_, keyIn_0_13 );
nand g123 ( new_n325_, new_n320_, new_n324_, new_n321_ );
nand g124 ( new_n326_, new_n315_, new_n323_, new_n317_, new_n325_ );
nand g125 ( new_n327_, new_n315_, new_n317_ );
nand g126 ( new_n328_, new_n323_, new_n325_ );
nand g127 ( new_n329_, new_n327_, new_n328_ );
nand g128 ( new_n330_, new_n329_, keyIn_0_46, new_n326_ );
not g129 ( new_n331_, keyIn_0_46 );
nand g130 ( new_n332_, new_n329_, new_n326_ );
nand g131 ( new_n333_, new_n332_, new_n331_ );
nand g132 ( new_n334_, new_n251_, new_n333_, new_n252_, new_n330_ );
nand g133 ( new_n335_, new_n333_, new_n330_ );
nand g134 ( new_n336_, new_n255_, new_n335_ );
nand g135 ( new_n337_, new_n336_, new_n309_, new_n334_ );
nand g136 ( new_n338_, new_n336_, new_n334_ );
nand g137 ( new_n339_, new_n338_, keyIn_0_62 );
nand g138 ( new_n340_, N131, N137 );
nand g139 ( new_n341_, new_n340_, keyIn_0_18 );
not g140 ( new_n342_, keyIn_0_18 );
nand g141 ( new_n343_, new_n342_, N131, N137 );
nand g142 ( new_n344_, new_n339_, new_n337_, new_n341_, new_n343_ );
nand g143 ( new_n345_, new_n339_, new_n337_ );
nand g144 ( new_n346_, new_n341_, new_n343_ );
nand g145 ( new_n347_, new_n345_, new_n346_ );
nand g146 ( new_n348_, new_n347_, new_n344_ );
nand g147 ( new_n349_, new_n348_, new_n308_ );
nand g148 ( new_n350_, new_n347_, keyIn_0_66, new_n344_ );
nand g149 ( new_n351_, new_n349_, new_n350_ );
not g150 ( new_n352_, keyIn_0_50 );
not g151 ( new_n353_, N25 );
nand g152 ( new_n354_, new_n353_, N9 );
not g153 ( new_n355_, N9 );
nand g154 ( new_n356_, new_n355_, N25 );
nand g155 ( new_n357_, new_n354_, new_n356_ );
nand g156 ( new_n358_, new_n357_, keyIn_0_28 );
not g157 ( new_n359_, keyIn_0_28 );
nand g158 ( new_n360_, new_n354_, new_n356_, new_n359_ );
nand g159 ( new_n361_, new_n358_, new_n360_ );
nor g160 ( new_n362_, N41, N57 );
not g161 ( new_n363_, new_n362_ );
nand g162 ( new_n364_, N41, N57 );
nand g163 ( new_n365_, new_n363_, new_n364_ );
nand g164 ( new_n366_, new_n365_, keyIn_0_29 );
not g165 ( new_n367_, new_n366_ );
nor g166 ( new_n368_, new_n365_, keyIn_0_29 );
nor g167 ( new_n369_, new_n367_, new_n368_ );
not g168 ( new_n370_, new_n369_ );
nand g169 ( new_n371_, new_n370_, new_n361_ );
nand g170 ( new_n372_, new_n369_, new_n358_, new_n360_ );
nand g171 ( new_n373_, new_n371_, new_n372_ );
nand g172 ( new_n374_, new_n373_, new_n352_ );
nand g173 ( new_n375_, new_n371_, keyIn_0_50, new_n372_ );
nand g174 ( new_n376_, new_n374_, new_n375_ );
not g175 ( new_n377_, new_n376_ );
nand g176 ( new_n378_, new_n351_, new_n377_ );
nand g177 ( new_n379_, new_n349_, new_n350_, new_n376_ );
nand g178 ( new_n380_, new_n378_, new_n379_ );
nand g179 ( new_n381_, new_n380_, new_n307_ );
nand g180 ( new_n382_, new_n378_, keyIn_0_74, new_n379_ );
nand g181 ( new_n383_, new_n381_, new_n306_, new_n382_ );
not g182 ( new_n384_, keyIn_0_75 );
not g183 ( new_n385_, keyIn_0_63 );
not g184 ( new_n386_, keyIn_0_47 );
not g185 ( new_n387_, keyIn_0_14 );
not g186 ( new_n388_, N113 );
not g187 ( new_n389_, N117 );
nand g188 ( new_n390_, new_n388_, new_n389_ );
nand g189 ( new_n391_, N113, N117 );
nand g190 ( new_n392_, new_n390_, new_n391_ );
nand g191 ( new_n393_, new_n392_, new_n387_ );
nand g192 ( new_n394_, new_n390_, keyIn_0_14, new_n391_ );
not g193 ( new_n395_, N121 );
not g194 ( new_n396_, N125 );
nand g195 ( new_n397_, new_n395_, new_n396_ );
nand g196 ( new_n398_, N121, N125 );
nand g197 ( new_n399_, new_n397_, new_n398_ );
nand g198 ( new_n400_, new_n399_, keyIn_0_15 );
not g199 ( new_n401_, keyIn_0_15 );
nand g200 ( new_n402_, new_n397_, new_n401_, new_n398_ );
nand g201 ( new_n403_, new_n393_, new_n400_, new_n394_, new_n402_ );
nand g202 ( new_n404_, new_n393_, new_n394_ );
nand g203 ( new_n405_, new_n400_, new_n402_ );
nand g204 ( new_n406_, new_n404_, new_n405_ );
nand g205 ( new_n407_, new_n406_, new_n403_ );
nand g206 ( new_n408_, new_n407_, new_n386_ );
nand g207 ( new_n409_, new_n406_, keyIn_0_47, new_n403_ );
nand g208 ( new_n410_, new_n226_, new_n408_, new_n228_, new_n409_ );
nand g209 ( new_n411_, new_n408_, new_n409_ );
nand g210 ( new_n412_, new_n254_, new_n411_ );
nand g211 ( new_n413_, new_n412_, new_n385_, new_n410_ );
nand g212 ( new_n414_, new_n412_, new_n410_ );
nand g213 ( new_n415_, new_n414_, keyIn_0_63 );
nand g214 ( new_n416_, N132, N137 );
nand g215 ( new_n417_, new_n416_, keyIn_0_19 );
not g216 ( new_n418_, keyIn_0_19 );
nand g217 ( new_n419_, new_n418_, N132, N137 );
nand g218 ( new_n420_, new_n415_, new_n413_, new_n417_, new_n419_ );
nand g219 ( new_n421_, new_n415_, new_n413_ );
nand g220 ( new_n422_, new_n417_, new_n419_ );
nand g221 ( new_n423_, new_n421_, new_n422_ );
nand g222 ( new_n424_, new_n423_, new_n420_ );
nand g223 ( new_n425_, new_n424_, keyIn_0_67 );
not g224 ( new_n426_, keyIn_0_67 );
nand g225 ( new_n427_, new_n423_, new_n426_, new_n420_ );
nand g226 ( new_n428_, new_n425_, new_n427_ );
not g227 ( new_n429_, N29 );
nand g228 ( new_n430_, new_n429_, N13 );
not g229 ( new_n431_, N13 );
nand g230 ( new_n432_, new_n431_, N29 );
nand g231 ( new_n433_, new_n430_, new_n432_ );
nand g232 ( new_n434_, new_n433_, keyIn_0_30 );
not g233 ( new_n435_, keyIn_0_30 );
nand g234 ( new_n436_, new_n430_, new_n432_, new_n435_ );
nand g235 ( new_n437_, new_n434_, new_n436_ );
not g236 ( new_n438_, N61 );
nand g237 ( new_n439_, new_n438_, N45 );
not g238 ( new_n440_, N45 );
nand g239 ( new_n441_, new_n440_, N61 );
nand g240 ( new_n442_, new_n439_, new_n441_ );
nand g241 ( new_n443_, new_n442_, keyIn_0_31 );
not g242 ( new_n444_, keyIn_0_31 );
nand g243 ( new_n445_, new_n439_, new_n441_, new_n444_ );
nand g244 ( new_n446_, new_n443_, new_n445_ );
nand g245 ( new_n447_, new_n437_, new_n446_ );
nand g246 ( new_n448_, new_n434_, new_n443_, new_n436_, new_n445_ );
nand g247 ( new_n449_, new_n447_, new_n448_ );
nand g248 ( new_n450_, new_n449_, keyIn_0_51 );
not g249 ( new_n451_, keyIn_0_51 );
nand g250 ( new_n452_, new_n447_, new_n451_, new_n448_ );
nand g251 ( new_n453_, new_n450_, new_n452_ );
nand g252 ( new_n454_, new_n428_, new_n453_ );
nand g253 ( new_n455_, new_n425_, new_n427_, new_n450_, new_n452_ );
nand g254 ( new_n456_, new_n454_, new_n455_ );
nand g255 ( new_n457_, new_n456_, new_n384_ );
nand g256 ( new_n458_, new_n454_, keyIn_0_75, new_n455_ );
nand g257 ( new_n459_, new_n457_, new_n458_ );
not g258 ( new_n460_, new_n459_ );
nand g259 ( new_n461_, new_n381_, new_n382_ );
nand g260 ( new_n462_, new_n461_, keyIn_0_82 );
nand g261 ( new_n463_, new_n462_, new_n383_, new_n460_ );
not g262 ( new_n464_, new_n463_ );
not g263 ( new_n465_, keyIn_0_81 );
not g264 ( new_n466_, keyIn_0_61 );
nand g265 ( new_n467_, new_n333_, new_n408_, new_n330_, new_n409_ );
nand g266 ( new_n468_, new_n335_, new_n411_ );
nand g267 ( new_n469_, new_n468_, new_n466_, new_n467_ );
nand g268 ( new_n470_, new_n468_, new_n467_ );
nand g269 ( new_n471_, new_n470_, keyIn_0_61 );
nand g270 ( new_n472_, N130, N137 );
nand g271 ( new_n473_, new_n472_, keyIn_0_17 );
not g272 ( new_n474_, keyIn_0_17 );
nand g273 ( new_n475_, new_n474_, N130, N137 );
nand g274 ( new_n476_, new_n471_, new_n469_, new_n473_, new_n475_ );
nand g275 ( new_n477_, new_n471_, new_n469_ );
nand g276 ( new_n478_, new_n473_, new_n475_ );
nand g277 ( new_n479_, new_n477_, new_n478_ );
nand g278 ( new_n480_, new_n479_, keyIn_0_65, new_n476_ );
not g279 ( new_n481_, keyIn_0_65 );
nand g280 ( new_n482_, new_n479_, new_n476_ );
nand g281 ( new_n483_, new_n482_, new_n481_ );
nand g282 ( new_n484_, new_n483_, new_n480_ );
nor g283 ( new_n485_, N5, N21 );
not g284 ( new_n486_, new_n485_ );
nand g285 ( new_n487_, N5, N21 );
nand g286 ( new_n488_, new_n486_, new_n487_ );
nand g287 ( new_n489_, new_n488_, keyIn_0_26 );
not g288 ( new_n490_, new_n489_ );
nor g289 ( new_n491_, new_n488_, keyIn_0_26 );
nor g290 ( new_n492_, new_n490_, new_n491_ );
not g291 ( new_n493_, new_n492_ );
nor g292 ( new_n494_, N37, N53 );
not g293 ( new_n495_, new_n494_ );
nand g294 ( new_n496_, N37, N53 );
nand g295 ( new_n497_, new_n495_, new_n496_ );
nand g296 ( new_n498_, new_n497_, keyIn_0_27 );
not g297 ( new_n499_, new_n498_ );
nor g298 ( new_n500_, new_n497_, keyIn_0_27 );
nor g299 ( new_n501_, new_n499_, new_n500_ );
not g300 ( new_n502_, new_n501_ );
nand g301 ( new_n503_, new_n493_, new_n502_ );
nand g302 ( new_n504_, new_n492_, new_n501_ );
nand g303 ( new_n505_, new_n503_, new_n504_ );
nand g304 ( new_n506_, new_n505_, keyIn_0_49 );
not g305 ( new_n507_, keyIn_0_49 );
nand g306 ( new_n508_, new_n503_, new_n507_, new_n504_ );
nand g307 ( new_n509_, new_n506_, new_n508_ );
nand g308 ( new_n510_, new_n484_, new_n509_ );
nand g309 ( new_n511_, new_n483_, new_n480_, new_n506_, new_n508_ );
nand g310 ( new_n512_, new_n510_, keyIn_0_73, new_n511_ );
not g311 ( new_n513_, keyIn_0_73 );
nand g312 ( new_n514_, new_n510_, new_n511_ );
nand g313 ( new_n515_, new_n514_, new_n513_ );
nand g314 ( new_n516_, new_n515_, new_n465_, new_n512_ );
nand g315 ( new_n517_, new_n515_, new_n512_ );
nand g316 ( new_n518_, new_n517_, keyIn_0_81 );
nand g317 ( new_n519_, new_n518_, new_n516_ );
not g318 ( new_n520_, keyIn_0_80 );
nand g319 ( new_n521_, new_n303_, new_n520_, new_n300_ );
nand g320 ( new_n522_, new_n304_, keyIn_0_80 );
nand g321 ( new_n523_, new_n522_, new_n521_ );
nand g322 ( new_n524_, new_n464_, new_n519_, new_n523_ );
nand g323 ( new_n525_, new_n524_, keyIn_0_104 );
not g324 ( new_n526_, new_n461_ );
not g325 ( new_n527_, keyIn_0_84 );
nand g326 ( new_n528_, new_n515_, new_n527_, new_n512_ );
nand g327 ( new_n529_, new_n517_, keyIn_0_84 );
nand g328 ( new_n530_, new_n529_, new_n526_, new_n528_ );
not g329 ( new_n531_, new_n530_ );
not g330 ( new_n532_, keyIn_0_85 );
nand g331 ( new_n533_, new_n457_, new_n532_, new_n458_ );
nand g332 ( new_n534_, new_n459_, keyIn_0_85 );
nand g333 ( new_n535_, new_n534_, new_n533_ );
nand g334 ( new_n536_, new_n303_, keyIn_0_83, new_n300_ );
not g335 ( new_n537_, keyIn_0_83 );
nand g336 ( new_n538_, new_n304_, new_n537_ );
nand g337 ( new_n539_, new_n538_, new_n536_ );
nand g338 ( new_n540_, new_n531_, new_n535_, new_n539_ );
nand g339 ( new_n541_, new_n540_, keyIn_0_105 );
nand g340 ( new_n542_, new_n525_, new_n541_ );
not g341 ( new_n543_, keyIn_0_105 );
nand g342 ( new_n544_, new_n535_, new_n539_ );
nor g343 ( new_n545_, new_n544_, new_n530_ );
nand g344 ( new_n546_, new_n545_, new_n543_ );
not g345 ( new_n547_, keyIn_0_104 );
nand g346 ( new_n548_, new_n519_, new_n523_ );
nor g347 ( new_n549_, new_n548_, new_n463_ );
nand g348 ( new_n550_, new_n549_, new_n547_ );
nand g349 ( new_n551_, new_n546_, new_n550_ );
nor g350 ( new_n552_, new_n551_, new_n542_ );
not g351 ( new_n553_, keyIn_0_86 );
nand g352 ( new_n554_, new_n304_, new_n553_ );
not g353 ( new_n555_, keyIn_0_87 );
nand g354 ( new_n556_, new_n381_, new_n555_, new_n382_ );
not g355 ( new_n557_, keyIn_0_88 );
nand g356 ( new_n558_, new_n457_, new_n557_, new_n458_ );
nand g357 ( new_n559_, new_n556_, new_n558_ );
not g358 ( new_n560_, new_n559_ );
not g359 ( new_n561_, new_n517_ );
nand g360 ( new_n562_, new_n459_, keyIn_0_88 );
nand g361 ( new_n563_, new_n303_, keyIn_0_86, new_n300_ );
nand g362 ( new_n564_, new_n461_, keyIn_0_87 );
nand g363 ( new_n565_, new_n562_, new_n564_, new_n561_, new_n563_ );
not g364 ( new_n566_, new_n565_ );
nand g365 ( new_n567_, new_n566_, new_n554_, new_n560_ );
nand g366 ( new_n568_, new_n567_, keyIn_0_106 );
not g367 ( new_n569_, keyIn_0_106 );
nand g368 ( new_n570_, new_n566_, new_n569_, new_n554_, new_n560_ );
nand g369 ( new_n571_, new_n568_, new_n570_ );
not g370 ( new_n572_, keyIn_0_107 );
not g371 ( new_n573_, keyIn_0_91 );
nand g372 ( new_n574_, new_n459_, new_n573_ );
not g373 ( new_n575_, new_n574_ );
not g374 ( new_n576_, keyIn_0_90 );
nand g375 ( new_n577_, new_n381_, new_n576_, new_n382_ );
nand g376 ( new_n578_, new_n457_, keyIn_0_91, new_n458_ );
nand g377 ( new_n579_, new_n577_, new_n578_ );
nor g378 ( new_n580_, new_n575_, new_n579_ );
not g379 ( new_n581_, keyIn_0_89 );
nand g380 ( new_n582_, new_n517_, new_n581_ );
nand g381 ( new_n583_, new_n515_, keyIn_0_89, new_n512_ );
nand g382 ( new_n584_, new_n461_, keyIn_0_90 );
nand g383 ( new_n585_, new_n582_, new_n584_, new_n305_, new_n583_ );
not g384 ( new_n586_, new_n585_ );
nand g385 ( new_n587_, new_n586_, new_n572_, new_n580_ );
nand g386 ( new_n588_, new_n586_, new_n580_ );
nand g387 ( new_n589_, new_n588_, keyIn_0_107 );
nand g388 ( new_n590_, new_n589_, new_n587_ );
nand g389 ( new_n591_, new_n552_, keyIn_0_112, new_n571_, new_n590_ );
not g390 ( new_n592_, keyIn_0_112 );
nor g391 ( new_n593_, new_n549_, new_n547_ );
nor g392 ( new_n594_, new_n545_, new_n543_ );
nor g393 ( new_n595_, new_n593_, new_n594_ );
nor g394 ( new_n596_, new_n540_, keyIn_0_105 );
nor g395 ( new_n597_, new_n548_, keyIn_0_104, new_n463_ );
nor g396 ( new_n598_, new_n596_, new_n597_ );
nand g397 ( new_n599_, new_n595_, new_n598_, new_n571_, new_n590_ );
nand g398 ( new_n600_, new_n599_, new_n592_ );
nand g399 ( new_n601_, new_n600_, new_n591_ );
not g400 ( new_n602_, new_n601_ );
not g401 ( new_n603_, keyIn_0_78 );
not g402 ( new_n604_, keyIn_0_70 );
not g403 ( new_n605_, keyIn_0_58 );
not g404 ( new_n606_, N5 );
nand g405 ( new_n607_, new_n202_, new_n606_ );
nand g406 ( new_n608_, N1, N5 );
nand g407 ( new_n609_, new_n607_, new_n608_ );
nand g408 ( new_n610_, new_n609_, keyIn_0_0 );
not g409 ( new_n611_, keyIn_0_0 );
nand g410 ( new_n612_, new_n607_, new_n611_, new_n608_ );
nand g411 ( new_n613_, new_n355_, new_n431_ );
nand g412 ( new_n614_, N9, N13 );
nand g413 ( new_n615_, new_n613_, new_n614_ );
nand g414 ( new_n616_, new_n615_, keyIn_0_1 );
not g415 ( new_n617_, keyIn_0_1 );
nand g416 ( new_n618_, new_n613_, new_n617_, new_n614_ );
nand g417 ( new_n619_, new_n610_, new_n616_, new_n612_, new_n618_ );
nand g418 ( new_n620_, new_n610_, new_n612_ );
nand g419 ( new_n621_, new_n616_, new_n618_ );
nand g420 ( new_n622_, new_n620_, new_n621_ );
nand g421 ( new_n623_, new_n622_, keyIn_0_40, new_n619_ );
not g422 ( new_n624_, keyIn_0_40 );
nand g423 ( new_n625_, new_n622_, new_n619_ );
nand g424 ( new_n626_, new_n625_, new_n624_ );
not g425 ( new_n627_, keyIn_0_42 );
not g426 ( new_n628_, N33 );
not g427 ( new_n629_, N37 );
nand g428 ( new_n630_, new_n628_, new_n629_ );
nand g429 ( new_n631_, N33, N37 );
nand g430 ( new_n632_, new_n630_, new_n631_ );
nand g431 ( new_n633_, new_n632_, keyIn_0_4 );
not g432 ( new_n634_, keyIn_0_4 );
nand g433 ( new_n635_, new_n630_, new_n634_, new_n631_ );
not g434 ( new_n636_, N41 );
nand g435 ( new_n637_, new_n636_, new_n440_ );
nand g436 ( new_n638_, N41, N45 );
nand g437 ( new_n639_, new_n637_, new_n638_ );
nand g438 ( new_n640_, new_n639_, keyIn_0_5 );
not g439 ( new_n641_, keyIn_0_5 );
nand g440 ( new_n642_, new_n637_, new_n641_, new_n638_ );
nand g441 ( new_n643_, new_n633_, new_n640_, new_n635_, new_n642_ );
nand g442 ( new_n644_, new_n633_, new_n635_ );
nand g443 ( new_n645_, new_n640_, new_n642_ );
nand g444 ( new_n646_, new_n644_, new_n645_ );
nand g445 ( new_n647_, new_n646_, new_n643_ );
nand g446 ( new_n648_, new_n647_, new_n627_ );
nand g447 ( new_n649_, new_n646_, keyIn_0_42, new_n643_ );
nand g448 ( new_n650_, new_n626_, new_n648_, new_n623_, new_n649_ );
nand g449 ( new_n651_, new_n626_, new_n623_ );
nand g450 ( new_n652_, new_n648_, new_n649_ );
nand g451 ( new_n653_, new_n651_, new_n652_ );
nand g452 ( new_n654_, new_n653_, new_n605_, new_n650_ );
nand g453 ( new_n655_, new_n653_, new_n650_ );
nand g454 ( new_n656_, new_n655_, keyIn_0_58 );
nand g455 ( new_n657_, N135, N137 );
nand g456 ( new_n658_, new_n657_, keyIn_0_22 );
not g457 ( new_n659_, keyIn_0_22 );
nand g458 ( new_n660_, new_n659_, N135, N137 );
nand g459 ( new_n661_, new_n656_, new_n654_, new_n658_, new_n660_ );
nand g460 ( new_n662_, new_n656_, new_n654_ );
nand g461 ( new_n663_, new_n658_, new_n660_ );
nand g462 ( new_n664_, new_n662_, new_n663_ );
nand g463 ( new_n665_, new_n664_, new_n661_ );
nand g464 ( new_n666_, new_n665_, new_n604_ );
nand g465 ( new_n667_, new_n664_, keyIn_0_70, new_n661_ );
nand g466 ( new_n668_, new_n666_, new_n667_ );
nand g467 ( new_n669_, new_n213_, N73 );
nand g468 ( new_n670_, new_n238_, N89 );
nand g469 ( new_n671_, new_n669_, new_n670_ );
nand g470 ( new_n672_, new_n671_, keyIn_0_36 );
not g471 ( new_n673_, keyIn_0_36 );
nand g472 ( new_n674_, new_n669_, new_n670_, new_n673_ );
nand g473 ( new_n675_, new_n672_, new_n674_ );
nor g474 ( new_n676_, N105, N121 );
not g475 ( new_n677_, new_n676_ );
nand g476 ( new_n678_, N105, N121 );
nand g477 ( new_n679_, new_n677_, new_n678_ );
nand g478 ( new_n680_, new_n679_, keyIn_0_37 );
not g479 ( new_n681_, new_n680_ );
nor g480 ( new_n682_, new_n679_, keyIn_0_37 );
nor g481 ( new_n683_, new_n681_, new_n682_ );
not g482 ( new_n684_, new_n683_ );
nand g483 ( new_n685_, new_n684_, new_n675_ );
nand g484 ( new_n686_, new_n683_, new_n672_, new_n674_ );
nand g485 ( new_n687_, new_n685_, new_n686_ );
nand g486 ( new_n688_, new_n687_, keyIn_0_54 );
not g487 ( new_n689_, keyIn_0_54 );
nand g488 ( new_n690_, new_n685_, new_n689_, new_n686_ );
nand g489 ( new_n691_, new_n688_, new_n690_ );
nand g490 ( new_n692_, new_n668_, new_n691_ );
nand g491 ( new_n693_, new_n666_, new_n667_, new_n688_, new_n690_ );
nand g492 ( new_n694_, new_n692_, new_n693_ );
nand g493 ( new_n695_, new_n694_, new_n603_ );
nand g494 ( new_n696_, new_n692_, keyIn_0_78, new_n693_ );
nand g495 ( new_n697_, new_n695_, new_n696_ );
not g496 ( new_n698_, new_n697_ );
not g497 ( new_n699_, keyIn_0_71 );
not g498 ( new_n700_, keyIn_0_59 );
not g499 ( new_n701_, keyIn_0_41 );
not g500 ( new_n702_, keyIn_0_2 );
not g501 ( new_n703_, N17 );
not g502 ( new_n704_, N21 );
nand g503 ( new_n705_, new_n703_, new_n704_ );
nand g504 ( new_n706_, N17, N21 );
nand g505 ( new_n707_, new_n705_, new_n706_ );
nand g506 ( new_n708_, new_n707_, new_n702_ );
nand g507 ( new_n709_, new_n705_, keyIn_0_2, new_n706_ );
nand g508 ( new_n710_, new_n353_, new_n429_ );
nand g509 ( new_n711_, N25, N29 );
nand g510 ( new_n712_, new_n710_, new_n711_ );
nand g511 ( new_n713_, new_n712_, keyIn_0_3 );
not g512 ( new_n714_, keyIn_0_3 );
nand g513 ( new_n715_, new_n710_, new_n714_, new_n711_ );
nand g514 ( new_n716_, new_n708_, new_n713_, new_n709_, new_n715_ );
nand g515 ( new_n717_, new_n708_, new_n709_ );
nand g516 ( new_n718_, new_n713_, new_n715_ );
nand g517 ( new_n719_, new_n717_, new_n718_ );
nand g518 ( new_n720_, new_n719_, new_n716_ );
nand g519 ( new_n721_, new_n720_, new_n701_ );
nand g520 ( new_n722_, new_n719_, keyIn_0_41, new_n716_ );
not g521 ( new_n723_, N49 );
not g522 ( new_n724_, N53 );
nand g523 ( new_n725_, new_n723_, new_n724_ );
nand g524 ( new_n726_, N49, N53 );
nand g525 ( new_n727_, new_n725_, new_n726_ );
nand g526 ( new_n728_, new_n727_, keyIn_0_6 );
not g527 ( new_n729_, keyIn_0_6 );
nand g528 ( new_n730_, new_n725_, new_n729_, new_n726_ );
not g529 ( new_n731_, N57 );
nand g530 ( new_n732_, new_n731_, new_n438_ );
nand g531 ( new_n733_, N57, N61 );
nand g532 ( new_n734_, new_n732_, new_n733_ );
nand g533 ( new_n735_, new_n734_, keyIn_0_7 );
not g534 ( new_n736_, keyIn_0_7 );
nand g535 ( new_n737_, new_n732_, new_n736_, new_n733_ );
nand g536 ( new_n738_, new_n728_, new_n735_, new_n730_, new_n737_ );
nand g537 ( new_n739_, new_n728_, new_n730_ );
nand g538 ( new_n740_, new_n735_, new_n737_ );
nand g539 ( new_n741_, new_n739_, new_n740_ );
nand g540 ( new_n742_, new_n741_, new_n738_ );
nand g541 ( new_n743_, new_n742_, keyIn_0_43 );
not g542 ( new_n744_, keyIn_0_43 );
nand g543 ( new_n745_, new_n741_, new_n744_, new_n738_ );
nand g544 ( new_n746_, new_n721_, new_n743_, new_n722_, new_n745_ );
nand g545 ( new_n747_, new_n721_, new_n722_ );
nand g546 ( new_n748_, new_n743_, new_n745_ );
nand g547 ( new_n749_, new_n747_, new_n748_ );
nand g548 ( new_n750_, new_n749_, new_n700_, new_n746_ );
nand g549 ( new_n751_, new_n749_, new_n746_ );
nand g550 ( new_n752_, new_n751_, keyIn_0_59 );
nand g551 ( new_n753_, N136, N137 );
nand g552 ( new_n754_, new_n753_, keyIn_0_23 );
not g553 ( new_n755_, keyIn_0_23 );
nand g554 ( new_n756_, new_n755_, N136, N137 );
nand g555 ( new_n757_, new_n752_, new_n750_, new_n754_, new_n756_ );
nand g556 ( new_n758_, new_n752_, new_n750_ );
nand g557 ( new_n759_, new_n754_, new_n756_ );
nand g558 ( new_n760_, new_n758_, new_n759_ );
nand g559 ( new_n761_, new_n760_, new_n757_ );
nand g560 ( new_n762_, new_n761_, new_n699_ );
nand g561 ( new_n763_, new_n760_, keyIn_0_71, new_n757_ );
nand g562 ( new_n764_, new_n762_, new_n763_ );
not g563 ( new_n765_, keyIn_0_55 );
nor g564 ( new_n766_, N77, N93 );
not g565 ( new_n767_, new_n766_ );
nand g566 ( new_n768_, N77, N93 );
nand g567 ( new_n769_, new_n767_, new_n768_ );
nand g568 ( new_n770_, new_n769_, keyIn_0_38 );
not g569 ( new_n771_, new_n770_ );
nor g570 ( new_n772_, new_n769_, keyIn_0_38 );
nor g571 ( new_n773_, new_n771_, new_n772_ );
not g572 ( new_n774_, new_n773_ );
nor g573 ( new_n775_, N109, N125 );
not g574 ( new_n776_, new_n775_ );
nand g575 ( new_n777_, N109, N125 );
nand g576 ( new_n778_, new_n776_, new_n777_ );
nand g577 ( new_n779_, new_n778_, keyIn_0_39 );
not g578 ( new_n780_, new_n779_ );
nor g579 ( new_n781_, new_n778_, keyIn_0_39 );
nor g580 ( new_n782_, new_n780_, new_n781_ );
not g581 ( new_n783_, new_n782_ );
nand g582 ( new_n784_, new_n774_, new_n783_ );
nand g583 ( new_n785_, new_n773_, new_n782_ );
nand g584 ( new_n786_, new_n784_, new_n785_ );
nand g585 ( new_n787_, new_n786_, new_n765_ );
nand g586 ( new_n788_, new_n784_, keyIn_0_55, new_n785_ );
nand g587 ( new_n789_, new_n787_, new_n788_ );
not g588 ( new_n790_, new_n789_ );
nand g589 ( new_n791_, new_n764_, new_n790_ );
nand g590 ( new_n792_, new_n762_, new_n763_, new_n789_ );
nand g591 ( new_n793_, new_n791_, keyIn_0_79, new_n792_ );
not g592 ( new_n794_, keyIn_0_79 );
nand g593 ( new_n795_, new_n791_, new_n792_ );
nand g594 ( new_n796_, new_n795_, new_n794_ );
nand g595 ( new_n797_, new_n796_, new_n793_ );
nor g596 ( new_n798_, new_n698_, new_n797_ );
not g597 ( new_n799_, keyIn_0_76 );
not g598 ( new_n800_, keyIn_0_56 );
nand g599 ( new_n801_, new_n626_, new_n721_, new_n623_, new_n722_ );
nand g600 ( new_n802_, new_n651_, new_n747_ );
nand g601 ( new_n803_, new_n802_, new_n800_, new_n801_ );
nand g602 ( new_n804_, new_n802_, new_n801_ );
nand g603 ( new_n805_, new_n804_, keyIn_0_56 );
nand g604 ( new_n806_, N133, N137 );
nand g605 ( new_n807_, new_n806_, keyIn_0_20 );
not g606 ( new_n808_, keyIn_0_20 );
nand g607 ( new_n809_, new_n808_, N133, N137 );
nand g608 ( new_n810_, new_n805_, new_n803_, new_n807_, new_n809_ );
nand g609 ( new_n811_, new_n805_, new_n803_ );
nand g610 ( new_n812_, new_n807_, new_n809_ );
nand g611 ( new_n813_, new_n811_, new_n812_ );
nand g612 ( new_n814_, new_n813_, new_n810_ );
nand g613 ( new_n815_, new_n814_, keyIn_0_68 );
not g614 ( new_n816_, keyIn_0_68 );
nand g615 ( new_n817_, new_n813_, new_n816_, new_n810_ );
nand g616 ( new_n818_, new_n815_, new_n817_ );
not g617 ( new_n819_, keyIn_0_52 );
nand g618 ( new_n820_, new_n205_, N65 );
nand g619 ( new_n821_, new_n230_, N81 );
nand g620 ( new_n822_, new_n820_, new_n821_ );
nand g621 ( new_n823_, new_n822_, keyIn_0_32 );
not g622 ( new_n824_, keyIn_0_32 );
nand g623 ( new_n825_, new_n820_, new_n821_, new_n824_ );
nand g624 ( new_n826_, new_n823_, new_n825_ );
nor g625 ( new_n827_, N97, N113 );
not g626 ( new_n828_, new_n827_ );
nand g627 ( new_n829_, N97, N113 );
nand g628 ( new_n830_, new_n828_, new_n829_ );
nand g629 ( new_n831_, new_n830_, keyIn_0_33 );
not g630 ( new_n832_, new_n831_ );
nor g631 ( new_n833_, new_n830_, keyIn_0_33 );
nor g632 ( new_n834_, new_n832_, new_n833_ );
not g633 ( new_n835_, new_n834_ );
nand g634 ( new_n836_, new_n835_, new_n826_ );
nand g635 ( new_n837_, new_n834_, new_n823_, new_n825_ );
nand g636 ( new_n838_, new_n836_, new_n837_ );
nand g637 ( new_n839_, new_n838_, new_n819_ );
nand g638 ( new_n840_, new_n836_, keyIn_0_52, new_n837_ );
nand g639 ( new_n841_, new_n839_, new_n840_ );
nand g640 ( new_n842_, new_n818_, new_n841_ );
nand g641 ( new_n843_, new_n815_, new_n817_, new_n839_, new_n840_ );
nand g642 ( new_n844_, new_n842_, new_n843_ );
nand g643 ( new_n845_, new_n844_, new_n799_ );
nand g644 ( new_n846_, new_n842_, keyIn_0_76, new_n843_ );
nand g645 ( new_n847_, new_n845_, new_n846_ );
not g646 ( new_n848_, new_n847_ );
not g647 ( new_n849_, keyIn_0_57 );
nand g648 ( new_n850_, new_n648_, new_n743_, new_n649_, new_n745_ );
nand g649 ( new_n851_, new_n652_, new_n748_ );
nand g650 ( new_n852_, new_n851_, new_n849_, new_n850_ );
nand g651 ( new_n853_, new_n851_, new_n850_ );
nand g652 ( new_n854_, new_n853_, keyIn_0_57 );
nand g653 ( new_n855_, N134, N137 );
nand g654 ( new_n856_, new_n855_, keyIn_0_21 );
not g655 ( new_n857_, keyIn_0_21 );
nand g656 ( new_n858_, new_n857_, N134, N137 );
nand g657 ( new_n859_, new_n854_, new_n852_, new_n856_, new_n858_ );
nand g658 ( new_n860_, new_n854_, new_n852_ );
nand g659 ( new_n861_, new_n856_, new_n858_ );
nand g660 ( new_n862_, new_n860_, new_n861_ );
nand g661 ( new_n863_, new_n862_, new_n859_ );
nand g662 ( new_n864_, new_n863_, keyIn_0_69 );
not g663 ( new_n865_, keyIn_0_69 );
nand g664 ( new_n866_, new_n862_, new_n865_, new_n859_ );
nand g665 ( new_n867_, new_n864_, new_n866_ );
not g666 ( new_n868_, keyIn_0_53 );
nand g667 ( new_n869_, new_n389_, N101 );
nand g668 ( new_n870_, new_n311_, N117 );
nand g669 ( new_n871_, new_n869_, new_n870_ );
nand g670 ( new_n872_, new_n871_, keyIn_0_35 );
not g671 ( new_n873_, keyIn_0_35 );
nand g672 ( new_n874_, new_n869_, new_n870_, new_n873_ );
nand g673 ( new_n875_, new_n872_, new_n874_ );
nor g674 ( new_n876_, N69, N85 );
not g675 ( new_n877_, new_n876_ );
nand g676 ( new_n878_, N69, N85 );
nand g677 ( new_n879_, new_n877_, new_n878_ );
nand g678 ( new_n880_, new_n879_, keyIn_0_34 );
not g679 ( new_n881_, new_n880_ );
nor g680 ( new_n882_, new_n879_, keyIn_0_34 );
nor g681 ( new_n883_, new_n881_, new_n882_ );
not g682 ( new_n884_, new_n883_ );
nand g683 ( new_n885_, new_n884_, new_n875_ );
nand g684 ( new_n886_, new_n883_, new_n872_, new_n874_ );
nand g685 ( new_n887_, new_n885_, new_n886_ );
nand g686 ( new_n888_, new_n887_, new_n868_ );
nand g687 ( new_n889_, new_n885_, keyIn_0_53, new_n886_ );
nand g688 ( new_n890_, new_n888_, new_n889_ );
nand g689 ( new_n891_, new_n867_, new_n890_ );
nand g690 ( new_n892_, new_n864_, new_n866_, new_n888_, new_n889_ );
nand g691 ( new_n893_, new_n891_, keyIn_0_77, new_n892_ );
not g692 ( new_n894_, keyIn_0_77 );
nand g693 ( new_n895_, new_n891_, new_n892_ );
nand g694 ( new_n896_, new_n895_, new_n894_ );
nand g695 ( new_n897_, new_n896_, new_n893_ );
nor g696 ( new_n898_, new_n848_, new_n897_ );
nand g697 ( new_n899_, new_n602_, new_n798_, new_n898_ );
nand g698 ( new_n900_, new_n899_, keyIn_0_114 );
not g699 ( new_n901_, keyIn_0_114 );
nor g700 ( new_n902_, new_n601_, new_n698_, new_n797_ );
nand g701 ( new_n903_, new_n902_, new_n901_, new_n898_ );
nand g702 ( new_n904_, new_n900_, new_n903_ );
nand g703 ( new_n905_, new_n904_, new_n202_, new_n305_ );
nand g704 ( new_n906_, new_n904_, new_n305_ );
nand g705 ( new_n907_, new_n906_, N1 );
nand g706 ( N724, new_n907_, new_n905_ );
nand g707 ( new_n909_, new_n904_, new_n606_, new_n561_ );
nand g708 ( new_n910_, new_n904_, new_n561_ );
nand g709 ( new_n911_, new_n910_, N5 );
nand g710 ( N725, new_n911_, new_n909_ );
nand g711 ( new_n913_, new_n904_, new_n355_, new_n526_ );
nand g712 ( new_n914_, new_n904_, new_n526_ );
nand g713 ( new_n915_, new_n914_, N9 );
nand g714 ( N726, new_n915_, new_n913_ );
nand g715 ( new_n917_, new_n904_, new_n431_, new_n460_ );
nand g716 ( new_n918_, new_n904_, new_n460_ );
nand g717 ( new_n919_, new_n918_, N13 );
nand g718 ( N727, new_n919_, new_n917_ );
nand g719 ( new_n921_, new_n698_, new_n797_ );
nor g720 ( new_n922_, new_n921_, new_n848_, new_n897_ );
nand g721 ( new_n923_, new_n602_, keyIn_0_115, new_n922_ );
not g722 ( new_n924_, keyIn_0_115 );
nand g723 ( new_n925_, new_n602_, new_n922_ );
nand g724 ( new_n926_, new_n925_, new_n924_ );
nand g725 ( new_n927_, new_n926_, new_n923_ );
nand g726 ( new_n928_, new_n927_, new_n305_ );
nand g727 ( new_n929_, new_n928_, N17 );
nand g728 ( new_n930_, new_n927_, new_n703_, new_n305_ );
nand g729 ( N728, new_n929_, new_n930_ );
nand g730 ( new_n932_, new_n927_, new_n561_ );
nand g731 ( new_n933_, new_n932_, N21 );
nand g732 ( new_n934_, new_n927_, new_n704_, new_n561_ );
nand g733 ( N729, new_n933_, new_n934_ );
nand g734 ( new_n936_, new_n927_, new_n526_ );
nand g735 ( new_n937_, new_n936_, N25 );
nand g736 ( new_n938_, new_n927_, new_n353_, new_n526_ );
nand g737 ( N730, new_n937_, new_n938_ );
nand g738 ( new_n940_, new_n927_, new_n460_ );
nand g739 ( new_n941_, new_n940_, N29 );
nand g740 ( new_n942_, new_n927_, new_n429_, new_n460_ );
nand g741 ( N731, new_n941_, new_n942_ );
not g742 ( new_n944_, keyIn_0_116 );
not g743 ( new_n945_, new_n897_ );
nor g744 ( new_n946_, new_n945_, new_n847_ );
nand g745 ( new_n947_, new_n602_, new_n798_, new_n946_ );
nand g746 ( new_n948_, new_n947_, new_n944_ );
nand g747 ( new_n949_, new_n902_, keyIn_0_116, new_n946_ );
nand g748 ( new_n950_, new_n948_, new_n949_ );
nand g749 ( new_n951_, new_n950_, new_n305_ );
nand g750 ( new_n952_, new_n951_, N33 );
nand g751 ( new_n953_, new_n950_, new_n628_, new_n305_ );
nand g752 ( N732, new_n952_, new_n953_ );
nand g753 ( new_n955_, new_n950_, new_n561_ );
nand g754 ( new_n956_, new_n955_, N37 );
nand g755 ( new_n957_, new_n950_, new_n629_, new_n561_ );
nand g756 ( N733, new_n956_, new_n957_ );
nand g757 ( new_n959_, new_n950_, new_n526_ );
nand g758 ( new_n960_, new_n959_, N41 );
nand g759 ( new_n961_, new_n950_, new_n636_, new_n526_ );
nand g760 ( N734, new_n960_, new_n961_ );
nand g761 ( new_n963_, new_n950_, new_n460_ );
nand g762 ( new_n964_, new_n963_, N45 );
nand g763 ( new_n965_, new_n950_, new_n440_, new_n460_ );
nand g764 ( N735, new_n964_, new_n965_ );
not g765 ( new_n967_, keyIn_0_117 );
nor g766 ( new_n968_, new_n921_, new_n847_, new_n945_ );
nand g767 ( new_n969_, new_n600_, new_n591_, new_n968_ );
nand g768 ( new_n970_, new_n969_, new_n967_ );
nand g769 ( new_n971_, new_n600_, new_n591_, keyIn_0_117, new_n968_ );
nand g770 ( new_n972_, new_n970_, new_n971_ );
nand g771 ( new_n973_, new_n972_, new_n305_ );
nand g772 ( new_n974_, new_n973_, N49 );
nand g773 ( new_n975_, new_n972_, new_n723_, new_n305_ );
nand g774 ( N736, new_n974_, new_n975_ );
nand g775 ( new_n977_, new_n972_, new_n561_ );
nand g776 ( new_n978_, new_n977_, N53 );
nand g777 ( new_n979_, new_n972_, new_n724_, new_n561_ );
nand g778 ( N737, new_n978_, new_n979_ );
nand g779 ( new_n981_, new_n972_, new_n526_ );
nand g780 ( new_n982_, new_n981_, N57 );
nand g781 ( new_n983_, new_n972_, new_n731_, new_n526_ );
nand g782 ( N738, new_n982_, new_n983_ );
not g783 ( new_n985_, keyIn_0_122 );
nand g784 ( new_n986_, new_n972_, new_n460_ );
nand g785 ( new_n987_, new_n986_, new_n985_ );
nand g786 ( new_n988_, new_n972_, keyIn_0_122, new_n460_ );
nand g787 ( new_n989_, new_n987_, new_n988_ );
nand g788 ( new_n990_, new_n989_, N61 );
nand g789 ( new_n991_, new_n987_, new_n438_, new_n988_ );
nand g790 ( N739, new_n990_, new_n991_ );
not g791 ( new_n993_, keyIn_0_123 );
not g792 ( new_n994_, keyIn_0_118 );
not g793 ( new_n995_, keyIn_0_113 );
not g794 ( new_n996_, keyIn_0_100 );
nand g795 ( new_n997_, new_n796_, new_n996_, new_n793_ );
not g796 ( new_n998_, keyIn_0_99 );
nand g797 ( new_n999_, new_n697_, new_n998_ );
nand g798 ( new_n1000_, new_n695_, keyIn_0_99, new_n696_ );
nand g799 ( new_n1001_, new_n999_, new_n997_, new_n1000_ );
nand g800 ( new_n1002_, new_n845_, keyIn_0_98, new_n846_ );
not g801 ( new_n1003_, keyIn_0_98 );
nand g802 ( new_n1004_, new_n847_, new_n1003_ );
nand g803 ( new_n1005_, new_n1004_, new_n1002_ );
not g804 ( new_n1006_, new_n1005_ );
nand g805 ( new_n1007_, new_n797_, keyIn_0_100 );
nand g806 ( new_n1008_, new_n1007_, new_n897_ );
nor g807 ( new_n1009_, new_n1006_, new_n1001_, new_n1008_ );
nor g808 ( new_n1010_, new_n1009_, keyIn_0_110 );
not g809 ( new_n1011_, keyIn_0_109 );
nand g810 ( new_n1012_, new_n797_, keyIn_0_97 );
not g811 ( new_n1013_, keyIn_0_97 );
nand g812 ( new_n1014_, new_n796_, new_n1013_, new_n793_ );
nand g813 ( new_n1015_, new_n1014_, new_n697_ );
not g814 ( new_n1016_, new_n1015_ );
nand g815 ( new_n1017_, new_n896_, keyIn_0_96, new_n893_ );
not g816 ( new_n1018_, keyIn_0_96 );
nand g817 ( new_n1019_, new_n897_, new_n1018_ );
nand g818 ( new_n1020_, new_n1019_, new_n1017_ );
nand g819 ( new_n1021_, new_n845_, keyIn_0_95, new_n846_ );
not g820 ( new_n1022_, keyIn_0_95 );
nand g821 ( new_n1023_, new_n847_, new_n1022_ );
nand g822 ( new_n1024_, new_n1023_, new_n1021_ );
nand g823 ( new_n1025_, new_n1016_, new_n1020_, new_n1024_, new_n1012_ );
nand g824 ( new_n1026_, new_n1025_, new_n1011_ );
not g825 ( new_n1027_, new_n1026_ );
nor g826 ( new_n1028_, new_n1010_, new_n1027_ );
not g827 ( new_n1029_, new_n1012_ );
nor g828 ( new_n1030_, new_n1029_, new_n1015_ );
nand g829 ( new_n1031_, new_n1030_, keyIn_0_109, new_n1020_, new_n1024_ );
not g830 ( new_n1032_, new_n1031_ );
not g831 ( new_n1033_, keyIn_0_110 );
not g832 ( new_n1034_, new_n1001_ );
not g833 ( new_n1035_, new_n1008_ );
nand g834 ( new_n1036_, new_n1034_, new_n1005_, new_n1035_ );
nor g835 ( new_n1037_, new_n1036_, new_n1033_ );
nor g836 ( new_n1038_, new_n1037_, new_n1032_ );
not g837 ( new_n1039_, keyIn_0_103 );
nand g838 ( new_n1040_, new_n796_, new_n1039_, new_n793_ );
nand g839 ( new_n1041_, new_n897_, keyIn_0_101 );
not g840 ( new_n1042_, keyIn_0_101 );
nand g841 ( new_n1043_, new_n896_, new_n1042_, new_n893_ );
nand g842 ( new_n1044_, new_n1041_, new_n1040_, new_n1043_ );
not g843 ( new_n1045_, new_n1044_ );
not g844 ( new_n1046_, keyIn_0_102 );
nand g845 ( new_n1047_, new_n698_, new_n1046_ );
nand g846 ( new_n1048_, new_n697_, keyIn_0_102 );
nand g847 ( new_n1049_, new_n1047_, new_n1048_ );
nand g848 ( new_n1050_, new_n797_, keyIn_0_103 );
nand g849 ( new_n1051_, new_n1050_, new_n847_ );
not g850 ( new_n1052_, new_n1051_ );
nand g851 ( new_n1053_, new_n1045_, new_n1049_, new_n1052_, keyIn_0_111 );
not g852 ( new_n1054_, keyIn_0_111 );
nand g853 ( new_n1055_, new_n1045_, new_n1049_, new_n1052_ );
nand g854 ( new_n1056_, new_n1055_, new_n1054_ );
nand g855 ( new_n1057_, new_n1056_, new_n1053_ );
not g856 ( new_n1058_, keyIn_0_92 );
nand g857 ( new_n1059_, new_n847_, new_n1058_ );
not g858 ( new_n1060_, new_n1059_ );
nand g859 ( new_n1061_, new_n845_, keyIn_0_92, new_n846_ );
nand g860 ( new_n1062_, new_n1061_, new_n797_ );
nor g861 ( new_n1063_, new_n1060_, new_n1062_ );
not g862 ( new_n1064_, keyIn_0_93 );
nand g863 ( new_n1065_, new_n945_, new_n1064_ );
nand g864 ( new_n1066_, new_n897_, keyIn_0_93 );
nand g865 ( new_n1067_, new_n1065_, new_n1066_ );
nand g866 ( new_n1068_, new_n698_, keyIn_0_94 );
not g867 ( new_n1069_, keyIn_0_94 );
nand g868 ( new_n1070_, new_n697_, new_n1069_ );
nand g869 ( new_n1071_, new_n1068_, new_n1070_ );
nand g870 ( new_n1072_, new_n1063_, new_n1067_, new_n1071_ );
nand g871 ( new_n1073_, new_n1072_, keyIn_0_108 );
not g872 ( new_n1074_, keyIn_0_108 );
nand g873 ( new_n1075_, new_n1063_, new_n1067_, new_n1071_, new_n1074_ );
nand g874 ( new_n1076_, new_n1073_, new_n1075_ );
nand g875 ( new_n1077_, new_n1028_, new_n1038_, new_n1057_, new_n1076_ );
nand g876 ( new_n1078_, new_n1077_, new_n995_ );
nand g877 ( new_n1079_, new_n1036_, new_n1033_ );
nand g878 ( new_n1080_, new_n1079_, new_n1026_ );
nand g879 ( new_n1081_, new_n1009_, keyIn_0_110 );
nand g880 ( new_n1082_, new_n1081_, new_n1031_ );
nor g881 ( new_n1083_, new_n1082_, new_n1080_ );
nand g882 ( new_n1084_, new_n1083_, keyIn_0_113, new_n1057_, new_n1076_ );
nand g883 ( new_n1085_, new_n305_, new_n517_ );
nand g884 ( new_n1086_, new_n526_, new_n459_ );
nor g885 ( new_n1087_, new_n1085_, new_n1086_ );
nand g886 ( new_n1088_, new_n1078_, new_n1084_, new_n994_, new_n1087_ );
nand g887 ( new_n1089_, new_n1078_, new_n1084_, new_n1087_ );
nand g888 ( new_n1090_, new_n1089_, keyIn_0_118 );
nand g889 ( new_n1091_, new_n1090_, new_n1088_ );
nand g890 ( new_n1092_, new_n1091_, new_n847_ );
nand g891 ( new_n1093_, new_n1092_, new_n993_ );
nand g892 ( new_n1094_, new_n1091_, keyIn_0_123, new_n847_ );
nand g893 ( new_n1095_, new_n1093_, new_n1094_ );
nand g894 ( new_n1096_, new_n1095_, new_n230_ );
nand g895 ( new_n1097_, new_n1093_, N65, new_n1094_ );
nand g896 ( N740, new_n1096_, new_n1097_ );
nand g897 ( new_n1099_, new_n1091_, new_n897_ );
nand g898 ( new_n1100_, new_n1099_, keyIn_0_124 );
not g899 ( new_n1101_, keyIn_0_124 );
nand g900 ( new_n1102_, new_n1091_, new_n1101_, new_n897_ );
nand g901 ( new_n1103_, new_n1100_, new_n1102_ );
nand g902 ( new_n1104_, new_n1103_, N69 );
nand g903 ( new_n1105_, new_n1100_, new_n231_, new_n1102_ );
nand g904 ( N741, new_n1104_, new_n1105_ );
not g905 ( new_n1107_, keyIn_0_125 );
nand g906 ( new_n1108_, new_n1091_, new_n697_ );
nand g907 ( new_n1109_, new_n1108_, new_n1107_ );
nand g908 ( new_n1110_, new_n1091_, keyIn_0_125, new_n697_ );
nand g909 ( new_n1111_, new_n1109_, new_n1110_ );
nand g910 ( new_n1112_, new_n1111_, N73 );
nand g911 ( new_n1113_, new_n1109_, new_n238_, new_n1110_ );
nand g912 ( N742, new_n1112_, new_n1113_ );
nand g913 ( new_n1115_, new_n1091_, new_n797_ );
nand g914 ( new_n1116_, new_n1115_, keyIn_0_126 );
not g915 ( new_n1117_, keyIn_0_126 );
nand g916 ( new_n1118_, new_n1091_, new_n1117_, new_n797_ );
nand g917 ( new_n1119_, new_n1116_, new_n1118_ );
nand g918 ( new_n1120_, new_n1119_, N77 );
nand g919 ( new_n1121_, new_n1116_, new_n239_, new_n1118_ );
nand g920 ( N743, new_n1120_, new_n1121_ );
not g921 ( new_n1123_, keyIn_0_127 );
not g922 ( new_n1124_, keyIn_0_119 );
nand g923 ( new_n1125_, new_n460_, new_n461_ );
nor g924 ( new_n1126_, new_n1085_, new_n1125_ );
nand g925 ( new_n1127_, new_n1078_, new_n1084_, new_n1124_, new_n1126_ );
nand g926 ( new_n1128_, new_n1078_, new_n1084_, new_n1126_ );
nand g927 ( new_n1129_, new_n1128_, keyIn_0_119 );
nand g928 ( new_n1130_, new_n1129_, new_n1127_ );
nand g929 ( new_n1131_, new_n1130_, new_n847_ );
nand g930 ( new_n1132_, new_n1131_, new_n1123_ );
nand g931 ( new_n1133_, new_n1130_, keyIn_0_127, new_n847_ );
nand g932 ( new_n1134_, new_n1132_, new_n1133_ );
nand g933 ( new_n1135_, new_n1134_, new_n205_ );
nand g934 ( new_n1136_, new_n1132_, N81, new_n1133_ );
nand g935 ( N744, new_n1135_, new_n1136_ );
nand g936 ( new_n1138_, new_n1130_, new_n897_ );
nand g937 ( new_n1139_, new_n1138_, N85 );
nand g938 ( new_n1140_, new_n1130_, new_n206_, new_n897_ );
nand g939 ( N745, new_n1139_, new_n1140_ );
nand g940 ( new_n1142_, new_n1130_, new_n697_ );
nand g941 ( new_n1143_, new_n1142_, N89 );
nand g942 ( new_n1144_, new_n1130_, new_n213_, new_n697_ );
nand g943 ( N746, new_n1143_, new_n1144_ );
nand g944 ( new_n1146_, new_n1130_, new_n797_ );
nand g945 ( new_n1147_, new_n1146_, N93 );
nand g946 ( new_n1148_, new_n1130_, new_n214_, new_n797_ );
nand g947 ( N747, new_n1147_, new_n1148_ );
nand g948 ( new_n1150_, new_n561_, new_n304_ );
nor g949 ( new_n1151_, new_n1086_, new_n1150_ );
nand g950 ( new_n1152_, new_n1078_, new_n1084_, keyIn_0_120, new_n1151_ );
not g951 ( new_n1153_, keyIn_0_120 );
nand g952 ( new_n1154_, new_n1078_, new_n1084_, new_n1151_ );
nand g953 ( new_n1155_, new_n1154_, new_n1153_ );
nand g954 ( new_n1156_, new_n1155_, new_n1152_ );
nand g955 ( new_n1157_, new_n1156_, new_n847_ );
nand g956 ( new_n1158_, new_n1157_, N97 );
nand g957 ( new_n1159_, new_n1156_, new_n310_, new_n847_ );
nand g958 ( N748, new_n1158_, new_n1159_ );
nand g959 ( new_n1161_, new_n1156_, new_n897_ );
nand g960 ( new_n1162_, new_n1161_, N101 );
nand g961 ( new_n1163_, new_n1156_, new_n311_, new_n897_ );
nand g962 ( N749, new_n1162_, new_n1163_ );
nand g963 ( new_n1165_, new_n1156_, new_n697_ );
nand g964 ( new_n1166_, new_n1165_, N105 );
nand g965 ( new_n1167_, new_n1156_, new_n318_, new_n697_ );
nand g966 ( N750, new_n1166_, new_n1167_ );
nand g967 ( new_n1169_, new_n1156_, new_n797_ );
nand g968 ( new_n1170_, new_n1169_, N109 );
nand g969 ( new_n1171_, new_n1156_, new_n319_, new_n797_ );
nand g970 ( N751, new_n1170_, new_n1171_ );
not g971 ( new_n1173_, keyIn_0_121 );
nor g972 ( new_n1174_, new_n1125_, new_n1150_ );
nand g973 ( new_n1175_, new_n1078_, new_n1084_, new_n1173_, new_n1174_ );
nand g974 ( new_n1176_, new_n1078_, new_n1084_, new_n1174_ );
nand g975 ( new_n1177_, new_n1176_, keyIn_0_121 );
nand g976 ( new_n1178_, new_n1177_, new_n1175_ );
nand g977 ( new_n1179_, new_n1178_, new_n847_ );
nand g978 ( new_n1180_, new_n1179_, N113 );
nand g979 ( new_n1181_, new_n1178_, new_n388_, new_n847_ );
nand g980 ( N752, new_n1180_, new_n1181_ );
nand g981 ( new_n1183_, new_n1178_, new_n897_ );
nand g982 ( new_n1184_, new_n1183_, N117 );
nand g983 ( new_n1185_, new_n1178_, new_n389_, new_n897_ );
nand g984 ( N753, new_n1184_, new_n1185_ );
nand g985 ( new_n1187_, new_n1178_, new_n697_ );
nand g986 ( new_n1188_, new_n1187_, N121 );
nand g987 ( new_n1189_, new_n1178_, new_n395_, new_n697_ );
nand g988 ( N754, new_n1188_, new_n1189_ );
nand g989 ( new_n1191_, new_n1178_, new_n797_ );
nand g990 ( new_n1192_, new_n1191_, N125 );
nand g991 ( new_n1193_, new_n1178_, new_n396_, new_n797_ );
nand g992 ( N755, new_n1192_, new_n1193_ );
endmodule