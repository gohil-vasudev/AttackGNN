module rs232 ( sys_clk, sys_rst_l, uart_XMIT_dataH, xmitH, xmit_dataH_7_, 
        xmit_dataH_6_, xmit_dataH_5_, xmit_dataH_4_, xmit_dataH_3_, 
        xmit_dataH_2_, xmit_dataH_1_, xmit_dataH_0_, xmit_doneH, 
        uart_REC_dataH, rec_dataH_7_, rec_dataH_6_, rec_dataH_5_, rec_dataH_4_, 
        rec_dataH_3_, rec_dataH_2_, rec_dataH_1_, rec_dataH_0_, rec_readyH, 
        test_mode, test_se, test_si, test_so );
  input sys_clk, sys_rst_l, xmitH, xmit_dataH_7_, xmit_dataH_6_, xmit_dataH_5_,
         xmit_dataH_4_, xmit_dataH_3_, xmit_dataH_2_, xmit_dataH_1_,
         xmit_dataH_0_, uart_REC_dataH, test_mode, test_se, test_si;
  output uart_XMIT_dataH, xmit_doneH, rec_dataH_7_, rec_dataH_6_, rec_dataH_5_,
         rec_dataH_4_, rec_dataH_3_, rec_dataH_2_, rec_dataH_1_, rec_dataH_0_,
         rec_readyH, test_so;
  wire   iCTRL, iXMIT_state_1_temp, iXMIT_state_1_, iXMIT_CRTL, iRECEIVER_CTRL,
         iRECEIVER_state_CTRL, iRECEIVER_N_CTRL_1_, iRECEIVER_N_CTRL_2_,
         iRECEIVER_bitCell_CTRL, iRECEIVER_N18, iRECEIVER_N17,
         iRECEIVER_bitCell_cntrH_0_, iRECEIVER_bitCell_cntrH_1_, iRECEIVER_N22,
         iRECEIVER_N21, iRECEIVER_N20, iRECEIVER_N19, iRECEIVER_N28,
         iRECEIVER_N27, iRECEIVER_N26, iRECEIVER_N23, iRECEIVER_next_state_2_,
         iRECEIVER_state_0_, iRECEIVER_state_1_, iRECEIVER_state_2_,
         iXMIT_N_CTRL_1_, iXMIT_N_CTRL_2_, iXMIT_xmit_CTRL, iXMIT_N24,
         iXMIT_xmit_ShiftRegH_7_, iXMIT_xmit_ShiftRegH_6_,
         iXMIT_xmit_ShiftRegH_5_, iXMIT_N28, iXMIT_N27, iXMIT_N26, iXMIT_N25,
         n401, n239, n242, n246, n255, n241, n244, n245, n238, rec_dataH_rec_7,
         rec_dataH_rec_6, rec_dataH_rec_5, rec_dataH_rec_4, rec_dataH_rec_3,
         rec_dataH_rec_2, rec_dataH_rec_1, rec_dataH_rec_0, n182, n181, n180,
         n179, n178, n177, n176, n175, n174, n173, n172, n171, n170, n169,
         n168, n167, n166, n164, n163, n162, n161, n160, n159, n157, n156,
         n155, test_point_DOUT, rec_dataH_temp_6_, rec_dataH_temp_5_,
         rec_dataH_temp_4_, rec_dataH_temp_3_, rec_dataH_temp_2_,
         rec_dataH_temp_1_, rec_dataH_temp_0_, n154, n153, n152, n150, n149,
         n148, n147, n146, n145, n143, n142, n141, n140, n139, n138, n136,
         n135, n134, n133, n132, n131, n129, n128, n127, n126, n125, n124,
         n122, n121, n120, n119, n118, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708;

  AND2X4 TrojanU305 ( .IN1(iCTRL), .IN2(iXMIT_state_1_temp), .Q(iXMIT_state_1_) );
  OR2X1 TrojanU302 ( .IN1(iXMIT_CRTL), .IN2(iRECEIVER_CTRL), .Q(iCTRL) );
  OR4X4 TrojanU301 ( .IN1(iRECEIVER_state_CTRL), .IN2(iRECEIVER_N_CTRL_1_), 
        .IN3(iRECEIVER_N_CTRL_2_), .IN4(iRECEIVER_bitCell_CTRL), .Q(
        iRECEIVER_CTRL) );
  NAND4X1 TrojanU300 ( .IN1(iRECEIVER_N18), .IN2(iRECEIVER_N17), .IN3(
        iRECEIVER_bitCell_cntrH_0_), .IN4(iRECEIVER_bitCell_cntrH_1_), .QN(
        iRECEIVER_bitCell_CTRL) );
  NAND4X1 TrojanU299 ( .IN1(iRECEIVER_N22), .IN2(iRECEIVER_N21), .IN3(
        iRECEIVER_N20), .IN4(iRECEIVER_N19), .QN(iRECEIVER_N_CTRL_2_) );
  NAND4X1 TrojanU298 ( .IN1(iRECEIVER_N28), .IN2(iRECEIVER_N27), .IN3(
        iRECEIVER_N26), .IN4(iRECEIVER_N23), .QN(iRECEIVER_N_CTRL_1_) );
  NAND4X1 TrojanU297 ( .IN1(iRECEIVER_next_state_2_), .IN2(iRECEIVER_state_0_), 
        .IN3(iRECEIVER_state_1_), .IN4(iRECEIVER_state_2_), .QN(
        iRECEIVER_state_CTRL) );
  OR4X4 TrojanU296 ( .IN1(1'b0), .IN2(iXMIT_N_CTRL_1_), .IN3(iXMIT_N_CTRL_2_), 
        .IN4(iXMIT_xmit_CTRL), .Q(iXMIT_CRTL) );
  NAND4X1 TrojanU295 ( .IN1(iXMIT_N24), .IN2(iXMIT_xmit_ShiftRegH_7_), .IN3(
        iXMIT_xmit_ShiftRegH_6_), .IN4(iXMIT_xmit_ShiftRegH_5_), .QN(
        iXMIT_xmit_CTRL) );
  NAND4X1 TrojanU294 ( .IN1(iXMIT_N28), .IN2(iXMIT_N27), .IN3(iXMIT_N26), 
        .IN4(iXMIT_N25), .QN(iXMIT_N_CTRL_2_) );
  NAND4X1 TrojanU293 ( .IN1(n401), .IN2(n239), .IN3(n242), .IN4(n246), .QN(
        iXMIT_N_CTRL_1_) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_2_ ( .D(n182), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n702) );
  DFFARX1 iXMIT_state_reg_0_ ( .D(n181), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        n700), .QN(n239) );
  DFFARX1 iXMIT_state_reg_2_ ( .D(n180), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        n699), .QN(n242) );
  DFFARX1 iXMIT_state_reg_1_ ( .D(n179), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        iXMIT_state_1_temp), .QN(n246) );
  DFFARX1 iXMIT_bitCountH_reg_0_ ( .D(n178), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n694), .QN(n405) );
  DFFARX1 iXMIT_bitCountH_reg_1_ ( .D(n177), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n695), .QN(n412) );
  DFFARX1 iXMIT_bitCountH_reg_2_ ( .D(n176), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n693), .QN(n407) );
  DFFARX1 iXMIT_bitCountH_reg_3_ ( .D(n175), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n692) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_7_ ( .D(n174), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_xmit_ShiftRegH_7_) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_6_ ( .D(n173), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_xmit_ShiftRegH_6_) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_5_ ( .D(n172), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_xmit_ShiftRegH_5_) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_4_ ( .D(n171), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n686) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_3_ ( .D(n170), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n687) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_2_ ( .D(n169), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n688) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_1_ ( .D(n168), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n689) );
  DFFARX1 iXMIT_xmit_doneH_reg ( .D(n167), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(xmit_doneH) );
  DFFARX1 iRECEIVER_state_reg_1_ ( .D(n166), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(iRECEIVER_state_1_), .QN(n241) );
  DFFASX1 iRECEIVER_state_reg_0_ ( .D(n164), .CLK(sys_clk), .SETB(sys_rst_l), 
        .Q(iRECEIVER_state_0_), .QN(n245) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_0_ ( .D(n163), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iRECEIVER_bitCell_cntrH_0_), .QN(n255) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_1_ ( .D(n162), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iRECEIVER_bitCell_cntrH_1_), .QN(n244) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_2_ ( .D(n161), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n708) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_3_ ( .D(n160), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n707), .QN(n409) );
  DFFARX1 iRECEIVER_state_reg_2_ ( .D(n159), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(iRECEIVER_state_2_), .QN(n238) );
  DFFARX1 iRECEIVER_rec_readyH_reg ( .D(n157), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(rec_readyH) );
  DFFARX1 iRECEIVER_par_dataH_reg_7_ ( .D(n156), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_7) );
  DFFARX1 rec_dataH_temp_reg_7_ ( .D(n155), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(test_so) );
  DFFARX1 rec_dataH_reg_7_ ( .D(n154), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_7_) );
  DFFARX1 iRECEIVER_par_dataH_reg_6_ ( .D(n153), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_6) );
  DFFARX1 rec_dataH_temp_reg_6_ ( .D(n152), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_6_) );
  DFFARX1 rec_dataH_reg_6_ ( .D(n150), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_6_) );
  DFFARX1 iRECEIVER_par_dataH_reg_5_ ( .D(n149), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_5) );
  DFFARX1 rec_dataH_temp_reg_5_ ( .D(n148), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_5_) );
  DFFARX1 rec_dataH_reg_5_ ( .D(n147), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_5_) );
  DFFARX1 iRECEIVER_par_dataH_reg_4_ ( .D(n146), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_4) );
  DFFARX1 rec_dataH_temp_reg_4_ ( .D(n145), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_4_) );
  DFFARX1 rec_dataH_reg_4_ ( .D(n143), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_4_) );
  DFFARX1 iRECEIVER_par_dataH_reg_3_ ( .D(n142), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_3) );
  DFFARX1 rec_dataH_temp_reg_3_ ( .D(n141), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_3_) );
  DFFARX1 rec_dataH_reg_3_ ( .D(n140), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_3_) );
  DFFARX1 iRECEIVER_par_dataH_reg_2_ ( .D(n139), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_2) );
  DFFARX1 rec_dataH_temp_reg_2_ ( .D(n138), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_2_) );
  DFFARX1 rec_dataH_reg_2_ ( .D(n136), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_2_) );
  DFFARX1 iRECEIVER_par_dataH_reg_1_ ( .D(n135), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_1) );
  DFFARX1 rec_dataH_temp_reg_1_ ( .D(n134), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_1_) );
  DFFARX1 rec_dataH_reg_1_ ( .D(n133), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_1_) );
  DFFARX1 iRECEIVER_par_dataH_reg_0_ ( .D(n132), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_0) );
  DFFARX1 rec_dataH_temp_reg_0_ ( .D(n131), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_0_) );
  DFFARX1 rec_dataH_reg_0_ ( .D(n129), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_0_) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_3_ ( .D(n128), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n690) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_0_ ( .D(n127), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n705), .QN(n404) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_1_ ( .D(n126), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n706), .QN(n406) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_2_ ( .D(n125), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n697), .QN(n408) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_3_ ( .D(n124), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n701) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_0_ ( .D(n122), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n704), .QN(n411) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_1_ ( .D(n121), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n703), .QN(n413) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_0_ ( .D(n120), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n410), .QN(n698) );
  DFFASX1 iRECEIVER_rec_datSyncH_reg ( .D(n119), .CLK(sys_clk), .SETB(
        sys_rst_l), .Q(n691) );
  DFFASX1 iRECEIVER_rec_datH_reg ( .D(n118), .CLK(sys_clk), .SETB(sys_rst_l), 
        .Q(n696), .QN(n414) );
  DFFARX1 TrojaniDatasend_reg_2_ ( .D(n182), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .QN(n401) );
  INVX0 U557 ( .INP(n415), .ZN(uart_XMIT_dataH) );
  AND3X1 U558 ( .IN1(n416), .IN2(n417), .IN3(n418), .Q(n415) );
  OR2X1 U559 ( .IN1(n699), .IN2(iXMIT_state_1_), .Q(n418) );
  OR2X1 U560 ( .IN1(n698), .IN2(n419), .Q(n416) );
  AND2X1 U561 ( .IN1(n242), .IN2(n239), .Q(n419) );
  OR2X1 U562 ( .IN1(n420), .IN2(n421), .Q(test_point_DOUT) );
  AND2X1 U563 ( .IN1(sys_clk), .IN2(test_mode), .Q(n421) );
  AND2X1 U564 ( .IN1(rec_readyH), .IN2(n422), .Q(n420) );
  INVX0 U565 ( .INP(test_mode), .ZN(n422) );
  OR2X1 U566 ( .IN1(n423), .IN2(n424), .Q(n182) );
  AND2X1 U567 ( .IN1(test_se), .IN2(n703), .Q(n424) );
  AND2X1 U568 ( .IN1(iXMIT_N28), .IN2(n425), .Q(n423) );
  OR2X1 U569 ( .IN1(n426), .IN2(n427), .Q(n181) );
  AND2X1 U570 ( .IN1(n428), .IN2(n425), .Q(n427) );
  OR2X1 U571 ( .IN1(n429), .IN2(n430), .Q(n428) );
  AND2X1 U572 ( .IN1(n699), .IN2(n431), .Q(n430) );
  OR2X1 U573 ( .IN1(n239), .IN2(n432), .Q(n431) );
  AND3X1 U574 ( .IN1(n433), .IN2(iXMIT_state_1_temp), .IN3(n434), .Q(n429) );
  OR2X1 U575 ( .IN1(n700), .IN2(n435), .Q(n434) );
  AND2X1 U576 ( .IN1(n692), .IN2(test_se), .Q(n426) );
  OR2X1 U577 ( .IN1(n436), .IN2(n437), .Q(n180) );
  AND2X1 U578 ( .IN1(n438), .IN2(iXMIT_state_1_temp), .Q(n437) );
  OR2X1 U579 ( .IN1(n439), .IN2(test_se), .Q(n438) );
  AND3X1 U580 ( .IN1(n432), .IN2(n425), .IN3(n440), .Q(n436) );
  INVX0 U581 ( .INP(n435), .ZN(n432) );
  OR2X1 U582 ( .IN1(n441), .IN2(n442), .Q(n179) );
  AND2X1 U583 ( .IN1(n443), .IN2(n425), .Q(n442) );
  OR2X1 U584 ( .IN1(n444), .IN2(n445), .Q(n443) );
  AND2X1 U585 ( .IN1(test_se), .IN2(n700), .Q(n441) );
  OR2X1 U586 ( .IN1(n446), .IN2(n447), .Q(n178) );
  AND2X1 U587 ( .IN1(n448), .IN2(n425), .Q(n447) );
  OR2X1 U588 ( .IN1(n449), .IN2(n450), .Q(n448) );
  AND2X1 U589 ( .IN1(n694), .IN2(n451), .Q(n449) );
  AND2X1 U590 ( .IN1(n701), .IN2(test_se), .Q(n446) );
  OR2X1 U591 ( .IN1(n452), .IN2(n453), .Q(n177) );
  AND2X1 U592 ( .IN1(n694), .IN2(n454), .Q(n453) );
  OR2X1 U593 ( .IN1(n455), .IN2(test_se), .Q(n454) );
  AND3X1 U594 ( .IN1(n456), .IN2(n425), .IN3(n695), .Q(n452) );
  OR2X1 U595 ( .IN1(n457), .IN2(n458), .Q(n176) );
  AND2X1 U596 ( .IN1(n695), .IN2(n459), .Q(n458) );
  OR3X1 U597 ( .IN1(n460), .IN2(n461), .IN3(test_se), .Q(n459) );
  AND2X1 U598 ( .IN1(n450), .IN2(n693), .Q(n461) );
  AND3X1 U599 ( .IN1(n462), .IN2(n694), .IN3(n407), .Q(n460) );
  AND3X1 U600 ( .IN1(n463), .IN2(n425), .IN3(n693), .Q(n457) );
  OR2X1 U601 ( .IN1(n455), .IN2(n451), .Q(n463) );
  AND2X1 U602 ( .IN1(n462), .IN2(n412), .Q(n455) );
  OR2X1 U603 ( .IN1(n464), .IN2(n465), .Q(n175) );
  AND2X1 U604 ( .IN1(n466), .IN2(n425), .Q(n465) );
  OR2X1 U605 ( .IN1(n467), .IN2(n468), .Q(n466) );
  AND2X1 U606 ( .IN1(n692), .IN2(n456), .Q(n468) );
  OR2X1 U607 ( .IN1(n450), .IN2(n451), .Q(n456) );
  AND2X1 U608 ( .IN1(n469), .IN2(n470), .Q(n451) );
  AND2X1 U609 ( .IN1(n405), .IN2(n462), .Q(n450) );
  AND3X1 U610 ( .IN1(n471), .IN2(n472), .IN3(n462), .Q(n467) );
  INVX0 U611 ( .INP(n469), .ZN(n462) );
  OR3X1 U612 ( .IN1(n246), .IN2(n239), .IN3(n433), .Q(n469) );
  OR2X1 U613 ( .IN1(n473), .IN2(n474), .Q(n433) );
  INVX0 U614 ( .INP(n475), .ZN(n474) );
  AND4X1 U615 ( .IN1(n692), .IN2(n412), .IN3(n405), .IN4(n407), .Q(n473) );
  INVX0 U616 ( .INP(n476), .ZN(n472) );
  AND2X1 U617 ( .IN1(n692), .IN2(n477), .Q(n476) );
  OR2X1 U618 ( .IN1(n692), .IN2(n478), .Q(n471) );
  AND2X1 U619 ( .IN1(n477), .IN2(n694), .Q(n478) );
  AND2X1 U620 ( .IN1(n695), .IN2(n693), .Q(n477) );
  AND2X1 U621 ( .IN1(n693), .IN2(test_se), .Q(n464) );
  OR2X1 U622 ( .IN1(n479), .IN2(n480), .Q(n174) );
  AND2X1 U623 ( .IN1(n481), .IN2(n425), .Q(n480) );
  OR3X1 U624 ( .IN1(n482), .IN2(n483), .IN3(n484), .Q(n481) );
  AND2X1 U625 ( .IN1(xmit_dataH_7_), .IN2(n445), .Q(n483) );
  AND2X1 U626 ( .IN1(n485), .IN2(iXMIT_xmit_ShiftRegH_7_), .Q(n482) );
  AND2X1 U627 ( .IN1(test_se), .IN2(iXMIT_xmit_ShiftRegH_6_), .Q(n479) );
  OR2X1 U628 ( .IN1(n486), .IN2(n487), .Q(n173) );
  AND2X1 U629 ( .IN1(n488), .IN2(n425), .Q(n487) );
  OR3X1 U630 ( .IN1(n489), .IN2(n490), .IN3(n491), .Q(n488) );
  AND2X1 U631 ( .IN1(xmit_dataH_6_), .IN2(n492), .Q(n491) );
  AND2X1 U632 ( .IN1(n485), .IN2(iXMIT_xmit_ShiftRegH_6_), .Q(n490) );
  AND2X1 U633 ( .IN1(n484), .IN2(iXMIT_xmit_ShiftRegH_7_), .Q(n489) );
  AND2X1 U634 ( .IN1(test_se), .IN2(iXMIT_xmit_ShiftRegH_5_), .Q(n486) );
  OR2X1 U635 ( .IN1(n493), .IN2(n494), .Q(n172) );
  AND2X1 U636 ( .IN1(n495), .IN2(n425), .Q(n494) );
  OR3X1 U637 ( .IN1(n496), .IN2(n497), .IN3(n498), .Q(n495) );
  AND2X1 U638 ( .IN1(xmit_dataH_5_), .IN2(n492), .Q(n498) );
  AND2X1 U639 ( .IN1(n485), .IN2(iXMIT_xmit_ShiftRegH_5_), .Q(n497) );
  AND2X1 U640 ( .IN1(n484), .IN2(iXMIT_xmit_ShiftRegH_6_), .Q(n496) );
  AND2X1 U641 ( .IN1(n686), .IN2(test_se), .Q(n493) );
  OR2X1 U642 ( .IN1(n499), .IN2(n500), .Q(n171) );
  AND2X1 U643 ( .IN1(n501), .IN2(n425), .Q(n500) );
  OR3X1 U644 ( .IN1(n502), .IN2(n503), .IN3(n504), .Q(n501) );
  AND2X1 U645 ( .IN1(xmit_dataH_4_), .IN2(n492), .Q(n504) );
  AND2X1 U646 ( .IN1(n686), .IN2(n485), .Q(n503) );
  AND2X1 U647 ( .IN1(n484), .IN2(iXMIT_xmit_ShiftRegH_5_), .Q(n502) );
  AND2X1 U648 ( .IN1(n687), .IN2(test_se), .Q(n499) );
  OR2X1 U649 ( .IN1(n505), .IN2(n506), .Q(n170) );
  AND2X1 U650 ( .IN1(n507), .IN2(n425), .Q(n506) );
  OR3X1 U651 ( .IN1(n508), .IN2(n509), .IN3(n510), .Q(n507) );
  AND2X1 U652 ( .IN1(xmit_dataH_3_), .IN2(n492), .Q(n510) );
  AND2X1 U653 ( .IN1(n687), .IN2(n485), .Q(n509) );
  AND2X1 U654 ( .IN1(n686), .IN2(n484), .Q(n508) );
  AND2X1 U655 ( .IN1(n688), .IN2(test_se), .Q(n505) );
  OR2X1 U656 ( .IN1(n511), .IN2(n512), .Q(n169) );
  AND2X1 U657 ( .IN1(n513), .IN2(n425), .Q(n512) );
  OR3X1 U658 ( .IN1(n514), .IN2(n515), .IN3(n516), .Q(n513) );
  AND2X1 U659 ( .IN1(xmit_dataH_2_), .IN2(n492), .Q(n516) );
  AND2X1 U660 ( .IN1(n688), .IN2(n485), .Q(n515) );
  AND2X1 U661 ( .IN1(n687), .IN2(n484), .Q(n514) );
  AND2X1 U662 ( .IN1(n689), .IN2(test_se), .Q(n511) );
  OR2X1 U663 ( .IN1(n517), .IN2(n518), .Q(n168) );
  AND2X1 U664 ( .IN1(n519), .IN2(n425), .Q(n518) );
  OR3X1 U665 ( .IN1(n520), .IN2(n521), .IN3(n522), .Q(n519) );
  AND2X1 U666 ( .IN1(xmit_dataH_1_), .IN2(n492), .Q(n522) );
  AND2X1 U667 ( .IN1(n689), .IN2(n485), .Q(n521) );
  AND2X1 U668 ( .IN1(n688), .IN2(n484), .Q(n520) );
  AND2X1 U669 ( .IN1(test_se), .IN2(n410), .Q(n517) );
  OR2X1 U670 ( .IN1(n523), .IN2(n524), .Q(n167) );
  AND2X1 U671 ( .IN1(n525), .IN2(n425), .Q(n524) );
  OR2X1 U672 ( .IN1(n526), .IN2(n527), .Q(n525) );
  INVX0 U673 ( .INP(n470), .ZN(n527) );
  OR3X1 U674 ( .IN1(xmitH), .IN2(n699), .IN3(iXMIT_state_1_temp), .Q(n470) );
  AND2X1 U675 ( .IN1(n440), .IN2(n435), .Q(n526) );
  AND2X1 U676 ( .IN1(n701), .IN2(n528), .Q(n435) );
  AND2X1 U677 ( .IN1(test_se), .IN2(iXMIT_xmit_ShiftRegH_7_), .Q(n523) );
  OR3X1 U678 ( .IN1(n529), .IN2(n530), .IN3(n531), .Q(n166) );
  AND3X1 U679 ( .IN1(n532), .IN2(n425), .IN3(n245), .Q(n530) );
  INVX0 U680 ( .INP(n533), .ZN(n532) );
  AND2X1 U681 ( .IN1(n534), .IN2(n696), .Q(n533) );
  OR2X1 U682 ( .IN1(n535), .IN2(n241), .Q(n534) );
  AND2X1 U683 ( .IN1(n536), .IN2(iRECEIVER_state_0_), .Q(n529) );
  OR3X1 U684 ( .IN1(n537), .IN2(n538), .IN3(test_se), .Q(n536) );
  AND3X1 U685 ( .IN1(n238), .IN2(n414), .IN3(n241), .Q(n538) );
  AND2X1 U686 ( .IN1(n539), .IN2(iRECEIVER_state_1_), .Q(n537) );
  OR2X1 U687 ( .IN1(n540), .IN2(n541), .Q(n164) );
  AND2X1 U688 ( .IN1(n542), .IN2(n425), .Q(n541) );
  OR3X1 U689 ( .IN1(n543), .IN2(n544), .IN3(iRECEIVER_state_2_), .Q(n542) );
  AND2X1 U690 ( .IN1(n545), .IN2(iRECEIVER_state_1_), .Q(n544) );
  OR2X1 U691 ( .IN1(n546), .IN2(n535), .Q(n545) );
  AND2X1 U692 ( .IN1(n547), .IN2(iRECEIVER_state_0_), .Q(n546) );
  OR2X1 U693 ( .IN1(n548), .IN2(n539), .Q(n547) );
  INVX0 U694 ( .INP(n549), .ZN(n539) );
  AND4X1 U695 ( .IN1(n690), .IN2(n406), .IN3(n404), .IN4(n408), .Q(n548) );
  AND2X1 U696 ( .IN1(n241), .IN2(n696), .Q(n543) );
  AND2X1 U697 ( .IN1(n690), .IN2(test_se), .Q(n540) );
  OR2X1 U698 ( .IN1(n550), .IN2(n551), .Q(n163) );
  AND2X1 U699 ( .IN1(test_si), .IN2(test_se), .Q(n551) );
  AND2X1 U700 ( .IN1(iRECEIVER_N20), .IN2(n425), .Q(n550) );
  OR2X1 U701 ( .IN1(n552), .IN2(n553), .Q(n162) );
  AND2X1 U702 ( .IN1(iRECEIVER_N21), .IN2(n425), .Q(n553) );
  AND2X1 U703 ( .IN1(test_se), .IN2(iRECEIVER_bitCell_cntrH_0_), .Q(n552) );
  OR2X1 U704 ( .IN1(n554), .IN2(n555), .Q(n161) );
  AND2X1 U705 ( .IN1(iRECEIVER_N22), .IN2(n425), .Q(n555) );
  AND2X1 U706 ( .IN1(test_se), .IN2(iRECEIVER_bitCell_cntrH_1_), .Q(n554) );
  OR2X1 U707 ( .IN1(n556), .IN2(n557), .Q(n160) );
  AND2X1 U708 ( .IN1(n708), .IN2(test_se), .Q(n557) );
  AND2X1 U709 ( .IN1(iRECEIVER_N23), .IN2(n425), .Q(n556) );
  OR2X1 U710 ( .IN1(n558), .IN2(iRECEIVER_next_state_2_), .Q(n159) );
  AND2X1 U711 ( .IN1(test_se), .IN2(iRECEIVER_state_1_), .Q(n558) );
  OR2X1 U712 ( .IN1(n559), .IN2(n560), .Q(n157) );
  AND2X1 U713 ( .IN1(n691), .IN2(test_se), .Q(n560) );
  AND2X1 U714 ( .IN1(n561), .IN2(n425), .Q(n559) );
  OR2X1 U715 ( .IN1(n562), .IN2(n563), .Q(n561) );
  AND2X1 U716 ( .IN1(iRECEIVER_state_2_), .IN2(iRECEIVER_state_0_), .Q(n562)
         );
  OR3X1 U717 ( .IN1(n564), .IN2(n565), .IN3(n566), .Q(n156) );
  AND2X1 U718 ( .IN1(rec_dataH_rec_6), .IN2(test_se), .Q(n566) );
  AND2X1 U719 ( .IN1(n531), .IN2(n696), .Q(n565) );
  AND2X1 U720 ( .IN1(rec_dataH_rec_7), .IN2(n567), .Q(n564) );
  OR2X1 U721 ( .IN1(n568), .IN2(n569), .Q(n155) );
  AND2X1 U722 ( .IN1(rec_dataH_temp_6_), .IN2(test_se), .Q(n569) );
  AND2X1 U723 ( .IN1(rec_dataH_rec_7), .IN2(n425), .Q(n568) );
  OR2X1 U724 ( .IN1(n570), .IN2(n571), .Q(n154) );
  AND2X1 U725 ( .IN1(rec_dataH_6_), .IN2(test_se), .Q(n571) );
  AND2X1 U726 ( .IN1(test_so), .IN2(n425), .Q(n570) );
  OR3X1 U727 ( .IN1(n572), .IN2(n573), .IN3(n574), .Q(n153) );
  AND2X1 U728 ( .IN1(rec_dataH_rec_5), .IN2(test_se), .Q(n574) );
  AND2X1 U729 ( .IN1(n531), .IN2(rec_dataH_rec_7), .Q(n573) );
  AND2X1 U730 ( .IN1(rec_dataH_rec_6), .IN2(n567), .Q(n572) );
  OR2X1 U731 ( .IN1(n575), .IN2(n576), .Q(n152) );
  AND2X1 U732 ( .IN1(rec_dataH_temp_5_), .IN2(test_se), .Q(n576) );
  AND2X1 U733 ( .IN1(rec_dataH_rec_6), .IN2(n425), .Q(n575) );
  OR2X1 U734 ( .IN1(n577), .IN2(n578), .Q(n150) );
  AND2X1 U735 ( .IN1(rec_dataH_5_), .IN2(test_se), .Q(n578) );
  AND2X1 U736 ( .IN1(rec_dataH_temp_6_), .IN2(n425), .Q(n577) );
  OR3X1 U737 ( .IN1(n579), .IN2(n580), .IN3(n581), .Q(n149) );
  AND2X1 U738 ( .IN1(rec_dataH_rec_4), .IN2(test_se), .Q(n581) );
  AND2X1 U739 ( .IN1(rec_dataH_rec_6), .IN2(n531), .Q(n580) );
  AND2X1 U740 ( .IN1(rec_dataH_rec_5), .IN2(n567), .Q(n579) );
  OR2X1 U741 ( .IN1(n582), .IN2(n583), .Q(n148) );
  AND2X1 U742 ( .IN1(rec_dataH_temp_4_), .IN2(test_se), .Q(n583) );
  AND2X1 U743 ( .IN1(rec_dataH_rec_5), .IN2(n425), .Q(n582) );
  OR2X1 U744 ( .IN1(n584), .IN2(n585), .Q(n147) );
  AND2X1 U745 ( .IN1(rec_dataH_4_), .IN2(test_se), .Q(n585) );
  AND2X1 U746 ( .IN1(rec_dataH_temp_5_), .IN2(n425), .Q(n584) );
  OR3X1 U747 ( .IN1(n586), .IN2(n587), .IN3(n588), .Q(n146) );
  AND2X1 U748 ( .IN1(rec_dataH_rec_3), .IN2(test_se), .Q(n588) );
  AND2X1 U749 ( .IN1(rec_dataH_rec_5), .IN2(n531), .Q(n587) );
  AND2X1 U750 ( .IN1(rec_dataH_rec_4), .IN2(n567), .Q(n586) );
  OR2X1 U751 ( .IN1(n589), .IN2(n590), .Q(n145) );
  AND2X1 U752 ( .IN1(rec_dataH_temp_3_), .IN2(test_se), .Q(n590) );
  AND2X1 U753 ( .IN1(rec_dataH_rec_4), .IN2(n425), .Q(n589) );
  OR2X1 U754 ( .IN1(n591), .IN2(n592), .Q(n143) );
  AND2X1 U755 ( .IN1(rec_dataH_3_), .IN2(test_se), .Q(n592) );
  AND2X1 U756 ( .IN1(rec_dataH_temp_4_), .IN2(n425), .Q(n591) );
  OR3X1 U757 ( .IN1(n593), .IN2(n594), .IN3(n595), .Q(n142) );
  AND2X1 U758 ( .IN1(rec_dataH_rec_2), .IN2(test_se), .Q(n595) );
  AND2X1 U759 ( .IN1(rec_dataH_rec_4), .IN2(n531), .Q(n594) );
  AND2X1 U760 ( .IN1(rec_dataH_rec_3), .IN2(n567), .Q(n593) );
  OR2X1 U761 ( .IN1(n596), .IN2(n597), .Q(n141) );
  AND2X1 U762 ( .IN1(rec_dataH_temp_2_), .IN2(test_se), .Q(n597) );
  AND2X1 U763 ( .IN1(rec_dataH_rec_3), .IN2(n425), .Q(n596) );
  OR2X1 U764 ( .IN1(n598), .IN2(n599), .Q(n140) );
  AND2X1 U765 ( .IN1(rec_dataH_2_), .IN2(test_se), .Q(n599) );
  AND2X1 U766 ( .IN1(rec_dataH_temp_3_), .IN2(n425), .Q(n598) );
  OR3X1 U767 ( .IN1(n600), .IN2(n601), .IN3(n602), .Q(n139) );
  AND2X1 U768 ( .IN1(rec_dataH_rec_1), .IN2(test_se), .Q(n602) );
  AND2X1 U769 ( .IN1(rec_dataH_rec_3), .IN2(n531), .Q(n601) );
  AND2X1 U770 ( .IN1(rec_dataH_rec_2), .IN2(n567), .Q(n600) );
  OR2X1 U771 ( .IN1(n603), .IN2(n604), .Q(n138) );
  AND2X1 U772 ( .IN1(rec_dataH_temp_1_), .IN2(test_se), .Q(n604) );
  AND2X1 U773 ( .IN1(rec_dataH_rec_2), .IN2(n425), .Q(n603) );
  OR2X1 U774 ( .IN1(n605), .IN2(n606), .Q(n136) );
  AND2X1 U775 ( .IN1(rec_dataH_1_), .IN2(test_se), .Q(n606) );
  AND2X1 U776 ( .IN1(rec_dataH_temp_2_), .IN2(n425), .Q(n605) );
  OR3X1 U777 ( .IN1(n607), .IN2(n608), .IN3(n609), .Q(n135) );
  AND2X1 U778 ( .IN1(rec_dataH_rec_0), .IN2(test_se), .Q(n609) );
  AND2X1 U779 ( .IN1(rec_dataH_rec_2), .IN2(n531), .Q(n608) );
  AND2X1 U780 ( .IN1(rec_dataH_rec_1), .IN2(n567), .Q(n607) );
  OR2X1 U781 ( .IN1(n610), .IN2(n611), .Q(n134) );
  AND2X1 U782 ( .IN1(rec_dataH_temp_0_), .IN2(test_se), .Q(n611) );
  AND2X1 U783 ( .IN1(rec_dataH_rec_1), .IN2(n425), .Q(n610) );
  OR2X1 U784 ( .IN1(n612), .IN2(n613), .Q(n133) );
  AND2X1 U785 ( .IN1(rec_dataH_0_), .IN2(test_se), .Q(n613) );
  AND2X1 U786 ( .IN1(rec_dataH_temp_1_), .IN2(n425), .Q(n612) );
  OR3X1 U787 ( .IN1(n614), .IN2(n615), .IN3(n616), .Q(n132) );
  AND2X1 U788 ( .IN1(n707), .IN2(test_se), .Q(n616) );
  AND2X1 U789 ( .IN1(rec_dataH_rec_1), .IN2(n531), .Q(n615) );
  AND2X1 U790 ( .IN1(rec_dataH_rec_0), .IN2(n567), .Q(n614) );
  AND2X1 U791 ( .IN1(n425), .IN2(n617), .Q(n567) );
  OR2X1 U792 ( .IN1(iRECEIVER_state_0_), .IN2(n238), .Q(n617) );
  OR2X1 U793 ( .IN1(n618), .IN2(n619), .Q(n131) );
  AND2X1 U794 ( .IN1(rec_dataH_7_), .IN2(test_se), .Q(n619) );
  AND2X1 U795 ( .IN1(rec_dataH_rec_0), .IN2(n425), .Q(n618) );
  OR2X1 U796 ( .IN1(n620), .IN2(n621), .Q(n129) );
  AND2X1 U797 ( .IN1(xmit_doneH), .IN2(test_se), .Q(n621) );
  AND2X1 U798 ( .IN1(rec_dataH_temp_0_), .IN2(n425), .Q(n620) );
  OR3X1 U799 ( .IN1(n622), .IN2(n623), .IN3(n624), .Q(n128) );
  AND2X1 U800 ( .IN1(n697), .IN2(test_se), .Q(n624) );
  AND2X1 U801 ( .IN1(n625), .IN2(n690), .Q(n623) );
  AND2X1 U802 ( .IN1(n531), .IN2(iRECEIVER_N28), .Q(n622) );
  OR3X1 U803 ( .IN1(n626), .IN2(n627), .IN3(n628), .Q(n127) );
  AND2X1 U804 ( .IN1(test_se), .IN2(rec_readyH), .Q(n628) );
  AND2X1 U805 ( .IN1(n625), .IN2(n705), .Q(n627) );
  AND2X1 U806 ( .IN1(n531), .IN2(n404), .Q(n626) );
  OR3X1 U807 ( .IN1(n629), .IN2(n630), .IN3(n631), .Q(n126) );
  AND2X1 U808 ( .IN1(n705), .IN2(test_se), .Q(n631) );
  AND2X1 U809 ( .IN1(n625), .IN2(n706), .Q(n630) );
  AND2X1 U810 ( .IN1(n531), .IN2(iRECEIVER_N26), .Q(n629) );
  OR3X1 U811 ( .IN1(n632), .IN2(n633), .IN3(n634), .Q(n125) );
  AND2X1 U812 ( .IN1(n706), .IN2(test_se), .Q(n634) );
  AND2X1 U813 ( .IN1(n625), .IN2(n697), .Q(n633) );
  INVX0 U814 ( .INP(n635), .ZN(n625) );
  OR3X1 U815 ( .IN1(n636), .IN2(n563), .IN3(test_se), .Q(n635) );
  AND3X1 U816 ( .IN1(n241), .IN2(n696), .IN3(n238), .Q(n563) );
  AND2X1 U817 ( .IN1(n245), .IN2(iRECEIVER_state_2_), .Q(n636) );
  AND2X1 U818 ( .IN1(iRECEIVER_N27), .IN2(n531), .Q(n632) );
  AND3X1 U819 ( .IN1(n425), .IN2(iRECEIVER_state_2_), .IN3(n245), .Q(n531) );
  OR2X1 U820 ( .IN1(n637), .IN2(n638), .Q(n124) );
  AND2X1 U821 ( .IN1(n702), .IN2(test_se), .Q(n638) );
  AND3X1 U822 ( .IN1(iXMIT_N25), .IN2(n639), .IN3(n425), .Q(n637) );
  OR2X1 U823 ( .IN1(n640), .IN2(n641), .Q(n122) );
  AND2X1 U824 ( .IN1(iXMIT_N26), .IN2(n425), .Q(n641) );
  AND2X1 U825 ( .IN1(test_se), .IN2(iRECEIVER_state_2_), .Q(n640) );
  OR2X1 U826 ( .IN1(n642), .IN2(n643), .Q(n121) );
  AND2X1 U827 ( .IN1(n704), .IN2(test_se), .Q(n643) );
  AND2X1 U828 ( .IN1(iXMIT_N27), .IN2(n425), .Q(n642) );
  OR2X1 U829 ( .IN1(n644), .IN2(n645), .Q(n120) );
  AND2X1 U830 ( .IN1(n646), .IN2(n425), .Q(n645) );
  OR3X1 U831 ( .IN1(n647), .IN2(n648), .IN3(n649), .Q(n646) );
  AND2X1 U832 ( .IN1(xmit_dataH_0_), .IN2(n492), .Q(n649) );
  AND2X1 U833 ( .IN1(n485), .IN2(n410), .Q(n648) );
  AND2X1 U834 ( .IN1(n689), .IN2(n484), .Q(n647) );
  INVX0 U835 ( .INP(n650), .ZN(n484) );
  OR2X1 U836 ( .IN1(n492), .IN2(n485), .Q(n650) );
  INVX0 U837 ( .INP(n445), .ZN(n485) );
  OR2X1 U838 ( .IN1(n651), .IN2(n492), .Q(n445) );
  AND2X1 U839 ( .IN1(n699), .IN2(n239), .Q(n651) );
  AND3X1 U840 ( .IN1(n242), .IN2(n246), .IN3(xmitH), .Q(n492) );
  AND2X1 U841 ( .IN1(test_se), .IN2(n699), .Q(n644) );
  OR2X1 U842 ( .IN1(n652), .IN2(n653), .Q(n119) );
  AND2X1 U843 ( .IN1(n696), .IN2(test_se), .Q(n653) );
  AND2X1 U844 ( .IN1(uart_REC_dataH), .IN2(n425), .Q(n652) );
  OR2X1 U845 ( .IN1(n654), .IN2(n655), .Q(n118) );
  AND2X1 U846 ( .IN1(rec_dataH_rec_7), .IN2(test_se), .Q(n655) );
  AND2X1 U847 ( .IN1(n691), .IN2(n425), .Q(n654) );
  INVX0 U848 ( .INP(test_se), .ZN(n425) );
  AND2X1 U849 ( .IN1(n639), .IN2(iXMIT_N24), .Q(iXMIT_N28) );
  OR2X1 U850 ( .IN1(n656), .IN2(n657), .Q(iXMIT_N27) );
  AND2X1 U851 ( .IN1(iXMIT_N26), .IN2(n703), .Q(n657) );
  AND3X1 U852 ( .IN1(n704), .IN2(n639), .IN3(n413), .Q(n656) );
  AND2X1 U853 ( .IN1(n411), .IN2(n639), .Q(iXMIT_N26) );
  OR2X1 U854 ( .IN1(n444), .IN2(n440), .Q(n639) );
  INVX0 U855 ( .INP(n417), .ZN(n440) );
  OR2X1 U856 ( .IN1(n239), .IN2(n242), .Q(n417) );
  AND2X1 U857 ( .IN1(n658), .IN2(iXMIT_state_1_temp), .Q(n444) );
  INVX0 U858 ( .INP(n439), .ZN(n658) );
  AND2X1 U859 ( .IN1(n700), .IN2(n475), .Q(n439) );
  AND4X1 U860 ( .IN1(n702), .IN2(n701), .IN3(n411), .IN4(n703), .Q(n475) );
  OR2X1 U861 ( .IN1(n659), .IN2(n660), .Q(iXMIT_N25) );
  INVX0 U862 ( .INP(n661), .ZN(n660) );
  OR2X1 U863 ( .IN1(n662), .IN2(n701), .Q(n661) );
  AND2X1 U864 ( .IN1(n701), .IN2(n662), .Q(n659) );
  AND2X1 U865 ( .IN1(n662), .IN2(n663), .Q(iXMIT_N24) );
  OR2X1 U866 ( .IN1(n702), .IN2(n664), .Q(n663) );
  AND2X1 U867 ( .IN1(n703), .IN2(n704), .Q(n664) );
  INVX0 U868 ( .INP(n528), .ZN(n662) );
  AND3X1 U869 ( .IN1(n703), .IN2(n704), .IN3(n702), .Q(n528) );
  AND2X1 U870 ( .IN1(iRECEIVER_state_1_), .IN2(n665), .Q(
        iRECEIVER_next_state_2_) );
  OR2X1 U871 ( .IN1(n666), .IN2(n667), .Q(iRECEIVER_N28) );
  INVX0 U872 ( .INP(n668), .ZN(n667) );
  OR2X1 U873 ( .IN1(n669), .IN2(n690), .Q(n668) );
  AND2X1 U874 ( .IN1(n690), .IN2(n669), .Q(n666) );
  AND2X1 U875 ( .IN1(n669), .IN2(n670), .Q(iRECEIVER_N27) );
  OR2X1 U876 ( .IN1(n697), .IN2(n671), .Q(n670) );
  AND2X1 U877 ( .IN1(n706), .IN2(n705), .Q(n671) );
  OR3X1 U878 ( .IN1(n406), .IN2(n404), .IN3(n408), .Q(n669) );
  OR2X1 U879 ( .IN1(n672), .IN2(n673), .Q(iRECEIVER_N26) );
  AND2X1 U880 ( .IN1(n706), .IN2(n404), .Q(n673) );
  AND2X1 U881 ( .IN1(n705), .IN2(n406), .Q(n672) );
  AND2X1 U882 ( .IN1(iRECEIVER_N19), .IN2(n674), .Q(iRECEIVER_N23) );
  AND2X1 U883 ( .IN1(n674), .IN2(iRECEIVER_N18), .Q(iRECEIVER_N22) );
  AND2X1 U884 ( .IN1(iRECEIVER_N17), .IN2(n674), .Q(iRECEIVER_N21) );
  AND2X1 U885 ( .IN1(n255), .IN2(n674), .Q(iRECEIVER_N20) );
  INVX0 U886 ( .INP(n675), .ZN(n674) );
  OR4X1 U887 ( .IN1(n676), .IN2(iRECEIVER_state_2_), .IN3(n241), .IN4(n665), 
        .Q(n675) );
  AND2X1 U888 ( .IN1(iRECEIVER_state_0_), .IN2(n549), .Q(n665) );
  AND4X1 U889 ( .IN1(n708), .IN2(n707), .IN3(iRECEIVER_bitCell_cntrH_1_), 
        .IN4(n255), .Q(n549) );
  AND2X1 U890 ( .IN1(n535), .IN2(n245), .Q(n676) );
  AND4X1 U891 ( .IN1(n255), .IN2(n708), .IN3(n409), .IN4(n244), .Q(n535) );
  INVX0 U892 ( .INP(n677), .ZN(iRECEIVER_N19) );
  AND2X1 U893 ( .IN1(n678), .IN2(n679), .Q(n677) );
  OR2X1 U894 ( .IN1(n680), .IN2(n707), .Q(n679) );
  OR2X1 U895 ( .IN1(n409), .IN2(n681), .Q(n678) );
  AND2X1 U896 ( .IN1(n680), .IN2(n682), .Q(iRECEIVER_N18) );
  OR2X1 U897 ( .IN1(n708), .IN2(n683), .Q(n682) );
  AND2X1 U898 ( .IN1(iRECEIVER_bitCell_cntrH_0_), .IN2(
        iRECEIVER_bitCell_cntrH_1_), .Q(n683) );
  INVX0 U899 ( .INP(n681), .ZN(n680) );
  AND3X1 U900 ( .IN1(iRECEIVER_bitCell_cntrH_0_), .IN2(
        iRECEIVER_bitCell_cntrH_1_), .IN3(n708), .Q(n681) );
  OR2X1 U901 ( .IN1(n684), .IN2(n685), .Q(iRECEIVER_N17) );
  AND2X1 U902 ( .IN1(n244), .IN2(iRECEIVER_bitCell_cntrH_0_), .Q(n685) );
  AND2X1 U903 ( .IN1(n255), .IN2(iRECEIVER_bitCell_cntrH_1_), .Q(n684) );
endmodule

