module add_mul_comp_sub_16_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, 
        a_7_, a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, 
        b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, 
        b_13_, b_14_, b_15_, Result_0_, Result_1_, Result_2_, Result_3_, 
        Result_4_, Result_5_, Result_6_, Result_7_, Result_8_, Result_9_, 
        Result_10_, Result_11_, Result_12_, Result_13_, Result_14_, Result_15_, 
        Result_16_, Result_17_, Result_18_, Result_19_, Result_20_, Result_21_, 
        Result_22_, Result_23_, Result_24_, Result_25_, Result_26_, Result_27_, 
        Result_28_, Result_29_, Result_30_, Result_31_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_,
         b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_;
  wire   Result_9_, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501;
  assign Result_8_ = Result_9_;
  assign Result_6_ = Result_9_;
  assign Result_4_ = Result_9_;
  assign Result_2_ = Result_9_;
  assign Result_15_ = Result_9_;
  assign Result_13_ = Result_9_;
  assign Result_11_ = Result_9_;
  assign Result_0_ = Result_9_;
  assign Result_10_ = Result_9_;
  assign Result_12_ = Result_9_;
  assign Result_14_ = Result_9_;
  assign Result_1_ = Result_9_;
  assign Result_3_ = Result_9_;
  assign Result_5_ = Result_9_;
  assign Result_7_ = Result_9_;

  NOR2_X1 U269 ( .A1(n252), .A2(n253), .ZN(Result_9_) );
  NOR2_X1 U270 ( .A1(n254), .A2(n255), .ZN(n253) );
  INV_X1 U271 ( .A(n256), .ZN(n255) );
  AND2_X1 U272 ( .A1(n257), .A2(n258), .ZN(n254) );
  XOR2_X1 U273 ( .A(b_15_), .B(a_15_), .Z(Result_31_) );
  NAND2_X1 U274 ( .A1(n259), .A2(n260), .ZN(Result_30_) );
  NAND4_X1 U275 ( .A1(n261), .A2(a_15_), .A3(n262), .A4(n263), .ZN(n260) );
  NOR2_X1 U276 ( .A1(n264), .A2(n265), .ZN(n261) );
  NOR2_X1 U277 ( .A1(b_15_), .A2(n266), .ZN(n265) );
  NOR2_X1 U278 ( .A1(n267), .A2(n268), .ZN(n264) );
  NAND3_X1 U279 ( .A1(n269), .A2(n270), .A3(n271), .ZN(n259) );
  XOR2_X1 U280 ( .A(b_14_), .B(a_14_), .Z(n271) );
  NAND3_X1 U281 ( .A1(n272), .A2(n268), .A3(a_15_), .ZN(n270) );
  NAND2_X1 U282 ( .A1(n273), .A2(n274), .ZN(n269) );
  NAND2_X1 U283 ( .A1(n275), .A2(n276), .ZN(Result_29_) );
  NAND2_X1 U284 ( .A1(n267), .A2(n277), .ZN(n276) );
  XOR2_X1 U285 ( .A(n278), .B(n279), .Z(n277) );
  NAND2_X1 U286 ( .A1(n280), .A2(n266), .ZN(n275) );
  XNOR2_X1 U287 ( .A(n281), .B(n278), .ZN(n280) );
  NAND2_X1 U288 ( .A1(n282), .A2(n283), .ZN(n278) );
  NAND2_X1 U289 ( .A1(n284), .A2(n285), .ZN(Result_28_) );
  NAND2_X1 U290 ( .A1(n267), .A2(n286), .ZN(n285) );
  XNOR2_X1 U291 ( .A(n287), .B(n288), .ZN(n286) );
  NAND2_X1 U292 ( .A1(n289), .A2(n266), .ZN(n284) );
  XOR2_X1 U293 ( .A(n290), .B(n287), .Z(n289) );
  AND2_X1 U294 ( .A1(n291), .A2(n292), .ZN(n287) );
  NAND2_X1 U295 ( .A1(n293), .A2(n294), .ZN(Result_27_) );
  NAND2_X1 U296 ( .A1(n267), .A2(n295), .ZN(n294) );
  XOR2_X1 U297 ( .A(n296), .B(n297), .Z(n295) );
  NAND2_X1 U298 ( .A1(n298), .A2(n266), .ZN(n293) );
  XNOR2_X1 U299 ( .A(n299), .B(n296), .ZN(n298) );
  NAND2_X1 U300 ( .A1(n300), .A2(n301), .ZN(n296) );
  NAND2_X1 U301 ( .A1(n302), .A2(n303), .ZN(Result_26_) );
  NAND2_X1 U302 ( .A1(n267), .A2(n304), .ZN(n303) );
  XNOR2_X1 U303 ( .A(n305), .B(n306), .ZN(n304) );
  NAND2_X1 U304 ( .A1(n307), .A2(n266), .ZN(n302) );
  XOR2_X1 U305 ( .A(n308), .B(n305), .Z(n307) );
  AND2_X1 U306 ( .A1(n309), .A2(n310), .ZN(n305) );
  NAND2_X1 U307 ( .A1(n311), .A2(n312), .ZN(Result_25_) );
  NAND2_X1 U308 ( .A1(n267), .A2(n313), .ZN(n312) );
  XOR2_X1 U309 ( .A(n314), .B(n315), .Z(n313) );
  NAND2_X1 U310 ( .A1(n316), .A2(n266), .ZN(n311) );
  XNOR2_X1 U311 ( .A(n317), .B(n314), .ZN(n316) );
  NAND2_X1 U312 ( .A1(n318), .A2(n319), .ZN(n314) );
  NAND2_X1 U313 ( .A1(n320), .A2(n321), .ZN(Result_24_) );
  NAND2_X1 U314 ( .A1(n267), .A2(n322), .ZN(n321) );
  XNOR2_X1 U315 ( .A(n323), .B(n324), .ZN(n322) );
  NAND2_X1 U316 ( .A1(n325), .A2(n266), .ZN(n320) );
  XOR2_X1 U317 ( .A(n326), .B(n323), .Z(n325) );
  AND2_X1 U318 ( .A1(n327), .A2(n328), .ZN(n323) );
  NAND2_X1 U319 ( .A1(n329), .A2(n330), .ZN(Result_23_) );
  NAND2_X1 U320 ( .A1(n267), .A2(n331), .ZN(n330) );
  XOR2_X1 U321 ( .A(n332), .B(n333), .Z(n331) );
  NAND2_X1 U322 ( .A1(n334), .A2(n266), .ZN(n329) );
  XNOR2_X1 U323 ( .A(n335), .B(n332), .ZN(n334) );
  NAND2_X1 U324 ( .A1(n336), .A2(n337), .ZN(n332) );
  NAND2_X1 U325 ( .A1(n338), .A2(n339), .ZN(Result_22_) );
  NAND2_X1 U326 ( .A1(n267), .A2(n340), .ZN(n339) );
  XNOR2_X1 U327 ( .A(n341), .B(n342), .ZN(n340) );
  NAND2_X1 U328 ( .A1(n343), .A2(n266), .ZN(n338) );
  XOR2_X1 U329 ( .A(n344), .B(n341), .Z(n343) );
  AND2_X1 U330 ( .A1(n345), .A2(n346), .ZN(n341) );
  NAND2_X1 U331 ( .A1(n347), .A2(n348), .ZN(Result_21_) );
  NAND2_X1 U332 ( .A1(n267), .A2(n349), .ZN(n348) );
  XOR2_X1 U333 ( .A(n350), .B(n351), .Z(n349) );
  NAND2_X1 U334 ( .A1(n352), .A2(n266), .ZN(n347) );
  XNOR2_X1 U335 ( .A(n353), .B(n350), .ZN(n352) );
  NAND2_X1 U336 ( .A1(n354), .A2(n355), .ZN(n350) );
  NAND2_X1 U337 ( .A1(n356), .A2(n357), .ZN(Result_20_) );
  NAND2_X1 U338 ( .A1(n267), .A2(n358), .ZN(n357) );
  XNOR2_X1 U339 ( .A(n359), .B(n360), .ZN(n358) );
  NAND2_X1 U340 ( .A1(n361), .A2(n266), .ZN(n356) );
  XOR2_X1 U341 ( .A(n362), .B(n359), .Z(n361) );
  AND2_X1 U342 ( .A1(n363), .A2(n364), .ZN(n359) );
  NAND2_X1 U343 ( .A1(n365), .A2(n366), .ZN(Result_19_) );
  NAND2_X1 U344 ( .A1(n267), .A2(n367), .ZN(n366) );
  XOR2_X1 U345 ( .A(n368), .B(n369), .Z(n367) );
  NAND2_X1 U346 ( .A1(n370), .A2(n266), .ZN(n365) );
  XNOR2_X1 U347 ( .A(n371), .B(n368), .ZN(n370) );
  NAND2_X1 U348 ( .A1(n372), .A2(n373), .ZN(n368) );
  NAND2_X1 U349 ( .A1(n374), .A2(n375), .ZN(Result_18_) );
  NAND2_X1 U350 ( .A1(n267), .A2(n376), .ZN(n375) );
  XNOR2_X1 U351 ( .A(n377), .B(n378), .ZN(n376) );
  NAND2_X1 U352 ( .A1(n379), .A2(n266), .ZN(n374) );
  XOR2_X1 U353 ( .A(n380), .B(n377), .Z(n379) );
  AND2_X1 U354 ( .A1(n381), .A2(n382), .ZN(n377) );
  NAND2_X1 U355 ( .A1(n383), .A2(n384), .ZN(Result_17_) );
  NAND2_X1 U356 ( .A1(n267), .A2(n385), .ZN(n384) );
  XOR2_X1 U357 ( .A(n386), .B(n387), .Z(n385) );
  NAND2_X1 U358 ( .A1(n388), .A2(n266), .ZN(n383) );
  XNOR2_X1 U359 ( .A(n389), .B(n386), .ZN(n388) );
  NAND2_X1 U360 ( .A1(n257), .A2(n390), .ZN(n386) );
  NAND2_X1 U361 ( .A1(n391), .A2(n392), .ZN(Result_16_) );
  NAND2_X1 U362 ( .A1(n267), .A2(n393), .ZN(n392) );
  XNOR2_X1 U363 ( .A(n394), .B(n395), .ZN(n393) );
  NOR2_X1 U364 ( .A1(n396), .A2(n397), .ZN(n395) );
  AND2_X1 U365 ( .A1(n387), .A2(a_1_), .ZN(n397) );
  NOR2_X1 U366 ( .A1(n398), .A2(n399), .ZN(n396) );
  NOR2_X1 U367 ( .A1(a_1_), .A2(n387), .ZN(n398) );
  NAND2_X1 U368 ( .A1(n400), .A2(n401), .ZN(n387) );
  NAND2_X1 U369 ( .A1(b_2_), .A2(n402), .ZN(n401) );
  OR2_X1 U370 ( .A1(n378), .A2(a_2_), .ZN(n402) );
  NAND2_X1 U371 ( .A1(a_2_), .A2(n378), .ZN(n400) );
  NAND2_X1 U372 ( .A1(n403), .A2(n404), .ZN(n378) );
  NAND2_X1 U373 ( .A1(b_3_), .A2(n405), .ZN(n404) );
  OR2_X1 U374 ( .A1(n369), .A2(a_3_), .ZN(n405) );
  NAND2_X1 U375 ( .A1(a_3_), .A2(n369), .ZN(n403) );
  NAND2_X1 U376 ( .A1(n406), .A2(n407), .ZN(n369) );
  NAND2_X1 U377 ( .A1(b_4_), .A2(n408), .ZN(n407) );
  OR2_X1 U378 ( .A1(n360), .A2(a_4_), .ZN(n408) );
  NAND2_X1 U379 ( .A1(a_4_), .A2(n360), .ZN(n406) );
  NAND2_X1 U380 ( .A1(n409), .A2(n410), .ZN(n360) );
  NAND2_X1 U381 ( .A1(b_5_), .A2(n411), .ZN(n410) );
  OR2_X1 U382 ( .A1(n351), .A2(a_5_), .ZN(n411) );
  NAND2_X1 U383 ( .A1(a_5_), .A2(n351), .ZN(n409) );
  NAND2_X1 U384 ( .A1(n412), .A2(n413), .ZN(n351) );
  NAND2_X1 U385 ( .A1(b_6_), .A2(n414), .ZN(n413) );
  OR2_X1 U386 ( .A1(n342), .A2(a_6_), .ZN(n414) );
  NAND2_X1 U387 ( .A1(a_6_), .A2(n342), .ZN(n412) );
  NAND2_X1 U388 ( .A1(n415), .A2(n416), .ZN(n342) );
  NAND2_X1 U389 ( .A1(b_7_), .A2(n417), .ZN(n416) );
  OR2_X1 U390 ( .A1(n333), .A2(a_7_), .ZN(n417) );
  NAND2_X1 U391 ( .A1(a_7_), .A2(n333), .ZN(n415) );
  NAND2_X1 U392 ( .A1(n418), .A2(n419), .ZN(n333) );
  NAND2_X1 U393 ( .A1(b_8_), .A2(n420), .ZN(n419) );
  OR2_X1 U394 ( .A1(n324), .A2(a_8_), .ZN(n420) );
  NAND2_X1 U395 ( .A1(a_8_), .A2(n324), .ZN(n418) );
  NAND2_X1 U396 ( .A1(n421), .A2(n422), .ZN(n324) );
  NAND2_X1 U397 ( .A1(b_9_), .A2(n423), .ZN(n422) );
  OR2_X1 U398 ( .A1(n315), .A2(a_9_), .ZN(n423) );
  NAND2_X1 U399 ( .A1(a_9_), .A2(n315), .ZN(n421) );
  NAND2_X1 U400 ( .A1(n424), .A2(n425), .ZN(n315) );
  NAND2_X1 U401 ( .A1(b_10_), .A2(n426), .ZN(n425) );
  OR2_X1 U402 ( .A1(n306), .A2(a_10_), .ZN(n426) );
  NAND2_X1 U403 ( .A1(a_10_), .A2(n306), .ZN(n424) );
  NAND2_X1 U404 ( .A1(n427), .A2(n428), .ZN(n306) );
  NAND2_X1 U405 ( .A1(b_11_), .A2(n429), .ZN(n428) );
  OR2_X1 U406 ( .A1(n297), .A2(a_11_), .ZN(n429) );
  NAND2_X1 U407 ( .A1(a_11_), .A2(n297), .ZN(n427) );
  NAND2_X1 U408 ( .A1(n430), .A2(n431), .ZN(n297) );
  NAND2_X1 U409 ( .A1(b_12_), .A2(n432), .ZN(n431) );
  OR2_X1 U410 ( .A1(n288), .A2(a_12_), .ZN(n432) );
  NAND2_X1 U411 ( .A1(a_12_), .A2(n288), .ZN(n430) );
  NAND2_X1 U412 ( .A1(n433), .A2(n434), .ZN(n288) );
  NAND2_X1 U413 ( .A1(b_13_), .A2(n435), .ZN(n434) );
  OR2_X1 U414 ( .A1(n279), .A2(a_13_), .ZN(n435) );
  NAND2_X1 U415 ( .A1(a_13_), .A2(n279), .ZN(n433) );
  NAND2_X1 U416 ( .A1(n436), .A2(n437), .ZN(n279) );
  NAND2_X1 U417 ( .A1(b_14_), .A2(n438), .ZN(n437) );
  OR2_X1 U418 ( .A1(a_14_), .A2(n273), .ZN(n438) );
  NAND2_X1 U419 ( .A1(n273), .A2(a_14_), .ZN(n436) );
  AND2_X1 U420 ( .A1(b_15_), .A2(a_15_), .ZN(n273) );
  INV_X1 U421 ( .A(n272), .ZN(n267) );
  NAND2_X1 U422 ( .A1(n274), .A2(n439), .ZN(n272) );
  NAND4_X1 U423 ( .A1(n440), .A2(n441), .A3(n442), .A4(n443), .ZN(n439) );
  NOR4_X1 U424 ( .A1(n444), .A2(n445), .A3(n446), .A4(n447), .ZN(n443) );
  NOR4_X1 U425 ( .A1(n448), .A2(n449), .A3(n450), .A4(n451), .ZN(n442) );
  NOR4_X1 U426 ( .A1(n452), .A2(n453), .A3(n454), .A4(n455), .ZN(n441) );
  NOR4_X1 U427 ( .A1(n456), .A2(n252), .A3(n457), .A4(n458), .ZN(n440) );
  NOR2_X1 U428 ( .A1(a_15_), .A2(n268), .ZN(n458) );
  INV_X1 U429 ( .A(n266), .ZN(n274) );
  NAND2_X1 U430 ( .A1(n459), .A2(n266), .ZN(n391) );
  NAND2_X1 U431 ( .A1(n256), .A2(n460), .ZN(n266) );
  NAND2_X1 U432 ( .A1(n461), .A2(n462), .ZN(n460) );
  NAND2_X1 U433 ( .A1(n390), .A2(n463), .ZN(n461) );
  NAND3_X1 U434 ( .A1(n257), .A2(n381), .A3(n464), .ZN(n463) );
  NAND3_X1 U435 ( .A1(n382), .A2(n465), .A3(n373), .ZN(n464) );
  NAND3_X1 U436 ( .A1(n363), .A2(n372), .A3(n466), .ZN(n465) );
  NAND3_X1 U437 ( .A1(n364), .A2(n467), .A3(n355), .ZN(n466) );
  NAND3_X1 U438 ( .A1(n345), .A2(n354), .A3(n468), .ZN(n467) );
  NAND3_X1 U439 ( .A1(n346), .A2(n469), .A3(n337), .ZN(n468) );
  NAND3_X1 U440 ( .A1(n327), .A2(n336), .A3(n470), .ZN(n469) );
  NAND3_X1 U441 ( .A1(n328), .A2(n471), .A3(n319), .ZN(n470) );
  NAND3_X1 U442 ( .A1(n309), .A2(n318), .A3(n472), .ZN(n471) );
  NAND3_X1 U443 ( .A1(n310), .A2(n473), .A3(n301), .ZN(n472) );
  OR2_X1 U444 ( .A1(n299), .A2(n453), .ZN(n473) );
  NAND3_X1 U445 ( .A1(n258), .A2(n257), .A3(n394), .ZN(n459) );
  NAND2_X1 U446 ( .A1(n462), .A2(n256), .ZN(n394) );
  NAND2_X1 U447 ( .A1(a_0_), .A2(n474), .ZN(n256) );
  INV_X1 U448 ( .A(n252), .ZN(n462) );
  NOR2_X1 U449 ( .A1(n474), .A2(a_0_), .ZN(n252) );
  INV_X1 U450 ( .A(b_0_), .ZN(n474) );
  INV_X1 U451 ( .A(n457), .ZN(n257) );
  NOR2_X1 U452 ( .A1(n399), .A2(a_1_), .ZN(n457) );
  NAND2_X1 U453 ( .A1(n389), .A2(n390), .ZN(n258) );
  NAND2_X1 U454 ( .A1(a_1_), .A2(n399), .ZN(n390) );
  INV_X1 U455 ( .A(b_1_), .ZN(n399) );
  NAND2_X1 U456 ( .A1(n381), .A2(n475), .ZN(n389) );
  NAND2_X1 U457 ( .A1(n382), .A2(n380), .ZN(n475) );
  NAND2_X1 U458 ( .A1(n372), .A2(n476), .ZN(n380) );
  NAND2_X1 U459 ( .A1(n373), .A2(n371), .ZN(n476) );
  NAND2_X1 U460 ( .A1(n363), .A2(n477), .ZN(n371) );
  NAND2_X1 U461 ( .A1(n364), .A2(n362), .ZN(n477) );
  NAND2_X1 U462 ( .A1(n354), .A2(n478), .ZN(n362) );
  NAND2_X1 U463 ( .A1(n355), .A2(n353), .ZN(n478) );
  NAND2_X1 U464 ( .A1(n345), .A2(n479), .ZN(n353) );
  NAND2_X1 U465 ( .A1(n346), .A2(n344), .ZN(n479) );
  NAND2_X1 U466 ( .A1(n336), .A2(n480), .ZN(n344) );
  NAND2_X1 U467 ( .A1(n337), .A2(n335), .ZN(n480) );
  NAND2_X1 U468 ( .A1(n327), .A2(n481), .ZN(n335) );
  NAND2_X1 U469 ( .A1(n328), .A2(n326), .ZN(n481) );
  NAND2_X1 U470 ( .A1(n318), .A2(n482), .ZN(n326) );
  NAND2_X1 U471 ( .A1(n319), .A2(n317), .ZN(n482) );
  NAND2_X1 U472 ( .A1(n309), .A2(n483), .ZN(n317) );
  NAND2_X1 U473 ( .A1(n310), .A2(n308), .ZN(n483) );
  NAND2_X1 U474 ( .A1(n300), .A2(n484), .ZN(n308) );
  NAND2_X1 U475 ( .A1(n301), .A2(n299), .ZN(n484) );
  NAND2_X1 U476 ( .A1(n291), .A2(n485), .ZN(n299) );
  NAND2_X1 U477 ( .A1(n292), .A2(n290), .ZN(n485) );
  NAND2_X1 U478 ( .A1(n282), .A2(n486), .ZN(n290) );
  NAND2_X1 U479 ( .A1(n283), .A2(n281), .ZN(n486) );
  NAND2_X1 U480 ( .A1(n263), .A2(n487), .ZN(n281) );
  NAND2_X1 U481 ( .A1(n488), .A2(n262), .ZN(n487) );
  NAND2_X1 U482 ( .A1(a_14_), .A2(n489), .ZN(n262) );
  NAND2_X1 U483 ( .A1(a_15_), .A2(n268), .ZN(n488) );
  INV_X1 U484 ( .A(b_15_), .ZN(n268) );
  INV_X1 U485 ( .A(n455), .ZN(n263) );
  NOR2_X1 U486 ( .A1(n489), .A2(a_14_), .ZN(n455) );
  INV_X1 U487 ( .A(b_14_), .ZN(n489) );
  NAND2_X1 U488 ( .A1(a_13_), .A2(n490), .ZN(n283) );
  INV_X1 U489 ( .A(n456), .ZN(n282) );
  NOR2_X1 U490 ( .A1(n490), .A2(a_13_), .ZN(n456) );
  INV_X1 U491 ( .A(b_13_), .ZN(n490) );
  NAND2_X1 U492 ( .A1(a_12_), .A2(n491), .ZN(n292) );
  INV_X1 U493 ( .A(n454), .ZN(n291) );
  NOR2_X1 U494 ( .A1(n491), .A2(a_12_), .ZN(n454) );
  INV_X1 U495 ( .A(b_12_), .ZN(n491) );
  NAND2_X1 U496 ( .A1(a_11_), .A2(n492), .ZN(n301) );
  INV_X1 U497 ( .A(n453), .ZN(n300) );
  NOR2_X1 U498 ( .A1(n492), .A2(a_11_), .ZN(n453) );
  INV_X1 U499 ( .A(b_11_), .ZN(n492) );
  NAND2_X1 U500 ( .A1(a_10_), .A2(n493), .ZN(n310) );
  INV_X1 U501 ( .A(n452), .ZN(n309) );
  NOR2_X1 U502 ( .A1(n493), .A2(a_10_), .ZN(n452) );
  INV_X1 U503 ( .A(b_10_), .ZN(n493) );
  NAND2_X1 U504 ( .A1(a_9_), .A2(n494), .ZN(n319) );
  INV_X1 U505 ( .A(n451), .ZN(n318) );
  NOR2_X1 U506 ( .A1(n494), .A2(a_9_), .ZN(n451) );
  INV_X1 U507 ( .A(b_9_), .ZN(n494) );
  NAND2_X1 U508 ( .A1(a_8_), .A2(n495), .ZN(n328) );
  INV_X1 U509 ( .A(n450), .ZN(n327) );
  NOR2_X1 U510 ( .A1(n495), .A2(a_8_), .ZN(n450) );
  INV_X1 U511 ( .A(b_8_), .ZN(n495) );
  NAND2_X1 U512 ( .A1(a_7_), .A2(n496), .ZN(n337) );
  INV_X1 U513 ( .A(n449), .ZN(n336) );
  NOR2_X1 U514 ( .A1(n496), .A2(a_7_), .ZN(n449) );
  INV_X1 U515 ( .A(b_7_), .ZN(n496) );
  NAND2_X1 U516 ( .A1(a_6_), .A2(n497), .ZN(n346) );
  INV_X1 U517 ( .A(n448), .ZN(n345) );
  NOR2_X1 U518 ( .A1(n497), .A2(a_6_), .ZN(n448) );
  INV_X1 U519 ( .A(b_6_), .ZN(n497) );
  NAND2_X1 U520 ( .A1(a_5_), .A2(n498), .ZN(n355) );
  INV_X1 U521 ( .A(n447), .ZN(n354) );
  NOR2_X1 U522 ( .A1(n498), .A2(a_5_), .ZN(n447) );
  INV_X1 U523 ( .A(b_5_), .ZN(n498) );
  NAND2_X1 U524 ( .A1(a_4_), .A2(n499), .ZN(n364) );
  INV_X1 U525 ( .A(n446), .ZN(n363) );
  NOR2_X1 U526 ( .A1(n499), .A2(a_4_), .ZN(n446) );
  INV_X1 U527 ( .A(b_4_), .ZN(n499) );
  NAND2_X1 U528 ( .A1(a_3_), .A2(n500), .ZN(n373) );
  INV_X1 U529 ( .A(n445), .ZN(n372) );
  NOR2_X1 U530 ( .A1(n500), .A2(a_3_), .ZN(n445) );
  INV_X1 U531 ( .A(b_3_), .ZN(n500) );
  NAND2_X1 U532 ( .A1(a_2_), .A2(n501), .ZN(n382) );
  INV_X1 U533 ( .A(n444), .ZN(n381) );
  NOR2_X1 U534 ( .A1(n501), .A2(a_2_), .ZN(n444) );
  INV_X1 U535 ( .A(b_2_), .ZN(n501) );
endmodule

