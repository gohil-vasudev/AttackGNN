module add_mul_comp_sub_32_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, 
        a_7_, a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, 
        a_17_, a_18_, a_19_, a_20_, a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, 
        a_27_, a_28_, a_29_, a_30_, a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, 
        b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, 
        b_16_, b_17_, b_18_, b_19_, b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, 
        b_26_, b_27_, b_28_, b_29_, b_30_, b_31_, Result_0_, Result_1_, 
        Result_2_, Result_3_, Result_4_, Result_5_, Result_6_, Result_7_, 
        Result_8_, Result_9_, Result_10_, Result_11_, Result_12_, Result_13_, 
        Result_14_, Result_15_, Result_16_, Result_17_, Result_18_, Result_19_, 
        Result_20_, Result_21_, Result_22_, Result_23_, Result_24_, Result_25_, 
        Result_26_, Result_27_, Result_28_, Result_29_, Result_30_, Result_31_, 
        Result_32_, Result_33_, Result_34_, Result_35_, Result_36_, Result_37_, 
        Result_38_, Result_39_, Result_40_, Result_41_, Result_42_, Result_43_, 
        Result_44_, Result_45_, Result_46_, Result_47_, Result_48_, Result_49_, 
        Result_50_, Result_51_, Result_52_, Result_53_, Result_54_, Result_55_, 
        Result_56_, Result_57_, Result_58_, Result_59_, Result_60_, Result_61_, 
        Result_62_, Result_63_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, a_19_, a_20_,
         a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, a_29_, a_30_,
         a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_,
         b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, b_18_, b_19_,
         b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, b_28_, b_29_,
         b_30_, b_31_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_,
         Result_32_, Result_33_, Result_34_, Result_35_, Result_36_,
         Result_37_, Result_38_, Result_39_, Result_40_, Result_41_,
         Result_42_, Result_43_, Result_44_, Result_45_, Result_46_,
         Result_47_, Result_48_, Result_49_, Result_50_, Result_51_,
         Result_52_, Result_53_, Result_54_, Result_55_, Result_56_,
         Result_57_, Result_58_, Result_59_, Result_60_, Result_61_,
         Result_62_, Result_63_;
  wire   Result_9_, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095;
  assign Result_8_ = Result_9_;
  assign Result_6_ = Result_9_;
  assign Result_4_ = Result_9_;
  assign Result_31_ = Result_9_;
  assign Result_2_ = Result_9_;
  assign Result_28_ = Result_9_;
  assign Result_26_ = Result_9_;
  assign Result_24_ = Result_9_;
  assign Result_22_ = Result_9_;
  assign Result_20_ = Result_9_;
  assign Result_19_ = Result_9_;
  assign Result_17_ = Result_9_;
  assign Result_15_ = Result_9_;
  assign Result_13_ = Result_9_;
  assign Result_11_ = Result_9_;
  assign Result_0_ = Result_9_;
  assign Result_10_ = Result_9_;
  assign Result_12_ = Result_9_;
  assign Result_14_ = Result_9_;
  assign Result_16_ = Result_9_;
  assign Result_18_ = Result_9_;
  assign Result_1_ = Result_9_;
  assign Result_21_ = Result_9_;
  assign Result_23_ = Result_9_;
  assign Result_25_ = Result_9_;
  assign Result_27_ = Result_9_;
  assign Result_29_ = Result_9_;
  assign Result_30_ = Result_9_;
  assign Result_3_ = Result_9_;
  assign Result_5_ = Result_9_;
  assign Result_7_ = Result_9_;

  OR2_X2 U582 ( .A1(n908), .A2(n909), .ZN(Result_9_) );
  OR2_X1 U583 ( .A1(n549), .A2(n550), .ZN(Result_63_) );
  OR2_X1 U584 ( .A1(n551), .A2(n552), .ZN(Result_62_) );
  AND2_X1 U585 ( .A1(n553), .A2(n554), .ZN(n552) );
  OR2_X1 U586 ( .A1(n555), .A2(n556), .ZN(n554) );
  AND2_X1 U587 ( .A1(Result_9_), .A2(n557), .ZN(n556) );
  AND2_X1 U588 ( .A1(n558), .A2(n559), .ZN(n555) );
  OR2_X1 U589 ( .A1(n560), .A2(n561), .ZN(n559) );
  INV_X1 U590 ( .A(b_31_), .ZN(n561) );
  AND2_X1 U591 ( .A1(n562), .A2(n563), .ZN(n551) );
  OR2_X1 U592 ( .A1(n564), .A2(n565), .ZN(n563) );
  AND2_X1 U593 ( .A1(n549), .A2(Result_9_), .ZN(n565) );
  AND3_X1 U594 ( .A1(b_31_), .A2(a_31_), .A3(n558), .ZN(n564) );
  INV_X1 U595 ( .A(n553), .ZN(n562) );
  OR2_X1 U596 ( .A1(n566), .A2(n567), .ZN(n553) );
  INV_X1 U597 ( .A(n568), .ZN(n567) );
  OR2_X1 U598 ( .A1(n569), .A2(n570), .ZN(Result_61_) );
  AND2_X1 U599 ( .A1(n571), .A2(Result_9_), .ZN(n570) );
  XOR2_X1 U600 ( .A(n572), .B(n573), .Z(n571) );
  AND2_X1 U601 ( .A1(n558), .A2(n574), .ZN(n569) );
  XOR2_X1 U602 ( .A(n573), .B(n575), .Z(n574) );
  OR2_X1 U603 ( .A1(n576), .A2(n577), .ZN(n573) );
  INV_X1 U604 ( .A(n578), .ZN(n577) );
  OR2_X1 U605 ( .A1(n579), .A2(n580), .ZN(Result_60_) );
  AND2_X1 U606 ( .A1(n581), .A2(Result_9_), .ZN(n580) );
  XOR2_X1 U607 ( .A(n582), .B(n583), .Z(n581) );
  AND2_X1 U608 ( .A1(n584), .A2(n558), .ZN(n579) );
  XNOR2_X1 U609 ( .A(n583), .B(n585), .ZN(n584) );
  OR2_X1 U610 ( .A1(n586), .A2(n587), .ZN(n583) );
  INV_X1 U611 ( .A(n588), .ZN(n587) );
  OR2_X1 U612 ( .A1(n589), .A2(n590), .ZN(Result_59_) );
  AND2_X1 U613 ( .A1(n591), .A2(Result_9_), .ZN(n590) );
  XOR2_X1 U614 ( .A(n592), .B(n593), .Z(n591) );
  AND2_X1 U615 ( .A1(n594), .A2(n558), .ZN(n589) );
  XNOR2_X1 U616 ( .A(n593), .B(n595), .ZN(n594) );
  OR2_X1 U617 ( .A1(n596), .A2(n597), .ZN(n593) );
  INV_X1 U618 ( .A(n598), .ZN(n597) );
  OR2_X1 U619 ( .A1(n599), .A2(n600), .ZN(Result_58_) );
  AND2_X1 U620 ( .A1(n601), .A2(Result_9_), .ZN(n600) );
  XOR2_X1 U621 ( .A(n602), .B(n603), .Z(n601) );
  AND2_X1 U622 ( .A1(n604), .A2(n558), .ZN(n599) );
  XNOR2_X1 U623 ( .A(n603), .B(n605), .ZN(n604) );
  OR2_X1 U624 ( .A1(n606), .A2(n607), .ZN(n603) );
  INV_X1 U625 ( .A(n608), .ZN(n607) );
  OR2_X1 U626 ( .A1(n609), .A2(n610), .ZN(Result_57_) );
  AND2_X1 U627 ( .A1(n611), .A2(Result_9_), .ZN(n610) );
  XOR2_X1 U628 ( .A(n612), .B(n613), .Z(n611) );
  AND2_X1 U629 ( .A1(n614), .A2(n558), .ZN(n609) );
  XNOR2_X1 U630 ( .A(n613), .B(n615), .ZN(n614) );
  OR2_X1 U631 ( .A1(n616), .A2(n617), .ZN(n613) );
  INV_X1 U632 ( .A(n618), .ZN(n617) );
  OR2_X1 U633 ( .A1(n619), .A2(n620), .ZN(Result_56_) );
  AND2_X1 U634 ( .A1(n621), .A2(Result_9_), .ZN(n620) );
  XOR2_X1 U635 ( .A(n622), .B(n623), .Z(n621) );
  AND2_X1 U636 ( .A1(n624), .A2(n558), .ZN(n619) );
  XNOR2_X1 U637 ( .A(n623), .B(n625), .ZN(n624) );
  OR2_X1 U638 ( .A1(n626), .A2(n627), .ZN(n623) );
  INV_X1 U639 ( .A(n628), .ZN(n627) );
  OR2_X1 U640 ( .A1(n629), .A2(n630), .ZN(Result_55_) );
  AND2_X1 U641 ( .A1(n631), .A2(Result_9_), .ZN(n630) );
  XOR2_X1 U642 ( .A(n632), .B(n633), .Z(n631) );
  AND2_X1 U643 ( .A1(n634), .A2(n558), .ZN(n629) );
  XNOR2_X1 U644 ( .A(n633), .B(n635), .ZN(n634) );
  OR2_X1 U645 ( .A1(n636), .A2(n637), .ZN(n633) );
  INV_X1 U646 ( .A(n638), .ZN(n637) );
  OR2_X1 U647 ( .A1(n639), .A2(n640), .ZN(Result_54_) );
  AND2_X1 U648 ( .A1(n641), .A2(Result_9_), .ZN(n640) );
  XOR2_X1 U649 ( .A(n642), .B(n643), .Z(n641) );
  AND2_X1 U650 ( .A1(n644), .A2(n558), .ZN(n639) );
  XNOR2_X1 U651 ( .A(n643), .B(n645), .ZN(n644) );
  OR2_X1 U652 ( .A1(n646), .A2(n647), .ZN(n643) );
  INV_X1 U653 ( .A(n648), .ZN(n647) );
  OR2_X1 U654 ( .A1(n649), .A2(n650), .ZN(Result_53_) );
  AND2_X1 U655 ( .A1(n651), .A2(Result_9_), .ZN(n650) );
  XOR2_X1 U656 ( .A(n652), .B(n653), .Z(n651) );
  AND2_X1 U657 ( .A1(n654), .A2(n558), .ZN(n649) );
  XNOR2_X1 U658 ( .A(n653), .B(n655), .ZN(n654) );
  OR2_X1 U659 ( .A1(n656), .A2(n657), .ZN(n653) );
  INV_X1 U660 ( .A(n658), .ZN(n657) );
  OR2_X1 U661 ( .A1(n659), .A2(n660), .ZN(Result_52_) );
  AND2_X1 U662 ( .A1(n661), .A2(Result_9_), .ZN(n660) );
  XOR2_X1 U663 ( .A(n662), .B(n663), .Z(n661) );
  AND2_X1 U664 ( .A1(n664), .A2(n558), .ZN(n659) );
  XNOR2_X1 U665 ( .A(n663), .B(n665), .ZN(n664) );
  OR2_X1 U666 ( .A1(n666), .A2(n667), .ZN(n663) );
  INV_X1 U667 ( .A(n668), .ZN(n667) );
  OR2_X1 U668 ( .A1(n669), .A2(n670), .ZN(Result_51_) );
  AND2_X1 U669 ( .A1(n671), .A2(Result_9_), .ZN(n670) );
  XOR2_X1 U670 ( .A(n672), .B(n673), .Z(n671) );
  AND2_X1 U671 ( .A1(n674), .A2(n558), .ZN(n669) );
  XNOR2_X1 U672 ( .A(n673), .B(n675), .ZN(n674) );
  OR2_X1 U673 ( .A1(n676), .A2(n677), .ZN(n673) );
  INV_X1 U674 ( .A(n678), .ZN(n677) );
  OR2_X1 U675 ( .A1(n679), .A2(n680), .ZN(Result_50_) );
  AND2_X1 U676 ( .A1(n681), .A2(Result_9_), .ZN(n680) );
  XOR2_X1 U677 ( .A(n682), .B(n683), .Z(n681) );
  AND2_X1 U678 ( .A1(n684), .A2(n558), .ZN(n679) );
  XNOR2_X1 U679 ( .A(n683), .B(n685), .ZN(n684) );
  OR2_X1 U680 ( .A1(n686), .A2(n687), .ZN(n683) );
  INV_X1 U681 ( .A(n688), .ZN(n687) );
  OR2_X1 U682 ( .A1(n689), .A2(n690), .ZN(Result_49_) );
  AND2_X1 U683 ( .A1(n691), .A2(Result_9_), .ZN(n690) );
  XOR2_X1 U684 ( .A(n692), .B(n693), .Z(n691) );
  AND2_X1 U685 ( .A1(n694), .A2(n558), .ZN(n689) );
  XNOR2_X1 U686 ( .A(n693), .B(n695), .ZN(n694) );
  OR2_X1 U687 ( .A1(n696), .A2(n697), .ZN(n693) );
  INV_X1 U688 ( .A(n698), .ZN(n697) );
  OR2_X1 U689 ( .A1(n699), .A2(n700), .ZN(Result_48_) );
  AND2_X1 U690 ( .A1(n701), .A2(Result_9_), .ZN(n700) );
  XOR2_X1 U691 ( .A(n702), .B(n703), .Z(n701) );
  AND2_X1 U692 ( .A1(n704), .A2(n558), .ZN(n699) );
  XNOR2_X1 U693 ( .A(n703), .B(n705), .ZN(n704) );
  OR2_X1 U694 ( .A1(n706), .A2(n707), .ZN(n703) );
  INV_X1 U695 ( .A(n708), .ZN(n707) );
  OR2_X1 U696 ( .A1(n709), .A2(n710), .ZN(Result_47_) );
  AND2_X1 U697 ( .A1(n711), .A2(Result_9_), .ZN(n710) );
  XOR2_X1 U698 ( .A(n712), .B(n713), .Z(n711) );
  AND2_X1 U699 ( .A1(n714), .A2(n558), .ZN(n709) );
  XNOR2_X1 U700 ( .A(n713), .B(n715), .ZN(n714) );
  OR2_X1 U701 ( .A1(n716), .A2(n717), .ZN(n713) );
  INV_X1 U702 ( .A(n718), .ZN(n717) );
  OR2_X1 U703 ( .A1(n719), .A2(n720), .ZN(Result_46_) );
  AND2_X1 U704 ( .A1(n721), .A2(Result_9_), .ZN(n720) );
  XOR2_X1 U705 ( .A(n722), .B(n723), .Z(n721) );
  AND2_X1 U706 ( .A1(n724), .A2(n558), .ZN(n719) );
  XNOR2_X1 U707 ( .A(n723), .B(n725), .ZN(n724) );
  OR2_X1 U708 ( .A1(n726), .A2(n727), .ZN(n723) );
  INV_X1 U709 ( .A(n728), .ZN(n727) );
  OR2_X1 U710 ( .A1(n729), .A2(n730), .ZN(Result_45_) );
  AND2_X1 U711 ( .A1(n731), .A2(Result_9_), .ZN(n730) );
  XOR2_X1 U712 ( .A(n732), .B(n733), .Z(n731) );
  AND2_X1 U713 ( .A1(n734), .A2(n558), .ZN(n729) );
  XNOR2_X1 U714 ( .A(n733), .B(n735), .ZN(n734) );
  OR2_X1 U715 ( .A1(n736), .A2(n737), .ZN(n733) );
  INV_X1 U716 ( .A(n738), .ZN(n737) );
  OR2_X1 U717 ( .A1(n739), .A2(n740), .ZN(Result_44_) );
  AND2_X1 U718 ( .A1(n741), .A2(Result_9_), .ZN(n740) );
  XOR2_X1 U719 ( .A(n742), .B(n743), .Z(n741) );
  AND2_X1 U720 ( .A1(n744), .A2(n558), .ZN(n739) );
  XNOR2_X1 U721 ( .A(n743), .B(n745), .ZN(n744) );
  OR2_X1 U722 ( .A1(n746), .A2(n747), .ZN(n743) );
  INV_X1 U723 ( .A(n748), .ZN(n747) );
  OR2_X1 U724 ( .A1(n749), .A2(n750), .ZN(Result_43_) );
  AND2_X1 U725 ( .A1(n751), .A2(Result_9_), .ZN(n750) );
  XOR2_X1 U726 ( .A(n752), .B(n753), .Z(n751) );
  AND2_X1 U727 ( .A1(n754), .A2(n558), .ZN(n749) );
  XNOR2_X1 U728 ( .A(n753), .B(n755), .ZN(n754) );
  OR2_X1 U729 ( .A1(n756), .A2(n757), .ZN(n753) );
  INV_X1 U730 ( .A(n758), .ZN(n757) );
  OR2_X1 U731 ( .A1(n759), .A2(n760), .ZN(Result_42_) );
  AND2_X1 U732 ( .A1(n761), .A2(Result_9_), .ZN(n760) );
  XOR2_X1 U733 ( .A(n762), .B(n763), .Z(n761) );
  AND2_X1 U734 ( .A1(n764), .A2(n558), .ZN(n759) );
  XNOR2_X1 U735 ( .A(n763), .B(n765), .ZN(n764) );
  OR2_X1 U736 ( .A1(n766), .A2(n767), .ZN(n763) );
  INV_X1 U737 ( .A(n768), .ZN(n767) );
  OR2_X1 U738 ( .A1(n769), .A2(n770), .ZN(Result_41_) );
  AND2_X1 U739 ( .A1(n771), .A2(Result_9_), .ZN(n770) );
  XOR2_X1 U740 ( .A(n772), .B(n773), .Z(n771) );
  AND2_X1 U741 ( .A1(n774), .A2(n558), .ZN(n769) );
  XNOR2_X1 U742 ( .A(n773), .B(n775), .ZN(n774) );
  OR2_X1 U743 ( .A1(n776), .A2(n777), .ZN(n773) );
  INV_X1 U744 ( .A(n778), .ZN(n777) );
  OR2_X1 U745 ( .A1(n779), .A2(n780), .ZN(Result_40_) );
  AND2_X1 U746 ( .A1(n781), .A2(Result_9_), .ZN(n780) );
  XOR2_X1 U747 ( .A(n782), .B(n783), .Z(n781) );
  AND2_X1 U748 ( .A1(n784), .A2(n558), .ZN(n779) );
  XNOR2_X1 U749 ( .A(n783), .B(n785), .ZN(n784) );
  OR2_X1 U750 ( .A1(n786), .A2(n787), .ZN(n783) );
  INV_X1 U751 ( .A(n788), .ZN(n787) );
  OR2_X1 U752 ( .A1(n789), .A2(n790), .ZN(Result_39_) );
  AND2_X1 U753 ( .A1(n791), .A2(Result_9_), .ZN(n790) );
  XOR2_X1 U754 ( .A(n792), .B(n793), .Z(n791) );
  AND2_X1 U755 ( .A1(n794), .A2(n558), .ZN(n789) );
  XNOR2_X1 U756 ( .A(n793), .B(n795), .ZN(n794) );
  OR2_X1 U757 ( .A1(n796), .A2(n797), .ZN(n793) );
  INV_X1 U758 ( .A(n798), .ZN(n797) );
  OR2_X1 U759 ( .A1(n799), .A2(n800), .ZN(Result_38_) );
  AND2_X1 U760 ( .A1(n801), .A2(Result_9_), .ZN(n800) );
  XOR2_X1 U761 ( .A(n802), .B(n803), .Z(n801) );
  AND2_X1 U762 ( .A1(n804), .A2(n558), .ZN(n799) );
  XNOR2_X1 U763 ( .A(n803), .B(n805), .ZN(n804) );
  OR2_X1 U764 ( .A1(n806), .A2(n807), .ZN(n803) );
  INV_X1 U765 ( .A(n808), .ZN(n807) );
  OR2_X1 U766 ( .A1(n809), .A2(n810), .ZN(Result_37_) );
  AND2_X1 U767 ( .A1(n811), .A2(Result_9_), .ZN(n810) );
  XOR2_X1 U768 ( .A(n812), .B(n813), .Z(n811) );
  AND2_X1 U769 ( .A1(n814), .A2(n558), .ZN(n809) );
  XNOR2_X1 U770 ( .A(n813), .B(n815), .ZN(n814) );
  OR2_X1 U771 ( .A1(n816), .A2(n817), .ZN(n813) );
  INV_X1 U772 ( .A(n818), .ZN(n817) );
  OR2_X1 U773 ( .A1(n819), .A2(n820), .ZN(Result_36_) );
  AND2_X1 U774 ( .A1(n821), .A2(Result_9_), .ZN(n820) );
  XOR2_X1 U775 ( .A(n822), .B(n823), .Z(n821) );
  AND2_X1 U776 ( .A1(n824), .A2(n558), .ZN(n819) );
  XNOR2_X1 U777 ( .A(n823), .B(n825), .ZN(n824) );
  OR2_X1 U778 ( .A1(n826), .A2(n827), .ZN(n823) );
  INV_X1 U779 ( .A(n828), .ZN(n827) );
  OR2_X1 U780 ( .A1(n829), .A2(n830), .ZN(Result_35_) );
  AND2_X1 U781 ( .A1(n831), .A2(Result_9_), .ZN(n830) );
  XOR2_X1 U782 ( .A(n832), .B(n833), .Z(n831) );
  AND2_X1 U783 ( .A1(n834), .A2(n558), .ZN(n829) );
  XNOR2_X1 U784 ( .A(n833), .B(n835), .ZN(n834) );
  OR2_X1 U785 ( .A1(n836), .A2(n837), .ZN(n833) );
  INV_X1 U786 ( .A(n838), .ZN(n837) );
  OR2_X1 U787 ( .A1(n839), .A2(n840), .ZN(Result_34_) );
  AND2_X1 U788 ( .A1(n841), .A2(Result_9_), .ZN(n840) );
  XOR2_X1 U789 ( .A(n842), .B(n843), .Z(n841) );
  AND2_X1 U790 ( .A1(n844), .A2(n558), .ZN(n839) );
  XNOR2_X1 U791 ( .A(n843), .B(n845), .ZN(n844) );
  OR2_X1 U792 ( .A1(n846), .A2(n847), .ZN(n843) );
  INV_X1 U793 ( .A(n848), .ZN(n847) );
  OR2_X1 U794 ( .A1(n849), .A2(n850), .ZN(Result_33_) );
  AND2_X1 U795 ( .A1(n851), .A2(Result_9_), .ZN(n850) );
  XOR2_X1 U796 ( .A(n852), .B(n853), .Z(n851) );
  AND2_X1 U797 ( .A1(n854), .A2(n558), .ZN(n849) );
  XOR2_X1 U798 ( .A(n853), .B(n855), .Z(n854) );
  OR2_X1 U799 ( .A1(n856), .A2(n857), .ZN(n853) );
  INV_X1 U800 ( .A(n858), .ZN(n857) );
  OR2_X1 U801 ( .A1(n859), .A2(n860), .ZN(Result_32_) );
  AND2_X1 U802 ( .A1(n861), .A2(Result_9_), .ZN(n860) );
  OR2_X1 U803 ( .A1(n862), .A2(n863), .ZN(n861) );
  INV_X1 U804 ( .A(n864), .ZN(n862) );
  OR2_X1 U805 ( .A1(n856), .A2(n865), .ZN(n864) );
  AND2_X1 U806 ( .A1(n852), .A2(n858), .ZN(n865) );
  OR2_X1 U807 ( .A1(n866), .A2(n846), .ZN(n852) );
  AND2_X1 U808 ( .A1(n842), .A2(n848), .ZN(n866) );
  OR2_X1 U809 ( .A1(n867), .A2(n836), .ZN(n842) );
  AND2_X1 U810 ( .A1(n832), .A2(n838), .ZN(n867) );
  OR2_X1 U811 ( .A1(n868), .A2(n826), .ZN(n832) );
  AND2_X1 U812 ( .A1(n822), .A2(n828), .ZN(n868) );
  OR2_X1 U813 ( .A1(n869), .A2(n816), .ZN(n822) );
  AND2_X1 U814 ( .A1(n812), .A2(n818), .ZN(n869) );
  OR2_X1 U815 ( .A1(n870), .A2(n806), .ZN(n812) );
  AND2_X1 U816 ( .A1(n802), .A2(n808), .ZN(n870) );
  OR2_X1 U817 ( .A1(n871), .A2(n796), .ZN(n802) );
  AND2_X1 U818 ( .A1(n792), .A2(n798), .ZN(n871) );
  OR2_X1 U819 ( .A1(n872), .A2(n786), .ZN(n792) );
  AND2_X1 U820 ( .A1(n782), .A2(n788), .ZN(n872) );
  OR2_X1 U821 ( .A1(n873), .A2(n776), .ZN(n782) );
  AND2_X1 U822 ( .A1(n772), .A2(n778), .ZN(n873) );
  OR2_X1 U823 ( .A1(n874), .A2(n766), .ZN(n772) );
  AND2_X1 U824 ( .A1(n762), .A2(n768), .ZN(n874) );
  OR2_X1 U825 ( .A1(n875), .A2(n756), .ZN(n762) );
  AND2_X1 U826 ( .A1(n752), .A2(n758), .ZN(n875) );
  OR2_X1 U827 ( .A1(n876), .A2(n746), .ZN(n752) );
  AND2_X1 U828 ( .A1(n742), .A2(n748), .ZN(n876) );
  OR2_X1 U829 ( .A1(n877), .A2(n736), .ZN(n742) );
  AND2_X1 U830 ( .A1(n732), .A2(n738), .ZN(n877) );
  OR2_X1 U831 ( .A1(n878), .A2(n726), .ZN(n732) );
  AND2_X1 U832 ( .A1(n722), .A2(n728), .ZN(n878) );
  OR2_X1 U833 ( .A1(n879), .A2(n716), .ZN(n722) );
  AND2_X1 U834 ( .A1(n712), .A2(n718), .ZN(n879) );
  OR2_X1 U835 ( .A1(n880), .A2(n706), .ZN(n712) );
  AND2_X1 U836 ( .A1(n702), .A2(n708), .ZN(n880) );
  OR2_X1 U837 ( .A1(n881), .A2(n696), .ZN(n702) );
  AND2_X1 U838 ( .A1(n692), .A2(n698), .ZN(n881) );
  OR2_X1 U839 ( .A1(n882), .A2(n686), .ZN(n692) );
  AND2_X1 U840 ( .A1(n682), .A2(n688), .ZN(n882) );
  OR2_X1 U841 ( .A1(n883), .A2(n676), .ZN(n682) );
  AND2_X1 U842 ( .A1(n672), .A2(n678), .ZN(n883) );
  OR2_X1 U843 ( .A1(n884), .A2(n666), .ZN(n672) );
  AND2_X1 U844 ( .A1(n662), .A2(n668), .ZN(n884) );
  OR2_X1 U845 ( .A1(n885), .A2(n656), .ZN(n662) );
  AND2_X1 U846 ( .A1(n652), .A2(n658), .ZN(n885) );
  OR2_X1 U847 ( .A1(n886), .A2(n646), .ZN(n652) );
  AND2_X1 U848 ( .A1(n642), .A2(n648), .ZN(n886) );
  OR2_X1 U849 ( .A1(n887), .A2(n636), .ZN(n642) );
  AND2_X1 U850 ( .A1(n632), .A2(n638), .ZN(n887) );
  OR2_X1 U851 ( .A1(n888), .A2(n626), .ZN(n632) );
  AND2_X1 U852 ( .A1(n622), .A2(n628), .ZN(n888) );
  OR2_X1 U853 ( .A1(n889), .A2(n616), .ZN(n622) );
  AND2_X1 U854 ( .A1(n612), .A2(n618), .ZN(n889) );
  OR2_X1 U855 ( .A1(n890), .A2(n606), .ZN(n612) );
  AND2_X1 U856 ( .A1(n602), .A2(n608), .ZN(n890) );
  OR2_X1 U857 ( .A1(n891), .A2(n596), .ZN(n602) );
  AND2_X1 U858 ( .A1(n592), .A2(n598), .ZN(n891) );
  OR2_X1 U859 ( .A1(n892), .A2(n586), .ZN(n592) );
  AND2_X1 U860 ( .A1(n582), .A2(n588), .ZN(n892) );
  AND2_X1 U861 ( .A1(n893), .A2(n558), .ZN(n859) );
  INV_X1 U862 ( .A(n894), .ZN(n558) );
  OR2_X1 U863 ( .A1(Result_9_), .A2(n895), .ZN(n894) );
  AND2_X1 U864 ( .A1(n896), .A2(n897), .ZN(n895) );
  AND4_X1 U865 ( .A1(n898), .A2(n899), .A3(n900), .A4(n901), .ZN(n897) );
  AND4_X1 U866 ( .A1(n808), .A2(n818), .A3(n828), .A4(n838), .ZN(n901) );
  AND4_X1 U867 ( .A1(n768), .A2(n778), .A3(n788), .A4(n798), .ZN(n900) );
  AND4_X1 U868 ( .A1(n728), .A2(n738), .A3(n748), .A4(n758), .ZN(n899) );
  AND4_X1 U869 ( .A1(n688), .A2(n698), .A3(n708), .A4(n718), .ZN(n898) );
  AND4_X1 U870 ( .A1(n902), .A2(n903), .A3(n904), .A4(n905), .ZN(n896) );
  AND4_X1 U871 ( .A1(n648), .A2(n658), .A3(n668), .A4(n678), .ZN(n905) );
  AND4_X1 U872 ( .A1(n608), .A2(n618), .A3(n628), .A4(n638), .ZN(n904) );
  AND4_X1 U873 ( .A1(n848), .A2(n578), .A3(n588), .A4(n598), .ZN(n903) );
  AND4_X1 U874 ( .A1(n906), .A2(n568), .A3(n907), .A4(n858), .ZN(n902) );
  INV_X1 U875 ( .A(n550), .ZN(n906) );
  AND2_X1 U876 ( .A1(n560), .A2(b_31_), .ZN(n550) );
  AND2_X1 U877 ( .A1(n910), .A2(n907), .ZN(n908) );
  OR2_X1 U878 ( .A1(n911), .A2(n856), .ZN(n910) );
  AND2_X1 U879 ( .A1(n912), .A2(a_1_), .ZN(n856) );
  AND2_X1 U880 ( .A1(n913), .A2(n858), .ZN(n911) );
  OR2_X1 U881 ( .A1(a_1_), .A2(n912), .ZN(n858) );
  INV_X1 U882 ( .A(b_1_), .ZN(n912) );
  OR2_X1 U883 ( .A1(n914), .A2(n846), .ZN(n913) );
  AND2_X1 U884 ( .A1(n915), .A2(a_2_), .ZN(n846) );
  AND2_X1 U885 ( .A1(n916), .A2(n848), .ZN(n914) );
  OR2_X1 U886 ( .A1(a_2_), .A2(n915), .ZN(n848) );
  OR2_X1 U887 ( .A1(n917), .A2(n836), .ZN(n916) );
  AND2_X1 U888 ( .A1(n918), .A2(a_3_), .ZN(n836) );
  AND3_X1 U889 ( .A1(n828), .A2(n838), .A3(n919), .ZN(n917) );
  OR3_X1 U890 ( .A1(n816), .A2(n826), .A3(n920), .ZN(n919) );
  AND3_X1 U891 ( .A1(n808), .A2(n818), .A3(n921), .ZN(n920) );
  OR3_X1 U892 ( .A1(n796), .A2(n806), .A3(n922), .ZN(n921) );
  AND3_X1 U893 ( .A1(n788), .A2(n798), .A3(n923), .ZN(n922) );
  OR3_X1 U894 ( .A1(n776), .A2(n786), .A3(n924), .ZN(n923) );
  AND3_X1 U895 ( .A1(n768), .A2(n778), .A3(n925), .ZN(n924) );
  OR3_X1 U896 ( .A1(n756), .A2(n766), .A3(n926), .ZN(n925) );
  AND3_X1 U897 ( .A1(n748), .A2(n758), .A3(n927), .ZN(n926) );
  OR3_X1 U898 ( .A1(n736), .A2(n746), .A3(n928), .ZN(n927) );
  AND3_X1 U899 ( .A1(n728), .A2(n738), .A3(n929), .ZN(n928) );
  OR3_X1 U900 ( .A1(n716), .A2(n726), .A3(n930), .ZN(n929) );
  AND3_X1 U901 ( .A1(n708), .A2(n718), .A3(n931), .ZN(n930) );
  OR3_X1 U902 ( .A1(n696), .A2(n706), .A3(n932), .ZN(n931) );
  AND3_X1 U903 ( .A1(n688), .A2(n698), .A3(n933), .ZN(n932) );
  OR3_X1 U904 ( .A1(n676), .A2(n686), .A3(n934), .ZN(n933) );
  AND3_X1 U905 ( .A1(n668), .A2(n678), .A3(n935), .ZN(n934) );
  OR3_X1 U906 ( .A1(n656), .A2(n666), .A3(n936), .ZN(n935) );
  AND3_X1 U907 ( .A1(n648), .A2(n658), .A3(n937), .ZN(n936) );
  OR3_X1 U908 ( .A1(n636), .A2(n646), .A3(n938), .ZN(n937) );
  AND3_X1 U909 ( .A1(n628), .A2(n638), .A3(n939), .ZN(n938) );
  OR3_X1 U910 ( .A1(n616), .A2(n626), .A3(n940), .ZN(n939) );
  AND3_X1 U911 ( .A1(n608), .A2(n618), .A3(n941), .ZN(n940) );
  OR3_X1 U912 ( .A1(n596), .A2(n606), .A3(n942), .ZN(n941) );
  AND3_X1 U913 ( .A1(n588), .A2(n598), .A3(n943), .ZN(n942) );
  OR2_X1 U914 ( .A1(n586), .A2(n582), .ZN(n943) );
  OR2_X1 U915 ( .A1(n944), .A2(n576), .ZN(n582) );
  AND2_X1 U916 ( .A1(a_29_), .A2(n945), .ZN(n576) );
  AND2_X1 U917 ( .A1(n572), .A2(n578), .ZN(n944) );
  OR2_X1 U918 ( .A1(a_29_), .A2(n945), .ZN(n578) );
  OR2_X1 U919 ( .A1(n946), .A2(n566), .ZN(n572) );
  AND2_X1 U920 ( .A1(n947), .A2(a_30_), .ZN(n566) );
  AND2_X1 U921 ( .A1(n549), .A2(n568), .ZN(n946) );
  OR2_X1 U922 ( .A1(a_30_), .A2(n947), .ZN(n568) );
  INV_X1 U923 ( .A(b_30_), .ZN(n947) );
  INV_X1 U924 ( .A(n557), .ZN(n549) );
  OR2_X1 U925 ( .A1(b_31_), .A2(n560), .ZN(n557) );
  INV_X1 U926 ( .A(a_31_), .ZN(n560) );
  AND2_X1 U927 ( .A1(n948), .A2(a_28_), .ZN(n586) );
  OR2_X1 U928 ( .A1(a_27_), .A2(n949), .ZN(n598) );
  OR2_X1 U929 ( .A1(a_28_), .A2(n948), .ZN(n588) );
  AND2_X1 U930 ( .A1(n950), .A2(a_26_), .ZN(n606) );
  AND2_X1 U931 ( .A1(n949), .A2(a_27_), .ZN(n596) );
  OR2_X1 U932 ( .A1(a_25_), .A2(n951), .ZN(n618) );
  OR2_X1 U933 ( .A1(a_26_), .A2(n950), .ZN(n608) );
  AND2_X1 U934 ( .A1(n952), .A2(a_24_), .ZN(n626) );
  AND2_X1 U935 ( .A1(n951), .A2(a_25_), .ZN(n616) );
  OR2_X1 U936 ( .A1(a_23_), .A2(n953), .ZN(n638) );
  OR2_X1 U937 ( .A1(a_24_), .A2(n952), .ZN(n628) );
  AND2_X1 U938 ( .A1(n954), .A2(a_22_), .ZN(n646) );
  AND2_X1 U939 ( .A1(n953), .A2(a_23_), .ZN(n636) );
  OR2_X1 U940 ( .A1(a_21_), .A2(n955), .ZN(n658) );
  OR2_X1 U941 ( .A1(a_22_), .A2(n954), .ZN(n648) );
  AND2_X1 U942 ( .A1(n956), .A2(a_20_), .ZN(n666) );
  AND2_X1 U943 ( .A1(n955), .A2(a_21_), .ZN(n656) );
  OR2_X1 U944 ( .A1(a_19_), .A2(n957), .ZN(n678) );
  OR2_X1 U945 ( .A1(a_20_), .A2(n956), .ZN(n668) );
  AND2_X1 U946 ( .A1(n958), .A2(a_18_), .ZN(n686) );
  AND2_X1 U947 ( .A1(n957), .A2(a_19_), .ZN(n676) );
  OR2_X1 U948 ( .A1(a_17_), .A2(n959), .ZN(n698) );
  OR2_X1 U949 ( .A1(a_18_), .A2(n958), .ZN(n688) );
  AND2_X1 U950 ( .A1(n960), .A2(a_16_), .ZN(n706) );
  AND2_X1 U951 ( .A1(n959), .A2(a_17_), .ZN(n696) );
  OR2_X1 U952 ( .A1(a_15_), .A2(n961), .ZN(n718) );
  OR2_X1 U953 ( .A1(a_16_), .A2(n960), .ZN(n708) );
  AND2_X1 U954 ( .A1(n962), .A2(a_14_), .ZN(n726) );
  AND2_X1 U955 ( .A1(n961), .A2(a_15_), .ZN(n716) );
  OR2_X1 U956 ( .A1(a_13_), .A2(n963), .ZN(n738) );
  OR2_X1 U957 ( .A1(a_14_), .A2(n962), .ZN(n728) );
  AND2_X1 U958 ( .A1(n964), .A2(a_12_), .ZN(n746) );
  AND2_X1 U959 ( .A1(n963), .A2(a_13_), .ZN(n736) );
  OR2_X1 U960 ( .A1(a_11_), .A2(n965), .ZN(n758) );
  OR2_X1 U961 ( .A1(a_12_), .A2(n964), .ZN(n748) );
  AND2_X1 U962 ( .A1(n966), .A2(a_10_), .ZN(n766) );
  AND2_X1 U963 ( .A1(n965), .A2(a_11_), .ZN(n756) );
  OR2_X1 U964 ( .A1(a_9_), .A2(n967), .ZN(n778) );
  OR2_X1 U965 ( .A1(a_10_), .A2(n966), .ZN(n768) );
  AND2_X1 U966 ( .A1(n968), .A2(a_8_), .ZN(n786) );
  AND2_X1 U967 ( .A1(n967), .A2(a_9_), .ZN(n776) );
  OR2_X1 U968 ( .A1(a_7_), .A2(n969), .ZN(n798) );
  OR2_X1 U969 ( .A1(a_8_), .A2(n968), .ZN(n788) );
  AND2_X1 U970 ( .A1(n970), .A2(a_6_), .ZN(n806) );
  AND2_X1 U971 ( .A1(n969), .A2(a_7_), .ZN(n796) );
  OR2_X1 U972 ( .A1(a_5_), .A2(n971), .ZN(n818) );
  OR2_X1 U973 ( .A1(a_6_), .A2(n970), .ZN(n808) );
  AND2_X1 U974 ( .A1(n972), .A2(a_4_), .ZN(n826) );
  AND2_X1 U975 ( .A1(n971), .A2(a_5_), .ZN(n816) );
  OR2_X1 U976 ( .A1(a_3_), .A2(n918), .ZN(n838) );
  OR2_X1 U977 ( .A1(a_4_), .A2(n972), .ZN(n828) );
  XNOR2_X1 U978 ( .A(n863), .B(n973), .ZN(n893) );
  AND2_X1 U979 ( .A1(n974), .A2(n975), .ZN(n973) );
  OR2_X1 U980 ( .A1(b_1_), .A2(n976), .ZN(n975) );
  AND2_X1 U981 ( .A1(n855), .A2(a_1_), .ZN(n976) );
  OR2_X1 U982 ( .A1(a_1_), .A2(n855), .ZN(n974) );
  INV_X1 U983 ( .A(n977), .ZN(n855) );
  OR2_X1 U984 ( .A1(n978), .A2(n979), .ZN(n977) );
  AND2_X1 U985 ( .A1(n845), .A2(n980), .ZN(n979) );
  AND2_X1 U986 ( .A1(n981), .A2(n915), .ZN(n978) );
  INV_X1 U987 ( .A(b_2_), .ZN(n915) );
  OR2_X1 U988 ( .A1(n980), .A2(n845), .ZN(n981) );
  OR2_X1 U989 ( .A1(n982), .A2(n983), .ZN(n845) );
  AND2_X1 U990 ( .A1(n835), .A2(n984), .ZN(n983) );
  AND2_X1 U991 ( .A1(n985), .A2(n918), .ZN(n982) );
  INV_X1 U992 ( .A(b_3_), .ZN(n918) );
  OR2_X1 U993 ( .A1(n984), .A2(n835), .ZN(n985) );
  OR2_X1 U994 ( .A1(n986), .A2(n987), .ZN(n835) );
  AND2_X1 U995 ( .A1(n825), .A2(n988), .ZN(n987) );
  AND2_X1 U996 ( .A1(n989), .A2(n972), .ZN(n986) );
  INV_X1 U997 ( .A(b_4_), .ZN(n972) );
  OR2_X1 U998 ( .A1(n988), .A2(n825), .ZN(n989) );
  OR2_X1 U999 ( .A1(n990), .A2(n991), .ZN(n825) );
  AND2_X1 U1000 ( .A1(n815), .A2(n992), .ZN(n991) );
  AND2_X1 U1001 ( .A1(n993), .A2(n971), .ZN(n990) );
  INV_X1 U1002 ( .A(b_5_), .ZN(n971) );
  OR2_X1 U1003 ( .A1(n992), .A2(n815), .ZN(n993) );
  OR2_X1 U1004 ( .A1(n994), .A2(n995), .ZN(n815) );
  AND2_X1 U1005 ( .A1(n805), .A2(n996), .ZN(n995) );
  AND2_X1 U1006 ( .A1(n997), .A2(n970), .ZN(n994) );
  INV_X1 U1007 ( .A(b_6_), .ZN(n970) );
  OR2_X1 U1008 ( .A1(n996), .A2(n805), .ZN(n997) );
  OR2_X1 U1009 ( .A1(n998), .A2(n999), .ZN(n805) );
  AND2_X1 U1010 ( .A1(n795), .A2(n1000), .ZN(n999) );
  AND2_X1 U1011 ( .A1(n1001), .A2(n969), .ZN(n998) );
  INV_X1 U1012 ( .A(b_7_), .ZN(n969) );
  OR2_X1 U1013 ( .A1(n1000), .A2(n795), .ZN(n1001) );
  OR2_X1 U1014 ( .A1(n1002), .A2(n1003), .ZN(n795) );
  AND2_X1 U1015 ( .A1(n785), .A2(n1004), .ZN(n1003) );
  AND2_X1 U1016 ( .A1(n1005), .A2(n968), .ZN(n1002) );
  INV_X1 U1017 ( .A(b_8_), .ZN(n968) );
  OR2_X1 U1018 ( .A1(n1004), .A2(n785), .ZN(n1005) );
  OR2_X1 U1019 ( .A1(n1006), .A2(n1007), .ZN(n785) );
  AND2_X1 U1020 ( .A1(n775), .A2(n1008), .ZN(n1007) );
  AND2_X1 U1021 ( .A1(n1009), .A2(n967), .ZN(n1006) );
  INV_X1 U1022 ( .A(b_9_), .ZN(n967) );
  OR2_X1 U1023 ( .A1(n1008), .A2(n775), .ZN(n1009) );
  OR2_X1 U1024 ( .A1(n1010), .A2(n1011), .ZN(n775) );
  AND2_X1 U1025 ( .A1(n765), .A2(n1012), .ZN(n1011) );
  AND2_X1 U1026 ( .A1(n1013), .A2(n966), .ZN(n1010) );
  INV_X1 U1027 ( .A(b_10_), .ZN(n966) );
  OR2_X1 U1028 ( .A1(n1012), .A2(n765), .ZN(n1013) );
  OR2_X1 U1029 ( .A1(n1014), .A2(n1015), .ZN(n765) );
  AND2_X1 U1030 ( .A1(n755), .A2(n1016), .ZN(n1015) );
  AND2_X1 U1031 ( .A1(n1017), .A2(n965), .ZN(n1014) );
  INV_X1 U1032 ( .A(b_11_), .ZN(n965) );
  OR2_X1 U1033 ( .A1(n1016), .A2(n755), .ZN(n1017) );
  OR2_X1 U1034 ( .A1(n1018), .A2(n1019), .ZN(n755) );
  AND2_X1 U1035 ( .A1(n745), .A2(n1020), .ZN(n1019) );
  AND2_X1 U1036 ( .A1(n1021), .A2(n964), .ZN(n1018) );
  INV_X1 U1037 ( .A(b_12_), .ZN(n964) );
  OR2_X1 U1038 ( .A1(n1020), .A2(n745), .ZN(n1021) );
  OR2_X1 U1039 ( .A1(n1022), .A2(n1023), .ZN(n745) );
  AND2_X1 U1040 ( .A1(n735), .A2(n1024), .ZN(n1023) );
  AND2_X1 U1041 ( .A1(n1025), .A2(n963), .ZN(n1022) );
  INV_X1 U1042 ( .A(b_13_), .ZN(n963) );
  OR2_X1 U1043 ( .A1(n1024), .A2(n735), .ZN(n1025) );
  OR2_X1 U1044 ( .A1(n1026), .A2(n1027), .ZN(n735) );
  AND2_X1 U1045 ( .A1(n725), .A2(n1028), .ZN(n1027) );
  AND2_X1 U1046 ( .A1(n1029), .A2(n962), .ZN(n1026) );
  INV_X1 U1047 ( .A(b_14_), .ZN(n962) );
  OR2_X1 U1048 ( .A1(n1028), .A2(n725), .ZN(n1029) );
  OR2_X1 U1049 ( .A1(n1030), .A2(n1031), .ZN(n725) );
  AND2_X1 U1050 ( .A1(n715), .A2(n1032), .ZN(n1031) );
  AND2_X1 U1051 ( .A1(n1033), .A2(n961), .ZN(n1030) );
  INV_X1 U1052 ( .A(b_15_), .ZN(n961) );
  OR2_X1 U1053 ( .A1(n1032), .A2(n715), .ZN(n1033) );
  OR2_X1 U1054 ( .A1(n1034), .A2(n1035), .ZN(n715) );
  AND2_X1 U1055 ( .A1(n705), .A2(n1036), .ZN(n1035) );
  AND2_X1 U1056 ( .A1(n1037), .A2(n960), .ZN(n1034) );
  INV_X1 U1057 ( .A(b_16_), .ZN(n960) );
  OR2_X1 U1058 ( .A1(n1036), .A2(n705), .ZN(n1037) );
  OR2_X1 U1059 ( .A1(n1038), .A2(n1039), .ZN(n705) );
  AND2_X1 U1060 ( .A1(n695), .A2(n1040), .ZN(n1039) );
  AND2_X1 U1061 ( .A1(n1041), .A2(n959), .ZN(n1038) );
  INV_X1 U1062 ( .A(b_17_), .ZN(n959) );
  OR2_X1 U1063 ( .A1(n1040), .A2(n695), .ZN(n1041) );
  OR2_X1 U1064 ( .A1(n1042), .A2(n1043), .ZN(n695) );
  AND2_X1 U1065 ( .A1(n685), .A2(n1044), .ZN(n1043) );
  AND2_X1 U1066 ( .A1(n1045), .A2(n958), .ZN(n1042) );
  INV_X1 U1067 ( .A(b_18_), .ZN(n958) );
  OR2_X1 U1068 ( .A1(n1044), .A2(n685), .ZN(n1045) );
  OR2_X1 U1069 ( .A1(n1046), .A2(n1047), .ZN(n685) );
  AND2_X1 U1070 ( .A1(n675), .A2(n1048), .ZN(n1047) );
  AND2_X1 U1071 ( .A1(n1049), .A2(n957), .ZN(n1046) );
  INV_X1 U1072 ( .A(b_19_), .ZN(n957) );
  OR2_X1 U1073 ( .A1(n1048), .A2(n675), .ZN(n1049) );
  OR2_X1 U1074 ( .A1(n1050), .A2(n1051), .ZN(n675) );
  AND2_X1 U1075 ( .A1(n665), .A2(n1052), .ZN(n1051) );
  AND2_X1 U1076 ( .A1(n1053), .A2(n956), .ZN(n1050) );
  INV_X1 U1077 ( .A(b_20_), .ZN(n956) );
  OR2_X1 U1078 ( .A1(n1052), .A2(n665), .ZN(n1053) );
  OR2_X1 U1079 ( .A1(n1054), .A2(n1055), .ZN(n665) );
  AND2_X1 U1080 ( .A1(n655), .A2(n1056), .ZN(n1055) );
  AND2_X1 U1081 ( .A1(n1057), .A2(n955), .ZN(n1054) );
  INV_X1 U1082 ( .A(b_21_), .ZN(n955) );
  OR2_X1 U1083 ( .A1(n1056), .A2(n655), .ZN(n1057) );
  OR2_X1 U1084 ( .A1(n1058), .A2(n1059), .ZN(n655) );
  AND2_X1 U1085 ( .A1(n645), .A2(n1060), .ZN(n1059) );
  AND2_X1 U1086 ( .A1(n1061), .A2(n954), .ZN(n1058) );
  INV_X1 U1087 ( .A(b_22_), .ZN(n954) );
  OR2_X1 U1088 ( .A1(n1060), .A2(n645), .ZN(n1061) );
  OR2_X1 U1089 ( .A1(n1062), .A2(n1063), .ZN(n645) );
  AND2_X1 U1090 ( .A1(n635), .A2(n1064), .ZN(n1063) );
  AND2_X1 U1091 ( .A1(n1065), .A2(n953), .ZN(n1062) );
  INV_X1 U1092 ( .A(b_23_), .ZN(n953) );
  OR2_X1 U1093 ( .A1(n1064), .A2(n635), .ZN(n1065) );
  OR2_X1 U1094 ( .A1(n1066), .A2(n1067), .ZN(n635) );
  AND2_X1 U1095 ( .A1(n625), .A2(n1068), .ZN(n1067) );
  AND2_X1 U1096 ( .A1(n1069), .A2(n952), .ZN(n1066) );
  INV_X1 U1097 ( .A(b_24_), .ZN(n952) );
  OR2_X1 U1098 ( .A1(n1068), .A2(n625), .ZN(n1069) );
  OR2_X1 U1099 ( .A1(n1070), .A2(n1071), .ZN(n625) );
  AND2_X1 U1100 ( .A1(n615), .A2(n1072), .ZN(n1071) );
  AND2_X1 U1101 ( .A1(n1073), .A2(n951), .ZN(n1070) );
  INV_X1 U1102 ( .A(b_25_), .ZN(n951) );
  OR2_X1 U1103 ( .A1(n1072), .A2(n615), .ZN(n1073) );
  OR2_X1 U1104 ( .A1(n1074), .A2(n1075), .ZN(n615) );
  AND2_X1 U1105 ( .A1(n605), .A2(n1076), .ZN(n1075) );
  AND2_X1 U1106 ( .A1(n1077), .A2(n950), .ZN(n1074) );
  INV_X1 U1107 ( .A(b_26_), .ZN(n950) );
  OR2_X1 U1108 ( .A1(n1076), .A2(n605), .ZN(n1077) );
  OR2_X1 U1109 ( .A1(n1078), .A2(n1079), .ZN(n605) );
  AND2_X1 U1110 ( .A1(n595), .A2(n1080), .ZN(n1079) );
  AND2_X1 U1111 ( .A1(n1081), .A2(n949), .ZN(n1078) );
  INV_X1 U1112 ( .A(b_27_), .ZN(n949) );
  OR2_X1 U1113 ( .A1(n1080), .A2(n595), .ZN(n1081) );
  OR2_X1 U1114 ( .A1(n1082), .A2(n1083), .ZN(n595) );
  AND2_X1 U1115 ( .A1(n585), .A2(n1084), .ZN(n1083) );
  AND2_X1 U1116 ( .A1(n1085), .A2(n948), .ZN(n1082) );
  INV_X1 U1117 ( .A(b_28_), .ZN(n948) );
  OR2_X1 U1118 ( .A1(n1084), .A2(n585), .ZN(n1085) );
  OR2_X1 U1119 ( .A1(n1086), .A2(n1087), .ZN(n585) );
  AND2_X1 U1120 ( .A1(n1088), .A2(n1089), .ZN(n1087) );
  AND2_X1 U1121 ( .A1(n1090), .A2(n945), .ZN(n1086) );
  INV_X1 U1122 ( .A(b_29_), .ZN(n945) );
  OR2_X1 U1123 ( .A1(n1088), .A2(n1089), .ZN(n1090) );
  INV_X1 U1124 ( .A(a_29_), .ZN(n1089) );
  INV_X1 U1125 ( .A(n575), .ZN(n1088) );
  OR2_X1 U1126 ( .A1(n1091), .A2(n1092), .ZN(n575) );
  AND2_X1 U1127 ( .A1(a_30_), .A2(b_30_), .ZN(n1092) );
  AND3_X1 U1128 ( .A1(a_31_), .A2(n1093), .A3(b_31_), .ZN(n1091) );
  OR2_X1 U1129 ( .A1(a_30_), .A2(b_30_), .ZN(n1093) );
  INV_X1 U1130 ( .A(a_28_), .ZN(n1084) );
  INV_X1 U1131 ( .A(a_27_), .ZN(n1080) );
  INV_X1 U1132 ( .A(a_26_), .ZN(n1076) );
  INV_X1 U1133 ( .A(a_25_), .ZN(n1072) );
  INV_X1 U1134 ( .A(a_24_), .ZN(n1068) );
  INV_X1 U1135 ( .A(a_23_), .ZN(n1064) );
  INV_X1 U1136 ( .A(a_22_), .ZN(n1060) );
  INV_X1 U1137 ( .A(a_21_), .ZN(n1056) );
  INV_X1 U1138 ( .A(a_20_), .ZN(n1052) );
  INV_X1 U1139 ( .A(a_19_), .ZN(n1048) );
  INV_X1 U1140 ( .A(a_18_), .ZN(n1044) );
  INV_X1 U1141 ( .A(a_17_), .ZN(n1040) );
  INV_X1 U1142 ( .A(a_16_), .ZN(n1036) );
  INV_X1 U1143 ( .A(a_15_), .ZN(n1032) );
  INV_X1 U1144 ( .A(a_14_), .ZN(n1028) );
  INV_X1 U1145 ( .A(a_13_), .ZN(n1024) );
  INV_X1 U1146 ( .A(a_12_), .ZN(n1020) );
  INV_X1 U1147 ( .A(a_11_), .ZN(n1016) );
  INV_X1 U1148 ( .A(a_10_), .ZN(n1012) );
  INV_X1 U1149 ( .A(a_9_), .ZN(n1008) );
  INV_X1 U1150 ( .A(a_8_), .ZN(n1004) );
  INV_X1 U1151 ( .A(a_7_), .ZN(n1000) );
  INV_X1 U1152 ( .A(a_6_), .ZN(n996) );
  INV_X1 U1153 ( .A(a_5_), .ZN(n992) );
  INV_X1 U1154 ( .A(a_4_), .ZN(n988) );
  INV_X1 U1155 ( .A(a_3_), .ZN(n984) );
  INV_X1 U1156 ( .A(a_2_), .ZN(n980) );
  AND2_X1 U1157 ( .A1(n907), .A2(n1094), .ZN(n863) );
  INV_X1 U1158 ( .A(n909), .ZN(n1094) );
  AND2_X1 U1159 ( .A1(a_0_), .A2(n1095), .ZN(n909) );
  OR2_X1 U1160 ( .A1(a_0_), .A2(n1095), .ZN(n907) );
  INV_X1 U1161 ( .A(b_0_), .ZN(n1095) );
endmodule

