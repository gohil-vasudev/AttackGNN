module add_mul_16_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, 
        a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, 
        b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, 
        b_15_, operation, Result_0_, Result_1_, Result_2_, Result_3_, 
        Result_4_, Result_5_, Result_6_, Result_7_, Result_8_, Result_9_, 
        Result_10_, Result_11_, Result_12_, Result_13_, Result_14_, Result_15_, 
        Result_16_, Result_17_, Result_18_, Result_19_, Result_20_, Result_21_, 
        Result_22_, Result_23_, Result_24_, Result_25_, Result_26_, Result_27_, 
        Result_28_, Result_29_, Result_30_, Result_31_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_,
         b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_,
         operation;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_;
  wire   n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842;

  AND2_X1 U1946 ( .A1(n1914), .A2(operation), .ZN(Result_9_) );
  XOR2_X1 U1947 ( .A(n1915), .B(n1916), .Z(n1914) );
  AND2_X1 U1948 ( .A1(n1917), .A2(n1918), .ZN(n1916) );
  OR2_X1 U1949 ( .A1(n1919), .A2(n1920), .ZN(n1918) );
  AND2_X1 U1950 ( .A1(n1921), .A2(n1922), .ZN(n1920) );
  INV_X1 U1951 ( .A(n1923), .ZN(n1917) );
  AND2_X1 U1952 ( .A1(n1924), .A2(operation), .ZN(Result_8_) );
  XOR2_X1 U1953 ( .A(n1925), .B(n1926), .Z(n1924) );
  AND2_X1 U1954 ( .A1(operation), .A2(n1927), .ZN(Result_7_) );
  XOR2_X1 U1955 ( .A(n1928), .B(n1929), .Z(n1927) );
  AND2_X1 U1956 ( .A1(n1930), .A2(n1931), .ZN(n1929) );
  OR2_X1 U1957 ( .A1(n1932), .A2(n1933), .ZN(n1931) );
  AND2_X1 U1958 ( .A1(n1934), .A2(n1935), .ZN(n1933) );
  INV_X1 U1959 ( .A(n1936), .ZN(n1930) );
  AND2_X1 U1960 ( .A1(n1937), .A2(operation), .ZN(Result_6_) );
  XOR2_X1 U1961 ( .A(n1938), .B(n1939), .Z(n1937) );
  AND2_X1 U1962 ( .A1(operation), .A2(n1940), .ZN(Result_5_) );
  XOR2_X1 U1963 ( .A(n1941), .B(n1942), .Z(n1940) );
  AND2_X1 U1964 ( .A1(n1943), .A2(n1944), .ZN(n1942) );
  OR2_X1 U1965 ( .A1(n1945), .A2(n1946), .ZN(n1944) );
  AND2_X1 U1966 ( .A1(n1947), .A2(n1948), .ZN(n1946) );
  INV_X1 U1967 ( .A(n1949), .ZN(n1943) );
  AND2_X1 U1968 ( .A1(n1950), .A2(operation), .ZN(Result_4_) );
  XOR2_X1 U1969 ( .A(n1951), .B(n1952), .Z(n1950) );
  AND2_X1 U1970 ( .A1(operation), .A2(n1953), .ZN(Result_3_) );
  XOR2_X1 U1971 ( .A(n1954), .B(n1955), .Z(n1953) );
  AND2_X1 U1972 ( .A1(n1956), .A2(n1957), .ZN(n1955) );
  OR2_X1 U1973 ( .A1(n1958), .A2(n1959), .ZN(n1957) );
  AND2_X1 U1974 ( .A1(n1960), .A2(n1961), .ZN(n1959) );
  INV_X1 U1975 ( .A(n1962), .ZN(n1956) );
  OR2_X1 U1976 ( .A1(n1963), .A2(n1964), .ZN(Result_31_) );
  AND2_X1 U1977 ( .A1(n1965), .A2(operation), .ZN(n1964) );
  INV_X1 U1978 ( .A(n1966), .ZN(n1965) );
  AND2_X1 U1979 ( .A1(n1967), .A2(n1968), .ZN(n1963) );
  XNOR2_X1 U1980 ( .A(n1969), .B(a_15_), .ZN(n1967) );
  OR2_X1 U1981 ( .A1(n1970), .A2(n1971), .ZN(Result_30_) );
  AND2_X1 U1982 ( .A1(n1972), .A2(n1968), .ZN(n1971) );
  XNOR2_X1 U1983 ( .A(n1966), .B(n1973), .ZN(n1972) );
  XNOR2_X1 U1984 ( .A(n1974), .B(a_14_), .ZN(n1973) );
  AND2_X1 U1985 ( .A1(operation), .A2(n1975), .ZN(n1970) );
  OR2_X1 U1986 ( .A1(n1976), .A2(n1977), .ZN(n1975) );
  AND2_X1 U1987 ( .A1(b_15_), .A2(n1978), .ZN(n1977) );
  OR2_X1 U1988 ( .A1(n1979), .A2(n1980), .ZN(n1978) );
  AND2_X1 U1989 ( .A1(a_14_), .A2(n1974), .ZN(n1979) );
  AND2_X1 U1990 ( .A1(b_14_), .A2(n1981), .ZN(n1976) );
  OR2_X1 U1991 ( .A1(n1982), .A2(n1983), .ZN(n1981) );
  AND2_X1 U1992 ( .A1(a_15_), .A2(n1969), .ZN(n1982) );
  AND2_X1 U1993 ( .A1(n1984), .A2(operation), .ZN(Result_2_) );
  XOR2_X1 U1994 ( .A(n1985), .B(n1986), .Z(n1984) );
  OR2_X1 U1995 ( .A1(n1987), .A2(n1988), .ZN(Result_29_) );
  AND2_X1 U1996 ( .A1(n1989), .A2(operation), .ZN(n1988) );
  XOR2_X1 U1997 ( .A(n1990), .B(n1991), .Z(n1989) );
  XNOR2_X1 U1998 ( .A(n1992), .B(n1993), .ZN(n1991) );
  AND2_X1 U1999 ( .A1(n1994), .A2(n1968), .ZN(n1987) );
  OR3_X1 U2000 ( .A1(n1995), .A2(n1996), .A3(n1997), .ZN(n1994) );
  INV_X1 U2001 ( .A(n1998), .ZN(n1997) );
  OR2_X1 U2002 ( .A1(n1999), .A2(n2000), .ZN(n1998) );
  AND2_X1 U2003 ( .A1(n2001), .A2(n2002), .ZN(n1996) );
  XNOR2_X1 U2004 ( .A(n2000), .B(a_13_), .ZN(n2001) );
  AND3_X1 U2005 ( .A1(n2000), .A2(n2003), .A3(b_13_), .ZN(n1995) );
  OR2_X1 U2006 ( .A1(n2004), .A2(n2005), .ZN(Result_28_) );
  AND2_X1 U2007 ( .A1(n2006), .A2(operation), .ZN(n2005) );
  XNOR2_X1 U2008 ( .A(n2007), .B(n2008), .ZN(n2006) );
  XOR2_X1 U2009 ( .A(n2009), .B(n2010), .Z(n2008) );
  AND2_X1 U2010 ( .A1(n2011), .A2(n1968), .ZN(n2004) );
  XOR2_X1 U2011 ( .A(n2012), .B(n2013), .Z(n2011) );
  OR2_X1 U2012 ( .A1(n2014), .A2(n2015), .ZN(n2013) );
  OR2_X1 U2013 ( .A1(n2016), .A2(n2017), .ZN(Result_27_) );
  AND2_X1 U2014 ( .A1(n2018), .A2(operation), .ZN(n2017) );
  XNOR2_X1 U2015 ( .A(n2019), .B(n2020), .ZN(n2018) );
  XOR2_X1 U2016 ( .A(n2021), .B(n2022), .Z(n2020) );
  AND2_X1 U2017 ( .A1(n2023), .A2(n1968), .ZN(n2016) );
  OR3_X1 U2018 ( .A1(n2024), .A2(n2025), .A3(n2026), .ZN(n2023) );
  INV_X1 U2019 ( .A(n2027), .ZN(n2026) );
  OR2_X1 U2020 ( .A1(n2028), .A2(n2029), .ZN(n2027) );
  AND2_X1 U2021 ( .A1(n2030), .A2(n2031), .ZN(n2025) );
  XNOR2_X1 U2022 ( .A(a_11_), .B(n2028), .ZN(n2030) );
  AND3_X1 U2023 ( .A1(n2028), .A2(n2032), .A3(b_11_), .ZN(n2024) );
  OR2_X1 U2024 ( .A1(n2033), .A2(n2034), .ZN(Result_26_) );
  AND2_X1 U2025 ( .A1(n2035), .A2(operation), .ZN(n2034) );
  XNOR2_X1 U2026 ( .A(n2036), .B(n2037), .ZN(n2035) );
  XOR2_X1 U2027 ( .A(n2038), .B(n2039), .Z(n2037) );
  AND2_X1 U2028 ( .A1(n2040), .A2(n1968), .ZN(n2033) );
  XOR2_X1 U2029 ( .A(n2041), .B(n2042), .Z(n2040) );
  OR2_X1 U2030 ( .A1(n2043), .A2(n2044), .ZN(n2042) );
  OR2_X1 U2031 ( .A1(n2045), .A2(n2046), .ZN(Result_25_) );
  AND2_X1 U2032 ( .A1(n2047), .A2(operation), .ZN(n2046) );
  XNOR2_X1 U2033 ( .A(n2048), .B(n2049), .ZN(n2047) );
  XOR2_X1 U2034 ( .A(n2050), .B(n2051), .Z(n2049) );
  AND2_X1 U2035 ( .A1(n2052), .A2(n1968), .ZN(n2045) );
  OR3_X1 U2036 ( .A1(n2053), .A2(n2054), .A3(n2055), .ZN(n2052) );
  INV_X1 U2037 ( .A(n2056), .ZN(n2055) );
  OR2_X1 U2038 ( .A1(n2057), .A2(n2058), .ZN(n2056) );
  AND2_X1 U2039 ( .A1(n2059), .A2(n2060), .ZN(n2054) );
  XNOR2_X1 U2040 ( .A(a_9_), .B(n2057), .ZN(n2059) );
  AND3_X1 U2041 ( .A1(n2057), .A2(n2061), .A3(b_9_), .ZN(n2053) );
  OR2_X1 U2042 ( .A1(n2062), .A2(n2063), .ZN(Result_24_) );
  AND2_X1 U2043 ( .A1(n2064), .A2(operation), .ZN(n2063) );
  XNOR2_X1 U2044 ( .A(n2065), .B(n2066), .ZN(n2064) );
  XOR2_X1 U2045 ( .A(n2067), .B(n2068), .Z(n2066) );
  AND2_X1 U2046 ( .A1(n2069), .A2(n1968), .ZN(n2062) );
  XOR2_X1 U2047 ( .A(n2070), .B(n2071), .Z(n2069) );
  OR2_X1 U2048 ( .A1(n2072), .A2(n2073), .ZN(n2071) );
  OR2_X1 U2049 ( .A1(n2074), .A2(n2075), .ZN(Result_23_) );
  AND2_X1 U2050 ( .A1(n2076), .A2(operation), .ZN(n2075) );
  XNOR2_X1 U2051 ( .A(n2077), .B(n2078), .ZN(n2076) );
  XOR2_X1 U2052 ( .A(n2079), .B(n2080), .Z(n2078) );
  AND2_X1 U2053 ( .A1(n2081), .A2(n1968), .ZN(n2074) );
  OR3_X1 U2054 ( .A1(n2082), .A2(n2083), .A3(n2084), .ZN(n2081) );
  INV_X1 U2055 ( .A(n2085), .ZN(n2084) );
  OR2_X1 U2056 ( .A1(n2086), .A2(n2087), .ZN(n2085) );
  AND2_X1 U2057 ( .A1(n2088), .A2(n2089), .ZN(n2083) );
  XNOR2_X1 U2058 ( .A(a_7_), .B(n2086), .ZN(n2088) );
  AND3_X1 U2059 ( .A1(n2086), .A2(n2090), .A3(b_7_), .ZN(n2082) );
  OR2_X1 U2060 ( .A1(n2091), .A2(n2092), .ZN(Result_22_) );
  AND2_X1 U2061 ( .A1(n2093), .A2(operation), .ZN(n2092) );
  XNOR2_X1 U2062 ( .A(n2094), .B(n2095), .ZN(n2093) );
  XOR2_X1 U2063 ( .A(n2096), .B(n2097), .Z(n2095) );
  AND2_X1 U2064 ( .A1(n2098), .A2(n1968), .ZN(n2091) );
  XOR2_X1 U2065 ( .A(n2099), .B(n2100), .Z(n2098) );
  OR2_X1 U2066 ( .A1(n2101), .A2(n2102), .ZN(n2100) );
  OR2_X1 U2067 ( .A1(n2103), .A2(n2104), .ZN(Result_21_) );
  AND2_X1 U2068 ( .A1(n2105), .A2(operation), .ZN(n2104) );
  XNOR2_X1 U2069 ( .A(n2106), .B(n2107), .ZN(n2105) );
  XOR2_X1 U2070 ( .A(n2108), .B(n2109), .Z(n2107) );
  AND2_X1 U2071 ( .A1(n2110), .A2(n1968), .ZN(n2103) );
  OR3_X1 U2072 ( .A1(n2111), .A2(n2112), .A3(n2113), .ZN(n2110) );
  INV_X1 U2073 ( .A(n2114), .ZN(n2113) );
  OR2_X1 U2074 ( .A1(n2115), .A2(n2116), .ZN(n2114) );
  AND2_X1 U2075 ( .A1(n2117), .A2(n2118), .ZN(n2112) );
  XNOR2_X1 U2076 ( .A(a_5_), .B(n2115), .ZN(n2117) );
  AND3_X1 U2077 ( .A1(n2115), .A2(n2119), .A3(b_5_), .ZN(n2111) );
  OR2_X1 U2078 ( .A1(n2120), .A2(n2121), .ZN(Result_20_) );
  AND2_X1 U2079 ( .A1(n2122), .A2(operation), .ZN(n2121) );
  XNOR2_X1 U2080 ( .A(n2123), .B(n2124), .ZN(n2122) );
  XOR2_X1 U2081 ( .A(n2125), .B(n2126), .Z(n2124) );
  AND2_X1 U2082 ( .A1(n2127), .A2(n1968), .ZN(n2120) );
  XOR2_X1 U2083 ( .A(n2128), .B(n2129), .Z(n2127) );
  OR2_X1 U2084 ( .A1(n2130), .A2(n2131), .ZN(n2129) );
  AND2_X1 U2085 ( .A1(operation), .A2(n2132), .ZN(Result_1_) );
  XOR2_X1 U2086 ( .A(n2133), .B(n2134), .Z(n2132) );
  AND2_X1 U2087 ( .A1(n2135), .A2(n2136), .ZN(n2134) );
  OR2_X1 U2088 ( .A1(n2137), .A2(n2138), .ZN(n2136) );
  AND2_X1 U2089 ( .A1(n2139), .A2(n2140), .ZN(n2137) );
  INV_X1 U2090 ( .A(n2141), .ZN(n2135) );
  OR2_X1 U2091 ( .A1(n2142), .A2(n2143), .ZN(Result_19_) );
  AND2_X1 U2092 ( .A1(n2144), .A2(operation), .ZN(n2143) );
  XNOR2_X1 U2093 ( .A(n2145), .B(n2146), .ZN(n2144) );
  XOR2_X1 U2094 ( .A(n2147), .B(n2148), .Z(n2146) );
  AND2_X1 U2095 ( .A1(n2149), .A2(n1968), .ZN(n2142) );
  OR3_X1 U2096 ( .A1(n2150), .A2(n2151), .A3(n2152), .ZN(n2149) );
  INV_X1 U2097 ( .A(n2153), .ZN(n2152) );
  OR2_X1 U2098 ( .A1(n2154), .A2(n2155), .ZN(n2153) );
  AND2_X1 U2099 ( .A1(n2156), .A2(n2157), .ZN(n2151) );
  XNOR2_X1 U2100 ( .A(a_3_), .B(n2154), .ZN(n2156) );
  AND3_X1 U2101 ( .A1(n2154), .A2(n2158), .A3(b_3_), .ZN(n2150) );
  OR2_X1 U2102 ( .A1(n2159), .A2(n2160), .ZN(Result_18_) );
  AND2_X1 U2103 ( .A1(n2161), .A2(operation), .ZN(n2160) );
  XNOR2_X1 U2104 ( .A(n2162), .B(n2163), .ZN(n2161) );
  XOR2_X1 U2105 ( .A(n2164), .B(n2165), .Z(n2163) );
  AND2_X1 U2106 ( .A1(n2166), .A2(n1968), .ZN(n2159) );
  XOR2_X1 U2107 ( .A(n2167), .B(n2168), .Z(n2166) );
  OR2_X1 U2108 ( .A1(n2169), .A2(n2170), .ZN(n2168) );
  OR2_X1 U2109 ( .A1(n2171), .A2(n2172), .ZN(Result_17_) );
  AND2_X1 U2110 ( .A1(n2173), .A2(operation), .ZN(n2172) );
  XNOR2_X1 U2111 ( .A(n2174), .B(n2175), .ZN(n2173) );
  XOR2_X1 U2112 ( .A(n2176), .B(n2177), .Z(n2175) );
  AND2_X1 U2113 ( .A1(n2178), .A2(n1968), .ZN(n2171) );
  OR3_X1 U2114 ( .A1(n2179), .A2(n2180), .A3(n2181), .ZN(n2178) );
  INV_X1 U2115 ( .A(n2182), .ZN(n2181) );
  OR2_X1 U2116 ( .A1(n2183), .A2(n2184), .ZN(n2182) );
  AND2_X1 U2117 ( .A1(n2185), .A2(n2186), .ZN(n2180) );
  XNOR2_X1 U2118 ( .A(a_1_), .B(n2183), .ZN(n2185) );
  AND3_X1 U2119 ( .A1(n2183), .A2(n2187), .A3(b_1_), .ZN(n2179) );
  OR2_X1 U2120 ( .A1(n2188), .A2(n2189), .ZN(Result_16_) );
  AND2_X1 U2121 ( .A1(n2190), .A2(operation), .ZN(n2189) );
  XNOR2_X1 U2122 ( .A(n2191), .B(n2192), .ZN(n2190) );
  XOR2_X1 U2123 ( .A(n2193), .B(n2194), .Z(n2192) );
  AND2_X1 U2124 ( .A1(n2195), .A2(n1968), .ZN(n2188) );
  INV_X1 U2125 ( .A(operation), .ZN(n1968) );
  XOR2_X1 U2126 ( .A(n2196), .B(n2197), .Z(n2195) );
  XNOR2_X1 U2127 ( .A(a_0_), .B(b_0_), .ZN(n2197) );
  OR2_X1 U2128 ( .A1(n2198), .A2(n2199), .ZN(n2196) );
  AND2_X1 U2129 ( .A1(n2187), .A2(n2186), .ZN(n2199) );
  AND2_X1 U2130 ( .A1(n2183), .A2(n2184), .ZN(n2198) );
  OR2_X1 U2131 ( .A1(n2200), .A2(n2169), .ZN(n2183) );
  AND2_X1 U2132 ( .A1(n2201), .A2(n2202), .ZN(n2169) );
  AND2_X1 U2133 ( .A1(n2167), .A2(n2203), .ZN(n2200) );
  OR2_X1 U2134 ( .A1(n2204), .A2(n2205), .ZN(n2167) );
  AND2_X1 U2135 ( .A1(n2158), .A2(n2157), .ZN(n2205) );
  AND2_X1 U2136 ( .A1(n2154), .A2(n2155), .ZN(n2204) );
  OR2_X1 U2137 ( .A1(n2206), .A2(n2130), .ZN(n2154) );
  AND2_X1 U2138 ( .A1(n2207), .A2(n2208), .ZN(n2130) );
  AND2_X1 U2139 ( .A1(n2128), .A2(n2209), .ZN(n2206) );
  OR2_X1 U2140 ( .A1(n2210), .A2(n2211), .ZN(n2128) );
  AND2_X1 U2141 ( .A1(n2119), .A2(n2118), .ZN(n2211) );
  AND2_X1 U2142 ( .A1(n2115), .A2(n2116), .ZN(n2210) );
  OR2_X1 U2143 ( .A1(n2212), .A2(n2101), .ZN(n2115) );
  AND2_X1 U2144 ( .A1(n2213), .A2(n2214), .ZN(n2101) );
  AND2_X1 U2145 ( .A1(n2099), .A2(n2215), .ZN(n2212) );
  OR2_X1 U2146 ( .A1(n2216), .A2(n2217), .ZN(n2099) );
  AND2_X1 U2147 ( .A1(n2090), .A2(n2089), .ZN(n2217) );
  AND2_X1 U2148 ( .A1(n2086), .A2(n2087), .ZN(n2216) );
  OR2_X1 U2149 ( .A1(n2218), .A2(n2072), .ZN(n2086) );
  AND2_X1 U2150 ( .A1(n2219), .A2(n2220), .ZN(n2072) );
  AND2_X1 U2151 ( .A1(n2070), .A2(n2221), .ZN(n2218) );
  OR2_X1 U2152 ( .A1(n2222), .A2(n2223), .ZN(n2070) );
  AND2_X1 U2153 ( .A1(n2061), .A2(n2060), .ZN(n2223) );
  AND2_X1 U2154 ( .A1(n2057), .A2(n2058), .ZN(n2222) );
  OR2_X1 U2155 ( .A1(n2224), .A2(n2043), .ZN(n2057) );
  AND2_X1 U2156 ( .A1(n2225), .A2(n2226), .ZN(n2043) );
  AND2_X1 U2157 ( .A1(n2041), .A2(n2227), .ZN(n2224) );
  OR2_X1 U2158 ( .A1(n2228), .A2(n2229), .ZN(n2041) );
  AND2_X1 U2159 ( .A1(n2032), .A2(n2031), .ZN(n2229) );
  AND2_X1 U2160 ( .A1(n2028), .A2(n2029), .ZN(n2228) );
  OR2_X1 U2161 ( .A1(n2230), .A2(n2015), .ZN(n2028) );
  AND2_X1 U2162 ( .A1(n2231), .A2(n2232), .ZN(n2015) );
  AND2_X1 U2163 ( .A1(n2012), .A2(n2233), .ZN(n2230) );
  OR2_X1 U2164 ( .A1(n2234), .A2(n2235), .ZN(n2012) );
  AND2_X1 U2165 ( .A1(n2003), .A2(n2002), .ZN(n2235) );
  AND2_X1 U2166 ( .A1(n2000), .A2(n1999), .ZN(n2234) );
  AND2_X1 U2167 ( .A1(n2236), .A2(n2237), .ZN(n2000) );
  OR2_X1 U2168 ( .A1(n1974), .A2(n2238), .ZN(n2237) );
  AND2_X1 U2169 ( .A1(n2239), .A2(n1966), .ZN(n2238) );
  OR2_X1 U2170 ( .A1(n2240), .A2(n1969), .ZN(n1966) );
  AND2_X1 U2171 ( .A1(operation), .A2(n2241), .ZN(Result_15_) );
  XNOR2_X1 U2172 ( .A(n2242), .B(n2243), .ZN(n2241) );
  AND3_X1 U2173 ( .A1(n2244), .A2(n2245), .A3(operation), .ZN(Result_14_) );
  OR2_X1 U2174 ( .A1(n2246), .A2(n2247), .ZN(n2244) );
  AND2_X1 U2175 ( .A1(n2248), .A2(n2243), .ZN(n2246) );
  AND2_X1 U2176 ( .A1(operation), .A2(n2249), .ZN(Result_13_) );
  XNOR2_X1 U2177 ( .A(n2250), .B(n2251), .ZN(n2249) );
  OR2_X1 U2178 ( .A1(n2252), .A2(n2253), .ZN(n2251) );
  AND2_X1 U2179 ( .A1(n2254), .A2(n2255), .ZN(n2252) );
  OR2_X1 U2180 ( .A1(n2256), .A2(n2257), .ZN(n2254) );
  AND2_X1 U2181 ( .A1(n2258), .A2(operation), .ZN(Result_12_) );
  XOR2_X1 U2182 ( .A(n2259), .B(n2260), .Z(n2258) );
  AND2_X1 U2183 ( .A1(n2261), .A2(n2262), .ZN(n2260) );
  OR2_X1 U2184 ( .A1(n2263), .A2(n2264), .ZN(n2262) );
  INV_X1 U2185 ( .A(n2265), .ZN(n2261) );
  AND2_X1 U2186 ( .A1(n2266), .A2(operation), .ZN(Result_11_) );
  XOR2_X1 U2187 ( .A(n2267), .B(n2268), .Z(n2266) );
  AND2_X1 U2188 ( .A1(n2269), .A2(n2270), .ZN(n2268) );
  OR2_X1 U2189 ( .A1(n2271), .A2(n2272), .ZN(n2270) );
  AND2_X1 U2190 ( .A1(n2273), .A2(n2274), .ZN(n2271) );
  INV_X1 U2191 ( .A(n2275), .ZN(n2269) );
  AND2_X1 U2192 ( .A1(n2276), .A2(operation), .ZN(Result_10_) );
  XOR2_X1 U2193 ( .A(n2277), .B(n2278), .Z(n2276) );
  AND2_X1 U2194 ( .A1(n2279), .A2(n2280), .ZN(n2278) );
  OR2_X1 U2195 ( .A1(n2281), .A2(n2282), .ZN(n2280) );
  AND2_X1 U2196 ( .A1(n2283), .A2(n2284), .ZN(n2281) );
  INV_X1 U2197 ( .A(n2285), .ZN(n2279) );
  AND2_X1 U2198 ( .A1(operation), .A2(n2286), .ZN(Result_0_) );
  OR3_X1 U2199 ( .A1(n2141), .A2(n2287), .A3(n2288), .ZN(n2286) );
  INV_X1 U2200 ( .A(n2289), .ZN(n2288) );
  OR2_X1 U2201 ( .A1(n2290), .A2(n2291), .ZN(n2289) );
  AND2_X1 U2202 ( .A1(n2133), .A2(n2138), .ZN(n2287) );
  AND2_X1 U2203 ( .A1(n1985), .A2(n1986), .ZN(n2133) );
  XNOR2_X1 U2204 ( .A(n2140), .B(n2292), .ZN(n1986) );
  OR2_X1 U2205 ( .A1(n2293), .A2(n2294), .ZN(n1985) );
  OR2_X1 U2206 ( .A1(n2295), .A2(n1962), .ZN(n2293) );
  AND3_X1 U2207 ( .A1(n1961), .A2(n1960), .A3(n1958), .ZN(n1962) );
  INV_X1 U2208 ( .A(n2296), .ZN(n1960) );
  AND2_X1 U2209 ( .A1(n1954), .A2(n1958), .ZN(n2295) );
  INV_X1 U2210 ( .A(n2297), .ZN(n1958) );
  OR2_X1 U2211 ( .A1(n2298), .A2(n2294), .ZN(n2297) );
  INV_X1 U2212 ( .A(n2299), .ZN(n2294) );
  OR2_X1 U2213 ( .A1(n2300), .A2(n2301), .ZN(n2299) );
  AND2_X1 U2214 ( .A1(n2300), .A2(n2301), .ZN(n2298) );
  OR2_X1 U2215 ( .A1(n2302), .A2(n2303), .ZN(n2301) );
  AND2_X1 U2216 ( .A1(n2304), .A2(n2305), .ZN(n2303) );
  AND2_X1 U2217 ( .A1(n2306), .A2(n2307), .ZN(n2302) );
  OR2_X1 U2218 ( .A1(n2305), .A2(n2304), .ZN(n2307) );
  XOR2_X1 U2219 ( .A(n2308), .B(n2309), .Z(n2300) );
  XOR2_X1 U2220 ( .A(n2310), .B(n2311), .Z(n2309) );
  AND2_X1 U2221 ( .A1(n1951), .A2(n1952), .ZN(n1954) );
  XNOR2_X1 U2222 ( .A(n1961), .B(n2296), .ZN(n1952) );
  OR2_X1 U2223 ( .A1(n2312), .A2(n2313), .ZN(n2296) );
  AND2_X1 U2224 ( .A1(n2314), .A2(n2315), .ZN(n2313) );
  AND2_X1 U2225 ( .A1(n2316), .A2(n2317), .ZN(n2312) );
  OR2_X1 U2226 ( .A1(n2315), .A2(n2314), .ZN(n2317) );
  XNOR2_X1 U2227 ( .A(n2306), .B(n2318), .ZN(n1961) );
  XOR2_X1 U2228 ( .A(n2305), .B(n2304), .Z(n2318) );
  OR2_X1 U2229 ( .A1(n2157), .A2(n2291), .ZN(n2304) );
  OR2_X1 U2230 ( .A1(n2319), .A2(n2320), .ZN(n2305) );
  AND2_X1 U2231 ( .A1(n2321), .A2(n2322), .ZN(n2320) );
  AND2_X1 U2232 ( .A1(n2323), .A2(n2324), .ZN(n2319) );
  OR2_X1 U2233 ( .A1(n2322), .A2(n2321), .ZN(n2324) );
  XOR2_X1 U2234 ( .A(n2325), .B(n2326), .Z(n2306) );
  XOR2_X1 U2235 ( .A(n2327), .B(n2328), .Z(n2326) );
  OR2_X1 U2236 ( .A1(n2329), .A2(n2330), .ZN(n1951) );
  OR2_X1 U2237 ( .A1(n2331), .A2(n1949), .ZN(n2329) );
  AND3_X1 U2238 ( .A1(n1948), .A2(n1947), .A3(n1945), .ZN(n1949) );
  INV_X1 U2239 ( .A(n2332), .ZN(n1947) );
  AND2_X1 U2240 ( .A1(n1941), .A2(n1945), .ZN(n2331) );
  INV_X1 U2241 ( .A(n2333), .ZN(n1945) );
  OR2_X1 U2242 ( .A1(n2334), .A2(n2330), .ZN(n2333) );
  INV_X1 U2243 ( .A(n2335), .ZN(n2330) );
  OR2_X1 U2244 ( .A1(n2336), .A2(n2337), .ZN(n2335) );
  AND2_X1 U2245 ( .A1(n2336), .A2(n2337), .ZN(n2334) );
  OR2_X1 U2246 ( .A1(n2338), .A2(n2339), .ZN(n2337) );
  AND2_X1 U2247 ( .A1(n2340), .A2(n2341), .ZN(n2339) );
  AND2_X1 U2248 ( .A1(n2342), .A2(n2343), .ZN(n2338) );
  OR2_X1 U2249 ( .A1(n2341), .A2(n2340), .ZN(n2343) );
  XOR2_X1 U2250 ( .A(n2316), .B(n2344), .Z(n2336) );
  XOR2_X1 U2251 ( .A(n2315), .B(n2314), .Z(n2344) );
  OR2_X1 U2252 ( .A1(n2208), .A2(n2291), .ZN(n2314) );
  OR2_X1 U2253 ( .A1(n2345), .A2(n2346), .ZN(n2315) );
  AND2_X1 U2254 ( .A1(n2347), .A2(n2348), .ZN(n2346) );
  AND2_X1 U2255 ( .A1(n2349), .A2(n2350), .ZN(n2345) );
  OR2_X1 U2256 ( .A1(n2348), .A2(n2347), .ZN(n2350) );
  XOR2_X1 U2257 ( .A(n2323), .B(n2351), .Z(n2316) );
  XOR2_X1 U2258 ( .A(n2322), .B(n2321), .Z(n2351) );
  OR2_X1 U2259 ( .A1(n2157), .A2(n2187), .ZN(n2321) );
  OR2_X1 U2260 ( .A1(n2352), .A2(n2353), .ZN(n2322) );
  AND2_X1 U2261 ( .A1(n2354), .A2(n2355), .ZN(n2353) );
  AND2_X1 U2262 ( .A1(n2356), .A2(n2357), .ZN(n2352) );
  OR2_X1 U2263 ( .A1(n2355), .A2(n2354), .ZN(n2357) );
  XNOR2_X1 U2264 ( .A(n2358), .B(n2359), .ZN(n2323) );
  XNOR2_X1 U2265 ( .A(n2203), .B(n2360), .ZN(n2358) );
  AND2_X1 U2266 ( .A1(n1938), .A2(n1939), .ZN(n1941) );
  XNOR2_X1 U2267 ( .A(n1948), .B(n2332), .ZN(n1939) );
  OR2_X1 U2268 ( .A1(n2361), .A2(n2362), .ZN(n2332) );
  AND2_X1 U2269 ( .A1(n2363), .A2(n2364), .ZN(n2362) );
  AND2_X1 U2270 ( .A1(n2365), .A2(n2366), .ZN(n2361) );
  OR2_X1 U2271 ( .A1(n2364), .A2(n2363), .ZN(n2366) );
  XNOR2_X1 U2272 ( .A(n2342), .B(n2367), .ZN(n1948) );
  XOR2_X1 U2273 ( .A(n2341), .B(n2340), .Z(n2367) );
  OR2_X1 U2274 ( .A1(n2118), .A2(n2291), .ZN(n2340) );
  OR2_X1 U2275 ( .A1(n2368), .A2(n2369), .ZN(n2341) );
  AND2_X1 U2276 ( .A1(n2370), .A2(n2371), .ZN(n2369) );
  AND2_X1 U2277 ( .A1(n2372), .A2(n2373), .ZN(n2368) );
  OR2_X1 U2278 ( .A1(n2371), .A2(n2370), .ZN(n2373) );
  XOR2_X1 U2279 ( .A(n2349), .B(n2374), .Z(n2342) );
  XOR2_X1 U2280 ( .A(n2348), .B(n2347), .Z(n2374) );
  OR2_X1 U2281 ( .A1(n2208), .A2(n2187), .ZN(n2347) );
  OR2_X1 U2282 ( .A1(n2375), .A2(n2376), .ZN(n2348) );
  AND2_X1 U2283 ( .A1(n2377), .A2(n2378), .ZN(n2376) );
  AND2_X1 U2284 ( .A1(n2379), .A2(n2380), .ZN(n2375) );
  OR2_X1 U2285 ( .A1(n2378), .A2(n2377), .ZN(n2380) );
  XOR2_X1 U2286 ( .A(n2356), .B(n2381), .Z(n2349) );
  XOR2_X1 U2287 ( .A(n2355), .B(n2354), .Z(n2381) );
  OR2_X1 U2288 ( .A1(n2157), .A2(n2201), .ZN(n2354) );
  OR2_X1 U2289 ( .A1(n2382), .A2(n2383), .ZN(n2355) );
  AND2_X1 U2290 ( .A1(n2155), .A2(n2384), .ZN(n2383) );
  AND2_X1 U2291 ( .A1(n2385), .A2(n2386), .ZN(n2382) );
  OR2_X1 U2292 ( .A1(n2384), .A2(n2155), .ZN(n2386) );
  XOR2_X1 U2293 ( .A(n2387), .B(n2388), .Z(n2356) );
  XOR2_X1 U2294 ( .A(n2389), .B(n2390), .Z(n2388) );
  OR2_X1 U2295 ( .A1(n2391), .A2(n2392), .ZN(n1938) );
  OR2_X1 U2296 ( .A1(n2393), .A2(n1936), .ZN(n2391) );
  AND3_X1 U2297 ( .A1(n1935), .A2(n1934), .A3(n1932), .ZN(n1936) );
  INV_X1 U2298 ( .A(n2394), .ZN(n1934) );
  AND2_X1 U2299 ( .A1(n1928), .A2(n1932), .ZN(n2393) );
  INV_X1 U2300 ( .A(n2395), .ZN(n1932) );
  OR2_X1 U2301 ( .A1(n2396), .A2(n2392), .ZN(n2395) );
  INV_X1 U2302 ( .A(n2397), .ZN(n2392) );
  OR2_X1 U2303 ( .A1(n2398), .A2(n2399), .ZN(n2397) );
  AND2_X1 U2304 ( .A1(n2398), .A2(n2399), .ZN(n2396) );
  OR2_X1 U2305 ( .A1(n2400), .A2(n2401), .ZN(n2399) );
  AND2_X1 U2306 ( .A1(n2402), .A2(n2403), .ZN(n2401) );
  AND2_X1 U2307 ( .A1(n2404), .A2(n2405), .ZN(n2400) );
  OR2_X1 U2308 ( .A1(n2403), .A2(n2402), .ZN(n2405) );
  XOR2_X1 U2309 ( .A(n2365), .B(n2406), .Z(n2398) );
  XOR2_X1 U2310 ( .A(n2364), .B(n2363), .Z(n2406) );
  OR2_X1 U2311 ( .A1(n2214), .A2(n2291), .ZN(n2363) );
  OR2_X1 U2312 ( .A1(n2407), .A2(n2408), .ZN(n2364) );
  AND2_X1 U2313 ( .A1(n2409), .A2(n2410), .ZN(n2408) );
  AND2_X1 U2314 ( .A1(n2411), .A2(n2412), .ZN(n2407) );
  OR2_X1 U2315 ( .A1(n2410), .A2(n2409), .ZN(n2412) );
  XOR2_X1 U2316 ( .A(n2372), .B(n2413), .Z(n2365) );
  XOR2_X1 U2317 ( .A(n2371), .B(n2370), .Z(n2413) );
  OR2_X1 U2318 ( .A1(n2118), .A2(n2187), .ZN(n2370) );
  OR2_X1 U2319 ( .A1(n2414), .A2(n2415), .ZN(n2371) );
  AND2_X1 U2320 ( .A1(n2416), .A2(n2417), .ZN(n2415) );
  AND2_X1 U2321 ( .A1(n2418), .A2(n2419), .ZN(n2414) );
  OR2_X1 U2322 ( .A1(n2417), .A2(n2416), .ZN(n2419) );
  XOR2_X1 U2323 ( .A(n2379), .B(n2420), .Z(n2372) );
  XOR2_X1 U2324 ( .A(n2378), .B(n2377), .Z(n2420) );
  OR2_X1 U2325 ( .A1(n2208), .A2(n2201), .ZN(n2377) );
  OR2_X1 U2326 ( .A1(n2421), .A2(n2422), .ZN(n2378) );
  AND2_X1 U2327 ( .A1(n2423), .A2(n2424), .ZN(n2422) );
  AND2_X1 U2328 ( .A1(n2425), .A2(n2426), .ZN(n2421) );
  OR2_X1 U2329 ( .A1(n2424), .A2(n2423), .ZN(n2426) );
  XOR2_X1 U2330 ( .A(n2385), .B(n2427), .Z(n2379) );
  XOR2_X1 U2331 ( .A(n2384), .B(n2155), .Z(n2427) );
  OR2_X1 U2332 ( .A1(n2158), .A2(n2157), .ZN(n2155) );
  OR2_X1 U2333 ( .A1(n2428), .A2(n2429), .ZN(n2384) );
  AND2_X1 U2334 ( .A1(n2430), .A2(n2431), .ZN(n2429) );
  AND2_X1 U2335 ( .A1(n2432), .A2(n2433), .ZN(n2428) );
  OR2_X1 U2336 ( .A1(n2431), .A2(n2430), .ZN(n2433) );
  XOR2_X1 U2337 ( .A(n2434), .B(n2435), .Z(n2385) );
  XOR2_X1 U2338 ( .A(n2436), .B(n2437), .Z(n2435) );
  AND2_X1 U2339 ( .A1(n1925), .A2(n1926), .ZN(n1928) );
  XNOR2_X1 U2340 ( .A(n1935), .B(n2394), .ZN(n1926) );
  OR2_X1 U2341 ( .A1(n2438), .A2(n2439), .ZN(n2394) );
  AND2_X1 U2342 ( .A1(n2440), .A2(n2441), .ZN(n2439) );
  AND2_X1 U2343 ( .A1(n2442), .A2(n2443), .ZN(n2438) );
  OR2_X1 U2344 ( .A1(n2441), .A2(n2440), .ZN(n2443) );
  XNOR2_X1 U2345 ( .A(n2404), .B(n2444), .ZN(n1935) );
  XOR2_X1 U2346 ( .A(n2403), .B(n2402), .Z(n2444) );
  OR2_X1 U2347 ( .A1(n2089), .A2(n2291), .ZN(n2402) );
  OR2_X1 U2348 ( .A1(n2445), .A2(n2446), .ZN(n2403) );
  AND2_X1 U2349 ( .A1(n2447), .A2(n2448), .ZN(n2446) );
  AND2_X1 U2350 ( .A1(n2449), .A2(n2450), .ZN(n2445) );
  OR2_X1 U2351 ( .A1(n2448), .A2(n2447), .ZN(n2450) );
  XOR2_X1 U2352 ( .A(n2411), .B(n2451), .Z(n2404) );
  XOR2_X1 U2353 ( .A(n2410), .B(n2409), .Z(n2451) );
  OR2_X1 U2354 ( .A1(n2214), .A2(n2187), .ZN(n2409) );
  OR2_X1 U2355 ( .A1(n2452), .A2(n2453), .ZN(n2410) );
  AND2_X1 U2356 ( .A1(n2454), .A2(n2455), .ZN(n2453) );
  AND2_X1 U2357 ( .A1(n2456), .A2(n2457), .ZN(n2452) );
  OR2_X1 U2358 ( .A1(n2455), .A2(n2454), .ZN(n2457) );
  XOR2_X1 U2359 ( .A(n2418), .B(n2458), .Z(n2411) );
  XOR2_X1 U2360 ( .A(n2417), .B(n2416), .Z(n2458) );
  OR2_X1 U2361 ( .A1(n2118), .A2(n2201), .ZN(n2416) );
  OR2_X1 U2362 ( .A1(n2459), .A2(n2460), .ZN(n2417) );
  AND2_X1 U2363 ( .A1(n2461), .A2(n2462), .ZN(n2460) );
  AND2_X1 U2364 ( .A1(n2463), .A2(n2464), .ZN(n2459) );
  OR2_X1 U2365 ( .A1(n2462), .A2(n2461), .ZN(n2464) );
  XOR2_X1 U2366 ( .A(n2425), .B(n2465), .Z(n2418) );
  XOR2_X1 U2367 ( .A(n2424), .B(n2423), .Z(n2465) );
  OR2_X1 U2368 ( .A1(n2208), .A2(n2158), .ZN(n2423) );
  OR2_X1 U2369 ( .A1(n2466), .A2(n2467), .ZN(n2424) );
  AND2_X1 U2370 ( .A1(n2468), .A2(n2209), .ZN(n2467) );
  AND2_X1 U2371 ( .A1(n2469), .A2(n2470), .ZN(n2466) );
  OR2_X1 U2372 ( .A1(n2209), .A2(n2468), .ZN(n2470) );
  XOR2_X1 U2373 ( .A(n2432), .B(n2471), .Z(n2425) );
  XOR2_X1 U2374 ( .A(n2431), .B(n2430), .Z(n2471) );
  OR2_X1 U2375 ( .A1(n2207), .A2(n2157), .ZN(n2430) );
  OR2_X1 U2376 ( .A1(n2472), .A2(n2473), .ZN(n2431) );
  AND2_X1 U2377 ( .A1(n2474), .A2(n2475), .ZN(n2473) );
  AND2_X1 U2378 ( .A1(n2476), .A2(n2477), .ZN(n2472) );
  OR2_X1 U2379 ( .A1(n2475), .A2(n2474), .ZN(n2477) );
  XOR2_X1 U2380 ( .A(n2478), .B(n2479), .Z(n2432) );
  XOR2_X1 U2381 ( .A(n2480), .B(n2481), .Z(n2479) );
  OR2_X1 U2382 ( .A1(n2482), .A2(n2483), .ZN(n1925) );
  OR2_X1 U2383 ( .A1(n2484), .A2(n1923), .ZN(n2482) );
  AND3_X1 U2384 ( .A1(n1922), .A2(n1921), .A3(n1919), .ZN(n1923) );
  INV_X1 U2385 ( .A(n2485), .ZN(n1921) );
  AND2_X1 U2386 ( .A1(n1919), .A2(n1915), .ZN(n2484) );
  OR2_X1 U2387 ( .A1(n2486), .A2(n2285), .ZN(n1915) );
  AND3_X1 U2388 ( .A1(n2284), .A2(n2282), .A3(n2283), .ZN(n2285) );
  INV_X1 U2389 ( .A(n2487), .ZN(n2283) );
  AND2_X1 U2390 ( .A1(n2282), .A2(n2277), .ZN(n2486) );
  OR2_X1 U2391 ( .A1(n2488), .A2(n2275), .ZN(n2277) );
  AND3_X1 U2392 ( .A1(n2274), .A2(n2272), .A3(n2273), .ZN(n2275) );
  INV_X1 U2393 ( .A(n2489), .ZN(n2273) );
  AND2_X1 U2394 ( .A1(n2272), .A2(n2267), .ZN(n2488) );
  OR2_X1 U2395 ( .A1(n2490), .A2(n2265), .ZN(n2267) );
  AND2_X1 U2396 ( .A1(n2264), .A2(n2263), .ZN(n2265) );
  AND2_X1 U2397 ( .A1(n2264), .A2(n2259), .ZN(n2490) );
  OR2_X1 U2398 ( .A1(n2491), .A2(n2253), .ZN(n2259) );
  INV_X1 U2399 ( .A(n2492), .ZN(n2253) );
  OR3_X1 U2400 ( .A1(n2257), .A2(n2256), .A3(n2255), .ZN(n2492) );
  INV_X1 U2401 ( .A(n2493), .ZN(n2491) );
  OR2_X1 U2402 ( .A1(n2245), .A2(n2255), .ZN(n2493) );
  OR2_X1 U2403 ( .A1(n2494), .A2(n2263), .ZN(n2255) );
  INV_X1 U2404 ( .A(n2495), .ZN(n2263) );
  OR2_X1 U2405 ( .A1(n2496), .A2(n2497), .ZN(n2495) );
  AND2_X1 U2406 ( .A1(n2496), .A2(n2497), .ZN(n2494) );
  OR2_X1 U2407 ( .A1(n2498), .A2(n2499), .ZN(n2497) );
  AND2_X1 U2408 ( .A1(n2500), .A2(n2501), .ZN(n2499) );
  AND2_X1 U2409 ( .A1(n2502), .A2(n2503), .ZN(n2498) );
  OR2_X1 U2410 ( .A1(n2501), .A2(n2500), .ZN(n2503) );
  XOR2_X1 U2411 ( .A(n2504), .B(n2505), .Z(n2496) );
  XOR2_X1 U2412 ( .A(n2506), .B(n2507), .Z(n2505) );
  INV_X1 U2413 ( .A(n2250), .ZN(n2245) );
  AND3_X1 U2414 ( .A1(n2243), .A2(n2247), .A3(n2248), .ZN(n2250) );
  INV_X1 U2415 ( .A(n2242), .ZN(n2248) );
  OR2_X1 U2416 ( .A1(n2508), .A2(n2509), .ZN(n2242) );
  AND2_X1 U2417 ( .A1(n2194), .A2(n2193), .ZN(n2509) );
  AND2_X1 U2418 ( .A1(n2191), .A2(n2510), .ZN(n2508) );
  OR2_X1 U2419 ( .A1(n2194), .A2(n2193), .ZN(n2510) );
  OR2_X1 U2420 ( .A1(n2511), .A2(n2512), .ZN(n2193) );
  AND2_X1 U2421 ( .A1(n2177), .A2(n2176), .ZN(n2512) );
  AND2_X1 U2422 ( .A1(n2174), .A2(n2513), .ZN(n2511) );
  OR2_X1 U2423 ( .A1(n2177), .A2(n2176), .ZN(n2513) );
  OR2_X1 U2424 ( .A1(n2514), .A2(n2515), .ZN(n2176) );
  AND2_X1 U2425 ( .A1(n2165), .A2(n2164), .ZN(n2515) );
  AND2_X1 U2426 ( .A1(n2162), .A2(n2516), .ZN(n2514) );
  OR2_X1 U2427 ( .A1(n2165), .A2(n2164), .ZN(n2516) );
  OR2_X1 U2428 ( .A1(n2517), .A2(n2518), .ZN(n2164) );
  AND2_X1 U2429 ( .A1(n2148), .A2(n2147), .ZN(n2518) );
  AND2_X1 U2430 ( .A1(n2145), .A2(n2519), .ZN(n2517) );
  OR2_X1 U2431 ( .A1(n2148), .A2(n2147), .ZN(n2519) );
  OR2_X1 U2432 ( .A1(n2520), .A2(n2521), .ZN(n2147) );
  AND2_X1 U2433 ( .A1(n2126), .A2(n2125), .ZN(n2521) );
  AND2_X1 U2434 ( .A1(n2123), .A2(n2522), .ZN(n2520) );
  OR2_X1 U2435 ( .A1(n2126), .A2(n2125), .ZN(n2522) );
  OR2_X1 U2436 ( .A1(n2523), .A2(n2524), .ZN(n2125) );
  AND2_X1 U2437 ( .A1(n2109), .A2(n2108), .ZN(n2524) );
  AND2_X1 U2438 ( .A1(n2106), .A2(n2525), .ZN(n2523) );
  OR2_X1 U2439 ( .A1(n2109), .A2(n2108), .ZN(n2525) );
  OR2_X1 U2440 ( .A1(n2526), .A2(n2527), .ZN(n2108) );
  AND2_X1 U2441 ( .A1(n2097), .A2(n2096), .ZN(n2527) );
  AND2_X1 U2442 ( .A1(n2094), .A2(n2528), .ZN(n2526) );
  OR2_X1 U2443 ( .A1(n2097), .A2(n2096), .ZN(n2528) );
  OR2_X1 U2444 ( .A1(n2529), .A2(n2530), .ZN(n2096) );
  AND2_X1 U2445 ( .A1(n2080), .A2(n2079), .ZN(n2530) );
  AND2_X1 U2446 ( .A1(n2077), .A2(n2531), .ZN(n2529) );
  OR2_X1 U2447 ( .A1(n2080), .A2(n2079), .ZN(n2531) );
  OR2_X1 U2448 ( .A1(n2532), .A2(n2533), .ZN(n2079) );
  AND2_X1 U2449 ( .A1(n2068), .A2(n2067), .ZN(n2533) );
  AND2_X1 U2450 ( .A1(n2065), .A2(n2534), .ZN(n2532) );
  OR2_X1 U2451 ( .A1(n2068), .A2(n2067), .ZN(n2534) );
  OR2_X1 U2452 ( .A1(n2535), .A2(n2536), .ZN(n2067) );
  AND2_X1 U2453 ( .A1(n2051), .A2(n2050), .ZN(n2536) );
  AND2_X1 U2454 ( .A1(n2048), .A2(n2537), .ZN(n2535) );
  OR2_X1 U2455 ( .A1(n2051), .A2(n2050), .ZN(n2537) );
  OR2_X1 U2456 ( .A1(n2538), .A2(n2539), .ZN(n2050) );
  AND2_X1 U2457 ( .A1(n2039), .A2(n2038), .ZN(n2539) );
  AND2_X1 U2458 ( .A1(n2036), .A2(n2540), .ZN(n2538) );
  OR2_X1 U2459 ( .A1(n2039), .A2(n2038), .ZN(n2540) );
  OR2_X1 U2460 ( .A1(n2541), .A2(n2542), .ZN(n2038) );
  AND2_X1 U2461 ( .A1(n2022), .A2(n2021), .ZN(n2542) );
  AND2_X1 U2462 ( .A1(n2019), .A2(n2543), .ZN(n2541) );
  OR2_X1 U2463 ( .A1(n2022), .A2(n2021), .ZN(n2543) );
  OR2_X1 U2464 ( .A1(n2544), .A2(n2545), .ZN(n2021) );
  AND2_X1 U2465 ( .A1(n2010), .A2(n2009), .ZN(n2545) );
  AND2_X1 U2466 ( .A1(n2007), .A2(n2546), .ZN(n2544) );
  OR2_X1 U2467 ( .A1(n2010), .A2(n2009), .ZN(n2546) );
  OR2_X1 U2468 ( .A1(n2547), .A2(n2548), .ZN(n2009) );
  AND2_X1 U2469 ( .A1(n1990), .A2(n1993), .ZN(n2548) );
  AND2_X1 U2470 ( .A1(n1992), .A2(n2549), .ZN(n2547) );
  OR2_X1 U2471 ( .A1(n1990), .A2(n1993), .ZN(n2549) );
  OR2_X1 U2472 ( .A1(n2003), .A2(n1969), .ZN(n1993) );
  OR2_X1 U2473 ( .A1(n1974), .A2(n2236), .ZN(n1990) );
  OR2_X1 U2474 ( .A1(n1969), .A2(n2550), .ZN(n2236) );
  INV_X1 U2475 ( .A(n2551), .ZN(n1992) );
  OR2_X1 U2476 ( .A1(n2552), .A2(n2553), .ZN(n2551) );
  AND2_X1 U2477 ( .A1(b_14_), .A2(n2554), .ZN(n2553) );
  OR2_X1 U2478 ( .A1(n2555), .A2(n1980), .ZN(n2554) );
  AND2_X1 U2479 ( .A1(a_14_), .A2(n2002), .ZN(n2555) );
  AND2_X1 U2480 ( .A1(b_13_), .A2(n2556), .ZN(n2552) );
  OR2_X1 U2481 ( .A1(n2557), .A2(n1983), .ZN(n2556) );
  AND2_X1 U2482 ( .A1(a_15_), .A2(n1974), .ZN(n2557) );
  OR2_X1 U2483 ( .A1(n1969), .A2(n2231), .ZN(n2010) );
  XNOR2_X1 U2484 ( .A(n2558), .B(n2559), .ZN(n2007) );
  XNOR2_X1 U2485 ( .A(n2560), .B(n2561), .ZN(n2559) );
  OR2_X1 U2486 ( .A1(n1969), .A2(n2032), .ZN(n2022) );
  XOR2_X1 U2487 ( .A(n2562), .B(n2563), .Z(n2019) );
  XOR2_X1 U2488 ( .A(n2564), .B(n2565), .Z(n2563) );
  OR2_X1 U2489 ( .A1(n1969), .A2(n2225), .ZN(n2039) );
  XOR2_X1 U2490 ( .A(n2566), .B(n2567), .Z(n2036) );
  XOR2_X1 U2491 ( .A(n2568), .B(n2569), .Z(n2567) );
  OR2_X1 U2492 ( .A1(n1969), .A2(n2061), .ZN(n2051) );
  XOR2_X1 U2493 ( .A(n2570), .B(n2571), .Z(n2048) );
  XOR2_X1 U2494 ( .A(n2572), .B(n2573), .Z(n2571) );
  OR2_X1 U2495 ( .A1(n1969), .A2(n2219), .ZN(n2068) );
  XOR2_X1 U2496 ( .A(n2574), .B(n2575), .Z(n2065) );
  XOR2_X1 U2497 ( .A(n2576), .B(n2577), .Z(n2575) );
  OR2_X1 U2498 ( .A1(n1969), .A2(n2090), .ZN(n2080) );
  XOR2_X1 U2499 ( .A(n2578), .B(n2579), .Z(n2077) );
  XOR2_X1 U2500 ( .A(n2580), .B(n2581), .Z(n2579) );
  OR2_X1 U2501 ( .A1(n1969), .A2(n2213), .ZN(n2097) );
  XOR2_X1 U2502 ( .A(n2582), .B(n2583), .Z(n2094) );
  XOR2_X1 U2503 ( .A(n2584), .B(n2585), .Z(n2583) );
  OR2_X1 U2504 ( .A1(n1969), .A2(n2119), .ZN(n2109) );
  XOR2_X1 U2505 ( .A(n2586), .B(n2587), .Z(n2106) );
  XOR2_X1 U2506 ( .A(n2588), .B(n2589), .Z(n2587) );
  OR2_X1 U2507 ( .A1(n1969), .A2(n2207), .ZN(n2126) );
  XOR2_X1 U2508 ( .A(n2590), .B(n2591), .Z(n2123) );
  XOR2_X1 U2509 ( .A(n2592), .B(n2593), .Z(n2591) );
  OR2_X1 U2510 ( .A1(n1969), .A2(n2158), .ZN(n2148) );
  XOR2_X1 U2511 ( .A(n2594), .B(n2595), .Z(n2145) );
  XOR2_X1 U2512 ( .A(n2596), .B(n2597), .Z(n2595) );
  OR2_X1 U2513 ( .A1(n1969), .A2(n2201), .ZN(n2165) );
  XOR2_X1 U2514 ( .A(n2598), .B(n2599), .Z(n2162) );
  XOR2_X1 U2515 ( .A(n2600), .B(n2601), .Z(n2599) );
  OR2_X1 U2516 ( .A1(n1969), .A2(n2187), .ZN(n2177) );
  XOR2_X1 U2517 ( .A(n2602), .B(n2603), .Z(n2174) );
  XOR2_X1 U2518 ( .A(n2604), .B(n2605), .Z(n2603) );
  OR2_X1 U2519 ( .A1(n1969), .A2(n2291), .ZN(n2194) );
  INV_X1 U2520 ( .A(b_15_), .ZN(n1969) );
  XOR2_X1 U2521 ( .A(n2606), .B(n2607), .Z(n2191) );
  XOR2_X1 U2522 ( .A(n2608), .B(n2609), .Z(n2607) );
  XOR2_X1 U2523 ( .A(n2256), .B(n2257), .Z(n2247) );
  OR2_X1 U2524 ( .A1(n2610), .A2(n2611), .ZN(n2257) );
  AND2_X1 U2525 ( .A1(n2612), .A2(n2613), .ZN(n2611) );
  AND2_X1 U2526 ( .A1(n2614), .A2(n2615), .ZN(n2610) );
  OR2_X1 U2527 ( .A1(n2612), .A2(n2613), .ZN(n2615) );
  XOR2_X1 U2528 ( .A(n2502), .B(n2616), .Z(n2256) );
  XOR2_X1 U2529 ( .A(n2501), .B(n2500), .Z(n2616) );
  OR2_X1 U2530 ( .A1(n2002), .A2(n2291), .ZN(n2500) );
  OR2_X1 U2531 ( .A1(n2617), .A2(n2618), .ZN(n2501) );
  AND2_X1 U2532 ( .A1(n2619), .A2(n2620), .ZN(n2618) );
  AND2_X1 U2533 ( .A1(n2621), .A2(n2622), .ZN(n2617) );
  OR2_X1 U2534 ( .A1(n2620), .A2(n2619), .ZN(n2622) );
  XOR2_X1 U2535 ( .A(n2623), .B(n2624), .Z(n2502) );
  XOR2_X1 U2536 ( .A(n2625), .B(n2626), .Z(n2624) );
  XNOR2_X1 U2537 ( .A(n2614), .B(n2627), .ZN(n2243) );
  XOR2_X1 U2538 ( .A(n2613), .B(n2612), .Z(n2627) );
  OR2_X1 U2539 ( .A1(n1974), .A2(n2291), .ZN(n2612) );
  OR2_X1 U2540 ( .A1(n2628), .A2(n2629), .ZN(n2613) );
  AND2_X1 U2541 ( .A1(n2609), .A2(n2608), .ZN(n2629) );
  AND2_X1 U2542 ( .A1(n2606), .A2(n2630), .ZN(n2628) );
  OR2_X1 U2543 ( .A1(n2608), .A2(n2609), .ZN(n2630) );
  OR2_X1 U2544 ( .A1(n1974), .A2(n2187), .ZN(n2609) );
  OR2_X1 U2545 ( .A1(n2631), .A2(n2632), .ZN(n2608) );
  AND2_X1 U2546 ( .A1(n2605), .A2(n2604), .ZN(n2632) );
  AND2_X1 U2547 ( .A1(n2602), .A2(n2633), .ZN(n2631) );
  OR2_X1 U2548 ( .A1(n2604), .A2(n2605), .ZN(n2633) );
  OR2_X1 U2549 ( .A1(n1974), .A2(n2201), .ZN(n2605) );
  OR2_X1 U2550 ( .A1(n2634), .A2(n2635), .ZN(n2604) );
  AND2_X1 U2551 ( .A1(n2601), .A2(n2600), .ZN(n2635) );
  AND2_X1 U2552 ( .A1(n2598), .A2(n2636), .ZN(n2634) );
  OR2_X1 U2553 ( .A1(n2600), .A2(n2601), .ZN(n2636) );
  OR2_X1 U2554 ( .A1(n1974), .A2(n2158), .ZN(n2601) );
  OR2_X1 U2555 ( .A1(n2637), .A2(n2638), .ZN(n2600) );
  AND2_X1 U2556 ( .A1(n2597), .A2(n2596), .ZN(n2638) );
  AND2_X1 U2557 ( .A1(n2594), .A2(n2639), .ZN(n2637) );
  OR2_X1 U2558 ( .A1(n2596), .A2(n2597), .ZN(n2639) );
  OR2_X1 U2559 ( .A1(n1974), .A2(n2207), .ZN(n2597) );
  OR2_X1 U2560 ( .A1(n2640), .A2(n2641), .ZN(n2596) );
  AND2_X1 U2561 ( .A1(n2593), .A2(n2592), .ZN(n2641) );
  AND2_X1 U2562 ( .A1(n2590), .A2(n2642), .ZN(n2640) );
  OR2_X1 U2563 ( .A1(n2592), .A2(n2593), .ZN(n2642) );
  OR2_X1 U2564 ( .A1(n1974), .A2(n2119), .ZN(n2593) );
  OR2_X1 U2565 ( .A1(n2643), .A2(n2644), .ZN(n2592) );
  AND2_X1 U2566 ( .A1(n2589), .A2(n2588), .ZN(n2644) );
  AND2_X1 U2567 ( .A1(n2586), .A2(n2645), .ZN(n2643) );
  OR2_X1 U2568 ( .A1(n2588), .A2(n2589), .ZN(n2645) );
  OR2_X1 U2569 ( .A1(n1974), .A2(n2213), .ZN(n2589) );
  OR2_X1 U2570 ( .A1(n2646), .A2(n2647), .ZN(n2588) );
  AND2_X1 U2571 ( .A1(n2585), .A2(n2584), .ZN(n2647) );
  AND2_X1 U2572 ( .A1(n2582), .A2(n2648), .ZN(n2646) );
  OR2_X1 U2573 ( .A1(n2584), .A2(n2585), .ZN(n2648) );
  OR2_X1 U2574 ( .A1(n1974), .A2(n2090), .ZN(n2585) );
  OR2_X1 U2575 ( .A1(n2649), .A2(n2650), .ZN(n2584) );
  AND2_X1 U2576 ( .A1(n2581), .A2(n2580), .ZN(n2650) );
  AND2_X1 U2577 ( .A1(n2578), .A2(n2651), .ZN(n2649) );
  OR2_X1 U2578 ( .A1(n2580), .A2(n2581), .ZN(n2651) );
  OR2_X1 U2579 ( .A1(n1974), .A2(n2219), .ZN(n2581) );
  OR2_X1 U2580 ( .A1(n2652), .A2(n2653), .ZN(n2580) );
  AND2_X1 U2581 ( .A1(n2577), .A2(n2576), .ZN(n2653) );
  AND2_X1 U2582 ( .A1(n2574), .A2(n2654), .ZN(n2652) );
  OR2_X1 U2583 ( .A1(n2576), .A2(n2577), .ZN(n2654) );
  OR2_X1 U2584 ( .A1(n1974), .A2(n2061), .ZN(n2577) );
  OR2_X1 U2585 ( .A1(n2655), .A2(n2656), .ZN(n2576) );
  AND2_X1 U2586 ( .A1(n2573), .A2(n2572), .ZN(n2656) );
  AND2_X1 U2587 ( .A1(n2570), .A2(n2657), .ZN(n2655) );
  OR2_X1 U2588 ( .A1(n2572), .A2(n2573), .ZN(n2657) );
  OR2_X1 U2589 ( .A1(n1974), .A2(n2225), .ZN(n2573) );
  OR2_X1 U2590 ( .A1(n2658), .A2(n2659), .ZN(n2572) );
  AND2_X1 U2591 ( .A1(n2569), .A2(n2568), .ZN(n2659) );
  AND2_X1 U2592 ( .A1(n2566), .A2(n2660), .ZN(n2658) );
  OR2_X1 U2593 ( .A1(n2568), .A2(n2569), .ZN(n2660) );
  OR2_X1 U2594 ( .A1(n1974), .A2(n2032), .ZN(n2569) );
  OR2_X1 U2595 ( .A1(n2661), .A2(n2662), .ZN(n2568) );
  AND2_X1 U2596 ( .A1(n2565), .A2(n2564), .ZN(n2662) );
  AND2_X1 U2597 ( .A1(n2562), .A2(n2663), .ZN(n2661) );
  OR2_X1 U2598 ( .A1(n2564), .A2(n2565), .ZN(n2663) );
  OR2_X1 U2599 ( .A1(n1974), .A2(n2231), .ZN(n2565) );
  OR2_X1 U2600 ( .A1(n2664), .A2(n2665), .ZN(n2564) );
  AND2_X1 U2601 ( .A1(n2558), .A2(n2561), .ZN(n2665) );
  AND2_X1 U2602 ( .A1(n2560), .A2(n2666), .ZN(n2664) );
  OR2_X1 U2603 ( .A1(n2561), .A2(n2558), .ZN(n2666) );
  OR2_X1 U2604 ( .A1(n1974), .A2(n2003), .ZN(n2558) );
  OR3_X1 U2605 ( .A1(n2002), .A2(n1974), .A3(n2550), .ZN(n2561) );
  INV_X1 U2606 ( .A(b_14_), .ZN(n1974) );
  INV_X1 U2607 ( .A(n2667), .ZN(n2560) );
  OR2_X1 U2608 ( .A1(n2668), .A2(n2669), .ZN(n2667) );
  AND2_X1 U2609 ( .A1(b_13_), .A2(n2670), .ZN(n2669) );
  OR2_X1 U2610 ( .A1(n2671), .A2(n1980), .ZN(n2670) );
  AND2_X1 U2611 ( .A1(a_14_), .A2(n2232), .ZN(n2671) );
  AND2_X1 U2612 ( .A1(b_12_), .A2(n2672), .ZN(n2668) );
  OR2_X1 U2613 ( .A1(n2673), .A2(n1983), .ZN(n2672) );
  AND2_X1 U2614 ( .A1(a_15_), .A2(n2002), .ZN(n2673) );
  XNOR2_X1 U2615 ( .A(n1999), .B(n2674), .ZN(n2562) );
  XNOR2_X1 U2616 ( .A(n2675), .B(n2676), .ZN(n2674) );
  XOR2_X1 U2617 ( .A(n2677), .B(n2678), .Z(n2566) );
  XOR2_X1 U2618 ( .A(n2679), .B(n2680), .Z(n2678) );
  XOR2_X1 U2619 ( .A(n2681), .B(n2682), .Z(n2570) );
  XOR2_X1 U2620 ( .A(n2683), .B(n2684), .Z(n2682) );
  XOR2_X1 U2621 ( .A(n2685), .B(n2686), .Z(n2574) );
  XOR2_X1 U2622 ( .A(n2687), .B(n2688), .Z(n2686) );
  XOR2_X1 U2623 ( .A(n2689), .B(n2690), .Z(n2578) );
  XOR2_X1 U2624 ( .A(n2691), .B(n2692), .Z(n2690) );
  XOR2_X1 U2625 ( .A(n2693), .B(n2694), .Z(n2582) );
  XOR2_X1 U2626 ( .A(n2695), .B(n2696), .Z(n2694) );
  XOR2_X1 U2627 ( .A(n2697), .B(n2698), .Z(n2586) );
  XOR2_X1 U2628 ( .A(n2699), .B(n2700), .Z(n2698) );
  XOR2_X1 U2629 ( .A(n2701), .B(n2702), .Z(n2590) );
  XOR2_X1 U2630 ( .A(n2703), .B(n2704), .Z(n2702) );
  XOR2_X1 U2631 ( .A(n2705), .B(n2706), .Z(n2594) );
  XOR2_X1 U2632 ( .A(n2707), .B(n2708), .Z(n2706) );
  XOR2_X1 U2633 ( .A(n2709), .B(n2710), .Z(n2598) );
  XOR2_X1 U2634 ( .A(n2711), .B(n2712), .Z(n2710) );
  XOR2_X1 U2635 ( .A(n2713), .B(n2714), .Z(n2602) );
  XOR2_X1 U2636 ( .A(n2715), .B(n2716), .Z(n2714) );
  XOR2_X1 U2637 ( .A(n2717), .B(n2718), .Z(n2606) );
  XOR2_X1 U2638 ( .A(n2719), .B(n2720), .Z(n2718) );
  XOR2_X1 U2639 ( .A(n2621), .B(n2721), .Z(n2614) );
  XOR2_X1 U2640 ( .A(n2620), .B(n2619), .Z(n2721) );
  OR2_X1 U2641 ( .A1(n2002), .A2(n2187), .ZN(n2619) );
  OR2_X1 U2642 ( .A1(n2722), .A2(n2723), .ZN(n2620) );
  AND2_X1 U2643 ( .A1(n2720), .A2(n2719), .ZN(n2723) );
  AND2_X1 U2644 ( .A1(n2717), .A2(n2724), .ZN(n2722) );
  OR2_X1 U2645 ( .A1(n2719), .A2(n2720), .ZN(n2724) );
  OR2_X1 U2646 ( .A1(n2002), .A2(n2201), .ZN(n2720) );
  OR2_X1 U2647 ( .A1(n2725), .A2(n2726), .ZN(n2719) );
  AND2_X1 U2648 ( .A1(n2716), .A2(n2715), .ZN(n2726) );
  AND2_X1 U2649 ( .A1(n2713), .A2(n2727), .ZN(n2725) );
  OR2_X1 U2650 ( .A1(n2715), .A2(n2716), .ZN(n2727) );
  OR2_X1 U2651 ( .A1(n2002), .A2(n2158), .ZN(n2716) );
  OR2_X1 U2652 ( .A1(n2728), .A2(n2729), .ZN(n2715) );
  AND2_X1 U2653 ( .A1(n2712), .A2(n2711), .ZN(n2729) );
  AND2_X1 U2654 ( .A1(n2709), .A2(n2730), .ZN(n2728) );
  OR2_X1 U2655 ( .A1(n2711), .A2(n2712), .ZN(n2730) );
  OR2_X1 U2656 ( .A1(n2002), .A2(n2207), .ZN(n2712) );
  OR2_X1 U2657 ( .A1(n2731), .A2(n2732), .ZN(n2711) );
  AND2_X1 U2658 ( .A1(n2708), .A2(n2707), .ZN(n2732) );
  AND2_X1 U2659 ( .A1(n2705), .A2(n2733), .ZN(n2731) );
  OR2_X1 U2660 ( .A1(n2707), .A2(n2708), .ZN(n2733) );
  OR2_X1 U2661 ( .A1(n2002), .A2(n2119), .ZN(n2708) );
  OR2_X1 U2662 ( .A1(n2734), .A2(n2735), .ZN(n2707) );
  AND2_X1 U2663 ( .A1(n2704), .A2(n2703), .ZN(n2735) );
  AND2_X1 U2664 ( .A1(n2701), .A2(n2736), .ZN(n2734) );
  OR2_X1 U2665 ( .A1(n2703), .A2(n2704), .ZN(n2736) );
  OR2_X1 U2666 ( .A1(n2002), .A2(n2213), .ZN(n2704) );
  OR2_X1 U2667 ( .A1(n2737), .A2(n2738), .ZN(n2703) );
  AND2_X1 U2668 ( .A1(n2700), .A2(n2699), .ZN(n2738) );
  AND2_X1 U2669 ( .A1(n2697), .A2(n2739), .ZN(n2737) );
  OR2_X1 U2670 ( .A1(n2699), .A2(n2700), .ZN(n2739) );
  OR2_X1 U2671 ( .A1(n2002), .A2(n2090), .ZN(n2700) );
  OR2_X1 U2672 ( .A1(n2740), .A2(n2741), .ZN(n2699) );
  AND2_X1 U2673 ( .A1(n2696), .A2(n2695), .ZN(n2741) );
  AND2_X1 U2674 ( .A1(n2693), .A2(n2742), .ZN(n2740) );
  OR2_X1 U2675 ( .A1(n2695), .A2(n2696), .ZN(n2742) );
  OR2_X1 U2676 ( .A1(n2002), .A2(n2219), .ZN(n2696) );
  OR2_X1 U2677 ( .A1(n2743), .A2(n2744), .ZN(n2695) );
  AND2_X1 U2678 ( .A1(n2692), .A2(n2691), .ZN(n2744) );
  AND2_X1 U2679 ( .A1(n2689), .A2(n2745), .ZN(n2743) );
  OR2_X1 U2680 ( .A1(n2691), .A2(n2692), .ZN(n2745) );
  OR2_X1 U2681 ( .A1(n2002), .A2(n2061), .ZN(n2692) );
  OR2_X1 U2682 ( .A1(n2746), .A2(n2747), .ZN(n2691) );
  AND2_X1 U2683 ( .A1(n2688), .A2(n2687), .ZN(n2747) );
  AND2_X1 U2684 ( .A1(n2685), .A2(n2748), .ZN(n2746) );
  OR2_X1 U2685 ( .A1(n2687), .A2(n2688), .ZN(n2748) );
  OR2_X1 U2686 ( .A1(n2002), .A2(n2225), .ZN(n2688) );
  OR2_X1 U2687 ( .A1(n2749), .A2(n2750), .ZN(n2687) );
  AND2_X1 U2688 ( .A1(n2684), .A2(n2683), .ZN(n2750) );
  AND2_X1 U2689 ( .A1(n2681), .A2(n2751), .ZN(n2749) );
  OR2_X1 U2690 ( .A1(n2683), .A2(n2684), .ZN(n2751) );
  OR2_X1 U2691 ( .A1(n2002), .A2(n2032), .ZN(n2684) );
  OR2_X1 U2692 ( .A1(n2752), .A2(n2753), .ZN(n2683) );
  AND2_X1 U2693 ( .A1(n2680), .A2(n2679), .ZN(n2753) );
  AND2_X1 U2694 ( .A1(n2677), .A2(n2754), .ZN(n2752) );
  OR2_X1 U2695 ( .A1(n2679), .A2(n2680), .ZN(n2754) );
  OR2_X1 U2696 ( .A1(n2002), .A2(n2231), .ZN(n2680) );
  OR2_X1 U2697 ( .A1(n2755), .A2(n2756), .ZN(n2679) );
  AND2_X1 U2698 ( .A1(n1999), .A2(n2676), .ZN(n2756) );
  AND2_X1 U2699 ( .A1(n2675), .A2(n2757), .ZN(n2755) );
  OR2_X1 U2700 ( .A1(n2676), .A2(n1999), .ZN(n2757) );
  OR2_X1 U2701 ( .A1(n2002), .A2(n2003), .ZN(n1999) );
  OR3_X1 U2702 ( .A1(n2002), .A2(n2550), .A3(n2232), .ZN(n2676) );
  INV_X1 U2703 ( .A(b_13_), .ZN(n2002) );
  INV_X1 U2704 ( .A(n2758), .ZN(n2675) );
  OR2_X1 U2705 ( .A1(n2759), .A2(n2760), .ZN(n2758) );
  AND2_X1 U2706 ( .A1(b_12_), .A2(n2761), .ZN(n2760) );
  OR2_X1 U2707 ( .A1(n2762), .A2(n1980), .ZN(n2761) );
  AND2_X1 U2708 ( .A1(a_14_), .A2(n2031), .ZN(n2762) );
  AND2_X1 U2709 ( .A1(b_11_), .A2(n2763), .ZN(n2759) );
  OR2_X1 U2710 ( .A1(n2764), .A2(n1983), .ZN(n2763) );
  AND2_X1 U2711 ( .A1(a_15_), .A2(n2232), .ZN(n2764) );
  XNOR2_X1 U2712 ( .A(n2765), .B(n2766), .ZN(n2677) );
  XNOR2_X1 U2713 ( .A(n2767), .B(n2768), .ZN(n2766) );
  XOR2_X1 U2714 ( .A(n2769), .B(n2770), .Z(n2681) );
  XNOR2_X1 U2715 ( .A(n2771), .B(n2014), .ZN(n2770) );
  XOR2_X1 U2716 ( .A(n2772), .B(n2773), .Z(n2685) );
  XOR2_X1 U2717 ( .A(n2774), .B(n2775), .Z(n2773) );
  XOR2_X1 U2718 ( .A(n2776), .B(n2777), .Z(n2689) );
  XOR2_X1 U2719 ( .A(n2778), .B(n2779), .Z(n2777) );
  XOR2_X1 U2720 ( .A(n2780), .B(n2781), .Z(n2693) );
  XOR2_X1 U2721 ( .A(n2782), .B(n2783), .Z(n2781) );
  XOR2_X1 U2722 ( .A(n2784), .B(n2785), .Z(n2697) );
  XOR2_X1 U2723 ( .A(n2786), .B(n2787), .Z(n2785) );
  XOR2_X1 U2724 ( .A(n2788), .B(n2789), .Z(n2701) );
  XOR2_X1 U2725 ( .A(n2790), .B(n2791), .Z(n2789) );
  XOR2_X1 U2726 ( .A(n2792), .B(n2793), .Z(n2705) );
  XOR2_X1 U2727 ( .A(n2794), .B(n2795), .Z(n2793) );
  XOR2_X1 U2728 ( .A(n2796), .B(n2797), .Z(n2709) );
  XOR2_X1 U2729 ( .A(n2798), .B(n2799), .Z(n2797) );
  XOR2_X1 U2730 ( .A(n2800), .B(n2801), .Z(n2713) );
  XOR2_X1 U2731 ( .A(n2802), .B(n2803), .Z(n2801) );
  XOR2_X1 U2732 ( .A(n2804), .B(n2805), .Z(n2717) );
  XOR2_X1 U2733 ( .A(n2806), .B(n2807), .Z(n2805) );
  XOR2_X1 U2734 ( .A(n2808), .B(n2809), .Z(n2621) );
  XOR2_X1 U2735 ( .A(n2810), .B(n2811), .Z(n2809) );
  XNOR2_X1 U2736 ( .A(n2274), .B(n2489), .ZN(n2264) );
  OR2_X1 U2737 ( .A1(n2812), .A2(n2813), .ZN(n2489) );
  AND2_X1 U2738 ( .A1(n2507), .A2(n2506), .ZN(n2813) );
  AND2_X1 U2739 ( .A1(n2504), .A2(n2814), .ZN(n2812) );
  OR2_X1 U2740 ( .A1(n2506), .A2(n2507), .ZN(n2814) );
  OR2_X1 U2741 ( .A1(n2232), .A2(n2291), .ZN(n2507) );
  OR2_X1 U2742 ( .A1(n2815), .A2(n2816), .ZN(n2506) );
  AND2_X1 U2743 ( .A1(n2626), .A2(n2625), .ZN(n2816) );
  AND2_X1 U2744 ( .A1(n2623), .A2(n2817), .ZN(n2815) );
  OR2_X1 U2745 ( .A1(n2625), .A2(n2626), .ZN(n2817) );
  OR2_X1 U2746 ( .A1(n2232), .A2(n2187), .ZN(n2626) );
  OR2_X1 U2747 ( .A1(n2818), .A2(n2819), .ZN(n2625) );
  AND2_X1 U2748 ( .A1(n2811), .A2(n2810), .ZN(n2819) );
  AND2_X1 U2749 ( .A1(n2808), .A2(n2820), .ZN(n2818) );
  OR2_X1 U2750 ( .A1(n2810), .A2(n2811), .ZN(n2820) );
  OR2_X1 U2751 ( .A1(n2232), .A2(n2201), .ZN(n2811) );
  OR2_X1 U2752 ( .A1(n2821), .A2(n2822), .ZN(n2810) );
  AND2_X1 U2753 ( .A1(n2807), .A2(n2806), .ZN(n2822) );
  AND2_X1 U2754 ( .A1(n2804), .A2(n2823), .ZN(n2821) );
  OR2_X1 U2755 ( .A1(n2806), .A2(n2807), .ZN(n2823) );
  OR2_X1 U2756 ( .A1(n2232), .A2(n2158), .ZN(n2807) );
  OR2_X1 U2757 ( .A1(n2824), .A2(n2825), .ZN(n2806) );
  AND2_X1 U2758 ( .A1(n2803), .A2(n2802), .ZN(n2825) );
  AND2_X1 U2759 ( .A1(n2800), .A2(n2826), .ZN(n2824) );
  OR2_X1 U2760 ( .A1(n2802), .A2(n2803), .ZN(n2826) );
  OR2_X1 U2761 ( .A1(n2232), .A2(n2207), .ZN(n2803) );
  OR2_X1 U2762 ( .A1(n2827), .A2(n2828), .ZN(n2802) );
  AND2_X1 U2763 ( .A1(n2799), .A2(n2798), .ZN(n2828) );
  AND2_X1 U2764 ( .A1(n2796), .A2(n2829), .ZN(n2827) );
  OR2_X1 U2765 ( .A1(n2798), .A2(n2799), .ZN(n2829) );
  OR2_X1 U2766 ( .A1(n2232), .A2(n2119), .ZN(n2799) );
  OR2_X1 U2767 ( .A1(n2830), .A2(n2831), .ZN(n2798) );
  AND2_X1 U2768 ( .A1(n2795), .A2(n2794), .ZN(n2831) );
  AND2_X1 U2769 ( .A1(n2792), .A2(n2832), .ZN(n2830) );
  OR2_X1 U2770 ( .A1(n2794), .A2(n2795), .ZN(n2832) );
  OR2_X1 U2771 ( .A1(n2232), .A2(n2213), .ZN(n2795) );
  OR2_X1 U2772 ( .A1(n2833), .A2(n2834), .ZN(n2794) );
  AND2_X1 U2773 ( .A1(n2791), .A2(n2790), .ZN(n2834) );
  AND2_X1 U2774 ( .A1(n2788), .A2(n2835), .ZN(n2833) );
  OR2_X1 U2775 ( .A1(n2790), .A2(n2791), .ZN(n2835) );
  OR2_X1 U2776 ( .A1(n2232), .A2(n2090), .ZN(n2791) );
  OR2_X1 U2777 ( .A1(n2836), .A2(n2837), .ZN(n2790) );
  AND2_X1 U2778 ( .A1(n2787), .A2(n2786), .ZN(n2837) );
  AND2_X1 U2779 ( .A1(n2784), .A2(n2838), .ZN(n2836) );
  OR2_X1 U2780 ( .A1(n2786), .A2(n2787), .ZN(n2838) );
  OR2_X1 U2781 ( .A1(n2232), .A2(n2219), .ZN(n2787) );
  OR2_X1 U2782 ( .A1(n2839), .A2(n2840), .ZN(n2786) );
  AND2_X1 U2783 ( .A1(n2783), .A2(n2782), .ZN(n2840) );
  AND2_X1 U2784 ( .A1(n2780), .A2(n2841), .ZN(n2839) );
  OR2_X1 U2785 ( .A1(n2782), .A2(n2783), .ZN(n2841) );
  OR2_X1 U2786 ( .A1(n2232), .A2(n2061), .ZN(n2783) );
  OR2_X1 U2787 ( .A1(n2842), .A2(n2843), .ZN(n2782) );
  AND2_X1 U2788 ( .A1(n2779), .A2(n2778), .ZN(n2843) );
  AND2_X1 U2789 ( .A1(n2776), .A2(n2844), .ZN(n2842) );
  OR2_X1 U2790 ( .A1(n2778), .A2(n2779), .ZN(n2844) );
  OR2_X1 U2791 ( .A1(n2232), .A2(n2225), .ZN(n2779) );
  OR2_X1 U2792 ( .A1(n2845), .A2(n2846), .ZN(n2778) );
  AND2_X1 U2793 ( .A1(n2775), .A2(n2774), .ZN(n2846) );
  AND2_X1 U2794 ( .A1(n2772), .A2(n2847), .ZN(n2845) );
  OR2_X1 U2795 ( .A1(n2774), .A2(n2775), .ZN(n2847) );
  OR2_X1 U2796 ( .A1(n2232), .A2(n2032), .ZN(n2775) );
  OR2_X1 U2797 ( .A1(n2848), .A2(n2849), .ZN(n2774) );
  AND2_X1 U2798 ( .A1(n2233), .A2(n2771), .ZN(n2849) );
  AND2_X1 U2799 ( .A1(n2769), .A2(n2850), .ZN(n2848) );
  OR2_X1 U2800 ( .A1(n2771), .A2(n2233), .ZN(n2850) );
  INV_X1 U2801 ( .A(n2014), .ZN(n2233) );
  AND2_X1 U2802 ( .A1(a_12_), .A2(b_12_), .ZN(n2014) );
  OR2_X1 U2803 ( .A1(n2851), .A2(n2852), .ZN(n2771) );
  AND2_X1 U2804 ( .A1(n2765), .A2(n2768), .ZN(n2852) );
  AND2_X1 U2805 ( .A1(n2767), .A2(n2853), .ZN(n2851) );
  OR2_X1 U2806 ( .A1(n2768), .A2(n2765), .ZN(n2853) );
  OR2_X1 U2807 ( .A1(n2003), .A2(n2232), .ZN(n2765) );
  OR3_X1 U2808 ( .A1(n2550), .A2(n2232), .A3(n2031), .ZN(n2768) );
  INV_X1 U2809 ( .A(b_12_), .ZN(n2232) );
  INV_X1 U2810 ( .A(n2854), .ZN(n2767) );
  OR2_X1 U2811 ( .A1(n2855), .A2(n2856), .ZN(n2854) );
  AND2_X1 U2812 ( .A1(b_11_), .A2(n2857), .ZN(n2856) );
  OR2_X1 U2813 ( .A1(n2858), .A2(n1980), .ZN(n2857) );
  AND2_X1 U2814 ( .A1(a_14_), .A2(n2226), .ZN(n2858) );
  AND2_X1 U2815 ( .A1(b_10_), .A2(n2859), .ZN(n2855) );
  OR2_X1 U2816 ( .A1(n2860), .A2(n1983), .ZN(n2859) );
  AND2_X1 U2817 ( .A1(a_15_), .A2(n2031), .ZN(n2860) );
  XNOR2_X1 U2818 ( .A(n2861), .B(n2862), .ZN(n2769) );
  XNOR2_X1 U2819 ( .A(n2863), .B(n2864), .ZN(n2862) );
  XNOR2_X1 U2820 ( .A(n2865), .B(n2866), .ZN(n2772) );
  XNOR2_X1 U2821 ( .A(n2867), .B(n2868), .ZN(n2865) );
  XOR2_X1 U2822 ( .A(n2869), .B(n2870), .Z(n2776) );
  XOR2_X1 U2823 ( .A(n2871), .B(n2029), .Z(n2870) );
  XOR2_X1 U2824 ( .A(n2872), .B(n2873), .Z(n2780) );
  XOR2_X1 U2825 ( .A(n2874), .B(n2875), .Z(n2873) );
  XOR2_X1 U2826 ( .A(n2876), .B(n2877), .Z(n2784) );
  XOR2_X1 U2827 ( .A(n2878), .B(n2879), .Z(n2877) );
  XOR2_X1 U2828 ( .A(n2880), .B(n2881), .Z(n2788) );
  XOR2_X1 U2829 ( .A(n2882), .B(n2883), .Z(n2881) );
  XOR2_X1 U2830 ( .A(n2884), .B(n2885), .Z(n2792) );
  XOR2_X1 U2831 ( .A(n2886), .B(n2887), .Z(n2885) );
  XOR2_X1 U2832 ( .A(n2888), .B(n2889), .Z(n2796) );
  XOR2_X1 U2833 ( .A(n2890), .B(n2891), .Z(n2889) );
  XOR2_X1 U2834 ( .A(n2892), .B(n2893), .Z(n2800) );
  XOR2_X1 U2835 ( .A(n2894), .B(n2895), .Z(n2893) );
  XOR2_X1 U2836 ( .A(n2896), .B(n2897), .Z(n2804) );
  XOR2_X1 U2837 ( .A(n2898), .B(n2899), .Z(n2897) );
  XOR2_X1 U2838 ( .A(n2900), .B(n2901), .Z(n2808) );
  XOR2_X1 U2839 ( .A(n2902), .B(n2903), .Z(n2901) );
  XOR2_X1 U2840 ( .A(n2904), .B(n2905), .Z(n2623) );
  XOR2_X1 U2841 ( .A(n2906), .B(n2907), .Z(n2905) );
  XOR2_X1 U2842 ( .A(n2908), .B(n2909), .Z(n2504) );
  XOR2_X1 U2843 ( .A(n2910), .B(n2911), .Z(n2909) );
  XNOR2_X1 U2844 ( .A(n2912), .B(n2913), .ZN(n2274) );
  XOR2_X1 U2845 ( .A(n2914), .B(n2915), .Z(n2913) );
  XNOR2_X1 U2846 ( .A(n2284), .B(n2487), .ZN(n2272) );
  OR2_X1 U2847 ( .A1(n2916), .A2(n2917), .ZN(n2487) );
  AND2_X1 U2848 ( .A1(n2915), .A2(n2914), .ZN(n2917) );
  AND2_X1 U2849 ( .A1(n2912), .A2(n2918), .ZN(n2916) );
  OR2_X1 U2850 ( .A1(n2914), .A2(n2915), .ZN(n2918) );
  OR2_X1 U2851 ( .A1(n2031), .A2(n2291), .ZN(n2915) );
  OR2_X1 U2852 ( .A1(n2919), .A2(n2920), .ZN(n2914) );
  AND2_X1 U2853 ( .A1(n2911), .A2(n2910), .ZN(n2920) );
  AND2_X1 U2854 ( .A1(n2908), .A2(n2921), .ZN(n2919) );
  OR2_X1 U2855 ( .A1(n2910), .A2(n2911), .ZN(n2921) );
  OR2_X1 U2856 ( .A1(n2031), .A2(n2187), .ZN(n2911) );
  OR2_X1 U2857 ( .A1(n2922), .A2(n2923), .ZN(n2910) );
  AND2_X1 U2858 ( .A1(n2907), .A2(n2906), .ZN(n2923) );
  AND2_X1 U2859 ( .A1(n2904), .A2(n2924), .ZN(n2922) );
  OR2_X1 U2860 ( .A1(n2906), .A2(n2907), .ZN(n2924) );
  OR2_X1 U2861 ( .A1(n2031), .A2(n2201), .ZN(n2907) );
  OR2_X1 U2862 ( .A1(n2925), .A2(n2926), .ZN(n2906) );
  AND2_X1 U2863 ( .A1(n2903), .A2(n2902), .ZN(n2926) );
  AND2_X1 U2864 ( .A1(n2900), .A2(n2927), .ZN(n2925) );
  OR2_X1 U2865 ( .A1(n2902), .A2(n2903), .ZN(n2927) );
  OR2_X1 U2866 ( .A1(n2031), .A2(n2158), .ZN(n2903) );
  OR2_X1 U2867 ( .A1(n2928), .A2(n2929), .ZN(n2902) );
  AND2_X1 U2868 ( .A1(n2899), .A2(n2898), .ZN(n2929) );
  AND2_X1 U2869 ( .A1(n2896), .A2(n2930), .ZN(n2928) );
  OR2_X1 U2870 ( .A1(n2898), .A2(n2899), .ZN(n2930) );
  OR2_X1 U2871 ( .A1(n2031), .A2(n2207), .ZN(n2899) );
  OR2_X1 U2872 ( .A1(n2931), .A2(n2932), .ZN(n2898) );
  AND2_X1 U2873 ( .A1(n2895), .A2(n2894), .ZN(n2932) );
  AND2_X1 U2874 ( .A1(n2892), .A2(n2933), .ZN(n2931) );
  OR2_X1 U2875 ( .A1(n2894), .A2(n2895), .ZN(n2933) );
  OR2_X1 U2876 ( .A1(n2031), .A2(n2119), .ZN(n2895) );
  OR2_X1 U2877 ( .A1(n2934), .A2(n2935), .ZN(n2894) );
  AND2_X1 U2878 ( .A1(n2891), .A2(n2890), .ZN(n2935) );
  AND2_X1 U2879 ( .A1(n2888), .A2(n2936), .ZN(n2934) );
  OR2_X1 U2880 ( .A1(n2890), .A2(n2891), .ZN(n2936) );
  OR2_X1 U2881 ( .A1(n2031), .A2(n2213), .ZN(n2891) );
  OR2_X1 U2882 ( .A1(n2937), .A2(n2938), .ZN(n2890) );
  AND2_X1 U2883 ( .A1(n2887), .A2(n2886), .ZN(n2938) );
  AND2_X1 U2884 ( .A1(n2884), .A2(n2939), .ZN(n2937) );
  OR2_X1 U2885 ( .A1(n2886), .A2(n2887), .ZN(n2939) );
  OR2_X1 U2886 ( .A1(n2031), .A2(n2090), .ZN(n2887) );
  OR2_X1 U2887 ( .A1(n2940), .A2(n2941), .ZN(n2886) );
  AND2_X1 U2888 ( .A1(n2883), .A2(n2882), .ZN(n2941) );
  AND2_X1 U2889 ( .A1(n2880), .A2(n2942), .ZN(n2940) );
  OR2_X1 U2890 ( .A1(n2882), .A2(n2883), .ZN(n2942) );
  OR2_X1 U2891 ( .A1(n2031), .A2(n2219), .ZN(n2883) );
  OR2_X1 U2892 ( .A1(n2943), .A2(n2944), .ZN(n2882) );
  AND2_X1 U2893 ( .A1(n2879), .A2(n2878), .ZN(n2944) );
  AND2_X1 U2894 ( .A1(n2876), .A2(n2945), .ZN(n2943) );
  OR2_X1 U2895 ( .A1(n2878), .A2(n2879), .ZN(n2945) );
  OR2_X1 U2896 ( .A1(n2031), .A2(n2061), .ZN(n2879) );
  OR2_X1 U2897 ( .A1(n2946), .A2(n2947), .ZN(n2878) );
  AND2_X1 U2898 ( .A1(n2875), .A2(n2874), .ZN(n2947) );
  AND2_X1 U2899 ( .A1(n2872), .A2(n2948), .ZN(n2946) );
  OR2_X1 U2900 ( .A1(n2874), .A2(n2875), .ZN(n2948) );
  OR2_X1 U2901 ( .A1(n2031), .A2(n2225), .ZN(n2875) );
  OR2_X1 U2902 ( .A1(n2949), .A2(n2950), .ZN(n2874) );
  AND2_X1 U2903 ( .A1(n2029), .A2(n2871), .ZN(n2950) );
  AND2_X1 U2904 ( .A1(n2869), .A2(n2951), .ZN(n2949) );
  OR2_X1 U2905 ( .A1(n2871), .A2(n2029), .ZN(n2951) );
  OR2_X1 U2906 ( .A1(n2032), .A2(n2031), .ZN(n2029) );
  OR2_X1 U2907 ( .A1(n2952), .A2(n2953), .ZN(n2871) );
  AND2_X1 U2908 ( .A1(n2868), .A2(n2867), .ZN(n2953) );
  AND2_X1 U2909 ( .A1(n2866), .A2(n2954), .ZN(n2952) );
  OR2_X1 U2910 ( .A1(n2867), .A2(n2868), .ZN(n2954) );
  OR2_X1 U2911 ( .A1(n2231), .A2(n2031), .ZN(n2868) );
  OR2_X1 U2912 ( .A1(n2955), .A2(n2956), .ZN(n2867) );
  AND2_X1 U2913 ( .A1(n2861), .A2(n2864), .ZN(n2956) );
  AND2_X1 U2914 ( .A1(n2863), .A2(n2957), .ZN(n2955) );
  OR2_X1 U2915 ( .A1(n2864), .A2(n2861), .ZN(n2957) );
  OR2_X1 U2916 ( .A1(n2003), .A2(n2031), .ZN(n2861) );
  OR3_X1 U2917 ( .A1(n2550), .A2(n2031), .A3(n2226), .ZN(n2864) );
  INV_X1 U2918 ( .A(b_11_), .ZN(n2031) );
  INV_X1 U2919 ( .A(n2958), .ZN(n2863) );
  OR2_X1 U2920 ( .A1(n2959), .A2(n2960), .ZN(n2958) );
  AND2_X1 U2921 ( .A1(b_9_), .A2(n2961), .ZN(n2960) );
  OR2_X1 U2922 ( .A1(n2962), .A2(n1983), .ZN(n2961) );
  AND2_X1 U2923 ( .A1(a_15_), .A2(n2226), .ZN(n2962) );
  AND2_X1 U2924 ( .A1(b_10_), .A2(n2963), .ZN(n2959) );
  OR2_X1 U2925 ( .A1(n2964), .A2(n1980), .ZN(n2963) );
  AND2_X1 U2926 ( .A1(a_14_), .A2(n2060), .ZN(n2964) );
  XNOR2_X1 U2927 ( .A(n2965), .B(n2966), .ZN(n2866) );
  XNOR2_X1 U2928 ( .A(n2967), .B(n2968), .ZN(n2966) );
  XOR2_X1 U2929 ( .A(n2969), .B(n2970), .Z(n2869) );
  XOR2_X1 U2930 ( .A(n2971), .B(n2972), .Z(n2970) );
  XOR2_X1 U2931 ( .A(n2973), .B(n2974), .Z(n2872) );
  XOR2_X1 U2932 ( .A(n2975), .B(n2976), .Z(n2974) );
  XOR2_X1 U2933 ( .A(n2977), .B(n2978), .Z(n2876) );
  XNOR2_X1 U2934 ( .A(n2979), .B(n2044), .ZN(n2978) );
  XOR2_X1 U2935 ( .A(n2980), .B(n2981), .Z(n2880) );
  XOR2_X1 U2936 ( .A(n2982), .B(n2983), .Z(n2981) );
  XOR2_X1 U2937 ( .A(n2984), .B(n2985), .Z(n2884) );
  XOR2_X1 U2938 ( .A(n2986), .B(n2987), .Z(n2985) );
  XOR2_X1 U2939 ( .A(n2988), .B(n2989), .Z(n2888) );
  XOR2_X1 U2940 ( .A(n2990), .B(n2991), .Z(n2989) );
  XOR2_X1 U2941 ( .A(n2992), .B(n2993), .Z(n2892) );
  XOR2_X1 U2942 ( .A(n2994), .B(n2995), .Z(n2993) );
  XOR2_X1 U2943 ( .A(n2996), .B(n2997), .Z(n2896) );
  XOR2_X1 U2944 ( .A(n2998), .B(n2999), .Z(n2997) );
  XOR2_X1 U2945 ( .A(n3000), .B(n3001), .Z(n2900) );
  XOR2_X1 U2946 ( .A(n3002), .B(n3003), .Z(n3001) );
  XOR2_X1 U2947 ( .A(n3004), .B(n3005), .Z(n2904) );
  XOR2_X1 U2948 ( .A(n3006), .B(n3007), .Z(n3005) );
  XOR2_X1 U2949 ( .A(n3008), .B(n3009), .Z(n2908) );
  XOR2_X1 U2950 ( .A(n3010), .B(n3011), .Z(n3009) );
  XOR2_X1 U2951 ( .A(n3012), .B(n3013), .Z(n2912) );
  XOR2_X1 U2952 ( .A(n3014), .B(n3015), .Z(n3013) );
  XNOR2_X1 U2953 ( .A(n3016), .B(n3017), .ZN(n2284) );
  XOR2_X1 U2954 ( .A(n3018), .B(n3019), .Z(n3017) );
  XNOR2_X1 U2955 ( .A(n1922), .B(n2485), .ZN(n2282) );
  OR2_X1 U2956 ( .A1(n3020), .A2(n3021), .ZN(n2485) );
  AND2_X1 U2957 ( .A1(n3019), .A2(n3018), .ZN(n3021) );
  AND2_X1 U2958 ( .A1(n3016), .A2(n3022), .ZN(n3020) );
  OR2_X1 U2959 ( .A1(n3018), .A2(n3019), .ZN(n3022) );
  OR2_X1 U2960 ( .A1(n2226), .A2(n2291), .ZN(n3019) );
  OR2_X1 U2961 ( .A1(n3023), .A2(n3024), .ZN(n3018) );
  AND2_X1 U2962 ( .A1(n3015), .A2(n3014), .ZN(n3024) );
  AND2_X1 U2963 ( .A1(n3012), .A2(n3025), .ZN(n3023) );
  OR2_X1 U2964 ( .A1(n3014), .A2(n3015), .ZN(n3025) );
  OR2_X1 U2965 ( .A1(n2226), .A2(n2187), .ZN(n3015) );
  OR2_X1 U2966 ( .A1(n3026), .A2(n3027), .ZN(n3014) );
  AND2_X1 U2967 ( .A1(n3011), .A2(n3010), .ZN(n3027) );
  AND2_X1 U2968 ( .A1(n3008), .A2(n3028), .ZN(n3026) );
  OR2_X1 U2969 ( .A1(n3010), .A2(n3011), .ZN(n3028) );
  OR2_X1 U2970 ( .A1(n2226), .A2(n2201), .ZN(n3011) );
  OR2_X1 U2971 ( .A1(n3029), .A2(n3030), .ZN(n3010) );
  AND2_X1 U2972 ( .A1(n3004), .A2(n3007), .ZN(n3030) );
  AND2_X1 U2973 ( .A1(n3031), .A2(n3006), .ZN(n3029) );
  OR2_X1 U2974 ( .A1(n3032), .A2(n3033), .ZN(n3006) );
  AND2_X1 U2975 ( .A1(n3003), .A2(n3002), .ZN(n3033) );
  AND2_X1 U2976 ( .A1(n3000), .A2(n3034), .ZN(n3032) );
  OR2_X1 U2977 ( .A1(n3002), .A2(n3003), .ZN(n3034) );
  OR2_X1 U2978 ( .A1(n2226), .A2(n2207), .ZN(n3003) );
  OR2_X1 U2979 ( .A1(n3035), .A2(n3036), .ZN(n3002) );
  AND2_X1 U2980 ( .A1(n2996), .A2(n2999), .ZN(n3036) );
  AND2_X1 U2981 ( .A1(n3037), .A2(n2998), .ZN(n3035) );
  OR2_X1 U2982 ( .A1(n3038), .A2(n3039), .ZN(n2998) );
  AND2_X1 U2983 ( .A1(n2992), .A2(n2995), .ZN(n3039) );
  AND2_X1 U2984 ( .A1(n3040), .A2(n2994), .ZN(n3038) );
  OR2_X1 U2985 ( .A1(n3041), .A2(n3042), .ZN(n2994) );
  AND2_X1 U2986 ( .A1(n2988), .A2(n2991), .ZN(n3042) );
  AND2_X1 U2987 ( .A1(n3043), .A2(n2990), .ZN(n3041) );
  OR2_X1 U2988 ( .A1(n3044), .A2(n3045), .ZN(n2990) );
  AND2_X1 U2989 ( .A1(n2984), .A2(n2987), .ZN(n3045) );
  AND2_X1 U2990 ( .A1(n3046), .A2(n2986), .ZN(n3044) );
  OR2_X1 U2991 ( .A1(n3047), .A2(n3048), .ZN(n2986) );
  AND2_X1 U2992 ( .A1(n2980), .A2(n2983), .ZN(n3048) );
  AND2_X1 U2993 ( .A1(n3049), .A2(n2982), .ZN(n3047) );
  OR2_X1 U2994 ( .A1(n3050), .A2(n3051), .ZN(n2982) );
  AND2_X1 U2995 ( .A1(n2977), .A2(n2227), .ZN(n3051) );
  AND2_X1 U2996 ( .A1(n3052), .A2(n2979), .ZN(n3050) );
  OR2_X1 U2997 ( .A1(n3053), .A2(n3054), .ZN(n2979) );
  AND2_X1 U2998 ( .A1(n2973), .A2(n2976), .ZN(n3054) );
  AND2_X1 U2999 ( .A1(n3055), .A2(n2975), .ZN(n3053) );
  OR2_X1 U3000 ( .A1(n3056), .A2(n3057), .ZN(n2975) );
  AND2_X1 U3001 ( .A1(n2969), .A2(n2972), .ZN(n3057) );
  AND2_X1 U3002 ( .A1(n3058), .A2(n2971), .ZN(n3056) );
  OR2_X1 U3003 ( .A1(n3059), .A2(n3060), .ZN(n2971) );
  AND2_X1 U3004 ( .A1(n2965), .A2(n2968), .ZN(n3060) );
  AND2_X1 U3005 ( .A1(n2967), .A2(n3061), .ZN(n3059) );
  OR2_X1 U3006 ( .A1(n2968), .A2(n2965), .ZN(n3061) );
  OR2_X1 U3007 ( .A1(n2003), .A2(n2226), .ZN(n2965) );
  OR3_X1 U3008 ( .A1(n2550), .A2(n2226), .A3(n2060), .ZN(n2968) );
  INV_X1 U3009 ( .A(n3062), .ZN(n2967) );
  OR2_X1 U3010 ( .A1(n3063), .A2(n3064), .ZN(n3062) );
  AND2_X1 U3011 ( .A1(b_9_), .A2(n3065), .ZN(n3064) );
  OR2_X1 U3012 ( .A1(n3066), .A2(n1980), .ZN(n3065) );
  AND2_X1 U3013 ( .A1(a_14_), .A2(n2220), .ZN(n3066) );
  AND2_X1 U3014 ( .A1(b_8_), .A2(n3067), .ZN(n3063) );
  OR2_X1 U3015 ( .A1(n3068), .A2(n1983), .ZN(n3067) );
  AND2_X1 U3016 ( .A1(a_15_), .A2(n2060), .ZN(n3068) );
  OR2_X1 U3017 ( .A1(n2972), .A2(n2969), .ZN(n3058) );
  XNOR2_X1 U3018 ( .A(n3069), .B(n3070), .ZN(n2969) );
  XNOR2_X1 U3019 ( .A(n3071), .B(n3072), .ZN(n3070) );
  OR2_X1 U3020 ( .A1(n2231), .A2(n2226), .ZN(n2972) );
  OR2_X1 U3021 ( .A1(n2976), .A2(n2973), .ZN(n3055) );
  XOR2_X1 U3022 ( .A(n3073), .B(n3074), .Z(n2973) );
  XOR2_X1 U3023 ( .A(n3075), .B(n3076), .Z(n3074) );
  OR2_X1 U3024 ( .A1(n2032), .A2(n2226), .ZN(n2976) );
  OR2_X1 U3025 ( .A1(n2227), .A2(n2977), .ZN(n3052) );
  XOR2_X1 U3026 ( .A(n3077), .B(n3078), .Z(n2977) );
  XOR2_X1 U3027 ( .A(n3079), .B(n3080), .Z(n3078) );
  INV_X1 U3028 ( .A(n2044), .ZN(n2227) );
  AND2_X1 U3029 ( .A1(a_10_), .A2(b_10_), .ZN(n2044) );
  OR2_X1 U3030 ( .A1(n2983), .A2(n2980), .ZN(n3049) );
  XOR2_X1 U3031 ( .A(n3081), .B(n3082), .Z(n2980) );
  XOR2_X1 U3032 ( .A(n3083), .B(n3084), .Z(n3082) );
  OR2_X1 U3033 ( .A1(n2226), .A2(n2061), .ZN(n2983) );
  OR2_X1 U3034 ( .A1(n2987), .A2(n2984), .ZN(n3046) );
  XOR2_X1 U3035 ( .A(n3085), .B(n3086), .Z(n2984) );
  XOR2_X1 U3036 ( .A(n3087), .B(n2058), .Z(n3086) );
  OR2_X1 U3037 ( .A1(n2226), .A2(n2219), .ZN(n2987) );
  OR2_X1 U3038 ( .A1(n2991), .A2(n2988), .ZN(n3043) );
  XOR2_X1 U3039 ( .A(n3088), .B(n3089), .Z(n2988) );
  XOR2_X1 U3040 ( .A(n3090), .B(n3091), .Z(n3089) );
  OR2_X1 U3041 ( .A1(n2226), .A2(n2090), .ZN(n2991) );
  OR2_X1 U3042 ( .A1(n2995), .A2(n2992), .ZN(n3040) );
  XOR2_X1 U3043 ( .A(n3092), .B(n3093), .Z(n2992) );
  XOR2_X1 U3044 ( .A(n3094), .B(n3095), .Z(n3093) );
  OR2_X1 U3045 ( .A1(n2226), .A2(n2213), .ZN(n2995) );
  OR2_X1 U3046 ( .A1(n2999), .A2(n2996), .ZN(n3037) );
  XOR2_X1 U3047 ( .A(n3096), .B(n3097), .Z(n2996) );
  XOR2_X1 U3048 ( .A(n3098), .B(n3099), .Z(n3097) );
  OR2_X1 U3049 ( .A1(n2226), .A2(n2119), .ZN(n2999) );
  XOR2_X1 U3050 ( .A(n3100), .B(n3101), .Z(n3000) );
  XOR2_X1 U3051 ( .A(n3102), .B(n3103), .Z(n3101) );
  OR2_X1 U3052 ( .A1(n3007), .A2(n3004), .ZN(n3031) );
  XOR2_X1 U3053 ( .A(n3104), .B(n3105), .Z(n3004) );
  XOR2_X1 U3054 ( .A(n3106), .B(n3107), .Z(n3105) );
  OR2_X1 U3055 ( .A1(n2226), .A2(n2158), .ZN(n3007) );
  INV_X1 U3056 ( .A(b_10_), .ZN(n2226) );
  XOR2_X1 U3057 ( .A(n3108), .B(n3109), .Z(n3008) );
  XOR2_X1 U3058 ( .A(n3110), .B(n3111), .Z(n3109) );
  XOR2_X1 U3059 ( .A(n3112), .B(n3113), .Z(n3012) );
  XOR2_X1 U3060 ( .A(n3114), .B(n3115), .Z(n3113) );
  XOR2_X1 U3061 ( .A(n3116), .B(n3117), .Z(n3016) );
  XOR2_X1 U3062 ( .A(n3118), .B(n3119), .Z(n3117) );
  XNOR2_X1 U3063 ( .A(n3120), .B(n3121), .ZN(n1922) );
  XOR2_X1 U3064 ( .A(n3122), .B(n3123), .Z(n3121) );
  INV_X1 U3065 ( .A(n3124), .ZN(n1919) );
  OR2_X1 U3066 ( .A1(n3125), .A2(n2483), .ZN(n3124) );
  INV_X1 U3067 ( .A(n3126), .ZN(n2483) );
  OR2_X1 U3068 ( .A1(n3127), .A2(n3128), .ZN(n3126) );
  AND2_X1 U3069 ( .A1(n3127), .A2(n3128), .ZN(n3125) );
  OR2_X1 U3070 ( .A1(n3129), .A2(n3130), .ZN(n3128) );
  AND2_X1 U3071 ( .A1(n3123), .A2(n3122), .ZN(n3130) );
  AND2_X1 U3072 ( .A1(n3120), .A2(n3131), .ZN(n3129) );
  OR2_X1 U3073 ( .A1(n3122), .A2(n3123), .ZN(n3131) );
  OR2_X1 U3074 ( .A1(n2060), .A2(n2291), .ZN(n3123) );
  OR2_X1 U3075 ( .A1(n3132), .A2(n3133), .ZN(n3122) );
  AND2_X1 U3076 ( .A1(n3119), .A2(n3118), .ZN(n3133) );
  AND2_X1 U3077 ( .A1(n3116), .A2(n3134), .ZN(n3132) );
  OR2_X1 U3078 ( .A1(n3118), .A2(n3119), .ZN(n3134) );
  OR2_X1 U3079 ( .A1(n2060), .A2(n2187), .ZN(n3119) );
  OR2_X1 U3080 ( .A1(n3135), .A2(n3136), .ZN(n3118) );
  AND2_X1 U3081 ( .A1(n3115), .A2(n3114), .ZN(n3136) );
  AND2_X1 U3082 ( .A1(n3112), .A2(n3137), .ZN(n3135) );
  OR2_X1 U3083 ( .A1(n3114), .A2(n3115), .ZN(n3137) );
  OR2_X1 U3084 ( .A1(n2060), .A2(n2201), .ZN(n3115) );
  OR2_X1 U3085 ( .A1(n3138), .A2(n3139), .ZN(n3114) );
  AND2_X1 U3086 ( .A1(n3111), .A2(n3110), .ZN(n3139) );
  AND2_X1 U3087 ( .A1(n3108), .A2(n3140), .ZN(n3138) );
  OR2_X1 U3088 ( .A1(n3110), .A2(n3111), .ZN(n3140) );
  OR2_X1 U3089 ( .A1(n2060), .A2(n2158), .ZN(n3111) );
  OR2_X1 U3090 ( .A1(n3141), .A2(n3142), .ZN(n3110) );
  AND2_X1 U3091 ( .A1(n3104), .A2(n3107), .ZN(n3142) );
  AND2_X1 U3092 ( .A1(n3143), .A2(n3106), .ZN(n3141) );
  OR2_X1 U3093 ( .A1(n3144), .A2(n3145), .ZN(n3106) );
  AND2_X1 U3094 ( .A1(n3103), .A2(n3102), .ZN(n3145) );
  AND2_X1 U3095 ( .A1(n3100), .A2(n3146), .ZN(n3144) );
  OR2_X1 U3096 ( .A1(n3102), .A2(n3103), .ZN(n3146) );
  OR2_X1 U3097 ( .A1(n2060), .A2(n2119), .ZN(n3103) );
  OR2_X1 U3098 ( .A1(n3147), .A2(n3148), .ZN(n3102) );
  AND2_X1 U3099 ( .A1(n3096), .A2(n3099), .ZN(n3148) );
  AND2_X1 U3100 ( .A1(n3149), .A2(n3098), .ZN(n3147) );
  OR2_X1 U3101 ( .A1(n3150), .A2(n3151), .ZN(n3098) );
  AND2_X1 U3102 ( .A1(n3092), .A2(n3095), .ZN(n3151) );
  AND2_X1 U3103 ( .A1(n3152), .A2(n3094), .ZN(n3150) );
  OR2_X1 U3104 ( .A1(n3153), .A2(n3154), .ZN(n3094) );
  AND2_X1 U3105 ( .A1(n3088), .A2(n3091), .ZN(n3154) );
  AND2_X1 U3106 ( .A1(n3155), .A2(n3090), .ZN(n3153) );
  OR2_X1 U3107 ( .A1(n3156), .A2(n3157), .ZN(n3090) );
  AND2_X1 U3108 ( .A1(n3085), .A2(n2058), .ZN(n3157) );
  AND2_X1 U3109 ( .A1(n3158), .A2(n3087), .ZN(n3156) );
  OR2_X1 U3110 ( .A1(n3159), .A2(n3160), .ZN(n3087) );
  AND2_X1 U3111 ( .A1(n3081), .A2(n3084), .ZN(n3160) );
  AND2_X1 U3112 ( .A1(n3161), .A2(n3083), .ZN(n3159) );
  OR2_X1 U3113 ( .A1(n3162), .A2(n3163), .ZN(n3083) );
  AND2_X1 U3114 ( .A1(n3077), .A2(n3080), .ZN(n3163) );
  AND2_X1 U3115 ( .A1(n3164), .A2(n3079), .ZN(n3162) );
  OR2_X1 U3116 ( .A1(n3165), .A2(n3166), .ZN(n3079) );
  AND2_X1 U3117 ( .A1(n3073), .A2(n3076), .ZN(n3166) );
  AND2_X1 U3118 ( .A1(n3167), .A2(n3075), .ZN(n3165) );
  OR2_X1 U3119 ( .A1(n3168), .A2(n3169), .ZN(n3075) );
  AND2_X1 U3120 ( .A1(n3069), .A2(n3072), .ZN(n3169) );
  AND2_X1 U3121 ( .A1(n3071), .A2(n3170), .ZN(n3168) );
  OR2_X1 U3122 ( .A1(n3072), .A2(n3069), .ZN(n3170) );
  OR2_X1 U3123 ( .A1(n2003), .A2(n2060), .ZN(n3069) );
  OR3_X1 U3124 ( .A1(n2550), .A2(n2060), .A3(n2220), .ZN(n3072) );
  INV_X1 U3125 ( .A(n3171), .ZN(n3071) );
  OR2_X1 U3126 ( .A1(n3172), .A2(n3173), .ZN(n3171) );
  AND2_X1 U3127 ( .A1(b_8_), .A2(n3174), .ZN(n3173) );
  OR2_X1 U3128 ( .A1(n3175), .A2(n1980), .ZN(n3174) );
  AND2_X1 U3129 ( .A1(a_14_), .A2(n2089), .ZN(n3175) );
  AND2_X1 U3130 ( .A1(b_7_), .A2(n3176), .ZN(n3172) );
  OR2_X1 U3131 ( .A1(n3177), .A2(n1983), .ZN(n3176) );
  AND2_X1 U3132 ( .A1(a_15_), .A2(n2220), .ZN(n3177) );
  OR2_X1 U3133 ( .A1(n3076), .A2(n3073), .ZN(n3167) );
  XNOR2_X1 U3134 ( .A(n3178), .B(n3179), .ZN(n3073) );
  XNOR2_X1 U3135 ( .A(n3180), .B(n3181), .ZN(n3179) );
  OR2_X1 U3136 ( .A1(n2231), .A2(n2060), .ZN(n3076) );
  OR2_X1 U3137 ( .A1(n3080), .A2(n3077), .ZN(n3164) );
  XOR2_X1 U3138 ( .A(n3182), .B(n3183), .Z(n3077) );
  XOR2_X1 U3139 ( .A(n3184), .B(n3185), .Z(n3183) );
  OR2_X1 U3140 ( .A1(n2032), .A2(n2060), .ZN(n3080) );
  OR2_X1 U3141 ( .A1(n3084), .A2(n3081), .ZN(n3161) );
  XOR2_X1 U3142 ( .A(n3186), .B(n3187), .Z(n3081) );
  XOR2_X1 U3143 ( .A(n3188), .B(n3189), .Z(n3187) );
  OR2_X1 U3144 ( .A1(n2225), .A2(n2060), .ZN(n3084) );
  OR2_X1 U3145 ( .A1(n2058), .A2(n3085), .ZN(n3158) );
  XOR2_X1 U3146 ( .A(n3190), .B(n3191), .Z(n3085) );
  XOR2_X1 U3147 ( .A(n3192), .B(n3193), .Z(n3191) );
  OR2_X1 U3148 ( .A1(n2061), .A2(n2060), .ZN(n2058) );
  OR2_X1 U3149 ( .A1(n3091), .A2(n3088), .ZN(n3155) );
  XOR2_X1 U3150 ( .A(n3194), .B(n3195), .Z(n3088) );
  XOR2_X1 U3151 ( .A(n3196), .B(n3197), .Z(n3195) );
  OR2_X1 U3152 ( .A1(n2060), .A2(n2219), .ZN(n3091) );
  OR2_X1 U3153 ( .A1(n3095), .A2(n3092), .ZN(n3152) );
  XNOR2_X1 U3154 ( .A(n3198), .B(n3199), .ZN(n3092) );
  XNOR2_X1 U3155 ( .A(n2221), .B(n3200), .ZN(n3198) );
  OR2_X1 U3156 ( .A1(n2060), .A2(n2090), .ZN(n3095) );
  OR2_X1 U3157 ( .A1(n3099), .A2(n3096), .ZN(n3149) );
  XOR2_X1 U3158 ( .A(n3201), .B(n3202), .Z(n3096) );
  XOR2_X1 U3159 ( .A(n3203), .B(n3204), .Z(n3202) );
  OR2_X1 U3160 ( .A1(n2060), .A2(n2213), .ZN(n3099) );
  XOR2_X1 U3161 ( .A(n3205), .B(n3206), .Z(n3100) );
  XOR2_X1 U3162 ( .A(n3207), .B(n3208), .Z(n3206) );
  OR2_X1 U3163 ( .A1(n3107), .A2(n3104), .ZN(n3143) );
  XOR2_X1 U3164 ( .A(n3209), .B(n3210), .Z(n3104) );
  XOR2_X1 U3165 ( .A(n3211), .B(n3212), .Z(n3210) );
  OR2_X1 U3166 ( .A1(n2060), .A2(n2207), .ZN(n3107) );
  INV_X1 U3167 ( .A(b_9_), .ZN(n2060) );
  XOR2_X1 U3168 ( .A(n3213), .B(n3214), .Z(n3108) );
  XOR2_X1 U3169 ( .A(n3215), .B(n3216), .Z(n3214) );
  XOR2_X1 U3170 ( .A(n3217), .B(n3218), .Z(n3112) );
  XOR2_X1 U3171 ( .A(n3219), .B(n3220), .Z(n3218) );
  XOR2_X1 U3172 ( .A(n3221), .B(n3222), .Z(n3116) );
  XOR2_X1 U3173 ( .A(n3223), .B(n3224), .Z(n3222) );
  XOR2_X1 U3174 ( .A(n3225), .B(n3226), .Z(n3120) );
  XOR2_X1 U3175 ( .A(n3227), .B(n3228), .Z(n3226) );
  XOR2_X1 U3176 ( .A(n2442), .B(n3229), .Z(n3127) );
  XOR2_X1 U3177 ( .A(n2441), .B(n2440), .Z(n3229) );
  OR2_X1 U3178 ( .A1(n2220), .A2(n2291), .ZN(n2440) );
  OR2_X1 U3179 ( .A1(n3230), .A2(n3231), .ZN(n2441) );
  AND2_X1 U3180 ( .A1(n3228), .A2(n3227), .ZN(n3231) );
  AND2_X1 U3181 ( .A1(n3225), .A2(n3232), .ZN(n3230) );
  OR2_X1 U3182 ( .A1(n3227), .A2(n3228), .ZN(n3232) );
  OR2_X1 U3183 ( .A1(n2220), .A2(n2187), .ZN(n3228) );
  OR2_X1 U3184 ( .A1(n3233), .A2(n3234), .ZN(n3227) );
  AND2_X1 U3185 ( .A1(n3224), .A2(n3223), .ZN(n3234) );
  AND2_X1 U3186 ( .A1(n3221), .A2(n3235), .ZN(n3233) );
  OR2_X1 U3187 ( .A1(n3223), .A2(n3224), .ZN(n3235) );
  OR2_X1 U3188 ( .A1(n2220), .A2(n2201), .ZN(n3224) );
  OR2_X1 U3189 ( .A1(n3236), .A2(n3237), .ZN(n3223) );
  AND2_X1 U3190 ( .A1(n3220), .A2(n3219), .ZN(n3237) );
  AND2_X1 U3191 ( .A1(n3217), .A2(n3238), .ZN(n3236) );
  OR2_X1 U3192 ( .A1(n3219), .A2(n3220), .ZN(n3238) );
  OR2_X1 U3193 ( .A1(n2220), .A2(n2158), .ZN(n3220) );
  OR2_X1 U3194 ( .A1(n3239), .A2(n3240), .ZN(n3219) );
  AND2_X1 U3195 ( .A1(n3216), .A2(n3215), .ZN(n3240) );
  AND2_X1 U3196 ( .A1(n3213), .A2(n3241), .ZN(n3239) );
  OR2_X1 U3197 ( .A1(n3215), .A2(n3216), .ZN(n3241) );
  OR2_X1 U3198 ( .A1(n2220), .A2(n2207), .ZN(n3216) );
  OR2_X1 U3199 ( .A1(n3242), .A2(n3243), .ZN(n3215) );
  AND2_X1 U3200 ( .A1(n3209), .A2(n3212), .ZN(n3243) );
  AND2_X1 U3201 ( .A1(n3244), .A2(n3211), .ZN(n3242) );
  OR2_X1 U3202 ( .A1(n3245), .A2(n3246), .ZN(n3211) );
  AND2_X1 U3203 ( .A1(n3208), .A2(n3207), .ZN(n3246) );
  AND2_X1 U3204 ( .A1(n3205), .A2(n3247), .ZN(n3245) );
  OR2_X1 U3205 ( .A1(n3207), .A2(n3208), .ZN(n3247) );
  OR2_X1 U3206 ( .A1(n2220), .A2(n2213), .ZN(n3208) );
  OR2_X1 U3207 ( .A1(n3248), .A2(n3249), .ZN(n3207) );
  AND2_X1 U3208 ( .A1(n3201), .A2(n3204), .ZN(n3249) );
  AND2_X1 U3209 ( .A1(n3250), .A2(n3203), .ZN(n3248) );
  OR2_X1 U3210 ( .A1(n3251), .A2(n3252), .ZN(n3203) );
  AND2_X1 U3211 ( .A1(n3199), .A2(n2221), .ZN(n3252) );
  AND2_X1 U3212 ( .A1(n3253), .A2(n3200), .ZN(n3251) );
  OR2_X1 U3213 ( .A1(n3254), .A2(n3255), .ZN(n3200) );
  AND2_X1 U3214 ( .A1(n3194), .A2(n3197), .ZN(n3255) );
  AND2_X1 U3215 ( .A1(n3256), .A2(n3196), .ZN(n3254) );
  OR2_X1 U3216 ( .A1(n3257), .A2(n3258), .ZN(n3196) );
  AND2_X1 U3217 ( .A1(n3190), .A2(n3193), .ZN(n3258) );
  AND2_X1 U3218 ( .A1(n3259), .A2(n3192), .ZN(n3257) );
  OR2_X1 U3219 ( .A1(n3260), .A2(n3261), .ZN(n3192) );
  AND2_X1 U3220 ( .A1(n3186), .A2(n3189), .ZN(n3261) );
  AND2_X1 U3221 ( .A1(n3262), .A2(n3188), .ZN(n3260) );
  OR2_X1 U3222 ( .A1(n3263), .A2(n3264), .ZN(n3188) );
  AND2_X1 U3223 ( .A1(n3182), .A2(n3185), .ZN(n3264) );
  AND2_X1 U3224 ( .A1(n3265), .A2(n3184), .ZN(n3263) );
  OR2_X1 U3225 ( .A1(n3266), .A2(n3267), .ZN(n3184) );
  AND2_X1 U3226 ( .A1(n3178), .A2(n3181), .ZN(n3267) );
  AND2_X1 U3227 ( .A1(n3180), .A2(n3268), .ZN(n3266) );
  OR2_X1 U3228 ( .A1(n3181), .A2(n3178), .ZN(n3268) );
  OR2_X1 U3229 ( .A1(n2003), .A2(n2220), .ZN(n3178) );
  OR3_X1 U3230 ( .A1(n2550), .A2(n2220), .A3(n2089), .ZN(n3181) );
  INV_X1 U3231 ( .A(n3269), .ZN(n3180) );
  OR2_X1 U3232 ( .A1(n3270), .A2(n3271), .ZN(n3269) );
  AND2_X1 U3233 ( .A1(b_7_), .A2(n3272), .ZN(n3271) );
  OR2_X1 U3234 ( .A1(n3273), .A2(n1980), .ZN(n3272) );
  AND2_X1 U3235 ( .A1(a_14_), .A2(n2214), .ZN(n3273) );
  AND2_X1 U3236 ( .A1(b_6_), .A2(n3274), .ZN(n3270) );
  OR2_X1 U3237 ( .A1(n3275), .A2(n1983), .ZN(n3274) );
  AND2_X1 U3238 ( .A1(a_15_), .A2(n2089), .ZN(n3275) );
  OR2_X1 U3239 ( .A1(n3185), .A2(n3182), .ZN(n3265) );
  XNOR2_X1 U3240 ( .A(n3276), .B(n3277), .ZN(n3182) );
  XNOR2_X1 U3241 ( .A(n3278), .B(n3279), .ZN(n3277) );
  OR2_X1 U3242 ( .A1(n2231), .A2(n2220), .ZN(n3185) );
  OR2_X1 U3243 ( .A1(n3189), .A2(n3186), .ZN(n3262) );
  XOR2_X1 U3244 ( .A(n3280), .B(n3281), .Z(n3186) );
  XOR2_X1 U3245 ( .A(n3282), .B(n3283), .Z(n3281) );
  OR2_X1 U3246 ( .A1(n2032), .A2(n2220), .ZN(n3189) );
  OR2_X1 U3247 ( .A1(n3193), .A2(n3190), .ZN(n3259) );
  XOR2_X1 U3248 ( .A(n3284), .B(n3285), .Z(n3190) );
  XOR2_X1 U3249 ( .A(n3286), .B(n3287), .Z(n3285) );
  OR2_X1 U3250 ( .A1(n2225), .A2(n2220), .ZN(n3193) );
  OR2_X1 U3251 ( .A1(n3197), .A2(n3194), .ZN(n3256) );
  XOR2_X1 U3252 ( .A(n3288), .B(n3289), .Z(n3194) );
  XOR2_X1 U3253 ( .A(n3290), .B(n3291), .Z(n3289) );
  OR2_X1 U3254 ( .A1(n2061), .A2(n2220), .ZN(n3197) );
  OR2_X1 U3255 ( .A1(n2221), .A2(n3199), .ZN(n3253) );
  XOR2_X1 U3256 ( .A(n3292), .B(n3293), .Z(n3199) );
  XOR2_X1 U3257 ( .A(n3294), .B(n3295), .Z(n3293) );
  INV_X1 U3258 ( .A(n2073), .ZN(n2221) );
  AND2_X1 U3259 ( .A1(a_8_), .A2(b_8_), .ZN(n2073) );
  OR2_X1 U3260 ( .A1(n3204), .A2(n3201), .ZN(n3250) );
  XOR2_X1 U3261 ( .A(n3296), .B(n3297), .Z(n3201) );
  XOR2_X1 U3262 ( .A(n3298), .B(n3299), .Z(n3297) );
  OR2_X1 U3263 ( .A1(n2220), .A2(n2090), .ZN(n3204) );
  XOR2_X1 U3264 ( .A(n3300), .B(n3301), .Z(n3205) );
  XOR2_X1 U3265 ( .A(n3302), .B(n2087), .Z(n3301) );
  OR2_X1 U3266 ( .A1(n3212), .A2(n3209), .ZN(n3244) );
  XOR2_X1 U3267 ( .A(n3303), .B(n3304), .Z(n3209) );
  XOR2_X1 U3268 ( .A(n3305), .B(n3306), .Z(n3304) );
  OR2_X1 U3269 ( .A1(n2220), .A2(n2119), .ZN(n3212) );
  INV_X1 U3270 ( .A(b_8_), .ZN(n2220) );
  XOR2_X1 U3271 ( .A(n3307), .B(n3308), .Z(n3213) );
  XOR2_X1 U3272 ( .A(n3309), .B(n3310), .Z(n3308) );
  XOR2_X1 U3273 ( .A(n3311), .B(n3312), .Z(n3217) );
  XOR2_X1 U3274 ( .A(n3313), .B(n3314), .Z(n3312) );
  XOR2_X1 U3275 ( .A(n3315), .B(n3316), .Z(n3221) );
  XOR2_X1 U3276 ( .A(n3317), .B(n3318), .Z(n3316) );
  XOR2_X1 U3277 ( .A(n3319), .B(n3320), .Z(n3225) );
  XOR2_X1 U3278 ( .A(n3321), .B(n3322), .Z(n3320) );
  XOR2_X1 U3279 ( .A(n2449), .B(n3323), .Z(n2442) );
  XOR2_X1 U3280 ( .A(n2448), .B(n2447), .Z(n3323) );
  OR2_X1 U3281 ( .A1(n2089), .A2(n2187), .ZN(n2447) );
  OR2_X1 U3282 ( .A1(n3324), .A2(n3325), .ZN(n2448) );
  AND2_X1 U3283 ( .A1(n3322), .A2(n3321), .ZN(n3325) );
  AND2_X1 U3284 ( .A1(n3319), .A2(n3326), .ZN(n3324) );
  OR2_X1 U3285 ( .A1(n3321), .A2(n3322), .ZN(n3326) );
  OR2_X1 U3286 ( .A1(n2089), .A2(n2201), .ZN(n3322) );
  OR2_X1 U3287 ( .A1(n3327), .A2(n3328), .ZN(n3321) );
  AND2_X1 U3288 ( .A1(n3318), .A2(n3317), .ZN(n3328) );
  AND2_X1 U3289 ( .A1(n3315), .A2(n3329), .ZN(n3327) );
  OR2_X1 U3290 ( .A1(n3317), .A2(n3318), .ZN(n3329) );
  OR2_X1 U3291 ( .A1(n2089), .A2(n2158), .ZN(n3318) );
  OR2_X1 U3292 ( .A1(n3330), .A2(n3331), .ZN(n3317) );
  AND2_X1 U3293 ( .A1(n3314), .A2(n3313), .ZN(n3331) );
  AND2_X1 U3294 ( .A1(n3311), .A2(n3332), .ZN(n3330) );
  OR2_X1 U3295 ( .A1(n3313), .A2(n3314), .ZN(n3332) );
  OR2_X1 U3296 ( .A1(n2089), .A2(n2207), .ZN(n3314) );
  OR2_X1 U3297 ( .A1(n3333), .A2(n3334), .ZN(n3313) );
  AND2_X1 U3298 ( .A1(n3310), .A2(n3309), .ZN(n3334) );
  AND2_X1 U3299 ( .A1(n3307), .A2(n3335), .ZN(n3333) );
  OR2_X1 U3300 ( .A1(n3309), .A2(n3310), .ZN(n3335) );
  OR2_X1 U3301 ( .A1(n2089), .A2(n2119), .ZN(n3310) );
  OR2_X1 U3302 ( .A1(n3336), .A2(n3337), .ZN(n3309) );
  AND2_X1 U3303 ( .A1(n3303), .A2(n3306), .ZN(n3337) );
  AND2_X1 U3304 ( .A1(n3338), .A2(n3305), .ZN(n3336) );
  OR2_X1 U3305 ( .A1(n3339), .A2(n3340), .ZN(n3305) );
  AND2_X1 U3306 ( .A1(n2087), .A2(n3302), .ZN(n3340) );
  AND2_X1 U3307 ( .A1(n3300), .A2(n3341), .ZN(n3339) );
  OR2_X1 U3308 ( .A1(n3302), .A2(n2087), .ZN(n3341) );
  OR2_X1 U3309 ( .A1(n2090), .A2(n2089), .ZN(n2087) );
  OR2_X1 U3310 ( .A1(n3342), .A2(n3343), .ZN(n3302) );
  AND2_X1 U3311 ( .A1(n3296), .A2(n3299), .ZN(n3343) );
  AND2_X1 U3312 ( .A1(n3344), .A2(n3298), .ZN(n3342) );
  OR2_X1 U3313 ( .A1(n3345), .A2(n3346), .ZN(n3298) );
  AND2_X1 U3314 ( .A1(n3292), .A2(n3295), .ZN(n3346) );
  AND2_X1 U3315 ( .A1(n3347), .A2(n3294), .ZN(n3345) );
  OR2_X1 U3316 ( .A1(n3348), .A2(n3349), .ZN(n3294) );
  AND2_X1 U3317 ( .A1(n3288), .A2(n3291), .ZN(n3349) );
  AND2_X1 U3318 ( .A1(n3350), .A2(n3290), .ZN(n3348) );
  OR2_X1 U3319 ( .A1(n3351), .A2(n3352), .ZN(n3290) );
  AND2_X1 U3320 ( .A1(n3284), .A2(n3287), .ZN(n3352) );
  AND2_X1 U3321 ( .A1(n3353), .A2(n3286), .ZN(n3351) );
  OR2_X1 U3322 ( .A1(n3354), .A2(n3355), .ZN(n3286) );
  AND2_X1 U3323 ( .A1(n3280), .A2(n3283), .ZN(n3355) );
  AND2_X1 U3324 ( .A1(n3356), .A2(n3282), .ZN(n3354) );
  OR2_X1 U3325 ( .A1(n3357), .A2(n3358), .ZN(n3282) );
  AND2_X1 U3326 ( .A1(n3276), .A2(n3279), .ZN(n3358) );
  AND2_X1 U3327 ( .A1(n3278), .A2(n3359), .ZN(n3357) );
  OR2_X1 U3328 ( .A1(n3279), .A2(n3276), .ZN(n3359) );
  OR2_X1 U3329 ( .A1(n2003), .A2(n2089), .ZN(n3276) );
  OR3_X1 U3330 ( .A1(n2550), .A2(n2089), .A3(n2214), .ZN(n3279) );
  INV_X1 U3331 ( .A(n3360), .ZN(n3278) );
  OR2_X1 U3332 ( .A1(n3361), .A2(n3362), .ZN(n3360) );
  AND2_X1 U3333 ( .A1(b_6_), .A2(n3363), .ZN(n3362) );
  OR2_X1 U3334 ( .A1(n3364), .A2(n1980), .ZN(n3363) );
  AND2_X1 U3335 ( .A1(a_14_), .A2(n2118), .ZN(n3364) );
  AND2_X1 U3336 ( .A1(b_5_), .A2(n3365), .ZN(n3361) );
  OR2_X1 U3337 ( .A1(n3366), .A2(n1983), .ZN(n3365) );
  AND2_X1 U3338 ( .A1(a_15_), .A2(n2214), .ZN(n3366) );
  OR2_X1 U3339 ( .A1(n3283), .A2(n3280), .ZN(n3356) );
  XNOR2_X1 U3340 ( .A(n3367), .B(n3368), .ZN(n3280) );
  XNOR2_X1 U3341 ( .A(n3369), .B(n3370), .ZN(n3368) );
  OR2_X1 U3342 ( .A1(n2231), .A2(n2089), .ZN(n3283) );
  OR2_X1 U3343 ( .A1(n3287), .A2(n3284), .ZN(n3353) );
  XOR2_X1 U3344 ( .A(n3371), .B(n3372), .Z(n3284) );
  XOR2_X1 U3345 ( .A(n3373), .B(n3374), .Z(n3372) );
  OR2_X1 U3346 ( .A1(n2032), .A2(n2089), .ZN(n3287) );
  OR2_X1 U3347 ( .A1(n3291), .A2(n3288), .ZN(n3350) );
  XOR2_X1 U3348 ( .A(n3375), .B(n3376), .Z(n3288) );
  XOR2_X1 U3349 ( .A(n3377), .B(n3378), .Z(n3376) );
  OR2_X1 U3350 ( .A1(n2225), .A2(n2089), .ZN(n3291) );
  OR2_X1 U3351 ( .A1(n3295), .A2(n3292), .ZN(n3347) );
  XOR2_X1 U3352 ( .A(n3379), .B(n3380), .Z(n3292) );
  XOR2_X1 U3353 ( .A(n3381), .B(n3382), .Z(n3380) );
  OR2_X1 U3354 ( .A1(n2061), .A2(n2089), .ZN(n3295) );
  OR2_X1 U3355 ( .A1(n3299), .A2(n3296), .ZN(n3344) );
  XOR2_X1 U3356 ( .A(n3383), .B(n3384), .Z(n3296) );
  XOR2_X1 U3357 ( .A(n3385), .B(n3386), .Z(n3384) );
  OR2_X1 U3358 ( .A1(n2219), .A2(n2089), .ZN(n3299) );
  XOR2_X1 U3359 ( .A(n3387), .B(n3388), .Z(n3300) );
  XOR2_X1 U3360 ( .A(n3389), .B(n3390), .Z(n3388) );
  OR2_X1 U3361 ( .A1(n3306), .A2(n3303), .ZN(n3338) );
  XOR2_X1 U3362 ( .A(n3391), .B(n3392), .Z(n3303) );
  XOR2_X1 U3363 ( .A(n3393), .B(n3394), .Z(n3392) );
  OR2_X1 U3364 ( .A1(n2089), .A2(n2213), .ZN(n3306) );
  INV_X1 U3365 ( .A(b_7_), .ZN(n2089) );
  XNOR2_X1 U3366 ( .A(n3395), .B(n3396), .ZN(n3307) );
  XNOR2_X1 U3367 ( .A(n2215), .B(n3397), .ZN(n3395) );
  XOR2_X1 U3368 ( .A(n3398), .B(n3399), .Z(n3311) );
  XOR2_X1 U3369 ( .A(n3400), .B(n3401), .Z(n3399) );
  XOR2_X1 U3370 ( .A(n3402), .B(n3403), .Z(n3315) );
  XOR2_X1 U3371 ( .A(n3404), .B(n3405), .Z(n3403) );
  XOR2_X1 U3372 ( .A(n3406), .B(n3407), .Z(n3319) );
  XOR2_X1 U3373 ( .A(n3408), .B(n3409), .Z(n3407) );
  XOR2_X1 U3374 ( .A(n2456), .B(n3410), .Z(n2449) );
  XOR2_X1 U3375 ( .A(n2455), .B(n2454), .Z(n3410) );
  OR2_X1 U3376 ( .A1(n2214), .A2(n2201), .ZN(n2454) );
  OR2_X1 U3377 ( .A1(n3411), .A2(n3412), .ZN(n2455) );
  AND2_X1 U3378 ( .A1(n3409), .A2(n3408), .ZN(n3412) );
  AND2_X1 U3379 ( .A1(n3406), .A2(n3413), .ZN(n3411) );
  OR2_X1 U3380 ( .A1(n3408), .A2(n3409), .ZN(n3413) );
  OR2_X1 U3381 ( .A1(n2214), .A2(n2158), .ZN(n3409) );
  OR2_X1 U3382 ( .A1(n3414), .A2(n3415), .ZN(n3408) );
  AND2_X1 U3383 ( .A1(n3405), .A2(n3404), .ZN(n3415) );
  AND2_X1 U3384 ( .A1(n3402), .A2(n3416), .ZN(n3414) );
  OR2_X1 U3385 ( .A1(n3404), .A2(n3405), .ZN(n3416) );
  OR2_X1 U3386 ( .A1(n2214), .A2(n2207), .ZN(n3405) );
  OR2_X1 U3387 ( .A1(n3417), .A2(n3418), .ZN(n3404) );
  AND2_X1 U3388 ( .A1(n3401), .A2(n3400), .ZN(n3418) );
  AND2_X1 U3389 ( .A1(n3398), .A2(n3419), .ZN(n3417) );
  OR2_X1 U3390 ( .A1(n3400), .A2(n3401), .ZN(n3419) );
  OR2_X1 U3391 ( .A1(n2214), .A2(n2119), .ZN(n3401) );
  OR2_X1 U3392 ( .A1(n3420), .A2(n3421), .ZN(n3400) );
  AND2_X1 U3393 ( .A1(n3397), .A2(n2215), .ZN(n3421) );
  AND2_X1 U3394 ( .A1(n3396), .A2(n3422), .ZN(n3420) );
  OR2_X1 U3395 ( .A1(n2215), .A2(n3397), .ZN(n3422) );
  OR2_X1 U3396 ( .A1(n3423), .A2(n3424), .ZN(n3397) );
  AND2_X1 U3397 ( .A1(n3391), .A2(n3394), .ZN(n3424) );
  AND2_X1 U3398 ( .A1(n3425), .A2(n3393), .ZN(n3423) );
  OR2_X1 U3399 ( .A1(n3426), .A2(n3427), .ZN(n3393) );
  AND2_X1 U3400 ( .A1(n3390), .A2(n3389), .ZN(n3427) );
  AND2_X1 U3401 ( .A1(n3387), .A2(n3428), .ZN(n3426) );
  OR2_X1 U3402 ( .A1(n3389), .A2(n3390), .ZN(n3428) );
  OR2_X1 U3403 ( .A1(n2219), .A2(n2214), .ZN(n3390) );
  OR2_X1 U3404 ( .A1(n3429), .A2(n3430), .ZN(n3389) );
  AND2_X1 U3405 ( .A1(n3383), .A2(n3386), .ZN(n3430) );
  AND2_X1 U3406 ( .A1(n3431), .A2(n3385), .ZN(n3429) );
  OR2_X1 U3407 ( .A1(n3432), .A2(n3433), .ZN(n3385) );
  AND2_X1 U3408 ( .A1(n3379), .A2(n3382), .ZN(n3433) );
  AND2_X1 U3409 ( .A1(n3434), .A2(n3381), .ZN(n3432) );
  OR2_X1 U3410 ( .A1(n3435), .A2(n3436), .ZN(n3381) );
  AND2_X1 U3411 ( .A1(n3375), .A2(n3378), .ZN(n3436) );
  AND2_X1 U3412 ( .A1(n3437), .A2(n3377), .ZN(n3435) );
  OR2_X1 U3413 ( .A1(n3438), .A2(n3439), .ZN(n3377) );
  AND2_X1 U3414 ( .A1(n3371), .A2(n3374), .ZN(n3439) );
  AND2_X1 U3415 ( .A1(n3440), .A2(n3373), .ZN(n3438) );
  OR2_X1 U3416 ( .A1(n3441), .A2(n3442), .ZN(n3373) );
  AND2_X1 U3417 ( .A1(n3367), .A2(n3370), .ZN(n3442) );
  AND2_X1 U3418 ( .A1(n3369), .A2(n3443), .ZN(n3441) );
  OR2_X1 U3419 ( .A1(n3370), .A2(n3367), .ZN(n3443) );
  OR2_X1 U3420 ( .A1(n2003), .A2(n2214), .ZN(n3367) );
  OR3_X1 U3421 ( .A1(n2550), .A2(n2214), .A3(n2118), .ZN(n3370) );
  INV_X1 U3422 ( .A(n3444), .ZN(n3369) );
  OR2_X1 U3423 ( .A1(n3445), .A2(n3446), .ZN(n3444) );
  AND2_X1 U3424 ( .A1(b_5_), .A2(n3447), .ZN(n3446) );
  OR2_X1 U3425 ( .A1(n3448), .A2(n1980), .ZN(n3447) );
  AND2_X1 U3426 ( .A1(a_14_), .A2(n2208), .ZN(n3448) );
  AND2_X1 U3427 ( .A1(b_4_), .A2(n3449), .ZN(n3445) );
  OR2_X1 U3428 ( .A1(n3450), .A2(n1983), .ZN(n3449) );
  AND2_X1 U3429 ( .A1(a_15_), .A2(n2118), .ZN(n3450) );
  OR2_X1 U3430 ( .A1(n3374), .A2(n3371), .ZN(n3440) );
  XNOR2_X1 U3431 ( .A(n3451), .B(n3452), .ZN(n3371) );
  XNOR2_X1 U3432 ( .A(n3453), .B(n3454), .ZN(n3452) );
  OR2_X1 U3433 ( .A1(n2231), .A2(n2214), .ZN(n3374) );
  OR2_X1 U3434 ( .A1(n3378), .A2(n3375), .ZN(n3437) );
  XOR2_X1 U3435 ( .A(n3455), .B(n3456), .Z(n3375) );
  XOR2_X1 U3436 ( .A(n3457), .B(n3458), .Z(n3456) );
  OR2_X1 U3437 ( .A1(n2032), .A2(n2214), .ZN(n3378) );
  OR2_X1 U3438 ( .A1(n3382), .A2(n3379), .ZN(n3434) );
  XOR2_X1 U3439 ( .A(n3459), .B(n3460), .Z(n3379) );
  XOR2_X1 U3440 ( .A(n3461), .B(n3462), .Z(n3460) );
  OR2_X1 U3441 ( .A1(n2225), .A2(n2214), .ZN(n3382) );
  OR2_X1 U3442 ( .A1(n3386), .A2(n3383), .ZN(n3431) );
  XOR2_X1 U3443 ( .A(n3463), .B(n3464), .Z(n3383) );
  XOR2_X1 U3444 ( .A(n3465), .B(n3466), .Z(n3464) );
  OR2_X1 U3445 ( .A1(n2061), .A2(n2214), .ZN(n3386) );
  XOR2_X1 U3446 ( .A(n3467), .B(n3468), .Z(n3387) );
  XOR2_X1 U3447 ( .A(n3469), .B(n3470), .Z(n3468) );
  OR2_X1 U3448 ( .A1(n3394), .A2(n3391), .ZN(n3425) );
  XOR2_X1 U3449 ( .A(n3471), .B(n3472), .Z(n3391) );
  XOR2_X1 U3450 ( .A(n3473), .B(n3474), .Z(n3472) );
  OR2_X1 U3451 ( .A1(n2090), .A2(n2214), .ZN(n3394) );
  INV_X1 U3452 ( .A(b_6_), .ZN(n2214) );
  INV_X1 U3453 ( .A(n2102), .ZN(n2215) );
  AND2_X1 U3454 ( .A1(a_6_), .A2(b_6_), .ZN(n2102) );
  XOR2_X1 U3455 ( .A(n3475), .B(n3476), .Z(n3396) );
  XOR2_X1 U3456 ( .A(n3477), .B(n3478), .Z(n3476) );
  XOR2_X1 U3457 ( .A(n3479), .B(n3480), .Z(n3398) );
  XOR2_X1 U3458 ( .A(n3481), .B(n3482), .Z(n3480) );
  XOR2_X1 U3459 ( .A(n3483), .B(n3484), .Z(n3402) );
  XOR2_X1 U3460 ( .A(n3485), .B(n2116), .Z(n3484) );
  XOR2_X1 U3461 ( .A(n3486), .B(n3487), .Z(n3406) );
  XOR2_X1 U3462 ( .A(n3488), .B(n3489), .Z(n3487) );
  XOR2_X1 U3463 ( .A(n2463), .B(n3490), .Z(n2456) );
  XOR2_X1 U3464 ( .A(n2462), .B(n2461), .Z(n3490) );
  OR2_X1 U3465 ( .A1(n2118), .A2(n2158), .ZN(n2461) );
  OR2_X1 U3466 ( .A1(n3491), .A2(n3492), .ZN(n2462) );
  AND2_X1 U3467 ( .A1(n3489), .A2(n3488), .ZN(n3492) );
  AND2_X1 U3468 ( .A1(n3486), .A2(n3493), .ZN(n3491) );
  OR2_X1 U3469 ( .A1(n3488), .A2(n3489), .ZN(n3493) );
  OR2_X1 U3470 ( .A1(n2118), .A2(n2207), .ZN(n3489) );
  OR2_X1 U3471 ( .A1(n3494), .A2(n3495), .ZN(n3488) );
  AND2_X1 U3472 ( .A1(n2116), .A2(n3485), .ZN(n3495) );
  AND2_X1 U3473 ( .A1(n3483), .A2(n3496), .ZN(n3494) );
  OR2_X1 U3474 ( .A1(n3485), .A2(n2116), .ZN(n3496) );
  OR2_X1 U3475 ( .A1(n2119), .A2(n2118), .ZN(n2116) );
  OR2_X1 U3476 ( .A1(n3497), .A2(n3498), .ZN(n3485) );
  AND2_X1 U3477 ( .A1(n3482), .A2(n3481), .ZN(n3498) );
  AND2_X1 U3478 ( .A1(n3479), .A2(n3499), .ZN(n3497) );
  OR2_X1 U3479 ( .A1(n3481), .A2(n3482), .ZN(n3499) );
  OR2_X1 U3480 ( .A1(n2213), .A2(n2118), .ZN(n3482) );
  OR2_X1 U3481 ( .A1(n3500), .A2(n3501), .ZN(n3481) );
  AND2_X1 U3482 ( .A1(n3478), .A2(n3477), .ZN(n3501) );
  AND2_X1 U3483 ( .A1(n3475), .A2(n3502), .ZN(n3500) );
  OR2_X1 U3484 ( .A1(n3477), .A2(n3478), .ZN(n3502) );
  OR2_X1 U3485 ( .A1(n2090), .A2(n2118), .ZN(n3478) );
  OR2_X1 U3486 ( .A1(n3503), .A2(n3504), .ZN(n3477) );
  AND2_X1 U3487 ( .A1(n3471), .A2(n3474), .ZN(n3504) );
  AND2_X1 U3488 ( .A1(n3505), .A2(n3473), .ZN(n3503) );
  OR2_X1 U3489 ( .A1(n3506), .A2(n3507), .ZN(n3473) );
  AND2_X1 U3490 ( .A1(n3470), .A2(n3469), .ZN(n3507) );
  AND2_X1 U3491 ( .A1(n3467), .A2(n3508), .ZN(n3506) );
  OR2_X1 U3492 ( .A1(n3469), .A2(n3470), .ZN(n3508) );
  OR2_X1 U3493 ( .A1(n2061), .A2(n2118), .ZN(n3470) );
  OR2_X1 U3494 ( .A1(n3509), .A2(n3510), .ZN(n3469) );
  AND2_X1 U3495 ( .A1(n3463), .A2(n3466), .ZN(n3510) );
  AND2_X1 U3496 ( .A1(n3511), .A2(n3465), .ZN(n3509) );
  OR2_X1 U3497 ( .A1(n3512), .A2(n3513), .ZN(n3465) );
  AND2_X1 U3498 ( .A1(n3459), .A2(n3462), .ZN(n3513) );
  AND2_X1 U3499 ( .A1(n3514), .A2(n3461), .ZN(n3512) );
  OR2_X1 U3500 ( .A1(n3515), .A2(n3516), .ZN(n3461) );
  AND2_X1 U3501 ( .A1(n3455), .A2(n3458), .ZN(n3516) );
  AND2_X1 U3502 ( .A1(n3517), .A2(n3457), .ZN(n3515) );
  OR2_X1 U3503 ( .A1(n3518), .A2(n3519), .ZN(n3457) );
  AND2_X1 U3504 ( .A1(n3451), .A2(n3454), .ZN(n3519) );
  AND2_X1 U3505 ( .A1(n3453), .A2(n3520), .ZN(n3518) );
  OR2_X1 U3506 ( .A1(n3454), .A2(n3451), .ZN(n3520) );
  OR2_X1 U3507 ( .A1(n2003), .A2(n2118), .ZN(n3451) );
  OR3_X1 U3508 ( .A1(n2550), .A2(n2118), .A3(n2208), .ZN(n3454) );
  INV_X1 U3509 ( .A(n3521), .ZN(n3453) );
  OR2_X1 U3510 ( .A1(n3522), .A2(n3523), .ZN(n3521) );
  AND2_X1 U3511 ( .A1(b_4_), .A2(n3524), .ZN(n3523) );
  OR2_X1 U3512 ( .A1(n3525), .A2(n1980), .ZN(n3524) );
  AND2_X1 U3513 ( .A1(a_14_), .A2(n2157), .ZN(n3525) );
  AND2_X1 U3514 ( .A1(b_3_), .A2(n3526), .ZN(n3522) );
  OR2_X1 U3515 ( .A1(n3527), .A2(n1983), .ZN(n3526) );
  AND2_X1 U3516 ( .A1(a_15_), .A2(n2208), .ZN(n3527) );
  OR2_X1 U3517 ( .A1(n3458), .A2(n3455), .ZN(n3517) );
  XNOR2_X1 U3518 ( .A(n3528), .B(n3529), .ZN(n3455) );
  XNOR2_X1 U3519 ( .A(n3530), .B(n3531), .ZN(n3529) );
  OR2_X1 U3520 ( .A1(n2231), .A2(n2118), .ZN(n3458) );
  OR2_X1 U3521 ( .A1(n3462), .A2(n3459), .ZN(n3514) );
  XOR2_X1 U3522 ( .A(n3532), .B(n3533), .Z(n3459) );
  XOR2_X1 U3523 ( .A(n3534), .B(n3535), .Z(n3533) );
  OR2_X1 U3524 ( .A1(n2032), .A2(n2118), .ZN(n3462) );
  OR2_X1 U3525 ( .A1(n3466), .A2(n3463), .ZN(n3511) );
  XOR2_X1 U3526 ( .A(n3536), .B(n3537), .Z(n3463) );
  XOR2_X1 U3527 ( .A(n3538), .B(n3539), .Z(n3537) );
  OR2_X1 U3528 ( .A1(n2225), .A2(n2118), .ZN(n3466) );
  XOR2_X1 U3529 ( .A(n3540), .B(n3541), .Z(n3467) );
  XOR2_X1 U3530 ( .A(n3542), .B(n3543), .Z(n3541) );
  OR2_X1 U3531 ( .A1(n3474), .A2(n3471), .ZN(n3505) );
  XOR2_X1 U3532 ( .A(n3544), .B(n3545), .Z(n3471) );
  XOR2_X1 U3533 ( .A(n3546), .B(n3547), .Z(n3545) );
  OR2_X1 U3534 ( .A1(n2219), .A2(n2118), .ZN(n3474) );
  INV_X1 U3535 ( .A(b_5_), .ZN(n2118) );
  XOR2_X1 U3536 ( .A(n3548), .B(n3549), .Z(n3475) );
  XOR2_X1 U3537 ( .A(n3550), .B(n3551), .Z(n3549) );
  XOR2_X1 U3538 ( .A(n3552), .B(n3553), .Z(n3479) );
  XOR2_X1 U3539 ( .A(n3554), .B(n3555), .Z(n3553) );
  XOR2_X1 U3540 ( .A(n3556), .B(n3557), .Z(n3483) );
  XOR2_X1 U3541 ( .A(n3558), .B(n3559), .Z(n3557) );
  XOR2_X1 U3542 ( .A(n3560), .B(n3561), .Z(n3486) );
  XOR2_X1 U3543 ( .A(n3562), .B(n3563), .Z(n3561) );
  XNOR2_X1 U3544 ( .A(n3564), .B(n2469), .ZN(n2463) );
  XOR2_X1 U3545 ( .A(n2476), .B(n3565), .Z(n2469) );
  XOR2_X1 U3546 ( .A(n2475), .B(n2474), .Z(n3565) );
  OR2_X1 U3547 ( .A1(n2119), .A2(n2157), .ZN(n2474) );
  OR2_X1 U3548 ( .A1(n3566), .A2(n3567), .ZN(n2475) );
  AND2_X1 U3549 ( .A1(n3568), .A2(n3569), .ZN(n3567) );
  AND2_X1 U3550 ( .A1(n3570), .A2(n3571), .ZN(n3566) );
  OR2_X1 U3551 ( .A1(n3569), .A2(n3568), .ZN(n3571) );
  XOR2_X1 U3552 ( .A(n3572), .B(n3573), .Z(n2476) );
  XOR2_X1 U3553 ( .A(n3574), .B(n3575), .Z(n3573) );
  XNOR2_X1 U3554 ( .A(n2209), .B(n2468), .ZN(n3564) );
  OR2_X1 U3555 ( .A1(n3576), .A2(n3577), .ZN(n2468) );
  AND2_X1 U3556 ( .A1(n3563), .A2(n3562), .ZN(n3577) );
  AND2_X1 U3557 ( .A1(n3560), .A2(n3578), .ZN(n3576) );
  OR2_X1 U3558 ( .A1(n3562), .A2(n3563), .ZN(n3578) );
  OR2_X1 U3559 ( .A1(n2119), .A2(n2208), .ZN(n3563) );
  OR2_X1 U3560 ( .A1(n3579), .A2(n3580), .ZN(n3562) );
  AND2_X1 U3561 ( .A1(n3559), .A2(n3558), .ZN(n3580) );
  AND2_X1 U3562 ( .A1(n3556), .A2(n3581), .ZN(n3579) );
  OR2_X1 U3563 ( .A1(n3558), .A2(n3559), .ZN(n3581) );
  OR2_X1 U3564 ( .A1(n2213), .A2(n2208), .ZN(n3559) );
  OR2_X1 U3565 ( .A1(n3582), .A2(n3583), .ZN(n3558) );
  AND2_X1 U3566 ( .A1(n3555), .A2(n3554), .ZN(n3583) );
  AND2_X1 U3567 ( .A1(n3552), .A2(n3584), .ZN(n3582) );
  OR2_X1 U3568 ( .A1(n3554), .A2(n3555), .ZN(n3584) );
  OR2_X1 U3569 ( .A1(n2090), .A2(n2208), .ZN(n3555) );
  OR2_X1 U3570 ( .A1(n3585), .A2(n3586), .ZN(n3554) );
  AND2_X1 U3571 ( .A1(n3551), .A2(n3550), .ZN(n3586) );
  AND2_X1 U3572 ( .A1(n3548), .A2(n3587), .ZN(n3585) );
  OR2_X1 U3573 ( .A1(n3550), .A2(n3551), .ZN(n3587) );
  OR2_X1 U3574 ( .A1(n2219), .A2(n2208), .ZN(n3551) );
  OR2_X1 U3575 ( .A1(n3588), .A2(n3589), .ZN(n3550) );
  AND2_X1 U3576 ( .A1(n3544), .A2(n3547), .ZN(n3589) );
  AND2_X1 U3577 ( .A1(n3590), .A2(n3546), .ZN(n3588) );
  OR2_X1 U3578 ( .A1(n3591), .A2(n3592), .ZN(n3546) );
  AND2_X1 U3579 ( .A1(n3543), .A2(n3542), .ZN(n3592) );
  AND2_X1 U3580 ( .A1(n3540), .A2(n3593), .ZN(n3591) );
  OR2_X1 U3581 ( .A1(n3542), .A2(n3543), .ZN(n3593) );
  OR2_X1 U3582 ( .A1(n2225), .A2(n2208), .ZN(n3543) );
  OR2_X1 U3583 ( .A1(n3594), .A2(n3595), .ZN(n3542) );
  AND2_X1 U3584 ( .A1(n3536), .A2(n3539), .ZN(n3595) );
  AND2_X1 U3585 ( .A1(n3596), .A2(n3538), .ZN(n3594) );
  OR2_X1 U3586 ( .A1(n3597), .A2(n3598), .ZN(n3538) );
  AND2_X1 U3587 ( .A1(n3532), .A2(n3535), .ZN(n3598) );
  AND2_X1 U3588 ( .A1(n3599), .A2(n3534), .ZN(n3597) );
  OR2_X1 U3589 ( .A1(n3600), .A2(n3601), .ZN(n3534) );
  AND2_X1 U3590 ( .A1(n3528), .A2(n3531), .ZN(n3601) );
  AND2_X1 U3591 ( .A1(n3530), .A2(n3602), .ZN(n3600) );
  OR2_X1 U3592 ( .A1(n3531), .A2(n3528), .ZN(n3602) );
  OR2_X1 U3593 ( .A1(n2003), .A2(n2208), .ZN(n3528) );
  OR3_X1 U3594 ( .A1(n2550), .A2(n2208), .A3(n2157), .ZN(n3531) );
  INV_X1 U3595 ( .A(n3603), .ZN(n3530) );
  OR2_X1 U3596 ( .A1(n3604), .A2(n3605), .ZN(n3603) );
  AND2_X1 U3597 ( .A1(b_3_), .A2(n3606), .ZN(n3605) );
  OR2_X1 U3598 ( .A1(n3607), .A2(n1980), .ZN(n3606) );
  AND2_X1 U3599 ( .A1(a_14_), .A2(n2202), .ZN(n3607) );
  AND2_X1 U3600 ( .A1(b_2_), .A2(n3608), .ZN(n3604) );
  OR2_X1 U3601 ( .A1(n3609), .A2(n1983), .ZN(n3608) );
  AND2_X1 U3602 ( .A1(a_15_), .A2(n2157), .ZN(n3609) );
  OR2_X1 U3603 ( .A1(n3535), .A2(n3532), .ZN(n3599) );
  XNOR2_X1 U3604 ( .A(n3610), .B(n3611), .ZN(n3532) );
  XNOR2_X1 U3605 ( .A(n3612), .B(n3613), .ZN(n3611) );
  OR2_X1 U3606 ( .A1(n2231), .A2(n2208), .ZN(n3535) );
  OR2_X1 U3607 ( .A1(n3539), .A2(n3536), .ZN(n3596) );
  XOR2_X1 U3608 ( .A(n3614), .B(n3615), .Z(n3536) );
  XOR2_X1 U3609 ( .A(n3616), .B(n3617), .Z(n3615) );
  OR2_X1 U3610 ( .A1(n2032), .A2(n2208), .ZN(n3539) );
  XOR2_X1 U3611 ( .A(n3618), .B(n3619), .Z(n3540) );
  XOR2_X1 U3612 ( .A(n3620), .B(n3621), .Z(n3619) );
  OR2_X1 U3613 ( .A1(n3547), .A2(n3544), .ZN(n3590) );
  XOR2_X1 U3614 ( .A(n3622), .B(n3623), .Z(n3544) );
  XOR2_X1 U3615 ( .A(n3624), .B(n3625), .Z(n3623) );
  OR2_X1 U3616 ( .A1(n2061), .A2(n2208), .ZN(n3547) );
  INV_X1 U3617 ( .A(b_4_), .ZN(n2208) );
  XOR2_X1 U3618 ( .A(n3626), .B(n3627), .Z(n3548) );
  XOR2_X1 U3619 ( .A(n3628), .B(n3629), .Z(n3627) );
  XOR2_X1 U3620 ( .A(n3630), .B(n3631), .Z(n3552) );
  XOR2_X1 U3621 ( .A(n3632), .B(n3633), .Z(n3631) );
  XOR2_X1 U3622 ( .A(n3634), .B(n3635), .Z(n3556) );
  XOR2_X1 U3623 ( .A(n3636), .B(n3637), .Z(n3635) );
  XOR2_X1 U3624 ( .A(n3570), .B(n3638), .Z(n3560) );
  XOR2_X1 U3625 ( .A(n3569), .B(n3568), .Z(n3638) );
  OR2_X1 U3626 ( .A1(n2213), .A2(n2157), .ZN(n3568) );
  OR2_X1 U3627 ( .A1(n3639), .A2(n3640), .ZN(n3569) );
  AND2_X1 U3628 ( .A1(n3637), .A2(n3636), .ZN(n3640) );
  AND2_X1 U3629 ( .A1(n3634), .A2(n3641), .ZN(n3639) );
  OR2_X1 U3630 ( .A1(n3636), .A2(n3637), .ZN(n3641) );
  OR2_X1 U3631 ( .A1(n2090), .A2(n2157), .ZN(n3637) );
  OR2_X1 U3632 ( .A1(n3642), .A2(n3643), .ZN(n3636) );
  AND2_X1 U3633 ( .A1(n3633), .A2(n3632), .ZN(n3643) );
  AND2_X1 U3634 ( .A1(n3630), .A2(n3644), .ZN(n3642) );
  OR2_X1 U3635 ( .A1(n3632), .A2(n3633), .ZN(n3644) );
  OR2_X1 U3636 ( .A1(n2219), .A2(n2157), .ZN(n3633) );
  OR2_X1 U3637 ( .A1(n3645), .A2(n3646), .ZN(n3632) );
  AND2_X1 U3638 ( .A1(n3629), .A2(n3628), .ZN(n3646) );
  AND2_X1 U3639 ( .A1(n3626), .A2(n3647), .ZN(n3645) );
  OR2_X1 U3640 ( .A1(n3628), .A2(n3629), .ZN(n3647) );
  OR2_X1 U3641 ( .A1(n2061), .A2(n2157), .ZN(n3629) );
  OR2_X1 U3642 ( .A1(n3648), .A2(n3649), .ZN(n3628) );
  AND2_X1 U3643 ( .A1(n3622), .A2(n3625), .ZN(n3649) );
  AND2_X1 U3644 ( .A1(n3650), .A2(n3624), .ZN(n3648) );
  OR2_X1 U3645 ( .A1(n3651), .A2(n3652), .ZN(n3624) );
  AND2_X1 U3646 ( .A1(n3621), .A2(n3620), .ZN(n3652) );
  AND2_X1 U3647 ( .A1(n3618), .A2(n3653), .ZN(n3651) );
  OR2_X1 U3648 ( .A1(n3620), .A2(n3621), .ZN(n3653) );
  OR2_X1 U3649 ( .A1(n2032), .A2(n2157), .ZN(n3621) );
  OR2_X1 U3650 ( .A1(n3654), .A2(n3655), .ZN(n3620) );
  AND2_X1 U3651 ( .A1(n3614), .A2(n3617), .ZN(n3655) );
  AND2_X1 U3652 ( .A1(n3656), .A2(n3616), .ZN(n3654) );
  OR2_X1 U3653 ( .A1(n3657), .A2(n3658), .ZN(n3616) );
  AND2_X1 U3654 ( .A1(n3610), .A2(n3613), .ZN(n3658) );
  AND2_X1 U3655 ( .A1(n3612), .A2(n3659), .ZN(n3657) );
  OR2_X1 U3656 ( .A1(n3613), .A2(n3610), .ZN(n3659) );
  OR2_X1 U3657 ( .A1(n2003), .A2(n2157), .ZN(n3610) );
  OR3_X1 U3658 ( .A1(n2550), .A2(n2157), .A3(n2202), .ZN(n3613) );
  INV_X1 U3659 ( .A(n3660), .ZN(n3612) );
  OR2_X1 U3660 ( .A1(n3661), .A2(n3662), .ZN(n3660) );
  AND2_X1 U3661 ( .A1(b_2_), .A2(n3663), .ZN(n3662) );
  OR2_X1 U3662 ( .A1(n3664), .A2(n1980), .ZN(n3663) );
  AND2_X1 U3663 ( .A1(a_14_), .A2(n2186), .ZN(n3664) );
  AND2_X1 U3664 ( .A1(b_1_), .A2(n3665), .ZN(n3661) );
  OR2_X1 U3665 ( .A1(n3666), .A2(n1983), .ZN(n3665) );
  AND2_X1 U3666 ( .A1(a_15_), .A2(n2202), .ZN(n3666) );
  OR2_X1 U3667 ( .A1(n3617), .A2(n3614), .ZN(n3656) );
  XNOR2_X1 U3668 ( .A(n3667), .B(n3668), .ZN(n3614) );
  XNOR2_X1 U3669 ( .A(n3669), .B(n3670), .ZN(n3668) );
  OR2_X1 U3670 ( .A1(n2231), .A2(n2157), .ZN(n3617) );
  XOR2_X1 U3671 ( .A(n3671), .B(n3672), .Z(n3618) );
  XOR2_X1 U3672 ( .A(n3673), .B(n3674), .Z(n3672) );
  OR2_X1 U3673 ( .A1(n3625), .A2(n3622), .ZN(n3650) );
  XOR2_X1 U3674 ( .A(n3675), .B(n3676), .Z(n3622) );
  XOR2_X1 U3675 ( .A(n3677), .B(n3678), .Z(n3676) );
  OR2_X1 U3676 ( .A1(n2225), .A2(n2157), .ZN(n3625) );
  INV_X1 U3677 ( .A(b_3_), .ZN(n2157) );
  XOR2_X1 U3678 ( .A(n3679), .B(n3680), .Z(n3626) );
  XOR2_X1 U3679 ( .A(n3681), .B(n3682), .Z(n3680) );
  XOR2_X1 U3680 ( .A(n3683), .B(n3684), .Z(n3630) );
  XOR2_X1 U3681 ( .A(n3685), .B(n3686), .Z(n3684) );
  XOR2_X1 U3682 ( .A(n3687), .B(n3688), .Z(n3634) );
  XOR2_X1 U3683 ( .A(n3689), .B(n3690), .Z(n3688) );
  XOR2_X1 U3684 ( .A(n3691), .B(n3692), .Z(n3570) );
  XOR2_X1 U3685 ( .A(n3693), .B(n3694), .Z(n3692) );
  INV_X1 U3686 ( .A(n2131), .ZN(n2209) );
  AND2_X1 U3687 ( .A1(a_4_), .A2(b_4_), .ZN(n2131) );
  AND3_X1 U3688 ( .A1(n2140), .A2(n2138), .A3(n2139), .ZN(n2141) );
  INV_X1 U3689 ( .A(n2292), .ZN(n2139) );
  OR2_X1 U3690 ( .A1(n3695), .A2(n3696), .ZN(n2292) );
  AND2_X1 U3691 ( .A1(n2311), .A2(n2310), .ZN(n3696) );
  AND2_X1 U3692 ( .A1(n2308), .A2(n3697), .ZN(n3695) );
  OR2_X1 U3693 ( .A1(n2310), .A2(n2311), .ZN(n3697) );
  OR2_X1 U3694 ( .A1(n2202), .A2(n2291), .ZN(n2311) );
  OR2_X1 U3695 ( .A1(n3698), .A2(n3699), .ZN(n2310) );
  AND2_X1 U3696 ( .A1(n2328), .A2(n2327), .ZN(n3699) );
  AND2_X1 U3697 ( .A1(n2325), .A2(n3700), .ZN(n3698) );
  OR2_X1 U3698 ( .A1(n2327), .A2(n2328), .ZN(n3700) );
  OR2_X1 U3699 ( .A1(n2202), .A2(n2187), .ZN(n2328) );
  OR2_X1 U3700 ( .A1(n3701), .A2(n3702), .ZN(n2327) );
  AND2_X1 U3701 ( .A1(n2360), .A2(n2203), .ZN(n3702) );
  AND2_X1 U3702 ( .A1(n2359), .A2(n3703), .ZN(n3701) );
  OR2_X1 U3703 ( .A1(n2203), .A2(n2360), .ZN(n3703) );
  OR2_X1 U3704 ( .A1(n3704), .A2(n3705), .ZN(n2360) );
  AND2_X1 U3705 ( .A1(n2390), .A2(n2389), .ZN(n3705) );
  AND2_X1 U3706 ( .A1(n2387), .A2(n3706), .ZN(n3704) );
  OR2_X1 U3707 ( .A1(n2389), .A2(n2390), .ZN(n3706) );
  OR2_X1 U3708 ( .A1(n2158), .A2(n2202), .ZN(n2390) );
  OR2_X1 U3709 ( .A1(n3707), .A2(n3708), .ZN(n2389) );
  AND2_X1 U3710 ( .A1(n2437), .A2(n2436), .ZN(n3708) );
  AND2_X1 U3711 ( .A1(n2434), .A2(n3709), .ZN(n3707) );
  OR2_X1 U3712 ( .A1(n2436), .A2(n2437), .ZN(n3709) );
  OR2_X1 U3713 ( .A1(n2207), .A2(n2202), .ZN(n2437) );
  OR2_X1 U3714 ( .A1(n3710), .A2(n3711), .ZN(n2436) );
  AND2_X1 U3715 ( .A1(n2481), .A2(n2480), .ZN(n3711) );
  AND2_X1 U3716 ( .A1(n2478), .A2(n3712), .ZN(n3710) );
  OR2_X1 U3717 ( .A1(n2480), .A2(n2481), .ZN(n3712) );
  OR2_X1 U3718 ( .A1(n2119), .A2(n2202), .ZN(n2481) );
  OR2_X1 U3719 ( .A1(n3713), .A2(n3714), .ZN(n2480) );
  AND2_X1 U3720 ( .A1(n3575), .A2(n3574), .ZN(n3714) );
  AND2_X1 U3721 ( .A1(n3572), .A2(n3715), .ZN(n3713) );
  OR2_X1 U3722 ( .A1(n3574), .A2(n3575), .ZN(n3715) );
  OR2_X1 U3723 ( .A1(n2213), .A2(n2202), .ZN(n3575) );
  OR2_X1 U3724 ( .A1(n3716), .A2(n3717), .ZN(n3574) );
  AND2_X1 U3725 ( .A1(n3694), .A2(n3693), .ZN(n3717) );
  AND2_X1 U3726 ( .A1(n3691), .A2(n3718), .ZN(n3716) );
  OR2_X1 U3727 ( .A1(n3693), .A2(n3694), .ZN(n3718) );
  OR2_X1 U3728 ( .A1(n2090), .A2(n2202), .ZN(n3694) );
  OR2_X1 U3729 ( .A1(n3719), .A2(n3720), .ZN(n3693) );
  AND2_X1 U3730 ( .A1(n3690), .A2(n3689), .ZN(n3720) );
  AND2_X1 U3731 ( .A1(n3687), .A2(n3721), .ZN(n3719) );
  OR2_X1 U3732 ( .A1(n3689), .A2(n3690), .ZN(n3721) );
  OR2_X1 U3733 ( .A1(n2219), .A2(n2202), .ZN(n3690) );
  OR2_X1 U3734 ( .A1(n3722), .A2(n3723), .ZN(n3689) );
  AND2_X1 U3735 ( .A1(n3686), .A2(n3685), .ZN(n3723) );
  AND2_X1 U3736 ( .A1(n3683), .A2(n3724), .ZN(n3722) );
  OR2_X1 U3737 ( .A1(n3685), .A2(n3686), .ZN(n3724) );
  OR2_X1 U3738 ( .A1(n2061), .A2(n2202), .ZN(n3686) );
  OR2_X1 U3739 ( .A1(n3725), .A2(n3726), .ZN(n3685) );
  AND2_X1 U3740 ( .A1(n3682), .A2(n3681), .ZN(n3726) );
  AND2_X1 U3741 ( .A1(n3679), .A2(n3727), .ZN(n3725) );
  OR2_X1 U3742 ( .A1(n3681), .A2(n3682), .ZN(n3727) );
  OR2_X1 U3743 ( .A1(n2225), .A2(n2202), .ZN(n3682) );
  OR2_X1 U3744 ( .A1(n3728), .A2(n3729), .ZN(n3681) );
  AND2_X1 U3745 ( .A1(n3675), .A2(n3678), .ZN(n3729) );
  AND2_X1 U3746 ( .A1(n3730), .A2(n3677), .ZN(n3728) );
  OR2_X1 U3747 ( .A1(n3731), .A2(n3732), .ZN(n3677) );
  AND2_X1 U3748 ( .A1(n3674), .A2(n3673), .ZN(n3732) );
  AND2_X1 U3749 ( .A1(n3671), .A2(n3733), .ZN(n3731) );
  OR2_X1 U3750 ( .A1(n3673), .A2(n3674), .ZN(n3733) );
  OR2_X1 U3751 ( .A1(n2231), .A2(n2202), .ZN(n3674) );
  OR2_X1 U3752 ( .A1(n3734), .A2(n3735), .ZN(n3673) );
  AND2_X1 U3753 ( .A1(n3667), .A2(n3670), .ZN(n3735) );
  AND2_X1 U3754 ( .A1(n3669), .A2(n3736), .ZN(n3734) );
  OR2_X1 U3755 ( .A1(n3670), .A2(n3667), .ZN(n3736) );
  OR2_X1 U3756 ( .A1(n2003), .A2(n2202), .ZN(n3667) );
  OR3_X1 U3757 ( .A1(n2550), .A2(n2202), .A3(n2186), .ZN(n3670) );
  INV_X1 U3758 ( .A(n3737), .ZN(n3669) );
  OR2_X1 U3759 ( .A1(n3738), .A2(n3739), .ZN(n3737) );
  AND2_X1 U3760 ( .A1(b_1_), .A2(n3740), .ZN(n3739) );
  OR2_X1 U3761 ( .A1(n3741), .A2(n1980), .ZN(n3740) );
  AND2_X1 U3762 ( .A1(n2240), .A2(a_14_), .ZN(n1980) );
  AND2_X1 U3763 ( .A1(a_14_), .A2(n3742), .ZN(n3741) );
  AND2_X1 U3764 ( .A1(b_0_), .A2(n3743), .ZN(n3738) );
  OR2_X1 U3765 ( .A1(n3744), .A2(n1983), .ZN(n3743) );
  AND2_X1 U3766 ( .A1(n2239), .A2(a_15_), .ZN(n1983) );
  AND2_X1 U3767 ( .A1(a_15_), .A2(n2186), .ZN(n3744) );
  XNOR2_X1 U3768 ( .A(n3745), .B(n3746), .ZN(n3671) );
  OR2_X1 U3769 ( .A1(n3747), .A2(n3748), .ZN(n3745) );
  INV_X1 U3770 ( .A(n3749), .ZN(n3748) );
  AND2_X1 U3771 ( .A1(n3750), .A2(n3751), .ZN(n3747) );
  OR2_X1 U3772 ( .A1(n2239), .A2(n3742), .ZN(n3750) );
  OR2_X1 U3773 ( .A1(n3678), .A2(n3675), .ZN(n3730) );
  XOR2_X1 U3774 ( .A(n3752), .B(n3753), .Z(n3675) );
  XOR2_X1 U3775 ( .A(n3754), .B(n3755), .Z(n3752) );
  OR2_X1 U3776 ( .A1(n2032), .A2(n2202), .ZN(n3678) );
  INV_X1 U3777 ( .A(b_2_), .ZN(n2202) );
  XNOR2_X1 U3778 ( .A(n3756), .B(n3757), .ZN(n3679) );
  XNOR2_X1 U3779 ( .A(n3758), .B(n3759), .ZN(n3756) );
  XNOR2_X1 U3780 ( .A(n3760), .B(n3761), .ZN(n3683) );
  XNOR2_X1 U3781 ( .A(n3762), .B(n3763), .ZN(n3760) );
  XNOR2_X1 U3782 ( .A(n3764), .B(n3765), .ZN(n3687) );
  XNOR2_X1 U3783 ( .A(n3766), .B(n3767), .ZN(n3764) );
  XOR2_X1 U3784 ( .A(n3768), .B(n3769), .Z(n3691) );
  XOR2_X1 U3785 ( .A(n3770), .B(n3771), .Z(n3769) );
  XOR2_X1 U3786 ( .A(n3772), .B(n3773), .Z(n3572) );
  XOR2_X1 U3787 ( .A(n3774), .B(n3775), .Z(n3773) );
  XOR2_X1 U3788 ( .A(n3776), .B(n3777), .Z(n2478) );
  XOR2_X1 U3789 ( .A(n3778), .B(n3779), .Z(n3777) );
  XOR2_X1 U3790 ( .A(n3780), .B(n3781), .Z(n2434) );
  XOR2_X1 U3791 ( .A(n3782), .B(n3783), .Z(n3781) );
  XOR2_X1 U3792 ( .A(n3784), .B(n3785), .Z(n2387) );
  XOR2_X1 U3793 ( .A(n3786), .B(n3787), .Z(n3785) );
  INV_X1 U3794 ( .A(n2170), .ZN(n2203) );
  AND2_X1 U3795 ( .A1(a_2_), .A2(b_2_), .ZN(n2170) );
  XOR2_X1 U3796 ( .A(n3788), .B(n3789), .Z(n2359) );
  XOR2_X1 U3797 ( .A(n3790), .B(n3791), .Z(n3789) );
  XOR2_X1 U3798 ( .A(n3792), .B(n3793), .Z(n2325) );
  XOR2_X1 U3799 ( .A(n3794), .B(n3795), .Z(n3793) );
  XOR2_X1 U3800 ( .A(n3796), .B(n3797), .Z(n2308) );
  XOR2_X1 U3801 ( .A(n3798), .B(n2184), .Z(n3797) );
  XOR2_X1 U3802 ( .A(n3799), .B(n2290), .Z(n2138) );
  OR2_X1 U3803 ( .A1(n3800), .A2(n3801), .ZN(n2290) );
  AND2_X1 U3804 ( .A1(n3802), .A2(n3803), .ZN(n3801) );
  AND2_X1 U3805 ( .A1(n3804), .A2(n3805), .ZN(n3800) );
  OR2_X1 U3806 ( .A1(n3803), .A2(n3802), .ZN(n3804) );
  OR2_X1 U3807 ( .A1(n2291), .A2(n3742), .ZN(n3799) );
  XNOR2_X1 U3808 ( .A(n3802), .B(n3806), .ZN(n2140) );
  XOR2_X1 U3809 ( .A(n3803), .B(n3805), .Z(n3806) );
  OR2_X1 U3810 ( .A1(n2186), .A2(n2291), .ZN(n3805) );
  INV_X1 U3811 ( .A(a_0_), .ZN(n2291) );
  OR2_X1 U3812 ( .A1(n3807), .A2(n3808), .ZN(n3803) );
  AND2_X1 U3813 ( .A1(n3796), .A2(n3798), .ZN(n3808) );
  AND2_X1 U3814 ( .A1(n3809), .A2(n2184), .ZN(n3807) );
  OR2_X1 U3815 ( .A1(n2187), .A2(n2186), .ZN(n2184) );
  OR2_X1 U3816 ( .A1(n3798), .A2(n3796), .ZN(n3809) );
  OR2_X1 U3817 ( .A1(n2201), .A2(n3742), .ZN(n3796) );
  OR2_X1 U3818 ( .A1(n3810), .A2(n3811), .ZN(n3798) );
  AND2_X1 U3819 ( .A1(n3792), .A2(n3794), .ZN(n3811) );
  AND2_X1 U3820 ( .A1(n3812), .A2(n3795), .ZN(n3810) );
  OR2_X1 U3821 ( .A1(n2158), .A2(n3742), .ZN(n3795) );
  OR2_X1 U3822 ( .A1(n3794), .A2(n3792), .ZN(n3812) );
  OR2_X1 U3823 ( .A1(n2201), .A2(n2186), .ZN(n3792) );
  INV_X1 U3824 ( .A(a_2_), .ZN(n2201) );
  OR2_X1 U3825 ( .A1(n3813), .A2(n3814), .ZN(n3794) );
  AND2_X1 U3826 ( .A1(n3788), .A2(n3790), .ZN(n3814) );
  AND2_X1 U3827 ( .A1(n3815), .A2(n3791), .ZN(n3813) );
  OR2_X1 U3828 ( .A1(n2207), .A2(n3742), .ZN(n3791) );
  OR2_X1 U3829 ( .A1(n3790), .A2(n3788), .ZN(n3815) );
  OR2_X1 U3830 ( .A1(n2158), .A2(n2186), .ZN(n3788) );
  INV_X1 U3831 ( .A(a_3_), .ZN(n2158) );
  OR2_X1 U3832 ( .A1(n3816), .A2(n3817), .ZN(n3790) );
  AND2_X1 U3833 ( .A1(n3784), .A2(n3786), .ZN(n3817) );
  AND2_X1 U3834 ( .A1(n3818), .A2(n3787), .ZN(n3816) );
  OR2_X1 U3835 ( .A1(n2119), .A2(n3742), .ZN(n3787) );
  OR2_X1 U3836 ( .A1(n3786), .A2(n3784), .ZN(n3818) );
  OR2_X1 U3837 ( .A1(n2207), .A2(n2186), .ZN(n3784) );
  INV_X1 U3838 ( .A(a_4_), .ZN(n2207) );
  OR2_X1 U3839 ( .A1(n3819), .A2(n3820), .ZN(n3786) );
  AND2_X1 U3840 ( .A1(n3780), .A2(n3782), .ZN(n3820) );
  AND2_X1 U3841 ( .A1(n3821), .A2(n3783), .ZN(n3819) );
  OR2_X1 U3842 ( .A1(n2213), .A2(n3742), .ZN(n3783) );
  OR2_X1 U3843 ( .A1(n3782), .A2(n3780), .ZN(n3821) );
  OR2_X1 U3844 ( .A1(n2119), .A2(n2186), .ZN(n3780) );
  INV_X1 U3845 ( .A(a_5_), .ZN(n2119) );
  OR2_X1 U3846 ( .A1(n3822), .A2(n3823), .ZN(n3782) );
  AND2_X1 U3847 ( .A1(n3776), .A2(n3778), .ZN(n3823) );
  AND2_X1 U3848 ( .A1(n3824), .A2(n3779), .ZN(n3822) );
  OR2_X1 U3849 ( .A1(n2090), .A2(n3742), .ZN(n3779) );
  OR2_X1 U3850 ( .A1(n3778), .A2(n3776), .ZN(n3824) );
  OR2_X1 U3851 ( .A1(n2213), .A2(n2186), .ZN(n3776) );
  INV_X1 U3852 ( .A(a_6_), .ZN(n2213) );
  OR2_X1 U3853 ( .A1(n3825), .A2(n3826), .ZN(n3778) );
  AND2_X1 U3854 ( .A1(n3772), .A2(n3774), .ZN(n3826) );
  AND2_X1 U3855 ( .A1(n3827), .A2(n3775), .ZN(n3825) );
  OR2_X1 U3856 ( .A1(n2219), .A2(n3742), .ZN(n3775) );
  OR2_X1 U3857 ( .A1(n3774), .A2(n3772), .ZN(n3827) );
  OR2_X1 U3858 ( .A1(n2090), .A2(n2186), .ZN(n3772) );
  INV_X1 U3859 ( .A(a_7_), .ZN(n2090) );
  OR2_X1 U3860 ( .A1(n3828), .A2(n3829), .ZN(n3774) );
  AND2_X1 U3861 ( .A1(n3768), .A2(n3770), .ZN(n3829) );
  AND2_X1 U3862 ( .A1(n3830), .A2(n3771), .ZN(n3828) );
  OR2_X1 U3863 ( .A1(n2061), .A2(n3742), .ZN(n3771) );
  OR2_X1 U3864 ( .A1(n3770), .A2(n3768), .ZN(n3830) );
  OR2_X1 U3865 ( .A1(n2219), .A2(n2186), .ZN(n3768) );
  INV_X1 U3866 ( .A(a_8_), .ZN(n2219) );
  OR2_X1 U3867 ( .A1(n3831), .A2(n3832), .ZN(n3770) );
  AND2_X1 U3868 ( .A1(n3765), .A2(n3767), .ZN(n3832) );
  AND2_X1 U3869 ( .A1(n3833), .A2(n3766), .ZN(n3831) );
  OR2_X1 U3870 ( .A1(n2225), .A2(n3742), .ZN(n3766) );
  OR2_X1 U3871 ( .A1(n3767), .A2(n3765), .ZN(n3833) );
  OR2_X1 U3872 ( .A1(n2061), .A2(n2186), .ZN(n3765) );
  INV_X1 U3873 ( .A(a_9_), .ZN(n2061) );
  OR2_X1 U3874 ( .A1(n3834), .A2(n3835), .ZN(n3767) );
  AND2_X1 U3875 ( .A1(n3761), .A2(n3763), .ZN(n3835) );
  AND2_X1 U3876 ( .A1(n3836), .A2(n3762), .ZN(n3834) );
  OR2_X1 U3877 ( .A1(n2032), .A2(n3742), .ZN(n3762) );
  OR2_X1 U3878 ( .A1(n3763), .A2(n3761), .ZN(n3836) );
  OR2_X1 U3879 ( .A1(n2225), .A2(n2186), .ZN(n3761) );
  INV_X1 U3880 ( .A(a_10_), .ZN(n2225) );
  OR2_X1 U3881 ( .A1(n3837), .A2(n3838), .ZN(n3763) );
  AND2_X1 U3882 ( .A1(n3757), .A2(n3759), .ZN(n3838) );
  AND2_X1 U3883 ( .A1(n3839), .A2(n3758), .ZN(n3837) );
  OR2_X1 U3884 ( .A1(n2231), .A2(n3742), .ZN(n3758) );
  OR2_X1 U3885 ( .A1(n3759), .A2(n3757), .ZN(n3839) );
  OR2_X1 U3886 ( .A1(n2032), .A2(n2186), .ZN(n3757) );
  INV_X1 U3887 ( .A(a_11_), .ZN(n2032) );
  OR2_X1 U3888 ( .A1(n3840), .A2(n3841), .ZN(n3759) );
  AND2_X1 U3889 ( .A1(n3753), .A2(n3755), .ZN(n3841) );
  AND2_X1 U3890 ( .A1(n3754), .A2(n3842), .ZN(n3840) );
  OR2_X1 U3891 ( .A1(n3755), .A2(n3753), .ZN(n3842) );
  OR2_X1 U3892 ( .A1(n2231), .A2(n2186), .ZN(n3753) );
  INV_X1 U3893 ( .A(a_12_), .ZN(n2231) );
  OR2_X1 U3894 ( .A1(n2003), .A2(n3742), .ZN(n3755) );
  AND2_X1 U3895 ( .A1(n3749), .A2(n3746), .ZN(n3754) );
  OR3_X1 U3896 ( .A1(n2550), .A2(n2186), .A3(n3742), .ZN(n3746) );
  OR2_X1 U3897 ( .A1(n2240), .A2(n2239), .ZN(n2550) );
  INV_X1 U3898 ( .A(a_15_), .ZN(n2240) );
  OR3_X1 U3899 ( .A1(n2239), .A2(n3742), .A3(n3751), .ZN(n3749) );
  OR2_X1 U3900 ( .A1(n2003), .A2(n2186), .ZN(n3751) );
  INV_X1 U3901 ( .A(b_1_), .ZN(n2186) );
  INV_X1 U3902 ( .A(a_13_), .ZN(n2003) );
  INV_X1 U3903 ( .A(a_14_), .ZN(n2239) );
  OR2_X1 U3904 ( .A1(n2187), .A2(n3742), .ZN(n3802) );
  INV_X1 U3905 ( .A(b_0_), .ZN(n3742) );
  INV_X1 U3906 ( .A(a_1_), .ZN(n2187) );
endmodule

