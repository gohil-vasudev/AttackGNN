module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n595_, new_n614_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n439_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n170_, new_n246_, new_n682_, new_n812_, new_n679_, new_n266_, new_n667_, new_n367_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n602_, new_n114_, new_n188_, new_n240_, new_n660_, new_n413_, new_n695_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n649_, new_n678_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n735_, new_n500_, new_n786_, new_n799_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n742_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n774_, new_n157_, new_n716_, new_n153_, new_n701_, new_n792_, new_n133_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n766_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n110_, new_n315_, new_n685_, new_n124_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n796_, new_n248_, new_n350_, new_n117_, new_n655_, new_n630_, new_n759_, new_n167_, new_n385_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n764_, new_n150_, new_n683_, new_n108_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n622_, new_n629_, new_n702_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n158_, new_n763_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n816_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n650_, new_n708_, new_n750_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n506_, new_n680_, new_n256_, new_n778_, new_n452_, new_n381_, new_n656_, new_n771_, new_n388_, new_n508_, new_n714_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n657_, new_n652_, new_n314_, new_n582_, new_n118_, new_n363_, new_n165_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n790_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n805_, new_n559_, new_n762_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n794_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n688_, new_n155_, new_n384_, new_n410_, new_n543_, new_n113_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n809_, new_n654_, new_n713_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n130_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n138_, new_n749_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n562_, new_n578_, new_n126_, new_n808_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n800_, new_n379_, new_n719_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n143_, new_n520_, new_n125_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n237_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n748_, new_n182_, new_n407_, new_n666_, new_n813_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n191_, new_n755_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n112_, new_n121_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n782_, new_n354_, new_n444_, new_n518_, new_n737_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n801_, new_n789_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n662_, new_n440_, new_n733_, new_n122_, new_n531_, new_n593_, new_n111_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n115_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n134_, new_n769_, new_n651_, new_n433_, new_n435_, new_n109_, new_n776_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n815_, new_n278_, new_n304_, new_n523_, new_n638_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n129_, new_n711_, new_n644_, new_n731_, new_n599_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n196_, new_n818_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n754_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n803_, new_n330_, new_n727_, new_n375_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n791_, new_n357_, new_n320_, new_n780_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n128_, new_n358_, new_n348_, new_n610_, new_n159_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n802_, new_n697_, new_n185_, new_n709_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n120_, new_n521_, new_n793_, new_n406_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n135_, new_n573_, new_n765_, new_n405_;

or g000 ( new_n108_, keyIn_0_5, N89 );
not g001 ( new_n109_, N95 );
and g002 ( new_n110_, keyIn_0_5, N89 );
or g003 ( new_n111_, new_n110_, new_n109_ );
not g004 ( new_n112_, new_n111_ );
and g005 ( new_n113_, new_n112_, new_n108_ );
not g006 ( new_n114_, keyIn_0_9 );
not g007 ( new_n115_, N69 );
or g008 ( new_n116_, new_n115_, N63 );
and g009 ( new_n117_, new_n116_, new_n114_ );
not g010 ( new_n118_, N63 );
and g011 ( new_n119_, new_n118_, keyIn_0_9 );
and g012 ( new_n120_, new_n119_, N69 );
or g013 ( new_n121_, new_n117_, new_n120_ );
not g014 ( new_n122_, keyIn_0_8 );
not g015 ( new_n123_, N24 );
and g016 ( new_n124_, new_n123_, N30 );
or g017 ( new_n125_, new_n124_, new_n122_ );
not g018 ( new_n126_, N30 );
or g019 ( new_n127_, keyIn_0_8, N24 );
or g020 ( new_n128_, new_n127_, new_n126_ );
and g021 ( new_n129_, new_n125_, new_n128_ );
or g022 ( new_n130_, new_n121_, new_n129_ );
or g023 ( new_n131_, new_n130_, new_n113_ );
not g024 ( new_n132_, keyIn_0_10 );
not g025 ( new_n133_, N108 );
or g026 ( new_n134_, new_n133_, N102 );
and g027 ( new_n135_, new_n134_, new_n132_ );
not g028 ( new_n136_, N102 );
and g029 ( new_n137_, new_n136_, keyIn_0_10 );
and g030 ( new_n138_, new_n137_, N108 );
or g031 ( new_n139_, new_n135_, new_n138_ );
not g032 ( new_n140_, N50 );
and g033 ( new_n141_, new_n140_, N56 );
not g034 ( new_n142_, N76 );
and g035 ( new_n143_, new_n142_, N82 );
not g036 ( new_n144_, N1 );
and g037 ( new_n145_, new_n144_, N4 );
or g038 ( new_n146_, new_n143_, new_n145_ );
or g039 ( new_n147_, new_n146_, new_n141_ );
or g040 ( new_n148_, new_n147_, new_n139_ );
not g041 ( new_n149_, N17 );
not g042 ( new_n150_, keyIn_0_7 );
or g043 ( new_n151_, new_n150_, N11 );
or g044 ( new_n152_, new_n151_, new_n149_ );
not g045 ( new_n153_, N11 );
and g046 ( new_n154_, new_n153_, N17 );
or g047 ( new_n155_, new_n154_, keyIn_0_7 );
and g048 ( new_n156_, new_n152_, new_n155_ );
not g049 ( new_n157_, keyIn_0_2 );
not g050 ( new_n158_, N37 );
and g051 ( new_n159_, new_n157_, new_n158_ );
and g052 ( new_n160_, keyIn_0_2, N37 );
or g053 ( new_n161_, new_n159_, new_n160_ );
and g054 ( new_n162_, new_n161_, N43 );
or g055 ( new_n163_, new_n156_, new_n162_ );
or g056 ( new_n164_, new_n148_, new_n163_ );
or g057 ( new_n165_, new_n164_, new_n131_ );
and g058 ( new_n166_, new_n165_, keyIn_0_20 );
not g059 ( new_n167_, keyIn_0_20 );
not g060 ( new_n168_, new_n113_ );
and g061 ( new_n169_, new_n118_, N69 );
or g062 ( new_n170_, new_n169_, keyIn_0_9 );
or g063 ( new_n171_, new_n114_, N63 );
or g064 ( new_n172_, new_n171_, new_n115_ );
and g065 ( new_n173_, new_n172_, new_n170_ );
or g066 ( new_n174_, new_n126_, N24 );
and g067 ( new_n175_, new_n174_, keyIn_0_8 );
and g068 ( new_n176_, new_n122_, new_n123_ );
and g069 ( new_n177_, new_n176_, N30 );
or g070 ( new_n178_, new_n175_, new_n177_ );
and g071 ( new_n179_, new_n178_, new_n173_ );
and g072 ( new_n180_, new_n179_, new_n168_ );
and g073 ( new_n181_, new_n136_, N108 );
or g074 ( new_n182_, new_n181_, keyIn_0_10 );
or g075 ( new_n183_, new_n132_, N102 );
or g076 ( new_n184_, new_n183_, new_n133_ );
and g077 ( new_n185_, new_n184_, new_n182_ );
not g078 ( new_n186_, new_n141_ );
not g079 ( new_n187_, N82 );
or g080 ( new_n188_, new_n187_, N76 );
not g081 ( new_n189_, N4 );
or g082 ( new_n190_, new_n189_, N1 );
and g083 ( new_n191_, new_n188_, new_n190_ );
and g084 ( new_n192_, new_n191_, new_n186_ );
and g085 ( new_n193_, new_n185_, new_n192_ );
and g086 ( new_n194_, new_n153_, keyIn_0_7 );
and g087 ( new_n195_, new_n194_, N17 );
or g088 ( new_n196_, new_n149_, N11 );
and g089 ( new_n197_, new_n196_, new_n150_ );
or g090 ( new_n198_, new_n197_, new_n195_ );
not g091 ( new_n199_, N43 );
or g092 ( new_n200_, keyIn_0_2, N37 );
not g093 ( new_n201_, new_n160_ );
and g094 ( new_n202_, new_n201_, new_n200_ );
or g095 ( new_n203_, new_n202_, new_n199_ );
and g096 ( new_n204_, new_n198_, new_n203_ );
and g097 ( new_n205_, new_n204_, new_n193_ );
and g098 ( new_n206_, new_n180_, new_n205_ );
and g099 ( new_n207_, new_n206_, new_n167_ );
or g100 ( N223, new_n166_, new_n207_ );
not g101 ( new_n209_, keyIn_0_21 );
and g102 ( new_n210_, new_n165_, keyIn_0_18 );
not g103 ( new_n211_, keyIn_0_18 );
and g104 ( new_n212_, new_n206_, new_n211_ );
or g105 ( new_n213_, new_n210_, new_n212_ );
and g106 ( new_n214_, new_n213_, new_n198_ );
or g107 ( new_n215_, new_n206_, new_n211_ );
not g108 ( new_n216_, new_n212_ );
and g109 ( new_n217_, new_n216_, new_n215_ );
and g110 ( new_n218_, new_n217_, new_n156_ );
or g111 ( new_n219_, new_n214_, new_n218_ );
and g112 ( new_n220_, new_n219_, new_n209_ );
or g113 ( new_n221_, new_n217_, new_n156_ );
or g114 ( new_n222_, new_n213_, new_n198_ );
and g115 ( new_n223_, new_n222_, new_n221_ );
and g116 ( new_n224_, new_n223_, keyIn_0_21 );
or g117 ( new_n225_, new_n220_, new_n224_ );
not g118 ( new_n226_, N21 );
and g119 ( new_n227_, new_n226_, N17 );
not g120 ( new_n228_, new_n227_ );
or g121 ( new_n229_, new_n225_, new_n228_ );
or g122 ( new_n230_, new_n229_, keyIn_0_29 );
not g123 ( new_n231_, keyIn_0_29 );
or g124 ( new_n232_, new_n223_, keyIn_0_21 );
or g125 ( new_n233_, new_n219_, new_n209_ );
and g126 ( new_n234_, new_n233_, new_n232_ );
and g127 ( new_n235_, new_n234_, new_n227_ );
or g128 ( new_n236_, new_n235_, new_n231_ );
and g129 ( new_n237_, new_n230_, new_n236_ );
and g130 ( new_n238_, new_n213_, new_n185_ );
and g131 ( new_n239_, new_n217_, new_n139_ );
or g132 ( new_n240_, new_n238_, new_n239_ );
not g133 ( new_n241_, N112 );
and g134 ( new_n242_, new_n241_, N108 );
and g135 ( new_n243_, new_n242_, keyIn_0_17 );
not g136 ( new_n244_, new_n243_ );
or g137 ( new_n245_, new_n242_, keyIn_0_17 );
and g138 ( new_n246_, new_n244_, new_n245_ );
not g139 ( new_n247_, new_n246_ );
and g140 ( new_n248_, new_n240_, new_n247_ );
not g141 ( new_n249_, new_n248_ );
and g142 ( new_n250_, new_n213_, new_n168_ );
and g143 ( new_n251_, new_n113_, new_n211_ );
or g144 ( new_n252_, new_n250_, new_n251_ );
not g145 ( new_n253_, N99 );
and g146 ( new_n254_, new_n253_, N95 );
and g147 ( new_n255_, new_n252_, new_n254_ );
not g148 ( new_n256_, new_n255_ );
and g149 ( new_n257_, new_n249_, new_n256_ );
not g150 ( new_n258_, new_n257_ );
and g151 ( new_n259_, new_n213_, new_n186_ );
and g152 ( new_n260_, new_n217_, new_n141_ );
or g153 ( new_n261_, new_n259_, new_n260_ );
not g154 ( new_n262_, keyIn_0_13 );
not g155 ( new_n263_, N60 );
and g156 ( new_n264_, new_n263_, N56 );
and g157 ( new_n265_, new_n264_, new_n262_ );
not g158 ( new_n266_, new_n265_ );
or g159 ( new_n267_, new_n264_, new_n262_ );
and g160 ( new_n268_, new_n266_, new_n267_ );
not g161 ( new_n269_, new_n268_ );
and g162 ( new_n270_, new_n261_, new_n269_ );
and g163 ( new_n271_, new_n213_, new_n178_ );
and g164 ( new_n272_, new_n129_, new_n211_ );
or g165 ( new_n273_, new_n271_, new_n272_ );
not g166 ( new_n274_, N34 );
and g167 ( new_n275_, new_n126_, keyIn_0_1 );
not g168 ( new_n276_, new_n275_ );
or g169 ( new_n277_, new_n126_, keyIn_0_1 );
and g170 ( new_n278_, new_n276_, new_n277_ );
and g171 ( new_n279_, new_n278_, new_n274_ );
and g172 ( new_n280_, new_n273_, new_n279_ );
or g173 ( new_n281_, new_n270_, new_n280_ );
and g174 ( new_n282_, new_n213_, new_n188_ );
and g175 ( new_n283_, new_n217_, new_n143_ );
or g176 ( new_n284_, new_n282_, new_n283_ );
not g177 ( new_n285_, N86 );
and g178 ( new_n286_, new_n285_, N82 );
and g179 ( new_n287_, new_n284_, new_n286_ );
and g180 ( new_n288_, new_n213_, new_n173_ );
and g181 ( new_n289_, new_n217_, new_n121_ );
or g182 ( new_n290_, new_n288_, new_n289_ );
not g183 ( new_n291_, N73 );
and g184 ( new_n292_, keyIn_0_4, N69 );
not g185 ( new_n293_, new_n292_ );
or g186 ( new_n294_, keyIn_0_4, N69 );
and g187 ( new_n295_, new_n293_, new_n294_ );
not g188 ( new_n296_, new_n295_ );
and g189 ( new_n297_, new_n296_, new_n291_ );
and g190 ( new_n298_, new_n290_, new_n297_ );
or g191 ( new_n299_, new_n287_, new_n298_ );
or g192 ( new_n300_, new_n299_, new_n281_ );
or g193 ( new_n301_, new_n300_, new_n258_ );
not g194 ( new_n302_, keyIn_0_27 );
or g195 ( new_n303_, new_n213_, new_n190_ );
or g196 ( new_n304_, new_n217_, new_n145_ );
and g197 ( new_n305_, new_n303_, new_n304_ );
not g198 ( new_n306_, keyIn_0_6 );
not g199 ( new_n307_, N8 );
and g200 ( new_n308_, new_n189_, keyIn_0_0 );
not g201 ( new_n309_, new_n308_ );
or g202 ( new_n310_, new_n189_, keyIn_0_0 );
and g203 ( new_n311_, new_n309_, new_n310_ );
not g204 ( new_n312_, new_n311_ );
and g205 ( new_n313_, new_n312_, new_n307_ );
not g206 ( new_n314_, new_n313_ );
and g207 ( new_n315_, new_n314_, new_n306_ );
and g208 ( new_n316_, new_n313_, keyIn_0_6 );
or g209 ( new_n317_, new_n315_, new_n316_ );
not g210 ( new_n318_, new_n317_ );
or g211 ( new_n319_, new_n305_, new_n318_ );
or g212 ( new_n320_, new_n319_, new_n302_ );
and g213 ( new_n321_, new_n217_, new_n145_ );
and g214 ( new_n322_, new_n213_, new_n190_ );
or g215 ( new_n323_, new_n322_, new_n321_ );
and g216 ( new_n324_, new_n323_, new_n317_ );
or g217 ( new_n325_, new_n324_, keyIn_0_27 );
and g218 ( new_n326_, new_n320_, new_n325_ );
not g219 ( new_n327_, keyIn_0_30 );
or g220 ( new_n328_, new_n213_, new_n203_ );
or g221 ( new_n329_, new_n217_, new_n162_ );
and g222 ( new_n330_, new_n328_, new_n329_ );
not g223 ( new_n331_, keyIn_0_12 );
not g224 ( new_n332_, N47 );
and g225 ( new_n333_, new_n199_, keyIn_0_3 );
not g226 ( new_n334_, new_n333_ );
or g227 ( new_n335_, new_n199_, keyIn_0_3 );
and g228 ( new_n336_, new_n334_, new_n335_ );
not g229 ( new_n337_, new_n336_ );
and g230 ( new_n338_, new_n337_, new_n332_ );
not g231 ( new_n339_, new_n338_ );
and g232 ( new_n340_, new_n339_, new_n331_ );
and g233 ( new_n341_, new_n338_, keyIn_0_12 );
or g234 ( new_n342_, new_n340_, new_n341_ );
not g235 ( new_n343_, new_n342_ );
or g236 ( new_n344_, new_n330_, new_n343_ );
or g237 ( new_n345_, new_n344_, new_n327_ );
and g238 ( new_n346_, new_n217_, new_n162_ );
and g239 ( new_n347_, new_n213_, new_n203_ );
or g240 ( new_n348_, new_n347_, new_n346_ );
and g241 ( new_n349_, new_n348_, new_n342_ );
or g242 ( new_n350_, new_n349_, keyIn_0_30 );
and g243 ( new_n351_, new_n345_, new_n350_ );
or g244 ( new_n352_, new_n326_, new_n351_ );
or g245 ( new_n353_, new_n301_, new_n352_ );
or g246 ( new_n354_, new_n353_, new_n237_ );
or g247 ( new_n355_, new_n354_, keyIn_0_32 );
not g248 ( new_n356_, keyIn_0_32 );
and g249 ( new_n357_, new_n235_, new_n231_ );
and g250 ( new_n358_, new_n229_, keyIn_0_29 );
or g251 ( new_n359_, new_n358_, new_n357_ );
not g252 ( new_n360_, new_n259_ );
not g253 ( new_n361_, new_n260_ );
and g254 ( new_n362_, new_n360_, new_n361_ );
or g255 ( new_n363_, new_n362_, new_n268_ );
not g256 ( new_n364_, new_n280_ );
and g257 ( new_n365_, new_n363_, new_n364_ );
not g258 ( new_n366_, new_n287_ );
not g259 ( new_n367_, new_n288_ );
not g260 ( new_n368_, new_n289_ );
and g261 ( new_n369_, new_n367_, new_n368_ );
not g262 ( new_n370_, new_n297_ );
or g263 ( new_n371_, new_n369_, new_n370_ );
and g264 ( new_n372_, new_n366_, new_n371_ );
and g265 ( new_n373_, new_n372_, new_n365_ );
and g266 ( new_n374_, new_n373_, new_n257_ );
and g267 ( new_n375_, new_n324_, keyIn_0_27 );
and g268 ( new_n376_, new_n319_, new_n302_ );
or g269 ( new_n377_, new_n376_, new_n375_ );
and g270 ( new_n378_, new_n349_, keyIn_0_30 );
and g271 ( new_n379_, new_n344_, new_n327_ );
or g272 ( new_n380_, new_n379_, new_n378_ );
and g273 ( new_n381_, new_n377_, new_n380_ );
and g274 ( new_n382_, new_n374_, new_n381_ );
and g275 ( new_n383_, new_n382_, new_n359_ );
or g276 ( new_n384_, new_n383_, new_n356_ );
and g277 ( new_n385_, new_n355_, new_n384_ );
and g278 ( new_n386_, new_n385_, keyIn_0_38 );
not g279 ( new_n387_, keyIn_0_38 );
and g280 ( new_n388_, new_n383_, new_n356_ );
and g281 ( new_n389_, new_n354_, keyIn_0_32 );
or g282 ( new_n390_, new_n389_, new_n388_ );
and g283 ( new_n391_, new_n390_, new_n387_ );
or g284 ( N329, new_n386_, new_n391_ );
not g285 ( new_n393_, keyIn_0_48 );
not g286 ( new_n394_, keyIn_0_42 );
and g287 ( new_n395_, new_n385_, keyIn_0_37 );
not g288 ( new_n396_, keyIn_0_37 );
and g289 ( new_n397_, new_n390_, new_n396_ );
or g290 ( new_n398_, new_n395_, new_n397_ );
and g291 ( new_n399_, new_n398_, new_n371_ );
or g292 ( new_n400_, new_n390_, new_n396_ );
or g293 ( new_n401_, new_n385_, keyIn_0_37 );
and g294 ( new_n402_, new_n400_, new_n401_ );
and g295 ( new_n403_, new_n402_, new_n298_ );
or g296 ( new_n404_, new_n399_, new_n403_ );
or g297 ( new_n405_, new_n404_, new_n394_ );
or g298 ( new_n406_, new_n402_, new_n298_ );
or g299 ( new_n407_, new_n398_, new_n371_ );
and g300 ( new_n408_, new_n407_, new_n406_ );
or g301 ( new_n409_, new_n408_, keyIn_0_42 );
and g302 ( new_n410_, new_n405_, new_n409_ );
not g303 ( new_n411_, keyIn_0_14 );
not g304 ( new_n412_, N79 );
and g305 ( new_n413_, new_n296_, new_n412_ );
and g306 ( new_n414_, new_n413_, new_n411_ );
not g307 ( new_n415_, new_n414_ );
or g308 ( new_n416_, new_n413_, new_n411_ );
and g309 ( new_n417_, new_n415_, new_n416_ );
or g310 ( new_n418_, new_n369_, new_n417_ );
and g311 ( new_n419_, new_n418_, keyIn_0_35 );
not g312 ( new_n420_, new_n419_ );
or g313 ( new_n421_, new_n418_, keyIn_0_35 );
and g314 ( new_n422_, new_n420_, new_n421_ );
or g315 ( new_n423_, new_n410_, new_n422_ );
and g316 ( new_n424_, new_n423_, keyIn_0_46 );
not g317 ( new_n425_, new_n424_ );
not g318 ( new_n426_, keyIn_0_45 );
and g319 ( new_n427_, new_n398_, new_n351_ );
and g320 ( new_n428_, new_n402_, new_n380_ );
or g321 ( new_n429_, new_n427_, new_n428_ );
and g322 ( new_n430_, new_n429_, keyIn_0_41 );
not g323 ( new_n431_, keyIn_0_41 );
or g324 ( new_n432_, new_n402_, new_n380_ );
or g325 ( new_n433_, new_n398_, new_n351_ );
and g326 ( new_n434_, new_n433_, new_n432_ );
and g327 ( new_n435_, new_n434_, new_n431_ );
or g328 ( new_n436_, new_n430_, new_n435_ );
not g329 ( new_n437_, N53 );
and g330 ( new_n438_, new_n337_, new_n437_ );
and g331 ( new_n439_, new_n348_, new_n438_ );
and g332 ( new_n440_, new_n436_, new_n439_ );
or g333 ( new_n441_, new_n440_, new_n426_ );
or g334 ( new_n442_, new_n434_, new_n431_ );
or g335 ( new_n443_, new_n429_, keyIn_0_41 );
and g336 ( new_n444_, new_n443_, new_n442_ );
not g337 ( new_n445_, new_n439_ );
or g338 ( new_n446_, new_n444_, new_n445_ );
or g339 ( new_n447_, new_n446_, keyIn_0_45 );
and g340 ( new_n448_, new_n447_, new_n441_ );
and g341 ( new_n449_, new_n448_, new_n425_ );
not g342 ( new_n450_, keyIn_0_40 );
and g343 ( new_n451_, new_n398_, new_n359_ );
and g344 ( new_n452_, new_n402_, new_n237_ );
or g345 ( new_n453_, new_n451_, new_n452_ );
and g346 ( new_n454_, new_n453_, new_n450_ );
not g347 ( new_n455_, new_n454_ );
or g348 ( new_n456_, new_n453_, new_n450_ );
not g349 ( new_n457_, N27 );
and g350 ( new_n458_, new_n457_, N17 );
and g351 ( new_n459_, new_n234_, new_n458_ );
and g352 ( new_n460_, new_n459_, keyIn_0_33 );
not g353 ( new_n461_, new_n460_ );
or g354 ( new_n462_, new_n459_, keyIn_0_33 );
and g355 ( new_n463_, new_n461_, new_n462_ );
and g356 ( new_n464_, new_n456_, new_n463_ );
and g357 ( new_n465_, new_n464_, new_n455_ );
not g358 ( new_n466_, new_n465_ );
or g359 ( new_n467_, new_n402_, new_n377_ );
or g360 ( new_n468_, new_n398_, new_n326_ );
and g361 ( new_n469_, new_n468_, new_n467_ );
and g362 ( new_n470_, new_n469_, keyIn_0_39 );
not g363 ( new_n471_, keyIn_0_39 );
and g364 ( new_n472_, new_n398_, new_n326_ );
and g365 ( new_n473_, new_n402_, new_n377_ );
or g366 ( new_n474_, new_n472_, new_n473_ );
and g367 ( new_n475_, new_n474_, new_n471_ );
not g368 ( new_n476_, keyIn_0_28 );
not g369 ( new_n477_, N14 );
and g370 ( new_n478_, new_n312_, new_n477_ );
and g371 ( new_n479_, new_n323_, new_n478_ );
not g372 ( new_n480_, new_n479_ );
and g373 ( new_n481_, new_n480_, new_n476_ );
and g374 ( new_n482_, new_n479_, keyIn_0_28 );
or g375 ( new_n483_, new_n481_, new_n482_ );
not g376 ( new_n484_, new_n483_ );
or g377 ( new_n485_, new_n475_, new_n484_ );
or g378 ( new_n486_, new_n485_, new_n470_ );
or g379 ( new_n487_, new_n402_, new_n249_ );
or g380 ( new_n488_, new_n398_, new_n248_ );
and g381 ( new_n489_, new_n488_, new_n487_ );
and g382 ( new_n490_, new_n489_, keyIn_0_43 );
not g383 ( new_n491_, keyIn_0_43 );
and g384 ( new_n492_, new_n398_, new_n248_ );
and g385 ( new_n493_, new_n402_, new_n249_ );
or g386 ( new_n494_, new_n492_, new_n493_ );
and g387 ( new_n495_, new_n494_, new_n491_ );
not g388 ( new_n496_, keyIn_0_31 );
not g389 ( new_n497_, N115 );
and g390 ( new_n498_, new_n497_, N108 );
and g391 ( new_n499_, new_n240_, new_n498_ );
not g392 ( new_n500_, new_n499_ );
and g393 ( new_n501_, new_n500_, new_n496_ );
and g394 ( new_n502_, new_n499_, keyIn_0_31 );
or g395 ( new_n503_, new_n501_, new_n502_ );
not g396 ( new_n504_, new_n503_ );
or g397 ( new_n505_, new_n495_, new_n504_ );
or g398 ( new_n506_, new_n505_, new_n490_ );
and g399 ( new_n507_, new_n486_, new_n506_ );
and g400 ( new_n508_, new_n507_, new_n466_ );
or g401 ( new_n509_, new_n423_, keyIn_0_46 );
and g402 ( new_n510_, new_n402_, new_n270_ );
not g403 ( new_n511_, new_n510_ );
and g404 ( new_n512_, new_n398_, new_n363_ );
not g405 ( new_n513_, new_n512_ );
not g406 ( new_n514_, N66 );
and g407 ( new_n515_, new_n514_, N56 );
and g408 ( new_n516_, new_n261_, new_n515_ );
and g409 ( new_n517_, new_n513_, new_n516_ );
and g410 ( new_n518_, new_n517_, new_n511_ );
not g411 ( new_n519_, new_n518_ );
or g412 ( new_n520_, new_n398_, new_n287_ );
or g413 ( new_n521_, new_n402_, new_n366_ );
and g414 ( new_n522_, new_n520_, new_n521_ );
not g415 ( new_n523_, keyIn_0_36 );
not g416 ( new_n524_, new_n282_ );
not g417 ( new_n525_, new_n283_ );
and g418 ( new_n526_, new_n524_, new_n525_ );
not g419 ( new_n527_, keyIn_0_15 );
not g420 ( new_n528_, N92 );
and g421 ( new_n529_, new_n528_, N82 );
and g422 ( new_n530_, new_n529_, new_n527_ );
not g423 ( new_n531_, new_n530_ );
or g424 ( new_n532_, new_n529_, new_n527_ );
and g425 ( new_n533_, new_n531_, new_n532_ );
or g426 ( new_n534_, new_n526_, new_n533_ );
and g427 ( new_n535_, new_n534_, new_n523_ );
not g428 ( new_n536_, new_n535_ );
or g429 ( new_n537_, new_n534_, new_n523_ );
and g430 ( new_n538_, new_n536_, new_n537_ );
or g431 ( new_n539_, new_n522_, new_n538_ );
or g432 ( new_n540_, new_n398_, new_n280_ );
or g433 ( new_n541_, new_n402_, new_n364_ );
and g434 ( new_n542_, new_n540_, new_n541_ );
not g435 ( new_n543_, keyIn_0_34 );
not g436 ( new_n544_, new_n271_ );
not g437 ( new_n545_, new_n272_ );
and g438 ( new_n546_, new_n544_, new_n545_ );
not g439 ( new_n547_, keyIn_0_11 );
not g440 ( new_n548_, N40 );
and g441 ( new_n549_, new_n278_, new_n548_ );
and g442 ( new_n550_, new_n549_, new_n547_ );
not g443 ( new_n551_, new_n550_ );
or g444 ( new_n552_, new_n549_, new_n547_ );
and g445 ( new_n553_, new_n551_, new_n552_ );
or g446 ( new_n554_, new_n546_, new_n553_ );
and g447 ( new_n555_, new_n554_, new_n543_ );
not g448 ( new_n556_, new_n555_ );
or g449 ( new_n557_, new_n554_, new_n543_ );
and g450 ( new_n558_, new_n556_, new_n557_ );
or g451 ( new_n559_, new_n542_, new_n558_ );
and g452 ( new_n560_, new_n539_, new_n559_ );
and g453 ( new_n561_, new_n560_, new_n519_ );
or g454 ( new_n562_, new_n398_, new_n255_ );
or g455 ( new_n563_, new_n402_, new_n256_ );
and g456 ( new_n564_, new_n562_, new_n563_ );
not g457 ( new_n565_, N105 );
and g458 ( new_n566_, new_n565_, N95 );
and g459 ( new_n567_, new_n566_, keyIn_0_16 );
not g460 ( new_n568_, new_n567_ );
or g461 ( new_n569_, new_n566_, keyIn_0_16 );
and g462 ( new_n570_, new_n568_, new_n569_ );
and g463 ( new_n571_, new_n252_, new_n570_ );
not g464 ( new_n572_, new_n571_ );
or g465 ( new_n573_, new_n564_, new_n572_ );
or g466 ( new_n574_, new_n573_, keyIn_0_47 );
not g467 ( new_n575_, keyIn_0_47 );
and g468 ( new_n576_, new_n402_, new_n256_ );
and g469 ( new_n577_, new_n398_, new_n255_ );
or g470 ( new_n578_, new_n577_, new_n576_ );
and g471 ( new_n579_, new_n578_, new_n571_ );
or g472 ( new_n580_, new_n579_, new_n575_ );
and g473 ( new_n581_, new_n574_, new_n580_ );
and g474 ( new_n582_, new_n581_, new_n561_ );
and g475 ( new_n583_, new_n509_, new_n582_ );
and g476 ( new_n584_, new_n583_, new_n508_ );
and g477 ( new_n585_, new_n449_, new_n584_ );
not g478 ( new_n586_, new_n585_ );
and g479 ( new_n587_, new_n586_, new_n393_ );
and g480 ( new_n588_, new_n585_, keyIn_0_48 );
or g481 ( N370, new_n587_, new_n588_ );
not g482 ( new_n590_, keyIn_0_58 );
not g483 ( new_n591_, keyIn_0_49 );
or g484 ( new_n592_, new_n585_, keyIn_0_48 );
not g485 ( new_n593_, new_n588_ );
and g486 ( new_n594_, new_n593_, new_n592_ );
and g487 ( new_n595_, new_n594_, new_n591_ );
not g488 ( new_n596_, new_n595_ );
or g489 ( new_n597_, new_n594_, new_n591_ );
and g490 ( new_n598_, new_n597_, N105 );
and g491 ( new_n599_, new_n598_, new_n596_ );
not g492 ( new_n600_, new_n599_ );
and g493 ( new_n601_, new_n600_, keyIn_0_52 );
not g494 ( new_n602_, keyIn_0_52 );
and g495 ( new_n603_, new_n599_, new_n602_ );
and g496 ( new_n604_, new_n390_, N99 );
and g497 ( new_n605_, new_n206_, keyIn_0_19 );
not g498 ( new_n606_, new_n605_ );
or g499 ( new_n607_, new_n206_, keyIn_0_19 );
and g500 ( new_n608_, new_n606_, new_n607_ );
not g501 ( new_n609_, new_n608_ );
and g502 ( new_n610_, new_n609_, N89 );
or g503 ( new_n611_, new_n610_, new_n109_ );
or g504 ( new_n612_, new_n604_, new_n611_ );
or g505 ( new_n613_, new_n603_, new_n612_ );
or g506 ( new_n614_, new_n613_, new_n601_ );
and g507 ( new_n615_, new_n614_, keyIn_0_55 );
not g508 ( new_n616_, new_n615_ );
or g509 ( new_n617_, new_n614_, keyIn_0_55 );
and g510 ( new_n618_, new_n616_, new_n617_ );
not g511 ( new_n619_, keyIn_0_50 );
and g512 ( new_n620_, new_n597_, N66 );
and g513 ( new_n621_, new_n620_, new_n596_ );
and g514 ( new_n622_, new_n621_, new_n619_ );
and g515 ( new_n623_, N370, keyIn_0_49 );
or g516 ( new_n624_, new_n623_, new_n514_ );
or g517 ( new_n625_, new_n624_, new_n595_ );
and g518 ( new_n626_, new_n625_, keyIn_0_50 );
and g519 ( new_n627_, new_n390_, N60 );
not g520 ( new_n628_, new_n627_ );
not g521 ( new_n629_, keyIn_0_24 );
and g522 ( new_n630_, new_n609_, N50 );
and g523 ( new_n631_, new_n630_, new_n629_ );
not g524 ( new_n632_, new_n631_ );
or g525 ( new_n633_, new_n630_, new_n629_ );
and g526 ( new_n634_, new_n633_, N56 );
and g527 ( new_n635_, new_n634_, new_n632_ );
and g528 ( new_n636_, new_n628_, new_n635_ );
not g529 ( new_n637_, new_n636_ );
or g530 ( new_n638_, new_n626_, new_n637_ );
or g531 ( new_n639_, new_n638_, new_n622_ );
or g532 ( new_n640_, new_n623_, new_n437_ );
or g533 ( new_n641_, new_n640_, new_n595_ );
and g534 ( new_n642_, new_n390_, N47 );
and g535 ( new_n643_, new_n609_, N37 );
not g536 ( new_n644_, new_n643_ );
and g537 ( new_n645_, new_n644_, keyIn_0_23 );
not g538 ( new_n646_, new_n645_ );
or g539 ( new_n647_, new_n644_, keyIn_0_23 );
and g540 ( new_n648_, new_n646_, new_n647_ );
or g541 ( new_n649_, new_n648_, new_n199_ );
or g542 ( new_n650_, new_n642_, new_n649_ );
not g543 ( new_n651_, new_n650_ );
and g544 ( new_n652_, new_n641_, new_n651_ );
not g545 ( new_n653_, new_n652_ );
and g546 ( new_n654_, new_n639_, new_n653_ );
and g547 ( new_n655_, new_n597_, N115 );
and g548 ( new_n656_, new_n655_, new_n596_ );
not g549 ( new_n657_, new_n656_ );
not g550 ( new_n658_, keyIn_0_44 );
and g551 ( new_n659_, new_n390_, N112 );
not g552 ( new_n660_, new_n659_ );
and g553 ( new_n661_, new_n660_, new_n658_ );
and g554 ( new_n662_, new_n659_, keyIn_0_44 );
or g555 ( new_n663_, new_n661_, new_n662_ );
and g556 ( new_n664_, new_n609_, N102 );
or g557 ( new_n665_, new_n664_, new_n133_ );
not g558 ( new_n666_, new_n665_ );
and g559 ( new_n667_, new_n663_, new_n666_ );
and g560 ( new_n668_, new_n657_, new_n667_ );
not g561 ( new_n669_, new_n668_ );
and g562 ( new_n670_, new_n669_, keyIn_0_56 );
not g563 ( new_n671_, keyIn_0_56 );
and g564 ( new_n672_, new_n668_, new_n671_ );
or g565 ( new_n673_, new_n670_, new_n672_ );
and g566 ( new_n674_, new_n597_, N27 );
and g567 ( new_n675_, new_n674_, new_n596_ );
and g568 ( new_n676_, new_n390_, N21 );
not g569 ( new_n677_, new_n676_ );
not g570 ( new_n678_, keyIn_0_22 );
and g571 ( new_n679_, new_n609_, N11 );
and g572 ( new_n680_, new_n679_, new_n678_ );
not g573 ( new_n681_, new_n680_ );
or g574 ( new_n682_, new_n679_, new_n678_ );
and g575 ( new_n683_, new_n682_, N17 );
and g576 ( new_n684_, new_n683_, new_n681_ );
and g577 ( new_n685_, new_n677_, new_n684_ );
not g578 ( new_n686_, new_n685_ );
or g579 ( new_n687_, new_n675_, new_n686_ );
and g580 ( new_n688_, new_n597_, N40 );
and g581 ( new_n689_, new_n688_, new_n596_ );
and g582 ( new_n690_, new_n390_, N34 );
and g583 ( new_n691_, new_n609_, N24 );
or g584 ( new_n692_, new_n691_, new_n126_ );
or g585 ( new_n693_, new_n690_, new_n692_ );
or g586 ( new_n694_, new_n689_, new_n693_ );
and g587 ( new_n695_, new_n687_, new_n694_ );
and g588 ( new_n696_, new_n673_, new_n695_ );
not g589 ( new_n697_, keyIn_0_51 );
and g590 ( new_n698_, new_n597_, N79 );
and g591 ( new_n699_, new_n698_, new_n596_ );
and g592 ( new_n700_, new_n699_, new_n697_ );
not g593 ( new_n701_, new_n700_ );
or g594 ( new_n702_, new_n699_, new_n697_ );
and g595 ( new_n703_, new_n701_, new_n702_ );
and g596 ( new_n704_, new_n390_, N73 );
not g597 ( new_n705_, new_n704_ );
not g598 ( new_n706_, keyIn_0_25 );
and g599 ( new_n707_, new_n609_, N63 );
and g600 ( new_n708_, new_n707_, new_n706_ );
not g601 ( new_n709_, new_n708_ );
or g602 ( new_n710_, new_n707_, new_n706_ );
and g603 ( new_n711_, new_n710_, N69 );
and g604 ( new_n712_, new_n711_, new_n709_ );
and g605 ( new_n713_, new_n705_, new_n712_ );
not g606 ( new_n714_, new_n713_ );
or g607 ( new_n715_, new_n703_, new_n714_ );
not g608 ( new_n716_, keyIn_0_54 );
or g609 ( new_n717_, new_n623_, new_n528_ );
or g610 ( new_n718_, new_n717_, new_n595_ );
and g611 ( new_n719_, new_n390_, N86 );
not g612 ( new_n720_, new_n719_ );
not g613 ( new_n721_, keyIn_0_26 );
and g614 ( new_n722_, new_n609_, N76 );
and g615 ( new_n723_, new_n722_, new_n721_ );
not g616 ( new_n724_, new_n723_ );
or g617 ( new_n725_, new_n722_, new_n721_ );
and g618 ( new_n726_, new_n725_, N82 );
and g619 ( new_n727_, new_n726_, new_n724_ );
and g620 ( new_n728_, new_n720_, new_n727_ );
and g621 ( new_n729_, new_n718_, new_n728_ );
and g622 ( new_n730_, new_n729_, new_n716_ );
and g623 ( new_n731_, new_n597_, N92 );
and g624 ( new_n732_, new_n731_, new_n596_ );
not g625 ( new_n733_, new_n728_ );
or g626 ( new_n734_, new_n732_, new_n733_ );
and g627 ( new_n735_, new_n734_, keyIn_0_54 );
or g628 ( new_n736_, new_n730_, new_n735_ );
and g629 ( new_n737_, new_n715_, new_n736_ );
and g630 ( new_n738_, new_n696_, new_n737_ );
and g631 ( new_n739_, new_n738_, new_n654_ );
and g632 ( new_n740_, new_n739_, new_n618_ );
or g633 ( new_n741_, new_n740_, new_n590_ );
and g634 ( new_n742_, new_n740_, new_n590_ );
not g635 ( new_n743_, new_n742_ );
not g636 ( new_n744_, keyIn_0_57 );
and g637 ( new_n745_, new_n597_, N14 );
and g638 ( new_n746_, new_n745_, new_n596_ );
and g639 ( new_n747_, new_n390_, N8 );
and g640 ( new_n748_, new_n609_, N1 );
or g641 ( new_n749_, new_n748_, new_n189_ );
or g642 ( new_n750_, new_n747_, new_n749_ );
or g643 ( new_n751_, new_n746_, new_n750_ );
and g644 ( new_n752_, new_n751_, keyIn_0_53 );
not g645 ( new_n753_, new_n752_ );
or g646 ( new_n754_, new_n751_, keyIn_0_53 );
and g647 ( new_n755_, new_n753_, new_n754_ );
not g648 ( new_n756_, new_n755_ );
or g649 ( new_n757_, new_n756_, new_n744_ );
or g650 ( new_n758_, new_n755_, keyIn_0_57 );
and g651 ( new_n759_, new_n757_, new_n758_ );
and g652 ( new_n760_, new_n743_, new_n759_ );
and g653 ( N421, new_n760_, new_n741_ );
and g654 ( new_n762_, new_n652_, new_n694_ );
not g655 ( new_n763_, new_n762_ );
and g656 ( new_n764_, new_n763_, keyIn_0_60 );
not g657 ( new_n765_, new_n764_ );
or g658 ( new_n766_, new_n763_, keyIn_0_60 );
and g659 ( new_n767_, new_n765_, new_n766_ );
not g660 ( new_n768_, new_n767_ );
and g661 ( new_n769_, new_n639_, new_n695_ );
and g662 ( new_n770_, new_n768_, new_n769_ );
not g663 ( new_n771_, new_n770_ );
and g664 ( new_n772_, new_n771_, keyIn_0_62 );
not g665 ( new_n773_, keyIn_0_62 );
and g666 ( new_n774_, new_n770_, new_n773_ );
or g667 ( N430, new_n772_, new_n774_ );
not g668 ( new_n776_, keyIn_0_63 );
not g669 ( new_n777_, keyIn_0_59 );
or g670 ( new_n778_, new_n734_, keyIn_0_54 );
or g671 ( new_n779_, new_n729_, new_n716_ );
and g672 ( new_n780_, new_n779_, new_n778_ );
and g673 ( new_n781_, new_n780_, new_n777_ );
not g674 ( new_n782_, new_n781_ );
or g675 ( new_n783_, new_n780_, new_n777_ );
and g676 ( new_n784_, new_n783_, new_n654_ );
and g677 ( new_n785_, new_n784_, new_n782_ );
and g678 ( new_n786_, new_n785_, keyIn_0_61 );
not g679 ( new_n787_, keyIn_0_61 );
not g680 ( new_n788_, new_n622_ );
or g681 ( new_n789_, new_n621_, new_n619_ );
and g682 ( new_n790_, new_n789_, new_n636_ );
and g683 ( new_n791_, new_n790_, new_n788_ );
or g684 ( new_n792_, new_n791_, new_n652_ );
and g685 ( new_n793_, new_n736_, keyIn_0_59 );
or g686 ( new_n794_, new_n793_, new_n792_ );
or g687 ( new_n795_, new_n794_, new_n781_ );
and g688 ( new_n796_, new_n795_, new_n787_ );
not g689 ( new_n797_, new_n694_ );
or g690 ( new_n798_, new_n715_, new_n797_ );
or g691 ( new_n799_, new_n798_, new_n792_ );
and g692 ( new_n800_, new_n799_, new_n695_ );
not g693 ( new_n801_, new_n800_ );
or g694 ( new_n802_, new_n796_, new_n801_ );
or g695 ( new_n803_, new_n802_, new_n786_ );
and g696 ( new_n804_, new_n803_, new_n776_ );
not g697 ( new_n805_, new_n786_ );
or g698 ( new_n806_, new_n785_, keyIn_0_61 );
and g699 ( new_n807_, new_n806_, new_n800_ );
and g700 ( new_n808_, new_n807_, new_n805_ );
and g701 ( new_n809_, new_n808_, keyIn_0_63 );
or g702 ( N431, new_n804_, new_n809_ );
not g703 ( new_n811_, new_n618_ );
and g704 ( new_n812_, new_n653_, new_n694_ );
and g705 ( new_n813_, new_n736_, new_n812_ );
and g706 ( new_n814_, new_n811_, new_n813_ );
not g707 ( new_n815_, new_n799_ );
not g708 ( new_n816_, new_n687_ );
or g709 ( new_n817_, new_n767_, new_n816_ );
or g710 ( new_n818_, new_n817_, new_n815_ );
or g711 ( N432, new_n818_, new_n814_ );
endmodule