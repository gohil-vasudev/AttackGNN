module locked_c3540 (  G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698, G2897, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,  G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698, G2897, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1409_, new_n1410_, new_n1411_, new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1453_, new_n1454_, new_n1455_, new_n1456_;
  INV_X1 g0000 ( .A(G58), .ZN(new_n137_) );
  INV_X1 g0001 ( .A(G68), .ZN(new_n138_) );
  AND2_X1 g0002 ( .A1(new_n137_), .A2(new_n138_), .ZN(new_n139_) );
  INV_X1 g0003 ( .A(G50), .ZN(new_n140_) );
  INV_X1 g0004 ( .A(G77), .ZN(new_n141_) );
  AND2_X1 g0005 ( .A1(new_n140_), .A2(new_n141_), .ZN(new_n142_) );
  AND2_X1 g0006 ( .A1(new_n139_), .A2(new_n142_), .ZN(G353) );
  INV_X1 g0007 ( .A(G97), .ZN(new_n144_) );
  INV_X1 g0008 ( .A(G107), .ZN(new_n145_) );
  AND2_X1 g0009 ( .A1(new_n144_), .A2(new_n145_), .ZN(new_n146_) );
  INV_X1 g0010 ( .A(new_n146_), .ZN(new_n147_) );
  AND2_X1 g0011 ( .A1(new_n147_), .A2(G87), .ZN(new_n148_) );
  INV_X1 g0012 ( .A(new_n148_), .ZN(G355) );
  AND2_X1 g0013 ( .A1(G1), .A2(G20), .ZN(new_n150_) );
  INV_X1 g0014 ( .A(KEYINPUT49), .ZN(new_n151_) );
  AND2_X1 g0015 ( .A1(G50), .A2(G226), .ZN(new_n152_) );
  AND2_X1 g0016 ( .A1(G58), .A2(G232), .ZN(new_n153_) );
  AND2_X1 g0017 ( .A1(G77), .A2(G244), .ZN(new_n154_) );
  AND2_X1 g0018 ( .A1(G68), .A2(G238), .ZN(new_n155_) );
  OR4_X1 g0019 ( .A1(new_n152_), .A2(new_n153_), .A3(new_n154_), .A4(new_n155_), .ZN(new_n156_) );
  OR2_X1 g0020 ( .A1(new_n156_), .A2(new_n151_), .ZN(new_n157_) );
  INV_X1 g0021 ( .A(new_n156_), .ZN(new_n158_) );
  OR2_X1 g0022 ( .A1(new_n158_), .A2(KEYINPUT49), .ZN(new_n159_) );
  INV_X1 g0023 ( .A(KEYINPUT50), .ZN(new_n160_) );
  AND2_X1 g0024 ( .A1(G107), .A2(G264), .ZN(new_n161_) );
  AND2_X1 g0025 ( .A1(new_n161_), .A2(new_n160_), .ZN(new_n162_) );
  INV_X1 g0026 ( .A(new_n161_), .ZN(new_n163_) );
  AND2_X1 g0027 ( .A1(new_n163_), .A2(KEYINPUT50), .ZN(new_n164_) );
  OR2_X1 g0028 ( .A1(new_n164_), .A2(new_n162_), .ZN(new_n165_) );
  AND2_X1 g0029 ( .A1(G97), .A2(G257), .ZN(new_n166_) );
  INV_X1 g0030 ( .A(new_n166_), .ZN(new_n167_) );
  AND2_X1 g0031 ( .A1(G87), .A2(G250), .ZN(new_n168_) );
  INV_X1 g0032 ( .A(new_n168_), .ZN(new_n169_) );
  AND2_X1 g0033 ( .A1(G116), .A2(G270), .ZN(new_n170_) );
  INV_X1 g0034 ( .A(new_n170_), .ZN(new_n171_) );
  AND3_X1 g0035 ( .A1(new_n167_), .A2(new_n169_), .A3(new_n171_), .ZN(new_n172_) );
  AND4_X1 g0036 ( .A1(new_n159_), .A2(new_n157_), .A3(new_n165_), .A4(new_n172_), .ZN(new_n173_) );
  OR2_X1 g0037 ( .A1(new_n173_), .A2(new_n150_), .ZN(new_n174_) );
  INV_X1 g0038 ( .A(G20), .ZN(new_n175_) );
  AND3_X1 g0039 ( .A1(G1), .A2(G13), .A3(KEYINPUT2), .ZN(new_n176_) );
  INV_X1 g0040 ( .A(new_n176_), .ZN(new_n177_) );
  AND2_X1 g0041 ( .A1(G1), .A2(G13), .ZN(new_n178_) );
  OR2_X1 g0042 ( .A1(new_n178_), .A2(KEYINPUT2), .ZN(new_n179_) );
  AND2_X1 g0043 ( .A1(new_n179_), .A2(new_n177_), .ZN(new_n180_) );
  OR2_X1 g0044 ( .A1(new_n180_), .A2(new_n175_), .ZN(new_n181_) );
  OR3_X1 g0045 ( .A1(new_n181_), .A2(new_n140_), .A3(new_n139_), .ZN(new_n182_) );
  INV_X1 g0046 ( .A(G13), .ZN(new_n183_) );
  AND2_X1 g0047 ( .A1(new_n150_), .A2(new_n183_), .ZN(new_n184_) );
  OR2_X1 g0048 ( .A1(G257), .A2(G264), .ZN(new_n185_) );
  AND3_X1 g0049 ( .A1(new_n184_), .A2(G250), .A3(new_n185_), .ZN(new_n186_) );
  INV_X1 g0050 ( .A(new_n186_), .ZN(new_n187_) );
  AND3_X1 g0051 ( .A1(new_n174_), .A2(new_n182_), .A3(new_n187_), .ZN(G361) );
  INV_X1 g0052 ( .A(G238), .ZN(new_n189_) );
  INV_X1 g0053 ( .A(G232), .ZN(new_n190_) );
  INV_X1 g0054 ( .A(G244), .ZN(new_n191_) );
  AND2_X1 g0055 ( .A1(new_n190_), .A2(new_n191_), .ZN(new_n192_) );
  AND2_X1 g0056 ( .A1(G232), .A2(G244), .ZN(new_n193_) );
  OR2_X1 g0057 ( .A1(new_n192_), .A2(new_n193_), .ZN(new_n194_) );
  INV_X1 g0058 ( .A(new_n194_), .ZN(new_n195_) );
  AND2_X1 g0059 ( .A1(new_n195_), .A2(G226), .ZN(new_n196_) );
  INV_X1 g0060 ( .A(G226), .ZN(new_n197_) );
  AND2_X1 g0061 ( .A1(new_n194_), .A2(new_n197_), .ZN(new_n198_) );
  OR2_X1 g0062 ( .A1(new_n196_), .A2(new_n198_), .ZN(new_n199_) );
  INV_X1 g0063 ( .A(new_n199_), .ZN(new_n200_) );
  AND2_X1 g0064 ( .A1(new_n200_), .A2(new_n189_), .ZN(new_n201_) );
  AND2_X1 g0065 ( .A1(new_n199_), .A2(G238), .ZN(new_n202_) );
  OR2_X1 g0066 ( .A1(new_n201_), .A2(new_n202_), .ZN(new_n203_) );
  OR2_X1 g0067 ( .A1(G264), .A2(G270), .ZN(new_n204_) );
  AND2_X1 g0068 ( .A1(G264), .A2(G270), .ZN(new_n205_) );
  INV_X1 g0069 ( .A(new_n205_), .ZN(new_n206_) );
  AND2_X1 g0070 ( .A1(new_n206_), .A2(new_n204_), .ZN(new_n207_) );
  INV_X1 g0071 ( .A(G250), .ZN(new_n208_) );
  INV_X1 g0072 ( .A(G257), .ZN(new_n209_) );
  AND2_X1 g0073 ( .A1(new_n208_), .A2(new_n209_), .ZN(new_n210_) );
  AND2_X1 g0074 ( .A1(G250), .A2(G257), .ZN(new_n211_) );
  OR2_X1 g0075 ( .A1(new_n210_), .A2(new_n211_), .ZN(new_n212_) );
  INV_X1 g0076 ( .A(new_n212_), .ZN(new_n213_) );
  AND2_X1 g0077 ( .A1(new_n213_), .A2(new_n207_), .ZN(new_n214_) );
  INV_X1 g0078 ( .A(new_n214_), .ZN(new_n215_) );
  OR2_X1 g0079 ( .A1(new_n213_), .A2(new_n207_), .ZN(new_n216_) );
  AND2_X1 g0080 ( .A1(new_n215_), .A2(new_n216_), .ZN(new_n217_) );
  AND2_X1 g0081 ( .A1(new_n203_), .A2(new_n217_), .ZN(new_n218_) );
  INV_X1 g0082 ( .A(new_n203_), .ZN(new_n219_) );
  INV_X1 g0083 ( .A(new_n217_), .ZN(new_n220_) );
  AND2_X1 g0084 ( .A1(new_n219_), .A2(new_n220_), .ZN(new_n221_) );
  OR2_X1 g0085 ( .A1(new_n221_), .A2(new_n218_), .ZN(G358) );
  INV_X1 g0086 ( .A(KEYINPUT51), .ZN(new_n223_) );
  AND2_X1 g0087 ( .A1(G97), .A2(G107), .ZN(new_n224_) );
  OR2_X1 g0088 ( .A1(new_n146_), .A2(new_n224_), .ZN(new_n225_) );
  AND2_X1 g0089 ( .A1(new_n225_), .A2(new_n223_), .ZN(new_n226_) );
  INV_X1 g0090 ( .A(new_n225_), .ZN(new_n227_) );
  AND2_X1 g0091 ( .A1(new_n227_), .A2(KEYINPUT51), .ZN(new_n228_) );
  OR2_X1 g0092 ( .A1(new_n228_), .A2(new_n226_), .ZN(new_n229_) );
  INV_X1 g0093 ( .A(new_n229_), .ZN(new_n230_) );
  INV_X1 g0094 ( .A(G87), .ZN(new_n231_) );
  INV_X1 g0095 ( .A(G116), .ZN(new_n232_) );
  AND2_X1 g0096 ( .A1(new_n231_), .A2(new_n232_), .ZN(new_n233_) );
  AND2_X1 g0097 ( .A1(G87), .A2(G116), .ZN(new_n234_) );
  OR2_X1 g0098 ( .A1(new_n233_), .A2(new_n234_), .ZN(new_n235_) );
  INV_X1 g0099 ( .A(new_n235_), .ZN(new_n236_) );
  AND2_X1 g0100 ( .A1(new_n230_), .A2(new_n236_), .ZN(new_n237_) );
  AND2_X1 g0101 ( .A1(new_n229_), .A2(new_n235_), .ZN(new_n238_) );
  OR2_X1 g0102 ( .A1(new_n237_), .A2(new_n238_), .ZN(new_n239_) );
  INV_X1 g0103 ( .A(new_n239_), .ZN(new_n240_) );
  AND2_X1 g0104 ( .A1(G50), .A2(G77), .ZN(new_n241_) );
  OR2_X1 g0105 ( .A1(new_n142_), .A2(new_n241_), .ZN(new_n242_) );
  INV_X1 g0106 ( .A(new_n242_), .ZN(new_n243_) );
  AND2_X1 g0107 ( .A1(G58), .A2(G68), .ZN(new_n244_) );
  OR2_X1 g0108 ( .A1(new_n139_), .A2(new_n244_), .ZN(new_n245_) );
  INV_X1 g0109 ( .A(new_n245_), .ZN(new_n246_) );
  AND2_X1 g0110 ( .A1(new_n243_), .A2(new_n246_), .ZN(new_n247_) );
  AND2_X1 g0111 ( .A1(new_n242_), .A2(new_n245_), .ZN(new_n248_) );
  OR2_X1 g0112 ( .A1(new_n247_), .A2(new_n248_), .ZN(new_n249_) );
  INV_X1 g0113 ( .A(new_n249_), .ZN(new_n250_) );
  AND2_X1 g0114 ( .A1(new_n240_), .A2(new_n250_), .ZN(new_n251_) );
  AND2_X1 g0115 ( .A1(new_n239_), .A2(new_n249_), .ZN(new_n252_) );
  OR2_X1 g0116 ( .A1(new_n251_), .A2(new_n252_), .ZN(G351) );
  INV_X1 g0117 ( .A(KEYINPUT30), .ZN(new_n254_) );
  AND3_X1 g0118 ( .A1(G1), .A2(G20), .A3(G33), .ZN(new_n255_) );
  OR2_X1 g0119 ( .A1(new_n255_), .A2(KEYINPUT3), .ZN(new_n256_) );
  AND4_X1 g0120 ( .A1(G1), .A2(G20), .A3(G33), .A4(KEYINPUT3), .ZN(new_n257_) );
  INV_X1 g0121 ( .A(new_n257_), .ZN(new_n258_) );
  AND2_X1 g0122 ( .A1(new_n256_), .A2(new_n258_), .ZN(new_n259_) );
  INV_X1 g0123 ( .A(new_n259_), .ZN(new_n260_) );
  AND2_X1 g0124 ( .A1(new_n260_), .A2(new_n180_), .ZN(new_n261_) );
  OR3_X1 g0125 ( .A1(new_n261_), .A2(new_n175_), .A3(KEYINPUT4), .ZN(new_n262_) );
  INV_X1 g0126 ( .A(KEYINPUT4), .ZN(new_n263_) );
  INV_X1 g0127 ( .A(new_n180_), .ZN(new_n264_) );
  OR2_X1 g0128 ( .A1(new_n264_), .A2(new_n259_), .ZN(new_n265_) );
  AND2_X1 g0129 ( .A1(new_n265_), .A2(G20), .ZN(new_n266_) );
  OR2_X1 g0130 ( .A1(new_n266_), .A2(new_n263_), .ZN(new_n267_) );
  AND2_X1 g0131 ( .A1(new_n267_), .A2(new_n262_), .ZN(new_n268_) );
  AND2_X1 g0132 ( .A1(new_n268_), .A2(new_n245_), .ZN(new_n269_) );
  INV_X1 g0133 ( .A(G1), .ZN(new_n270_) );
  AND2_X1 g0134 ( .A1(new_n270_), .A2(G20), .ZN(new_n271_) );
  OR2_X1 g0135 ( .A1(new_n265_), .A2(new_n271_), .ZN(new_n272_) );
  INV_X1 g0136 ( .A(new_n272_), .ZN(new_n273_) );
  AND2_X1 g0137 ( .A1(new_n273_), .A2(G58), .ZN(new_n274_) );
  INV_X1 g0138 ( .A(G33), .ZN(new_n275_) );
  AND3_X1 g0139 ( .A1(new_n264_), .A2(new_n175_), .A3(new_n275_), .ZN(new_n276_) );
  AND2_X1 g0140 ( .A1(new_n276_), .A2(G159), .ZN(new_n277_) );
  OR2_X1 g0141 ( .A1(new_n275_), .A2(G20), .ZN(new_n278_) );
  OR2_X1 g0142 ( .A1(new_n180_), .A2(new_n278_), .ZN(new_n279_) );
  INV_X1 g0143 ( .A(new_n279_), .ZN(new_n280_) );
  AND2_X1 g0144 ( .A1(new_n280_), .A2(G68), .ZN(new_n281_) );
  AND2_X1 g0145 ( .A1(new_n271_), .A2(G13), .ZN(new_n282_) );
  AND2_X1 g0146 ( .A1(new_n282_), .A2(new_n137_), .ZN(new_n283_) );
  OR4_X1 g0147 ( .A1(new_n274_), .A2(new_n277_), .A3(new_n281_), .A4(new_n283_), .ZN(new_n284_) );
  OR2_X1 g0148 ( .A1(new_n284_), .A2(new_n269_), .ZN(new_n285_) );
  AND2_X1 g0149 ( .A1(new_n285_), .A2(new_n254_), .ZN(new_n286_) );
  INV_X1 g0150 ( .A(new_n286_), .ZN(new_n287_) );
  OR2_X1 g0151 ( .A1(new_n285_), .A2(new_n254_), .ZN(new_n288_) );
  AND2_X1 g0152 ( .A1(new_n287_), .A2(new_n288_), .ZN(new_n289_) );
  INV_X1 g0153 ( .A(new_n289_), .ZN(new_n290_) );
  INV_X1 g0154 ( .A(KEYINPUT33), .ZN(new_n291_) );
  INV_X1 g0155 ( .A(G1698), .ZN(new_n292_) );
  OR3_X1 g0156 ( .A1(new_n180_), .A2(G33), .A3(new_n292_), .ZN(new_n293_) );
  INV_X1 g0157 ( .A(new_n293_), .ZN(new_n294_) );
  AND2_X1 g0158 ( .A1(new_n294_), .A2(G226), .ZN(new_n295_) );
  OR2_X1 g0159 ( .A1(new_n295_), .A2(KEYINPUT32), .ZN(new_n296_) );
  INV_X1 g0160 ( .A(new_n296_), .ZN(new_n297_) );
  OR3_X1 g0161 ( .A1(new_n180_), .A2(G33), .A3(G1698), .ZN(new_n298_) );
  INV_X1 g0162 ( .A(new_n298_), .ZN(new_n299_) );
  AND2_X1 g0163 ( .A1(new_n299_), .A2(G223), .ZN(new_n300_) );
  AND2_X1 g0164 ( .A1(new_n295_), .A2(KEYINPUT32), .ZN(new_n301_) );
  OR3_X1 g0165 ( .A1(new_n297_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_) );
  AND2_X1 g0166 ( .A1(new_n302_), .A2(new_n291_), .ZN(new_n303_) );
  INV_X1 g0167 ( .A(new_n303_), .ZN(new_n304_) );
  OR2_X1 g0168 ( .A1(new_n302_), .A2(new_n291_), .ZN(new_n305_) );
  OR3_X1 g0169 ( .A1(new_n180_), .A2(new_n275_), .A3(G41), .ZN(new_n306_) );
  INV_X1 g0170 ( .A(new_n306_), .ZN(new_n307_) );
  AND2_X1 g0171 ( .A1(new_n307_), .A2(G87), .ZN(new_n308_) );
  OR2_X1 g0172 ( .A1(new_n308_), .A2(KEYINPUT31), .ZN(new_n309_) );
  AND2_X1 g0173 ( .A1(new_n308_), .A2(KEYINPUT31), .ZN(new_n310_) );
  INV_X1 g0174 ( .A(new_n310_), .ZN(new_n311_) );
  AND2_X1 g0175 ( .A1(new_n311_), .A2(new_n309_), .ZN(new_n312_) );
  INV_X1 g0176 ( .A(new_n312_), .ZN(new_n313_) );
  INV_X1 g0177 ( .A(G41), .ZN(new_n314_) );
  INV_X1 g0178 ( .A(G45), .ZN(new_n315_) );
  AND2_X1 g0179 ( .A1(new_n314_), .A2(new_n315_), .ZN(new_n316_) );
  INV_X1 g0180 ( .A(new_n316_), .ZN(new_n317_) );
  AND3_X1 g0181 ( .A1(new_n317_), .A2(new_n270_), .A3(G274), .ZN(new_n318_) );
  INV_X1 g0182 ( .A(new_n318_), .ZN(new_n319_) );
  OR2_X1 g0183 ( .A1(new_n316_), .A2(G1), .ZN(new_n320_) );
  AND2_X1 g0184 ( .A1(G33), .A2(G41), .ZN(new_n321_) );
  OR2_X1 g0185 ( .A1(new_n180_), .A2(new_n321_), .ZN(new_n322_) );
  AND2_X1 g0186 ( .A1(new_n322_), .A2(new_n320_), .ZN(new_n323_) );
  AND2_X1 g0187 ( .A1(new_n323_), .A2(G232), .ZN(new_n324_) );
  INV_X1 g0188 ( .A(new_n324_), .ZN(new_n325_) );
  AND3_X1 g0189 ( .A1(new_n313_), .A2(new_n319_), .A3(new_n325_), .ZN(new_n326_) );
  AND3_X1 g0190 ( .A1(new_n304_), .A2(new_n305_), .A3(new_n326_), .ZN(new_n327_) );
  AND2_X1 g0191 ( .A1(new_n327_), .A2(G179), .ZN(new_n328_) );
  OR2_X1 g0192 ( .A1(new_n328_), .A2(KEYINPUT34), .ZN(new_n329_) );
  INV_X1 g0193 ( .A(G169), .ZN(new_n330_) );
  OR2_X1 g0194 ( .A1(new_n327_), .A2(new_n330_), .ZN(new_n331_) );
  INV_X1 g0195 ( .A(KEYINPUT34), .ZN(new_n332_) );
  INV_X1 g0196 ( .A(new_n328_), .ZN(new_n333_) );
  OR2_X1 g0197 ( .A1(new_n333_), .A2(new_n332_), .ZN(new_n334_) );
  AND3_X1 g0198 ( .A1(new_n334_), .A2(new_n329_), .A3(new_n331_), .ZN(new_n335_) );
  OR2_X1 g0199 ( .A1(new_n335_), .A2(new_n290_), .ZN(new_n336_) );
  INV_X1 g0200 ( .A(G200), .ZN(new_n337_) );
  AND2_X1 g0201 ( .A1(new_n294_), .A2(G238), .ZN(new_n338_) );
  OR2_X1 g0202 ( .A1(new_n338_), .A2(KEYINPUT6), .ZN(new_n339_) );
  INV_X1 g0203 ( .A(KEYINPUT6), .ZN(new_n340_) );
  OR3_X1 g0204 ( .A1(new_n293_), .A2(new_n189_), .A3(new_n340_), .ZN(new_n341_) );
  OR2_X1 g0205 ( .A1(new_n298_), .A2(new_n190_), .ZN(new_n342_) );
  OR2_X1 g0206 ( .A1(new_n306_), .A2(new_n145_), .ZN(new_n343_) );
  AND3_X1 g0207 ( .A1(new_n342_), .A2(new_n343_), .A3(new_n319_), .ZN(new_n344_) );
  AND3_X1 g0208 ( .A1(new_n339_), .A2(new_n344_), .A3(new_n341_), .ZN(new_n345_) );
  OR2_X1 g0209 ( .A1(new_n345_), .A2(KEYINPUT7), .ZN(new_n346_) );
  AND2_X1 g0210 ( .A1(new_n345_), .A2(KEYINPUT7), .ZN(new_n347_) );
  INV_X1 g0211 ( .A(new_n347_), .ZN(new_n348_) );
  AND2_X1 g0212 ( .A1(new_n323_), .A2(G244), .ZN(new_n349_) );
  INV_X1 g0213 ( .A(new_n349_), .ZN(new_n350_) );
  AND3_X1 g0214 ( .A1(new_n348_), .A2(new_n346_), .A3(new_n350_), .ZN(new_n351_) );
  OR2_X1 g0215 ( .A1(new_n351_), .A2(new_n337_), .ZN(new_n352_) );
  AND2_X1 g0216 ( .A1(new_n351_), .A2(G190), .ZN(new_n353_) );
  INV_X1 g0217 ( .A(new_n353_), .ZN(new_n354_) );
  OR2_X1 g0218 ( .A1(new_n268_), .A2(new_n273_), .ZN(new_n355_) );
  AND2_X1 g0219 ( .A1(new_n355_), .A2(G77), .ZN(new_n356_) );
  AND2_X1 g0220 ( .A1(new_n276_), .A2(G58), .ZN(new_n357_) );
  AND2_X1 g0221 ( .A1(new_n280_), .A2(G87), .ZN(new_n358_) );
  AND2_X1 g0222 ( .A1(new_n282_), .A2(new_n141_), .ZN(new_n359_) );
  OR4_X1 g0223 ( .A1(new_n356_), .A2(new_n357_), .A3(new_n358_), .A4(new_n359_), .ZN(new_n360_) );
  INV_X1 g0224 ( .A(new_n360_), .ZN(new_n361_) );
  AND3_X1 g0225 ( .A1(new_n354_), .A2(new_n352_), .A3(new_n361_), .ZN(new_n362_) );
  INV_X1 g0226 ( .A(new_n362_), .ZN(new_n363_) );
  AND2_X1 g0227 ( .A1(new_n351_), .A2(G179), .ZN(new_n364_) );
  INV_X1 g0228 ( .A(new_n364_), .ZN(new_n365_) );
  OR2_X1 g0229 ( .A1(new_n351_), .A2(new_n330_), .ZN(new_n366_) );
  AND2_X1 g0230 ( .A1(new_n365_), .A2(new_n366_), .ZN(new_n367_) );
  INV_X1 g0231 ( .A(new_n367_), .ZN(new_n368_) );
  AND2_X1 g0232 ( .A1(new_n368_), .A2(new_n360_), .ZN(new_n369_) );
  INV_X1 g0233 ( .A(new_n369_), .ZN(new_n370_) );
  AND2_X1 g0234 ( .A1(new_n370_), .A2(new_n363_), .ZN(new_n371_) );
  OR2_X1 g0235 ( .A1(new_n327_), .A2(new_n337_), .ZN(new_n372_) );
  AND2_X1 g0236 ( .A1(new_n372_), .A2(KEYINPUT35), .ZN(new_n373_) );
  OR2_X1 g0237 ( .A1(new_n372_), .A2(KEYINPUT35), .ZN(new_n374_) );
  INV_X1 g0238 ( .A(new_n374_), .ZN(new_n375_) );
  AND2_X1 g0239 ( .A1(new_n327_), .A2(G190), .ZN(new_n376_) );
  OR4_X1 g0240 ( .A1(new_n375_), .A2(new_n289_), .A3(new_n373_), .A4(new_n376_), .ZN(new_n377_) );
  INV_X1 g0241 ( .A(KEYINPUT37), .ZN(new_n378_) );
  AND2_X1 g0242 ( .A1(new_n355_), .A2(G50), .ZN(new_n379_) );
  INV_X1 g0243 ( .A(new_n139_), .ZN(new_n380_) );
  AND2_X1 g0244 ( .A1(new_n268_), .A2(new_n380_), .ZN(new_n381_) );
  AND2_X1 g0245 ( .A1(new_n276_), .A2(G150), .ZN(new_n382_) );
  AND2_X1 g0246 ( .A1(new_n280_), .A2(G58), .ZN(new_n383_) );
  AND2_X1 g0247 ( .A1(new_n282_), .A2(new_n140_), .ZN(new_n384_) );
  OR3_X1 g0248 ( .A1(new_n382_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_) );
  OR3_X1 g0249 ( .A1(new_n379_), .A2(new_n381_), .A3(new_n385_), .ZN(new_n386_) );
  INV_X1 g0250 ( .A(G179), .ZN(new_n387_) );
  INV_X1 g0251 ( .A(KEYINPUT36), .ZN(new_n388_) );
  AND2_X1 g0252 ( .A1(new_n299_), .A2(G222), .ZN(new_n389_) );
  AND2_X1 g0253 ( .A1(new_n389_), .A2(new_n388_), .ZN(new_n390_) );
  INV_X1 g0254 ( .A(new_n390_), .ZN(new_n391_) );
  OR2_X1 g0255 ( .A1(new_n389_), .A2(new_n388_), .ZN(new_n392_) );
  AND2_X1 g0256 ( .A1(new_n391_), .A2(new_n392_), .ZN(new_n393_) );
  AND2_X1 g0257 ( .A1(new_n294_), .A2(G223), .ZN(new_n394_) );
  AND2_X1 g0258 ( .A1(new_n323_), .A2(G226), .ZN(new_n395_) );
  AND2_X1 g0259 ( .A1(new_n307_), .A2(G77), .ZN(new_n396_) );
  OR4_X1 g0260 ( .A1(new_n395_), .A2(new_n394_), .A3(new_n396_), .A4(new_n318_), .ZN(new_n397_) );
  OR2_X1 g0261 ( .A1(new_n393_), .A2(new_n397_), .ZN(new_n398_) );
  INV_X1 g0262 ( .A(new_n398_), .ZN(new_n399_) );
  AND2_X1 g0263 ( .A1(new_n399_), .A2(new_n387_), .ZN(new_n400_) );
  INV_X1 g0264 ( .A(new_n400_), .ZN(new_n401_) );
  AND2_X1 g0265 ( .A1(new_n398_), .A2(new_n330_), .ZN(new_n402_) );
  INV_X1 g0266 ( .A(new_n402_), .ZN(new_n403_) );
  AND3_X1 g0267 ( .A1(new_n401_), .A2(new_n386_), .A3(new_n403_), .ZN(new_n404_) );
  INV_X1 g0268 ( .A(new_n404_), .ZN(new_n405_) );
  AND2_X1 g0269 ( .A1(new_n399_), .A2(G190), .ZN(new_n406_) );
  AND2_X1 g0270 ( .A1(new_n398_), .A2(G200), .ZN(new_n407_) );
  OR3_X1 g0271 ( .A1(new_n386_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_) );
  AND2_X1 g0272 ( .A1(new_n405_), .A2(new_n408_), .ZN(new_n409_) );
  AND2_X1 g0273 ( .A1(new_n409_), .A2(new_n378_), .ZN(new_n410_) );
  INV_X1 g0274 ( .A(new_n409_), .ZN(new_n411_) );
  AND2_X1 g0275 ( .A1(new_n411_), .A2(KEYINPUT37), .ZN(new_n412_) );
  OR2_X1 g0276 ( .A1(new_n412_), .A2(new_n410_), .ZN(new_n413_) );
  OR2_X1 g0277 ( .A1(new_n268_), .A2(new_n282_), .ZN(new_n414_) );
  AND2_X1 g0278 ( .A1(new_n414_), .A2(new_n138_), .ZN(new_n415_) );
  AND2_X1 g0279 ( .A1(new_n273_), .A2(G68), .ZN(new_n416_) );
  AND2_X1 g0280 ( .A1(new_n276_), .A2(G50), .ZN(new_n417_) );
  AND2_X1 g0281 ( .A1(new_n280_), .A2(G77), .ZN(new_n418_) );
  OR3_X1 g0282 ( .A1(new_n416_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_) );
  OR2_X1 g0283 ( .A1(new_n415_), .A2(new_n419_), .ZN(new_n420_) );
  INV_X1 g0284 ( .A(KEYINPUT28), .ZN(new_n421_) );
  OR2_X1 g0285 ( .A1(new_n298_), .A2(new_n197_), .ZN(new_n422_) );
  OR2_X1 g0286 ( .A1(new_n306_), .A2(new_n144_), .ZN(new_n423_) );
  AND3_X1 g0287 ( .A1(new_n422_), .A2(new_n423_), .A3(new_n319_), .ZN(new_n424_) );
  AND2_X1 g0288 ( .A1(new_n323_), .A2(G238), .ZN(new_n425_) );
  INV_X1 g0289 ( .A(new_n425_), .ZN(new_n426_) );
  AND2_X1 g0290 ( .A1(new_n294_), .A2(G232), .ZN(new_n427_) );
  INV_X1 g0291 ( .A(new_n427_), .ZN(new_n428_) );
  AND3_X1 g0292 ( .A1(new_n424_), .A2(new_n426_), .A3(new_n428_), .ZN(new_n429_) );
  AND2_X1 g0293 ( .A1(new_n429_), .A2(G190), .ZN(new_n430_) );
  INV_X1 g0294 ( .A(new_n430_), .ZN(new_n431_) );
  AND2_X1 g0295 ( .A1(new_n431_), .A2(new_n421_), .ZN(new_n432_) );
  AND2_X1 g0296 ( .A1(new_n430_), .A2(KEYINPUT28), .ZN(new_n433_) );
  OR2_X1 g0297 ( .A1(new_n432_), .A2(new_n433_), .ZN(new_n434_) );
  INV_X1 g0298 ( .A(KEYINPUT27), .ZN(new_n435_) );
  INV_X1 g0299 ( .A(new_n429_), .ZN(new_n436_) );
  AND2_X1 g0300 ( .A1(new_n436_), .A2(G200), .ZN(new_n437_) );
  AND2_X1 g0301 ( .A1(new_n437_), .A2(new_n435_), .ZN(new_n438_) );
  OR2_X1 g0302 ( .A1(new_n437_), .A2(new_n435_), .ZN(new_n439_) );
  INV_X1 g0303 ( .A(new_n439_), .ZN(new_n440_) );
  OR4_X1 g0304 ( .A1(new_n434_), .A2(new_n420_), .A3(new_n440_), .A4(new_n438_), .ZN(new_n441_) );
  INV_X1 g0305 ( .A(new_n420_), .ZN(new_n442_) );
  AND2_X1 g0306 ( .A1(new_n429_), .A2(new_n387_), .ZN(new_n443_) );
  AND2_X1 g0307 ( .A1(new_n436_), .A2(new_n330_), .ZN(new_n444_) );
  OR3_X1 g0308 ( .A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_) );
  AND2_X1 g0309 ( .A1(new_n441_), .A2(new_n445_), .ZN(new_n446_) );
  AND4_X1 g0310 ( .A1(new_n413_), .A2(new_n371_), .A3(new_n377_), .A4(new_n446_), .ZN(new_n447_) );
  AND2_X1 g0311 ( .A1(new_n447_), .A2(new_n336_), .ZN(new_n448_) );
  INV_X1 g0312 ( .A(KEYINPUT16), .ZN(new_n449_) );
  INV_X1 g0313 ( .A(new_n278_), .ZN(new_n450_) );
  AND3_X1 g0314 ( .A1(new_n264_), .A2(G116), .A3(new_n450_), .ZN(new_n451_) );
  OR2_X1 g0315 ( .A1(new_n451_), .A2(new_n449_), .ZN(new_n452_) );
  AND4_X1 g0316 ( .A1(new_n264_), .A2(G116), .A3(new_n449_), .A4(new_n450_), .ZN(new_n453_) );
  INV_X1 g0317 ( .A(new_n453_), .ZN(new_n454_) );
  AND2_X1 g0318 ( .A1(new_n452_), .A2(new_n454_), .ZN(new_n455_) );
  INV_X1 g0319 ( .A(new_n282_), .ZN(new_n456_) );
  AND2_X1 g0320 ( .A1(new_n270_), .A2(G33), .ZN(new_n457_) );
  INV_X1 g0321 ( .A(new_n457_), .ZN(new_n458_) );
  AND4_X1 g0322 ( .A1(new_n260_), .A2(new_n180_), .A3(new_n456_), .A4(new_n458_), .ZN(new_n459_) );
  AND2_X1 g0323 ( .A1(new_n459_), .A2(G107), .ZN(new_n460_) );
  OR3_X1 g0324 ( .A1(new_n455_), .A2(new_n460_), .A3(KEYINPUT17), .ZN(new_n461_) );
  INV_X1 g0325 ( .A(new_n461_), .ZN(new_n462_) );
  OR2_X1 g0326 ( .A1(new_n455_), .A2(new_n460_), .ZN(new_n463_) );
  AND2_X1 g0327 ( .A1(new_n463_), .A2(KEYINPUT17), .ZN(new_n464_) );
  OR2_X1 g0328 ( .A1(new_n464_), .A2(new_n462_), .ZN(new_n465_) );
  INV_X1 g0329 ( .A(new_n262_), .ZN(new_n466_) );
  OR2_X1 g0330 ( .A1(new_n261_), .A2(new_n175_), .ZN(new_n467_) );
  AND2_X1 g0331 ( .A1(new_n467_), .A2(KEYINPUT4), .ZN(new_n468_) );
  OR2_X1 g0332 ( .A1(new_n468_), .A2(new_n466_), .ZN(new_n469_) );
  AND2_X1 g0333 ( .A1(new_n469_), .A2(new_n456_), .ZN(new_n470_) );
  OR2_X1 g0334 ( .A1(new_n470_), .A2(G107), .ZN(new_n471_) );
  AND2_X1 g0335 ( .A1(new_n276_), .A2(G87), .ZN(new_n472_) );
  INV_X1 g0336 ( .A(new_n472_), .ZN(new_n473_) );
  AND3_X1 g0337 ( .A1(new_n471_), .A2(new_n465_), .A3(new_n473_), .ZN(new_n474_) );
  AND2_X1 g0338 ( .A1(new_n270_), .A2(G45), .ZN(new_n475_) );
  AND3_X1 g0339 ( .A1(new_n475_), .A2(new_n314_), .A3(G274), .ZN(new_n476_) );
  INV_X1 g0340 ( .A(new_n475_), .ZN(new_n477_) );
  OR2_X1 g0341 ( .A1(new_n477_), .A2(G41), .ZN(new_n478_) );
  AND3_X1 g0342 ( .A1(new_n322_), .A2(G264), .A3(new_n478_), .ZN(new_n479_) );
  OR2_X1 g0343 ( .A1(new_n479_), .A2(new_n476_), .ZN(new_n480_) );
  AND4_X1 g0344 ( .A1(new_n264_), .A2(G33), .A3(new_n314_), .A4(G294), .ZN(new_n481_) );
  AND2_X1 g0345 ( .A1(new_n481_), .A2(KEYINPUT14), .ZN(new_n482_) );
  INV_X1 g0346 ( .A(KEYINPUT14), .ZN(new_n483_) );
  INV_X1 g0347 ( .A(G294), .ZN(new_n484_) );
  OR4_X1 g0348 ( .A1(new_n180_), .A2(new_n275_), .A3(G41), .A4(new_n484_), .ZN(new_n485_) );
  AND2_X1 g0349 ( .A1(new_n485_), .A2(new_n483_), .ZN(new_n486_) );
  OR2_X1 g0350 ( .A1(new_n482_), .A2(new_n486_), .ZN(new_n487_) );
  AND4_X1 g0351 ( .A1(new_n264_), .A2(new_n275_), .A3(G250), .A4(new_n292_), .ZN(new_n488_) );
  AND4_X1 g0352 ( .A1(new_n264_), .A2(new_n275_), .A3(G257), .A4(G1698), .ZN(new_n489_) );
  OR2_X1 g0353 ( .A1(new_n488_), .A2(new_n489_), .ZN(new_n490_) );
  OR4_X1 g0354 ( .A1(new_n487_), .A2(G179), .A3(new_n480_), .A4(new_n490_), .ZN(new_n491_) );
  AND2_X1 g0355 ( .A1(new_n491_), .A2(KEYINPUT15), .ZN(new_n492_) );
  INV_X1 g0356 ( .A(KEYINPUT15), .ZN(new_n493_) );
  INV_X1 g0357 ( .A(new_n480_), .ZN(new_n494_) );
  OR2_X1 g0358 ( .A1(new_n485_), .A2(new_n483_), .ZN(new_n495_) );
  OR2_X1 g0359 ( .A1(new_n481_), .A2(KEYINPUT14), .ZN(new_n496_) );
  INV_X1 g0360 ( .A(new_n488_), .ZN(new_n497_) );
  INV_X1 g0361 ( .A(new_n489_), .ZN(new_n498_) );
  AND4_X1 g0362 ( .A1(new_n496_), .A2(new_n495_), .A3(new_n497_), .A4(new_n498_), .ZN(new_n499_) );
  AND3_X1 g0363 ( .A1(new_n499_), .A2(new_n387_), .A3(new_n494_), .ZN(new_n500_) );
  AND2_X1 g0364 ( .A1(new_n500_), .A2(new_n493_), .ZN(new_n501_) );
  OR3_X1 g0365 ( .A1(new_n487_), .A2(new_n480_), .A3(new_n490_), .ZN(new_n502_) );
  AND2_X1 g0366 ( .A1(new_n502_), .A2(new_n330_), .ZN(new_n503_) );
  OR3_X1 g0367 ( .A1(new_n492_), .A2(new_n501_), .A3(new_n503_), .ZN(new_n504_) );
  OR2_X1 g0368 ( .A1(new_n474_), .A2(new_n504_), .ZN(new_n505_) );
  INV_X1 g0369 ( .A(KEYINPUT17), .ZN(new_n506_) );
  OR3_X1 g0370 ( .A1(new_n180_), .A2(new_n232_), .A3(new_n278_), .ZN(new_n507_) );
  AND2_X1 g0371 ( .A1(new_n507_), .A2(KEYINPUT16), .ZN(new_n508_) );
  OR2_X1 g0372 ( .A1(new_n508_), .A2(new_n453_), .ZN(new_n509_) );
  OR4_X1 g0373 ( .A1(new_n265_), .A2(new_n145_), .A3(new_n282_), .A4(new_n457_), .ZN(new_n510_) );
  AND2_X1 g0374 ( .A1(new_n509_), .A2(new_n510_), .ZN(new_n511_) );
  OR2_X1 g0375 ( .A1(new_n511_), .A2(new_n506_), .ZN(new_n512_) );
  AND2_X1 g0376 ( .A1(new_n512_), .A2(new_n461_), .ZN(new_n513_) );
  AND2_X1 g0377 ( .A1(new_n414_), .A2(new_n145_), .ZN(new_n514_) );
  OR3_X1 g0378 ( .A1(new_n514_), .A2(new_n513_), .A3(new_n472_), .ZN(new_n515_) );
  AND2_X1 g0379 ( .A1(new_n499_), .A2(new_n494_), .ZN(new_n516_) );
  OR2_X1 g0380 ( .A1(new_n516_), .A2(new_n337_), .ZN(new_n517_) );
  AND2_X1 g0381 ( .A1(new_n516_), .A2(G190), .ZN(new_n518_) );
  INV_X1 g0382 ( .A(new_n518_), .ZN(new_n519_) );
  AND2_X1 g0383 ( .A1(new_n519_), .A2(new_n517_), .ZN(new_n520_) );
  INV_X1 g0384 ( .A(new_n520_), .ZN(new_n521_) );
  OR2_X1 g0385 ( .A1(new_n515_), .A2(new_n521_), .ZN(new_n522_) );
  AND3_X1 g0386 ( .A1(new_n522_), .A2(new_n505_), .A3(KEYINPUT0), .ZN(new_n523_) );
  INV_X1 g0387 ( .A(KEYINPUT0), .ZN(new_n524_) );
  OR2_X1 g0388 ( .A1(new_n500_), .A2(new_n493_), .ZN(new_n525_) );
  INV_X1 g0389 ( .A(new_n501_), .ZN(new_n526_) );
  INV_X1 g0390 ( .A(new_n503_), .ZN(new_n527_) );
  AND3_X1 g0391 ( .A1(new_n526_), .A2(new_n527_), .A3(new_n525_), .ZN(new_n528_) );
  AND2_X1 g0392 ( .A1(new_n515_), .A2(new_n528_), .ZN(new_n529_) );
  AND4_X1 g0393 ( .A1(new_n520_), .A2(new_n465_), .A3(new_n471_), .A4(new_n473_), .ZN(new_n530_) );
  OR2_X1 g0394 ( .A1(new_n529_), .A2(new_n530_), .ZN(new_n531_) );
  AND2_X1 g0395 ( .A1(new_n531_), .A2(new_n524_), .ZN(new_n532_) );
  OR2_X1 g0396 ( .A1(new_n532_), .A2(new_n523_), .ZN(new_n533_) );
  INV_X1 g0397 ( .A(KEYINPUT12), .ZN(new_n534_) );
  INV_X1 g0398 ( .A(new_n476_), .ZN(new_n535_) );
  OR2_X1 g0399 ( .A1(new_n293_), .A2(new_n208_), .ZN(new_n536_) );
  OR2_X1 g0400 ( .A1(new_n298_), .A2(new_n191_), .ZN(new_n537_) );
  INV_X1 g0401 ( .A(G283), .ZN(new_n538_) );
  OR2_X1 g0402 ( .A1(new_n306_), .A2(new_n538_), .ZN(new_n539_) );
  AND4_X1 g0403 ( .A1(new_n536_), .A2(new_n537_), .A3(new_n539_), .A4(new_n535_), .ZN(new_n540_) );
  AND2_X1 g0404 ( .A1(new_n540_), .A2(new_n534_), .ZN(new_n541_) );
  INV_X1 g0405 ( .A(new_n541_), .ZN(new_n542_) );
  OR2_X1 g0406 ( .A1(new_n540_), .A2(new_n534_), .ZN(new_n543_) );
  AND2_X1 g0407 ( .A1(new_n322_), .A2(new_n478_), .ZN(new_n544_) );
  AND2_X1 g0408 ( .A1(new_n544_), .A2(G257), .ZN(new_n545_) );
  INV_X1 g0409 ( .A(new_n545_), .ZN(new_n546_) );
  AND3_X1 g0410 ( .A1(new_n542_), .A2(new_n543_), .A3(new_n546_), .ZN(new_n547_) );
  OR2_X1 g0411 ( .A1(new_n547_), .A2(G169), .ZN(new_n548_) );
  AND2_X1 g0412 ( .A1(new_n547_), .A2(new_n387_), .ZN(new_n549_) );
  INV_X1 g0413 ( .A(new_n549_), .ZN(new_n550_) );
  AND2_X1 g0414 ( .A1(new_n268_), .A2(new_n225_), .ZN(new_n551_) );
  INV_X1 g0415 ( .A(KEYINPUT13), .ZN(new_n552_) );
  AND2_X1 g0416 ( .A1(new_n280_), .A2(G107), .ZN(new_n553_) );
  AND2_X1 g0417 ( .A1(new_n282_), .A2(new_n144_), .ZN(new_n554_) );
  OR2_X1 g0418 ( .A1(new_n553_), .A2(new_n554_), .ZN(new_n555_) );
  INV_X1 g0419 ( .A(new_n555_), .ZN(new_n556_) );
  AND2_X1 g0420 ( .A1(new_n556_), .A2(new_n552_), .ZN(new_n557_) );
  AND2_X1 g0421 ( .A1(new_n555_), .A2(KEYINPUT13), .ZN(new_n558_) );
  OR2_X1 g0422 ( .A1(new_n557_), .A2(new_n558_), .ZN(new_n559_) );
  INV_X1 g0423 ( .A(new_n559_), .ZN(new_n560_) );
  AND2_X1 g0424 ( .A1(new_n459_), .A2(G97), .ZN(new_n561_) );
  AND2_X1 g0425 ( .A1(new_n276_), .A2(G77), .ZN(new_n562_) );
  OR4_X1 g0426 ( .A1(new_n560_), .A2(new_n551_), .A3(new_n561_), .A4(new_n562_), .ZN(new_n563_) );
  AND3_X1 g0427 ( .A1(new_n563_), .A2(new_n548_), .A3(new_n550_), .ZN(new_n564_) );
  INV_X1 g0428 ( .A(new_n563_), .ZN(new_n565_) );
  OR2_X1 g0429 ( .A1(new_n547_), .A2(new_n337_), .ZN(new_n566_) );
  AND2_X1 g0430 ( .A1(new_n547_), .A2(G190), .ZN(new_n567_) );
  INV_X1 g0431 ( .A(new_n567_), .ZN(new_n568_) );
  AND3_X1 g0432 ( .A1(new_n565_), .A2(new_n566_), .A3(new_n568_), .ZN(new_n569_) );
  OR2_X1 g0433 ( .A1(new_n569_), .A2(new_n564_), .ZN(new_n570_) );
  INV_X1 g0434 ( .A(new_n570_), .ZN(new_n571_) );
  INV_X1 g0435 ( .A(KEYINPUT9), .ZN(new_n572_) );
  AND2_X1 g0436 ( .A1(new_n459_), .A2(G87), .ZN(new_n573_) );
  OR2_X1 g0437 ( .A1(new_n268_), .A2(new_n573_), .ZN(new_n574_) );
  AND2_X1 g0438 ( .A1(new_n146_), .A2(new_n231_), .ZN(new_n575_) );
  INV_X1 g0439 ( .A(new_n575_), .ZN(new_n576_) );
  AND2_X1 g0440 ( .A1(new_n574_), .A2(new_n576_), .ZN(new_n577_) );
  OR2_X1 g0441 ( .A1(new_n577_), .A2(new_n572_), .ZN(new_n578_) );
  INV_X1 g0442 ( .A(new_n578_), .ZN(new_n579_) );
  AND2_X1 g0443 ( .A1(new_n577_), .A2(new_n572_), .ZN(new_n580_) );
  AND2_X1 g0444 ( .A1(new_n276_), .A2(G68), .ZN(new_n581_) );
  AND2_X1 g0445 ( .A1(new_n280_), .A2(G97), .ZN(new_n582_) );
  AND2_X1 g0446 ( .A1(new_n282_), .A2(new_n231_), .ZN(new_n583_) );
  OR3_X1 g0447 ( .A1(new_n581_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_) );
  OR3_X1 g0448 ( .A1(new_n579_), .A2(new_n580_), .A3(new_n584_), .ZN(new_n585_) );
  INV_X1 g0449 ( .A(KEYINPUT8), .ZN(new_n586_) );
  AND2_X1 g0450 ( .A1(new_n294_), .A2(G244), .ZN(new_n587_) );
  AND2_X1 g0451 ( .A1(new_n299_), .A2(G238), .ZN(new_n588_) );
  OR2_X1 g0452 ( .A1(new_n587_), .A2(new_n588_), .ZN(new_n589_) );
  INV_X1 g0453 ( .A(new_n589_), .ZN(new_n590_) );
  AND2_X1 g0454 ( .A1(new_n590_), .A2(new_n586_), .ZN(new_n591_) );
  INV_X1 g0455 ( .A(new_n591_), .ZN(new_n592_) );
  AND2_X1 g0456 ( .A1(new_n589_), .A2(KEYINPUT8), .ZN(new_n593_) );
  INV_X1 g0457 ( .A(new_n593_), .ZN(new_n594_) );
  AND3_X1 g0458 ( .A1(new_n322_), .A2(G250), .A3(new_n477_), .ZN(new_n595_) );
  AND2_X1 g0459 ( .A1(new_n307_), .A2(G116), .ZN(new_n596_) );
  AND2_X1 g0460 ( .A1(new_n475_), .A2(G274), .ZN(new_n597_) );
  OR3_X1 g0461 ( .A1(new_n596_), .A2(new_n595_), .A3(new_n597_), .ZN(new_n598_) );
  INV_X1 g0462 ( .A(new_n598_), .ZN(new_n599_) );
  AND3_X1 g0463 ( .A1(new_n592_), .A2(new_n594_), .A3(new_n599_), .ZN(new_n600_) );
  AND2_X1 g0464 ( .A1(new_n600_), .A2(G190), .ZN(new_n601_) );
  INV_X1 g0465 ( .A(new_n600_), .ZN(new_n602_) );
  AND2_X1 g0466 ( .A1(new_n602_), .A2(G200), .ZN(new_n603_) );
  OR3_X1 g0467 ( .A1(new_n585_), .A2(new_n601_), .A3(new_n603_), .ZN(new_n604_) );
  INV_X1 g0468 ( .A(new_n585_), .ZN(new_n605_) );
  OR2_X1 g0469 ( .A1(new_n600_), .A2(new_n330_), .ZN(new_n606_) );
  AND2_X1 g0470 ( .A1(new_n600_), .A2(G179), .ZN(new_n607_) );
  INV_X1 g0471 ( .A(new_n607_), .ZN(new_n608_) );
  AND2_X1 g0472 ( .A1(new_n608_), .A2(new_n606_), .ZN(new_n609_) );
  OR2_X1 g0473 ( .A1(new_n605_), .A2(new_n609_), .ZN(new_n610_) );
  AND2_X1 g0474 ( .A1(new_n610_), .A2(new_n604_), .ZN(new_n611_) );
  INV_X1 g0475 ( .A(KEYINPUT11), .ZN(new_n612_) );
  OR2_X1 g0476 ( .A1(new_n268_), .A2(new_n459_), .ZN(new_n613_) );
  AND2_X1 g0477 ( .A1(new_n613_), .A2(G116), .ZN(new_n614_) );
  AND2_X1 g0478 ( .A1(new_n276_), .A2(G97), .ZN(new_n615_) );
  AND2_X1 g0479 ( .A1(new_n280_), .A2(G283), .ZN(new_n616_) );
  AND2_X1 g0480 ( .A1(new_n282_), .A2(new_n232_), .ZN(new_n617_) );
  OR3_X1 g0481 ( .A1(new_n615_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n618_) );
  OR2_X1 g0482 ( .A1(new_n614_), .A2(new_n618_), .ZN(new_n619_) );
  OR2_X1 g0483 ( .A1(new_n298_), .A2(new_n209_), .ZN(new_n620_) );
  INV_X1 g0484 ( .A(G264), .ZN(new_n621_) );
  OR2_X1 g0485 ( .A1(new_n293_), .A2(new_n621_), .ZN(new_n622_) );
  INV_X1 g0486 ( .A(G303), .ZN(new_n623_) );
  OR2_X1 g0487 ( .A1(new_n306_), .A2(new_n623_), .ZN(new_n624_) );
  AND4_X1 g0488 ( .A1(new_n620_), .A2(new_n622_), .A3(new_n624_), .A4(new_n535_), .ZN(new_n625_) );
  AND2_X1 g0489 ( .A1(new_n544_), .A2(G270), .ZN(new_n626_) );
  OR2_X1 g0490 ( .A1(new_n626_), .A2(KEYINPUT10), .ZN(new_n627_) );
  AND2_X1 g0491 ( .A1(new_n626_), .A2(KEYINPUT10), .ZN(new_n628_) );
  INV_X1 g0492 ( .A(new_n628_), .ZN(new_n629_) );
  AND3_X1 g0493 ( .A1(new_n629_), .A2(new_n625_), .A3(new_n627_), .ZN(new_n630_) );
  AND2_X1 g0494 ( .A1(new_n630_), .A2(G190), .ZN(new_n631_) );
  INV_X1 g0495 ( .A(new_n630_), .ZN(new_n632_) );
  AND2_X1 g0496 ( .A1(new_n632_), .A2(G200), .ZN(new_n633_) );
  OR3_X1 g0497 ( .A1(new_n619_), .A2(new_n631_), .A3(new_n633_), .ZN(new_n634_) );
  INV_X1 g0498 ( .A(new_n619_), .ZN(new_n635_) );
  OR2_X1 g0499 ( .A1(new_n630_), .A2(new_n330_), .ZN(new_n636_) );
  AND2_X1 g0500 ( .A1(new_n630_), .A2(G179), .ZN(new_n637_) );
  INV_X1 g0501 ( .A(new_n637_), .ZN(new_n638_) );
  AND2_X1 g0502 ( .A1(new_n638_), .A2(new_n636_), .ZN(new_n639_) );
  OR2_X1 g0503 ( .A1(new_n635_), .A2(new_n639_), .ZN(new_n640_) );
  AND3_X1 g0504 ( .A1(new_n640_), .A2(new_n634_), .A3(new_n612_), .ZN(new_n641_) );
  INV_X1 g0505 ( .A(new_n631_), .ZN(new_n642_) );
  INV_X1 g0506 ( .A(new_n633_), .ZN(new_n643_) );
  AND3_X1 g0507 ( .A1(new_n635_), .A2(new_n642_), .A3(new_n643_), .ZN(new_n644_) );
  INV_X1 g0508 ( .A(new_n639_), .ZN(new_n645_) );
  AND2_X1 g0509 ( .A1(new_n645_), .A2(new_n619_), .ZN(new_n646_) );
  OR2_X1 g0510 ( .A1(new_n646_), .A2(new_n644_), .ZN(new_n647_) );
  AND2_X1 g0511 ( .A1(new_n647_), .A2(KEYINPUT11), .ZN(new_n648_) );
  OR2_X1 g0512 ( .A1(new_n648_), .A2(new_n641_), .ZN(new_n649_) );
  AND2_X1 g0513 ( .A1(new_n649_), .A2(new_n611_), .ZN(new_n650_) );
  AND4_X1 g0514 ( .A1(new_n448_), .A2(new_n533_), .A3(new_n571_), .A4(new_n650_), .ZN(G372) );
  INV_X1 g0515 ( .A(new_n336_), .ZN(new_n652_) );
  INV_X1 g0516 ( .A(new_n445_), .ZN(new_n653_) );
  AND2_X1 g0517 ( .A1(new_n369_), .A2(new_n446_), .ZN(new_n654_) );
  OR2_X1 g0518 ( .A1(new_n654_), .A2(new_n653_), .ZN(new_n655_) );
  AND2_X1 g0519 ( .A1(new_n655_), .A2(new_n377_), .ZN(new_n656_) );
  OR2_X1 g0520 ( .A1(new_n656_), .A2(new_n652_), .ZN(new_n657_) );
  AND2_X1 g0521 ( .A1(new_n657_), .A2(new_n413_), .ZN(new_n658_) );
  OR2_X1 g0522 ( .A1(new_n658_), .A2(new_n404_), .ZN(new_n659_) );
  AND2_X1 g0523 ( .A1(new_n533_), .A2(new_n646_), .ZN(new_n660_) );
  OR2_X1 g0524 ( .A1(new_n660_), .A2(new_n529_), .ZN(new_n661_) );
  AND2_X1 g0525 ( .A1(new_n661_), .A2(new_n571_), .ZN(new_n662_) );
  INV_X1 g0526 ( .A(new_n610_), .ZN(new_n663_) );
  OR2_X1 g0527 ( .A1(new_n663_), .A2(new_n564_), .ZN(new_n664_) );
  OR2_X1 g0528 ( .A1(new_n662_), .A2(new_n664_), .ZN(new_n665_) );
  AND2_X1 g0529 ( .A1(new_n665_), .A2(new_n604_), .ZN(new_n666_) );
  AND2_X1 g0530 ( .A1(new_n666_), .A2(new_n448_), .ZN(new_n667_) );
  OR2_X1 g0531 ( .A1(new_n667_), .A2(new_n659_), .ZN(G369) );
  AND4_X1 g0532 ( .A1(new_n270_), .A2(new_n175_), .A3(G13), .A4(G213), .ZN(new_n669_) );
  AND2_X1 g0533 ( .A1(new_n669_), .A2(G343), .ZN(new_n670_) );
  AND2_X1 g0534 ( .A1(new_n515_), .A2(new_n670_), .ZN(new_n671_) );
  INV_X1 g0535 ( .A(new_n671_), .ZN(new_n672_) );
  AND2_X1 g0536 ( .A1(new_n533_), .A2(new_n672_), .ZN(new_n673_) );
  AND2_X1 g0537 ( .A1(new_n529_), .A2(new_n670_), .ZN(new_n674_) );
  OR2_X1 g0538 ( .A1(new_n673_), .A2(new_n674_), .ZN(new_n675_) );
  AND2_X1 g0539 ( .A1(new_n619_), .A2(new_n670_), .ZN(new_n676_) );
  INV_X1 g0540 ( .A(new_n676_), .ZN(new_n677_) );
  AND2_X1 g0541 ( .A1(new_n649_), .A2(new_n677_), .ZN(new_n678_) );
  AND2_X1 g0542 ( .A1(new_n646_), .A2(new_n670_), .ZN(new_n679_) );
  OR2_X1 g0543 ( .A1(new_n678_), .A2(new_n679_), .ZN(new_n680_) );
  AND2_X1 g0544 ( .A1(new_n680_), .A2(G330), .ZN(new_n681_) );
  AND2_X1 g0545 ( .A1(new_n681_), .A2(new_n675_), .ZN(new_n682_) );
  INV_X1 g0546 ( .A(new_n670_), .ZN(new_n683_) );
  AND2_X1 g0547 ( .A1(new_n661_), .A2(new_n683_), .ZN(new_n684_) );
  OR2_X1 g0548 ( .A1(new_n682_), .A2(new_n684_), .ZN(G399) );
  AND4_X1 g0549 ( .A1(new_n650_), .A2(new_n533_), .A3(new_n571_), .A4(new_n683_), .ZN(new_n686_) );
  INV_X1 g0550 ( .A(KEYINPUT18), .ZN(new_n687_) );
  AND2_X1 g0551 ( .A1(new_n600_), .A2(new_n547_), .ZN(new_n688_) );
  AND2_X1 g0552 ( .A1(new_n688_), .A2(new_n687_), .ZN(new_n689_) );
  INV_X1 g0553 ( .A(new_n689_), .ZN(new_n690_) );
  OR2_X1 g0554 ( .A1(new_n688_), .A2(new_n687_), .ZN(new_n691_) );
  AND4_X1 g0555 ( .A1(new_n690_), .A2(new_n516_), .A3(new_n637_), .A4(new_n691_), .ZN(new_n692_) );
  INV_X1 g0556 ( .A(new_n547_), .ZN(new_n693_) );
  AND2_X1 g0557 ( .A1(new_n632_), .A2(new_n387_), .ZN(new_n694_) );
  AND4_X1 g0558 ( .A1(new_n602_), .A2(new_n502_), .A3(new_n693_), .A4(new_n694_), .ZN(new_n695_) );
  OR2_X1 g0559 ( .A1(new_n692_), .A2(new_n695_), .ZN(new_n696_) );
  AND2_X1 g0560 ( .A1(new_n696_), .A2(new_n670_), .ZN(new_n697_) );
  OR2_X1 g0561 ( .A1(new_n686_), .A2(new_n697_), .ZN(new_n698_) );
  AND2_X1 g0562 ( .A1(new_n698_), .A2(G330), .ZN(new_n699_) );
  AND2_X1 g0563 ( .A1(new_n666_), .A2(new_n683_), .ZN(new_n700_) );
  OR2_X1 g0564 ( .A1(new_n700_), .A2(new_n699_), .ZN(new_n701_) );
  AND2_X1 g0565 ( .A1(new_n701_), .A2(new_n270_), .ZN(new_n702_) );
  AND2_X1 g0566 ( .A1(new_n575_), .A2(new_n232_), .ZN(new_n703_) );
  AND2_X1 g0567 ( .A1(new_n184_), .A2(new_n314_), .ZN(new_n704_) );
  INV_X1 g0568 ( .A(new_n704_), .ZN(new_n705_) );
  AND3_X1 g0569 ( .A1(new_n703_), .A2(new_n705_), .A3(G1), .ZN(new_n706_) );
  AND3_X1 g0570 ( .A1(new_n704_), .A2(G50), .A3(new_n380_), .ZN(new_n707_) );
  OR3_X1 g0571 ( .A1(new_n702_), .A2(new_n706_), .A3(new_n707_), .ZN(G364) );
  INV_X1 g0572 ( .A(new_n680_), .ZN(new_n709_) );
  AND2_X1 g0573 ( .A1(new_n183_), .A2(new_n275_), .ZN(new_n710_) );
  AND2_X1 g0574 ( .A1(new_n710_), .A2(new_n175_), .ZN(new_n711_) );
  AND2_X1 g0575 ( .A1(new_n709_), .A2(new_n711_), .ZN(new_n712_) );
  AND2_X1 g0576 ( .A1(new_n712_), .A2(KEYINPUT62), .ZN(new_n713_) );
  INV_X1 g0577 ( .A(new_n713_), .ZN(new_n714_) );
  OR2_X1 g0578 ( .A1(new_n712_), .A2(KEYINPUT62), .ZN(new_n715_) );
  INV_X1 g0579 ( .A(G190), .ZN(new_n716_) );
  AND2_X1 g0580 ( .A1(new_n387_), .A2(G20), .ZN(new_n717_) );
  AND2_X1 g0581 ( .A1(new_n717_), .A2(new_n716_), .ZN(new_n718_) );
  AND2_X1 g0582 ( .A1(new_n718_), .A2(new_n337_), .ZN(new_n719_) );
  AND2_X1 g0583 ( .A1(new_n719_), .A2(G159), .ZN(new_n720_) );
  AND2_X1 g0584 ( .A1(G20), .A2(G179), .ZN(new_n721_) );
  AND3_X1 g0585 ( .A1(new_n721_), .A2(new_n716_), .A3(G200), .ZN(new_n722_) );
  AND2_X1 g0586 ( .A1(new_n722_), .A2(G68), .ZN(new_n723_) );
  AND3_X1 g0587 ( .A1(new_n387_), .A2(new_n337_), .A3(G190), .ZN(new_n724_) );
  OR2_X1 g0588 ( .A1(new_n724_), .A2(new_n175_), .ZN(new_n725_) );
  AND2_X1 g0589 ( .A1(new_n725_), .A2(G97), .ZN(new_n726_) );
  AND3_X1 g0590 ( .A1(new_n721_), .A2(new_n716_), .A3(new_n337_), .ZN(new_n727_) );
  AND2_X1 g0591 ( .A1(new_n727_), .A2(G77), .ZN(new_n728_) );
  OR4_X1 g0592 ( .A1(new_n720_), .A2(new_n723_), .A3(new_n726_), .A4(new_n728_), .ZN(new_n729_) );
  INV_X1 g0593 ( .A(new_n729_), .ZN(new_n730_) );
  AND2_X1 g0594 ( .A1(new_n730_), .A2(KEYINPUT61), .ZN(new_n731_) );
  OR2_X1 g0595 ( .A1(new_n730_), .A2(KEYINPUT61), .ZN(new_n732_) );
  INV_X1 g0596 ( .A(new_n732_), .ZN(new_n733_) );
  AND2_X1 g0597 ( .A1(new_n330_), .A2(G20), .ZN(new_n734_) );
  OR2_X1 g0598 ( .A1(new_n180_), .A2(new_n734_), .ZN(new_n735_) );
  INV_X1 g0599 ( .A(new_n735_), .ZN(new_n736_) );
  AND2_X1 g0600 ( .A1(new_n736_), .A2(new_n275_), .ZN(new_n737_) );
  INV_X1 g0601 ( .A(new_n737_), .ZN(new_n738_) );
  AND2_X1 g0602 ( .A1(new_n718_), .A2(G200), .ZN(new_n739_) );
  AND2_X1 g0603 ( .A1(new_n739_), .A2(G107), .ZN(new_n740_) );
  AND2_X1 g0604 ( .A1(G190), .A2(G200), .ZN(new_n741_) );
  AND2_X1 g0605 ( .A1(new_n721_), .A2(new_n741_), .ZN(new_n742_) );
  AND2_X1 g0606 ( .A1(new_n742_), .A2(G50), .ZN(new_n743_) );
  AND3_X1 g0607 ( .A1(new_n721_), .A2(G190), .A3(new_n337_), .ZN(new_n744_) );
  AND2_X1 g0608 ( .A1(new_n744_), .A2(G58), .ZN(new_n745_) );
  AND2_X1 g0609 ( .A1(new_n717_), .A2(new_n741_), .ZN(new_n746_) );
  AND2_X1 g0610 ( .A1(new_n746_), .A2(G87), .ZN(new_n747_) );
  OR4_X1 g0611 ( .A1(new_n740_), .A2(new_n743_), .A3(new_n745_), .A4(new_n747_), .ZN(new_n748_) );
  OR4_X1 g0612 ( .A1(new_n733_), .A2(new_n731_), .A3(new_n738_), .A4(new_n748_), .ZN(new_n749_) );
  INV_X1 g0613 ( .A(KEYINPUT24), .ZN(new_n750_) );
  AND2_X1 g0614 ( .A1(new_n184_), .A2(G33), .ZN(new_n751_) );
  AND2_X1 g0615 ( .A1(new_n751_), .A2(new_n750_), .ZN(new_n752_) );
  INV_X1 g0616 ( .A(new_n752_), .ZN(new_n753_) );
  OR2_X1 g0617 ( .A1(new_n751_), .A2(new_n750_), .ZN(new_n754_) );
  AND2_X1 g0618 ( .A1(new_n753_), .A2(new_n754_), .ZN(new_n755_) );
  INV_X1 g0619 ( .A(new_n755_), .ZN(new_n756_) );
  AND2_X1 g0620 ( .A1(new_n249_), .A2(G45), .ZN(new_n757_) );
  AND3_X1 g0621 ( .A1(new_n380_), .A2(new_n315_), .A3(G50), .ZN(new_n758_) );
  OR3_X1 g0622 ( .A1(new_n757_), .A2(new_n756_), .A3(new_n758_), .ZN(new_n759_) );
  INV_X1 g0623 ( .A(new_n184_), .ZN(new_n760_) );
  AND2_X1 g0624 ( .A1(new_n760_), .A2(new_n232_), .ZN(new_n761_) );
  AND2_X1 g0625 ( .A1(new_n761_), .A2(KEYINPUT60), .ZN(new_n762_) );
  INV_X1 g0626 ( .A(new_n762_), .ZN(new_n763_) );
  OR2_X1 g0627 ( .A1(new_n761_), .A2(KEYINPUT60), .ZN(new_n764_) );
  AND2_X1 g0628 ( .A1(G355), .A2(new_n710_), .ZN(new_n765_) );
  INV_X1 g0629 ( .A(new_n765_), .ZN(new_n766_) );
  AND4_X1 g0630 ( .A1(new_n759_), .A2(new_n763_), .A3(new_n764_), .A4(new_n766_), .ZN(new_n767_) );
  INV_X1 g0631 ( .A(new_n711_), .ZN(new_n768_) );
  AND2_X1 g0632 ( .A1(new_n735_), .A2(new_n768_), .ZN(new_n769_) );
  INV_X1 g0633 ( .A(new_n769_), .ZN(new_n770_) );
  OR2_X1 g0634 ( .A1(new_n767_), .A2(new_n770_), .ZN(new_n771_) );
  AND2_X1 g0635 ( .A1(new_n739_), .A2(G283), .ZN(new_n772_) );
  AND2_X1 g0636 ( .A1(new_n725_), .A2(G294), .ZN(new_n773_) );
  AND2_X1 g0637 ( .A1(new_n722_), .A2(G317), .ZN(new_n774_) );
  OR3_X1 g0638 ( .A1(new_n772_), .A2(new_n773_), .A3(new_n774_), .ZN(new_n775_) );
  AND2_X1 g0639 ( .A1(new_n736_), .A2(G33), .ZN(new_n776_) );
  INV_X1 g0640 ( .A(new_n776_), .ZN(new_n777_) );
  AND2_X1 g0641 ( .A1(new_n742_), .A2(G326), .ZN(new_n778_) );
  AND2_X1 g0642 ( .A1(new_n746_), .A2(G303), .ZN(new_n779_) );
  AND2_X1 g0643 ( .A1(new_n744_), .A2(G322), .ZN(new_n780_) );
  OR3_X1 g0644 ( .A1(new_n779_), .A2(new_n780_), .A3(new_n778_), .ZN(new_n781_) );
  AND2_X1 g0645 ( .A1(new_n719_), .A2(G329), .ZN(new_n782_) );
  AND2_X1 g0646 ( .A1(new_n727_), .A2(G311), .ZN(new_n783_) );
  OR2_X1 g0647 ( .A1(new_n782_), .A2(new_n783_), .ZN(new_n784_) );
  OR4_X1 g0648 ( .A1(new_n777_), .A2(new_n775_), .A3(new_n781_), .A4(new_n784_), .ZN(new_n785_) );
  INV_X1 g0649 ( .A(KEYINPUT1), .ZN(new_n786_) );
  AND3_X1 g0650 ( .A1(new_n175_), .A2(G13), .A3(G45), .ZN(new_n787_) );
  OR2_X1 g0651 ( .A1(new_n787_), .A2(new_n270_), .ZN(new_n788_) );
  AND2_X1 g0652 ( .A1(new_n788_), .A2(new_n786_), .ZN(new_n789_) );
  INV_X1 g0653 ( .A(new_n789_), .ZN(new_n790_) );
  OR2_X1 g0654 ( .A1(new_n788_), .A2(new_n786_), .ZN(new_n791_) );
  AND2_X1 g0655 ( .A1(new_n790_), .A2(new_n791_), .ZN(new_n792_) );
  AND2_X1 g0656 ( .A1(new_n792_), .A2(new_n705_), .ZN(new_n793_) );
  AND4_X1 g0657 ( .A1(new_n771_), .A2(new_n749_), .A3(new_n785_), .A4(new_n793_), .ZN(new_n794_) );
  AND3_X1 g0658 ( .A1(new_n714_), .A2(new_n715_), .A3(new_n794_), .ZN(new_n795_) );
  INV_X1 g0659 ( .A(new_n681_), .ZN(new_n796_) );
  INV_X1 g0660 ( .A(new_n793_), .ZN(new_n797_) );
  OR2_X1 g0661 ( .A1(new_n680_), .A2(G330), .ZN(new_n798_) );
  AND3_X1 g0662 ( .A1(new_n796_), .A2(new_n797_), .A3(new_n798_), .ZN(new_n799_) );
  OR2_X1 g0663 ( .A1(new_n795_), .A2(new_n799_), .ZN(G396) );
  INV_X1 g0664 ( .A(new_n701_), .ZN(new_n801_) );
  INV_X1 g0665 ( .A(KEYINPUT5), .ZN(new_n802_) );
  AND2_X1 g0666 ( .A1(new_n360_), .A2(new_n670_), .ZN(new_n803_) );
  INV_X1 g0667 ( .A(new_n803_), .ZN(new_n804_) );
  AND2_X1 g0668 ( .A1(new_n804_), .A2(new_n802_), .ZN(new_n805_) );
  AND2_X1 g0669 ( .A1(new_n803_), .A2(KEYINPUT5), .ZN(new_n806_) );
  OR2_X1 g0670 ( .A1(new_n805_), .A2(new_n806_), .ZN(new_n807_) );
  AND2_X1 g0671 ( .A1(new_n371_), .A2(new_n807_), .ZN(new_n808_) );
  INV_X1 g0672 ( .A(new_n805_), .ZN(new_n809_) );
  INV_X1 g0673 ( .A(new_n806_), .ZN(new_n810_) );
  AND3_X1 g0674 ( .A1(new_n809_), .A2(new_n368_), .A3(new_n810_), .ZN(new_n811_) );
  OR2_X1 g0675 ( .A1(new_n808_), .A2(new_n811_), .ZN(new_n812_) );
  INV_X1 g0676 ( .A(new_n812_), .ZN(new_n813_) );
  AND2_X1 g0677 ( .A1(new_n801_), .A2(new_n813_), .ZN(new_n814_) );
  AND2_X1 g0678 ( .A1(new_n701_), .A2(new_n812_), .ZN(new_n815_) );
  OR3_X1 g0679 ( .A1(new_n814_), .A2(new_n793_), .A3(new_n815_), .ZN(new_n816_) );
  AND2_X1 g0680 ( .A1(new_n813_), .A2(new_n710_), .ZN(new_n817_) );
  AND2_X1 g0681 ( .A1(new_n722_), .A2(G150), .ZN(new_n818_) );
  AND2_X1 g0682 ( .A1(new_n739_), .A2(G68), .ZN(new_n819_) );
  AND2_X1 g0683 ( .A1(new_n744_), .A2(G143), .ZN(new_n820_) );
  OR3_X1 g0684 ( .A1(new_n819_), .A2(new_n818_), .A3(new_n820_), .ZN(new_n821_) );
  INV_X1 g0685 ( .A(KEYINPUT19), .ZN(new_n822_) );
  AND2_X1 g0686 ( .A1(new_n719_), .A2(G132), .ZN(new_n823_) );
  OR2_X1 g0687 ( .A1(new_n823_), .A2(new_n822_), .ZN(new_n824_) );
  INV_X1 g0688 ( .A(new_n824_), .ZN(new_n825_) );
  AND2_X1 g0689 ( .A1(new_n823_), .A2(new_n822_), .ZN(new_n826_) );
  OR4_X1 g0690 ( .A1(new_n738_), .A2(new_n825_), .A3(new_n821_), .A4(new_n826_), .ZN(new_n827_) );
  INV_X1 g0691 ( .A(KEYINPUT20), .ZN(new_n828_) );
  AND2_X1 g0692 ( .A1(new_n725_), .A2(G58), .ZN(new_n829_) );
  AND2_X1 g0693 ( .A1(new_n727_), .A2(G159), .ZN(new_n830_) );
  AND2_X1 g0694 ( .A1(new_n746_), .A2(G50), .ZN(new_n831_) );
  AND2_X1 g0695 ( .A1(new_n742_), .A2(G137), .ZN(new_n832_) );
  OR3_X1 g0696 ( .A1(new_n831_), .A2(new_n830_), .A3(new_n832_), .ZN(new_n833_) );
  OR2_X1 g0697 ( .A1(new_n833_), .A2(new_n829_), .ZN(new_n834_) );
  INV_X1 g0698 ( .A(new_n834_), .ZN(new_n835_) );
  AND2_X1 g0699 ( .A1(new_n835_), .A2(new_n828_), .ZN(new_n836_) );
  AND2_X1 g0700 ( .A1(new_n834_), .A2(KEYINPUT20), .ZN(new_n837_) );
  OR3_X1 g0701 ( .A1(new_n827_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_) );
  INV_X1 g0702 ( .A(new_n838_), .ZN(new_n839_) );
  INV_X1 g0703 ( .A(KEYINPUT21), .ZN(new_n840_) );
  AND2_X1 g0704 ( .A1(new_n727_), .A2(G116), .ZN(new_n841_) );
  OR2_X1 g0705 ( .A1(new_n841_), .A2(new_n840_), .ZN(new_n842_) );
  AND2_X1 g0706 ( .A1(new_n841_), .A2(new_n840_), .ZN(new_n843_) );
  INV_X1 g0707 ( .A(new_n843_), .ZN(new_n844_) );
  AND2_X1 g0708 ( .A1(new_n744_), .A2(G294), .ZN(new_n845_) );
  INV_X1 g0709 ( .A(new_n845_), .ZN(new_n846_) );
  AND2_X1 g0710 ( .A1(new_n846_), .A2(G33), .ZN(new_n847_) );
  AND2_X1 g0711 ( .A1(new_n746_), .A2(G107), .ZN(new_n848_) );
  INV_X1 g0712 ( .A(new_n848_), .ZN(new_n849_) );
  AND2_X1 g0713 ( .A1(new_n742_), .A2(G303), .ZN(new_n850_) );
  INV_X1 g0714 ( .A(new_n850_), .ZN(new_n851_) );
  AND2_X1 g0715 ( .A1(new_n849_), .A2(new_n851_), .ZN(new_n852_) );
  AND4_X1 g0716 ( .A1(new_n852_), .A2(new_n842_), .A3(new_n844_), .A4(new_n847_), .ZN(new_n853_) );
  AND2_X1 g0717 ( .A1(new_n739_), .A2(G87), .ZN(new_n854_) );
  OR2_X1 g0718 ( .A1(new_n854_), .A2(KEYINPUT22), .ZN(new_n855_) );
  AND2_X1 g0719 ( .A1(new_n854_), .A2(KEYINPUT22), .ZN(new_n856_) );
  INV_X1 g0720 ( .A(new_n856_), .ZN(new_n857_) );
  AND2_X1 g0721 ( .A1(new_n857_), .A2(new_n855_), .ZN(new_n858_) );
  INV_X1 g0722 ( .A(new_n726_), .ZN(new_n859_) );
  AND2_X1 g0723 ( .A1(new_n736_), .A2(new_n859_), .ZN(new_n860_) );
  INV_X1 g0724 ( .A(G311), .ZN(new_n861_) );
  INV_X1 g0725 ( .A(new_n719_), .ZN(new_n862_) );
  OR2_X1 g0726 ( .A1(new_n862_), .A2(new_n861_), .ZN(new_n863_) );
  AND2_X1 g0727 ( .A1(new_n722_), .A2(G283), .ZN(new_n864_) );
  INV_X1 g0728 ( .A(new_n864_), .ZN(new_n865_) );
  AND2_X1 g0729 ( .A1(new_n863_), .A2(new_n865_), .ZN(new_n866_) );
  AND4_X1 g0730 ( .A1(new_n858_), .A2(new_n853_), .A3(new_n860_), .A4(new_n866_), .ZN(new_n867_) );
  INV_X1 g0731 ( .A(new_n710_), .ZN(new_n868_) );
  AND3_X1 g0732 ( .A1(new_n735_), .A2(new_n141_), .A3(new_n868_), .ZN(new_n869_) );
  OR4_X1 g0733 ( .A1(new_n839_), .A2(new_n797_), .A3(new_n867_), .A4(new_n869_), .ZN(new_n870_) );
  OR2_X1 g0734 ( .A1(new_n817_), .A2(new_n870_), .ZN(new_n871_) );
  AND2_X1 g0735 ( .A1(new_n816_), .A2(new_n871_), .ZN(new_n872_) );
  INV_X1 g0736 ( .A(new_n872_), .ZN(G384) );
  INV_X1 g0737 ( .A(new_n669_), .ZN(new_n874_) );
  AND2_X1 g0738 ( .A1(new_n652_), .A2(new_n874_), .ZN(new_n875_) );
  AND3_X1 g0739 ( .A1(new_n665_), .A2(new_n363_), .A3(new_n604_), .ZN(new_n876_) );
  OR2_X1 g0740 ( .A1(new_n876_), .A2(new_n369_), .ZN(new_n877_) );
  INV_X1 g0741 ( .A(KEYINPUT29), .ZN(new_n878_) );
  AND2_X1 g0742 ( .A1(new_n420_), .A2(new_n670_), .ZN(new_n879_) );
  INV_X1 g0743 ( .A(new_n879_), .ZN(new_n880_) );
  AND2_X1 g0744 ( .A1(new_n446_), .A2(new_n880_), .ZN(new_n881_) );
  AND2_X1 g0745 ( .A1(new_n653_), .A2(new_n670_), .ZN(new_n882_) );
  OR2_X1 g0746 ( .A1(new_n881_), .A2(new_n882_), .ZN(new_n883_) );
  AND2_X1 g0747 ( .A1(new_n883_), .A2(new_n878_), .ZN(new_n884_) );
  INV_X1 g0748 ( .A(new_n881_), .ZN(new_n885_) );
  INV_X1 g0749 ( .A(new_n882_), .ZN(new_n886_) );
  AND3_X1 g0750 ( .A1(new_n885_), .A2(KEYINPUT29), .A3(new_n886_), .ZN(new_n887_) );
  OR2_X1 g0751 ( .A1(new_n884_), .A2(new_n887_), .ZN(new_n888_) );
  AND3_X1 g0752 ( .A1(new_n877_), .A2(new_n683_), .A3(new_n888_), .ZN(new_n889_) );
  INV_X1 g0753 ( .A(new_n889_), .ZN(new_n890_) );
  AND2_X1 g0754 ( .A1(new_n653_), .A2(new_n683_), .ZN(new_n891_) );
  INV_X1 g0755 ( .A(new_n891_), .ZN(new_n892_) );
  AND2_X1 g0756 ( .A1(new_n890_), .A2(new_n892_), .ZN(new_n893_) );
  INV_X1 g0757 ( .A(new_n893_), .ZN(new_n894_) );
  INV_X1 g0758 ( .A(new_n875_), .ZN(new_n895_) );
  AND2_X1 g0759 ( .A1(new_n289_), .A2(new_n669_), .ZN(new_n896_) );
  INV_X1 g0760 ( .A(new_n896_), .ZN(new_n897_) );
  AND2_X1 g0761 ( .A1(new_n377_), .A2(new_n897_), .ZN(new_n898_) );
  OR2_X1 g0762 ( .A1(new_n898_), .A2(new_n652_), .ZN(new_n899_) );
  AND2_X1 g0763 ( .A1(new_n895_), .A2(new_n899_), .ZN(new_n900_) );
  AND2_X1 g0764 ( .A1(new_n894_), .A2(new_n900_), .ZN(new_n901_) );
  OR2_X1 g0765 ( .A1(new_n901_), .A2(new_n875_), .ZN(new_n902_) );
  INV_X1 g0766 ( .A(new_n902_), .ZN(new_n903_) );
  INV_X1 g0767 ( .A(new_n659_), .ZN(new_n904_) );
  AND3_X1 g0768 ( .A1(new_n666_), .A2(new_n448_), .A3(new_n683_), .ZN(new_n905_) );
  INV_X1 g0769 ( .A(new_n905_), .ZN(new_n906_) );
  AND2_X1 g0770 ( .A1(new_n906_), .A2(new_n904_), .ZN(new_n907_) );
  AND2_X1 g0771 ( .A1(new_n903_), .A2(new_n907_), .ZN(new_n908_) );
  INV_X1 g0772 ( .A(new_n907_), .ZN(new_n909_) );
  AND2_X1 g0773 ( .A1(new_n902_), .A2(new_n909_), .ZN(new_n910_) );
  OR2_X1 g0774 ( .A1(new_n908_), .A2(new_n910_), .ZN(new_n911_) );
  INV_X1 g0775 ( .A(new_n911_), .ZN(new_n912_) );
  AND2_X1 g0776 ( .A1(new_n888_), .A2(new_n812_), .ZN(new_n913_) );
  AND2_X1 g0777 ( .A1(new_n913_), .A2(new_n900_), .ZN(new_n914_) );
  AND2_X1 g0778 ( .A1(new_n914_), .A2(new_n448_), .ZN(new_n915_) );
  INV_X1 g0779 ( .A(new_n915_), .ZN(new_n916_) );
  OR2_X1 g0780 ( .A1(new_n914_), .A2(new_n448_), .ZN(new_n917_) );
  AND2_X1 g0781 ( .A1(new_n917_), .A2(new_n699_), .ZN(new_n918_) );
  AND2_X1 g0782 ( .A1(new_n918_), .A2(new_n916_), .ZN(new_n919_) );
  INV_X1 g0783 ( .A(new_n919_), .ZN(new_n920_) );
  AND2_X1 g0784 ( .A1(new_n912_), .A2(new_n920_), .ZN(new_n921_) );
  AND2_X1 g0785 ( .A1(new_n911_), .A2(new_n919_), .ZN(new_n922_) );
  OR2_X1 g0786 ( .A1(new_n921_), .A2(new_n922_), .ZN(new_n923_) );
  AND2_X1 g0787 ( .A1(new_n923_), .A2(new_n181_), .ZN(new_n924_) );
  AND2_X1 g0788 ( .A1(new_n183_), .A2(G1), .ZN(new_n925_) );
  OR2_X1 g0789 ( .A1(new_n924_), .A2(new_n925_), .ZN(new_n926_) );
  AND2_X1 g0790 ( .A1(G50), .A2(G58), .ZN(new_n927_) );
  AND2_X1 g0791 ( .A1(new_n927_), .A2(new_n138_), .ZN(new_n928_) );
  INV_X1 g0792 ( .A(new_n927_), .ZN(new_n929_) );
  AND2_X1 g0793 ( .A1(new_n929_), .A2(G68), .ZN(new_n930_) );
  OR2_X1 g0794 ( .A1(new_n930_), .A2(new_n928_), .ZN(new_n931_) );
  OR2_X1 g0795 ( .A1(new_n140_), .A2(G77), .ZN(new_n932_) );
  AND2_X1 g0796 ( .A1(new_n931_), .A2(new_n932_), .ZN(new_n933_) );
  OR3_X1 g0797 ( .A1(new_n933_), .A2(new_n270_), .A3(G13), .ZN(new_n934_) );
  AND2_X1 g0798 ( .A1(new_n926_), .A2(new_n934_), .ZN(new_n935_) );
  AND4_X1 g0799 ( .A1(new_n264_), .A2(G20), .A3(G116), .A4(new_n227_), .ZN(new_n936_) );
  OR2_X1 g0800 ( .A1(new_n935_), .A2(new_n936_), .ZN(G367) );
  OR2_X1 g0801 ( .A1(new_n662_), .A2(new_n564_), .ZN(new_n938_) );
  OR2_X1 g0802 ( .A1(new_n938_), .A2(new_n611_), .ZN(new_n939_) );
  INV_X1 g0803 ( .A(new_n611_), .ZN(new_n940_) );
  INV_X1 g0804 ( .A(new_n564_), .ZN(new_n941_) );
  INV_X1 g0805 ( .A(new_n523_), .ZN(new_n942_) );
  AND2_X1 g0806 ( .A1(new_n522_), .A2(new_n505_), .ZN(new_n943_) );
  OR2_X1 g0807 ( .A1(new_n943_), .A2(KEYINPUT0), .ZN(new_n944_) );
  AND2_X1 g0808 ( .A1(new_n944_), .A2(new_n942_), .ZN(new_n945_) );
  OR2_X1 g0809 ( .A1(new_n945_), .A2(new_n640_), .ZN(new_n946_) );
  AND2_X1 g0810 ( .A1(new_n946_), .A2(new_n505_), .ZN(new_n947_) );
  OR2_X1 g0811 ( .A1(new_n947_), .A2(new_n570_), .ZN(new_n948_) );
  AND2_X1 g0812 ( .A1(new_n948_), .A2(new_n941_), .ZN(new_n949_) );
  OR2_X1 g0813 ( .A1(new_n949_), .A2(new_n940_), .ZN(new_n950_) );
  AND3_X1 g0814 ( .A1(new_n950_), .A2(new_n939_), .A3(new_n683_), .ZN(new_n951_) );
  AND2_X1 g0815 ( .A1(new_n604_), .A2(new_n670_), .ZN(new_n952_) );
  OR2_X1 g0816 ( .A1(new_n951_), .A2(new_n952_), .ZN(new_n953_) );
  AND2_X1 g0817 ( .A1(new_n953_), .A2(KEYINPUT53), .ZN(new_n954_) );
  INV_X1 g0818 ( .A(KEYINPUT53), .ZN(new_n955_) );
  AND2_X1 g0819 ( .A1(new_n949_), .A2(new_n940_), .ZN(new_n956_) );
  AND2_X1 g0820 ( .A1(new_n938_), .A2(new_n611_), .ZN(new_n957_) );
  OR3_X1 g0821 ( .A1(new_n956_), .A2(new_n957_), .A3(new_n670_), .ZN(new_n958_) );
  INV_X1 g0822 ( .A(new_n952_), .ZN(new_n959_) );
  AND3_X1 g0823 ( .A1(new_n958_), .A2(new_n955_), .A3(new_n959_), .ZN(new_n960_) );
  AND3_X1 g0824 ( .A1(new_n585_), .A2(new_n609_), .A3(new_n670_), .ZN(new_n961_) );
  OR3_X1 g0825 ( .A1(new_n954_), .A2(new_n960_), .A3(new_n961_), .ZN(new_n962_) );
  AND2_X1 g0826 ( .A1(new_n563_), .A2(new_n670_), .ZN(new_n963_) );
  INV_X1 g0827 ( .A(new_n963_), .ZN(new_n964_) );
  AND2_X1 g0828 ( .A1(new_n571_), .A2(new_n964_), .ZN(new_n965_) );
  AND2_X1 g0829 ( .A1(new_n564_), .A2(new_n670_), .ZN(new_n966_) );
  OR2_X1 g0830 ( .A1(new_n965_), .A2(new_n966_), .ZN(new_n967_) );
  AND2_X1 g0831 ( .A1(new_n682_), .A2(new_n967_), .ZN(new_n968_) );
  AND2_X1 g0832 ( .A1(new_n962_), .A2(new_n968_), .ZN(new_n969_) );
  INV_X1 g0833 ( .A(new_n954_), .ZN(new_n970_) );
  INV_X1 g0834 ( .A(new_n960_), .ZN(new_n971_) );
  INV_X1 g0835 ( .A(new_n961_), .ZN(new_n972_) );
  AND3_X1 g0836 ( .A1(new_n970_), .A2(new_n971_), .A3(new_n972_), .ZN(new_n973_) );
  INV_X1 g0837 ( .A(new_n968_), .ZN(new_n974_) );
  AND2_X1 g0838 ( .A1(new_n973_), .A2(new_n974_), .ZN(new_n975_) );
  OR2_X1 g0839 ( .A1(new_n975_), .A2(new_n969_), .ZN(new_n976_) );
  INV_X1 g0840 ( .A(new_n682_), .ZN(new_n977_) );
  OR2_X1 g0841 ( .A1(new_n947_), .A2(new_n670_), .ZN(new_n978_) );
  AND2_X1 g0842 ( .A1(new_n978_), .A2(new_n964_), .ZN(new_n979_) );
  AND2_X1 g0843 ( .A1(new_n979_), .A2(new_n570_), .ZN(new_n980_) );
  OR2_X1 g0844 ( .A1(new_n684_), .A2(new_n963_), .ZN(new_n981_) );
  AND2_X1 g0845 ( .A1(new_n981_), .A2(new_n571_), .ZN(new_n982_) );
  OR2_X1 g0846 ( .A1(new_n980_), .A2(new_n982_), .ZN(new_n983_) );
  OR2_X1 g0847 ( .A1(new_n983_), .A2(new_n977_), .ZN(new_n984_) );
  OR2_X1 g0848 ( .A1(new_n981_), .A2(new_n571_), .ZN(new_n985_) );
  OR2_X1 g0849 ( .A1(new_n979_), .A2(new_n570_), .ZN(new_n986_) );
  AND2_X1 g0850 ( .A1(new_n986_), .A2(new_n985_), .ZN(new_n987_) );
  OR2_X1 g0851 ( .A1(new_n987_), .A2(new_n682_), .ZN(new_n988_) );
  AND2_X1 g0852 ( .A1(new_n646_), .A2(new_n683_), .ZN(new_n989_) );
  OR2_X1 g0853 ( .A1(new_n989_), .A2(new_n671_), .ZN(new_n990_) );
  AND2_X1 g0854 ( .A1(new_n533_), .A2(new_n990_), .ZN(new_n991_) );
  INV_X1 g0855 ( .A(new_n991_), .ZN(new_n992_) );
  OR2_X1 g0856 ( .A1(new_n533_), .A2(new_n990_), .ZN(new_n993_) );
  AND2_X1 g0857 ( .A1(new_n992_), .A2(new_n993_), .ZN(new_n994_) );
  AND2_X1 g0858 ( .A1(new_n796_), .A2(new_n994_), .ZN(new_n995_) );
  INV_X1 g0859 ( .A(new_n994_), .ZN(new_n996_) );
  AND2_X1 g0860 ( .A1(new_n681_), .A2(new_n996_), .ZN(new_n997_) );
  OR2_X1 g0861 ( .A1(new_n995_), .A2(new_n997_), .ZN(new_n998_) );
  AND3_X1 g0862 ( .A1(new_n984_), .A2(new_n988_), .A3(new_n998_), .ZN(new_n999_) );
  OR2_X1 g0863 ( .A1(new_n999_), .A2(KEYINPUT52), .ZN(new_n1000_) );
  INV_X1 g0864 ( .A(KEYINPUT52), .ZN(new_n1001_) );
  AND2_X1 g0865 ( .A1(new_n987_), .A2(new_n682_), .ZN(new_n1002_) );
  AND2_X1 g0866 ( .A1(new_n983_), .A2(new_n977_), .ZN(new_n1003_) );
  OR2_X1 g0867 ( .A1(new_n1003_), .A2(new_n1002_), .ZN(new_n1004_) );
  INV_X1 g0868 ( .A(new_n998_), .ZN(new_n1005_) );
  OR3_X1 g0869 ( .A1(new_n1004_), .A2(new_n1001_), .A3(new_n1005_), .ZN(new_n1006_) );
  AND2_X1 g0870 ( .A1(new_n801_), .A2(new_n792_), .ZN(new_n1007_) );
  AND3_X1 g0871 ( .A1(new_n1006_), .A2(new_n1000_), .A3(new_n1007_), .ZN(new_n1008_) );
  INV_X1 g0872 ( .A(new_n1008_), .ZN(new_n1009_) );
  AND3_X1 g0873 ( .A1(new_n976_), .A2(new_n797_), .A3(new_n1009_), .ZN(new_n1010_) );
  AND2_X1 g0874 ( .A1(new_n940_), .A2(new_n711_), .ZN(new_n1011_) );
  INV_X1 g0875 ( .A(new_n1011_), .ZN(new_n1012_) );
  AND2_X1 g0876 ( .A1(new_n719_), .A2(G317), .ZN(new_n1013_) );
  AND2_X1 g0877 ( .A1(new_n722_), .A2(G294), .ZN(new_n1014_) );
  AND2_X1 g0878 ( .A1(new_n739_), .A2(G97), .ZN(new_n1015_) );
  AND2_X1 g0879 ( .A1(new_n727_), .A2(G283), .ZN(new_n1016_) );
  OR4_X1 g0880 ( .A1(new_n1013_), .A2(new_n1015_), .A3(new_n1014_), .A4(new_n1016_), .ZN(new_n1017_) );
  INV_X1 g0881 ( .A(KEYINPUT54), .ZN(new_n1018_) );
  AND2_X1 g0882 ( .A1(new_n742_), .A2(G311), .ZN(new_n1019_) );
  AND2_X1 g0883 ( .A1(new_n1019_), .A2(new_n1018_), .ZN(new_n1020_) );
  INV_X1 g0884 ( .A(new_n1020_), .ZN(new_n1021_) );
  OR2_X1 g0885 ( .A1(new_n1019_), .A2(new_n1018_), .ZN(new_n1022_) );
  AND2_X1 g0886 ( .A1(new_n1021_), .A2(new_n1022_), .ZN(new_n1023_) );
  AND2_X1 g0887 ( .A1(new_n725_), .A2(G107), .ZN(new_n1024_) );
  AND2_X1 g0888 ( .A1(new_n744_), .A2(G303), .ZN(new_n1025_) );
  AND2_X1 g0889 ( .A1(new_n746_), .A2(G116), .ZN(new_n1026_) );
  OR3_X1 g0890 ( .A1(new_n1024_), .A2(new_n1025_), .A3(new_n1026_), .ZN(new_n1027_) );
  OR4_X1 g0891 ( .A1(new_n1017_), .A2(new_n777_), .A3(new_n1023_), .A4(new_n1027_), .ZN(new_n1028_) );
  AND2_X1 g0892 ( .A1(new_n727_), .A2(G50), .ZN(new_n1029_) );
  AND2_X1 g0893 ( .A1(new_n719_), .A2(G137), .ZN(new_n1030_) );
  AND2_X1 g0894 ( .A1(new_n722_), .A2(G159), .ZN(new_n1031_) );
  OR3_X1 g0895 ( .A1(new_n1030_), .A2(new_n1029_), .A3(new_n1031_), .ZN(new_n1032_) );
  AND2_X1 g0896 ( .A1(new_n742_), .A2(G143), .ZN(new_n1033_) );
  AND2_X1 g0897 ( .A1(new_n746_), .A2(G58), .ZN(new_n1034_) );
  AND2_X1 g0898 ( .A1(new_n744_), .A2(G150), .ZN(new_n1035_) );
  OR3_X1 g0899 ( .A1(new_n1034_), .A2(new_n1035_), .A3(new_n1033_), .ZN(new_n1036_) );
  AND2_X1 g0900 ( .A1(new_n739_), .A2(G77), .ZN(new_n1037_) );
  INV_X1 g0901 ( .A(new_n1037_), .ZN(new_n1038_) );
  AND2_X1 g0902 ( .A1(new_n725_), .A2(G68), .ZN(new_n1039_) );
  INV_X1 g0903 ( .A(new_n1039_), .ZN(new_n1040_) );
  AND2_X1 g0904 ( .A1(new_n1038_), .A2(new_n1040_), .ZN(new_n1041_) );
  INV_X1 g0905 ( .A(new_n1041_), .ZN(new_n1042_) );
  OR4_X1 g0906 ( .A1(new_n1042_), .A2(new_n738_), .A3(new_n1032_), .A4(new_n1036_), .ZN(new_n1043_) );
  AND2_X1 g0907 ( .A1(new_n220_), .A2(new_n755_), .ZN(new_n1044_) );
  AND2_X1 g0908 ( .A1(new_n760_), .A2(G87), .ZN(new_n1045_) );
  OR3_X1 g0909 ( .A1(new_n1044_), .A2(new_n770_), .A3(new_n1045_), .ZN(new_n1046_) );
  AND4_X1 g0910 ( .A1(new_n1046_), .A2(new_n793_), .A3(new_n1028_), .A4(new_n1043_), .ZN(new_n1047_) );
  AND2_X1 g0911 ( .A1(new_n1012_), .A2(new_n1047_), .ZN(new_n1048_) );
  OR3_X1 g0912 ( .A1(new_n1010_), .A2(KEYINPUT55), .A3(new_n1048_), .ZN(new_n1049_) );
  INV_X1 g0913 ( .A(KEYINPUT55), .ZN(new_n1050_) );
  OR2_X1 g0914 ( .A1(new_n973_), .A2(new_n974_), .ZN(new_n1051_) );
  OR2_X1 g0915 ( .A1(new_n962_), .A2(new_n968_), .ZN(new_n1052_) );
  AND2_X1 g0916 ( .A1(new_n1051_), .A2(new_n1052_), .ZN(new_n1053_) );
  OR2_X1 g0917 ( .A1(new_n1008_), .A2(new_n793_), .ZN(new_n1054_) );
  OR2_X1 g0918 ( .A1(new_n1053_), .A2(new_n1054_), .ZN(new_n1055_) );
  INV_X1 g0919 ( .A(new_n1048_), .ZN(new_n1056_) );
  AND2_X1 g0920 ( .A1(new_n1055_), .A2(new_n1056_), .ZN(new_n1057_) );
  OR2_X1 g0921 ( .A1(new_n1057_), .A2(new_n1050_), .ZN(new_n1058_) );
  AND2_X1 g0922 ( .A1(new_n1058_), .A2(new_n1049_), .ZN(G387) );
  INV_X1 g0923 ( .A(new_n1007_), .ZN(new_n1060_) );
  AND3_X1 g0924 ( .A1(new_n1060_), .A2(new_n797_), .A3(new_n998_), .ZN(new_n1061_) );
  AND3_X1 g0925 ( .A1(new_n801_), .A2(new_n704_), .A3(new_n1005_), .ZN(new_n1062_) );
  OR2_X1 g0926 ( .A1(new_n675_), .A2(new_n768_), .ZN(new_n1063_) );
  AND2_X1 g0927 ( .A1(new_n203_), .A2(G45), .ZN(new_n1064_) );
  INV_X1 g0928 ( .A(KEYINPUT23), .ZN(new_n1065_) );
  AND2_X1 g0929 ( .A1(G68), .A2(G77), .ZN(new_n1066_) );
  INV_X1 g0930 ( .A(new_n1066_), .ZN(new_n1067_) );
  AND4_X1 g0931 ( .A1(new_n703_), .A2(new_n140_), .A3(G58), .A4(new_n1067_), .ZN(new_n1068_) );
  OR2_X1 g0932 ( .A1(new_n1068_), .A2(G45), .ZN(new_n1069_) );
  AND2_X1 g0933 ( .A1(new_n1069_), .A2(new_n1065_), .ZN(new_n1070_) );
  INV_X1 g0934 ( .A(new_n1070_), .ZN(new_n1071_) );
  OR2_X1 g0935 ( .A1(new_n1069_), .A2(new_n1065_), .ZN(new_n1072_) );
  AND2_X1 g0936 ( .A1(new_n1071_), .A2(new_n1072_), .ZN(new_n1073_) );
  OR2_X1 g0937 ( .A1(new_n1064_), .A2(new_n1073_), .ZN(new_n1074_) );
  AND2_X1 g0938 ( .A1(new_n1074_), .A2(new_n755_), .ZN(new_n1075_) );
  OR2_X1 g0939 ( .A1(new_n703_), .A2(new_n868_), .ZN(new_n1076_) );
  INV_X1 g0940 ( .A(new_n1076_), .ZN(new_n1077_) );
  AND2_X1 g0941 ( .A1(new_n760_), .A2(new_n145_), .ZN(new_n1078_) );
  OR3_X1 g0942 ( .A1(new_n1075_), .A2(new_n1077_), .A3(new_n1078_), .ZN(new_n1079_) );
  AND2_X1 g0943 ( .A1(new_n1079_), .A2(new_n769_), .ZN(new_n1080_) );
  INV_X1 g0944 ( .A(new_n1080_), .ZN(new_n1081_) );
  AND2_X1 g0945 ( .A1(new_n725_), .A2(G87), .ZN(new_n1082_) );
  AND2_X1 g0946 ( .A1(new_n722_), .A2(G58), .ZN(new_n1083_) );
  AND2_X1 g0947 ( .A1(new_n727_), .A2(G68), .ZN(new_n1084_) );
  OR3_X1 g0948 ( .A1(new_n1082_), .A2(new_n1083_), .A3(new_n1084_), .ZN(new_n1085_) );
  AND2_X1 g0949 ( .A1(new_n744_), .A2(G50), .ZN(new_n1086_) );
  AND2_X1 g0950 ( .A1(new_n746_), .A2(G77), .ZN(new_n1087_) );
  AND2_X1 g0951 ( .A1(new_n742_), .A2(G159), .ZN(new_n1088_) );
  OR2_X1 g0952 ( .A1(new_n1087_), .A2(new_n1088_), .ZN(new_n1089_) );
  AND2_X1 g0953 ( .A1(new_n719_), .A2(G150), .ZN(new_n1090_) );
  OR4_X1 g0954 ( .A1(new_n1015_), .A2(new_n1089_), .A3(new_n1090_), .A4(new_n1086_), .ZN(new_n1091_) );
  OR3_X1 g0955 ( .A1(new_n1091_), .A2(new_n738_), .A3(new_n1085_), .ZN(new_n1092_) );
  INV_X1 g0956 ( .A(KEYINPUT25), .ZN(new_n1093_) );
  AND2_X1 g0957 ( .A1(new_n739_), .A2(G116), .ZN(new_n1094_) );
  AND2_X1 g0958 ( .A1(new_n1094_), .A2(new_n1093_), .ZN(new_n1095_) );
  OR2_X1 g0959 ( .A1(new_n1094_), .A2(new_n1093_), .ZN(new_n1096_) );
  INV_X1 g0960 ( .A(new_n1096_), .ZN(new_n1097_) );
  INV_X1 g0961 ( .A(KEYINPUT26), .ZN(new_n1098_) );
  AND2_X1 g0962 ( .A1(new_n746_), .A2(G294), .ZN(new_n1099_) );
  AND2_X1 g0963 ( .A1(new_n742_), .A2(G322), .ZN(new_n1100_) );
  OR2_X1 g0964 ( .A1(new_n1099_), .A2(new_n1100_), .ZN(new_n1101_) );
  INV_X1 g0965 ( .A(new_n1101_), .ZN(new_n1102_) );
  AND2_X1 g0966 ( .A1(new_n1102_), .A2(new_n1098_), .ZN(new_n1103_) );
  AND2_X1 g0967 ( .A1(new_n1101_), .A2(KEYINPUT26), .ZN(new_n1104_) );
  OR2_X1 g0968 ( .A1(new_n1103_), .A2(new_n1104_), .ZN(new_n1105_) );
  AND2_X1 g0969 ( .A1(new_n727_), .A2(G303), .ZN(new_n1106_) );
  AND2_X1 g0970 ( .A1(new_n725_), .A2(G283), .ZN(new_n1107_) );
  AND2_X1 g0971 ( .A1(new_n722_), .A2(G311), .ZN(new_n1108_) );
  OR3_X1 g0972 ( .A1(new_n1107_), .A2(new_n1106_), .A3(new_n1108_), .ZN(new_n1109_) );
  AND2_X1 g0973 ( .A1(new_n719_), .A2(G326), .ZN(new_n1110_) );
  AND2_X1 g0974 ( .A1(new_n744_), .A2(G317), .ZN(new_n1111_) );
  OR3_X1 g0975 ( .A1(new_n777_), .A2(new_n1110_), .A3(new_n1111_), .ZN(new_n1112_) );
  OR2_X1 g0976 ( .A1(new_n1112_), .A2(new_n1109_), .ZN(new_n1113_) );
  OR4_X1 g0977 ( .A1(new_n1113_), .A2(new_n1095_), .A3(new_n1097_), .A4(new_n1105_), .ZN(new_n1114_) );
  AND4_X1 g0978 ( .A1(new_n1081_), .A2(new_n793_), .A3(new_n1092_), .A4(new_n1114_), .ZN(new_n1115_) );
  AND2_X1 g0979 ( .A1(new_n1063_), .A2(new_n1115_), .ZN(new_n1116_) );
  OR3_X1 g0980 ( .A1(new_n1061_), .A2(new_n1062_), .A3(new_n1116_), .ZN(G393) );
  AND2_X1 g0981 ( .A1(new_n801_), .A2(new_n998_), .ZN(new_n1118_) );
  INV_X1 g0982 ( .A(new_n1118_), .ZN(new_n1119_) );
  AND2_X1 g0983 ( .A1(new_n1119_), .A2(new_n1004_), .ZN(new_n1120_) );
  INV_X1 g0984 ( .A(new_n1120_), .ZN(new_n1121_) );
  AND4_X1 g0985 ( .A1(new_n1121_), .A2(new_n704_), .A3(new_n1000_), .A4(new_n1006_), .ZN(new_n1122_) );
  INV_X1 g0986 ( .A(new_n1122_), .ZN(new_n1123_) );
  OR3_X1 g0987 ( .A1(new_n1007_), .A2(new_n1004_), .A3(new_n793_), .ZN(new_n1124_) );
  OR2_X1 g0988 ( .A1(new_n967_), .A2(new_n768_), .ZN(new_n1125_) );
  INV_X1 g0989 ( .A(KEYINPUT58), .ZN(new_n1126_) );
  AND2_X1 g0990 ( .A1(new_n744_), .A2(G311), .ZN(new_n1127_) );
  OR3_X1 g0991 ( .A1(new_n740_), .A2(new_n275_), .A3(new_n1127_), .ZN(new_n1128_) );
  AND2_X1 g0992 ( .A1(new_n719_), .A2(G322), .ZN(new_n1129_) );
  AND2_X1 g0993 ( .A1(new_n727_), .A2(G294), .ZN(new_n1130_) );
  OR2_X1 g0994 ( .A1(new_n1129_), .A2(new_n1130_), .ZN(new_n1131_) );
  AND2_X1 g0995 ( .A1(new_n725_), .A2(G116), .ZN(new_n1132_) );
  AND2_X1 g0996 ( .A1(new_n722_), .A2(G303), .ZN(new_n1133_) );
  OR4_X1 g0997 ( .A1(new_n1128_), .A2(new_n1131_), .A3(new_n1132_), .A4(new_n1133_), .ZN(new_n1134_) );
  INV_X1 g0998 ( .A(new_n1134_), .ZN(new_n1135_) );
  AND2_X1 g0999 ( .A1(new_n1135_), .A2(new_n1126_), .ZN(new_n1136_) );
  AND2_X1 g1000 ( .A1(new_n1134_), .A2(KEYINPUT58), .ZN(new_n1137_) );
  INV_X1 g1001 ( .A(KEYINPUT59), .ZN(new_n1138_) );
  AND2_X1 g1002 ( .A1(new_n746_), .A2(G283), .ZN(new_n1139_) );
  AND2_X1 g1003 ( .A1(new_n742_), .A2(G317), .ZN(new_n1140_) );
  OR2_X1 g1004 ( .A1(new_n1139_), .A2(new_n1140_), .ZN(new_n1141_) );
  INV_X1 g1005 ( .A(new_n1141_), .ZN(new_n1142_) );
  AND2_X1 g1006 ( .A1(new_n1142_), .A2(new_n1138_), .ZN(new_n1143_) );
  AND2_X1 g1007 ( .A1(new_n1141_), .A2(KEYINPUT59), .ZN(new_n1144_) );
  OR2_X1 g1008 ( .A1(new_n1143_), .A2(new_n1144_), .ZN(new_n1145_) );
  INV_X1 g1009 ( .A(new_n1145_), .ZN(new_n1146_) );
  OR3_X1 g1010 ( .A1(new_n1136_), .A2(new_n1137_), .A3(new_n1146_), .ZN(new_n1147_) );
  INV_X1 g1011 ( .A(KEYINPUT57), .ZN(new_n1148_) );
  AND2_X1 g1012 ( .A1(new_n742_), .A2(G150), .ZN(new_n1149_) );
  OR2_X1 g1013 ( .A1(new_n1149_), .A2(KEYINPUT56), .ZN(new_n1150_) );
  INV_X1 g1014 ( .A(new_n1150_), .ZN(new_n1151_) );
  AND2_X1 g1015 ( .A1(new_n746_), .A2(G68), .ZN(new_n1152_) );
  AND2_X1 g1016 ( .A1(new_n1149_), .A2(KEYINPUT56), .ZN(new_n1153_) );
  OR3_X1 g1017 ( .A1(new_n1151_), .A2(new_n1152_), .A3(new_n1153_), .ZN(new_n1154_) );
  INV_X1 g1018 ( .A(new_n1154_), .ZN(new_n1155_) );
  AND2_X1 g1019 ( .A1(new_n1155_), .A2(new_n1148_), .ZN(new_n1156_) );
  AND2_X1 g1020 ( .A1(new_n1154_), .A2(KEYINPUT57), .ZN(new_n1157_) );
  OR2_X1 g1021 ( .A1(new_n1156_), .A2(new_n1157_), .ZN(new_n1158_) );
  AND2_X1 g1022 ( .A1(new_n719_), .A2(G143), .ZN(new_n1159_) );
  AND2_X1 g1023 ( .A1(new_n744_), .A2(G159), .ZN(new_n1160_) );
  OR3_X1 g1024 ( .A1(new_n1159_), .A2(G33), .A3(new_n1160_), .ZN(new_n1161_) );
  INV_X1 g1025 ( .A(new_n1161_), .ZN(new_n1162_) );
  AND2_X1 g1026 ( .A1(new_n725_), .A2(G77), .ZN(new_n1163_) );
  AND2_X1 g1027 ( .A1(new_n722_), .A2(G50), .ZN(new_n1164_) );
  AND2_X1 g1028 ( .A1(new_n727_), .A2(G58), .ZN(new_n1165_) );
  OR3_X1 g1029 ( .A1(new_n1163_), .A2(new_n1164_), .A3(new_n1165_), .ZN(new_n1166_) );
  INV_X1 g1030 ( .A(new_n1166_), .ZN(new_n1167_) );
  AND4_X1 g1031 ( .A1(new_n1158_), .A2(new_n858_), .A3(new_n1162_), .A4(new_n1167_), .ZN(new_n1168_) );
  INV_X1 g1032 ( .A(new_n1168_), .ZN(new_n1169_) );
  AND2_X1 g1033 ( .A1(new_n1147_), .A2(new_n1169_), .ZN(new_n1170_) );
  OR2_X1 g1034 ( .A1(new_n1170_), .A2(new_n735_), .ZN(new_n1171_) );
  AND2_X1 g1035 ( .A1(new_n239_), .A2(new_n755_), .ZN(new_n1172_) );
  AND2_X1 g1036 ( .A1(new_n760_), .A2(G97), .ZN(new_n1173_) );
  OR3_X1 g1037 ( .A1(new_n1172_), .A2(new_n770_), .A3(new_n1173_), .ZN(new_n1174_) );
  AND4_X1 g1038 ( .A1(new_n1125_), .A2(new_n793_), .A3(new_n1171_), .A4(new_n1174_), .ZN(new_n1175_) );
  INV_X1 g1039 ( .A(new_n1175_), .ZN(new_n1176_) );
  AND2_X1 g1040 ( .A1(new_n1124_), .A2(new_n1176_), .ZN(new_n1177_) );
  AND2_X1 g1041 ( .A1(new_n1123_), .A2(new_n1177_), .ZN(new_n1178_) );
  INV_X1 g1042 ( .A(new_n1178_), .ZN(G390) );
  INV_X1 g1043 ( .A(KEYINPUT39), .ZN(new_n1180_) );
  AND3_X1 g1044 ( .A1(new_n913_), .A2(new_n698_), .A3(G330), .ZN(new_n1181_) );
  AND2_X1 g1045 ( .A1(new_n1181_), .A2(new_n1180_), .ZN(new_n1182_) );
  OR2_X1 g1046 ( .A1(new_n1181_), .A2(new_n1180_), .ZN(new_n1183_) );
  INV_X1 g1047 ( .A(new_n1183_), .ZN(new_n1184_) );
  OR2_X1 g1048 ( .A1(new_n1184_), .A2(new_n1182_), .ZN(new_n1185_) );
  OR3_X1 g1049 ( .A1(new_n1185_), .A2(new_n889_), .A3(new_n891_), .ZN(new_n1186_) );
  INV_X1 g1050 ( .A(KEYINPUT40), .ZN(new_n1187_) );
  AND2_X1 g1051 ( .A1(new_n900_), .A2(new_n1187_), .ZN(new_n1188_) );
  INV_X1 g1052 ( .A(new_n900_), .ZN(new_n1189_) );
  AND2_X1 g1053 ( .A1(new_n1189_), .A2(KEYINPUT40), .ZN(new_n1190_) );
  OR2_X1 g1054 ( .A1(new_n1190_), .A2(new_n1188_), .ZN(new_n1191_) );
  AND2_X1 g1055 ( .A1(new_n1186_), .A2(new_n1191_), .ZN(new_n1192_) );
  INV_X1 g1056 ( .A(new_n1182_), .ZN(new_n1193_) );
  AND2_X1 g1057 ( .A1(new_n1193_), .A2(new_n1183_), .ZN(new_n1194_) );
  AND3_X1 g1058 ( .A1(new_n890_), .A2(new_n892_), .A3(new_n1194_), .ZN(new_n1195_) );
  INV_X1 g1059 ( .A(new_n1191_), .ZN(new_n1196_) );
  AND2_X1 g1060 ( .A1(new_n1195_), .A2(new_n1196_), .ZN(new_n1197_) );
  OR2_X1 g1061 ( .A1(new_n1197_), .A2(new_n1192_), .ZN(new_n1198_) );
  INV_X1 g1062 ( .A(KEYINPUT38), .ZN(new_n1199_) );
  AND2_X1 g1063 ( .A1(new_n699_), .A2(new_n448_), .ZN(new_n1200_) );
  OR3_X1 g1064 ( .A1(new_n905_), .A2(new_n659_), .A3(new_n1200_), .ZN(new_n1201_) );
  AND2_X1 g1065 ( .A1(new_n1201_), .A2(new_n1199_), .ZN(new_n1202_) );
  INV_X1 g1066 ( .A(new_n1201_), .ZN(new_n1203_) );
  AND2_X1 g1067 ( .A1(new_n1203_), .A2(KEYINPUT38), .ZN(new_n1204_) );
  OR2_X1 g1068 ( .A1(new_n1204_), .A2(new_n1202_), .ZN(new_n1205_) );
  AND2_X1 g1069 ( .A1(new_n877_), .A2(new_n683_), .ZN(new_n1206_) );
  INV_X1 g1070 ( .A(new_n1206_), .ZN(new_n1207_) );
  INV_X1 g1071 ( .A(new_n888_), .ZN(new_n1208_) );
  AND2_X1 g1072 ( .A1(new_n699_), .A2(new_n812_), .ZN(new_n1209_) );
  INV_X1 g1073 ( .A(new_n1209_), .ZN(new_n1210_) );
  AND3_X1 g1074 ( .A1(new_n1207_), .A2(new_n1208_), .A3(new_n1210_), .ZN(new_n1211_) );
  INV_X1 g1075 ( .A(new_n1211_), .ZN(new_n1212_) );
  OR2_X1 g1076 ( .A1(new_n1206_), .A2(new_n1209_), .ZN(new_n1213_) );
  AND2_X1 g1077 ( .A1(new_n1213_), .A2(new_n888_), .ZN(new_n1214_) );
  INV_X1 g1078 ( .A(new_n1214_), .ZN(new_n1215_) );
  AND3_X1 g1079 ( .A1(new_n1205_), .A2(new_n1212_), .A3(new_n1215_), .ZN(new_n1216_) );
  AND2_X1 g1080 ( .A1(new_n1216_), .A2(new_n1198_), .ZN(new_n1217_) );
  INV_X1 g1081 ( .A(new_n1217_), .ZN(new_n1218_) );
  OR2_X1 g1082 ( .A1(new_n1216_), .A2(new_n1198_), .ZN(new_n1219_) );
  AND3_X1 g1083 ( .A1(new_n1218_), .A2(new_n704_), .A3(new_n1219_), .ZN(new_n1220_) );
  INV_X1 g1084 ( .A(new_n792_), .ZN(new_n1221_) );
  AND2_X1 g1085 ( .A1(new_n1198_), .A2(new_n1221_), .ZN(new_n1222_) );
  AND2_X1 g1086 ( .A1(new_n1189_), .A2(new_n710_), .ZN(new_n1223_) );
  AND2_X1 g1087 ( .A1(new_n725_), .A2(G159), .ZN(new_n1224_) );
  AND2_X1 g1088 ( .A1(new_n739_), .A2(G50), .ZN(new_n1225_) );
  AND2_X1 g1089 ( .A1(new_n727_), .A2(G143), .ZN(new_n1226_) );
  OR3_X1 g1090 ( .A1(new_n1225_), .A2(new_n1224_), .A3(new_n1226_), .ZN(new_n1227_) );
  AND2_X1 g1091 ( .A1(new_n742_), .A2(G128), .ZN(new_n1228_) );
  AND2_X1 g1092 ( .A1(new_n746_), .A2(G150), .ZN(new_n1229_) );
  AND2_X1 g1093 ( .A1(new_n744_), .A2(G132), .ZN(new_n1230_) );
  OR3_X1 g1094 ( .A1(new_n1229_), .A2(new_n1230_), .A3(new_n1228_), .ZN(new_n1231_) );
  AND2_X1 g1095 ( .A1(new_n719_), .A2(G125), .ZN(new_n1232_) );
  AND2_X1 g1096 ( .A1(new_n722_), .A2(G137), .ZN(new_n1233_) );
  OR2_X1 g1097 ( .A1(new_n1232_), .A2(new_n1233_), .ZN(new_n1234_) );
  OR4_X1 g1098 ( .A1(new_n738_), .A2(new_n1227_), .A3(new_n1231_), .A4(new_n1234_), .ZN(new_n1235_) );
  INV_X1 g1099 ( .A(new_n1235_), .ZN(new_n1236_) );
  INV_X1 g1100 ( .A(KEYINPUT48), .ZN(new_n1237_) );
  AND2_X1 g1101 ( .A1(new_n719_), .A2(G294), .ZN(new_n1238_) );
  AND2_X1 g1102 ( .A1(new_n727_), .A2(G97), .ZN(new_n1239_) );
  OR2_X1 g1103 ( .A1(new_n1238_), .A2(new_n1239_), .ZN(new_n1240_) );
  AND2_X1 g1104 ( .A1(new_n1240_), .A2(new_n1237_), .ZN(new_n1241_) );
  INV_X1 g1105 ( .A(new_n1240_), .ZN(new_n1242_) );
  AND2_X1 g1106 ( .A1(new_n1242_), .A2(KEYINPUT48), .ZN(new_n1243_) );
  OR2_X1 g1107 ( .A1(new_n1243_), .A2(new_n1241_), .ZN(new_n1244_) );
  INV_X1 g1108 ( .A(new_n819_), .ZN(new_n1245_) );
  INV_X1 g1109 ( .A(new_n1163_), .ZN(new_n1246_) );
  INV_X1 g1110 ( .A(new_n747_), .ZN(new_n1247_) );
  AND2_X1 g1111 ( .A1(new_n742_), .A2(G283), .ZN(new_n1248_) );
  INV_X1 g1112 ( .A(new_n1248_), .ZN(new_n1249_) );
  AND2_X1 g1113 ( .A1(new_n1247_), .A2(new_n1249_), .ZN(new_n1250_) );
  AND2_X1 g1114 ( .A1(new_n722_), .A2(G107), .ZN(new_n1251_) );
  INV_X1 g1115 ( .A(new_n1251_), .ZN(new_n1252_) );
  AND4_X1 g1116 ( .A1(new_n1245_), .A2(new_n1250_), .A3(new_n1246_), .A4(new_n1252_), .ZN(new_n1253_) );
  INV_X1 g1117 ( .A(KEYINPUT47), .ZN(new_n1254_) );
  AND2_X1 g1118 ( .A1(new_n744_), .A2(G116), .ZN(new_n1255_) );
  INV_X1 g1119 ( .A(new_n1255_), .ZN(new_n1256_) );
  AND2_X1 g1120 ( .A1(new_n1256_), .A2(new_n1254_), .ZN(new_n1257_) );
  AND2_X1 g1121 ( .A1(new_n1255_), .A2(KEYINPUT47), .ZN(new_n1258_) );
  OR2_X1 g1122 ( .A1(new_n1257_), .A2(new_n1258_), .ZN(new_n1259_) );
  AND4_X1 g1123 ( .A1(new_n1244_), .A2(new_n776_), .A3(new_n1253_), .A4(new_n1259_), .ZN(new_n1260_) );
  AND3_X1 g1124 ( .A1(new_n735_), .A2(new_n137_), .A3(new_n868_), .ZN(new_n1261_) );
  OR4_X1 g1125 ( .A1(new_n1260_), .A2(new_n797_), .A3(new_n1236_), .A4(new_n1261_), .ZN(new_n1262_) );
  OR2_X1 g1126 ( .A1(new_n1223_), .A2(new_n1262_), .ZN(new_n1263_) );
  INV_X1 g1127 ( .A(new_n1263_), .ZN(new_n1264_) );
  OR3_X1 g1128 ( .A1(new_n1220_), .A2(new_n1222_), .A3(new_n1264_), .ZN(G378) );
  AND2_X1 g1129 ( .A1(new_n1215_), .A2(new_n1212_), .ZN(new_n1266_) );
  AND2_X1 g1130 ( .A1(new_n1198_), .A2(new_n1266_), .ZN(new_n1267_) );
  AND2_X1 g1131 ( .A1(new_n1267_), .A2(KEYINPUT41), .ZN(new_n1268_) );
  INV_X1 g1132 ( .A(KEYINPUT41), .ZN(new_n1269_) );
  OR2_X1 g1133 ( .A1(new_n1195_), .A2(new_n1196_), .ZN(new_n1270_) );
  OR2_X1 g1134 ( .A1(new_n1186_), .A2(new_n1191_), .ZN(new_n1271_) );
  AND2_X1 g1135 ( .A1(new_n1270_), .A2(new_n1271_), .ZN(new_n1272_) );
  OR2_X1 g1136 ( .A1(new_n1214_), .A2(new_n1211_), .ZN(new_n1273_) );
  OR2_X1 g1137 ( .A1(new_n1272_), .A2(new_n1273_), .ZN(new_n1274_) );
  AND2_X1 g1138 ( .A1(new_n1274_), .A2(new_n1269_), .ZN(new_n1275_) );
  OR2_X1 g1139 ( .A1(new_n1275_), .A2(new_n1268_), .ZN(new_n1276_) );
  AND2_X1 g1140 ( .A1(new_n1205_), .A2(new_n792_), .ZN(new_n1277_) );
  AND2_X1 g1141 ( .A1(new_n1276_), .A2(new_n1277_), .ZN(new_n1278_) );
  AND2_X1 g1142 ( .A1(new_n914_), .A2(new_n699_), .ZN(new_n1279_) );
  INV_X1 g1143 ( .A(new_n1279_), .ZN(new_n1280_) );
  AND2_X1 g1144 ( .A1(new_n386_), .A2(new_n669_), .ZN(new_n1281_) );
  INV_X1 g1145 ( .A(new_n1281_), .ZN(new_n1282_) );
  AND2_X1 g1146 ( .A1(new_n413_), .A2(new_n1282_), .ZN(new_n1283_) );
  AND2_X1 g1147 ( .A1(new_n404_), .A2(new_n669_), .ZN(new_n1284_) );
  OR2_X1 g1148 ( .A1(new_n1283_), .A2(new_n1284_), .ZN(new_n1285_) );
  INV_X1 g1149 ( .A(new_n1285_), .ZN(new_n1286_) );
  AND3_X1 g1150 ( .A1(new_n903_), .A2(new_n1280_), .A3(new_n1286_), .ZN(new_n1287_) );
  OR2_X1 g1151 ( .A1(new_n902_), .A2(new_n1279_), .ZN(new_n1288_) );
  AND2_X1 g1152 ( .A1(new_n1288_), .A2(new_n1285_), .ZN(new_n1289_) );
  OR3_X1 g1153 ( .A1(new_n1289_), .A2(new_n793_), .A3(new_n1287_), .ZN(new_n1290_) );
  OR2_X1 g1154 ( .A1(new_n1278_), .A2(new_n1290_), .ZN(new_n1291_) );
  AND2_X1 g1155 ( .A1(new_n1286_), .A2(new_n710_), .ZN(new_n1292_) );
  AND2_X1 g1156 ( .A1(new_n739_), .A2(G159), .ZN(new_n1293_) );
  AND2_X1 g1157 ( .A1(new_n722_), .A2(G132), .ZN(new_n1294_) );
  OR2_X1 g1158 ( .A1(new_n1293_), .A2(new_n1294_), .ZN(new_n1295_) );
  OR2_X1 g1159 ( .A1(new_n1295_), .A2(KEYINPUT44), .ZN(new_n1296_) );
  AND2_X1 g1160 ( .A1(new_n744_), .A2(G128), .ZN(new_n1297_) );
  INV_X1 g1161 ( .A(new_n1297_), .ZN(new_n1298_) );
  AND2_X1 g1162 ( .A1(new_n746_), .A2(G143), .ZN(new_n1299_) );
  INV_X1 g1163 ( .A(new_n1299_), .ZN(new_n1300_) );
  AND2_X1 g1164 ( .A1(new_n742_), .A2(G125), .ZN(new_n1301_) );
  INV_X1 g1165 ( .A(new_n1301_), .ZN(new_n1302_) );
  AND3_X1 g1166 ( .A1(new_n1300_), .A2(new_n1298_), .A3(new_n1302_), .ZN(new_n1303_) );
  INV_X1 g1167 ( .A(G124), .ZN(new_n1304_) );
  OR2_X1 g1168 ( .A1(new_n862_), .A2(new_n1304_), .ZN(new_n1305_) );
  INV_X1 g1169 ( .A(G150), .ZN(new_n1306_) );
  INV_X1 g1170 ( .A(new_n725_), .ZN(new_n1307_) );
  OR2_X1 g1171 ( .A1(new_n1307_), .A2(new_n1306_), .ZN(new_n1308_) );
  AND3_X1 g1172 ( .A1(new_n1303_), .A2(new_n1305_), .A3(new_n1308_), .ZN(new_n1309_) );
  INV_X1 g1173 ( .A(KEYINPUT44), .ZN(new_n1310_) );
  INV_X1 g1174 ( .A(new_n1295_), .ZN(new_n1311_) );
  OR2_X1 g1175 ( .A1(new_n1311_), .A2(new_n1310_), .ZN(new_n1312_) );
  INV_X1 g1176 ( .A(KEYINPUT43), .ZN(new_n1313_) );
  AND2_X1 g1177 ( .A1(new_n727_), .A2(G137), .ZN(new_n1314_) );
  INV_X1 g1178 ( .A(new_n1314_), .ZN(new_n1315_) );
  AND2_X1 g1179 ( .A1(new_n1315_), .A2(new_n1313_), .ZN(new_n1316_) );
  AND2_X1 g1180 ( .A1(new_n1314_), .A2(KEYINPUT43), .ZN(new_n1317_) );
  OR2_X1 g1181 ( .A1(new_n1316_), .A2(new_n1317_), .ZN(new_n1318_) );
  AND4_X1 g1182 ( .A1(new_n1312_), .A2(new_n1296_), .A3(new_n1309_), .A4(new_n1318_), .ZN(new_n1319_) );
  OR2_X1 g1183 ( .A1(new_n1319_), .A2(G33), .ZN(new_n1320_) );
  AND2_X1 g1184 ( .A1(new_n744_), .A2(G107), .ZN(new_n1321_) );
  AND2_X1 g1185 ( .A1(new_n1321_), .A2(KEYINPUT42), .ZN(new_n1322_) );
  INV_X1 g1186 ( .A(new_n1322_), .ZN(new_n1323_) );
  AND2_X1 g1187 ( .A1(new_n727_), .A2(G87), .ZN(new_n1324_) );
  INV_X1 g1188 ( .A(new_n1324_), .ZN(new_n1325_) );
  OR2_X1 g1189 ( .A1(new_n862_), .A2(new_n538_), .ZN(new_n1326_) );
  AND2_X1 g1190 ( .A1(new_n722_), .A2(G97), .ZN(new_n1327_) );
  INV_X1 g1191 ( .A(new_n1327_), .ZN(new_n1328_) );
  AND4_X1 g1192 ( .A1(new_n1326_), .A2(new_n1323_), .A3(new_n1325_), .A4(new_n1328_), .ZN(new_n1329_) );
  INV_X1 g1193 ( .A(new_n1087_), .ZN(new_n1330_) );
  AND2_X1 g1194 ( .A1(new_n742_), .A2(G116), .ZN(new_n1331_) );
  INV_X1 g1195 ( .A(new_n1331_), .ZN(new_n1332_) );
  AND3_X1 g1196 ( .A1(new_n1040_), .A2(new_n1330_), .A3(new_n1332_), .ZN(new_n1333_) );
  OR2_X1 g1197 ( .A1(new_n1321_), .A2(KEYINPUT42), .ZN(new_n1334_) );
  AND2_X1 g1198 ( .A1(new_n739_), .A2(G58), .ZN(new_n1335_) );
  INV_X1 g1199 ( .A(new_n1335_), .ZN(new_n1336_) );
  AND4_X1 g1200 ( .A1(new_n1329_), .A2(new_n1333_), .A3(new_n1334_), .A4(new_n1336_), .ZN(new_n1337_) );
  OR2_X1 g1201 ( .A1(new_n1337_), .A2(new_n275_), .ZN(new_n1338_) );
  AND2_X1 g1202 ( .A1(new_n736_), .A2(new_n314_), .ZN(new_n1339_) );
  AND3_X1 g1203 ( .A1(new_n1320_), .A2(new_n1338_), .A3(new_n1339_), .ZN(new_n1340_) );
  OR3_X1 g1204 ( .A1(new_n1339_), .A2(G50), .A3(new_n710_), .ZN(new_n1341_) );
  INV_X1 g1205 ( .A(new_n1341_), .ZN(new_n1342_) );
  OR4_X1 g1206 ( .A1(new_n1292_), .A2(new_n797_), .A3(new_n1340_), .A4(new_n1342_), .ZN(new_n1343_) );
  AND2_X1 g1207 ( .A1(new_n1291_), .A2(new_n1343_), .ZN(new_n1344_) );
  INV_X1 g1208 ( .A(new_n1344_), .ZN(G375) );
  INV_X1 g1209 ( .A(new_n1216_), .ZN(new_n1346_) );
  INV_X1 g1210 ( .A(new_n1202_), .ZN(new_n1347_) );
  OR2_X1 g1211 ( .A1(new_n1201_), .A2(new_n1199_), .ZN(new_n1348_) );
  AND2_X1 g1212 ( .A1(new_n1347_), .A2(new_n1348_), .ZN(new_n1349_) );
  AND2_X1 g1213 ( .A1(new_n1273_), .A2(new_n1349_), .ZN(new_n1350_) );
  INV_X1 g1214 ( .A(new_n1350_), .ZN(new_n1351_) );
  AND3_X1 g1215 ( .A1(new_n1351_), .A2(KEYINPUT46), .A3(new_n1346_), .ZN(new_n1352_) );
  INV_X1 g1216 ( .A(KEYINPUT46), .ZN(new_n1353_) );
  OR2_X1 g1217 ( .A1(new_n1350_), .A2(new_n1216_), .ZN(new_n1354_) );
  AND2_X1 g1218 ( .A1(new_n1354_), .A2(new_n1353_), .ZN(new_n1355_) );
  OR2_X1 g1219 ( .A1(new_n1355_), .A2(new_n1352_), .ZN(new_n1356_) );
  AND2_X1 g1220 ( .A1(new_n1356_), .A2(new_n704_), .ZN(new_n1357_) );
  AND2_X1 g1221 ( .A1(new_n1266_), .A2(new_n1221_), .ZN(new_n1358_) );
  INV_X1 g1222 ( .A(new_n1358_), .ZN(new_n1359_) );
  AND2_X1 g1223 ( .A1(new_n1208_), .A2(new_n710_), .ZN(new_n1360_) );
  INV_X1 g1224 ( .A(KEYINPUT45), .ZN(new_n1361_) );
  AND2_X1 g1225 ( .A1(new_n725_), .A2(G50), .ZN(new_n1362_) );
  AND2_X1 g1226 ( .A1(new_n727_), .A2(G150), .ZN(new_n1363_) );
  AND2_X1 g1227 ( .A1(new_n722_), .A2(G143), .ZN(new_n1364_) );
  OR3_X1 g1228 ( .A1(new_n1362_), .A2(new_n1363_), .A3(new_n1364_), .ZN(new_n1365_) );
  AND2_X1 g1229 ( .A1(new_n746_), .A2(G159), .ZN(new_n1366_) );
  AND2_X1 g1230 ( .A1(new_n744_), .A2(G137), .ZN(new_n1367_) );
  AND2_X1 g1231 ( .A1(new_n742_), .A2(G132), .ZN(new_n1368_) );
  OR2_X1 g1232 ( .A1(new_n1367_), .A2(new_n1368_), .ZN(new_n1369_) );
  AND2_X1 g1233 ( .A1(new_n719_), .A2(G128), .ZN(new_n1370_) );
  OR4_X1 g1234 ( .A1(new_n1335_), .A2(new_n1370_), .A3(new_n1369_), .A4(new_n1366_), .ZN(new_n1371_) );
  OR3_X1 g1235 ( .A1(new_n1371_), .A2(new_n738_), .A3(new_n1365_), .ZN(new_n1372_) );
  AND2_X1 g1236 ( .A1(new_n727_), .A2(G107), .ZN(new_n1373_) );
  AND2_X1 g1237 ( .A1(new_n719_), .A2(G303), .ZN(new_n1374_) );
  AND2_X1 g1238 ( .A1(new_n722_), .A2(G116), .ZN(new_n1375_) );
  OR3_X1 g1239 ( .A1(new_n1374_), .A2(new_n1373_), .A3(new_n1375_), .ZN(new_n1376_) );
  AND2_X1 g1240 ( .A1(new_n744_), .A2(G283), .ZN(new_n1377_) );
  AND2_X1 g1241 ( .A1(new_n746_), .A2(G97), .ZN(new_n1378_) );
  AND2_X1 g1242 ( .A1(new_n742_), .A2(G294), .ZN(new_n1379_) );
  OR3_X1 g1243 ( .A1(new_n1378_), .A2(new_n1377_), .A3(new_n1379_), .ZN(new_n1380_) );
  OR2_X1 g1244 ( .A1(new_n1037_), .A2(new_n1082_), .ZN(new_n1381_) );
  OR4_X1 g1245 ( .A1(new_n777_), .A2(new_n1376_), .A3(new_n1380_), .A4(new_n1381_), .ZN(new_n1382_) );
  AND3_X1 g1246 ( .A1(new_n735_), .A2(new_n138_), .A3(new_n868_), .ZN(new_n1383_) );
  INV_X1 g1247 ( .A(new_n1383_), .ZN(new_n1384_) );
  AND4_X1 g1248 ( .A1(new_n1382_), .A2(new_n1372_), .A3(new_n793_), .A4(new_n1384_), .ZN(new_n1385_) );
  AND2_X1 g1249 ( .A1(new_n1385_), .A2(new_n1361_), .ZN(new_n1386_) );
  INV_X1 g1250 ( .A(new_n1386_), .ZN(new_n1387_) );
  OR2_X1 g1251 ( .A1(new_n1385_), .A2(new_n1361_), .ZN(new_n1388_) );
  AND2_X1 g1252 ( .A1(new_n1387_), .A2(new_n1388_), .ZN(new_n1389_) );
  OR2_X1 g1253 ( .A1(new_n1360_), .A2(new_n1389_), .ZN(new_n1390_) );
  AND2_X1 g1254 ( .A1(new_n1359_), .A2(new_n1390_), .ZN(new_n1391_) );
  INV_X1 g1255 ( .A(new_n1391_), .ZN(new_n1392_) );
  OR2_X1 g1256 ( .A1(new_n1357_), .A2(new_n1392_), .ZN(G381) );
  INV_X1 g1257 ( .A(new_n1049_), .ZN(new_n1394_) );
  OR2_X1 g1258 ( .A1(new_n1010_), .A2(new_n1048_), .ZN(new_n1395_) );
  AND2_X1 g1259 ( .A1(new_n1395_), .A2(KEYINPUT55), .ZN(new_n1396_) );
  OR2_X1 g1260 ( .A1(new_n1396_), .A2(new_n1394_), .ZN(new_n1397_) );
  INV_X1 g1261 ( .A(new_n1357_), .ZN(new_n1398_) );
  AND2_X1 g1262 ( .A1(new_n1398_), .A2(new_n1391_), .ZN(new_n1399_) );
  INV_X1 g1263 ( .A(new_n1291_), .ZN(new_n1400_) );
  INV_X1 g1264 ( .A(new_n1343_), .ZN(new_n1401_) );
  OR3_X1 g1265 ( .A1(new_n1400_), .A2(G378), .A3(new_n1401_), .ZN(new_n1402_) );
  INV_X1 g1266 ( .A(new_n1402_), .ZN(new_n1403_) );
  INV_X1 g1267 ( .A(G396), .ZN(new_n1404_) );
  INV_X1 g1268 ( .A(G393), .ZN(new_n1405_) );
  AND4_X1 g1269 ( .A1(new_n1178_), .A2(new_n1404_), .A3(new_n872_), .A4(new_n1405_), .ZN(new_n1406_) );
  AND4_X1 g1270 ( .A1(new_n1403_), .A2(new_n1397_), .A3(new_n1399_), .A4(new_n1406_), .ZN(new_n1407_) );
  INV_X1 g1271 ( .A(new_n1407_), .ZN(G407) );
  INV_X1 g1272 ( .A(G213), .ZN(new_n1409_) );
  INV_X1 g1273 ( .A(G343), .ZN(new_n1410_) );
  AND2_X1 g1274 ( .A1(new_n1403_), .A2(new_n1410_), .ZN(new_n1411_) );
  OR3_X1 g1275 ( .A1(new_n1407_), .A2(new_n1409_), .A3(new_n1411_), .ZN(G409) );
  AND2_X1 g1276 ( .A1(new_n1410_), .A2(G213), .ZN(new_n1413_) );
  AND2_X1 g1277 ( .A1(new_n1413_), .A2(G2897), .ZN(new_n1414_) );
  OR2_X1 g1278 ( .A1(new_n1414_), .A2(KEYINPUT63), .ZN(new_n1415_) );
  AND2_X1 g1279 ( .A1(new_n1414_), .A2(KEYINPUT63), .ZN(new_n1416_) );
  INV_X1 g1280 ( .A(new_n1416_), .ZN(new_n1417_) );
  AND2_X1 g1281 ( .A1(new_n1417_), .A2(new_n1415_), .ZN(new_n1418_) );
  INV_X1 g1282 ( .A(new_n1418_), .ZN(new_n1419_) );
  INV_X1 g1283 ( .A(new_n1413_), .ZN(new_n1420_) );
  INV_X1 g1284 ( .A(G378), .ZN(new_n1421_) );
  OR2_X1 g1285 ( .A1(new_n1344_), .A2(new_n1421_), .ZN(new_n1422_) );
  AND3_X1 g1286 ( .A1(new_n1422_), .A2(new_n1402_), .A3(new_n1420_), .ZN(new_n1423_) );
  INV_X1 g1287 ( .A(new_n1423_), .ZN(new_n1424_) );
  AND2_X1 g1288 ( .A1(new_n1178_), .A2(G396), .ZN(new_n1425_) );
  AND2_X1 g1289 ( .A1(G390), .A2(new_n1404_), .ZN(new_n1426_) );
  OR2_X1 g1290 ( .A1(new_n1426_), .A2(new_n1425_), .ZN(new_n1427_) );
  INV_X1 g1291 ( .A(new_n1427_), .ZN(new_n1428_) );
  AND3_X1 g1292 ( .A1(new_n1428_), .A2(new_n1398_), .A3(new_n1391_), .ZN(new_n1429_) );
  INV_X1 g1293 ( .A(new_n1429_), .ZN(new_n1430_) );
  AND2_X1 g1294 ( .A1(G381), .A2(new_n1427_), .ZN(new_n1431_) );
  INV_X1 g1295 ( .A(new_n1431_), .ZN(new_n1432_) );
  AND2_X1 g1296 ( .A1(G393), .A2(new_n872_), .ZN(new_n1433_) );
  AND2_X1 g1297 ( .A1(new_n1405_), .A2(G384), .ZN(new_n1434_) );
  OR2_X1 g1298 ( .A1(new_n1434_), .A2(new_n1433_), .ZN(new_n1435_) );
  OR3_X1 g1299 ( .A1(new_n1396_), .A2(new_n1394_), .A3(new_n1435_), .ZN(new_n1436_) );
  INV_X1 g1300 ( .A(new_n1435_), .ZN(new_n1437_) );
  OR2_X1 g1301 ( .A1(G387), .A2(new_n1437_), .ZN(new_n1438_) );
  AND2_X1 g1302 ( .A1(new_n1438_), .A2(new_n1436_), .ZN(new_n1439_) );
  AND3_X1 g1303 ( .A1(new_n1439_), .A2(new_n1430_), .A3(new_n1432_), .ZN(new_n1440_) );
  INV_X1 g1304 ( .A(new_n1440_), .ZN(new_n1441_) );
  OR2_X1 g1305 ( .A1(new_n1431_), .A2(new_n1429_), .ZN(new_n1442_) );
  INV_X1 g1306 ( .A(new_n1436_), .ZN(new_n1443_) );
  AND2_X1 g1307 ( .A1(new_n1397_), .A2(new_n1435_), .ZN(new_n1444_) );
  OR2_X1 g1308 ( .A1(new_n1444_), .A2(new_n1443_), .ZN(new_n1445_) );
  AND2_X1 g1309 ( .A1(new_n1442_), .A2(new_n1445_), .ZN(new_n1446_) );
  INV_X1 g1310 ( .A(new_n1446_), .ZN(new_n1447_) );
  AND4_X1 g1311 ( .A1(new_n1447_), .A2(new_n1424_), .A3(new_n1419_), .A4(new_n1441_), .ZN(new_n1448_) );
  OR2_X1 g1312 ( .A1(new_n1423_), .A2(new_n1418_), .ZN(new_n1449_) );
  OR2_X1 g1313 ( .A1(new_n1446_), .A2(new_n1440_), .ZN(new_n1450_) );
  AND2_X1 g1314 ( .A1(new_n1450_), .A2(new_n1449_), .ZN(new_n1451_) );
  OR2_X1 g1315 ( .A1(new_n1451_), .A2(new_n1448_), .ZN(G405) );
  AND2_X1 g1316 ( .A1(new_n1422_), .A2(new_n1402_), .ZN(new_n1453_) );
  AND2_X1 g1317 ( .A1(new_n1450_), .A2(new_n1453_), .ZN(new_n1454_) );
  INV_X1 g1318 ( .A(new_n1453_), .ZN(new_n1455_) );
  AND3_X1 g1319 ( .A1(new_n1447_), .A2(new_n1455_), .A3(new_n1441_), .ZN(new_n1456_) );
  OR2_X1 g1320 ( .A1(new_n1454_), .A2(new_n1456_), .ZN(G402) );
endmodule


