module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n155_, new_n384_, new_n595_, new_n410_, new_n614_, new_n445_, new_n236_, new_n238_, new_n479_, new_n543_, new_n250_, new_n501_, new_n288_, new_n371_, new_n509_, new_n454_, new_n421_, new_n202_, new_n296_, new_n308_, new_n620_, new_n368_, new_n232_, new_n258_, new_n439_, new_n283_, new_n223_, new_n156_, new_n306_, new_n291_, new_n366_, new_n261_, new_n241_, new_n309_, new_n566_, new_n186_, new_n339_, new_n365_, new_n616_, new_n197_, new_n529_, new_n386_, new_n323_, new_n401_, new_n389_, new_n259_, new_n362_, new_n514_, new_n601_, new_n604_, new_n556_, new_n227_, new_n416_, new_n222_, new_n456_, new_n170_, new_n246_, new_n571_, new_n400_, new_n328_, new_n460_, new_n266_, new_n367_, new_n542_, new_n548_, new_n173_, new_n220_, new_n130_, new_n505_, new_n619_, new_n419_, new_n471_, new_n624_, new_n268_, new_n374_, new_n577_, new_n534_, new_n376_, new_n380_, new_n214_, new_n451_, new_n489_, new_n424_, new_n138_, new_n310_, new_n602_, new_n144_, new_n275_, new_n188_, new_n240_, new_n413_, new_n526_, new_n352_, new_n442_, new_n575_, new_n485_, new_n525_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n562_, new_n578_, new_n462_, new_n603_, new_n564_, new_n177_, new_n493_, new_n547_, new_n264_, new_n379_, new_n500_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n317_, new_n344_, new_n143_, new_n520_, new_n287_, new_n125_, new_n253_, new_n504_, new_n403_, new_n475_, new_n237_, new_n427_, new_n234_, new_n532_, new_n472_, new_n557_, new_n393_, new_n260_, new_n418_, new_n251_, new_n189_, new_n300_, new_n292_, new_n411_, new_n215_, new_n507_, new_n152_, new_n605_, new_n157_, new_n182_, new_n407_, new_n153_, new_n480_, new_n625_, new_n133_, new_n257_, new_n481_, new_n212_, new_n151_, new_n513_, new_n592_, new_n364_, new_n449_, new_n580_, new_n484_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n282_, new_n583_, new_n617_, new_n522_, new_n588_, new_n201_, new_n428_, new_n192_, new_n414_, new_n199_, new_n487_, new_n360_, new_n546_, new_n612_, new_n315_, new_n302_, new_n191_, new_n326_, new_n554_, new_n225_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n387_, new_n606_, new_n544_, new_n476_, new_n615_, new_n589_, new_n248_, new_n350_, new_n415_, new_n537_, new_n221_, new_n385_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n478_, new_n461_, new_n459_, new_n569_, new_n555_, new_n174_, new_n297_, new_n361_, new_n565_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n340_, new_n147_, new_n510_, new_n285_, new_n502_, new_n613_, new_n351_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n517_, new_n325_, new_n609_, new_n417_, new_n591_, new_n180_, new_n515_, new_n530_, new_n332_, new_n318_, new_n622_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n321_, new_n440_, new_n443_, new_n324_, new_n122_, new_n531_, new_n593_, new_n252_, new_n585_, new_n486_, new_n491_, new_n549_, new_n466_, new_n262_, new_n160_, new_n312_, new_n271_, new_n535_, new_n274_, new_n372_, new_n242_, new_n503_, new_n527_, new_n218_, new_n497_, new_n307_, new_n190_, new_n305_, new_n420_, new_n568_, new_n597_, new_n408_, new_n470_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n213_, new_n433_, new_n435_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n265_, new_n506_, new_n370_, new_n256_, new_n584_, new_n452_, new_n278_, new_n304_, new_n381_, new_n523_, new_n388_, new_n550_, new_n217_, new_n269_, new_n508_, new_n512_, new_n194_, new_n483_, new_n394_, new_n299_, new_n129_, new_n599_, new_n314_, new_n582_, new_n412_, new_n607_, new_n441_, new_n477_, new_n327_, new_n216_, new_n600_, new_n594_, new_n561_, new_n495_, new_n431_, new_n196_, new_n280_, new_n574_, new_n426_, new_n319_, new_n235_, new_n398_, new_n301_, new_n169_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n338_, new_n207_, new_n267_, new_n473_, new_n140_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n187_, new_n311_, new_n587_, new_n465_, new_n195_, new_n567_, new_n263_, new_n334_, new_n331_, new_n576_, new_n341_, new_n378_, new_n621_, new_n357_, new_n320_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n245_, new_n402_, new_n474_, new_n579_, new_n467_, new_n286_, new_n404_, new_n335_, new_n347_, new_n193_, new_n490_, new_n560_, new_n346_, new_n396_, new_n198_, new_n438_, new_n358_, new_n208_, new_n348_, new_n610_, new_n159_, new_n322_, new_n228_, new_n545_, new_n611_, new_n289_, new_n528_, new_n179_, new_n425_, new_n436_, new_n175_, new_n226_, new_n397_, new_n399_, new_n596_, new_n373_, new_n171_, new_n559_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n233_, new_n136_, new_n469_, new_n284_, new_n119_, new_n391_, new_n293_, new_n178_, new_n437_, new_n551_, new_n168_, new_n279_, new_n455_, new_n295_, new_n359_, new_n132_, new_n618_, new_n120_, new_n521_, new_n166_, new_n162_, new_n457_, new_n553_, new_n406_, new_n356_, new_n333_, new_n229_, new_n536_, new_n290_, new_n464_, new_n204_, new_n369_, new_n181_, new_n135_, new_n448_, new_n573_, new_n276_, new_n405_;

not g000 ( new_n119_, N75 );
nand g001 ( new_n120_, N29, N42 );
nor g002 ( N388, new_n120_, new_n119_ );
not g003 ( new_n122_, N80 );
nand g004 ( new_n123_, N29, N36 );
nor g005 ( N389, new_n123_, new_n122_ );
not g006 ( new_n125_, N42 );
nor g007 ( N390, new_n123_, new_n125_ );
nand g008 ( new_n127_, N85, N86 );
not g009 ( N391, new_n127_ );
not g010 ( new_n129_, N17 );
not g011 ( new_n130_, N13 );
nand g012 ( new_n131_, N1, N8 );
nor g013 ( new_n132_, new_n131_, new_n130_ );
not g014 ( new_n133_, new_n132_ );
nor g015 ( N418, new_n133_, new_n129_ );
not g016 ( new_n135_, N390 );
nand g017 ( new_n136_, N1, N26 );
nand g018 ( new_n137_, N13, N17 );
nor g019 ( new_n138_, new_n136_, new_n137_ );
nand g020 ( N419, new_n135_, new_n138_ );
nand g021 ( new_n140_, N59, N75 );
not g022 ( new_n141_, new_n140_ );
nand g023 ( N420, new_n141_, N80 );
nand g024 ( new_n143_, N36, N59 );
not g025 ( new_n144_, new_n143_ );
nand g026 ( N421, new_n144_, N80 );
nand g027 ( N422, new_n144_, N42 );
not g028 ( new_n147_, N90 );
nor g029 ( new_n148_, N87, N88 );
nor g030 ( N423, new_n148_, new_n147_ );
nand g031 ( N446, new_n138_, N390 );
not g032 ( new_n151_, keyIn_0_0 );
not g033 ( new_n152_, new_n136_ );
nand g034 ( new_n153_, new_n152_, N51 );
nand g035 ( new_n154_, new_n153_, new_n151_ );
not g036 ( new_n155_, N51 );
nor g037 ( new_n156_, new_n136_, new_n155_ );
nand g038 ( new_n157_, new_n156_, keyIn_0_0 );
nand g039 ( N447, new_n154_, new_n157_ );
nand g040 ( new_n159_, new_n132_, N55 );
nand g041 ( new_n160_, N29, N68 );
nor g042 ( N448, new_n159_, new_n160_ );
nand g043 ( new_n162_, N59, N68 );
not g044 ( new_n163_, new_n162_ );
nand g045 ( new_n164_, new_n163_, N74 );
nor g046 ( N449, new_n159_, new_n164_ );
not g047 ( new_n166_, N89 );
nor g048 ( N450, new_n148_, new_n166_ );
xor g049 ( new_n168_, N111, N116 );
xnor g050 ( new_n169_, N121, N126 );
xnor g051 ( new_n170_, new_n168_, new_n169_ );
xnor g052 ( new_n171_, new_n170_, N135 );
xnor g053 ( new_n172_, N91, N96 );
xnor g054 ( new_n173_, N101, N106 );
xnor g055 ( new_n174_, new_n172_, new_n173_ );
xnor g056 ( new_n175_, new_n174_, N130 );
xnor g057 ( N767, new_n171_, new_n175_ );
xor g058 ( new_n177_, N183, N189 );
xnor g059 ( new_n178_, N195, N201 );
xnor g060 ( new_n179_, new_n177_, new_n178_ );
xnor g061 ( new_n180_, new_n179_, N207 );
xnor g062 ( new_n181_, N159, N165 );
xnor g063 ( new_n182_, N171, N177 );
xnor g064 ( new_n183_, new_n181_, new_n182_ );
xnor g065 ( new_n184_, new_n183_, N130 );
xnor g066 ( N768, new_n180_, new_n184_ );
not g067 ( new_n186_, N261 );
not g068 ( new_n187_, N201 );
not g069 ( new_n188_, keyIn_0_9 );
not g070 ( new_n189_, keyIn_0_4 );
nand g071 ( new_n190_, N447, new_n189_ );
xnor g072 ( new_n191_, new_n156_, new_n151_ );
nand g073 ( new_n192_, new_n191_, keyIn_0_4 );
nand g074 ( new_n193_, new_n192_, new_n190_ );
xnor g075 ( new_n194_, new_n193_, keyIn_0_7 );
nand g076 ( new_n195_, N17, N42 );
xnor g077 ( new_n196_, new_n195_, keyIn_0_3 );
nor g078 ( new_n197_, N17, N42 );
xnor g079 ( new_n198_, new_n197_, keyIn_0_2 );
nor g080 ( new_n199_, new_n198_, new_n196_ );
nor g081 ( new_n200_, new_n199_, keyIn_0_6 );
nand g082 ( new_n201_, new_n199_, keyIn_0_6 );
nand g083 ( new_n202_, N59, N156 );
not g084 ( new_n203_, new_n202_ );
nand g085 ( new_n204_, new_n201_, new_n203_ );
nor g086 ( new_n205_, new_n204_, new_n200_ );
nand g087 ( new_n206_, new_n194_, new_n205_ );
nand g088 ( new_n207_, new_n206_, new_n188_ );
not g089 ( new_n208_, keyIn_0_7 );
xnor g090 ( new_n209_, new_n193_, new_n208_ );
not g091 ( new_n210_, new_n205_ );
nor g092 ( new_n211_, new_n209_, new_n210_ );
nand g093 ( new_n212_, new_n211_, keyIn_0_9 );
nand g094 ( new_n213_, new_n212_, new_n207_ );
not g095 ( new_n214_, keyIn_0_5 );
nand g096 ( new_n215_, N17, N51 );
nor g097 ( new_n216_, new_n131_, new_n215_ );
xnor g098 ( new_n217_, new_n216_, keyIn_0_1 );
nor g099 ( new_n218_, new_n217_, new_n214_ );
nand g100 ( new_n219_, new_n217_, new_n214_ );
nand g101 ( new_n220_, new_n141_, N42 );
nand g102 ( new_n221_, new_n219_, new_n220_ );
nor g103 ( new_n222_, new_n221_, new_n218_ );
xnor g104 ( new_n223_, new_n222_, keyIn_0_8 );
not g105 ( new_n224_, new_n223_ );
nand g106 ( new_n225_, new_n213_, new_n224_ );
nor g107 ( new_n226_, new_n225_, keyIn_0_10 );
nand g108 ( new_n227_, new_n225_, keyIn_0_10 );
nand g109 ( new_n228_, new_n227_, N126 );
nor g110 ( new_n229_, new_n228_, new_n226_ );
nand g111 ( new_n230_, N29, N75 );
nor g112 ( new_n231_, new_n230_, new_n122_ );
nand g113 ( new_n232_, new_n194_, new_n231_ );
not g114 ( new_n233_, N268 );
nand g115 ( new_n234_, new_n233_, N55 );
nor g116 ( new_n235_, new_n232_, new_n234_ );
not g117 ( new_n236_, new_n235_ );
nand g118 ( new_n237_, new_n202_, N17 );
not g119 ( new_n238_, new_n237_ );
nand g120 ( new_n239_, new_n194_, new_n238_ );
nand g121 ( new_n240_, new_n239_, N1 );
nand g122 ( new_n241_, new_n240_, N153 );
nand g123 ( new_n242_, new_n241_, new_n236_ );
nor g124 ( new_n243_, new_n229_, new_n242_ );
nor g125 ( new_n244_, new_n243_, new_n187_ );
not g126 ( new_n245_, new_n244_ );
nand g127 ( new_n246_, new_n243_, new_n187_ );
nand g128 ( new_n247_, new_n245_, new_n246_ );
nand g129 ( new_n248_, new_n247_, new_n186_ );
not g130 ( new_n249_, N219 );
nor g131 ( new_n250_, new_n247_, new_n186_ );
nor g132 ( new_n251_, new_n250_, new_n249_ );
nand g133 ( new_n252_, new_n251_, new_n248_ );
not g134 ( new_n253_, N228 );
nor g135 ( new_n254_, new_n247_, new_n253_ );
nand g136 ( new_n255_, new_n244_, N237 );
not g137 ( new_n256_, N246 );
nor g138 ( new_n257_, new_n243_, new_n256_ );
not g139 ( new_n258_, N73 );
nand g140 ( new_n259_, N42, N72 );
nor g141 ( new_n260_, new_n259_, new_n258_ );
nand g142 ( new_n261_, new_n260_, new_n163_ );
nor g143 ( new_n262_, new_n159_, new_n261_ );
nand g144 ( new_n263_, new_n262_, N201 );
nand g145 ( new_n264_, N255, N267 );
nand g146 ( new_n265_, N121, N210 );
nand g147 ( new_n266_, new_n264_, new_n265_ );
not g148 ( new_n267_, new_n266_ );
nand g149 ( new_n268_, new_n263_, new_n267_ );
nor g150 ( new_n269_, new_n257_, new_n268_ );
nand g151 ( new_n270_, new_n269_, new_n255_ );
nor g152 ( new_n271_, new_n254_, new_n270_ );
nand g153 ( N850, new_n252_, new_n271_ );
not g154 ( new_n273_, keyIn_0_14 );
not g155 ( new_n274_, keyIn_0_13 );
not g156 ( new_n275_, keyIn_0_12 );
nand g157 ( new_n276_, new_n227_, N111 );
nor g158 ( new_n277_, new_n276_, new_n226_ );
nand g159 ( new_n278_, new_n277_, keyIn_0_11 );
nand g160 ( new_n279_, new_n240_, N143 );
not g161 ( new_n280_, new_n279_ );
nor g162 ( new_n281_, new_n277_, keyIn_0_11 );
nor g163 ( new_n282_, new_n281_, new_n280_ );
nand g164 ( new_n283_, new_n282_, new_n278_ );
nor g165 ( new_n284_, new_n283_, new_n275_ );
nand g166 ( new_n285_, new_n283_, new_n275_ );
nand g167 ( new_n286_, new_n285_, new_n236_ );
nor g168 ( new_n287_, new_n286_, new_n284_ );
xnor g169 ( new_n288_, new_n287_, new_n274_ );
nand g170 ( new_n289_, new_n288_, N183 );
xnor g171 ( new_n290_, new_n289_, new_n273_ );
not g172 ( new_n291_, keyIn_0_15 );
not g173 ( new_n292_, N183 );
not g174 ( new_n293_, new_n284_ );
not g175 ( new_n294_, new_n278_ );
not g176 ( new_n295_, keyIn_0_11 );
not g177 ( new_n296_, new_n226_ );
not g178 ( new_n297_, new_n276_ );
nand g179 ( new_n298_, new_n297_, new_n296_ );
nand g180 ( new_n299_, new_n298_, new_n295_ );
nand g181 ( new_n300_, new_n299_, new_n279_ );
nor g182 ( new_n301_, new_n300_, new_n294_ );
nor g183 ( new_n302_, new_n301_, keyIn_0_12 );
nor g184 ( new_n303_, new_n302_, new_n235_ );
nand g185 ( new_n304_, new_n303_, new_n293_ );
nand g186 ( new_n305_, new_n304_, new_n274_ );
nand g187 ( new_n306_, new_n287_, keyIn_0_13 );
nand g188 ( new_n307_, new_n305_, new_n306_ );
nand g189 ( new_n308_, new_n307_, new_n292_ );
xnor g190 ( new_n309_, new_n308_, new_n291_ );
nor g191 ( new_n310_, new_n290_, new_n309_ );
xor g192 ( new_n311_, new_n225_, keyIn_0_10 );
nand g193 ( new_n312_, new_n311_, N116 );
nand g194 ( new_n313_, new_n240_, N146 );
nand g195 ( new_n314_, new_n313_, new_n236_ );
not g196 ( new_n315_, new_n314_ );
nand g197 ( new_n316_, new_n312_, new_n315_ );
nor g198 ( new_n317_, new_n316_, N189 );
not g199 ( new_n318_, new_n317_ );
not g200 ( new_n319_, N195 );
nand g201 ( new_n320_, new_n227_, N121 );
nor g202 ( new_n321_, new_n320_, new_n226_ );
nand g203 ( new_n322_, new_n240_, N149 );
nand g204 ( new_n323_, new_n322_, new_n236_ );
nor g205 ( new_n324_, new_n321_, new_n323_ );
nor g206 ( new_n325_, new_n324_, new_n319_ );
not g207 ( new_n326_, new_n325_ );
nand g208 ( new_n327_, new_n324_, new_n319_ );
xnor g209 ( new_n328_, new_n327_, keyIn_0_16 );
not g210 ( new_n329_, keyIn_0_18 );
nand g211 ( new_n330_, new_n246_, N261 );
not g212 ( new_n331_, new_n330_ );
nand g213 ( new_n332_, new_n331_, new_n329_ );
nand g214 ( new_n333_, new_n332_, new_n245_ );
nand g215 ( new_n334_, new_n333_, new_n328_ );
nand g216 ( new_n335_, new_n334_, new_n326_ );
nand g217 ( new_n336_, new_n335_, new_n318_ );
nand g218 ( new_n337_, new_n316_, N189 );
nor g219 ( new_n338_, new_n330_, new_n317_ );
nand g220 ( new_n339_, new_n328_, new_n338_ );
nand g221 ( new_n340_, new_n339_, keyIn_0_18 );
nand g222 ( new_n341_, new_n340_, new_n337_ );
not g223 ( new_n342_, new_n341_ );
nand g224 ( new_n343_, new_n336_, new_n342_ );
nand g225 ( new_n344_, new_n310_, new_n343_ );
nor g226 ( new_n345_, new_n310_, new_n343_ );
nor g227 ( new_n346_, new_n345_, new_n249_ );
nand g228 ( new_n347_, new_n346_, new_n344_ );
not g229 ( new_n348_, N237 );
nand g230 ( new_n349_, new_n289_, keyIn_0_14 );
nor g231 ( new_n350_, new_n307_, new_n292_ );
nand g232 ( new_n351_, new_n350_, new_n273_ );
nand g233 ( new_n352_, new_n351_, new_n349_ );
xnor g234 ( new_n353_, new_n352_, keyIn_0_17 );
nor g235 ( new_n354_, new_n353_, new_n348_ );
nand g236 ( new_n355_, new_n310_, N228 );
nor g237 ( new_n356_, new_n307_, new_n256_ );
nand g238 ( new_n357_, new_n262_, N183 );
nand g239 ( new_n358_, N106, N210 );
nand g240 ( new_n359_, new_n357_, new_n358_ );
nor g241 ( new_n360_, new_n356_, new_n359_ );
nand g242 ( new_n361_, new_n355_, new_n360_ );
nor g243 ( new_n362_, new_n354_, new_n361_ );
nand g244 ( N863, new_n347_, new_n362_ );
not g245 ( new_n364_, new_n337_ );
nor g246 ( new_n365_, new_n364_, new_n317_ );
not g247 ( new_n366_, new_n365_ );
nand g248 ( new_n367_, new_n330_, new_n245_ );
nand g249 ( new_n368_, new_n328_, new_n367_ );
nand g250 ( new_n369_, new_n368_, new_n326_ );
not g251 ( new_n370_, new_n369_ );
nand g252 ( new_n371_, new_n370_, new_n366_ );
nand g253 ( new_n372_, new_n369_, new_n365_ );
nand g254 ( new_n373_, new_n372_, N219 );
not g255 ( new_n374_, new_n373_ );
nand g256 ( new_n375_, new_n374_, new_n371_ );
nor g257 ( new_n376_, new_n366_, new_n253_ );
nand g258 ( new_n377_, new_n364_, N237 );
nand g259 ( new_n378_, new_n316_, N246 );
nand g260 ( new_n379_, new_n262_, N189 );
nand g261 ( new_n380_, N255, N259 );
nand g262 ( new_n381_, N111, N210 );
nand g263 ( new_n382_, new_n380_, new_n381_ );
not g264 ( new_n383_, new_n382_ );
nand g265 ( new_n384_, new_n379_, new_n383_ );
not g266 ( new_n385_, new_n384_ );
nand g267 ( new_n386_, new_n378_, new_n385_ );
not g268 ( new_n387_, new_n386_ );
nand g269 ( new_n388_, new_n387_, new_n377_ );
nor g270 ( new_n389_, new_n376_, new_n388_ );
nand g271 ( N864, new_n375_, new_n389_ );
not g272 ( new_n391_, new_n367_ );
nand g273 ( new_n392_, new_n328_, new_n326_ );
nand g274 ( new_n393_, new_n392_, new_n391_ );
nor g275 ( new_n394_, new_n392_, new_n391_ );
nor g276 ( new_n395_, new_n394_, new_n249_ );
nand g277 ( new_n396_, new_n395_, new_n393_ );
nor g278 ( new_n397_, new_n392_, new_n253_ );
nand g279 ( new_n398_, new_n325_, N237 );
nor g280 ( new_n399_, new_n324_, new_n256_ );
nand g281 ( new_n400_, new_n262_, N195 );
nand g282 ( new_n401_, N255, N260 );
nand g283 ( new_n402_, N116, N210 );
nand g284 ( new_n403_, new_n401_, new_n402_ );
not g285 ( new_n404_, new_n403_ );
nand g286 ( new_n405_, new_n400_, new_n404_ );
nor g287 ( new_n406_, new_n399_, new_n405_ );
nand g288 ( new_n407_, new_n406_, new_n398_ );
nor g289 ( new_n408_, new_n397_, new_n407_ );
nand g290 ( N865, new_n396_, new_n408_ );
not g291 ( new_n410_, keyIn_0_21 );
not g292 ( new_n411_, keyIn_0_17 );
nand g293 ( new_n412_, new_n352_, new_n411_ );
nand g294 ( new_n413_, new_n290_, keyIn_0_17 );
nand g295 ( new_n414_, new_n413_, new_n412_ );
nor g296 ( new_n415_, new_n414_, new_n410_ );
not g297 ( new_n416_, new_n415_ );
not g298 ( new_n417_, keyIn_0_22 );
nor g299 ( new_n418_, new_n308_, new_n291_ );
nand g300 ( new_n419_, new_n308_, new_n291_ );
nand g301 ( new_n420_, new_n419_, new_n343_ );
nor g302 ( new_n421_, new_n420_, new_n418_ );
xnor g303 ( new_n422_, new_n421_, new_n417_ );
nor g304 ( new_n423_, new_n353_, keyIn_0_21 );
nor g305 ( new_n424_, new_n423_, new_n422_ );
nand g306 ( new_n425_, new_n424_, new_n416_ );
nand g307 ( new_n426_, new_n425_, keyIn_0_23 );
not g308 ( new_n427_, keyIn_0_23 );
xnor g309 ( new_n428_, new_n421_, keyIn_0_22 );
nand g310 ( new_n429_, new_n414_, new_n410_ );
nand g311 ( new_n430_, new_n428_, new_n429_ );
nor g312 ( new_n431_, new_n430_, new_n415_ );
nand g313 ( new_n432_, new_n431_, new_n427_ );
nand g314 ( new_n433_, new_n426_, new_n432_ );
not g315 ( new_n434_, N177 );
nand g316 ( new_n435_, new_n311_, N106 );
nand g317 ( new_n436_, new_n202_, N55 );
nor g318 ( new_n437_, new_n209_, new_n436_ );
nand g319 ( new_n438_, new_n437_, N153 );
not g320 ( new_n439_, new_n438_ );
nand g321 ( new_n440_, N138, N152 );
nor g322 ( new_n441_, new_n129_, N268 );
not g323 ( new_n442_, new_n441_ );
nor g324 ( new_n443_, new_n232_, new_n442_ );
not g325 ( new_n444_, new_n443_ );
nand g326 ( new_n445_, new_n444_, new_n440_ );
nor g327 ( new_n446_, new_n445_, new_n439_ );
nand g328 ( new_n447_, new_n435_, new_n446_ );
not g329 ( new_n448_, new_n447_ );
nand g330 ( new_n449_, new_n448_, new_n434_ );
nand g331 ( new_n450_, new_n433_, new_n449_ );
nor g332 ( new_n451_, new_n448_, new_n434_ );
not g333 ( new_n452_, new_n451_ );
nand g334 ( new_n453_, new_n450_, new_n452_ );
not g335 ( new_n454_, N171 );
nand g336 ( new_n455_, new_n311_, N101 );
nand g337 ( new_n456_, new_n437_, N149 );
not g338 ( new_n457_, new_n456_ );
nand g339 ( new_n458_, N17, N138 );
nand g340 ( new_n459_, new_n444_, new_n458_ );
nor g341 ( new_n460_, new_n459_, new_n457_ );
nand g342 ( new_n461_, new_n455_, new_n460_ );
not g343 ( new_n462_, new_n461_ );
nand g344 ( new_n463_, new_n462_, new_n454_ );
nand g345 ( new_n464_, new_n453_, new_n463_ );
nand g346 ( new_n465_, new_n461_, N171 );
nand g347 ( new_n466_, new_n464_, new_n465_ );
not g348 ( new_n467_, N165 );
nand g349 ( new_n468_, new_n311_, N96 );
nand g350 ( new_n469_, new_n437_, N146 );
not g351 ( new_n470_, new_n469_ );
nand g352 ( new_n471_, N51, N138 );
nand g353 ( new_n472_, new_n444_, new_n471_ );
nor g354 ( new_n473_, new_n472_, new_n470_ );
nand g355 ( new_n474_, new_n468_, new_n473_ );
not g356 ( new_n475_, new_n474_ );
nand g357 ( new_n476_, new_n475_, new_n467_ );
nand g358 ( new_n477_, new_n466_, new_n476_ );
nor g359 ( new_n478_, new_n475_, new_n467_ );
not g360 ( new_n479_, new_n478_ );
nand g361 ( new_n480_, new_n477_, new_n479_ );
not g362 ( new_n481_, N159 );
nand g363 ( new_n482_, new_n311_, N91 );
nand g364 ( new_n483_, new_n437_, N143 );
not g365 ( new_n484_, new_n483_ );
nand g366 ( new_n485_, N8, N138 );
nand g367 ( new_n486_, new_n444_, new_n485_ );
nor g368 ( new_n487_, new_n486_, new_n484_ );
nand g369 ( new_n488_, new_n482_, new_n487_ );
not g370 ( new_n489_, new_n488_ );
nand g371 ( new_n490_, new_n489_, new_n481_ );
nand g372 ( new_n491_, new_n480_, new_n490_ );
nor g373 ( new_n492_, new_n489_, new_n481_ );
not g374 ( new_n493_, new_n492_ );
nand g375 ( N866, new_n491_, new_n493_ );
not g376 ( new_n495_, keyIn_0_29 );
not g377 ( new_n496_, keyIn_0_28 );
nand g378 ( new_n497_, new_n452_, new_n449_ );
not g379 ( new_n498_, new_n497_ );
nand g380 ( new_n499_, new_n433_, new_n498_ );
nand g381 ( new_n500_, new_n499_, keyIn_0_25 );
not g382 ( new_n501_, new_n500_ );
nor g383 ( new_n502_, new_n433_, new_n498_ );
nor g384 ( new_n503_, new_n502_, keyIn_0_24 );
nor g385 ( new_n504_, new_n501_, new_n503_ );
not g386 ( new_n505_, keyIn_0_24 );
xnor g387 ( new_n506_, new_n431_, keyIn_0_23 );
nand g388 ( new_n507_, new_n506_, new_n497_ );
nor g389 ( new_n508_, new_n507_, new_n505_ );
nor g390 ( new_n509_, new_n499_, keyIn_0_25 );
nor g391 ( new_n510_, new_n508_, new_n509_ );
nand g392 ( new_n511_, new_n504_, new_n510_ );
nor g393 ( new_n512_, new_n511_, keyIn_0_26 );
not g394 ( new_n513_, new_n512_ );
not g395 ( new_n514_, keyIn_0_26 );
nand g396 ( new_n515_, new_n507_, new_n505_ );
nand g397 ( new_n516_, new_n515_, new_n500_ );
nand g398 ( new_n517_, new_n502_, keyIn_0_24 );
not g399 ( new_n518_, keyIn_0_25 );
nor g400 ( new_n519_, new_n506_, new_n497_ );
nand g401 ( new_n520_, new_n519_, new_n518_ );
nand g402 ( new_n521_, new_n520_, new_n517_ );
nor g403 ( new_n522_, new_n521_, new_n516_ );
nor g404 ( new_n523_, new_n522_, new_n514_ );
nor g405 ( new_n524_, new_n523_, new_n249_ );
nand g406 ( new_n525_, new_n524_, new_n513_ );
nor g407 ( new_n526_, new_n525_, keyIn_0_27 );
not g408 ( new_n527_, new_n526_ );
not g409 ( new_n528_, keyIn_0_27 );
nand g410 ( new_n529_, new_n511_, keyIn_0_26 );
nand g411 ( new_n530_, new_n529_, N219 );
nor g412 ( new_n531_, new_n530_, new_n512_ );
nor g413 ( new_n532_, new_n531_, new_n528_ );
nand g414 ( new_n533_, N101, N210 );
not g415 ( new_n534_, new_n533_ );
nor g416 ( new_n535_, new_n532_, new_n534_ );
nand g417 ( new_n536_, new_n535_, new_n527_ );
nor g418 ( new_n537_, new_n536_, new_n496_ );
not g419 ( new_n538_, new_n537_ );
nand g420 ( new_n539_, new_n525_, keyIn_0_27 );
nand g421 ( new_n540_, new_n539_, new_n533_ );
nor g422 ( new_n541_, new_n540_, new_n526_ );
nor g423 ( new_n542_, new_n541_, keyIn_0_28 );
nor g424 ( new_n543_, new_n497_, new_n253_ );
not g425 ( new_n544_, new_n543_ );
nor g426 ( new_n545_, new_n544_, keyIn_0_20 );
nand g427 ( new_n546_, new_n544_, keyIn_0_20 );
nor g428 ( new_n547_, new_n452_, new_n348_ );
nand g429 ( new_n548_, new_n447_, N246 );
nand g430 ( new_n549_, new_n262_, N177 );
nand g431 ( new_n550_, new_n548_, new_n549_ );
nor g432 ( new_n551_, new_n547_, new_n550_ );
nand g433 ( new_n552_, new_n546_, new_n551_ );
nor g434 ( new_n553_, new_n552_, new_n545_ );
not g435 ( new_n554_, new_n553_ );
nor g436 ( new_n555_, new_n542_, new_n554_ );
nand g437 ( new_n556_, new_n555_, new_n538_ );
nand g438 ( new_n557_, new_n556_, new_n495_ );
nand g439 ( new_n558_, new_n536_, new_n496_ );
nand g440 ( new_n559_, new_n558_, new_n553_ );
nor g441 ( new_n560_, new_n559_, new_n537_ );
nand g442 ( new_n561_, new_n560_, keyIn_0_29 );
nand g443 ( new_n562_, new_n557_, new_n561_ );
nand g444 ( new_n563_, new_n562_, keyIn_0_30 );
not g445 ( new_n564_, keyIn_0_30 );
xnor g446 ( new_n565_, new_n560_, new_n495_ );
nand g447 ( new_n566_, new_n565_, new_n564_ );
nand g448 ( new_n567_, new_n566_, new_n563_ );
nand g449 ( new_n568_, new_n567_, keyIn_0_31 );
not g450 ( new_n569_, keyIn_0_31 );
xnor g451 ( new_n570_, new_n562_, new_n564_ );
nand g452 ( new_n571_, new_n570_, new_n569_ );
nand g453 ( N874, new_n571_, new_n568_ );
nand g454 ( new_n573_, new_n493_, new_n490_ );
not g455 ( new_n574_, new_n573_ );
nand g456 ( new_n575_, new_n480_, new_n574_ );
nor g457 ( new_n576_, new_n480_, new_n574_ );
nor g458 ( new_n577_, new_n576_, new_n249_ );
nand g459 ( new_n578_, new_n577_, new_n575_ );
nor g460 ( new_n579_, new_n573_, new_n253_ );
nand g461 ( new_n580_, new_n492_, N237 );
nand g462 ( new_n581_, new_n488_, N246 );
nand g463 ( new_n582_, new_n262_, N159 );
nand g464 ( new_n583_, N210, N268 );
nand g465 ( new_n584_, new_n582_, new_n583_ );
not g466 ( new_n585_, new_n584_ );
nand g467 ( new_n586_, new_n581_, new_n585_ );
not g468 ( new_n587_, new_n586_ );
nand g469 ( new_n588_, new_n580_, new_n587_ );
nor g470 ( new_n589_, new_n579_, new_n588_ );
nand g471 ( N878, new_n578_, new_n589_ );
nand g472 ( new_n591_, new_n479_, new_n476_ );
not g473 ( new_n592_, new_n591_ );
nand g474 ( new_n593_, new_n466_, new_n592_ );
nor g475 ( new_n594_, new_n466_, new_n592_ );
nor g476 ( new_n595_, new_n594_, new_n249_ );
nand g477 ( new_n596_, new_n595_, new_n593_ );
nor g478 ( new_n597_, new_n591_, new_n253_ );
nand g479 ( new_n598_, new_n478_, N237 );
nand g480 ( new_n599_, new_n474_, N246 );
nand g481 ( new_n600_, new_n262_, N165 );
nand g482 ( new_n601_, N91, N210 );
nand g483 ( new_n602_, new_n600_, new_n601_ );
not g484 ( new_n603_, new_n602_ );
nand g485 ( new_n604_, new_n599_, new_n603_ );
not g486 ( new_n605_, new_n604_ );
nand g487 ( new_n606_, new_n598_, new_n605_ );
nor g488 ( new_n607_, new_n597_, new_n606_ );
nand g489 ( N879, new_n596_, new_n607_ );
xnor g490 ( new_n609_, new_n461_, new_n454_ );
nand g491 ( new_n610_, new_n453_, new_n609_ );
nor g492 ( new_n611_, new_n453_, new_n609_ );
nor g493 ( new_n612_, new_n611_, new_n249_ );
nand g494 ( new_n613_, new_n612_, new_n610_ );
nor g495 ( new_n614_, new_n465_, new_n348_ );
xor g496 ( new_n615_, new_n614_, keyIn_0_19 );
nand g497 ( new_n616_, new_n609_, N228 );
nand g498 ( new_n617_, new_n461_, N246 );
nand g499 ( new_n618_, new_n262_, N171 );
nand g500 ( new_n619_, N96, N210 );
nand g501 ( new_n620_, new_n618_, new_n619_ );
not g502 ( new_n621_, new_n620_ );
nand g503 ( new_n622_, new_n617_, new_n621_ );
not g504 ( new_n623_, new_n622_ );
nand g505 ( new_n624_, new_n616_, new_n623_ );
nor g506 ( new_n625_, new_n615_, new_n624_ );
nand g507 ( N880, new_n613_, new_n625_ );
endmodule