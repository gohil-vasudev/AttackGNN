module locked_c1355 (  G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,  G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT  );
  input  G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n303_, new_n305_, new_n306_, new_n308_, new_n309_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n321_, new_n323_, new_n324_, new_n326_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n336_, new_n338_, new_n340_, new_n341_, new_n343_, new_n344_, new_n346_, new_n348_, new_n350_, new_n351_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n381_, new_n382_, new_n384_, new_n385_, new_n387_, new_n388_, new_n389_, new_n391_, new_n392_, new_n394_, new_n395_, new_n396_, new_n398_, new_n400_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n416_, new_n417_, new_n418_, new_n420_, new_n422_, new_n423_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n431_, new_n432_, new_n434_, new_n436_, new_n437_;
  INV_X1 g000 ( .A(G1GAT), .ZN(new_n138_) );
  XOR2_X1 g001 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(new_n139_) );
  XNOR2_X1 g002 ( .A(G148GAT), .B(KEYINPUT6), .ZN(new_n140_) );
  XNOR2_X1 g003 ( .A(new_n139_), .B(new_n140_), .ZN(new_n141_) );
  XOR2_X1 g004 ( .A(G155GAT), .B(KEYINPUT3), .Z(new_n142_) );
  XNOR2_X1 g005 ( .A(G141GAT), .B(KEYINPUT2), .ZN(new_n143_) );
  XNOR2_X1 g006 ( .A(new_n142_), .B(new_n143_), .ZN(new_n144_) );
  XNOR2_X1 g007 ( .A(G57GAT), .B(KEYINPUT1), .ZN(new_n145_) );
  AND2_X1 g008 ( .A1(G225GAT), .A2(G233GAT), .ZN(new_n146_) );
  XNOR2_X1 g009 ( .A(new_n145_), .B(new_n146_), .ZN(new_n147_) );
  XNOR2_X1 g010 ( .A(new_n144_), .B(new_n147_), .ZN(new_n148_) );
  XNOR2_X1 g011 ( .A(G120GAT), .B(G127GAT), .ZN(new_n149_) );
  XNOR2_X1 g012 ( .A(G113GAT), .B(KEYINPUT0), .ZN(new_n150_) );
  XNOR2_X1 g013 ( .A(new_n149_), .B(new_n150_), .ZN(new_n151_) );
  XNOR2_X1 g014 ( .A(new_n151_), .B(new_n138_), .ZN(new_n152_) );
  XNOR2_X1 g015 ( .A(new_n148_), .B(new_n152_), .ZN(new_n153_) );
  XOR2_X1 g016 ( .A(G29GAT), .B(G134GAT), .Z(new_n154_) );
  XNOR2_X1 g017 ( .A(new_n153_), .B(new_n154_), .ZN(new_n155_) );
  XOR2_X1 g018 ( .A(G85GAT), .B(G162GAT), .Z(new_n156_) );
  XNOR2_X1 g019 ( .A(new_n155_), .B(new_n156_), .ZN(new_n157_) );
  XOR2_X1 g020 ( .A(new_n157_), .B(new_n141_), .Z(new_n158_) );
  INV_X1 g021 ( .A(new_n158_), .ZN(new_n159_) );
  XNOR2_X1 g022 ( .A(G211GAT), .B(G218GAT), .ZN(new_n160_) );
  XNOR2_X1 g023 ( .A(G204GAT), .B(KEYINPUT21), .ZN(new_n161_) );
  XNOR2_X1 g024 ( .A(new_n160_), .B(new_n161_), .ZN(new_n162_) );
  XNOR2_X1 g025 ( .A(new_n162_), .B(G197GAT), .ZN(new_n163_) );
  XOR2_X1 g026 ( .A(new_n163_), .B(new_n144_), .Z(new_n164_) );
  XOR2_X1 g027 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(new_n165_) );
  XNOR2_X1 g028 ( .A(G22GAT), .B(KEYINPUT22), .ZN(new_n166_) );
  XNOR2_X1 g029 ( .A(new_n165_), .B(new_n166_), .ZN(new_n167_) );
  XNOR2_X1 g030 ( .A(G78GAT), .B(G106GAT), .ZN(new_n168_) );
  AND2_X1 g031 ( .A1(new_n168_), .A2(G148GAT), .ZN(new_n169_) );
  AND2_X1 g032 ( .A1(G78GAT), .A2(G106GAT), .ZN(new_n170_) );
  INV_X1 g033 ( .A(new_n170_), .ZN(new_n171_) );
  INV_X1 g034 ( .A(G148GAT), .ZN(new_n172_) );
  OR2_X1 g035 ( .A1(G78GAT), .A2(G106GAT), .ZN(new_n173_) );
  AND2_X1 g036 ( .A1(new_n173_), .A2(new_n172_), .ZN(new_n174_) );
  AND2_X1 g037 ( .A1(new_n174_), .A2(new_n171_), .ZN(new_n175_) );
  OR2_X1 g038 ( .A1(new_n175_), .A2(new_n169_), .ZN(new_n176_) );
  XOR2_X1 g039 ( .A(new_n176_), .B(new_n167_), .Z(new_n177_) );
  XNOR2_X1 g040 ( .A(new_n164_), .B(new_n177_), .ZN(new_n178_) );
  XNOR2_X1 g041 ( .A(G50GAT), .B(G162GAT), .ZN(new_n179_) );
  INV_X1 g042 ( .A(new_n179_), .ZN(new_n180_) );
  XNOR2_X1 g043 ( .A(new_n178_), .B(new_n180_), .ZN(new_n181_) );
  AND2_X1 g044 ( .A1(G228GAT), .A2(G233GAT), .ZN(new_n182_) );
  XOR2_X1 g045 ( .A(new_n181_), .B(new_n182_), .Z(new_n183_) );
  XOR2_X1 g046 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(new_n184_) );
  XNOR2_X1 g047 ( .A(G169GAT), .B(KEYINPUT19), .ZN(new_n185_) );
  XNOR2_X1 g048 ( .A(new_n184_), .B(new_n185_), .ZN(new_n186_) );
  XNOR2_X1 g049 ( .A(G134GAT), .B(G190GAT), .ZN(new_n187_) );
  XNOR2_X1 g050 ( .A(G43GAT), .B(G99GAT), .ZN(new_n188_) );
  XOR2_X1 g051 ( .A(new_n187_), .B(new_n188_), .Z(new_n189_) );
  XNOR2_X1 g052 ( .A(new_n189_), .B(new_n186_), .ZN(new_n190_) );
  XOR2_X1 g053 ( .A(new_n151_), .B(G15GAT), .Z(new_n191_) );
  AND2_X1 g054 ( .A1(G227GAT), .A2(G233GAT), .ZN(new_n192_) );
  XNOR2_X1 g055 ( .A(new_n191_), .B(new_n192_), .ZN(new_n193_) );
  XOR2_X1 g056 ( .A(G176GAT), .B(G183GAT), .Z(new_n194_) );
  XNOR2_X1 g057 ( .A(G71GAT), .B(KEYINPUT20), .ZN(new_n195_) );
  XNOR2_X1 g058 ( .A(new_n194_), .B(new_n195_), .ZN(new_n196_) );
  XNOR2_X1 g059 ( .A(new_n193_), .B(new_n196_), .ZN(new_n197_) );
  XNOR2_X1 g060 ( .A(new_n197_), .B(new_n190_), .ZN(new_n198_) );
  OR2_X1 g061 ( .A1(new_n183_), .A2(new_n198_), .ZN(new_n199_) );
  XOR2_X1 g062 ( .A(new_n199_), .B(KEYINPUT26), .Z(new_n200_) );
  XOR2_X1 g063 ( .A(G36GAT), .B(G190GAT), .Z(new_n201_) );
  XNOR2_X1 g064 ( .A(new_n163_), .B(new_n201_), .ZN(new_n202_) );
  INV_X1 g065 ( .A(G92GAT), .ZN(new_n203_) );
  XNOR2_X1 g066 ( .A(G64GAT), .B(G176GAT), .ZN(new_n204_) );
  XNOR2_X1 g067 ( .A(new_n204_), .B(new_n203_), .ZN(new_n205_) );
  AND2_X1 g068 ( .A1(G226GAT), .A2(G233GAT), .ZN(new_n206_) );
  XNOR2_X1 g069 ( .A(new_n205_), .B(new_n206_), .ZN(new_n207_) );
  XNOR2_X1 g070 ( .A(G8GAT), .B(G183GAT), .ZN(new_n208_) );
  XNOR2_X1 g071 ( .A(new_n207_), .B(new_n208_), .ZN(new_n209_) );
  XNOR2_X1 g072 ( .A(new_n202_), .B(new_n209_), .ZN(new_n210_) );
  XNOR2_X1 g073 ( .A(new_n210_), .B(new_n186_), .ZN(new_n211_) );
  XNOR2_X1 g074 ( .A(new_n211_), .B(KEYINPUT27), .ZN(new_n212_) );
  AND2_X1 g075 ( .A1(new_n200_), .A2(new_n212_), .ZN(new_n213_) );
  INV_X1 g076 ( .A(new_n198_), .ZN(new_n214_) );
  INV_X1 g077 ( .A(new_n211_), .ZN(new_n215_) );
  OR2_X1 g078 ( .A1(new_n214_), .A2(new_n215_), .ZN(new_n216_) );
  AND2_X1 g079 ( .A1(new_n183_), .A2(new_n216_), .ZN(new_n217_) );
  XOR2_X1 g080 ( .A(new_n217_), .B(KEYINPUT25), .Z(new_n218_) );
  OR2_X1 g081 ( .A1(new_n213_), .A2(new_n218_), .ZN(new_n219_) );
  AND2_X1 g082 ( .A1(new_n219_), .A2(new_n158_), .ZN(new_n220_) );
  XNOR2_X1 g083 ( .A(new_n183_), .B(KEYINPUT28), .ZN(new_n221_) );
  AND2_X1 g084 ( .A1(new_n159_), .A2(new_n212_), .ZN(new_n222_) );
  AND2_X1 g085 ( .A1(new_n222_), .A2(new_n214_), .ZN(new_n223_) );
  AND2_X1 g086 ( .A1(new_n223_), .A2(new_n221_), .ZN(new_n224_) );
  OR2_X1 g087 ( .A1(new_n220_), .A2(new_n224_), .ZN(new_n225_) );
  XNOR2_X1 g088 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(new_n226_) );
  XNOR2_X1 g089 ( .A(G64GAT), .B(KEYINPUT15), .ZN(new_n227_) );
  XOR2_X1 g090 ( .A(new_n226_), .B(new_n227_), .Z(new_n228_) );
  XNOR2_X1 g091 ( .A(G78GAT), .B(G155GAT), .ZN(new_n229_) );
  XNOR2_X1 g092 ( .A(G127GAT), .B(G211GAT), .ZN(new_n230_) );
  XNOR2_X1 g093 ( .A(new_n229_), .B(new_n230_), .ZN(new_n231_) );
  XNOR2_X1 g094 ( .A(new_n228_), .B(new_n231_), .ZN(new_n232_) );
  XOR2_X1 g095 ( .A(G57GAT), .B(G71GAT), .Z(new_n233_) );
  XNOR2_X1 g096 ( .A(new_n233_), .B(KEYINPUT13), .ZN(new_n234_) );
  XNOR2_X1 g097 ( .A(G15GAT), .B(G22GAT), .ZN(new_n235_) );
  XNOR2_X1 g098 ( .A(new_n235_), .B(new_n138_), .ZN(new_n236_) );
  XNOR2_X1 g099 ( .A(new_n234_), .B(new_n236_), .ZN(new_n237_) );
  XNOR2_X1 g100 ( .A(new_n232_), .B(new_n237_), .ZN(new_n238_) );
  XOR2_X1 g101 ( .A(new_n238_), .B(new_n208_), .Z(new_n239_) );
  AND2_X1 g102 ( .A1(G231GAT), .A2(G233GAT), .ZN(new_n240_) );
  XNOR2_X1 g103 ( .A(new_n239_), .B(new_n240_), .ZN(new_n241_) );
  XNOR2_X1 g104 ( .A(KEYINPUT11), .B(KEYINPUT10), .ZN(new_n242_) );
  AND2_X1 g105 ( .A1(G232GAT), .A2(G233GAT), .ZN(new_n243_) );
  XNOR2_X1 g106 ( .A(new_n242_), .B(new_n243_), .ZN(new_n244_) );
  XOR2_X1 g107 ( .A(new_n244_), .B(KEYINPUT9), .Z(new_n245_) );
  XNOR2_X1 g108 ( .A(G43GAT), .B(KEYINPUT8), .ZN(new_n246_) );
  AND2_X1 g109 ( .A1(new_n246_), .A2(KEYINPUT7), .ZN(new_n247_) );
  AND2_X1 g110 ( .A1(G43GAT), .A2(KEYINPUT8), .ZN(new_n248_) );
  INV_X1 g111 ( .A(new_n248_), .ZN(new_n249_) );
  INV_X1 g112 ( .A(KEYINPUT7), .ZN(new_n250_) );
  OR2_X1 g113 ( .A1(G43GAT), .A2(KEYINPUT8), .ZN(new_n251_) );
  AND2_X1 g114 ( .A1(new_n251_), .A2(new_n250_), .ZN(new_n252_) );
  AND2_X1 g115 ( .A1(new_n252_), .A2(new_n249_), .ZN(new_n253_) );
  OR2_X1 g116 ( .A1(new_n253_), .A2(new_n247_), .ZN(new_n254_) );
  XOR2_X1 g117 ( .A(G85GAT), .B(G99GAT), .Z(new_n255_) );
  OR2_X1 g118 ( .A1(new_n255_), .A2(new_n203_), .ZN(new_n256_) );
  INV_X1 g119 ( .A(G85GAT), .ZN(new_n257_) );
  INV_X1 g120 ( .A(G99GAT), .ZN(new_n258_) );
  AND2_X1 g121 ( .A1(new_n257_), .A2(new_n258_), .ZN(new_n259_) );
  AND2_X1 g122 ( .A1(G85GAT), .A2(G99GAT), .ZN(new_n260_) );
  OR2_X1 g123 ( .A1(new_n260_), .A2(G92GAT), .ZN(new_n261_) );
  OR2_X1 g124 ( .A1(new_n261_), .A2(new_n259_), .ZN(new_n262_) );
  AND2_X1 g125 ( .A1(new_n262_), .A2(new_n256_), .ZN(new_n263_) );
  XNOR2_X1 g126 ( .A(new_n254_), .B(new_n263_), .ZN(new_n264_) );
  XNOR2_X1 g127 ( .A(new_n264_), .B(new_n245_), .ZN(new_n265_) );
  XNOR2_X1 g128 ( .A(G106GAT), .B(G218GAT), .ZN(new_n266_) );
  XNOR2_X1 g129 ( .A(new_n154_), .B(new_n266_), .ZN(new_n267_) );
  XNOR2_X1 g130 ( .A(new_n265_), .B(new_n267_), .ZN(new_n268_) );
  XNOR2_X1 g131 ( .A(new_n268_), .B(new_n180_), .ZN(new_n269_) );
  XOR2_X1 g132 ( .A(new_n269_), .B(new_n201_), .Z(new_n270_) );
  AND2_X1 g133 ( .A1(new_n270_), .A2(new_n241_), .ZN(new_n271_) );
  XNOR2_X1 g134 ( .A(new_n271_), .B(KEYINPUT16), .ZN(new_n272_) );
  AND2_X1 g135 ( .A1(new_n225_), .A2(new_n272_), .ZN(new_n273_) );
  XNOR2_X1 g136 ( .A(new_n176_), .B(new_n263_), .ZN(new_n274_) );
  XNOR2_X1 g137 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(new_n275_) );
  AND2_X1 g138 ( .A1(G230GAT), .A2(G233GAT), .ZN(new_n276_) );
  XNOR2_X1 g139 ( .A(new_n275_), .B(new_n276_), .ZN(new_n277_) );
  XNOR2_X1 g140 ( .A(new_n277_), .B(KEYINPUT32), .ZN(new_n278_) );
  XNOR2_X1 g141 ( .A(new_n274_), .B(new_n278_), .ZN(new_n279_) );
  XNOR2_X1 g142 ( .A(new_n279_), .B(new_n204_), .ZN(new_n280_) );
  XOR2_X1 g143 ( .A(G120GAT), .B(G204GAT), .Z(new_n281_) );
  XNOR2_X1 g144 ( .A(new_n280_), .B(new_n281_), .ZN(new_n282_) );
  XNOR2_X1 g145 ( .A(new_n282_), .B(new_n234_), .ZN(new_n283_) );
  INV_X1 g146 ( .A(new_n283_), .ZN(new_n284_) );
  XOR2_X1 g147 ( .A(G113GAT), .B(G197GAT), .Z(new_n285_) );
  XNOR2_X1 g148 ( .A(G29GAT), .B(G141GAT), .ZN(new_n286_) );
  XNOR2_X1 g149 ( .A(new_n285_), .B(new_n286_), .ZN(new_n287_) );
  XNOR2_X1 g150 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(new_n288_) );
  XNOR2_X1 g151 ( .A(G8GAT), .B(G169GAT), .ZN(new_n289_) );
  XNOR2_X1 g152 ( .A(new_n288_), .B(new_n289_), .ZN(new_n290_) );
  XNOR2_X1 g153 ( .A(new_n287_), .B(new_n290_), .ZN(new_n291_) );
  XNOR2_X1 g154 ( .A(new_n254_), .B(new_n236_), .ZN(new_n292_) );
  XOR2_X1 g155 ( .A(new_n292_), .B(new_n291_), .Z(new_n293_) );
  XNOR2_X1 g156 ( .A(G36GAT), .B(G50GAT), .ZN(new_n294_) );
  AND2_X1 g157 ( .A1(G229GAT), .A2(G233GAT), .ZN(new_n295_) );
  XNOR2_X1 g158 ( .A(new_n294_), .B(new_n295_), .ZN(new_n296_) );
  XOR2_X1 g159 ( .A(new_n293_), .B(new_n296_), .Z(new_n297_) );
  AND2_X1 g160 ( .A1(new_n284_), .A2(new_n297_), .ZN(new_n298_) );
  AND2_X1 g161 ( .A1(new_n273_), .A2(new_n298_), .ZN(new_n299_) );
  AND2_X1 g162 ( .A1(new_n299_), .A2(new_n159_), .ZN(new_n300_) );
  XNOR2_X1 g163 ( .A(new_n300_), .B(KEYINPUT34), .ZN(new_n301_) );
  XNOR2_X1 g164 ( .A(new_n301_), .B(new_n138_), .ZN(G1324GAT) );
  AND2_X1 g165 ( .A1(new_n299_), .A2(new_n211_), .ZN(new_n303_) );
  XOR2_X1 g166 ( .A(new_n303_), .B(G8GAT), .Z(G1325GAT) );
  AND2_X1 g167 ( .A1(new_n299_), .A2(new_n198_), .ZN(new_n305_) );
  XNOR2_X1 g168 ( .A(G15GAT), .B(KEYINPUT35), .ZN(new_n306_) );
  XNOR2_X1 g169 ( .A(new_n305_), .B(new_n306_), .ZN(G1326GAT) );
  INV_X1 g170 ( .A(new_n221_), .ZN(new_n308_) );
  AND2_X1 g171 ( .A1(new_n299_), .A2(new_n308_), .ZN(new_n309_) );
  XOR2_X1 g172 ( .A(new_n309_), .B(G22GAT), .Z(G1327GAT) );
  INV_X1 g173 ( .A(new_n241_), .ZN(new_n311_) );
  XOR2_X1 g174 ( .A(new_n270_), .B(KEYINPUT36), .Z(new_n312_) );
  AND2_X1 g175 ( .A1(new_n312_), .A2(new_n311_), .ZN(new_n313_) );
  AND2_X1 g176 ( .A1(new_n225_), .A2(new_n313_), .ZN(new_n314_) );
  XOR2_X1 g177 ( .A(new_n314_), .B(KEYINPUT37), .Z(new_n315_) );
  AND2_X1 g178 ( .A1(new_n315_), .A2(new_n298_), .ZN(new_n316_) );
  XNOR2_X1 g179 ( .A(new_n316_), .B(KEYINPUT38), .ZN(new_n317_) );
  AND2_X1 g180 ( .A1(new_n317_), .A2(new_n159_), .ZN(new_n318_) );
  XNOR2_X1 g181 ( .A(G29GAT), .B(KEYINPUT39), .ZN(new_n319_) );
  XNOR2_X1 g182 ( .A(new_n318_), .B(new_n319_), .ZN(G1328GAT) );
  AND2_X1 g183 ( .A1(new_n317_), .A2(new_n211_), .ZN(new_n321_) );
  XOR2_X1 g184 ( .A(new_n321_), .B(G36GAT), .Z(G1329GAT) );
  AND2_X1 g185 ( .A1(new_n317_), .A2(new_n198_), .ZN(new_n323_) );
  XOR2_X1 g186 ( .A(new_n323_), .B(KEYINPUT40), .Z(new_n324_) );
  XNOR2_X1 g187 ( .A(new_n324_), .B(G43GAT), .ZN(G1330GAT) );
  AND2_X1 g188 ( .A1(new_n317_), .A2(new_n308_), .ZN(new_n326_) );
  XOR2_X1 g189 ( .A(new_n326_), .B(G50GAT), .Z(G1331GAT) );
  INV_X1 g190 ( .A(new_n297_), .ZN(new_n328_) );
  INV_X1 g191 ( .A(KEYINPUT41), .ZN(new_n329_) );
  XNOR2_X1 g192 ( .A(new_n283_), .B(new_n329_), .ZN(new_n330_) );
  AND2_X1 g193 ( .A1(new_n330_), .A2(new_n328_), .ZN(new_n331_) );
  AND2_X1 g194 ( .A1(new_n273_), .A2(new_n331_), .ZN(new_n332_) );
  AND2_X1 g195 ( .A1(new_n332_), .A2(new_n159_), .ZN(new_n333_) );
  XOR2_X1 g196 ( .A(G57GAT), .B(KEYINPUT42), .Z(new_n334_) );
  XNOR2_X1 g197 ( .A(new_n333_), .B(new_n334_), .ZN(G1332GAT) );
  AND2_X1 g198 ( .A1(new_n332_), .A2(new_n211_), .ZN(new_n336_) );
  XOR2_X1 g199 ( .A(new_n336_), .B(G64GAT), .Z(G1333GAT) );
  AND2_X1 g200 ( .A1(new_n332_), .A2(new_n198_), .ZN(new_n338_) );
  XOR2_X1 g201 ( .A(new_n338_), .B(G71GAT), .Z(G1334GAT) );
  AND2_X1 g202 ( .A1(new_n332_), .A2(new_n308_), .ZN(new_n340_) );
  XNOR2_X1 g203 ( .A(G78GAT), .B(KEYINPUT43), .ZN(new_n341_) );
  XNOR2_X1 g204 ( .A(new_n340_), .B(new_n341_), .ZN(G1335GAT) );
  AND2_X1 g205 ( .A1(new_n315_), .A2(new_n331_), .ZN(new_n343_) );
  AND2_X1 g206 ( .A1(new_n343_), .A2(new_n159_), .ZN(new_n344_) );
  XNOR2_X1 g207 ( .A(new_n344_), .B(new_n257_), .ZN(G1336GAT) );
  AND2_X1 g208 ( .A1(new_n343_), .A2(new_n211_), .ZN(new_n346_) );
  XNOR2_X1 g209 ( .A(new_n346_), .B(new_n203_), .ZN(G1337GAT) );
  AND2_X1 g210 ( .A1(new_n343_), .A2(new_n198_), .ZN(new_n348_) );
  XNOR2_X1 g211 ( .A(new_n348_), .B(new_n258_), .ZN(G1338GAT) );
  AND2_X1 g212 ( .A1(new_n343_), .A2(new_n308_), .ZN(new_n350_) );
  XNOR2_X1 g213 ( .A(new_n350_), .B(KEYINPUT44), .ZN(new_n351_) );
  XOR2_X1 g214 ( .A(new_n351_), .B(G106GAT), .Z(G1339GAT) );
  INV_X1 g215 ( .A(KEYINPUT48), .ZN(new_n353_) );
  INV_X1 g216 ( .A(KEYINPUT47), .ZN(new_n354_) );
  AND2_X1 g217 ( .A1(new_n330_), .A2(new_n297_), .ZN(new_n355_) );
  AND2_X1 g218 ( .A1(new_n355_), .A2(KEYINPUT46), .ZN(new_n356_) );
  INV_X1 g219 ( .A(new_n356_), .ZN(new_n357_) );
  OR2_X1 g220 ( .A1(new_n355_), .A2(KEYINPUT46), .ZN(new_n358_) );
  AND2_X1 g221 ( .A1(new_n270_), .A2(new_n311_), .ZN(new_n359_) );
  AND2_X1 g222 ( .A1(new_n358_), .A2(new_n359_), .ZN(new_n360_) );
  AND2_X1 g223 ( .A1(new_n360_), .A2(new_n357_), .ZN(new_n361_) );
  AND2_X1 g224 ( .A1(new_n361_), .A2(new_n354_), .ZN(new_n362_) );
  INV_X1 g225 ( .A(new_n362_), .ZN(new_n363_) );
  OR2_X1 g226 ( .A1(new_n361_), .A2(new_n354_), .ZN(new_n364_) );
  AND2_X1 g227 ( .A1(new_n312_), .A2(new_n241_), .ZN(new_n365_) );
  XOR2_X1 g228 ( .A(new_n365_), .B(KEYINPUT45), .Z(new_n366_) );
  AND2_X1 g229 ( .A1(new_n284_), .A2(new_n328_), .ZN(new_n367_) );
  INV_X1 g230 ( .A(new_n367_), .ZN(new_n368_) );
  OR2_X1 g231 ( .A1(new_n366_), .A2(new_n368_), .ZN(new_n369_) );
  AND2_X1 g232 ( .A1(new_n364_), .A2(new_n369_), .ZN(new_n370_) );
  AND2_X1 g233 ( .A1(new_n370_), .A2(new_n363_), .ZN(new_n371_) );
  INV_X1 g234 ( .A(new_n371_), .ZN(new_n372_) );
  OR2_X1 g235 ( .A1(new_n372_), .A2(new_n353_), .ZN(new_n373_) );
  OR2_X1 g236 ( .A1(new_n371_), .A2(KEYINPUT48), .ZN(new_n374_) );
  AND2_X1 g237 ( .A1(new_n374_), .A2(new_n222_), .ZN(new_n375_) );
  AND2_X1 g238 ( .A1(new_n375_), .A2(new_n373_), .ZN(new_n376_) );
  AND2_X1 g239 ( .A1(new_n221_), .A2(new_n198_), .ZN(new_n377_) );
  AND2_X1 g240 ( .A1(new_n376_), .A2(new_n377_), .ZN(new_n378_) );
  AND2_X1 g241 ( .A1(new_n378_), .A2(new_n297_), .ZN(new_n379_) );
  XOR2_X1 g242 ( .A(new_n379_), .B(G113GAT), .Z(G1340GAT) );
  AND2_X1 g243 ( .A1(new_n378_), .A2(new_n330_), .ZN(new_n381_) );
  XNOR2_X1 g244 ( .A(G120GAT), .B(KEYINPUT49), .ZN(new_n382_) );
  XNOR2_X1 g245 ( .A(new_n381_), .B(new_n382_), .ZN(G1341GAT) );
  AND2_X1 g246 ( .A1(new_n378_), .A2(new_n241_), .ZN(new_n384_) );
  XNOR2_X1 g247 ( .A(new_n384_), .B(KEYINPUT50), .ZN(new_n385_) );
  XOR2_X1 g248 ( .A(new_n385_), .B(G127GAT), .Z(G1342GAT) );
  INV_X1 g249 ( .A(new_n270_), .ZN(new_n387_) );
  AND2_X1 g250 ( .A1(new_n378_), .A2(new_n387_), .ZN(new_n388_) );
  XNOR2_X1 g251 ( .A(G134GAT), .B(KEYINPUT51), .ZN(new_n389_) );
  XNOR2_X1 g252 ( .A(new_n388_), .B(new_n389_), .ZN(G1343GAT) );
  AND2_X1 g253 ( .A1(new_n376_), .A2(new_n200_), .ZN(new_n391_) );
  AND2_X1 g254 ( .A1(new_n391_), .A2(new_n297_), .ZN(new_n392_) );
  XOR2_X1 g255 ( .A(new_n392_), .B(G141GAT), .Z(G1344GAT) );
  AND2_X1 g256 ( .A1(new_n391_), .A2(new_n330_), .ZN(new_n394_) );
  XNOR2_X1 g257 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(new_n395_) );
  XNOR2_X1 g258 ( .A(new_n394_), .B(new_n395_), .ZN(new_n396_) );
  XNOR2_X1 g259 ( .A(new_n396_), .B(G148GAT), .ZN(G1345GAT) );
  AND2_X1 g260 ( .A1(new_n391_), .A2(new_n241_), .ZN(new_n398_) );
  XOR2_X1 g261 ( .A(new_n398_), .B(G155GAT), .Z(G1346GAT) );
  AND2_X1 g262 ( .A1(new_n391_), .A2(new_n387_), .ZN(new_n400_) );
  XOR2_X1 g263 ( .A(new_n400_), .B(G162GAT), .Z(G1347GAT) );
  INV_X1 g264 ( .A(KEYINPUT55), .ZN(new_n402_) );
  INV_X1 g265 ( .A(KEYINPUT54), .ZN(new_n403_) );
  AND2_X1 g266 ( .A1(new_n374_), .A2(new_n211_), .ZN(new_n404_) );
  AND2_X1 g267 ( .A1(new_n404_), .A2(new_n373_), .ZN(new_n405_) );
  OR2_X1 g268 ( .A1(new_n405_), .A2(new_n403_), .ZN(new_n406_) );
  AND2_X1 g269 ( .A1(new_n406_), .A2(new_n158_), .ZN(new_n407_) );
  AND2_X1 g270 ( .A1(new_n405_), .A2(new_n403_), .ZN(new_n408_) );
  INV_X1 g271 ( .A(new_n408_), .ZN(new_n409_) );
  AND2_X1 g272 ( .A1(new_n409_), .A2(new_n183_), .ZN(new_n410_) );
  AND2_X1 g273 ( .A1(new_n410_), .A2(new_n407_), .ZN(new_n411_) );
  XNOR2_X1 g274 ( .A(new_n411_), .B(new_n402_), .ZN(new_n412_) );
  AND2_X1 g275 ( .A1(new_n412_), .A2(new_n198_), .ZN(new_n413_) );
  AND2_X1 g276 ( .A1(new_n413_), .A2(new_n297_), .ZN(new_n414_) );
  XOR2_X1 g277 ( .A(new_n414_), .B(G169GAT), .Z(G1348GAT) );
  AND2_X1 g278 ( .A1(new_n413_), .A2(new_n330_), .ZN(new_n416_) );
  XNOR2_X1 g279 ( .A(KEYINPUT57), .B(KEYINPUT56), .ZN(new_n417_) );
  XNOR2_X1 g280 ( .A(new_n416_), .B(new_n417_), .ZN(new_n418_) );
  XNOR2_X1 g281 ( .A(new_n418_), .B(G176GAT), .ZN(G1349GAT) );
  AND2_X1 g282 ( .A1(new_n413_), .A2(new_n241_), .ZN(new_n420_) );
  XOR2_X1 g283 ( .A(new_n420_), .B(G183GAT), .Z(G1350GAT) );
  AND2_X1 g284 ( .A1(new_n413_), .A2(new_n387_), .ZN(new_n422_) );
  XOR2_X1 g285 ( .A(G190GAT), .B(KEYINPUT58), .Z(new_n423_) );
  XNOR2_X1 g286 ( .A(new_n422_), .B(new_n423_), .ZN(G1351GAT) );
  AND2_X1 g287 ( .A1(new_n409_), .A2(new_n200_), .ZN(new_n425_) );
  AND2_X1 g288 ( .A1(new_n425_), .A2(new_n407_), .ZN(new_n426_) );
  AND2_X1 g289 ( .A1(new_n426_), .A2(new_n297_), .ZN(new_n427_) );
  XNOR2_X1 g290 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(new_n428_) );
  XNOR2_X1 g291 ( .A(new_n427_), .B(new_n428_), .ZN(new_n429_) );
  XNOR2_X1 g292 ( .A(new_n429_), .B(G197GAT), .ZN(G1352GAT) );
  XNOR2_X1 g293 ( .A(G204GAT), .B(KEYINPUT61), .ZN(new_n431_) );
  AND2_X1 g294 ( .A1(new_n426_), .A2(new_n283_), .ZN(new_n432_) );
  XNOR2_X1 g295 ( .A(new_n432_), .B(new_n431_), .ZN(G1353GAT) );
  AND2_X1 g296 ( .A1(new_n426_), .A2(new_n241_), .ZN(new_n434_) );
  XOR2_X1 g297 ( .A(new_n434_), .B(G211GAT), .Z(G1354GAT) );
  AND2_X1 g298 ( .A1(new_n426_), .A2(new_n312_), .ZN(new_n436_) );
  XNOR2_X1 g299 ( .A(new_n436_), .B(KEYINPUT62), .ZN(new_n437_) );
  XOR2_X1 g300 ( .A(new_n437_), .B(G218GAT), .Z(G1355GAT) );
endmodule


