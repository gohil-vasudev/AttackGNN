module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n614_, new_n445_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n421_, new_n439_, new_n283_, new_n223_, new_n390_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n456_, new_n246_, new_n170_, new_n266_, new_n367_, new_n542_, new_n173_, new_n220_, new_n419_, new_n534_, new_n214_, new_n489_, new_n424_, new_n602_, new_n188_, new_n240_, new_n413_, new_n526_, new_n442_, new_n211_, new_n552_, new_n342_, new_n462_, new_n603_, new_n564_, new_n500_, new_n317_, new_n287_, new_n504_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n152_, new_n157_, new_n153_, new_n257_, new_n481_, new_n212_, new_n449_, new_n484_, new_n272_, new_n282_, new_n201_, new_n192_, new_n414_, new_n315_, new_n326_, new_n554_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n589_, new_n248_, new_n167_, new_n385_, new_n478_, new_n461_, new_n297_, new_n361_, new_n565_, new_n150_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n180_, new_n530_, new_n318_, new_n321_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n549_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n506_, new_n256_, new_n452_, new_n381_, new_n388_, new_n508_, new_n194_, new_n483_, new_n394_, new_n299_, new_n142_, new_n139_, new_n314_, new_n582_, new_n363_, new_n165_, new_n441_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n187_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n402_, new_n579_, new_n286_, new_n335_, new_n347_, new_n396_, new_n198_, new_n438_, new_n208_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n399_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n553_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n155_, new_n384_, new_n410_, new_n543_, new_n371_, new_n454_, new_n202_, new_n296_, new_n308_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n309_, new_n529_, new_n323_, new_n259_, new_n362_, new_n604_, new_n227_, new_n416_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n505_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n138_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n562_, new_n578_, new_n177_, new_n493_, new_n547_, new_n264_, new_n273_, new_n224_, new_n586_, new_n270_, new_n598_, new_n570_, new_n143_, new_n520_, new_n145_, new_n253_, new_n403_, new_n475_, new_n237_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n605_, new_n182_, new_n407_, new_n480_, new_n151_, new_n513_, new_n592_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n588_, new_n428_, new_n199_, new_n146_, new_n487_, new_n546_, new_n612_, new_n302_, new_n191_, new_n225_, new_n387_, new_n544_, new_n476_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n444_, new_n392_, new_n518_, new_n340_, new_n147_, new_n285_, new_n502_, new_n209_, new_n337_, new_n446_, new_n203_, new_n316_, new_n590_, new_n417_, new_n591_, new_n515_, new_n332_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n440_, new_n531_, new_n252_, new_n585_, new_n160_, new_n312_, new_n372_, new_n242_, new_n503_, new_n527_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n433_, new_n435_, new_n265_, new_n584_, new_n278_, new_n304_, new_n523_, new_n550_, new_n217_, new_n269_, new_n512_, new_n599_, new_n412_, new_n607_, new_n327_, new_n594_, new_n561_, new_n495_, new_n431_, new_n196_, new_n574_, new_n319_, new_n338_, new_n336_, new_n247_, new_n539_, new_n330_, new_n294_, new_n195_, new_n576_, new_n357_, new_n320_, new_n245_, new_n474_, new_n467_, new_n404_, new_n193_, new_n560_, new_n610_, new_n159_, new_n322_, new_n228_, new_n545_, new_n289_, new_n425_, new_n175_, new_n226_, new_n185_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n551_, new_n168_, new_n279_, new_n455_, new_n521_, new_n406_, new_n229_, new_n536_, new_n204_, new_n181_, new_n573_, new_n405_;

xnor g000 ( new_n138_, N65, N69 );
xnor g001 ( new_n139_, N73, N77 );
xnor g002 ( new_n140_, new_n138_, new_n139_ );
xnor g003 ( new_n141_, N81, N85 );
xnor g004 ( new_n142_, N89, N93 );
xnor g005 ( new_n143_, new_n141_, new_n142_ );
xnor g006 ( new_n144_, new_n140_, new_n143_ );
nand g007 ( new_n145_, N129, N137 );
xnor g008 ( new_n146_, new_n144_, new_n145_ );
xor g009 ( new_n147_, N1, N17 );
xnor g010 ( new_n148_, N33, N49 );
xnor g011 ( new_n149_, new_n147_, new_n148_ );
xor g012 ( new_n150_, new_n146_, new_n149_ );
not g013 ( new_n151_, new_n150_ );
xor g014 ( new_n152_, N65, N81 );
xnor g015 ( new_n153_, new_n152_, keyIn_0_8 );
xnor g016 ( new_n154_, N97, N113 );
xnor g017 ( new_n155_, new_n154_, keyIn_0_9 );
xnor g018 ( new_n156_, new_n153_, new_n155_ );
xnor g019 ( new_n157_, new_n156_, keyIn_0_16 );
not g020 ( new_n158_, new_n157_ );
not g021 ( new_n159_, keyIn_0_20 );
not g022 ( new_n160_, keyIn_0_18 );
nand g023 ( new_n161_, N1, N5 );
or g024 ( new_n162_, N1, N5 );
nand g025 ( new_n163_, new_n162_, new_n161_ );
nand g026 ( new_n164_, new_n163_, keyIn_0_0 );
not g027 ( new_n165_, keyIn_0_0 );
nand g028 ( new_n166_, new_n162_, new_n165_, new_n161_ );
xnor g029 ( new_n167_, N9, N13 );
nand g030 ( new_n168_, new_n167_, keyIn_0_1 );
not g031 ( new_n169_, keyIn_0_1 );
nand g032 ( new_n170_, N9, N13 );
or g033 ( new_n171_, N9, N13 );
nand g034 ( new_n172_, new_n171_, new_n169_, new_n170_ );
nand g035 ( new_n173_, new_n164_, new_n168_, new_n166_, new_n172_ );
nand g036 ( new_n174_, new_n164_, new_n166_ );
nand g037 ( new_n175_, new_n168_, new_n172_ );
nand g038 ( new_n176_, new_n174_, new_n175_ );
nand g039 ( new_n177_, new_n176_, keyIn_0_12, new_n173_ );
not g040 ( new_n178_, keyIn_0_12 );
nand g041 ( new_n179_, new_n176_, new_n173_ );
nand g042 ( new_n180_, new_n179_, new_n178_ );
not g043 ( new_n181_, keyIn_0_13 );
nand g044 ( new_n182_, N17, N21 );
or g045 ( new_n183_, N17, N21 );
nand g046 ( new_n184_, new_n183_, new_n182_ );
nand g047 ( new_n185_, new_n184_, keyIn_0_2 );
not g048 ( new_n186_, keyIn_0_2 );
nand g049 ( new_n187_, new_n183_, new_n186_, new_n182_ );
nand g050 ( new_n188_, N25, N29 );
or g051 ( new_n189_, N25, N29 );
nand g052 ( new_n190_, new_n189_, new_n188_ );
nand g053 ( new_n191_, new_n190_, keyIn_0_3 );
not g054 ( new_n192_, keyIn_0_3 );
nand g055 ( new_n193_, new_n189_, new_n192_, new_n188_ );
nand g056 ( new_n194_, new_n185_, new_n191_, new_n187_, new_n193_ );
nand g057 ( new_n195_, new_n185_, new_n187_ );
nand g058 ( new_n196_, new_n191_, new_n193_ );
nand g059 ( new_n197_, new_n195_, new_n196_ );
nand g060 ( new_n198_, new_n197_, new_n181_, new_n194_ );
nand g061 ( new_n199_, new_n197_, new_n194_ );
nand g062 ( new_n200_, new_n199_, keyIn_0_13 );
nand g063 ( new_n201_, new_n200_, new_n198_ );
nand g064 ( new_n202_, new_n201_, new_n177_, new_n180_ );
nand g065 ( new_n203_, new_n180_, new_n177_ );
nand g066 ( new_n204_, new_n203_, new_n198_, new_n200_ );
nand g067 ( new_n205_, new_n202_, new_n204_ );
nand g068 ( new_n206_, new_n205_, new_n160_ );
nand g069 ( new_n207_, new_n202_, new_n204_, keyIn_0_18 );
nand g070 ( new_n208_, N133, N137 );
xor g071 ( new_n209_, new_n208_, keyIn_0_6 );
nand g072 ( new_n210_, new_n206_, new_n207_, new_n209_ );
nand g073 ( new_n211_, new_n206_, new_n207_ );
not g074 ( new_n212_, new_n209_ );
nand g075 ( new_n213_, new_n211_, new_n212_ );
nand g076 ( new_n214_, new_n213_, new_n159_, new_n210_ );
nand g077 ( new_n215_, new_n213_, new_n210_ );
nand g078 ( new_n216_, new_n215_, keyIn_0_20 );
nand g079 ( new_n217_, new_n216_, new_n214_ );
nand g080 ( new_n218_, new_n217_, new_n158_ );
nand g081 ( new_n219_, new_n216_, new_n157_, new_n214_ );
nand g082 ( new_n220_, new_n218_, keyIn_0_22, new_n219_ );
not g083 ( new_n221_, keyIn_0_22 );
nand g084 ( new_n222_, new_n218_, new_n219_ );
nand g085 ( new_n223_, new_n222_, new_n221_ );
nand g086 ( new_n224_, new_n223_, new_n220_ );
nand g087 ( new_n225_, N33, N37 );
or g088 ( new_n226_, N33, N37 );
nand g089 ( new_n227_, new_n226_, new_n225_ );
nand g090 ( new_n228_, new_n227_, keyIn_0_4 );
not g091 ( new_n229_, keyIn_0_4 );
nand g092 ( new_n230_, new_n226_, new_n229_, new_n225_ );
nand g093 ( new_n231_, N41, N45 );
or g094 ( new_n232_, N41, N45 );
nand g095 ( new_n233_, new_n232_, new_n231_ );
nand g096 ( new_n234_, new_n233_, keyIn_0_5 );
not g097 ( new_n235_, keyIn_0_5 );
nand g098 ( new_n236_, new_n232_, new_n235_, new_n231_ );
nand g099 ( new_n237_, new_n228_, new_n234_, new_n230_, new_n236_ );
nand g100 ( new_n238_, new_n228_, new_n230_ );
nand g101 ( new_n239_, new_n234_, new_n236_ );
nand g102 ( new_n240_, new_n238_, new_n239_ );
nand g103 ( new_n241_, new_n240_, keyIn_0_14, new_n237_ );
not g104 ( new_n242_, keyIn_0_14 );
nand g105 ( new_n243_, new_n240_, new_n237_ );
nand g106 ( new_n244_, new_n243_, new_n242_ );
nand g107 ( new_n245_, new_n244_, new_n241_ );
xor g108 ( new_n246_, N49, N53 );
xnor g109 ( new_n247_, N57, N61 );
xnor g110 ( new_n248_, new_n246_, new_n247_ );
xnor g111 ( new_n249_, new_n245_, new_n248_ );
nand g112 ( new_n250_, N134, N137 );
xnor g113 ( new_n251_, new_n249_, new_n250_ );
xnor g114 ( new_n252_, N69, N85 );
xnor g115 ( new_n253_, N101, N117 );
xnor g116 ( new_n254_, new_n252_, new_n253_ );
not g117 ( new_n255_, new_n254_ );
nand g118 ( new_n256_, new_n251_, new_n255_ );
or g119 ( new_n257_, new_n251_, new_n255_ );
nand g120 ( new_n258_, new_n257_, new_n256_ );
not g121 ( new_n259_, new_n258_ );
and g122 ( new_n260_, new_n224_, new_n259_ );
not g123 ( new_n261_, keyIn_0_23 );
xor g124 ( new_n262_, N73, N89 );
xnor g125 ( new_n263_, new_n262_, keyIn_0_10 );
xnor g126 ( new_n264_, N105, N121 );
xnor g127 ( new_n265_, new_n264_, keyIn_0_11 );
xnor g128 ( new_n266_, new_n263_, new_n265_ );
xor g129 ( new_n267_, new_n266_, keyIn_0_17 );
not g130 ( new_n268_, new_n267_ );
not g131 ( new_n269_, keyIn_0_21 );
and g132 ( new_n270_, N135, N137 );
or g133 ( new_n271_, new_n270_, keyIn_0_7 );
nand g134 ( new_n272_, keyIn_0_7, N135, N137 );
not g135 ( new_n273_, keyIn_0_19 );
nand g136 ( new_n274_, new_n245_, new_n177_, new_n180_ );
nand g137 ( new_n275_, new_n203_, new_n241_, new_n244_ );
nand g138 ( new_n276_, new_n274_, new_n275_ );
nand g139 ( new_n277_, new_n276_, new_n273_ );
nand g140 ( new_n278_, new_n274_, new_n275_, keyIn_0_19 );
nand g141 ( new_n279_, new_n277_, new_n271_, new_n272_, new_n278_ );
nand g142 ( new_n280_, new_n271_, new_n272_ );
nand g143 ( new_n281_, new_n277_, new_n278_ );
nand g144 ( new_n282_, new_n281_, new_n280_ );
nand g145 ( new_n283_, new_n282_, new_n269_, new_n279_ );
nand g146 ( new_n284_, new_n282_, new_n279_ );
nand g147 ( new_n285_, new_n284_, keyIn_0_21 );
nand g148 ( new_n286_, new_n285_, new_n268_, new_n283_ );
nand g149 ( new_n287_, new_n285_, new_n283_ );
nand g150 ( new_n288_, new_n287_, new_n267_ );
nand g151 ( new_n289_, new_n288_, new_n286_ );
nand g152 ( new_n290_, new_n289_, new_n261_ );
nand g153 ( new_n291_, new_n288_, keyIn_0_23, new_n286_ );
nand g154 ( new_n292_, new_n290_, new_n291_ );
xnor g155 ( new_n293_, N97, N101 );
xnor g156 ( new_n294_, N105, N109 );
xnor g157 ( new_n295_, new_n293_, new_n294_ );
xnor g158 ( new_n296_, new_n140_, new_n295_ );
nand g159 ( new_n297_, N131, N137 );
xnor g160 ( new_n298_, new_n296_, new_n297_ );
xor g161 ( new_n299_, N9, N25 );
xnor g162 ( new_n300_, N41, N57 );
xnor g163 ( new_n301_, new_n299_, new_n300_ );
xor g164 ( new_n302_, new_n298_, new_n301_ );
not g165 ( new_n303_, new_n302_ );
nand g166 ( new_n304_, new_n151_, new_n303_, keyIn_0_24 );
nand g167 ( new_n305_, new_n303_, keyIn_0_24 );
nand g168 ( new_n306_, new_n305_, new_n150_ );
xnor g169 ( new_n307_, N113, N117 );
xnor g170 ( new_n308_, N121, N125 );
xnor g171 ( new_n309_, new_n307_, new_n308_ );
xnor g172 ( new_n310_, new_n295_, new_n309_ );
nand g173 ( new_n311_, N130, N137 );
xnor g174 ( new_n312_, new_n310_, new_n311_ );
xor g175 ( new_n313_, N5, N21 );
xnor g176 ( new_n314_, N37, N53 );
xnor g177 ( new_n315_, new_n313_, new_n314_ );
xor g178 ( new_n316_, new_n312_, new_n315_ );
nand g179 ( new_n317_, new_n306_, new_n304_, new_n316_ );
not g180 ( new_n318_, new_n316_ );
nand g181 ( new_n319_, new_n318_, new_n150_, new_n302_ );
nand g182 ( new_n320_, new_n317_, new_n319_ );
xnor g183 ( new_n321_, new_n143_, new_n309_ );
nand g184 ( new_n322_, N132, N137 );
xnor g185 ( new_n323_, new_n321_, new_n322_ );
xor g186 ( new_n324_, N13, N29 );
xnor g187 ( new_n325_, N45, N61 );
xnor g188 ( new_n326_, new_n324_, new_n325_ );
xor g189 ( new_n327_, new_n326_, keyIn_0_15 );
xnor g190 ( new_n328_, new_n323_, new_n327_ );
nand g191 ( new_n329_, new_n320_, new_n328_ );
not g192 ( new_n330_, new_n328_ );
nand g193 ( new_n331_, new_n150_, new_n330_, new_n302_, new_n316_ );
nand g194 ( new_n332_, new_n329_, new_n331_ );
xnor g195 ( new_n333_, new_n201_, new_n248_ );
nand g196 ( new_n334_, N136, N137 );
xnor g197 ( new_n335_, new_n333_, new_n334_ );
xor g198 ( new_n336_, N77, N93 );
xnor g199 ( new_n337_, N109, N125 );
xnor g200 ( new_n338_, new_n336_, new_n337_ );
xnor g201 ( new_n339_, new_n335_, new_n338_ );
not g202 ( new_n340_, new_n339_ );
and g203 ( new_n341_, new_n292_, new_n332_, new_n340_ );
and g204 ( new_n342_, new_n341_, new_n260_ );
nand g205 ( new_n343_, new_n342_, new_n151_ );
xnor g206 ( N724, new_n343_, N1 );
nand g207 ( new_n345_, new_n342_, new_n318_ );
xnor g208 ( N725, new_n345_, N5 );
nand g209 ( new_n347_, new_n342_, new_n303_ );
xnor g210 ( N726, new_n347_, N9 );
nand g211 ( new_n349_, new_n342_, new_n330_ );
xnor g212 ( N727, new_n349_, N13 );
and g213 ( new_n351_, new_n290_, new_n332_, new_n291_, new_n339_ );
and g214 ( new_n352_, new_n351_, new_n260_ );
nand g215 ( new_n353_, new_n352_, new_n151_ );
xnor g216 ( N728, new_n353_, N17 );
nand g217 ( new_n355_, new_n352_, new_n318_ );
xnor g218 ( N729, new_n355_, N21 );
nand g219 ( new_n357_, new_n352_, new_n303_ );
xnor g220 ( N730, new_n357_, N25 );
nand g221 ( new_n359_, new_n352_, new_n330_ );
xnor g222 ( N731, new_n359_, N29 );
nor g223 ( new_n361_, new_n224_, new_n259_ );
and g224 ( new_n362_, new_n341_, new_n361_ );
nand g225 ( new_n363_, new_n362_, new_n151_ );
xnor g226 ( N732, new_n363_, N33 );
nand g227 ( new_n365_, new_n362_, new_n318_ );
xnor g228 ( N733, new_n365_, N37 );
nand g229 ( new_n367_, new_n362_, new_n303_ );
xnor g230 ( N734, new_n367_, N41 );
nand g231 ( new_n369_, new_n362_, new_n330_ );
xnor g232 ( N735, new_n369_, N45 );
and g233 ( new_n371_, new_n351_, new_n361_ );
nand g234 ( new_n372_, new_n371_, new_n151_ );
xnor g235 ( N736, new_n372_, N49 );
nand g236 ( new_n374_, new_n371_, new_n318_ );
xnor g237 ( N737, new_n374_, N53 );
nand g238 ( new_n376_, new_n371_, new_n303_ );
xnor g239 ( N738, new_n376_, N57 );
nand g240 ( new_n378_, new_n371_, new_n330_ );
xnor g241 ( N739, new_n378_, N61 );
not g242 ( new_n380_, keyIn_0_52 );
not g243 ( new_n381_, N65 );
nand g244 ( new_n382_, new_n223_, keyIn_0_25, new_n220_ );
and g245 ( new_n383_, new_n258_, keyIn_0_26 );
nor g246 ( new_n384_, new_n258_, keyIn_0_26 );
nor g247 ( new_n385_, new_n383_, new_n384_, new_n340_ );
and g248 ( new_n386_, new_n382_, new_n385_ );
not g249 ( new_n387_, keyIn_0_25 );
nand g250 ( new_n388_, new_n224_, new_n387_ );
not g251 ( new_n389_, keyIn_0_27 );
nand g252 ( new_n390_, new_n292_, new_n389_ );
nand g253 ( new_n391_, new_n290_, keyIn_0_27, new_n291_ );
nand g254 ( new_n392_, new_n386_, new_n388_, new_n390_, new_n391_ );
xnor g255 ( new_n393_, new_n392_, keyIn_0_32 );
not g256 ( new_n394_, keyIn_0_34 );
nand g257 ( new_n395_, new_n223_, keyIn_0_29, new_n220_ );
not g258 ( new_n396_, keyIn_0_29 );
nand g259 ( new_n397_, new_n224_, new_n396_ );
nand g260 ( new_n398_, new_n397_, new_n395_ );
nand g261 ( new_n399_, new_n292_, keyIn_0_30 );
not g262 ( new_n400_, keyIn_0_30 );
nand g263 ( new_n401_, new_n290_, new_n400_, new_n291_ );
nor g264 ( new_n402_, new_n259_, new_n339_ );
and g265 ( new_n403_, new_n401_, new_n402_ );
nand g266 ( new_n404_, new_n398_, new_n403_, new_n399_ );
nand g267 ( new_n405_, new_n404_, new_n394_ );
nand g268 ( new_n406_, new_n398_, new_n403_, keyIn_0_34, new_n399_ );
and g269 ( new_n407_, new_n405_, new_n406_ );
not g270 ( new_n408_, keyIn_0_33 );
nand g271 ( new_n409_, new_n224_, keyIn_0_28 );
not g272 ( new_n410_, keyIn_0_28 );
nand g273 ( new_n411_, new_n223_, new_n410_, new_n220_ );
nor g274 ( new_n412_, new_n258_, new_n339_ );
nand g275 ( new_n413_, new_n409_, new_n292_, new_n411_, new_n412_ );
xnor g276 ( new_n414_, new_n413_, new_n408_ );
nand g277 ( new_n415_, new_n290_, keyIn_0_31, new_n291_ );
not g278 ( new_n416_, keyIn_0_31 );
nand g279 ( new_n417_, new_n292_, new_n416_ );
nand g280 ( new_n418_, new_n417_, new_n415_ );
and g281 ( new_n419_, new_n224_, new_n259_, new_n340_ );
nand g282 ( new_n420_, new_n418_, new_n419_ );
nand g283 ( new_n421_, new_n420_, keyIn_0_35 );
not g284 ( new_n422_, keyIn_0_35 );
nand g285 ( new_n423_, new_n418_, new_n419_, new_n422_ );
nand g286 ( new_n424_, new_n339_, keyIn_0_35 );
nand g287 ( new_n425_, new_n421_, new_n423_, new_n424_ );
nand g288 ( new_n426_, new_n393_, new_n407_, new_n414_, new_n425_ );
nand g289 ( new_n427_, new_n426_, keyIn_0_36 );
nand g290 ( new_n428_, new_n421_, new_n423_ );
not g291 ( new_n429_, keyIn_0_36 );
and g292 ( new_n430_, new_n414_, new_n429_ );
nand g293 ( new_n431_, new_n430_, new_n393_, new_n407_, new_n428_ );
nand g294 ( new_n432_, new_n427_, new_n431_ );
nand g295 ( new_n433_, new_n151_, new_n316_ );
nand g296 ( new_n434_, new_n303_, new_n328_ );
nor g297 ( new_n435_, new_n433_, new_n434_ );
nand g298 ( new_n436_, new_n432_, new_n435_ );
nand g299 ( new_n437_, new_n436_, keyIn_0_37 );
not g300 ( new_n438_, keyIn_0_37 );
nand g301 ( new_n439_, new_n432_, new_n438_, new_n435_ );
nand g302 ( new_n440_, new_n437_, new_n439_ );
nand g303 ( new_n441_, new_n440_, new_n224_ );
nand g304 ( new_n442_, new_n441_, keyIn_0_40 );
not g305 ( new_n443_, keyIn_0_40 );
nand g306 ( new_n444_, new_n440_, new_n443_, new_n224_ );
nand g307 ( new_n445_, new_n442_, new_n444_ );
nand g308 ( new_n446_, new_n445_, new_n381_ );
nand g309 ( new_n447_, new_n442_, N65, new_n444_ );
nand g310 ( new_n448_, new_n446_, new_n380_, new_n447_ );
nand g311 ( new_n449_, new_n446_, new_n447_ );
nand g312 ( new_n450_, new_n449_, keyIn_0_52 );
nand g313 ( N740, new_n450_, new_n448_ );
not g314 ( new_n452_, keyIn_0_53 );
not g315 ( new_n453_, N69 );
nand g316 ( new_n454_, new_n440_, new_n258_ );
nand g317 ( new_n455_, new_n454_, keyIn_0_41 );
not g318 ( new_n456_, keyIn_0_41 );
nand g319 ( new_n457_, new_n440_, new_n456_, new_n258_ );
nand g320 ( new_n458_, new_n455_, new_n457_ );
nand g321 ( new_n459_, new_n458_, new_n453_ );
nand g322 ( new_n460_, new_n455_, N69, new_n457_ );
nand g323 ( new_n461_, new_n459_, new_n452_, new_n460_ );
nand g324 ( new_n462_, new_n459_, new_n460_ );
nand g325 ( new_n463_, new_n462_, keyIn_0_53 );
nand g326 ( N741, new_n463_, new_n461_ );
not g327 ( new_n465_, keyIn_0_54 );
not g328 ( new_n466_, N73 );
nand g329 ( new_n467_, new_n440_, new_n292_ );
nand g330 ( new_n468_, new_n467_, keyIn_0_42 );
not g331 ( new_n469_, keyIn_0_42 );
nand g332 ( new_n470_, new_n440_, new_n469_, new_n292_ );
nand g333 ( new_n471_, new_n468_, new_n470_ );
nand g334 ( new_n472_, new_n471_, new_n466_ );
nand g335 ( new_n473_, new_n468_, N73, new_n470_ );
nand g336 ( new_n474_, new_n472_, new_n465_, new_n473_ );
nand g337 ( new_n475_, new_n472_, new_n473_ );
nand g338 ( new_n476_, new_n475_, keyIn_0_54 );
nand g339 ( N742, new_n476_, new_n474_ );
not g340 ( new_n478_, keyIn_0_55 );
not g341 ( new_n479_, N77 );
nand g342 ( new_n480_, new_n440_, new_n339_ );
nand g343 ( new_n481_, new_n480_, keyIn_0_43 );
not g344 ( new_n482_, keyIn_0_43 );
nand g345 ( new_n483_, new_n440_, new_n482_, new_n339_ );
nand g346 ( new_n484_, new_n481_, new_n483_ );
nand g347 ( new_n485_, new_n484_, new_n479_ );
nand g348 ( new_n486_, new_n481_, N77, new_n483_ );
nand g349 ( new_n487_, new_n485_, new_n478_, new_n486_ );
nand g350 ( new_n488_, new_n485_, new_n486_ );
nand g351 ( new_n489_, new_n488_, keyIn_0_55 );
nand g352 ( N743, new_n489_, new_n487_ );
not g353 ( new_n491_, N81 );
not g354 ( new_n492_, keyIn_0_38 );
nor g355 ( new_n493_, new_n433_, new_n303_, new_n328_ );
nand g356 ( new_n494_, new_n432_, new_n493_ );
nand g357 ( new_n495_, new_n494_, new_n492_ );
nand g358 ( new_n496_, new_n432_, keyIn_0_38, new_n493_ );
nand g359 ( new_n497_, new_n495_, new_n496_ );
nand g360 ( new_n498_, new_n497_, new_n224_ );
nand g361 ( new_n499_, new_n498_, keyIn_0_44 );
not g362 ( new_n500_, keyIn_0_44 );
nand g363 ( new_n501_, new_n497_, new_n500_, new_n224_ );
nand g364 ( new_n502_, new_n499_, new_n501_ );
nand g365 ( new_n503_, new_n502_, new_n491_ );
nand g366 ( new_n504_, new_n499_, N81, new_n501_ );
nand g367 ( new_n505_, new_n503_, keyIn_0_56, new_n504_ );
not g368 ( new_n506_, keyIn_0_56 );
nand g369 ( new_n507_, new_n503_, new_n504_ );
nand g370 ( new_n508_, new_n507_, new_n506_ );
nand g371 ( N744, new_n508_, new_n505_ );
not g372 ( new_n510_, keyIn_0_57 );
not g373 ( new_n511_, N85 );
nand g374 ( new_n512_, new_n497_, new_n258_ );
nand g375 ( new_n513_, new_n512_, keyIn_0_45 );
not g376 ( new_n514_, keyIn_0_45 );
nand g377 ( new_n515_, new_n497_, new_n514_, new_n258_ );
nand g378 ( new_n516_, new_n513_, new_n515_ );
nand g379 ( new_n517_, new_n516_, new_n511_ );
nand g380 ( new_n518_, new_n513_, N85, new_n515_ );
nand g381 ( new_n519_, new_n517_, new_n510_, new_n518_ );
nand g382 ( new_n520_, new_n517_, new_n518_ );
nand g383 ( new_n521_, new_n520_, keyIn_0_57 );
nand g384 ( N745, new_n521_, new_n519_ );
not g385 ( new_n523_, N89 );
nand g386 ( new_n524_, new_n497_, new_n292_ );
nand g387 ( new_n525_, new_n524_, keyIn_0_46 );
not g388 ( new_n526_, keyIn_0_46 );
nand g389 ( new_n527_, new_n497_, new_n526_, new_n292_ );
nand g390 ( new_n528_, new_n525_, new_n527_ );
nand g391 ( new_n529_, new_n528_, new_n523_ );
nand g392 ( new_n530_, new_n525_, N89, new_n527_ );
nand g393 ( new_n531_, new_n529_, keyIn_0_58, new_n530_ );
not g394 ( new_n532_, keyIn_0_58 );
nand g395 ( new_n533_, new_n529_, new_n530_ );
nand g396 ( new_n534_, new_n533_, new_n532_ );
nand g397 ( N746, new_n534_, new_n531_ );
not g398 ( new_n536_, keyIn_0_59 );
not g399 ( new_n537_, N93 );
nand g400 ( new_n538_, new_n497_, new_n339_ );
nand g401 ( new_n539_, new_n538_, keyIn_0_47 );
not g402 ( new_n540_, keyIn_0_47 );
nand g403 ( new_n541_, new_n497_, new_n540_, new_n339_ );
nand g404 ( new_n542_, new_n539_, new_n541_ );
nand g405 ( new_n543_, new_n542_, new_n537_ );
nand g406 ( new_n544_, new_n539_, N93, new_n541_ );
nand g407 ( new_n545_, new_n543_, new_n536_, new_n544_ );
nand g408 ( new_n546_, new_n543_, new_n544_ );
nand g409 ( new_n547_, new_n546_, keyIn_0_59 );
nand g410 ( N747, new_n547_, new_n545_ );
not g411 ( new_n549_, N97 );
nor g412 ( new_n550_, new_n434_, new_n151_, new_n316_ );
nand g413 ( new_n551_, new_n432_, new_n550_ );
nand g414 ( new_n552_, new_n551_, keyIn_0_39 );
not g415 ( new_n553_, keyIn_0_39 );
nand g416 ( new_n554_, new_n432_, new_n553_, new_n550_ );
nand g417 ( new_n555_, new_n552_, new_n554_ );
nand g418 ( new_n556_, new_n555_, new_n224_ );
nand g419 ( new_n557_, new_n556_, keyIn_0_48 );
not g420 ( new_n558_, keyIn_0_48 );
nand g421 ( new_n559_, new_n555_, new_n558_, new_n224_ );
nand g422 ( new_n560_, new_n557_, new_n559_ );
nand g423 ( new_n561_, new_n560_, new_n549_ );
nand g424 ( new_n562_, new_n557_, N97, new_n559_ );
nand g425 ( new_n563_, new_n561_, keyIn_0_60, new_n562_ );
not g426 ( new_n564_, keyIn_0_60 );
nand g427 ( new_n565_, new_n561_, new_n562_ );
nand g428 ( new_n566_, new_n565_, new_n564_ );
nand g429 ( N748, new_n566_, new_n563_ );
not g430 ( new_n568_, N101 );
nand g431 ( new_n569_, new_n555_, new_n258_ );
nand g432 ( new_n570_, new_n569_, keyIn_0_49 );
not g433 ( new_n571_, keyIn_0_49 );
nand g434 ( new_n572_, new_n555_, new_n571_, new_n258_ );
nand g435 ( new_n573_, new_n570_, new_n572_ );
nand g436 ( new_n574_, new_n573_, new_n568_ );
nand g437 ( new_n575_, new_n570_, N101, new_n572_ );
nand g438 ( new_n576_, new_n574_, keyIn_0_61, new_n575_ );
not g439 ( new_n577_, keyIn_0_61 );
nand g440 ( new_n578_, new_n574_, new_n575_ );
nand g441 ( new_n579_, new_n578_, new_n577_ );
nand g442 ( N749, new_n579_, new_n576_ );
not g443 ( new_n581_, N105 );
nand g444 ( new_n582_, new_n555_, new_n292_ );
nand g445 ( new_n583_, new_n582_, keyIn_0_50 );
not g446 ( new_n584_, keyIn_0_50 );
nand g447 ( new_n585_, new_n555_, new_n584_, new_n292_ );
nand g448 ( new_n586_, new_n583_, new_n585_ );
nand g449 ( new_n587_, new_n586_, new_n581_ );
nand g450 ( new_n588_, new_n583_, N105, new_n585_ );
nand g451 ( new_n589_, new_n587_, keyIn_0_62, new_n588_ );
not g452 ( new_n590_, keyIn_0_62 );
nand g453 ( new_n591_, new_n587_, new_n588_ );
nand g454 ( new_n592_, new_n591_, new_n590_ );
nand g455 ( N750, new_n592_, new_n589_ );
not g456 ( new_n594_, N109 );
nand g457 ( new_n595_, new_n555_, keyIn_0_51, new_n339_ );
not g458 ( new_n596_, keyIn_0_51 );
nand g459 ( new_n597_, new_n555_, new_n339_ );
nand g460 ( new_n598_, new_n597_, new_n596_ );
nand g461 ( new_n599_, new_n598_, new_n595_ );
nand g462 ( new_n600_, new_n599_, new_n594_ );
nand g463 ( new_n601_, new_n598_, N109, new_n595_ );
nand g464 ( new_n602_, new_n600_, new_n601_ );
nand g465 ( new_n603_, new_n602_, keyIn_0_63 );
not g466 ( new_n604_, keyIn_0_63 );
nand g467 ( new_n605_, new_n600_, new_n604_, new_n601_ );
nand g468 ( N751, new_n603_, new_n605_ );
nor g469 ( new_n607_, new_n319_, new_n328_ );
nand g470 ( new_n608_, new_n432_, new_n224_, new_n607_ );
xnor g471 ( N752, new_n608_, N113 );
nand g472 ( new_n610_, new_n432_, new_n258_, new_n607_ );
xnor g473 ( N753, new_n610_, N117 );
nand g474 ( new_n612_, new_n432_, new_n292_, new_n607_ );
xnor g475 ( N754, new_n612_, N121 );
nand g476 ( new_n614_, new_n432_, new_n339_, new_n607_ );
xnor g477 ( N755, new_n614_, N125 );
endmodule