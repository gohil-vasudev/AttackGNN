module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n595_, new_n614_, new_n445_, new_n699_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n421_, new_n720_, new_n620_, new_n368_, new_n738_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n566_, new_n641_, new_n339_, new_n365_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n246_, new_n682_, new_n679_, new_n266_, new_n667_, new_n367_, new_n542_, new_n548_, new_n669_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n637_, new_n451_, new_n489_, new_n424_, new_n602_, new_n695_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n642_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n735_, new_n500_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n427_, new_n532_, new_n472_, new_n393_, new_n418_, new_n292_, new_n626_, new_n716_, new_n701_, new_n257_, new_n481_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n272_, new_n282_, new_n634_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n655_, new_n630_, new_n385_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n683_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n318_, new_n622_, new_n629_, new_n702_, new_n321_, new_n715_, new_n443_, new_n324_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n498_, new_n492_, new_n496_, new_n650_, new_n708_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n506_, new_n680_, new_n256_, new_n452_, new_n381_, new_n656_, new_n388_, new_n508_, new_n714_, new_n483_, new_n394_, new_n299_, new_n657_, new_n652_, new_n314_, new_n582_, new_n363_, new_n441_, new_n477_, new_n664_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n541_, new_n458_, new_n447_, new_n267_, new_n473_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n488_, new_n524_, new_n705_, new_n277_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n438_, new_n632_, new_n671_, new_n528_, new_n572_, new_n436_, new_n397_, new_n729_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n437_, new_n295_, new_n359_, new_n628_, new_n409_, new_n457_, new_n553_, new_n668_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n688_, new_n384_, new_n410_, new_n543_, new_n371_, new_n509_, new_n454_, new_n296_, new_n661_, new_n308_, new_n633_, new_n232_, new_n258_, new_n724_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n654_, new_n713_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n310_, new_n275_, new_n352_, new_n575_, new_n562_, new_n578_, new_n525_, new_n493_, new_n547_, new_n264_, new_n665_, new_n379_, new_n719_, new_n273_, new_n586_, new_n270_, new_n570_, new_n598_, new_n520_, new_n253_, new_n717_, new_n403_, new_n475_, new_n237_, new_n557_, new_n260_, new_n300_, new_n411_, new_n673_, new_n407_, new_n666_, new_n480_, new_n625_, new_n730_, new_n736_, new_n513_, new_n592_, new_n726_, new_n558_, new_n231_, new_n313_, new_n382_, new_n583_, new_n239_, new_n617_, new_n718_, new_n522_, new_n588_, new_n428_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n415_, new_n537_, new_n243_, new_n450_, new_n345_, new_n298_, new_n499_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n737_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n337_, new_n446_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n519_, new_n563_, new_n440_, new_n733_, new_n531_, new_n593_, new_n252_, new_n585_, new_n312_, new_n535_, new_n372_, new_n725_, new_n242_, new_n503_, new_n527_, new_n307_, new_n597_, new_n408_, new_n470_, new_n651_, new_n433_, new_n435_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n278_, new_n304_, new_n523_, new_n638_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n711_, new_n644_, new_n731_, new_n599_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n431_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n653_, new_n336_, new_n377_, new_n539_, new_n727_, new_n375_, new_n294_, new_n627_, new_n704_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n490_, new_n560_, new_n358_, new_n348_, new_n610_, new_n322_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n226_, new_n697_, new_n709_, new_n373_, new_n540_, new_n434_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n551_, new_n279_, new_n455_, new_n618_, new_n521_, new_n406_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n573_, new_n405_;

and g000 ( N388, N29, N42, N75 );
and g001 ( N389, N29, N36, N80 );
nand g002 ( new_n217_, N29, N36, N42 );
xnor g003 ( N390, new_n217_, keyIn_0_6 );
and g004 ( N391, N85, N86 );
and g005 ( new_n220_, N1, N8 );
and g006 ( N418, new_n220_, N13, N17 );
xnor g007 ( new_n222_, new_n217_, keyIn_0_0 );
and g008 ( new_n223_, N1, N13, N17, N26 );
nand g009 ( N419, new_n222_, new_n223_ );
nand g010 ( N420, N59, N75, N80 );
nand g011 ( new_n226_, N36, N59, N80 );
xnor g012 ( new_n227_, new_n226_, keyIn_0_8 );
xor g013 ( N421, new_n227_, keyIn_0_19 );
nand g014 ( new_n229_, N36, N42, N59 );
xor g015 ( N422, new_n229_, keyIn_0_9 );
not g016 ( new_n231_, N90 );
nor g017 ( new_n232_, N87, N88 );
nor g018 ( new_n233_, new_n232_, new_n231_ );
xor g019 ( N423, new_n233_, keyIn_0_20 );
not g020 ( new_n235_, new_n222_ );
nand g021 ( N446, new_n235_, new_n223_ );
not g022 ( new_n237_, keyIn_0_1 );
nand g023 ( new_n238_, N1, N26, N51 );
nand g024 ( new_n239_, new_n238_, new_n237_ );
nand g025 ( new_n240_, keyIn_0_1, N1, N26, N51 );
nand g026 ( N447, new_n239_, new_n240_ );
nand g027 ( new_n242_, new_n220_, N13, N55 );
xor g028 ( new_n243_, new_n242_, keyIn_0_3 );
nand g029 ( new_n244_, N29, N68 );
xor g030 ( new_n245_, new_n244_, keyIn_0_4 );
nand g031 ( new_n246_, new_n243_, new_n245_ );
xor g032 ( N448, new_n246_, keyIn_0_27 );
nand g033 ( new_n248_, N59, N68, N74 );
xor g034 ( new_n249_, new_n248_, keyIn_0_5 );
nand g035 ( new_n250_, new_n243_, new_n249_ );
xnor g036 ( N449, new_n250_, keyIn_0_28 );
not g037 ( new_n252_, N89 );
nor g038 ( new_n253_, new_n232_, new_n252_ );
xor g039 ( N450, new_n253_, keyIn_0_29 );
not g040 ( new_n255_, keyIn_0_63 );
not g041 ( new_n256_, N130 );
nand g042 ( new_n257_, N101, N106 );
nand g043 ( new_n258_, new_n257_, keyIn_0_10 );
or g044 ( new_n259_, N101, N106 );
nand g045 ( new_n260_, new_n259_, keyIn_0_11 );
or g046 ( new_n261_, new_n257_, keyIn_0_10 );
or g047 ( new_n262_, new_n259_, keyIn_0_11 );
nand g048 ( new_n263_, new_n262_, new_n258_, new_n260_, new_n261_ );
xor g049 ( new_n264_, new_n263_, keyIn_0_22 );
xnor g050 ( new_n265_, N91, N96 );
xnor g051 ( new_n266_, new_n265_, keyIn_0_21 );
or g052 ( new_n267_, new_n264_, new_n266_ );
nand g053 ( new_n268_, new_n267_, keyIn_0_30 );
nand g054 ( new_n269_, new_n264_, new_n266_ );
or g055 ( new_n270_, new_n267_, keyIn_0_30 );
nand g056 ( new_n271_, new_n270_, new_n268_, new_n269_ );
and g057 ( new_n272_, new_n271_, new_n256_ );
or g058 ( new_n273_, new_n272_, keyIn_0_45 );
or g059 ( new_n274_, new_n271_, new_n256_ );
or g060 ( new_n275_, new_n274_, keyIn_0_44 );
nand g061 ( new_n276_, new_n272_, keyIn_0_45 );
nand g062 ( new_n277_, new_n274_, keyIn_0_44 );
nand g063 ( new_n278_, new_n275_, new_n273_, new_n276_, new_n277_ );
nand g064 ( new_n279_, new_n278_, keyIn_0_57 );
xnor g065 ( new_n280_, N111, N116 );
xnor g066 ( new_n281_, new_n280_, keyIn_0_23 );
not g067 ( new_n282_, N121 );
not g068 ( new_n283_, N126 );
nand g069 ( new_n284_, new_n282_, new_n283_ );
nor g070 ( new_n285_, new_n284_, keyIn_0_12 );
and g071 ( new_n286_, new_n284_, keyIn_0_12 );
nor g072 ( new_n287_, new_n282_, new_n283_ );
nor g073 ( new_n288_, new_n286_, new_n285_, keyIn_0_31, new_n287_ );
xnor g074 ( new_n289_, new_n288_, new_n281_ );
nor g075 ( new_n290_, new_n289_, N135 );
xnor g076 ( new_n291_, new_n290_, keyIn_0_46 );
nand g077 ( new_n292_, new_n289_, N135 );
nand g078 ( new_n293_, new_n291_, new_n292_ );
xnor g079 ( new_n294_, new_n293_, keyIn_0_53 );
or g080 ( new_n295_, new_n278_, keyIn_0_57 );
nand g081 ( new_n296_, new_n295_, new_n279_, new_n294_ );
and g082 ( new_n297_, new_n296_, new_n255_ );
not g083 ( new_n298_, new_n294_ );
and g084 ( new_n299_, new_n278_, new_n298_ );
nor g085 ( new_n300_, new_n296_, new_n255_ );
nor g086 ( N767, new_n297_, new_n300_, new_n299_ );
not g087 ( new_n302_, keyIn_0_64 );
not g088 ( new_n303_, keyIn_0_51 );
not g089 ( new_n304_, N207 );
xor g090 ( new_n305_, N183, N189 );
xnor g091 ( new_n306_, new_n305_, keyIn_0_25 );
xnor g092 ( new_n307_, N195, N201 );
xnor g093 ( new_n308_, new_n307_, keyIn_0_26 );
xnor g094 ( new_n309_, new_n306_, new_n308_ );
nor g095 ( new_n310_, new_n309_, new_n304_ );
or g096 ( new_n311_, new_n310_, new_n303_ );
nand g097 ( new_n312_, new_n309_, new_n304_ );
nand g098 ( new_n313_, new_n310_, new_n303_ );
nand g099 ( new_n314_, new_n311_, new_n312_, new_n313_ );
nand g100 ( new_n315_, new_n314_, keyIn_0_62 );
nand g101 ( new_n316_, N159, N165 );
or g102 ( new_n317_, new_n316_, keyIn_0_15 );
or g103 ( new_n318_, N159, N165 );
nand g104 ( new_n319_, new_n316_, keyIn_0_15 );
nand g105 ( new_n320_, new_n317_, new_n318_, new_n319_ );
xnor g106 ( new_n321_, N171, N177 );
xnor g107 ( new_n322_, new_n320_, new_n321_ );
xnor g108 ( new_n323_, new_n322_, new_n256_ );
xor g109 ( new_n324_, new_n323_, keyIn_0_61 );
or g110 ( new_n325_, new_n314_, keyIn_0_62 );
nand g111 ( new_n326_, new_n325_, new_n315_, new_n324_ );
nor g112 ( new_n327_, new_n326_, new_n302_ );
and g113 ( new_n328_, new_n326_, new_n302_ );
and g114 ( new_n329_, new_n314_, new_n323_ );
nor g115 ( N768, new_n328_, new_n327_, new_n329_ );
not g116 ( new_n331_, keyIn_0_50 );
not g117 ( new_n332_, keyIn_0_36 );
not g118 ( new_n333_, keyIn_0_2 );
nand g119 ( new_n334_, new_n220_, new_n333_, N17, N51 );
nand g120 ( new_n335_, N1, N8, N17, N51 );
nand g121 ( new_n336_, new_n335_, keyIn_0_2 );
nand g122 ( new_n337_, new_n334_, new_n336_ );
not g123 ( new_n338_, keyIn_0_7 );
nand g124 ( new_n339_, N42, N59, N75 );
xnor g125 ( new_n340_, new_n339_, new_n338_ );
nand g126 ( new_n341_, new_n337_, new_n340_ );
nand g127 ( new_n342_, N17, N42 );
nand g128 ( new_n343_, N59, N156 );
nor g129 ( new_n344_, N17, N42 );
nor g130 ( new_n345_, new_n344_, new_n343_ );
nand g131 ( new_n346_, N447, new_n342_, new_n345_ );
nand g132 ( new_n347_, new_n341_, new_n332_, new_n346_ );
nand g133 ( new_n348_, new_n341_, new_n346_ );
nand g134 ( new_n349_, new_n348_, keyIn_0_36 );
nand g135 ( new_n350_, new_n349_, N126, new_n347_ );
nand g136 ( new_n351_, new_n350_, new_n331_ );
nand g137 ( new_n352_, new_n349_, keyIn_0_50, N126, new_n347_ );
nand g138 ( new_n353_, new_n351_, new_n352_ );
not g139 ( new_n354_, keyIn_0_35 );
nand g140 ( new_n355_, new_n343_, keyIn_0_14 );
not g141 ( new_n356_, keyIn_0_14 );
nand g142 ( new_n357_, new_n356_, N59, N156 );
nand g143 ( new_n358_, new_n355_, new_n357_ );
nand g144 ( new_n359_, N447, N17, new_n358_ );
nand g145 ( new_n360_, new_n359_, new_n354_ );
nand g146 ( new_n361_, N447, keyIn_0_35, new_n358_, N17 );
nand g147 ( new_n362_, new_n360_, new_n361_ );
nand g148 ( new_n363_, new_n362_, N1 );
nand g149 ( new_n364_, new_n363_, N153 );
nand g150 ( new_n365_, new_n353_, keyIn_0_56, new_n364_ );
not g151 ( new_n366_, keyIn_0_56 );
nand g152 ( new_n367_, new_n353_, new_n364_ );
nand g153 ( new_n368_, new_n367_, new_n366_ );
nand g154 ( new_n369_, N447, N55 );
xor g155 ( new_n370_, keyIn_0_24, N268 );
nand g156 ( new_n371_, N29, N75, N80 );
nor g157 ( new_n372_, new_n369_, new_n370_, new_n371_ );
not g158 ( new_n373_, new_n372_ );
nand g159 ( new_n374_, new_n368_, new_n365_, new_n373_ );
nand g160 ( new_n375_, new_n374_, N201 );
not g161 ( new_n376_, N201 );
nand g162 ( new_n377_, new_n368_, new_n376_, new_n365_, new_n373_ );
nand g163 ( new_n378_, new_n375_, new_n377_ );
xnor g164 ( new_n379_, new_n378_, keyIn_0_82 );
and g165 ( new_n380_, new_n379_, N261 );
nand g166 ( new_n381_, new_n380_, keyIn_0_93 );
or g167 ( new_n382_, new_n380_, keyIn_0_93 );
or g168 ( new_n383_, new_n379_, N261 );
nand g169 ( new_n384_, new_n382_, N219, new_n381_, new_n383_ );
nand g170 ( new_n385_, new_n379_, N228 );
not g171 ( new_n386_, N237 );
nor g172 ( new_n387_, new_n375_, new_n386_ );
and g173 ( new_n388_, new_n374_, N246 );
and g174 ( new_n389_, N42, N72, N73 );
nand g175 ( new_n390_, new_n243_, N59, N68, new_n389_ );
xor g176 ( new_n391_, new_n390_, keyIn_0_33 );
nand g177 ( new_n392_, new_n391_, N201 );
and g178 ( new_n393_, N255, N267 );
nand g179 ( new_n394_, new_n393_, keyIn_0_18 );
or g180 ( new_n395_, new_n393_, keyIn_0_18 );
nand g181 ( new_n396_, N121, N210 );
nand g182 ( new_n397_, new_n392_, new_n394_, new_n395_, new_n396_ );
nor g183 ( new_n398_, new_n387_, new_n388_, new_n397_ );
nand g184 ( N850, new_n384_, new_n385_, new_n398_ );
nand g185 ( new_n400_, new_n363_, N143 );
xnor g186 ( new_n401_, new_n372_, keyIn_0_42 );
nand g187 ( new_n402_, new_n349_, new_n347_ );
not g188 ( new_n403_, new_n402_ );
nand g189 ( new_n404_, new_n403_, N111 );
nand g190 ( new_n405_, new_n404_, new_n400_, new_n401_ );
nand g191 ( new_n406_, new_n405_, N183 );
or g192 ( new_n407_, new_n405_, N183 );
nand g193 ( new_n408_, new_n407_, new_n406_ );
xnor g194 ( new_n409_, new_n408_, keyIn_0_79 );
not g195 ( new_n410_, N189 );
not g196 ( new_n411_, keyIn_0_60 );
nand g197 ( new_n412_, new_n363_, N146 );
nand g198 ( new_n413_, new_n412_, keyIn_0_48 );
not g199 ( new_n414_, keyIn_0_48 );
nand g200 ( new_n415_, new_n363_, new_n414_, N146 );
nand g201 ( new_n416_, new_n413_, new_n415_ );
and g202 ( new_n417_, new_n349_, N116, new_n347_ );
nor g203 ( new_n418_, new_n417_, new_n372_ );
nand g204 ( new_n419_, new_n416_, new_n418_ );
nand g205 ( new_n420_, new_n419_, new_n411_ );
nand g206 ( new_n421_, new_n416_, new_n418_, keyIn_0_60 );
nand g207 ( new_n422_, new_n420_, new_n410_, new_n421_ );
nand g208 ( new_n423_, new_n422_, keyIn_0_70 );
not g209 ( new_n424_, keyIn_0_70 );
nand g210 ( new_n425_, new_n420_, new_n424_, new_n410_, new_n421_ );
nand g211 ( new_n426_, new_n423_, new_n425_ );
not g212 ( new_n427_, keyIn_0_72 );
not g213 ( new_n428_, N195 );
not g214 ( new_n429_, keyIn_0_49 );
nand g215 ( new_n430_, new_n363_, N149 );
nand g216 ( new_n431_, new_n430_, new_n429_ );
nand g217 ( new_n432_, new_n363_, keyIn_0_49, N149 );
nand g218 ( new_n433_, new_n431_, new_n432_ );
nand g219 ( new_n434_, new_n349_, N121, new_n347_ );
xnor g220 ( new_n435_, new_n372_, keyIn_0_43 );
and g221 ( new_n436_, new_n435_, new_n434_ );
nand g222 ( new_n437_, new_n433_, new_n428_, new_n436_ );
nand g223 ( new_n438_, new_n437_, new_n427_ );
nand g224 ( new_n439_, new_n433_, keyIn_0_72, new_n428_, new_n436_ );
nand g225 ( new_n440_, new_n438_, new_n439_ );
and g226 ( new_n441_, new_n440_, N201, new_n374_ );
nand g227 ( new_n442_, new_n426_, new_n441_, keyIn_0_95 );
not g228 ( new_n443_, keyIn_0_90 );
nand g229 ( new_n444_, new_n420_, new_n421_ );
nand g230 ( new_n445_, new_n444_, N189 );
nand g231 ( new_n446_, new_n445_, new_n443_ );
nand g232 ( new_n447_, new_n444_, keyIn_0_90, N189 );
nand g233 ( new_n448_, new_n446_, new_n447_ );
and g234 ( new_n449_, new_n442_, new_n448_ );
not g235 ( new_n450_, keyIn_0_95 );
nand g236 ( new_n451_, new_n426_, new_n441_ );
nand g237 ( new_n452_, new_n451_, new_n450_ );
not g238 ( new_n453_, keyIn_0_80 );
nand g239 ( new_n454_, new_n433_, new_n436_ );
nand g240 ( new_n455_, new_n454_, N195 );
nand g241 ( new_n456_, new_n455_, keyIn_0_71 );
not g242 ( new_n457_, keyIn_0_71 );
nand g243 ( new_n458_, new_n454_, new_n457_, N195 );
nand g244 ( new_n459_, new_n456_, new_n458_ );
nand g245 ( new_n460_, new_n459_, new_n453_ );
nand g246 ( new_n461_, new_n456_, keyIn_0_80, new_n458_ );
nand g247 ( new_n462_, new_n460_, new_n461_ );
nand g248 ( new_n463_, new_n440_, new_n377_, N261 );
nand g249 ( new_n464_, new_n462_, new_n463_ );
nand g250 ( new_n465_, new_n464_, new_n426_ );
nand g251 ( new_n466_, new_n449_, new_n465_, new_n452_ );
xnor g252 ( new_n467_, new_n466_, new_n409_ );
or g253 ( new_n468_, new_n467_, keyIn_0_103 );
nand g254 ( new_n469_, new_n467_, keyIn_0_103 );
nand g255 ( new_n470_, new_n468_, N219, new_n469_ );
xnor g256 ( new_n471_, new_n470_, keyIn_0_106 );
nand g257 ( new_n472_, new_n409_, N228 );
or g258 ( new_n473_, new_n472_, keyIn_0_89 );
xnor g259 ( new_n474_, new_n406_, keyIn_0_78 );
nand g260 ( new_n475_, new_n474_, N237 );
nand g261 ( new_n476_, new_n472_, keyIn_0_89 );
nand g262 ( new_n477_, new_n473_, new_n475_, new_n476_ );
or g263 ( new_n478_, new_n477_, keyIn_0_98 );
nand g264 ( new_n479_, new_n477_, keyIn_0_98 );
nand g265 ( new_n480_, new_n405_, N246 );
nand g266 ( new_n481_, N106, N210 );
nand g267 ( new_n482_, new_n391_, N183 );
and g268 ( new_n483_, new_n480_, new_n481_, new_n482_ );
nand g269 ( new_n484_, new_n471_, new_n478_, new_n479_, new_n483_ );
xor g270 ( N863, new_n484_, keyIn_0_120 );
and g271 ( new_n486_, new_n426_, new_n445_ );
xor g272 ( new_n487_, new_n462_, keyIn_0_91 );
not g273 ( new_n488_, new_n463_ );
nand g274 ( new_n489_, new_n488_, keyIn_0_83 );
xor g275 ( new_n490_, new_n441_, keyIn_0_94 );
or g276 ( new_n491_, new_n488_, keyIn_0_83 );
nand g277 ( new_n492_, new_n487_, new_n489_, new_n490_, new_n491_ );
xnor g278 ( new_n493_, new_n492_, keyIn_0_99 );
nand g279 ( new_n494_, new_n493_, new_n486_ );
or g280 ( new_n495_, new_n493_, new_n486_ );
nand g281 ( new_n496_, new_n495_, N219, new_n494_ );
nand g282 ( new_n497_, N111, N210 );
nand g283 ( new_n498_, new_n496_, new_n497_ );
nand g284 ( new_n499_, new_n498_, keyIn_0_111 );
or g285 ( new_n500_, new_n498_, keyIn_0_111 );
nand g286 ( new_n501_, new_n486_, N228 );
nand g287 ( new_n502_, new_n444_, N189, N237 );
nand g288 ( new_n503_, new_n444_, N246 );
nand g289 ( new_n504_, new_n391_, N189 );
nand g290 ( new_n505_, N255, N259 );
and g291 ( new_n506_, new_n502_, new_n503_, new_n504_, new_n505_ );
nand g292 ( N864, new_n500_, new_n499_, new_n501_, new_n506_ );
nand g293 ( new_n508_, new_n460_, N237, new_n461_ );
not g294 ( new_n509_, N228 );
nand g295 ( new_n510_, new_n459_, new_n440_ );
nor g296 ( new_n511_, new_n510_, new_n509_ );
xnor g297 ( new_n512_, new_n511_, keyIn_0_92 );
nand g298 ( new_n513_, new_n512_, new_n508_ );
xor g299 ( new_n514_, new_n513_, keyIn_0_100 );
nand g300 ( new_n515_, new_n377_, N261 );
nand g301 ( new_n516_, new_n515_, new_n375_ );
xor g302 ( new_n517_, new_n516_, new_n510_ );
xnor g303 ( new_n518_, new_n517_, keyIn_0_104 );
nand g304 ( new_n519_, new_n518_, N219 );
nand g305 ( new_n520_, new_n454_, N246 );
nand g306 ( new_n521_, N255, N260 );
and g307 ( new_n522_, new_n520_, new_n521_ );
and g308 ( new_n523_, new_n522_, keyIn_0_81 );
nor g309 ( new_n524_, new_n522_, keyIn_0_81 );
and g310 ( new_n525_, new_n391_, N195 );
nand g311 ( new_n526_, N116, N210 );
xor g312 ( new_n527_, new_n526_, keyIn_0_17 );
nor g313 ( new_n528_, new_n523_, new_n524_, new_n525_, new_n527_ );
nand g314 ( new_n529_, new_n514_, new_n519_, new_n528_ );
xor g315 ( N865, new_n529_, keyIn_0_117 );
nand g316 ( new_n531_, N447, N55, new_n358_ );
xnor g317 ( new_n532_, new_n531_, keyIn_0_34 );
not g318 ( new_n533_, new_n532_ );
nand g319 ( new_n534_, new_n533_, N146 );
xor g320 ( new_n535_, new_n534_, keyIn_0_39 );
nand g321 ( new_n536_, new_n403_, N96 );
nand g322 ( new_n537_, N51, N138 );
nor g323 ( new_n538_, new_n371_, N268 );
nand g324 ( new_n539_, N447, N17, new_n538_ );
xnor g325 ( new_n540_, new_n539_, keyIn_0_40 );
nand g326 ( new_n541_, new_n535_, new_n536_, new_n537_, new_n540_ );
nor g327 ( new_n542_, new_n541_, N165 );
xnor g328 ( new_n543_, new_n542_, keyIn_0_66 );
nand g329 ( new_n544_, new_n403_, N101 );
nand g330 ( new_n545_, N17, N138 );
nand g331 ( new_n546_, new_n544_, new_n545_ );
xor g332 ( new_n547_, new_n546_, keyIn_0_55 );
nand g333 ( new_n548_, new_n533_, N149 );
or g334 ( new_n549_, new_n548_, keyIn_0_41 );
nand g335 ( new_n550_, new_n548_, keyIn_0_41 );
nand g336 ( new_n551_, new_n547_, new_n539_, new_n549_, new_n550_ );
nor g337 ( new_n552_, new_n551_, N171 );
xor g338 ( new_n553_, new_n552_, keyIn_0_68 );
not g339 ( new_n554_, new_n474_ );
not g340 ( new_n555_, keyIn_0_101 );
nand g341 ( new_n556_, new_n466_, new_n407_ );
nand g342 ( new_n557_, new_n556_, new_n555_ );
nand g343 ( new_n558_, new_n466_, keyIn_0_101, new_n407_ );
nand g344 ( new_n559_, new_n557_, new_n558_ );
nand g345 ( new_n560_, new_n559_, new_n554_ );
nand g346 ( new_n561_, new_n560_, keyIn_0_102 );
not g347 ( new_n562_, keyIn_0_102 );
nand g348 ( new_n563_, new_n559_, new_n562_, new_n554_ );
nand g349 ( new_n564_, new_n561_, new_n563_ );
nand g350 ( new_n565_, new_n533_, N153 );
nand g351 ( new_n566_, new_n565_, new_n539_ );
nand g352 ( new_n567_, new_n566_, keyIn_0_47 );
or g353 ( new_n568_, new_n566_, keyIn_0_47 );
nand g354 ( new_n569_, new_n403_, N106 );
nand g355 ( new_n570_, N138, N152 );
xor g356 ( new_n571_, new_n570_, keyIn_0_13 );
nand g357 ( new_n572_, new_n568_, new_n567_, new_n569_, new_n571_ );
xnor g358 ( new_n573_, new_n572_, keyIn_0_59 );
nor g359 ( new_n574_, new_n573_, N177 );
xnor g360 ( new_n575_, new_n574_, keyIn_0_69 );
nand g361 ( new_n576_, new_n564_, new_n543_, new_n553_, new_n575_ );
nand g362 ( new_n577_, new_n573_, N177 );
not g363 ( new_n578_, new_n577_ );
nand g364 ( new_n579_, new_n553_, new_n578_ );
nand g365 ( new_n580_, new_n551_, N171 );
xnor g366 ( new_n581_, new_n580_, keyIn_0_67 );
nand g367 ( new_n582_, new_n579_, new_n581_ );
nand g368 ( new_n583_, new_n582_, new_n543_ );
nand g369 ( new_n584_, new_n541_, N165 );
and g370 ( new_n585_, new_n583_, new_n584_ );
nand g371 ( new_n586_, new_n576_, new_n585_ );
nand g372 ( new_n587_, new_n403_, N91 );
nand g373 ( new_n588_, N8, N138 );
nand g374 ( new_n589_, new_n587_, new_n588_ );
xor g375 ( new_n590_, new_n589_, keyIn_0_54 );
nand g376 ( new_n591_, new_n533_, keyIn_0_37, N143 );
xnor g377 ( new_n592_, new_n539_, keyIn_0_38 );
not g378 ( new_n593_, keyIn_0_37 );
nand g379 ( new_n594_, new_n533_, N143 );
nand g380 ( new_n595_, new_n594_, new_n593_ );
nand g381 ( new_n596_, new_n590_, new_n591_, new_n592_, new_n595_ );
xor g382 ( new_n597_, new_n596_, keyIn_0_58 );
nor g383 ( new_n598_, new_n597_, N159 );
xor g384 ( new_n599_, new_n598_, keyIn_0_65 );
nand g385 ( new_n600_, new_n586_, new_n599_ );
xnor g386 ( new_n601_, new_n600_, keyIn_0_114 );
nand g387 ( new_n602_, new_n597_, N159 );
xnor g388 ( new_n603_, new_n602_, keyIn_0_73 );
nand g389 ( new_n604_, new_n601_, new_n603_ );
xnor g390 ( N866, new_n604_, keyIn_0_118 );
nand g391 ( new_n606_, new_n575_, new_n577_ );
not g392 ( new_n607_, new_n606_ );
nor g393 ( new_n608_, new_n564_, new_n607_ );
nand g394 ( new_n609_, new_n608_, keyIn_0_105 );
or g395 ( new_n610_, new_n608_, keyIn_0_105 );
nand g396 ( new_n611_, new_n564_, new_n607_ );
nand g397 ( new_n612_, new_n610_, new_n609_, new_n611_ );
xnor g398 ( new_n613_, new_n612_, keyIn_0_110 );
nand g399 ( new_n614_, new_n613_, N219 );
nand g400 ( new_n615_, new_n607_, N228 );
nand g401 ( new_n616_, new_n578_, N237 );
nand g402 ( new_n617_, new_n573_, N246 );
nand g403 ( new_n618_, new_n391_, N177 );
xnor g404 ( new_n619_, new_n618_, keyIn_0_52 );
nand g405 ( new_n620_, N101, N210 );
and g406 ( new_n621_, new_n616_, new_n617_, new_n619_, new_n620_ );
nand g407 ( new_n622_, new_n614_, new_n615_, new_n621_ );
xnor g408 ( N874, new_n622_, keyIn_0_123 );
not g409 ( new_n624_, keyIn_0_125 );
not g410 ( new_n625_, keyIn_0_112 );
nand g411 ( new_n626_, new_n599_, new_n602_ );
xor g412 ( new_n627_, new_n626_, keyIn_0_74 );
nand g413 ( new_n628_, new_n576_, new_n627_, new_n625_, new_n585_ );
nand g414 ( new_n629_, new_n576_, new_n585_, new_n627_ );
nand g415 ( new_n630_, new_n629_, keyIn_0_112 );
not g416 ( new_n631_, new_n627_ );
nand g417 ( new_n632_, new_n586_, new_n631_ );
nand g418 ( new_n633_, new_n630_, new_n628_, new_n632_ );
nand g419 ( new_n634_, new_n633_, keyIn_0_115 );
not g420 ( new_n635_, keyIn_0_115 );
nand g421 ( new_n636_, new_n630_, new_n632_, new_n635_, new_n628_ );
nand g422 ( new_n637_, new_n634_, new_n636_ );
nand g423 ( new_n638_, new_n637_, N219 );
nand g424 ( new_n639_, new_n370_, N210 );
xor g425 ( new_n640_, new_n639_, keyIn_0_32 );
nand g426 ( new_n641_, new_n638_, new_n640_ );
nand g427 ( new_n642_, new_n641_, keyIn_0_121 );
not g428 ( new_n643_, keyIn_0_121 );
nand g429 ( new_n644_, new_n638_, new_n643_, new_n640_ );
nand g430 ( new_n645_, new_n642_, new_n644_ );
nor g431 ( new_n646_, new_n627_, new_n509_ );
nor g432 ( new_n647_, new_n603_, new_n386_ );
not g433 ( new_n648_, new_n647_ );
nor g434 ( new_n649_, new_n648_, keyIn_0_84 );
nand g435 ( new_n650_, new_n648_, keyIn_0_84 );
nand g436 ( new_n651_, new_n597_, N246 );
nand g437 ( new_n652_, new_n391_, N159 );
nand g438 ( new_n653_, new_n650_, new_n651_, new_n652_ );
nor g439 ( new_n654_, new_n646_, new_n649_, new_n653_ );
nand g440 ( new_n655_, new_n645_, new_n654_ );
nand g441 ( new_n656_, new_n655_, keyIn_0_124 );
not g442 ( new_n657_, keyIn_0_124 );
nand g443 ( new_n658_, new_n645_, new_n657_, new_n654_ );
nand g444 ( new_n659_, new_n656_, new_n658_ );
nand g445 ( new_n660_, new_n659_, new_n624_ );
nand g446 ( new_n661_, new_n656_, keyIn_0_125, new_n658_ );
nand g447 ( N878, new_n660_, new_n661_ );
not g448 ( new_n663_, keyIn_0_126 );
nand g449 ( new_n664_, new_n543_, new_n584_ );
not g450 ( new_n665_, keyIn_0_108 );
not g451 ( new_n666_, keyIn_0_107 );
and g452 ( new_n667_, new_n564_, new_n553_, new_n575_ );
or g453 ( new_n668_, new_n667_, new_n666_ );
nand g454 ( new_n669_, new_n667_, new_n666_ );
xnor g455 ( new_n670_, new_n579_, keyIn_0_96 );
xor g456 ( new_n671_, new_n581_, keyIn_0_86 );
nand g457 ( new_n672_, new_n668_, new_n669_, new_n670_, new_n671_ );
xnor g458 ( new_n673_, new_n672_, new_n665_ );
nand g459 ( new_n674_, new_n673_, new_n664_ );
or g460 ( new_n675_, new_n673_, new_n664_ );
nand g461 ( new_n676_, new_n675_, N219, new_n674_ );
or g462 ( new_n677_, new_n676_, keyIn_0_119 );
nand g463 ( new_n678_, new_n676_, keyIn_0_119 );
nor g464 ( new_n679_, new_n664_, new_n509_ );
not g465 ( new_n680_, new_n679_ );
nor g466 ( new_n681_, new_n680_, keyIn_0_85 );
and g467 ( new_n682_, new_n680_, keyIn_0_85 );
nand g468 ( new_n683_, new_n541_, N246 );
nand g469 ( new_n684_, new_n391_, N165 );
and g470 ( new_n685_, new_n683_, new_n684_ );
nand g471 ( new_n686_, new_n685_, keyIn_0_75 );
or g472 ( new_n687_, new_n685_, keyIn_0_75 );
nand g473 ( new_n688_, new_n541_, N165, N237 );
nand g474 ( new_n689_, N91, N210 );
xor g475 ( new_n690_, new_n689_, keyIn_0_16 );
nand g476 ( new_n691_, new_n687_, new_n686_, new_n688_, new_n690_ );
nor g477 ( new_n692_, new_n682_, new_n681_, new_n691_ );
nand g478 ( new_n693_, new_n677_, new_n678_, new_n692_ );
nand g479 ( new_n694_, new_n693_, new_n663_ );
nand g480 ( new_n695_, new_n677_, keyIn_0_126, new_n678_, new_n692_ );
nand g481 ( N879, new_n694_, new_n695_ );
not g482 ( new_n697_, keyIn_0_122 );
nand g483 ( new_n698_, new_n553_, new_n581_ );
xnor g484 ( new_n699_, new_n698_, keyIn_0_76 );
not g485 ( new_n700_, new_n699_ );
nand g486 ( new_n701_, new_n564_, new_n575_ );
xnor g487 ( new_n702_, new_n577_, keyIn_0_88 );
nand g488 ( new_n703_, new_n701_, new_n702_ );
nand g489 ( new_n704_, new_n703_, keyIn_0_109 );
not g490 ( new_n705_, keyIn_0_109 );
nand g491 ( new_n706_, new_n701_, new_n705_, new_n702_ );
nand g492 ( new_n707_, new_n704_, keyIn_0_113, new_n700_, new_n706_ );
not g493 ( new_n708_, keyIn_0_113 );
nand g494 ( new_n709_, new_n704_, new_n700_, new_n706_ );
nand g495 ( new_n710_, new_n709_, new_n708_ );
nand g496 ( new_n711_, new_n710_, new_n707_ );
nand g497 ( new_n712_, new_n704_, new_n706_ );
nand g498 ( new_n713_, new_n712_, new_n699_ );
nand g499 ( new_n714_, new_n711_, new_n713_ );
nand g500 ( new_n715_, new_n714_, keyIn_0_116 );
not g501 ( new_n716_, keyIn_0_116 );
nand g502 ( new_n717_, new_n711_, new_n716_, new_n713_ );
nand g503 ( new_n718_, new_n715_, new_n717_ );
nand g504 ( new_n719_, new_n718_, N219 );
nand g505 ( new_n720_, N96, N210 );
nand g506 ( new_n721_, new_n719_, new_n720_ );
nand g507 ( new_n722_, new_n721_, new_n697_ );
nand g508 ( new_n723_, new_n719_, keyIn_0_122, new_n720_ );
nand g509 ( new_n724_, new_n699_, N228 );
xnor g510 ( new_n725_, new_n724_, keyIn_0_87 );
or g511 ( new_n726_, new_n581_, new_n386_ );
nand g512 ( new_n727_, new_n725_, new_n726_ );
and g513 ( new_n728_, new_n727_, keyIn_0_97 );
nor g514 ( new_n729_, new_n727_, keyIn_0_97 );
nand g515 ( new_n730_, new_n551_, N246 );
nand g516 ( new_n731_, new_n391_, N171 );
nand g517 ( new_n732_, new_n730_, new_n731_ );
xor g518 ( new_n733_, new_n732_, keyIn_0_77 );
nor g519 ( new_n734_, new_n728_, new_n729_, new_n733_ );
nand g520 ( new_n735_, new_n722_, new_n723_, new_n734_ );
nand g521 ( new_n736_, new_n735_, keyIn_0_127 );
not g522 ( new_n737_, keyIn_0_127 );
nand g523 ( new_n738_, new_n722_, new_n737_, new_n723_, new_n734_ );
and g524 ( N880, new_n736_, new_n738_ );
endmodule