module add_mul_sub_16_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, 
        b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, 
        b_14_, b_15_, operation_0_, operation_1_, Result_0_, Result_1_, 
        Result_2_, Result_3_, Result_4_, Result_5_, Result_6_, Result_7_, 
        Result_8_, Result_9_, Result_10_, Result_11_, Result_12_, Result_13_, 
        Result_14_, Result_15_, Result_16_, Result_17_, Result_18_, Result_19_, 
        Result_20_, Result_21_, Result_22_, Result_23_, Result_24_, Result_25_, 
        Result_26_, Result_27_, Result_28_, Result_29_, Result_30_, Result_31_
 );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_,
         b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_,
         operation_0_, operation_1_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_;
  wire   n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455;

  OR2_X1 U2202 ( .A1(n2170), .A2(n2171), .ZN(Result_9_) );
  AND2_X1 U2203 ( .A1(n2172), .A2(n2173), .ZN(n2170) );
  XOR2_X1 U2204 ( .A(n2174), .B(n2175), .Z(n2172) );
  OR2_X1 U2205 ( .A1(n2176), .A2(n2171), .ZN(Result_8_) );
  AND2_X1 U2206 ( .A1(n2173), .A2(n2177), .ZN(n2176) );
  XOR2_X1 U2207 ( .A(n2178), .B(n2179), .Z(n2177) );
  OR2_X1 U2208 ( .A1(n2180), .A2(n2171), .ZN(Result_7_) );
  AND2_X1 U2209 ( .A1(n2173), .A2(n2181), .ZN(n2180) );
  XOR2_X1 U2210 ( .A(n2182), .B(n2183), .Z(n2181) );
  OR2_X1 U2211 ( .A1(n2184), .A2(n2171), .ZN(Result_6_) );
  AND2_X1 U2212 ( .A1(n2173), .A2(n2185), .ZN(n2184) );
  XOR2_X1 U2213 ( .A(n2186), .B(n2187), .Z(n2185) );
  OR2_X1 U2214 ( .A1(n2188), .A2(n2171), .ZN(Result_5_) );
  AND2_X1 U2215 ( .A1(n2173), .A2(n2189), .ZN(n2188) );
  XOR2_X1 U2216 ( .A(n2190), .B(n2191), .Z(n2189) );
  OR2_X1 U2217 ( .A1(n2192), .A2(n2171), .ZN(Result_4_) );
  AND2_X1 U2218 ( .A1(n2173), .A2(n2193), .ZN(n2192) );
  XOR2_X1 U2219 ( .A(n2194), .B(n2195), .Z(n2193) );
  OR2_X1 U2220 ( .A1(n2196), .A2(n2171), .ZN(Result_3_) );
  AND2_X1 U2221 ( .A1(n2173), .A2(n2197), .ZN(n2196) );
  XOR2_X1 U2222 ( .A(n2198), .B(n2199), .Z(n2197) );
  OR2_X1 U2223 ( .A1(n2200), .A2(n2201), .ZN(Result_31_) );
  AND2_X1 U2224 ( .A1(n2202), .A2(n2173), .ZN(n2201) );
  AND2_X1 U2225 ( .A1(n2203), .A2(n2204), .ZN(n2200) );
  OR2_X1 U2226 ( .A1(n2205), .A2(n2206), .ZN(n2204) );
  OR2_X1 U2227 ( .A1(n2207), .A2(n2208), .ZN(n2206) );
  OR2_X1 U2228 ( .A1(n2209), .A2(n2210), .ZN(n2203) );
  OR2_X1 U2229 ( .A1(n2211), .A2(n2212), .ZN(Result_30_) );
  OR2_X1 U2230 ( .A1(n2213), .A2(n2214), .ZN(n2212) );
  AND2_X1 U2231 ( .A1(n2215), .A2(n2173), .ZN(n2214) );
  AND2_X1 U2232 ( .A1(b_14_), .A2(n2216), .ZN(n2215) );
  OR2_X1 U2233 ( .A1(n2209), .A2(n2217), .ZN(n2216) );
  AND2_X1 U2234 ( .A1(n2218), .A2(n2219), .ZN(n2213) );
  OR2_X1 U2235 ( .A1(n2220), .A2(n2221), .ZN(n2211) );
  AND2_X1 U2236 ( .A1(a_14_), .A2(n2222), .ZN(n2221) );
  OR2_X1 U2237 ( .A1(n2223), .A2(n2224), .ZN(n2222) );
  OR2_X1 U2238 ( .A1(n2225), .A2(n2226), .ZN(n2224) );
  AND2_X1 U2239 ( .A1(n2227), .A2(n2228), .ZN(n2226) );
  OR2_X1 U2240 ( .A1(n2229), .A2(n2219), .ZN(n2227) );
  OR2_X1 U2241 ( .A1(n2230), .A2(n2231), .ZN(n2219) );
  OR2_X1 U2242 ( .A1(n2232), .A2(n2233), .ZN(n2231) );
  AND2_X1 U2243 ( .A1(n2208), .A2(n2234), .ZN(n2233) );
  AND2_X1 U2244 ( .A1(n2205), .A2(n2235), .ZN(n2232) );
  AND2_X1 U2245 ( .A1(n2207), .A2(n2236), .ZN(n2230) );
  INV_X1 U2246 ( .A(n2210), .ZN(n2236) );
  AND2_X1 U2247 ( .A1(n2173), .A2(b_15_), .ZN(n2229) );
  AND2_X1 U2248 ( .A1(b_14_), .A2(n2237), .ZN(n2225) );
  AND2_X1 U2249 ( .A1(n2173), .A2(n2210), .ZN(n2223) );
  AND2_X1 U2250 ( .A1(n2238), .A2(n2239), .ZN(n2220) );
  AND2_X1 U2251 ( .A1(n2237), .A2(n2228), .ZN(n2238) );
  OR2_X1 U2252 ( .A1(n2240), .A2(n2241), .ZN(n2237) );
  OR2_X1 U2253 ( .A1(n2242), .A2(n2243), .ZN(n2241) );
  AND2_X1 U2254 ( .A1(n2208), .A2(n2209), .ZN(n2243) );
  AND2_X1 U2255 ( .A1(n2205), .A2(n2202), .ZN(n2242) );
  AND2_X1 U2256 ( .A1(n2207), .A2(n2210), .ZN(n2240) );
  OR2_X1 U2257 ( .A1(n2244), .A2(n2171), .ZN(Result_2_) );
  AND2_X1 U2258 ( .A1(n2173), .A2(n2245), .ZN(n2244) );
  XOR2_X1 U2259 ( .A(n2246), .B(n2247), .Z(n2245) );
  OR2_X1 U2260 ( .A1(n2248), .A2(n2249), .ZN(Result_29_) );
  OR2_X1 U2261 ( .A1(n2250), .A2(n2251), .ZN(n2249) );
  AND2_X1 U2262 ( .A1(n2252), .A2(n2253), .ZN(n2251) );
  OR2_X1 U2263 ( .A1(n2254), .A2(n2255), .ZN(n2253) );
  OR2_X1 U2264 ( .A1(n2256), .A2(n2257), .ZN(n2255) );
  AND2_X1 U2265 ( .A1(n2208), .A2(n2258), .ZN(n2257) );
  AND2_X1 U2266 ( .A1(n2205), .A2(n2259), .ZN(n2256) );
  INV_X1 U2267 ( .A(n2260), .ZN(n2259) );
  AND2_X1 U2268 ( .A1(n2207), .A2(n2261), .ZN(n2254) );
  INV_X1 U2269 ( .A(n2262), .ZN(n2252) );
  AND2_X1 U2270 ( .A1(n2262), .A2(n2263), .ZN(n2250) );
  OR2_X1 U2271 ( .A1(n2264), .A2(n2265), .ZN(n2263) );
  OR2_X1 U2272 ( .A1(n2266), .A2(n2267), .ZN(n2265) );
  AND2_X1 U2273 ( .A1(n2208), .A2(n2268), .ZN(n2267) );
  AND2_X1 U2274 ( .A1(n2260), .A2(n2205), .ZN(n2266) );
  AND2_X1 U2275 ( .A1(n2207), .A2(n2269), .ZN(n2264) );
  INV_X1 U2276 ( .A(n2261), .ZN(n2269) );
  XNOR2_X1 U2277 ( .A(a_13_), .B(n2270), .ZN(n2262) );
  AND2_X1 U2278 ( .A1(n2271), .A2(n2173), .ZN(n2248) );
  XOR2_X1 U2279 ( .A(n2272), .B(n2273), .Z(n2271) );
  XNOR2_X1 U2280 ( .A(n2274), .B(n2275), .ZN(n2273) );
  OR2_X1 U2281 ( .A1(n2276), .A2(n2277), .ZN(Result_28_) );
  OR2_X1 U2282 ( .A1(n2278), .A2(n2279), .ZN(n2277) );
  AND2_X1 U2283 ( .A1(n2280), .A2(n2281), .ZN(n2279) );
  OR2_X1 U2284 ( .A1(n2282), .A2(n2283), .ZN(n2281) );
  OR2_X1 U2285 ( .A1(n2284), .A2(n2285), .ZN(n2283) );
  AND2_X1 U2286 ( .A1(n2208), .A2(n2286), .ZN(n2285) );
  AND2_X1 U2287 ( .A1(n2287), .A2(n2205), .ZN(n2284) );
  INV_X1 U2288 ( .A(n2288), .ZN(n2287) );
  AND2_X1 U2289 ( .A1(n2207), .A2(n2289), .ZN(n2282) );
  INV_X1 U2290 ( .A(n2290), .ZN(n2280) );
  AND2_X1 U2291 ( .A1(n2290), .A2(n2291), .ZN(n2278) );
  OR2_X1 U2292 ( .A1(n2292), .A2(n2293), .ZN(n2291) );
  OR2_X1 U2293 ( .A1(n2294), .A2(n2295), .ZN(n2293) );
  AND2_X1 U2294 ( .A1(n2208), .A2(n2296), .ZN(n2295) );
  INV_X1 U2295 ( .A(n2286), .ZN(n2296) );
  AND2_X1 U2296 ( .A1(n2205), .A2(n2288), .ZN(n2294) );
  AND2_X1 U2297 ( .A1(n2207), .A2(n2297), .ZN(n2292) );
  INV_X1 U2298 ( .A(n2289), .ZN(n2297) );
  XNOR2_X1 U2299 ( .A(a_12_), .B(n2298), .ZN(n2290) );
  AND2_X1 U2300 ( .A1(n2299), .A2(n2173), .ZN(n2276) );
  XNOR2_X1 U2301 ( .A(n2300), .B(n2301), .ZN(n2299) );
  XOR2_X1 U2302 ( .A(n2302), .B(n2303), .Z(n2301) );
  OR2_X1 U2303 ( .A1(n2304), .A2(n2305), .ZN(Result_27_) );
  OR2_X1 U2304 ( .A1(n2306), .A2(n2307), .ZN(n2305) );
  AND2_X1 U2305 ( .A1(n2308), .A2(n2309), .ZN(n2307) );
  OR2_X1 U2306 ( .A1(n2310), .A2(n2311), .ZN(n2309) );
  OR2_X1 U2307 ( .A1(n2312), .A2(n2313), .ZN(n2311) );
  AND2_X1 U2308 ( .A1(n2208), .A2(n2314), .ZN(n2313) );
  AND2_X1 U2309 ( .A1(n2315), .A2(n2205), .ZN(n2312) );
  INV_X1 U2310 ( .A(n2316), .ZN(n2315) );
  AND2_X1 U2311 ( .A1(n2207), .A2(n2317), .ZN(n2310) );
  INV_X1 U2312 ( .A(n2318), .ZN(n2308) );
  AND2_X1 U2313 ( .A1(n2318), .A2(n2319), .ZN(n2306) );
  OR2_X1 U2314 ( .A1(n2320), .A2(n2321), .ZN(n2319) );
  OR2_X1 U2315 ( .A1(n2322), .A2(n2323), .ZN(n2321) );
  AND2_X1 U2316 ( .A1(n2208), .A2(n2324), .ZN(n2323) );
  INV_X1 U2317 ( .A(n2314), .ZN(n2324) );
  AND2_X1 U2318 ( .A1(n2205), .A2(n2316), .ZN(n2322) );
  AND2_X1 U2319 ( .A1(n2207), .A2(n2325), .ZN(n2320) );
  INV_X1 U2320 ( .A(n2317), .ZN(n2325) );
  XNOR2_X1 U2321 ( .A(a_11_), .B(n2326), .ZN(n2318) );
  AND2_X1 U2322 ( .A1(n2327), .A2(n2173), .ZN(n2304) );
  XNOR2_X1 U2323 ( .A(n2328), .B(n2329), .ZN(n2327) );
  XOR2_X1 U2324 ( .A(n2330), .B(n2331), .Z(n2329) );
  OR2_X1 U2325 ( .A1(n2332), .A2(n2333), .ZN(Result_26_) );
  OR2_X1 U2326 ( .A1(n2334), .A2(n2335), .ZN(n2333) );
  AND2_X1 U2327 ( .A1(n2336), .A2(n2337), .ZN(n2335) );
  OR2_X1 U2328 ( .A1(n2338), .A2(n2339), .ZN(n2337) );
  OR2_X1 U2329 ( .A1(n2340), .A2(n2341), .ZN(n2339) );
  AND2_X1 U2330 ( .A1(n2208), .A2(n2342), .ZN(n2341) );
  AND2_X1 U2331 ( .A1(n2343), .A2(n2205), .ZN(n2340) );
  INV_X1 U2332 ( .A(n2344), .ZN(n2343) );
  AND2_X1 U2333 ( .A1(n2207), .A2(n2345), .ZN(n2338) );
  INV_X1 U2334 ( .A(n2346), .ZN(n2336) );
  AND2_X1 U2335 ( .A1(n2346), .A2(n2347), .ZN(n2334) );
  OR2_X1 U2336 ( .A1(n2348), .A2(n2349), .ZN(n2347) );
  OR2_X1 U2337 ( .A1(n2350), .A2(n2351), .ZN(n2349) );
  AND2_X1 U2338 ( .A1(n2208), .A2(n2352), .ZN(n2351) );
  INV_X1 U2339 ( .A(n2342), .ZN(n2352) );
  AND2_X1 U2340 ( .A1(n2205), .A2(n2344), .ZN(n2350) );
  AND2_X1 U2341 ( .A1(n2207), .A2(n2353), .ZN(n2348) );
  INV_X1 U2342 ( .A(n2345), .ZN(n2353) );
  XNOR2_X1 U2343 ( .A(a_10_), .B(n2354), .ZN(n2346) );
  AND2_X1 U2344 ( .A1(n2355), .A2(n2173), .ZN(n2332) );
  XNOR2_X1 U2345 ( .A(n2356), .B(n2357), .ZN(n2355) );
  XOR2_X1 U2346 ( .A(n2358), .B(n2359), .Z(n2357) );
  OR2_X1 U2347 ( .A1(n2360), .A2(n2361), .ZN(Result_25_) );
  OR2_X1 U2348 ( .A1(n2362), .A2(n2363), .ZN(n2361) );
  AND2_X1 U2349 ( .A1(n2364), .A2(n2365), .ZN(n2363) );
  OR2_X1 U2350 ( .A1(n2366), .A2(n2367), .ZN(n2365) );
  OR2_X1 U2351 ( .A1(n2368), .A2(n2369), .ZN(n2367) );
  AND2_X1 U2352 ( .A1(n2208), .A2(n2370), .ZN(n2369) );
  AND2_X1 U2353 ( .A1(n2371), .A2(n2205), .ZN(n2368) );
  INV_X1 U2354 ( .A(n2372), .ZN(n2371) );
  AND2_X1 U2355 ( .A1(n2207), .A2(n2373), .ZN(n2366) );
  INV_X1 U2356 ( .A(n2374), .ZN(n2364) );
  AND2_X1 U2357 ( .A1(n2374), .A2(n2375), .ZN(n2362) );
  OR2_X1 U2358 ( .A1(n2376), .A2(n2377), .ZN(n2375) );
  OR2_X1 U2359 ( .A1(n2378), .A2(n2379), .ZN(n2377) );
  AND2_X1 U2360 ( .A1(n2208), .A2(n2380), .ZN(n2379) );
  INV_X1 U2361 ( .A(n2370), .ZN(n2380) );
  AND2_X1 U2362 ( .A1(n2205), .A2(n2372), .ZN(n2378) );
  AND2_X1 U2363 ( .A1(n2207), .A2(n2381), .ZN(n2376) );
  INV_X1 U2364 ( .A(n2373), .ZN(n2381) );
  XNOR2_X1 U2365 ( .A(a_9_), .B(n2382), .ZN(n2374) );
  AND2_X1 U2366 ( .A1(n2383), .A2(n2173), .ZN(n2360) );
  XNOR2_X1 U2367 ( .A(n2384), .B(n2385), .ZN(n2383) );
  XOR2_X1 U2368 ( .A(n2386), .B(n2387), .Z(n2385) );
  OR2_X1 U2369 ( .A1(n2388), .A2(n2389), .ZN(Result_24_) );
  OR2_X1 U2370 ( .A1(n2390), .A2(n2391), .ZN(n2389) );
  AND2_X1 U2371 ( .A1(n2392), .A2(n2393), .ZN(n2391) );
  OR2_X1 U2372 ( .A1(n2394), .A2(n2395), .ZN(n2393) );
  OR2_X1 U2373 ( .A1(n2396), .A2(n2397), .ZN(n2395) );
  AND2_X1 U2374 ( .A1(n2208), .A2(n2398), .ZN(n2397) );
  INV_X1 U2375 ( .A(n2399), .ZN(n2398) );
  AND2_X1 U2376 ( .A1(n2205), .A2(n2400), .ZN(n2396) );
  AND2_X1 U2377 ( .A1(n2207), .A2(n2401), .ZN(n2394) );
  INV_X1 U2378 ( .A(n2402), .ZN(n2401) );
  AND2_X1 U2379 ( .A1(n2403), .A2(n2404), .ZN(n2390) );
  INV_X1 U2380 ( .A(n2392), .ZN(n2404) );
  AND2_X1 U2381 ( .A1(n2405), .A2(n2406), .ZN(n2392) );
  OR2_X1 U2382 ( .A1(a_8_), .A2(b_8_), .ZN(n2405) );
  OR2_X1 U2383 ( .A1(n2407), .A2(n2408), .ZN(n2403) );
  OR2_X1 U2384 ( .A1(n2409), .A2(n2410), .ZN(n2408) );
  AND2_X1 U2385 ( .A1(n2208), .A2(n2399), .ZN(n2410) );
  AND2_X1 U2386 ( .A1(n2411), .A2(n2205), .ZN(n2409) );
  INV_X1 U2387 ( .A(n2400), .ZN(n2411) );
  AND2_X1 U2388 ( .A1(n2207), .A2(n2402), .ZN(n2407) );
  AND2_X1 U2389 ( .A1(n2412), .A2(n2173), .ZN(n2388) );
  XNOR2_X1 U2390 ( .A(n2413), .B(n2414), .ZN(n2412) );
  XOR2_X1 U2391 ( .A(n2415), .B(n2416), .Z(n2414) );
  OR2_X1 U2392 ( .A1(n2417), .A2(n2418), .ZN(Result_23_) );
  OR2_X1 U2393 ( .A1(n2419), .A2(n2420), .ZN(n2418) );
  AND2_X1 U2394 ( .A1(n2421), .A2(n2422), .ZN(n2420) );
  OR2_X1 U2395 ( .A1(n2423), .A2(n2424), .ZN(n2422) );
  OR2_X1 U2396 ( .A1(n2425), .A2(n2426), .ZN(n2424) );
  AND2_X1 U2397 ( .A1(n2208), .A2(n2427), .ZN(n2426) );
  INV_X1 U2398 ( .A(n2428), .ZN(n2427) );
  AND2_X1 U2399 ( .A1(n2205), .A2(n2429), .ZN(n2425) );
  AND2_X1 U2400 ( .A1(n2207), .A2(n2430), .ZN(n2423) );
  INV_X1 U2401 ( .A(n2431), .ZN(n2430) );
  AND2_X1 U2402 ( .A1(n2432), .A2(n2433), .ZN(n2419) );
  INV_X1 U2403 ( .A(n2421), .ZN(n2433) );
  AND2_X1 U2404 ( .A1(n2434), .A2(n2435), .ZN(n2421) );
  OR2_X1 U2405 ( .A1(a_7_), .A2(b_7_), .ZN(n2434) );
  OR2_X1 U2406 ( .A1(n2436), .A2(n2437), .ZN(n2432) );
  OR2_X1 U2407 ( .A1(n2438), .A2(n2439), .ZN(n2437) );
  AND2_X1 U2408 ( .A1(n2208), .A2(n2428), .ZN(n2439) );
  AND2_X1 U2409 ( .A1(n2440), .A2(n2205), .ZN(n2438) );
  INV_X1 U2410 ( .A(n2429), .ZN(n2440) );
  AND2_X1 U2411 ( .A1(n2207), .A2(n2431), .ZN(n2436) );
  AND2_X1 U2412 ( .A1(n2441), .A2(n2173), .ZN(n2417) );
  XNOR2_X1 U2413 ( .A(n2442), .B(n2443), .ZN(n2441) );
  XOR2_X1 U2414 ( .A(n2444), .B(n2445), .Z(n2443) );
  OR2_X1 U2415 ( .A1(n2446), .A2(n2447), .ZN(Result_22_) );
  OR2_X1 U2416 ( .A1(n2448), .A2(n2449), .ZN(n2447) );
  AND2_X1 U2417 ( .A1(n2450), .A2(n2451), .ZN(n2449) );
  OR2_X1 U2418 ( .A1(n2452), .A2(n2453), .ZN(n2451) );
  OR2_X1 U2419 ( .A1(n2454), .A2(n2455), .ZN(n2453) );
  AND2_X1 U2420 ( .A1(n2208), .A2(n2456), .ZN(n2455) );
  INV_X1 U2421 ( .A(n2457), .ZN(n2456) );
  AND2_X1 U2422 ( .A1(n2205), .A2(n2458), .ZN(n2454) );
  AND2_X1 U2423 ( .A1(n2207), .A2(n2459), .ZN(n2452) );
  INV_X1 U2424 ( .A(n2460), .ZN(n2459) );
  AND2_X1 U2425 ( .A1(n2461), .A2(n2462), .ZN(n2448) );
  INV_X1 U2426 ( .A(n2450), .ZN(n2462) );
  AND2_X1 U2427 ( .A1(n2463), .A2(n2464), .ZN(n2450) );
  OR2_X1 U2428 ( .A1(a_6_), .A2(b_6_), .ZN(n2463) );
  OR2_X1 U2429 ( .A1(n2465), .A2(n2466), .ZN(n2461) );
  OR2_X1 U2430 ( .A1(n2467), .A2(n2468), .ZN(n2466) );
  AND2_X1 U2431 ( .A1(n2208), .A2(n2457), .ZN(n2468) );
  AND2_X1 U2432 ( .A1(n2469), .A2(n2205), .ZN(n2467) );
  INV_X1 U2433 ( .A(n2458), .ZN(n2469) );
  AND2_X1 U2434 ( .A1(n2207), .A2(n2460), .ZN(n2465) );
  AND2_X1 U2435 ( .A1(n2470), .A2(n2173), .ZN(n2446) );
  XNOR2_X1 U2436 ( .A(n2471), .B(n2472), .ZN(n2470) );
  XOR2_X1 U2437 ( .A(n2473), .B(n2474), .Z(n2472) );
  OR2_X1 U2438 ( .A1(n2475), .A2(n2476), .ZN(Result_21_) );
  OR2_X1 U2439 ( .A1(n2477), .A2(n2478), .ZN(n2476) );
  AND2_X1 U2440 ( .A1(n2479), .A2(n2480), .ZN(n2478) );
  OR2_X1 U2441 ( .A1(n2481), .A2(n2482), .ZN(n2480) );
  OR2_X1 U2442 ( .A1(n2483), .A2(n2484), .ZN(n2482) );
  AND2_X1 U2443 ( .A1(n2208), .A2(n2485), .ZN(n2484) );
  INV_X1 U2444 ( .A(n2486), .ZN(n2485) );
  AND2_X1 U2445 ( .A1(n2205), .A2(n2487), .ZN(n2483) );
  AND2_X1 U2446 ( .A1(n2207), .A2(n2488), .ZN(n2481) );
  INV_X1 U2447 ( .A(n2489), .ZN(n2488) );
  AND2_X1 U2448 ( .A1(n2490), .A2(n2491), .ZN(n2477) );
  INV_X1 U2449 ( .A(n2479), .ZN(n2491) );
  AND2_X1 U2450 ( .A1(n2492), .A2(n2493), .ZN(n2479) );
  OR2_X1 U2451 ( .A1(a_5_), .A2(b_5_), .ZN(n2492) );
  OR2_X1 U2452 ( .A1(n2494), .A2(n2495), .ZN(n2490) );
  OR2_X1 U2453 ( .A1(n2496), .A2(n2497), .ZN(n2495) );
  AND2_X1 U2454 ( .A1(n2208), .A2(n2486), .ZN(n2497) );
  AND2_X1 U2455 ( .A1(n2498), .A2(n2205), .ZN(n2496) );
  INV_X1 U2456 ( .A(n2487), .ZN(n2498) );
  AND2_X1 U2457 ( .A1(n2207), .A2(n2489), .ZN(n2494) );
  AND2_X1 U2458 ( .A1(n2499), .A2(n2173), .ZN(n2475) );
  XNOR2_X1 U2459 ( .A(n2500), .B(n2501), .ZN(n2499) );
  XOR2_X1 U2460 ( .A(n2502), .B(n2503), .Z(n2501) );
  OR2_X1 U2461 ( .A1(n2504), .A2(n2505), .ZN(Result_20_) );
  OR2_X1 U2462 ( .A1(n2506), .A2(n2507), .ZN(n2505) );
  AND2_X1 U2463 ( .A1(n2508), .A2(n2509), .ZN(n2507) );
  OR2_X1 U2464 ( .A1(n2510), .A2(n2511), .ZN(n2509) );
  OR2_X1 U2465 ( .A1(n2512), .A2(n2513), .ZN(n2511) );
  AND2_X1 U2466 ( .A1(n2208), .A2(n2514), .ZN(n2513) );
  INV_X1 U2467 ( .A(n2515), .ZN(n2514) );
  AND2_X1 U2468 ( .A1(n2205), .A2(n2516), .ZN(n2512) );
  AND2_X1 U2469 ( .A1(n2207), .A2(n2517), .ZN(n2510) );
  INV_X1 U2470 ( .A(n2518), .ZN(n2517) );
  AND2_X1 U2471 ( .A1(n2519), .A2(n2520), .ZN(n2506) );
  INV_X1 U2472 ( .A(n2508), .ZN(n2520) );
  AND2_X1 U2473 ( .A1(n2521), .A2(n2522), .ZN(n2508) );
  OR2_X1 U2474 ( .A1(a_4_), .A2(b_4_), .ZN(n2521) );
  OR2_X1 U2475 ( .A1(n2523), .A2(n2524), .ZN(n2519) );
  OR2_X1 U2476 ( .A1(n2525), .A2(n2526), .ZN(n2524) );
  AND2_X1 U2477 ( .A1(n2208), .A2(n2515), .ZN(n2526) );
  AND2_X1 U2478 ( .A1(n2527), .A2(n2205), .ZN(n2525) );
  INV_X1 U2479 ( .A(n2516), .ZN(n2527) );
  AND2_X1 U2480 ( .A1(n2207), .A2(n2518), .ZN(n2523) );
  AND2_X1 U2481 ( .A1(n2528), .A2(n2173), .ZN(n2504) );
  XNOR2_X1 U2482 ( .A(n2529), .B(n2530), .ZN(n2528) );
  XOR2_X1 U2483 ( .A(n2531), .B(n2532), .Z(n2530) );
  OR2_X1 U2484 ( .A1(n2533), .A2(n2171), .ZN(Result_1_) );
  AND2_X1 U2485 ( .A1(n2173), .A2(n2534), .ZN(n2533) );
  XOR2_X1 U2486 ( .A(n2535), .B(n2536), .Z(n2534) );
  AND2_X1 U2487 ( .A1(n2537), .A2(n2538), .ZN(n2536) );
  OR2_X1 U2488 ( .A1(n2539), .A2(n2540), .ZN(n2538) );
  AND2_X1 U2489 ( .A1(n2541), .A2(n2542), .ZN(n2539) );
  INV_X1 U2490 ( .A(n2543), .ZN(n2537) );
  OR2_X1 U2491 ( .A1(n2544), .A2(n2545), .ZN(Result_19_) );
  OR2_X1 U2492 ( .A1(n2546), .A2(n2547), .ZN(n2545) );
  AND2_X1 U2493 ( .A1(n2548), .A2(n2549), .ZN(n2547) );
  OR2_X1 U2494 ( .A1(n2550), .A2(n2551), .ZN(n2549) );
  OR2_X1 U2495 ( .A1(n2552), .A2(n2553), .ZN(n2551) );
  AND2_X1 U2496 ( .A1(n2208), .A2(n2554), .ZN(n2553) );
  INV_X1 U2497 ( .A(n2555), .ZN(n2554) );
  AND2_X1 U2498 ( .A1(n2205), .A2(n2556), .ZN(n2552) );
  AND2_X1 U2499 ( .A1(n2207), .A2(n2557), .ZN(n2550) );
  INV_X1 U2500 ( .A(n2558), .ZN(n2557) );
  AND2_X1 U2501 ( .A1(n2559), .A2(n2560), .ZN(n2546) );
  INV_X1 U2502 ( .A(n2548), .ZN(n2560) );
  AND2_X1 U2503 ( .A1(n2561), .A2(n2562), .ZN(n2548) );
  OR2_X1 U2504 ( .A1(a_3_), .A2(b_3_), .ZN(n2561) );
  OR2_X1 U2505 ( .A1(n2563), .A2(n2564), .ZN(n2559) );
  OR2_X1 U2506 ( .A1(n2565), .A2(n2566), .ZN(n2564) );
  AND2_X1 U2507 ( .A1(n2208), .A2(n2555), .ZN(n2566) );
  AND2_X1 U2508 ( .A1(n2567), .A2(n2205), .ZN(n2565) );
  INV_X1 U2509 ( .A(n2556), .ZN(n2567) );
  AND2_X1 U2510 ( .A1(n2207), .A2(n2558), .ZN(n2563) );
  AND2_X1 U2511 ( .A1(n2568), .A2(n2173), .ZN(n2544) );
  XNOR2_X1 U2512 ( .A(n2569), .B(n2570), .ZN(n2568) );
  XOR2_X1 U2513 ( .A(n2571), .B(n2572), .Z(n2570) );
  OR2_X1 U2514 ( .A1(n2573), .A2(n2574), .ZN(Result_18_) );
  OR2_X1 U2515 ( .A1(n2575), .A2(n2576), .ZN(n2574) );
  AND2_X1 U2516 ( .A1(n2577), .A2(n2578), .ZN(n2576) );
  OR2_X1 U2517 ( .A1(n2579), .A2(n2580), .ZN(n2578) );
  OR2_X1 U2518 ( .A1(n2581), .A2(n2582), .ZN(n2580) );
  AND2_X1 U2519 ( .A1(n2208), .A2(n2583), .ZN(n2582) );
  INV_X1 U2520 ( .A(n2584), .ZN(n2583) );
  AND2_X1 U2521 ( .A1(n2205), .A2(n2585), .ZN(n2581) );
  AND2_X1 U2522 ( .A1(n2207), .A2(n2586), .ZN(n2579) );
  INV_X1 U2523 ( .A(n2587), .ZN(n2586) );
  AND2_X1 U2524 ( .A1(n2588), .A2(n2589), .ZN(n2575) );
  INV_X1 U2525 ( .A(n2577), .ZN(n2589) );
  AND2_X1 U2526 ( .A1(n2590), .A2(n2591), .ZN(n2577) );
  OR2_X1 U2527 ( .A1(a_2_), .A2(b_2_), .ZN(n2590) );
  OR2_X1 U2528 ( .A1(n2592), .A2(n2593), .ZN(n2588) );
  OR2_X1 U2529 ( .A1(n2594), .A2(n2595), .ZN(n2593) );
  AND2_X1 U2530 ( .A1(n2208), .A2(n2584), .ZN(n2595) );
  AND2_X1 U2531 ( .A1(n2596), .A2(n2205), .ZN(n2594) );
  INV_X1 U2532 ( .A(n2585), .ZN(n2596) );
  AND2_X1 U2533 ( .A1(n2207), .A2(n2587), .ZN(n2592) );
  AND2_X1 U2534 ( .A1(n2597), .A2(n2173), .ZN(n2573) );
  XNOR2_X1 U2535 ( .A(n2598), .B(n2599), .ZN(n2597) );
  XOR2_X1 U2536 ( .A(n2600), .B(n2601), .Z(n2599) );
  OR2_X1 U2537 ( .A1(n2602), .A2(n2603), .ZN(Result_17_) );
  OR2_X1 U2538 ( .A1(n2604), .A2(n2605), .ZN(n2603) );
  AND2_X1 U2539 ( .A1(n2606), .A2(n2607), .ZN(n2605) );
  OR2_X1 U2540 ( .A1(n2608), .A2(n2609), .ZN(n2607) );
  OR2_X1 U2541 ( .A1(n2610), .A2(n2611), .ZN(n2609) );
  AND2_X1 U2542 ( .A1(n2208), .A2(n2612), .ZN(n2611) );
  INV_X1 U2543 ( .A(n2613), .ZN(n2612) );
  AND2_X1 U2544 ( .A1(n2205), .A2(n2614), .ZN(n2610) );
  AND2_X1 U2545 ( .A1(n2207), .A2(n2615), .ZN(n2608) );
  INV_X1 U2546 ( .A(n2616), .ZN(n2615) );
  AND2_X1 U2547 ( .A1(n2617), .A2(n2618), .ZN(n2604) );
  INV_X1 U2548 ( .A(n2606), .ZN(n2618) );
  AND2_X1 U2549 ( .A1(n2619), .A2(n2620), .ZN(n2606) );
  OR2_X1 U2550 ( .A1(a_1_), .A2(b_1_), .ZN(n2619) );
  OR2_X1 U2551 ( .A1(n2621), .A2(n2622), .ZN(n2617) );
  OR2_X1 U2552 ( .A1(n2623), .A2(n2624), .ZN(n2622) );
  AND2_X1 U2553 ( .A1(n2208), .A2(n2613), .ZN(n2624) );
  AND2_X1 U2554 ( .A1(n2625), .A2(n2205), .ZN(n2623) );
  INV_X1 U2555 ( .A(n2614), .ZN(n2625) );
  AND2_X1 U2556 ( .A1(n2207), .A2(n2616), .ZN(n2621) );
  AND2_X1 U2557 ( .A1(n2626), .A2(n2173), .ZN(n2602) );
  XNOR2_X1 U2558 ( .A(n2627), .B(n2628), .ZN(n2626) );
  XOR2_X1 U2559 ( .A(n2629), .B(n2630), .Z(n2628) );
  OR2_X1 U2560 ( .A1(n2631), .A2(n2632), .ZN(Result_16_) );
  OR2_X1 U2561 ( .A1(n2633), .A2(n2634), .ZN(n2632) );
  AND2_X1 U2562 ( .A1(n2635), .A2(n2636), .ZN(n2634) );
  INV_X1 U2563 ( .A(n2637), .ZN(n2636) );
  OR2_X1 U2564 ( .A1(n2638), .A2(n2639), .ZN(n2635) );
  OR2_X1 U2565 ( .A1(n2640), .A2(n2641), .ZN(n2639) );
  AND2_X1 U2566 ( .A1(n2208), .A2(n2642), .ZN(n2641) );
  AND2_X1 U2567 ( .A1(n2205), .A2(n2643), .ZN(n2640) );
  AND2_X1 U2568 ( .A1(n2644), .A2(n2207), .ZN(n2638) );
  INV_X1 U2569 ( .A(n2645), .ZN(n2644) );
  AND2_X1 U2570 ( .A1(n2637), .A2(n2646), .ZN(n2633) );
  OR2_X1 U2571 ( .A1(n2647), .A2(n2648), .ZN(n2646) );
  OR2_X1 U2572 ( .A1(n2649), .A2(n2650), .ZN(n2648) );
  AND2_X1 U2573 ( .A1(n2208), .A2(n2651), .ZN(n2650) );
  AND2_X1 U2574 ( .A1(n2652), .A2(n2205), .ZN(n2649) );
  AND2_X1 U2575 ( .A1(n2653), .A2(n2654), .ZN(n2205) );
  INV_X1 U2576 ( .A(n2643), .ZN(n2652) );
  OR2_X1 U2577 ( .A1(n2655), .A2(n2656), .ZN(n2643) );
  AND2_X1 U2578 ( .A1(n2657), .A2(n2658), .ZN(n2656) );
  AND2_X1 U2579 ( .A1(n2614), .A2(n2620), .ZN(n2655) );
  OR2_X1 U2580 ( .A1(n2659), .A2(n2660), .ZN(n2614) );
  AND2_X1 U2581 ( .A1(n2661), .A2(n2662), .ZN(n2660) );
  AND2_X1 U2582 ( .A1(n2585), .A2(n2591), .ZN(n2659) );
  OR2_X1 U2583 ( .A1(n2663), .A2(n2664), .ZN(n2585) );
  AND2_X1 U2584 ( .A1(n2665), .A2(n2666), .ZN(n2664) );
  AND2_X1 U2585 ( .A1(n2556), .A2(n2562), .ZN(n2663) );
  OR2_X1 U2586 ( .A1(n2667), .A2(n2668), .ZN(n2556) );
  AND2_X1 U2587 ( .A1(n2669), .A2(n2670), .ZN(n2668) );
  AND2_X1 U2588 ( .A1(n2516), .A2(n2522), .ZN(n2667) );
  OR2_X1 U2589 ( .A1(n2671), .A2(n2672), .ZN(n2516) );
  AND2_X1 U2590 ( .A1(n2673), .A2(n2674), .ZN(n2672) );
  AND2_X1 U2591 ( .A1(n2487), .A2(n2493), .ZN(n2671) );
  OR2_X1 U2592 ( .A1(n2675), .A2(n2676), .ZN(n2487) );
  AND2_X1 U2593 ( .A1(n2677), .A2(n2678), .ZN(n2676) );
  AND2_X1 U2594 ( .A1(n2458), .A2(n2464), .ZN(n2675) );
  OR2_X1 U2595 ( .A1(n2679), .A2(n2680), .ZN(n2458) );
  AND2_X1 U2596 ( .A1(n2681), .A2(n2682), .ZN(n2680) );
  AND2_X1 U2597 ( .A1(n2429), .A2(n2435), .ZN(n2679) );
  OR2_X1 U2598 ( .A1(n2683), .A2(n2684), .ZN(n2429) );
  AND2_X1 U2599 ( .A1(n2685), .A2(n2686), .ZN(n2684) );
  AND2_X1 U2600 ( .A1(n2400), .A2(n2406), .ZN(n2683) );
  OR2_X1 U2601 ( .A1(n2687), .A2(n2688), .ZN(n2400) );
  AND2_X1 U2602 ( .A1(n2689), .A2(n2382), .ZN(n2688) );
  AND2_X1 U2603 ( .A1(n2372), .A2(n2690), .ZN(n2687) );
  OR2_X1 U2604 ( .A1(n2691), .A2(n2692), .ZN(n2372) );
  AND2_X1 U2605 ( .A1(n2693), .A2(n2354), .ZN(n2692) );
  AND2_X1 U2606 ( .A1(n2344), .A2(n2694), .ZN(n2691) );
  OR2_X1 U2607 ( .A1(n2695), .A2(n2696), .ZN(n2344) );
  AND2_X1 U2608 ( .A1(n2697), .A2(n2326), .ZN(n2696) );
  AND2_X1 U2609 ( .A1(n2316), .A2(n2698), .ZN(n2695) );
  OR2_X1 U2610 ( .A1(n2699), .A2(n2700), .ZN(n2316) );
  AND2_X1 U2611 ( .A1(n2701), .A2(n2298), .ZN(n2700) );
  AND2_X1 U2612 ( .A1(n2288), .A2(n2702), .ZN(n2699) );
  OR2_X1 U2613 ( .A1(n2703), .A2(n2704), .ZN(n2288) );
  AND2_X1 U2614 ( .A1(n2705), .A2(n2270), .ZN(n2704) );
  AND2_X1 U2615 ( .A1(n2260), .A2(n2706), .ZN(n2703) );
  AND2_X1 U2616 ( .A1(n2707), .A2(n2708), .ZN(n2260) );
  OR2_X1 U2617 ( .A1(n2228), .A2(n2709), .ZN(n2708) );
  AND2_X1 U2618 ( .A1(n2239), .A2(n2235), .ZN(n2709) );
  INV_X1 U2619 ( .A(n2202), .ZN(n2235) );
  AND2_X1 U2620 ( .A1(a_15_), .A2(b_15_), .ZN(n2202) );
  AND2_X1 U2621 ( .A1(n2207), .A2(n2645), .ZN(n2647) );
  AND2_X1 U2622 ( .A1(n2710), .A2(n2711), .ZN(n2637) );
  AND2_X1 U2623 ( .A1(n2712), .A2(n2173), .ZN(n2631) );
  XNOR2_X1 U2624 ( .A(n2713), .B(n2714), .ZN(n2712) );
  XOR2_X1 U2625 ( .A(n2715), .B(n2716), .Z(n2714) );
  OR2_X1 U2626 ( .A1(n2717), .A2(n2171), .ZN(Result_15_) );
  AND2_X1 U2627 ( .A1(n2173), .A2(n2718), .ZN(n2717) );
  XNOR2_X1 U2628 ( .A(n2719), .B(n2720), .ZN(n2718) );
  OR2_X1 U2629 ( .A1(n2721), .A2(n2171), .ZN(Result_14_) );
  AND2_X1 U2630 ( .A1(n2722), .A2(n2173), .ZN(n2721) );
  AND2_X1 U2631 ( .A1(n2723), .A2(n2724), .ZN(n2722) );
  OR2_X1 U2632 ( .A1(n2725), .A2(n2726), .ZN(n2723) );
  AND2_X1 U2633 ( .A1(n2727), .A2(n2720), .ZN(n2725) );
  OR2_X1 U2634 ( .A1(n2728), .A2(n2171), .ZN(Result_13_) );
  AND2_X1 U2635 ( .A1(n2173), .A2(n2729), .ZN(n2728) );
  XOR2_X1 U2636 ( .A(n2724), .B(n2730), .Z(n2729) );
  OR2_X1 U2637 ( .A1(n2731), .A2(n2732), .ZN(n2730) );
  AND2_X1 U2638 ( .A1(n2733), .A2(n2734), .ZN(n2732) );
  INV_X1 U2639 ( .A(n2735), .ZN(n2724) );
  OR2_X1 U2640 ( .A1(n2736), .A2(n2171), .ZN(Result_12_) );
  AND2_X1 U2641 ( .A1(n2737), .A2(n2173), .ZN(n2736) );
  XOR2_X1 U2642 ( .A(n2738), .B(n2739), .Z(n2737) );
  AND2_X1 U2643 ( .A1(n2740), .A2(n2741), .ZN(n2739) );
  OR2_X1 U2644 ( .A1(n2742), .A2(n2743), .ZN(n2741) );
  INV_X1 U2645 ( .A(n2744), .ZN(n2740) );
  OR2_X1 U2646 ( .A1(n2745), .A2(n2171), .ZN(Result_11_) );
  AND2_X1 U2647 ( .A1(n2746), .A2(n2173), .ZN(n2745) );
  XOR2_X1 U2648 ( .A(n2747), .B(n2748), .Z(n2746) );
  AND2_X1 U2649 ( .A1(n2749), .A2(n2750), .ZN(n2748) );
  OR2_X1 U2650 ( .A1(n2751), .A2(n2752), .ZN(n2750) );
  AND2_X1 U2651 ( .A1(n2753), .A2(n2754), .ZN(n2751) );
  INV_X1 U2652 ( .A(n2755), .ZN(n2749) );
  OR2_X1 U2653 ( .A1(n2756), .A2(n2171), .ZN(Result_10_) );
  AND2_X1 U2654 ( .A1(n2757), .A2(n2173), .ZN(n2756) );
  XOR2_X1 U2655 ( .A(n2758), .B(n2759), .Z(n2757) );
  AND2_X1 U2656 ( .A1(n2760), .A2(n2761), .ZN(n2759) );
  OR2_X1 U2657 ( .A1(n2762), .A2(n2763), .ZN(n2761) );
  INV_X1 U2658 ( .A(n2764), .ZN(n2760) );
  OR2_X1 U2659 ( .A1(n2765), .A2(n2171), .ZN(Result_0_) );
  OR2_X1 U2660 ( .A1(n2766), .A2(n2767), .ZN(n2171) );
  AND2_X1 U2661 ( .A1(n2207), .A2(n2768), .ZN(n2767) );
  OR2_X1 U2662 ( .A1(n2769), .A2(n2770), .ZN(n2768) );
  AND2_X1 U2663 ( .A1(n2645), .A2(n2711), .ZN(n2769) );
  OR2_X1 U2664 ( .A1(n2771), .A2(n2772), .ZN(n2645) );
  AND2_X1 U2665 ( .A1(n2616), .A2(n2657), .ZN(n2772) );
  AND2_X1 U2666 ( .A1(b_1_), .A2(n2773), .ZN(n2771) );
  OR2_X1 U2667 ( .A1(n2657), .A2(n2616), .ZN(n2773) );
  OR2_X1 U2668 ( .A1(n2774), .A2(n2775), .ZN(n2616) );
  AND2_X1 U2669 ( .A1(n2587), .A2(n2661), .ZN(n2775) );
  AND2_X1 U2670 ( .A1(b_2_), .A2(n2776), .ZN(n2774) );
  OR2_X1 U2671 ( .A1(n2661), .A2(n2587), .ZN(n2776) );
  OR2_X1 U2672 ( .A1(n2777), .A2(n2778), .ZN(n2587) );
  AND2_X1 U2673 ( .A1(n2558), .A2(n2665), .ZN(n2778) );
  AND2_X1 U2674 ( .A1(b_3_), .A2(n2779), .ZN(n2777) );
  OR2_X1 U2675 ( .A1(n2665), .A2(n2558), .ZN(n2779) );
  OR2_X1 U2676 ( .A1(n2780), .A2(n2781), .ZN(n2558) );
  AND2_X1 U2677 ( .A1(n2518), .A2(n2669), .ZN(n2781) );
  AND2_X1 U2678 ( .A1(b_4_), .A2(n2782), .ZN(n2780) );
  OR2_X1 U2679 ( .A1(n2669), .A2(n2518), .ZN(n2782) );
  OR2_X1 U2680 ( .A1(n2783), .A2(n2784), .ZN(n2518) );
  AND2_X1 U2681 ( .A1(n2489), .A2(n2673), .ZN(n2784) );
  AND2_X1 U2682 ( .A1(b_5_), .A2(n2785), .ZN(n2783) );
  OR2_X1 U2683 ( .A1(n2673), .A2(n2489), .ZN(n2785) );
  OR2_X1 U2684 ( .A1(n2786), .A2(n2787), .ZN(n2489) );
  AND2_X1 U2685 ( .A1(n2460), .A2(n2677), .ZN(n2787) );
  AND2_X1 U2686 ( .A1(b_6_), .A2(n2788), .ZN(n2786) );
  OR2_X1 U2687 ( .A1(n2677), .A2(n2460), .ZN(n2788) );
  OR2_X1 U2688 ( .A1(n2789), .A2(n2790), .ZN(n2460) );
  AND2_X1 U2689 ( .A1(n2431), .A2(n2681), .ZN(n2790) );
  AND2_X1 U2690 ( .A1(b_7_), .A2(n2791), .ZN(n2789) );
  OR2_X1 U2691 ( .A1(n2681), .A2(n2431), .ZN(n2791) );
  OR2_X1 U2692 ( .A1(n2792), .A2(n2793), .ZN(n2431) );
  AND2_X1 U2693 ( .A1(n2402), .A2(n2685), .ZN(n2793) );
  AND2_X1 U2694 ( .A1(b_8_), .A2(n2794), .ZN(n2792) );
  OR2_X1 U2695 ( .A1(n2685), .A2(n2402), .ZN(n2794) );
  OR2_X1 U2696 ( .A1(n2795), .A2(n2796), .ZN(n2402) );
  AND2_X1 U2697 ( .A1(n2373), .A2(n2689), .ZN(n2796) );
  AND2_X1 U2698 ( .A1(b_9_), .A2(n2797), .ZN(n2795) );
  OR2_X1 U2699 ( .A1(n2689), .A2(n2373), .ZN(n2797) );
  OR2_X1 U2700 ( .A1(n2798), .A2(n2799), .ZN(n2373) );
  AND2_X1 U2701 ( .A1(n2345), .A2(n2693), .ZN(n2799) );
  AND2_X1 U2702 ( .A1(b_10_), .A2(n2800), .ZN(n2798) );
  OR2_X1 U2703 ( .A1(n2693), .A2(n2345), .ZN(n2800) );
  OR2_X1 U2704 ( .A1(n2801), .A2(n2802), .ZN(n2345) );
  AND2_X1 U2705 ( .A1(n2317), .A2(n2697), .ZN(n2802) );
  AND2_X1 U2706 ( .A1(b_11_), .A2(n2803), .ZN(n2801) );
  OR2_X1 U2707 ( .A1(n2697), .A2(n2317), .ZN(n2803) );
  OR2_X1 U2708 ( .A1(n2804), .A2(n2805), .ZN(n2317) );
  AND2_X1 U2709 ( .A1(n2289), .A2(n2701), .ZN(n2805) );
  AND2_X1 U2710 ( .A1(b_12_), .A2(n2806), .ZN(n2804) );
  OR2_X1 U2711 ( .A1(n2701), .A2(n2289), .ZN(n2806) );
  OR2_X1 U2712 ( .A1(n2807), .A2(n2808), .ZN(n2289) );
  AND2_X1 U2713 ( .A1(n2261), .A2(n2705), .ZN(n2808) );
  AND2_X1 U2714 ( .A1(b_13_), .A2(n2809), .ZN(n2807) );
  OR2_X1 U2715 ( .A1(n2705), .A2(n2261), .ZN(n2809) );
  OR2_X1 U2716 ( .A1(n2218), .A2(n2810), .ZN(n2261) );
  AND2_X1 U2717 ( .A1(n2210), .A2(n2811), .ZN(n2810) );
  AND2_X1 U2718 ( .A1(n2812), .A2(b_15_), .ZN(n2210) );
  AND2_X1 U2719 ( .A1(n2654), .A2(operation_1_), .ZN(n2207) );
  INV_X1 U2720 ( .A(operation_0_), .ZN(n2654) );
  AND2_X1 U2721 ( .A1(n2813), .A2(n2208), .ZN(n2766) );
  AND2_X1 U2722 ( .A1(n2653), .A2(operation_0_), .ZN(n2208) );
  INV_X1 U2723 ( .A(operation_1_), .ZN(n2653) );
  AND2_X1 U2724 ( .A1(n2814), .A2(n2710), .ZN(n2813) );
  INV_X1 U2725 ( .A(n2770), .ZN(n2710) );
  AND2_X1 U2726 ( .A1(n2815), .A2(b_0_), .ZN(n2770) );
  INV_X1 U2727 ( .A(n2816), .ZN(n2814) );
  AND2_X1 U2728 ( .A1(n2711), .A2(n2642), .ZN(n2816) );
  INV_X1 U2729 ( .A(n2651), .ZN(n2642) );
  OR2_X1 U2730 ( .A1(n2817), .A2(n2818), .ZN(n2651) );
  AND2_X1 U2731 ( .A1(a_1_), .A2(n2613), .ZN(n2818) );
  AND2_X1 U2732 ( .A1(n2819), .A2(n2658), .ZN(n2817) );
  OR2_X1 U2733 ( .A1(a_1_), .A2(n2613), .ZN(n2819) );
  OR2_X1 U2734 ( .A1(n2820), .A2(n2821), .ZN(n2613) );
  AND2_X1 U2735 ( .A1(a_2_), .A2(n2584), .ZN(n2821) );
  AND2_X1 U2736 ( .A1(n2822), .A2(n2662), .ZN(n2820) );
  OR2_X1 U2737 ( .A1(a_2_), .A2(n2584), .ZN(n2822) );
  OR2_X1 U2738 ( .A1(n2823), .A2(n2824), .ZN(n2584) );
  AND2_X1 U2739 ( .A1(a_3_), .A2(n2555), .ZN(n2824) );
  AND2_X1 U2740 ( .A1(n2825), .A2(n2666), .ZN(n2823) );
  OR2_X1 U2741 ( .A1(a_3_), .A2(n2555), .ZN(n2825) );
  OR2_X1 U2742 ( .A1(n2826), .A2(n2827), .ZN(n2555) );
  AND2_X1 U2743 ( .A1(a_4_), .A2(n2515), .ZN(n2827) );
  AND2_X1 U2744 ( .A1(n2828), .A2(n2670), .ZN(n2826) );
  OR2_X1 U2745 ( .A1(a_4_), .A2(n2515), .ZN(n2828) );
  OR2_X1 U2746 ( .A1(n2829), .A2(n2830), .ZN(n2515) );
  AND2_X1 U2747 ( .A1(a_5_), .A2(n2486), .ZN(n2830) );
  AND2_X1 U2748 ( .A1(n2831), .A2(n2674), .ZN(n2829) );
  OR2_X1 U2749 ( .A1(a_5_), .A2(n2486), .ZN(n2831) );
  OR2_X1 U2750 ( .A1(n2832), .A2(n2833), .ZN(n2486) );
  AND2_X1 U2751 ( .A1(a_6_), .A2(n2457), .ZN(n2833) );
  AND2_X1 U2752 ( .A1(n2834), .A2(n2678), .ZN(n2832) );
  OR2_X1 U2753 ( .A1(a_6_), .A2(n2457), .ZN(n2834) );
  OR2_X1 U2754 ( .A1(n2835), .A2(n2836), .ZN(n2457) );
  AND2_X1 U2755 ( .A1(a_7_), .A2(n2428), .ZN(n2836) );
  AND2_X1 U2756 ( .A1(n2837), .A2(n2682), .ZN(n2835) );
  OR2_X1 U2757 ( .A1(a_7_), .A2(n2428), .ZN(n2837) );
  OR2_X1 U2758 ( .A1(n2838), .A2(n2839), .ZN(n2428) );
  AND2_X1 U2759 ( .A1(a_8_), .A2(n2399), .ZN(n2839) );
  AND2_X1 U2760 ( .A1(n2840), .A2(n2686), .ZN(n2838) );
  OR2_X1 U2761 ( .A1(a_8_), .A2(n2399), .ZN(n2840) );
  OR2_X1 U2762 ( .A1(n2841), .A2(n2842), .ZN(n2399) );
  AND2_X1 U2763 ( .A1(a_9_), .A2(n2370), .ZN(n2842) );
  AND2_X1 U2764 ( .A1(n2843), .A2(n2382), .ZN(n2841) );
  OR2_X1 U2765 ( .A1(a_9_), .A2(n2370), .ZN(n2843) );
  OR2_X1 U2766 ( .A1(n2844), .A2(n2845), .ZN(n2370) );
  AND2_X1 U2767 ( .A1(a_10_), .A2(n2342), .ZN(n2845) );
  AND2_X1 U2768 ( .A1(n2846), .A2(n2354), .ZN(n2844) );
  OR2_X1 U2769 ( .A1(a_10_), .A2(n2342), .ZN(n2846) );
  OR2_X1 U2770 ( .A1(n2847), .A2(n2848), .ZN(n2342) );
  AND2_X1 U2771 ( .A1(a_11_), .A2(n2314), .ZN(n2848) );
  AND2_X1 U2772 ( .A1(n2849), .A2(n2326), .ZN(n2847) );
  OR2_X1 U2773 ( .A1(a_11_), .A2(n2314), .ZN(n2849) );
  OR2_X1 U2774 ( .A1(n2850), .A2(n2851), .ZN(n2314) );
  AND2_X1 U2775 ( .A1(a_12_), .A2(n2286), .ZN(n2851) );
  AND2_X1 U2776 ( .A1(n2852), .A2(n2298), .ZN(n2850) );
  OR2_X1 U2777 ( .A1(a_12_), .A2(n2286), .ZN(n2852) );
  OR2_X1 U2778 ( .A1(n2853), .A2(n2854), .ZN(n2286) );
  AND2_X1 U2779 ( .A1(a_13_), .A2(n2258), .ZN(n2854) );
  AND2_X1 U2780 ( .A1(n2855), .A2(n2270), .ZN(n2853) );
  OR2_X1 U2781 ( .A1(a_13_), .A2(n2258), .ZN(n2855) );
  INV_X1 U2782 ( .A(n2268), .ZN(n2258) );
  AND2_X1 U2783 ( .A1(n2856), .A2(n2811), .ZN(n2268) );
  OR2_X1 U2784 ( .A1(b_14_), .A2(n2239), .ZN(n2811) );
  OR2_X1 U2785 ( .A1(n2234), .A2(n2218), .ZN(n2856) );
  AND2_X1 U2786 ( .A1(n2239), .A2(b_14_), .ZN(n2218) );
  INV_X1 U2787 ( .A(n2209), .ZN(n2234) );
  AND2_X1 U2788 ( .A1(n2857), .A2(a_15_), .ZN(n2209) );
  OR2_X1 U2789 ( .A1(b_0_), .A2(n2815), .ZN(n2711) );
  AND2_X1 U2790 ( .A1(n2173), .A2(n2858), .ZN(n2765) );
  OR2_X1 U2791 ( .A1(n2859), .A2(n2860), .ZN(n2858) );
  OR2_X1 U2792 ( .A1(n2543), .A2(n2861), .ZN(n2860) );
  AND2_X1 U2793 ( .A1(n2535), .A2(n2540), .ZN(n2861) );
  AND2_X1 U2794 ( .A1(n2246), .A2(n2247), .ZN(n2535) );
  XNOR2_X1 U2795 ( .A(n2542), .B(n2862), .ZN(n2247) );
  OR2_X1 U2796 ( .A1(n2863), .A2(n2864), .ZN(n2246) );
  AND2_X1 U2797 ( .A1(n2198), .A2(n2199), .ZN(n2864) );
  INV_X1 U2798 ( .A(n2865), .ZN(n2199) );
  OR2_X1 U2799 ( .A1(n2866), .A2(n2863), .ZN(n2865) );
  AND2_X1 U2800 ( .A1(n2867), .A2(n2868), .ZN(n2866) );
  OR2_X1 U2801 ( .A1(n2869), .A2(n2870), .ZN(n2198) );
  AND2_X1 U2802 ( .A1(n2194), .A2(n2195), .ZN(n2869) );
  INV_X1 U2803 ( .A(n2871), .ZN(n2195) );
  OR2_X1 U2804 ( .A1(n2872), .A2(n2870), .ZN(n2871) );
  INV_X1 U2805 ( .A(n2873), .ZN(n2870) );
  OR2_X1 U2806 ( .A1(n2874), .A2(n2875), .ZN(n2873) );
  AND2_X1 U2807 ( .A1(n2874), .A2(n2875), .ZN(n2872) );
  OR2_X1 U2808 ( .A1(n2876), .A2(n2877), .ZN(n2875) );
  AND2_X1 U2809 ( .A1(n2878), .A2(n2879), .ZN(n2877) );
  AND2_X1 U2810 ( .A1(n2880), .A2(n2881), .ZN(n2876) );
  OR2_X1 U2811 ( .A1(n2879), .A2(n2878), .ZN(n2881) );
  XOR2_X1 U2812 ( .A(n2882), .B(n2883), .Z(n2874) );
  XOR2_X1 U2813 ( .A(n2884), .B(n2885), .Z(n2883) );
  OR2_X1 U2814 ( .A1(n2886), .A2(n2887), .ZN(n2194) );
  AND2_X1 U2815 ( .A1(n2190), .A2(n2191), .ZN(n2887) );
  INV_X1 U2816 ( .A(n2888), .ZN(n2191) );
  OR2_X1 U2817 ( .A1(n2889), .A2(n2886), .ZN(n2888) );
  AND2_X1 U2818 ( .A1(n2890), .A2(n2891), .ZN(n2889) );
  OR2_X1 U2819 ( .A1(n2892), .A2(n2893), .ZN(n2190) );
  AND2_X1 U2820 ( .A1(n2186), .A2(n2187), .ZN(n2892) );
  INV_X1 U2821 ( .A(n2894), .ZN(n2187) );
  OR2_X1 U2822 ( .A1(n2895), .A2(n2893), .ZN(n2894) );
  INV_X1 U2823 ( .A(n2896), .ZN(n2893) );
  OR2_X1 U2824 ( .A1(n2897), .A2(n2898), .ZN(n2896) );
  AND2_X1 U2825 ( .A1(n2897), .A2(n2898), .ZN(n2895) );
  OR2_X1 U2826 ( .A1(n2899), .A2(n2900), .ZN(n2898) );
  AND2_X1 U2827 ( .A1(n2901), .A2(n2902), .ZN(n2900) );
  AND2_X1 U2828 ( .A1(n2903), .A2(n2904), .ZN(n2899) );
  OR2_X1 U2829 ( .A1(n2902), .A2(n2901), .ZN(n2904) );
  XOR2_X1 U2830 ( .A(n2905), .B(n2906), .Z(n2897) );
  XOR2_X1 U2831 ( .A(n2907), .B(n2908), .Z(n2906) );
  OR2_X1 U2832 ( .A1(n2909), .A2(n2910), .ZN(n2186) );
  AND2_X1 U2833 ( .A1(n2182), .A2(n2183), .ZN(n2910) );
  INV_X1 U2834 ( .A(n2911), .ZN(n2183) );
  OR2_X1 U2835 ( .A1(n2912), .A2(n2909), .ZN(n2911) );
  AND2_X1 U2836 ( .A1(n2913), .A2(n2914), .ZN(n2912) );
  OR2_X1 U2837 ( .A1(n2915), .A2(n2916), .ZN(n2182) );
  AND2_X1 U2838 ( .A1(n2178), .A2(n2179), .ZN(n2915) );
  INV_X1 U2839 ( .A(n2917), .ZN(n2179) );
  OR2_X1 U2840 ( .A1(n2918), .A2(n2916), .ZN(n2917) );
  INV_X1 U2841 ( .A(n2919), .ZN(n2916) );
  OR2_X1 U2842 ( .A1(n2920), .A2(n2921), .ZN(n2919) );
  AND2_X1 U2843 ( .A1(n2920), .A2(n2921), .ZN(n2918) );
  OR2_X1 U2844 ( .A1(n2922), .A2(n2923), .ZN(n2921) );
  AND2_X1 U2845 ( .A1(n2924), .A2(n2925), .ZN(n2923) );
  AND2_X1 U2846 ( .A1(n2926), .A2(n2927), .ZN(n2922) );
  OR2_X1 U2847 ( .A1(n2925), .A2(n2924), .ZN(n2927) );
  XOR2_X1 U2848 ( .A(n2928), .B(n2929), .Z(n2920) );
  XOR2_X1 U2849 ( .A(n2930), .B(n2931), .Z(n2929) );
  OR2_X1 U2850 ( .A1(n2932), .A2(n2933), .ZN(n2178) );
  AND2_X1 U2851 ( .A1(n2174), .A2(n2175), .ZN(n2933) );
  INV_X1 U2852 ( .A(n2934), .ZN(n2175) );
  OR2_X1 U2853 ( .A1(n2935), .A2(n2932), .ZN(n2934) );
  AND2_X1 U2854 ( .A1(n2936), .A2(n2937), .ZN(n2935) );
  OR2_X1 U2855 ( .A1(n2938), .A2(n2939), .ZN(n2174) );
  OR2_X1 U2856 ( .A1(n2940), .A2(n2764), .ZN(n2938) );
  AND2_X1 U2857 ( .A1(n2762), .A2(n2763), .ZN(n2764) );
  AND2_X1 U2858 ( .A1(n2941), .A2(n2942), .ZN(n2763) );
  INV_X1 U2859 ( .A(n2943), .ZN(n2941) );
  AND2_X1 U2860 ( .A1(n2762), .A2(n2758), .ZN(n2940) );
  OR2_X1 U2861 ( .A1(n2944), .A2(n2755), .ZN(n2758) );
  AND2_X1 U2862 ( .A1(n2753), .A2(n2945), .ZN(n2755) );
  AND2_X1 U2863 ( .A1(n2754), .A2(n2752), .ZN(n2945) );
  INV_X1 U2864 ( .A(n2946), .ZN(n2753) );
  AND2_X1 U2865 ( .A1(n2752), .A2(n2747), .ZN(n2944) );
  OR2_X1 U2866 ( .A1(n2947), .A2(n2744), .ZN(n2747) );
  AND2_X1 U2867 ( .A1(n2743), .A2(n2742), .ZN(n2744) );
  AND2_X1 U2868 ( .A1(n2743), .A2(n2738), .ZN(n2947) );
  OR2_X1 U2869 ( .A1(n2948), .A2(n2731), .ZN(n2738) );
  AND2_X1 U2870 ( .A1(n2949), .A2(n2950), .ZN(n2731) );
  INV_X1 U2871 ( .A(n2734), .ZN(n2950) );
  OR2_X1 U2872 ( .A1(n2951), .A2(n2952), .ZN(n2734) );
  AND2_X1 U2873 ( .A1(n2735), .A2(n2949), .ZN(n2948) );
  INV_X1 U2874 ( .A(n2733), .ZN(n2949) );
  OR2_X1 U2875 ( .A1(n2953), .A2(n2742), .ZN(n2733) );
  INV_X1 U2876 ( .A(n2954), .ZN(n2742) );
  OR2_X1 U2877 ( .A1(n2955), .A2(n2956), .ZN(n2954) );
  AND2_X1 U2878 ( .A1(n2955), .A2(n2956), .ZN(n2953) );
  OR2_X1 U2879 ( .A1(n2957), .A2(n2958), .ZN(n2956) );
  AND2_X1 U2880 ( .A1(n2959), .A2(n2960), .ZN(n2958) );
  AND2_X1 U2881 ( .A1(n2961), .A2(n2962), .ZN(n2957) );
  OR2_X1 U2882 ( .A1(n2960), .A2(n2959), .ZN(n2962) );
  XOR2_X1 U2883 ( .A(n2963), .B(n2964), .Z(n2955) );
  XOR2_X1 U2884 ( .A(n2965), .B(n2966), .Z(n2964) );
  AND2_X1 U2885 ( .A1(n2727), .A2(n2967), .ZN(n2735) );
  AND2_X1 U2886 ( .A1(n2720), .A2(n2726), .ZN(n2967) );
  XOR2_X1 U2887 ( .A(n2952), .B(n2951), .Z(n2726) );
  OR2_X1 U2888 ( .A1(n2968), .A2(n2969), .ZN(n2951) );
  AND2_X1 U2889 ( .A1(n2970), .A2(n2971), .ZN(n2969) );
  AND2_X1 U2890 ( .A1(n2972), .A2(n2973), .ZN(n2968) );
  OR2_X1 U2891 ( .A1(n2970), .A2(n2971), .ZN(n2973) );
  XOR2_X1 U2892 ( .A(n2961), .B(n2974), .Z(n2952) );
  XOR2_X1 U2893 ( .A(n2960), .B(n2959), .Z(n2974) );
  OR2_X1 U2894 ( .A1(n2815), .A2(n2270), .ZN(n2959) );
  OR2_X1 U2895 ( .A1(n2975), .A2(n2976), .ZN(n2960) );
  AND2_X1 U2896 ( .A1(n2977), .A2(n2978), .ZN(n2976) );
  AND2_X1 U2897 ( .A1(n2979), .A2(n2980), .ZN(n2975) );
  OR2_X1 U2898 ( .A1(n2978), .A2(n2977), .ZN(n2980) );
  XOR2_X1 U2899 ( .A(n2981), .B(n2982), .Z(n2961) );
  XOR2_X1 U2900 ( .A(n2983), .B(n2984), .Z(n2982) );
  XNOR2_X1 U2901 ( .A(n2972), .B(n2985), .ZN(n2720) );
  XOR2_X1 U2902 ( .A(n2971), .B(n2970), .Z(n2985) );
  OR2_X1 U2903 ( .A1(n2228), .A2(n2815), .ZN(n2970) );
  OR2_X1 U2904 ( .A1(n2986), .A2(n2987), .ZN(n2971) );
  AND2_X1 U2905 ( .A1(n2988), .A2(n2989), .ZN(n2987) );
  AND2_X1 U2906 ( .A1(n2990), .A2(n2991), .ZN(n2986) );
  OR2_X1 U2907 ( .A1(n2989), .A2(n2988), .ZN(n2991) );
  XOR2_X1 U2908 ( .A(n2979), .B(n2992), .Z(n2972) );
  XOR2_X1 U2909 ( .A(n2978), .B(n2977), .Z(n2992) );
  OR2_X1 U2910 ( .A1(n2657), .A2(n2270), .ZN(n2977) );
  OR2_X1 U2911 ( .A1(n2993), .A2(n2994), .ZN(n2978) );
  AND2_X1 U2912 ( .A1(n2995), .A2(n2996), .ZN(n2994) );
  AND2_X1 U2913 ( .A1(n2997), .A2(n2998), .ZN(n2993) );
  OR2_X1 U2914 ( .A1(n2996), .A2(n2995), .ZN(n2998) );
  XOR2_X1 U2915 ( .A(n2999), .B(n3000), .Z(n2979) );
  XOR2_X1 U2916 ( .A(n3001), .B(n3002), .Z(n3000) );
  INV_X1 U2917 ( .A(n2719), .ZN(n2727) );
  OR2_X1 U2918 ( .A1(n3003), .A2(n3004), .ZN(n2719) );
  AND2_X1 U2919 ( .A1(n2716), .A2(n2715), .ZN(n3004) );
  AND2_X1 U2920 ( .A1(n2713), .A2(n3005), .ZN(n3003) );
  OR2_X1 U2921 ( .A1(n2716), .A2(n2715), .ZN(n3005) );
  OR2_X1 U2922 ( .A1(n3006), .A2(n3007), .ZN(n2715) );
  AND2_X1 U2923 ( .A1(n2630), .A2(n2629), .ZN(n3007) );
  AND2_X1 U2924 ( .A1(n2627), .A2(n3008), .ZN(n3006) );
  OR2_X1 U2925 ( .A1(n2630), .A2(n2629), .ZN(n3008) );
  OR2_X1 U2926 ( .A1(n3009), .A2(n3010), .ZN(n2629) );
  AND2_X1 U2927 ( .A1(n2601), .A2(n2600), .ZN(n3010) );
  AND2_X1 U2928 ( .A1(n2598), .A2(n3011), .ZN(n3009) );
  OR2_X1 U2929 ( .A1(n2601), .A2(n2600), .ZN(n3011) );
  OR2_X1 U2930 ( .A1(n3012), .A2(n3013), .ZN(n2600) );
  AND2_X1 U2931 ( .A1(n2572), .A2(n2571), .ZN(n3013) );
  AND2_X1 U2932 ( .A1(n2569), .A2(n3014), .ZN(n3012) );
  OR2_X1 U2933 ( .A1(n2572), .A2(n2571), .ZN(n3014) );
  OR2_X1 U2934 ( .A1(n3015), .A2(n3016), .ZN(n2571) );
  AND2_X1 U2935 ( .A1(n2532), .A2(n2531), .ZN(n3016) );
  AND2_X1 U2936 ( .A1(n2529), .A2(n3017), .ZN(n3015) );
  OR2_X1 U2937 ( .A1(n2532), .A2(n2531), .ZN(n3017) );
  OR2_X1 U2938 ( .A1(n3018), .A2(n3019), .ZN(n2531) );
  AND2_X1 U2939 ( .A1(n2503), .A2(n2502), .ZN(n3019) );
  AND2_X1 U2940 ( .A1(n2500), .A2(n3020), .ZN(n3018) );
  OR2_X1 U2941 ( .A1(n2503), .A2(n2502), .ZN(n3020) );
  OR2_X1 U2942 ( .A1(n3021), .A2(n3022), .ZN(n2502) );
  AND2_X1 U2943 ( .A1(n2474), .A2(n2473), .ZN(n3022) );
  AND2_X1 U2944 ( .A1(n2471), .A2(n3023), .ZN(n3021) );
  OR2_X1 U2945 ( .A1(n2474), .A2(n2473), .ZN(n3023) );
  OR2_X1 U2946 ( .A1(n3024), .A2(n3025), .ZN(n2473) );
  AND2_X1 U2947 ( .A1(n2445), .A2(n2444), .ZN(n3025) );
  AND2_X1 U2948 ( .A1(n2442), .A2(n3026), .ZN(n3024) );
  OR2_X1 U2949 ( .A1(n2445), .A2(n2444), .ZN(n3026) );
  OR2_X1 U2950 ( .A1(n3027), .A2(n3028), .ZN(n2444) );
  AND2_X1 U2951 ( .A1(n2416), .A2(n2415), .ZN(n3028) );
  AND2_X1 U2952 ( .A1(n2413), .A2(n3029), .ZN(n3027) );
  OR2_X1 U2953 ( .A1(n2416), .A2(n2415), .ZN(n3029) );
  OR2_X1 U2954 ( .A1(n3030), .A2(n3031), .ZN(n2415) );
  AND2_X1 U2955 ( .A1(n2387), .A2(n2386), .ZN(n3031) );
  AND2_X1 U2956 ( .A1(n2384), .A2(n3032), .ZN(n3030) );
  OR2_X1 U2957 ( .A1(n2387), .A2(n2386), .ZN(n3032) );
  OR2_X1 U2958 ( .A1(n3033), .A2(n3034), .ZN(n2386) );
  AND2_X1 U2959 ( .A1(n2359), .A2(n2358), .ZN(n3034) );
  AND2_X1 U2960 ( .A1(n2356), .A2(n3035), .ZN(n3033) );
  OR2_X1 U2961 ( .A1(n2359), .A2(n2358), .ZN(n3035) );
  OR2_X1 U2962 ( .A1(n3036), .A2(n3037), .ZN(n2358) );
  AND2_X1 U2963 ( .A1(n2331), .A2(n2330), .ZN(n3037) );
  AND2_X1 U2964 ( .A1(n2328), .A2(n3038), .ZN(n3036) );
  OR2_X1 U2965 ( .A1(n2331), .A2(n2330), .ZN(n3038) );
  OR2_X1 U2966 ( .A1(n3039), .A2(n3040), .ZN(n2330) );
  AND2_X1 U2967 ( .A1(n2303), .A2(n2302), .ZN(n3040) );
  AND2_X1 U2968 ( .A1(n2300), .A2(n3041), .ZN(n3039) );
  OR2_X1 U2969 ( .A1(n2303), .A2(n2302), .ZN(n3041) );
  OR2_X1 U2970 ( .A1(n3042), .A2(n3043), .ZN(n2302) );
  AND2_X1 U2971 ( .A1(n2272), .A2(n2275), .ZN(n3043) );
  AND2_X1 U2972 ( .A1(n2274), .A2(n3044), .ZN(n3042) );
  OR2_X1 U2973 ( .A1(n2272), .A2(n2275), .ZN(n3044) );
  OR2_X1 U2974 ( .A1(n2705), .A2(n2857), .ZN(n2275) );
  OR2_X1 U2975 ( .A1(n2228), .A2(n2707), .ZN(n2272) );
  OR2_X1 U2976 ( .A1(n2857), .A2(n3045), .ZN(n2707) );
  INV_X1 U2977 ( .A(n3046), .ZN(n2274) );
  OR2_X1 U2978 ( .A1(n3047), .A2(n3048), .ZN(n3046) );
  AND2_X1 U2979 ( .A1(b_14_), .A2(n3049), .ZN(n3048) );
  OR2_X1 U2980 ( .A1(n3050), .A2(n3051), .ZN(n3049) );
  AND2_X1 U2981 ( .A1(a_14_), .A2(n2270), .ZN(n3050) );
  AND2_X1 U2982 ( .A1(b_13_), .A2(n3052), .ZN(n3047) );
  OR2_X1 U2983 ( .A1(n3053), .A2(n2217), .ZN(n3052) );
  AND2_X1 U2984 ( .A1(a_15_), .A2(n2228), .ZN(n3053) );
  OR2_X1 U2985 ( .A1(n2701), .A2(n2857), .ZN(n2303) );
  XNOR2_X1 U2986 ( .A(n3054), .B(n3055), .ZN(n2300) );
  XNOR2_X1 U2987 ( .A(n3056), .B(n3057), .ZN(n3055) );
  OR2_X1 U2988 ( .A1(n2697), .A2(n2857), .ZN(n2331) );
  XNOR2_X1 U2989 ( .A(n3058), .B(n3059), .ZN(n2328) );
  XNOR2_X1 U2990 ( .A(n3060), .B(n3061), .ZN(n3058) );
  OR2_X1 U2991 ( .A1(n2693), .A2(n2857), .ZN(n2359) );
  XOR2_X1 U2992 ( .A(n3062), .B(n3063), .Z(n2356) );
  XOR2_X1 U2993 ( .A(n3064), .B(n3065), .Z(n3063) );
  OR2_X1 U2994 ( .A1(n2689), .A2(n2857), .ZN(n2387) );
  XOR2_X1 U2995 ( .A(n3066), .B(n3067), .Z(n2384) );
  XOR2_X1 U2996 ( .A(n3068), .B(n3069), .Z(n3067) );
  OR2_X1 U2997 ( .A1(n2685), .A2(n2857), .ZN(n2416) );
  XOR2_X1 U2998 ( .A(n3070), .B(n3071), .Z(n2413) );
  XOR2_X1 U2999 ( .A(n3072), .B(n3073), .Z(n3071) );
  OR2_X1 U3000 ( .A1(n2681), .A2(n2857), .ZN(n2445) );
  XOR2_X1 U3001 ( .A(n3074), .B(n3075), .Z(n2442) );
  XOR2_X1 U3002 ( .A(n3076), .B(n3077), .Z(n3075) );
  OR2_X1 U3003 ( .A1(n2677), .A2(n2857), .ZN(n2474) );
  XOR2_X1 U3004 ( .A(n3078), .B(n3079), .Z(n2471) );
  XOR2_X1 U3005 ( .A(n3080), .B(n3081), .Z(n3079) );
  OR2_X1 U3006 ( .A1(n2673), .A2(n2857), .ZN(n2503) );
  XOR2_X1 U3007 ( .A(n3082), .B(n3083), .Z(n2500) );
  XOR2_X1 U3008 ( .A(n3084), .B(n3085), .Z(n3083) );
  OR2_X1 U3009 ( .A1(n2669), .A2(n2857), .ZN(n2532) );
  XOR2_X1 U3010 ( .A(n3086), .B(n3087), .Z(n2529) );
  XOR2_X1 U3011 ( .A(n3088), .B(n3089), .Z(n3087) );
  OR2_X1 U3012 ( .A1(n2665), .A2(n2857), .ZN(n2572) );
  XOR2_X1 U3013 ( .A(n3090), .B(n3091), .Z(n2569) );
  XOR2_X1 U3014 ( .A(n3092), .B(n3093), .Z(n3091) );
  OR2_X1 U3015 ( .A1(n2661), .A2(n2857), .ZN(n2601) );
  XOR2_X1 U3016 ( .A(n3094), .B(n3095), .Z(n2598) );
  XOR2_X1 U3017 ( .A(n3096), .B(n3097), .Z(n3095) );
  OR2_X1 U3018 ( .A1(n2657), .A2(n2857), .ZN(n2630) );
  XOR2_X1 U3019 ( .A(n3098), .B(n3099), .Z(n2627) );
  XOR2_X1 U3020 ( .A(n3100), .B(n3101), .Z(n3099) );
  OR2_X1 U3021 ( .A1(n2815), .A2(n2857), .ZN(n2716) );
  INV_X1 U3022 ( .A(b_15_), .ZN(n2857) );
  XOR2_X1 U3023 ( .A(n2990), .B(n3102), .Z(n2713) );
  XOR2_X1 U3024 ( .A(n2989), .B(n2988), .Z(n3102) );
  OR2_X1 U3025 ( .A1(n2228), .A2(n2657), .ZN(n2988) );
  OR2_X1 U3026 ( .A1(n3103), .A2(n3104), .ZN(n2989) );
  AND2_X1 U3027 ( .A1(n3101), .A2(n3100), .ZN(n3104) );
  AND2_X1 U3028 ( .A1(n3098), .A2(n3105), .ZN(n3103) );
  OR2_X1 U3029 ( .A1(n3100), .A2(n3101), .ZN(n3105) );
  OR2_X1 U3030 ( .A1(n2228), .A2(n2661), .ZN(n3101) );
  OR2_X1 U3031 ( .A1(n3106), .A2(n3107), .ZN(n3100) );
  AND2_X1 U3032 ( .A1(n3097), .A2(n3096), .ZN(n3107) );
  AND2_X1 U3033 ( .A1(n3094), .A2(n3108), .ZN(n3106) );
  OR2_X1 U3034 ( .A1(n3096), .A2(n3097), .ZN(n3108) );
  OR2_X1 U3035 ( .A1(n2228), .A2(n2665), .ZN(n3097) );
  OR2_X1 U3036 ( .A1(n3109), .A2(n3110), .ZN(n3096) );
  AND2_X1 U3037 ( .A1(n3093), .A2(n3092), .ZN(n3110) );
  AND2_X1 U3038 ( .A1(n3090), .A2(n3111), .ZN(n3109) );
  OR2_X1 U3039 ( .A1(n3092), .A2(n3093), .ZN(n3111) );
  OR2_X1 U3040 ( .A1(n2228), .A2(n2669), .ZN(n3093) );
  OR2_X1 U3041 ( .A1(n3112), .A2(n3113), .ZN(n3092) );
  AND2_X1 U3042 ( .A1(n3089), .A2(n3088), .ZN(n3113) );
  AND2_X1 U3043 ( .A1(n3086), .A2(n3114), .ZN(n3112) );
  OR2_X1 U3044 ( .A1(n3088), .A2(n3089), .ZN(n3114) );
  OR2_X1 U3045 ( .A1(n2228), .A2(n2673), .ZN(n3089) );
  OR2_X1 U3046 ( .A1(n3115), .A2(n3116), .ZN(n3088) );
  AND2_X1 U3047 ( .A1(n3085), .A2(n3084), .ZN(n3116) );
  AND2_X1 U3048 ( .A1(n3082), .A2(n3117), .ZN(n3115) );
  OR2_X1 U3049 ( .A1(n3084), .A2(n3085), .ZN(n3117) );
  OR2_X1 U3050 ( .A1(n2228), .A2(n2677), .ZN(n3085) );
  OR2_X1 U3051 ( .A1(n3118), .A2(n3119), .ZN(n3084) );
  AND2_X1 U3052 ( .A1(n3081), .A2(n3080), .ZN(n3119) );
  AND2_X1 U3053 ( .A1(n3078), .A2(n3120), .ZN(n3118) );
  OR2_X1 U3054 ( .A1(n3080), .A2(n3081), .ZN(n3120) );
  OR2_X1 U3055 ( .A1(n2228), .A2(n2681), .ZN(n3081) );
  OR2_X1 U3056 ( .A1(n3121), .A2(n3122), .ZN(n3080) );
  AND2_X1 U3057 ( .A1(n3077), .A2(n3076), .ZN(n3122) );
  AND2_X1 U3058 ( .A1(n3074), .A2(n3123), .ZN(n3121) );
  OR2_X1 U3059 ( .A1(n3076), .A2(n3077), .ZN(n3123) );
  OR2_X1 U3060 ( .A1(n2228), .A2(n2685), .ZN(n3077) );
  OR2_X1 U3061 ( .A1(n3124), .A2(n3125), .ZN(n3076) );
  AND2_X1 U3062 ( .A1(n3073), .A2(n3072), .ZN(n3125) );
  AND2_X1 U3063 ( .A1(n3070), .A2(n3126), .ZN(n3124) );
  OR2_X1 U3064 ( .A1(n3072), .A2(n3073), .ZN(n3126) );
  OR2_X1 U3065 ( .A1(n2228), .A2(n2689), .ZN(n3073) );
  OR2_X1 U3066 ( .A1(n3127), .A2(n3128), .ZN(n3072) );
  AND2_X1 U3067 ( .A1(n3069), .A2(n3068), .ZN(n3128) );
  AND2_X1 U3068 ( .A1(n3066), .A2(n3129), .ZN(n3127) );
  OR2_X1 U3069 ( .A1(n3068), .A2(n3069), .ZN(n3129) );
  OR2_X1 U3070 ( .A1(n2228), .A2(n2693), .ZN(n3069) );
  OR2_X1 U3071 ( .A1(n3130), .A2(n3131), .ZN(n3068) );
  AND2_X1 U3072 ( .A1(n3065), .A2(n3064), .ZN(n3131) );
  AND2_X1 U3073 ( .A1(n3062), .A2(n3132), .ZN(n3130) );
  OR2_X1 U3074 ( .A1(n3064), .A2(n3065), .ZN(n3132) );
  OR2_X1 U3075 ( .A1(n2228), .A2(n2697), .ZN(n3065) );
  OR2_X1 U3076 ( .A1(n3133), .A2(n3134), .ZN(n3064) );
  AND2_X1 U3077 ( .A1(n3061), .A2(n3060), .ZN(n3134) );
  AND2_X1 U3078 ( .A1(n3059), .A2(n3135), .ZN(n3133) );
  OR2_X1 U3079 ( .A1(n3060), .A2(n3061), .ZN(n3135) );
  OR2_X1 U3080 ( .A1(n2228), .A2(n2701), .ZN(n3061) );
  OR2_X1 U3081 ( .A1(n3136), .A2(n3137), .ZN(n3060) );
  AND2_X1 U3082 ( .A1(n3054), .A2(n3057), .ZN(n3137) );
  AND2_X1 U3083 ( .A1(n3056), .A2(n3138), .ZN(n3136) );
  OR2_X1 U3084 ( .A1(n3057), .A2(n3054), .ZN(n3138) );
  OR2_X1 U3085 ( .A1(n2228), .A2(n2705), .ZN(n3054) );
  OR2_X1 U3086 ( .A1(n3045), .A2(n3139), .ZN(n3057) );
  OR2_X1 U3087 ( .A1(n2228), .A2(n2270), .ZN(n3139) );
  INV_X1 U3088 ( .A(b_14_), .ZN(n2228) );
  INV_X1 U3089 ( .A(n3140), .ZN(n3056) );
  OR2_X1 U3090 ( .A1(n3141), .A2(n3142), .ZN(n3140) );
  AND2_X1 U3091 ( .A1(b_13_), .A2(n3143), .ZN(n3142) );
  OR2_X1 U3092 ( .A1(n3144), .A2(n3051), .ZN(n3143) );
  AND2_X1 U3093 ( .A1(a_14_), .A2(n2298), .ZN(n3144) );
  AND2_X1 U3094 ( .A1(b_12_), .A2(n3145), .ZN(n3141) );
  OR2_X1 U3095 ( .A1(n3146), .A2(n2217), .ZN(n3145) );
  AND2_X1 U3096 ( .A1(a_15_), .A2(n2270), .ZN(n3146) );
  XNOR2_X1 U3097 ( .A(n2706), .B(n3147), .ZN(n3059) );
  XNOR2_X1 U3098 ( .A(n3148), .B(n3149), .ZN(n3147) );
  XNOR2_X1 U3099 ( .A(n3150), .B(n3151), .ZN(n3062) );
  XNOR2_X1 U3100 ( .A(n3152), .B(n3153), .ZN(n3150) );
  XOR2_X1 U3101 ( .A(n3154), .B(n3155), .Z(n3066) );
  XOR2_X1 U3102 ( .A(n3156), .B(n3157), .Z(n3155) );
  XOR2_X1 U3103 ( .A(n3158), .B(n3159), .Z(n3070) );
  XOR2_X1 U3104 ( .A(n3160), .B(n3161), .Z(n3159) );
  XOR2_X1 U3105 ( .A(n3162), .B(n3163), .Z(n3074) );
  XOR2_X1 U3106 ( .A(n3164), .B(n3165), .Z(n3163) );
  XOR2_X1 U3107 ( .A(n3166), .B(n3167), .Z(n3078) );
  XOR2_X1 U3108 ( .A(n3168), .B(n3169), .Z(n3167) );
  XOR2_X1 U3109 ( .A(n3170), .B(n3171), .Z(n3082) );
  XOR2_X1 U3110 ( .A(n3172), .B(n3173), .Z(n3171) );
  XOR2_X1 U3111 ( .A(n3174), .B(n3175), .Z(n3086) );
  XOR2_X1 U3112 ( .A(n3176), .B(n3177), .Z(n3175) );
  XOR2_X1 U3113 ( .A(n3178), .B(n3179), .Z(n3090) );
  XOR2_X1 U3114 ( .A(n3180), .B(n3181), .Z(n3179) );
  XOR2_X1 U3115 ( .A(n3182), .B(n3183), .Z(n3094) );
  XOR2_X1 U3116 ( .A(n3184), .B(n3185), .Z(n3183) );
  XOR2_X1 U3117 ( .A(n3186), .B(n3187), .Z(n3098) );
  XOR2_X1 U3118 ( .A(n3188), .B(n3189), .Z(n3187) );
  XOR2_X1 U3119 ( .A(n2997), .B(n3190), .Z(n2990) );
  XOR2_X1 U3120 ( .A(n2996), .B(n2995), .Z(n3190) );
  OR2_X1 U3121 ( .A1(n2661), .A2(n2270), .ZN(n2995) );
  OR2_X1 U3122 ( .A1(n3191), .A2(n3192), .ZN(n2996) );
  AND2_X1 U3123 ( .A1(n3189), .A2(n3188), .ZN(n3192) );
  AND2_X1 U3124 ( .A1(n3186), .A2(n3193), .ZN(n3191) );
  OR2_X1 U3125 ( .A1(n3188), .A2(n3189), .ZN(n3193) );
  OR2_X1 U3126 ( .A1(n2665), .A2(n2270), .ZN(n3189) );
  OR2_X1 U3127 ( .A1(n3194), .A2(n3195), .ZN(n3188) );
  AND2_X1 U3128 ( .A1(n3185), .A2(n3184), .ZN(n3195) );
  AND2_X1 U3129 ( .A1(n3182), .A2(n3196), .ZN(n3194) );
  OR2_X1 U3130 ( .A1(n3184), .A2(n3185), .ZN(n3196) );
  OR2_X1 U3131 ( .A1(n2669), .A2(n2270), .ZN(n3185) );
  OR2_X1 U3132 ( .A1(n3197), .A2(n3198), .ZN(n3184) );
  AND2_X1 U3133 ( .A1(n3181), .A2(n3180), .ZN(n3198) );
  AND2_X1 U3134 ( .A1(n3178), .A2(n3199), .ZN(n3197) );
  OR2_X1 U3135 ( .A1(n3180), .A2(n3181), .ZN(n3199) );
  OR2_X1 U3136 ( .A1(n2673), .A2(n2270), .ZN(n3181) );
  OR2_X1 U3137 ( .A1(n3200), .A2(n3201), .ZN(n3180) );
  AND2_X1 U3138 ( .A1(n3177), .A2(n3176), .ZN(n3201) );
  AND2_X1 U3139 ( .A1(n3174), .A2(n3202), .ZN(n3200) );
  OR2_X1 U3140 ( .A1(n3176), .A2(n3177), .ZN(n3202) );
  OR2_X1 U3141 ( .A1(n2677), .A2(n2270), .ZN(n3177) );
  OR2_X1 U3142 ( .A1(n3203), .A2(n3204), .ZN(n3176) );
  AND2_X1 U3143 ( .A1(n3173), .A2(n3172), .ZN(n3204) );
  AND2_X1 U3144 ( .A1(n3170), .A2(n3205), .ZN(n3203) );
  OR2_X1 U3145 ( .A1(n3172), .A2(n3173), .ZN(n3205) );
  OR2_X1 U3146 ( .A1(n2681), .A2(n2270), .ZN(n3173) );
  OR2_X1 U3147 ( .A1(n3206), .A2(n3207), .ZN(n3172) );
  AND2_X1 U3148 ( .A1(n3169), .A2(n3168), .ZN(n3207) );
  AND2_X1 U3149 ( .A1(n3166), .A2(n3208), .ZN(n3206) );
  OR2_X1 U3150 ( .A1(n3168), .A2(n3169), .ZN(n3208) );
  OR2_X1 U3151 ( .A1(n2685), .A2(n2270), .ZN(n3169) );
  OR2_X1 U3152 ( .A1(n3209), .A2(n3210), .ZN(n3168) );
  AND2_X1 U3153 ( .A1(n3165), .A2(n3164), .ZN(n3210) );
  AND2_X1 U3154 ( .A1(n3162), .A2(n3211), .ZN(n3209) );
  OR2_X1 U3155 ( .A1(n3164), .A2(n3165), .ZN(n3211) );
  OR2_X1 U3156 ( .A1(n2689), .A2(n2270), .ZN(n3165) );
  OR2_X1 U3157 ( .A1(n3212), .A2(n3213), .ZN(n3164) );
  AND2_X1 U3158 ( .A1(n3161), .A2(n3160), .ZN(n3213) );
  AND2_X1 U3159 ( .A1(n3158), .A2(n3214), .ZN(n3212) );
  OR2_X1 U3160 ( .A1(n3160), .A2(n3161), .ZN(n3214) );
  OR2_X1 U3161 ( .A1(n2693), .A2(n2270), .ZN(n3161) );
  OR2_X1 U3162 ( .A1(n3215), .A2(n3216), .ZN(n3160) );
  AND2_X1 U3163 ( .A1(n3157), .A2(n3156), .ZN(n3216) );
  AND2_X1 U3164 ( .A1(n3154), .A2(n3217), .ZN(n3215) );
  OR2_X1 U3165 ( .A1(n3156), .A2(n3157), .ZN(n3217) );
  OR2_X1 U3166 ( .A1(n2697), .A2(n2270), .ZN(n3157) );
  OR2_X1 U3167 ( .A1(n3218), .A2(n3219), .ZN(n3156) );
  AND2_X1 U3168 ( .A1(n3153), .A2(n3152), .ZN(n3219) );
  AND2_X1 U3169 ( .A1(n3151), .A2(n3220), .ZN(n3218) );
  OR2_X1 U3170 ( .A1(n3152), .A2(n3153), .ZN(n3220) );
  OR2_X1 U3171 ( .A1(n2701), .A2(n2270), .ZN(n3153) );
  OR2_X1 U3172 ( .A1(n3221), .A2(n3222), .ZN(n3152) );
  AND2_X1 U3173 ( .A1(n2706), .A2(n3149), .ZN(n3222) );
  AND2_X1 U3174 ( .A1(n3148), .A2(n3223), .ZN(n3221) );
  OR2_X1 U3175 ( .A1(n3149), .A2(n2706), .ZN(n3223) );
  OR2_X1 U3176 ( .A1(n2705), .A2(n2270), .ZN(n2706) );
  OR2_X1 U3177 ( .A1(n3045), .A2(n3224), .ZN(n3149) );
  OR2_X1 U3178 ( .A1(n2270), .A2(n2298), .ZN(n3224) );
  INV_X1 U3179 ( .A(b_13_), .ZN(n2270) );
  INV_X1 U3180 ( .A(n3225), .ZN(n3148) );
  OR2_X1 U3181 ( .A1(n3226), .A2(n3227), .ZN(n3225) );
  AND2_X1 U3182 ( .A1(b_12_), .A2(n3228), .ZN(n3227) );
  OR2_X1 U3183 ( .A1(n3229), .A2(n3051), .ZN(n3228) );
  AND2_X1 U3184 ( .A1(a_14_), .A2(n2326), .ZN(n3229) );
  AND2_X1 U3185 ( .A1(b_11_), .A2(n3230), .ZN(n3226) );
  OR2_X1 U3186 ( .A1(n3231), .A2(n2217), .ZN(n3230) );
  AND2_X1 U3187 ( .A1(a_15_), .A2(n2298), .ZN(n3231) );
  XNOR2_X1 U3188 ( .A(n3232), .B(n3233), .ZN(n3151) );
  XNOR2_X1 U3189 ( .A(n3234), .B(n3235), .ZN(n3233) );
  XNOR2_X1 U3190 ( .A(n3236), .B(n3237), .ZN(n3154) );
  XNOR2_X1 U3191 ( .A(n3238), .B(n2702), .ZN(n3236) );
  XOR2_X1 U3192 ( .A(n3239), .B(n3240), .Z(n3158) );
  XOR2_X1 U3193 ( .A(n3241), .B(n3242), .Z(n3240) );
  XOR2_X1 U3194 ( .A(n3243), .B(n3244), .Z(n3162) );
  XOR2_X1 U3195 ( .A(n3245), .B(n3246), .Z(n3244) );
  XOR2_X1 U3196 ( .A(n3247), .B(n3248), .Z(n3166) );
  XOR2_X1 U3197 ( .A(n3249), .B(n3250), .Z(n3248) );
  XOR2_X1 U3198 ( .A(n3251), .B(n3252), .Z(n3170) );
  XOR2_X1 U3199 ( .A(n3253), .B(n3254), .Z(n3252) );
  XOR2_X1 U3200 ( .A(n3255), .B(n3256), .Z(n3174) );
  XOR2_X1 U3201 ( .A(n3257), .B(n3258), .Z(n3256) );
  XOR2_X1 U3202 ( .A(n3259), .B(n3260), .Z(n3178) );
  XOR2_X1 U3203 ( .A(n3261), .B(n3262), .Z(n3260) );
  XOR2_X1 U3204 ( .A(n3263), .B(n3264), .Z(n3182) );
  XOR2_X1 U3205 ( .A(n3265), .B(n3266), .Z(n3264) );
  XOR2_X1 U3206 ( .A(n3267), .B(n3268), .Z(n3186) );
  XOR2_X1 U3207 ( .A(n3269), .B(n3270), .Z(n3268) );
  XOR2_X1 U3208 ( .A(n3271), .B(n3272), .Z(n2997) );
  XOR2_X1 U3209 ( .A(n3273), .B(n3274), .Z(n3272) );
  XNOR2_X1 U3210 ( .A(n2754), .B(n2946), .ZN(n2743) );
  OR2_X1 U3211 ( .A1(n3275), .A2(n3276), .ZN(n2946) );
  AND2_X1 U3212 ( .A1(n2966), .A2(n2965), .ZN(n3276) );
  AND2_X1 U3213 ( .A1(n2963), .A2(n3277), .ZN(n3275) );
  OR2_X1 U3214 ( .A1(n2965), .A2(n2966), .ZN(n3277) );
  OR2_X1 U3215 ( .A1(n2815), .A2(n2298), .ZN(n2966) );
  OR2_X1 U3216 ( .A1(n3278), .A2(n3279), .ZN(n2965) );
  AND2_X1 U3217 ( .A1(n2984), .A2(n2983), .ZN(n3279) );
  AND2_X1 U3218 ( .A1(n2981), .A2(n3280), .ZN(n3278) );
  OR2_X1 U3219 ( .A1(n2983), .A2(n2984), .ZN(n3280) );
  OR2_X1 U3220 ( .A1(n2657), .A2(n2298), .ZN(n2984) );
  OR2_X1 U3221 ( .A1(n3281), .A2(n3282), .ZN(n2983) );
  AND2_X1 U3222 ( .A1(n3002), .A2(n3001), .ZN(n3282) );
  AND2_X1 U3223 ( .A1(n2999), .A2(n3283), .ZN(n3281) );
  OR2_X1 U3224 ( .A1(n3001), .A2(n3002), .ZN(n3283) );
  OR2_X1 U3225 ( .A1(n2661), .A2(n2298), .ZN(n3002) );
  OR2_X1 U3226 ( .A1(n3284), .A2(n3285), .ZN(n3001) );
  AND2_X1 U3227 ( .A1(n3274), .A2(n3273), .ZN(n3285) );
  AND2_X1 U3228 ( .A1(n3271), .A2(n3286), .ZN(n3284) );
  OR2_X1 U3229 ( .A1(n3273), .A2(n3274), .ZN(n3286) );
  OR2_X1 U3230 ( .A1(n2665), .A2(n2298), .ZN(n3274) );
  OR2_X1 U3231 ( .A1(n3287), .A2(n3288), .ZN(n3273) );
  AND2_X1 U3232 ( .A1(n3270), .A2(n3269), .ZN(n3288) );
  AND2_X1 U3233 ( .A1(n3267), .A2(n3289), .ZN(n3287) );
  OR2_X1 U3234 ( .A1(n3269), .A2(n3270), .ZN(n3289) );
  OR2_X1 U3235 ( .A1(n2669), .A2(n2298), .ZN(n3270) );
  OR2_X1 U3236 ( .A1(n3290), .A2(n3291), .ZN(n3269) );
  AND2_X1 U3237 ( .A1(n3266), .A2(n3265), .ZN(n3291) );
  AND2_X1 U3238 ( .A1(n3263), .A2(n3292), .ZN(n3290) );
  OR2_X1 U3239 ( .A1(n3265), .A2(n3266), .ZN(n3292) );
  OR2_X1 U3240 ( .A1(n2673), .A2(n2298), .ZN(n3266) );
  OR2_X1 U3241 ( .A1(n3293), .A2(n3294), .ZN(n3265) );
  AND2_X1 U3242 ( .A1(n3262), .A2(n3261), .ZN(n3294) );
  AND2_X1 U3243 ( .A1(n3259), .A2(n3295), .ZN(n3293) );
  OR2_X1 U3244 ( .A1(n3261), .A2(n3262), .ZN(n3295) );
  OR2_X1 U3245 ( .A1(n2677), .A2(n2298), .ZN(n3262) );
  OR2_X1 U3246 ( .A1(n3296), .A2(n3297), .ZN(n3261) );
  AND2_X1 U3247 ( .A1(n3258), .A2(n3257), .ZN(n3297) );
  AND2_X1 U3248 ( .A1(n3255), .A2(n3298), .ZN(n3296) );
  OR2_X1 U3249 ( .A1(n3257), .A2(n3258), .ZN(n3298) );
  OR2_X1 U3250 ( .A1(n2681), .A2(n2298), .ZN(n3258) );
  OR2_X1 U3251 ( .A1(n3299), .A2(n3300), .ZN(n3257) );
  AND2_X1 U3252 ( .A1(n3254), .A2(n3253), .ZN(n3300) );
  AND2_X1 U3253 ( .A1(n3251), .A2(n3301), .ZN(n3299) );
  OR2_X1 U3254 ( .A1(n3253), .A2(n3254), .ZN(n3301) );
  OR2_X1 U3255 ( .A1(n2685), .A2(n2298), .ZN(n3254) );
  OR2_X1 U3256 ( .A1(n3302), .A2(n3303), .ZN(n3253) );
  AND2_X1 U3257 ( .A1(n3250), .A2(n3249), .ZN(n3303) );
  AND2_X1 U3258 ( .A1(n3247), .A2(n3304), .ZN(n3302) );
  OR2_X1 U3259 ( .A1(n3249), .A2(n3250), .ZN(n3304) );
  OR2_X1 U3260 ( .A1(n2689), .A2(n2298), .ZN(n3250) );
  OR2_X1 U3261 ( .A1(n3305), .A2(n3306), .ZN(n3249) );
  AND2_X1 U3262 ( .A1(n3246), .A2(n3245), .ZN(n3306) );
  AND2_X1 U3263 ( .A1(n3243), .A2(n3307), .ZN(n3305) );
  OR2_X1 U3264 ( .A1(n3245), .A2(n3246), .ZN(n3307) );
  OR2_X1 U3265 ( .A1(n2693), .A2(n2298), .ZN(n3246) );
  OR2_X1 U3266 ( .A1(n3308), .A2(n3309), .ZN(n3245) );
  AND2_X1 U3267 ( .A1(n3242), .A2(n3241), .ZN(n3309) );
  AND2_X1 U3268 ( .A1(n3239), .A2(n3310), .ZN(n3308) );
  OR2_X1 U3269 ( .A1(n3241), .A2(n3242), .ZN(n3310) );
  OR2_X1 U3270 ( .A1(n2697), .A2(n2298), .ZN(n3242) );
  OR2_X1 U3271 ( .A1(n3311), .A2(n3312), .ZN(n3241) );
  AND2_X1 U3272 ( .A1(n2702), .A2(n3238), .ZN(n3312) );
  AND2_X1 U3273 ( .A1(n3237), .A2(n3313), .ZN(n3311) );
  OR2_X1 U3274 ( .A1(n3238), .A2(n2702), .ZN(n3313) );
  OR2_X1 U3275 ( .A1(n2701), .A2(n2298), .ZN(n2702) );
  OR2_X1 U3276 ( .A1(n3314), .A2(n3315), .ZN(n3238) );
  AND2_X1 U3277 ( .A1(n3232), .A2(n3235), .ZN(n3315) );
  AND2_X1 U3278 ( .A1(n3234), .A2(n3316), .ZN(n3314) );
  OR2_X1 U3279 ( .A1(n3235), .A2(n3232), .ZN(n3316) );
  OR2_X1 U3280 ( .A1(n2705), .A2(n2298), .ZN(n3232) );
  OR2_X1 U3281 ( .A1(n3045), .A2(n3317), .ZN(n3235) );
  OR2_X1 U3282 ( .A1(n2298), .A2(n2326), .ZN(n3317) );
  INV_X1 U3283 ( .A(b_12_), .ZN(n2298) );
  INV_X1 U3284 ( .A(n3318), .ZN(n3234) );
  OR2_X1 U3285 ( .A1(n3319), .A2(n3320), .ZN(n3318) );
  AND2_X1 U3286 ( .A1(b_11_), .A2(n3321), .ZN(n3320) );
  OR2_X1 U3287 ( .A1(n3322), .A2(n3051), .ZN(n3321) );
  AND2_X1 U3288 ( .A1(a_14_), .A2(n2354), .ZN(n3322) );
  AND2_X1 U3289 ( .A1(b_10_), .A2(n3323), .ZN(n3319) );
  OR2_X1 U3290 ( .A1(n3324), .A2(n2217), .ZN(n3323) );
  AND2_X1 U3291 ( .A1(a_15_), .A2(n2326), .ZN(n3324) );
  XNOR2_X1 U3292 ( .A(n3325), .B(n3326), .ZN(n3237) );
  XNOR2_X1 U3293 ( .A(n3327), .B(n3328), .ZN(n3326) );
  XNOR2_X1 U3294 ( .A(n3329), .B(n3330), .ZN(n3239) );
  XNOR2_X1 U3295 ( .A(n3331), .B(n3332), .ZN(n3329) );
  XOR2_X1 U3296 ( .A(n3333), .B(n3334), .Z(n3243) );
  XOR2_X1 U3297 ( .A(n3335), .B(n2698), .Z(n3334) );
  XOR2_X1 U3298 ( .A(n3336), .B(n3337), .Z(n3247) );
  XOR2_X1 U3299 ( .A(n3338), .B(n3339), .Z(n3337) );
  XOR2_X1 U3300 ( .A(n3340), .B(n3341), .Z(n3251) );
  XOR2_X1 U3301 ( .A(n3342), .B(n3343), .Z(n3341) );
  XOR2_X1 U3302 ( .A(n3344), .B(n3345), .Z(n3255) );
  XOR2_X1 U3303 ( .A(n3346), .B(n3347), .Z(n3345) );
  XOR2_X1 U3304 ( .A(n3348), .B(n3349), .Z(n3259) );
  XOR2_X1 U3305 ( .A(n3350), .B(n3351), .Z(n3349) );
  XOR2_X1 U3306 ( .A(n3352), .B(n3353), .Z(n3263) );
  XOR2_X1 U3307 ( .A(n3354), .B(n3355), .Z(n3353) );
  XOR2_X1 U3308 ( .A(n3356), .B(n3357), .Z(n3267) );
  XOR2_X1 U3309 ( .A(n3358), .B(n3359), .Z(n3357) );
  XOR2_X1 U3310 ( .A(n3360), .B(n3361), .Z(n3271) );
  XOR2_X1 U3311 ( .A(n3362), .B(n3363), .Z(n3361) );
  XOR2_X1 U3312 ( .A(n3364), .B(n3365), .Z(n2999) );
  XOR2_X1 U3313 ( .A(n3366), .B(n3367), .Z(n3365) );
  XOR2_X1 U3314 ( .A(n3368), .B(n3369), .Z(n2981) );
  XOR2_X1 U3315 ( .A(n3370), .B(n3371), .Z(n3369) );
  XOR2_X1 U3316 ( .A(n3372), .B(n3373), .Z(n2963) );
  XOR2_X1 U3317 ( .A(n3374), .B(n3375), .Z(n3373) );
  XNOR2_X1 U3318 ( .A(n3376), .B(n3377), .ZN(n2754) );
  XOR2_X1 U3319 ( .A(n3378), .B(n3379), .Z(n3377) );
  XNOR2_X1 U3320 ( .A(n2942), .B(n2943), .ZN(n2752) );
  OR2_X1 U3321 ( .A1(n3380), .A2(n3381), .ZN(n2943) );
  AND2_X1 U3322 ( .A1(n3379), .A2(n3378), .ZN(n3381) );
  AND2_X1 U3323 ( .A1(n3376), .A2(n3382), .ZN(n3380) );
  OR2_X1 U3324 ( .A1(n3378), .A2(n3379), .ZN(n3382) );
  OR2_X1 U3325 ( .A1(n2815), .A2(n2326), .ZN(n3379) );
  OR2_X1 U3326 ( .A1(n3383), .A2(n3384), .ZN(n3378) );
  AND2_X1 U3327 ( .A1(n3375), .A2(n3374), .ZN(n3384) );
  AND2_X1 U3328 ( .A1(n3372), .A2(n3385), .ZN(n3383) );
  OR2_X1 U3329 ( .A1(n3374), .A2(n3375), .ZN(n3385) );
  OR2_X1 U3330 ( .A1(n2657), .A2(n2326), .ZN(n3375) );
  OR2_X1 U3331 ( .A1(n3386), .A2(n3387), .ZN(n3374) );
  AND2_X1 U3332 ( .A1(n3371), .A2(n3370), .ZN(n3387) );
  AND2_X1 U3333 ( .A1(n3368), .A2(n3388), .ZN(n3386) );
  OR2_X1 U3334 ( .A1(n3370), .A2(n3371), .ZN(n3388) );
  OR2_X1 U3335 ( .A1(n2661), .A2(n2326), .ZN(n3371) );
  OR2_X1 U3336 ( .A1(n3389), .A2(n3390), .ZN(n3370) );
  AND2_X1 U3337 ( .A1(n3367), .A2(n3366), .ZN(n3390) );
  AND2_X1 U3338 ( .A1(n3364), .A2(n3391), .ZN(n3389) );
  OR2_X1 U3339 ( .A1(n3366), .A2(n3367), .ZN(n3391) );
  OR2_X1 U3340 ( .A1(n2665), .A2(n2326), .ZN(n3367) );
  OR2_X1 U3341 ( .A1(n3392), .A2(n3393), .ZN(n3366) );
  AND2_X1 U3342 ( .A1(n3363), .A2(n3362), .ZN(n3393) );
  AND2_X1 U3343 ( .A1(n3360), .A2(n3394), .ZN(n3392) );
  OR2_X1 U3344 ( .A1(n3362), .A2(n3363), .ZN(n3394) );
  OR2_X1 U3345 ( .A1(n2669), .A2(n2326), .ZN(n3363) );
  OR2_X1 U3346 ( .A1(n3395), .A2(n3396), .ZN(n3362) );
  AND2_X1 U3347 ( .A1(n3359), .A2(n3358), .ZN(n3396) );
  AND2_X1 U3348 ( .A1(n3356), .A2(n3397), .ZN(n3395) );
  OR2_X1 U3349 ( .A1(n3358), .A2(n3359), .ZN(n3397) );
  OR2_X1 U3350 ( .A1(n2673), .A2(n2326), .ZN(n3359) );
  OR2_X1 U3351 ( .A1(n3398), .A2(n3399), .ZN(n3358) );
  AND2_X1 U3352 ( .A1(n3355), .A2(n3354), .ZN(n3399) );
  AND2_X1 U3353 ( .A1(n3352), .A2(n3400), .ZN(n3398) );
  OR2_X1 U3354 ( .A1(n3354), .A2(n3355), .ZN(n3400) );
  OR2_X1 U3355 ( .A1(n2677), .A2(n2326), .ZN(n3355) );
  OR2_X1 U3356 ( .A1(n3401), .A2(n3402), .ZN(n3354) );
  AND2_X1 U3357 ( .A1(n3351), .A2(n3350), .ZN(n3402) );
  AND2_X1 U3358 ( .A1(n3348), .A2(n3403), .ZN(n3401) );
  OR2_X1 U3359 ( .A1(n3350), .A2(n3351), .ZN(n3403) );
  OR2_X1 U3360 ( .A1(n2681), .A2(n2326), .ZN(n3351) );
  OR2_X1 U3361 ( .A1(n3404), .A2(n3405), .ZN(n3350) );
  AND2_X1 U3362 ( .A1(n3347), .A2(n3346), .ZN(n3405) );
  AND2_X1 U3363 ( .A1(n3344), .A2(n3406), .ZN(n3404) );
  OR2_X1 U3364 ( .A1(n3346), .A2(n3347), .ZN(n3406) );
  OR2_X1 U3365 ( .A1(n2685), .A2(n2326), .ZN(n3347) );
  OR2_X1 U3366 ( .A1(n3407), .A2(n3408), .ZN(n3346) );
  AND2_X1 U3367 ( .A1(n3343), .A2(n3342), .ZN(n3408) );
  AND2_X1 U3368 ( .A1(n3340), .A2(n3409), .ZN(n3407) );
  OR2_X1 U3369 ( .A1(n3342), .A2(n3343), .ZN(n3409) );
  OR2_X1 U3370 ( .A1(n2689), .A2(n2326), .ZN(n3343) );
  OR2_X1 U3371 ( .A1(n3410), .A2(n3411), .ZN(n3342) );
  AND2_X1 U3372 ( .A1(n3339), .A2(n3338), .ZN(n3411) );
  AND2_X1 U3373 ( .A1(n3336), .A2(n3412), .ZN(n3410) );
  OR2_X1 U3374 ( .A1(n3338), .A2(n3339), .ZN(n3412) );
  OR2_X1 U3375 ( .A1(n2693), .A2(n2326), .ZN(n3339) );
  OR2_X1 U3376 ( .A1(n3413), .A2(n3414), .ZN(n3338) );
  AND2_X1 U3377 ( .A1(n2698), .A2(n3335), .ZN(n3414) );
  AND2_X1 U3378 ( .A1(n3333), .A2(n3415), .ZN(n3413) );
  OR2_X1 U3379 ( .A1(n3335), .A2(n2698), .ZN(n3415) );
  OR2_X1 U3380 ( .A1(n2697), .A2(n2326), .ZN(n2698) );
  OR2_X1 U3381 ( .A1(n3416), .A2(n3417), .ZN(n3335) );
  AND2_X1 U3382 ( .A1(n3332), .A2(n3331), .ZN(n3417) );
  AND2_X1 U3383 ( .A1(n3330), .A2(n3418), .ZN(n3416) );
  OR2_X1 U3384 ( .A1(n3331), .A2(n3332), .ZN(n3418) );
  OR2_X1 U3385 ( .A1(n2701), .A2(n2326), .ZN(n3332) );
  OR2_X1 U3386 ( .A1(n3419), .A2(n3420), .ZN(n3331) );
  AND2_X1 U3387 ( .A1(n3325), .A2(n3328), .ZN(n3420) );
  AND2_X1 U3388 ( .A1(n3327), .A2(n3421), .ZN(n3419) );
  OR2_X1 U3389 ( .A1(n3328), .A2(n3325), .ZN(n3421) );
  OR2_X1 U3390 ( .A1(n2705), .A2(n2326), .ZN(n3325) );
  OR2_X1 U3391 ( .A1(n3045), .A2(n3422), .ZN(n3328) );
  OR2_X1 U3392 ( .A1(n2326), .A2(n2354), .ZN(n3422) );
  INV_X1 U3393 ( .A(b_11_), .ZN(n2326) );
  INV_X1 U3394 ( .A(n3423), .ZN(n3327) );
  OR2_X1 U3395 ( .A1(n3424), .A2(n3425), .ZN(n3423) );
  AND2_X1 U3396 ( .A1(b_9_), .A2(n3426), .ZN(n3425) );
  OR2_X1 U3397 ( .A1(n3427), .A2(n2217), .ZN(n3426) );
  AND2_X1 U3398 ( .A1(a_15_), .A2(n2354), .ZN(n3427) );
  AND2_X1 U3399 ( .A1(b_10_), .A2(n3428), .ZN(n3424) );
  OR2_X1 U3400 ( .A1(n3429), .A2(n3051), .ZN(n3428) );
  AND2_X1 U3401 ( .A1(a_14_), .A2(n2382), .ZN(n3429) );
  XNOR2_X1 U3402 ( .A(n3430), .B(n3431), .ZN(n3330) );
  XNOR2_X1 U3403 ( .A(n3432), .B(n3433), .ZN(n3431) );
  XNOR2_X1 U3404 ( .A(n3434), .B(n3435), .ZN(n3333) );
  XNOR2_X1 U3405 ( .A(n3436), .B(n3437), .ZN(n3434) );
  XOR2_X1 U3406 ( .A(n3438), .B(n3439), .Z(n3336) );
  XOR2_X1 U3407 ( .A(n3440), .B(n3441), .Z(n3439) );
  XOR2_X1 U3408 ( .A(n3442), .B(n3443), .Z(n3340) );
  XOR2_X1 U3409 ( .A(n3444), .B(n2694), .Z(n3443) );
  XOR2_X1 U3410 ( .A(n3445), .B(n3446), .Z(n3344) );
  XOR2_X1 U3411 ( .A(n3447), .B(n3448), .Z(n3446) );
  XOR2_X1 U3412 ( .A(n3449), .B(n3450), .Z(n3348) );
  XOR2_X1 U3413 ( .A(n3451), .B(n3452), .Z(n3450) );
  XOR2_X1 U3414 ( .A(n3453), .B(n3454), .Z(n3352) );
  XOR2_X1 U3415 ( .A(n3455), .B(n3456), .Z(n3454) );
  XOR2_X1 U3416 ( .A(n3457), .B(n3458), .Z(n3356) );
  XOR2_X1 U3417 ( .A(n3459), .B(n3460), .Z(n3458) );
  XOR2_X1 U3418 ( .A(n3461), .B(n3462), .Z(n3360) );
  XOR2_X1 U3419 ( .A(n3463), .B(n3464), .Z(n3462) );
  XOR2_X1 U3420 ( .A(n3465), .B(n3466), .Z(n3364) );
  XOR2_X1 U3421 ( .A(n3467), .B(n3468), .Z(n3466) );
  XOR2_X1 U3422 ( .A(n3469), .B(n3470), .Z(n3368) );
  XOR2_X1 U3423 ( .A(n3471), .B(n3472), .Z(n3470) );
  XOR2_X1 U3424 ( .A(n3473), .B(n3474), .Z(n3372) );
  XOR2_X1 U3425 ( .A(n3475), .B(n3476), .Z(n3474) );
  XOR2_X1 U3426 ( .A(n3477), .B(n3478), .Z(n3376) );
  XOR2_X1 U3427 ( .A(n3479), .B(n3480), .Z(n3478) );
  XNOR2_X1 U3428 ( .A(n3481), .B(n3482), .ZN(n2942) );
  XOR2_X1 U3429 ( .A(n3483), .B(n3484), .Z(n3482) );
  INV_X1 U3430 ( .A(n3485), .ZN(n2762) );
  OR2_X1 U3431 ( .A1(n3486), .A2(n2939), .ZN(n3485) );
  INV_X1 U3432 ( .A(n3487), .ZN(n2939) );
  OR2_X1 U3433 ( .A1(n3488), .A2(n3489), .ZN(n3487) );
  AND2_X1 U3434 ( .A1(n3488), .A2(n3489), .ZN(n3486) );
  OR2_X1 U3435 ( .A1(n3490), .A2(n3491), .ZN(n3489) );
  AND2_X1 U3436 ( .A1(n3484), .A2(n3483), .ZN(n3491) );
  AND2_X1 U3437 ( .A1(n3481), .A2(n3492), .ZN(n3490) );
  OR2_X1 U3438 ( .A1(n3484), .A2(n3483), .ZN(n3492) );
  OR2_X1 U3439 ( .A1(n3493), .A2(n3494), .ZN(n3483) );
  AND2_X1 U3440 ( .A1(n3480), .A2(n3479), .ZN(n3494) );
  AND2_X1 U3441 ( .A1(n3477), .A2(n3495), .ZN(n3493) );
  OR2_X1 U3442 ( .A1(n3480), .A2(n3479), .ZN(n3495) );
  OR2_X1 U3443 ( .A1(n3496), .A2(n3497), .ZN(n3479) );
  AND2_X1 U3444 ( .A1(n3476), .A2(n3475), .ZN(n3497) );
  AND2_X1 U3445 ( .A1(n3473), .A2(n3498), .ZN(n3496) );
  OR2_X1 U3446 ( .A1(n3476), .A2(n3475), .ZN(n3498) );
  OR2_X1 U3447 ( .A1(n3499), .A2(n3500), .ZN(n3475) );
  AND2_X1 U3448 ( .A1(n3469), .A2(n3472), .ZN(n3500) );
  AND2_X1 U3449 ( .A1(n3501), .A2(n3471), .ZN(n3499) );
  OR2_X1 U3450 ( .A1(n3502), .A2(n3503), .ZN(n3471) );
  AND2_X1 U3451 ( .A1(n3468), .A2(n3467), .ZN(n3503) );
  AND2_X1 U3452 ( .A1(n3465), .A2(n3504), .ZN(n3502) );
  OR2_X1 U3453 ( .A1(n3468), .A2(n3467), .ZN(n3504) );
  OR2_X1 U3454 ( .A1(n3505), .A2(n3506), .ZN(n3467) );
  AND2_X1 U3455 ( .A1(n3461), .A2(n3464), .ZN(n3506) );
  AND2_X1 U3456 ( .A1(n3507), .A2(n3463), .ZN(n3505) );
  OR2_X1 U3457 ( .A1(n3508), .A2(n3509), .ZN(n3463) );
  AND2_X1 U3458 ( .A1(n3457), .A2(n3460), .ZN(n3509) );
  AND2_X1 U3459 ( .A1(n3510), .A2(n3459), .ZN(n3508) );
  OR2_X1 U3460 ( .A1(n3511), .A2(n3512), .ZN(n3459) );
  AND2_X1 U3461 ( .A1(n3453), .A2(n3456), .ZN(n3512) );
  AND2_X1 U3462 ( .A1(n3513), .A2(n3455), .ZN(n3511) );
  OR2_X1 U3463 ( .A1(n3514), .A2(n3515), .ZN(n3455) );
  AND2_X1 U3464 ( .A1(n3449), .A2(n3452), .ZN(n3515) );
  AND2_X1 U3465 ( .A1(n3516), .A2(n3451), .ZN(n3514) );
  OR2_X1 U3466 ( .A1(n3517), .A2(n3518), .ZN(n3451) );
  AND2_X1 U3467 ( .A1(n3445), .A2(n3448), .ZN(n3518) );
  AND2_X1 U3468 ( .A1(n3519), .A2(n3447), .ZN(n3517) );
  OR2_X1 U3469 ( .A1(n3520), .A2(n3521), .ZN(n3447) );
  AND2_X1 U3470 ( .A1(n3442), .A2(n2694), .ZN(n3521) );
  AND2_X1 U3471 ( .A1(n3522), .A2(n3444), .ZN(n3520) );
  OR2_X1 U3472 ( .A1(n3523), .A2(n3524), .ZN(n3444) );
  AND2_X1 U3473 ( .A1(n3438), .A2(n3441), .ZN(n3524) );
  AND2_X1 U3474 ( .A1(n3525), .A2(n3440), .ZN(n3523) );
  OR2_X1 U3475 ( .A1(n3526), .A2(n3527), .ZN(n3440) );
  AND2_X1 U3476 ( .A1(n3435), .A2(n3437), .ZN(n3527) );
  AND2_X1 U3477 ( .A1(n3528), .A2(n3436), .ZN(n3526) );
  OR2_X1 U3478 ( .A1(n3529), .A2(n3530), .ZN(n3436) );
  AND2_X1 U3479 ( .A1(n3430), .A2(n3433), .ZN(n3530) );
  AND2_X1 U3480 ( .A1(n3432), .A2(n3531), .ZN(n3529) );
  OR2_X1 U3481 ( .A1(n3430), .A2(n3433), .ZN(n3531) );
  OR2_X1 U3482 ( .A1(n3045), .A2(n3532), .ZN(n3433) );
  OR2_X1 U3483 ( .A1(n2354), .A2(n2382), .ZN(n3532) );
  OR2_X1 U3484 ( .A1(n2705), .A2(n2354), .ZN(n3430) );
  INV_X1 U3485 ( .A(n3533), .ZN(n3432) );
  OR2_X1 U3486 ( .A1(n3534), .A2(n3535), .ZN(n3533) );
  AND2_X1 U3487 ( .A1(b_9_), .A2(n3536), .ZN(n3535) );
  OR2_X1 U3488 ( .A1(n3537), .A2(n3051), .ZN(n3536) );
  AND2_X1 U3489 ( .A1(a_14_), .A2(n2686), .ZN(n3537) );
  AND2_X1 U3490 ( .A1(b_8_), .A2(n3538), .ZN(n3534) );
  OR2_X1 U3491 ( .A1(n3539), .A2(n2217), .ZN(n3538) );
  AND2_X1 U3492 ( .A1(a_15_), .A2(n2382), .ZN(n3539) );
  OR2_X1 U3493 ( .A1(n3435), .A2(n3437), .ZN(n3528) );
  OR2_X1 U3494 ( .A1(n2701), .A2(n2354), .ZN(n3437) );
  XNOR2_X1 U3495 ( .A(n3540), .B(n3541), .ZN(n3435) );
  XNOR2_X1 U3496 ( .A(n3542), .B(n3543), .ZN(n3541) );
  OR2_X1 U3497 ( .A1(n3438), .A2(n3441), .ZN(n3525) );
  OR2_X1 U3498 ( .A1(n2697), .A2(n2354), .ZN(n3441) );
  XNOR2_X1 U3499 ( .A(n3544), .B(n3545), .ZN(n3438) );
  XNOR2_X1 U3500 ( .A(n3546), .B(n3547), .ZN(n3544) );
  OR2_X1 U3501 ( .A1(n3442), .A2(n2694), .ZN(n3522) );
  OR2_X1 U3502 ( .A1(n2693), .A2(n2354), .ZN(n2694) );
  XOR2_X1 U3503 ( .A(n3548), .B(n3549), .Z(n3442) );
  XOR2_X1 U3504 ( .A(n3550), .B(n3551), .Z(n3549) );
  OR2_X1 U3505 ( .A1(n3445), .A2(n3448), .ZN(n3519) );
  OR2_X1 U3506 ( .A1(n2689), .A2(n2354), .ZN(n3448) );
  XOR2_X1 U3507 ( .A(n3552), .B(n3553), .Z(n3445) );
  XOR2_X1 U3508 ( .A(n3554), .B(n3555), .Z(n3553) );
  OR2_X1 U3509 ( .A1(n3449), .A2(n3452), .ZN(n3516) );
  OR2_X1 U3510 ( .A1(n2685), .A2(n2354), .ZN(n3452) );
  XOR2_X1 U3511 ( .A(n3556), .B(n3557), .Z(n3449) );
  XOR2_X1 U3512 ( .A(n3558), .B(n2690), .Z(n3557) );
  OR2_X1 U3513 ( .A1(n3453), .A2(n3456), .ZN(n3513) );
  OR2_X1 U3514 ( .A1(n2681), .A2(n2354), .ZN(n3456) );
  XOR2_X1 U3515 ( .A(n3559), .B(n3560), .Z(n3453) );
  XOR2_X1 U3516 ( .A(n3561), .B(n3562), .Z(n3560) );
  OR2_X1 U3517 ( .A1(n3457), .A2(n3460), .ZN(n3510) );
  OR2_X1 U3518 ( .A1(n2677), .A2(n2354), .ZN(n3460) );
  XOR2_X1 U3519 ( .A(n3563), .B(n3564), .Z(n3457) );
  XOR2_X1 U3520 ( .A(n3565), .B(n3566), .Z(n3564) );
  OR2_X1 U3521 ( .A1(n3461), .A2(n3464), .ZN(n3507) );
  OR2_X1 U3522 ( .A1(n2673), .A2(n2354), .ZN(n3464) );
  XOR2_X1 U3523 ( .A(n3567), .B(n3568), .Z(n3461) );
  XOR2_X1 U3524 ( .A(n3569), .B(n3570), .Z(n3568) );
  OR2_X1 U3525 ( .A1(n2669), .A2(n2354), .ZN(n3468) );
  XOR2_X1 U3526 ( .A(n3571), .B(n3572), .Z(n3465) );
  XOR2_X1 U3527 ( .A(n3573), .B(n3574), .Z(n3572) );
  OR2_X1 U3528 ( .A1(n3469), .A2(n3472), .ZN(n3501) );
  OR2_X1 U3529 ( .A1(n2665), .A2(n2354), .ZN(n3472) );
  XOR2_X1 U3530 ( .A(n3575), .B(n3576), .Z(n3469) );
  XOR2_X1 U3531 ( .A(n3577), .B(n3578), .Z(n3576) );
  OR2_X1 U3532 ( .A1(n2661), .A2(n2354), .ZN(n3476) );
  XOR2_X1 U3533 ( .A(n3579), .B(n3580), .Z(n3473) );
  XOR2_X1 U3534 ( .A(n3581), .B(n3582), .Z(n3580) );
  OR2_X1 U3535 ( .A1(n2657), .A2(n2354), .ZN(n3480) );
  XOR2_X1 U3536 ( .A(n3583), .B(n3584), .Z(n3477) );
  XOR2_X1 U3537 ( .A(n3585), .B(n3586), .Z(n3584) );
  OR2_X1 U3538 ( .A1(n2815), .A2(n2354), .ZN(n3484) );
  INV_X1 U3539 ( .A(b_10_), .ZN(n2354) );
  XOR2_X1 U3540 ( .A(n3587), .B(n3588), .Z(n3481) );
  XOR2_X1 U3541 ( .A(n3589), .B(n3590), .Z(n3588) );
  XOR2_X1 U3542 ( .A(n3591), .B(n3592), .Z(n3488) );
  XOR2_X1 U3543 ( .A(n3593), .B(n3594), .Z(n3592) );
  INV_X1 U3544 ( .A(n3595), .ZN(n2932) );
  OR2_X1 U3545 ( .A1(n2936), .A2(n2937), .ZN(n3595) );
  OR2_X1 U3546 ( .A1(n3596), .A2(n3597), .ZN(n2937) );
  AND2_X1 U3547 ( .A1(n3594), .A2(n3593), .ZN(n3597) );
  AND2_X1 U3548 ( .A1(n3591), .A2(n3598), .ZN(n3596) );
  OR2_X1 U3549 ( .A1(n3594), .A2(n3593), .ZN(n3598) );
  OR2_X1 U3550 ( .A1(n3599), .A2(n3600), .ZN(n3593) );
  AND2_X1 U3551 ( .A1(n3590), .A2(n3589), .ZN(n3600) );
  AND2_X1 U3552 ( .A1(n3587), .A2(n3601), .ZN(n3599) );
  OR2_X1 U3553 ( .A1(n3590), .A2(n3589), .ZN(n3601) );
  OR2_X1 U3554 ( .A1(n3602), .A2(n3603), .ZN(n3589) );
  AND2_X1 U3555 ( .A1(n3586), .A2(n3585), .ZN(n3603) );
  AND2_X1 U3556 ( .A1(n3583), .A2(n3604), .ZN(n3602) );
  OR2_X1 U3557 ( .A1(n3586), .A2(n3585), .ZN(n3604) );
  OR2_X1 U3558 ( .A1(n3605), .A2(n3606), .ZN(n3585) );
  AND2_X1 U3559 ( .A1(n3582), .A2(n3581), .ZN(n3606) );
  AND2_X1 U3560 ( .A1(n3579), .A2(n3607), .ZN(n3605) );
  OR2_X1 U3561 ( .A1(n3582), .A2(n3581), .ZN(n3607) );
  OR2_X1 U3562 ( .A1(n3608), .A2(n3609), .ZN(n3581) );
  AND2_X1 U3563 ( .A1(n3575), .A2(n3578), .ZN(n3609) );
  AND2_X1 U3564 ( .A1(n3610), .A2(n3577), .ZN(n3608) );
  OR2_X1 U3565 ( .A1(n3611), .A2(n3612), .ZN(n3577) );
  AND2_X1 U3566 ( .A1(n3574), .A2(n3573), .ZN(n3612) );
  AND2_X1 U3567 ( .A1(n3571), .A2(n3613), .ZN(n3611) );
  OR2_X1 U3568 ( .A1(n3574), .A2(n3573), .ZN(n3613) );
  OR2_X1 U3569 ( .A1(n3614), .A2(n3615), .ZN(n3573) );
  AND2_X1 U3570 ( .A1(n3567), .A2(n3570), .ZN(n3615) );
  AND2_X1 U3571 ( .A1(n3616), .A2(n3569), .ZN(n3614) );
  OR2_X1 U3572 ( .A1(n3617), .A2(n3618), .ZN(n3569) );
  AND2_X1 U3573 ( .A1(n3563), .A2(n3566), .ZN(n3618) );
  AND2_X1 U3574 ( .A1(n3619), .A2(n3565), .ZN(n3617) );
  OR2_X1 U3575 ( .A1(n3620), .A2(n3621), .ZN(n3565) );
  AND2_X1 U3576 ( .A1(n3559), .A2(n3562), .ZN(n3621) );
  AND2_X1 U3577 ( .A1(n3622), .A2(n3561), .ZN(n3620) );
  OR2_X1 U3578 ( .A1(n3623), .A2(n3624), .ZN(n3561) );
  AND2_X1 U3579 ( .A1(n3556), .A2(n2690), .ZN(n3624) );
  AND2_X1 U3580 ( .A1(n3625), .A2(n3558), .ZN(n3623) );
  OR2_X1 U3581 ( .A1(n3626), .A2(n3627), .ZN(n3558) );
  AND2_X1 U3582 ( .A1(n3552), .A2(n3555), .ZN(n3627) );
  AND2_X1 U3583 ( .A1(n3628), .A2(n3554), .ZN(n3626) );
  OR2_X1 U3584 ( .A1(n3629), .A2(n3630), .ZN(n3554) );
  AND2_X1 U3585 ( .A1(n3548), .A2(n3551), .ZN(n3630) );
  AND2_X1 U3586 ( .A1(n3631), .A2(n3550), .ZN(n3629) );
  OR2_X1 U3587 ( .A1(n3632), .A2(n3633), .ZN(n3550) );
  AND2_X1 U3588 ( .A1(n3545), .A2(n3547), .ZN(n3633) );
  AND2_X1 U3589 ( .A1(n3634), .A2(n3546), .ZN(n3632) );
  OR2_X1 U3590 ( .A1(n3635), .A2(n3636), .ZN(n3546) );
  AND2_X1 U3591 ( .A1(n3540), .A2(n3543), .ZN(n3636) );
  AND2_X1 U3592 ( .A1(n3542), .A2(n3637), .ZN(n3635) );
  OR2_X1 U3593 ( .A1(n3540), .A2(n3543), .ZN(n3637) );
  OR2_X1 U3594 ( .A1(n3045), .A2(n3638), .ZN(n3543) );
  OR2_X1 U3595 ( .A1(n2382), .A2(n2686), .ZN(n3638) );
  OR2_X1 U3596 ( .A1(n2705), .A2(n2382), .ZN(n3540) );
  INV_X1 U3597 ( .A(n3639), .ZN(n3542) );
  OR2_X1 U3598 ( .A1(n3640), .A2(n3641), .ZN(n3639) );
  AND2_X1 U3599 ( .A1(b_8_), .A2(n3642), .ZN(n3641) );
  OR2_X1 U3600 ( .A1(n3643), .A2(n3051), .ZN(n3642) );
  AND2_X1 U3601 ( .A1(a_14_), .A2(n2682), .ZN(n3643) );
  AND2_X1 U3602 ( .A1(b_7_), .A2(n3644), .ZN(n3640) );
  OR2_X1 U3603 ( .A1(n3645), .A2(n2217), .ZN(n3644) );
  AND2_X1 U3604 ( .A1(a_15_), .A2(n2686), .ZN(n3645) );
  OR2_X1 U3605 ( .A1(n3545), .A2(n3547), .ZN(n3634) );
  OR2_X1 U3606 ( .A1(n2701), .A2(n2382), .ZN(n3547) );
  XNOR2_X1 U3607 ( .A(n3646), .B(n3647), .ZN(n3545) );
  XNOR2_X1 U3608 ( .A(n3648), .B(n3649), .ZN(n3647) );
  OR2_X1 U3609 ( .A1(n3548), .A2(n3551), .ZN(n3631) );
  OR2_X1 U3610 ( .A1(n2697), .A2(n2382), .ZN(n3551) );
  XNOR2_X1 U3611 ( .A(n3650), .B(n3651), .ZN(n3548) );
  XNOR2_X1 U3612 ( .A(n3652), .B(n3653), .ZN(n3650) );
  OR2_X1 U3613 ( .A1(n3552), .A2(n3555), .ZN(n3628) );
  OR2_X1 U3614 ( .A1(n2693), .A2(n2382), .ZN(n3555) );
  XOR2_X1 U3615 ( .A(n3654), .B(n3655), .Z(n3552) );
  XOR2_X1 U3616 ( .A(n3656), .B(n3657), .Z(n3655) );
  OR2_X1 U3617 ( .A1(n3556), .A2(n2690), .ZN(n3625) );
  OR2_X1 U3618 ( .A1(n2689), .A2(n2382), .ZN(n2690) );
  XOR2_X1 U3619 ( .A(n3658), .B(n3659), .Z(n3556) );
  XOR2_X1 U3620 ( .A(n3660), .B(n3661), .Z(n3659) );
  OR2_X1 U3621 ( .A1(n3559), .A2(n3562), .ZN(n3622) );
  OR2_X1 U3622 ( .A1(n2685), .A2(n2382), .ZN(n3562) );
  XOR2_X1 U3623 ( .A(n3662), .B(n3663), .Z(n3559) );
  XOR2_X1 U3624 ( .A(n3664), .B(n3665), .Z(n3663) );
  OR2_X1 U3625 ( .A1(n3563), .A2(n3566), .ZN(n3619) );
  OR2_X1 U3626 ( .A1(n2681), .A2(n2382), .ZN(n3566) );
  XOR2_X1 U3627 ( .A(n3666), .B(n3667), .Z(n3563) );
  XOR2_X1 U3628 ( .A(n3668), .B(n2406), .Z(n3667) );
  OR2_X1 U3629 ( .A1(n3567), .A2(n3570), .ZN(n3616) );
  OR2_X1 U3630 ( .A1(n2677), .A2(n2382), .ZN(n3570) );
  XOR2_X1 U3631 ( .A(n3669), .B(n3670), .Z(n3567) );
  XOR2_X1 U3632 ( .A(n3671), .B(n3672), .Z(n3670) );
  OR2_X1 U3633 ( .A1(n2673), .A2(n2382), .ZN(n3574) );
  XOR2_X1 U3634 ( .A(n3673), .B(n3674), .Z(n3571) );
  XOR2_X1 U3635 ( .A(n3675), .B(n3676), .Z(n3674) );
  OR2_X1 U3636 ( .A1(n3575), .A2(n3578), .ZN(n3610) );
  OR2_X1 U3637 ( .A1(n2669), .A2(n2382), .ZN(n3578) );
  XOR2_X1 U3638 ( .A(n3677), .B(n3678), .Z(n3575) );
  XOR2_X1 U3639 ( .A(n3679), .B(n3680), .Z(n3678) );
  OR2_X1 U3640 ( .A1(n2665), .A2(n2382), .ZN(n3582) );
  XOR2_X1 U3641 ( .A(n3681), .B(n3682), .Z(n3579) );
  XOR2_X1 U3642 ( .A(n3683), .B(n3684), .Z(n3682) );
  OR2_X1 U3643 ( .A1(n2661), .A2(n2382), .ZN(n3586) );
  XOR2_X1 U3644 ( .A(n3685), .B(n3686), .Z(n3583) );
  XOR2_X1 U3645 ( .A(n3687), .B(n3688), .Z(n3686) );
  OR2_X1 U3646 ( .A1(n2657), .A2(n2382), .ZN(n3590) );
  XOR2_X1 U3647 ( .A(n3689), .B(n3690), .Z(n3587) );
  XOR2_X1 U3648 ( .A(n3691), .B(n3692), .Z(n3690) );
  OR2_X1 U3649 ( .A1(n2815), .A2(n2382), .ZN(n3594) );
  INV_X1 U3650 ( .A(b_9_), .ZN(n2382) );
  XOR2_X1 U3651 ( .A(n3693), .B(n3694), .Z(n3591) );
  XOR2_X1 U3652 ( .A(n3695), .B(n3696), .Z(n3694) );
  XOR2_X1 U3653 ( .A(n2926), .B(n3697), .Z(n2936) );
  XOR2_X1 U3654 ( .A(n2925), .B(n2924), .Z(n3697) );
  OR2_X1 U3655 ( .A1(n2815), .A2(n2686), .ZN(n2924) );
  OR2_X1 U3656 ( .A1(n3698), .A2(n3699), .ZN(n2925) );
  AND2_X1 U3657 ( .A1(n3696), .A2(n3695), .ZN(n3699) );
  AND2_X1 U3658 ( .A1(n3693), .A2(n3700), .ZN(n3698) );
  OR2_X1 U3659 ( .A1(n3695), .A2(n3696), .ZN(n3700) );
  OR2_X1 U3660 ( .A1(n2657), .A2(n2686), .ZN(n3696) );
  OR2_X1 U3661 ( .A1(n3701), .A2(n3702), .ZN(n3695) );
  AND2_X1 U3662 ( .A1(n3692), .A2(n3691), .ZN(n3702) );
  AND2_X1 U3663 ( .A1(n3689), .A2(n3703), .ZN(n3701) );
  OR2_X1 U3664 ( .A1(n3691), .A2(n3692), .ZN(n3703) );
  OR2_X1 U3665 ( .A1(n2661), .A2(n2686), .ZN(n3692) );
  OR2_X1 U3666 ( .A1(n3704), .A2(n3705), .ZN(n3691) );
  AND2_X1 U3667 ( .A1(n3688), .A2(n3687), .ZN(n3705) );
  AND2_X1 U3668 ( .A1(n3685), .A2(n3706), .ZN(n3704) );
  OR2_X1 U3669 ( .A1(n3687), .A2(n3688), .ZN(n3706) );
  OR2_X1 U3670 ( .A1(n2665), .A2(n2686), .ZN(n3688) );
  OR2_X1 U3671 ( .A1(n3707), .A2(n3708), .ZN(n3687) );
  AND2_X1 U3672 ( .A1(n3684), .A2(n3683), .ZN(n3708) );
  AND2_X1 U3673 ( .A1(n3681), .A2(n3709), .ZN(n3707) );
  OR2_X1 U3674 ( .A1(n3683), .A2(n3684), .ZN(n3709) );
  OR2_X1 U3675 ( .A1(n2669), .A2(n2686), .ZN(n3684) );
  OR2_X1 U3676 ( .A1(n3710), .A2(n3711), .ZN(n3683) );
  AND2_X1 U3677 ( .A1(n3677), .A2(n3680), .ZN(n3711) );
  AND2_X1 U3678 ( .A1(n3712), .A2(n3679), .ZN(n3710) );
  OR2_X1 U3679 ( .A1(n3713), .A2(n3714), .ZN(n3679) );
  AND2_X1 U3680 ( .A1(n3676), .A2(n3675), .ZN(n3714) );
  AND2_X1 U3681 ( .A1(n3673), .A2(n3715), .ZN(n3713) );
  OR2_X1 U3682 ( .A1(n3675), .A2(n3676), .ZN(n3715) );
  OR2_X1 U3683 ( .A1(n2677), .A2(n2686), .ZN(n3676) );
  OR2_X1 U3684 ( .A1(n3716), .A2(n3717), .ZN(n3675) );
  AND2_X1 U3685 ( .A1(n3669), .A2(n3672), .ZN(n3717) );
  AND2_X1 U3686 ( .A1(n3718), .A2(n3671), .ZN(n3716) );
  OR2_X1 U3687 ( .A1(n3719), .A2(n3720), .ZN(n3671) );
  AND2_X1 U3688 ( .A1(n3666), .A2(n2406), .ZN(n3720) );
  AND2_X1 U3689 ( .A1(n3721), .A2(n3668), .ZN(n3719) );
  OR2_X1 U3690 ( .A1(n3722), .A2(n3723), .ZN(n3668) );
  AND2_X1 U3691 ( .A1(n3662), .A2(n3665), .ZN(n3723) );
  AND2_X1 U3692 ( .A1(n3724), .A2(n3664), .ZN(n3722) );
  OR2_X1 U3693 ( .A1(n3725), .A2(n3726), .ZN(n3664) );
  AND2_X1 U3694 ( .A1(n3658), .A2(n3661), .ZN(n3726) );
  AND2_X1 U3695 ( .A1(n3727), .A2(n3660), .ZN(n3725) );
  OR2_X1 U3696 ( .A1(n3728), .A2(n3729), .ZN(n3660) );
  AND2_X1 U3697 ( .A1(n3654), .A2(n3657), .ZN(n3729) );
  AND2_X1 U3698 ( .A1(n3730), .A2(n3656), .ZN(n3728) );
  OR2_X1 U3699 ( .A1(n3731), .A2(n3732), .ZN(n3656) );
  AND2_X1 U3700 ( .A1(n3651), .A2(n3653), .ZN(n3732) );
  AND2_X1 U3701 ( .A1(n3733), .A2(n3652), .ZN(n3731) );
  OR2_X1 U3702 ( .A1(n3734), .A2(n3735), .ZN(n3652) );
  AND2_X1 U3703 ( .A1(n3646), .A2(n3649), .ZN(n3735) );
  AND2_X1 U3704 ( .A1(n3648), .A2(n3736), .ZN(n3734) );
  OR2_X1 U3705 ( .A1(n3649), .A2(n3646), .ZN(n3736) );
  OR2_X1 U3706 ( .A1(n2705), .A2(n2686), .ZN(n3646) );
  OR2_X1 U3707 ( .A1(n3045), .A2(n3737), .ZN(n3649) );
  OR2_X1 U3708 ( .A1(n2686), .A2(n2682), .ZN(n3737) );
  INV_X1 U3709 ( .A(n3738), .ZN(n3648) );
  OR2_X1 U3710 ( .A1(n3739), .A2(n3740), .ZN(n3738) );
  AND2_X1 U3711 ( .A1(b_7_), .A2(n3741), .ZN(n3740) );
  OR2_X1 U3712 ( .A1(n3742), .A2(n3051), .ZN(n3741) );
  AND2_X1 U3713 ( .A1(a_14_), .A2(n2678), .ZN(n3742) );
  AND2_X1 U3714 ( .A1(b_6_), .A2(n3743), .ZN(n3739) );
  OR2_X1 U3715 ( .A1(n3744), .A2(n2217), .ZN(n3743) );
  AND2_X1 U3716 ( .A1(a_15_), .A2(n2682), .ZN(n3744) );
  OR2_X1 U3717 ( .A1(n3653), .A2(n3651), .ZN(n3733) );
  XNOR2_X1 U3718 ( .A(n3745), .B(n3746), .ZN(n3651) );
  XNOR2_X1 U3719 ( .A(n3747), .B(n3748), .ZN(n3746) );
  OR2_X1 U3720 ( .A1(n2701), .A2(n2686), .ZN(n3653) );
  OR2_X1 U3721 ( .A1(n3657), .A2(n3654), .ZN(n3730) );
  XNOR2_X1 U3722 ( .A(n3749), .B(n3750), .ZN(n3654) );
  XNOR2_X1 U3723 ( .A(n3751), .B(n3752), .ZN(n3749) );
  OR2_X1 U3724 ( .A1(n2697), .A2(n2686), .ZN(n3657) );
  OR2_X1 U3725 ( .A1(n3661), .A2(n3658), .ZN(n3727) );
  XOR2_X1 U3726 ( .A(n3753), .B(n3754), .Z(n3658) );
  XOR2_X1 U3727 ( .A(n3755), .B(n3756), .Z(n3754) );
  OR2_X1 U3728 ( .A1(n2693), .A2(n2686), .ZN(n3661) );
  OR2_X1 U3729 ( .A1(n3665), .A2(n3662), .ZN(n3724) );
  XOR2_X1 U3730 ( .A(n3757), .B(n3758), .Z(n3662) );
  XOR2_X1 U3731 ( .A(n3759), .B(n3760), .Z(n3758) );
  OR2_X1 U3732 ( .A1(n2689), .A2(n2686), .ZN(n3665) );
  OR2_X1 U3733 ( .A1(n2406), .A2(n3666), .ZN(n3721) );
  XOR2_X1 U3734 ( .A(n3761), .B(n3762), .Z(n3666) );
  XOR2_X1 U3735 ( .A(n3763), .B(n3764), .Z(n3762) );
  OR2_X1 U3736 ( .A1(n2685), .A2(n2686), .ZN(n2406) );
  OR2_X1 U3737 ( .A1(n3672), .A2(n3669), .ZN(n3718) );
  XOR2_X1 U3738 ( .A(n3765), .B(n3766), .Z(n3669) );
  XOR2_X1 U3739 ( .A(n3767), .B(n3768), .Z(n3766) );
  OR2_X1 U3740 ( .A1(n2681), .A2(n2686), .ZN(n3672) );
  XOR2_X1 U3741 ( .A(n3769), .B(n3770), .Z(n3673) );
  XOR2_X1 U3742 ( .A(n3771), .B(n2435), .Z(n3770) );
  OR2_X1 U3743 ( .A1(n3680), .A2(n3677), .ZN(n3712) );
  XOR2_X1 U3744 ( .A(n3772), .B(n3773), .Z(n3677) );
  XOR2_X1 U3745 ( .A(n3774), .B(n3775), .Z(n3773) );
  OR2_X1 U3746 ( .A1(n2673), .A2(n2686), .ZN(n3680) );
  INV_X1 U3747 ( .A(b_8_), .ZN(n2686) );
  XOR2_X1 U3748 ( .A(n3776), .B(n3777), .Z(n3681) );
  XOR2_X1 U3749 ( .A(n3778), .B(n3779), .Z(n3777) );
  XOR2_X1 U3750 ( .A(n3780), .B(n3781), .Z(n3685) );
  XOR2_X1 U3751 ( .A(n3782), .B(n3783), .Z(n3781) );
  XOR2_X1 U3752 ( .A(n3784), .B(n3785), .Z(n3689) );
  XOR2_X1 U3753 ( .A(n3786), .B(n3787), .Z(n3785) );
  XOR2_X1 U3754 ( .A(n3788), .B(n3789), .Z(n3693) );
  XOR2_X1 U3755 ( .A(n3790), .B(n3791), .Z(n3789) );
  XOR2_X1 U3756 ( .A(n3792), .B(n3793), .Z(n2926) );
  XOR2_X1 U3757 ( .A(n3794), .B(n3795), .Z(n3793) );
  INV_X1 U3758 ( .A(n3796), .ZN(n2909) );
  OR2_X1 U3759 ( .A1(n2913), .A2(n2914), .ZN(n3796) );
  OR2_X1 U3760 ( .A1(n3797), .A2(n3798), .ZN(n2914) );
  AND2_X1 U3761 ( .A1(n2931), .A2(n2930), .ZN(n3798) );
  AND2_X1 U3762 ( .A1(n2928), .A2(n3799), .ZN(n3797) );
  OR2_X1 U3763 ( .A1(n2930), .A2(n2931), .ZN(n3799) );
  OR2_X1 U3764 ( .A1(n2815), .A2(n2682), .ZN(n2931) );
  OR2_X1 U3765 ( .A1(n3800), .A2(n3801), .ZN(n2930) );
  AND2_X1 U3766 ( .A1(n3795), .A2(n3794), .ZN(n3801) );
  AND2_X1 U3767 ( .A1(n3792), .A2(n3802), .ZN(n3800) );
  OR2_X1 U3768 ( .A1(n3794), .A2(n3795), .ZN(n3802) );
  OR2_X1 U3769 ( .A1(n2657), .A2(n2682), .ZN(n3795) );
  OR2_X1 U3770 ( .A1(n3803), .A2(n3804), .ZN(n3794) );
  AND2_X1 U3771 ( .A1(n3791), .A2(n3790), .ZN(n3804) );
  AND2_X1 U3772 ( .A1(n3788), .A2(n3805), .ZN(n3803) );
  OR2_X1 U3773 ( .A1(n3790), .A2(n3791), .ZN(n3805) );
  OR2_X1 U3774 ( .A1(n2661), .A2(n2682), .ZN(n3791) );
  OR2_X1 U3775 ( .A1(n3806), .A2(n3807), .ZN(n3790) );
  AND2_X1 U3776 ( .A1(n3787), .A2(n3786), .ZN(n3807) );
  AND2_X1 U3777 ( .A1(n3784), .A2(n3808), .ZN(n3806) );
  OR2_X1 U3778 ( .A1(n3786), .A2(n3787), .ZN(n3808) );
  OR2_X1 U3779 ( .A1(n2665), .A2(n2682), .ZN(n3787) );
  OR2_X1 U3780 ( .A1(n3809), .A2(n3810), .ZN(n3786) );
  AND2_X1 U3781 ( .A1(n3783), .A2(n3782), .ZN(n3810) );
  AND2_X1 U3782 ( .A1(n3780), .A2(n3811), .ZN(n3809) );
  OR2_X1 U3783 ( .A1(n3782), .A2(n3783), .ZN(n3811) );
  OR2_X1 U3784 ( .A1(n2669), .A2(n2682), .ZN(n3783) );
  OR2_X1 U3785 ( .A1(n3812), .A2(n3813), .ZN(n3782) );
  AND2_X1 U3786 ( .A1(n3779), .A2(n3778), .ZN(n3813) );
  AND2_X1 U3787 ( .A1(n3776), .A2(n3814), .ZN(n3812) );
  OR2_X1 U3788 ( .A1(n3778), .A2(n3779), .ZN(n3814) );
  OR2_X1 U3789 ( .A1(n2673), .A2(n2682), .ZN(n3779) );
  OR2_X1 U3790 ( .A1(n3815), .A2(n3816), .ZN(n3778) );
  AND2_X1 U3791 ( .A1(n3772), .A2(n3775), .ZN(n3816) );
  AND2_X1 U3792 ( .A1(n3817), .A2(n3774), .ZN(n3815) );
  OR2_X1 U3793 ( .A1(n3818), .A2(n3819), .ZN(n3774) );
  AND2_X1 U3794 ( .A1(n2435), .A2(n3771), .ZN(n3819) );
  AND2_X1 U3795 ( .A1(n3769), .A2(n3820), .ZN(n3818) );
  OR2_X1 U3796 ( .A1(n3771), .A2(n2435), .ZN(n3820) );
  OR2_X1 U3797 ( .A1(n2681), .A2(n2682), .ZN(n2435) );
  OR2_X1 U3798 ( .A1(n3821), .A2(n3822), .ZN(n3771) );
  AND2_X1 U3799 ( .A1(n3765), .A2(n3768), .ZN(n3822) );
  AND2_X1 U3800 ( .A1(n3823), .A2(n3767), .ZN(n3821) );
  OR2_X1 U3801 ( .A1(n3824), .A2(n3825), .ZN(n3767) );
  AND2_X1 U3802 ( .A1(n3761), .A2(n3764), .ZN(n3825) );
  AND2_X1 U3803 ( .A1(n3826), .A2(n3763), .ZN(n3824) );
  OR2_X1 U3804 ( .A1(n3827), .A2(n3828), .ZN(n3763) );
  AND2_X1 U3805 ( .A1(n3757), .A2(n3760), .ZN(n3828) );
  AND2_X1 U3806 ( .A1(n3829), .A2(n3759), .ZN(n3827) );
  OR2_X1 U3807 ( .A1(n3830), .A2(n3831), .ZN(n3759) );
  AND2_X1 U3808 ( .A1(n3753), .A2(n3756), .ZN(n3831) );
  AND2_X1 U3809 ( .A1(n3832), .A2(n3755), .ZN(n3830) );
  OR2_X1 U3810 ( .A1(n3833), .A2(n3834), .ZN(n3755) );
  AND2_X1 U3811 ( .A1(n3750), .A2(n3752), .ZN(n3834) );
  AND2_X1 U3812 ( .A1(n3835), .A2(n3751), .ZN(n3833) );
  OR2_X1 U3813 ( .A1(n3836), .A2(n3837), .ZN(n3751) );
  AND2_X1 U3814 ( .A1(n3745), .A2(n3748), .ZN(n3837) );
  AND2_X1 U3815 ( .A1(n3747), .A2(n3838), .ZN(n3836) );
  OR2_X1 U3816 ( .A1(n3748), .A2(n3745), .ZN(n3838) );
  OR2_X1 U3817 ( .A1(n2705), .A2(n2682), .ZN(n3745) );
  OR2_X1 U3818 ( .A1(n3045), .A2(n3839), .ZN(n3748) );
  OR2_X1 U3819 ( .A1(n2682), .A2(n2678), .ZN(n3839) );
  INV_X1 U3820 ( .A(n3840), .ZN(n3747) );
  OR2_X1 U3821 ( .A1(n3841), .A2(n3842), .ZN(n3840) );
  AND2_X1 U3822 ( .A1(b_6_), .A2(n3843), .ZN(n3842) );
  OR2_X1 U3823 ( .A1(n3844), .A2(n3051), .ZN(n3843) );
  AND2_X1 U3824 ( .A1(a_14_), .A2(n2674), .ZN(n3844) );
  AND2_X1 U3825 ( .A1(b_5_), .A2(n3845), .ZN(n3841) );
  OR2_X1 U3826 ( .A1(n3846), .A2(n2217), .ZN(n3845) );
  AND2_X1 U3827 ( .A1(a_15_), .A2(n2678), .ZN(n3846) );
  OR2_X1 U3828 ( .A1(n3752), .A2(n3750), .ZN(n3835) );
  XNOR2_X1 U3829 ( .A(n3847), .B(n3848), .ZN(n3750) );
  XNOR2_X1 U3830 ( .A(n3849), .B(n3850), .ZN(n3848) );
  OR2_X1 U3831 ( .A1(n2701), .A2(n2682), .ZN(n3752) );
  OR2_X1 U3832 ( .A1(n3756), .A2(n3753), .ZN(n3832) );
  XNOR2_X1 U3833 ( .A(n3851), .B(n3852), .ZN(n3753) );
  XNOR2_X1 U3834 ( .A(n3853), .B(n3854), .ZN(n3851) );
  OR2_X1 U3835 ( .A1(n2697), .A2(n2682), .ZN(n3756) );
  OR2_X1 U3836 ( .A1(n3760), .A2(n3757), .ZN(n3829) );
  XOR2_X1 U3837 ( .A(n3855), .B(n3856), .Z(n3757) );
  XOR2_X1 U3838 ( .A(n3857), .B(n3858), .Z(n3856) );
  OR2_X1 U3839 ( .A1(n2693), .A2(n2682), .ZN(n3760) );
  OR2_X1 U3840 ( .A1(n3764), .A2(n3761), .ZN(n3826) );
  XOR2_X1 U3841 ( .A(n3859), .B(n3860), .Z(n3761) );
  XOR2_X1 U3842 ( .A(n3861), .B(n3862), .Z(n3860) );
  OR2_X1 U3843 ( .A1(n2689), .A2(n2682), .ZN(n3764) );
  OR2_X1 U3844 ( .A1(n3768), .A2(n3765), .ZN(n3823) );
  XOR2_X1 U3845 ( .A(n3863), .B(n3864), .Z(n3765) );
  XOR2_X1 U3846 ( .A(n3865), .B(n3866), .Z(n3864) );
  OR2_X1 U3847 ( .A1(n2685), .A2(n2682), .ZN(n3768) );
  XOR2_X1 U3848 ( .A(n3867), .B(n3868), .Z(n3769) );
  XOR2_X1 U3849 ( .A(n3869), .B(n3870), .Z(n3868) );
  OR2_X1 U3850 ( .A1(n3775), .A2(n3772), .ZN(n3817) );
  XOR2_X1 U3851 ( .A(n3871), .B(n3872), .Z(n3772) );
  XOR2_X1 U3852 ( .A(n3873), .B(n3874), .Z(n3872) );
  OR2_X1 U3853 ( .A1(n2677), .A2(n2682), .ZN(n3775) );
  INV_X1 U3854 ( .A(b_7_), .ZN(n2682) );
  XOR2_X1 U3855 ( .A(n3875), .B(n3876), .Z(n3776) );
  XOR2_X1 U3856 ( .A(n3877), .B(n2464), .Z(n3876) );
  XOR2_X1 U3857 ( .A(n3878), .B(n3879), .Z(n3780) );
  XOR2_X1 U3858 ( .A(n3880), .B(n3881), .Z(n3879) );
  XOR2_X1 U3859 ( .A(n3882), .B(n3883), .Z(n3784) );
  XOR2_X1 U3860 ( .A(n3884), .B(n3885), .Z(n3883) );
  XOR2_X1 U3861 ( .A(n3886), .B(n3887), .Z(n3788) );
  XOR2_X1 U3862 ( .A(n3888), .B(n3889), .Z(n3887) );
  XOR2_X1 U3863 ( .A(n3890), .B(n3891), .Z(n3792) );
  XOR2_X1 U3864 ( .A(n3892), .B(n3893), .Z(n3891) );
  XOR2_X1 U3865 ( .A(n3894), .B(n3895), .Z(n2928) );
  XOR2_X1 U3866 ( .A(n3896), .B(n3897), .Z(n3895) );
  XOR2_X1 U3867 ( .A(n2903), .B(n3898), .Z(n2913) );
  XOR2_X1 U3868 ( .A(n2902), .B(n2901), .Z(n3898) );
  OR2_X1 U3869 ( .A1(n2815), .A2(n2678), .ZN(n2901) );
  OR2_X1 U3870 ( .A1(n3899), .A2(n3900), .ZN(n2902) );
  AND2_X1 U3871 ( .A1(n3897), .A2(n3896), .ZN(n3900) );
  AND2_X1 U3872 ( .A1(n3894), .A2(n3901), .ZN(n3899) );
  OR2_X1 U3873 ( .A1(n3896), .A2(n3897), .ZN(n3901) );
  OR2_X1 U3874 ( .A1(n2657), .A2(n2678), .ZN(n3897) );
  OR2_X1 U3875 ( .A1(n3902), .A2(n3903), .ZN(n3896) );
  AND2_X1 U3876 ( .A1(n3893), .A2(n3892), .ZN(n3903) );
  AND2_X1 U3877 ( .A1(n3890), .A2(n3904), .ZN(n3902) );
  OR2_X1 U3878 ( .A1(n3892), .A2(n3893), .ZN(n3904) );
  OR2_X1 U3879 ( .A1(n2661), .A2(n2678), .ZN(n3893) );
  OR2_X1 U3880 ( .A1(n3905), .A2(n3906), .ZN(n3892) );
  AND2_X1 U3881 ( .A1(n3889), .A2(n3888), .ZN(n3906) );
  AND2_X1 U3882 ( .A1(n3886), .A2(n3907), .ZN(n3905) );
  OR2_X1 U3883 ( .A1(n3888), .A2(n3889), .ZN(n3907) );
  OR2_X1 U3884 ( .A1(n2665), .A2(n2678), .ZN(n3889) );
  OR2_X1 U3885 ( .A1(n3908), .A2(n3909), .ZN(n3888) );
  AND2_X1 U3886 ( .A1(n3885), .A2(n3884), .ZN(n3909) );
  AND2_X1 U3887 ( .A1(n3882), .A2(n3910), .ZN(n3908) );
  OR2_X1 U3888 ( .A1(n3884), .A2(n3885), .ZN(n3910) );
  OR2_X1 U3889 ( .A1(n2669), .A2(n2678), .ZN(n3885) );
  OR2_X1 U3890 ( .A1(n3911), .A2(n3912), .ZN(n3884) );
  AND2_X1 U3891 ( .A1(n3881), .A2(n3880), .ZN(n3912) );
  AND2_X1 U3892 ( .A1(n3878), .A2(n3913), .ZN(n3911) );
  OR2_X1 U3893 ( .A1(n3880), .A2(n3881), .ZN(n3913) );
  OR2_X1 U3894 ( .A1(n2673), .A2(n2678), .ZN(n3881) );
  OR2_X1 U3895 ( .A1(n3914), .A2(n3915), .ZN(n3880) );
  AND2_X1 U3896 ( .A1(n2464), .A2(n3877), .ZN(n3915) );
  AND2_X1 U3897 ( .A1(n3875), .A2(n3916), .ZN(n3914) );
  OR2_X1 U3898 ( .A1(n3877), .A2(n2464), .ZN(n3916) );
  OR2_X1 U3899 ( .A1(n2677), .A2(n2678), .ZN(n2464) );
  OR2_X1 U3900 ( .A1(n3917), .A2(n3918), .ZN(n3877) );
  AND2_X1 U3901 ( .A1(n3871), .A2(n3874), .ZN(n3918) );
  AND2_X1 U3902 ( .A1(n3919), .A2(n3873), .ZN(n3917) );
  OR2_X1 U3903 ( .A1(n3920), .A2(n3921), .ZN(n3873) );
  AND2_X1 U3904 ( .A1(n3870), .A2(n3869), .ZN(n3921) );
  AND2_X1 U3905 ( .A1(n3867), .A2(n3922), .ZN(n3920) );
  OR2_X1 U3906 ( .A1(n3869), .A2(n3870), .ZN(n3922) );
  OR2_X1 U3907 ( .A1(n2685), .A2(n2678), .ZN(n3870) );
  OR2_X1 U3908 ( .A1(n3923), .A2(n3924), .ZN(n3869) );
  AND2_X1 U3909 ( .A1(n3863), .A2(n3866), .ZN(n3924) );
  AND2_X1 U3910 ( .A1(n3925), .A2(n3865), .ZN(n3923) );
  OR2_X1 U3911 ( .A1(n3926), .A2(n3927), .ZN(n3865) );
  AND2_X1 U3912 ( .A1(n3859), .A2(n3862), .ZN(n3927) );
  AND2_X1 U3913 ( .A1(n3928), .A2(n3861), .ZN(n3926) );
  OR2_X1 U3914 ( .A1(n3929), .A2(n3930), .ZN(n3861) );
  AND2_X1 U3915 ( .A1(n3855), .A2(n3858), .ZN(n3930) );
  AND2_X1 U3916 ( .A1(n3931), .A2(n3857), .ZN(n3929) );
  OR2_X1 U3917 ( .A1(n3932), .A2(n3933), .ZN(n3857) );
  AND2_X1 U3918 ( .A1(n3852), .A2(n3854), .ZN(n3933) );
  AND2_X1 U3919 ( .A1(n3934), .A2(n3853), .ZN(n3932) );
  OR2_X1 U3920 ( .A1(n3935), .A2(n3936), .ZN(n3853) );
  AND2_X1 U3921 ( .A1(n3847), .A2(n3850), .ZN(n3936) );
  AND2_X1 U3922 ( .A1(n3849), .A2(n3937), .ZN(n3935) );
  OR2_X1 U3923 ( .A1(n3850), .A2(n3847), .ZN(n3937) );
  OR2_X1 U3924 ( .A1(n2705), .A2(n2678), .ZN(n3847) );
  OR2_X1 U3925 ( .A1(n3045), .A2(n3938), .ZN(n3850) );
  OR2_X1 U3926 ( .A1(n2678), .A2(n2674), .ZN(n3938) );
  INV_X1 U3927 ( .A(n3939), .ZN(n3849) );
  OR2_X1 U3928 ( .A1(n3940), .A2(n3941), .ZN(n3939) );
  AND2_X1 U3929 ( .A1(b_5_), .A2(n3942), .ZN(n3941) );
  OR2_X1 U3930 ( .A1(n3943), .A2(n3051), .ZN(n3942) );
  AND2_X1 U3931 ( .A1(a_14_), .A2(n2670), .ZN(n3943) );
  AND2_X1 U3932 ( .A1(b_4_), .A2(n3944), .ZN(n3940) );
  OR2_X1 U3933 ( .A1(n3945), .A2(n2217), .ZN(n3944) );
  AND2_X1 U3934 ( .A1(a_15_), .A2(n2674), .ZN(n3945) );
  OR2_X1 U3935 ( .A1(n3854), .A2(n3852), .ZN(n3934) );
  XNOR2_X1 U3936 ( .A(n3946), .B(n3947), .ZN(n3852) );
  XNOR2_X1 U3937 ( .A(n3948), .B(n3949), .ZN(n3947) );
  OR2_X1 U3938 ( .A1(n2701), .A2(n2678), .ZN(n3854) );
  OR2_X1 U3939 ( .A1(n3858), .A2(n3855), .ZN(n3931) );
  XNOR2_X1 U3940 ( .A(n3950), .B(n3951), .ZN(n3855) );
  XNOR2_X1 U3941 ( .A(n3952), .B(n3953), .ZN(n3950) );
  OR2_X1 U3942 ( .A1(n2697), .A2(n2678), .ZN(n3858) );
  OR2_X1 U3943 ( .A1(n3862), .A2(n3859), .ZN(n3928) );
  XOR2_X1 U3944 ( .A(n3954), .B(n3955), .Z(n3859) );
  XOR2_X1 U3945 ( .A(n3956), .B(n3957), .Z(n3955) );
  OR2_X1 U3946 ( .A1(n2693), .A2(n2678), .ZN(n3862) );
  OR2_X1 U3947 ( .A1(n3866), .A2(n3863), .ZN(n3925) );
  XOR2_X1 U3948 ( .A(n3958), .B(n3959), .Z(n3863) );
  XOR2_X1 U3949 ( .A(n3960), .B(n3961), .Z(n3959) );
  OR2_X1 U3950 ( .A1(n2689), .A2(n2678), .ZN(n3866) );
  XOR2_X1 U3951 ( .A(n3962), .B(n3963), .Z(n3867) );
  XOR2_X1 U3952 ( .A(n3964), .B(n3965), .Z(n3963) );
  OR2_X1 U3953 ( .A1(n3874), .A2(n3871), .ZN(n3919) );
  XOR2_X1 U3954 ( .A(n3966), .B(n3967), .Z(n3871) );
  XOR2_X1 U3955 ( .A(n3968), .B(n3969), .Z(n3967) );
  OR2_X1 U3956 ( .A1(n2681), .A2(n2678), .ZN(n3874) );
  INV_X1 U3957 ( .A(b_6_), .ZN(n2678) );
  XOR2_X1 U3958 ( .A(n3970), .B(n3971), .Z(n3875) );
  XOR2_X1 U3959 ( .A(n3972), .B(n3973), .Z(n3971) );
  XOR2_X1 U3960 ( .A(n3974), .B(n3975), .Z(n3878) );
  XOR2_X1 U3961 ( .A(n3976), .B(n3977), .Z(n3975) );
  XOR2_X1 U3962 ( .A(n3978), .B(n3979), .Z(n3882) );
  XOR2_X1 U3963 ( .A(n3980), .B(n2493), .Z(n3979) );
  XOR2_X1 U3964 ( .A(n3981), .B(n3982), .Z(n3886) );
  XOR2_X1 U3965 ( .A(n3983), .B(n3984), .Z(n3982) );
  XOR2_X1 U3966 ( .A(n3985), .B(n3986), .Z(n3890) );
  XOR2_X1 U3967 ( .A(n3987), .B(n3988), .Z(n3986) );
  XOR2_X1 U3968 ( .A(n3989), .B(n3990), .Z(n3894) );
  XOR2_X1 U3969 ( .A(n3991), .B(n3992), .Z(n3990) );
  XOR2_X1 U3970 ( .A(n3993), .B(n3994), .Z(n2903) );
  XOR2_X1 U3971 ( .A(n3995), .B(n3996), .Z(n3994) );
  INV_X1 U3972 ( .A(n3997), .ZN(n2886) );
  OR2_X1 U3973 ( .A1(n2890), .A2(n2891), .ZN(n3997) );
  OR2_X1 U3974 ( .A1(n3998), .A2(n3999), .ZN(n2891) );
  AND2_X1 U3975 ( .A1(n2908), .A2(n2907), .ZN(n3999) );
  AND2_X1 U3976 ( .A1(n2905), .A2(n4000), .ZN(n3998) );
  OR2_X1 U3977 ( .A1(n2907), .A2(n2908), .ZN(n4000) );
  OR2_X1 U3978 ( .A1(n2815), .A2(n2674), .ZN(n2908) );
  OR2_X1 U3979 ( .A1(n4001), .A2(n4002), .ZN(n2907) );
  AND2_X1 U3980 ( .A1(n3996), .A2(n3995), .ZN(n4002) );
  AND2_X1 U3981 ( .A1(n3993), .A2(n4003), .ZN(n4001) );
  OR2_X1 U3982 ( .A1(n3995), .A2(n3996), .ZN(n4003) );
  OR2_X1 U3983 ( .A1(n2657), .A2(n2674), .ZN(n3996) );
  OR2_X1 U3984 ( .A1(n4004), .A2(n4005), .ZN(n3995) );
  AND2_X1 U3985 ( .A1(n3992), .A2(n3991), .ZN(n4005) );
  AND2_X1 U3986 ( .A1(n3989), .A2(n4006), .ZN(n4004) );
  OR2_X1 U3987 ( .A1(n3991), .A2(n3992), .ZN(n4006) );
  OR2_X1 U3988 ( .A1(n2661), .A2(n2674), .ZN(n3992) );
  OR2_X1 U3989 ( .A1(n4007), .A2(n4008), .ZN(n3991) );
  AND2_X1 U3990 ( .A1(n3988), .A2(n3987), .ZN(n4008) );
  AND2_X1 U3991 ( .A1(n3985), .A2(n4009), .ZN(n4007) );
  OR2_X1 U3992 ( .A1(n3987), .A2(n3988), .ZN(n4009) );
  OR2_X1 U3993 ( .A1(n2665), .A2(n2674), .ZN(n3988) );
  OR2_X1 U3994 ( .A1(n4010), .A2(n4011), .ZN(n3987) );
  AND2_X1 U3995 ( .A1(n3984), .A2(n3983), .ZN(n4011) );
  AND2_X1 U3996 ( .A1(n3981), .A2(n4012), .ZN(n4010) );
  OR2_X1 U3997 ( .A1(n3983), .A2(n3984), .ZN(n4012) );
  OR2_X1 U3998 ( .A1(n2669), .A2(n2674), .ZN(n3984) );
  OR2_X1 U3999 ( .A1(n4013), .A2(n4014), .ZN(n3983) );
  AND2_X1 U4000 ( .A1(n2493), .A2(n3980), .ZN(n4014) );
  AND2_X1 U4001 ( .A1(n3978), .A2(n4015), .ZN(n4013) );
  OR2_X1 U4002 ( .A1(n3980), .A2(n2493), .ZN(n4015) );
  OR2_X1 U4003 ( .A1(n2673), .A2(n2674), .ZN(n2493) );
  OR2_X1 U4004 ( .A1(n4016), .A2(n4017), .ZN(n3980) );
  AND2_X1 U4005 ( .A1(n3977), .A2(n3976), .ZN(n4017) );
  AND2_X1 U4006 ( .A1(n3974), .A2(n4018), .ZN(n4016) );
  OR2_X1 U4007 ( .A1(n3976), .A2(n3977), .ZN(n4018) );
  OR2_X1 U4008 ( .A1(n2677), .A2(n2674), .ZN(n3977) );
  OR2_X1 U4009 ( .A1(n4019), .A2(n4020), .ZN(n3976) );
  AND2_X1 U4010 ( .A1(n3973), .A2(n3972), .ZN(n4020) );
  AND2_X1 U4011 ( .A1(n3970), .A2(n4021), .ZN(n4019) );
  OR2_X1 U4012 ( .A1(n3972), .A2(n3973), .ZN(n4021) );
  OR2_X1 U4013 ( .A1(n2681), .A2(n2674), .ZN(n3973) );
  OR2_X1 U4014 ( .A1(n4022), .A2(n4023), .ZN(n3972) );
  AND2_X1 U4015 ( .A1(n3966), .A2(n3969), .ZN(n4023) );
  AND2_X1 U4016 ( .A1(n4024), .A2(n3968), .ZN(n4022) );
  OR2_X1 U4017 ( .A1(n4025), .A2(n4026), .ZN(n3968) );
  AND2_X1 U4018 ( .A1(n3965), .A2(n3964), .ZN(n4026) );
  AND2_X1 U4019 ( .A1(n3962), .A2(n4027), .ZN(n4025) );
  OR2_X1 U4020 ( .A1(n3964), .A2(n3965), .ZN(n4027) );
  OR2_X1 U4021 ( .A1(n2689), .A2(n2674), .ZN(n3965) );
  OR2_X1 U4022 ( .A1(n4028), .A2(n4029), .ZN(n3964) );
  AND2_X1 U4023 ( .A1(n3958), .A2(n3961), .ZN(n4029) );
  AND2_X1 U4024 ( .A1(n4030), .A2(n3960), .ZN(n4028) );
  OR2_X1 U4025 ( .A1(n4031), .A2(n4032), .ZN(n3960) );
  AND2_X1 U4026 ( .A1(n3954), .A2(n3957), .ZN(n4032) );
  AND2_X1 U4027 ( .A1(n4033), .A2(n3956), .ZN(n4031) );
  OR2_X1 U4028 ( .A1(n4034), .A2(n4035), .ZN(n3956) );
  AND2_X1 U4029 ( .A1(n3951), .A2(n3953), .ZN(n4035) );
  AND2_X1 U4030 ( .A1(n4036), .A2(n3952), .ZN(n4034) );
  OR2_X1 U4031 ( .A1(n4037), .A2(n4038), .ZN(n3952) );
  AND2_X1 U4032 ( .A1(n3946), .A2(n3949), .ZN(n4038) );
  AND2_X1 U4033 ( .A1(n3948), .A2(n4039), .ZN(n4037) );
  OR2_X1 U4034 ( .A1(n3949), .A2(n3946), .ZN(n4039) );
  OR2_X1 U4035 ( .A1(n2705), .A2(n2674), .ZN(n3946) );
  OR2_X1 U4036 ( .A1(n3045), .A2(n4040), .ZN(n3949) );
  OR2_X1 U4037 ( .A1(n2674), .A2(n2670), .ZN(n4040) );
  INV_X1 U4038 ( .A(n4041), .ZN(n3948) );
  OR2_X1 U4039 ( .A1(n4042), .A2(n4043), .ZN(n4041) );
  AND2_X1 U4040 ( .A1(b_4_), .A2(n4044), .ZN(n4043) );
  OR2_X1 U4041 ( .A1(n4045), .A2(n3051), .ZN(n4044) );
  AND2_X1 U4042 ( .A1(a_14_), .A2(n2666), .ZN(n4045) );
  AND2_X1 U4043 ( .A1(b_3_), .A2(n4046), .ZN(n4042) );
  OR2_X1 U4044 ( .A1(n4047), .A2(n2217), .ZN(n4046) );
  AND2_X1 U4045 ( .A1(a_15_), .A2(n2670), .ZN(n4047) );
  OR2_X1 U4046 ( .A1(n3953), .A2(n3951), .ZN(n4036) );
  XNOR2_X1 U4047 ( .A(n4048), .B(n4049), .ZN(n3951) );
  XNOR2_X1 U4048 ( .A(n4050), .B(n4051), .ZN(n4049) );
  OR2_X1 U4049 ( .A1(n2701), .A2(n2674), .ZN(n3953) );
  OR2_X1 U4050 ( .A1(n3957), .A2(n3954), .ZN(n4033) );
  XNOR2_X1 U4051 ( .A(n4052), .B(n4053), .ZN(n3954) );
  XNOR2_X1 U4052 ( .A(n4054), .B(n4055), .ZN(n4052) );
  OR2_X1 U4053 ( .A1(n2697), .A2(n2674), .ZN(n3957) );
  OR2_X1 U4054 ( .A1(n3961), .A2(n3958), .ZN(n4030) );
  XOR2_X1 U4055 ( .A(n4056), .B(n4057), .Z(n3958) );
  XOR2_X1 U4056 ( .A(n4058), .B(n4059), .Z(n4057) );
  OR2_X1 U4057 ( .A1(n2693), .A2(n2674), .ZN(n3961) );
  XOR2_X1 U4058 ( .A(n4060), .B(n4061), .Z(n3962) );
  XOR2_X1 U4059 ( .A(n4062), .B(n4063), .Z(n4061) );
  OR2_X1 U4060 ( .A1(n3969), .A2(n3966), .ZN(n4024) );
  XOR2_X1 U4061 ( .A(n4064), .B(n4065), .Z(n3966) );
  XOR2_X1 U4062 ( .A(n4066), .B(n4067), .Z(n4065) );
  OR2_X1 U4063 ( .A1(n2685), .A2(n2674), .ZN(n3969) );
  INV_X1 U4064 ( .A(b_5_), .ZN(n2674) );
  XOR2_X1 U4065 ( .A(n4068), .B(n4069), .Z(n3970) );
  XOR2_X1 U4066 ( .A(n4070), .B(n4071), .Z(n4069) );
  XOR2_X1 U4067 ( .A(n4072), .B(n4073), .Z(n3974) );
  XOR2_X1 U4068 ( .A(n4074), .B(n4075), .Z(n4073) );
  XOR2_X1 U4069 ( .A(n4076), .B(n4077), .Z(n3978) );
  XOR2_X1 U4070 ( .A(n4078), .B(n4079), .Z(n4077) );
  XOR2_X1 U4071 ( .A(n4080), .B(n4081), .Z(n3981) );
  XOR2_X1 U4072 ( .A(n4082), .B(n4083), .Z(n4081) );
  XOR2_X1 U4073 ( .A(n4084), .B(n4085), .Z(n3985) );
  XOR2_X1 U4074 ( .A(n4086), .B(n2522), .Z(n4085) );
  XOR2_X1 U4075 ( .A(n4087), .B(n4088), .Z(n3989) );
  XOR2_X1 U4076 ( .A(n4089), .B(n4090), .Z(n4088) );
  XOR2_X1 U4077 ( .A(n4091), .B(n4092), .Z(n3993) );
  XOR2_X1 U4078 ( .A(n4093), .B(n4094), .Z(n4092) );
  XOR2_X1 U4079 ( .A(n4095), .B(n4096), .Z(n2905) );
  XOR2_X1 U4080 ( .A(n4097), .B(n4098), .Z(n4096) );
  XOR2_X1 U4081 ( .A(n2880), .B(n4099), .Z(n2890) );
  XOR2_X1 U4082 ( .A(n2879), .B(n2878), .Z(n4099) );
  OR2_X1 U4083 ( .A1(n2815), .A2(n2670), .ZN(n2878) );
  OR2_X1 U4084 ( .A1(n4100), .A2(n4101), .ZN(n2879) );
  AND2_X1 U4085 ( .A1(n4098), .A2(n4097), .ZN(n4101) );
  AND2_X1 U4086 ( .A1(n4095), .A2(n4102), .ZN(n4100) );
  OR2_X1 U4087 ( .A1(n4097), .A2(n4098), .ZN(n4102) );
  OR2_X1 U4088 ( .A1(n2657), .A2(n2670), .ZN(n4098) );
  OR2_X1 U4089 ( .A1(n4103), .A2(n4104), .ZN(n4097) );
  AND2_X1 U4090 ( .A1(n4094), .A2(n4093), .ZN(n4104) );
  AND2_X1 U4091 ( .A1(n4091), .A2(n4105), .ZN(n4103) );
  OR2_X1 U4092 ( .A1(n4093), .A2(n4094), .ZN(n4105) );
  OR2_X1 U4093 ( .A1(n2661), .A2(n2670), .ZN(n4094) );
  OR2_X1 U4094 ( .A1(n4106), .A2(n4107), .ZN(n4093) );
  AND2_X1 U4095 ( .A1(n4090), .A2(n4089), .ZN(n4107) );
  AND2_X1 U4096 ( .A1(n4087), .A2(n4108), .ZN(n4106) );
  OR2_X1 U4097 ( .A1(n4089), .A2(n4090), .ZN(n4108) );
  OR2_X1 U4098 ( .A1(n2665), .A2(n2670), .ZN(n4090) );
  OR2_X1 U4099 ( .A1(n4109), .A2(n4110), .ZN(n4089) );
  AND2_X1 U4100 ( .A1(n2522), .A2(n4086), .ZN(n4110) );
  AND2_X1 U4101 ( .A1(n4084), .A2(n4111), .ZN(n4109) );
  OR2_X1 U4102 ( .A1(n4086), .A2(n2522), .ZN(n4111) );
  OR2_X1 U4103 ( .A1(n2669), .A2(n2670), .ZN(n2522) );
  OR2_X1 U4104 ( .A1(n4112), .A2(n4113), .ZN(n4086) );
  AND2_X1 U4105 ( .A1(n4083), .A2(n4082), .ZN(n4113) );
  AND2_X1 U4106 ( .A1(n4080), .A2(n4114), .ZN(n4112) );
  OR2_X1 U4107 ( .A1(n4082), .A2(n4083), .ZN(n4114) );
  OR2_X1 U4108 ( .A1(n2673), .A2(n2670), .ZN(n4083) );
  OR2_X1 U4109 ( .A1(n4115), .A2(n4116), .ZN(n4082) );
  AND2_X1 U4110 ( .A1(n4079), .A2(n4078), .ZN(n4116) );
  AND2_X1 U4111 ( .A1(n4076), .A2(n4117), .ZN(n4115) );
  OR2_X1 U4112 ( .A1(n4078), .A2(n4079), .ZN(n4117) );
  OR2_X1 U4113 ( .A1(n2677), .A2(n2670), .ZN(n4079) );
  OR2_X1 U4114 ( .A1(n4118), .A2(n4119), .ZN(n4078) );
  AND2_X1 U4115 ( .A1(n4075), .A2(n4074), .ZN(n4119) );
  AND2_X1 U4116 ( .A1(n4072), .A2(n4120), .ZN(n4118) );
  OR2_X1 U4117 ( .A1(n4074), .A2(n4075), .ZN(n4120) );
  OR2_X1 U4118 ( .A1(n2681), .A2(n2670), .ZN(n4075) );
  OR2_X1 U4119 ( .A1(n4121), .A2(n4122), .ZN(n4074) );
  AND2_X1 U4120 ( .A1(n4071), .A2(n4070), .ZN(n4122) );
  AND2_X1 U4121 ( .A1(n4068), .A2(n4123), .ZN(n4121) );
  OR2_X1 U4122 ( .A1(n4070), .A2(n4071), .ZN(n4123) );
  OR2_X1 U4123 ( .A1(n2685), .A2(n2670), .ZN(n4071) );
  OR2_X1 U4124 ( .A1(n4124), .A2(n4125), .ZN(n4070) );
  AND2_X1 U4125 ( .A1(n4064), .A2(n4067), .ZN(n4125) );
  AND2_X1 U4126 ( .A1(n4126), .A2(n4066), .ZN(n4124) );
  OR2_X1 U4127 ( .A1(n4127), .A2(n4128), .ZN(n4066) );
  AND2_X1 U4128 ( .A1(n4063), .A2(n4062), .ZN(n4128) );
  AND2_X1 U4129 ( .A1(n4060), .A2(n4129), .ZN(n4127) );
  OR2_X1 U4130 ( .A1(n4062), .A2(n4063), .ZN(n4129) );
  OR2_X1 U4131 ( .A1(n2693), .A2(n2670), .ZN(n4063) );
  OR2_X1 U4132 ( .A1(n4130), .A2(n4131), .ZN(n4062) );
  AND2_X1 U4133 ( .A1(n4056), .A2(n4059), .ZN(n4131) );
  AND2_X1 U4134 ( .A1(n4132), .A2(n4058), .ZN(n4130) );
  OR2_X1 U4135 ( .A1(n4133), .A2(n4134), .ZN(n4058) );
  AND2_X1 U4136 ( .A1(n4053), .A2(n4055), .ZN(n4134) );
  AND2_X1 U4137 ( .A1(n4135), .A2(n4054), .ZN(n4133) );
  OR2_X1 U4138 ( .A1(n4136), .A2(n4137), .ZN(n4054) );
  AND2_X1 U4139 ( .A1(n4048), .A2(n4051), .ZN(n4137) );
  AND2_X1 U4140 ( .A1(n4050), .A2(n4138), .ZN(n4136) );
  OR2_X1 U4141 ( .A1(n4051), .A2(n4048), .ZN(n4138) );
  OR2_X1 U4142 ( .A1(n2705), .A2(n2670), .ZN(n4048) );
  OR2_X1 U4143 ( .A1(n3045), .A2(n4139), .ZN(n4051) );
  OR2_X1 U4144 ( .A1(n2670), .A2(n2666), .ZN(n4139) );
  INV_X1 U4145 ( .A(n4140), .ZN(n4050) );
  OR2_X1 U4146 ( .A1(n4141), .A2(n4142), .ZN(n4140) );
  AND2_X1 U4147 ( .A1(b_3_), .A2(n4143), .ZN(n4142) );
  OR2_X1 U4148 ( .A1(n4144), .A2(n3051), .ZN(n4143) );
  AND2_X1 U4149 ( .A1(a_14_), .A2(n2662), .ZN(n4144) );
  AND2_X1 U4150 ( .A1(b_2_), .A2(n4145), .ZN(n4141) );
  OR2_X1 U4151 ( .A1(n4146), .A2(n2217), .ZN(n4145) );
  AND2_X1 U4152 ( .A1(a_15_), .A2(n2666), .ZN(n4146) );
  OR2_X1 U4153 ( .A1(n4055), .A2(n4053), .ZN(n4135) );
  XNOR2_X1 U4154 ( .A(n4147), .B(n4148), .ZN(n4053) );
  XNOR2_X1 U4155 ( .A(n4149), .B(n4150), .ZN(n4148) );
  OR2_X1 U4156 ( .A1(n2701), .A2(n2670), .ZN(n4055) );
  OR2_X1 U4157 ( .A1(n4059), .A2(n4056), .ZN(n4132) );
  XNOR2_X1 U4158 ( .A(n4151), .B(n4152), .ZN(n4056) );
  XNOR2_X1 U4159 ( .A(n4153), .B(n4154), .ZN(n4151) );
  OR2_X1 U4160 ( .A1(n2697), .A2(n2670), .ZN(n4059) );
  XOR2_X1 U4161 ( .A(n4155), .B(n4156), .Z(n4060) );
  XOR2_X1 U4162 ( .A(n4157), .B(n4158), .Z(n4156) );
  OR2_X1 U4163 ( .A1(n4067), .A2(n4064), .ZN(n4126) );
  XOR2_X1 U4164 ( .A(n4159), .B(n4160), .Z(n4064) );
  XOR2_X1 U4165 ( .A(n4161), .B(n4162), .Z(n4160) );
  OR2_X1 U4166 ( .A1(n2689), .A2(n2670), .ZN(n4067) );
  INV_X1 U4167 ( .A(b_4_), .ZN(n2670) );
  XOR2_X1 U4168 ( .A(n4163), .B(n4164), .Z(n4068) );
  XOR2_X1 U4169 ( .A(n4165), .B(n4166), .Z(n4164) );
  XOR2_X1 U4170 ( .A(n4167), .B(n4168), .Z(n4072) );
  XOR2_X1 U4171 ( .A(n4169), .B(n4170), .Z(n4168) );
  XOR2_X1 U4172 ( .A(n4171), .B(n4172), .Z(n4076) );
  XOR2_X1 U4173 ( .A(n4173), .B(n4174), .Z(n4172) );
  XOR2_X1 U4174 ( .A(n4175), .B(n4176), .Z(n4080) );
  XOR2_X1 U4175 ( .A(n4177), .B(n4178), .Z(n4176) );
  XOR2_X1 U4176 ( .A(n4179), .B(n4180), .Z(n4084) );
  XOR2_X1 U4177 ( .A(n4181), .B(n4182), .Z(n4180) );
  XOR2_X1 U4178 ( .A(n4183), .B(n4184), .Z(n4087) );
  XOR2_X1 U4179 ( .A(n4185), .B(n4186), .Z(n4184) );
  XOR2_X1 U4180 ( .A(n4187), .B(n4188), .Z(n4091) );
  XOR2_X1 U4181 ( .A(n4189), .B(n2562), .Z(n4188) );
  XOR2_X1 U4182 ( .A(n4190), .B(n4191), .Z(n4095) );
  XOR2_X1 U4183 ( .A(n4192), .B(n4193), .Z(n4191) );
  XOR2_X1 U4184 ( .A(n4194), .B(n4195), .Z(n2880) );
  XOR2_X1 U4185 ( .A(n4196), .B(n4197), .Z(n4195) );
  INV_X1 U4186 ( .A(n4198), .ZN(n2863) );
  OR2_X1 U4187 ( .A1(n2867), .A2(n2868), .ZN(n4198) );
  OR2_X1 U4188 ( .A1(n4199), .A2(n4200), .ZN(n2868) );
  AND2_X1 U4189 ( .A1(n2885), .A2(n2884), .ZN(n4200) );
  AND2_X1 U4190 ( .A1(n2882), .A2(n4201), .ZN(n4199) );
  OR2_X1 U4191 ( .A1(n2884), .A2(n2885), .ZN(n4201) );
  OR2_X1 U4192 ( .A1(n2815), .A2(n2666), .ZN(n2885) );
  OR2_X1 U4193 ( .A1(n4202), .A2(n4203), .ZN(n2884) );
  AND2_X1 U4194 ( .A1(n4197), .A2(n4196), .ZN(n4203) );
  AND2_X1 U4195 ( .A1(n4194), .A2(n4204), .ZN(n4202) );
  OR2_X1 U4196 ( .A1(n4196), .A2(n4197), .ZN(n4204) );
  OR2_X1 U4197 ( .A1(n2657), .A2(n2666), .ZN(n4197) );
  OR2_X1 U4198 ( .A1(n4205), .A2(n4206), .ZN(n4196) );
  AND2_X1 U4199 ( .A1(n4193), .A2(n4192), .ZN(n4206) );
  AND2_X1 U4200 ( .A1(n4190), .A2(n4207), .ZN(n4205) );
  OR2_X1 U4201 ( .A1(n4192), .A2(n4193), .ZN(n4207) );
  OR2_X1 U4202 ( .A1(n2661), .A2(n2666), .ZN(n4193) );
  OR2_X1 U4203 ( .A1(n4208), .A2(n4209), .ZN(n4192) );
  AND2_X1 U4204 ( .A1(n2562), .A2(n4189), .ZN(n4209) );
  AND2_X1 U4205 ( .A1(n4187), .A2(n4210), .ZN(n4208) );
  OR2_X1 U4206 ( .A1(n4189), .A2(n2562), .ZN(n4210) );
  OR2_X1 U4207 ( .A1(n2665), .A2(n2666), .ZN(n2562) );
  OR2_X1 U4208 ( .A1(n4211), .A2(n4212), .ZN(n4189) );
  AND2_X1 U4209 ( .A1(n4186), .A2(n4185), .ZN(n4212) );
  AND2_X1 U4210 ( .A1(n4183), .A2(n4213), .ZN(n4211) );
  OR2_X1 U4211 ( .A1(n4185), .A2(n4186), .ZN(n4213) );
  OR2_X1 U4212 ( .A1(n2669), .A2(n2666), .ZN(n4186) );
  OR2_X1 U4213 ( .A1(n4214), .A2(n4215), .ZN(n4185) );
  AND2_X1 U4214 ( .A1(n4182), .A2(n4181), .ZN(n4215) );
  AND2_X1 U4215 ( .A1(n4179), .A2(n4216), .ZN(n4214) );
  OR2_X1 U4216 ( .A1(n4181), .A2(n4182), .ZN(n4216) );
  OR2_X1 U4217 ( .A1(n2673), .A2(n2666), .ZN(n4182) );
  OR2_X1 U4218 ( .A1(n4217), .A2(n4218), .ZN(n4181) );
  AND2_X1 U4219 ( .A1(n4178), .A2(n4177), .ZN(n4218) );
  AND2_X1 U4220 ( .A1(n4175), .A2(n4219), .ZN(n4217) );
  OR2_X1 U4221 ( .A1(n4177), .A2(n4178), .ZN(n4219) );
  OR2_X1 U4222 ( .A1(n2677), .A2(n2666), .ZN(n4178) );
  OR2_X1 U4223 ( .A1(n4220), .A2(n4221), .ZN(n4177) );
  AND2_X1 U4224 ( .A1(n4174), .A2(n4173), .ZN(n4221) );
  AND2_X1 U4225 ( .A1(n4171), .A2(n4222), .ZN(n4220) );
  OR2_X1 U4226 ( .A1(n4173), .A2(n4174), .ZN(n4222) );
  OR2_X1 U4227 ( .A1(n2681), .A2(n2666), .ZN(n4174) );
  OR2_X1 U4228 ( .A1(n4223), .A2(n4224), .ZN(n4173) );
  AND2_X1 U4229 ( .A1(n4170), .A2(n4169), .ZN(n4224) );
  AND2_X1 U4230 ( .A1(n4167), .A2(n4225), .ZN(n4223) );
  OR2_X1 U4231 ( .A1(n4169), .A2(n4170), .ZN(n4225) );
  OR2_X1 U4232 ( .A1(n2685), .A2(n2666), .ZN(n4170) );
  OR2_X1 U4233 ( .A1(n4226), .A2(n4227), .ZN(n4169) );
  AND2_X1 U4234 ( .A1(n4166), .A2(n4165), .ZN(n4227) );
  AND2_X1 U4235 ( .A1(n4163), .A2(n4228), .ZN(n4226) );
  OR2_X1 U4236 ( .A1(n4165), .A2(n4166), .ZN(n4228) );
  OR2_X1 U4237 ( .A1(n2689), .A2(n2666), .ZN(n4166) );
  OR2_X1 U4238 ( .A1(n4229), .A2(n4230), .ZN(n4165) );
  AND2_X1 U4239 ( .A1(n4159), .A2(n4162), .ZN(n4230) );
  AND2_X1 U4240 ( .A1(n4231), .A2(n4161), .ZN(n4229) );
  OR2_X1 U4241 ( .A1(n4232), .A2(n4233), .ZN(n4161) );
  AND2_X1 U4242 ( .A1(n4158), .A2(n4157), .ZN(n4233) );
  AND2_X1 U4243 ( .A1(n4155), .A2(n4234), .ZN(n4232) );
  OR2_X1 U4244 ( .A1(n4157), .A2(n4158), .ZN(n4234) );
  OR2_X1 U4245 ( .A1(n2697), .A2(n2666), .ZN(n4158) );
  OR2_X1 U4246 ( .A1(n4235), .A2(n4236), .ZN(n4157) );
  AND2_X1 U4247 ( .A1(n4152), .A2(n4154), .ZN(n4236) );
  AND2_X1 U4248 ( .A1(n4237), .A2(n4153), .ZN(n4235) );
  OR2_X1 U4249 ( .A1(n4238), .A2(n4239), .ZN(n4153) );
  AND2_X1 U4250 ( .A1(n4147), .A2(n4150), .ZN(n4239) );
  AND2_X1 U4251 ( .A1(n4149), .A2(n4240), .ZN(n4238) );
  OR2_X1 U4252 ( .A1(n4150), .A2(n4147), .ZN(n4240) );
  OR2_X1 U4253 ( .A1(n2705), .A2(n2666), .ZN(n4147) );
  OR2_X1 U4254 ( .A1(n3045), .A2(n4241), .ZN(n4150) );
  OR2_X1 U4255 ( .A1(n2666), .A2(n2662), .ZN(n4241) );
  INV_X1 U4256 ( .A(n4242), .ZN(n4149) );
  OR2_X1 U4257 ( .A1(n4243), .A2(n4244), .ZN(n4242) );
  AND2_X1 U4258 ( .A1(b_2_), .A2(n4245), .ZN(n4244) );
  OR2_X1 U4259 ( .A1(n4246), .A2(n3051), .ZN(n4245) );
  AND2_X1 U4260 ( .A1(a_14_), .A2(n2658), .ZN(n4246) );
  AND2_X1 U4261 ( .A1(b_1_), .A2(n4247), .ZN(n4243) );
  OR2_X1 U4262 ( .A1(n4248), .A2(n2217), .ZN(n4247) );
  AND2_X1 U4263 ( .A1(a_15_), .A2(n2662), .ZN(n4248) );
  OR2_X1 U4264 ( .A1(n4154), .A2(n4152), .ZN(n4237) );
  XNOR2_X1 U4265 ( .A(n4249), .B(n4250), .ZN(n4152) );
  XNOR2_X1 U4266 ( .A(n4251), .B(n4252), .ZN(n4250) );
  OR2_X1 U4267 ( .A1(n2701), .A2(n2666), .ZN(n4154) );
  XNOR2_X1 U4268 ( .A(n4253), .B(n4254), .ZN(n4155) );
  XNOR2_X1 U4269 ( .A(n4255), .B(n4256), .ZN(n4253) );
  OR2_X1 U4270 ( .A1(n4162), .A2(n4159), .ZN(n4231) );
  XOR2_X1 U4271 ( .A(n4257), .B(n4258), .Z(n4159) );
  XOR2_X1 U4272 ( .A(n4259), .B(n4260), .Z(n4258) );
  OR2_X1 U4273 ( .A1(n2693), .A2(n2666), .ZN(n4162) );
  INV_X1 U4274 ( .A(b_3_), .ZN(n2666) );
  XOR2_X1 U4275 ( .A(n4261), .B(n4262), .Z(n4163) );
  XOR2_X1 U4276 ( .A(n4263), .B(n4264), .Z(n4262) );
  XOR2_X1 U4277 ( .A(n4265), .B(n4266), .Z(n4167) );
  XOR2_X1 U4278 ( .A(n4267), .B(n4268), .Z(n4266) );
  XOR2_X1 U4279 ( .A(n4269), .B(n4270), .Z(n4171) );
  XOR2_X1 U4280 ( .A(n4271), .B(n4272), .Z(n4270) );
  XOR2_X1 U4281 ( .A(n4273), .B(n4274), .Z(n4175) );
  XOR2_X1 U4282 ( .A(n4275), .B(n4276), .Z(n4274) );
  XOR2_X1 U4283 ( .A(n4277), .B(n4278), .Z(n4179) );
  XOR2_X1 U4284 ( .A(n4279), .B(n4280), .Z(n4278) );
  XOR2_X1 U4285 ( .A(n4281), .B(n4282), .Z(n4183) );
  XOR2_X1 U4286 ( .A(n4283), .B(n4284), .Z(n4282) );
  XOR2_X1 U4287 ( .A(n4285), .B(n4286), .Z(n4187) );
  XOR2_X1 U4288 ( .A(n4287), .B(n4288), .Z(n4286) );
  XOR2_X1 U4289 ( .A(n4289), .B(n4290), .Z(n4190) );
  XOR2_X1 U4290 ( .A(n4291), .B(n4292), .Z(n4290) );
  XOR2_X1 U4291 ( .A(n4293), .B(n4294), .Z(n4194) );
  XOR2_X1 U4292 ( .A(n4295), .B(n2591), .Z(n4294) );
  XOR2_X1 U4293 ( .A(n4296), .B(n4297), .Z(n2882) );
  XOR2_X1 U4294 ( .A(n4298), .B(n4299), .Z(n4297) );
  XOR2_X1 U4295 ( .A(n4300), .B(n4301), .Z(n2867) );
  XOR2_X1 U4296 ( .A(n4302), .B(n4303), .Z(n4301) );
  AND2_X1 U4297 ( .A1(n2541), .A2(n4304), .ZN(n2543) );
  AND2_X1 U4298 ( .A1(n2542), .A2(n2540), .ZN(n4304) );
  XOR2_X1 U4299 ( .A(n4305), .B(n4306), .Z(n2540) );
  OR2_X1 U4300 ( .A1(n4307), .A2(n2815), .ZN(n4305) );
  XNOR2_X1 U4301 ( .A(n4308), .B(n4309), .ZN(n2542) );
  XOR2_X1 U4302 ( .A(n4310), .B(n4311), .Z(n4309) );
  INV_X1 U4303 ( .A(n2862), .ZN(n2541) );
  OR2_X1 U4304 ( .A1(n4312), .A2(n4313), .ZN(n2862) );
  AND2_X1 U4305 ( .A1(n4303), .A2(n4302), .ZN(n4313) );
  AND2_X1 U4306 ( .A1(n4300), .A2(n4314), .ZN(n4312) );
  OR2_X1 U4307 ( .A1(n4302), .A2(n4303), .ZN(n4314) );
  OR2_X1 U4308 ( .A1(n2815), .A2(n2662), .ZN(n4303) );
  OR2_X1 U4309 ( .A1(n4315), .A2(n4316), .ZN(n4302) );
  AND2_X1 U4310 ( .A1(n4299), .A2(n4298), .ZN(n4316) );
  AND2_X1 U4311 ( .A1(n4296), .A2(n4317), .ZN(n4315) );
  OR2_X1 U4312 ( .A1(n4298), .A2(n4299), .ZN(n4317) );
  OR2_X1 U4313 ( .A1(n2657), .A2(n2662), .ZN(n4299) );
  OR2_X1 U4314 ( .A1(n4318), .A2(n4319), .ZN(n4298) );
  AND2_X1 U4315 ( .A1(n2591), .A2(n4295), .ZN(n4319) );
  AND2_X1 U4316 ( .A1(n4293), .A2(n4320), .ZN(n4318) );
  OR2_X1 U4317 ( .A1(n4295), .A2(n2591), .ZN(n4320) );
  OR2_X1 U4318 ( .A1(n2661), .A2(n2662), .ZN(n2591) );
  OR2_X1 U4319 ( .A1(n4321), .A2(n4322), .ZN(n4295) );
  AND2_X1 U4320 ( .A1(n4292), .A2(n4291), .ZN(n4322) );
  AND2_X1 U4321 ( .A1(n4289), .A2(n4323), .ZN(n4321) );
  OR2_X1 U4322 ( .A1(n4291), .A2(n4292), .ZN(n4323) );
  OR2_X1 U4323 ( .A1(n2665), .A2(n2662), .ZN(n4292) );
  OR2_X1 U4324 ( .A1(n4324), .A2(n4325), .ZN(n4291) );
  AND2_X1 U4325 ( .A1(n4288), .A2(n4287), .ZN(n4325) );
  AND2_X1 U4326 ( .A1(n4285), .A2(n4326), .ZN(n4324) );
  OR2_X1 U4327 ( .A1(n4287), .A2(n4288), .ZN(n4326) );
  OR2_X1 U4328 ( .A1(n2669), .A2(n2662), .ZN(n4288) );
  OR2_X1 U4329 ( .A1(n4327), .A2(n4328), .ZN(n4287) );
  AND2_X1 U4330 ( .A1(n4284), .A2(n4283), .ZN(n4328) );
  AND2_X1 U4331 ( .A1(n4281), .A2(n4329), .ZN(n4327) );
  OR2_X1 U4332 ( .A1(n4283), .A2(n4284), .ZN(n4329) );
  OR2_X1 U4333 ( .A1(n2673), .A2(n2662), .ZN(n4284) );
  OR2_X1 U4334 ( .A1(n4330), .A2(n4331), .ZN(n4283) );
  AND2_X1 U4335 ( .A1(n4280), .A2(n4279), .ZN(n4331) );
  AND2_X1 U4336 ( .A1(n4277), .A2(n4332), .ZN(n4330) );
  OR2_X1 U4337 ( .A1(n4279), .A2(n4280), .ZN(n4332) );
  OR2_X1 U4338 ( .A1(n2677), .A2(n2662), .ZN(n4280) );
  OR2_X1 U4339 ( .A1(n4333), .A2(n4334), .ZN(n4279) );
  AND2_X1 U4340 ( .A1(n4276), .A2(n4275), .ZN(n4334) );
  AND2_X1 U4341 ( .A1(n4273), .A2(n4335), .ZN(n4333) );
  OR2_X1 U4342 ( .A1(n4275), .A2(n4276), .ZN(n4335) );
  OR2_X1 U4343 ( .A1(n2681), .A2(n2662), .ZN(n4276) );
  OR2_X1 U4344 ( .A1(n4336), .A2(n4337), .ZN(n4275) );
  AND2_X1 U4345 ( .A1(n4272), .A2(n4271), .ZN(n4337) );
  AND2_X1 U4346 ( .A1(n4269), .A2(n4338), .ZN(n4336) );
  OR2_X1 U4347 ( .A1(n4271), .A2(n4272), .ZN(n4338) );
  OR2_X1 U4348 ( .A1(n2685), .A2(n2662), .ZN(n4272) );
  OR2_X1 U4349 ( .A1(n4339), .A2(n4340), .ZN(n4271) );
  AND2_X1 U4350 ( .A1(n4268), .A2(n4267), .ZN(n4340) );
  AND2_X1 U4351 ( .A1(n4265), .A2(n4341), .ZN(n4339) );
  OR2_X1 U4352 ( .A1(n4267), .A2(n4268), .ZN(n4341) );
  OR2_X1 U4353 ( .A1(n2689), .A2(n2662), .ZN(n4268) );
  OR2_X1 U4354 ( .A1(n4342), .A2(n4343), .ZN(n4267) );
  AND2_X1 U4355 ( .A1(n4264), .A2(n4263), .ZN(n4343) );
  AND2_X1 U4356 ( .A1(n4261), .A2(n4344), .ZN(n4342) );
  OR2_X1 U4357 ( .A1(n4263), .A2(n4264), .ZN(n4344) );
  OR2_X1 U4358 ( .A1(n2693), .A2(n2662), .ZN(n4264) );
  OR2_X1 U4359 ( .A1(n4345), .A2(n4346), .ZN(n4263) );
  AND2_X1 U4360 ( .A1(n4257), .A2(n4260), .ZN(n4346) );
  AND2_X1 U4361 ( .A1(n4347), .A2(n4259), .ZN(n4345) );
  OR2_X1 U4362 ( .A1(n4348), .A2(n4349), .ZN(n4259) );
  AND2_X1 U4363 ( .A1(n4256), .A2(n4255), .ZN(n4349) );
  AND2_X1 U4364 ( .A1(n4254), .A2(n4350), .ZN(n4348) );
  OR2_X1 U4365 ( .A1(n4255), .A2(n4256), .ZN(n4350) );
  OR2_X1 U4366 ( .A1(n2701), .A2(n2662), .ZN(n4256) );
  OR2_X1 U4367 ( .A1(n4351), .A2(n4352), .ZN(n4255) );
  AND2_X1 U4368 ( .A1(n4249), .A2(n4252), .ZN(n4352) );
  AND2_X1 U4369 ( .A1(n4251), .A2(n4353), .ZN(n4351) );
  OR2_X1 U4370 ( .A1(n4252), .A2(n4249), .ZN(n4353) );
  OR2_X1 U4371 ( .A1(n2705), .A2(n2662), .ZN(n4249) );
  OR2_X1 U4372 ( .A1(n3045), .A2(n4354), .ZN(n4252) );
  OR2_X1 U4373 ( .A1(n2662), .A2(n2658), .ZN(n4354) );
  INV_X1 U4374 ( .A(n4355), .ZN(n4251) );
  OR2_X1 U4375 ( .A1(n4356), .A2(n4357), .ZN(n4355) );
  AND2_X1 U4376 ( .A1(b_1_), .A2(n4358), .ZN(n4357) );
  OR2_X1 U4377 ( .A1(n4359), .A2(n3051), .ZN(n4358) );
  AND2_X1 U4378 ( .A1(n2812), .A2(a_14_), .ZN(n3051) );
  AND2_X1 U4379 ( .A1(a_14_), .A2(n4307), .ZN(n4359) );
  AND2_X1 U4380 ( .A1(b_0_), .A2(n4360), .ZN(n4356) );
  OR2_X1 U4381 ( .A1(n4361), .A2(n2217), .ZN(n4360) );
  AND2_X1 U4382 ( .A1(n2239), .A2(a_15_), .ZN(n2217) );
  AND2_X1 U4383 ( .A1(a_15_), .A2(n2658), .ZN(n4361) );
  XOR2_X1 U4384 ( .A(n4362), .B(n4363), .Z(n4254) );
  XOR2_X1 U4385 ( .A(n4364), .B(n4365), .Z(n4362) );
  OR2_X1 U4386 ( .A1(n4260), .A2(n4257), .ZN(n4347) );
  XOR2_X1 U4387 ( .A(n4366), .B(n4367), .Z(n4257) );
  XOR2_X1 U4388 ( .A(n4368), .B(n4369), .Z(n4366) );
  OR2_X1 U4389 ( .A1(n2697), .A2(n2662), .ZN(n4260) );
  INV_X1 U4390 ( .A(b_2_), .ZN(n2662) );
  XNOR2_X1 U4391 ( .A(n4370), .B(n4371), .ZN(n4261) );
  XNOR2_X1 U4392 ( .A(n4372), .B(n4373), .ZN(n4370) );
  XNOR2_X1 U4393 ( .A(n4374), .B(n4375), .ZN(n4265) );
  XNOR2_X1 U4394 ( .A(n4376), .B(n4377), .ZN(n4374) );
  XNOR2_X1 U4395 ( .A(n4378), .B(n4379), .ZN(n4269) );
  XNOR2_X1 U4396 ( .A(n4380), .B(n4381), .ZN(n4378) );
  XOR2_X1 U4397 ( .A(n4382), .B(n4383), .Z(n4273) );
  XOR2_X1 U4398 ( .A(n4384), .B(n4385), .Z(n4383) );
  XOR2_X1 U4399 ( .A(n4386), .B(n4387), .Z(n4277) );
  XOR2_X1 U4400 ( .A(n4388), .B(n4389), .Z(n4387) );
  XOR2_X1 U4401 ( .A(n4390), .B(n4391), .Z(n4281) );
  XOR2_X1 U4402 ( .A(n4392), .B(n4393), .Z(n4391) );
  XOR2_X1 U4403 ( .A(n4394), .B(n4395), .Z(n4285) );
  XOR2_X1 U4404 ( .A(n4396), .B(n4397), .Z(n4395) );
  XOR2_X1 U4405 ( .A(n4398), .B(n4399), .Z(n4289) );
  XOR2_X1 U4406 ( .A(n4400), .B(n4401), .Z(n4399) );
  XOR2_X1 U4407 ( .A(n4402), .B(n4403), .Z(n4293) );
  XOR2_X1 U4408 ( .A(n4404), .B(n4405), .Z(n4403) );
  XOR2_X1 U4409 ( .A(n4406), .B(n4407), .Z(n4296) );
  XOR2_X1 U4410 ( .A(n4408), .B(n4409), .Z(n4407) );
  XOR2_X1 U4411 ( .A(n4410), .B(n4411), .Z(n4300) );
  XOR2_X1 U4412 ( .A(n4412), .B(n2620), .Z(n4411) );
  AND2_X1 U4413 ( .A1(n4413), .A2(a_0_), .ZN(n2859) );
  INV_X1 U4414 ( .A(n4306), .ZN(n4413) );
  OR2_X1 U4415 ( .A1(n4414), .A2(n4415), .ZN(n4306) );
  AND2_X1 U4416 ( .A1(n4308), .A2(n4310), .ZN(n4415) );
  AND2_X1 U4417 ( .A1(n4416), .A2(n4311), .ZN(n4414) );
  OR2_X1 U4418 ( .A1(n2815), .A2(n2658), .ZN(n4311) );
  INV_X1 U4419 ( .A(a_0_), .ZN(n2815) );
  OR2_X1 U4420 ( .A1(n4310), .A2(n4308), .ZN(n4416) );
  OR2_X1 U4421 ( .A1(n4307), .A2(n2657), .ZN(n4308) );
  OR2_X1 U4422 ( .A1(n4417), .A2(n4418), .ZN(n4310) );
  AND2_X1 U4423 ( .A1(n4410), .A2(n4412), .ZN(n4418) );
  AND2_X1 U4424 ( .A1(n4419), .A2(n2620), .ZN(n4417) );
  OR2_X1 U4425 ( .A1(n2657), .A2(n2658), .ZN(n2620) );
  INV_X1 U4426 ( .A(a_1_), .ZN(n2657) );
  OR2_X1 U4427 ( .A1(n4412), .A2(n4410), .ZN(n4419) );
  OR2_X1 U4428 ( .A1(n4307), .A2(n2661), .ZN(n4410) );
  OR2_X1 U4429 ( .A1(n4420), .A2(n4421), .ZN(n4412) );
  AND2_X1 U4430 ( .A1(n4406), .A2(n4408), .ZN(n4421) );
  AND2_X1 U4431 ( .A1(n4422), .A2(n4409), .ZN(n4420) );
  OR2_X1 U4432 ( .A1(n4307), .A2(n2665), .ZN(n4409) );
  OR2_X1 U4433 ( .A1(n4408), .A2(n4406), .ZN(n4422) );
  OR2_X1 U4434 ( .A1(n2661), .A2(n2658), .ZN(n4406) );
  INV_X1 U4435 ( .A(a_2_), .ZN(n2661) );
  OR2_X1 U4436 ( .A1(n4423), .A2(n4424), .ZN(n4408) );
  AND2_X1 U4437 ( .A1(n4402), .A2(n4404), .ZN(n4424) );
  AND2_X1 U4438 ( .A1(n4425), .A2(n4405), .ZN(n4423) );
  OR2_X1 U4439 ( .A1(n4307), .A2(n2669), .ZN(n4405) );
  OR2_X1 U4440 ( .A1(n4404), .A2(n4402), .ZN(n4425) );
  OR2_X1 U4441 ( .A1(n2665), .A2(n2658), .ZN(n4402) );
  INV_X1 U4442 ( .A(a_3_), .ZN(n2665) );
  OR2_X1 U4443 ( .A1(n4426), .A2(n4427), .ZN(n4404) );
  AND2_X1 U4444 ( .A1(n4398), .A2(n4400), .ZN(n4427) );
  AND2_X1 U4445 ( .A1(n4428), .A2(n4401), .ZN(n4426) );
  OR2_X1 U4446 ( .A1(n4307), .A2(n2673), .ZN(n4401) );
  OR2_X1 U4447 ( .A1(n4400), .A2(n4398), .ZN(n4428) );
  OR2_X1 U4448 ( .A1(n2669), .A2(n2658), .ZN(n4398) );
  INV_X1 U4449 ( .A(a_4_), .ZN(n2669) );
  OR2_X1 U4450 ( .A1(n4429), .A2(n4430), .ZN(n4400) );
  AND2_X1 U4451 ( .A1(n4394), .A2(n4396), .ZN(n4430) );
  AND2_X1 U4452 ( .A1(n4431), .A2(n4397), .ZN(n4429) );
  OR2_X1 U4453 ( .A1(n4307), .A2(n2677), .ZN(n4397) );
  OR2_X1 U4454 ( .A1(n4396), .A2(n4394), .ZN(n4431) );
  OR2_X1 U4455 ( .A1(n2673), .A2(n2658), .ZN(n4394) );
  INV_X1 U4456 ( .A(a_5_), .ZN(n2673) );
  OR2_X1 U4457 ( .A1(n4432), .A2(n4433), .ZN(n4396) );
  AND2_X1 U4458 ( .A1(n4390), .A2(n4392), .ZN(n4433) );
  AND2_X1 U4459 ( .A1(n4434), .A2(n4393), .ZN(n4432) );
  OR2_X1 U4460 ( .A1(n4307), .A2(n2681), .ZN(n4393) );
  OR2_X1 U4461 ( .A1(n4392), .A2(n4390), .ZN(n4434) );
  OR2_X1 U4462 ( .A1(n2677), .A2(n2658), .ZN(n4390) );
  INV_X1 U4463 ( .A(a_6_), .ZN(n2677) );
  OR2_X1 U4464 ( .A1(n4435), .A2(n4436), .ZN(n4392) );
  AND2_X1 U4465 ( .A1(n4386), .A2(n4388), .ZN(n4436) );
  AND2_X1 U4466 ( .A1(n4437), .A2(n4389), .ZN(n4435) );
  OR2_X1 U4467 ( .A1(n4307), .A2(n2685), .ZN(n4389) );
  OR2_X1 U4468 ( .A1(n4388), .A2(n4386), .ZN(n4437) );
  OR2_X1 U4469 ( .A1(n2681), .A2(n2658), .ZN(n4386) );
  INV_X1 U4470 ( .A(a_7_), .ZN(n2681) );
  OR2_X1 U4471 ( .A1(n4438), .A2(n4439), .ZN(n4388) );
  AND2_X1 U4472 ( .A1(n4382), .A2(n4384), .ZN(n4439) );
  AND2_X1 U4473 ( .A1(n4440), .A2(n4385), .ZN(n4438) );
  OR2_X1 U4474 ( .A1(n4307), .A2(n2689), .ZN(n4385) );
  OR2_X1 U4475 ( .A1(n4384), .A2(n4382), .ZN(n4440) );
  OR2_X1 U4476 ( .A1(n2685), .A2(n2658), .ZN(n4382) );
  INV_X1 U4477 ( .A(a_8_), .ZN(n2685) );
  OR2_X1 U4478 ( .A1(n4441), .A2(n4442), .ZN(n4384) );
  AND2_X1 U4479 ( .A1(n4379), .A2(n4381), .ZN(n4442) );
  AND2_X1 U4480 ( .A1(n4443), .A2(n4380), .ZN(n4441) );
  OR2_X1 U4481 ( .A1(n4307), .A2(n2693), .ZN(n4380) );
  OR2_X1 U4482 ( .A1(n4381), .A2(n4379), .ZN(n4443) );
  OR2_X1 U4483 ( .A1(n2689), .A2(n2658), .ZN(n4379) );
  INV_X1 U4484 ( .A(a_9_), .ZN(n2689) );
  OR2_X1 U4485 ( .A1(n4444), .A2(n4445), .ZN(n4381) );
  AND2_X1 U4486 ( .A1(n4375), .A2(n4377), .ZN(n4445) );
  AND2_X1 U4487 ( .A1(n4446), .A2(n4376), .ZN(n4444) );
  OR2_X1 U4488 ( .A1(n4307), .A2(n2697), .ZN(n4376) );
  OR2_X1 U4489 ( .A1(n4377), .A2(n4375), .ZN(n4446) );
  OR2_X1 U4490 ( .A1(n2693), .A2(n2658), .ZN(n4375) );
  INV_X1 U4491 ( .A(a_10_), .ZN(n2693) );
  OR2_X1 U4492 ( .A1(n4447), .A2(n4448), .ZN(n4377) );
  AND2_X1 U4493 ( .A1(n4371), .A2(n4373), .ZN(n4448) );
  AND2_X1 U4494 ( .A1(n4449), .A2(n4372), .ZN(n4447) );
  OR2_X1 U4495 ( .A1(n4307), .A2(n2701), .ZN(n4372) );
  OR2_X1 U4496 ( .A1(n4373), .A2(n4371), .ZN(n4449) );
  OR2_X1 U4497 ( .A1(n2697), .A2(n2658), .ZN(n4371) );
  INV_X1 U4498 ( .A(a_11_), .ZN(n2697) );
  OR2_X1 U4499 ( .A1(n4450), .A2(n4451), .ZN(n4373) );
  AND2_X1 U4500 ( .A1(n4367), .A2(n4369), .ZN(n4451) );
  AND2_X1 U4501 ( .A1(n4368), .A2(n4452), .ZN(n4450) );
  OR2_X1 U4502 ( .A1(n4369), .A2(n4367), .ZN(n4452) );
  OR2_X1 U4503 ( .A1(n2701), .A2(n2658), .ZN(n4367) );
  INV_X1 U4504 ( .A(a_12_), .ZN(n2701) );
  OR2_X1 U4505 ( .A1(n4307), .A2(n2705), .ZN(n4369) );
  INV_X1 U4506 ( .A(a_13_), .ZN(n2705) );
  AND2_X1 U4507 ( .A1(n4453), .A2(n4365), .ZN(n4368) );
  OR2_X1 U4508 ( .A1(n3045), .A2(n4454), .ZN(n4365) );
  OR2_X1 U4509 ( .A1(n4307), .A2(n2658), .ZN(n4454) );
  INV_X1 U4510 ( .A(b_1_), .ZN(n2658) );
  INV_X1 U4511 ( .A(b_0_), .ZN(n4307) );
  OR2_X1 U4512 ( .A1(n2812), .A2(n2239), .ZN(n3045) );
  INV_X1 U4513 ( .A(a_14_), .ZN(n2239) );
  INV_X1 U4514 ( .A(a_15_), .ZN(n2812) );
  INV_X1 U4515 ( .A(n4455), .ZN(n4453) );
  AND2_X1 U4516 ( .A1(n4363), .A2(n4364), .ZN(n4455) );
  AND2_X1 U4517 ( .A1(a_13_), .A2(b_1_), .ZN(n4364) );
  AND2_X1 U4518 ( .A1(a_14_), .A2(b_0_), .ZN(n4363) );
  AND2_X1 U4519 ( .A1(operation_0_), .A2(operation_1_), .ZN(n2173) );
endmodule

