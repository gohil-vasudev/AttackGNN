module add_mul_sub_4_bit ( a_0_, a_1_, a_2_, a_3_, b_0_, b_1_, b_2_, b_3_, 
        operation_0_, operation_1_, Result_0_, Result_1_, Result_2_, Result_3_, 
        Result_4_, Result_5_, Result_6_, Result_7_ );
  input a_0_, a_1_, a_2_, a_3_, b_0_, b_1_, b_2_, b_3_, operation_0_,
         operation_1_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_;
  wire   n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386;

  OR2_X1 U186 ( .A1(n178), .A2(n179), .ZN(Result_7_) );
  AND2_X1 U187 ( .A1(n180), .A2(n181), .ZN(n179) );
  INV_X1 U188 ( .A(n182), .ZN(n181) );
  OR2_X1 U189 ( .A1(n183), .A2(n184), .ZN(n180) );
  AND2_X1 U190 ( .A1(n182), .A2(n185), .ZN(n178) );
  OR2_X1 U191 ( .A1(n186), .A2(n187), .ZN(Result_6_) );
  OR2_X1 U192 ( .A1(n188), .A2(n189), .ZN(n187) );
  AND2_X1 U193 ( .A1(n190), .A2(n191), .ZN(n189) );
  OR2_X1 U194 ( .A1(n192), .A2(n193), .ZN(n190) );
  AND2_X1 U195 ( .A1(a_2_), .A2(n194), .ZN(n193) );
  OR2_X1 U196 ( .A1(n195), .A2(n196), .ZN(n194) );
  AND2_X1 U197 ( .A1(n182), .A2(b_3_), .ZN(n195) );
  AND2_X1 U198 ( .A1(n197), .A2(n198), .ZN(n192) );
  AND2_X1 U199 ( .A1(b_2_), .A2(n199), .ZN(n188) );
  OR2_X1 U200 ( .A1(n200), .A2(n201), .ZN(n199) );
  OR2_X1 U201 ( .A1(n202), .A2(n203), .ZN(n201) );
  AND2_X1 U202 ( .A1(n204), .A2(n198), .ZN(n203) );
  OR2_X1 U203 ( .A1(n205), .A2(n196), .ZN(n204) );
  OR2_X1 U204 ( .A1(n206), .A2(n207), .ZN(n196) );
  OR2_X1 U205 ( .A1(n208), .A2(n209), .ZN(n207) );
  AND2_X1 U206 ( .A1(n210), .A2(n211), .ZN(n209) );
  INV_X1 U207 ( .A(n183), .ZN(n211) );
  AND2_X1 U208 ( .A1(n212), .A2(n213), .ZN(n208) );
  AND2_X1 U209 ( .A1(n214), .A2(n215), .ZN(n206) );
  INV_X1 U210 ( .A(n184), .ZN(n215) );
  AND2_X1 U211 ( .A1(n182), .A2(a_3_), .ZN(n205) );
  AND2_X1 U212 ( .A1(a_2_), .A2(n197), .ZN(n202) );
  OR2_X1 U213 ( .A1(n216), .A2(n217), .ZN(n197) );
  OR2_X1 U214 ( .A1(n218), .A2(n219), .ZN(n217) );
  AND2_X1 U215 ( .A1(n183), .A2(n210), .ZN(n219) );
  AND2_X1 U216 ( .A1(n212), .A2(n185), .ZN(n218) );
  AND2_X1 U217 ( .A1(n214), .A2(n184), .ZN(n216) );
  AND2_X1 U218 ( .A1(n183), .A2(n182), .ZN(n200) );
  AND2_X1 U219 ( .A1(n220), .A2(a_2_), .ZN(n186) );
  AND2_X1 U220 ( .A1(n184), .A2(n182), .ZN(n220) );
  OR2_X1 U221 ( .A1(n221), .A2(n222), .ZN(Result_5_) );
  OR2_X1 U222 ( .A1(n223), .A2(n224), .ZN(n222) );
  AND2_X1 U223 ( .A1(n225), .A2(n226), .ZN(n224) );
  OR2_X1 U224 ( .A1(n227), .A2(n228), .ZN(n226) );
  OR2_X1 U225 ( .A1(n229), .A2(n230), .ZN(n228) );
  AND2_X1 U226 ( .A1(n210), .A2(n231), .ZN(n230) );
  AND2_X1 U227 ( .A1(n212), .A2(n232), .ZN(n229) );
  AND2_X1 U228 ( .A1(n214), .A2(n233), .ZN(n227) );
  INV_X1 U229 ( .A(n234), .ZN(n225) );
  AND2_X1 U230 ( .A1(n234), .A2(n235), .ZN(n223) );
  OR2_X1 U231 ( .A1(n236), .A2(n237), .ZN(n235) );
  OR2_X1 U232 ( .A1(n238), .A2(n239), .ZN(n237) );
  AND2_X1 U233 ( .A1(n240), .A2(n210), .ZN(n239) );
  INV_X1 U234 ( .A(n231), .ZN(n240) );
  AND2_X1 U235 ( .A1(n241), .A2(n212), .ZN(n238) );
  INV_X1 U236 ( .A(n232), .ZN(n241) );
  AND2_X1 U237 ( .A1(n242), .A2(n214), .ZN(n236) );
  INV_X1 U238 ( .A(n233), .ZN(n242) );
  XNOR2_X1 U239 ( .A(b_1_), .B(n243), .ZN(n234) );
  AND2_X1 U240 ( .A1(n182), .A2(n244), .ZN(n221) );
  XOR2_X1 U241 ( .A(n245), .B(n246), .Z(n244) );
  XNOR2_X1 U242 ( .A(n247), .B(n248), .ZN(n246) );
  OR2_X1 U243 ( .A1(n249), .A2(n250), .ZN(Result_4_) );
  OR2_X1 U244 ( .A1(n251), .A2(n252), .ZN(n250) );
  AND2_X1 U245 ( .A1(n253), .A2(n254), .ZN(n252) );
  INV_X1 U246 ( .A(n255), .ZN(n254) );
  OR2_X1 U247 ( .A1(n256), .A2(n257), .ZN(n253) );
  OR2_X1 U248 ( .A1(n258), .A2(n259), .ZN(n257) );
  AND2_X1 U249 ( .A1(n260), .A2(n210), .ZN(n259) );
  INV_X1 U250 ( .A(n261), .ZN(n260) );
  AND2_X1 U251 ( .A1(n262), .A2(n212), .ZN(n258) );
  INV_X1 U252 ( .A(n263), .ZN(n262) );
  AND2_X1 U253 ( .A1(n264), .A2(n214), .ZN(n256) );
  INV_X1 U254 ( .A(n265), .ZN(n264) );
  AND2_X1 U255 ( .A1(n255), .A2(n266), .ZN(n251) );
  OR2_X1 U256 ( .A1(n267), .A2(n268), .ZN(n266) );
  OR2_X1 U257 ( .A1(n269), .A2(n270), .ZN(n268) );
  AND2_X1 U258 ( .A1(n210), .A2(n261), .ZN(n270) );
  AND2_X1 U259 ( .A1(n212), .A2(n263), .ZN(n269) );
  OR2_X1 U260 ( .A1(n271), .A2(n272), .ZN(n263) );
  AND2_X1 U261 ( .A1(a_1_), .A2(n232), .ZN(n272) );
  AND2_X1 U262 ( .A1(b_1_), .A2(n273), .ZN(n271) );
  OR2_X1 U263 ( .A1(a_1_), .A2(n232), .ZN(n273) );
  OR2_X1 U264 ( .A1(n274), .A2(n275), .ZN(n232) );
  AND2_X1 U265 ( .A1(a_2_), .A2(n185), .ZN(n275) );
  AND2_X1 U266 ( .A1(b_2_), .A2(n276), .ZN(n274) );
  OR2_X1 U267 ( .A1(n185), .A2(a_2_), .ZN(n276) );
  AND2_X1 U268 ( .A1(n277), .A2(n278), .ZN(n212) );
  AND2_X1 U269 ( .A1(n214), .A2(n265), .ZN(n267) );
  AND2_X1 U270 ( .A1(n279), .A2(n280), .ZN(n255) );
  AND2_X1 U271 ( .A1(n182), .A2(n281), .ZN(n249) );
  XNOR2_X1 U272 ( .A(n282), .B(n283), .ZN(n281) );
  XOR2_X1 U273 ( .A(n284), .B(n285), .Z(n283) );
  OR2_X1 U274 ( .A1(n286), .A2(n287), .ZN(Result_3_) );
  AND2_X1 U275 ( .A1(n182), .A2(n288), .ZN(n286) );
  XNOR2_X1 U276 ( .A(n289), .B(n290), .ZN(n288) );
  OR2_X1 U277 ( .A1(n291), .A2(n287), .ZN(Result_2_) );
  AND2_X1 U278 ( .A1(n292), .A2(n182), .ZN(n291) );
  XOR2_X1 U279 ( .A(n293), .B(n294), .Z(n292) );
  OR2_X1 U280 ( .A1(n295), .A2(n287), .ZN(Result_1_) );
  AND2_X1 U281 ( .A1(n182), .A2(n296), .ZN(n295) );
  XNOR2_X1 U282 ( .A(n297), .B(n298), .ZN(n296) );
  OR2_X1 U283 ( .A1(n299), .A2(n287), .ZN(Result_0_) );
  OR2_X1 U284 ( .A1(n300), .A2(n301), .ZN(n287) );
  AND2_X1 U285 ( .A1(n214), .A2(n302), .ZN(n301) );
  OR2_X1 U286 ( .A1(n303), .A2(n304), .ZN(n302) );
  AND2_X1 U287 ( .A1(n265), .A2(n279), .ZN(n303) );
  INV_X1 U288 ( .A(n305), .ZN(n279) );
  OR2_X1 U289 ( .A1(n306), .A2(n307), .ZN(n265) );
  AND2_X1 U290 ( .A1(n233), .A2(n243), .ZN(n307) );
  AND2_X1 U291 ( .A1(b_1_), .A2(n308), .ZN(n306) );
  OR2_X1 U292 ( .A1(n243), .A2(n233), .ZN(n308) );
  OR2_X1 U293 ( .A1(n309), .A2(n310), .ZN(n233) );
  AND2_X1 U294 ( .A1(n184), .A2(n198), .ZN(n310) );
  AND2_X1 U295 ( .A1(b_2_), .A2(n311), .ZN(n309) );
  OR2_X1 U296 ( .A1(n184), .A2(n198), .ZN(n311) );
  AND2_X1 U297 ( .A1(n312), .A2(b_3_), .ZN(n184) );
  AND2_X1 U298 ( .A1(n278), .A2(operation_1_), .ZN(n214) );
  INV_X1 U299 ( .A(operation_0_), .ZN(n278) );
  AND2_X1 U300 ( .A1(n313), .A2(n210), .ZN(n300) );
  AND2_X1 U301 ( .A1(n277), .A2(operation_0_), .ZN(n210) );
  INV_X1 U302 ( .A(operation_1_), .ZN(n277) );
  AND2_X1 U303 ( .A1(n314), .A2(n280), .ZN(n313) );
  INV_X1 U304 ( .A(n304), .ZN(n280) );
  AND2_X1 U305 ( .A1(n315), .A2(b_0_), .ZN(n304) );
  OR2_X1 U306 ( .A1(n305), .A2(n261), .ZN(n314) );
  OR2_X1 U307 ( .A1(n316), .A2(n317), .ZN(n261) );
  AND2_X1 U308 ( .A1(a_1_), .A2(n231), .ZN(n317) );
  AND2_X1 U309 ( .A1(n318), .A2(n319), .ZN(n316) );
  OR2_X1 U310 ( .A1(a_1_), .A2(n231), .ZN(n318) );
  OR2_X1 U311 ( .A1(n320), .A2(n321), .ZN(n231) );
  AND2_X1 U312 ( .A1(n183), .A2(a_2_), .ZN(n321) );
  AND2_X1 U313 ( .A1(n322), .A2(n191), .ZN(n320) );
  OR2_X1 U314 ( .A1(n183), .A2(a_2_), .ZN(n322) );
  AND2_X1 U315 ( .A1(n323), .A2(a_3_), .ZN(n183) );
  AND2_X1 U316 ( .A1(n324), .A2(a_0_), .ZN(n305) );
  AND2_X1 U317 ( .A1(n182), .A2(n325), .ZN(n299) );
  OR2_X1 U318 ( .A1(n326), .A2(n327), .ZN(n325) );
  OR2_X1 U319 ( .A1(n328), .A2(n329), .ZN(n327) );
  AND2_X1 U320 ( .A1(n298), .A2(n330), .ZN(n329) );
  INV_X1 U321 ( .A(n297), .ZN(n330) );
  OR2_X1 U322 ( .A1(n331), .A2(n328), .ZN(n297) );
  AND2_X1 U323 ( .A1(n332), .A2(n333), .ZN(n331) );
  AND2_X1 U324 ( .A1(n293), .A2(n294), .ZN(n298) );
  AND2_X1 U325 ( .A1(n290), .A2(n334), .ZN(n294) );
  INV_X1 U326 ( .A(n289), .ZN(n334) );
  OR2_X1 U327 ( .A1(n335), .A2(n336), .ZN(n289) );
  AND2_X1 U328 ( .A1(n285), .A2(n284), .ZN(n336) );
  AND2_X1 U329 ( .A1(n282), .A2(n337), .ZN(n335) );
  OR2_X1 U330 ( .A1(n284), .A2(n285), .ZN(n337) );
  OR2_X1 U331 ( .A1(n323), .A2(n315), .ZN(n285) );
  OR2_X1 U332 ( .A1(n338), .A2(n339), .ZN(n284) );
  AND2_X1 U333 ( .A1(n245), .A2(n248), .ZN(n339) );
  AND2_X1 U334 ( .A1(n340), .A2(n247), .ZN(n338) );
  OR2_X1 U335 ( .A1(n341), .A2(n342), .ZN(n247) );
  INV_X1 U336 ( .A(n343), .ZN(n342) );
  AND2_X1 U337 ( .A1(n344), .A2(n345), .ZN(n341) );
  OR2_X1 U338 ( .A1(n312), .A2(n319), .ZN(n345) );
  OR2_X1 U339 ( .A1(n198), .A2(n191), .ZN(n344) );
  OR2_X1 U340 ( .A1(n248), .A2(n245), .ZN(n340) );
  OR2_X1 U341 ( .A1(n323), .A2(n243), .ZN(n245) );
  INV_X1 U342 ( .A(b_3_), .ZN(n323) );
  OR2_X1 U343 ( .A1(n191), .A2(n346), .ZN(n248) );
  OR2_X1 U344 ( .A1(n213), .A2(n198), .ZN(n346) );
  INV_X1 U345 ( .A(n185), .ZN(n213) );
  AND2_X1 U346 ( .A1(a_3_), .A2(b_3_), .ZN(n185) );
  XNOR2_X1 U347 ( .A(n347), .B(n348), .ZN(n282) );
  XNOR2_X1 U348 ( .A(n349), .B(n343), .ZN(n347) );
  XOR2_X1 U349 ( .A(n350), .B(n351), .Z(n290) );
  XNOR2_X1 U350 ( .A(n352), .B(n353), .ZN(n350) );
  XOR2_X1 U351 ( .A(n354), .B(n355), .Z(n293) );
  INV_X1 U352 ( .A(n356), .ZN(n328) );
  OR2_X1 U353 ( .A1(n332), .A2(n333), .ZN(n356) );
  OR2_X1 U354 ( .A1(n354), .A2(n355), .ZN(n333) );
  XOR2_X1 U355 ( .A(n357), .B(n358), .Z(n355) );
  XOR2_X1 U356 ( .A(n359), .B(n360), .Z(n357) );
  OR2_X1 U357 ( .A1(n361), .A2(n362), .ZN(n354) );
  AND2_X1 U358 ( .A1(n352), .A2(n353), .ZN(n362) );
  AND2_X1 U359 ( .A1(n351), .A2(n363), .ZN(n361) );
  OR2_X1 U360 ( .A1(n353), .A2(n352), .ZN(n363) );
  OR2_X1 U361 ( .A1(n364), .A2(n365), .ZN(n352) );
  AND2_X1 U362 ( .A1(n348), .A2(n343), .ZN(n365) );
  AND2_X1 U363 ( .A1(n366), .A2(n349), .ZN(n364) );
  OR2_X1 U364 ( .A1(n367), .A2(n368), .ZN(n349) );
  INV_X1 U365 ( .A(n369), .ZN(n368) );
  AND2_X1 U366 ( .A1(n370), .A2(n371), .ZN(n367) );
  OR2_X1 U367 ( .A1(n312), .A2(n324), .ZN(n370) );
  OR2_X1 U368 ( .A1(n343), .A2(n348), .ZN(n366) );
  OR2_X1 U369 ( .A1(n191), .A2(n243), .ZN(n348) );
  OR2_X1 U370 ( .A1(n371), .A2(n372), .ZN(n343) );
  OR2_X1 U371 ( .A1(n312), .A2(n191), .ZN(n372) );
  OR2_X1 U372 ( .A1(n191), .A2(n315), .ZN(n353) );
  INV_X1 U373 ( .A(b_2_), .ZN(n191) );
  XNOR2_X1 U374 ( .A(n373), .B(n369), .ZN(n351) );
  OR2_X1 U375 ( .A1(n374), .A2(n375), .ZN(n373) );
  INV_X1 U376 ( .A(n376), .ZN(n375) );
  AND2_X1 U377 ( .A1(n377), .A2(n378), .ZN(n374) );
  OR2_X1 U378 ( .A1(n326), .A2(n379), .ZN(n332) );
  AND2_X1 U379 ( .A1(n380), .A2(n381), .ZN(n379) );
  OR2_X1 U380 ( .A1(n324), .A2(n315), .ZN(n380) );
  AND2_X1 U381 ( .A1(n382), .A2(a_0_), .ZN(n326) );
  INV_X1 U382 ( .A(n381), .ZN(n382) );
  OR2_X1 U383 ( .A1(n383), .A2(n384), .ZN(n381) );
  AND2_X1 U384 ( .A1(n358), .A2(n360), .ZN(n384) );
  AND2_X1 U385 ( .A1(n359), .A2(n385), .ZN(n383) );
  OR2_X1 U386 ( .A1(n360), .A2(n358), .ZN(n385) );
  OR2_X1 U387 ( .A1(n243), .A2(n324), .ZN(n358) );
  OR2_X1 U388 ( .A1(n319), .A2(n315), .ZN(n360) );
  INV_X1 U389 ( .A(a_0_), .ZN(n315) );
  AND2_X1 U390 ( .A1(n376), .A2(n369), .ZN(n359) );
  OR2_X1 U391 ( .A1(n324), .A2(n386), .ZN(n369) );
  OR2_X1 U392 ( .A1(n312), .A2(n371), .ZN(n386) );
  OR2_X1 U393 ( .A1(n198), .A2(n319), .ZN(n371) );
  INV_X1 U394 ( .A(a_3_), .ZN(n312) );
  OR2_X1 U395 ( .A1(n378), .A2(n377), .ZN(n376) );
  OR2_X1 U396 ( .A1(n243), .A2(n319), .ZN(n377) );
  INV_X1 U397 ( .A(b_1_), .ZN(n319) );
  INV_X1 U398 ( .A(a_1_), .ZN(n243) );
  OR2_X1 U399 ( .A1(n198), .A2(n324), .ZN(n378) );
  INV_X1 U400 ( .A(b_0_), .ZN(n324) );
  INV_X1 U401 ( .A(a_2_), .ZN(n198) );
  AND2_X1 U402 ( .A1(operation_0_), .A2(operation_1_), .ZN(n182) );
endmodule

