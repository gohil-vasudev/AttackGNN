module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n595_, new_n614_, new_n445_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n421_, new_n620_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n636_, new_n670_, new_n456_, new_n246_, new_n170_, new_n682_, new_n679_, new_n266_, new_n667_, new_n367_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n624_, new_n534_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n602_, new_n240_, new_n413_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n462_, new_n603_, new_n564_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n626_, new_n152_, new_n153_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n655_, new_n630_, new_n167_, new_n385_, new_n478_, new_n461_, new_n297_, new_n361_, new_n565_, new_n683_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n530_, new_n318_, new_n622_, new_n629_, new_n321_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n549_, new_n676_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n650_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n506_, new_n680_, new_n256_, new_n452_, new_n381_, new_n656_, new_n388_, new_n508_, new_n194_, new_n483_, new_n394_, new_n299_, new_n657_, new_n652_, new_n314_, new_n582_, new_n363_, new_n165_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n187_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n488_, new_n524_, new_n277_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n346_, new_n396_, new_n438_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n399_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n437_, new_n295_, new_n359_, new_n628_, new_n162_, new_n409_, new_n457_, new_n553_, new_n668_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n155_, new_n384_, new_n410_, new_n543_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n654_, new_n604_, new_n227_, new_n416_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n310_, new_n275_, new_n575_, new_n562_, new_n525_, new_n578_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n379_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n520_, new_n253_, new_n403_, new_n475_, new_n237_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n605_, new_n182_, new_n407_, new_n666_, new_n480_, new_n625_, new_n151_, new_n513_, new_n592_, new_n558_, new_n231_, new_n219_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n522_, new_n588_, new_n428_, new_n199_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n225_, new_n387_, new_n544_, new_n476_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n499_, new_n533_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n285_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n662_, new_n440_, new_n531_, new_n252_, new_n585_, new_n160_, new_n312_, new_n535_, new_n372_, new_n242_, new_n503_, new_n527_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n651_, new_n433_, new_n435_, new_n265_, new_n370_, new_n584_, new_n278_, new_n304_, new_n523_, new_n638_, new_n550_, new_n217_, new_n269_, new_n512_, new_n644_, new_n599_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n594_, new_n561_, new_n495_, new_n431_, new_n196_, new_n319_, new_n640_, new_n684_, new_n338_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n627_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n358_, new_n348_, new_n610_, new_n322_, new_n545_, new_n611_, new_n289_, new_n425_, new_n226_, new_n185_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n551_, new_n168_, new_n279_, new_n455_, new_n618_, new_n521_, new_n406_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n573_, new_n405_;

not g000 ( new_n151_, N42 );
nand g001 ( new_n152_, N29, N75 );
nor g002 ( new_n153_, new_n152_, new_n151_ );
xnor g003 ( N388, new_n153_, keyIn_0_3 );
not g004 ( new_n155_, N80 );
nand g005 ( new_n156_, N29, N36 );
nor g006 ( N389, new_n156_, new_n155_ );
nor g007 ( new_n158_, new_n156_, new_n151_ );
xor g008 ( N390, new_n158_, keyIn_0_4 );
nand g009 ( new_n160_, N85, N86 );
not g010 ( N391, new_n160_ );
not g011 ( new_n162_, N13 );
nand g012 ( new_n163_, N1, N8 );
nor g013 ( new_n164_, new_n163_, new_n162_ );
nand g014 ( new_n165_, new_n164_, N17 );
xnor g015 ( N418, new_n165_, keyIn_0_0 );
xnor g016 ( new_n167_, new_n158_, keyIn_0_1 );
not g017 ( new_n168_, new_n167_ );
nand g018 ( new_n169_, N1, N26 );
nand g019 ( new_n170_, N13, N17 );
nor g020 ( new_n171_, new_n169_, new_n170_ );
nand g021 ( N419, new_n168_, new_n171_ );
nand g022 ( new_n173_, N59, N75 );
not g023 ( new_n174_, new_n173_ );
nand g024 ( N420, new_n174_, N80 );
nand g025 ( new_n176_, N36, N59 );
not g026 ( new_n177_, new_n176_ );
nand g027 ( N421, new_n177_, N80 );
nor g028 ( new_n179_, new_n176_, new_n151_ );
xnor g029 ( N422, new_n179_, keyIn_0_5 );
not g030 ( new_n181_, N90 );
nor g031 ( new_n182_, N87, N88 );
nor g032 ( N423, new_n182_, new_n181_ );
nand g033 ( N446, new_n167_, new_n171_ );
not g034 ( new_n185_, keyIn_0_2 );
not g035 ( new_n186_, N51 );
nor g036 ( new_n187_, new_n169_, new_n186_ );
xnor g037 ( N447, new_n187_, new_n185_ );
nand g038 ( new_n189_, new_n164_, N55 );
nand g039 ( new_n190_, N29, N68 );
nor g040 ( N448, new_n189_, new_n190_ );
nand g041 ( new_n192_, N59, N68 );
nor g042 ( new_n193_, new_n189_, new_n192_ );
nand g043 ( new_n194_, new_n193_, N74 );
xor g044 ( N449, new_n194_, keyIn_0_12 );
not g045 ( new_n196_, N89 );
nor g046 ( new_n197_, new_n182_, new_n196_ );
xnor g047 ( N450, new_n197_, keyIn_0_9 );
nor g048 ( new_n199_, N111, N116 );
nor g049 ( new_n200_, new_n199_, keyIn_0_6 );
not g050 ( new_n201_, N111 );
nand g051 ( new_n202_, new_n201_, keyIn_0_6 );
nor g052 ( new_n203_, new_n202_, N116 );
nor g053 ( new_n204_, new_n203_, new_n200_ );
nand g054 ( new_n205_, N111, N116 );
not g055 ( new_n206_, new_n205_ );
nor g056 ( new_n207_, new_n204_, new_n206_ );
xnor g057 ( new_n208_, N121, N126 );
xnor g058 ( new_n209_, new_n207_, new_n208_ );
nor g059 ( new_n210_, new_n209_, N135 );
not g060 ( new_n211_, new_n210_ );
nor g061 ( new_n212_, new_n211_, keyIn_0_19 );
nand g062 ( new_n213_, new_n211_, keyIn_0_19 );
nand g063 ( new_n214_, new_n209_, N135 );
nand g064 ( new_n215_, new_n213_, new_n214_ );
nor g065 ( new_n216_, new_n215_, new_n212_ );
xnor g066 ( new_n217_, N91, N96 );
xnor g067 ( new_n218_, N101, N106 );
xnor g068 ( new_n219_, new_n217_, new_n218_ );
xnor g069 ( new_n220_, new_n219_, N130 );
nand g070 ( new_n221_, new_n216_, new_n220_ );
nor g071 ( new_n222_, new_n221_, keyIn_0_32 );
nand g072 ( new_n223_, new_n221_, keyIn_0_32 );
not g073 ( new_n224_, new_n216_ );
not g074 ( new_n225_, new_n220_ );
nand g075 ( new_n226_, new_n224_, new_n225_ );
nand g076 ( new_n227_, new_n223_, new_n226_ );
nor g077 ( N767, new_n227_, new_n222_ );
not g078 ( new_n229_, keyIn_0_25 );
xnor g079 ( new_n230_, N171, N177 );
nor g080 ( new_n231_, N159, N165 );
not g081 ( new_n232_, keyIn_0_13 );
nand g082 ( new_n233_, N159, N165 );
nand g083 ( new_n234_, new_n233_, new_n232_ );
nor g084 ( new_n235_, new_n234_, new_n231_ );
xnor g085 ( new_n236_, new_n235_, new_n230_ );
nor g086 ( new_n237_, new_n236_, N130 );
nand g087 ( new_n238_, new_n237_, new_n229_ );
nor g088 ( new_n239_, new_n237_, new_n229_ );
nand g089 ( new_n240_, new_n236_, N130 );
nand g090 ( new_n241_, new_n240_, keyIn_0_31 );
nor g091 ( new_n242_, new_n239_, new_n241_ );
nand g092 ( new_n243_, new_n242_, new_n238_ );
not g093 ( new_n244_, N207 );
xnor g094 ( new_n245_, N183, N189 );
xnor g095 ( new_n246_, N195, N201 );
xnor g096 ( new_n247_, new_n245_, new_n246_ );
nand g097 ( new_n248_, new_n247_, new_n244_ );
nor g098 ( new_n249_, new_n248_, keyIn_0_26 );
not g099 ( new_n250_, new_n247_ );
nand g100 ( new_n251_, new_n250_, N207 );
nand g101 ( new_n252_, new_n248_, keyIn_0_26 );
nand g102 ( new_n253_, new_n252_, new_n251_ );
nor g103 ( new_n254_, new_n253_, new_n249_ );
xnor g104 ( N768, new_n243_, new_n254_ );
nor g105 ( new_n256_, new_n152_, new_n155_ );
not g106 ( new_n257_, new_n256_ );
nand g107 ( new_n258_, N447, N55 );
nor g108 ( new_n259_, new_n258_, new_n257_ );
not g109 ( new_n260_, new_n259_ );
nor g110 ( new_n261_, new_n260_, keyIn_0_15 );
not g111 ( new_n262_, new_n261_ );
not g112 ( new_n263_, keyIn_0_15 );
nor g113 ( new_n264_, new_n259_, new_n263_ );
xor g114 ( new_n265_, keyIn_0_10, N268 );
not g115 ( new_n266_, new_n265_ );
nor g116 ( new_n267_, new_n264_, new_n266_ );
nand g117 ( new_n268_, new_n262_, new_n267_ );
not g118 ( new_n269_, keyIn_0_24 );
nor g119 ( new_n270_, N17, N42 );
nand g120 ( new_n271_, N59, N156 );
not g121 ( new_n272_, new_n271_ );
nand g122 ( new_n273_, N17, N42 );
nand g123 ( new_n274_, new_n272_, new_n273_ );
nor g124 ( new_n275_, new_n274_, new_n270_ );
nand g125 ( new_n276_, N447, new_n275_ );
nand g126 ( new_n277_, N42, N59 );
not g127 ( new_n278_, new_n277_ );
nand g128 ( new_n279_, new_n278_, N75 );
nand g129 ( new_n280_, N17, N51 );
nor g130 ( new_n281_, new_n163_, new_n280_ );
nand g131 ( new_n282_, new_n279_, new_n281_ );
nand g132 ( new_n283_, new_n276_, new_n282_ );
nand g133 ( new_n284_, new_n283_, N126 );
nor g134 ( new_n285_, new_n284_, new_n269_ );
not g135 ( new_n286_, N17 );
not g136 ( new_n287_, new_n169_ );
nand g137 ( new_n288_, new_n287_, N51 );
nand g138 ( new_n289_, new_n288_, new_n185_ );
nand g139 ( new_n290_, new_n187_, keyIn_0_2 );
nand g140 ( new_n291_, new_n289_, new_n290_ );
nor g141 ( new_n292_, new_n291_, new_n286_ );
nand g142 ( new_n293_, new_n292_, new_n271_ );
nand g143 ( new_n294_, new_n293_, N1 );
nand g144 ( new_n295_, new_n294_, N153 );
nand g145 ( new_n296_, new_n284_, new_n269_ );
nand g146 ( new_n297_, new_n295_, new_n296_ );
nor g147 ( new_n298_, new_n297_, new_n285_ );
nand g148 ( new_n299_, new_n298_, new_n268_ );
nand g149 ( new_n300_, new_n299_, N201 );
xnor g150 ( new_n301_, new_n300_, keyIn_0_37 );
not g151 ( new_n302_, N201 );
not g152 ( new_n303_, new_n267_ );
nor g153 ( new_n304_, new_n303_, new_n261_ );
not g154 ( new_n305_, new_n285_ );
not g155 ( new_n306_, new_n297_ );
nand g156 ( new_n307_, new_n306_, new_n305_ );
nor g157 ( new_n308_, new_n307_, new_n304_ );
nand g158 ( new_n309_, new_n308_, new_n302_ );
nand g159 ( new_n310_, new_n309_, keyIn_0_38 );
not g160 ( new_n311_, new_n310_ );
nor g161 ( new_n312_, new_n309_, keyIn_0_38 );
nor g162 ( new_n313_, new_n311_, new_n312_ );
nand g163 ( new_n314_, new_n313_, new_n301_ );
xor g164 ( new_n315_, new_n314_, N261 );
nor g165 ( new_n316_, new_n315_, keyIn_0_52 );
nand g166 ( new_n317_, new_n315_, keyIn_0_52 );
nand g167 ( new_n318_, new_n317_, N219 );
nor g168 ( new_n319_, new_n318_, new_n316_ );
nand g169 ( new_n320_, N121, N210 );
not g170 ( new_n321_, new_n320_ );
nor g171 ( new_n322_, new_n319_, new_n321_ );
xor g172 ( new_n323_, new_n322_, keyIn_0_56 );
not g173 ( new_n324_, keyIn_0_8 );
nand g174 ( new_n325_, N42, N72 );
not g175 ( new_n326_, new_n325_ );
nand g176 ( new_n327_, new_n193_, new_n326_ );
nor g177 ( new_n328_, new_n327_, new_n324_ );
nand g178 ( new_n329_, new_n327_, new_n324_ );
nand g179 ( new_n330_, new_n329_, N73 );
nor g180 ( new_n331_, new_n330_, new_n328_ );
xnor g181 ( new_n332_, new_n331_, keyIn_0_11 );
xnor g182 ( new_n333_, new_n332_, keyIn_0_14 );
xnor g183 ( new_n334_, new_n333_, keyIn_0_16 );
nor g184 ( new_n335_, new_n334_, new_n302_ );
xnor g185 ( new_n336_, new_n335_, keyIn_0_28 );
not g186 ( new_n337_, keyIn_0_50 );
not g187 ( new_n338_, N237 );
nor g188 ( new_n339_, new_n301_, new_n338_ );
nor g189 ( new_n340_, new_n339_, new_n337_ );
nand g190 ( new_n341_, new_n299_, N246 );
nand g191 ( new_n342_, N255, N267 );
nand g192 ( new_n343_, new_n341_, new_n342_ );
nor g193 ( new_n344_, new_n340_, new_n343_ );
not g194 ( new_n345_, N228 );
nor g195 ( new_n346_, new_n314_, new_n345_ );
not g196 ( new_n347_, new_n339_ );
nor g197 ( new_n348_, new_n347_, keyIn_0_50 );
nor g198 ( new_n349_, new_n346_, new_n348_ );
nand g199 ( new_n350_, new_n349_, new_n344_ );
nor g200 ( new_n351_, new_n350_, new_n336_ );
nand g201 ( N850, new_n323_, new_n351_ );
not g202 ( new_n353_, keyIn_0_53 );
not g203 ( new_n354_, keyIn_0_29 );
nand g204 ( new_n355_, new_n283_, N111 );
nor g205 ( new_n356_, new_n355_, keyIn_0_22 );
nand g206 ( new_n357_, new_n294_, N143 );
nand g207 ( new_n358_, new_n355_, keyIn_0_22 );
nand g208 ( new_n359_, new_n357_, new_n358_ );
nor g209 ( new_n360_, new_n359_, new_n356_ );
nand g210 ( new_n361_, new_n360_, new_n268_ );
xnor g211 ( new_n362_, new_n361_, new_n354_ );
nand g212 ( new_n363_, new_n362_, N183 );
xnor g213 ( new_n364_, new_n363_, keyIn_0_36 );
nor g214 ( new_n365_, new_n362_, N183 );
nor g215 ( new_n366_, new_n364_, new_n365_ );
not g216 ( new_n367_, keyIn_0_30 );
not g217 ( new_n368_, keyIn_0_23 );
nand g218 ( new_n369_, new_n283_, N116 );
nor g219 ( new_n370_, new_n369_, new_n368_ );
nand g220 ( new_n371_, new_n294_, N146 );
nand g221 ( new_n372_, new_n369_, new_n368_ );
nand g222 ( new_n373_, new_n371_, new_n372_ );
nor g223 ( new_n374_, new_n373_, new_n370_ );
nand g224 ( new_n375_, new_n374_, new_n268_ );
xnor g225 ( new_n376_, new_n375_, new_n367_ );
nor g226 ( new_n377_, new_n376_, N189 );
not g227 ( new_n378_, new_n377_ );
nand g228 ( new_n379_, new_n294_, N149 );
nand g229 ( new_n380_, new_n283_, N121 );
nand g230 ( new_n381_, new_n379_, new_n380_ );
nor g231 ( new_n382_, new_n304_, new_n381_ );
not g232 ( new_n383_, new_n382_ );
nor g233 ( new_n384_, new_n383_, N195 );
nor g234 ( new_n385_, new_n301_, new_n384_ );
nand g235 ( new_n386_, new_n385_, new_n378_ );
xor g236 ( new_n387_, new_n386_, keyIn_0_51 );
nand g237 ( new_n388_, new_n310_, N261 );
nor g238 ( new_n389_, new_n388_, new_n312_ );
nor g239 ( new_n390_, new_n377_, new_n384_ );
nand g240 ( new_n391_, new_n390_, new_n389_ );
nor g241 ( new_n392_, new_n391_, keyIn_0_42 );
nand g242 ( new_n393_, new_n391_, keyIn_0_42 );
not g243 ( new_n394_, N195 );
nor g244 ( new_n395_, new_n382_, new_n394_ );
not g245 ( new_n396_, new_n395_ );
nor g246 ( new_n397_, new_n377_, new_n396_ );
not g247 ( new_n398_, N189 );
not g248 ( new_n399_, new_n376_ );
nor g249 ( new_n400_, new_n399_, new_n398_ );
nor g250 ( new_n401_, new_n397_, new_n400_ );
nand g251 ( new_n402_, new_n393_, new_n401_ );
nor g252 ( new_n403_, new_n402_, new_n392_ );
nand g253 ( new_n404_, new_n403_, new_n387_ );
nand g254 ( new_n405_, new_n404_, new_n366_ );
nor g255 ( new_n406_, new_n405_, new_n353_ );
not g256 ( new_n407_, new_n366_ );
not g257 ( new_n408_, new_n404_ );
nand g258 ( new_n409_, new_n408_, new_n407_ );
nand g259 ( new_n410_, new_n405_, new_n353_ );
nand g260 ( new_n411_, new_n410_, new_n409_ );
nor g261 ( new_n412_, new_n411_, new_n406_ );
nand g262 ( new_n413_, new_n412_, keyIn_0_55 );
not g263 ( new_n414_, N219 );
nor g264 ( new_n415_, new_n412_, keyIn_0_55 );
nor g265 ( new_n416_, new_n415_, new_n414_ );
nand g266 ( new_n417_, new_n416_, new_n413_ );
not g267 ( new_n418_, keyIn_0_47 );
nor g268 ( new_n419_, new_n407_, new_n345_ );
not g269 ( new_n420_, new_n419_ );
nand g270 ( new_n421_, new_n420_, new_n418_ );
not g271 ( new_n422_, keyIn_0_27 );
not g272 ( new_n423_, new_n334_ );
nand g273 ( new_n424_, new_n423_, N183 );
nor g274 ( new_n425_, new_n424_, new_n422_ );
nand g275 ( new_n426_, new_n424_, new_n422_ );
not g276 ( new_n427_, N246 );
not g277 ( new_n428_, new_n362_ );
nor g278 ( new_n429_, new_n428_, new_n427_ );
nand g279 ( new_n430_, N106, N210 );
not g280 ( new_n431_, new_n430_ );
nor g281 ( new_n432_, new_n429_, new_n431_ );
nand g282 ( new_n433_, new_n426_, new_n432_ );
nor g283 ( new_n434_, new_n433_, new_n425_ );
nand g284 ( new_n435_, new_n421_, new_n434_ );
nand g285 ( new_n436_, new_n419_, keyIn_0_47 );
xnor g286 ( new_n437_, new_n364_, keyIn_0_40 );
nand g287 ( new_n438_, new_n437_, N237 );
nand g288 ( new_n439_, new_n436_, new_n438_ );
nor g289 ( new_n440_, new_n435_, new_n439_ );
nand g290 ( N863, new_n417_, new_n440_ );
nor g291 ( new_n442_, new_n400_, new_n377_ );
not g292 ( new_n443_, new_n301_ );
nor g293 ( new_n444_, new_n389_, new_n443_ );
nor g294 ( new_n445_, new_n444_, new_n384_ );
not g295 ( new_n446_, new_n445_ );
xor g296 ( new_n447_, new_n395_, keyIn_0_49 );
nand g297 ( new_n448_, new_n446_, new_n447_ );
nand g298 ( new_n449_, new_n448_, new_n442_ );
nor g299 ( new_n450_, new_n448_, new_n442_ );
nor g300 ( new_n451_, new_n450_, new_n414_ );
nand g301 ( new_n452_, new_n451_, new_n449_ );
nor g302 ( new_n453_, new_n334_, new_n398_ );
nand g303 ( new_n454_, new_n400_, N237 );
nand g304 ( new_n455_, N111, N210 );
nand g305 ( new_n456_, new_n454_, new_n455_ );
nor g306 ( new_n457_, new_n456_, new_n453_ );
nand g307 ( new_n458_, new_n376_, N246 );
nand g308 ( new_n459_, N255, N259 );
nand g309 ( new_n460_, new_n458_, new_n459_ );
xnor g310 ( new_n461_, new_n460_, keyIn_0_41 );
nand g311 ( new_n462_, new_n457_, new_n461_ );
nand g312 ( new_n463_, new_n442_, N228 );
xor g313 ( new_n464_, new_n463_, keyIn_0_48 );
nor g314 ( new_n465_, new_n464_, new_n462_ );
nand g315 ( N864, new_n452_, new_n465_ );
nand g316 ( new_n467_, new_n445_, new_n396_ );
not g317 ( new_n468_, new_n444_ );
nor g318 ( new_n469_, new_n384_, new_n395_ );
nor g319 ( new_n470_, new_n468_, new_n469_ );
nor g320 ( new_n471_, new_n470_, new_n414_ );
nand g321 ( new_n472_, new_n471_, new_n467_ );
nor g322 ( new_n473_, new_n334_, new_n394_ );
nand g323 ( new_n474_, new_n469_, N228 );
nor g324 ( new_n475_, new_n396_, new_n338_ );
nand g325 ( new_n476_, new_n383_, N246 );
nand g326 ( new_n477_, N255, N260 );
nand g327 ( new_n478_, N116, N210 );
nand g328 ( new_n479_, new_n477_, new_n478_ );
not g329 ( new_n480_, new_n479_ );
nand g330 ( new_n481_, new_n476_, new_n480_ );
nor g331 ( new_n482_, new_n475_, new_n481_ );
nand g332 ( new_n483_, new_n482_, new_n474_ );
nor g333 ( new_n484_, new_n483_, new_n473_ );
nand g334 ( N865, new_n472_, new_n484_ );
not g335 ( new_n486_, N177 );
not g336 ( new_n487_, keyIn_0_18 );
nor g337 ( new_n488_, new_n257_, N268 );
nand g338 ( new_n489_, new_n292_, new_n488_ );
not g339 ( new_n490_, new_n489_ );
nor g340 ( new_n491_, new_n490_, new_n487_ );
nand g341 ( new_n492_, N138, N152 );
not g342 ( new_n493_, new_n492_ );
nor g343 ( new_n494_, new_n491_, new_n493_ );
not g344 ( new_n495_, new_n494_ );
nand g345 ( new_n496_, new_n283_, N106 );
nor g346 ( new_n497_, new_n258_, new_n272_ );
nand g347 ( new_n498_, new_n497_, N153 );
not g348 ( new_n499_, new_n498_ );
nor g349 ( new_n500_, new_n489_, keyIn_0_18 );
nor g350 ( new_n501_, new_n499_, new_n500_ );
nand g351 ( new_n502_, new_n501_, new_n496_ );
nor g352 ( new_n503_, new_n502_, new_n495_ );
nor g353 ( new_n504_, new_n503_, new_n486_ );
not g354 ( new_n505_, new_n504_ );
not g355 ( new_n506_, new_n503_ );
nor g356 ( new_n507_, new_n506_, N177 );
not g357 ( new_n508_, new_n507_ );
not g358 ( new_n509_, keyIn_0_46 );
nand g359 ( new_n510_, new_n437_, new_n509_ );
not g360 ( new_n511_, keyIn_0_40 );
xnor g361 ( new_n512_, new_n364_, new_n511_ );
nand g362 ( new_n513_, new_n512_, keyIn_0_46 );
nand g363 ( new_n514_, new_n510_, new_n513_ );
not g364 ( new_n515_, new_n365_ );
nand g365 ( new_n516_, new_n404_, new_n515_ );
nand g366 ( new_n517_, new_n516_, new_n514_ );
xnor g367 ( new_n518_, new_n517_, keyIn_0_54 );
nand g368 ( new_n519_, new_n518_, new_n508_ );
nand g369 ( new_n520_, new_n519_, new_n505_ );
nand g370 ( new_n521_, new_n497_, N149 );
nor g371 ( new_n522_, new_n521_, keyIn_0_17 );
nand g372 ( new_n523_, new_n521_, keyIn_0_17 );
nand g373 ( new_n524_, new_n283_, N101 );
not g374 ( new_n525_, new_n524_ );
nand g375 ( new_n526_, N17, N138 );
nand g376 ( new_n527_, new_n489_, new_n526_ );
nor g377 ( new_n528_, new_n525_, new_n527_ );
nand g378 ( new_n529_, new_n528_, new_n523_ );
nor g379 ( new_n530_, new_n529_, new_n522_ );
not g380 ( new_n531_, new_n530_ );
nor g381 ( new_n532_, new_n531_, N171 );
not g382 ( new_n533_, new_n532_ );
nand g383 ( new_n534_, new_n520_, new_n533_ );
nand g384 ( new_n535_, new_n531_, N171 );
xnor g385 ( new_n536_, new_n535_, keyIn_0_35 );
nand g386 ( new_n537_, new_n534_, new_n536_ );
not g387 ( new_n538_, N165 );
nand g388 ( new_n539_, new_n497_, N146 );
nand g389 ( new_n540_, new_n539_, new_n489_ );
not g390 ( new_n541_, new_n540_ );
nor g391 ( new_n542_, new_n541_, keyIn_0_21 );
nand g392 ( new_n543_, new_n541_, keyIn_0_21 );
not g393 ( new_n544_, new_n543_ );
nand g394 ( new_n545_, new_n283_, N96 );
nand g395 ( new_n546_, N51, N138 );
nand g396 ( new_n547_, new_n545_, new_n546_ );
nor g397 ( new_n548_, new_n544_, new_n547_ );
not g398 ( new_n549_, new_n548_ );
nor g399 ( new_n550_, new_n549_, new_n542_ );
nand g400 ( new_n551_, new_n550_, new_n538_ );
nand g401 ( new_n552_, new_n537_, new_n551_ );
not g402 ( new_n553_, new_n550_ );
nand g403 ( new_n554_, new_n553_, N165 );
nand g404 ( new_n555_, new_n552_, new_n554_ );
not g405 ( new_n556_, N159 );
nand g406 ( new_n557_, new_n497_, N143 );
nand g407 ( new_n558_, new_n557_, new_n489_ );
nor g408 ( new_n559_, new_n558_, keyIn_0_20 );
nand g409 ( new_n560_, new_n558_, keyIn_0_20 );
nand g410 ( new_n561_, new_n283_, N91 );
nand g411 ( new_n562_, N8, N138 );
nand g412 ( new_n563_, new_n561_, new_n562_ );
not g413 ( new_n564_, new_n563_ );
nand g414 ( new_n565_, new_n560_, new_n564_ );
nor g415 ( new_n566_, new_n565_, new_n559_ );
nand g416 ( new_n567_, new_n566_, new_n556_ );
xor g417 ( new_n568_, new_n567_, keyIn_0_33 );
not g418 ( new_n569_, new_n568_ );
nand g419 ( new_n570_, new_n555_, new_n569_ );
nor g420 ( new_n571_, new_n566_, new_n556_ );
xor g421 ( new_n572_, new_n571_, keyIn_0_43 );
nand g422 ( new_n573_, new_n570_, new_n572_ );
xnor g423 ( N866, new_n573_, keyIn_0_59 );
nor g424 ( new_n575_, new_n507_, new_n504_ );
nor g425 ( new_n576_, new_n518_, new_n575_ );
nand g426 ( new_n577_, new_n576_, keyIn_0_57 );
nor g427 ( new_n578_, new_n576_, keyIn_0_57 );
nand g428 ( new_n579_, new_n518_, new_n575_ );
nand g429 ( new_n580_, new_n579_, N219 );
nor g430 ( new_n581_, new_n578_, new_n580_ );
nand g431 ( new_n582_, new_n581_, new_n577_ );
nor g432 ( new_n583_, new_n334_, new_n486_ );
nand g433 ( new_n584_, new_n575_, N228 );
nor g434 ( new_n585_, new_n505_, new_n338_ );
nand g435 ( new_n586_, new_n506_, N246 );
nand g436 ( new_n587_, N101, N210 );
nand g437 ( new_n588_, new_n586_, new_n587_ );
nor g438 ( new_n589_, new_n585_, new_n588_ );
nand g439 ( new_n590_, new_n589_, new_n584_ );
nor g440 ( new_n591_, new_n590_, new_n583_ );
nand g441 ( new_n592_, new_n582_, new_n591_ );
xor g442 ( N874, new_n592_, keyIn_0_62 );
not g443 ( new_n594_, new_n570_ );
not g444 ( new_n595_, new_n571_ );
nand g445 ( new_n596_, new_n594_, new_n595_ );
nor g446 ( new_n597_, new_n568_, new_n571_ );
nor g447 ( new_n598_, new_n555_, new_n597_ );
nor g448 ( new_n599_, new_n598_, new_n414_ );
nand g449 ( new_n600_, new_n596_, new_n599_ );
nand g450 ( new_n601_, new_n423_, N159 );
nor g451 ( new_n602_, new_n566_, new_n427_ );
xnor g452 ( new_n603_, new_n602_, keyIn_0_34 );
nand g453 ( new_n604_, new_n601_, new_n603_ );
nor g454 ( new_n605_, new_n604_, keyIn_0_39 );
nand g455 ( new_n606_, new_n604_, keyIn_0_39 );
not g456 ( new_n607_, new_n597_ );
nor g457 ( new_n608_, new_n607_, new_n345_ );
nand g458 ( new_n609_, new_n266_, N210 );
nand g459 ( new_n610_, new_n571_, N237 );
nand g460 ( new_n611_, new_n610_, new_n609_ );
nor g461 ( new_n612_, new_n608_, new_n611_ );
nand g462 ( new_n613_, new_n612_, new_n606_ );
nor g463 ( new_n614_, new_n613_, new_n605_ );
nand g464 ( N878, new_n600_, new_n614_ );
not g465 ( new_n616_, keyIn_0_60 );
nand g466 ( new_n617_, new_n554_, new_n551_ );
nor g467 ( new_n618_, new_n519_, new_n532_ );
not g468 ( new_n619_, keyIn_0_44 );
nor g469 ( new_n620_, new_n536_, new_n619_ );
not g470 ( new_n621_, new_n536_ );
nor g471 ( new_n622_, new_n621_, keyIn_0_44 );
nor g472 ( new_n623_, new_n505_, new_n532_ );
nor g473 ( new_n624_, new_n622_, new_n623_ );
not g474 ( new_n625_, new_n624_ );
nor g475 ( new_n626_, new_n625_, new_n620_ );
not g476 ( new_n627_, new_n626_ );
nor g477 ( new_n628_, new_n618_, new_n627_ );
nand g478 ( new_n629_, new_n628_, new_n617_ );
nand g479 ( new_n630_, new_n629_, keyIn_0_58 );
not g480 ( new_n631_, keyIn_0_58 );
not g481 ( new_n632_, new_n617_ );
not g482 ( new_n633_, keyIn_0_54 );
xnor g483 ( new_n634_, new_n517_, new_n633_ );
nor g484 ( new_n635_, new_n634_, new_n507_ );
nand g485 ( new_n636_, new_n635_, new_n533_ );
nand g486 ( new_n637_, new_n636_, new_n626_ );
nor g487 ( new_n638_, new_n637_, new_n632_ );
nand g488 ( new_n639_, new_n638_, new_n631_ );
nand g489 ( new_n640_, new_n630_, new_n639_ );
nor g490 ( new_n641_, new_n628_, new_n617_ );
nor g491 ( new_n642_, new_n641_, new_n414_ );
nand g492 ( new_n643_, new_n640_, new_n642_ );
not g493 ( new_n644_, keyIn_0_7 );
nand g494 ( new_n645_, N91, N210 );
nand g495 ( new_n646_, new_n645_, new_n644_ );
nand g496 ( new_n647_, keyIn_0_7, N91 );
not g497 ( new_n648_, new_n647_ );
nand g498 ( new_n649_, new_n648_, N210 );
nand g499 ( new_n650_, new_n649_, new_n646_ );
nand g500 ( new_n651_, new_n643_, new_n650_ );
xnor g501 ( new_n652_, new_n651_, new_n616_ );
nor g502 ( new_n653_, new_n334_, new_n538_ );
nand g503 ( new_n654_, new_n632_, N228 );
nor g504 ( new_n655_, new_n554_, new_n338_ );
nor g505 ( new_n656_, new_n550_, new_n427_ );
nor g506 ( new_n657_, new_n655_, new_n656_ );
nand g507 ( new_n658_, new_n654_, new_n657_ );
nor g508 ( new_n659_, new_n658_, new_n653_ );
nand g509 ( N879, new_n652_, new_n659_ );
not g510 ( new_n661_, keyIn_0_61 );
nor g511 ( new_n662_, new_n621_, new_n532_ );
nand g512 ( new_n663_, new_n520_, new_n662_ );
nor g513 ( new_n664_, new_n520_, new_n662_ );
nor g514 ( new_n665_, new_n664_, new_n414_ );
nand g515 ( new_n666_, new_n665_, new_n663_ );
nand g516 ( new_n667_, N96, N210 );
nand g517 ( new_n668_, new_n666_, new_n667_ );
xnor g518 ( new_n669_, new_n668_, new_n661_ );
nor g519 ( new_n670_, new_n536_, new_n338_ );
xnor g520 ( new_n671_, new_n670_, keyIn_0_45 );
nand g521 ( new_n672_, new_n662_, N228 );
nand g522 ( new_n673_, new_n423_, N171 );
not g523 ( new_n674_, new_n673_ );
nor g524 ( new_n675_, new_n530_, new_n427_ );
nor g525 ( new_n676_, new_n674_, new_n675_ );
nand g526 ( new_n677_, new_n676_, new_n672_ );
nor g527 ( new_n678_, new_n677_, new_n671_ );
nand g528 ( new_n679_, new_n669_, new_n678_ );
nand g529 ( new_n680_, new_n679_, keyIn_0_63 );
not g530 ( new_n681_, keyIn_0_63 );
xnor g531 ( new_n682_, new_n668_, keyIn_0_61 );
not g532 ( new_n683_, new_n678_ );
nor g533 ( new_n684_, new_n682_, new_n683_ );
nand g534 ( new_n685_, new_n684_, new_n681_ );
nand g535 ( N880, new_n685_, new_n680_ );
endmodule