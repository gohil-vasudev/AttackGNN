module add_mul_combine_8_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, Result_mul_0_, 
        Result_mul_1_, Result_mul_2_, Result_mul_3_, Result_mul_4_, 
        Result_mul_5_, Result_mul_6_, Result_mul_7_, Result_mul_8_, 
        Result_mul_9_, Result_mul_10_, Result_mul_11_, Result_mul_12_, 
        Result_mul_13_, Result_mul_14_, Result_mul_15_, Result_add_0_, 
        Result_add_1_, Result_add_2_, Result_add_3_, Result_add_4_, 
        Result_add_5_, Result_add_6_, Result_add_7_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_,
         b_4_, b_5_, b_6_, b_7_;
  output Result_mul_0_, Result_mul_1_, Result_mul_2_, Result_mul_3_,
         Result_mul_4_, Result_mul_5_, Result_mul_6_, Result_mul_7_,
         Result_mul_8_, Result_mul_9_, Result_mul_10_, Result_mul_11_,
         Result_mul_12_, Result_mul_13_, Result_mul_14_, Result_mul_15_,
         Result_add_0_, Result_add_1_, Result_add_2_, Result_add_3_,
         Result_add_4_, Result_add_5_, Result_add_6_, Result_add_7_;
  wire   n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874;

  XNOR2_X1 U448 ( .A(n424), .B(n425), .ZN(Result_mul_9_) );
  XOR2_X1 U449 ( .A(n426), .B(n427), .Z(n425) );
  XNOR2_X1 U450 ( .A(n428), .B(n429), .ZN(Result_mul_8_) );
  XOR2_X1 U451 ( .A(n430), .B(n431), .Z(n429) );
  XOR2_X1 U452 ( .A(n432), .B(n433), .Z(Result_mul_7_) );
  AND2_X1 U453 ( .A1(n434), .A2(n435), .ZN(Result_mul_6_) );
  OR2_X1 U454 ( .A1(n436), .A2(n437), .ZN(n434) );
  XOR2_X1 U455 ( .A(n438), .B(n439), .Z(n437) );
  INV_X1 U456 ( .A(n440), .ZN(n436) );
  XOR2_X1 U457 ( .A(n441), .B(n442), .Z(Result_mul_5_) );
  AND2_X1 U458 ( .A1(n435), .A2(n443), .ZN(n442) );
  XNOR2_X1 U459 ( .A(n444), .B(n445), .ZN(Result_mul_4_) );
  AND2_X1 U460 ( .A1(n446), .A2(n447), .ZN(n444) );
  XOR2_X1 U461 ( .A(n448), .B(n449), .Z(Result_mul_3_) );
  AND2_X1 U462 ( .A1(n450), .A2(n451), .ZN(n449) );
  OR2_X1 U463 ( .A1(n452), .A2(n453), .ZN(n451) );
  INV_X1 U464 ( .A(n454), .ZN(n450) );
  XOR2_X1 U465 ( .A(n455), .B(n456), .Z(Result_mul_2_) );
  XOR2_X1 U466 ( .A(n457), .B(n458), .Z(Result_mul_1_) );
  AND2_X1 U467 ( .A1(n459), .A2(n460), .ZN(n458) );
  OR2_X1 U468 ( .A1(n461), .A2(n462), .ZN(n460) );
  AND2_X1 U469 ( .A1(n463), .A2(n464), .ZN(n461) );
  INV_X1 U470 ( .A(n465), .ZN(n459) );
  XNOR2_X1 U471 ( .A(n466), .B(n467), .ZN(Result_mul_14_) );
  AND2_X1 U472 ( .A1(b_7_), .A2(a_6_), .ZN(n467) );
  XOR2_X1 U473 ( .A(n468), .B(n469), .Z(Result_mul_13_) );
  XNOR2_X1 U474 ( .A(n470), .B(n471), .ZN(n469) );
  XNOR2_X1 U475 ( .A(n472), .B(n473), .ZN(Result_mul_12_) );
  XOR2_X1 U476 ( .A(n474), .B(n475), .Z(n473) );
  XNOR2_X1 U477 ( .A(n476), .B(n477), .ZN(Result_mul_11_) );
  XOR2_X1 U478 ( .A(n478), .B(n479), .Z(n477) );
  XNOR2_X1 U479 ( .A(n480), .B(n481), .ZN(Result_mul_10_) );
  XOR2_X1 U480 ( .A(n482), .B(n483), .Z(n481) );
  OR2_X1 U481 ( .A1(n484), .A2(n485), .ZN(Result_mul_0_) );
  OR2_X1 U482 ( .A1(n465), .A2(n486), .ZN(n485) );
  AND2_X1 U483 ( .A1(n457), .A2(n462), .ZN(n486) );
  AND2_X1 U484 ( .A1(n455), .A2(n456), .ZN(n457) );
  XNOR2_X1 U485 ( .A(n464), .B(n487), .ZN(n456) );
  OR2_X1 U486 ( .A1(n488), .A2(n489), .ZN(n455) );
  OR2_X1 U487 ( .A1(n490), .A2(n454), .ZN(n488) );
  AND2_X1 U488 ( .A1(n452), .A2(n453), .ZN(n454) );
  AND2_X1 U489 ( .A1(n491), .A2(n492), .ZN(n453) );
  INV_X1 U490 ( .A(n493), .ZN(n491) );
  AND2_X1 U491 ( .A1(n448), .A2(n452), .ZN(n490) );
  INV_X1 U492 ( .A(n494), .ZN(n452) );
  OR2_X1 U493 ( .A1(n495), .A2(n489), .ZN(n494) );
  INV_X1 U494 ( .A(n496), .ZN(n489) );
  OR2_X1 U495 ( .A1(n497), .A2(n498), .ZN(n496) );
  AND2_X1 U496 ( .A1(n497), .A2(n498), .ZN(n495) );
  OR2_X1 U497 ( .A1(n499), .A2(n500), .ZN(n498) );
  AND2_X1 U498 ( .A1(n501), .A2(n502), .ZN(n500) );
  AND2_X1 U499 ( .A1(n503), .A2(n504), .ZN(n499) );
  OR2_X1 U500 ( .A1(n502), .A2(n501), .ZN(n504) );
  XOR2_X1 U501 ( .A(n505), .B(n506), .Z(n497) );
  XOR2_X1 U502 ( .A(n507), .B(n508), .Z(n506) );
  AND2_X1 U503 ( .A1(n509), .A2(n445), .ZN(n448) );
  XNOR2_X1 U504 ( .A(n492), .B(n493), .ZN(n445) );
  OR2_X1 U505 ( .A1(n510), .A2(n511), .ZN(n493) );
  AND2_X1 U506 ( .A1(n512), .A2(n513), .ZN(n511) );
  AND2_X1 U507 ( .A1(n514), .A2(n515), .ZN(n510) );
  OR2_X1 U508 ( .A1(n513), .A2(n512), .ZN(n515) );
  XOR2_X1 U509 ( .A(n516), .B(n503), .Z(n492) );
  XOR2_X1 U510 ( .A(n517), .B(n518), .Z(n503) );
  XOR2_X1 U511 ( .A(n519), .B(n520), .Z(n518) );
  XNOR2_X1 U512 ( .A(n502), .B(n501), .ZN(n516) );
  OR2_X1 U513 ( .A1(n521), .A2(n522), .ZN(n501) );
  AND2_X1 U514 ( .A1(n523), .A2(n524), .ZN(n522) );
  AND2_X1 U515 ( .A1(n525), .A2(n526), .ZN(n521) );
  OR2_X1 U516 ( .A1(n524), .A2(n523), .ZN(n526) );
  OR2_X1 U517 ( .A1(n527), .A2(n528), .ZN(n502) );
  OR2_X1 U518 ( .A1(n529), .A2(n530), .ZN(n509) );
  INV_X1 U519 ( .A(n447), .ZN(n529) );
  AND2_X1 U520 ( .A1(n531), .A2(n532), .ZN(n447) );
  OR2_X1 U521 ( .A1(n443), .A2(n441), .ZN(n532) );
  OR2_X1 U522 ( .A1(n435), .A2(n441), .ZN(n531) );
  OR2_X1 U523 ( .A1(n533), .A2(n530), .ZN(n441) );
  INV_X1 U524 ( .A(n446), .ZN(n530) );
  OR2_X1 U525 ( .A1(n534), .A2(n535), .ZN(n446) );
  AND2_X1 U526 ( .A1(n534), .A2(n535), .ZN(n533) );
  OR2_X1 U527 ( .A1(n536), .A2(n537), .ZN(n535) );
  AND2_X1 U528 ( .A1(n538), .A2(n539), .ZN(n537) );
  AND2_X1 U529 ( .A1(n540), .A2(n541), .ZN(n536) );
  OR2_X1 U530 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U531 ( .A(n514), .B(n542), .Z(n534) );
  XOR2_X1 U532 ( .A(n513), .B(n512), .Z(n542) );
  OR2_X1 U533 ( .A1(n543), .A2(n528), .ZN(n512) );
  OR2_X1 U534 ( .A1(n544), .A2(n545), .ZN(n513) );
  AND2_X1 U535 ( .A1(n546), .A2(n547), .ZN(n545) );
  AND2_X1 U536 ( .A1(n548), .A2(n549), .ZN(n544) );
  OR2_X1 U537 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U538 ( .A(n550), .B(n525), .ZN(n514) );
  XNOR2_X1 U539 ( .A(n551), .B(n552), .ZN(n525) );
  XNOR2_X1 U540 ( .A(n553), .B(n554), .ZN(n551) );
  XNOR2_X1 U541 ( .A(n524), .B(n523), .ZN(n550) );
  OR2_X1 U542 ( .A1(n555), .A2(n556), .ZN(n523) );
  AND2_X1 U543 ( .A1(n557), .A2(n558), .ZN(n556) );
  AND2_X1 U544 ( .A1(n559), .A2(n560), .ZN(n555) );
  OR2_X1 U545 ( .A1(n558), .A2(n557), .ZN(n560) );
  OR2_X1 U546 ( .A1(n527), .A2(n561), .ZN(n524) );
  OR2_X1 U547 ( .A1(n562), .A2(n440), .ZN(n435) );
  OR2_X1 U548 ( .A1(n433), .A2(n432), .ZN(n440) );
  OR2_X1 U549 ( .A1(n563), .A2(n564), .ZN(n432) );
  AND2_X1 U550 ( .A1(n431), .A2(n430), .ZN(n564) );
  AND2_X1 U551 ( .A1(n428), .A2(n565), .ZN(n563) );
  OR2_X1 U552 ( .A1(n430), .A2(n431), .ZN(n565) );
  OR2_X1 U553 ( .A1(n566), .A2(n528), .ZN(n431) );
  OR2_X1 U554 ( .A1(n567), .A2(n568), .ZN(n430) );
  AND2_X1 U555 ( .A1(n427), .A2(n426), .ZN(n568) );
  AND2_X1 U556 ( .A1(n424), .A2(n569), .ZN(n567) );
  OR2_X1 U557 ( .A1(n426), .A2(n427), .ZN(n569) );
  OR2_X1 U558 ( .A1(n566), .A2(n561), .ZN(n427) );
  OR2_X1 U559 ( .A1(n570), .A2(n571), .ZN(n426) );
  AND2_X1 U560 ( .A1(n483), .A2(n482), .ZN(n571) );
  AND2_X1 U561 ( .A1(n480), .A2(n572), .ZN(n570) );
  OR2_X1 U562 ( .A1(n483), .A2(n482), .ZN(n572) );
  OR2_X1 U563 ( .A1(n573), .A2(n574), .ZN(n482) );
  AND2_X1 U564 ( .A1(n479), .A2(n478), .ZN(n574) );
  AND2_X1 U565 ( .A1(n476), .A2(n575), .ZN(n573) );
  OR2_X1 U566 ( .A1(n479), .A2(n478), .ZN(n575) );
  OR2_X1 U567 ( .A1(n576), .A2(n577), .ZN(n478) );
  AND2_X1 U568 ( .A1(n475), .A2(n474), .ZN(n577) );
  AND2_X1 U569 ( .A1(n472), .A2(n578), .ZN(n576) );
  OR2_X1 U570 ( .A1(n475), .A2(n474), .ZN(n578) );
  OR2_X1 U571 ( .A1(n579), .A2(n580), .ZN(n474) );
  AND2_X1 U572 ( .A1(n470), .A2(n471), .ZN(n580) );
  AND2_X1 U573 ( .A1(n468), .A2(n581), .ZN(n579) );
  OR2_X1 U574 ( .A1(n470), .A2(n471), .ZN(n581) );
  INV_X1 U575 ( .A(n582), .ZN(n471) );
  OR2_X1 U576 ( .A1(n583), .A2(n566), .ZN(n470) );
  XOR2_X1 U577 ( .A(n584), .B(n585), .Z(n468) );
  OR2_X1 U578 ( .A1(n586), .A2(n587), .ZN(n584) );
  OR2_X1 U579 ( .A1(n588), .A2(n566), .ZN(n475) );
  XNOR2_X1 U580 ( .A(n589), .B(n590), .ZN(n472) );
  XNOR2_X1 U581 ( .A(n591), .B(n592), .ZN(n589) );
  OR2_X1 U582 ( .A1(n593), .A2(n566), .ZN(n479) );
  XOR2_X1 U583 ( .A(n594), .B(n595), .Z(n476) );
  XOR2_X1 U584 ( .A(n596), .B(n597), .Z(n595) );
  OR2_X1 U585 ( .A1(n598), .A2(n566), .ZN(n483) );
  XOR2_X1 U586 ( .A(n599), .B(n600), .Z(n480) );
  XOR2_X1 U587 ( .A(n601), .B(n602), .Z(n600) );
  XOR2_X1 U588 ( .A(n603), .B(n604), .Z(n424) );
  XOR2_X1 U589 ( .A(n605), .B(n606), .Z(n604) );
  XOR2_X1 U590 ( .A(n607), .B(n608), .Z(n428) );
  XOR2_X1 U591 ( .A(n609), .B(n610), .Z(n608) );
  XOR2_X1 U592 ( .A(n611), .B(n612), .Z(n433) );
  XOR2_X1 U593 ( .A(n613), .B(n614), .Z(n612) );
  OR2_X1 U594 ( .A1(n615), .A2(n616), .ZN(n562) );
  AND2_X1 U595 ( .A1(n438), .A2(n439), .ZN(n616) );
  INV_X1 U596 ( .A(n443), .ZN(n615) );
  OR2_X1 U597 ( .A1(n438), .A2(n439), .ZN(n443) );
  OR2_X1 U598 ( .A1(n617), .A2(n618), .ZN(n439) );
  AND2_X1 U599 ( .A1(n614), .A2(n613), .ZN(n618) );
  AND2_X1 U600 ( .A1(n611), .A2(n619), .ZN(n617) );
  OR2_X1 U601 ( .A1(n613), .A2(n614), .ZN(n619) );
  OR2_X1 U602 ( .A1(n620), .A2(n528), .ZN(n614) );
  OR2_X1 U603 ( .A1(n621), .A2(n622), .ZN(n613) );
  AND2_X1 U604 ( .A1(n610), .A2(n609), .ZN(n622) );
  AND2_X1 U605 ( .A1(n607), .A2(n623), .ZN(n621) );
  OR2_X1 U606 ( .A1(n609), .A2(n610), .ZN(n623) );
  OR2_X1 U607 ( .A1(n620), .A2(n561), .ZN(n610) );
  OR2_X1 U608 ( .A1(n624), .A2(n625), .ZN(n609) );
  AND2_X1 U609 ( .A1(n606), .A2(n605), .ZN(n625) );
  AND2_X1 U610 ( .A1(n603), .A2(n626), .ZN(n624) );
  OR2_X1 U611 ( .A1(n605), .A2(n606), .ZN(n626) );
  OR2_X1 U612 ( .A1(n620), .A2(n598), .ZN(n606) );
  OR2_X1 U613 ( .A1(n627), .A2(n628), .ZN(n605) );
  AND2_X1 U614 ( .A1(n602), .A2(n601), .ZN(n628) );
  AND2_X1 U615 ( .A1(n599), .A2(n629), .ZN(n627) );
  OR2_X1 U616 ( .A1(n602), .A2(n601), .ZN(n629) );
  OR2_X1 U617 ( .A1(n630), .A2(n631), .ZN(n601) );
  AND2_X1 U618 ( .A1(n597), .A2(n596), .ZN(n631) );
  AND2_X1 U619 ( .A1(n594), .A2(n632), .ZN(n630) );
  OR2_X1 U620 ( .A1(n597), .A2(n596), .ZN(n632) );
  OR2_X1 U621 ( .A1(n633), .A2(n634), .ZN(n596) );
  AND2_X1 U622 ( .A1(n591), .A2(n592), .ZN(n634) );
  AND2_X1 U623 ( .A1(n590), .A2(n635), .ZN(n633) );
  OR2_X1 U624 ( .A1(n591), .A2(n592), .ZN(n635) );
  OR2_X1 U625 ( .A1(n466), .A2(n636), .ZN(n592) );
  OR2_X1 U626 ( .A1(n586), .A2(n620), .ZN(n466) );
  OR2_X1 U627 ( .A1(n583), .A2(n620), .ZN(n591) );
  XNOR2_X1 U628 ( .A(n637), .B(n636), .ZN(n590) );
  OR2_X1 U629 ( .A1(n638), .A2(n587), .ZN(n636) );
  OR2_X1 U630 ( .A1(n586), .A2(n543), .ZN(n637) );
  OR2_X1 U631 ( .A1(n588), .A2(n620), .ZN(n597) );
  XOR2_X1 U632 ( .A(n639), .B(n640), .Z(n594) );
  XOR2_X1 U633 ( .A(n641), .B(n642), .Z(n640) );
  OR2_X1 U634 ( .A1(n593), .A2(n620), .ZN(n602) );
  XOR2_X1 U635 ( .A(n643), .B(n644), .Z(n599) );
  XOR2_X1 U636 ( .A(n645), .B(n646), .Z(n644) );
  XOR2_X1 U637 ( .A(n647), .B(n648), .Z(n603) );
  XOR2_X1 U638 ( .A(n649), .B(n650), .Z(n648) );
  XOR2_X1 U639 ( .A(n651), .B(n652), .Z(n607) );
  XOR2_X1 U640 ( .A(n653), .B(n654), .Z(n652) );
  XOR2_X1 U641 ( .A(n655), .B(n656), .Z(n611) );
  XOR2_X1 U642 ( .A(n657), .B(n658), .Z(n656) );
  XOR2_X1 U643 ( .A(n538), .B(n659), .Z(n438) );
  XOR2_X1 U644 ( .A(n541), .B(n539), .Z(n659) );
  OR2_X1 U645 ( .A1(n587), .A2(n528), .ZN(n539) );
  OR2_X1 U646 ( .A1(n660), .A2(n661), .ZN(n541) );
  AND2_X1 U647 ( .A1(n658), .A2(n657), .ZN(n661) );
  AND2_X1 U648 ( .A1(n655), .A2(n662), .ZN(n660) );
  OR2_X1 U649 ( .A1(n657), .A2(n658), .ZN(n662) );
  OR2_X1 U650 ( .A1(n587), .A2(n561), .ZN(n658) );
  OR2_X1 U651 ( .A1(n663), .A2(n664), .ZN(n657) );
  AND2_X1 U652 ( .A1(n654), .A2(n653), .ZN(n664) );
  AND2_X1 U653 ( .A1(n651), .A2(n665), .ZN(n663) );
  OR2_X1 U654 ( .A1(n653), .A2(n654), .ZN(n665) );
  OR2_X1 U655 ( .A1(n587), .A2(n598), .ZN(n654) );
  OR2_X1 U656 ( .A1(n666), .A2(n667), .ZN(n653) );
  AND2_X1 U657 ( .A1(n650), .A2(n649), .ZN(n667) );
  AND2_X1 U658 ( .A1(n647), .A2(n668), .ZN(n666) );
  OR2_X1 U659 ( .A1(n649), .A2(n650), .ZN(n668) );
  OR2_X1 U660 ( .A1(n587), .A2(n593), .ZN(n650) );
  OR2_X1 U661 ( .A1(n669), .A2(n670), .ZN(n649) );
  AND2_X1 U662 ( .A1(n646), .A2(n645), .ZN(n670) );
  AND2_X1 U663 ( .A1(n643), .A2(n671), .ZN(n669) );
  OR2_X1 U664 ( .A1(n646), .A2(n645), .ZN(n671) );
  OR2_X1 U665 ( .A1(n672), .A2(n673), .ZN(n645) );
  AND2_X1 U666 ( .A1(n639), .A2(n641), .ZN(n673) );
  AND2_X1 U667 ( .A1(n674), .A2(n642), .ZN(n672) );
  OR2_X1 U668 ( .A1(n639), .A2(n641), .ZN(n674) );
  OR2_X1 U669 ( .A1(n587), .A2(n675), .ZN(n641) );
  OR2_X1 U670 ( .A1(n586), .A2(n676), .ZN(n675) );
  OR2_X1 U671 ( .A1(n677), .A2(n678), .ZN(n639) );
  INV_X1 U672 ( .A(n679), .ZN(n678) );
  AND2_X1 U673 ( .A1(n680), .A2(n676), .ZN(n677) );
  OR2_X1 U674 ( .A1(n588), .A2(n587), .ZN(n646) );
  XNOR2_X1 U675 ( .A(n681), .B(n682), .ZN(n643) );
  XNOR2_X1 U676 ( .A(n683), .B(n679), .ZN(n681) );
  XNOR2_X1 U677 ( .A(n684), .B(n685), .ZN(n647) );
  XNOR2_X1 U678 ( .A(n686), .B(n687), .ZN(n684) );
  XOR2_X1 U679 ( .A(n688), .B(n689), .Z(n651) );
  XOR2_X1 U680 ( .A(n690), .B(n691), .Z(n689) );
  XOR2_X1 U681 ( .A(n692), .B(n693), .Z(n655) );
  XOR2_X1 U682 ( .A(n694), .B(n695), .Z(n693) );
  XOR2_X1 U683 ( .A(n546), .B(n696), .Z(n538) );
  XOR2_X1 U684 ( .A(n549), .B(n547), .Z(n696) );
  OR2_X1 U685 ( .A1(n543), .A2(n561), .ZN(n547) );
  OR2_X1 U686 ( .A1(n697), .A2(n698), .ZN(n549) );
  AND2_X1 U687 ( .A1(n695), .A2(n694), .ZN(n698) );
  AND2_X1 U688 ( .A1(n692), .A2(n699), .ZN(n697) );
  OR2_X1 U689 ( .A1(n694), .A2(n695), .ZN(n699) );
  OR2_X1 U690 ( .A1(n543), .A2(n598), .ZN(n695) );
  OR2_X1 U691 ( .A1(n700), .A2(n701), .ZN(n694) );
  AND2_X1 U692 ( .A1(n691), .A2(n690), .ZN(n701) );
  AND2_X1 U693 ( .A1(n688), .A2(n702), .ZN(n700) );
  OR2_X1 U694 ( .A1(n690), .A2(n691), .ZN(n702) );
  OR2_X1 U695 ( .A1(n543), .A2(n593), .ZN(n691) );
  OR2_X1 U696 ( .A1(n703), .A2(n704), .ZN(n690) );
  AND2_X1 U697 ( .A1(n685), .A2(n687), .ZN(n704) );
  AND2_X1 U698 ( .A1(n705), .A2(n686), .ZN(n703) );
  OR2_X1 U699 ( .A1(n685), .A2(n687), .ZN(n705) );
  OR2_X1 U700 ( .A1(n706), .A2(n707), .ZN(n687) );
  AND2_X1 U701 ( .A1(n682), .A2(n679), .ZN(n707) );
  AND2_X1 U702 ( .A1(n708), .A2(n683), .ZN(n706) );
  OR2_X1 U703 ( .A1(n709), .A2(n710), .ZN(n683) );
  AND2_X1 U704 ( .A1(n711), .A2(n712), .ZN(n709) );
  OR2_X1 U705 ( .A1(n682), .A2(n679), .ZN(n708) );
  OR2_X1 U706 ( .A1(n680), .A2(n676), .ZN(n679) );
  OR2_X1 U707 ( .A1(n638), .A2(n543), .ZN(n676) );
  OR2_X1 U708 ( .A1(n586), .A2(n527), .ZN(n680) );
  OR2_X1 U709 ( .A1(n583), .A2(n543), .ZN(n682) );
  XOR2_X1 U710 ( .A(n713), .B(n710), .Z(n685) );
  INV_X1 U711 ( .A(n714), .ZN(n710) );
  XNOR2_X1 U712 ( .A(n715), .B(n716), .ZN(n713) );
  XNOR2_X1 U713 ( .A(n717), .B(n718), .ZN(n688) );
  XNOR2_X1 U714 ( .A(n719), .B(n720), .ZN(n717) );
  XNOR2_X1 U715 ( .A(n721), .B(n722), .ZN(n692) );
  XNOR2_X1 U716 ( .A(n723), .B(n724), .ZN(n721) );
  XNOR2_X1 U717 ( .A(n725), .B(n559), .ZN(n546) );
  XNOR2_X1 U718 ( .A(n726), .B(n727), .ZN(n559) );
  XNOR2_X1 U719 ( .A(n728), .B(n729), .ZN(n726) );
  XNOR2_X1 U720 ( .A(n558), .B(n557), .ZN(n725) );
  OR2_X1 U721 ( .A1(n730), .A2(n731), .ZN(n557) );
  AND2_X1 U722 ( .A1(n722), .A2(n724), .ZN(n731) );
  AND2_X1 U723 ( .A1(n732), .A2(n723), .ZN(n730) );
  OR2_X1 U724 ( .A1(n722), .A2(n724), .ZN(n732) );
  OR2_X1 U725 ( .A1(n733), .A2(n734), .ZN(n724) );
  AND2_X1 U726 ( .A1(n720), .A2(n719), .ZN(n734) );
  AND2_X1 U727 ( .A1(n718), .A2(n735), .ZN(n733) );
  OR2_X1 U728 ( .A1(n719), .A2(n720), .ZN(n735) );
  OR2_X1 U729 ( .A1(n736), .A2(n737), .ZN(n720) );
  AND2_X1 U730 ( .A1(n714), .A2(n716), .ZN(n737) );
  AND2_X1 U731 ( .A1(n738), .A2(n715), .ZN(n736) );
  OR2_X1 U732 ( .A1(n739), .A2(n740), .ZN(n715) );
  INV_X1 U733 ( .A(n741), .ZN(n740) );
  AND2_X1 U734 ( .A1(n742), .A2(n743), .ZN(n739) );
  OR2_X1 U735 ( .A1(n716), .A2(n714), .ZN(n738) );
  OR2_X1 U736 ( .A1(n711), .A2(n712), .ZN(n714) );
  OR2_X1 U737 ( .A1(n586), .A2(n744), .ZN(n712) );
  OR2_X1 U738 ( .A1(n638), .A2(n527), .ZN(n711) );
  OR2_X1 U739 ( .A1(n527), .A2(n583), .ZN(n716) );
  OR2_X1 U740 ( .A1(n527), .A2(n588), .ZN(n719) );
  XNOR2_X1 U741 ( .A(n745), .B(n746), .ZN(n718) );
  XNOR2_X1 U742 ( .A(n747), .B(n741), .ZN(n745) );
  XOR2_X1 U743 ( .A(n748), .B(n749), .Z(n722) );
  XOR2_X1 U744 ( .A(n750), .B(n751), .Z(n749) );
  OR2_X1 U745 ( .A1(n527), .A2(n598), .ZN(n558) );
  AND2_X1 U746 ( .A1(n463), .A2(n752), .ZN(n465) );
  AND2_X1 U747 ( .A1(n464), .A2(n462), .ZN(n752) );
  XOR2_X1 U748 ( .A(n753), .B(n754), .Z(n462) );
  OR2_X1 U749 ( .A1(n755), .A2(n528), .ZN(n753) );
  XNOR2_X1 U750 ( .A(n756), .B(n757), .ZN(n464) );
  XOR2_X1 U751 ( .A(n758), .B(n759), .Z(n757) );
  INV_X1 U752 ( .A(n487), .ZN(n463) );
  OR2_X1 U753 ( .A1(n760), .A2(n761), .ZN(n487) );
  AND2_X1 U754 ( .A1(n508), .A2(n507), .ZN(n761) );
  AND2_X1 U755 ( .A1(n505), .A2(n762), .ZN(n760) );
  OR2_X1 U756 ( .A1(n507), .A2(n508), .ZN(n762) );
  OR2_X1 U757 ( .A1(n744), .A2(n528), .ZN(n508) );
  OR2_X1 U758 ( .A1(n763), .A2(n764), .ZN(n507) );
  AND2_X1 U759 ( .A1(n520), .A2(n519), .ZN(n764) );
  AND2_X1 U760 ( .A1(n517), .A2(n765), .ZN(n763) );
  OR2_X1 U761 ( .A1(n519), .A2(n520), .ZN(n765) );
  OR2_X1 U762 ( .A1(n744), .A2(n561), .ZN(n520) );
  OR2_X1 U763 ( .A1(n766), .A2(n767), .ZN(n519) );
  AND2_X1 U764 ( .A1(n552), .A2(n554), .ZN(n767) );
  AND2_X1 U765 ( .A1(n768), .A2(n553), .ZN(n766) );
  OR2_X1 U766 ( .A1(n552), .A2(n554), .ZN(n768) );
  OR2_X1 U767 ( .A1(n769), .A2(n770), .ZN(n554) );
  AND2_X1 U768 ( .A1(n729), .A2(n728), .ZN(n770) );
  AND2_X1 U769 ( .A1(n727), .A2(n771), .ZN(n769) );
  OR2_X1 U770 ( .A1(n728), .A2(n729), .ZN(n771) );
  OR2_X1 U771 ( .A1(n772), .A2(n773), .ZN(n729) );
  AND2_X1 U772 ( .A1(n751), .A2(n750), .ZN(n773) );
  AND2_X1 U773 ( .A1(n748), .A2(n774), .ZN(n772) );
  OR2_X1 U774 ( .A1(n750), .A2(n751), .ZN(n774) );
  OR2_X1 U775 ( .A1(n744), .A2(n588), .ZN(n751) );
  OR2_X1 U776 ( .A1(n775), .A2(n776), .ZN(n750) );
  AND2_X1 U777 ( .A1(n746), .A2(n741), .ZN(n776) );
  AND2_X1 U778 ( .A1(n777), .A2(n747), .ZN(n775) );
  OR2_X1 U779 ( .A1(n778), .A2(n779), .ZN(n747) );
  INV_X1 U780 ( .A(n780), .ZN(n779) );
  AND2_X1 U781 ( .A1(n781), .A2(n782), .ZN(n778) );
  OR2_X1 U782 ( .A1(n741), .A2(n746), .ZN(n777) );
  OR2_X1 U783 ( .A1(n744), .A2(n583), .ZN(n746) );
  OR2_X1 U784 ( .A1(n742), .A2(n743), .ZN(n741) );
  OR2_X1 U785 ( .A1(n744), .A2(n638), .ZN(n743) );
  OR2_X1 U786 ( .A1(n586), .A2(n783), .ZN(n742) );
  XNOR2_X1 U787 ( .A(n784), .B(n780), .ZN(n748) );
  OR2_X1 U788 ( .A1(n785), .A2(n786), .ZN(n784) );
  INV_X1 U789 ( .A(n787), .ZN(n786) );
  AND2_X1 U790 ( .A1(n788), .A2(n789), .ZN(n785) );
  OR2_X1 U791 ( .A1(n744), .A2(n593), .ZN(n728) );
  XOR2_X1 U792 ( .A(n790), .B(n791), .Z(n727) );
  XOR2_X1 U793 ( .A(n792), .B(n793), .Z(n790) );
  XOR2_X1 U794 ( .A(n794), .B(n795), .Z(n552) );
  XOR2_X1 U795 ( .A(n796), .B(n797), .Z(n795) );
  XOR2_X1 U796 ( .A(n798), .B(n799), .Z(n517) );
  XOR2_X1 U797 ( .A(n800), .B(n801), .Z(n799) );
  XOR2_X1 U798 ( .A(n802), .B(n803), .Z(n505) );
  XOR2_X1 U799 ( .A(n804), .B(n805), .Z(n803) );
  AND2_X1 U800 ( .A1(n806), .A2(a_0_), .ZN(n484) );
  INV_X1 U801 ( .A(n754), .ZN(n806) );
  OR2_X1 U802 ( .A1(n807), .A2(n808), .ZN(n754) );
  AND2_X1 U803 ( .A1(n756), .A2(n758), .ZN(n808) );
  AND2_X1 U804 ( .A1(n809), .A2(n759), .ZN(n807) );
  OR2_X1 U805 ( .A1(n783), .A2(n528), .ZN(n759) );
  INV_X1 U806 ( .A(a_0_), .ZN(n528) );
  OR2_X1 U807 ( .A1(n758), .A2(n756), .ZN(n809) );
  OR2_X1 U808 ( .A1(n561), .A2(n755), .ZN(n756) );
  OR2_X1 U809 ( .A1(n810), .A2(n811), .ZN(n758) );
  AND2_X1 U810 ( .A1(n802), .A2(n804), .ZN(n811) );
  AND2_X1 U811 ( .A1(n812), .A2(n805), .ZN(n810) );
  OR2_X1 U812 ( .A1(n804), .A2(n802), .ZN(n812) );
  OR2_X1 U813 ( .A1(n598), .A2(n755), .ZN(n802) );
  OR2_X1 U814 ( .A1(n813), .A2(n814), .ZN(n804) );
  AND2_X1 U815 ( .A1(n798), .A2(n800), .ZN(n814) );
  AND2_X1 U816 ( .A1(n815), .A2(n801), .ZN(n813) );
  OR2_X1 U817 ( .A1(n593), .A2(n755), .ZN(n801) );
  OR2_X1 U818 ( .A1(n800), .A2(n798), .ZN(n815) );
  OR2_X1 U819 ( .A1(n783), .A2(n598), .ZN(n798) );
  OR2_X1 U820 ( .A1(n816), .A2(n817), .ZN(n800) );
  AND2_X1 U821 ( .A1(n794), .A2(n796), .ZN(n817) );
  AND2_X1 U822 ( .A1(n818), .A2(n797), .ZN(n816) );
  OR2_X1 U823 ( .A1(n783), .A2(n593), .ZN(n797) );
  OR2_X1 U824 ( .A1(n796), .A2(n794), .ZN(n818) );
  OR2_X1 U825 ( .A1(n588), .A2(n755), .ZN(n794) );
  OR2_X1 U826 ( .A1(n819), .A2(n820), .ZN(n796) );
  AND2_X1 U827 ( .A1(n791), .A2(n793), .ZN(n820) );
  AND2_X1 U828 ( .A1(n792), .A2(n821), .ZN(n819) );
  OR2_X1 U829 ( .A1(n793), .A2(n791), .ZN(n821) );
  OR2_X1 U830 ( .A1(n583), .A2(n755), .ZN(n791) );
  OR2_X1 U831 ( .A1(n783), .A2(n588), .ZN(n793) );
  AND2_X1 U832 ( .A1(n787), .A2(n780), .ZN(n792) );
  OR2_X1 U833 ( .A1(n782), .A2(n781), .ZN(n780) );
  OR2_X1 U834 ( .A1(n586), .A2(n755), .ZN(n781) );
  INV_X1 U835 ( .A(a_7_), .ZN(n586) );
  OR2_X1 U836 ( .A1(n638), .A2(n783), .ZN(n782) );
  OR2_X1 U837 ( .A1(n789), .A2(n788), .ZN(n787) );
  OR2_X1 U838 ( .A1(n638), .A2(n755), .ZN(n788) );
  INV_X1 U839 ( .A(b_0_), .ZN(n755) );
  OR2_X1 U840 ( .A1(n783), .A2(n583), .ZN(n789) );
  XNOR2_X1 U841 ( .A(n566), .B(a_7_), .ZN(Result_add_7_) );
  INV_X1 U842 ( .A(b_7_), .ZN(n566) );
  OR2_X1 U843 ( .A1(n582), .A2(n822), .ZN(Result_add_6_) );
  OR2_X1 U844 ( .A1(n823), .A2(n824), .ZN(n822) );
  INV_X1 U845 ( .A(n825), .ZN(n824) );
  OR2_X1 U846 ( .A1(n826), .A2(n620), .ZN(n825) );
  OR2_X1 U847 ( .A1(Result_mul_15_), .A2(a_6_), .ZN(n826) );
  AND2_X1 U848 ( .A1(n827), .A2(n620), .ZN(n823) );
  INV_X1 U849 ( .A(b_6_), .ZN(n620) );
  XNOR2_X1 U850 ( .A(n638), .B(Result_mul_15_), .ZN(n827) );
  INV_X1 U851 ( .A(a_6_), .ZN(n638) );
  AND2_X1 U852 ( .A1(n585), .A2(Result_mul_15_), .ZN(n582) );
  OR2_X1 U853 ( .A1(n828), .A2(n829), .ZN(Result_add_5_) );
  OR2_X1 U854 ( .A1(n830), .A2(n831), .ZN(n829) );
  AND2_X1 U855 ( .A1(n832), .A2(n587), .ZN(n831) );
  XNOR2_X1 U856 ( .A(n833), .B(a_5_), .ZN(n832) );
  AND2_X1 U857 ( .A1(n834), .A2(b_5_), .ZN(n830) );
  AND2_X1 U858 ( .A1(n833), .A2(n583), .ZN(n834) );
  INV_X1 U859 ( .A(n835), .ZN(n828) );
  OR2_X1 U860 ( .A1(n642), .A2(n833), .ZN(n835) );
  XNOR2_X1 U861 ( .A(n836), .B(n837), .ZN(Result_add_4_) );
  AND2_X1 U862 ( .A1(n686), .A2(n838), .ZN(n837) );
  OR2_X1 U863 ( .A1(n839), .A2(n840), .ZN(Result_add_3_) );
  OR2_X1 U864 ( .A1(n841), .A2(n842), .ZN(n840) );
  AND2_X1 U865 ( .A1(n843), .A2(n527), .ZN(n842) );
  XNOR2_X1 U866 ( .A(n593), .B(n844), .ZN(n843) );
  AND2_X1 U867 ( .A1(n845), .A2(b_3_), .ZN(n841) );
  AND2_X1 U868 ( .A1(n846), .A2(n593), .ZN(n845) );
  AND2_X1 U869 ( .A1(n844), .A2(n847), .ZN(n839) );
  XNOR2_X1 U870 ( .A(n848), .B(n849), .ZN(Result_add_2_) );
  AND2_X1 U871 ( .A1(n553), .A2(n850), .ZN(n849) );
  OR2_X1 U872 ( .A1(n851), .A2(n852), .ZN(Result_add_1_) );
  OR2_X1 U873 ( .A1(n853), .A2(n854), .ZN(n852) );
  AND2_X1 U874 ( .A1(n855), .A2(n783), .ZN(n854) );
  XNOR2_X1 U875 ( .A(n561), .B(n856), .ZN(n855) );
  AND2_X1 U876 ( .A1(n857), .A2(b_1_), .ZN(n853) );
  AND2_X1 U877 ( .A1(n858), .A2(n561), .ZN(n857) );
  INV_X1 U878 ( .A(n859), .ZN(n851) );
  OR2_X1 U879 ( .A1(n858), .A2(n805), .ZN(n859) );
  XOR2_X1 U880 ( .A(n860), .B(n861), .Z(Result_add_0_) );
  XNOR2_X1 U881 ( .A(a_0_), .B(b_0_), .ZN(n861) );
  OR2_X1 U882 ( .A1(n862), .A2(n863), .ZN(n860) );
  AND2_X1 U883 ( .A1(n561), .A2(n783), .ZN(n863) );
  AND2_X1 U884 ( .A1(n858), .A2(n805), .ZN(n862) );
  OR2_X1 U885 ( .A1(n783), .A2(n561), .ZN(n805) );
  INV_X1 U886 ( .A(a_1_), .ZN(n561) );
  INV_X1 U887 ( .A(b_1_), .ZN(n783) );
  INV_X1 U888 ( .A(n856), .ZN(n858) );
  AND2_X1 U889 ( .A1(n864), .A2(n850), .ZN(n856) );
  OR2_X1 U890 ( .A1(a_2_), .A2(b_2_), .ZN(n850) );
  INV_X1 U891 ( .A(n865), .ZN(n864) );
  AND2_X1 U892 ( .A1(n848), .A2(n553), .ZN(n865) );
  OR2_X1 U893 ( .A1(n744), .A2(n598), .ZN(n553) );
  INV_X1 U894 ( .A(a_2_), .ZN(n598) );
  INV_X1 U895 ( .A(b_2_), .ZN(n744) );
  OR2_X1 U896 ( .A1(n866), .A2(n867), .ZN(n848) );
  AND2_X1 U897 ( .A1(n593), .A2(n527), .ZN(n867) );
  INV_X1 U898 ( .A(b_3_), .ZN(n527) );
  INV_X1 U899 ( .A(a_3_), .ZN(n593) );
  AND2_X1 U900 ( .A1(n846), .A2(n723), .ZN(n866) );
  INV_X1 U901 ( .A(n847), .ZN(n723) );
  AND2_X1 U902 ( .A1(b_3_), .A2(a_3_), .ZN(n847) );
  INV_X1 U903 ( .A(n844), .ZN(n846) );
  AND2_X1 U904 ( .A1(n868), .A2(n838), .ZN(n844) );
  OR2_X1 U905 ( .A1(a_4_), .A2(b_4_), .ZN(n838) );
  INV_X1 U906 ( .A(n869), .ZN(n868) );
  AND2_X1 U907 ( .A1(n836), .A2(n686), .ZN(n869) );
  OR2_X1 U908 ( .A1(n588), .A2(n543), .ZN(n686) );
  INV_X1 U909 ( .A(b_4_), .ZN(n543) );
  INV_X1 U910 ( .A(a_4_), .ZN(n588) );
  OR2_X1 U911 ( .A1(n870), .A2(n871), .ZN(n836) );
  AND2_X1 U912 ( .A1(n583), .A2(n587), .ZN(n871) );
  AND2_X1 U913 ( .A1(n833), .A2(n642), .ZN(n870) );
  OR2_X1 U914 ( .A1(n583), .A2(n587), .ZN(n642) );
  INV_X1 U915 ( .A(b_5_), .ZN(n587) );
  INV_X1 U916 ( .A(a_5_), .ZN(n583) );
  INV_X1 U917 ( .A(n872), .ZN(n833) );
  OR2_X1 U918 ( .A1(n873), .A2(n585), .ZN(n872) );
  AND2_X1 U919 ( .A1(a_6_), .A2(b_6_), .ZN(n585) );
  AND2_X1 U920 ( .A1(Result_mul_15_), .A2(n874), .ZN(n873) );
  OR2_X1 U921 ( .A1(a_6_), .A2(b_6_), .ZN(n874) );
  AND2_X1 U922 ( .A1(a_7_), .A2(b_7_), .ZN(Result_mul_15_) );
endmodule

