module s35932 ( CK, CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_10, CRC_OUT_1_11, 
        CRC_OUT_1_12, CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, 
        CRC_OUT_1_17, CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_2, CRC_OUT_1_20, 
        CRC_OUT_1_21, CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, 
        CRC_OUT_1_26, CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_3, 
        CRC_OUT_1_30, CRC_OUT_1_31, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, 
        CRC_OUT_1_7, CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_2_0, CRC_OUT_2_1, 
        CRC_OUT_2_10, CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, 
        CRC_OUT_2_15, CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, 
        CRC_OUT_2_2, CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, 
        CRC_OUT_2_24, CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, 
        CRC_OUT_2_29, CRC_OUT_2_3, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_2_4, 
        CRC_OUT_2_5, CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, 
        CRC_OUT_3_0, CRC_OUT_3_1, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, 
        CRC_OUT_3_13, CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, 
        CRC_OUT_3_18, CRC_OUT_3_19, CRC_OUT_3_2, CRC_OUT_3_20, CRC_OUT_3_21, 
        CRC_OUT_3_22, CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, 
        CRC_OUT_3_27, CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_3, CRC_OUT_3_30, 
        CRC_OUT_3_31, CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, 
        CRC_OUT_3_8, CRC_OUT_3_9, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_10, 
        CRC_OUT_4_11, CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, 
        CRC_OUT_4_16, CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_2, 
        CRC_OUT_4_20, CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, 
        CRC_OUT_4_25, CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, 
        CRC_OUT_4_3, CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_4_4, CRC_OUT_4_5, 
        CRC_OUT_4_6, CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_5_0, 
        CRC_OUT_5_1, CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, 
        CRC_OUT_5_14, CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, 
        CRC_OUT_5_19, CRC_OUT_5_2, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, 
        CRC_OUT_5_23, CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, 
        CRC_OUT_5_28, CRC_OUT_5_29, CRC_OUT_5_3, CRC_OUT_5_30, CRC_OUT_5_31, 
        CRC_OUT_5_4, CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, 
        CRC_OUT_5_9, CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_10, CRC_OUT_6_11, 
        CRC_OUT_6_12, CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, 
        CRC_OUT_6_17, CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_2, CRC_OUT_6_20, 
        CRC_OUT_6_21, CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, 
        CRC_OUT_6_26, CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_3, 
        CRC_OUT_6_30, CRC_OUT_6_31, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, 
        CRC_OUT_6_7, CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_7_0, CRC_OUT_7_1, 
        CRC_OUT_7_10, CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, 
        CRC_OUT_7_15, CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, 
        CRC_OUT_7_2, CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, 
        CRC_OUT_7_24, CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, 
        CRC_OUT_7_29, CRC_OUT_7_3, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_7_4, 
        CRC_OUT_7_5, CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, 
        CRC_OUT_8_0, CRC_OUT_8_1, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, 
        CRC_OUT_8_13, CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, 
        CRC_OUT_8_18, CRC_OUT_8_19, CRC_OUT_8_2, CRC_OUT_8_20, CRC_OUT_8_21, 
        CRC_OUT_8_22, CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, 
        CRC_OUT_8_27, CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_3, CRC_OUT_8_30, 
        CRC_OUT_8_31, CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, 
        CRC_OUT_8_8, CRC_OUT_8_9, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_10, 
        CRC_OUT_9_11, CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, 
        CRC_OUT_9_16, CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_2, 
        CRC_OUT_9_20, CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, 
        CRC_OUT_9_25, CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, 
        CRC_OUT_9_3, CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_9_4, CRC_OUT_9_5, 
        CRC_OUT_9_6, CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, DATA_0_0, DATA_0_1, 
        DATA_0_10, DATA_0_11, DATA_0_12, DATA_0_13, DATA_0_14, DATA_0_15, 
        DATA_0_16, DATA_0_17, DATA_0_18, DATA_0_19, DATA_0_2, DATA_0_20, 
        DATA_0_21, DATA_0_22, DATA_0_23, DATA_0_24, DATA_0_25, DATA_0_26, 
        DATA_0_27, DATA_0_28, DATA_0_29, DATA_0_3, DATA_0_30, DATA_0_31, 
        DATA_0_4, DATA_0_5, DATA_0_6, DATA_0_7, DATA_0_8, DATA_0_9, DATA_9_0, 
        DATA_9_1, DATA_9_10, DATA_9_11, DATA_9_12, DATA_9_13, DATA_9_14, 
        DATA_9_15, DATA_9_16, DATA_9_17, DATA_9_18, DATA_9_19, DATA_9_2, 
        DATA_9_20, DATA_9_21, DATA_9_22, DATA_9_23, DATA_9_24, DATA_9_25, 
        DATA_9_26, DATA_9_27, DATA_9_28, DATA_9_29, DATA_9_3, DATA_9_30, 
        DATA_9_31, DATA_9_4, DATA_9_5, DATA_9_6, DATA_9_7, DATA_9_8, DATA_9_9, 
        RESET, TM0, TM1, test_se, test_si1, test_so1, test_si2, test_so2, 
        test_si3, test_so3, test_si4, test_so4, test_si5, test_so5, test_si6, 
        test_so6, test_si7, test_so7, test_si8, test_so8, test_si9, test_so9, 
        test_si10, test_so10, test_si11, test_so11, test_si12, test_so12, 
        test_si13, test_so13, test_si14, test_so14, test_si15, test_so15, 
        test_si16, test_so16, test_si17, test_so17, test_si18, test_so18, 
        test_si19, test_so19, test_si20, test_so20, test_si21, test_so21, 
        test_si22, test_so22, test_si23, test_so23, test_si24, test_so24, 
        test_si25, test_so25, test_si26, test_so26, test_si27, test_so27, 
        test_si28, test_so28, test_si29, test_so29, test_si30, test_so30, 
        test_si31, test_so31, test_si32, test_so32, test_si33, test_so33, 
        test_si34, test_so34, test_si35, test_so35, test_si36, test_so36, 
        test_si37, test_so37, test_si38, test_so38, test_si39, test_so39, 
        test_si40, test_so40, test_si41, test_so41, test_si42, test_so42, 
        test_si43, test_so43, test_si44, test_so44, test_si45, test_so45, 
        test_si46, test_so46, test_si47, test_so47, test_si48, test_so48, 
        test_si49, test_so49, test_si50, test_so50, test_si51, test_so51, 
        test_si52, test_so52, test_si53, test_so53, test_si54, test_so54, 
        test_si55, test_so55, test_si56, test_so56, test_si57, test_so57, 
        test_si58, test_so58, test_si59, test_so59, test_si60, test_so60, 
        test_si61, test_so61, test_si62, test_so62, test_si63, test_so63, 
        test_si64, test_so64, test_si65, test_so65, test_si66, test_so66, 
        test_si67, test_so67, test_si68, test_so68, test_si69, test_so69, 
        test_si70, test_so70, test_si71, test_so71, test_si72, test_so72, 
        test_si73, test_so73, test_si74, test_so74, test_si75, test_so75, 
        test_si76, test_so76, test_si77, test_so77, test_si78, test_so78, 
        test_si79, test_so79, test_si80, test_so80, test_si81, test_so81, 
        test_si82, test_so82, test_si83, test_so83, test_si84, test_so84, 
        test_si85, test_so85, test_si86, test_so86, test_si87, test_so87, 
        test_si88, test_so88, test_si89, test_so89, test_si90, test_so90, 
        test_si91, test_so91, test_si92, test_so92, test_si93, test_so93, 
        test_si94, test_so94, test_si95, test_so95, test_si96, test_so96, 
        test_si97, test_so97, test_si98, test_so98, test_si99, test_so99, 
        test_si100, test_so100 );
  input CK, DATA_0_0, DATA_0_1, DATA_0_10, DATA_0_11, DATA_0_12, DATA_0_13,
         DATA_0_14, DATA_0_15, DATA_0_16, DATA_0_17, DATA_0_18, DATA_0_19,
         DATA_0_2, DATA_0_20, DATA_0_21, DATA_0_22, DATA_0_23, DATA_0_24,
         DATA_0_25, DATA_0_26, DATA_0_27, DATA_0_28, DATA_0_29, DATA_0_3,
         DATA_0_30, DATA_0_31, DATA_0_4, DATA_0_5, DATA_0_6, DATA_0_7,
         DATA_0_8, DATA_0_9, RESET, TM0, TM1, test_se, test_si1, test_si2,
         test_si3, test_si4, test_si5, test_si6, test_si7, test_si8, test_si9,
         test_si10, test_si11, test_si12, test_si13, test_si14, test_si15,
         test_si16, test_si17, test_si18, test_si19, test_si20, test_si21,
         test_si22, test_si23, test_si24, test_si25, test_si26, test_si27,
         test_si28, test_si29, test_si30, test_si31, test_si32, test_si33,
         test_si34, test_si35, test_si36, test_si37, test_si38, test_si39,
         test_si40, test_si41, test_si42, test_si43, test_si44, test_si45,
         test_si46, test_si47, test_si48, test_si49, test_si50, test_si51,
         test_si52, test_si53, test_si54, test_si55, test_si56, test_si57,
         test_si58, test_si59, test_si60, test_si61, test_si62, test_si63,
         test_si64, test_si65, test_si66, test_si67, test_si68, test_si69,
         test_si70, test_si71, test_si72, test_si73, test_si74, test_si75,
         test_si76, test_si77, test_si78, test_si79, test_si80, test_si81,
         test_si82, test_si83, test_si84, test_si85, test_si86, test_si87,
         test_si88, test_si89, test_si90, test_si91, test_si92, test_si93,
         test_si94, test_si95, test_si96, test_si97, test_si98, test_si99,
         test_si100;
  output CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_10, CRC_OUT_1_11, CRC_OUT_1_12,
         CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, CRC_OUT_1_17,
         CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_2, CRC_OUT_1_20, CRC_OUT_1_21,
         CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, CRC_OUT_1_26,
         CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_3, CRC_OUT_1_30,
         CRC_OUT_1_31, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, CRC_OUT_1_7,
         CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_2_0, CRC_OUT_2_1, CRC_OUT_2_10,
         CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, CRC_OUT_2_15,
         CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, CRC_OUT_2_2,
         CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, CRC_OUT_2_24,
         CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, CRC_OUT_2_29,
         CRC_OUT_2_3, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_2_4, CRC_OUT_2_5,
         CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, CRC_OUT_3_0,
         CRC_OUT_3_1, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, CRC_OUT_3_13,
         CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, CRC_OUT_3_18,
         CRC_OUT_3_19, CRC_OUT_3_2, CRC_OUT_3_20, CRC_OUT_3_21, CRC_OUT_3_22,
         CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, CRC_OUT_3_27,
         CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_3, CRC_OUT_3_30, CRC_OUT_3_31,
         CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, CRC_OUT_3_8,
         CRC_OUT_3_9, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_10, CRC_OUT_4_11,
         CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, CRC_OUT_4_16,
         CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_2, CRC_OUT_4_20,
         CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, CRC_OUT_4_25,
         CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, CRC_OUT_4_3,
         CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_4_4, CRC_OUT_4_5, CRC_OUT_4_6,
         CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_5_0, CRC_OUT_5_1,
         CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, CRC_OUT_5_14,
         CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, CRC_OUT_5_19,
         CRC_OUT_5_2, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, CRC_OUT_5_23,
         CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, CRC_OUT_5_28,
         CRC_OUT_5_29, CRC_OUT_5_3, CRC_OUT_5_30, CRC_OUT_5_31, CRC_OUT_5_4,
         CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, CRC_OUT_5_9,
         CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_10, CRC_OUT_6_11, CRC_OUT_6_12,
         CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, CRC_OUT_6_17,
         CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_2, CRC_OUT_6_20, CRC_OUT_6_21,
         CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, CRC_OUT_6_26,
         CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_3, CRC_OUT_6_30,
         CRC_OUT_6_31, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, CRC_OUT_6_7,
         CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_7_0, CRC_OUT_7_1, CRC_OUT_7_10,
         CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, CRC_OUT_7_15,
         CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, CRC_OUT_7_2,
         CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, CRC_OUT_7_24,
         CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, CRC_OUT_7_29,
         CRC_OUT_7_3, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_7_4, CRC_OUT_7_5,
         CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, CRC_OUT_8_0,
         CRC_OUT_8_1, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, CRC_OUT_8_13,
         CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, CRC_OUT_8_18,
         CRC_OUT_8_19, CRC_OUT_8_2, CRC_OUT_8_20, CRC_OUT_8_21, CRC_OUT_8_22,
         CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, CRC_OUT_8_27,
         CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_3, CRC_OUT_8_30, CRC_OUT_8_31,
         CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, CRC_OUT_8_8,
         CRC_OUT_8_9, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_10, CRC_OUT_9_11,
         CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, CRC_OUT_9_16,
         CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_2, CRC_OUT_9_20,
         CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, CRC_OUT_9_25,
         CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, CRC_OUT_9_3,
         CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_9_4, CRC_OUT_9_5, CRC_OUT_9_6,
         CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, DATA_9_0, DATA_9_1, DATA_9_10,
         DATA_9_11, DATA_9_12, DATA_9_13, DATA_9_14, DATA_9_15, DATA_9_16,
         DATA_9_17, DATA_9_18, DATA_9_19, DATA_9_2, DATA_9_20, DATA_9_21,
         DATA_9_22, DATA_9_23, DATA_9_24, DATA_9_25, DATA_9_26, DATA_9_27,
         DATA_9_28, DATA_9_29, DATA_9_3, DATA_9_30, DATA_9_31, DATA_9_4,
         DATA_9_5, DATA_9_6, DATA_9_7, DATA_9_8, DATA_9_9, test_so1, test_so2,
         test_so3, test_so4, test_so5, test_so6, test_so7, test_so8, test_so9,
         test_so10, test_so11, test_so12, test_so13, test_so14, test_so15,
         test_so16, test_so17, test_so18, test_so19, test_so20, test_so21,
         test_so22, test_so23, test_so24, test_so25, test_so26, test_so27,
         test_so28, test_so29, test_so30, test_so31, test_so32, test_so33,
         test_so34, test_so35, test_so36, test_so37, test_so38, test_so39,
         test_so40, test_so41, test_so42, test_so43, test_so44, test_so45,
         test_so46, test_so47, test_so48, test_so49, test_so50, test_so51,
         test_so52, test_so53, test_so54, test_so55, test_so56, test_so57,
         test_so58, test_so59, test_so60, test_so61, test_so62, test_so63,
         test_so64, test_so65, test_so66, test_so67, test_so68, test_so69,
         test_so70, test_so71, test_so72, test_so73, test_so74, test_so75,
         test_so76, test_so77, test_so78, test_so79, test_so80, test_so81,
         test_so82, test_so83, test_so84, test_so85, test_so86, test_so87,
         test_so88, test_so89, test_so90, test_so91, test_so92, test_so93,
         test_so94, test_so95, test_so96, test_so97, test_so98, test_so99,
         test_so100;
  wire   test_so9, test_so10, test_so20, test_so21, test_so31, test_so32,
         test_so42, test_so43, test_so53, test_so54, test_so65, test_so66,
         test_so76, test_so77, test_so87, test_so88, test_so99, test_so100,
         WX484, WX485, WX486, WX487, WX488, WX489, WX490, WX491, WX492, WX493,
         WX494, WX495, WX496, WX497, WX498, WX499, WX500, WX501, WX502, WX503,
         WX504, WX505, WX506, WX507, WX508, WX509, WX510, WX511, WX512, WX513,
         WX514, WX515, WX516, WX517, WX518, WX520, WX521, WX522, WX523, WX524,
         WX525, WX526, WX527, WX528, WX529, WX530, WX531, WX532, WX533, WX534,
         WX535, WX536, WX537, WX538, WX539, WX540, WX541, WX542, WX543, WX544,
         WX545, WX546, WX547, WX644, WX645, n3529, WX646, WX647, n3527, WX648,
         WX649, n3525, WX650, WX652, WX653, n3521, WX654, WX655, n3519, WX656,
         WX657, n3517, WX658, WX659, n3515, WX660, WX661, n3513, WX662, WX663,
         n3511, WX664, WX665, n3509, WX666, WX667, n3507, WX668, WX669, n3505,
         WX670, WX671, n3503, WX672, WX673, n3501, WX674, WX675, n3499, WX676,
         WX677, n3497, WX678, WX679, n3495, WX680, WX681, n3493, WX682, WX683,
         n3491, WX684, WX685, n3489, WX686, WX688, WX689, n3485, WX690, WX691,
         n3483, WX692, WX693, n3481, WX694, WX695, n3479, WX696, WX697, n3477,
         WX698, WX699, n3475, WX700, WX701, n3473, WX702, WX703, n3471, WX704,
         WX705, n3469, WX706, WX707, n3467, WX708, WX709, WX710, WX711, WX712,
         WX713, WX714, WX715, WX716, WX717, WX718, WX719, WX720, WX721, WX722,
         WX724, WX725, WX726, WX727, WX728, WX729, WX730, WX731, WX732, WX733,
         WX734, WX735, WX736, WX737, WX738, WX739, WX740, WX741, WX742, WX743,
         WX744, WX745, WX746, WX747, WX748, WX749, WX750, WX751, WX752, WX753,
         WX754, WX755, WX756, WX757, WX758, WX760, WX761, WX762, WX763, WX764,
         WX765, WX766, WX767, WX768, WX769, WX770, WX771, WX772, WX773, WX774,
         WX775, WX776, WX777, WX778, WX779, WX780, WX781, WX782, WX783, WX784,
         WX785, WX786, WX787, WX788, WX789, WX790, WX791, WX792, WX793, WX794,
         WX796, WX797, WX798, WX799, WX800, WX801, WX802, WX803, WX804, WX805,
         WX806, WX807, WX808, WX809, WX810, WX811, WX812, WX813, WX814, WX815,
         WX816, WX817, WX818, WX819, WX820, WX821, WX822, WX823, WX824, WX825,
         WX826, WX827, WX828, WX829, WX830, WX832, WX833, WX834, WX835, WX836,
         WX837, WX838, WX839, WX840, WX841, WX842, WX843, WX844, WX845, WX846,
         WX847, WX848, WX849, WX850, WX851, WX852, WX853, WX854, WX855, WX856,
         WX857, WX858, WX859, WX860, WX861, WX862, WX863, WX864, WX865, WX866,
         WX868, WX869, WX870, WX871, WX872, WX873, WX874, WX875, WX876, WX877,
         WX878, WX879, WX880, WX881, WX882, WX883, WX884, WX885, WX886, WX887,
         WX888, WX889, WX890, WX891, WX892, WX893, WX894, WX895, WX896, WX897,
         WX898, WX899, WX1264, DFF_160_n1, WX1266, WX1268, DFF_162_n1, WX1270,
         WX1272, DFF_164_n1, WX1274, DFF_165_n1, WX1276, DFF_166_n1, WX1278,
         DFF_167_n1, WX1280, DFF_168_n1, WX1282, DFF_169_n1, WX1284, WX1286,
         DFF_171_n1, WX1288, DFF_172_n1, WX1290, DFF_173_n1, WX1292,
         DFF_174_n1, WX1294, DFF_175_n1, WX1296, DFF_176_n1, WX1298,
         DFF_177_n1, WX1300, DFF_178_n1, WX1302, WX1304, DFF_180_n1, WX1306,
         DFF_181_n1, WX1308, DFF_182_n1, WX1310, DFF_183_n1, WX1312,
         DFF_184_n1, WX1314, DFF_185_n1, WX1316, DFF_186_n1, WX1318,
         DFF_187_n1, WX1320, DFF_188_n1, WX1322, DFF_189_n1, WX1324,
         DFF_190_n1, WX1326, DFF_191_n1, WX1778, n8702, n8701, n8700, n8699,
         n8696, n8695, n8694, n8693, n8692, n8691, n8690, n8689, n8688, n8687,
         n8686, n8685, n8684, n8683, n8682, n8681, n8680, n8677, n8676, n8675,
         n8674, n8673, n8672, n8671, WX1839, n8670, WX1937, n8669, WX1939,
         n8668, WX1941, n8667, WX1943, n8666, WX1945, n8665, WX1947, n8664,
         WX1949, n8663, WX1951, n8662, WX1953, n8661, WX1955, WX1957, n8658,
         WX1959, n8657, WX1961, n8656, WX1963, n8655, WX1965, n8654, WX1967,
         n8653, WX1969, WX1970, WX1971, WX1972, WX1973, WX1974, WX1975, WX1976,
         WX1977, WX1978, WX1979, WX1980, WX1981, WX1982, WX1983, WX1984,
         WX1985, WX1986, WX1987, WX1988, WX1989, WX1990, WX1991, WX1993,
         WX1994, WX1995, WX1996, WX1997, WX1998, WX1999, WX2000, WX2001,
         WX2002, WX2003, WX2004, WX2005, WX2006, WX2008, WX2009, WX2010,
         WX2011, WX2012, WX2013, WX2014, WX2015, WX2016, WX2017, WX2018,
         WX2019, WX2020, WX2021, WX2022, WX2023, WX2024, WX2025, WX2026,
         WX2029, WX2030, WX2031, WX2032, WX2033, WX2034, n3785, WX2035, WX2036,
         n3783, WX2037, WX2038, n3781, WX2039, WX2040, n3779, WX2041, WX2042,
         WX2043, WX2044, n3775, WX2045, WX2046, n3773, WX2047, WX2048, n3771,
         WX2049, WX2050, n3769, WX2051, WX2052, n3767, WX2053, WX2054, n3765,
         WX2055, WX2056, n3763, WX2057, WX2058, n3761, WX2059, WX2060, n3759,
         WX2061, WX2062, n3757, WX2063, WX2065, WX2066, WX2067, WX2068, WX2069,
         WX2070, WX2071, WX2072, WX2073, WX2074, WX2075, WX2076, WX2077,
         WX2078, WX2079, WX2080, WX2081, WX2082, WX2083, WX2084, WX2085,
         WX2086, WX2087, WX2088, WX2089, WX2090, WX2091, WX2092, WX2093,
         WX2094, WX2095, WX2096, WX2097, WX2098, WX2099, WX2101, WX2102,
         WX2103, WX2104, WX2105, WX2106, WX2107, WX2108, WX2109, WX2110,
         WX2111, WX2112, WX2113, WX2114, WX2115, WX2116, WX2117, WX2118,
         WX2119, WX2120, WX2121, WX2122, WX2123, WX2124, WX2125, WX2126,
         WX2127, WX2128, WX2129, WX2130, WX2131, WX2132, WX2133, WX2134,
         WX2135, WX2137, WX2138, WX2139, WX2140, WX2141, WX2142, WX2143,
         WX2144, WX2145, WX2146, WX2147, WX2148, WX2149, WX2150, WX2151,
         WX2152, WX2153, WX2154, WX2155, WX2156, WX2157, WX2158, WX2159,
         WX2160, WX2161, WX2162, WX2163, WX2164, WX2165, WX2166, WX2167,
         WX2168, WX2169, WX2170, WX2171, WX2173, WX2174, WX2175, WX2176,
         WX2177, WX2178, WX2179, WX2180, WX2181, WX2182, WX2183, WX2184,
         WX2185, WX2186, WX2187, WX2188, WX2189, WX2190, WX2191, WX2192,
         WX2557, DFF_352_n1, WX2559, DFF_353_n1, WX2561, DFF_354_n1, WX2563,
         WX2565, DFF_356_n1, WX2567, DFF_357_n1, WX2569, DFF_358_n1, WX2571,
         WX2573, DFF_360_n1, WX2575, WX2577, WX2579, DFF_363_n1, WX2581,
         DFF_364_n1, WX2583, DFF_365_n1, WX2585, DFF_366_n1, WX2587, WX2589,
         DFF_368_n1, WX2591, DFF_369_n1, WX2593, DFF_370_n1, WX2595,
         DFF_371_n1, WX2597, DFF_372_n1, WX2599, DFF_373_n1, WX2601,
         DFF_374_n1, WX2603, DFF_375_n1, WX2605, DFF_376_n1, WX2607, WX2609,
         DFF_378_n1, WX2611, WX2613, DFF_380_n1, WX2615, DFF_381_n1, WX2617,
         DFF_382_n1, WX2619, DFF_383_n1, WX3071, n8644, n8643, n8642, n8641,
         n8640, n8639, n8638, n8637, n8636, n8635, n8632, n8631, n8630, n8629,
         n8628, n8627, n8626, n8625, n8624, n8623, n8622, n8621, n8620, n8619,
         n8618, n8617, n8616, n8613, WX3132, n8612, WX3230, n8611, WX3232,
         n8610, WX3234, n8609, WX3236, n8608, WX3238, n8607, WX3240, n8606,
         WX3242, n8605, WX3244, n8604, WX3246, n8603, WX3248, n8602, WX3250,
         n8601, WX3252, n8600, WX3254, n8599, WX3256, n8598, WX3258, n8597,
         WX3260, WX3262, WX3263, WX3264, WX3265, WX3266, WX3267, WX3268,
         WX3269, WX3270, WX3271, WX3272, WX3273, WX3274, WX3275, WX3276,
         WX3277, WX3278, WX3279, WX3280, WX3281, WX3282, WX3283, WX3284,
         WX3285, WX3286, WX3287, WX3288, WX3289, WX3290, WX3291, WX3292,
         WX3293, WX3295, WX3299, WX3301, WX3303, WX3305, WX3307, WX3309,
         WX3311, WX3313, WX3315, WX3317, WX3319, WX3321, WX3323, WX3325,
         WX3326, WX3327, WX3328, WX3329, WX3330, WX3331, n3749, WX3332, WX3334,
         WX3335, WX3336, WX3337, n3743, WX3338, WX3339, n3741, WX3340, WX3341,
         n3739, WX3342, WX3343, n3737, WX3344, WX3345, n3735, WX3346, WX3347,
         n3733, WX3348, WX3349, WX3350, WX3351, n3729, WX3352, WX3353, n3727,
         WX3354, WX3355, n3725, WX3356, WX3357, WX3358, WX3359, WX3360, WX3361,
         WX3362, WX3363, WX3364, WX3365, WX3366, WX3367, WX3368, WX3370,
         WX3371, WX3372, WX3373, WX3374, WX3375, WX3376, WX3377, WX3378,
         WX3379, WX3380, WX3381, WX3382, WX3383, WX3384, WX3385, WX3386,
         WX3387, WX3388, WX3389, WX3390, WX3391, WX3392, WX3393, WX3394,
         WX3395, WX3396, WX3397, WX3398, WX3399, WX3400, WX3401, WX3402,
         WX3403, WX3404, WX3406, WX3407, WX3408, WX3409, WX3410, WX3411,
         WX3412, WX3413, WX3414, WX3415, WX3416, WX3417, WX3418, WX3419,
         WX3420, WX3421, WX3422, WX3423, WX3424, WX3425, WX3426, WX3427,
         WX3428, WX3429, WX3430, WX3431, WX3432, WX3433, WX3434, WX3435,
         WX3436, WX3437, WX3438, WX3440, WX3441, WX3442, WX3443, WX3444,
         WX3445, WX3446, WX3447, WX3448, WX3449, WX3450, WX3451, WX3452,
         WX3453, WX3454, WX3455, WX3456, WX3457, WX3458, WX3459, WX3460,
         WX3461, WX3462, WX3463, WX3464, WX3465, WX3466, WX3467, WX3468,
         WX3469, WX3470, WX3471, WX3472, WX3474, WX3475, WX3476, WX3477,
         WX3478, WX3479, WX3480, WX3481, WX3482, WX3483, WX3484, WX3485,
         WX3850, DFF_544_n1, WX3852, DFF_545_n1, WX3854, DFF_546_n1, WX3856,
         WX3858, DFF_548_n1, WX3860, WX3862, DFF_550_n1, WX3864, DFF_551_n1,
         WX3866, DFF_552_n1, WX3868, DFF_553_n1, WX3870, WX3872, DFF_555_n1,
         WX3874, DFF_556_n1, WX3876, DFF_557_n1, WX3878, DFF_558_n1, WX3880,
         WX3882, DFF_560_n1, WX3884, DFF_561_n1, WX3886, DFF_562_n1, WX3888,
         DFF_563_n1, WX3890, DFF_564_n1, WX3892, DFF_565_n1, WX3894, WX3896,
         DFF_567_n1, WX3898, DFF_568_n1, WX3900, DFF_569_n1, WX3902,
         DFF_570_n1, WX3904, WX3906, DFF_572_n1, WX3908, DFF_573_n1, WX3910,
         DFF_574_n1, WX3912, DFF_575_n1, WX4364, n8586, n8585, n8584, n8583,
         n8582, n8581, n8580, n8579, n8578, n8577, n8576, n8573, n8572, n8571,
         n8570, n8569, n8568, n8567, n8566, n8565, n8564, n8563, n8562, n8561,
         n8560, n8559, n8558, n8555, WX4425, n8554, WX4523, n8553, WX4525,
         n8552, WX4527, n8551, WX4529, n8550, WX4531, n8549, WX4533, n8548,
         WX4535, n8547, WX4537, n8546, WX4539, n8545, WX4541, n8544, WX4543,
         n8543, WX4545, n8542, WX4547, n8541, WX4549, n8540, WX4551, WX4553,
         n8537, WX4555, WX4556, WX4557, WX4558, WX4559, WX4560, WX4561, WX4562,
         WX4563, WX4564, WX4565, WX4566, WX4567, WX4568, WX4569, WX4570,
         WX4571, WX4572, WX4573, WX4574, WX4575, WX4576, WX4577, WX4578,
         WX4579, WX4580, WX4581, WX4582, WX4583, WX4584, WX4585, WX4588,
         WX4590, WX4592, WX4594, WX4596, WX4598, WX4600, WX4602, WX4604,
         WX4606, WX4608, WX4610, WX4612, WX4614, WX4616, WX4618, WX4619,
         WX4621, WX4622, WX4623, WX4624, n3717, WX4625, WX4626, WX4627, WX4628,
         n3713, WX4629, WX4630, WX4631, WX4632, WX4633, WX4634, n3707, WX4635,
         WX4636, n3705, WX4637, WX4638, n3703, WX4639, WX4640, n3701, WX4641,
         WX4642, WX4643, WX4644, n3697, WX4645, WX4646, n3695, WX4647, WX4648,
         n3693, WX4649, WX4650, n3691, WX4651, WX4652, WX4653, WX4655, WX4656,
         WX4657, WX4658, WX4659, WX4660, WX4661, WX4662, WX4663, WX4664,
         WX4665, WX4666, WX4667, WX4668, WX4669, WX4670, WX4671, WX4672,
         WX4673, WX4674, WX4675, WX4676, WX4677, WX4678, WX4679, WX4680,
         WX4681, WX4682, WX4683, WX4684, WX4685, WX4686, WX4687, WX4689,
         WX4690, WX4691, WX4692, WX4693, WX4694, WX4695, WX4696, WX4697,
         WX4698, WX4699, WX4700, WX4701, WX4702, WX4703, WX4704, WX4705,
         WX4706, WX4707, WX4708, WX4709, WX4710, WX4711, WX4712, WX4713,
         WX4714, WX4715, WX4716, WX4717, WX4718, WX4719, WX4720, WX4721,
         WX4723, WX4724, WX4725, WX4726, WX4727, WX4728, WX4729, WX4730,
         WX4731, WX4732, WX4733, WX4734, WX4735, WX4736, WX4737, WX4738,
         WX4739, WX4740, WX4741, WX4742, WX4743, WX4744, WX4745, WX4746,
         WX4747, WX4748, WX4749, WX4750, WX4751, WX4752, WX4753, WX4754,
         WX4755, WX4757, WX4758, WX4759, WX4760, WX4761, WX4762, WX4763,
         WX4764, WX4765, WX4766, WX4767, WX4768, WX4769, WX4770, WX4771,
         WX4772, WX4773, WX4774, WX4775, WX4776, WX4777, WX4778, WX5143,
         DFF_736_n1, WX5145, DFF_737_n1, WX5147, DFF_738_n1, WX5149, WX5151,
         DFF_740_n1, WX5153, WX5155, DFF_742_n1, WX5157, DFF_743_n1, WX5159,
         DFF_744_n1, WX5161, DFF_745_n1, WX5163, DFF_746_n1, WX5165,
         DFF_747_n1, WX5167, DFF_748_n1, WX5169, DFF_749_n1, WX5171,
         DFF_750_n1, WX5173, WX5175, DFF_752_n1, WX5177, DFF_753_n1, WX5179,
         DFF_754_n1, WX5181, DFF_755_n1, WX5183, DFF_756_n1, WX5185,
         DFF_757_n1, WX5187, WX5189, DFF_759_n1, WX5191, DFF_760_n1, WX5193,
         DFF_761_n1, WX5195, DFF_762_n1, WX5197, WX5199, DFF_764_n1, WX5201,
         DFF_765_n1, WX5203, DFF_766_n1, WX5205, DFF_767_n1, WX5657, n8528,
         n8527, n8526, n8525, n8524, n8523, n8520, n8519, n8518, n8517, n8516,
         n8515, n8514, n8513, n8512, n8511, n8510, n8509, n8508, n8507, n8506,
         n8505, n8502, n8501, n8500, n8499, n8498, n8497, WX5718, n8496,
         WX5816, n8495, WX5818, n8494, WX5820, n8493, WX5822, n8492, WX5824,
         n8491, WX5826, n8490, WX5828, n8489, WX5830, n8488, WX5832, n8487,
         WX5834, WX5836, n8484, WX5838, n8483, WX5840, n8482, WX5842, n8481,
         WX5844, n8480, WX5846, n8479, WX5848, WX5849, WX5850, WX5851, WX5852,
         WX5853, WX5854, WX5855, WX5856, WX5857, WX5858, WX5859, WX5860,
         WX5861, WX5862, WX5863, WX5864, WX5865, WX5866, WX5867, WX5868,
         WX5870, WX5871, WX5872, WX5873, WX5874, WX5875, WX5876, WX5877,
         WX5878, WX5879, WX5881, WX5883, WX5885, WX5887, WX5889, WX5891,
         WX5893, WX5895, WX5897, WX5899, WX5901, WX5905, WX5907, WX5909,
         WX5911, WX5912, WX5913, WX5914, WX5915, WX5916, WX5917, WX5918,
         WX5919, WX5920, WX5921, WX5922, WX5923, WX5924, WX5925, WX5926,
         WX5927, WX5928, WX5929, WX5930, WX5931, WX5932, WX5933, n3669, WX5934,
         WX5935, WX5936, WX5938, WX5939, n3663, WX5940, WX5941, n3661, WX5942,
         WX5943, WX5944, WX5945, WX5946, WX5947, WX5948, WX5949, WX5950,
         WX5951, WX5952, WX5953, WX5954, WX5955, WX5956, WX5957, WX5958,
         WX5959, WX5960, WX5961, WX5962, WX5963, WX5964, WX5965, WX5966,
         WX5967, WX5968, WX5969, WX5970, WX5972, WX5973, WX5974, WX5975,
         WX5976, WX5977, WX5978, WX5979, WX5980, WX5981, WX5982, WX5983,
         WX5984, WX5985, WX5986, WX5987, WX5988, WX5989, WX5990, WX5991,
         WX5992, WX5993, WX5994, WX5995, WX5996, WX5997, WX5998, WX5999,
         WX6000, WX6001, WX6002, WX6003, WX6004, WX6006, WX6007, WX6008,
         WX6009, WX6010, WX6011, WX6012, WX6013, WX6014, WX6015, WX6016,
         WX6017, WX6018, WX6019, WX6020, WX6021, WX6022, WX6023, WX6024,
         WX6025, WX6026, WX6027, WX6028, WX6029, WX6030, WX6031, WX6032,
         WX6033, WX6034, WX6035, WX6036, WX6037, WX6038, WX6040, WX6041,
         WX6042, WX6043, WX6044, WX6045, WX6046, WX6047, WX6048, WX6049,
         WX6050, WX6051, WX6052, WX6053, WX6054, WX6055, WX6056, WX6057,
         WX6058, WX6059, WX6060, WX6061, WX6062, WX6063, WX6064, WX6065,
         WX6066, WX6067, WX6068, WX6069, WX6070, WX6071, WX6436, WX6438,
         DFF_929_n1, WX6440, DFF_930_n1, WX6442, WX6444, DFF_932_n1, WX6446,
         DFF_933_n1, WX6448, DFF_934_n1, WX6450, DFF_935_n1, WX6452,
         DFF_936_n1, WX6454, DFF_937_n1, WX6456, WX6458, DFF_939_n1, WX6460,
         DFF_940_n1, WX6462, DFF_941_n1, WX6464, DFF_942_n1, WX6466,
         DFF_943_n1, WX6468, DFF_944_n1, WX6470, WX6472, DFF_946_n1, WX6474,
         DFF_947_n1, WX6476, DFF_948_n1, WX6478, DFF_949_n1, WX6480,
         DFF_950_n1, WX6482, DFF_951_n1, WX6484, DFF_952_n1, WX6486,
         DFF_953_n1, WX6488, DFF_954_n1, WX6490, DFF_955_n1, WX6492,
         DFF_956_n1, WX6494, DFF_957_n1, WX6496, DFF_958_n1, WX6498,
         DFF_959_n1, WX6950, n8470, n8467, n8466, n8465, n8464, n8463, n8462,
         n8461, n8460, n8459, n8458, n8457, n8456, n8455, n8454, n8453, n8452,
         n8449, n8448, n8447, n8446, n8445, WX6999, n8444, n8443, n8442, n8441,
         n8440, n8439, WX7011, n8438, WX7109, n8437, WX7111, n8436, WX7113,
         n8435, WX7115, n8434, WX7117, WX7119, n8431, WX7121, n8430, WX7123,
         n8429, WX7125, n8428, WX7127, n8427, WX7129, n8426, WX7131, n8425,
         WX7133, n8424, WX7135, n8423, WX7137, n8422, WX7139, n8421, WX7141,
         WX7142, WX7143, WX7144, WX7145, WX7146, WX7147, WX7148, WX7149,
         WX7150, WX7151, WX7153, WX7154, WX7155, WX7156, WX7157, WX7158,
         WX7159, WX7160, WX7161, WX7162, WX7163, WX7164, WX7165, WX7166,
         WX7167, WX7168, WX7169, WX7170, WX7171, WX7172, WX7174, WX7176,
         WX7178, WX7180, WX7182, WX7184, WX7188, WX7190, WX7192, WX7194,
         WX7196, WX7198, WX7200, WX7202, WX7204, WX7205, WX7206, WX7207,
         WX7208, WX7209, WX7210, WX7211, WX7212, WX7213, WX7214, WX7215,
         WX7216, n3647, WX7217, WX7218, WX7219, WX7221, WX7222, WX7223, WX7224,
         n3639, WX7225, WX7226, WX7227, WX7228, n3635, WX7229, WX7230, WX7231,
         WX7232, WX7233, WX7234, WX7235, WX7236, WX7237, WX7238, WX7239,
         WX7240, WX7241, WX7242, WX7243, WX7244, WX7245, WX7246, WX7247,
         WX7248, WX7249, WX7250, WX7251, WX7252, WX7253, WX7255, WX7256,
         WX7257, WX7258, WX7259, WX7260, WX7261, WX7262, WX7263, WX7264,
         WX7265, WX7266, WX7267, WX7268, WX7269, WX7270, WX7271, WX7272,
         WX7273, WX7274, WX7275, WX7276, WX7277, WX7278, WX7279, WX7280,
         WX7281, WX7282, WX7283, WX7284, WX7285, WX7286, WX7287, WX7289,
         WX7290, WX7291, WX7292, WX7293, WX7294, WX7295, WX7296, WX7297,
         WX7298, WX7299, WX7300, WX7301, WX7302, WX7303, WX7304, WX7305,
         WX7306, WX7307, WX7308, WX7309, WX7310, WX7311, WX7312, WX7313,
         WX7314, WX7315, WX7316, WX7317, WX7318, WX7319, WX7320, WX7321,
         WX7323, WX7324, WX7325, WX7326, WX7327, WX7328, WX7329, WX7330,
         WX7331, WX7332, WX7333, WX7334, WX7335, WX7336, WX7337, WX7338,
         WX7339, WX7340, WX7341, WX7342, WX7343, WX7344, WX7345, WX7346,
         WX7347, WX7348, WX7349, WX7350, WX7351, WX7352, WX7353, WX7354,
         WX7355, WX7357, WX7358, WX7359, WX7360, WX7361, WX7362, WX7363,
         WX7364, WX7729, DFF_1120_n1, WX7731, DFF_1121_n1, WX7733, DFF_1122_n1,
         WX7735, DFF_1123_n1, WX7737, DFF_1124_n1, WX7739, DFF_1125_n1, WX7741,
         DFF_1126_n1, WX7743, DFF_1127_n1, WX7745, DFF_1128_n1, WX7747,
         DFF_1129_n1, WX7749, WX7751, DFF_1131_n1, WX7753, WX7755, DFF_1133_n1,
         WX7757, DFF_1134_n1, WX7759, WX7761, DFF_1136_n1, WX7763, DFF_1137_n1,
         WX7765, DFF_1138_n1, WX7767, DFF_1139_n1, WX7769, WX7771, DFF_1141_n1,
         WX7773, DFF_1142_n1, WX7775, DFF_1143_n1, WX7777, DFF_1144_n1, WX7779,
         DFF_1145_n1, WX7781, DFF_1146_n1, WX7783, DFF_1147_n1, WX7785,
         DFF_1148_n1, WX7787, WX7789, DFF_1150_n1, WX7791, DFF_1151_n1, WX8243,
         n8411, n8410, n8409, n8408, n8407, n8406, n8405, n8404, n8403, n8402,
         n8401, WX8266, n8400, n8399, n8396, n8395, n8394, n8393, n8392, n8391,
         n8390, n8389, n8388, n8387, n8386, n8385, n8384, n8383, n8382, n8381,
         WX8304, WX8402, n8378, WX8404, n8377, WX8406, n8376, WX8408, n8375,
         WX8410, n8374, WX8412, n8373, WX8414, n8372, WX8416, n8371, WX8418,
         n8370, WX8420, n8369, WX8422, n8368, WX8424, n8367, WX8426, n8366,
         WX8428, n8365, WX8430, n8364, WX8432, n8363, WX8434, WX8436, WX8437,
         WX8438, WX8439, WX8440, WX8441, WX8442, WX8443, WX8444, WX8445,
         WX8446, WX8447, WX8448, WX8449, WX8450, WX8451, WX8452, WX8453,
         WX8454, WX8455, WX8456, WX8457, WX8458, WX8459, WX8460, WX8461,
         WX8462, WX8463, WX8464, WX8465, WX8467, WX8471, WX8473, WX8475,
         WX8477, WX8479, WX8481, WX8483, WX8485, WX8487, WX8489, WX8491,
         WX8493, WX8495, WX8497, WX8498, WX8499, n3625, WX8500, WX8501, WX8502,
         WX8504, WX8505, WX8506, WX8507, n3617, WX8508, WX8509, WX8510, WX8511,
         n3613, WX8512, WX8513, WX8514, WX8515, WX8516, WX8517, WX8518, WX8519,
         WX8520, WX8521, WX8522, WX8523, WX8524, WX8525, WX8526, WX8527,
         WX8528, WX8529, WX8530, WX8531, WX8532, WX8533, WX8534, WX8535,
         WX8536, WX8538, WX8539, WX8540, WX8541, WX8542, WX8543, WX8544,
         WX8545, WX8546, WX8547, WX8548, WX8549, WX8550, WX8551, WX8552,
         WX8553, WX8554, WX8555, WX8556, WX8557, WX8558, WX8559, WX8560,
         WX8561, WX8562, WX8563, WX8564, WX8565, WX8566, WX8567, WX8568,
         WX8569, WX8570, WX8572, WX8573, WX8574, WX8575, WX8576, WX8577,
         WX8578, WX8579, WX8580, WX8581, WX8582, WX8583, WX8584, WX8585,
         WX8586, WX8587, WX8588, WX8589, WX8590, WX8591, WX8592, WX8593,
         WX8594, WX8595, WX8596, WX8597, WX8598, WX8599, WX8600, WX8601,
         WX8602, WX8603, WX8604, WX8606, WX8607, WX8608, WX8609, WX8610,
         WX8611, WX8612, WX8613, WX8614, WX8615, WX8616, WX8617, WX8618,
         WX8619, WX8620, WX8621, WX8622, WX8623, WX8624, WX8625, WX8626,
         WX8627, WX8628, WX8629, WX8630, WX8631, WX8632, WX8633, WX8634,
         WX8635, WX8636, WX8637, WX8638, WX8640, WX8641, WX8642, WX8643,
         WX8644, WX8645, WX8646, WX8647, WX8648, WX8649, WX8650, WX8651,
         WX8652, WX8653, WX8654, WX8655, WX8656, WX8657, WX9022, DFF_1312_n1,
         WX9024, DFF_1313_n1, WX9026, DFF_1314_n1, WX9028, WX9030, DFF_1316_n1,
         WX9032, DFF_1317_n1, WX9034, DFF_1318_n1, WX9036, WX9038, WX9040,
         DFF_1321_n1, WX9042, WX9044, DFF_1323_n1, WX9046, DFF_1324_n1, WX9048,
         DFF_1325_n1, WX9050, DFF_1326_n1, WX9052, WX9054, DFF_1328_n1, WX9056,
         DFF_1329_n1, WX9058, DFF_1330_n1, WX9060, DFF_1331_n1, WX9062,
         DFF_1332_n1, WX9064, DFF_1333_n1, WX9066, DFF_1334_n1, WX9068,
         DFF_1335_n1, WX9070, WX9072, WX9074, DFF_1338_n1, WX9076, DFF_1339_n1,
         WX9078, DFF_1340_n1, WX9080, DFF_1341_n1, WX9082, DFF_1342_n1, WX9084,
         DFF_1343_n1, WX9536, n8353, n8352, n8351, n8350, n8349, n8348, n8347,
         n8346, n8343, n8342, n8341, n8340, n8339, n8338, n8337, n8336, n8335,
         n8334, n8333, n8332, n8331, n8330, n8329, n8328, n8325, n8324, n8323,
         n8322, WX9597, n8321, WX9695, n8320, WX9697, n8319, WX9699, n8318,
         WX9701, n8317, WX9703, n8316, WX9705, n8315, WX9707, n8314, WX9709,
         n8313, WX9711, n8312, WX9713, n8311, WX9715, n8310, WX9717, WX9719,
         n8307, WX9721, n8306, WX9723, n8305, WX9725, n8304, WX9727, WX9728,
         WX9729, WX9730, WX9731, WX9732, WX9733, WX9734, WX9735, WX9736,
         WX9737, WX9738, WX9739, WX9740, WX9741, WX9742, WX9743, WX9744,
         WX9745, WX9746, WX9747, WX9748, WX9749, WX9750, WX9751, WX9753,
         WX9754, WX9755, WX9756, WX9757, WX9758, WX9760, WX9762, WX9764,
         WX9766, WX9768, WX9770, WX9772, WX9774, WX9776, WX9778, WX9780,
         WX9782, WX9784, WX9788, WX9790, WX9791, WX9792, WX9793, WX9794, n3591,
         WX9795, WX9796, WX9797, WX9798, WX9799, WX9800, WX9801, WX9802,
         WX9803, WX9804, WX9805, WX9806, WX9807, WX9808, WX9809, WX9810,
         WX9811, WX9812, WX9813, WX9814, WX9815, WX9816, n3569, WX9817, WX9818,
         WX9819, WX9821, WX9822, WX9823, WX9824, WX9825, WX9826, WX9827,
         WX9828, WX9829, WX9830, WX9831, WX9832, WX9833, WX9834, WX9835,
         WX9836, WX9837, WX9838, WX9839, WX9840, WX9841, WX9842, WX9843,
         WX9844, WX9845, WX9846, WX9847, WX9848, WX9849, WX9850, WX9851,
         WX9852, WX9853, WX9855, WX9856, WX9857, WX9858, WX9859, WX9860,
         WX9861, WX9862, WX9863, WX9864, WX9865, WX9866, WX9867, WX9868,
         WX9869, WX9870, WX9871, WX9872, WX9873, WX9874, WX9875, WX9876,
         WX9877, WX9878, WX9879, WX9880, WX9881, WX9882, WX9883, WX9884,
         WX9885, WX9886, WX9887, WX9889, WX9890, WX9891, WX9892, WX9893,
         WX9894, WX9895, WX9896, WX9897, WX9898, WX9899, WX9900, WX9901,
         WX9902, WX9903, WX9904, WX9905, WX9906, WX9907, WX9908, WX9909,
         WX9910, WX9911, WX9912, WX9913, WX9914, WX9915, WX9916, WX9917,
         WX9918, WX9919, WX9920, WX9921, WX9923, WX9924, WX9925, WX9926,
         WX9927, WX9928, WX9929, WX9930, WX9931, WX9932, WX9933, WX9934,
         WX9935, WX9936, WX9937, WX9938, WX9939, WX9940, WX9941, WX9942,
         WX9943, WX9944, WX9945, WX9946, WX9947, WX9948, WX9949, WX9950,
         WX10315, DFF_1504_n1, WX10317, DFF_1505_n1, WX10319, WX10321, WX10323,
         DFF_1508_n1, WX10325, DFF_1509_n1, WX10327, DFF_1510_n1, WX10329,
         DFF_1511_n1, WX10331, DFF_1512_n1, WX10333, DFF_1513_n1, WX10335,
         WX10337, DFF_1515_n1, WX10339, DFF_1516_n1, WX10341, WX10343,
         DFF_1518_n1, WX10345, WX10347, DFF_1520_n1, WX10349, DFF_1521_n1,
         WX10351, DFF_1522_n1, WX10353, WX10355, DFF_1524_n1, WX10357,
         DFF_1525_n1, WX10359, DFF_1526_n1, WX10361, DFF_1527_n1, WX10363,
         DFF_1528_n1, WX10365, DFF_1529_n1, WX10367, DFF_1530_n1, WX10369,
         DFF_1531_n1, WX10371, DFF_1532_n1, WX10373, DFF_1533_n1, WX10375,
         WX10377, DFF_1535_n1, WX10829, n8295, n8294, n8293, n8290, n8289,
         n8288, n8287, n8286, n8285, n8284, n8283, n8282, n8281, n8280, n8279,
         n8278, n8277, n8276, n8275, n8272, n8271, n8270, n8269, n8268, n8267,
         n8266, n8265, n8264, WX10890, n8263, WX10988, n8262, WX10990, n8261,
         WX10992, n8260, WX10994, n8259, WX10996, n8258, WX10998, n8257,
         WX11000, WX11002, n8254, WX11004, n8253, WX11006, n8252, WX11008,
         n8251, WX11010, n8250, WX11012, n8249, WX11014, n8248, WX11016, n8247,
         WX11018, n8246, WX11020, WX11021, WX11022, WX11023, WX11024, WX11025,
         WX11026, WX11027, WX11028, WX11029, WX11030, WX11031, WX11032,
         WX11033, WX11034, WX11036, WX11037, WX11038, WX11039, WX11040,
         WX11041, WX11042, WX11043, WX11044, WX11045, WX11046, WX11047,
         WX11048, WX11049, WX11050, WX11051, WX11052, WX11053, WX11054,
         WX11055, WX11056, WX11057, WX11058, WX11059, WX11060, WX11061,
         WX11062, WX11063, WX11064, WX11065, WX11066, WX11067, WX11070,
         WX11071, WX11073, WX11074, WX11075, WX11077, WX11078, WX11079,
         WX11080, WX11081, WX11082, WX11083, WX11084, WX11085, WX11086,
         WX11087, WX11088, WX11089, WX11090, WX11091, WX11092, WX11093,
         WX11094, WX11095, WX11096, WX11097, WX11098, WX11099, n3547, WX11100,
         WX11101, WX11102, WX11104, WX11105, WX11106, WX11107, n3539, WX11108,
         WX11109, WX11110, WX11111, n3535, WX11112, WX11113, WX11114, WX11115,
         WX11116, WX11117, WX11118, WX11119, WX11120, WX11121, WX11122,
         WX11123, WX11124, WX11125, WX11126, WX11127, WX11128, WX11129,
         WX11130, WX11131, WX11132, WX11133, WX11134, WX11135, WX11136,
         WX11138, WX11139, WX11140, WX11141, WX11142, WX11143, WX11144,
         WX11145, WX11146, WX11147, WX11148, WX11149, WX11150, WX11151,
         WX11152, WX11153, WX11154, WX11155, WX11156, WX11157, WX11158,
         WX11159, WX11160, WX11161, WX11162, WX11163, WX11164, WX11165,
         WX11166, WX11167, WX11168, WX11169, WX11170, WX11172, WX11173,
         WX11174, WX11175, WX11176, WX11177, WX11178, WX11179, WX11180,
         WX11181, WX11182, WX11183, WX11184, WX11185, WX11186, WX11187,
         WX11188, WX11189, WX11190, WX11191, WX11192, WX11193, WX11194,
         WX11195, WX11196, WX11197, WX11198, WX11199, WX11200, WX11201,
         WX11202, WX11203, WX11204, WX11206, WX11207, WX11208, WX11209,
         WX11210, WX11211, WX11212, WX11213, WX11214, WX11215, WX11216,
         WX11217, WX11218, WX11219, WX11220, WX11221, WX11222, WX11223,
         WX11224, WX11225, WX11226, WX11227, WX11228, WX11229, WX11230,
         WX11231, WX11232, WX11233, WX11234, WX11235, WX11236, WX11237,
         WX11238, WX11240, WX11241, WX11242, WX11243, WX11608, DFF_1696_n1,
         WX11610, WX11612, DFF_1698_n1, WX11614, DFF_1699_n1, WX11616,
         DFF_1700_n1, WX11618, DFF_1701_n1, WX11620, DFF_1702_n1, WX11622,
         DFF_1703_n1, WX11624, DFF_1704_n1, WX11626, DFF_1705_n1, WX11628,
         DFF_1706_n1, WX11630, DFF_1707_n1, WX11632, DFF_1708_n1, WX11634,
         DFF_1709_n1, WX11636, WX11638, DFF_1711_n1, WX11640, DFF_1712_n1,
         WX11642, DFF_1713_n1, WX11644, WX11646, DFF_1715_n1, WX11648,
         DFF_1716_n1, WX11650, DFF_1717_n1, WX11652, DFF_1718_n1, WX11654,
         DFF_1719_n1, WX11656, DFF_1720_n1, WX11658, DFF_1721_n1, WX11660,
         DFF_1722_n1, WX11662, DFF_1723_n1, WX11664, DFF_1724_n1, WX11666,
         DFF_1725_n1, WX11668, DFF_1726_n1, WX11670, n2245, n2153, n3278,
         n2152, n2148, Tj_Trigger, Tj_OUT1, Tj_OUT2, Tj_OUT3, Tj_OUT4,
         Tj_OUT1234, Tj_OUT5, Tj_OUT6, Tj_OUT7, Tj_OUT8, Tj_OUT5678,
         test_se_NOT, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n67, n77, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n619, n621,
         n623, n658, n3061, n3063, n3064, n3066, n3068, n3070, n3072, n3074,
         n3076, n3078, n3080, n3082, n3083, n3085, n3086, n3088, n3089, n3091,
         n3092, n3094, n3096, n3098, n3100, n3102, n3103, n3105, n3106, n3108,
         n3109, n3111, n3113, n3115, n3117, n3119, n3121, n3123, n3125, n3127,
         n3129, n3131, n3133, n3135, n3137, n3139, n3141, n3143, n3145, n3147,
         n3149, n3150, n3152, n3153, n3155, n3156, n3158, n3160, n3162, n3164,
         n3166, n3167, n3169, n3170, n3172, n3173, n3175, n3176, n3178, n3180,
         n3182, n3183, n3185, n3186, n3188, n3189, n3191, n3192, n3194, n3196,
         n3198, n3200, n3202, n3204, n3206, n3208, n3210, n3211, n3213, n3215,
         n3217, n3219, n3221, n3223, n3225, n3227, n3229, n3231, n3232, n3234,
         n3235, n3236, n3238, n3240, n3242, n3244, n3246, n3248, n3249, n3251,
         n3253, n3254, n3256, n3258, n3260, n3261, n3263, n3265, n3266, n3268,
         n3270, n3272, n3273, n3275, n3277, n3280, n3282, n3284, n3285, n3287,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3468,
         n3470, n3472, n3474, n3476, n3478, n3480, n3482, n3484, n3486, n3487,
         n3488, n3490, n3492, n3494, n3496, n3498, n3500, n3502, n3504, n3506,
         n3508, n3510, n3512, n3514, n3516, n3518, n3520, n3522, n3523, n3524,
         n3526, n3528, n3530, n3532, n3534, n3536, n3538, n3540, n3542, n3543,
         n3544, n3546, n3548, n3550, n3552, n3554, n3556, n3558, n3560, n3562,
         n3564, n3565, n3566, n3568, n3570, n3572, n3574, n3576, n3578, n3580,
         n3582, n3584, n3586, n3588, n3590, n3592, n3594, n3596, n3598, n3600,
         n3602, n3604, n3606, n3608, n3610, n3612, n3614, n3616, n3618, n3620,
         n3621, n3622, n3624, n3626, n3628, n3630, n3632, n3634, n3636, n3638,
         n3640, n3642, n3643, n3644, n3646, n3648, n3650, n3652, n3654, n3656,
         n3658, n3660, n3662, n3664, n3665, n3666, n3668, n3670, n3672, n3674,
         n3676, n3678, n3680, n3682, n3684, n3686, n3688, n3690, n3692, n3694,
         n3696, n3698, n3700, n3702, n3704, n3706, n3708, n3710, n3712, n3714,
         n3716, n3718, n3720, n3721, n3722, n3724, n3726, n3728, n3730, n3732,
         n3734, n3736, n3738, n3740, n3742, n3744, n3746, n3747, n3748, n3750,
         n3752, n3754, n3755, n3756, n3758, n3760, n3762, n3764, n3766, n3768,
         n3770, n3772, n3774, n3776, n3778, n3780, n3782, n3784, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3831, n3832, n3833, n3834, n3836, n3837, n3838, n3839, n3840,
         n3841, n3843, n3844, n3846, n3847, n3849, n3850, n3852, n3853, n3855,
         n3856, n3857, n3859, n3861, n3862, n3863, n3864, n3866, n3867, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         U3558_n1, U3871_n1, U3991_n1, U5716_n1, U5717_n1, U5718_n1, U5719_n1,
         U5720_n1, U5721_n1, U5722_n1, U5723_n1, U5724_n1, U5725_n1, U5726_n1,
         U5727_n1, U5728_n1, U5729_n1, U5730_n1, U5731_n1, U5732_n1, U5733_n1,
         U5734_n1, U5735_n1, U5736_n1, U5737_n1, U5738_n1, U5739_n1, U5740_n1,
         U5741_n1, U5742_n1, U5743_n1, U5744_n1, U5745_n1, U5746_n1, U5747_n1,
         U5748_n1, U5749_n1, U5750_n1, U5751_n1, U5752_n1, U5753_n1, U5754_n1,
         U5755_n1, U5756_n1, U5757_n1, U5758_n1, U5759_n1, U5760_n1, U5761_n1,
         U5762_n1, U5763_n1, U5764_n1, U5765_n1, U5766_n1, U5767_n1, U5768_n1,
         U5769_n1, U5770_n1, U5771_n1, U5772_n1, U5773_n1, U5774_n1, U5775_n1,
         U5776_n1, U5777_n1, U5778_n1, U5779_n1, U5780_n1, U5781_n1, U5782_n1,
         U5783_n1, U5784_n1, U5785_n1, U5786_n1, U5787_n1, U5788_n1, U5789_n1,
         U5790_n1, U5791_n1, U5792_n1, U5793_n1, U5794_n1, U5795_n1, U5796_n1,
         U5797_n1, U5798_n1, U5799_n1, U5800_n1, U5801_n1, U5802_n1, U5803_n1,
         U5804_n1, U5805_n1, U5806_n1, U5807_n1, U5808_n1, U5809_n1, U5810_n1,
         U5811_n1, U5812_n1, U5813_n1, U5814_n1, U5815_n1, U5816_n1, U5817_n1,
         U5818_n1, U5819_n1, U5820_n1, U5821_n1, U5822_n1, U5823_n1, U5824_n1,
         U5825_n1, U5826_n1, U5827_n1, U5828_n1, U5829_n1, U5830_n1, U5831_n1,
         U5832_n1, U5833_n1, U5834_n1, U5835_n1, U5836_n1, U5837_n1, U5838_n1,
         U5839_n1, U5840_n1, U5841_n1, U5842_n1, U5843_n1, U5844_n1, U5845_n1,
         U5846_n1, U5847_n1, U5848_n1, U5849_n1, U5850_n1, U5851_n1, U5852_n1,
         U5853_n1, U5854_n1, U5855_n1, U5856_n1, U5857_n1, U5858_n1, U5859_n1,
         U5860_n1, U5861_n1, U5862_n1, U5863_n1, U5864_n1, U5865_n1, U5866_n1,
         U5867_n1, U5868_n1, U5869_n1, U5870_n1, U5871_n1, U5872_n1, U5873_n1,
         U5874_n1, U5875_n1, U5876_n1, U5877_n1, U5878_n1, U5879_n1, U5880_n1,
         U5881_n1, U5882_n1, U5883_n1, U5884_n1, U5885_n1, U5886_n1, U5887_n1,
         U5888_n1, U5889_n1, U5890_n1, U5891_n1, U5892_n1, U5893_n1, U5894_n1,
         U5895_n1, U5896_n1, U5897_n1, U5898_n1, U5899_n1, U5900_n1, U5901_n1,
         U5902_n1, U5903_n1, U5904_n1, U5905_n1, U5906_n1, U5907_n1, U5908_n1,
         U5909_n1, U5910_n1, U5911_n1, U5912_n1, U5913_n1, U5914_n1, U5915_n1,
         U5916_n1, U5917_n1, U5918_n1, U5919_n1, U5920_n1, U5921_n1, U5922_n1,
         U5923_n1, U5924_n1, U5925_n1, U5926_n1, U5927_n1, U5928_n1, U5929_n1,
         U5930_n1, U5931_n1, U5932_n1, U5933_n1, U5934_n1, U5935_n1, U5936_n1,
         U5937_n1, U5938_n1, U5939_n1, U5940_n1, U5941_n1, U5942_n1, U5943_n1,
         U5944_n1, U5945_n1, U5946_n1, U5947_n1, U5948_n1, U5949_n1, U5950_n1,
         U5951_n1, U5952_n1, U5953_n1, U5954_n1, U5955_n1, U5956_n1, U5957_n1,
         U5958_n1, U5959_n1, U5960_n1, U5961_n1, U5962_n1, U5963_n1, U5964_n1,
         U5965_n1, U5966_n1, U5967_n1, U5968_n1, U5969_n1, U5970_n1, U5971_n1,
         U5972_n1, U5973_n1, U5974_n1, U5975_n1, U5976_n1, U5977_n1, U5978_n1,
         U5979_n1, U5980_n1, U5981_n1, U5982_n1, U5983_n1, U5984_n1, U5985_n1,
         U5986_n1, U5987_n1, U5988_n1, U5989_n1, U5990_n1, U5991_n1, U5992_n1,
         U5993_n1, U5994_n1, U5995_n1, U5996_n1, U5997_n1, U5998_n1, U5999_n1,
         U6000_n1, U6001_n1, U6002_n1, U6003_n1, U6004_n1, U6005_n1, U6006_n1,
         U6007_n1, U6008_n1, U6009_n1, U6010_n1, U6011_n1, U6012_n1, U6013_n1,
         U6014_n1, U6015_n1, U6016_n1, U6017_n1, U6018_n1, U6019_n1, U6020_n1,
         U6021_n1, U6022_n1, U6023_n1, U6024_n1, U6025_n1, U6026_n1, U6027_n1,
         U6028_n1, U6029_n1, U6030_n1, U6031_n1, U6032_n1, U6033_n1, U6034_n1,
         U6035_n1, U6036_n1, U6037_n1, U6038_n1, U6039_n1, U6040_n1, U6041_n1,
         U6042_n1, U6043_n1, U6044_n1, U6045_n1, U6046_n1, U6047_n1, U6048_n1,
         U6049_n1, U6050_n1, U6051_n1, U6052_n1, U6053_n1, U6054_n1, U6055_n1,
         U6056_n1, U6057_n1, U6058_n1, U6059_n1, U6060_n1, U6061_n1, U6062_n1,
         U6063_n1, U6064_n1, U6065_n1, U6066_n1, U6067_n1, U6068_n1, U6069_n1,
         U6070_n1, U6071_n1, U6072_n1, U6073_n1, U6074_n1, U6075_n1, U6076_n1,
         U6077_n1, U6078_n1, U6079_n1, U6080_n1, U6081_n1, U6082_n1, U6083_n1,
         U6084_n1, U6085_n1, U6086_n1, U6087_n1, U6088_n1, U6089_n1, U6090_n1,
         U6091_n1, U6092_n1, U6093_n1, U6094_n1, U6095_n1, U6096_n1, U6097_n1,
         U6098_n1, U6099_n1, U6100_n1, U6101_n1, U6102_n1, U6103_n1, U6104_n1,
         U6105_n1, U6106_n1, U6107_n1, U6108_n1, U6109_n1, U6110_n1, U6111_n1,
         U6112_n1, U6113_n1, U6114_n1, U6115_n1, U6116_n1, U6117_n1, U6118_n1,
         U6119_n1, U6120_n1, U6121_n1, U6122_n1, U6123_n1, U6124_n1, U6125_n1,
         U6126_n1, U6127_n1, U6128_n1, U6129_n1, U6130_n1, U6131_n1, U6132_n1,
         U6133_n1, U6134_n1, U6135_n1, U6136_n1, U6137_n1, U6138_n1, U6139_n1,
         U6140_n1, U6141_n1, U6142_n1, U6143_n1, U6144_n1, U6145_n1, U6146_n1,
         U6147_n1, U6148_n1, U6149_n1, U6150_n1, U6151_n1, U6152_n1, U6153_n1,
         U6154_n1, U6155_n1, U6156_n1, U6157_n1, U6158_n1, U6159_n1, U6160_n1,
         U6161_n1, U6162_n1, U6163_n1, U6164_n1, U6165_n1, U6166_n1, U6167_n1,
         U6168_n1, U6169_n1, U6170_n1, U6171_n1, U6172_n1, U6173_n1, U6174_n1,
         U6175_n1, U6176_n1, U6177_n1, U6178_n1, U6179_n1, U6180_n1, U6181_n1,
         U6182_n1, U6183_n1, U6184_n1, U6185_n1, U6186_n1, U6187_n1, U6188_n1,
         U6189_n1, U6190_n1, U6191_n1, U6192_n1, U6193_n1, U6194_n1, U6195_n1,
         U6196_n1, U6197_n1, U6198_n1, U6199_n1, U6200_n1, U6201_n1, U6202_n1,
         U6203_n1, U6204_n1, U6205_n1, U6206_n1, U6207_n1, U6208_n1, U6209_n1,
         U6210_n1, U6211_n1, U6212_n1, U6213_n1, U6214_n1, U6215_n1, U6216_n1,
         U6217_n1, U6218_n1, U6219_n1, U6220_n1, U6221_n1, U6222_n1, U6223_n1,
         U6224_n1, U6225_n1, U6226_n1, U6227_n1, U6228_n1, U6229_n1, U6230_n1,
         U6231_n1, U6232_n1, U6233_n1, U6234_n1, U6235_n1, U6236_n1, U6237_n1,
         U6238_n1, U6239_n1, U6240_n1, U6241_n1, U6242_n1, U6243_n1, U6244_n1,
         U6245_n1, U6246_n1, U6247_n1, U6248_n1, U6249_n1, U6250_n1, U6251_n1,
         U6252_n1, U6253_n1, U6254_n1, U6255_n1, U6256_n1, U6257_n1, U6258_n1,
         U6259_n1, U6260_n1, U6261_n1, U6262_n1, U6263_n1, U6264_n1, U6265_n1,
         U6266_n1, U6267_n1, U6268_n1, U6269_n1, U6270_n1, U6271_n1, U6272_n1,
         U6273_n1, U6274_n1, U6275_n1, U6276_n1, U6277_n1, U6278_n1, U6279_n1,
         U6280_n1, U6281_n1, U6282_n1, U6283_n1, U6284_n1, U6285_n1, U6286_n1,
         U6287_n1, U6288_n1, U6289_n1, U6290_n1, U6291_n1, U6292_n1, U6293_n1,
         U6294_n1, U6295_n1, U6296_n1, U6297_n1, U6298_n1, U6299_n1, U6300_n1,
         U6301_n1, U6302_n1, U6303_n1, U6304_n1, U6305_n1, U6306_n1, U6307_n1,
         U6308_n1, U6309_n1, U6310_n1, U6311_n1, U6312_n1, U6313_n1, U6314_n1,
         U6315_n1, U6316_n1, U6317_n1, U6318_n1, U6319_n1, U6320_n1, U6321_n1,
         U6322_n1, U6323_n1, U6324_n1, U6325_n1, U6326_n1, U6327_n1, U6328_n1,
         U6329_n1, U6330_n1, U6331_n1, U6332_n1, U6333_n1, U6334_n1, U6335_n1,
         U6336_n1, U6337_n1, U6338_n1, U6339_n1, U6340_n1, U6341_n1, U6342_n1,
         U6343_n1, U6344_n1, U6345_n1, U6346_n1, U6347_n1, U6348_n1, U6349_n1,
         U6350_n1, U6351_n1, U6352_n1, U6353_n1, U6354_n1, U6355_n1, U6356_n1,
         U6357_n1, U6358_n1, U6359_n1, U6360_n1, U6361_n1, U6362_n1, U6363_n1,
         U6364_n1, U6365_n1, U6366_n1, U6367_n1, U6368_n1, U6369_n1, U6370_n1,
         U6371_n1, U6372_n1, U6373_n1, U6374_n1, U6375_n1, U6376_n1, U6377_n1,
         U6378_n1, U6379_n1, U6380_n1, U6381_n1, U6382_n1, U6383_n1, U6384_n1,
         U6385_n1, U6386_n1, U6387_n1, U6388_n1, U6389_n1, U6390_n1, U6391_n1,
         U6392_n1, U6393_n1, U6394_n1, U6395_n1, U6396_n1, U6397_n1, U6398_n1,
         U6399_n1, U6400_n1, U6401_n1, U6402_n1, U6403_n1, U6404_n1, U6405_n1,
         U6406_n1, U6407_n1, U6408_n1, U6409_n1, U6410_n1, U6411_n1, U6412_n1,
         U6413_n1, U6414_n1, U6415_n1, U6416_n1, U6417_n1, U6418_n1, U6419_n1,
         U6420_n1, U6421_n1, U6422_n1, U6423_n1, U6424_n1, U6425_n1, U6426_n1,
         U6427_n1, U6428_n1, U6429_n1, U6430_n1, U6431_n1, U6432_n1, U6433_n1,
         U6434_n1, U6435_n1, U6436_n1, U6437_n1, U6438_n1, U6439_n1, U6440_n1,
         U6441_n1, U6442_n1, U6443_n1, U6444_n1, U6445_n1, U6446_n1, U6447_n1,
         U6448_n1, U6449_n1, U6450_n1, U6451_n1, U6452_n1, U6453_n1, U6454_n1,
         U6455_n1, U6456_n1, U6457_n1, U6458_n1, U6459_n1, U6460_n1, U6461_n1,
         U6462_n1, U6463_n1, U6464_n1, U6465_n1, U6466_n1, U6467_n1, U6468_n1,
         U6469_n1, U6470_n1, U6471_n1, U6472_n1, U6473_n1, U6474_n1, U6475_n1,
         U6476_n1, U6477_n1, U6478_n1, U6479_n1, U6480_n1, U6481_n1, U6482_n1;
  assign CRC_OUT_9_1 = test_so9;
  assign CRC_OUT_9_19 = test_so10;
  assign CRC_OUT_8_7 = test_so20;
  assign CRC_OUT_8_25 = test_so21;
  assign CRC_OUT_7_10 = test_so31;
  assign CRC_OUT_7_27 = test_so32;
  assign CRC_OUT_6_5 = test_so42;
  assign CRC_OUT_6_22 = test_so43;
  assign CRC_OUT_5_0 = test_so53;
  assign CRC_OUT_5_17 = test_so54;
  assign CRC_OUT_4_12 = test_so65;
  assign CRC_OUT_4_29 = test_so66;
  assign CRC_OUT_3_7 = test_so76;
  assign CRC_OUT_3_24 = test_so77;
  assign CRC_OUT_2_2 = test_so87;
  assign CRC_OUT_2_19 = test_so88;
  assign CRC_OUT_1_14 = test_so99;
  assign CRC_OUT_1_31 = test_so100;

  SDFFX1 DFF_0_Q_reg ( .D(WX484), .SI(test_si1), .SE(n4280), .CLK(n4569), .Q(
        WX485) );
  SDFFX1 DFF_1_Q_reg ( .D(WX486), .SI(WX485), .SE(n4275), .CLK(n4571), .Q(
        WX487) );
  SDFFX1 DFF_2_Q_reg ( .D(WX488), .SI(WX487), .SE(n4275), .CLK(n4571), .Q(
        WX489) );
  SDFFX1 DFF_3_Q_reg ( .D(WX490), .SI(WX489), .SE(n4276), .CLK(n4571), .Q(
        WX491) );
  SDFFX1 DFF_4_Q_reg ( .D(WX492), .SI(WX491), .SE(n4276), .CLK(n4571), .Q(
        WX493) );
  SDFFX1 DFF_5_Q_reg ( .D(WX494), .SI(WX493), .SE(n4276), .CLK(n4571), .Q(
        WX495) );
  SDFFX1 DFF_6_Q_reg ( .D(WX496), .SI(WX495), .SE(n4276), .CLK(n4571), .Q(
        WX497) );
  SDFFX1 DFF_7_Q_reg ( .D(WX498), .SI(WX497), .SE(n4276), .CLK(n4571), .Q(
        WX499) );
  SDFFX1 DFF_8_Q_reg ( .D(WX500), .SI(WX499), .SE(n4276), .CLK(n4571), .Q(
        WX501) );
  SDFFX1 DFF_9_Q_reg ( .D(WX502), .SI(WX501), .SE(n4277), .CLK(n4570), .Q(
        WX503) );
  SDFFX1 DFF_10_Q_reg ( .D(WX504), .SI(WX503), .SE(n4277), .CLK(n4570), .Q(
        WX505) );
  SDFFX1 DFF_11_Q_reg ( .D(WX506), .SI(WX505), .SE(n4277), .CLK(n4570), .Q(
        WX507) );
  SDFFX1 DFF_12_Q_reg ( .D(WX508), .SI(WX507), .SE(n4277), .CLK(n4570), .Q(
        WX509) );
  SDFFX1 DFF_13_Q_reg ( .D(WX510), .SI(WX509), .SE(n4277), .CLK(n4570), .Q(
        WX511) );
  SDFFX1 DFF_14_Q_reg ( .D(WX512), .SI(WX511), .SE(n4277), .CLK(n4570), .Q(
        WX513) );
  SDFFX1 DFF_15_Q_reg ( .D(WX514), .SI(WX513), .SE(n4278), .CLK(n4570), .Q(
        WX515) );
  SDFFX1 DFF_16_Q_reg ( .D(WX516), .SI(WX515), .SE(n4278), .CLK(n4570), .Q(
        WX517) );
  SDFFX1 DFF_17_Q_reg ( .D(WX518), .SI(WX517), .SE(n4278), .CLK(n4570), .Q(
        test_so1) );
  SDFFX1 DFF_18_Q_reg ( .D(WX520), .SI(test_si2), .SE(n4278), .CLK(n4570), .Q(
        WX521) );
  SDFFX1 DFF_19_Q_reg ( .D(WX522), .SI(WX521), .SE(n4278), .CLK(n4570), .Q(
        WX523) );
  SDFFX1 DFF_20_Q_reg ( .D(WX524), .SI(WX523), .SE(n4278), .CLK(n4570), .Q(
        WX525) );
  SDFFX1 DFF_21_Q_reg ( .D(WX526), .SI(WX525), .SE(n4279), .CLK(n4569), .Q(
        WX527) );
  SDFFX1 DFF_22_Q_reg ( .D(WX528), .SI(WX527), .SE(n4279), .CLK(n4569), .Q(
        WX529) );
  SDFFX1 DFF_23_Q_reg ( .D(WX530), .SI(WX529), .SE(n4279), .CLK(n4569), .Q(
        WX531) );
  SDFFX1 DFF_24_Q_reg ( .D(WX532), .SI(WX531), .SE(n4279), .CLK(n4569), .Q(
        WX533) );
  SDFFX1 DFF_25_Q_reg ( .D(WX534), .SI(WX533), .SE(n4279), .CLK(n4569), .Q(
        WX535) );
  SDFFX1 DFF_26_Q_reg ( .D(WX536), .SI(WX535), .SE(n4279), .CLK(n4569), .Q(
        WX537) );
  SDFFX1 DFF_27_Q_reg ( .D(WX538), .SI(WX537), .SE(n4280), .CLK(n4569), .Q(
        WX539) );
  SDFFX1 DFF_28_Q_reg ( .D(WX540), .SI(WX539), .SE(n4280), .CLK(n4569), .Q(
        WX541) );
  SDFFX1 DFF_29_Q_reg ( .D(WX542), .SI(WX541), .SE(n4280), .CLK(n4569), .Q(
        WX543) );
  SDFFX1 DFF_30_Q_reg ( .D(WX544), .SI(WX543), .SE(n4280), .CLK(n4569), .Q(
        WX545) );
  SDFFX1 DFF_31_Q_reg ( .D(WX546), .SI(WX545), .SE(n4280), .CLK(n4569), .Q(
        WX547) );
  SDFFX1 DFF_32_Q_reg ( .D(WX644), .SI(WX547), .SE(n4275), .CLK(n4571), .Q(
        WX645), .QN(n3529) );
  SDFFX1 DFF_33_Q_reg ( .D(WX646), .SI(WX645), .SE(n4275), .CLK(n4571), .Q(
        WX647), .QN(n3527) );
  SDFFX1 DFF_34_Q_reg ( .D(WX648), .SI(WX647), .SE(n4275), .CLK(n4571), .Q(
        WX649), .QN(n3525) );
  SDFFX1 DFF_35_Q_reg ( .D(WX650), .SI(WX649), .SE(n4275), .CLK(n4571), .Q(
        test_so2) );
  SDFFX1 DFF_36_Q_reg ( .D(WX652), .SI(test_si3), .SE(n4274), .CLK(n4572), .Q(
        WX653), .QN(n3521) );
  SDFFX1 DFF_37_Q_reg ( .D(WX654), .SI(WX653), .SE(n4274), .CLK(n4572), .Q(
        WX655), .QN(n3519) );
  SDFFX1 DFF_38_Q_reg ( .D(WX656), .SI(WX655), .SE(n4274), .CLK(n4572), .Q(
        WX657), .QN(n3517) );
  SDFFX1 DFF_39_Q_reg ( .D(WX658), .SI(WX657), .SE(n4273), .CLK(n4572), .Q(
        WX659), .QN(n3515) );
  SDFFX1 DFF_40_Q_reg ( .D(WX660), .SI(WX659), .SE(n4273), .CLK(n4572), .Q(
        WX661), .QN(n3513) );
  SDFFX1 DFF_41_Q_reg ( .D(WX662), .SI(WX661), .SE(n4273), .CLK(n4572), .Q(
        WX663), .QN(n3511) );
  SDFFX1 DFF_42_Q_reg ( .D(WX664), .SI(WX663), .SE(n4272), .CLK(n4573), .Q(
        WX665), .QN(n3509) );
  SDFFX1 DFF_43_Q_reg ( .D(WX666), .SI(WX665), .SE(n4272), .CLK(n4573), .Q(
        WX667), .QN(n3507) );
  SDFFX1 DFF_44_Q_reg ( .D(WX668), .SI(WX667), .SE(n4272), .CLK(n4573), .Q(
        WX669), .QN(n3505) );
  SDFFX1 DFF_45_Q_reg ( .D(WX670), .SI(WX669), .SE(n4271), .CLK(n4573), .Q(
        WX671), .QN(n3503) );
  SDFFX1 DFF_46_Q_reg ( .D(WX672), .SI(WX671), .SE(n4271), .CLK(n4573), .Q(
        WX673), .QN(n3501) );
  SDFFX1 DFF_47_Q_reg ( .D(WX674), .SI(WX673), .SE(n4270), .CLK(n4574), .Q(
        WX675), .QN(n3499) );
  SDFFX1 DFF_48_Q_reg ( .D(WX676), .SI(WX675), .SE(n4270), .CLK(n4574), .Q(
        WX677), .QN(n3497) );
  SDFFX1 DFF_49_Q_reg ( .D(WX678), .SI(WX677), .SE(n4269), .CLK(n4574), .Q(
        WX679), .QN(n3495) );
  SDFFX1 DFF_50_Q_reg ( .D(WX680), .SI(WX679), .SE(n4268), .CLK(n4575), .Q(
        WX681), .QN(n3493) );
  SDFFX1 DFF_51_Q_reg ( .D(WX682), .SI(WX681), .SE(n4268), .CLK(n4575), .Q(
        WX683), .QN(n3491) );
  SDFFX1 DFF_52_Q_reg ( .D(WX684), .SI(WX683), .SE(n4267), .CLK(n4575), .Q(
        WX685), .QN(n3489) );
  SDFFX1 DFF_53_Q_reg ( .D(WX686), .SI(WX685), .SE(n4266), .CLK(n4576), .Q(
        test_so3) );
  SDFFX1 DFF_54_Q_reg ( .D(WX688), .SI(test_si4), .SE(n4265), .CLK(n4576), .Q(
        WX689), .QN(n3485) );
  SDFFX1 DFF_55_Q_reg ( .D(WX690), .SI(WX689), .SE(n4265), .CLK(n4576), .Q(
        WX691), .QN(n3483) );
  SDFFX1 DFF_56_Q_reg ( .D(WX692), .SI(WX691), .SE(n4264), .CLK(n4577), .Q(
        WX693), .QN(n3481) );
  SDFFX1 DFF_57_Q_reg ( .D(WX694), .SI(WX693), .SE(n4264), .CLK(n4577), .Q(
        WX695), .QN(n3479) );
  SDFFX1 DFF_58_Q_reg ( .D(WX696), .SI(WX695), .SE(n4263), .CLK(n4577), .Q(
        WX697), .QN(n3477) );
  SDFFX1 DFF_59_Q_reg ( .D(WX698), .SI(WX697), .SE(n4262), .CLK(n4578), .Q(
        WX699), .QN(n3475) );
  SDFFX1 DFF_60_Q_reg ( .D(WX700), .SI(WX699), .SE(n4262), .CLK(n4578), .Q(
        WX701), .QN(n3473) );
  SDFFX1 DFF_61_Q_reg ( .D(WX702), .SI(WX701), .SE(n4261), .CLK(n4578), .Q(
        WX703), .QN(n3471) );
  SDFFX1 DFF_62_Q_reg ( .D(WX704), .SI(WX703), .SE(n4260), .CLK(n4579), .Q(
        WX705), .QN(n3469) );
  SDFFX1 DFF_63_Q_reg ( .D(WX706), .SI(WX705), .SE(n4260), .CLK(n4579), .Q(
        WX707), .QN(n3467) );
  SDFFX1 DFF_64_Q_reg ( .D(WX708), .SI(WX707), .SE(n4259), .CLK(n4579), .Q(
        WX709), .QN(n7260) );
  SDFFX1 DFF_65_Q_reg ( .D(WX710), .SI(WX709), .SE(n4258), .CLK(n4580), .Q(
        WX711) );
  SDFFX1 DFF_66_Q_reg ( .D(WX712), .SI(WX711), .SE(n4258), .CLK(n4580), .Q(
        WX713), .QN(n3811) );
  SDFFX1 DFF_67_Q_reg ( .D(WX714), .SI(WX713), .SE(n4274), .CLK(n4572), .Q(
        WX715), .QN(n7263) );
  SDFFX1 DFF_68_Q_reg ( .D(WX716), .SI(WX715), .SE(n4274), .CLK(n4572), .Q(
        WX717), .QN(n3820) );
  SDFFX1 DFF_69_Q_reg ( .D(WX718), .SI(WX717), .SE(n4274), .CLK(n4572), .Q(
        WX719), .QN(n3822) );
  SDFFX1 DFF_70_Q_reg ( .D(WX720), .SI(WX719), .SE(n4273), .CLK(n4572), .Q(
        WX721), .QN(n3827) );
  SDFFX1 DFF_71_Q_reg ( .D(WX722), .SI(WX721), .SE(n4273), .CLK(n4572), .Q(
        test_so4) );
  SDFFX1 DFF_72_Q_reg ( .D(WX724), .SI(test_si5), .SE(n4273), .CLK(n4572), .Q(
        WX725), .QN(n3834) );
  SDFFX1 DFF_73_Q_reg ( .D(WX726), .SI(WX725), .SE(n4272), .CLK(n4573), .Q(
        WX727) );
  SDFFX1 DFF_74_Q_reg ( .D(WX728), .SI(WX727), .SE(n4272), .CLK(n4573), .Q(
        WX729) );
  SDFFX1 DFF_75_Q_reg ( .D(WX730), .SI(WX729), .SE(n4272), .CLK(n4573), .Q(
        WX731), .QN(n7269) );
  SDFFX1 DFF_76_Q_reg ( .D(WX732), .SI(WX731), .SE(n4271), .CLK(n4573), .Q(
        WX733), .QN(n3809) );
  SDFFX1 DFF_77_Q_reg ( .D(WX734), .SI(WX733), .SE(n4271), .CLK(n4573), .Q(
        WX735), .QN(n3818) );
  SDFFX1 DFF_78_Q_reg ( .D(WX736), .SI(WX735), .SE(n4270), .CLK(n4574), .Q(
        WX737), .QN(n3825) );
  SDFFX1 DFF_79_Q_reg ( .D(WX738), .SI(WX737), .SE(n4270), .CLK(n4574), .Q(
        WX739) );
  SDFFX1 DFF_80_Q_reg ( .D(WX740), .SI(WX739), .SE(n4269), .CLK(n4574), .Q(
        WX741) );
  SDFFX1 DFF_81_Q_reg ( .D(WX742), .SI(WX741), .SE(n4269), .CLK(n4574), .Q(
        WX743), .QN(n3857) );
  SDFFX1 DFF_82_Q_reg ( .D(WX744), .SI(WX743), .SE(n4268), .CLK(n4575), .Q(
        WX745), .QN(n3813) );
  SDFFX1 DFF_83_Q_reg ( .D(WX746), .SI(WX745), .SE(n4267), .CLK(n4575), .Q(
        WX747), .QN(n3829) );
  SDFFX1 DFF_84_Q_reg ( .D(WX748), .SI(WX747), .SE(n4267), .CLK(n4575), .Q(
        WX749), .QN(n3864) );
  SDFFX1 DFF_85_Q_reg ( .D(WX750), .SI(WX749), .SE(n4266), .CLK(n4576), .Q(
        WX751), .QN(n7278) );
  SDFFX1 DFF_86_Q_reg ( .D(WX752), .SI(WX751), .SE(n4266), .CLK(n4576), .Q(
        WX753), .QN(n7256) );
  SDFFX1 DFF_87_Q_reg ( .D(WX754), .SI(WX753), .SE(n4265), .CLK(n4576), .Q(
        WX755), .QN(n3837) );
  SDFFX1 DFF_88_Q_reg ( .D(WX756), .SI(WX755), .SE(n4264), .CLK(n4577), .Q(
        WX757) );
  SDFFX1 DFF_89_Q_reg ( .D(WX758), .SI(WX757), .SE(n4263), .CLK(n4577), .Q(
        test_so5) );
  SDFFX1 DFF_90_Q_reg ( .D(WX760), .SI(test_si6), .SE(n4263), .CLK(n4577), .Q(
        WX761), .QN(n3839) );
  SDFFX1 DFF_91_Q_reg ( .D(WX762), .SI(WX761), .SE(n4262), .CLK(n4578), .Q(
        WX763), .QN(n3841) );
  SDFFX1 DFF_92_Q_reg ( .D(WX764), .SI(WX763), .SE(n4261), .CLK(n4578), .Q(
        WX765), .QN(n3807) );
  SDFFX1 DFF_93_Q_reg ( .D(WX766), .SI(WX765), .SE(n4261), .CLK(n4578), .Q(
        WX767) );
  SDFFX1 DFF_94_Q_reg ( .D(WX768), .SI(WX767), .SE(n4260), .CLK(n4579), .Q(
        WX769), .QN(n3815) );
  SDFFX1 DFF_95_Q_reg ( .D(WX770), .SI(WX769), .SE(n4259), .CLK(n4579), .Q(
        WX771) );
  SDFFX1 DFF_96_Q_reg ( .D(WX772), .SI(WX771), .SE(n4259), .CLK(n4579), .Q(
        WX773) );
  SDFFX1 DFF_97_Q_reg ( .D(WX774), .SI(WX773), .SE(n4258), .CLK(n4580), .Q(
        WX775), .QN(n3804) );
  SDFFX1 DFF_98_Q_reg ( .D(WX776), .SI(WX775), .SE(n4258), .CLK(n4580), .Q(
        WX777), .QN(n7262) );
  SDFFX1 DFF_99_Q_reg ( .D(WX778), .SI(WX777), .SE(n4257), .CLK(n4580), .Q(
        WX779) );
  SDFFX1 DFF_100_Q_reg ( .D(WX780), .SI(WX779), .SE(n4257), .CLK(n4580), .Q(
        WX781), .QN(n7264) );
  SDFFX1 DFF_101_Q_reg ( .D(WX782), .SI(WX781), .SE(n4257), .CLK(n4580), .Q(
        WX783), .QN(n7265) );
  SDFFX1 DFF_102_Q_reg ( .D(WX784), .SI(WX783), .SE(n4256), .CLK(n4581), .Q(
        WX785), .QN(n7266) );
  SDFFX1 DFF_103_Q_reg ( .D(WX786), .SI(WX785), .SE(n4256), .CLK(n4581), .Q(
        WX787), .QN(n7267) );
  SDFFX1 DFF_104_Q_reg ( .D(WX788), .SI(WX787), .SE(n4256), .CLK(n4581), .Q(
        WX789), .QN(n7268) );
  SDFFX1 DFF_105_Q_reg ( .D(WX790), .SI(WX789), .SE(n4255), .CLK(n4581), .Q(
        WX791), .QN(n3843) );
  SDFFX1 DFF_106_Q_reg ( .D(WX792), .SI(WX791), .SE(n4255), .CLK(n4581), .Q(
        WX793), .QN(n3849) );
  SDFFX1 DFF_107_Q_reg ( .D(WX794), .SI(WX793), .SE(n4255), .CLK(n4581), .Q(
        test_so6) );
  SDFFX1 DFF_108_Q_reg ( .D(WX796), .SI(test_si7), .SE(n4271), .CLK(n4573), 
        .Q(WX797), .QN(n7270) );
  SDFFX1 DFF_109_Q_reg ( .D(WX798), .SI(WX797), .SE(n4271), .CLK(n4573), .Q(
        WX799), .QN(n7271) );
  SDFFX1 DFF_110_Q_reg ( .D(WX800), .SI(WX799), .SE(n4270), .CLK(n4574), .Q(
        WX801), .QN(n7272) );
  SDFFX1 DFF_111_Q_reg ( .D(WX802), .SI(WX801), .SE(n4270), .CLK(n4574), .Q(
        WX803), .QN(n7273) );
  SDFFX1 DFF_112_Q_reg ( .D(WX804), .SI(WX803), .SE(n4269), .CLK(n4574), .Q(
        WX805), .QN(n3846) );
  SDFFX1 DFF_113_Q_reg ( .D(WX806), .SI(WX805), .SE(n4269), .CLK(n4574), .Q(
        WX807), .QN(n7274) );
  SDFFX1 DFF_114_Q_reg ( .D(WX808), .SI(WX807), .SE(n4268), .CLK(n4575), .Q(
        WX809), .QN(n7275) );
  SDFFX1 DFF_115_Q_reg ( .D(WX810), .SI(WX809), .SE(n4267), .CLK(n4575), .Q(
        WX811), .QN(n7276) );
  SDFFX1 DFF_116_Q_reg ( .D(WX812), .SI(WX811), .SE(n4267), .CLK(n4575), .Q(
        WX813), .QN(n7277) );
  SDFFX1 DFF_117_Q_reg ( .D(WX814), .SI(WX813), .SE(n4266), .CLK(n4576), .Q(
        WX815) );
  SDFFX1 DFF_118_Q_reg ( .D(WX816), .SI(WX815), .SE(n4265), .CLK(n4576), .Q(
        WX817) );
  SDFFX1 DFF_119_Q_reg ( .D(WX818), .SI(WX817), .SE(n4265), .CLK(n4576), .Q(
        WX819), .QN(n7257) );
  SDFFX1 DFF_120_Q_reg ( .D(WX820), .SI(WX819), .SE(n4264), .CLK(n4577), .Q(
        WX821), .QN(n3861) );
  SDFFX1 DFF_121_Q_reg ( .D(WX822), .SI(WX821), .SE(n4263), .CLK(n4577), .Q(
        WX823) );
  SDFFX1 DFF_122_Q_reg ( .D(WX824), .SI(WX823), .SE(n4263), .CLK(n4577), .Q(
        WX825), .QN(n7258) );
  SDFFX1 DFF_123_Q_reg ( .D(WX826), .SI(WX825), .SE(n4262), .CLK(n4578), .Q(
        WX827), .QN(n7259) );
  SDFFX1 DFF_124_Q_reg ( .D(WX828), .SI(WX827), .SE(n4261), .CLK(n4578), .Q(
        WX829), .QN(n7261) );
  SDFFX1 DFF_125_Q_reg ( .D(WX830), .SI(WX829), .SE(n4261), .CLK(n4578), .Q(
        test_so7) );
  SDFFX1 DFF_126_Q_reg ( .D(WX832), .SI(test_si8), .SE(n4260), .CLK(n4579), 
        .Q(WX833), .QN(n7279) );
  SDFFX1 DFF_127_Q_reg ( .D(WX834), .SI(WX833), .SE(n4259), .CLK(n4579), .Q(
        WX835), .QN(n3866) );
  SDFFX1 DFF_128_Q_reg ( .D(WX836), .SI(WX835), .SE(n4259), .CLK(n4579), .Q(
        WX837), .QN(n3855) );
  SDFFX1 DFF_129_Q_reg ( .D(WX838), .SI(WX837), .SE(n4258), .CLK(n4580), .Q(
        WX839), .QN(n3805) );
  SDFFX1 DFF_130_Q_reg ( .D(WX840), .SI(WX839), .SE(n4258), .CLK(n4580), .Q(
        WX841), .QN(n3810) );
  SDFFX1 DFF_131_Q_reg ( .D(WX842), .SI(WX841), .SE(n4257), .CLK(n4580), .Q(
        WX843), .QN(n3816) );
  SDFFX1 DFF_132_Q_reg ( .D(WX844), .SI(WX843), .SE(n4257), .CLK(n4580), .Q(
        WX845), .QN(n3819) );
  SDFFX1 DFF_133_Q_reg ( .D(WX846), .SI(WX845), .SE(n4257), .CLK(n4580), .Q(
        WX847), .QN(n3821) );
  SDFFX1 DFF_134_Q_reg ( .D(WX848), .SI(WX847), .SE(n4256), .CLK(n4581), .Q(
        WX849), .QN(n3826) );
  SDFFX1 DFF_135_Q_reg ( .D(WX850), .SI(WX849), .SE(n4256), .CLK(n4581), .Q(
        WX851), .QN(n3832) );
  SDFFX1 DFF_136_Q_reg ( .D(WX852), .SI(WX851), .SE(n4256), .CLK(n4581), .Q(
        WX853), .QN(n3833) );
  SDFFX1 DFF_137_Q_reg ( .D(WX854), .SI(WX853), .SE(n4255), .CLK(n4581), .Q(
        WX855), .QN(n3844) );
  SDFFX1 DFF_138_Q_reg ( .D(WX856), .SI(WX855), .SE(n4255), .CLK(n4581), .Q(
        WX857), .QN(n3850) );
  SDFFX1 DFF_139_Q_reg ( .D(WX858), .SI(WX857), .SE(n4255), .CLK(n4581), .Q(
        WX859), .QN(n3853) );
  SDFFX1 DFF_140_Q_reg ( .D(WX860), .SI(WX859), .SE(n4254), .CLK(n4582), .Q(
        WX861), .QN(n3808) );
  SDFFX1 DFF_141_Q_reg ( .D(WX862), .SI(WX861), .SE(n4254), .CLK(n4582), .Q(
        WX863), .QN(n3817) );
  SDFFX1 DFF_142_Q_reg ( .D(WX864), .SI(WX863), .SE(n4254), .CLK(n4582), .Q(
        WX865), .QN(n3824) );
  SDFFX1 DFF_143_Q_reg ( .D(WX866), .SI(WX865), .SE(n4254), .CLK(n4582), .Q(
        test_so8) );
  SDFFX1 DFF_144_Q_reg ( .D(WX868), .SI(test_si9), .SE(n4269), .CLK(n4574), 
        .Q(WX869), .QN(n3847) );
  SDFFX1 DFF_145_Q_reg ( .D(WX870), .SI(WX869), .SE(n4268), .CLK(n4575), .Q(
        WX871), .QN(n3856) );
  SDFFX1 DFF_146_Q_reg ( .D(WX872), .SI(WX871), .SE(n4268), .CLK(n4575), .Q(
        WX873), .QN(n3812) );
  SDFFX1 DFF_147_Q_reg ( .D(WX874), .SI(WX873), .SE(n4267), .CLK(n4575), .Q(
        WX875), .QN(n3828) );
  SDFFX1 DFF_148_Q_reg ( .D(WX876), .SI(WX875), .SE(n4266), .CLK(n4576), .Q(
        WX877), .QN(n3863) );
  SDFFX1 DFF_149_Q_reg ( .D(WX878), .SI(WX877), .SE(n4266), .CLK(n4576), .Q(
        WX879), .QN(n3823) );
  SDFFX1 DFF_150_Q_reg ( .D(WX880), .SI(WX879), .SE(n4265), .CLK(n4576), .Q(
        WX881), .QN(n3831) );
  SDFFX1 DFF_151_Q_reg ( .D(WX882), .SI(WX881), .SE(n4264), .CLK(n4577), .Q(
        WX883), .QN(n3836) );
  SDFFX1 DFF_152_Q_reg ( .D(WX884), .SI(WX883), .SE(n4264), .CLK(n4577), .Q(
        WX885), .QN(n3862) );
  SDFFX1 DFF_153_Q_reg ( .D(WX886), .SI(WX885), .SE(n4263), .CLK(n4577), .Q(
        WX887), .QN(n3852) );
  SDFFX1 DFF_154_Q_reg ( .D(WX888), .SI(WX887), .SE(n4262), .CLK(n4578), .Q(
        WX889), .QN(n3838) );
  SDFFX1 DFF_155_Q_reg ( .D(WX890), .SI(WX889), .SE(n4262), .CLK(n4578), .Q(
        WX891), .QN(n3840) );
  SDFFX1 DFF_156_Q_reg ( .D(WX892), .SI(WX891), .SE(n4261), .CLK(n4578), .Q(
        WX893), .QN(n3806) );
  SDFFX1 DFF_157_Q_reg ( .D(WX894), .SI(WX893), .SE(n4260), .CLK(n4579), .Q(
        WX895), .QN(n3859) );
  SDFFX1 DFF_158_Q_reg ( .D(WX896), .SI(WX895), .SE(n4260), .CLK(n4579), .Q(
        WX897), .QN(n3814) );
  SDFFX1 DFF_159_Q_reg ( .D(WX898), .SI(WX897), .SE(n4259), .CLK(n4579), .Q(
        WX899), .QN(n3867) );
  SDFFX1 DFF_160_Q_reg ( .D(WX1264), .SI(WX899), .SE(n3996), .CLK(n4711), .Q(
        CRC_OUT_9_0), .QN(DFF_160_n1) );
  SDFFX1 DFF_161_Q_reg ( .D(WX1266), .SI(CRC_OUT_9_0), .SE(n3996), .CLK(n4711), 
        .Q(test_so9) );
  SDFFX1 DFF_162_Q_reg ( .D(WX1268), .SI(test_si10), .SE(n3995), .CLK(n4711), 
        .Q(CRC_OUT_9_2), .QN(DFF_162_n1) );
  SDFFX1 DFF_163_Q_reg ( .D(WX1270), .SI(CRC_OUT_9_2), .SE(n3995), .CLK(n4711), 
        .Q(CRC_OUT_9_3) );
  SDFFX1 DFF_164_Q_reg ( .D(WX1272), .SI(CRC_OUT_9_3), .SE(n3995), .CLK(n4711), 
        .Q(CRC_OUT_9_4), .QN(DFF_164_n1) );
  SDFFX1 DFF_165_Q_reg ( .D(WX1274), .SI(CRC_OUT_9_4), .SE(n3995), .CLK(n4711), 
        .Q(CRC_OUT_9_5), .QN(DFF_165_n1) );
  SDFFX1 DFF_166_Q_reg ( .D(WX1276), .SI(CRC_OUT_9_5), .SE(n3995), .CLK(n4711), 
        .Q(CRC_OUT_9_6), .QN(DFF_166_n1) );
  SDFFX1 DFF_167_Q_reg ( .D(WX1278), .SI(CRC_OUT_9_6), .SE(n3995), .CLK(n4711), 
        .Q(CRC_OUT_9_7), .QN(DFF_167_n1) );
  SDFFX1 DFF_168_Q_reg ( .D(WX1280), .SI(CRC_OUT_9_7), .SE(n3994), .CLK(n4712), 
        .Q(CRC_OUT_9_8), .QN(DFF_168_n1) );
  SDFFX1 DFF_169_Q_reg ( .D(WX1282), .SI(CRC_OUT_9_8), .SE(n3994), .CLK(n4712), 
        .Q(CRC_OUT_9_9), .QN(DFF_169_n1) );
  SDFFX1 DFF_170_Q_reg ( .D(WX1284), .SI(CRC_OUT_9_9), .SE(n3994), .CLK(n4712), 
        .Q(CRC_OUT_9_10) );
  SDFFX1 DFF_171_Q_reg ( .D(WX1286), .SI(CRC_OUT_9_10), .SE(n3994), .CLK(n4712), .Q(CRC_OUT_9_11), .QN(DFF_171_n1) );
  SDFFX1 DFF_172_Q_reg ( .D(WX1288), .SI(CRC_OUT_9_11), .SE(n3994), .CLK(n4712), .Q(CRC_OUT_9_12), .QN(DFF_172_n1) );
  SDFFX1 DFF_173_Q_reg ( .D(WX1290), .SI(CRC_OUT_9_12), .SE(n3994), .CLK(n4712), .Q(CRC_OUT_9_13), .QN(DFF_173_n1) );
  SDFFX1 DFF_174_Q_reg ( .D(WX1292), .SI(CRC_OUT_9_13), .SE(n3993), .CLK(n4712), .Q(CRC_OUT_9_14), .QN(DFF_174_n1) );
  SDFFX1 DFF_175_Q_reg ( .D(WX1294), .SI(CRC_OUT_9_14), .SE(n3993), .CLK(n4712), .Q(CRC_OUT_9_15), .QN(DFF_175_n1) );
  SDFFX1 DFF_176_Q_reg ( .D(WX1296), .SI(CRC_OUT_9_15), .SE(n3993), .CLK(n4712), .Q(CRC_OUT_9_16), .QN(DFF_176_n1) );
  SDFFX1 DFF_177_Q_reg ( .D(WX1298), .SI(CRC_OUT_9_16), .SE(n3993), .CLK(n4712), .Q(CRC_OUT_9_17), .QN(DFF_177_n1) );
  SDFFX1 DFF_178_Q_reg ( .D(WX1300), .SI(CRC_OUT_9_17), .SE(n3993), .CLK(n4712), .Q(CRC_OUT_9_18), .QN(DFF_178_n1) );
  SDFFX1 DFF_179_Q_reg ( .D(WX1302), .SI(CRC_OUT_9_18), .SE(n3993), .CLK(n4712), .Q(test_so10) );
  SDFFX1 DFF_180_Q_reg ( .D(WX1304), .SI(test_si11), .SE(n4254), .CLK(n4582), 
        .Q(CRC_OUT_9_20), .QN(DFF_180_n1) );
  SDFFX1 DFF_181_Q_reg ( .D(WX1306), .SI(CRC_OUT_9_20), .SE(n4254), .CLK(n4582), .Q(CRC_OUT_9_21), .QN(DFF_181_n1) );
  SDFFX1 DFF_182_Q_reg ( .D(WX1308), .SI(CRC_OUT_9_21), .SE(n4253), .CLK(n4582), .Q(CRC_OUT_9_22), .QN(DFF_182_n1) );
  SDFFX1 DFF_183_Q_reg ( .D(WX1310), .SI(CRC_OUT_9_22), .SE(n4253), .CLK(n4582), .Q(CRC_OUT_9_23), .QN(DFF_183_n1) );
  SDFFX1 DFF_184_Q_reg ( .D(WX1312), .SI(CRC_OUT_9_23), .SE(n4253), .CLK(n4582), .Q(CRC_OUT_9_24), .QN(DFF_184_n1) );
  SDFFX1 DFF_185_Q_reg ( .D(WX1314), .SI(CRC_OUT_9_24), .SE(n4253), .CLK(n4582), .Q(CRC_OUT_9_25), .QN(DFF_185_n1) );
  SDFFX1 DFF_186_Q_reg ( .D(WX1316), .SI(CRC_OUT_9_25), .SE(n4253), .CLK(n4582), .Q(CRC_OUT_9_26), .QN(DFF_186_n1) );
  SDFFX1 DFF_187_Q_reg ( .D(WX1318), .SI(CRC_OUT_9_26), .SE(n4253), .CLK(n4582), .Q(CRC_OUT_9_27), .QN(DFF_187_n1) );
  SDFFX1 DFF_188_Q_reg ( .D(WX1320), .SI(CRC_OUT_9_27), .SE(n4252), .CLK(n4583), .Q(CRC_OUT_9_28), .QN(DFF_188_n1) );
  SDFFX1 DFF_189_Q_reg ( .D(WX1322), .SI(CRC_OUT_9_28), .SE(n4252), .CLK(n4583), .Q(CRC_OUT_9_29), .QN(DFF_189_n1) );
  SDFFX1 DFF_190_Q_reg ( .D(WX1324), .SI(CRC_OUT_9_29), .SE(n4252), .CLK(n4583), .Q(CRC_OUT_9_30), .QN(DFF_190_n1) );
  SDFFX1 DFF_191_Q_reg ( .D(WX1326), .SI(CRC_OUT_9_30), .SE(n4252), .CLK(n4583), .Q(CRC_OUT_9_31), .QN(DFF_191_n1) );
  SDFFX1 DFF_192_Q_reg ( .D(n33), .SI(CRC_OUT_9_31), .SE(n4252), .CLK(n4583), 
        .Q(WX1778) );
  SDFFX1 DFF_193_Q_reg ( .D(n34), .SI(WX1778), .SE(n4247), .CLK(n4585), .Q(
        n8702) );
  SDFFX1 DFF_194_Q_reg ( .D(n35), .SI(n8702), .SE(n4247), .CLK(n4585), .Q(
        n8701) );
  SDFFX1 DFF_195_Q_reg ( .D(n36), .SI(n8701), .SE(n4247), .CLK(n4585), .Q(
        n8700) );
  SDFFX1 DFF_196_Q_reg ( .D(n37), .SI(n8700), .SE(n4247), .CLK(n4585), .Q(
        n8699) );
  SDFFX1 DFF_197_Q_reg ( .D(n38), .SI(n8699), .SE(n4247), .CLK(n4585), .Q(
        test_so11) );
  SDFFX1 DFF_198_Q_reg ( .D(n39), .SI(test_si12), .SE(n4247), .CLK(n4585), .Q(
        n8696) );
  SDFFX1 DFF_199_Q_reg ( .D(n40), .SI(n8696), .SE(n4248), .CLK(n4585), .Q(
        n8695) );
  SDFFX1 DFF_200_Q_reg ( .D(n41), .SI(n8695), .SE(n4248), .CLK(n4585), .Q(
        n8694) );
  SDFFX1 DFF_201_Q_reg ( .D(n42), .SI(n8694), .SE(n4248), .CLK(n4585), .Q(
        n8693) );
  SDFFX1 DFF_202_Q_reg ( .D(n43), .SI(n8693), .SE(n4248), .CLK(n4585), .Q(
        n8692) );
  SDFFX1 DFF_203_Q_reg ( .D(n44), .SI(n8692), .SE(n4248), .CLK(n4585), .Q(
        n8691) );
  SDFFX1 DFF_204_Q_reg ( .D(n45), .SI(n8691), .SE(n4248), .CLK(n4585), .Q(
        n8690) );
  SDFFX1 DFF_205_Q_reg ( .D(n46), .SI(n8690), .SE(n4249), .CLK(n4584), .Q(
        n8689) );
  SDFFX1 DFF_206_Q_reg ( .D(n47), .SI(n8689), .SE(n4249), .CLK(n4584), .Q(
        n8688) );
  SDFFX1 DFF_207_Q_reg ( .D(n48), .SI(n8688), .SE(n4249), .CLK(n4584), .Q(
        n8687) );
  SDFFX1 DFF_208_Q_reg ( .D(n49), .SI(n8687), .SE(n4249), .CLK(n4584), .Q(
        n8686) );
  SDFFX1 DFF_209_Q_reg ( .D(n50), .SI(n8686), .SE(n4249), .CLK(n4584), .Q(
        n8685) );
  SDFFX1 DFF_210_Q_reg ( .D(n51), .SI(n8685), .SE(n4249), .CLK(n4584), .Q(
        n8684) );
  SDFFX1 DFF_211_Q_reg ( .D(n52), .SI(n8684), .SE(n4250), .CLK(n4584), .Q(
        n8683) );
  SDFFX1 DFF_212_Q_reg ( .D(n53), .SI(n8683), .SE(n4250), .CLK(n4584), .Q(
        n8682) );
  SDFFX1 DFF_213_Q_reg ( .D(n54), .SI(n8682), .SE(n4250), .CLK(n4584), .Q(
        n8681) );
  SDFFX1 DFF_214_Q_reg ( .D(n55), .SI(n8681), .SE(n4250), .CLK(n4584), .Q(
        n8680) );
  SDFFX1 DFF_215_Q_reg ( .D(n56), .SI(n8680), .SE(n4250), .CLK(n4584), .Q(
        test_so12) );
  SDFFX1 DFF_216_Q_reg ( .D(n57), .SI(test_si13), .SE(n4250), .CLK(n4584), .Q(
        n8677) );
  SDFFX1 DFF_217_Q_reg ( .D(n58), .SI(n8677), .SE(n4251), .CLK(n4583), .Q(
        n8676) );
  SDFFX1 DFF_218_Q_reg ( .D(n59), .SI(n8676), .SE(n4251), .CLK(n4583), .Q(
        n8675) );
  SDFFX1 DFF_219_Q_reg ( .D(n60), .SI(n8675), .SE(n4251), .CLK(n4583), .Q(
        n8674) );
  SDFFX1 DFF_220_Q_reg ( .D(n61), .SI(n8674), .SE(n4251), .CLK(n4583), .Q(
        n8673) );
  SDFFX1 DFF_221_Q_reg ( .D(n62), .SI(n8673), .SE(n4251), .CLK(n4583), .Q(
        n8672) );
  SDFFX1 DFF_222_Q_reg ( .D(n63), .SI(n8672), .SE(n4251), .CLK(n4583), .Q(
        n8671) );
  SDFFX1 DFF_223_Q_reg ( .D(WX1839), .SI(n8671), .SE(n4252), .CLK(n4583), .Q(
        n8670) );
  SDFFX1 DFF_224_Q_reg ( .D(WX1937), .SI(n8670), .SE(n4246), .CLK(n4586), .Q(
        n8669), .QN(n7056) );
  SDFFX1 DFF_225_Q_reg ( .D(WX1939), .SI(n8669), .SE(n4246), .CLK(n4586), .Q(
        n8668), .QN(n7057) );
  SDFFX1 DFF_226_Q_reg ( .D(WX1941), .SI(n8668), .SE(n4245), .CLK(n4586), .Q(
        n8667), .QN(n7058) );
  SDFFX1 DFF_227_Q_reg ( .D(WX1943), .SI(n8667), .SE(n4245), .CLK(n4586), .Q(
        n8666), .QN(n7236) );
  SDFFX1 DFF_228_Q_reg ( .D(WX1945), .SI(n8666), .SE(n4244), .CLK(n4587), .Q(
        n8665), .QN(n7059) );
  SDFFX1 DFF_229_Q_reg ( .D(WX1947), .SI(n8665), .SE(n4243), .CLK(n4587), .Q(
        n8664), .QN(n7060) );
  SDFFX1 DFF_230_Q_reg ( .D(WX1949), .SI(n8664), .SE(n4243), .CLK(n4587), .Q(
        n8663), .QN(n7061) );
  SDFFX1 DFF_231_Q_reg ( .D(WX1951), .SI(n8663), .SE(n4242), .CLK(n4588), .Q(
        n8662), .QN(n7062) );
  SDFFX1 DFF_232_Q_reg ( .D(WX1953), .SI(n8662), .SE(n4242), .CLK(n4588), .Q(
        n8661), .QN(n7063) );
  SDFFX1 DFF_233_Q_reg ( .D(WX1955), .SI(n8661), .SE(n3996), .CLK(n4711), .Q(
        test_so13) );
  SDFFX1 DFF_234_Q_reg ( .D(WX1957), .SI(test_si14), .SE(n4240), .CLK(n4589), 
        .Q(n8658), .QN(n7064) );
  SDFFX1 DFF_235_Q_reg ( .D(WX1959), .SI(n8658), .SE(n4240), .CLK(n4589), .Q(
        n8657), .QN(n7065) );
  SDFFX1 DFF_236_Q_reg ( .D(WX1961), .SI(n8657), .SE(n4239), .CLK(n4589), .Q(
        n8656), .QN(n7066) );
  SDFFX1 DFF_237_Q_reg ( .D(WX1963), .SI(n8656), .SE(n4239), .CLK(n4589), .Q(
        n8655), .QN(n7224) );
  SDFFX1 DFF_238_Q_reg ( .D(WX1965), .SI(n8655), .SE(n4003), .CLK(n4707), .Q(
        n8654), .QN(n7067) );
  SDFFX1 DFF_239_Q_reg ( .D(WX1967), .SI(n8654), .SE(n4003), .CLK(n4707), .Q(
        n8653), .QN(n7068) );
  SDFFX1 DFF_240_Q_reg ( .D(WX1969), .SI(n8653), .SE(n3996), .CLK(n4711), .Q(
        WX1970), .QN(n3402) );
  SDFFX1 DFF_241_Q_reg ( .D(WX1971), .SI(WX1970), .SE(n4237), .CLK(n4590), .Q(
        WX1972) );
  SDFFX1 DFF_242_Q_reg ( .D(WX1973), .SI(WX1972), .SE(n4236), .CLK(n4591), .Q(
        WX1974), .QN(n3401) );
  SDFFX1 DFF_243_Q_reg ( .D(WX1975), .SI(WX1974), .SE(n4236), .CLK(n4591), .Q(
        WX1976), .QN(n3400) );
  SDFFX1 DFF_244_Q_reg ( .D(WX1977), .SI(WX1976), .SE(n4236), .CLK(n4591), .Q(
        WX1978), .QN(n3399) );
  SDFFX1 DFF_245_Q_reg ( .D(WX1979), .SI(WX1978), .SE(n4236), .CLK(n4591), .Q(
        WX1980) );
  SDFFX1 DFF_246_Q_reg ( .D(WX1981), .SI(WX1980), .SE(n4236), .CLK(n4591), .Q(
        WX1982), .QN(n3397) );
  SDFFX1 DFF_247_Q_reg ( .D(WX1983), .SI(WX1982), .SE(n4236), .CLK(n4591), .Q(
        WX1984), .QN(n3396) );
  SDFFX1 DFF_248_Q_reg ( .D(WX1985), .SI(WX1984), .SE(n4235), .CLK(n4591), .Q(
        WX1986), .QN(n3395) );
  SDFFX1 DFF_249_Q_reg ( .D(WX1987), .SI(WX1986), .SE(n4235), .CLK(n4591), .Q(
        WX1988), .QN(n3394) );
  SDFFX1 DFF_250_Q_reg ( .D(WX1989), .SI(WX1988), .SE(n4235), .CLK(n4591), .Q(
        WX1990), .QN(n3393) );
  SDFFX1 DFF_251_Q_reg ( .D(WX1991), .SI(WX1990), .SE(n4235), .CLK(n4591), .Q(
        test_so14) );
  SDFFX1 DFF_252_Q_reg ( .D(WX1993), .SI(test_si15), .SE(n4234), .CLK(n4592), 
        .Q(WX1994), .QN(n3392) );
  SDFFX1 DFF_253_Q_reg ( .D(WX1995), .SI(WX1994), .SE(n4234), .CLK(n4592), .Q(
        WX1996), .QN(n3391) );
  SDFFX1 DFF_254_Q_reg ( .D(WX1997), .SI(WX1996), .SE(n4234), .CLK(n4592), .Q(
        WX1998), .QN(n3390) );
  SDFFX1 DFF_255_Q_reg ( .D(WX1999), .SI(WX1998), .SE(n4234), .CLK(n4592), .Q(
        WX2000) );
  SDFFX1 DFF_256_Q_reg ( .D(WX2001), .SI(WX2000), .SE(n4246), .CLK(n4586), .Q(
        WX2002), .QN(n3074) );
  SDFFX1 DFF_257_Q_reg ( .D(WX2003), .SI(WX2002), .SE(n4246), .CLK(n4586), .Q(
        WX2004), .QN(n3287) );
  SDFFX1 DFF_258_Q_reg ( .D(WX2005), .SI(WX2004), .SE(n4245), .CLK(n4586), .Q(
        WX2006), .QN(n3285) );
  SDFFX1 DFF_259_Q_reg ( .D(n67), .SI(WX2006), .SE(n4245), .CLK(n4586), .Q(
        WX2008), .QN(n3284) );
  SDFFX1 DFF_260_Q_reg ( .D(WX2009), .SI(WX2008), .SE(n4244), .CLK(n4587), .Q(
        WX2010), .QN(n3282) );
  SDFFX1 DFF_261_Q_reg ( .D(WX2011), .SI(WX2010), .SE(n4244), .CLK(n4587), .Q(
        WX2012), .QN(n3280) );
  SDFFX1 DFF_262_Q_reg ( .D(WX2013), .SI(WX2012), .SE(n4243), .CLK(n4587), .Q(
        WX2014), .QN(n3277) );
  SDFFX1 DFF_263_Q_reg ( .D(WX2015), .SI(WX2014), .SE(n4242), .CLK(n4588), .Q(
        WX2016), .QN(n3275) );
  SDFFX1 DFF_264_Q_reg ( .D(WX2017), .SI(WX2016), .SE(n4242), .CLK(n4588), .Q(
        WX2018), .QN(n3273) );
  SDFFX1 DFF_265_Q_reg ( .D(WX2019), .SI(WX2018), .SE(n4241), .CLK(n4588), .Q(
        WX2020), .QN(n3272) );
  SDFFX1 DFF_266_Q_reg ( .D(WX2021), .SI(WX2020), .SE(n4241), .CLK(n4588), .Q(
        WX2022), .QN(n3270) );
  SDFFX1 DFF_267_Q_reg ( .D(WX2023), .SI(WX2022), .SE(n4240), .CLK(n4589), .Q(
        WX2024), .QN(n3268) );
  SDFFX1 DFF_268_Q_reg ( .D(WX2025), .SI(WX2024), .SE(n4239), .CLK(n4589), .Q(
        WX2026), .QN(n3266) );
  SDFFX1 DFF_269_Q_reg ( .D(n77), .SI(WX2026), .SE(n4238), .CLK(n4590), .Q(
        test_so15) );
  SDFFX1 DFF_270_Q_reg ( .D(WX2029), .SI(test_si16), .SE(n4003), .CLK(n4707), 
        .Q(WX2030), .QN(n3263) );
  SDFFX1 DFF_271_Q_reg ( .D(WX2031), .SI(WX2030), .SE(n4003), .CLK(n4707), .Q(
        WX2032), .QN(n3261) );
  SDFFX1 DFF_272_Q_reg ( .D(WX2033), .SI(WX2032), .SE(n4002), .CLK(n4708), .Q(
        WX2034), .QN(n3785) );
  SDFFX1 DFF_273_Q_reg ( .D(WX2035), .SI(WX2034), .SE(n4002), .CLK(n4708), .Q(
        WX2036), .QN(n3783) );
  SDFFX1 DFF_274_Q_reg ( .D(WX2037), .SI(WX2036), .SE(n4002), .CLK(n4708), .Q(
        WX2038), .QN(n3781) );
  SDFFX1 DFF_275_Q_reg ( .D(WX2039), .SI(WX2038), .SE(n4002), .CLK(n4708), .Q(
        WX2040), .QN(n3779) );
  SDFFX1 DFF_276_Q_reg ( .D(WX2041), .SI(WX2040), .SE(n4001), .CLK(n4708), .Q(
        WX2042) );
  SDFFX1 DFF_277_Q_reg ( .D(WX2043), .SI(WX2042), .SE(n4001), .CLK(n4708), .Q(
        WX2044), .QN(n3775) );
  SDFFX1 DFF_278_Q_reg ( .D(WX2045), .SI(WX2044), .SE(n4000), .CLK(n4709), .Q(
        WX2046), .QN(n3773) );
  SDFFX1 DFF_279_Q_reg ( .D(WX2047), .SI(WX2046), .SE(n4000), .CLK(n4709), .Q(
        WX2048), .QN(n3771) );
  SDFFX1 DFF_280_Q_reg ( .D(WX2049), .SI(WX2048), .SE(n3999), .CLK(n4709), .Q(
        WX2050), .QN(n3769) );
  SDFFX1 DFF_281_Q_reg ( .D(WX2051), .SI(WX2050), .SE(n3999), .CLK(n4709), .Q(
        WX2052), .QN(n3767) );
  SDFFX1 DFF_282_Q_reg ( .D(WX2053), .SI(WX2052), .SE(n3998), .CLK(n4710), .Q(
        WX2054), .QN(n3765) );
  SDFFX1 DFF_283_Q_reg ( .D(WX2055), .SI(WX2054), .SE(n4235), .CLK(n4591), .Q(
        WX2056), .QN(n3763) );
  SDFFX1 DFF_284_Q_reg ( .D(WX2057), .SI(WX2056), .SE(n4235), .CLK(n4591), .Q(
        WX2058), .QN(n3761) );
  SDFFX1 DFF_285_Q_reg ( .D(WX2059), .SI(WX2058), .SE(n4234), .CLK(n4592), .Q(
        WX2060), .QN(n3759) );
  SDFFX1 DFF_286_Q_reg ( .D(WX2061), .SI(WX2060), .SE(n4234), .CLK(n4592), .Q(
        WX2062), .QN(n3757) );
  SDFFX1 DFF_287_Q_reg ( .D(WX2063), .SI(WX2062), .SE(n4233), .CLK(n4592), .Q(
        test_so16) );
  SDFFX1 DFF_288_Q_reg ( .D(WX2065), .SI(test_si17), .SE(n4246), .CLK(n4586), 
        .Q(WX2066) );
  SDFFX1 DFF_289_Q_reg ( .D(WX2067), .SI(WX2066), .SE(n4246), .CLK(n4586), .Q(
        WX2068) );
  SDFFX1 DFF_290_Q_reg ( .D(WX2069), .SI(WX2068), .SE(n4245), .CLK(n4586), .Q(
        WX2070) );
  SDFFX1 DFF_291_Q_reg ( .D(WX2071), .SI(WX2070), .SE(n4245), .CLK(n4586), .Q(
        WX2072) );
  SDFFX1 DFF_292_Q_reg ( .D(WX2073), .SI(WX2072), .SE(n4244), .CLK(n4587), .Q(
        WX2074) );
  SDFFX1 DFF_293_Q_reg ( .D(WX2075), .SI(WX2074), .SE(n4244), .CLK(n4587), .Q(
        WX2076) );
  SDFFX1 DFF_294_Q_reg ( .D(WX2077), .SI(WX2076), .SE(n4243), .CLK(n4587), .Q(
        WX2078) );
  SDFFX1 DFF_295_Q_reg ( .D(WX2079), .SI(WX2078), .SE(n4242), .CLK(n4588), .Q(
        WX2080) );
  SDFFX1 DFF_296_Q_reg ( .D(WX2081), .SI(WX2080), .SE(n4241), .CLK(n4588), .Q(
        WX2082) );
  SDFFX1 DFF_297_Q_reg ( .D(WX2083), .SI(WX2082), .SE(n4241), .CLK(n4588), .Q(
        WX2084), .QN(n7229) );
  SDFFX1 DFF_298_Q_reg ( .D(WX2085), .SI(WX2084), .SE(n4240), .CLK(n4589), .Q(
        WX2086) );
  SDFFX1 DFF_299_Q_reg ( .D(WX2087), .SI(WX2086), .SE(n4240), .CLK(n4589), .Q(
        WX2088) );
  SDFFX1 DFF_300_Q_reg ( .D(WX2089), .SI(WX2088), .SE(n4239), .CLK(n4589), .Q(
        WX2090) );
  SDFFX1 DFF_301_Q_reg ( .D(WX2091), .SI(WX2090), .SE(n4238), .CLK(n4590), .Q(
        WX2092), .QN(n3265) );
  SDFFX1 DFF_302_Q_reg ( .D(WX2093), .SI(WX2092), .SE(n4238), .CLK(n4590), .Q(
        WX2094) );
  SDFFX1 DFF_303_Q_reg ( .D(WX2095), .SI(WX2094), .SE(n4238), .CLK(n4590), .Q(
        WX2096) );
  SDFFX1 DFF_304_Q_reg ( .D(WX2097), .SI(WX2096), .SE(n4237), .CLK(n4590), .Q(
        WX2098) );
  SDFFX1 DFF_305_Q_reg ( .D(WX2099), .SI(WX2098), .SE(n4237), .CLK(n4590), .Q(
        test_so17) );
  SDFFX1 DFF_306_Q_reg ( .D(WX2101), .SI(test_si18), .SE(n4002), .CLK(n4708), 
        .Q(WX2102) );
  SDFFX1 DFF_307_Q_reg ( .D(WX2103), .SI(WX2102), .SE(n4001), .CLK(n4708), .Q(
        WX2104) );
  SDFFX1 DFF_308_Q_reg ( .D(WX2105), .SI(WX2104), .SE(n4001), .CLK(n4708), .Q(
        WX2106), .QN(n7218) );
  SDFFX1 DFF_309_Q_reg ( .D(WX2107), .SI(WX2106), .SE(n4000), .CLK(n4709), .Q(
        WX2108), .QN(n3398) );
  SDFFX1 DFF_310_Q_reg ( .D(WX2109), .SI(WX2108), .SE(n4000), .CLK(n4709), .Q(
        WX2110) );
  SDFFX1 DFF_311_Q_reg ( .D(WX2111), .SI(WX2110), .SE(n3999), .CLK(n4709), .Q(
        WX2112) );
  SDFFX1 DFF_312_Q_reg ( .D(WX2113), .SI(WX2112), .SE(n3999), .CLK(n4709), .Q(
        WX2114) );
  SDFFX1 DFF_313_Q_reg ( .D(WX2115), .SI(WX2114), .SE(n3998), .CLK(n4710), .Q(
        WX2116) );
  SDFFX1 DFF_314_Q_reg ( .D(WX2117), .SI(WX2116), .SE(n3998), .CLK(n4710), .Q(
        WX2118) );
  SDFFX1 DFF_315_Q_reg ( .D(WX2119), .SI(WX2118), .SE(n3998), .CLK(n4710), .Q(
        WX2120) );
  SDFFX1 DFF_316_Q_reg ( .D(WX2121), .SI(WX2120), .SE(n3997), .CLK(n4710), .Q(
        WX2122) );
  SDFFX1 DFF_317_Q_reg ( .D(WX2123), .SI(WX2122), .SE(n3997), .CLK(n4710), .Q(
        WX2124) );
  SDFFX1 DFF_318_Q_reg ( .D(WX2125), .SI(WX2124), .SE(n3997), .CLK(n4710), .Q(
        WX2126) );
  SDFFX1 DFF_319_Q_reg ( .D(WX2127), .SI(WX2126), .SE(n4233), .CLK(n4592), .Q(
        WX2128), .QN(n3389) );
  SDFFX1 DFF_320_Q_reg ( .D(WX2129), .SI(WX2128), .SE(n4233), .CLK(n4592), .Q(
        WX2130), .QN(n3768) );
  SDFFX1 DFF_321_Q_reg ( .D(WX2131), .SI(WX2130), .SE(n4233), .CLK(n4592), .Q(
        WX2132), .QN(n3770) );
  SDFFX1 DFF_322_Q_reg ( .D(WX2133), .SI(WX2132), .SE(n4233), .CLK(n4592), .Q(
        WX2134), .QN(n3772) );
  SDFFX1 DFF_323_Q_reg ( .D(WX2135), .SI(WX2134), .SE(n4233), .CLK(n4592), .Q(
        test_so18) );
  SDFFX1 DFF_324_Q_reg ( .D(WX2137), .SI(test_si19), .SE(n4244), .CLK(n4587), 
        .Q(WX2138), .QN(n3774) );
  SDFFX1 DFF_325_Q_reg ( .D(WX2139), .SI(WX2138), .SE(n4243), .CLK(n4587), .Q(
        WX2140), .QN(n3776) );
  SDFFX1 DFF_326_Q_reg ( .D(WX2141), .SI(WX2140), .SE(n4243), .CLK(n4587), .Q(
        WX2142), .QN(n3778) );
  SDFFX1 DFF_327_Q_reg ( .D(WX2143), .SI(WX2142), .SE(n4242), .CLK(n4588), .Q(
        WX2144), .QN(n3780) );
  SDFFX1 DFF_328_Q_reg ( .D(WX2145), .SI(WX2144), .SE(n4241), .CLK(n4588), .Q(
        WX2146), .QN(n3782) );
  SDFFX1 DFF_329_Q_reg ( .D(WX2147), .SI(WX2146), .SE(n4241), .CLK(n4588), .Q(
        WX2148), .QN(n3784) );
  SDFFX1 DFF_330_Q_reg ( .D(WX2149), .SI(WX2148), .SE(n4240), .CLK(n4589), .Q(
        WX2150), .QN(n3786) );
  SDFFX1 DFF_331_Q_reg ( .D(WX2151), .SI(WX2150), .SE(n4239), .CLK(n4589), .Q(
        WX2152), .QN(n3787) );
  SDFFX1 DFF_332_Q_reg ( .D(WX2153), .SI(WX2152), .SE(n4239), .CLK(n4589), .Q(
        WX2154), .QN(n3788) );
  SDFFX1 DFF_333_Q_reg ( .D(WX2155), .SI(WX2154), .SE(n4238), .CLK(n4590), .Q(
        WX2156), .QN(n3789) );
  SDFFX1 DFF_334_Q_reg ( .D(WX2157), .SI(WX2156), .SE(n4238), .CLK(n4590), .Q(
        WX2158), .QN(n3790) );
  SDFFX1 DFF_335_Q_reg ( .D(WX2159), .SI(WX2158), .SE(n4237), .CLK(n4590), .Q(
        WX2160), .QN(n3430) );
  SDFFX1 DFF_336_Q_reg ( .D(WX2161), .SI(WX2160), .SE(n4237), .CLK(n4590), .Q(
        WX2162), .QN(n3791) );
  SDFFX1 DFF_337_Q_reg ( .D(WX2163), .SI(WX2162), .SE(n4237), .CLK(n4590), .Q(
        WX2164), .QN(n3792) );
  SDFFX1 DFF_338_Q_reg ( .D(WX2165), .SI(WX2164), .SE(n4002), .CLK(n4708), .Q(
        WX2166), .QN(n3793) );
  SDFFX1 DFF_339_Q_reg ( .D(WX2167), .SI(WX2166), .SE(n4001), .CLK(n4708), .Q(
        WX2168), .QN(n3794) );
  SDFFX1 DFF_340_Q_reg ( .D(WX2169), .SI(WX2168), .SE(n4001), .CLK(n4708), .Q(
        WX2170), .QN(n3431) );
  SDFFX1 DFF_341_Q_reg ( .D(WX2171), .SI(WX2170), .SE(n4000), .CLK(n4709), .Q(
        test_so19) );
  SDFFX1 DFF_342_Q_reg ( .D(WX2173), .SI(test_si20), .SE(n4000), .CLK(n4709), 
        .Q(WX2174), .QN(n3795) );
  SDFFX1 DFF_343_Q_reg ( .D(WX2175), .SI(WX2174), .SE(n3999), .CLK(n4709), .Q(
        WX2176), .QN(n3796) );
  SDFFX1 DFF_344_Q_reg ( .D(WX2177), .SI(WX2176), .SE(n3999), .CLK(n4709), .Q(
        WX2178), .QN(n3797) );
  SDFFX1 DFF_345_Q_reg ( .D(WX2179), .SI(WX2178), .SE(n3998), .CLK(n4710), .Q(
        WX2180), .QN(n3798) );
  SDFFX1 DFF_346_Q_reg ( .D(WX2181), .SI(WX2180), .SE(n3998), .CLK(n4710), .Q(
        WX2182), .QN(n3799) );
  SDFFX1 DFF_347_Q_reg ( .D(WX2183), .SI(WX2182), .SE(n3997), .CLK(n4710), .Q(
        WX2184), .QN(n3432) );
  SDFFX1 DFF_348_Q_reg ( .D(WX2185), .SI(WX2184), .SE(n3997), .CLK(n4710), .Q(
        WX2186), .QN(n3800) );
  SDFFX1 DFF_349_Q_reg ( .D(WX2187), .SI(WX2186), .SE(n3997), .CLK(n4710), .Q(
        WX2188), .QN(n3801) );
  SDFFX1 DFF_350_Q_reg ( .D(WX2189), .SI(WX2188), .SE(n3996), .CLK(n4711), .Q(
        WX2190), .QN(n3802) );
  SDFFX1 DFF_351_Q_reg ( .D(WX2191), .SI(WX2190), .SE(n3996), .CLK(n4711), .Q(
        WX2192), .QN(n3440) );
  SDFFX1 DFF_352_Q_reg ( .D(WX2557), .SI(WX2192), .SE(n4008), .CLK(n4705), .Q(
        CRC_OUT_8_0), .QN(DFF_352_n1) );
  SDFFX1 DFF_353_Q_reg ( .D(WX2559), .SI(CRC_OUT_8_0), .SE(n4008), .CLK(n4705), 
        .Q(CRC_OUT_8_1), .QN(DFF_353_n1) );
  SDFFX1 DFF_354_Q_reg ( .D(WX2561), .SI(CRC_OUT_8_1), .SE(n4008), .CLK(n4705), 
        .Q(CRC_OUT_8_2), .QN(DFF_354_n1) );
  SDFFX1 DFF_355_Q_reg ( .D(WX2563), .SI(CRC_OUT_8_2), .SE(n4008), .CLK(n4705), 
        .Q(CRC_OUT_8_3) );
  SDFFX1 DFF_356_Q_reg ( .D(WX2565), .SI(CRC_OUT_8_3), .SE(n4008), .CLK(n4705), 
        .Q(CRC_OUT_8_4), .QN(DFF_356_n1) );
  SDFFX1 DFF_357_Q_reg ( .D(WX2567), .SI(CRC_OUT_8_4), .SE(n4007), .CLK(n4705), 
        .Q(CRC_OUT_8_5), .QN(DFF_357_n1) );
  SDFFX1 DFF_358_Q_reg ( .D(WX2569), .SI(CRC_OUT_8_5), .SE(n4007), .CLK(n4705), 
        .Q(CRC_OUT_8_6), .QN(DFF_358_n1) );
  SDFFX1 DFF_359_Q_reg ( .D(WX2571), .SI(CRC_OUT_8_6), .SE(n4007), .CLK(n4705), 
        .Q(test_so20) );
  SDFFX1 DFF_360_Q_reg ( .D(WX2573), .SI(test_si21), .SE(n4007), .CLK(n4705), 
        .Q(CRC_OUT_8_8), .QN(DFF_360_n1) );
  SDFFX1 DFF_361_Q_reg ( .D(WX2575), .SI(CRC_OUT_8_8), .SE(n4007), .CLK(n4705), 
        .Q(CRC_OUT_8_9) );
  SDFFX1 DFF_362_Q_reg ( .D(WX2577), .SI(CRC_OUT_8_9), .SE(n4007), .CLK(n4705), 
        .Q(CRC_OUT_8_10) );
  SDFFX1 DFF_363_Q_reg ( .D(WX2579), .SI(CRC_OUT_8_10), .SE(n4006), .CLK(n4706), .Q(CRC_OUT_8_11), .QN(DFF_363_n1) );
  SDFFX1 DFF_364_Q_reg ( .D(WX2581), .SI(CRC_OUT_8_11), .SE(n4006), .CLK(n4706), .Q(CRC_OUT_8_12), .QN(DFF_364_n1) );
  SDFFX1 DFF_365_Q_reg ( .D(WX2583), .SI(CRC_OUT_8_12), .SE(n4006), .CLK(n4706), .Q(CRC_OUT_8_13), .QN(DFF_365_n1) );
  SDFFX1 DFF_366_Q_reg ( .D(WX2585), .SI(CRC_OUT_8_13), .SE(n4006), .CLK(n4706), .Q(CRC_OUT_8_14), .QN(DFF_366_n1) );
  SDFFX1 DFF_367_Q_reg ( .D(WX2587), .SI(CRC_OUT_8_14), .SE(n4006), .CLK(n4706), .Q(CRC_OUT_8_15) );
  SDFFX1 DFF_368_Q_reg ( .D(WX2589), .SI(CRC_OUT_8_15), .SE(n4006), .CLK(n4706), .Q(CRC_OUT_8_16), .QN(DFF_368_n1) );
  SDFFX1 DFF_369_Q_reg ( .D(WX2591), .SI(CRC_OUT_8_16), .SE(n4005), .CLK(n4706), .Q(CRC_OUT_8_17), .QN(DFF_369_n1) );
  SDFFX1 DFF_370_Q_reg ( .D(WX2593), .SI(CRC_OUT_8_17), .SE(n4005), .CLK(n4706), .Q(CRC_OUT_8_18), .QN(DFF_370_n1) );
  SDFFX1 DFF_371_Q_reg ( .D(WX2595), .SI(CRC_OUT_8_18), .SE(n4005), .CLK(n4706), .Q(CRC_OUT_8_19), .QN(DFF_371_n1) );
  SDFFX1 DFF_372_Q_reg ( .D(WX2597), .SI(CRC_OUT_8_19), .SE(n4005), .CLK(n4706), .Q(CRC_OUT_8_20), .QN(DFF_372_n1) );
  SDFFX1 DFF_373_Q_reg ( .D(WX2599), .SI(CRC_OUT_8_20), .SE(n4005), .CLK(n4706), .Q(CRC_OUT_8_21), .QN(DFF_373_n1) );
  SDFFX1 DFF_374_Q_reg ( .D(WX2601), .SI(CRC_OUT_8_21), .SE(n4005), .CLK(n4706), .Q(CRC_OUT_8_22), .QN(DFF_374_n1) );
  SDFFX1 DFF_375_Q_reg ( .D(WX2603), .SI(CRC_OUT_8_22), .SE(n4004), .CLK(n4707), .Q(CRC_OUT_8_23), .QN(DFF_375_n1) );
  SDFFX1 DFF_376_Q_reg ( .D(WX2605), .SI(CRC_OUT_8_23), .SE(n4004), .CLK(n4707), .Q(CRC_OUT_8_24), .QN(DFF_376_n1) );
  SDFFX1 DFF_377_Q_reg ( .D(WX2607), .SI(CRC_OUT_8_24), .SE(n4004), .CLK(n4707), .Q(test_so21) );
  SDFFX1 DFF_378_Q_reg ( .D(WX2609), .SI(test_si22), .SE(n4004), .CLK(n4707), 
        .Q(CRC_OUT_8_26), .QN(DFF_378_n1) );
  SDFFX1 DFF_379_Q_reg ( .D(WX2611), .SI(CRC_OUT_8_26), .SE(n4004), .CLK(n4707), .Q(CRC_OUT_8_27) );
  SDFFX1 DFF_380_Q_reg ( .D(WX2613), .SI(CRC_OUT_8_27), .SE(n4004), .CLK(n4707), .Q(CRC_OUT_8_28), .QN(DFF_380_n1) );
  SDFFX1 DFF_381_Q_reg ( .D(WX2615), .SI(CRC_OUT_8_28), .SE(n4003), .CLK(n4707), .Q(CRC_OUT_8_29), .QN(DFF_381_n1) );
  SDFFX1 DFF_382_Q_reg ( .D(WX2617), .SI(CRC_OUT_8_29), .SE(n4003), .CLK(n4707), .Q(CRC_OUT_8_30), .QN(DFF_382_n1) );
  SDFFX1 DFF_383_Q_reg ( .D(WX2619), .SI(CRC_OUT_8_30), .SE(n4232), .CLK(n4593), .Q(CRC_OUT_8_31), .QN(DFF_383_n1) );
  SDFFX1 DFF_384_Q_reg ( .D(n111), .SI(CRC_OUT_8_31), .SE(n4232), .CLK(n4593), 
        .Q(WX3071) );
  SDFFX1 DFF_385_Q_reg ( .D(n112), .SI(WX3071), .SE(n4227), .CLK(n4595), .Q(
        n8644) );
  SDFFX1 DFF_386_Q_reg ( .D(n113), .SI(n8644), .SE(n4227), .CLK(n4595), .Q(
        n8643) );
  SDFFX1 DFF_387_Q_reg ( .D(n114), .SI(n8643), .SE(n4227), .CLK(n4595), .Q(
        n8642) );
  SDFFX1 DFF_388_Q_reg ( .D(n115), .SI(n8642), .SE(n4228), .CLK(n4595), .Q(
        n8641) );
  SDFFX1 DFF_389_Q_reg ( .D(n116), .SI(n8641), .SE(n4228), .CLK(n4595), .Q(
        n8640) );
  SDFFX1 DFF_390_Q_reg ( .D(n117), .SI(n8640), .SE(n4228), .CLK(n4595), .Q(
        n8639) );
  SDFFX1 DFF_391_Q_reg ( .D(n118), .SI(n8639), .SE(n4228), .CLK(n4595), .Q(
        n8638) );
  SDFFX1 DFF_392_Q_reg ( .D(n119), .SI(n8638), .SE(n4228), .CLK(n4595), .Q(
        n8637) );
  SDFFX1 DFF_393_Q_reg ( .D(n120), .SI(n8637), .SE(n4228), .CLK(n4595), .Q(
        n8636) );
  SDFFX1 DFF_394_Q_reg ( .D(n121), .SI(n8636), .SE(n4229), .CLK(n4594), .Q(
        n8635) );
  SDFFX1 DFF_395_Q_reg ( .D(n122), .SI(n8635), .SE(n4229), .CLK(n4594), .Q(
        test_so22) );
  SDFFX1 DFF_396_Q_reg ( .D(n123), .SI(test_si23), .SE(n4229), .CLK(n4594), 
        .Q(n8632) );
  SDFFX1 DFF_397_Q_reg ( .D(n124), .SI(n8632), .SE(n4229), .CLK(n4594), .Q(
        n8631) );
  SDFFX1 DFF_398_Q_reg ( .D(n125), .SI(n8631), .SE(n4229), .CLK(n4594), .Q(
        n8630) );
  SDFFX1 DFF_399_Q_reg ( .D(n126), .SI(n8630), .SE(n4229), .CLK(n4594), .Q(
        n8629) );
  SDFFX1 DFF_400_Q_reg ( .D(n128), .SI(n8629), .SE(n4230), .CLK(n4594), .Q(
        n8628) );
  SDFFX1 DFF_401_Q_reg ( .D(n129), .SI(n8628), .SE(n4230), .CLK(n4594), .Q(
        n8627) );
  SDFFX1 DFF_402_Q_reg ( .D(n130), .SI(n8627), .SE(n4230), .CLK(n4594), .Q(
        n8626) );
  SDFFX1 DFF_403_Q_reg ( .D(n131), .SI(n8626), .SE(n4230), .CLK(n4594), .Q(
        n8625) );
  SDFFX1 DFF_404_Q_reg ( .D(n132), .SI(n8625), .SE(n4230), .CLK(n4594), .Q(
        n8624) );
  SDFFX1 DFF_405_Q_reg ( .D(n133), .SI(n8624), .SE(n4230), .CLK(n4594), .Q(
        n8623) );
  SDFFX1 DFF_406_Q_reg ( .D(n134), .SI(n8623), .SE(n4231), .CLK(n4593), .Q(
        n8622) );
  SDFFX1 DFF_407_Q_reg ( .D(n135), .SI(n8622), .SE(n4231), .CLK(n4593), .Q(
        n8621) );
  SDFFX1 DFF_408_Q_reg ( .D(n136), .SI(n8621), .SE(n4231), .CLK(n4593), .Q(
        n8620) );
  SDFFX1 DFF_409_Q_reg ( .D(n137), .SI(n8620), .SE(n4231), .CLK(n4593), .Q(
        n8619) );
  SDFFX1 DFF_410_Q_reg ( .D(n138), .SI(n8619), .SE(n4231), .CLK(n4593), .Q(
        n8618) );
  SDFFX1 DFF_411_Q_reg ( .D(n139), .SI(n8618), .SE(n4231), .CLK(n4593), .Q(
        n8617) );
  SDFFX1 DFF_412_Q_reg ( .D(n140), .SI(n8617), .SE(n4232), .CLK(n4593), .Q(
        n8616) );
  SDFFX1 DFF_413_Q_reg ( .D(n141), .SI(n8616), .SE(n4232), .CLK(n4593), .Q(
        test_so23) );
  SDFFX1 DFF_414_Q_reg ( .D(n142), .SI(test_si24), .SE(n4232), .CLK(n4593), 
        .Q(n8613) );
  SDFFX1 DFF_415_Q_reg ( .D(WX3132), .SI(n8613), .SE(n4232), .CLK(n4593), .Q(
        n8612) );
  SDFFX1 DFF_416_Q_reg ( .D(WX3230), .SI(n8612), .SE(n4227), .CLK(n4595), .Q(
        n8611), .QN(n7239) );
  SDFFX1 DFF_417_Q_reg ( .D(WX3232), .SI(n8611), .SE(n4226), .CLK(n4596), .Q(
        n8610), .QN(n7238) );
  SDFFX1 DFF_418_Q_reg ( .D(WX3234), .SI(n8610), .SE(n4226), .CLK(n4596), .Q(
        n8609), .QN(n7237) );
  SDFFX1 DFF_419_Q_reg ( .D(WX3236), .SI(n8609), .SE(n4226), .CLK(n4596), .Q(
        n8608), .QN(n7235) );
  SDFFX1 DFF_420_Q_reg ( .D(WX3238), .SI(n8608), .SE(n4226), .CLK(n4596), .Q(
        n8607), .QN(n7234) );
  SDFFX1 DFF_421_Q_reg ( .D(WX3240), .SI(n8607), .SE(n4225), .CLK(n4596), .Q(
        n8606), .QN(n7233) );
  SDFFX1 DFF_422_Q_reg ( .D(WX3242), .SI(n8606), .SE(n4225), .CLK(n4596), .Q(
        n8605), .QN(n7232) );
  SDFFX1 DFF_423_Q_reg ( .D(WX3244), .SI(n8605), .SE(n4224), .CLK(n4597), .Q(
        n8604), .QN(n7231) );
  SDFFX1 DFF_424_Q_reg ( .D(WX3246), .SI(n8604), .SE(n4224), .CLK(n4597), .Q(
        n8603), .QN(n7230) );
  SDFFX1 DFF_425_Q_reg ( .D(WX3248), .SI(n8603), .SE(n4223), .CLK(n4597), .Q(
        n8602), .QN(n7228) );
  SDFFX1 DFF_426_Q_reg ( .D(WX3250), .SI(n8602), .SE(n4223), .CLK(n4597), .Q(
        n8601), .QN(n7227) );
  SDFFX1 DFF_427_Q_reg ( .D(WX3252), .SI(n8601), .SE(n4222), .CLK(n4598), .Q(
        n8600), .QN(n7226) );
  SDFFX1 DFF_428_Q_reg ( .D(WX3254), .SI(n8600), .SE(n4221), .CLK(n4598), .Q(
        n8599), .QN(n7225) );
  SDFFX1 DFF_429_Q_reg ( .D(WX3256), .SI(n8599), .SE(n4220), .CLK(n4599), .Q(
        n8598), .QN(n7223) );
  SDFFX1 DFF_430_Q_reg ( .D(WX3258), .SI(n8598), .SE(n4220), .CLK(n4599), .Q(
        n8597), .QN(n7222) );
  SDFFX1 DFF_431_Q_reg ( .D(WX3260), .SI(n8597), .SE(n4219), .CLK(n4599), .Q(
        test_so24) );
  SDFFX1 DFF_432_Q_reg ( .D(WX3262), .SI(test_si25), .SE(n4014), .CLK(n4702), 
        .Q(WX3263), .QN(n3388) );
  SDFFX1 DFF_433_Q_reg ( .D(WX3264), .SI(WX3263), .SE(n4216), .CLK(n4601), .Q(
        WX3265), .QN(n3387) );
  SDFFX1 DFF_434_Q_reg ( .D(WX3266), .SI(WX3265), .SE(n4216), .CLK(n4601), .Q(
        WX3267), .QN(n3386) );
  SDFFX1 DFF_435_Q_reg ( .D(WX3268), .SI(WX3267), .SE(n4216), .CLK(n4601), .Q(
        WX3269) );
  SDFFX1 DFF_436_Q_reg ( .D(WX3270), .SI(WX3269), .SE(n4216), .CLK(n4601), .Q(
        WX3271), .QN(n3384) );
  SDFFX1 DFF_437_Q_reg ( .D(WX3272), .SI(WX3271), .SE(n4216), .CLK(n4601), .Q(
        WX3273), .QN(n3383) );
  SDFFX1 DFF_438_Q_reg ( .D(WX3274), .SI(WX3273), .SE(n4215), .CLK(n4601), .Q(
        WX3275), .QN(n3382) );
  SDFFX1 DFF_439_Q_reg ( .D(WX3276), .SI(WX3275), .SE(n4215), .CLK(n4601), .Q(
        WX3277) );
  SDFFX1 DFF_440_Q_reg ( .D(WX3278), .SI(WX3277), .SE(n4215), .CLK(n4601), .Q(
        WX3279), .QN(n3381) );
  SDFFX1 DFF_441_Q_reg ( .D(WX3280), .SI(WX3279), .SE(n4214), .CLK(n4602), .Q(
        WX3281) );
  SDFFX1 DFF_442_Q_reg ( .D(WX3282), .SI(WX3281), .SE(n4214), .CLK(n4602), .Q(
        WX3283), .QN(n3379) );
  SDFFX1 DFF_443_Q_reg ( .D(WX3284), .SI(WX3283), .SE(n4213), .CLK(n4602), .Q(
        WX3285), .QN(n3378) );
  SDFFX1 DFF_444_Q_reg ( .D(WX3286), .SI(WX3285), .SE(n4212), .CLK(n4603), .Q(
        WX3287), .QN(n3377) );
  SDFFX1 DFF_445_Q_reg ( .D(WX3288), .SI(WX3287), .SE(n4212), .CLK(n4603), .Q(
        WX3289), .QN(n3376) );
  SDFFX1 DFF_446_Q_reg ( .D(WX3290), .SI(WX3289), .SE(n4211), .CLK(n4603), .Q(
        WX3291), .QN(n3375) );
  SDFFX1 DFF_447_Q_reg ( .D(WX3292), .SI(WX3291), .SE(n4210), .CLK(n4604), .Q(
        WX3293), .QN(n3374) );
  SDFFX1 DFF_448_Q_reg ( .D(n143), .SI(WX3293), .SE(n4227), .CLK(n4595), .Q(
        WX3295), .QN(n3072) );
  SDFFX1 DFF_449_Q_reg ( .D(n144), .SI(WX3295), .SE(n4227), .CLK(n4595), .Q(
        test_so25) );
  SDFFX1 DFF_450_Q_reg ( .D(n145), .SI(test_si26), .SE(n4226), .CLK(n4596), 
        .Q(WX3299), .QN(n3258) );
  SDFFX1 DFF_451_Q_reg ( .D(n146), .SI(WX3299), .SE(n4226), .CLK(n4596), .Q(
        WX3301), .QN(n3256) );
  SDFFX1 DFF_452_Q_reg ( .D(n147), .SI(WX3301), .SE(n4225), .CLK(n4596), .Q(
        WX3303), .QN(n3254) );
  SDFFX1 DFF_453_Q_reg ( .D(n148), .SI(WX3303), .SE(n4225), .CLK(n4596), .Q(
        WX3305), .QN(n3253) );
  SDFFX1 DFF_454_Q_reg ( .D(n149), .SI(WX3305), .SE(n4225), .CLK(n4596), .Q(
        WX3307), .QN(n3251) );
  SDFFX1 DFF_455_Q_reg ( .D(n150), .SI(WX3307), .SE(n4224), .CLK(n4597), .Q(
        WX3309), .QN(n3249) );
  SDFFX1 DFF_456_Q_reg ( .D(n151), .SI(WX3309), .SE(n4224), .CLK(n4597), .Q(
        WX3311), .QN(n3248) );
  SDFFX1 DFF_457_Q_reg ( .D(n152), .SI(WX3311), .SE(n4223), .CLK(n4597), .Q(
        WX3313), .QN(n3246) );
  SDFFX1 DFF_458_Q_reg ( .D(n153), .SI(WX3313), .SE(n4223), .CLK(n4597), .Q(
        WX3315), .QN(n3244) );
  SDFFX1 DFF_459_Q_reg ( .D(n154), .SI(WX3315), .SE(n4222), .CLK(n4598), .Q(
        WX3317), .QN(n3242) );
  SDFFX1 DFF_460_Q_reg ( .D(n155), .SI(WX3317), .SE(n4221), .CLK(n4598), .Q(
        WX3319), .QN(n3240) );
  SDFFX1 DFF_461_Q_reg ( .D(n156), .SI(WX3319), .SE(n4221), .CLK(n4598), .Q(
        WX3321), .QN(n3238) );
  SDFFX1 DFF_462_Q_reg ( .D(n157), .SI(WX3321), .SE(n4220), .CLK(n4599), .Q(
        WX3323), .QN(n3236) );
  SDFFX1 DFF_463_Q_reg ( .D(n158), .SI(WX3323), .SE(n4219), .CLK(n4599), .Q(
        WX3325), .QN(n3235) );
  SDFFX1 DFF_464_Q_reg ( .D(WX3326), .SI(WX3325), .SE(n4014), .CLK(n4702), .Q(
        WX3327) );
  SDFFX1 DFF_465_Q_reg ( .D(WX3328), .SI(WX3327), .SE(n4013), .CLK(n4702), .Q(
        WX3329) );
  SDFFX1 DFF_466_Q_reg ( .D(WX3330), .SI(WX3329), .SE(n4013), .CLK(n4702), .Q(
        WX3331), .QN(n3749) );
  SDFFX1 DFF_467_Q_reg ( .D(WX3332), .SI(WX3331), .SE(n4012), .CLK(n4703), .Q(
        test_so26) );
  SDFFX1 DFF_468_Q_reg ( .D(WX3334), .SI(test_si27), .SE(n4216), .CLK(n4601), 
        .Q(WX3335) );
  SDFFX1 DFF_469_Q_reg ( .D(WX3336), .SI(WX3335), .SE(n4215), .CLK(n4601), .Q(
        WX3337), .QN(n3743) );
  SDFFX1 DFF_470_Q_reg ( .D(WX3338), .SI(WX3337), .SE(n4215), .CLK(n4601), .Q(
        WX3339), .QN(n3741) );
  SDFFX1 DFF_471_Q_reg ( .D(WX3340), .SI(WX3339), .SE(n4215), .CLK(n4601), .Q(
        WX3341), .QN(n3739) );
  SDFFX1 DFF_472_Q_reg ( .D(WX3342), .SI(WX3341), .SE(n4214), .CLK(n4602), .Q(
        WX3343), .QN(n3737) );
  SDFFX1 DFF_473_Q_reg ( .D(WX3344), .SI(WX3343), .SE(n4214), .CLK(n4602), .Q(
        WX3345), .QN(n3735) );
  SDFFX1 DFF_474_Q_reg ( .D(WX3346), .SI(WX3345), .SE(n4213), .CLK(n4602), .Q(
        WX3347), .QN(n3733) );
  SDFFX1 DFF_475_Q_reg ( .D(WX3348), .SI(WX3347), .SE(n4213), .CLK(n4602), .Q(
        WX3349) );
  SDFFX1 DFF_476_Q_reg ( .D(WX3350), .SI(WX3349), .SE(n4212), .CLK(n4603), .Q(
        WX3351), .QN(n3729) );
  SDFFX1 DFF_477_Q_reg ( .D(WX3352), .SI(WX3351), .SE(n4211), .CLK(n4603), .Q(
        WX3353), .QN(n3727) );
  SDFFX1 DFF_478_Q_reg ( .D(WX3354), .SI(WX3353), .SE(n4211), .CLK(n4603), .Q(
        WX3355), .QN(n3725) );
  SDFFX1 DFF_479_Q_reg ( .D(WX3356), .SI(WX3355), .SE(n4210), .CLK(n4604), .Q(
        WX3357) );
  SDFFX1 DFF_480_Q_reg ( .D(WX3358), .SI(WX3357), .SE(n4210), .CLK(n4604), .Q(
        WX3359) );
  SDFFX1 DFF_481_Q_reg ( .D(WX3360), .SI(WX3359), .SE(n4209), .CLK(n4604), .Q(
        WX3361), .QN(n3260) );
  SDFFX1 DFF_482_Q_reg ( .D(WX3362), .SI(WX3361), .SE(n4209), .CLK(n4604), .Q(
        WX3363) );
  SDFFX1 DFF_483_Q_reg ( .D(WX3364), .SI(WX3363), .SE(n4209), .CLK(n4604), .Q(
        WX3365) );
  SDFFX1 DFF_484_Q_reg ( .D(WX3366), .SI(WX3365), .SE(n4208), .CLK(n4605), .Q(
        WX3367) );
  SDFFX1 DFF_485_Q_reg ( .D(WX3368), .SI(WX3367), .SE(n4208), .CLK(n4605), .Q(
        test_so27) );
  SDFFX1 DFF_486_Q_reg ( .D(WX3370), .SI(test_si28), .SE(n4225), .CLK(n4596), 
        .Q(WX3371) );
  SDFFX1 DFF_487_Q_reg ( .D(WX3372), .SI(WX3371), .SE(n4224), .CLK(n4597), .Q(
        WX3373) );
  SDFFX1 DFF_488_Q_reg ( .D(WX3374), .SI(WX3373), .SE(n4224), .CLK(n4597), .Q(
        WX3375) );
  SDFFX1 DFF_489_Q_reg ( .D(WX3376), .SI(WX3375), .SE(n4223), .CLK(n4597), .Q(
        WX3377) );
  SDFFX1 DFF_490_Q_reg ( .D(WX3378), .SI(WX3377), .SE(n4222), .CLK(n4598), .Q(
        WX3379) );
  SDFFX1 DFF_491_Q_reg ( .D(WX3380), .SI(WX3379), .SE(n4222), .CLK(n4598), .Q(
        WX3381) );
  SDFFX1 DFF_492_Q_reg ( .D(WX3382), .SI(WX3381), .SE(n4221), .CLK(n4598), .Q(
        WX3383) );
  SDFFX1 DFF_493_Q_reg ( .D(WX3384), .SI(WX3383), .SE(n4221), .CLK(n4598), .Q(
        WX3385) );
  SDFFX1 DFF_494_Q_reg ( .D(WX3386), .SI(WX3385), .SE(n4220), .CLK(n4599), .Q(
        WX3387) );
  SDFFX1 DFF_495_Q_reg ( .D(WX3388), .SI(WX3387), .SE(n4219), .CLK(n4599), .Q(
        WX3389), .QN(n7221) );
  SDFFX1 DFF_496_Q_reg ( .D(WX3390), .SI(WX3389), .SE(n4013), .CLK(n4702), .Q(
        WX3391), .QN(n7220) );
  SDFFX1 DFF_497_Q_reg ( .D(WX3392), .SI(WX3391), .SE(n4013), .CLK(n4702), .Q(
        WX3393), .QN(n7219) );
  SDFFX1 DFF_498_Q_reg ( .D(WX3394), .SI(WX3393), .SE(n4012), .CLK(n4703), .Q(
        WX3395) );
  SDFFX1 DFF_499_Q_reg ( .D(WX3396), .SI(WX3395), .SE(n4012), .CLK(n4703), .Q(
        WX3397), .QN(n3385) );
  SDFFX1 DFF_500_Q_reg ( .D(WX3398), .SI(WX3397), .SE(n4012), .CLK(n4703), .Q(
        WX3399), .QN(n7217) );
  SDFFX1 DFF_501_Q_reg ( .D(WX3400), .SI(WX3399), .SE(n4011), .CLK(n4703), .Q(
        WX3401) );
  SDFFX1 DFF_502_Q_reg ( .D(WX3402), .SI(WX3401), .SE(n4011), .CLK(n4703), .Q(
        WX3403) );
  SDFFX1 DFF_503_Q_reg ( .D(WX3404), .SI(WX3403), .SE(n4011), .CLK(n4703), .Q(
        test_so28) );
  SDFFX1 DFF_504_Q_reg ( .D(WX3406), .SI(test_si29), .SE(n4214), .CLK(n4602), 
        .Q(WX3407) );
  SDFFX1 DFF_505_Q_reg ( .D(WX3408), .SI(WX3407), .SE(n4214), .CLK(n4602), .Q(
        WX3409), .QN(n3380) );
  SDFFX1 DFF_506_Q_reg ( .D(WX3410), .SI(WX3409), .SE(n4213), .CLK(n4602), .Q(
        WX3411) );
  SDFFX1 DFF_507_Q_reg ( .D(WX3412), .SI(WX3411), .SE(n4213), .CLK(n4602), .Q(
        WX3413), .QN(n7216) );
  SDFFX1 DFF_508_Q_reg ( .D(WX3414), .SI(WX3413), .SE(n4212), .CLK(n4603), .Q(
        WX3415) );
  SDFFX1 DFF_509_Q_reg ( .D(WX3416), .SI(WX3415), .SE(n4211), .CLK(n4603), .Q(
        WX3417) );
  SDFFX1 DFF_510_Q_reg ( .D(WX3418), .SI(WX3417), .SE(n4211), .CLK(n4603), .Q(
        WX3419) );
  SDFFX1 DFF_511_Q_reg ( .D(WX3420), .SI(WX3419), .SE(n4210), .CLK(n4604), .Q(
        WX3421), .QN(n7215) );
  SDFFX1 DFF_512_Q_reg ( .D(WX3422), .SI(WX3421), .SE(n4209), .CLK(n4604), .Q(
        WX3423), .QN(n3721) );
  SDFFX1 DFF_513_Q_reg ( .D(WX3424), .SI(WX3423), .SE(n4209), .CLK(n4604), .Q(
        WX3425), .QN(n3722) );
  SDFFX1 DFF_514_Q_reg ( .D(WX3426), .SI(WX3425), .SE(n4209), .CLK(n4604), .Q(
        WX3427), .QN(n3724) );
  SDFFX1 DFF_515_Q_reg ( .D(WX3428), .SI(WX3427), .SE(n4208), .CLK(n4605), .Q(
        WX3429), .QN(n3726) );
  SDFFX1 DFF_516_Q_reg ( .D(WX3430), .SI(WX3429), .SE(n4208), .CLK(n4605), .Q(
        WX3431), .QN(n3728) );
  SDFFX1 DFF_517_Q_reg ( .D(WX3432), .SI(WX3431), .SE(n4208), .CLK(n4605), .Q(
        WX3433), .QN(n3730) );
  SDFFX1 DFF_518_Q_reg ( .D(WX3434), .SI(WX3433), .SE(n4208), .CLK(n4605), .Q(
        WX3435), .QN(n3732) );
  SDFFX1 DFF_519_Q_reg ( .D(WX3436), .SI(WX3435), .SE(n4207), .CLK(n4605), .Q(
        WX3437), .QN(n3734) );
  SDFFX1 DFF_520_Q_reg ( .D(WX3438), .SI(WX3437), .SE(n4207), .CLK(n4605), .Q(
        test_so29) );
  SDFFX1 DFF_521_Q_reg ( .D(WX3440), .SI(test_si30), .SE(n4223), .CLK(n4597), 
        .Q(WX3441), .QN(n3736) );
  SDFFX1 DFF_522_Q_reg ( .D(WX3442), .SI(WX3441), .SE(n4222), .CLK(n4598), .Q(
        WX3443), .QN(n3738) );
  SDFFX1 DFF_523_Q_reg ( .D(WX3444), .SI(WX3443), .SE(n4222), .CLK(n4598), .Q(
        WX3445), .QN(n3740) );
  SDFFX1 DFF_524_Q_reg ( .D(WX3446), .SI(WX3445), .SE(n4221), .CLK(n4598), .Q(
        WX3447), .QN(n3742) );
  SDFFX1 DFF_525_Q_reg ( .D(WX3448), .SI(WX3447), .SE(n4220), .CLK(n4599), .Q(
        WX3449), .QN(n3744) );
  SDFFX1 DFF_526_Q_reg ( .D(WX3450), .SI(WX3449), .SE(n4220), .CLK(n4599), .Q(
        WX3451), .QN(n3746) );
  SDFFX1 DFF_527_Q_reg ( .D(WX3452), .SI(WX3451), .SE(n4219), .CLK(n4599), .Q(
        WX3453), .QN(n3427) );
  SDFFX1 DFF_528_Q_reg ( .D(WX3454), .SI(WX3453), .SE(n4013), .CLK(n4702), .Q(
        WX3455), .QN(n3747) );
  SDFFX1 DFF_529_Q_reg ( .D(WX3456), .SI(WX3455), .SE(n4013), .CLK(n4702), .Q(
        WX3457), .QN(n3748) );
  SDFFX1 DFF_530_Q_reg ( .D(WX3458), .SI(WX3457), .SE(n4012), .CLK(n4703), .Q(
        WX3459), .QN(n3750) );
  SDFFX1 DFF_531_Q_reg ( .D(WX3460), .SI(WX3459), .SE(n4012), .CLK(n4703), .Q(
        WX3461), .QN(n3752) );
  SDFFX1 DFF_532_Q_reg ( .D(WX3462), .SI(WX3461), .SE(n4011), .CLK(n4703), .Q(
        WX3463), .QN(n3428) );
  SDFFX1 DFF_533_Q_reg ( .D(WX3464), .SI(WX3463), .SE(n4011), .CLK(n4703), .Q(
        WX3465), .QN(n3754) );
  SDFFX1 DFF_534_Q_reg ( .D(WX3466), .SI(WX3465), .SE(n4011), .CLK(n4703), .Q(
        WX3467), .QN(n3755) );
  SDFFX1 DFF_535_Q_reg ( .D(WX3468), .SI(WX3467), .SE(n4010), .CLK(n4704), .Q(
        WX3469), .QN(n3756) );
  SDFFX1 DFF_536_Q_reg ( .D(WX3470), .SI(WX3469), .SE(n4010), .CLK(n4704), .Q(
        WX3471), .QN(n3758) );
  SDFFX1 DFF_537_Q_reg ( .D(WX3472), .SI(WX3471), .SE(n4010), .CLK(n4704), .Q(
        test_so30) );
  SDFFX1 DFF_538_Q_reg ( .D(WX3474), .SI(test_si31), .SE(n4213), .CLK(n4602), 
        .Q(WX3475), .QN(n3760) );
  SDFFX1 DFF_539_Q_reg ( .D(WX3476), .SI(WX3475), .SE(n4212), .CLK(n4603), .Q(
        WX3477), .QN(n3429) );
  SDFFX1 DFF_540_Q_reg ( .D(WX3478), .SI(WX3477), .SE(n4212), .CLK(n4603), .Q(
        WX3479), .QN(n3762) );
  SDFFX1 DFF_541_Q_reg ( .D(WX3480), .SI(WX3479), .SE(n4211), .CLK(n4603), .Q(
        WX3481), .QN(n3764) );
  SDFFX1 DFF_542_Q_reg ( .D(WX3482), .SI(WX3481), .SE(n4210), .CLK(n4604), .Q(
        WX3483), .QN(n3766) );
  SDFFX1 DFF_543_Q_reg ( .D(WX3484), .SI(WX3483), .SE(n4210), .CLK(n4604), .Q(
        WX3485), .QN(n3439) );
  SDFFX1 DFF_544_Q_reg ( .D(WX3850), .SI(WX3485), .SE(n4016), .CLK(n4701), .Q(
        CRC_OUT_7_0), .QN(DFF_544_n1) );
  SDFFX1 DFF_545_Q_reg ( .D(WX3852), .SI(CRC_OUT_7_0), .SE(n4016), .CLK(n4701), 
        .Q(CRC_OUT_7_1), .QN(DFF_545_n1) );
  SDFFX1 DFF_546_Q_reg ( .D(WX3854), .SI(CRC_OUT_7_1), .SE(n4016), .CLK(n4701), 
        .Q(CRC_OUT_7_2), .QN(DFF_546_n1) );
  SDFFX1 DFF_547_Q_reg ( .D(WX3856), .SI(CRC_OUT_7_2), .SE(n4016), .CLK(n4701), 
        .Q(CRC_OUT_7_3) );
  SDFFX1 DFF_548_Q_reg ( .D(WX3858), .SI(CRC_OUT_7_3), .SE(n4016), .CLK(n4701), 
        .Q(CRC_OUT_7_4), .QN(DFF_548_n1) );
  SDFFX1 DFF_549_Q_reg ( .D(WX3860), .SI(CRC_OUT_7_4), .SE(n4016), .CLK(n4701), 
        .Q(CRC_OUT_7_5) );
  SDFFX1 DFF_550_Q_reg ( .D(WX3862), .SI(CRC_OUT_7_5), .SE(n4015), .CLK(n4701), 
        .Q(CRC_OUT_7_6), .QN(DFF_550_n1) );
  SDFFX1 DFF_551_Q_reg ( .D(WX3864), .SI(CRC_OUT_7_6), .SE(n4015), .CLK(n4701), 
        .Q(CRC_OUT_7_7), .QN(DFF_551_n1) );
  SDFFX1 DFF_552_Q_reg ( .D(WX3866), .SI(CRC_OUT_7_7), .SE(n4015), .CLK(n4701), 
        .Q(CRC_OUT_7_8), .QN(DFF_552_n1) );
  SDFFX1 DFF_553_Q_reg ( .D(WX3868), .SI(CRC_OUT_7_8), .SE(n4015), .CLK(n4701), 
        .Q(CRC_OUT_7_9), .QN(DFF_553_n1) );
  SDFFX1 DFF_554_Q_reg ( .D(WX3870), .SI(CRC_OUT_7_9), .SE(n4015), .CLK(n4701), 
        .Q(test_so31) );
  SDFFX1 DFF_555_Q_reg ( .D(WX3872), .SI(test_si32), .SE(n4015), .CLK(n4701), 
        .Q(CRC_OUT_7_11), .QN(DFF_555_n1) );
  SDFFX1 DFF_556_Q_reg ( .D(WX3874), .SI(CRC_OUT_7_11), .SE(n4014), .CLK(n4702), .Q(CRC_OUT_7_12), .QN(DFF_556_n1) );
  SDFFX1 DFF_557_Q_reg ( .D(WX3876), .SI(CRC_OUT_7_12), .SE(n4014), .CLK(n4702), .Q(CRC_OUT_7_13), .QN(DFF_557_n1) );
  SDFFX1 DFF_558_Q_reg ( .D(WX3878), .SI(CRC_OUT_7_13), .SE(n4014), .CLK(n4702), .Q(CRC_OUT_7_14), .QN(DFF_558_n1) );
  SDFFX1 DFF_559_Q_reg ( .D(WX3880), .SI(CRC_OUT_7_14), .SE(n4014), .CLK(n4702), .Q(CRC_OUT_7_15) );
  SDFFX1 DFF_560_Q_reg ( .D(WX3882), .SI(CRC_OUT_7_15), .SE(n4010), .CLK(n4704), .Q(CRC_OUT_7_16), .QN(DFF_560_n1) );
  SDFFX1 DFF_561_Q_reg ( .D(WX3884), .SI(CRC_OUT_7_16), .SE(n4010), .CLK(n4704), .Q(CRC_OUT_7_17), .QN(DFF_561_n1) );
  SDFFX1 DFF_562_Q_reg ( .D(WX3886), .SI(CRC_OUT_7_17), .SE(n4010), .CLK(n4704), .Q(CRC_OUT_7_18), .QN(DFF_562_n1) );
  SDFFX1 DFF_563_Q_reg ( .D(WX3888), .SI(CRC_OUT_7_18), .SE(n4009), .CLK(n4704), .Q(CRC_OUT_7_19), .QN(DFF_563_n1) );
  SDFFX1 DFF_564_Q_reg ( .D(WX3890), .SI(CRC_OUT_7_19), .SE(n4009), .CLK(n4704), .Q(CRC_OUT_7_20), .QN(DFF_564_n1) );
  SDFFX1 DFF_565_Q_reg ( .D(WX3892), .SI(CRC_OUT_7_20), .SE(n4009), .CLK(n4704), .Q(CRC_OUT_7_21), .QN(DFF_565_n1) );
  SDFFX1 DFF_566_Q_reg ( .D(WX3894), .SI(CRC_OUT_7_21), .SE(n4009), .CLK(n4704), .Q(CRC_OUT_7_22) );
  SDFFX1 DFF_567_Q_reg ( .D(WX3896), .SI(CRC_OUT_7_22), .SE(n4009), .CLK(n4704), .Q(CRC_OUT_7_23), .QN(DFF_567_n1) );
  SDFFX1 DFF_568_Q_reg ( .D(WX3898), .SI(CRC_OUT_7_23), .SE(n4009), .CLK(n4704), .Q(CRC_OUT_7_24), .QN(DFF_568_n1) );
  SDFFX1 DFF_569_Q_reg ( .D(WX3900), .SI(CRC_OUT_7_24), .SE(n4008), .CLK(n4705), .Q(CRC_OUT_7_25), .QN(DFF_569_n1) );
  SDFFX1 DFF_570_Q_reg ( .D(WX3902), .SI(CRC_OUT_7_25), .SE(n4207), .CLK(n4605), .Q(CRC_OUT_7_26), .QN(DFF_570_n1) );
  SDFFX1 DFF_571_Q_reg ( .D(WX3904), .SI(CRC_OUT_7_26), .SE(n4207), .CLK(n4605), .Q(test_so32) );
  SDFFX1 DFF_572_Q_reg ( .D(WX3906), .SI(test_si33), .SE(n4207), .CLK(n4605), 
        .Q(CRC_OUT_7_28), .QN(DFF_572_n1) );
  SDFFX1 DFF_573_Q_reg ( .D(WX3908), .SI(CRC_OUT_7_28), .SE(n4207), .CLK(n4605), .Q(CRC_OUT_7_29), .QN(DFF_573_n1) );
  SDFFX1 DFF_574_Q_reg ( .D(WX3910), .SI(CRC_OUT_7_29), .SE(n4206), .CLK(n4606), .Q(CRC_OUT_7_30), .QN(DFF_574_n1) );
  SDFFX1 DFF_575_Q_reg ( .D(WX3912), .SI(CRC_OUT_7_30), .SE(n4206), .CLK(n4606), .Q(CRC_OUT_7_31), .QN(DFF_575_n1) );
  SDFFX1 DFF_576_Q_reg ( .D(n190), .SI(CRC_OUT_7_31), .SE(n4206), .CLK(n4606), 
        .Q(WX4364) );
  SDFFX1 DFF_577_Q_reg ( .D(n191), .SI(WX4364), .SE(n4201), .CLK(n4608), .Q(
        n8586) );
  SDFFX1 DFF_578_Q_reg ( .D(n192), .SI(n8586), .SE(n4201), .CLK(n4608), .Q(
        n8585) );
  SDFFX1 DFF_579_Q_reg ( .D(n193), .SI(n8585), .SE(n4201), .CLK(n4608), .Q(
        n8584) );
  SDFFX1 DFF_580_Q_reg ( .D(n194), .SI(n8584), .SE(n4201), .CLK(n4608), .Q(
        n8583) );
  SDFFX1 DFF_581_Q_reg ( .D(n195), .SI(n8583), .SE(n4202), .CLK(n4608), .Q(
        n8582) );
  SDFFX1 DFF_582_Q_reg ( .D(n196), .SI(n8582), .SE(n4202), .CLK(n4608), .Q(
        n8581) );
  SDFFX1 DFF_583_Q_reg ( .D(n197), .SI(n8581), .SE(n4202), .CLK(n4608), .Q(
        n8580) );
  SDFFX1 DFF_584_Q_reg ( .D(n198), .SI(n8580), .SE(n4202), .CLK(n4608), .Q(
        n8579) );
  SDFFX1 DFF_585_Q_reg ( .D(n199), .SI(n8579), .SE(n4202), .CLK(n4608), .Q(
        n8578) );
  SDFFX1 DFF_586_Q_reg ( .D(n200), .SI(n8578), .SE(n4202), .CLK(n4608), .Q(
        n8577) );
  SDFFX1 DFF_587_Q_reg ( .D(n201), .SI(n8577), .SE(n4203), .CLK(n4607), .Q(
        n8576) );
  SDFFX1 DFF_588_Q_reg ( .D(n202), .SI(n8576), .SE(n4203), .CLK(n4607), .Q(
        test_so33) );
  SDFFX1 DFF_589_Q_reg ( .D(n203), .SI(test_si34), .SE(n4203), .CLK(n4607), 
        .Q(n8573) );
  SDFFX1 DFF_590_Q_reg ( .D(n204), .SI(n8573), .SE(n4203), .CLK(n4607), .Q(
        n8572) );
  SDFFX1 DFF_591_Q_reg ( .D(n205), .SI(n8572), .SE(n4203), .CLK(n4607), .Q(
        n8571) );
  SDFFX1 DFF_592_Q_reg ( .D(n206), .SI(n8571), .SE(n4203), .CLK(n4607), .Q(
        n8570) );
  SDFFX1 DFF_593_Q_reg ( .D(n207), .SI(n8570), .SE(n4204), .CLK(n4607), .Q(
        n8569) );
  SDFFX1 DFF_594_Q_reg ( .D(n208), .SI(n8569), .SE(n4204), .CLK(n4607), .Q(
        n8568) );
  SDFFX1 DFF_595_Q_reg ( .D(n209), .SI(n8568), .SE(n4204), .CLK(n4607), .Q(
        n8567) );
  SDFFX1 DFF_596_Q_reg ( .D(n210), .SI(n8567), .SE(n4204), .CLK(n4607), .Q(
        n8566) );
  SDFFX1 DFF_597_Q_reg ( .D(n211), .SI(n8566), .SE(n4204), .CLK(n4607), .Q(
        n8565) );
  SDFFX1 DFF_598_Q_reg ( .D(n212), .SI(n8565), .SE(n4204), .CLK(n4607), .Q(
        n8564) );
  SDFFX1 DFF_599_Q_reg ( .D(n213), .SI(n8564), .SE(n4205), .CLK(n4606), .Q(
        n8563) );
  SDFFX1 DFF_600_Q_reg ( .D(n214), .SI(n8563), .SE(n4205), .CLK(n4606), .Q(
        n8562) );
  SDFFX1 DFF_601_Q_reg ( .D(n215), .SI(n8562), .SE(n4205), .CLK(n4606), .Q(
        n8561) );
  SDFFX1 DFF_602_Q_reg ( .D(n216), .SI(n8561), .SE(n4205), .CLK(n4606), .Q(
        n8560) );
  SDFFX1 DFF_603_Q_reg ( .D(n217), .SI(n8560), .SE(n4205), .CLK(n4606), .Q(
        n8559) );
  SDFFX1 DFF_604_Q_reg ( .D(n218), .SI(n8559), .SE(n4205), .CLK(n4606), .Q(
        n8558) );
  SDFFX1 DFF_605_Q_reg ( .D(n219), .SI(n8558), .SE(n4206), .CLK(n4606), .Q(
        test_so34) );
  SDFFX1 DFF_606_Q_reg ( .D(n220), .SI(test_si35), .SE(n4206), .CLK(n4606), 
        .Q(n8555) );
  SDFFX1 DFF_607_Q_reg ( .D(WX4425), .SI(n8555), .SE(n4206), .CLK(n4606), .Q(
        n8554) );
  SDFFX1 DFF_608_Q_reg ( .D(WX4523), .SI(n8554), .SE(n4201), .CLK(n4608), .Q(
        n8553), .QN(n7214) );
  SDFFX1 DFF_609_Q_reg ( .D(WX4525), .SI(n8553), .SE(n4200), .CLK(n4609), .Q(
        n8552), .QN(n7213) );
  SDFFX1 DFF_610_Q_reg ( .D(WX4527), .SI(n8552), .SE(n4200), .CLK(n4609), .Q(
        n8551), .QN(n7212) );
  SDFFX1 DFF_611_Q_reg ( .D(WX4529), .SI(n8551), .SE(n4199), .CLK(n4609), .Q(
        n8550), .QN(n7211) );
  SDFFX1 DFF_612_Q_reg ( .D(WX4531), .SI(n8550), .SE(n4199), .CLK(n4609), .Q(
        n8549), .QN(n7210) );
  SDFFX1 DFF_613_Q_reg ( .D(WX4533), .SI(n8549), .SE(n4198), .CLK(n4610), .Q(
        n8548), .QN(n7209) );
  SDFFX1 DFF_614_Q_reg ( .D(WX4535), .SI(n8548), .SE(n4198), .CLK(n4610), .Q(
        n8547), .QN(n7208) );
  SDFFX1 DFF_615_Q_reg ( .D(WX4537), .SI(n8547), .SE(n4197), .CLK(n4610), .Q(
        n8546), .QN(n7207) );
  SDFFX1 DFF_616_Q_reg ( .D(WX4539), .SI(n8546), .SE(n4196), .CLK(n4611), .Q(
        n8545), .QN(n7206) );
  SDFFX1 DFF_617_Q_reg ( .D(WX4541), .SI(n8545), .SE(n4195), .CLK(n4611), .Q(
        n8544), .QN(n7205) );
  SDFFX1 DFF_618_Q_reg ( .D(WX4543), .SI(n8544), .SE(n4195), .CLK(n4611), .Q(
        n8543), .QN(n7204) );
  SDFFX1 DFF_619_Q_reg ( .D(WX4545), .SI(n8543), .SE(n4194), .CLK(n4612), .Q(
        n8542), .QN(n7203) );
  SDFFX1 DFF_620_Q_reg ( .D(WX4547), .SI(n8542), .SE(n4194), .CLK(n4612), .Q(
        n8541), .QN(n7202) );
  SDFFX1 DFF_621_Q_reg ( .D(WX4549), .SI(n8541), .SE(n4017), .CLK(n4700), .Q(
        n8540), .QN(n7201) );
  SDFFX1 DFF_622_Q_reg ( .D(WX4551), .SI(n8540), .SE(n4218), .CLK(n4600), .Q(
        test_so35) );
  SDFFX1 DFF_623_Q_reg ( .D(WX4553), .SI(test_si36), .SE(n4217), .CLK(n4600), 
        .Q(n8537), .QN(n7199) );
  SDFFX1 DFF_624_Q_reg ( .D(WX4555), .SI(n8537), .SE(n4217), .CLK(n4600), .Q(
        WX4556) );
  SDFFX1 DFF_625_Q_reg ( .D(WX4557), .SI(WX4556), .SE(n4217), .CLK(n4600), .Q(
        WX4558), .QN(n3372) );
  SDFFX1 DFF_626_Q_reg ( .D(WX4559), .SI(WX4558), .SE(n4191), .CLK(n4613), .Q(
        WX4560) );
  SDFFX1 DFF_627_Q_reg ( .D(WX4561), .SI(WX4560), .SE(n4191), .CLK(n4613), .Q(
        WX4562), .QN(n3371) );
  SDFFX1 DFF_628_Q_reg ( .D(WX4563), .SI(WX4562), .SE(n4190), .CLK(n4614), .Q(
        WX4564) );
  SDFFX1 DFF_629_Q_reg ( .D(WX4565), .SI(WX4564), .SE(n4189), .CLK(n4614), .Q(
        WX4566), .QN(n3369) );
  SDFFX1 DFF_630_Q_reg ( .D(WX4567), .SI(WX4566), .SE(n4189), .CLK(n4614), .Q(
        WX4568), .QN(n3368) );
  SDFFX1 DFF_631_Q_reg ( .D(WX4569), .SI(WX4568), .SE(n4188), .CLK(n4615), .Q(
        WX4570), .QN(n3367) );
  SDFFX1 DFF_632_Q_reg ( .D(WX4571), .SI(WX4570), .SE(n4187), .CLK(n4615), .Q(
        WX4572), .QN(n3366) );
  SDFFX1 DFF_633_Q_reg ( .D(WX4573), .SI(WX4572), .SE(n4187), .CLK(n4615), .Q(
        WX4574), .QN(n3365) );
  SDFFX1 DFF_634_Q_reg ( .D(WX4575), .SI(WX4574), .SE(n4186), .CLK(n4616), .Q(
        WX4576), .QN(n3364) );
  SDFFX1 DFF_635_Q_reg ( .D(WX4577), .SI(WX4576), .SE(n4185), .CLK(n4616), .Q(
        WX4578), .QN(n3363) );
  SDFFX1 DFF_636_Q_reg ( .D(WX4579), .SI(WX4578), .SE(n4185), .CLK(n4616), .Q(
        WX4580), .QN(n3362) );
  SDFFX1 DFF_637_Q_reg ( .D(WX4581), .SI(WX4580), .SE(n4184), .CLK(n4617), .Q(
        WX4582), .QN(n3361) );
  SDFFX1 DFF_638_Q_reg ( .D(WX4583), .SI(WX4582), .SE(n4183), .CLK(n4617), .Q(
        WX4584), .QN(n3360) );
  SDFFX1 DFF_639_Q_reg ( .D(WX4585), .SI(WX4584), .SE(n4183), .CLK(n4617), .Q(
        test_so36) );
  SDFFX1 DFF_640_Q_reg ( .D(n221), .SI(test_si37), .SE(n4201), .CLK(n4608), 
        .Q(WX4588), .QN(n3070) );
  SDFFX1 DFF_641_Q_reg ( .D(n222), .SI(WX4588), .SE(n4200), .CLK(n4609), .Q(
        WX4590), .QN(n3234) );
  SDFFX1 DFF_642_Q_reg ( .D(n223), .SI(WX4590), .SE(n4200), .CLK(n4609), .Q(
        WX4592), .QN(n3232) );
  SDFFX1 DFF_643_Q_reg ( .D(n224), .SI(WX4592), .SE(n4200), .CLK(n4609), .Q(
        WX4594), .QN(n3231) );
  SDFFX1 DFF_644_Q_reg ( .D(n225), .SI(WX4594), .SE(n4199), .CLK(n4609), .Q(
        WX4596), .QN(n3229) );
  SDFFX1 DFF_645_Q_reg ( .D(n226), .SI(WX4596), .SE(n4198), .CLK(n4610), .Q(
        WX4598), .QN(n3227) );
  SDFFX1 DFF_646_Q_reg ( .D(n227), .SI(WX4598), .SE(n4198), .CLK(n4610), .Q(
        WX4600), .QN(n3225) );
  SDFFX1 DFF_647_Q_reg ( .D(n228), .SI(WX4600), .SE(n4197), .CLK(n4610), .Q(
        WX4602), .QN(n3223) );
  SDFFX1 DFF_648_Q_reg ( .D(n229), .SI(WX4602), .SE(n4196), .CLK(n4611), .Q(
        WX4604), .QN(n3221) );
  SDFFX1 DFF_649_Q_reg ( .D(n230), .SI(WX4604), .SE(n4196), .CLK(n4611), .Q(
        WX4606), .QN(n3219) );
  SDFFX1 DFF_650_Q_reg ( .D(n231), .SI(WX4606), .SE(n4195), .CLK(n4611), .Q(
        WX4608), .QN(n3217) );
  SDFFX1 DFF_651_Q_reg ( .D(n232), .SI(WX4608), .SE(n4194), .CLK(n4612), .Q(
        WX4610), .QN(n3215) );
  SDFFX1 DFF_652_Q_reg ( .D(n233), .SI(WX4610), .SE(n4194), .CLK(n4612), .Q(
        WX4612), .QN(n3213) );
  SDFFX1 DFF_653_Q_reg ( .D(n234), .SI(WX4612), .SE(n4193), .CLK(n4612), .Q(
        WX4614), .QN(n3211) );
  SDFFX1 DFF_654_Q_reg ( .D(n235), .SI(WX4614), .SE(n4218), .CLK(n4600), .Q(
        WX4616), .QN(n3210) );
  SDFFX1 DFF_655_Q_reg ( .D(n236), .SI(WX4616), .SE(n4217), .CLK(n4600), .Q(
        WX4618), .QN(n3208) );
  SDFFX1 DFF_656_Q_reg ( .D(WX4619), .SI(WX4618), .SE(n4217), .CLK(n4600), .Q(
        test_so37) );
  SDFFX1 DFF_657_Q_reg ( .D(WX4621), .SI(test_si38), .SE(n4217), .CLK(n4600), 
        .Q(WX4622) );
  SDFFX1 DFF_658_Q_reg ( .D(WX4623), .SI(WX4622), .SE(n4191), .CLK(n4613), .Q(
        WX4624), .QN(n3717) );
  SDFFX1 DFF_659_Q_reg ( .D(WX4625), .SI(WX4624), .SE(n4190), .CLK(n4614), .Q(
        WX4626) );
  SDFFX1 DFF_660_Q_reg ( .D(WX4627), .SI(WX4626), .SE(n4190), .CLK(n4614), .Q(
        WX4628), .QN(n3713) );
  SDFFX1 DFF_661_Q_reg ( .D(WX4629), .SI(WX4628), .SE(n4189), .CLK(n4614), .Q(
        WX4630) );
  SDFFX1 DFF_662_Q_reg ( .D(WX4631), .SI(WX4630), .SE(n4188), .CLK(n4615), .Q(
        WX4632) );
  SDFFX1 DFF_663_Q_reg ( .D(WX4633), .SI(WX4632), .SE(n4188), .CLK(n4615), .Q(
        WX4634), .QN(n3707) );
  SDFFX1 DFF_664_Q_reg ( .D(WX4635), .SI(WX4634), .SE(n4187), .CLK(n4615), .Q(
        WX4636), .QN(n3705) );
  SDFFX1 DFF_665_Q_reg ( .D(WX4637), .SI(WX4636), .SE(n4186), .CLK(n4616), .Q(
        WX4638), .QN(n3703) );
  SDFFX1 DFF_666_Q_reg ( .D(WX4639), .SI(WX4638), .SE(n4186), .CLK(n4616), .Q(
        WX4640), .QN(n3701) );
  SDFFX1 DFF_667_Q_reg ( .D(WX4641), .SI(WX4640), .SE(n4185), .CLK(n4616), .Q(
        WX4642) );
  SDFFX1 DFF_668_Q_reg ( .D(WX4643), .SI(WX4642), .SE(n4184), .CLK(n4617), .Q(
        WX4644), .QN(n3697) );
  SDFFX1 DFF_669_Q_reg ( .D(WX4645), .SI(WX4644), .SE(n4184), .CLK(n4617), .Q(
        WX4646), .QN(n3695) );
  SDFFX1 DFF_670_Q_reg ( .D(WX4647), .SI(WX4646), .SE(n4183), .CLK(n4617), .Q(
        WX4648), .QN(n3693) );
  SDFFX1 DFF_671_Q_reg ( .D(WX4649), .SI(WX4648), .SE(n4182), .CLK(n4618), .Q(
        WX4650), .QN(n3691) );
  SDFFX1 DFF_672_Q_reg ( .D(WX4651), .SI(WX4650), .SE(n4182), .CLK(n4618), .Q(
        WX4652) );
  SDFFX1 DFF_673_Q_reg ( .D(WX4653), .SI(WX4652), .SE(n4182), .CLK(n4618), .Q(
        test_so38) );
  SDFFX1 DFF_674_Q_reg ( .D(WX4655), .SI(test_si39), .SE(n4200), .CLK(n4609), 
        .Q(WX4656) );
  SDFFX1 DFF_675_Q_reg ( .D(WX4657), .SI(WX4656), .SE(n4199), .CLK(n4609), .Q(
        WX4658) );
  SDFFX1 DFF_676_Q_reg ( .D(WX4659), .SI(WX4658), .SE(n4199), .CLK(n4609), .Q(
        WX4660) );
  SDFFX1 DFF_677_Q_reg ( .D(WX4661), .SI(WX4660), .SE(n4198), .CLK(n4610), .Q(
        WX4662) );
  SDFFX1 DFF_678_Q_reg ( .D(WX4663), .SI(WX4662), .SE(n4197), .CLK(n4610), .Q(
        WX4664) );
  SDFFX1 DFF_679_Q_reg ( .D(WX4665), .SI(WX4664), .SE(n4197), .CLK(n4610), .Q(
        WX4666) );
  SDFFX1 DFF_680_Q_reg ( .D(WX4667), .SI(WX4666), .SE(n4196), .CLK(n4611), .Q(
        WX4668) );
  SDFFX1 DFF_681_Q_reg ( .D(WX4669), .SI(WX4668), .SE(n4196), .CLK(n4611), .Q(
        WX4670) );
  SDFFX1 DFF_682_Q_reg ( .D(WX4671), .SI(WX4670), .SE(n4195), .CLK(n4611), .Q(
        WX4672) );
  SDFFX1 DFF_683_Q_reg ( .D(WX4673), .SI(WX4672), .SE(n4194), .CLK(n4612), .Q(
        WX4674) );
  SDFFX1 DFF_684_Q_reg ( .D(WX4675), .SI(WX4674), .SE(n4193), .CLK(n4612), .Q(
        WX4676) );
  SDFFX1 DFF_685_Q_reg ( .D(WX4677), .SI(WX4676), .SE(n4193), .CLK(n4612), .Q(
        WX4678) );
  SDFFX1 DFF_686_Q_reg ( .D(WX4679), .SI(WX4678), .SE(n4193), .CLK(n4612), .Q(
        WX4680), .QN(n7200) );
  SDFFX1 DFF_687_Q_reg ( .D(WX4681), .SI(WX4680), .SE(n4192), .CLK(n4613), .Q(
        WX4682) );
  SDFFX1 DFF_688_Q_reg ( .D(WX4683), .SI(WX4682), .SE(n4192), .CLK(n4613), .Q(
        WX4684), .QN(n3373) );
  SDFFX1 DFF_689_Q_reg ( .D(WX4685), .SI(WX4684), .SE(n4192), .CLK(n4613), .Q(
        WX4686), .QN(n7198) );
  SDFFX1 DFF_690_Q_reg ( .D(WX4687), .SI(WX4686), .SE(n4191), .CLK(n4613), .Q(
        test_so39) );
  SDFFX1 DFF_691_Q_reg ( .D(WX4689), .SI(test_si40), .SE(n4190), .CLK(n4614), 
        .Q(WX4690), .QN(n7197) );
  SDFFX1 DFF_692_Q_reg ( .D(WX4691), .SI(WX4690), .SE(n4190), .CLK(n4614), .Q(
        WX4692), .QN(n3370) );
  SDFFX1 DFF_693_Q_reg ( .D(WX4693), .SI(WX4692), .SE(n4189), .CLK(n4614), .Q(
        WX4694), .QN(n7196) );
  SDFFX1 DFF_694_Q_reg ( .D(WX4695), .SI(WX4694), .SE(n4188), .CLK(n4615), .Q(
        WX4696), .QN(n7195) );
  SDFFX1 DFF_695_Q_reg ( .D(WX4697), .SI(WX4696), .SE(n4188), .CLK(n4615), .Q(
        WX4698) );
  SDFFX1 DFF_696_Q_reg ( .D(WX4699), .SI(WX4698), .SE(n4187), .CLK(n4615), .Q(
        WX4700) );
  SDFFX1 DFF_697_Q_reg ( .D(WX4701), .SI(WX4700), .SE(n4186), .CLK(n4616), .Q(
        WX4702) );
  SDFFX1 DFF_698_Q_reg ( .D(WX4703), .SI(WX4702), .SE(n4186), .CLK(n4616), .Q(
        WX4704) );
  SDFFX1 DFF_699_Q_reg ( .D(WX4705), .SI(WX4704), .SE(n4185), .CLK(n4616), .Q(
        WX4706), .QN(n7194) );
  SDFFX1 DFF_700_Q_reg ( .D(WX4707), .SI(WX4706), .SE(n4184), .CLK(n4617), .Q(
        WX4708) );
  SDFFX1 DFF_701_Q_reg ( .D(WX4709), .SI(WX4708), .SE(n4184), .CLK(n4617), .Q(
        WX4710) );
  SDFFX1 DFF_702_Q_reg ( .D(WX4711), .SI(WX4710), .SE(n4183), .CLK(n4617), .Q(
        WX4712) );
  SDFFX1 DFF_703_Q_reg ( .D(WX4713), .SI(WX4712), .SE(n4182), .CLK(n4618), .Q(
        WX4714) );
  SDFFX1 DFF_704_Q_reg ( .D(WX4715), .SI(WX4714), .SE(n4182), .CLK(n4618), .Q(
        WX4716), .QN(n3668) );
  SDFFX1 DFF_705_Q_reg ( .D(WX4717), .SI(WX4716), .SE(n4181), .CLK(n4618), .Q(
        WX4718), .QN(n3670) );
  SDFFX1 DFF_706_Q_reg ( .D(WX4719), .SI(WX4718), .SE(n4181), .CLK(n4618), .Q(
        WX4720), .QN(n3672) );
  SDFFX1 DFF_707_Q_reg ( .D(WX4721), .SI(WX4720), .SE(n4181), .CLK(n4618), .Q(
        test_so40) );
  SDFFX1 DFF_708_Q_reg ( .D(WX4723), .SI(test_si41), .SE(n4199), .CLK(n4609), 
        .Q(WX4724), .QN(n3674) );
  SDFFX1 DFF_709_Q_reg ( .D(WX4725), .SI(WX4724), .SE(n4198), .CLK(n4610), .Q(
        WX4726), .QN(n3676) );
  SDFFX1 DFF_710_Q_reg ( .D(WX4727), .SI(WX4726), .SE(n4197), .CLK(n4610), .Q(
        WX4728), .QN(n3678) );
  SDFFX1 DFF_711_Q_reg ( .D(WX4729), .SI(WX4728), .SE(n4197), .CLK(n4610), .Q(
        WX4730), .QN(n3680) );
  SDFFX1 DFF_712_Q_reg ( .D(WX4731), .SI(WX4730), .SE(n4196), .CLK(n4611), .Q(
        WX4732), .QN(n3682) );
  SDFFX1 DFF_713_Q_reg ( .D(WX4733), .SI(WX4732), .SE(n4195), .CLK(n4611), .Q(
        WX4734), .QN(n3684) );
  SDFFX1 DFF_714_Q_reg ( .D(WX4735), .SI(WX4734), .SE(n4195), .CLK(n4611), .Q(
        WX4736), .QN(n3686) );
  SDFFX1 DFF_715_Q_reg ( .D(WX4737), .SI(WX4736), .SE(n4194), .CLK(n4612), .Q(
        WX4738), .QN(n3688) );
  SDFFX1 DFF_716_Q_reg ( .D(WX4739), .SI(WX4738), .SE(n4193), .CLK(n4612), .Q(
        WX4740), .QN(n3690) );
  SDFFX1 DFF_717_Q_reg ( .D(WX4741), .SI(WX4740), .SE(n4193), .CLK(n4612), .Q(
        WX4742), .QN(n3692) );
  SDFFX1 DFF_718_Q_reg ( .D(WX4743), .SI(WX4742), .SE(n4192), .CLK(n4613), .Q(
        WX4744), .QN(n3694) );
  SDFFX1 DFF_719_Q_reg ( .D(WX4745), .SI(WX4744), .SE(n4192), .CLK(n4613), .Q(
        WX4746), .QN(n3425) );
  SDFFX1 DFF_720_Q_reg ( .D(WX4747), .SI(WX4746), .SE(n4192), .CLK(n4613), .Q(
        WX4748), .QN(n3696) );
  SDFFX1 DFF_721_Q_reg ( .D(WX4749), .SI(WX4748), .SE(n4191), .CLK(n4613), .Q(
        WX4750), .QN(n3698) );
  SDFFX1 DFF_722_Q_reg ( .D(WX4751), .SI(WX4750), .SE(n4191), .CLK(n4613), .Q(
        WX4752), .QN(n3700) );
  SDFFX1 DFF_723_Q_reg ( .D(WX4753), .SI(WX4752), .SE(n4190), .CLK(n4614), .Q(
        WX4754), .QN(n3702) );
  SDFFX1 DFF_724_Q_reg ( .D(WX4755), .SI(WX4754), .SE(n4189), .CLK(n4614), .Q(
        test_so41) );
  SDFFX1 DFF_725_Q_reg ( .D(WX4757), .SI(test_si42), .SE(n4189), .CLK(n4614), 
        .Q(WX4758), .QN(n3704) );
  SDFFX1 DFF_726_Q_reg ( .D(WX4759), .SI(WX4758), .SE(n4188), .CLK(n4615), .Q(
        WX4760), .QN(n3706) );
  SDFFX1 DFF_727_Q_reg ( .D(WX4761), .SI(WX4760), .SE(n4187), .CLK(n4615), .Q(
        WX4762), .QN(n3708) );
  SDFFX1 DFF_728_Q_reg ( .D(WX4763), .SI(WX4762), .SE(n4187), .CLK(n4615), .Q(
        WX4764), .QN(n3710) );
  SDFFX1 DFF_729_Q_reg ( .D(WX4765), .SI(WX4764), .SE(n4186), .CLK(n4616), .Q(
        WX4766), .QN(n3712) );
  SDFFX1 DFF_730_Q_reg ( .D(WX4767), .SI(WX4766), .SE(n4185), .CLK(n4616), .Q(
        WX4768), .QN(n3714) );
  SDFFX1 DFF_731_Q_reg ( .D(WX4769), .SI(WX4768), .SE(n4185), .CLK(n4616), .Q(
        WX4770), .QN(n3426) );
  SDFFX1 DFF_732_Q_reg ( .D(WX4771), .SI(WX4770), .SE(n4184), .CLK(n4617), .Q(
        WX4772), .QN(n3716) );
  SDFFX1 DFF_733_Q_reg ( .D(WX4773), .SI(WX4772), .SE(n4183), .CLK(n4617), .Q(
        WX4774), .QN(n3718) );
  SDFFX1 DFF_734_Q_reg ( .D(WX4775), .SI(WX4774), .SE(n4183), .CLK(n4617), .Q(
        WX4776), .QN(n3720) );
  SDFFX1 DFF_735_Q_reg ( .D(WX4777), .SI(WX4776), .SE(n4182), .CLK(n4618), .Q(
        WX4778), .QN(n3438) );
  SDFFX1 DFF_736_Q_reg ( .D(WX5143), .SI(WX4778), .SE(n4022), .CLK(n4698), .Q(
        CRC_OUT_6_0), .QN(DFF_736_n1) );
  SDFFX1 DFF_737_Q_reg ( .D(WX5145), .SI(CRC_OUT_6_0), .SE(n4021), .CLK(n4698), 
        .Q(CRC_OUT_6_1), .QN(DFF_737_n1) );
  SDFFX1 DFF_738_Q_reg ( .D(WX5147), .SI(CRC_OUT_6_1), .SE(n4021), .CLK(n4698), 
        .Q(CRC_OUT_6_2), .QN(DFF_738_n1) );
  SDFFX1 DFF_739_Q_reg ( .D(WX5149), .SI(CRC_OUT_6_2), .SE(n4021), .CLK(n4698), 
        .Q(CRC_OUT_6_3) );
  SDFFX1 DFF_740_Q_reg ( .D(WX5151), .SI(CRC_OUT_6_3), .SE(n4021), .CLK(n4698), 
        .Q(CRC_OUT_6_4), .QN(DFF_740_n1) );
  SDFFX1 DFF_741_Q_reg ( .D(WX5153), .SI(CRC_OUT_6_4), .SE(n4021), .CLK(n4698), 
        .Q(test_so42) );
  SDFFX1 DFF_742_Q_reg ( .D(WX5155), .SI(test_si43), .SE(n4021), .CLK(n4698), 
        .Q(CRC_OUT_6_6), .QN(DFF_742_n1) );
  SDFFX1 DFF_743_Q_reg ( .D(WX5157), .SI(CRC_OUT_6_6), .SE(n4020), .CLK(n4699), 
        .Q(CRC_OUT_6_7), .QN(DFF_743_n1) );
  SDFFX1 DFF_744_Q_reg ( .D(WX5159), .SI(CRC_OUT_6_7), .SE(n4020), .CLK(n4699), 
        .Q(CRC_OUT_6_8), .QN(DFF_744_n1) );
  SDFFX1 DFF_745_Q_reg ( .D(WX5161), .SI(CRC_OUT_6_8), .SE(n4020), .CLK(n4699), 
        .Q(CRC_OUT_6_9), .QN(DFF_745_n1) );
  SDFFX1 DFF_746_Q_reg ( .D(WX5163), .SI(CRC_OUT_6_9), .SE(n4020), .CLK(n4699), 
        .Q(CRC_OUT_6_10), .QN(DFF_746_n1) );
  SDFFX1 DFF_747_Q_reg ( .D(WX5165), .SI(CRC_OUT_6_10), .SE(n4020), .CLK(n4699), .Q(CRC_OUT_6_11), .QN(DFF_747_n1) );
  SDFFX1 DFF_748_Q_reg ( .D(WX5167), .SI(CRC_OUT_6_11), .SE(n4020), .CLK(n4699), .Q(CRC_OUT_6_12), .QN(DFF_748_n1) );
  SDFFX1 DFF_749_Q_reg ( .D(WX5169), .SI(CRC_OUT_6_12), .SE(n4019), .CLK(n4699), .Q(CRC_OUT_6_13), .QN(DFF_749_n1) );
  SDFFX1 DFF_750_Q_reg ( .D(WX5171), .SI(CRC_OUT_6_13), .SE(n4019), .CLK(n4699), .Q(CRC_OUT_6_14), .QN(DFF_750_n1) );
  SDFFX1 DFF_751_Q_reg ( .D(WX5173), .SI(CRC_OUT_6_14), .SE(n4019), .CLK(n4699), .Q(CRC_OUT_6_15) );
  SDFFX1 DFF_752_Q_reg ( .D(WX5175), .SI(CRC_OUT_6_15), .SE(n4019), .CLK(n4699), .Q(CRC_OUT_6_16), .QN(DFF_752_n1) );
  SDFFX1 DFF_753_Q_reg ( .D(WX5177), .SI(CRC_OUT_6_16), .SE(n4019), .CLK(n4699), .Q(CRC_OUT_6_17), .QN(DFF_753_n1) );
  SDFFX1 DFF_754_Q_reg ( .D(WX5179), .SI(CRC_OUT_6_17), .SE(n4019), .CLK(n4699), .Q(CRC_OUT_6_18), .QN(DFF_754_n1) );
  SDFFX1 DFF_755_Q_reg ( .D(WX5181), .SI(CRC_OUT_6_18), .SE(n4018), .CLK(n4700), .Q(CRC_OUT_6_19), .QN(DFF_755_n1) );
  SDFFX1 DFF_756_Q_reg ( .D(WX5183), .SI(CRC_OUT_6_19), .SE(n4018), .CLK(n4700), .Q(CRC_OUT_6_20), .QN(DFF_756_n1) );
  SDFFX1 DFF_757_Q_reg ( .D(WX5185), .SI(CRC_OUT_6_20), .SE(n4018), .CLK(n4700), .Q(CRC_OUT_6_21), .QN(DFF_757_n1) );
  SDFFX1 DFF_758_Q_reg ( .D(WX5187), .SI(CRC_OUT_6_21), .SE(n4018), .CLK(n4700), .Q(test_so43) );
  SDFFX1 DFF_759_Q_reg ( .D(WX5189), .SI(test_si44), .SE(n4018), .CLK(n4700), 
        .Q(CRC_OUT_6_23), .QN(DFF_759_n1) );
  SDFFX1 DFF_760_Q_reg ( .D(WX5191), .SI(CRC_OUT_6_23), .SE(n4018), .CLK(n4700), .Q(CRC_OUT_6_24), .QN(DFF_760_n1) );
  SDFFX1 DFF_761_Q_reg ( .D(WX5193), .SI(CRC_OUT_6_24), .SE(n4017), .CLK(n4700), .Q(CRC_OUT_6_25), .QN(DFF_761_n1) );
  SDFFX1 DFF_762_Q_reg ( .D(WX5195), .SI(CRC_OUT_6_25), .SE(n4017), .CLK(n4700), .Q(CRC_OUT_6_26), .QN(DFF_762_n1) );
  SDFFX1 DFF_763_Q_reg ( .D(WX5197), .SI(CRC_OUT_6_26), .SE(n4017), .CLK(n4700), .Q(CRC_OUT_6_27) );
  SDFFX1 DFF_764_Q_reg ( .D(WX5199), .SI(CRC_OUT_6_27), .SE(n4017), .CLK(n4700), .Q(CRC_OUT_6_28), .QN(DFF_764_n1) );
  SDFFX1 DFF_765_Q_reg ( .D(WX5201), .SI(CRC_OUT_6_28), .SE(n4017), .CLK(n4700), .Q(CRC_OUT_6_29), .QN(DFF_765_n1) );
  SDFFX1 DFF_766_Q_reg ( .D(WX5203), .SI(CRC_OUT_6_29), .SE(n4181), .CLK(n4618), .Q(CRC_OUT_6_30), .QN(DFF_766_n1) );
  SDFFX1 DFF_767_Q_reg ( .D(WX5205), .SI(CRC_OUT_6_30), .SE(n4181), .CLK(n4618), .Q(CRC_OUT_6_31), .QN(DFF_767_n1) );
  SDFFX1 DFF_768_Q_reg ( .D(n268), .SI(CRC_OUT_6_31), .SE(n4181), .CLK(n4618), 
        .Q(WX5657) );
  SDFFX1 DFF_769_Q_reg ( .D(n269), .SI(WX5657), .SE(n4175), .CLK(n4621), .Q(
        n8528) );
  SDFFX1 DFF_770_Q_reg ( .D(n270), .SI(n8528), .SE(n4176), .CLK(n4621), .Q(
        n8527) );
  SDFFX1 DFF_771_Q_reg ( .D(n271), .SI(n8527), .SE(n4176), .CLK(n4621), .Q(
        n8526) );
  SDFFX1 DFF_772_Q_reg ( .D(n272), .SI(n8526), .SE(n4176), .CLK(n4621), .Q(
        n8525) );
  SDFFX1 DFF_773_Q_reg ( .D(n273), .SI(n8525), .SE(n4176), .CLK(n4621), .Q(
        n8524) );
  SDFFX1 DFF_774_Q_reg ( .D(n274), .SI(n8524), .SE(n4176), .CLK(n4621), .Q(
        n8523) );
  SDFFX1 DFF_775_Q_reg ( .D(n275), .SI(n8523), .SE(n4176), .CLK(n4621), .Q(
        test_so44) );
  SDFFX1 DFF_776_Q_reg ( .D(n276), .SI(test_si45), .SE(n4177), .CLK(n4620), 
        .Q(n8520) );
  SDFFX1 DFF_777_Q_reg ( .D(n277), .SI(n8520), .SE(n4177), .CLK(n4620), .Q(
        n8519) );
  SDFFX1 DFF_778_Q_reg ( .D(n278), .SI(n8519), .SE(n4177), .CLK(n4620), .Q(
        n8518) );
  SDFFX1 DFF_779_Q_reg ( .D(n279), .SI(n8518), .SE(n4177), .CLK(n4620), .Q(
        n8517) );
  SDFFX1 DFF_780_Q_reg ( .D(n280), .SI(n8517), .SE(n4177), .CLK(n4620), .Q(
        n8516) );
  SDFFX1 DFF_781_Q_reg ( .D(n281), .SI(n8516), .SE(n4177), .CLK(n4620), .Q(
        n8515) );
  SDFFX1 DFF_782_Q_reg ( .D(n282), .SI(n8515), .SE(n4178), .CLK(n4620), .Q(
        n8514) );
  SDFFX1 DFF_783_Q_reg ( .D(n283), .SI(n8514), .SE(n4178), .CLK(n4620), .Q(
        n8513) );
  SDFFX1 DFF_784_Q_reg ( .D(n284), .SI(n8513), .SE(n4178), .CLK(n4620), .Q(
        n8512) );
  SDFFX1 DFF_785_Q_reg ( .D(n285), .SI(n8512), .SE(n4178), .CLK(n4620), .Q(
        n8511) );
  SDFFX1 DFF_786_Q_reg ( .D(n286), .SI(n8511), .SE(n4178), .CLK(n4620), .Q(
        n8510) );
  SDFFX1 DFF_787_Q_reg ( .D(n287), .SI(n8510), .SE(n4178), .CLK(n4620), .Q(
        n8509) );
  SDFFX1 DFF_788_Q_reg ( .D(n288), .SI(n8509), .SE(n4179), .CLK(n4619), .Q(
        n8508) );
  SDFFX1 DFF_789_Q_reg ( .D(n289), .SI(n8508), .SE(n4179), .CLK(n4619), .Q(
        n8507) );
  SDFFX1 DFF_790_Q_reg ( .D(n290), .SI(n8507), .SE(n4179), .CLK(n4619), .Q(
        n8506) );
  SDFFX1 DFF_791_Q_reg ( .D(n291), .SI(n8506), .SE(n4179), .CLK(n4619), .Q(
        n8505) );
  SDFFX1 DFF_792_Q_reg ( .D(n292), .SI(n8505), .SE(n4179), .CLK(n4619), .Q(
        test_so45) );
  SDFFX1 DFF_793_Q_reg ( .D(n293), .SI(test_si46), .SE(n4179), .CLK(n4619), 
        .Q(n8502) );
  SDFFX1 DFF_794_Q_reg ( .D(n294), .SI(n8502), .SE(n4180), .CLK(n4619), .Q(
        n8501) );
  SDFFX1 DFF_795_Q_reg ( .D(n295), .SI(n8501), .SE(n4180), .CLK(n4619), .Q(
        n8500) );
  SDFFX1 DFF_796_Q_reg ( .D(n296), .SI(n8500), .SE(n4180), .CLK(n4619), .Q(
        n8499) );
  SDFFX1 DFF_797_Q_reg ( .D(n297), .SI(n8499), .SE(n4180), .CLK(n4619), .Q(
        n8498) );
  SDFFX1 DFF_798_Q_reg ( .D(n298), .SI(n8498), .SE(n4180), .CLK(n4619), .Q(
        n8497) );
  SDFFX1 DFF_799_Q_reg ( .D(WX5718), .SI(n8497), .SE(n4180), .CLK(n4619), .Q(
        n8496) );
  SDFFX1 DFF_800_Q_reg ( .D(WX5816), .SI(n8496), .SE(n4175), .CLK(n4621), .Q(
        n8495), .QN(n7193) );
  SDFFX1 DFF_801_Q_reg ( .D(WX5818), .SI(n8495), .SE(n4175), .CLK(n4621), .Q(
        n8494), .QN(n7192) );
  SDFFX1 DFF_802_Q_reg ( .D(WX5820), .SI(n8494), .SE(n4175), .CLK(n4621), .Q(
        n8493), .QN(n7191) );
  SDFFX1 DFF_803_Q_reg ( .D(WX5822), .SI(n8493), .SE(n4174), .CLK(n4622), .Q(
        n8492), .QN(n7190) );
  SDFFX1 DFF_804_Q_reg ( .D(WX5824), .SI(n8492), .SE(n4174), .CLK(n4622), .Q(
        n8491), .QN(n7189) );
  SDFFX1 DFF_805_Q_reg ( .D(WX5826), .SI(n8491), .SE(n4173), .CLK(n4622), .Q(
        n8490), .QN(n7188) );
  SDFFX1 DFF_806_Q_reg ( .D(WX5828), .SI(n8490), .SE(n4173), .CLK(n4622), .Q(
        n8489), .QN(n7187) );
  SDFFX1 DFF_807_Q_reg ( .D(WX5830), .SI(n8489), .SE(n4173), .CLK(n4622), .Q(
        n8488), .QN(n7186) );
  SDFFX1 DFF_808_Q_reg ( .D(WX5832), .SI(n8488), .SE(n4173), .CLK(n4622), .Q(
        n8487), .QN(n7185) );
  SDFFX1 DFF_809_Q_reg ( .D(WX5834), .SI(n8487), .SE(n4022), .CLK(n4698), .Q(
        test_so46) );
  SDFFX1 DFF_810_Q_reg ( .D(WX5836), .SI(test_si47), .SE(n4172), .CLK(n4623), 
        .Q(n8484), .QN(n7183) );
  SDFFX1 DFF_811_Q_reg ( .D(WX5838), .SI(n8484), .SE(n4172), .CLK(n4623), .Q(
        n8483), .QN(n7182) );
  SDFFX1 DFF_812_Q_reg ( .D(WX5840), .SI(n8483), .SE(n4022), .CLK(n4698), .Q(
        n8482), .QN(n7181) );
  SDFFX1 DFF_813_Q_reg ( .D(WX5842), .SI(n8482), .SE(n4171), .CLK(n4623), .Q(
        n8481), .QN(n7180) );
  SDFFX1 DFF_814_Q_reg ( .D(WX5844), .SI(n8481), .SE(n4218), .CLK(n4600), .Q(
        n8480), .QN(n7179) );
  SDFFX1 DFF_815_Q_reg ( .D(WX5846), .SI(n8480), .SE(n4170), .CLK(n4624), .Q(
        n8479), .QN(n7178) );
  SDFFX1 DFF_816_Q_reg ( .D(WX5848), .SI(n8479), .SE(n4170), .CLK(n4624), .Q(
        WX5849), .QN(n3359) );
  SDFFX1 DFF_817_Q_reg ( .D(WX5850), .SI(WX5849), .SE(n4169), .CLK(n4624), .Q(
        WX5851), .QN(n3358) );
  SDFFX1 DFF_818_Q_reg ( .D(WX5852), .SI(WX5851), .SE(n4168), .CLK(n4625), .Q(
        WX5853), .QN(n3357) );
  SDFFX1 DFF_819_Q_reg ( .D(WX5854), .SI(WX5853), .SE(n4168), .CLK(n4625), .Q(
        WX5855), .QN(n3356) );
  SDFFX1 DFF_820_Q_reg ( .D(WX5856), .SI(WX5855), .SE(n4167), .CLK(n4625), .Q(
        WX5857), .QN(n3355) );
  SDFFX1 DFF_821_Q_reg ( .D(WX5858), .SI(WX5857), .SE(n4166), .CLK(n4626), .Q(
        WX5859), .QN(n3354) );
  SDFFX1 DFF_822_Q_reg ( .D(WX5860), .SI(WX5859), .SE(n4166), .CLK(n4626), .Q(
        WX5861), .QN(n3353) );
  SDFFX1 DFF_823_Q_reg ( .D(WX5862), .SI(WX5861), .SE(n4165), .CLK(n4626), .Q(
        WX5863), .QN(n3352) );
  SDFFX1 DFF_824_Q_reg ( .D(WX5864), .SI(WX5863), .SE(n4164), .CLK(n4627), .Q(
        WX5865), .QN(n3351) );
  SDFFX1 DFF_825_Q_reg ( .D(WX5866), .SI(WX5865), .SE(n4164), .CLK(n4627), .Q(
        WX5867), .QN(n3350) );
  SDFFX1 DFF_826_Q_reg ( .D(WX5868), .SI(WX5867), .SE(n4163), .CLK(n4627), .Q(
        test_so47) );
  SDFFX1 DFF_827_Q_reg ( .D(WX5870), .SI(test_si48), .SE(n4022), .CLK(n4698), 
        .Q(WX5871), .QN(n3349) );
  SDFFX1 DFF_828_Q_reg ( .D(WX5872), .SI(WX5871), .SE(n4161), .CLK(n4628), .Q(
        WX5873) );
  SDFFX1 DFF_829_Q_reg ( .D(WX5874), .SI(WX5873), .SE(n4161), .CLK(n4628), .Q(
        WX5875), .QN(n3347) );
  SDFFX1 DFF_830_Q_reg ( .D(WX5876), .SI(WX5875), .SE(n4161), .CLK(n4628), .Q(
        WX5877) );
  SDFFX1 DFF_831_Q_reg ( .D(WX5878), .SI(WX5877), .SE(n4160), .CLK(n4629), .Q(
        WX5879), .QN(n3346) );
  SDFFX1 DFF_832_Q_reg ( .D(n299), .SI(WX5879), .SE(n4175), .CLK(n4621), .Q(
        WX5881), .QN(n3068) );
  SDFFX1 DFF_833_Q_reg ( .D(n300), .SI(WX5881), .SE(n4175), .CLK(n4621), .Q(
        WX5883), .QN(n3206) );
  SDFFX1 DFF_834_Q_reg ( .D(n301), .SI(WX5883), .SE(n4174), .CLK(n4622), .Q(
        WX5885), .QN(n3204) );
  SDFFX1 DFF_835_Q_reg ( .D(n302), .SI(WX5885), .SE(n4174), .CLK(n4622), .Q(
        WX5887), .QN(n3202) );
  SDFFX1 DFF_836_Q_reg ( .D(n303), .SI(WX5887), .SE(n4174), .CLK(n4622), .Q(
        WX5889), .QN(n3200) );
  SDFFX1 DFF_837_Q_reg ( .D(n304), .SI(WX5889), .SE(n4174), .CLK(n4622), .Q(
        WX5891), .QN(n3198) );
  SDFFX1 DFF_838_Q_reg ( .D(n305), .SI(WX5891), .SE(n4173), .CLK(n4622), .Q(
        WX5893), .QN(n3196) );
  SDFFX1 DFF_839_Q_reg ( .D(n306), .SI(WX5893), .SE(n4173), .CLK(n4622), .Q(
        WX5895), .QN(n3194) );
  SDFFX1 DFF_840_Q_reg ( .D(n307), .SI(WX5895), .SE(n4172), .CLK(n4623), .Q(
        WX5897), .QN(n3192) );
  SDFFX1 DFF_841_Q_reg ( .D(n308), .SI(WX5897), .SE(n4172), .CLK(n4623), .Q(
        WX5899), .QN(n3191) );
  SDFFX1 DFF_842_Q_reg ( .D(n309), .SI(WX5899), .SE(n4172), .CLK(n4623), .Q(
        WX5901), .QN(n3189) );
  SDFFX1 DFF_843_Q_reg ( .D(n310), .SI(WX5901), .SE(n4172), .CLK(n4623), .Q(
        test_so48) );
  SDFFX1 DFF_844_Q_reg ( .D(n311), .SI(test_si49), .SE(n4022), .CLK(n4698), 
        .Q(WX5905), .QN(n3186) );
  SDFFX1 DFF_845_Q_reg ( .D(n312), .SI(WX5905), .SE(n4171), .CLK(n4623), .Q(
        WX5907), .QN(n3185) );
  SDFFX1 DFF_846_Q_reg ( .D(n313), .SI(WX5907), .SE(n4171), .CLK(n4623), .Q(
        WX5909), .QN(n3183) );
  SDFFX1 DFF_847_Q_reg ( .D(n314), .SI(WX5909), .SE(n4170), .CLK(n4624), .Q(
        WX5911), .QN(n3182) );
  SDFFX1 DFF_848_Q_reg ( .D(WX5912), .SI(WX5911), .SE(n4170), .CLK(n4624), .Q(
        WX5913) );
  SDFFX1 DFF_849_Q_reg ( .D(WX5914), .SI(WX5913), .SE(n4169), .CLK(n4624), .Q(
        WX5915) );
  SDFFX1 DFF_850_Q_reg ( .D(WX5916), .SI(WX5915), .SE(n4168), .CLK(n4625), .Q(
        WX5917) );
  SDFFX1 DFF_851_Q_reg ( .D(WX5918), .SI(WX5917), .SE(n4168), .CLK(n4625), .Q(
        WX5919) );
  SDFFX1 DFF_852_Q_reg ( .D(WX5920), .SI(WX5919), .SE(n4167), .CLK(n4625), .Q(
        WX5921) );
  SDFFX1 DFF_853_Q_reg ( .D(WX5922), .SI(WX5921), .SE(n4166), .CLK(n4626), .Q(
        WX5923) );
  SDFFX1 DFF_854_Q_reg ( .D(WX5924), .SI(WX5923), .SE(n4166), .CLK(n4626), .Q(
        WX5925) );
  SDFFX1 DFF_855_Q_reg ( .D(WX5926), .SI(WX5925), .SE(n4165), .CLK(n4626), .Q(
        WX5927) );
  SDFFX1 DFF_856_Q_reg ( .D(WX5928), .SI(WX5927), .SE(n4164), .CLK(n4627), .Q(
        WX5929) );
  SDFFX1 DFF_857_Q_reg ( .D(WX5930), .SI(WX5929), .SE(n4164), .CLK(n4627), .Q(
        WX5931) );
  SDFFX1 DFF_858_Q_reg ( .D(WX5932), .SI(WX5931), .SE(n4163), .CLK(n4627), .Q(
        WX5933), .QN(n3669) );
  SDFFX1 DFF_859_Q_reg ( .D(WX5934), .SI(WX5933), .SE(n4162), .CLK(n4628), .Q(
        WX5935) );
  SDFFX1 DFF_860_Q_reg ( .D(WX5936), .SI(WX5935), .SE(n4162), .CLK(n4628), .Q(
        test_so49) );
  SDFFX1 DFF_861_Q_reg ( .D(WX5938), .SI(test_si50), .SE(n4161), .CLK(n4628), 
        .Q(WX5939), .QN(n3663) );
  SDFFX1 DFF_862_Q_reg ( .D(WX5940), .SI(WX5939), .SE(n4160), .CLK(n4629), .Q(
        WX5941), .QN(n3661) );
  SDFFX1 DFF_863_Q_reg ( .D(WX5942), .SI(WX5941), .SE(n4160), .CLK(n4629), .Q(
        WX5943) );
  SDFFX1 DFF_864_Q_reg ( .D(WX5944), .SI(WX5943), .SE(n4159), .CLK(n4629), .Q(
        WX5945) );
  SDFFX1 DFF_865_Q_reg ( .D(WX5946), .SI(WX5945), .SE(n4159), .CLK(n4629), .Q(
        WX5947) );
  SDFFX1 DFF_866_Q_reg ( .D(WX5948), .SI(WX5947), .SE(n4159), .CLK(n4629), .Q(
        WX5949) );
  SDFFX1 DFF_867_Q_reg ( .D(WX5950), .SI(WX5949), .SE(n4158), .CLK(n4630), .Q(
        WX5951) );
  SDFFX1 DFF_868_Q_reg ( .D(WX5952), .SI(WX5951), .SE(n4158), .CLK(n4630), .Q(
        WX5953) );
  SDFFX1 DFF_869_Q_reg ( .D(WX5954), .SI(WX5953), .SE(n4158), .CLK(n4630), .Q(
        WX5955) );
  SDFFX1 DFF_870_Q_reg ( .D(WX5956), .SI(WX5955), .SE(n4157), .CLK(n4630), .Q(
        WX5957) );
  SDFFX1 DFF_871_Q_reg ( .D(WX5958), .SI(WX5957), .SE(n4157), .CLK(n4630), .Q(
        WX5959) );
  SDFFX1 DFF_872_Q_reg ( .D(WX5960), .SI(WX5959), .SE(n4157), .CLK(n4630), .Q(
        WX5961) );
  SDFFX1 DFF_873_Q_reg ( .D(WX5962), .SI(WX5961), .SE(n4156), .CLK(n4631), .Q(
        WX5963), .QN(n7184) );
  SDFFX1 DFF_874_Q_reg ( .D(WX5964), .SI(WX5963), .SE(n4156), .CLK(n4631), .Q(
        WX5965) );
  SDFFX1 DFF_875_Q_reg ( .D(WX5966), .SI(WX5965), .SE(n4171), .CLK(n4623), .Q(
        WX5967), .QN(n3188) );
  SDFFX1 DFF_876_Q_reg ( .D(WX5968), .SI(WX5967), .SE(n4171), .CLK(n4623), .Q(
        WX5969) );
  SDFFX1 DFF_877_Q_reg ( .D(WX5970), .SI(WX5969), .SE(n4171), .CLK(n4623), .Q(
        test_so50) );
  SDFFX1 DFF_878_Q_reg ( .D(WX5972), .SI(test_si51), .SE(n4170), .CLK(n4624), 
        .Q(WX5973) );
  SDFFX1 DFF_879_Q_reg ( .D(WX5974), .SI(WX5973), .SE(n4170), .CLK(n4624), .Q(
        WX5975) );
  SDFFX1 DFF_880_Q_reg ( .D(WX5976), .SI(WX5975), .SE(n4169), .CLK(n4624), .Q(
        WX5977), .QN(n7177) );
  SDFFX1 DFF_881_Q_reg ( .D(WX5978), .SI(WX5977), .SE(n4169), .CLK(n4624), .Q(
        WX5979), .QN(n7176) );
  SDFFX1 DFF_882_Q_reg ( .D(WX5980), .SI(WX5979), .SE(n4168), .CLK(n4625), .Q(
        WX5981), .QN(n7175) );
  SDFFX1 DFF_883_Q_reg ( .D(WX5982), .SI(WX5981), .SE(n4167), .CLK(n4625), .Q(
        WX5983), .QN(n7174) );
  SDFFX1 DFF_884_Q_reg ( .D(WX5984), .SI(WX5983), .SE(n4167), .CLK(n4625), .Q(
        WX5985), .QN(n7173) );
  SDFFX1 DFF_885_Q_reg ( .D(WX5986), .SI(WX5985), .SE(n4166), .CLK(n4626), .Q(
        WX5987), .QN(n7172) );
  SDFFX1 DFF_886_Q_reg ( .D(WX5988), .SI(WX5987), .SE(n4165), .CLK(n4626), .Q(
        WX5989), .QN(n7171) );
  SDFFX1 DFF_887_Q_reg ( .D(WX5990), .SI(WX5989), .SE(n4165), .CLK(n4626), .Q(
        WX5991), .QN(n7170) );
  SDFFX1 DFF_888_Q_reg ( .D(WX5992), .SI(WX5991), .SE(n4164), .CLK(n4627), .Q(
        WX5993), .QN(n7169) );
  SDFFX1 DFF_889_Q_reg ( .D(WX5994), .SI(WX5993), .SE(n4163), .CLK(n4627), .Q(
        WX5995), .QN(n7168) );
  SDFFX1 DFF_890_Q_reg ( .D(WX5996), .SI(WX5995), .SE(n4163), .CLK(n4627), .Q(
        WX5997) );
  SDFFX1 DFF_891_Q_reg ( .D(WX5998), .SI(WX5997), .SE(n4162), .CLK(n4628), .Q(
        WX5999), .QN(n7167) );
  SDFFX1 DFF_892_Q_reg ( .D(WX6000), .SI(WX5999), .SE(n4162), .CLK(n4628), .Q(
        WX6001), .QN(n3348) );
  SDFFX1 DFF_893_Q_reg ( .D(WX6002), .SI(WX6001), .SE(n4161), .CLK(n4628), .Q(
        WX6003) );
  SDFFX1 DFF_894_Q_reg ( .D(WX6004), .SI(WX6003), .SE(n4160), .CLK(n4629), .Q(
        test_so51) );
  SDFFX1 DFF_895_Q_reg ( .D(WX6006), .SI(test_si52), .SE(n4160), .CLK(n4629), 
        .Q(WX6007), .QN(n7166) );
  SDFFX1 DFF_896_Q_reg ( .D(WX6008), .SI(WX6007), .SE(n4159), .CLK(n4629), .Q(
        WX6009), .QN(n3618) );
  SDFFX1 DFF_897_Q_reg ( .D(WX6010), .SI(WX6009), .SE(n4159), .CLK(n4629), .Q(
        WX6011), .QN(n3620) );
  SDFFX1 DFF_898_Q_reg ( .D(WX6012), .SI(WX6011), .SE(n4158), .CLK(n4630), .Q(
        WX6013), .QN(n3621) );
  SDFFX1 DFF_899_Q_reg ( .D(WX6014), .SI(WX6013), .SE(n4158), .CLK(n4630), .Q(
        WX6015), .QN(n3622) );
  SDFFX1 DFF_900_Q_reg ( .D(WX6016), .SI(WX6015), .SE(n4158), .CLK(n4630), .Q(
        WX6017), .QN(n3624) );
  SDFFX1 DFF_901_Q_reg ( .D(WX6018), .SI(WX6017), .SE(n4157), .CLK(n4630), .Q(
        WX6019), .QN(n3626) );
  SDFFX1 DFF_902_Q_reg ( .D(WX6020), .SI(WX6019), .SE(n4157), .CLK(n4630), .Q(
        WX6021), .QN(n3628) );
  SDFFX1 DFF_903_Q_reg ( .D(WX6022), .SI(WX6021), .SE(n4157), .CLK(n4630), .Q(
        WX6023), .QN(n3630) );
  SDFFX1 DFF_904_Q_reg ( .D(WX6024), .SI(WX6023), .SE(n4156), .CLK(n4631), .Q(
        WX6025), .QN(n3632) );
  SDFFX1 DFF_905_Q_reg ( .D(WX6026), .SI(WX6025), .SE(n4156), .CLK(n4631), .Q(
        WX6027), .QN(n3634) );
  SDFFX1 DFF_906_Q_reg ( .D(WX6028), .SI(WX6027), .SE(n4156), .CLK(n4631), .Q(
        WX6029), .QN(n3636) );
  SDFFX1 DFF_907_Q_reg ( .D(WX6030), .SI(WX6029), .SE(n4156), .CLK(n4631), .Q(
        WX6031), .QN(n3638) );
  SDFFX1 DFF_908_Q_reg ( .D(WX6032), .SI(WX6031), .SE(n4155), .CLK(n4631), .Q(
        WX6033), .QN(n3640) );
  SDFFX1 DFF_909_Q_reg ( .D(WX6034), .SI(WX6033), .SE(n4155), .CLK(n4631), .Q(
        WX6035), .QN(n3642) );
  SDFFX1 DFF_910_Q_reg ( .D(WX6036), .SI(WX6035), .SE(n4155), .CLK(n4631), .Q(
        WX6037), .QN(n3643) );
  SDFFX1 DFF_911_Q_reg ( .D(WX6038), .SI(WX6037), .SE(n4155), .CLK(n4631), .Q(
        test_so52) );
  SDFFX1 DFF_912_Q_reg ( .D(WX6040), .SI(test_si53), .SE(n4169), .CLK(n4624), 
        .Q(WX6041), .QN(n3644) );
  SDFFX1 DFF_913_Q_reg ( .D(WX6042), .SI(WX6041), .SE(n4169), .CLK(n4624), .Q(
        WX6043), .QN(n3646) );
  SDFFX1 DFF_914_Q_reg ( .D(WX6044), .SI(WX6043), .SE(n4168), .CLK(n4625), .Q(
        WX6045), .QN(n3648) );
  SDFFX1 DFF_915_Q_reg ( .D(WX6046), .SI(WX6045), .SE(n4167), .CLK(n4625), .Q(
        WX6047), .QN(n3650) );
  SDFFX1 DFF_916_Q_reg ( .D(WX6048), .SI(WX6047), .SE(n4167), .CLK(n4625), .Q(
        WX6049), .QN(n3423) );
  SDFFX1 DFF_917_Q_reg ( .D(WX6050), .SI(WX6049), .SE(n4166), .CLK(n4626), .Q(
        WX6051), .QN(n3652) );
  SDFFX1 DFF_918_Q_reg ( .D(WX6052), .SI(WX6051), .SE(n4165), .CLK(n4626), .Q(
        WX6053), .QN(n3654) );
  SDFFX1 DFF_919_Q_reg ( .D(WX6054), .SI(WX6053), .SE(n4165), .CLK(n4626), .Q(
        WX6055), .QN(n3656) );
  SDFFX1 DFF_920_Q_reg ( .D(WX6056), .SI(WX6055), .SE(n4164), .CLK(n4627), .Q(
        WX6057), .QN(n3658) );
  SDFFX1 DFF_921_Q_reg ( .D(WX6058), .SI(WX6057), .SE(n4163), .CLK(n4627), .Q(
        WX6059), .QN(n3660) );
  SDFFX1 DFF_922_Q_reg ( .D(WX6060), .SI(WX6059), .SE(n4163), .CLK(n4627), .Q(
        WX6061), .QN(n3662) );
  SDFFX1 DFF_923_Q_reg ( .D(WX6062), .SI(WX6061), .SE(n4162), .CLK(n4628), .Q(
        WX6063), .QN(n3424) );
  SDFFX1 DFF_924_Q_reg ( .D(WX6064), .SI(WX6063), .SE(n4162), .CLK(n4628), .Q(
        WX6065), .QN(n3664) );
  SDFFX1 DFF_925_Q_reg ( .D(WX6066), .SI(WX6065), .SE(n4161), .CLK(n4628), .Q(
        WX6067), .QN(n3665) );
  SDFFX1 DFF_926_Q_reg ( .D(WX6068), .SI(WX6067), .SE(n4160), .CLK(n4629), .Q(
        WX6069), .QN(n3666) );
  SDFFX1 DFF_927_Q_reg ( .D(WX6070), .SI(WX6069), .SE(n4159), .CLK(n4629), .Q(
        WX6071), .QN(n3437) );
  SDFFX1 DFF_928_Q_reg ( .D(WX6436), .SI(WX6071), .SE(n4026), .CLK(n4696), .Q(
        test_so53) );
  SDFFX1 DFF_929_Q_reg ( .D(WX6438), .SI(test_si54), .SE(n4026), .CLK(n4696), 
        .Q(CRC_OUT_5_1), .QN(DFF_929_n1) );
  SDFFX1 DFF_930_Q_reg ( .D(WX6440), .SI(CRC_OUT_5_1), .SE(n4025), .CLK(n4696), 
        .Q(CRC_OUT_5_2), .QN(DFF_930_n1) );
  SDFFX1 DFF_931_Q_reg ( .D(WX6442), .SI(CRC_OUT_5_2), .SE(n4025), .CLK(n4696), 
        .Q(CRC_OUT_5_3) );
  SDFFX1 DFF_932_Q_reg ( .D(WX6444), .SI(CRC_OUT_5_3), .SE(n4025), .CLK(n4696), 
        .Q(CRC_OUT_5_4), .QN(DFF_932_n1) );
  SDFFX1 DFF_933_Q_reg ( .D(WX6446), .SI(CRC_OUT_5_4), .SE(n4025), .CLK(n4696), 
        .Q(CRC_OUT_5_5), .QN(DFF_933_n1) );
  SDFFX1 DFF_934_Q_reg ( .D(WX6448), .SI(CRC_OUT_5_5), .SE(n4025), .CLK(n4696), 
        .Q(CRC_OUT_5_6), .QN(DFF_934_n1) );
  SDFFX1 DFF_935_Q_reg ( .D(WX6450), .SI(CRC_OUT_5_6), .SE(n4025), .CLK(n4696), 
        .Q(CRC_OUT_5_7), .QN(DFF_935_n1) );
  SDFFX1 DFF_936_Q_reg ( .D(WX6452), .SI(CRC_OUT_5_7), .SE(n4024), .CLK(n4697), 
        .Q(CRC_OUT_5_8), .QN(DFF_936_n1) );
  SDFFX1 DFF_937_Q_reg ( .D(WX6454), .SI(CRC_OUT_5_8), .SE(n4024), .CLK(n4697), 
        .Q(CRC_OUT_5_9), .QN(DFF_937_n1) );
  SDFFX1 DFF_938_Q_reg ( .D(WX6456), .SI(CRC_OUT_5_9), .SE(n4024), .CLK(n4697), 
        .Q(CRC_OUT_5_10) );
  SDFFX1 DFF_939_Q_reg ( .D(WX6458), .SI(CRC_OUT_5_10), .SE(n4024), .CLK(n4697), .Q(CRC_OUT_5_11), .QN(DFF_939_n1) );
  SDFFX1 DFF_940_Q_reg ( .D(WX6460), .SI(CRC_OUT_5_11), .SE(n4024), .CLK(n4697), .Q(CRC_OUT_5_12), .QN(DFF_940_n1) );
  SDFFX1 DFF_941_Q_reg ( .D(WX6462), .SI(CRC_OUT_5_12), .SE(n4024), .CLK(n4697), .Q(CRC_OUT_5_13), .QN(DFF_941_n1) );
  SDFFX1 DFF_942_Q_reg ( .D(WX6464), .SI(CRC_OUT_5_13), .SE(n4023), .CLK(n4697), .Q(CRC_OUT_5_14), .QN(DFF_942_n1) );
  SDFFX1 DFF_943_Q_reg ( .D(WX6466), .SI(CRC_OUT_5_14), .SE(n4023), .CLK(n4697), .Q(CRC_OUT_5_15), .QN(DFF_943_n1) );
  SDFFX1 DFF_944_Q_reg ( .D(WX6468), .SI(CRC_OUT_5_15), .SE(n4023), .CLK(n4697), .Q(CRC_OUT_5_16), .QN(DFF_944_n1) );
  SDFFX1 DFF_945_Q_reg ( .D(WX6470), .SI(CRC_OUT_5_16), .SE(n4023), .CLK(n4697), .Q(test_so54) );
  SDFFX1 DFF_946_Q_reg ( .D(WX6472), .SI(test_si55), .SE(n4023), .CLK(n4697), 
        .Q(CRC_OUT_5_18), .QN(DFF_946_n1) );
  SDFFX1 DFF_947_Q_reg ( .D(WX6474), .SI(CRC_OUT_5_18), .SE(n4023), .CLK(n4697), .Q(CRC_OUT_5_19), .QN(DFF_947_n1) );
  SDFFX1 DFF_948_Q_reg ( .D(WX6476), .SI(CRC_OUT_5_19), .SE(n4022), .CLK(n4698), .Q(CRC_OUT_5_20), .QN(DFF_948_n1) );
  SDFFX1 DFF_949_Q_reg ( .D(WX6478), .SI(CRC_OUT_5_20), .SE(n4155), .CLK(n4631), .Q(CRC_OUT_5_21), .QN(DFF_949_n1) );
  SDFFX1 DFF_950_Q_reg ( .D(WX6480), .SI(CRC_OUT_5_21), .SE(n4155), .CLK(n4631), .Q(CRC_OUT_5_22), .QN(DFF_950_n1) );
  SDFFX1 DFF_951_Q_reg ( .D(WX6482), .SI(CRC_OUT_5_22), .SE(n4154), .CLK(n4632), .Q(CRC_OUT_5_23), .QN(DFF_951_n1) );
  SDFFX1 DFF_952_Q_reg ( .D(WX6484), .SI(CRC_OUT_5_23), .SE(n4154), .CLK(n4632), .Q(CRC_OUT_5_24), .QN(DFF_952_n1) );
  SDFFX1 DFF_953_Q_reg ( .D(WX6486), .SI(CRC_OUT_5_24), .SE(n4154), .CLK(n4632), .Q(CRC_OUT_5_25), .QN(DFF_953_n1) );
  SDFFX1 DFF_954_Q_reg ( .D(WX6488), .SI(CRC_OUT_5_25), .SE(n4154), .CLK(n4632), .Q(CRC_OUT_5_26), .QN(DFF_954_n1) );
  SDFFX1 DFF_955_Q_reg ( .D(WX6490), .SI(CRC_OUT_5_26), .SE(n4154), .CLK(n4632), .Q(CRC_OUT_5_27), .QN(DFF_955_n1) );
  SDFFX1 DFF_956_Q_reg ( .D(WX6492), .SI(CRC_OUT_5_27), .SE(n4154), .CLK(n4632), .Q(CRC_OUT_5_28), .QN(DFF_956_n1) );
  SDFFX1 DFF_957_Q_reg ( .D(WX6494), .SI(CRC_OUT_5_28), .SE(n4153), .CLK(n4632), .Q(CRC_OUT_5_29), .QN(DFF_957_n1) );
  SDFFX1 DFF_958_Q_reg ( .D(WX6496), .SI(CRC_OUT_5_29), .SE(n4153), .CLK(n4632), .Q(CRC_OUT_5_30), .QN(DFF_958_n1) );
  SDFFX1 DFF_959_Q_reg ( .D(WX6498), .SI(CRC_OUT_5_30), .SE(n4153), .CLK(n4632), .Q(CRC_OUT_5_31), .QN(DFF_959_n1) );
  SDFFX1 DFF_960_Q_reg ( .D(n346), .SI(CRC_OUT_5_31), .SE(n4153), .CLK(n4632), 
        .Q(WX6950) );
  SDFFX1 DFF_961_Q_reg ( .D(n347), .SI(WX6950), .SE(n4148), .CLK(n4635), .Q(
        n8470) );
  SDFFX1 DFF_962_Q_reg ( .D(n348), .SI(n8470), .SE(n4148), .CLK(n4635), .Q(
        test_so55) );
  SDFFX1 DFF_963_Q_reg ( .D(n349), .SI(test_si56), .SE(n4148), .CLK(n4635), 
        .Q(n8467) );
  SDFFX1 DFF_964_Q_reg ( .D(n350), .SI(n8467), .SE(n4148), .CLK(n4635), .Q(
        n8466) );
  SDFFX1 DFF_965_Q_reg ( .D(n351), .SI(n8466), .SE(n4148), .CLK(n4635), .Q(
        n8465) );
  SDFFX1 DFF_966_Q_reg ( .D(n352), .SI(n8465), .SE(n4149), .CLK(n4634), .Q(
        n8464) );
  SDFFX1 DFF_967_Q_reg ( .D(n353), .SI(n8464), .SE(n4149), .CLK(n4634), .Q(
        n8463) );
  SDFFX1 DFF_968_Q_reg ( .D(n354), .SI(n8463), .SE(n4149), .CLK(n4634), .Q(
        n8462) );
  SDFFX1 DFF_969_Q_reg ( .D(n355), .SI(n8462), .SE(n4149), .CLK(n4634), .Q(
        n8461) );
  SDFFX1 DFF_970_Q_reg ( .D(n356), .SI(n8461), .SE(n4149), .CLK(n4634), .Q(
        n8460) );
  SDFFX1 DFF_971_Q_reg ( .D(n357), .SI(n8460), .SE(n4149), .CLK(n4634), .Q(
        n8459) );
  SDFFX1 DFF_972_Q_reg ( .D(n358), .SI(n8459), .SE(n4150), .CLK(n4634), .Q(
        n8458) );
  SDFFX1 DFF_973_Q_reg ( .D(n359), .SI(n8458), .SE(n4150), .CLK(n4634), .Q(
        n8457) );
  SDFFX1 DFF_974_Q_reg ( .D(n360), .SI(n8457), .SE(n4150), .CLK(n4634), .Q(
        n8456) );
  SDFFX1 DFF_975_Q_reg ( .D(n361), .SI(n8456), .SE(n4150), .CLK(n4634), .Q(
        n8455) );
  SDFFX1 DFF_976_Q_reg ( .D(n362), .SI(n8455), .SE(n4150), .CLK(n4634), .Q(
        n8454) );
  SDFFX1 DFF_977_Q_reg ( .D(n363), .SI(n8454), .SE(n4150), .CLK(n4634), .Q(
        n8453) );
  SDFFX1 DFF_978_Q_reg ( .D(n364), .SI(n8453), .SE(n4151), .CLK(n4633), .Q(
        n8452) );
  SDFFX1 DFF_979_Q_reg ( .D(n365), .SI(n8452), .SE(n4151), .CLK(n4633), .Q(
        test_so56) );
  SDFFX1 DFF_980_Q_reg ( .D(n366), .SI(test_si57), .SE(n4151), .CLK(n4633), 
        .Q(n8449) );
  SDFFX1 DFF_981_Q_reg ( .D(n367), .SI(n8449), .SE(n4151), .CLK(n4633), .Q(
        n8448) );
  SDFFX1 DFF_982_Q_reg ( .D(n368), .SI(n8448), .SE(n4151), .CLK(n4633), .Q(
        n8447) );
  SDFFX1 DFF_983_Q_reg ( .D(n369), .SI(n8447), .SE(n4151), .CLK(n4633), .Q(
        n8446) );
  SDFFX1 DFF_984_Q_reg ( .D(n370), .SI(n8446), .SE(n4152), .CLK(n4633), .Q(
        n8445) );
  SDFFX1 DFF_985_Q_reg ( .D(WX6999), .SI(n8445), .SE(n4152), .CLK(n4633), .Q(
        n8444) );
  SDFFX1 DFF_986_Q_reg ( .D(n372), .SI(n8444), .SE(n4152), .CLK(n4633), .Q(
        n8443), .QN(n3871) );
  SDFFX1 DFF_987_Q_reg ( .D(n373), .SI(n8443), .SE(n4152), .CLK(n4633), .Q(
        n8442) );
  SDFFX1 DFF_988_Q_reg ( .D(n374), .SI(n8442), .SE(n4152), .CLK(n4633), .Q(
        n8441) );
  SDFFX1 DFF_989_Q_reg ( .D(n375), .SI(n8441), .SE(n4152), .CLK(n4633), .Q(
        n8440) );
  SDFFX1 DFF_990_Q_reg ( .D(n376), .SI(n8440), .SE(n4153), .CLK(n4632), .Q(
        n8439) );
  SDFFX1 DFF_991_Q_reg ( .D(WX7011), .SI(n8439), .SE(n4153), .CLK(n4632), .Q(
        n8438) );
  SDFFX1 DFF_992_Q_reg ( .D(WX7109), .SI(n8438), .SE(n4148), .CLK(n4635), .Q(
        n8437), .QN(n7165) );
  SDFFX1 DFF_993_Q_reg ( .D(WX7111), .SI(n8437), .SE(n4147), .CLK(n4635), .Q(
        n8436), .QN(n7164) );
  SDFFX1 DFF_994_Q_reg ( .D(WX7113), .SI(n8436), .SE(n4147), .CLK(n4635), .Q(
        n8435), .QN(n7163) );
  SDFFX1 DFF_995_Q_reg ( .D(WX7115), .SI(n8435), .SE(n4146), .CLK(n4636), .Q(
        n8434), .QN(n7162) );
  SDFFX1 DFF_996_Q_reg ( .D(WX7117), .SI(n8434), .SE(n4146), .CLK(n4636), .Q(
        test_so57) );
  SDFFX1 DFF_997_Q_reg ( .D(WX7119), .SI(test_si58), .SE(n4146), .CLK(n4636), 
        .Q(n8431), .QN(n7160) );
  SDFFX1 DFF_998_Q_reg ( .D(WX7121), .SI(n8431), .SE(n4146), .CLK(n4636), .Q(
        n8430), .QN(n7159) );
  SDFFX1 DFF_999_Q_reg ( .D(WX7123), .SI(n8430), .SE(n4026), .CLK(n4696), .Q(
        n8429), .QN(n7158) );
  SDFFX1 DFF_1000_Q_reg ( .D(WX7125), .SI(n8429), .SE(n4145), .CLK(n4636), .Q(
        n8428), .QN(n7157) );
  SDFFX1 DFF_1001_Q_reg ( .D(WX7127), .SI(n8428), .SE(n4144), .CLK(n4637), .Q(
        n8427), .QN(n7156) );
  SDFFX1 DFF_1002_Q_reg ( .D(WX7129), .SI(n8427), .SE(n4144), .CLK(n4637), .Q(
        n8426), .QN(n7155) );
  SDFFX1 DFF_1003_Q_reg ( .D(WX7131), .SI(n8426), .SE(n4143), .CLK(n4637), .Q(
        n8425), .QN(n7154) );
  SDFFX1 DFF_1004_Q_reg ( .D(WX7133), .SI(n8425), .SE(n4143), .CLK(n4637), .Q(
        n8424), .QN(n7153) );
  SDFFX1 DFF_1005_Q_reg ( .D(WX7135), .SI(n8424), .SE(n4026), .CLK(n4696), .Q(
        n8423), .QN(n7152) );
  SDFFX1 DFF_1006_Q_reg ( .D(WX7137), .SI(n8423), .SE(n4218), .CLK(n4600), .Q(
        n8422), .QN(n7151) );
  SDFFX1 DFF_1007_Q_reg ( .D(WX7139), .SI(n8422), .SE(n4141), .CLK(n4638), .Q(
        n8421), .QN(n7150) );
  SDFFX1 DFF_1008_Q_reg ( .D(WX7141), .SI(n8421), .SE(n4140), .CLK(n4639), .Q(
        WX7142), .QN(n3345) );
  SDFFX1 DFF_1009_Q_reg ( .D(WX7143), .SI(WX7142), .SE(n4140), .CLK(n4639), 
        .Q(WX7144), .QN(n3344) );
  SDFFX1 DFF_1010_Q_reg ( .D(WX7145), .SI(WX7144), .SE(n4139), .CLK(n4639), 
        .Q(WX7146), .QN(n3343) );
  SDFFX1 DFF_1011_Q_reg ( .D(WX7147), .SI(WX7146), .SE(n4138), .CLK(n4640), 
        .Q(WX7148), .QN(n3342) );
  SDFFX1 DFF_1012_Q_reg ( .D(WX7149), .SI(WX7148), .SE(n4138), .CLK(n4640), 
        .Q(WX7150), .QN(n3341) );
  SDFFX1 DFF_1013_Q_reg ( .D(WX7151), .SI(WX7150), .SE(n4137), .CLK(n4640), 
        .Q(test_so58) );
  SDFFX1 DFF_1014_Q_reg ( .D(WX7153), .SI(test_si59), .SE(n4026), .CLK(n4696), 
        .Q(WX7154), .QN(n3340) );
  SDFFX1 DFF_1015_Q_reg ( .D(WX7155), .SI(WX7154), .SE(n4135), .CLK(n4641), 
        .Q(WX7156) );
  SDFFX1 DFF_1016_Q_reg ( .D(WX7157), .SI(WX7156), .SE(n4135), .CLK(n4641), 
        .Q(WX7158), .QN(n3338) );
  SDFFX1 DFF_1017_Q_reg ( .D(WX7159), .SI(WX7158), .SE(n4135), .CLK(n4641), 
        .Q(WX7160) );
  SDFFX1 DFF_1018_Q_reg ( .D(WX7161), .SI(WX7160), .SE(n4134), .CLK(n4642), 
        .Q(WX7162), .QN(n3337) );
  SDFFX1 DFF_1019_Q_reg ( .D(WX7163), .SI(WX7162), .SE(n4133), .CLK(n4642), 
        .Q(WX7164) );
  SDFFX1 DFF_1020_Q_reg ( .D(WX7165), .SI(WX7164), .SE(n4133), .CLK(n4642), 
        .Q(WX7166), .QN(n3335) );
  SDFFX1 DFF_1021_Q_reg ( .D(WX7167), .SI(WX7166), .SE(n4132), .CLK(n4643), 
        .Q(WX7168), .QN(n3334) );
  SDFFX1 DFF_1022_Q_reg ( .D(WX7169), .SI(WX7168), .SE(n4131), .CLK(n4643), 
        .Q(WX7170), .QN(n3333) );
  SDFFX1 DFF_1023_Q_reg ( .D(WX7171), .SI(WX7170), .SE(n4131), .CLK(n4643), 
        .Q(WX7172), .QN(n3332) );
  SDFFX1 DFF_1024_Q_reg ( .D(n377), .SI(WX7172), .SE(n4147), .CLK(n4635), .Q(
        WX7174), .QN(n3066) );
  SDFFX1 DFF_1025_Q_reg ( .D(n378), .SI(WX7174), .SE(n4147), .CLK(n4635), .Q(
        WX7176), .QN(n3180) );
  SDFFX1 DFF_1026_Q_reg ( .D(n379), .SI(WX7176), .SE(n4147), .CLK(n4635), .Q(
        WX7178), .QN(n3178) );
  SDFFX1 DFF_1027_Q_reg ( .D(n380), .SI(WX7178), .SE(n4147), .CLK(n4635), .Q(
        WX7180), .QN(n3176) );
  SDFFX1 DFF_1028_Q_reg ( .D(n381), .SI(WX7180), .SE(n4146), .CLK(n4636), .Q(
        WX7182), .QN(n3175) );
  SDFFX1 DFF_1029_Q_reg ( .D(n382), .SI(WX7182), .SE(n4146), .CLK(n4636), .Q(
        WX7184), .QN(n3173) );
  SDFFX1 DFF_1030_Q_reg ( .D(n383), .SI(WX7184), .SE(n4145), .CLK(n4636), .Q(
        test_so59) );
  SDFFX1 DFF_1031_Q_reg ( .D(n384), .SI(test_si60), .SE(n4026), .CLK(n4696), 
        .Q(WX7188), .QN(n3170) );
  SDFFX1 DFF_1032_Q_reg ( .D(n385), .SI(WX7188), .SE(n4145), .CLK(n4636), .Q(
        WX7190), .QN(n3169) );
  SDFFX1 DFF_1033_Q_reg ( .D(n386), .SI(WX7190), .SE(n4144), .CLK(n4637), .Q(
        WX7192), .QN(n3167) );
  SDFFX1 DFF_1034_Q_reg ( .D(n387), .SI(WX7192), .SE(n4144), .CLK(n4637), .Q(
        WX7194), .QN(n3166) );
  SDFFX1 DFF_1035_Q_reg ( .D(n388), .SI(WX7194), .SE(n4143), .CLK(n4637), .Q(
        WX7196), .QN(n3164) );
  SDFFX1 DFF_1036_Q_reg ( .D(n389), .SI(WX7196), .SE(n4143), .CLK(n4637), .Q(
        WX7198), .QN(n3162) );
  SDFFX1 DFF_1037_Q_reg ( .D(n390), .SI(WX7198), .SE(n4142), .CLK(n4638), .Q(
        WX7200), .QN(n3160) );
  SDFFX1 DFF_1038_Q_reg ( .D(n391), .SI(WX7200), .SE(n4142), .CLK(n4638), .Q(
        WX7202), .QN(n3158) );
  SDFFX1 DFF_1039_Q_reg ( .D(n392), .SI(WX7202), .SE(n4141), .CLK(n4638), .Q(
        WX7204), .QN(n3156) );
  SDFFX1 DFF_1040_Q_reg ( .D(WX7205), .SI(WX7204), .SE(n4140), .CLK(n4639), 
        .Q(WX7206) );
  SDFFX1 DFF_1041_Q_reg ( .D(WX7207), .SI(WX7206), .SE(n4140), .CLK(n4639), 
        .Q(WX7208) );
  SDFFX1 DFF_1042_Q_reg ( .D(WX7209), .SI(WX7208), .SE(n4139), .CLK(n4639), 
        .Q(WX7210) );
  SDFFX1 DFF_1043_Q_reg ( .D(WX7211), .SI(WX7210), .SE(n4138), .CLK(n4640), 
        .Q(WX7212) );
  SDFFX1 DFF_1044_Q_reg ( .D(WX7213), .SI(WX7212), .SE(n4138), .CLK(n4640), 
        .Q(WX7214) );
  SDFFX1 DFF_1045_Q_reg ( .D(WX7215), .SI(WX7214), .SE(n4137), .CLK(n4640), 
        .Q(WX7216), .QN(n3647) );
  SDFFX1 DFF_1046_Q_reg ( .D(WX7217), .SI(WX7216), .SE(n4136), .CLK(n4641), 
        .Q(WX7218) );
  SDFFX1 DFF_1047_Q_reg ( .D(WX7219), .SI(WX7218), .SE(n4136), .CLK(n4641), 
        .Q(test_so60) );
  SDFFX1 DFF_1048_Q_reg ( .D(WX7221), .SI(test_si61), .SE(n4135), .CLK(n4641), 
        .Q(WX7222) );
  SDFFX1 DFF_1049_Q_reg ( .D(WX7223), .SI(WX7222), .SE(n4134), .CLK(n4642), 
        .Q(WX7224), .QN(n3639) );
  SDFFX1 DFF_1050_Q_reg ( .D(WX7225), .SI(WX7224), .SE(n4134), .CLK(n4642), 
        .Q(WX7226) );
  SDFFX1 DFF_1051_Q_reg ( .D(WX7227), .SI(WX7226), .SE(n4133), .CLK(n4642), 
        .Q(WX7228), .QN(n3635) );
  SDFFX1 DFF_1052_Q_reg ( .D(WX7229), .SI(WX7228), .SE(n4132), .CLK(n4643), 
        .Q(WX7230) );
  SDFFX1 DFF_1053_Q_reg ( .D(WX7231), .SI(WX7230), .SE(n4132), .CLK(n4643), 
        .Q(WX7232) );
  SDFFX1 DFF_1054_Q_reg ( .D(WX7233), .SI(WX7232), .SE(n4131), .CLK(n4643), 
        .Q(WX7234) );
  SDFFX1 DFF_1055_Q_reg ( .D(WX7235), .SI(WX7234), .SE(n4130), .CLK(n4644), 
        .Q(WX7236) );
  SDFFX1 DFF_1056_Q_reg ( .D(WX7237), .SI(WX7236), .SE(n4130), .CLK(n4644), 
        .Q(WX7238) );
  SDFFX1 DFF_1057_Q_reg ( .D(WX7239), .SI(WX7238), .SE(n4130), .CLK(n4644), 
        .Q(WX7240) );
  SDFFX1 DFF_1058_Q_reg ( .D(WX7241), .SI(WX7240), .SE(n4129), .CLK(n4644), 
        .Q(WX7242) );
  SDFFX1 DFF_1059_Q_reg ( .D(WX7243), .SI(WX7242), .SE(n4129), .CLK(n4644), 
        .Q(WX7244) );
  SDFFX1 DFF_1060_Q_reg ( .D(WX7245), .SI(WX7244), .SE(n4129), .CLK(n4644), 
        .Q(WX7246), .QN(n7161) );
  SDFFX1 DFF_1061_Q_reg ( .D(WX7247), .SI(WX7246), .SE(n4128), .CLK(n4645), 
        .Q(WX7248) );
  SDFFX1 DFF_1062_Q_reg ( .D(WX7249), .SI(WX7248), .SE(n4145), .CLK(n4636), 
        .Q(WX7250), .QN(n3172) );
  SDFFX1 DFF_1063_Q_reg ( .D(WX7251), .SI(WX7250), .SE(n4145), .CLK(n4636), 
        .Q(WX7252) );
  SDFFX1 DFF_1064_Q_reg ( .D(WX7253), .SI(WX7252), .SE(n4145), .CLK(n4636), 
        .Q(test_so61) );
  SDFFX1 DFF_1065_Q_reg ( .D(WX7255), .SI(test_si62), .SE(n4144), .CLK(n4637), 
        .Q(WX7256) );
  SDFFX1 DFF_1066_Q_reg ( .D(WX7257), .SI(WX7256), .SE(n4144), .CLK(n4637), 
        .Q(WX7258) );
  SDFFX1 DFF_1067_Q_reg ( .D(WX7259), .SI(WX7258), .SE(n4143), .CLK(n4637), 
        .Q(WX7260) );
  SDFFX1 DFF_1068_Q_reg ( .D(WX7261), .SI(WX7260), .SE(n4142), .CLK(n4638), 
        .Q(WX7262) );
  SDFFX1 DFF_1069_Q_reg ( .D(WX7263), .SI(WX7262), .SE(n4142), .CLK(n4638), 
        .Q(WX7264) );
  SDFFX1 DFF_1070_Q_reg ( .D(WX7265), .SI(WX7264), .SE(n4141), .CLK(n4638), 
        .Q(WX7266) );
  SDFFX1 DFF_1071_Q_reg ( .D(WX7267), .SI(WX7266), .SE(n4141), .CLK(n4638), 
        .Q(WX7268) );
  SDFFX1 DFF_1072_Q_reg ( .D(WX7269), .SI(WX7268), .SE(n4140), .CLK(n4639), 
        .Q(WX7270), .QN(n7149) );
  SDFFX1 DFF_1073_Q_reg ( .D(WX7271), .SI(WX7270), .SE(n4139), .CLK(n4639), 
        .Q(WX7272), .QN(n7148) );
  SDFFX1 DFF_1074_Q_reg ( .D(WX7273), .SI(WX7272), .SE(n4139), .CLK(n4639), 
        .Q(WX7274), .QN(n7147) );
  SDFFX1 DFF_1075_Q_reg ( .D(WX7275), .SI(WX7274), .SE(n4138), .CLK(n4640), 
        .Q(WX7276), .QN(n7146) );
  SDFFX1 DFF_1076_Q_reg ( .D(WX7277), .SI(WX7276), .SE(n4137), .CLK(n4640), 
        .Q(WX7278), .QN(n7145) );
  SDFFX1 DFF_1077_Q_reg ( .D(WX7279), .SI(WX7278), .SE(n4137), .CLK(n4640), 
        .Q(WX7280) );
  SDFFX1 DFF_1078_Q_reg ( .D(WX7281), .SI(WX7280), .SE(n4136), .CLK(n4641), 
        .Q(WX7282), .QN(n7144) );
  SDFFX1 DFF_1079_Q_reg ( .D(WX7283), .SI(WX7282), .SE(n4136), .CLK(n4641), 
        .Q(WX7284), .QN(n3339) );
  SDFFX1 DFF_1080_Q_reg ( .D(WX7285), .SI(WX7284), .SE(n4135), .CLK(n4641), 
        .Q(WX7286), .QN(n7143) );
  SDFFX1 DFF_1081_Q_reg ( .D(WX7287), .SI(WX7286), .SE(n4134), .CLK(n4642), 
        .Q(test_so62) );
  SDFFX1 DFF_1082_Q_reg ( .D(WX7289), .SI(test_si63), .SE(n4134), .CLK(n4642), 
        .Q(WX7290), .QN(n7142) );
  SDFFX1 DFF_1083_Q_reg ( .D(WX7291), .SI(WX7290), .SE(n4133), .CLK(n4642), 
        .Q(WX7292), .QN(n3336) );
  SDFFX1 DFF_1084_Q_reg ( .D(WX7293), .SI(WX7292), .SE(n4132), .CLK(n4643), 
        .Q(WX7294), .QN(n7141) );
  SDFFX1 DFF_1085_Q_reg ( .D(WX7295), .SI(WX7294), .SE(n4132), .CLK(n4643), 
        .Q(WX7296), .QN(n7140) );
  SDFFX1 DFF_1086_Q_reg ( .D(WX7297), .SI(WX7296), .SE(n4131), .CLK(n4643), 
        .Q(WX7298), .QN(n7139) );
  SDFFX1 DFF_1087_Q_reg ( .D(WX7299), .SI(WX7298), .SE(n4130), .CLK(n4644), 
        .Q(WX7300), .QN(n7138) );
  SDFFX1 DFF_1088_Q_reg ( .D(WX7301), .SI(WX7300), .SE(n4130), .CLK(n4644), 
        .Q(WX7302), .QN(n3565) );
  SDFFX1 DFF_1089_Q_reg ( .D(WX7303), .SI(WX7302), .SE(n4129), .CLK(n4644), 
        .Q(WX7304), .QN(n3566) );
  SDFFX1 DFF_1090_Q_reg ( .D(WX7305), .SI(WX7304), .SE(n4129), .CLK(n4644), 
        .Q(WX7306), .QN(n3568) );
  SDFFX1 DFF_1091_Q_reg ( .D(WX7307), .SI(WX7306), .SE(n4129), .CLK(n4644), 
        .Q(WX7308), .QN(n3570) );
  SDFFX1 DFF_1092_Q_reg ( .D(WX7309), .SI(WX7308), .SE(n4128), .CLK(n4645), 
        .Q(WX7310), .QN(n3572) );
  SDFFX1 DFF_1093_Q_reg ( .D(WX7311), .SI(WX7310), .SE(n4128), .CLK(n4645), 
        .Q(WX7312), .QN(n3574) );
  SDFFX1 DFF_1094_Q_reg ( .D(WX7313), .SI(WX7312), .SE(n4128), .CLK(n4645), 
        .Q(WX7314), .QN(n3576) );
  SDFFX1 DFF_1095_Q_reg ( .D(WX7315), .SI(WX7314), .SE(n4128), .CLK(n4645), 
        .Q(WX7316), .QN(n3578) );
  SDFFX1 DFF_1096_Q_reg ( .D(WX7317), .SI(WX7316), .SE(n4128), .CLK(n4645), 
        .Q(WX7318), .QN(n3580) );
  SDFFX1 DFF_1097_Q_reg ( .D(WX7319), .SI(WX7318), .SE(n4127), .CLK(n4645), 
        .Q(WX7320), .QN(n3582) );
  SDFFX1 DFF_1098_Q_reg ( .D(WX7321), .SI(WX7320), .SE(n4127), .CLK(n4645), 
        .Q(test_so63) );
  SDFFX1 DFF_1099_Q_reg ( .D(WX7323), .SI(test_si64), .SE(n4143), .CLK(n4637), 
        .Q(WX7324), .QN(n3584) );
  SDFFX1 DFF_1100_Q_reg ( .D(WX7325), .SI(WX7324), .SE(n4142), .CLK(n4638), 
        .Q(WX7326), .QN(n3586) );
  SDFFX1 DFF_1101_Q_reg ( .D(WX7327), .SI(WX7326), .SE(n4142), .CLK(n4638), 
        .Q(WX7328), .QN(n3588) );
  SDFFX1 DFF_1102_Q_reg ( .D(WX7329), .SI(WX7328), .SE(n4141), .CLK(n4638), 
        .Q(WX7330), .QN(n3590) );
  SDFFX1 DFF_1103_Q_reg ( .D(WX7331), .SI(WX7330), .SE(n4141), .CLK(n4638), 
        .Q(WX7332), .QN(n3421) );
  SDFFX1 DFF_1104_Q_reg ( .D(WX7333), .SI(WX7332), .SE(n4140), .CLK(n4639), 
        .Q(WX7334), .QN(n3592) );
  SDFFX1 DFF_1105_Q_reg ( .D(WX7335), .SI(WX7334), .SE(n4139), .CLK(n4639), 
        .Q(WX7336), .QN(n3594) );
  SDFFX1 DFF_1106_Q_reg ( .D(WX7337), .SI(WX7336), .SE(n4139), .CLK(n4639), 
        .Q(WX7338), .QN(n3596) );
  SDFFX1 DFF_1107_Q_reg ( .D(WX7339), .SI(WX7338), .SE(n4138), .CLK(n4640), 
        .Q(WX7340), .QN(n3598) );
  SDFFX1 DFF_1108_Q_reg ( .D(WX7341), .SI(WX7340), .SE(n4137), .CLK(n4640), 
        .Q(WX7342), .QN(n3422) );
  SDFFX1 DFF_1109_Q_reg ( .D(WX7343), .SI(WX7342), .SE(n4137), .CLK(n4640), 
        .Q(WX7344), .QN(n3600) );
  SDFFX1 DFF_1110_Q_reg ( .D(WX7345), .SI(WX7344), .SE(n4136), .CLK(n4641), 
        .Q(WX7346), .QN(n3602) );
  SDFFX1 DFF_1111_Q_reg ( .D(WX7347), .SI(WX7346), .SE(n4136), .CLK(n4641), 
        .Q(WX7348), .QN(n3604) );
  SDFFX1 DFF_1112_Q_reg ( .D(WX7349), .SI(WX7348), .SE(n4135), .CLK(n4641), 
        .Q(WX7350), .QN(n3606) );
  SDFFX1 DFF_1113_Q_reg ( .D(WX7351), .SI(WX7350), .SE(n4134), .CLK(n4642), 
        .Q(WX7352), .QN(n3608) );
  SDFFX1 DFF_1114_Q_reg ( .D(WX7353), .SI(WX7352), .SE(n4133), .CLK(n4642), 
        .Q(WX7354), .QN(n3610) );
  SDFFX1 DFF_1115_Q_reg ( .D(WX7355), .SI(WX7354), .SE(n4133), .CLK(n4642), 
        .Q(test_so64) );
  SDFFX1 DFF_1116_Q_reg ( .D(WX7357), .SI(test_si65), .SE(n4132), .CLK(n4643), 
        .Q(WX7358), .QN(n3612) );
  SDFFX1 DFF_1117_Q_reg ( .D(WX7359), .SI(WX7358), .SE(n4131), .CLK(n4643), 
        .Q(WX7360), .QN(n3614) );
  SDFFX1 DFF_1118_Q_reg ( .D(WX7361), .SI(WX7360), .SE(n4131), .CLK(n4643), 
        .Q(WX7362), .QN(n3616) );
  SDFFX1 DFF_1119_Q_reg ( .D(WX7363), .SI(WX7362), .SE(n4130), .CLK(n4644), 
        .Q(WX7364), .QN(n3436) );
  SDFFX1 DFF_1120_Q_reg ( .D(WX7729), .SI(WX7364), .SE(n4031), .CLK(n4693), 
        .Q(CRC_OUT_4_0), .QN(DFF_1120_n1) );
  SDFFX1 DFF_1121_Q_reg ( .D(WX7731), .SI(CRC_OUT_4_0), .SE(n4031), .CLK(n4693), .Q(CRC_OUT_4_1), .QN(DFF_1121_n1) );
  SDFFX1 DFF_1122_Q_reg ( .D(WX7733), .SI(CRC_OUT_4_1), .SE(n4030), .CLK(n4694), .Q(CRC_OUT_4_2), .QN(DFF_1122_n1) );
  SDFFX1 DFF_1123_Q_reg ( .D(WX7735), .SI(CRC_OUT_4_2), .SE(n4030), .CLK(n4694), .Q(CRC_OUT_4_3), .QN(DFF_1123_n1) );
  SDFFX1 DFF_1124_Q_reg ( .D(WX7737), .SI(CRC_OUT_4_3), .SE(n4030), .CLK(n4694), .Q(CRC_OUT_4_4), .QN(DFF_1124_n1) );
  SDFFX1 DFF_1125_Q_reg ( .D(WX7739), .SI(CRC_OUT_4_4), .SE(n4030), .CLK(n4694), .Q(CRC_OUT_4_5), .QN(DFF_1125_n1) );
  SDFFX1 DFF_1126_Q_reg ( .D(WX7741), .SI(CRC_OUT_4_5), .SE(n4030), .CLK(n4694), .Q(CRC_OUT_4_6), .QN(DFF_1126_n1) );
  SDFFX1 DFF_1127_Q_reg ( .D(WX7743), .SI(CRC_OUT_4_6), .SE(n4030), .CLK(n4694), .Q(CRC_OUT_4_7), .QN(DFF_1127_n1) );
  SDFFX1 DFF_1128_Q_reg ( .D(WX7745), .SI(CRC_OUT_4_7), .SE(n4029), .CLK(n4694), .Q(CRC_OUT_4_8), .QN(DFF_1128_n1) );
  SDFFX1 DFF_1129_Q_reg ( .D(WX7747), .SI(CRC_OUT_4_8), .SE(n4029), .CLK(n4694), .Q(CRC_OUT_4_9), .QN(DFF_1129_n1) );
  SDFFX1 DFF_1130_Q_reg ( .D(WX7749), .SI(CRC_OUT_4_9), .SE(n4029), .CLK(n4694), .Q(CRC_OUT_4_10) );
  SDFFX1 DFF_1131_Q_reg ( .D(WX7751), .SI(CRC_OUT_4_10), .SE(n4029), .CLK(
        n4694), .Q(CRC_OUT_4_11), .QN(DFF_1131_n1) );
  SDFFX1 DFF_1132_Q_reg ( .D(WX7753), .SI(CRC_OUT_4_11), .SE(n4029), .CLK(
        n4694), .Q(test_so65) );
  SDFFX1 DFF_1133_Q_reg ( .D(WX7755), .SI(test_si66), .SE(n4029), .CLK(n4694), 
        .Q(CRC_OUT_4_13), .QN(DFF_1133_n1) );
  SDFFX1 DFF_1134_Q_reg ( .D(WX7757), .SI(CRC_OUT_4_13), .SE(n4028), .CLK(
        n4695), .Q(CRC_OUT_4_14), .QN(DFF_1134_n1) );
  SDFFX1 DFF_1135_Q_reg ( .D(WX7759), .SI(CRC_OUT_4_14), .SE(n4028), .CLK(
        n4695), .Q(CRC_OUT_4_15) );
  SDFFX1 DFF_1136_Q_reg ( .D(WX7761), .SI(CRC_OUT_4_15), .SE(n4028), .CLK(
        n4695), .Q(CRC_OUT_4_16), .QN(DFF_1136_n1) );
  SDFFX1 DFF_1137_Q_reg ( .D(WX7763), .SI(CRC_OUT_4_16), .SE(n4028), .CLK(
        n4695), .Q(CRC_OUT_4_17), .QN(DFF_1137_n1) );
  SDFFX1 DFF_1138_Q_reg ( .D(WX7765), .SI(CRC_OUT_4_17), .SE(n4028), .CLK(
        n4695), .Q(CRC_OUT_4_18), .QN(DFF_1138_n1) );
  SDFFX1 DFF_1139_Q_reg ( .D(WX7767), .SI(CRC_OUT_4_18), .SE(n4028), .CLK(
        n4695), .Q(CRC_OUT_4_19), .QN(DFF_1139_n1) );
  SDFFX1 DFF_1140_Q_reg ( .D(WX7769), .SI(CRC_OUT_4_19), .SE(n4027), .CLK(
        n4695), .Q(CRC_OUT_4_20) );
  SDFFX1 DFF_1141_Q_reg ( .D(WX7771), .SI(CRC_OUT_4_20), .SE(n4027), .CLK(
        n4695), .Q(CRC_OUT_4_21), .QN(DFF_1141_n1) );
  SDFFX1 DFF_1142_Q_reg ( .D(WX7773), .SI(CRC_OUT_4_21), .SE(n4027), .CLK(
        n4695), .Q(CRC_OUT_4_22), .QN(DFF_1142_n1) );
  SDFFX1 DFF_1143_Q_reg ( .D(WX7775), .SI(CRC_OUT_4_22), .SE(n4027), .CLK(
        n4695), .Q(CRC_OUT_4_23), .QN(DFF_1143_n1) );
  SDFFX1 DFF_1144_Q_reg ( .D(WX7777), .SI(CRC_OUT_4_23), .SE(n4027), .CLK(
        n4695), .Q(CRC_OUT_4_24), .QN(DFF_1144_n1) );
  SDFFX1 DFF_1145_Q_reg ( .D(WX7779), .SI(CRC_OUT_4_24), .SE(n4027), .CLK(
        n4695), .Q(CRC_OUT_4_25), .QN(DFF_1145_n1) );
  SDFFX1 DFF_1146_Q_reg ( .D(WX7781), .SI(CRC_OUT_4_25), .SE(n4127), .CLK(
        n4645), .Q(CRC_OUT_4_26), .QN(DFF_1146_n1) );
  SDFFX1 DFF_1147_Q_reg ( .D(WX7783), .SI(CRC_OUT_4_26), .SE(n4127), .CLK(
        n4645), .Q(CRC_OUT_4_27), .QN(DFF_1147_n1) );
  SDFFX1 DFF_1148_Q_reg ( .D(WX7785), .SI(CRC_OUT_4_27), .SE(n4127), .CLK(
        n4645), .Q(CRC_OUT_4_28), .QN(DFF_1148_n1) );
  SDFFX1 DFF_1149_Q_reg ( .D(WX7787), .SI(CRC_OUT_4_28), .SE(n4127), .CLK(
        n4645), .Q(test_so66) );
  SDFFX1 DFF_1150_Q_reg ( .D(WX7789), .SI(test_si67), .SE(n4126), .CLK(n4646), 
        .Q(CRC_OUT_4_30), .QN(DFF_1150_n1) );
  SDFFX1 DFF_1151_Q_reg ( .D(WX7791), .SI(CRC_OUT_4_30), .SE(n4126), .CLK(
        n4646), .Q(CRC_OUT_4_31), .QN(DFF_1151_n1) );
  SDFFX1 DFF_1152_Q_reg ( .D(n424), .SI(CRC_OUT_4_31), .SE(n4126), .CLK(n4646), 
        .Q(WX8243) );
  SDFFX1 DFF_1153_Q_reg ( .D(n425), .SI(WX8243), .SE(n4126), .CLK(n4646), .Q(
        n8411) );
  SDFFX1 DFF_1154_Q_reg ( .D(n426), .SI(n8411), .SE(n4126), .CLK(n4646), .Q(
        n8410) );
  SDFFX1 DFF_1155_Q_reg ( .D(n427), .SI(n8410), .SE(n4126), .CLK(n4646), .Q(
        n8409) );
  SDFFX1 DFF_1156_Q_reg ( .D(n428), .SI(n8409), .SE(n4125), .CLK(n4646), .Q(
        n8408) );
  SDFFX1 DFF_1157_Q_reg ( .D(n429), .SI(n8408), .SE(n4125), .CLK(n4646), .Q(
        n8407) );
  SDFFX1 DFF_1158_Q_reg ( .D(n430), .SI(n8407), .SE(n4125), .CLK(n4646), .Q(
        n8406) );
  SDFFX1 DFF_1159_Q_reg ( .D(n431), .SI(n8406), .SE(n4125), .CLK(n4646), .Q(
        n8405) );
  SDFFX1 DFF_1160_Q_reg ( .D(n432), .SI(n8405), .SE(n4125), .CLK(n4646), .Q(
        n8404) );
  SDFFX1 DFF_1161_Q_reg ( .D(n433), .SI(n8404), .SE(n4125), .CLK(n4646), .Q(
        n8403) );
  SDFFX1 DFF_1162_Q_reg ( .D(n434), .SI(n8403), .SE(n4124), .CLK(n4647), .Q(
        n8402) );
  SDFFX1 DFF_1163_Q_reg ( .D(n435), .SI(n8402), .SE(n4124), .CLK(n4647), .Q(
        n8401) );
  SDFFX1 DFF_1164_Q_reg ( .D(WX8266), .SI(n8401), .SE(n4219), .CLK(n4599), .Q(
        n8400) );
  SDFFX1 DFF_1165_Q_reg ( .D(n437), .SI(n8400), .SE(n4219), .CLK(n4599), .Q(
        n8399), .QN(n3870) );
  SDFFX1 DFF_1166_Q_reg ( .D(n438), .SI(n8399), .SE(n4218), .CLK(n4600), .Q(
        test_so67) );
  SDFFX1 DFF_1167_Q_reg ( .D(n439), .SI(test_si68), .SE(n4121), .CLK(n4648), 
        .Q(n8396) );
  SDFFX1 DFF_1168_Q_reg ( .D(n440), .SI(n8396), .SE(n4122), .CLK(n4648), .Q(
        n8395) );
  SDFFX1 DFF_1169_Q_reg ( .D(n441), .SI(n8395), .SE(n4122), .CLK(n4648), .Q(
        n8394) );
  SDFFX1 DFF_1170_Q_reg ( .D(n442), .SI(n8394), .SE(n4122), .CLK(n4648), .Q(
        n8393) );
  SDFFX1 DFF_1171_Q_reg ( .D(n443), .SI(n8393), .SE(n4122), .CLK(n4648), .Q(
        n8392) );
  SDFFX1 DFF_1172_Q_reg ( .D(n444), .SI(n8392), .SE(n4122), .CLK(n4648), .Q(
        n8391) );
  SDFFX1 DFF_1173_Q_reg ( .D(n445), .SI(n8391), .SE(n4122), .CLK(n4648), .Q(
        n8390) );
  SDFFX1 DFF_1174_Q_reg ( .D(n446), .SI(n8390), .SE(n4123), .CLK(n4647), .Q(
        n8389) );
  SDFFX1 DFF_1175_Q_reg ( .D(n447), .SI(n8389), .SE(n4123), .CLK(n4647), .Q(
        n8388) );
  SDFFX1 DFF_1176_Q_reg ( .D(n448), .SI(n8388), .SE(n4123), .CLK(n4647), .Q(
        n8387) );
  SDFFX1 DFF_1177_Q_reg ( .D(n449), .SI(n8387), .SE(n4123), .CLK(n4647), .Q(
        n8386) );
  SDFFX1 DFF_1178_Q_reg ( .D(n450), .SI(n8386), .SE(n4123), .CLK(n4647), .Q(
        n8385) );
  SDFFX1 DFF_1179_Q_reg ( .D(n451), .SI(n8385), .SE(n4123), .CLK(n4647), .Q(
        n8384) );
  SDFFX1 DFF_1180_Q_reg ( .D(n452), .SI(n8384), .SE(n4124), .CLK(n4647), .Q(
        n8383) );
  SDFFX1 DFF_1181_Q_reg ( .D(n453), .SI(n8383), .SE(n4124), .CLK(n4647), .Q(
        n8382) );
  SDFFX1 DFF_1182_Q_reg ( .D(n454), .SI(n8382), .SE(n4124), .CLK(n4647), .Q(
        n8381) );
  SDFFX1 DFF_1183_Q_reg ( .D(WX8304), .SI(n8381), .SE(n4124), .CLK(n4647), .Q(
        test_so68) );
  SDFFX1 DFF_1184_Q_reg ( .D(WX8402), .SI(test_si69), .SE(n4121), .CLK(n4648), 
        .Q(n8378), .QN(n7137) );
  SDFFX1 DFF_1185_Q_reg ( .D(WX8404), .SI(n8378), .SE(n4121), .CLK(n4648), .Q(
        n8377), .QN(n7136) );
  SDFFX1 DFF_1186_Q_reg ( .D(WX8406), .SI(n8377), .SE(n4121), .CLK(n4648), .Q(
        n8376), .QN(n7135) );
  SDFFX1 DFF_1187_Q_reg ( .D(WX8408), .SI(n8376), .SE(n4120), .CLK(n4649), .Q(
        n8375), .QN(n7134) );
  SDFFX1 DFF_1188_Q_reg ( .D(WX8410), .SI(n8375), .SE(n4120), .CLK(n4649), .Q(
        n8374), .QN(n7133) );
  SDFFX1 DFF_1189_Q_reg ( .D(WX8412), .SI(n8374), .SE(n4119), .CLK(n4649), .Q(
        n8373), .QN(n7132) );
  SDFFX1 DFF_1190_Q_reg ( .D(WX8414), .SI(n8373), .SE(n4119), .CLK(n4649), .Q(
        n8372), .QN(n7131) );
  SDFFX1 DFF_1191_Q_reg ( .D(WX8416), .SI(n8372), .SE(n4118), .CLK(n4650), .Q(
        n8371), .QN(n7130) );
  SDFFX1 DFF_1192_Q_reg ( .D(WX8418), .SI(n8371), .SE(n4118), .CLK(n4650), .Q(
        n8370), .QN(n7129) );
  SDFFX1 DFF_1193_Q_reg ( .D(WX8420), .SI(n8370), .SE(n4116), .CLK(n4651), .Q(
        n8369), .QN(n7128) );
  SDFFX1 DFF_1194_Q_reg ( .D(WX8422), .SI(n8369), .SE(n4116), .CLK(n4651), .Q(
        n8368), .QN(n7127) );
  SDFFX1 DFF_1195_Q_reg ( .D(WX8424), .SI(n8368), .SE(n4115), .CLK(n4651), .Q(
        n8367), .QN(n7126) );
  SDFFX1 DFF_1196_Q_reg ( .D(WX8426), .SI(n8367), .SE(n4115), .CLK(n4651), .Q(
        n8366), .QN(n7125) );
  SDFFX1 DFF_1197_Q_reg ( .D(WX8428), .SI(n8366), .SE(n4031), .CLK(n4693), .Q(
        n8365), .QN(n7124) );
  SDFFX1 DFF_1198_Q_reg ( .D(WX8430), .SI(n8365), .SE(n4218), .CLK(n4600), .Q(
        n8364), .QN(n7123) );
  SDFFX1 DFF_1199_Q_reg ( .D(WX8432), .SI(n8364), .SE(n4113), .CLK(n4652), .Q(
        n8363), .QN(n7122) );
  SDFFX1 DFF_1200_Q_reg ( .D(WX8434), .SI(n8363), .SE(n4113), .CLK(n4652), .Q(
        test_so69) );
  SDFFX1 DFF_1201_Q_reg ( .D(WX8436), .SI(test_si70), .SE(n4031), .CLK(n4693), 
        .Q(WX8437), .QN(n3331) );
  SDFFX1 DFF_1202_Q_reg ( .D(WX8438), .SI(WX8437), .SE(n4111), .CLK(n4653), 
        .Q(WX8439) );
  SDFFX1 DFF_1203_Q_reg ( .D(WX8440), .SI(WX8439), .SE(n4111), .CLK(n4653), 
        .Q(WX8441), .QN(n3329) );
  SDFFX1 DFF_1204_Q_reg ( .D(WX8442), .SI(WX8441), .SE(n4110), .CLK(n4654), 
        .Q(WX8443) );
  SDFFX1 DFF_1205_Q_reg ( .D(WX8444), .SI(WX8443), .SE(n4109), .CLK(n4654), 
        .Q(WX8445), .QN(n3328) );
  SDFFX1 DFF_1206_Q_reg ( .D(WX8446), .SI(WX8445), .SE(n4109), .CLK(n4654), 
        .Q(WX8447) );
  SDFFX1 DFF_1207_Q_reg ( .D(WX8448), .SI(WX8447), .SE(n4108), .CLK(n4655), 
        .Q(WX8449), .QN(n3326) );
  SDFFX1 DFF_1208_Q_reg ( .D(WX8450), .SI(WX8449), .SE(n4107), .CLK(n4655), 
        .Q(WX8451), .QN(n3325) );
  SDFFX1 DFF_1209_Q_reg ( .D(WX8452), .SI(WX8451), .SE(n4107), .CLK(n4655), 
        .Q(WX8453), .QN(n3324) );
  SDFFX1 DFF_1210_Q_reg ( .D(WX8454), .SI(WX8453), .SE(n4106), .CLK(n4656), 
        .Q(WX8455), .QN(n3323) );
  SDFFX1 DFF_1211_Q_reg ( .D(WX8456), .SI(WX8455), .SE(n4105), .CLK(n4656), 
        .Q(WX8457), .QN(n3322) );
  SDFFX1 DFF_1212_Q_reg ( .D(WX8458), .SI(WX8457), .SE(n4105), .CLK(n4656), 
        .Q(WX8459), .QN(n3321) );
  SDFFX1 DFF_1213_Q_reg ( .D(WX8460), .SI(WX8459), .SE(n4104), .CLK(n4657), 
        .Q(WX8461), .QN(n3320) );
  SDFFX1 DFF_1214_Q_reg ( .D(WX8462), .SI(WX8461), .SE(n4103), .CLK(n4657), 
        .Q(WX8463), .QN(n3319) );
  SDFFX1 DFF_1215_Q_reg ( .D(WX8464), .SI(WX8463), .SE(n4103), .CLK(n4657), 
        .Q(WX8465), .QN(n3318) );
  SDFFX1 DFF_1216_Q_reg ( .D(n455), .SI(WX8465), .SE(n4121), .CLK(n4648), .Q(
        WX8467), .QN(n3064) );
  SDFFX1 DFF_1217_Q_reg ( .D(n456), .SI(WX8467), .SE(n4121), .CLK(n4648), .Q(
        test_so70) );
  SDFFX1 DFF_1218_Q_reg ( .D(n457), .SI(test_si71), .SE(n4120), .CLK(n4649), 
        .Q(WX8471), .QN(n3153) );
  SDFFX1 DFF_1219_Q_reg ( .D(n458), .SI(WX8471), .SE(n4120), .CLK(n4649), .Q(
        WX8473), .QN(n3152) );
  SDFFX1 DFF_1220_Q_reg ( .D(n459), .SI(WX8473), .SE(n4120), .CLK(n4649), .Q(
        WX8475), .QN(n3150) );
  SDFFX1 DFF_1221_Q_reg ( .D(n460), .SI(WX8475), .SE(n4119), .CLK(n4649), .Q(
        WX8477), .QN(n3149) );
  SDFFX1 DFF_1222_Q_reg ( .D(n461), .SI(WX8477), .SE(n4119), .CLK(n4649), .Q(
        WX8479), .QN(n3147) );
  SDFFX1 DFF_1223_Q_reg ( .D(n462), .SI(WX8479), .SE(n4118), .CLK(n4650), .Q(
        WX8481), .QN(n3145) );
  SDFFX1 DFF_1224_Q_reg ( .D(n463), .SI(WX8481), .SE(n4117), .CLK(n4650), .Q(
        WX8483), .QN(n3143) );
  SDFFX1 DFF_1225_Q_reg ( .D(n464), .SI(WX8483), .SE(n4117), .CLK(n4650), .Q(
        WX8485), .QN(n3141) );
  SDFFX1 DFF_1226_Q_reg ( .D(n465), .SI(WX8485), .SE(n4116), .CLK(n4651), .Q(
        WX8487), .QN(n3139) );
  SDFFX1 DFF_1227_Q_reg ( .D(n466), .SI(WX8487), .SE(n4116), .CLK(n4651), .Q(
        WX8489), .QN(n3137) );
  SDFFX1 DFF_1228_Q_reg ( .D(n467), .SI(WX8489), .SE(n4115), .CLK(n4651), .Q(
        WX8491), .QN(n3135) );
  SDFFX1 DFF_1229_Q_reg ( .D(n468), .SI(WX8491), .SE(n4114), .CLK(n4652), .Q(
        WX8493), .QN(n3133) );
  SDFFX1 DFF_1230_Q_reg ( .D(n469), .SI(WX8493), .SE(n4114), .CLK(n4652), .Q(
        WX8495), .QN(n3131) );
  SDFFX1 DFF_1231_Q_reg ( .D(n470), .SI(WX8495), .SE(n4113), .CLK(n4652), .Q(
        WX8497), .QN(n3129) );
  SDFFX1 DFF_1232_Q_reg ( .D(WX8498), .SI(WX8497), .SE(n4112), .CLK(n4653), 
        .Q(WX8499), .QN(n3625) );
  SDFFX1 DFF_1233_Q_reg ( .D(WX8500), .SI(WX8499), .SE(n4112), .CLK(n4653), 
        .Q(WX8501) );
  SDFFX1 DFF_1234_Q_reg ( .D(WX8502), .SI(WX8501), .SE(n4111), .CLK(n4653), 
        .Q(test_so71) );
  SDFFX1 DFF_1235_Q_reg ( .D(WX8504), .SI(test_si72), .SE(n4111), .CLK(n4653), 
        .Q(WX8505) );
  SDFFX1 DFF_1236_Q_reg ( .D(WX8506), .SI(WX8505), .SE(n4110), .CLK(n4654), 
        .Q(WX8507), .QN(n3617) );
  SDFFX1 DFF_1237_Q_reg ( .D(WX8508), .SI(WX8507), .SE(n4109), .CLK(n4654), 
        .Q(WX8509) );
  SDFFX1 DFF_1238_Q_reg ( .D(WX8510), .SI(WX8509), .SE(n4109), .CLK(n4654), 
        .Q(WX8511), .QN(n3613) );
  SDFFX1 DFF_1239_Q_reg ( .D(WX8512), .SI(WX8511), .SE(n4108), .CLK(n4655), 
        .Q(WX8513) );
  SDFFX1 DFF_1240_Q_reg ( .D(WX8514), .SI(WX8513), .SE(n4107), .CLK(n4655), 
        .Q(WX8515) );
  SDFFX1 DFF_1241_Q_reg ( .D(WX8516), .SI(WX8515), .SE(n4107), .CLK(n4655), 
        .Q(WX8517) );
  SDFFX1 DFF_1242_Q_reg ( .D(WX8518), .SI(WX8517), .SE(n4106), .CLK(n4656), 
        .Q(WX8519) );
  SDFFX1 DFF_1243_Q_reg ( .D(WX8520), .SI(WX8519), .SE(n4105), .CLK(n4656), 
        .Q(WX8521) );
  SDFFX1 DFF_1244_Q_reg ( .D(WX8522), .SI(WX8521), .SE(n4105), .CLK(n4656), 
        .Q(WX8523) );
  SDFFX1 DFF_1245_Q_reg ( .D(WX8524), .SI(WX8523), .SE(n4104), .CLK(n4657), 
        .Q(WX8525) );
  SDFFX1 DFF_1246_Q_reg ( .D(WX8526), .SI(WX8525), .SE(n4103), .CLK(n4657), 
        .Q(WX8527) );
  SDFFX1 DFF_1247_Q_reg ( .D(WX8528), .SI(WX8527), .SE(n4103), .CLK(n4657), 
        .Q(WX8529) );
  SDFFX1 DFF_1248_Q_reg ( .D(WX8530), .SI(WX8529), .SE(n4102), .CLK(n4658), 
        .Q(WX8531) );
  SDFFX1 DFF_1249_Q_reg ( .D(WX8532), .SI(WX8531), .SE(n4102), .CLK(n4658), 
        .Q(WX8533), .QN(n3155) );
  SDFFX1 DFF_1250_Q_reg ( .D(WX8534), .SI(WX8533), .SE(n4101), .CLK(n4658), 
        .Q(WX8535) );
  SDFFX1 DFF_1251_Q_reg ( .D(WX8536), .SI(WX8535), .SE(n4101), .CLK(n4658), 
        .Q(test_so72) );
  SDFFX1 DFF_1252_Q_reg ( .D(WX8538), .SI(test_si73), .SE(n4120), .CLK(n4649), 
        .Q(WX8539) );
  SDFFX1 DFF_1253_Q_reg ( .D(WX8540), .SI(WX8539), .SE(n4119), .CLK(n4649), 
        .Q(WX8541) );
  SDFFX1 DFF_1254_Q_reg ( .D(WX8542), .SI(WX8541), .SE(n4119), .CLK(n4649), 
        .Q(WX8543) );
  SDFFX1 DFF_1255_Q_reg ( .D(WX8544), .SI(WX8543), .SE(n4118), .CLK(n4650), 
        .Q(WX8545) );
  SDFFX1 DFF_1256_Q_reg ( .D(WX8546), .SI(WX8545), .SE(n4117), .CLK(n4650), 
        .Q(WX8547) );
  SDFFX1 DFF_1257_Q_reg ( .D(WX8548), .SI(WX8547), .SE(n4117), .CLK(n4650), 
        .Q(WX8549) );
  SDFFX1 DFF_1258_Q_reg ( .D(WX8550), .SI(WX8549), .SE(n4116), .CLK(n4651), 
        .Q(WX8551) );
  SDFFX1 DFF_1259_Q_reg ( .D(WX8552), .SI(WX8551), .SE(n4115), .CLK(n4651), 
        .Q(WX8553) );
  SDFFX1 DFF_1260_Q_reg ( .D(WX8554), .SI(WX8553), .SE(n4115), .CLK(n4651), 
        .Q(WX8555) );
  SDFFX1 DFF_1261_Q_reg ( .D(WX8556), .SI(WX8555), .SE(n4114), .CLK(n4652), 
        .Q(WX8557) );
  SDFFX1 DFF_1262_Q_reg ( .D(WX8558), .SI(WX8557), .SE(n4114), .CLK(n4652), 
        .Q(WX8559) );
  SDFFX1 DFF_1263_Q_reg ( .D(WX8560), .SI(WX8559), .SE(n4113), .CLK(n4652), 
        .Q(WX8561) );
  SDFFX1 DFF_1264_Q_reg ( .D(WX8562), .SI(WX8561), .SE(n4112), .CLK(n4653), 
        .Q(WX8563) );
  SDFFX1 DFF_1265_Q_reg ( .D(WX8564), .SI(WX8563), .SE(n4112), .CLK(n4653), 
        .Q(WX8565), .QN(n7121) );
  SDFFX1 DFF_1266_Q_reg ( .D(WX8566), .SI(WX8565), .SE(n4111), .CLK(n4653), 
        .Q(WX8567), .QN(n3330) );
  SDFFX1 DFF_1267_Q_reg ( .D(WX8568), .SI(WX8567), .SE(n4110), .CLK(n4654), 
        .Q(WX8569), .QN(n7120) );
  SDFFX1 DFF_1268_Q_reg ( .D(WX8570), .SI(WX8569), .SE(n4110), .CLK(n4654), 
        .Q(test_so73) );
  SDFFX1 DFF_1269_Q_reg ( .D(WX8572), .SI(test_si74), .SE(n4109), .CLK(n4654), 
        .Q(WX8573), .QN(n7119) );
  SDFFX1 DFF_1270_Q_reg ( .D(WX8574), .SI(WX8573), .SE(n4108), .CLK(n4655), 
        .Q(WX8575), .QN(n3327) );
  SDFFX1 DFF_1271_Q_reg ( .D(WX8576), .SI(WX8575), .SE(n4108), .CLK(n4655), 
        .Q(WX8577), .QN(n7118) );
  SDFFX1 DFF_1272_Q_reg ( .D(WX8578), .SI(WX8577), .SE(n4107), .CLK(n4655), 
        .Q(WX8579), .QN(n7117) );
  SDFFX1 DFF_1273_Q_reg ( .D(WX8580), .SI(WX8579), .SE(n4106), .CLK(n4656), 
        .Q(WX8581), .QN(n7116) );
  SDFFX1 DFF_1274_Q_reg ( .D(WX8582), .SI(WX8581), .SE(n4106), .CLK(n4656), 
        .Q(WX8583), .QN(n7115) );
  SDFFX1 DFF_1275_Q_reg ( .D(WX8584), .SI(WX8583), .SE(n4105), .CLK(n4656), 
        .Q(WX8585), .QN(n7114) );
  SDFFX1 DFF_1276_Q_reg ( .D(WX8586), .SI(WX8585), .SE(n4104), .CLK(n4657), 
        .Q(WX8587), .QN(n7113) );
  SDFFX1 DFF_1277_Q_reg ( .D(WX8588), .SI(WX8587), .SE(n4104), .CLK(n4657), 
        .Q(WX8589), .QN(n7112) );
  SDFFX1 DFF_1278_Q_reg ( .D(WX8590), .SI(WX8589), .SE(n4103), .CLK(n4657), 
        .Q(WX8591), .QN(n7111) );
  SDFFX1 DFF_1279_Q_reg ( .D(WX8592), .SI(WX8591), .SE(n4102), .CLK(n4658), 
        .Q(WX8593), .QN(n7110) );
  SDFFX1 DFF_1280_Q_reg ( .D(WX8594), .SI(WX8593), .SE(n4102), .CLK(n4658), 
        .Q(WX8595), .QN(n3518) );
  SDFFX1 DFF_1281_Q_reg ( .D(WX8596), .SI(WX8595), .SE(n4102), .CLK(n4658), 
        .Q(WX8597), .QN(n3520) );
  SDFFX1 DFF_1282_Q_reg ( .D(WX8598), .SI(WX8597), .SE(n4101), .CLK(n4658), 
        .Q(WX8599), .QN(n3522) );
  SDFFX1 DFF_1283_Q_reg ( .D(WX8600), .SI(WX8599), .SE(n4101), .CLK(n4658), 
        .Q(WX8601), .QN(n3523) );
  SDFFX1 DFF_1284_Q_reg ( .D(WX8602), .SI(WX8601), .SE(n4101), .CLK(n4658), 
        .Q(WX8603), .QN(n3524) );
  SDFFX1 DFF_1285_Q_reg ( .D(WX8604), .SI(WX8603), .SE(n4101), .CLK(n4658), 
        .Q(test_so74) );
  SDFFX1 DFF_1286_Q_reg ( .D(WX8606), .SI(test_si75), .SE(n4118), .CLK(n4650), 
        .Q(WX8607), .QN(n3526) );
  SDFFX1 DFF_1287_Q_reg ( .D(WX8608), .SI(WX8607), .SE(n4118), .CLK(n4650), 
        .Q(WX8609), .QN(n3528) );
  SDFFX1 DFF_1288_Q_reg ( .D(WX8610), .SI(WX8609), .SE(n4117), .CLK(n4650), 
        .Q(WX8611), .QN(n3530) );
  SDFFX1 DFF_1289_Q_reg ( .D(WX8612), .SI(WX8611), .SE(n4117), .CLK(n4650), 
        .Q(WX8613), .QN(n3532) );
  SDFFX1 DFF_1290_Q_reg ( .D(WX8614), .SI(WX8613), .SE(n4116), .CLK(n4651), 
        .Q(WX8615), .QN(n3534) );
  SDFFX1 DFF_1291_Q_reg ( .D(WX8616), .SI(WX8615), .SE(n4115), .CLK(n4651), 
        .Q(WX8617), .QN(n3536) );
  SDFFX1 DFF_1292_Q_reg ( .D(WX8618), .SI(WX8617), .SE(n4114), .CLK(n4652), 
        .Q(WX8619), .QN(n3538) );
  SDFFX1 DFF_1293_Q_reg ( .D(WX8620), .SI(WX8619), .SE(n4114), .CLK(n4652), 
        .Q(WX8621), .QN(n3540) );
  SDFFX1 DFF_1294_Q_reg ( .D(WX8622), .SI(WX8621), .SE(n4113), .CLK(n4652), 
        .Q(WX8623), .QN(n3542) );
  SDFFX1 DFF_1295_Q_reg ( .D(WX8624), .SI(WX8623), .SE(n4113), .CLK(n4652), 
        .Q(WX8625), .QN(n3418) );
  SDFFX1 DFF_1296_Q_reg ( .D(WX8626), .SI(WX8625), .SE(n4112), .CLK(n4653), 
        .Q(WX8627), .QN(n3543) );
  SDFFX1 DFF_1297_Q_reg ( .D(WX8628), .SI(WX8627), .SE(n4112), .CLK(n4653), 
        .Q(WX8629), .QN(n3544) );
  SDFFX1 DFF_1298_Q_reg ( .D(WX8630), .SI(WX8629), .SE(n4111), .CLK(n4653), 
        .Q(WX8631), .QN(n3546) );
  SDFFX1 DFF_1299_Q_reg ( .D(WX8632), .SI(WX8631), .SE(n4110), .CLK(n4654), 
        .Q(WX8633), .QN(n3548) );
  SDFFX1 DFF_1300_Q_reg ( .D(WX8634), .SI(WX8633), .SE(n4110), .CLK(n4654), 
        .Q(WX8635), .QN(n3419) );
  SDFFX1 DFF_1301_Q_reg ( .D(WX8636), .SI(WX8635), .SE(n4109), .CLK(n4654), 
        .Q(WX8637), .QN(n3550) );
  SDFFX1 DFF_1302_Q_reg ( .D(WX8638), .SI(WX8637), .SE(n4108), .CLK(n4655), 
        .Q(test_so75) );
  SDFFX1 DFF_1303_Q_reg ( .D(WX8640), .SI(test_si76), .SE(n4108), .CLK(n4655), 
        .Q(WX8641), .QN(n3552) );
  SDFFX1 DFF_1304_Q_reg ( .D(WX8642), .SI(WX8641), .SE(n4107), .CLK(n4655), 
        .Q(WX8643), .QN(n3554) );
  SDFFX1 DFF_1305_Q_reg ( .D(WX8644), .SI(WX8643), .SE(n4106), .CLK(n4656), 
        .Q(WX8645), .QN(n3556) );
  SDFFX1 DFF_1306_Q_reg ( .D(WX8646), .SI(WX8645), .SE(n4106), .CLK(n4656), 
        .Q(WX8647), .QN(n3558) );
  SDFFX1 DFF_1307_Q_reg ( .D(WX8648), .SI(WX8647), .SE(n4105), .CLK(n4656), 
        .Q(WX8649), .QN(n3420) );
  SDFFX1 DFF_1308_Q_reg ( .D(WX8650), .SI(WX8649), .SE(n4104), .CLK(n4657), 
        .Q(WX8651), .QN(n3560) );
  SDFFX1 DFF_1309_Q_reg ( .D(WX8652), .SI(WX8651), .SE(n4104), .CLK(n4657), 
        .Q(WX8653), .QN(n3562) );
  SDFFX1 DFF_1310_Q_reg ( .D(WX8654), .SI(WX8653), .SE(n4103), .CLK(n4657), 
        .Q(WX8655), .QN(n3564) );
  SDFFX1 DFF_1311_Q_reg ( .D(WX8656), .SI(WX8655), .SE(n4102), .CLK(n4658), 
        .Q(WX8657), .QN(n3435) );
  SDFFX1 DFF_1312_Q_reg ( .D(WX9022), .SI(WX8657), .SE(n4036), .CLK(n4691), 
        .Q(CRC_OUT_3_0), .QN(DFF_1312_n1) );
  SDFFX1 DFF_1313_Q_reg ( .D(WX9024), .SI(CRC_OUT_3_0), .SE(n4036), .CLK(n4691), .Q(CRC_OUT_3_1), .QN(DFF_1313_n1) );
  SDFFX1 DFF_1314_Q_reg ( .D(WX9026), .SI(CRC_OUT_3_1), .SE(n4035), .CLK(n4691), .Q(CRC_OUT_3_2), .QN(DFF_1314_n1) );
  SDFFX1 DFF_1315_Q_reg ( .D(WX9028), .SI(CRC_OUT_3_2), .SE(n4035), .CLK(n4691), .Q(CRC_OUT_3_3) );
  SDFFX1 DFF_1316_Q_reg ( .D(WX9030), .SI(CRC_OUT_3_3), .SE(n4035), .CLK(n4691), .Q(CRC_OUT_3_4), .QN(DFF_1316_n1) );
  SDFFX1 DFF_1317_Q_reg ( .D(WX9032), .SI(CRC_OUT_3_4), .SE(n4035), .CLK(n4691), .Q(CRC_OUT_3_5), .QN(DFF_1317_n1) );
  SDFFX1 DFF_1318_Q_reg ( .D(WX9034), .SI(CRC_OUT_3_5), .SE(n4035), .CLK(n4691), .Q(CRC_OUT_3_6), .QN(DFF_1318_n1) );
  SDFFX1 DFF_1319_Q_reg ( .D(WX9036), .SI(CRC_OUT_3_6), .SE(n4035), .CLK(n4691), .Q(test_so76) );
  SDFFX1 DFF_1320_Q_reg ( .D(WX9038), .SI(test_si77), .SE(n4034), .CLK(n4692), 
        .Q(CRC_OUT_3_8) );
  SDFFX1 DFF_1321_Q_reg ( .D(WX9040), .SI(CRC_OUT_3_8), .SE(n4034), .CLK(n4692), .Q(CRC_OUT_3_9), .QN(DFF_1321_n1) );
  SDFFX1 DFF_1322_Q_reg ( .D(WX9042), .SI(CRC_OUT_3_9), .SE(n4034), .CLK(n4692), .Q(CRC_OUT_3_10) );
  SDFFX1 DFF_1323_Q_reg ( .D(WX9044), .SI(CRC_OUT_3_10), .SE(n4034), .CLK(
        n4692), .Q(CRC_OUT_3_11), .QN(DFF_1323_n1) );
  SDFFX1 DFF_1324_Q_reg ( .D(WX9046), .SI(CRC_OUT_3_11), .SE(n4034), .CLK(
        n4692), .Q(CRC_OUT_3_12), .QN(DFF_1324_n1) );
  SDFFX1 DFF_1325_Q_reg ( .D(WX9048), .SI(CRC_OUT_3_12), .SE(n4034), .CLK(
        n4692), .Q(CRC_OUT_3_13), .QN(DFF_1325_n1) );
  SDFFX1 DFF_1326_Q_reg ( .D(WX9050), .SI(CRC_OUT_3_13), .SE(n4033), .CLK(
        n4692), .Q(CRC_OUT_3_14), .QN(DFF_1326_n1) );
  SDFFX1 DFF_1327_Q_reg ( .D(WX9052), .SI(CRC_OUT_3_14), .SE(n4033), .CLK(
        n4692), .Q(CRC_OUT_3_15) );
  SDFFX1 DFF_1328_Q_reg ( .D(WX9054), .SI(CRC_OUT_3_15), .SE(n4033), .CLK(
        n4692), .Q(CRC_OUT_3_16), .QN(DFF_1328_n1) );
  SDFFX1 DFF_1329_Q_reg ( .D(WX9056), .SI(CRC_OUT_3_16), .SE(n4033), .CLK(
        n4692), .Q(CRC_OUT_3_17), .QN(DFF_1329_n1) );
  SDFFX1 DFF_1330_Q_reg ( .D(WX9058), .SI(CRC_OUT_3_17), .SE(n4033), .CLK(
        n4692), .Q(CRC_OUT_3_18), .QN(DFF_1330_n1) );
  SDFFX1 DFF_1331_Q_reg ( .D(WX9060), .SI(CRC_OUT_3_18), .SE(n4033), .CLK(
        n4692), .Q(CRC_OUT_3_19), .QN(DFF_1331_n1) );
  SDFFX1 DFF_1332_Q_reg ( .D(WX9062), .SI(CRC_OUT_3_19), .SE(n4032), .CLK(
        n4693), .Q(CRC_OUT_3_20), .QN(DFF_1332_n1) );
  SDFFX1 DFF_1333_Q_reg ( .D(WX9064), .SI(CRC_OUT_3_20), .SE(n4032), .CLK(
        n4693), .Q(CRC_OUT_3_21), .QN(DFF_1333_n1) );
  SDFFX1 DFF_1334_Q_reg ( .D(WX9066), .SI(CRC_OUT_3_21), .SE(n4032), .CLK(
        n4693), .Q(CRC_OUT_3_22), .QN(DFF_1334_n1) );
  SDFFX1 DFF_1335_Q_reg ( .D(WX9068), .SI(CRC_OUT_3_22), .SE(n4032), .CLK(
        n4693), .Q(CRC_OUT_3_23), .QN(DFF_1335_n1) );
  SDFFX1 DFF_1336_Q_reg ( .D(WX9070), .SI(CRC_OUT_3_23), .SE(n4032), .CLK(
        n4693), .Q(test_so77) );
  SDFFX1 DFF_1337_Q_reg ( .D(WX9072), .SI(test_si78), .SE(n4032), .CLK(n4693), 
        .Q(CRC_OUT_3_25) );
  SDFFX1 DFF_1338_Q_reg ( .D(WX9074), .SI(CRC_OUT_3_25), .SE(n4031), .CLK(
        n4693), .Q(CRC_OUT_3_26), .QN(DFF_1338_n1) );
  SDFFX1 DFF_1339_Q_reg ( .D(WX9076), .SI(CRC_OUT_3_26), .SE(n4031), .CLK(
        n4693), .Q(CRC_OUT_3_27), .QN(DFF_1339_n1) );
  SDFFX1 DFF_1340_Q_reg ( .D(WX9078), .SI(CRC_OUT_3_27), .SE(n4100), .CLK(
        n4659), .Q(CRC_OUT_3_28), .QN(DFF_1340_n1) );
  SDFFX1 DFF_1341_Q_reg ( .D(WX9080), .SI(CRC_OUT_3_28), .SE(n4100), .CLK(
        n4659), .Q(CRC_OUT_3_29), .QN(DFF_1341_n1) );
  SDFFX1 DFF_1342_Q_reg ( .D(WX9082), .SI(CRC_OUT_3_29), .SE(n4100), .CLK(
        n4659), .Q(CRC_OUT_3_30), .QN(DFF_1342_n1) );
  SDFFX1 DFF_1343_Q_reg ( .D(WX9084), .SI(CRC_OUT_3_30), .SE(n4100), .CLK(
        n4659), .Q(CRC_OUT_3_31), .QN(DFF_1343_n1) );
  SDFFX1 DFF_1344_Q_reg ( .D(n502), .SI(CRC_OUT_3_31), .SE(n4100), .CLK(n4659), 
        .Q(WX9536) );
  SDFFX1 DFF_1345_Q_reg ( .D(n503), .SI(WX9536), .SE(n4095), .CLK(n4661), .Q(
        n8353) );
  SDFFX1 DFF_1346_Q_reg ( .D(n504), .SI(n8353), .SE(n4095), .CLK(n4661), .Q(
        n8352) );
  SDFFX1 DFF_1347_Q_reg ( .D(n505), .SI(n8352), .SE(n4095), .CLK(n4661), .Q(
        n8351) );
  SDFFX1 DFF_1348_Q_reg ( .D(n506), .SI(n8351), .SE(n4095), .CLK(n4661), .Q(
        n8350) );
  SDFFX1 DFF_1349_Q_reg ( .D(n507), .SI(n8350), .SE(n4095), .CLK(n4661), .Q(
        n8349) );
  SDFFX1 DFF_1350_Q_reg ( .D(n508), .SI(n8349), .SE(n4095), .CLK(n4661), .Q(
        n8348) );
  SDFFX1 DFF_1351_Q_reg ( .D(n509), .SI(n8348), .SE(n4096), .CLK(n4661), .Q(
        n8347) );
  SDFFX1 DFF_1352_Q_reg ( .D(n510), .SI(n8347), .SE(n4096), .CLK(n4661), .Q(
        n8346) );
  SDFFX1 DFF_1353_Q_reg ( .D(n511), .SI(n8346), .SE(n4096), .CLK(n4661), .Q(
        test_so78) );
  SDFFX1 DFF_1354_Q_reg ( .D(n512), .SI(test_si79), .SE(n4096), .CLK(n4661), 
        .Q(n8343) );
  SDFFX1 DFF_1355_Q_reg ( .D(n513), .SI(n8343), .SE(n4096), .CLK(n4661), .Q(
        n8342) );
  SDFFX1 DFF_1356_Q_reg ( .D(n514), .SI(n8342), .SE(n4096), .CLK(n4661), .Q(
        n8341) );
  SDFFX1 DFF_1357_Q_reg ( .D(n515), .SI(n8341), .SE(n4097), .CLK(n4660), .Q(
        n8340) );
  SDFFX1 DFF_1358_Q_reg ( .D(n516), .SI(n8340), .SE(n4097), .CLK(n4660), .Q(
        n8339) );
  SDFFX1 DFF_1359_Q_reg ( .D(n517), .SI(n8339), .SE(n4097), .CLK(n4660), .Q(
        n8338) );
  SDFFX1 DFF_1360_Q_reg ( .D(n518), .SI(n8338), .SE(n4097), .CLK(n4660), .Q(
        n8337) );
  SDFFX1 DFF_1361_Q_reg ( .D(n519), .SI(n8337), .SE(n4097), .CLK(n4660), .Q(
        n8336) );
  SDFFX1 DFF_1362_Q_reg ( .D(n520), .SI(n8336), .SE(n4097), .CLK(n4660), .Q(
        n8335) );
  SDFFX1 DFF_1363_Q_reg ( .D(n521), .SI(n8335), .SE(n4098), .CLK(n4660), .Q(
        n8334) );
  SDFFX1 DFF_1364_Q_reg ( .D(n522), .SI(n8334), .SE(n4098), .CLK(n4660), .Q(
        n8333) );
  SDFFX1 DFF_1365_Q_reg ( .D(n523), .SI(n8333), .SE(n4098), .CLK(n4660), .Q(
        n8332) );
  SDFFX1 DFF_1366_Q_reg ( .D(n524), .SI(n8332), .SE(n4098), .CLK(n4660), .Q(
        n8331) );
  SDFFX1 DFF_1367_Q_reg ( .D(n525), .SI(n8331), .SE(n4098), .CLK(n4660), .Q(
        n8330) );
  SDFFX1 DFF_1368_Q_reg ( .D(n526), .SI(n8330), .SE(n4098), .CLK(n4660), .Q(
        n8329) );
  SDFFX1 DFF_1369_Q_reg ( .D(n527), .SI(n8329), .SE(n4099), .CLK(n4659), .Q(
        n8328) );
  SDFFX1 DFF_1370_Q_reg ( .D(n528), .SI(n8328), .SE(n4099), .CLK(n4659), .Q(
        test_so79) );
  SDFFX1 DFF_1371_Q_reg ( .D(n529), .SI(test_si80), .SE(n4099), .CLK(n4659), 
        .Q(n8325) );
  SDFFX1 DFF_1372_Q_reg ( .D(n530), .SI(n8325), .SE(n4099), .CLK(n4659), .Q(
        n8324) );
  SDFFX1 DFF_1373_Q_reg ( .D(n531), .SI(n8324), .SE(n4099), .CLK(n4659), .Q(
        n8323) );
  SDFFX1 DFF_1374_Q_reg ( .D(n532), .SI(n8323), .SE(n4099), .CLK(n4659), .Q(
        n8322) );
  SDFFX1 DFF_1375_Q_reg ( .D(WX9597), .SI(n8322), .SE(n4100), .CLK(n4659), .Q(
        n8321) );
  SDFFX1 DFF_1376_Q_reg ( .D(WX9695), .SI(n8321), .SE(n4094), .CLK(n4662), .Q(
        n8320), .QN(n7109) );
  SDFFX1 DFF_1377_Q_reg ( .D(WX9697), .SI(n8320), .SE(n4094), .CLK(n4662), .Q(
        n8319), .QN(n7108) );
  SDFFX1 DFF_1378_Q_reg ( .D(WX9699), .SI(n8319), .SE(n4094), .CLK(n4662), .Q(
        n8318), .QN(n7107) );
  SDFFX1 DFF_1379_Q_reg ( .D(WX9701), .SI(n8318), .SE(n4093), .CLK(n4662), .Q(
        n8317), .QN(n7106) );
  SDFFX1 DFF_1380_Q_reg ( .D(WX9703), .SI(n8317), .SE(n4093), .CLK(n4662), .Q(
        n8316), .QN(n7105) );
  SDFFX1 DFF_1381_Q_reg ( .D(WX9705), .SI(n8316), .SE(n4093), .CLK(n4662), .Q(
        n8315), .QN(n7104) );
  SDFFX1 DFF_1382_Q_reg ( .D(WX9707), .SI(n8315), .SE(n4092), .CLK(n4663), .Q(
        n8314), .QN(n7103) );
  SDFFX1 DFF_1383_Q_reg ( .D(WX9709), .SI(n8314), .SE(n4092), .CLK(n4663), .Q(
        n8313), .QN(n7102) );
  SDFFX1 DFF_1384_Q_reg ( .D(WX9711), .SI(n8313), .SE(n4092), .CLK(n4663), .Q(
        n8312), .QN(n7101) );
  SDFFX1 DFF_1385_Q_reg ( .D(WX9713), .SI(n8312), .SE(n4091), .CLK(n4663), .Q(
        n8311), .QN(n7100) );
  SDFFX1 DFF_1386_Q_reg ( .D(WX9715), .SI(n8311), .SE(n4091), .CLK(n4663), .Q(
        n8310), .QN(n7099) );
  SDFFX1 DFF_1387_Q_reg ( .D(WX9717), .SI(n8310), .SE(n4036), .CLK(n4691), .Q(
        test_so80) );
  SDFFX1 DFF_1388_Q_reg ( .D(WX9719), .SI(test_si81), .SE(n4090), .CLK(n4664), 
        .Q(n8307), .QN(n7097) );
  SDFFX1 DFF_1389_Q_reg ( .D(WX9721), .SI(n8307), .SE(n4090), .CLK(n4664), .Q(
        n8306), .QN(n7096) );
  SDFFX1 DFF_1390_Q_reg ( .D(WX9723), .SI(n8306), .SE(n4037), .CLK(n4690), .Q(
        n8305), .QN(n7095) );
  SDFFX1 DFF_1391_Q_reg ( .D(WX9725), .SI(n8305), .SE(n4089), .CLK(n4664), .Q(
        n8304), .QN(n7094) );
  SDFFX1 DFF_1392_Q_reg ( .D(WX9727), .SI(n8304), .SE(n4036), .CLK(n4691), .Q(
        WX9728), .QN(n3317) );
  SDFFX1 DFF_1393_Q_reg ( .D(WX9729), .SI(WX9728), .SE(n4088), .CLK(n4665), 
        .Q(WX9730) );
  SDFFX1 DFF_1394_Q_reg ( .D(WX9731), .SI(WX9730), .SE(n4088), .CLK(n4665), 
        .Q(WX9732), .QN(n3315) );
  SDFFX1 DFF_1395_Q_reg ( .D(WX9733), .SI(WX9732), .SE(n4088), .CLK(n4665), 
        .Q(WX9734), .QN(n3314) );
  SDFFX1 DFF_1396_Q_reg ( .D(WX9735), .SI(WX9734), .SE(n4087), .CLK(n4665), 
        .Q(WX9736), .QN(n3313) );
  SDFFX1 DFF_1397_Q_reg ( .D(WX9737), .SI(WX9736), .SE(n4086), .CLK(n4666), 
        .Q(WX9738), .QN(n3312) );
  SDFFX1 DFF_1398_Q_reg ( .D(WX9739), .SI(WX9738), .SE(n4086), .CLK(n4666), 
        .Q(WX9740), .QN(n3311) );
  SDFFX1 DFF_1399_Q_reg ( .D(WX9741), .SI(WX9740), .SE(n4085), .CLK(n4666), 
        .Q(WX9742), .QN(n3310) );
  SDFFX1 DFF_1400_Q_reg ( .D(WX9743), .SI(WX9742), .SE(n4084), .CLK(n4667), 
        .Q(WX9744), .QN(n3309) );
  SDFFX1 DFF_1401_Q_reg ( .D(WX9745), .SI(WX9744), .SE(n4084), .CLK(n4667), 
        .Q(WX9746), .QN(n3308) );
  SDFFX1 DFF_1402_Q_reg ( .D(WX9747), .SI(WX9746), .SE(n4083), .CLK(n4667), 
        .Q(WX9748), .QN(n3307) );
  SDFFX1 DFF_1403_Q_reg ( .D(WX9749), .SI(WX9748), .SE(n4082), .CLK(n4668), 
        .Q(WX9750), .QN(n3306) );
  SDFFX1 DFF_1404_Q_reg ( .D(WX9751), .SI(WX9750), .SE(n4082), .CLK(n4668), 
        .Q(test_so81) );
  SDFFX1 DFF_1405_Q_reg ( .D(WX9753), .SI(test_si82), .SE(n4039), .CLK(n4689), 
        .Q(WX9754), .QN(n3305) );
  SDFFX1 DFF_1406_Q_reg ( .D(WX9755), .SI(WX9754), .SE(n4080), .CLK(n4669), 
        .Q(WX9756) );
  SDFFX1 DFF_1407_Q_reg ( .D(WX9757), .SI(WX9756), .SE(n4080), .CLK(n4669), 
        .Q(WX9758), .QN(n3303) );
  SDFFX1 DFF_1408_Q_reg ( .D(n533), .SI(WX9758), .SE(n4094), .CLK(n4662), .Q(
        WX9760), .QN(n3063) );
  SDFFX1 DFF_1409_Q_reg ( .D(n534), .SI(WX9760), .SE(n4094), .CLK(n4662), .Q(
        WX9762), .QN(n3127) );
  SDFFX1 DFF_1410_Q_reg ( .D(n535), .SI(WX9762), .SE(n4094), .CLK(n4662), .Q(
        WX9764), .QN(n3125) );
  SDFFX1 DFF_1411_Q_reg ( .D(n536), .SI(WX9764), .SE(n4093), .CLK(n4662), .Q(
        WX9766), .QN(n3123) );
  SDFFX1 DFF_1412_Q_reg ( .D(n537), .SI(WX9766), .SE(n4093), .CLK(n4662), .Q(
        WX9768), .QN(n3121) );
  SDFFX1 DFF_1413_Q_reg ( .D(n538), .SI(WX9768), .SE(n4093), .CLK(n4662), .Q(
        WX9770), .QN(n3119) );
  SDFFX1 DFF_1414_Q_reg ( .D(n539), .SI(WX9770), .SE(n4092), .CLK(n4663), .Q(
        WX9772), .QN(n3117) );
  SDFFX1 DFF_1415_Q_reg ( .D(n540), .SI(WX9772), .SE(n4092), .CLK(n4663), .Q(
        WX9774), .QN(n3115) );
  SDFFX1 DFF_1416_Q_reg ( .D(n541), .SI(WX9774), .SE(n4092), .CLK(n4663), .Q(
        WX9776), .QN(n3113) );
  SDFFX1 DFF_1417_Q_reg ( .D(n542), .SI(WX9776), .SE(n4091), .CLK(n4663), .Q(
        WX9778), .QN(n3111) );
  SDFFX1 DFF_1418_Q_reg ( .D(n543), .SI(WX9778), .SE(n4091), .CLK(n4663), .Q(
        WX9780), .QN(n3109) );
  SDFFX1 DFF_1419_Q_reg ( .D(n544), .SI(WX9780), .SE(n4091), .CLK(n4663), .Q(
        WX9782), .QN(n3108) );
  SDFFX1 DFF_1420_Q_reg ( .D(n545), .SI(WX9782), .SE(n4091), .CLK(n4663), .Q(
        WX9784), .QN(n3106) );
  SDFFX1 DFF_1421_Q_reg ( .D(n546), .SI(WX9784), .SE(n4090), .CLK(n4664), .Q(
        test_so82) );
  SDFFX1 DFF_1422_Q_reg ( .D(n547), .SI(test_si83), .SE(n4036), .CLK(n4691), 
        .Q(WX9788), .QN(n3103) );
  SDFFX1 DFF_1423_Q_reg ( .D(n548), .SI(WX9788), .SE(n4089), .CLK(n4664), .Q(
        WX9790), .QN(n3102) );
  SDFFX1 DFF_1424_Q_reg ( .D(WX9791), .SI(WX9790), .SE(n4089), .CLK(n4664), 
        .Q(WX9792) );
  SDFFX1 DFF_1425_Q_reg ( .D(WX9793), .SI(WX9792), .SE(n4089), .CLK(n4664), 
        .Q(WX9794), .QN(n3591) );
  SDFFX1 DFF_1426_Q_reg ( .D(WX9795), .SI(WX9794), .SE(n4088), .CLK(n4665), 
        .Q(WX9796) );
  SDFFX1 DFF_1427_Q_reg ( .D(WX9797), .SI(WX9796), .SE(n4087), .CLK(n4665), 
        .Q(WX9798) );
  SDFFX1 DFF_1428_Q_reg ( .D(WX9799), .SI(WX9798), .SE(n4087), .CLK(n4665), 
        .Q(WX9800) );
  SDFFX1 DFF_1429_Q_reg ( .D(WX9801), .SI(WX9800), .SE(n4086), .CLK(n4666), 
        .Q(WX9802) );
  SDFFX1 DFF_1430_Q_reg ( .D(WX9803), .SI(WX9802), .SE(n4085), .CLK(n4666), 
        .Q(WX9804) );
  SDFFX1 DFF_1431_Q_reg ( .D(WX9805), .SI(WX9804), .SE(n4085), .CLK(n4666), 
        .Q(WX9806) );
  SDFFX1 DFF_1432_Q_reg ( .D(WX9807), .SI(WX9806), .SE(n4084), .CLK(n4667), 
        .Q(WX9808) );
  SDFFX1 DFF_1433_Q_reg ( .D(WX9809), .SI(WX9808), .SE(n4083), .CLK(n4667), 
        .Q(WX9810) );
  SDFFX1 DFF_1434_Q_reg ( .D(WX9811), .SI(WX9810), .SE(n4083), .CLK(n4667), 
        .Q(WX9812) );
  SDFFX1 DFF_1435_Q_reg ( .D(WX9813), .SI(WX9812), .SE(n4082), .CLK(n4668), 
        .Q(WX9814) );
  SDFFX1 DFF_1436_Q_reg ( .D(WX9815), .SI(WX9814), .SE(n4081), .CLK(n4668), 
        .Q(WX9816), .QN(n3569) );
  SDFFX1 DFF_1437_Q_reg ( .D(WX9817), .SI(WX9816), .SE(n4081), .CLK(n4668), 
        .Q(WX9818) );
  SDFFX1 DFF_1438_Q_reg ( .D(WX9819), .SI(WX9818), .SE(n4080), .CLK(n4669), 
        .Q(test_so83) );
  SDFFX1 DFF_1439_Q_reg ( .D(WX9821), .SI(test_si84), .SE(n4080), .CLK(n4669), 
        .Q(WX9822) );
  SDFFX1 DFF_1440_Q_reg ( .D(WX9823), .SI(WX9822), .SE(n4079), .CLK(n4669), 
        .Q(WX9824) );
  SDFFX1 DFF_1441_Q_reg ( .D(WX9825), .SI(WX9824), .SE(n4079), .CLK(n4669), 
        .Q(WX9826) );
  SDFFX1 DFF_1442_Q_reg ( .D(WX9827), .SI(WX9826), .SE(n4078), .CLK(n4670), 
        .Q(WX9828) );
  SDFFX1 DFF_1443_Q_reg ( .D(WX9829), .SI(WX9828), .SE(n4078), .CLK(n4670), 
        .Q(WX9830) );
  SDFFX1 DFF_1444_Q_reg ( .D(WX9831), .SI(WX9830), .SE(n4078), .CLK(n4670), 
        .Q(WX9832) );
  SDFFX1 DFF_1445_Q_reg ( .D(WX9833), .SI(WX9832), .SE(n4077), .CLK(n4670), 
        .Q(WX9834) );
  SDFFX1 DFF_1446_Q_reg ( .D(WX9835), .SI(WX9834), .SE(n4077), .CLK(n4670), 
        .Q(WX9836) );
  SDFFX1 DFF_1447_Q_reg ( .D(WX9837), .SI(WX9836), .SE(n4077), .CLK(n4670), 
        .Q(WX9838) );
  SDFFX1 DFF_1448_Q_reg ( .D(WX9839), .SI(WX9838), .SE(n4076), .CLK(n4671), 
        .Q(WX9840) );
  SDFFX1 DFF_1449_Q_reg ( .D(WX9841), .SI(WX9840), .SE(n4076), .CLK(n4671), 
        .Q(WX9842) );
  SDFFX1 DFF_1450_Q_reg ( .D(WX9843), .SI(WX9842), .SE(n4076), .CLK(n4671), 
        .Q(WX9844) );
  SDFFX1 DFF_1451_Q_reg ( .D(WX9845), .SI(WX9844), .SE(n4075), .CLK(n4671), 
        .Q(WX9846), .QN(n7098) );
  SDFFX1 DFF_1452_Q_reg ( .D(WX9847), .SI(WX9846), .SE(n4075), .CLK(n4671), 
        .Q(WX9848) );
  SDFFX1 DFF_1453_Q_reg ( .D(WX9849), .SI(WX9848), .SE(n4090), .CLK(n4664), 
        .Q(WX9850), .QN(n3105) );
  SDFFX1 DFF_1454_Q_reg ( .D(WX9851), .SI(WX9850), .SE(n4090), .CLK(n4664), 
        .Q(WX9852) );
  SDFFX1 DFF_1455_Q_reg ( .D(WX9853), .SI(WX9852), .SE(n4090), .CLK(n4664), 
        .Q(test_so84) );
  SDFFX1 DFF_1456_Q_reg ( .D(WX9855), .SI(test_si85), .SE(n4089), .CLK(n4664), 
        .Q(WX9856), .QN(n7093) );
  SDFFX1 DFF_1457_Q_reg ( .D(WX9857), .SI(WX9856), .SE(n4089), .CLK(n4664), 
        .Q(WX9858), .QN(n3316) );
  SDFFX1 DFF_1458_Q_reg ( .D(WX9859), .SI(WX9858), .SE(n4088), .CLK(n4665), 
        .Q(WX9860), .QN(n7092) );
  SDFFX1 DFF_1459_Q_reg ( .D(WX9861), .SI(WX9860), .SE(n4087), .CLK(n4665), 
        .Q(WX9862), .QN(n7091) );
  SDFFX1 DFF_1460_Q_reg ( .D(WX9863), .SI(WX9862), .SE(n4087), .CLK(n4665), 
        .Q(WX9864), .QN(n7090) );
  SDFFX1 DFF_1461_Q_reg ( .D(WX9865), .SI(WX9864), .SE(n4086), .CLK(n4666), 
        .Q(WX9866), .QN(n7089) );
  SDFFX1 DFF_1462_Q_reg ( .D(WX9867), .SI(WX9866), .SE(n4085), .CLK(n4666), 
        .Q(WX9868), .QN(n7088) );
  SDFFX1 DFF_1463_Q_reg ( .D(WX9869), .SI(WX9868), .SE(n4085), .CLK(n4666), 
        .Q(WX9870), .QN(n7087) );
  SDFFX1 DFF_1464_Q_reg ( .D(WX9871), .SI(WX9870), .SE(n4084), .CLK(n4667), 
        .Q(WX9872), .QN(n7086) );
  SDFFX1 DFF_1465_Q_reg ( .D(WX9873), .SI(WX9872), .SE(n4083), .CLK(n4667), 
        .Q(WX9874), .QN(n7085) );
  SDFFX1 DFF_1466_Q_reg ( .D(WX9875), .SI(WX9874), .SE(n4083), .CLK(n4667), 
        .Q(WX9876), .QN(n7084) );
  SDFFX1 DFF_1467_Q_reg ( .D(WX9877), .SI(WX9876), .SE(n4082), .CLK(n4668), 
        .Q(WX9878), .QN(n7083) );
  SDFFX1 DFF_1468_Q_reg ( .D(WX9879), .SI(WX9878), .SE(n4081), .CLK(n4668), 
        .Q(WX9880) );
  SDFFX1 DFF_1469_Q_reg ( .D(WX9881), .SI(WX9880), .SE(n4081), .CLK(n4668), 
        .Q(WX9882), .QN(n7082) );
  SDFFX1 DFF_1470_Q_reg ( .D(WX9883), .SI(WX9882), .SE(n4080), .CLK(n4669), 
        .Q(WX9884), .QN(n3304) );
  SDFFX1 DFF_1471_Q_reg ( .D(WX9885), .SI(WX9884), .SE(n4079), .CLK(n4669), 
        .Q(WX9886), .QN(n7081) );
  SDFFX1 DFF_1472_Q_reg ( .D(WX9887), .SI(WX9886), .SE(n4079), .CLK(n4669), 
        .Q(test_so85) );
  SDFFX1 DFF_1473_Q_reg ( .D(WX9889), .SI(test_si86), .SE(n4079), .CLK(n4669), 
        .Q(WX9890), .QN(n3468) );
  SDFFX1 DFF_1474_Q_reg ( .D(WX9891), .SI(WX9890), .SE(n4078), .CLK(n4670), 
        .Q(WX9892), .QN(n3470) );
  SDFFX1 DFF_1475_Q_reg ( .D(WX9893), .SI(WX9892), .SE(n4078), .CLK(n4670), 
        .Q(WX9894), .QN(n3472) );
  SDFFX1 DFF_1476_Q_reg ( .D(WX9895), .SI(WX9894), .SE(n4078), .CLK(n4670), 
        .Q(WX9896), .QN(n3474) );
  SDFFX1 DFF_1477_Q_reg ( .D(WX9897), .SI(WX9896), .SE(n4077), .CLK(n4670), 
        .Q(WX9898), .QN(n3476) );
  SDFFX1 DFF_1478_Q_reg ( .D(WX9899), .SI(WX9898), .SE(n4077), .CLK(n4670), 
        .Q(WX9900), .QN(n3478) );
  SDFFX1 DFF_1479_Q_reg ( .D(WX9901), .SI(WX9900), .SE(n4077), .CLK(n4670), 
        .Q(WX9902), .QN(n3480) );
  SDFFX1 DFF_1480_Q_reg ( .D(WX9903), .SI(WX9902), .SE(n4076), .CLK(n4671), 
        .Q(WX9904), .QN(n3482) );
  SDFFX1 DFF_1481_Q_reg ( .D(WX9905), .SI(WX9904), .SE(n4076), .CLK(n4671), 
        .Q(WX9906), .QN(n3484) );
  SDFFX1 DFF_1482_Q_reg ( .D(WX9907), .SI(WX9906), .SE(n4076), .CLK(n4671), 
        .Q(WX9908), .QN(n3486) );
  SDFFX1 DFF_1483_Q_reg ( .D(WX9909), .SI(WX9908), .SE(n4075), .CLK(n4671), 
        .Q(WX9910), .QN(n3487) );
  SDFFX1 DFF_1484_Q_reg ( .D(WX9911), .SI(WX9910), .SE(n4075), .CLK(n4671), 
        .Q(WX9912), .QN(n3488) );
  SDFFX1 DFF_1485_Q_reg ( .D(WX9913), .SI(WX9912), .SE(n4075), .CLK(n4671), 
        .Q(WX9914), .QN(n3490) );
  SDFFX1 DFF_1486_Q_reg ( .D(WX9915), .SI(WX9914), .SE(n4075), .CLK(n4671), 
        .Q(WX9916), .QN(n3492) );
  SDFFX1 DFF_1487_Q_reg ( .D(WX9917), .SI(WX9916), .SE(n4074), .CLK(n4672), 
        .Q(WX9918), .QN(n3415) );
  SDFFX1 DFF_1488_Q_reg ( .D(WX9919), .SI(WX9918), .SE(n4074), .CLK(n4672), 
        .Q(WX9920), .QN(n3494) );
  SDFFX1 DFF_1489_Q_reg ( .D(WX9921), .SI(WX9920), .SE(n4074), .CLK(n4672), 
        .Q(test_so86) );
  SDFFX1 DFF_1490_Q_reg ( .D(WX9923), .SI(test_si87), .SE(n4088), .CLK(n4665), 
        .Q(WX9924), .QN(n3496) );
  SDFFX1 DFF_1491_Q_reg ( .D(WX9925), .SI(WX9924), .SE(n4087), .CLK(n4665), 
        .Q(WX9926), .QN(n3498) );
  SDFFX1 DFF_1492_Q_reg ( .D(WX9927), .SI(WX9926), .SE(n4086), .CLK(n4666), 
        .Q(WX9928), .QN(n3416) );
  SDFFX1 DFF_1493_Q_reg ( .D(WX9929), .SI(WX9928), .SE(n4086), .CLK(n4666), 
        .Q(WX9930), .QN(n3500) );
  SDFFX1 DFF_1494_Q_reg ( .D(WX9931), .SI(WX9930), .SE(n4085), .CLK(n4666), 
        .Q(WX9932), .QN(n3502) );
  SDFFX1 DFF_1495_Q_reg ( .D(WX9933), .SI(WX9932), .SE(n4084), .CLK(n4667), 
        .Q(WX9934), .QN(n3504) );
  SDFFX1 DFF_1496_Q_reg ( .D(WX9935), .SI(WX9934), .SE(n4084), .CLK(n4667), 
        .Q(WX9936), .QN(n3506) );
  SDFFX1 DFF_1497_Q_reg ( .D(WX9937), .SI(WX9936), .SE(n4083), .CLK(n4667), 
        .Q(WX9938), .QN(n3508) );
  SDFFX1 DFF_1498_Q_reg ( .D(WX9939), .SI(WX9938), .SE(n4082), .CLK(n4668), 
        .Q(WX9940), .QN(n3510) );
  SDFFX1 DFF_1499_Q_reg ( .D(WX9941), .SI(WX9940), .SE(n4082), .CLK(n4668), 
        .Q(WX9942), .QN(n3417) );
  SDFFX1 DFF_1500_Q_reg ( .D(WX9943), .SI(WX9942), .SE(n4081), .CLK(n4668), 
        .Q(WX9944), .QN(n3512) );
  SDFFX1 DFF_1501_Q_reg ( .D(WX9945), .SI(WX9944), .SE(n4081), .CLK(n4668), 
        .Q(WX9946), .QN(n3514) );
  SDFFX1 DFF_1502_Q_reg ( .D(WX9947), .SI(WX9946), .SE(n4080), .CLK(n4669), 
        .Q(WX9948), .QN(n3516) );
  SDFFX1 DFF_1503_Q_reg ( .D(WX9949), .SI(WX9948), .SE(n4079), .CLK(n4669), 
        .Q(WX9950), .QN(n3434) );
  SDFFX1 DFF_1504_Q_reg ( .D(WX10315), .SI(WX9950), .SE(n4040), .CLK(n4689), 
        .Q(CRC_OUT_2_0), .QN(DFF_1504_n1) );
  SDFFX1 DFF_1505_Q_reg ( .D(WX10317), .SI(CRC_OUT_2_0), .SE(n4040), .CLK(
        n4689), .Q(CRC_OUT_2_1), .QN(DFF_1505_n1) );
  SDFFX1 DFF_1506_Q_reg ( .D(WX10319), .SI(CRC_OUT_2_1), .SE(n4039), .CLK(
        n4689), .Q(test_so87) );
  SDFFX1 DFF_1507_Q_reg ( .D(WX10321), .SI(test_si88), .SE(n4039), .CLK(n4689), 
        .Q(CRC_OUT_2_3) );
  SDFFX1 DFF_1508_Q_reg ( .D(WX10323), .SI(CRC_OUT_2_3), .SE(n4039), .CLK(
        n4689), .Q(CRC_OUT_2_4), .QN(DFF_1508_n1) );
  SDFFX1 DFF_1509_Q_reg ( .D(WX10325), .SI(CRC_OUT_2_4), .SE(n4039), .CLK(
        n4689), .Q(CRC_OUT_2_5), .QN(DFF_1509_n1) );
  SDFFX1 DFF_1510_Q_reg ( .D(WX10327), .SI(CRC_OUT_2_5), .SE(n4039), .CLK(
        n4689), .Q(CRC_OUT_2_6), .QN(DFF_1510_n1) );
  SDFFX1 DFF_1511_Q_reg ( .D(WX10329), .SI(CRC_OUT_2_6), .SE(n4038), .CLK(
        n4690), .Q(CRC_OUT_2_7), .QN(DFF_1511_n1) );
  SDFFX1 DFF_1512_Q_reg ( .D(WX10331), .SI(CRC_OUT_2_7), .SE(n4038), .CLK(
        n4690), .Q(CRC_OUT_2_8), .QN(DFF_1512_n1) );
  SDFFX1 DFF_1513_Q_reg ( .D(WX10333), .SI(CRC_OUT_2_8), .SE(n4038), .CLK(
        n4690), .Q(CRC_OUT_2_9), .QN(DFF_1513_n1) );
  SDFFX1 DFF_1514_Q_reg ( .D(WX10335), .SI(CRC_OUT_2_9), .SE(n4038), .CLK(
        n4690), .Q(CRC_OUT_2_10) );
  SDFFX1 DFF_1515_Q_reg ( .D(WX10337), .SI(CRC_OUT_2_10), .SE(n4038), .CLK(
        n4690), .Q(CRC_OUT_2_11), .QN(DFF_1515_n1) );
  SDFFX1 DFF_1516_Q_reg ( .D(WX10339), .SI(CRC_OUT_2_11), .SE(n4038), .CLK(
        n4690), .Q(CRC_OUT_2_12), .QN(DFF_1516_n1) );
  SDFFX1 DFF_1517_Q_reg ( .D(WX10341), .SI(CRC_OUT_2_12), .SE(n4037), .CLK(
        n4690), .Q(CRC_OUT_2_13) );
  SDFFX1 DFF_1518_Q_reg ( .D(WX10343), .SI(CRC_OUT_2_13), .SE(n4037), .CLK(
        n4690), .Q(CRC_OUT_2_14), .QN(DFF_1518_n1) );
  SDFFX1 DFF_1519_Q_reg ( .D(WX10345), .SI(CRC_OUT_2_14), .SE(n4037), .CLK(
        n4690), .Q(CRC_OUT_2_15) );
  SDFFX1 DFF_1520_Q_reg ( .D(WX10347), .SI(CRC_OUT_2_15), .SE(n4037), .CLK(
        n4690), .Q(CRC_OUT_2_16), .QN(DFF_1520_n1) );
  SDFFX1 DFF_1521_Q_reg ( .D(WX10349), .SI(CRC_OUT_2_16), .SE(n4037), .CLK(
        n4690), .Q(CRC_OUT_2_17), .QN(DFF_1521_n1) );
  SDFFX1 DFF_1522_Q_reg ( .D(WX10351), .SI(CRC_OUT_2_17), .SE(n4036), .CLK(
        n4691), .Q(CRC_OUT_2_18), .QN(DFF_1522_n1) );
  SDFFX1 DFF_1523_Q_reg ( .D(WX10353), .SI(CRC_OUT_2_18), .SE(n4074), .CLK(
        n4672), .Q(test_so88) );
  SDFFX1 DFF_1524_Q_reg ( .D(WX10355), .SI(test_si89), .SE(n4074), .CLK(n4672), 
        .Q(CRC_OUT_2_20), .QN(DFF_1524_n1) );
  SDFFX1 DFF_1525_Q_reg ( .D(WX10357), .SI(CRC_OUT_2_20), .SE(n4074), .CLK(
        n4672), .Q(CRC_OUT_2_21), .QN(DFF_1525_n1) );
  SDFFX1 DFF_1526_Q_reg ( .D(WX10359), .SI(CRC_OUT_2_21), .SE(n4073), .CLK(
        n4672), .Q(CRC_OUT_2_22), .QN(DFF_1526_n1) );
  SDFFX1 DFF_1527_Q_reg ( .D(WX10361), .SI(CRC_OUT_2_22), .SE(n4073), .CLK(
        n4672), .Q(CRC_OUT_2_23), .QN(DFF_1527_n1) );
  SDFFX1 DFF_1528_Q_reg ( .D(WX10363), .SI(CRC_OUT_2_23), .SE(n4073), .CLK(
        n4672), .Q(CRC_OUT_2_24), .QN(DFF_1528_n1) );
  SDFFX1 DFF_1529_Q_reg ( .D(WX10365), .SI(CRC_OUT_2_24), .SE(n4073), .CLK(
        n4672), .Q(CRC_OUT_2_25), .QN(DFF_1529_n1) );
  SDFFX1 DFF_1530_Q_reg ( .D(WX10367), .SI(CRC_OUT_2_25), .SE(n4073), .CLK(
        n4672), .Q(CRC_OUT_2_26), .QN(DFF_1530_n1) );
  SDFFX1 DFF_1531_Q_reg ( .D(WX10369), .SI(CRC_OUT_2_26), .SE(n4073), .CLK(
        n4672), .Q(CRC_OUT_2_27), .QN(DFF_1531_n1) );
  SDFFX1 DFF_1532_Q_reg ( .D(WX10371), .SI(CRC_OUT_2_27), .SE(n4072), .CLK(
        n4673), .Q(CRC_OUT_2_28), .QN(DFF_1532_n1) );
  SDFFX1 DFF_1533_Q_reg ( .D(WX10373), .SI(CRC_OUT_2_28), .SE(n4072), .CLK(
        n4673), .Q(CRC_OUT_2_29), .QN(DFF_1533_n1) );
  SDFFX1 DFF_1534_Q_reg ( .D(WX10375), .SI(CRC_OUT_2_29), .SE(n4072), .CLK(
        n4673), .Q(CRC_OUT_2_30) );
  SDFFX1 DFF_1535_Q_reg ( .D(WX10377), .SI(CRC_OUT_2_30), .SE(n4072), .CLK(
        n4673), .Q(CRC_OUT_2_31), .QN(DFF_1535_n1) );
  SDFFX1 DFF_1536_Q_reg ( .D(n580), .SI(CRC_OUT_2_31), .SE(n4072), .CLK(n4673), 
        .Q(WX10829) );
  SDFFX1 DFF_1537_Q_reg ( .D(n581), .SI(WX10829), .SE(n4067), .CLK(n4675), .Q(
        n8295) );
  SDFFX1 DFF_1538_Q_reg ( .D(n582), .SI(n8295), .SE(n4067), .CLK(n4675), .Q(
        n8294) );
  SDFFX1 DFF_1539_Q_reg ( .D(n583), .SI(n8294), .SE(n4067), .CLK(n4675), .Q(
        n8293) );
  SDFFX1 DFF_1540_Q_reg ( .D(n584), .SI(n8293), .SE(n4067), .CLK(n4675), .Q(
        test_so89) );
  SDFFX1 DFF_1541_Q_reg ( .D(n585), .SI(test_si90), .SE(n4067), .CLK(n4675), 
        .Q(n8290) );
  SDFFX1 DFF_1542_Q_reg ( .D(n586), .SI(n8290), .SE(n4067), .CLK(n4675), .Q(
        n8289) );
  SDFFX1 DFF_1543_Q_reg ( .D(n587), .SI(n8289), .SE(n4068), .CLK(n4675), .Q(
        n8288) );
  SDFFX1 DFF_1544_Q_reg ( .D(n588), .SI(n8288), .SE(n4068), .CLK(n4675), .Q(
        n8287) );
  SDFFX1 DFF_1545_Q_reg ( .D(n589), .SI(n8287), .SE(n4068), .CLK(n4675), .Q(
        n8286) );
  SDFFX1 DFF_1546_Q_reg ( .D(n590), .SI(n8286), .SE(n4068), .CLK(n4675), .Q(
        n8285) );
  SDFFX1 DFF_1547_Q_reg ( .D(n591), .SI(n8285), .SE(n4068), .CLK(n4675), .Q(
        n8284) );
  SDFFX1 DFF_1548_Q_reg ( .D(n592), .SI(n8284), .SE(n4068), .CLK(n4675), .Q(
        n8283) );
  SDFFX1 DFF_1549_Q_reg ( .D(n593), .SI(n8283), .SE(n4069), .CLK(n4674), .Q(
        n8282) );
  SDFFX1 DFF_1550_Q_reg ( .D(n594), .SI(n8282), .SE(n4069), .CLK(n4674), .Q(
        n8281) );
  SDFFX1 DFF_1551_Q_reg ( .D(n595), .SI(n8281), .SE(n4069), .CLK(n4674), .Q(
        n8280) );
  SDFFX1 DFF_1552_Q_reg ( .D(n596), .SI(n8280), .SE(n4069), .CLK(n4674), .Q(
        n8279) );
  SDFFX1 DFF_1553_Q_reg ( .D(n597), .SI(n8279), .SE(n4069), .CLK(n4674), .Q(
        n8278) );
  SDFFX1 DFF_1554_Q_reg ( .D(n598), .SI(n8278), .SE(n4069), .CLK(n4674), .Q(
        n8277) );
  SDFFX1 DFF_1555_Q_reg ( .D(n599), .SI(n8277), .SE(n4070), .CLK(n4674), .Q(
        n8276) );
  SDFFX1 DFF_1556_Q_reg ( .D(n600), .SI(n8276), .SE(n4070), .CLK(n4674), .Q(
        n8275) );
  SDFFX1 DFF_1557_Q_reg ( .D(n601), .SI(n8275), .SE(n4070), .CLK(n4674), .Q(
        test_so90) );
  SDFFX1 DFF_1558_Q_reg ( .D(n602), .SI(test_si91), .SE(n4070), .CLK(n4674), 
        .Q(n8272) );
  SDFFX1 DFF_1559_Q_reg ( .D(n603), .SI(n8272), .SE(n4070), .CLK(n4674), .Q(
        n8271) );
  SDFFX1 DFF_1560_Q_reg ( .D(n604), .SI(n8271), .SE(n4070), .CLK(n4674), .Q(
        n8270) );
  SDFFX1 DFF_1561_Q_reg ( .D(n605), .SI(n8270), .SE(n4071), .CLK(n4673), .Q(
        n8269) );
  SDFFX1 DFF_1562_Q_reg ( .D(n606), .SI(n8269), .SE(n4071), .CLK(n4673), .Q(
        n8268) );
  SDFFX1 DFF_1563_Q_reg ( .D(n607), .SI(n8268), .SE(n4071), .CLK(n4673), .Q(
        n8267) );
  SDFFX1 DFF_1564_Q_reg ( .D(n608), .SI(n8267), .SE(n4071), .CLK(n4673), .Q(
        n8266) );
  SDFFX1 DFF_1565_Q_reg ( .D(n609), .SI(n8266), .SE(n4071), .CLK(n4673), .Q(
        n8265) );
  SDFFX1 DFF_1566_Q_reg ( .D(n610), .SI(n8265), .SE(n4071), .CLK(n4673), .Q(
        n8264) );
  SDFFX1 DFF_1567_Q_reg ( .D(WX10890), .SI(n8264), .SE(n4072), .CLK(n4673), 
        .Q(n8263) );
  SDFFX1 DFF_1568_Q_reg ( .D(WX10988), .SI(n8263), .SE(n4066), .CLK(n4676), 
        .Q(n8262), .QN(n7069) );
  SDFFX1 DFF_1569_Q_reg ( .D(WX10990), .SI(n8262), .SE(n4066), .CLK(n4676), 
        .Q(n8261), .QN(n7070) );
  SDFFX1 DFF_1570_Q_reg ( .D(WX10992), .SI(n8261), .SE(n4066), .CLK(n4676), 
        .Q(n8260), .QN(n7071) );
  SDFFX1 DFF_1571_Q_reg ( .D(WX10994), .SI(n8260), .SE(n4065), .CLK(n4676), 
        .Q(n8259), .QN(n7072) );
  SDFFX1 DFF_1572_Q_reg ( .D(WX10996), .SI(n8259), .SE(n4065), .CLK(n4676), 
        .Q(n8258), .QN(n7073) );
  SDFFX1 DFF_1573_Q_reg ( .D(WX10998), .SI(n8258), .SE(n4065), .CLK(n4676), 
        .Q(n8257), .QN(n7074) );
  SDFFX1 DFF_1574_Q_reg ( .D(WX11000), .SI(n8257), .SE(n4064), .CLK(n4677), 
        .Q(test_so91) );
  SDFFX1 DFF_1575_Q_reg ( .D(WX11002), .SI(test_si92), .SE(n4064), .CLK(n4677), 
        .Q(n8254), .QN(n7075) );
  SDFFX1 DFF_1576_Q_reg ( .D(WX11004), .SI(n8254), .SE(n4064), .CLK(n4677), 
        .Q(n8253), .QN(n7254) );
  SDFFX1 DFF_1577_Q_reg ( .D(WX11006), .SI(n8253), .SE(n4040), .CLK(n4689), 
        .Q(n8252), .QN(n7076) );
  SDFFX1 DFF_1578_Q_reg ( .D(WX11008), .SI(n8252), .SE(n4063), .CLK(n4677), 
        .Q(n8251), .QN(n7253) );
  SDFFX1 DFF_1579_Q_reg ( .D(WX11010), .SI(n8251), .SE(n4062), .CLK(n4678), 
        .Q(n8250), .QN(n7077) );
  SDFFX1 DFF_1580_Q_reg ( .D(WX11012), .SI(n8250), .SE(n4062), .CLK(n4678), 
        .Q(n8249), .QN(n7252) );
  SDFFX1 DFF_1581_Q_reg ( .D(WX11014), .SI(n8249), .SE(n4061), .CLK(n4678), 
        .Q(n8248), .QN(n7078) );
  SDFFX1 DFF_1582_Q_reg ( .D(WX11016), .SI(n8248), .SE(n4061), .CLK(n4678), 
        .Q(n8247), .QN(n7079) );
  SDFFX1 DFF_1583_Q_reg ( .D(WX11018), .SI(n8247), .SE(n4060), .CLK(n4679), 
        .Q(n8246), .QN(n7080) );
  SDFFX1 DFF_1584_Q_reg ( .D(WX11020), .SI(n8246), .SE(n4060), .CLK(n4679), 
        .Q(WX11021), .QN(n3302) );
  SDFFX1 DFF_1585_Q_reg ( .D(WX11022), .SI(WX11021), .SE(n4059), .CLK(n4679), 
        .Q(WX11023), .QN(n3301) );
  SDFFX1 DFF_1586_Q_reg ( .D(WX11024), .SI(WX11023), .SE(n4058), .CLK(n4680), 
        .Q(WX11025), .QN(n3300) );
  SDFFX1 DFF_1587_Q_reg ( .D(WX11026), .SI(WX11025), .SE(n4058), .CLK(n4680), 
        .Q(WX11027), .QN(n3299) );
  SDFFX1 DFF_1588_Q_reg ( .D(WX11028), .SI(WX11027), .SE(n4057), .CLK(n4680), 
        .Q(WX11029), .QN(n3298) );
  SDFFX1 DFF_1589_Q_reg ( .D(WX11030), .SI(WX11029), .SE(n4056), .CLK(n4681), 
        .Q(WX11031), .QN(n3297) );
  SDFFX1 DFF_1590_Q_reg ( .D(WX11032), .SI(WX11031), .SE(n4056), .CLK(n4681), 
        .Q(WX11033), .QN(n3296) );
  SDFFX1 DFF_1591_Q_reg ( .D(WX11034), .SI(WX11033), .SE(n4055), .CLK(n4681), 
        .Q(test_so92) );
  SDFFX1 DFF_1592_Q_reg ( .D(WX11036), .SI(test_si93), .SE(n4040), .CLK(n4689), 
        .Q(WX11037), .QN(n3295) );
  SDFFX1 DFF_1593_Q_reg ( .D(WX11038), .SI(WX11037), .SE(n4053), .CLK(n4682), 
        .Q(WX11039) );
  SDFFX1 DFF_1594_Q_reg ( .D(WX11040), .SI(WX11039), .SE(n4053), .CLK(n4682), 
        .Q(WX11041), .QN(n3293) );
  SDFFX1 DFF_1595_Q_reg ( .D(WX11042), .SI(WX11041), .SE(n4052), .CLK(n4683), 
        .Q(WX11043) );
  SDFFX1 DFF_1596_Q_reg ( .D(WX11044), .SI(WX11043), .SE(n4052), .CLK(n4683), 
        .Q(WX11045), .QN(n3292) );
  SDFFX1 DFF_1597_Q_reg ( .D(WX11046), .SI(WX11045), .SE(n4051), .CLK(n4683), 
        .Q(WX11047) );
  SDFFX1 DFF_1598_Q_reg ( .D(WX11048), .SI(WX11047), .SE(n4050), .CLK(n4684), 
        .Q(WX11049), .QN(n3290) );
  SDFFX1 DFF_1599_Q_reg ( .D(WX11050), .SI(WX11049), .SE(n4050), .CLK(n4684), 
        .Q(WX11051), .QN(n3289) );
  SDFFX1 DFF_1600_Q_reg ( .D(WX11052), .SI(WX11051), .SE(n4066), .CLK(n4676), 
        .Q(WX11053), .QN(n3061) );
  SDFFX1 DFF_1601_Q_reg ( .D(WX11054), .SI(WX11053), .SE(n4066), .CLK(n4676), 
        .Q(WX11055), .QN(n3100) );
  SDFFX1 DFF_1602_Q_reg ( .D(WX11056), .SI(WX11055), .SE(n4066), .CLK(n4676), 
        .Q(WX11057), .QN(n3098) );
  SDFFX1 DFF_1603_Q_reg ( .D(WX11058), .SI(WX11057), .SE(n4065), .CLK(n4676), 
        .Q(WX11059), .QN(n3096) );
  SDFFX1 DFF_1604_Q_reg ( .D(WX11060), .SI(WX11059), .SE(n4065), .CLK(n4676), 
        .Q(WX11061), .QN(n3094) );
  SDFFX1 DFF_1605_Q_reg ( .D(WX11062), .SI(WX11061), .SE(n4065), .CLK(n4676), 
        .Q(WX11063), .QN(n3092) );
  SDFFX1 DFF_1606_Q_reg ( .D(WX11064), .SI(WX11063), .SE(n4064), .CLK(n4677), 
        .Q(WX11065), .QN(n3091) );
  SDFFX1 DFF_1607_Q_reg ( .D(WX11066), .SI(WX11065), .SE(n4064), .CLK(n4677), 
        .Q(WX11067), .QN(n3089) );
  SDFFX1 DFF_1608_Q_reg ( .D(n619), .SI(WX11067), .SE(n4064), .CLK(n4677), .Q(
        test_so93) );
  SDFFX1 DFF_1609_Q_reg ( .D(WX11070), .SI(test_si94), .SE(n4040), .CLK(n4689), 
        .Q(WX11071), .QN(n3086) );
  SDFFX1 DFF_1610_Q_reg ( .D(n621), .SI(WX11071), .SE(n4063), .CLK(n4677), .Q(
        WX11073), .QN(n3085) );
  SDFFX1 DFF_1611_Q_reg ( .D(WX11074), .SI(WX11073), .SE(n4063), .CLK(n4677), 
        .Q(WX11075), .QN(n3083) );
  SDFFX1 DFF_1612_Q_reg ( .D(n623), .SI(WX11075), .SE(n4062), .CLK(n4678), .Q(
        WX11077), .QN(n3082) );
  SDFFX1 DFF_1613_Q_reg ( .D(WX11078), .SI(WX11077), .SE(n4062), .CLK(n4678), 
        .Q(WX11079), .QN(n3080) );
  SDFFX1 DFF_1614_Q_reg ( .D(WX11080), .SI(WX11079), .SE(n4061), .CLK(n4678), 
        .Q(WX11081), .QN(n3078) );
  SDFFX1 DFF_1615_Q_reg ( .D(WX11082), .SI(WX11081), .SE(n4060), .CLK(n4679), 
        .Q(WX11083), .QN(n3076) );
  SDFFX1 DFF_1616_Q_reg ( .D(WX11084), .SI(WX11083), .SE(n4059), .CLK(n4679), 
        .Q(WX11085) );
  SDFFX1 DFF_1617_Q_reg ( .D(WX11086), .SI(WX11085), .SE(n4059), .CLK(n4679), 
        .Q(WX11087) );
  SDFFX1 DFF_1618_Q_reg ( .D(WX11088), .SI(WX11087), .SE(n4058), .CLK(n4680), 
        .Q(WX11089) );
  SDFFX1 DFF_1619_Q_reg ( .D(WX11090), .SI(WX11089), .SE(n4057), .CLK(n4680), 
        .Q(WX11091) );
  SDFFX1 DFF_1620_Q_reg ( .D(WX11092), .SI(WX11091), .SE(n4057), .CLK(n4680), 
        .Q(WX11093) );
  SDFFX1 DFF_1621_Q_reg ( .D(WX11094), .SI(WX11093), .SE(n4056), .CLK(n4681), 
        .Q(WX11095) );
  SDFFX1 DFF_1622_Q_reg ( .D(WX11096), .SI(WX11095), .SE(n4055), .CLK(n4681), 
        .Q(WX11097) );
  SDFFX1 DFF_1623_Q_reg ( .D(WX11098), .SI(WX11097), .SE(n4055), .CLK(n4681), 
        .Q(WX11099), .QN(n3547) );
  SDFFX1 DFF_1624_Q_reg ( .D(WX11100), .SI(WX11099), .SE(n4054), .CLK(n4682), 
        .Q(WX11101) );
  SDFFX1 DFF_1625_Q_reg ( .D(WX11102), .SI(WX11101), .SE(n4054), .CLK(n4682), 
        .Q(test_so94) );
  SDFFX1 DFF_1626_Q_reg ( .D(WX11104), .SI(test_si95), .SE(n4053), .CLK(n4682), 
        .Q(WX11105) );
  SDFFX1 DFF_1627_Q_reg ( .D(WX11106), .SI(WX11105), .SE(n4052), .CLK(n4683), 
        .Q(WX11107), .QN(n3539) );
  SDFFX1 DFF_1628_Q_reg ( .D(WX11108), .SI(WX11107), .SE(n4052), .CLK(n4683), 
        .Q(WX11109) );
  SDFFX1 DFF_1629_Q_reg ( .D(WX11110), .SI(WX11109), .SE(n4051), .CLK(n4683), 
        .Q(WX11111), .QN(n3535) );
  SDFFX1 DFF_1630_Q_reg ( .D(WX11112), .SI(WX11111), .SE(n4050), .CLK(n4684), 
        .Q(WX11113) );
  SDFFX1 DFF_1631_Q_reg ( .D(WX11114), .SI(WX11113), .SE(n4050), .CLK(n4684), 
        .Q(WX11115) );
  SDFFX1 DFF_1632_Q_reg ( .D(WX11116), .SI(WX11115), .SE(n4049), .CLK(n4684), 
        .Q(WX11117) );
  SDFFX1 DFF_1633_Q_reg ( .D(WX11118), .SI(WX11117), .SE(n4049), .CLK(n4684), 
        .Q(WX11119) );
  SDFFX1 DFF_1634_Q_reg ( .D(WX11120), .SI(WX11119), .SE(n4048), .CLK(n4685), 
        .Q(WX11121) );
  SDFFX1 DFF_1635_Q_reg ( .D(WX11122), .SI(WX11121), .SE(n4048), .CLK(n4685), 
        .Q(WX11123) );
  SDFFX1 DFF_1636_Q_reg ( .D(WX11124), .SI(WX11123), .SE(n4048), .CLK(n4685), 
        .Q(WX11125) );
  SDFFX1 DFF_1637_Q_reg ( .D(WX11126), .SI(WX11125), .SE(n4047), .CLK(n4685), 
        .Q(WX11127) );
  SDFFX1 DFF_1638_Q_reg ( .D(WX11128), .SI(WX11127), .SE(n4047), .CLK(n4685), 
        .Q(WX11129), .QN(n7255) );
  SDFFX1 DFF_1639_Q_reg ( .D(WX11130), .SI(WX11129), .SE(n4047), .CLK(n4685), 
        .Q(WX11131) );
  SDFFX1 DFF_1640_Q_reg ( .D(WX11132), .SI(WX11131), .SE(n4063), .CLK(n4677), 
        .Q(WX11133), .QN(n3088) );
  SDFFX1 DFF_1641_Q_reg ( .D(WX11134), .SI(WX11133), .SE(n4063), .CLK(n4677), 
        .Q(WX11135) );
  SDFFX1 DFF_1642_Q_reg ( .D(WX11136), .SI(WX11135), .SE(n4063), .CLK(n4677), 
        .Q(test_so95) );
  SDFFX1 DFF_1643_Q_reg ( .D(WX11138), .SI(test_si96), .SE(n4062), .CLK(n4678), 
        .Q(WX11139) );
  SDFFX1 DFF_1644_Q_reg ( .D(WX11140), .SI(WX11139), .SE(n4062), .CLK(n4678), 
        .Q(WX11141) );
  SDFFX1 DFF_1645_Q_reg ( .D(WX11142), .SI(WX11141), .SE(n4061), .CLK(n4678), 
        .Q(WX11143) );
  SDFFX1 DFF_1646_Q_reg ( .D(WX11144), .SI(WX11143), .SE(n4061), .CLK(n4678), 
        .Q(WX11145) );
  SDFFX1 DFF_1647_Q_reg ( .D(WX11146), .SI(WX11145), .SE(n4060), .CLK(n4679), 
        .Q(WX11147) );
  SDFFX1 DFF_1648_Q_reg ( .D(WX11148), .SI(WX11147), .SE(n4059), .CLK(n4679), 
        .Q(WX11149), .QN(n7251) );
  SDFFX1 DFF_1649_Q_reg ( .D(WX11150), .SI(WX11149), .SE(n4059), .CLK(n4679), 
        .Q(WX11151), .QN(n7250) );
  SDFFX1 DFF_1650_Q_reg ( .D(WX11152), .SI(WX11151), .SE(n4058), .CLK(n4680), 
        .Q(WX11153), .QN(n7249) );
  SDFFX1 DFF_1651_Q_reg ( .D(WX11154), .SI(WX11153), .SE(n4057), .CLK(n4680), 
        .Q(WX11155), .QN(n7248) );
  SDFFX1 DFF_1652_Q_reg ( .D(WX11156), .SI(WX11155), .SE(n4057), .CLK(n4680), 
        .Q(WX11157), .QN(n7247) );
  SDFFX1 DFF_1653_Q_reg ( .D(WX11158), .SI(WX11157), .SE(n4056), .CLK(n4681), 
        .Q(WX11159), .QN(n7246) );
  SDFFX1 DFF_1654_Q_reg ( .D(WX11160), .SI(WX11159), .SE(n4055), .CLK(n4681), 
        .Q(WX11161), .QN(n7245) );
  SDFFX1 DFF_1655_Q_reg ( .D(WX11162), .SI(WX11161), .SE(n4055), .CLK(n4681), 
        .Q(WX11163) );
  SDFFX1 DFF_1656_Q_reg ( .D(WX11164), .SI(WX11163), .SE(n4054), .CLK(n4682), 
        .Q(WX11165), .QN(n7244) );
  SDFFX1 DFF_1657_Q_reg ( .D(WX11166), .SI(WX11165), .SE(n4054), .CLK(n4682), 
        .Q(WX11167), .QN(n3294) );
  SDFFX1 DFF_1658_Q_reg ( .D(WX11168), .SI(WX11167), .SE(n4053), .CLK(n4682), 
        .Q(WX11169), .QN(n7243) );
  SDFFX1 DFF_1659_Q_reg ( .D(WX11170), .SI(WX11169), .SE(n4052), .CLK(n4683), 
        .Q(test_so96) );
  SDFFX1 DFF_1660_Q_reg ( .D(WX11172), .SI(test_si97), .SE(n4051), .CLK(n4683), 
        .Q(WX11173), .QN(n7242) );
  SDFFX1 DFF_1661_Q_reg ( .D(WX11174), .SI(WX11173), .SE(n4051), .CLK(n4683), 
        .Q(WX11175), .QN(n3291) );
  SDFFX1 DFF_1662_Q_reg ( .D(WX11176), .SI(WX11175), .SE(n4050), .CLK(n4684), 
        .Q(WX11177), .QN(n7241) );
  SDFFX1 DFF_1663_Q_reg ( .D(WX11178), .SI(WX11177), .SE(n4049), .CLK(n4684), 
        .Q(WX11179), .QN(n7240) );
  SDFFX1 DFF_1664_Q_reg ( .D(WX11180), .SI(WX11179), .SE(n4049), .CLK(n4684), 
        .Q(WX11181), .QN(n3441) );
  SDFFX1 DFF_1665_Q_reg ( .D(WX11182), .SI(WX11181), .SE(n4049), .CLK(n4684), 
        .Q(WX11183), .QN(n3442) );
  SDFFX1 DFF_1666_Q_reg ( .D(WX11184), .SI(WX11183), .SE(n4048), .CLK(n4685), 
        .Q(WX11185), .QN(n3443) );
  SDFFX1 DFF_1667_Q_reg ( .D(WX11186), .SI(WX11185), .SE(n4048), .CLK(n4685), 
        .Q(WX11187), .QN(n3444) );
  SDFFX1 DFF_1668_Q_reg ( .D(WX11188), .SI(WX11187), .SE(n4048), .CLK(n4685), 
        .Q(WX11189), .QN(n3445) );
  SDFFX1 DFF_1669_Q_reg ( .D(WX11190), .SI(WX11189), .SE(n4047), .CLK(n4685), 
        .Q(WX11191), .QN(n3446) );
  SDFFX1 DFF_1670_Q_reg ( .D(WX11192), .SI(WX11191), .SE(n4047), .CLK(n4685), 
        .Q(WX11193), .QN(n3447) );
  SDFFX1 DFF_1671_Q_reg ( .D(WX11194), .SI(WX11193), .SE(n4047), .CLK(n4685), 
        .Q(WX11195), .QN(n3448) );
  SDFFX1 DFF_1672_Q_reg ( .D(WX11196), .SI(WX11195), .SE(n4046), .CLK(n4686), 
        .Q(WX11197), .QN(n3449) );
  SDFFX1 DFF_1673_Q_reg ( .D(WX11198), .SI(WX11197), .SE(n4046), .CLK(n4686), 
        .Q(WX11199), .QN(n3450) );
  SDFFX1 DFF_1674_Q_reg ( .D(WX11200), .SI(WX11199), .SE(n4046), .CLK(n4686), 
        .Q(WX11201), .QN(n3451) );
  SDFFX1 DFF_1675_Q_reg ( .D(WX11202), .SI(WX11201), .SE(n4046), .CLK(n4686), 
        .Q(WX11203), .QN(n3452) );
  SDFFX1 DFF_1676_Q_reg ( .D(WX11204), .SI(WX11203), .SE(n4046), .CLK(n4686), 
        .Q(test_so97) );
  SDFFX1 DFF_1677_Q_reg ( .D(WX11206), .SI(test_si98), .SE(n4061), .CLK(n4678), 
        .Q(WX11207), .QN(n3453) );
  SDFFX1 DFF_1678_Q_reg ( .D(WX11208), .SI(WX11207), .SE(n4060), .CLK(n4679), 
        .Q(WX11209), .QN(n3454) );
  SDFFX1 DFF_1679_Q_reg ( .D(WX11210), .SI(WX11209), .SE(n4060), .CLK(n4679), 
        .Q(WX11211), .QN(n3412) );
  SDFFX1 DFF_1680_Q_reg ( .D(WX11212), .SI(WX11211), .SE(n4059), .CLK(n4679), 
        .Q(WX11213), .QN(n3455) );
  SDFFX1 DFF_1681_Q_reg ( .D(WX11214), .SI(WX11213), .SE(n4058), .CLK(n4680), 
        .Q(WX11215), .QN(n3456) );
  SDFFX1 DFF_1682_Q_reg ( .D(WX11216), .SI(WX11215), .SE(n4058), .CLK(n4680), 
        .Q(WX11217), .QN(n3457) );
  SDFFX1 DFF_1683_Q_reg ( .D(WX11218), .SI(WX11217), .SE(n4057), .CLK(n4680), 
        .Q(WX11219), .QN(n3458) );
  SDFFX1 DFF_1684_Q_reg ( .D(WX11220), .SI(WX11219), .SE(n4056), .CLK(n4681), 
        .Q(WX11221), .QN(n3413) );
  SDFFX1 DFF_1685_Q_reg ( .D(WX11222), .SI(WX11221), .SE(n4056), .CLK(n4681), 
        .Q(WX11223), .QN(n3459) );
  SDFFX1 DFF_1686_Q_reg ( .D(WX11224), .SI(WX11223), .SE(n4055), .CLK(n4681), 
        .Q(WX11225), .QN(n3460) );
  SDFFX1 DFF_1687_Q_reg ( .D(WX11226), .SI(WX11225), .SE(n4054), .CLK(n4682), 
        .Q(WX11227), .QN(n3461) );
  SDFFX1 DFF_1688_Q_reg ( .D(WX11228), .SI(WX11227), .SE(n4054), .CLK(n4682), 
        .Q(WX11229), .QN(n3462) );
  SDFFX1 DFF_1689_Q_reg ( .D(WX11230), .SI(WX11229), .SE(n4053), .CLK(n4682), 
        .Q(WX11231), .QN(n3463) );
  SDFFX1 DFF_1690_Q_reg ( .D(WX11232), .SI(WX11231), .SE(n4053), .CLK(n4682), 
        .Q(WX11233), .QN(n3464) );
  SDFFX1 DFF_1691_Q_reg ( .D(WX11234), .SI(WX11233), .SE(n4052), .CLK(n4683), 
        .Q(WX11235), .QN(n3414) );
  SDFFX1 DFF_1692_Q_reg ( .D(WX11236), .SI(WX11235), .SE(n4051), .CLK(n4683), 
        .Q(WX11237), .QN(n3465) );
  SDFFX1 DFF_1693_Q_reg ( .D(WX11238), .SI(WX11237), .SE(n4051), .CLK(n4683), 
        .Q(test_so98) );
  SDFFX1 DFF_1694_Q_reg ( .D(WX11240), .SI(test_si99), .SE(n4050), .CLK(n4684), 
        .Q(WX11241), .QN(n3466) );
  SDFFX1 DFF_1695_Q_reg ( .D(WX11242), .SI(WX11241), .SE(n4049), .CLK(n4684), 
        .Q(WX11243), .QN(n3433) );
  SDFFX1 DFF_1696_Q_reg ( .D(WX11608), .SI(WX11243), .SE(n4044), .CLK(n4687), 
        .Q(CRC_OUT_1_0), .QN(DFF_1696_n1) );
  SDFFX1 DFF_1697_Q_reg ( .D(WX11610), .SI(CRC_OUT_1_0), .SE(n4044), .CLK(
        n4687), .Q(CRC_OUT_1_1) );
  SDFFX1 DFF_1698_Q_reg ( .D(WX11612), .SI(CRC_OUT_1_1), .SE(n4044), .CLK(
        n4687), .Q(CRC_OUT_1_2), .QN(DFF_1698_n1) );
  SDFFX1 DFF_1699_Q_reg ( .D(WX11614), .SI(CRC_OUT_1_2), .SE(n4044), .CLK(
        n4687), .Q(CRC_OUT_1_3), .QN(DFF_1699_n1) );
  SDFFX1 DFF_1700_Q_reg ( .D(WX11616), .SI(CRC_OUT_1_3), .SE(n4044), .CLK(
        n4687), .Q(CRC_OUT_1_4), .QN(DFF_1700_n1) );
  SDFFX1 DFF_1701_Q_reg ( .D(WX11618), .SI(CRC_OUT_1_4), .SE(n4043), .CLK(
        n4687), .Q(CRC_OUT_1_5), .QN(DFF_1701_n1) );
  SDFFX1 DFF_1702_Q_reg ( .D(WX11620), .SI(CRC_OUT_1_5), .SE(n4043), .CLK(
        n4687), .Q(CRC_OUT_1_6), .QN(DFF_1702_n1) );
  SDFFX1 DFF_1703_Q_reg ( .D(WX11622), .SI(CRC_OUT_1_6), .SE(n4043), .CLK(
        n4687), .Q(CRC_OUT_1_7), .QN(DFF_1703_n1) );
  SDFFX1 DFF_1704_Q_reg ( .D(WX11624), .SI(CRC_OUT_1_7), .SE(n4043), .CLK(
        n4687), .Q(CRC_OUT_1_8), .QN(DFF_1704_n1) );
  SDFFX1 DFF_1705_Q_reg ( .D(WX11626), .SI(CRC_OUT_1_8), .SE(n4043), .CLK(
        n4687), .Q(CRC_OUT_1_9), .QN(DFF_1705_n1) );
  SDFFX1 DFF_1706_Q_reg ( .D(WX11628), .SI(CRC_OUT_1_9), .SE(n4043), .CLK(
        n4687), .Q(CRC_OUT_1_10), .QN(DFF_1706_n1) );
  SDFFX1 DFF_1707_Q_reg ( .D(WX11630), .SI(CRC_OUT_1_10), .SE(n4042), .CLK(
        n4688), .Q(CRC_OUT_1_11), .QN(DFF_1707_n1) );
  SDFFX1 DFF_1708_Q_reg ( .D(WX11632), .SI(CRC_OUT_1_11), .SE(n4042), .CLK(
        n4688), .Q(CRC_OUT_1_12), .QN(DFF_1708_n1) );
  SDFFX1 DFF_1709_Q_reg ( .D(WX11634), .SI(CRC_OUT_1_12), .SE(n4042), .CLK(
        n4688), .Q(CRC_OUT_1_13), .QN(DFF_1709_n1) );
  SDFFX1 DFF_1710_Q_reg ( .D(WX11636), .SI(CRC_OUT_1_13), .SE(n4042), .CLK(
        n4688), .Q(test_so99) );
  SDFFX1 DFF_1711_Q_reg ( .D(WX11638), .SI(test_si100), .SE(n4042), .CLK(n4688), .Q(CRC_OUT_1_15), .QN(DFF_1711_n1) );
  SDFFX1 DFF_1712_Q_reg ( .D(WX11640), .SI(CRC_OUT_1_15), .SE(n4042), .CLK(
        n4688), .Q(CRC_OUT_1_16), .QN(DFF_1712_n1) );
  SDFFX1 DFF_1713_Q_reg ( .D(WX11642), .SI(CRC_OUT_1_16), .SE(n4041), .CLK(
        n4688), .Q(CRC_OUT_1_17), .QN(DFF_1713_n1) );
  SDFFX1 DFF_1714_Q_reg ( .D(WX11644), .SI(CRC_OUT_1_17), .SE(n4041), .CLK(
        n4688), .Q(CRC_OUT_1_18) );
  SDFFX1 DFF_1715_Q_reg ( .D(WX11646), .SI(CRC_OUT_1_18), .SE(n4041), .CLK(
        n4688), .Q(CRC_OUT_1_19), .QN(DFF_1715_n1) );
  SDFFX1 DFF_1716_Q_reg ( .D(WX11648), .SI(CRC_OUT_1_19), .SE(n4041), .CLK(
        n4688), .Q(CRC_OUT_1_20), .QN(DFF_1716_n1) );
  SDFFX1 DFF_1717_Q_reg ( .D(WX11650), .SI(CRC_OUT_1_20), .SE(n4041), .CLK(
        n4688), .Q(CRC_OUT_1_21), .QN(DFF_1717_n1) );
  SDFFX1 DFF_1718_Q_reg ( .D(WX11652), .SI(CRC_OUT_1_21), .SE(n4041), .CLK(
        n4688), .Q(CRC_OUT_1_22), .QN(DFF_1718_n1) );
  SDFFX1 DFF_1719_Q_reg ( .D(WX11654), .SI(CRC_OUT_1_22), .SE(n4040), .CLK(
        n4689), .Q(CRC_OUT_1_23), .QN(DFF_1719_n1) );
  SDFFX1 DFF_1720_Q_reg ( .D(WX11656), .SI(CRC_OUT_1_23), .SE(n4046), .CLK(
        n4686), .Q(CRC_OUT_1_24), .QN(DFF_1720_n1) );
  SDFFX1 DFF_1721_Q_reg ( .D(WX11658), .SI(CRC_OUT_1_24), .SE(n4045), .CLK(
        n4686), .Q(CRC_OUT_1_25), .QN(DFF_1721_n1) );
  SDFFX1 DFF_1722_Q_reg ( .D(WX11660), .SI(CRC_OUT_1_25), .SE(n4045), .CLK(
        n4686), .Q(CRC_OUT_1_26), .QN(DFF_1722_n1) );
  SDFFX1 DFF_1723_Q_reg ( .D(WX11662), .SI(CRC_OUT_1_26), .SE(n4045), .CLK(
        n4686), .Q(CRC_OUT_1_27), .QN(DFF_1723_n1) );
  SDFFX1 DFF_1724_Q_reg ( .D(WX11664), .SI(CRC_OUT_1_27), .SE(n4045), .CLK(
        n4686), .Q(CRC_OUT_1_28), .QN(DFF_1724_n1) );
  SDFFX1 DFF_1725_Q_reg ( .D(WX11666), .SI(CRC_OUT_1_28), .SE(n4045), .CLK(
        n4686), .Q(CRC_OUT_1_29), .QN(DFF_1725_n1) );
  SDFFX1 DFF_1726_Q_reg ( .D(WX11668), .SI(CRC_OUT_1_29), .SE(n4045), .CLK(
        n4686), .Q(CRC_OUT_1_30), .QN(DFF_1726_n1) );
  SDFFX1 DFF_1727_Q_reg ( .D(WX11670), .SI(CRC_OUT_1_30), .SE(n4044), .CLK(
        n4687), .Q(test_so100) );
  NOR2X0 Trojan1 ( .IN1(WX3442), .IN2(WX5974), .QN(Tj_OUT1) );
  NOR2X0 Trojan2 ( .IN1(WX806), .IN2(WX782), .QN(Tj_OUT2) );
  NOR2X0 Trojan3 ( .IN1(WX11632), .IN2(n128), .QN(Tj_OUT3) );
  NOR2X0 Trojan4 ( .IN1(WX5964), .IN2(n158), .QN(Tj_OUT4) );
  AND4X1 Trojan1234_NOT ( .IN1(Tj_OUT1), .IN2(Tj_OUT2), .IN3(Tj_OUT3), .IN4(
        Tj_OUT4), .Q(Tj_OUT1234) );
  NOR2X0 Trojan5 ( .IN1(WX8634), .IN2(WX3330), .QN(Tj_OUT5) );
  NOR2X0 Trojan6 ( .IN1(n140), .IN2(n132), .QN(Tj_OUT6) );
  NOR2X0 Trojan7 ( .IN1(WX862), .IN2(WX7227), .QN(Tj_OUT7) );
  NOR2X0 Trojan8 ( .IN1(WX11616), .IN2(n597), .QN(Tj_OUT8) );
  AND4X1 Trojan5678_NOT ( .IN1(Tj_OUT5), .IN2(Tj_OUT6), .IN3(Tj_OUT7), .IN4(
        Tj_OUT8), .Q(Tj_OUT5678) );
  INVX0 TrojanINVtest_se ( .INP(n4410), .ZN(test_se_NOT) );
  AND3X1 Trojan_Trigger ( .IN1(Tj_OUT1234), .IN2(Tj_OUT5678), .IN3(test_se_NOT), .Q(Tj_Trigger) );
  INVX0 U3706 ( .INP(TM1), .ZN(n3872) );
  INVX0 U3707 ( .INP(TM1), .ZN(n3873) );
  INVX0 U3708 ( .INP(TM1), .ZN(n3874) );
  INVX0 U3709 ( .INP(TM1), .ZN(n3875) );
  NBUFFX2 U3710 ( .INP(n3907), .Z(n3915) );
  NBUFFX2 U3711 ( .INP(n3912), .Z(n3930) );
  NBUFFX2 U3712 ( .INP(n3907), .Z(n3916) );
  NBUFFX2 U3713 ( .INP(n3907), .Z(n3917) );
  NBUFFX2 U3714 ( .INP(n3908), .Z(n3918) );
  NBUFFX2 U3715 ( .INP(n3908), .Z(n3919) );
  NBUFFX2 U3716 ( .INP(n3909), .Z(n3923) );
  NBUFFX2 U3717 ( .INP(n3910), .Z(n3924) );
  NBUFFX2 U3718 ( .INP(n3910), .Z(n3925) );
  NBUFFX2 U3719 ( .INP(n3910), .Z(n3926) );
  NBUFFX2 U3720 ( .INP(n3911), .Z(n3927) );
  NBUFFX2 U3721 ( .INP(n3911), .Z(n3928) );
  NBUFFX2 U3722 ( .INP(n3911), .Z(n3929) );
  NBUFFX2 U3723 ( .INP(n3908), .Z(n3920) );
  NBUFFX2 U3724 ( .INP(n3909), .Z(n3921) );
  NBUFFX2 U3725 ( .INP(n3909), .Z(n3922) );
  NBUFFX2 U3726 ( .INP(n3958), .Z(n3956) );
  NBUFFX2 U3727 ( .INP(n3962), .Z(n3934) );
  NBUFFX2 U3728 ( .INP(n3962), .Z(n3935) );
  NBUFFX2 U3729 ( .INP(n3962), .Z(n3936) );
  NBUFFX2 U3730 ( .INP(n3962), .Z(n3937) );
  NBUFFX2 U3731 ( .INP(n3960), .Z(n3944) );
  NBUFFX2 U3732 ( .INP(n3960), .Z(n3946) );
  NBUFFX2 U3733 ( .INP(n3960), .Z(n3947) );
  NBUFFX2 U3734 ( .INP(n3959), .Z(n3948) );
  NBUFFX2 U3735 ( .INP(n3959), .Z(n3949) );
  NBUFFX2 U3736 ( .INP(n3959), .Z(n3950) );
  NBUFFX2 U3737 ( .INP(n3961), .Z(n3938) );
  NBUFFX2 U3738 ( .INP(n3961), .Z(n3939) );
  NBUFFX2 U3739 ( .INP(n3960), .Z(n3945) );
  NBUFFX2 U3740 ( .INP(n3961), .Z(n3940) );
  NBUFFX2 U3741 ( .INP(n3961), .Z(n3941) );
  NBUFFX2 U3742 ( .INP(n3961), .Z(n3942) );
  NBUFFX2 U3743 ( .INP(n3960), .Z(n3943) );
  NBUFFX2 U3744 ( .INP(n3959), .Z(n3952) );
  NBUFFX2 U3745 ( .INP(n3959), .Z(n3951) );
  NBUFFX2 U3746 ( .INP(n3958), .Z(n3953) );
  NBUFFX2 U3747 ( .INP(n3958), .Z(n3954) );
  NBUFFX2 U3748 ( .INP(n3958), .Z(n3955) );
  NBUFFX2 U3749 ( .INP(n3958), .Z(n3957) );
  NBUFFX2 U3750 ( .INP(n4741), .Z(n4572) );
  NBUFFX2 U3751 ( .INP(n4741), .Z(n4570) );
  NBUFFX2 U3752 ( .INP(n4741), .Z(n4571) );
  NBUFFX2 U3753 ( .INP(n4741), .Z(n4569) );
  NBUFFX2 U3754 ( .INP(n4717), .Z(n4688) );
  NBUFFX2 U3755 ( .INP(n4718), .Z(n4687) );
  NBUFFX2 U3756 ( .INP(n4718), .Z(n4686) );
  NBUFFX2 U3757 ( .INP(n4718), .Z(n4685) );
  NBUFFX2 U3758 ( .INP(n4718), .Z(n4684) );
  NBUFFX2 U3759 ( .INP(n4718), .Z(n4683) );
  NBUFFX2 U3760 ( .INP(n4719), .Z(n4682) );
  NBUFFX2 U3761 ( .INP(n4719), .Z(n4681) );
  NBUFFX2 U3762 ( .INP(n4719), .Z(n4680) );
  NBUFFX2 U3763 ( .INP(n4719), .Z(n4679) );
  NBUFFX2 U3764 ( .INP(n4719), .Z(n4678) );
  NBUFFX2 U3765 ( .INP(n4720), .Z(n4677) );
  NBUFFX2 U3766 ( .INP(n4720), .Z(n4676) );
  NBUFFX2 U3767 ( .INP(n4720), .Z(n4674) );
  NBUFFX2 U3768 ( .INP(n4720), .Z(n4675) );
  NBUFFX2 U3769 ( .INP(n4720), .Z(n4673) );
  NBUFFX2 U3770 ( .INP(n4721), .Z(n4672) );
  NBUFFX2 U3771 ( .INP(n4721), .Z(n4671) );
  NBUFFX2 U3772 ( .INP(n4721), .Z(n4670) );
  NBUFFX2 U3773 ( .INP(n4721), .Z(n4669) );
  NBUFFX2 U3774 ( .INP(n4717), .Z(n4689) );
  NBUFFX2 U3775 ( .INP(n4721), .Z(n4668) );
  NBUFFX2 U3776 ( .INP(n4722), .Z(n4667) );
  NBUFFX2 U3777 ( .INP(n4722), .Z(n4666) );
  NBUFFX2 U3778 ( .INP(n4722), .Z(n4665) );
  NBUFFX2 U3779 ( .INP(n4717), .Z(n4690) );
  NBUFFX2 U3780 ( .INP(n4722), .Z(n4664) );
  NBUFFX2 U3781 ( .INP(n4722), .Z(n4663) );
  NBUFFX2 U3782 ( .INP(n4723), .Z(n4662) );
  NBUFFX2 U3783 ( .INP(n4723), .Z(n4660) );
  NBUFFX2 U3784 ( .INP(n4723), .Z(n4661) );
  NBUFFX2 U3785 ( .INP(n4723), .Z(n4659) );
  NBUFFX2 U3786 ( .INP(n4717), .Z(n4692) );
  NBUFFX2 U3787 ( .INP(n4717), .Z(n4691) );
  NBUFFX2 U3788 ( .INP(n4723), .Z(n4658) );
  NBUFFX2 U3789 ( .INP(n4724), .Z(n4657) );
  NBUFFX2 U3790 ( .INP(n4724), .Z(n4656) );
  NBUFFX2 U3791 ( .INP(n4724), .Z(n4655) );
  NBUFFX2 U3792 ( .INP(n4724), .Z(n4654) );
  NBUFFX2 U3793 ( .INP(n4724), .Z(n4653) );
  NBUFFX2 U3794 ( .INP(n4725), .Z(n4652) );
  NBUFFX2 U3795 ( .INP(n4725), .Z(n4651) );
  NBUFFX2 U3796 ( .INP(n4725), .Z(n4650) );
  NBUFFX2 U3797 ( .INP(n4725), .Z(n4649) );
  NBUFFX2 U3798 ( .INP(n4725), .Z(n4648) );
  NBUFFX2 U3799 ( .INP(n4726), .Z(n4647) );
  NBUFFX2 U3800 ( .INP(n4726), .Z(n4646) );
  NBUFFX2 U3801 ( .INP(n4716), .Z(n4695) );
  NBUFFX2 U3802 ( .INP(n4716), .Z(n4694) );
  NBUFFX2 U3803 ( .INP(n4716), .Z(n4693) );
  NBUFFX2 U3804 ( .INP(n4726), .Z(n4645) );
  NBUFFX2 U3805 ( .INP(n4726), .Z(n4644) );
  NBUFFX2 U3806 ( .INP(n4726), .Z(n4643) );
  NBUFFX2 U3807 ( .INP(n4727), .Z(n4642) );
  NBUFFX2 U3808 ( .INP(n4727), .Z(n4641) );
  NBUFFX2 U3809 ( .INP(n4727), .Z(n4640) );
  NBUFFX2 U3810 ( .INP(n4727), .Z(n4639) );
  NBUFFX2 U3811 ( .INP(n4727), .Z(n4638) );
  NBUFFX2 U3812 ( .INP(n4728), .Z(n4637) );
  NBUFFX2 U3813 ( .INP(n4728), .Z(n4636) );
  NBUFFX2 U3814 ( .INP(n4728), .Z(n4633) );
  NBUFFX2 U3815 ( .INP(n4728), .Z(n4634) );
  NBUFFX2 U3816 ( .INP(n4728), .Z(n4635) );
  NBUFFX2 U3817 ( .INP(n4729), .Z(n4632) );
  NBUFFX2 U3818 ( .INP(n4716), .Z(n4697) );
  NBUFFX2 U3819 ( .INP(n4716), .Z(n4696) );
  NBUFFX2 U3820 ( .INP(n4729), .Z(n4631) );
  NBUFFX2 U3821 ( .INP(n4729), .Z(n4630) );
  NBUFFX2 U3822 ( .INP(n4729), .Z(n4629) );
  NBUFFX2 U3823 ( .INP(n4729), .Z(n4628) );
  NBUFFX2 U3824 ( .INP(n4730), .Z(n4627) );
  NBUFFX2 U3825 ( .INP(n4730), .Z(n4626) );
  NBUFFX2 U3826 ( .INP(n4730), .Z(n4625) );
  NBUFFX2 U3827 ( .INP(n4730), .Z(n4624) );
  NBUFFX2 U3828 ( .INP(n4730), .Z(n4623) );
  NBUFFX2 U3829 ( .INP(n4731), .Z(n4622) );
  NBUFFX2 U3830 ( .INP(n4731), .Z(n4619) );
  NBUFFX2 U3831 ( .INP(n4731), .Z(n4620) );
  NBUFFX2 U3832 ( .INP(n4731), .Z(n4621) );
  NBUFFX2 U3833 ( .INP(n4715), .Z(n4699) );
  NBUFFX2 U3834 ( .INP(n4715), .Z(n4698) );
  NBUFFX2 U3835 ( .INP(n4731), .Z(n4618) );
  NBUFFX2 U3836 ( .INP(n4732), .Z(n4617) );
  NBUFFX2 U3837 ( .INP(n4732), .Z(n4616) );
  NBUFFX2 U3838 ( .INP(n4732), .Z(n4615) );
  NBUFFX2 U3839 ( .INP(n4732), .Z(n4614) );
  NBUFFX2 U3840 ( .INP(n4732), .Z(n4613) );
  NBUFFX2 U3841 ( .INP(n4735), .Z(n4600) );
  NBUFFX2 U3842 ( .INP(n4715), .Z(n4700) );
  NBUFFX2 U3843 ( .INP(n4733), .Z(n4612) );
  NBUFFX2 U3844 ( .INP(n4733), .Z(n4611) );
  NBUFFX2 U3845 ( .INP(n4733), .Z(n4610) );
  NBUFFX2 U3846 ( .INP(n4733), .Z(n4609) );
  NBUFFX2 U3847 ( .INP(n4734), .Z(n4607) );
  NBUFFX2 U3848 ( .INP(n4733), .Z(n4608) );
  NBUFFX2 U3849 ( .INP(n4734), .Z(n4606) );
  NBUFFX2 U3850 ( .INP(n4715), .Z(n4701) );
  NBUFFX2 U3851 ( .INP(n4714), .Z(n4704) );
  NBUFFX2 U3852 ( .INP(n4734), .Z(n4605) );
  NBUFFX2 U3853 ( .INP(n4714), .Z(n4703) );
  NBUFFX2 U3854 ( .INP(n4734), .Z(n4604) );
  NBUFFX2 U3855 ( .INP(n4734), .Z(n4603) );
  NBUFFX2 U3856 ( .INP(n4735), .Z(n4602) );
  NBUFFX2 U3857 ( .INP(n4735), .Z(n4601) );
  NBUFFX2 U3858 ( .INP(n4715), .Z(n4702) );
  NBUFFX2 U3859 ( .INP(n4735), .Z(n4599) );
  NBUFFX2 U3860 ( .INP(n4735), .Z(n4598) );
  NBUFFX2 U3861 ( .INP(n4736), .Z(n4597) );
  NBUFFX2 U3862 ( .INP(n4736), .Z(n4596) );
  NBUFFX2 U3863 ( .INP(n4736), .Z(n4594) );
  NBUFFX2 U3864 ( .INP(n4736), .Z(n4595) );
  NBUFFX2 U3865 ( .INP(n4736), .Z(n4593) );
  NBUFFX2 U3866 ( .INP(n4714), .Z(n4706) );
  NBUFFX2 U3867 ( .INP(n4714), .Z(n4705) );
  NBUFFX2 U3868 ( .INP(n4713), .Z(n4710) );
  NBUFFX2 U3869 ( .INP(n4713), .Z(n4709) );
  NBUFFX2 U3870 ( .INP(n4713), .Z(n4708) );
  NBUFFX2 U3872 ( .INP(n4737), .Z(n4592) );
  NBUFFX2 U3873 ( .INP(n4737), .Z(n4591) );
  NBUFFX2 U3874 ( .INP(n4737), .Z(n4590) );
  NBUFFX2 U3875 ( .INP(n4714), .Z(n4707) );
  NBUFFX2 U3876 ( .INP(n4737), .Z(n4589) );
  NBUFFX2 U3877 ( .INP(n4737), .Z(n4588) );
  NBUFFX2 U3878 ( .INP(n4738), .Z(n4587) );
  NBUFFX2 U3879 ( .INP(n4738), .Z(n4586) );
  NBUFFX2 U3880 ( .INP(n4738), .Z(n4584) );
  NBUFFX2 U3881 ( .INP(n4738), .Z(n4585) );
  NBUFFX2 U3882 ( .INP(n4738), .Z(n4583) );
  NBUFFX2 U3883 ( .INP(n4713), .Z(n4712) );
  NBUFFX2 U3884 ( .INP(n4713), .Z(n4711) );
  NBUFFX2 U3885 ( .INP(n4739), .Z(n4582) );
  NBUFFX2 U3886 ( .INP(n4739), .Z(n4581) );
  NBUFFX2 U3887 ( .INP(n4739), .Z(n4580) );
  NBUFFX2 U3888 ( .INP(n4739), .Z(n4579) );
  NBUFFX2 U3889 ( .INP(n4739), .Z(n4578) );
  NBUFFX2 U3890 ( .INP(n4740), .Z(n4577) );
  NBUFFX2 U3891 ( .INP(n4740), .Z(n4576) );
  NBUFFX2 U3892 ( .INP(n4740), .Z(n4575) );
  NBUFFX2 U3893 ( .INP(n4740), .Z(n4574) );
  NBUFFX2 U3894 ( .INP(n4740), .Z(n4573) );
  NBUFFX2 U3895 ( .INP(n3912), .Z(n3931) );
  NBUFFX2 U3896 ( .INP(n3989), .Z(n3982) );
  NBUFFX2 U3897 ( .INP(n3988), .Z(n3986) );
  NBUFFX2 U3898 ( .INP(n3988), .Z(n3985) );
  NBUFFX2 U3899 ( .INP(n3988), .Z(n3983) );
  NBUFFX2 U3900 ( .INP(n3988), .Z(n3984) );
  NBUFFX2 U3901 ( .INP(n3902), .Z(n3899) );
  NBUFFX2 U3902 ( .INP(n3902), .Z(n3897) );
  NBUFFX2 U3903 ( .INP(n3902), .Z(n3900) );
  NBUFFX2 U3904 ( .INP(n3902), .Z(n3898) );
  NBUFFX2 U3905 ( .INP(n3903), .Z(n3896) );
  NBUFFX2 U3906 ( .INP(n3989), .Z(n3981) );
  NBUFFX2 U3907 ( .INP(n3988), .Z(n3987) );
  NBUFFX2 U3908 ( .INP(n3992), .Z(n3967) );
  NBUFFX2 U3909 ( .INP(n3992), .Z(n3965) );
  NBUFFX2 U3910 ( .INP(n3992), .Z(n3966) );
  NBUFFX2 U3911 ( .INP(n3906), .Z(n3879) );
  NBUFFX2 U3912 ( .INP(n3906), .Z(n3878) );
  NBUFFX2 U3913 ( .INP(n3906), .Z(n3881) );
  NBUFFX2 U3914 ( .INP(n3906), .Z(n3880) );
  NBUFFX2 U3915 ( .INP(n3990), .Z(n3975) );
  NBUFFX2 U3916 ( .INP(n3990), .Z(n3976) );
  NBUFFX2 U3917 ( .INP(n3990), .Z(n3977) );
  NBUFFX2 U3918 ( .INP(n3989), .Z(n3978) );
  NBUFFX2 U3919 ( .INP(n3991), .Z(n3968) );
  NBUFFX2 U3920 ( .INP(n3991), .Z(n3970) );
  NBUFFX2 U3921 ( .INP(n3991), .Z(n3971) );
  NBUFFX2 U3922 ( .INP(n3991), .Z(n3972) );
  NBUFFX2 U3923 ( .INP(n3990), .Z(n3973) );
  NBUFFX2 U3924 ( .INP(n3990), .Z(n3974) );
  NBUFFX2 U3925 ( .INP(n3989), .Z(n3980) );
  NBUFFX2 U3926 ( .INP(n3989), .Z(n3979) );
  NBUFFX2 U3927 ( .INP(n3991), .Z(n3969) );
  NBUFFX2 U3928 ( .INP(n3905), .Z(n3886) );
  NBUFFX2 U3929 ( .INP(n3905), .Z(n3885) );
  NBUFFX2 U3930 ( .INP(n3905), .Z(n3884) );
  NBUFFX2 U3931 ( .INP(n3905), .Z(n3883) );
  NBUFFX2 U3932 ( .INP(n3905), .Z(n3882) );
  NBUFFX2 U3933 ( .INP(n3904), .Z(n3889) );
  NBUFFX2 U3934 ( .INP(n3904), .Z(n3887) );
  NBUFFX2 U3935 ( .INP(n3904), .Z(n3888) );
  NBUFFX2 U3936 ( .INP(n3903), .Z(n3894) );
  NBUFFX2 U3937 ( .INP(n3903), .Z(n3895) );
  NBUFFX2 U3938 ( .INP(n3903), .Z(n3893) );
  NBUFFX2 U3939 ( .INP(n3903), .Z(n3892) );
  NBUFFX2 U3940 ( .INP(n3904), .Z(n3891) );
  NBUFFX2 U3941 ( .INP(n3904), .Z(n3890) );
  NBUFFX2 U3942 ( .INP(n3914), .Z(n3907) );
  NBUFFX2 U3943 ( .INP(n3913), .Z(n3910) );
  NBUFFX2 U3944 ( .INP(n3913), .Z(n3911) );
  NBUFFX2 U3945 ( .INP(n3914), .Z(n3908) );
  NBUFFX2 U3946 ( .INP(n3914), .Z(n3909) );
  NBUFFX2 U3947 ( .INP(n3913), .Z(n3912) );
  NBUFFX2 U3948 ( .INP(n3902), .Z(n3901) );
  NBUFFX2 U3949 ( .INP(n2148), .Z(n3913) );
  NBUFFX2 U3950 ( .INP(n2148), .Z(n3914) );
  NBUFFX2 U3951 ( .INP(n4761), .Z(n3876) );
  NBUFFX2 U3952 ( .INP(n4761), .Z(n3877) );
  NBUFFX2 U3953 ( .INP(n3876), .Z(n3902) );
  NBUFFX2 U3954 ( .INP(n3876), .Z(n3903) );
  NBUFFX2 U3955 ( .INP(n3876), .Z(n3904) );
  NBUFFX2 U3956 ( .INP(n3877), .Z(n3905) );
  NBUFFX2 U3957 ( .INP(n3877), .Z(n3906) );
  NBUFFX2 U3958 ( .INP(n2152), .Z(n3932) );
  NBUFFX2 U3959 ( .INP(n2152), .Z(n3933) );
  NBUFFX2 U3960 ( .INP(n3932), .Z(n3958) );
  NBUFFX2 U3961 ( .INP(n3932), .Z(n3959) );
  NBUFFX2 U3962 ( .INP(n3932), .Z(n3960) );
  NBUFFX2 U3963 ( .INP(n3933), .Z(n3961) );
  NBUFFX2 U3964 ( .INP(n3933), .Z(n3962) );
  NBUFFX2 U3965 ( .INP(n2153), .Z(n3963) );
  NBUFFX2 U3966 ( .INP(n2153), .Z(n3964) );
  NBUFFX2 U3967 ( .INP(n3963), .Z(n3988) );
  NBUFFX2 U3968 ( .INP(n3963), .Z(n3989) );
  NBUFFX2 U3969 ( .INP(n3963), .Z(n3990) );
  NBUFFX2 U3970 ( .INP(n3964), .Z(n3991) );
  NBUFFX2 U3971 ( .INP(n3964), .Z(n3992) );
  NBUFFX2 U3972 ( .INP(n4377), .Z(n3993) );
  NBUFFX2 U3973 ( .INP(n4376), .Z(n3994) );
  NBUFFX2 U3974 ( .INP(n4376), .Z(n3995) );
  NBUFFX2 U3975 ( .INP(n4376), .Z(n3996) );
  NBUFFX2 U3976 ( .INP(n4375), .Z(n3997) );
  NBUFFX2 U3977 ( .INP(n4375), .Z(n3998) );
  NBUFFX2 U3978 ( .INP(n4375), .Z(n3999) );
  NBUFFX2 U3979 ( .INP(n4374), .Z(n4000) );
  NBUFFX2 U3980 ( .INP(n4374), .Z(n4001) );
  NBUFFX2 U3981 ( .INP(n4374), .Z(n4002) );
  NBUFFX2 U3982 ( .INP(n4373), .Z(n4003) );
  NBUFFX2 U3983 ( .INP(n4373), .Z(n4004) );
  NBUFFX2 U3984 ( .INP(n4373), .Z(n4005) );
  NBUFFX2 U3985 ( .INP(n4372), .Z(n4006) );
  NBUFFX2 U3986 ( .INP(n4372), .Z(n4007) );
  NBUFFX2 U3987 ( .INP(n4372), .Z(n4008) );
  NBUFFX2 U3988 ( .INP(n4371), .Z(n4009) );
  NBUFFX2 U3989 ( .INP(n4371), .Z(n4010) );
  NBUFFX2 U3990 ( .INP(n4371), .Z(n4011) );
  NBUFFX2 U3992 ( .INP(n4370), .Z(n4012) );
  NBUFFX2 U3993 ( .INP(n4370), .Z(n4013) );
  NBUFFX2 U3994 ( .INP(n4370), .Z(n4014) );
  NBUFFX2 U3995 ( .INP(n4369), .Z(n4015) );
  NBUFFX2 U3996 ( .INP(n4369), .Z(n4016) );
  NBUFFX2 U3997 ( .INP(n4369), .Z(n4017) );
  NBUFFX2 U3998 ( .INP(n4368), .Z(n4018) );
  NBUFFX2 U3999 ( .INP(n4368), .Z(n4019) );
  NBUFFX2 U4000 ( .INP(n4368), .Z(n4020) );
  NBUFFX2 U4001 ( .INP(n4367), .Z(n4021) );
  NBUFFX2 U4002 ( .INP(n4367), .Z(n4022) );
  NBUFFX2 U4003 ( .INP(n4367), .Z(n4023) );
  NBUFFX2 U4004 ( .INP(n4366), .Z(n4024) );
  NBUFFX2 U4005 ( .INP(n4366), .Z(n4025) );
  NBUFFX2 U4006 ( .INP(n4366), .Z(n4026) );
  NBUFFX2 U4007 ( .INP(n4365), .Z(n4027) );
  NBUFFX2 U4008 ( .INP(n4365), .Z(n4028) );
  NBUFFX2 U4009 ( .INP(n4365), .Z(n4029) );
  NBUFFX2 U4010 ( .INP(n4364), .Z(n4030) );
  NBUFFX2 U4011 ( .INP(n4364), .Z(n4031) );
  NBUFFX2 U4012 ( .INP(n4364), .Z(n4032) );
  NBUFFX2 U4013 ( .INP(n4363), .Z(n4033) );
  NBUFFX2 U4014 ( .INP(n4363), .Z(n4034) );
  NBUFFX2 U4015 ( .INP(n4363), .Z(n4035) );
  NBUFFX2 U4016 ( .INP(n4362), .Z(n4036) );
  NBUFFX2 U4017 ( .INP(n4362), .Z(n4037) );
  NBUFFX2 U4018 ( .INP(n4362), .Z(n4038) );
  NBUFFX2 U4019 ( .INP(n4361), .Z(n4039) );
  NBUFFX2 U4020 ( .INP(n4361), .Z(n4040) );
  NBUFFX2 U4021 ( .INP(n4361), .Z(n4041) );
  NBUFFX2 U4022 ( .INP(n4360), .Z(n4042) );
  NBUFFX2 U4023 ( .INP(n4360), .Z(n4043) );
  NBUFFX2 U4024 ( .INP(n4360), .Z(n4044) );
  NBUFFX2 U4025 ( .INP(n4359), .Z(n4045) );
  NBUFFX2 U4026 ( .INP(n4359), .Z(n4046) );
  NBUFFX2 U4027 ( .INP(n4359), .Z(n4047) );
  NBUFFX2 U4028 ( .INP(n4358), .Z(n4048) );
  NBUFFX2 U4029 ( .INP(n4358), .Z(n4049) );
  NBUFFX2 U4030 ( .INP(n4358), .Z(n4050) );
  NBUFFX2 U4031 ( .INP(n4357), .Z(n4051) );
  NBUFFX2 U4032 ( .INP(n4357), .Z(n4052) );
  NBUFFX2 U4033 ( .INP(n4357), .Z(n4053) );
  NBUFFX2 U4034 ( .INP(n4356), .Z(n4054) );
  NBUFFX2 U4035 ( .INP(n4356), .Z(n4055) );
  NBUFFX2 U4036 ( .INP(n4356), .Z(n4056) );
  NBUFFX2 U4037 ( .INP(n4355), .Z(n4057) );
  NBUFFX2 U4038 ( .INP(n4355), .Z(n4058) );
  NBUFFX2 U4039 ( .INP(n4355), .Z(n4059) );
  NBUFFX2 U4040 ( .INP(n4354), .Z(n4060) );
  NBUFFX2 U4041 ( .INP(n4354), .Z(n4061) );
  NBUFFX2 U4042 ( .INP(n4354), .Z(n4062) );
  NBUFFX2 U4043 ( .INP(n4353), .Z(n4063) );
  NBUFFX2 U4044 ( .INP(n4353), .Z(n4064) );
  NBUFFX2 U4045 ( .INP(n4353), .Z(n4065) );
  NBUFFX2 U4046 ( .INP(n4352), .Z(n4066) );
  NBUFFX2 U4047 ( .INP(n4352), .Z(n4067) );
  NBUFFX2 U4048 ( .INP(n4352), .Z(n4068) );
  NBUFFX2 U4049 ( .INP(n4351), .Z(n4069) );
  NBUFFX2 U4050 ( .INP(n4351), .Z(n4070) );
  NBUFFX2 U4051 ( .INP(n4351), .Z(n4071) );
  NBUFFX2 U4052 ( .INP(n4350), .Z(n4072) );
  NBUFFX2 U4053 ( .INP(n4350), .Z(n4073) );
  NBUFFX2 U4054 ( .INP(n4350), .Z(n4074) );
  NBUFFX2 U4055 ( .INP(n4349), .Z(n4075) );
  NBUFFX2 U4056 ( .INP(n4349), .Z(n4076) );
  NBUFFX2 U4057 ( .INP(n4349), .Z(n4077) );
  NBUFFX2 U4058 ( .INP(n4348), .Z(n4078) );
  NBUFFX2 U4059 ( .INP(n4348), .Z(n4079) );
  NBUFFX2 U4060 ( .INP(n4348), .Z(n4080) );
  NBUFFX2 U4061 ( .INP(n4347), .Z(n4081) );
  NBUFFX2 U4062 ( .INP(n4347), .Z(n4082) );
  NBUFFX2 U4063 ( .INP(n4347), .Z(n4083) );
  NBUFFX2 U4064 ( .INP(n4346), .Z(n4084) );
  NBUFFX2 U4065 ( .INP(n4346), .Z(n4085) );
  NBUFFX2 U4066 ( .INP(n4346), .Z(n4086) );
  NBUFFX2 U4067 ( .INP(n4345), .Z(n4087) );
  NBUFFX2 U4068 ( .INP(n4345), .Z(n4088) );
  NBUFFX2 U4069 ( .INP(n4345), .Z(n4089) );
  NBUFFX2 U4070 ( .INP(n4344), .Z(n4090) );
  NBUFFX2 U4071 ( .INP(n4344), .Z(n4091) );
  NBUFFX2 U4072 ( .INP(n4344), .Z(n4092) );
  NBUFFX2 U4073 ( .INP(n4343), .Z(n4093) );
  NBUFFX2 U4074 ( .INP(n4343), .Z(n4094) );
  NBUFFX2 U4075 ( .INP(n4343), .Z(n4095) );
  NBUFFX2 U4076 ( .INP(n4342), .Z(n4096) );
  NBUFFX2 U4077 ( .INP(n4342), .Z(n4097) );
  NBUFFX2 U4078 ( .INP(n4342), .Z(n4098) );
  NBUFFX2 U4079 ( .INP(n4341), .Z(n4099) );
  NBUFFX2 U4080 ( .INP(n4341), .Z(n4100) );
  NBUFFX2 U4081 ( .INP(n4341), .Z(n4101) );
  NBUFFX2 U4082 ( .INP(n4340), .Z(n4102) );
  NBUFFX2 U4083 ( .INP(n4340), .Z(n4103) );
  NBUFFX2 U4084 ( .INP(n4340), .Z(n4104) );
  NBUFFX2 U4085 ( .INP(n4339), .Z(n4105) );
  NBUFFX2 U4086 ( .INP(n4339), .Z(n4106) );
  NBUFFX2 U4087 ( .INP(n4339), .Z(n4107) );
  NBUFFX2 U4088 ( .INP(n4338), .Z(n4108) );
  NBUFFX2 U4089 ( .INP(n4338), .Z(n4109) );
  NBUFFX2 U4090 ( .INP(n4338), .Z(n4110) );
  NBUFFX2 U4091 ( .INP(n4337), .Z(n4111) );
  NBUFFX2 U4092 ( .INP(n4337), .Z(n4112) );
  NBUFFX2 U4093 ( .INP(n4337), .Z(n4113) );
  NBUFFX2 U4094 ( .INP(n4336), .Z(n4114) );
  NBUFFX2 U4095 ( .INP(n4336), .Z(n4115) );
  NBUFFX2 U4096 ( .INP(n4336), .Z(n4116) );
  NBUFFX2 U4097 ( .INP(n4335), .Z(n4117) );
  NBUFFX2 U4098 ( .INP(n4335), .Z(n4118) );
  NBUFFX2 U4099 ( .INP(n4335), .Z(n4119) );
  NBUFFX2 U4100 ( .INP(n4334), .Z(n4120) );
  NBUFFX2 U4101 ( .INP(n4334), .Z(n4121) );
  NBUFFX2 U4102 ( .INP(n4334), .Z(n4122) );
  NBUFFX2 U4103 ( .INP(n4333), .Z(n4123) );
  NBUFFX2 U4104 ( .INP(n4333), .Z(n4124) );
  NBUFFX2 U4105 ( .INP(n4333), .Z(n4125) );
  NBUFFX2 U4106 ( .INP(n4332), .Z(n4126) );
  NBUFFX2 U4107 ( .INP(n4332), .Z(n4127) );
  NBUFFX2 U4108 ( .INP(n4332), .Z(n4128) );
  NBUFFX2 U4109 ( .INP(n4331), .Z(n4129) );
  NBUFFX2 U4110 ( .INP(n4331), .Z(n4130) );
  NBUFFX2 U4111 ( .INP(n4331), .Z(n4131) );
  NBUFFX2 U4112 ( .INP(n4330), .Z(n4132) );
  NBUFFX2 U4113 ( .INP(n4330), .Z(n4133) );
  NBUFFX2 U4114 ( .INP(n4330), .Z(n4134) );
  NBUFFX2 U4115 ( .INP(n4329), .Z(n4135) );
  NBUFFX2 U4116 ( .INP(n4329), .Z(n4136) );
  NBUFFX2 U4117 ( .INP(n4329), .Z(n4137) );
  NBUFFX2 U4118 ( .INP(n4328), .Z(n4138) );
  NBUFFX2 U4119 ( .INP(n4328), .Z(n4139) );
  NBUFFX2 U4120 ( .INP(n4328), .Z(n4140) );
  NBUFFX2 U4121 ( .INP(n4327), .Z(n4141) );
  NBUFFX2 U4122 ( .INP(n4327), .Z(n4142) );
  NBUFFX2 U4123 ( .INP(n4327), .Z(n4143) );
  NBUFFX2 U4124 ( .INP(n4326), .Z(n4144) );
  NBUFFX2 U4125 ( .INP(n4326), .Z(n4145) );
  NBUFFX2 U4126 ( .INP(n4326), .Z(n4146) );
  NBUFFX2 U4127 ( .INP(n4325), .Z(n4147) );
  NBUFFX2 U4128 ( .INP(n4325), .Z(n4148) );
  NBUFFX2 U4129 ( .INP(n4325), .Z(n4149) );
  NBUFFX2 U4130 ( .INP(n4324), .Z(n4150) );
  NBUFFX2 U4131 ( .INP(n4324), .Z(n4151) );
  NBUFFX2 U4132 ( .INP(n4324), .Z(n4152) );
  NBUFFX2 U4133 ( .INP(n4323), .Z(n4153) );
  NBUFFX2 U4134 ( .INP(n4323), .Z(n4154) );
  NBUFFX2 U4135 ( .INP(n4323), .Z(n4155) );
  NBUFFX2 U4136 ( .INP(n4322), .Z(n4156) );
  NBUFFX2 U4137 ( .INP(n4322), .Z(n4157) );
  NBUFFX2 U4138 ( .INP(n4322), .Z(n4158) );
  NBUFFX2 U4139 ( .INP(n4321), .Z(n4159) );
  NBUFFX2 U4140 ( .INP(n4321), .Z(n4160) );
  NBUFFX2 U4141 ( .INP(n4321), .Z(n4161) );
  NBUFFX2 U4142 ( .INP(n4320), .Z(n4162) );
  NBUFFX2 U4143 ( .INP(n4320), .Z(n4163) );
  NBUFFX2 U4144 ( .INP(n4320), .Z(n4164) );
  NBUFFX2 U4145 ( .INP(n4319), .Z(n4165) );
  NBUFFX2 U4146 ( .INP(n4319), .Z(n4166) );
  NBUFFX2 U4147 ( .INP(n4319), .Z(n4167) );
  NBUFFX2 U4148 ( .INP(n4318), .Z(n4168) );
  NBUFFX2 U4149 ( .INP(n4318), .Z(n4169) );
  NBUFFX2 U4150 ( .INP(n4318), .Z(n4170) );
  NBUFFX2 U4151 ( .INP(n4317), .Z(n4171) );
  NBUFFX2 U4152 ( .INP(n4317), .Z(n4172) );
  NBUFFX2 U4153 ( .INP(n4317), .Z(n4173) );
  NBUFFX2 U4154 ( .INP(n4316), .Z(n4174) );
  NBUFFX2 U4155 ( .INP(n4316), .Z(n4175) );
  NBUFFX2 U4156 ( .INP(n4316), .Z(n4176) );
  NBUFFX2 U4157 ( .INP(n4315), .Z(n4177) );
  NBUFFX2 U4158 ( .INP(n4315), .Z(n4178) );
  NBUFFX2 U4159 ( .INP(n4315), .Z(n4179) );
  NBUFFX2 U4160 ( .INP(n4314), .Z(n4180) );
  NBUFFX2 U4161 ( .INP(n4314), .Z(n4181) );
  NBUFFX2 U4162 ( .INP(n4314), .Z(n4182) );
  NBUFFX2 U4163 ( .INP(n4313), .Z(n4183) );
  NBUFFX2 U4164 ( .INP(n4313), .Z(n4184) );
  NBUFFX2 U4165 ( .INP(n4313), .Z(n4185) );
  NBUFFX2 U4166 ( .INP(n4312), .Z(n4186) );
  NBUFFX2 U4167 ( .INP(n4312), .Z(n4187) );
  NBUFFX2 U4168 ( .INP(n4312), .Z(n4188) );
  NBUFFX2 U4169 ( .INP(n4311), .Z(n4189) );
  NBUFFX2 U4170 ( .INP(n4311), .Z(n4190) );
  NBUFFX2 U4171 ( .INP(n4311), .Z(n4191) );
  NBUFFX2 U4172 ( .INP(n4310), .Z(n4192) );
  NBUFFX2 U4173 ( .INP(n4310), .Z(n4193) );
  NBUFFX2 U4174 ( .INP(n4310), .Z(n4194) );
  NBUFFX2 U4175 ( .INP(n4309), .Z(n4195) );
  NBUFFX2 U4176 ( .INP(n4309), .Z(n4196) );
  NBUFFX2 U4177 ( .INP(n4309), .Z(n4197) );
  NBUFFX2 U4178 ( .INP(n4308), .Z(n4198) );
  NBUFFX2 U4179 ( .INP(n4308), .Z(n4199) );
  NBUFFX2 U4180 ( .INP(n4308), .Z(n4200) );
  NBUFFX2 U4181 ( .INP(n4307), .Z(n4201) );
  NBUFFX2 U4182 ( .INP(n4307), .Z(n4202) );
  NBUFFX2 U4183 ( .INP(n4307), .Z(n4203) );
  NBUFFX2 U4184 ( .INP(n4306), .Z(n4204) );
  NBUFFX2 U4185 ( .INP(n4306), .Z(n4205) );
  NBUFFX2 U4186 ( .INP(n4306), .Z(n4206) );
  NBUFFX2 U4187 ( .INP(n4305), .Z(n4207) );
  NBUFFX2 U4188 ( .INP(n4305), .Z(n4208) );
  NBUFFX2 U4189 ( .INP(n4305), .Z(n4209) );
  NBUFFX2 U4190 ( .INP(n4304), .Z(n4210) );
  NBUFFX2 U4191 ( .INP(n4304), .Z(n4211) );
  NBUFFX2 U4192 ( .INP(n4304), .Z(n4212) );
  NBUFFX2 U4193 ( .INP(n4303), .Z(n4213) );
  NBUFFX2 U4194 ( .INP(n4303), .Z(n4214) );
  NBUFFX2 U4195 ( .INP(n4303), .Z(n4215) );
  NBUFFX2 U4196 ( .INP(n4302), .Z(n4216) );
  NBUFFX2 U4197 ( .INP(n4302), .Z(n4217) );
  NBUFFX2 U4198 ( .INP(n4302), .Z(n4218) );
  NBUFFX2 U4199 ( .INP(n4301), .Z(n4219) );
  NBUFFX2 U4200 ( .INP(n4301), .Z(n4220) );
  NBUFFX2 U4201 ( .INP(n4301), .Z(n4221) );
  NBUFFX2 U4202 ( .INP(n4300), .Z(n4222) );
  NBUFFX2 U4203 ( .INP(n4300), .Z(n4223) );
  NBUFFX2 U4204 ( .INP(n4300), .Z(n4224) );
  NBUFFX2 U4205 ( .INP(n4299), .Z(n4225) );
  NBUFFX2 U4206 ( .INP(n4299), .Z(n4226) );
  NBUFFX2 U4207 ( .INP(n4299), .Z(n4227) );
  NBUFFX2 U4208 ( .INP(n4298), .Z(n4228) );
  NBUFFX2 U4209 ( .INP(n4298), .Z(n4229) );
  NBUFFX2 U4210 ( .INP(n4298), .Z(n4230) );
  NBUFFX2 U4211 ( .INP(n4297), .Z(n4231) );
  NBUFFX2 U4212 ( .INP(n4297), .Z(n4232) );
  NBUFFX2 U4213 ( .INP(n4297), .Z(n4233) );
  NBUFFX2 U4214 ( .INP(n4296), .Z(n4234) );
  NBUFFX2 U4215 ( .INP(n4296), .Z(n4235) );
  NBUFFX2 U4216 ( .INP(n4296), .Z(n4236) );
  NBUFFX2 U4217 ( .INP(n4295), .Z(n4237) );
  NBUFFX2 U4218 ( .INP(n4295), .Z(n4238) );
  NBUFFX2 U4219 ( .INP(n4295), .Z(n4239) );
  NBUFFX2 U4220 ( .INP(n4294), .Z(n4240) );
  NBUFFX2 U4221 ( .INP(n4294), .Z(n4241) );
  NBUFFX2 U4222 ( .INP(n4294), .Z(n4242) );
  NBUFFX2 U4223 ( .INP(n4293), .Z(n4243) );
  NBUFFX2 U4224 ( .INP(n4293), .Z(n4244) );
  NBUFFX2 U4225 ( .INP(n4293), .Z(n4245) );
  NBUFFX2 U4226 ( .INP(n4292), .Z(n4246) );
  NBUFFX2 U4227 ( .INP(n4292), .Z(n4247) );
  NBUFFX2 U4228 ( .INP(n4292), .Z(n4248) );
  NBUFFX2 U4229 ( .INP(n4291), .Z(n4249) );
  NBUFFX2 U4230 ( .INP(n4291), .Z(n4250) );
  NBUFFX2 U4231 ( .INP(n4291), .Z(n4251) );
  NBUFFX2 U4232 ( .INP(n4290), .Z(n4252) );
  NBUFFX2 U4233 ( .INP(n4290), .Z(n4253) );
  NBUFFX2 U4234 ( .INP(n4290), .Z(n4254) );
  NBUFFX2 U4235 ( .INP(n4289), .Z(n4255) );
  NBUFFX2 U4236 ( .INP(n4289), .Z(n4256) );
  NBUFFX2 U4237 ( .INP(n4289), .Z(n4257) );
  NBUFFX2 U4238 ( .INP(n4288), .Z(n4258) );
  NBUFFX2 U4239 ( .INP(n4288), .Z(n4259) );
  NBUFFX2 U4240 ( .INP(n4288), .Z(n4260) );
  NBUFFX2 U4241 ( .INP(n4287), .Z(n4261) );
  NBUFFX2 U4242 ( .INP(n4287), .Z(n4262) );
  NBUFFX2 U4243 ( .INP(n4287), .Z(n4263) );
  NBUFFX2 U4244 ( .INP(n4286), .Z(n4264) );
  NBUFFX2 U4245 ( .INP(n4286), .Z(n4265) );
  NBUFFX2 U4246 ( .INP(n4286), .Z(n4266) );
  NBUFFX2 U4247 ( .INP(n4285), .Z(n4267) );
  NBUFFX2 U4248 ( .INP(n4285), .Z(n4268) );
  NBUFFX2 U4249 ( .INP(n4285), .Z(n4269) );
  NBUFFX2 U4250 ( .INP(n4284), .Z(n4270) );
  NBUFFX2 U4251 ( .INP(n4284), .Z(n4271) );
  NBUFFX2 U4252 ( .INP(n4284), .Z(n4272) );
  NBUFFX2 U4253 ( .INP(n4283), .Z(n4273) );
  NBUFFX2 U4254 ( .INP(n4283), .Z(n4274) );
  NBUFFX2 U4255 ( .INP(n4283), .Z(n4275) );
  NBUFFX2 U4256 ( .INP(n4282), .Z(n4276) );
  NBUFFX2 U4257 ( .INP(n4282), .Z(n4277) );
  NBUFFX2 U4258 ( .INP(n4282), .Z(n4278) );
  NBUFFX2 U4259 ( .INP(n4281), .Z(n4279) );
  NBUFFX2 U4260 ( .INP(n4281), .Z(n4280) );
  NBUFFX2 U4261 ( .INP(n4410), .Z(n4281) );
  NBUFFX2 U4262 ( .INP(n4409), .Z(n4282) );
  NBUFFX2 U4263 ( .INP(n4409), .Z(n4283) );
  NBUFFX2 U4264 ( .INP(n4409), .Z(n4284) );
  NBUFFX2 U4265 ( .INP(n4408), .Z(n4285) );
  NBUFFX2 U4266 ( .INP(n4408), .Z(n4286) );
  NBUFFX2 U4267 ( .INP(n4408), .Z(n4287) );
  NBUFFX2 U4268 ( .INP(n4407), .Z(n4288) );
  NBUFFX2 U4269 ( .INP(n4407), .Z(n4289) );
  NBUFFX2 U4270 ( .INP(n4407), .Z(n4290) );
  NBUFFX2 U4271 ( .INP(n4406), .Z(n4291) );
  NBUFFX2 U4272 ( .INP(n4406), .Z(n4292) );
  NBUFFX2 U4273 ( .INP(n4406), .Z(n4293) );
  NBUFFX2 U4274 ( .INP(n4405), .Z(n4294) );
  NBUFFX2 U4275 ( .INP(n4405), .Z(n4295) );
  NBUFFX2 U4276 ( .INP(n4405), .Z(n4296) );
  NBUFFX2 U4277 ( .INP(n4404), .Z(n4297) );
  NBUFFX2 U4278 ( .INP(n4404), .Z(n4298) );
  NBUFFX2 U4279 ( .INP(n4404), .Z(n4299) );
  NBUFFX2 U4280 ( .INP(n4403), .Z(n4300) );
  NBUFFX2 U4281 ( .INP(n4403), .Z(n4301) );
  NBUFFX2 U4282 ( .INP(n4403), .Z(n4302) );
  NBUFFX2 U4283 ( .INP(n4402), .Z(n4303) );
  NBUFFX2 U4284 ( .INP(n4402), .Z(n4304) );
  NBUFFX2 U4285 ( .INP(n4402), .Z(n4305) );
  NBUFFX2 U4286 ( .INP(n4401), .Z(n4306) );
  NBUFFX2 U4287 ( .INP(n4401), .Z(n4307) );
  NBUFFX2 U4288 ( .INP(n4401), .Z(n4308) );
  NBUFFX2 U4289 ( .INP(n4400), .Z(n4309) );
  NBUFFX2 U4290 ( .INP(n4400), .Z(n4310) );
  NBUFFX2 U4291 ( .INP(n4400), .Z(n4311) );
  NBUFFX2 U4292 ( .INP(n4399), .Z(n4312) );
  NBUFFX2 U4293 ( .INP(n4399), .Z(n4313) );
  NBUFFX2 U4294 ( .INP(n4399), .Z(n4314) );
  NBUFFX2 U4295 ( .INP(n4398), .Z(n4315) );
  NBUFFX2 U4296 ( .INP(n4398), .Z(n4316) );
  NBUFFX2 U4297 ( .INP(n4398), .Z(n4317) );
  NBUFFX2 U4298 ( .INP(n4397), .Z(n4318) );
  NBUFFX2 U4299 ( .INP(n4397), .Z(n4319) );
  NBUFFX2 U4300 ( .INP(n4397), .Z(n4320) );
  NBUFFX2 U4301 ( .INP(n4396), .Z(n4321) );
  NBUFFX2 U4302 ( .INP(n4396), .Z(n4322) );
  NBUFFX2 U4303 ( .INP(n4396), .Z(n4323) );
  NBUFFX2 U4304 ( .INP(n4395), .Z(n4324) );
  NBUFFX2 U4305 ( .INP(n4395), .Z(n4325) );
  NBUFFX2 U4306 ( .INP(n4395), .Z(n4326) );
  NBUFFX2 U4307 ( .INP(n4394), .Z(n4327) );
  NBUFFX2 U4308 ( .INP(n4394), .Z(n4328) );
  NBUFFX2 U4309 ( .INP(n4394), .Z(n4329) );
  NBUFFX2 U4310 ( .INP(n4393), .Z(n4330) );
  NBUFFX2 U4311 ( .INP(n4393), .Z(n4331) );
  NBUFFX2 U4312 ( .INP(n4393), .Z(n4332) );
  NBUFFX2 U4313 ( .INP(n4392), .Z(n4333) );
  NBUFFX2 U4314 ( .INP(n4392), .Z(n4334) );
  NBUFFX2 U4315 ( .INP(n4392), .Z(n4335) );
  NBUFFX2 U4316 ( .INP(n4391), .Z(n4336) );
  NBUFFX2 U4317 ( .INP(n4391), .Z(n4337) );
  NBUFFX2 U4318 ( .INP(n4391), .Z(n4338) );
  NBUFFX2 U4319 ( .INP(n4390), .Z(n4339) );
  NBUFFX2 U4320 ( .INP(n4390), .Z(n4340) );
  NBUFFX2 U4321 ( .INP(n4390), .Z(n4341) );
  NBUFFX2 U4322 ( .INP(n4389), .Z(n4342) );
  NBUFFX2 U4323 ( .INP(n4389), .Z(n4343) );
  NBUFFX2 U4324 ( .INP(n4389), .Z(n4344) );
  NBUFFX2 U4325 ( .INP(n4388), .Z(n4345) );
  NBUFFX2 U4326 ( .INP(n4388), .Z(n4346) );
  NBUFFX2 U4327 ( .INP(n4388), .Z(n4347) );
  NBUFFX2 U4328 ( .INP(n4387), .Z(n4348) );
  NBUFFX2 U4329 ( .INP(n4387), .Z(n4349) );
  NBUFFX2 U4330 ( .INP(n4387), .Z(n4350) );
  NBUFFX2 U4331 ( .INP(n4386), .Z(n4351) );
  NBUFFX2 U4332 ( .INP(n4386), .Z(n4352) );
  NBUFFX2 U4333 ( .INP(n4386), .Z(n4353) );
  NBUFFX2 U4334 ( .INP(n4385), .Z(n4354) );
  NBUFFX2 U4335 ( .INP(n4385), .Z(n4355) );
  NBUFFX2 U4336 ( .INP(n4385), .Z(n4356) );
  NBUFFX2 U4337 ( .INP(n4384), .Z(n4357) );
  NBUFFX2 U4338 ( .INP(n4384), .Z(n4358) );
  NBUFFX2 U4339 ( .INP(n4384), .Z(n4359) );
  NBUFFX2 U4340 ( .INP(n4383), .Z(n4360) );
  NBUFFX2 U4341 ( .INP(n4383), .Z(n4361) );
  NBUFFX2 U4342 ( .INP(n4383), .Z(n4362) );
  NBUFFX2 U4343 ( .INP(n4382), .Z(n4363) );
  NBUFFX2 U4344 ( .INP(n4382), .Z(n4364) );
  NBUFFX2 U4345 ( .INP(n4382), .Z(n4365) );
  NBUFFX2 U4346 ( .INP(n4381), .Z(n4366) );
  NBUFFX2 U4347 ( .INP(n4381), .Z(n4367) );
  NBUFFX2 U4348 ( .INP(n4381), .Z(n4368) );
  NBUFFX2 U4349 ( .INP(n4380), .Z(n4369) );
  NBUFFX2 U4350 ( .INP(n4380), .Z(n4370) );
  NBUFFX2 U4351 ( .INP(n4380), .Z(n4371) );
  NBUFFX2 U4352 ( .INP(n4379), .Z(n4372) );
  NBUFFX2 U4353 ( .INP(n4379), .Z(n4373) );
  NBUFFX2 U4354 ( .INP(n4379), .Z(n4374) );
  NBUFFX2 U4355 ( .INP(n4378), .Z(n4375) );
  NBUFFX2 U4356 ( .INP(n4378), .Z(n4376) );
  NBUFFX2 U4357 ( .INP(n4378), .Z(n4377) );
  NBUFFX2 U4358 ( .INP(n4421), .Z(n4378) );
  NBUFFX2 U4359 ( .INP(n4421), .Z(n4379) );
  NBUFFX2 U4360 ( .INP(n4421), .Z(n4380) );
  NBUFFX2 U4361 ( .INP(n4420), .Z(n4381) );
  NBUFFX2 U4362 ( .INP(n4420), .Z(n4382) );
  NBUFFX2 U4363 ( .INP(n4420), .Z(n4383) );
  NBUFFX2 U4364 ( .INP(n4419), .Z(n4384) );
  NBUFFX2 U4365 ( .INP(n4419), .Z(n4385) );
  NBUFFX2 U4366 ( .INP(n4419), .Z(n4386) );
  NBUFFX2 U4367 ( .INP(n4418), .Z(n4387) );
  NBUFFX2 U4368 ( .INP(n4418), .Z(n4388) );
  NBUFFX2 U4369 ( .INP(n4418), .Z(n4389) );
  NBUFFX2 U4370 ( .INP(n4417), .Z(n4390) );
  NBUFFX2 U4371 ( .INP(n4417), .Z(n4391) );
  NBUFFX2 U4372 ( .INP(n4417), .Z(n4392) );
  NBUFFX2 U4373 ( .INP(n4416), .Z(n4393) );
  NBUFFX2 U4374 ( .INP(n4416), .Z(n4394) );
  NBUFFX2 U4375 ( .INP(n4416), .Z(n4395) );
  NBUFFX2 U4376 ( .INP(n4415), .Z(n4396) );
  NBUFFX2 U4377 ( .INP(n4415), .Z(n4397) );
  NBUFFX2 U4378 ( .INP(n4415), .Z(n4398) );
  NBUFFX2 U4379 ( .INP(n4414), .Z(n4399) );
  NBUFFX2 U4380 ( .INP(n4414), .Z(n4400) );
  NBUFFX2 U4381 ( .INP(n4414), .Z(n4401) );
  NBUFFX2 U4382 ( .INP(n4413), .Z(n4402) );
  NBUFFX2 U4383 ( .INP(n4413), .Z(n4403) );
  NBUFFX2 U4384 ( .INP(n4413), .Z(n4404) );
  NBUFFX2 U4385 ( .INP(n4412), .Z(n4405) );
  NBUFFX2 U4386 ( .INP(n4412), .Z(n4406) );
  NBUFFX2 U4387 ( .INP(n4412), .Z(n4407) );
  NBUFFX2 U4388 ( .INP(n4411), .Z(n4408) );
  NBUFFX2 U4389 ( .INP(n4411), .Z(n4409) );
  NBUFFX2 U4390 ( .INP(n4411), .Z(n4410) );
  NBUFFX2 U4391 ( .INP(n4425), .Z(n4411) );
  NBUFFX2 U4392 ( .INP(n4425), .Z(n4412) );
  NBUFFX2 U4393 ( .INP(n4424), .Z(n4413) );
  NBUFFX2 U4394 ( .INP(n4424), .Z(n4414) );
  NBUFFX2 U4395 ( .INP(n4424), .Z(n4415) );
  NBUFFX2 U4396 ( .INP(n4423), .Z(n4416) );
  NBUFFX2 U4397 ( .INP(n4423), .Z(n4417) );
  NBUFFX2 U4398 ( .INP(n4423), .Z(n4418) );
  NBUFFX2 U4399 ( .INP(n4422), .Z(n4419) );
  NBUFFX2 U4400 ( .INP(n4422), .Z(n4420) );
  NBUFFX2 U4401 ( .INP(n4422), .Z(n4421) );
  NBUFFX2 U4402 ( .INP(test_se), .Z(n4422) );
  NBUFFX2 U4403 ( .INP(test_se), .Z(n4423) );
  NBUFFX2 U4404 ( .INP(test_se), .Z(n4424) );
  NBUFFX2 U4405 ( .INP(test_se), .Z(n4425) );
  NBUFFX2 U4406 ( .INP(n4477), .Z(n4426) );
  NBUFFX2 U4407 ( .INP(n4477), .Z(n4427) );
  NBUFFX2 U4408 ( .INP(n4477), .Z(n4428) );
  NBUFFX2 U4409 ( .INP(n4476), .Z(n4429) );
  NBUFFX2 U4410 ( .INP(n4476), .Z(n4430) );
  NBUFFX2 U4411 ( .INP(n4476), .Z(n4431) );
  NBUFFX2 U4412 ( .INP(n4475), .Z(n4432) );
  NBUFFX2 U4413 ( .INP(n4475), .Z(n4433) );
  NBUFFX2 U4414 ( .INP(n4475), .Z(n4434) );
  NBUFFX2 U4415 ( .INP(n4474), .Z(n4435) );
  NBUFFX2 U4416 ( .INP(n4474), .Z(n4436) );
  NBUFFX2 U4417 ( .INP(n4474), .Z(n4437) );
  NBUFFX2 U4418 ( .INP(n4473), .Z(n4438) );
  NBUFFX2 U4419 ( .INP(n4473), .Z(n4439) );
  NBUFFX2 U4420 ( .INP(n4473), .Z(n4440) );
  NBUFFX2 U4421 ( .INP(n4472), .Z(n4441) );
  NBUFFX2 U4422 ( .INP(n4472), .Z(n4442) );
  NBUFFX2 U4423 ( .INP(n4472), .Z(n4443) );
  NBUFFX2 U4424 ( .INP(n4471), .Z(n4444) );
  NBUFFX2 U4425 ( .INP(n4471), .Z(n4445) );
  NBUFFX2 U4426 ( .INP(n4471), .Z(n4446) );
  NBUFFX2 U4427 ( .INP(n4470), .Z(n4447) );
  NBUFFX2 U4428 ( .INP(n4470), .Z(n4448) );
  NBUFFX2 U4429 ( .INP(n4470), .Z(n4449) );
  NBUFFX2 U4430 ( .INP(n4469), .Z(n4450) );
  NBUFFX2 U4431 ( .INP(n4469), .Z(n4451) );
  NBUFFX2 U4432 ( .INP(n4469), .Z(n4452) );
  NBUFFX2 U4433 ( .INP(n4468), .Z(n4453) );
  NBUFFX2 U4434 ( .INP(n4468), .Z(n4454) );
  NBUFFX2 U4435 ( .INP(n4468), .Z(n4455) );
  NBUFFX2 U4436 ( .INP(n4467), .Z(n4456) );
  NBUFFX2 U4437 ( .INP(n4467), .Z(n4457) );
  NBUFFX2 U4438 ( .INP(n4467), .Z(n4458) );
  NBUFFX2 U4439 ( .INP(n4466), .Z(n4459) );
  NBUFFX2 U4440 ( .INP(n4466), .Z(n4460) );
  NBUFFX2 U4441 ( .INP(n4466), .Z(n4461) );
  NBUFFX2 U4442 ( .INP(n4465), .Z(n4462) );
  NBUFFX2 U4443 ( .INP(n4465), .Z(n4463) );
  NBUFFX2 U4444 ( .INP(n4465), .Z(n4464) );
  NBUFFX2 U4445 ( .INP(n4482), .Z(n4465) );
  NBUFFX2 U4446 ( .INP(n4481), .Z(n4466) );
  NBUFFX2 U4447 ( .INP(n4481), .Z(n4467) );
  NBUFFX2 U4448 ( .INP(n4481), .Z(n4468) );
  NBUFFX2 U4449 ( .INP(n4480), .Z(n4469) );
  NBUFFX2 U4450 ( .INP(n4480), .Z(n4470) );
  NBUFFX2 U4451 ( .INP(n4480), .Z(n4471) );
  NBUFFX2 U4452 ( .INP(n4479), .Z(n4472) );
  NBUFFX2 U4453 ( .INP(n4479), .Z(n4473) );
  NBUFFX2 U4454 ( .INP(n4479), .Z(n4474) );
  NBUFFX2 U4455 ( .INP(n4478), .Z(n4475) );
  NBUFFX2 U4456 ( .INP(n4478), .Z(n4476) );
  NBUFFX2 U4457 ( .INP(n4478), .Z(n4477) );
  NBUFFX2 U4458 ( .INP(RESET), .Z(n4478) );
  NBUFFX2 U4459 ( .INP(RESET), .Z(n4479) );
  NBUFFX2 U4460 ( .INP(RESET), .Z(n4480) );
  NBUFFX2 U4461 ( .INP(RESET), .Z(n4481) );
  NBUFFX2 U4462 ( .INP(RESET), .Z(n4482) );
  INVX0 U4463 ( .INP(n4426), .ZN(n4483) );
  INVX0 U4464 ( .INP(n4426), .ZN(n4484) );
  INVX0 U4465 ( .INP(n4426), .ZN(n4485) );
  INVX0 U4466 ( .INP(n4426), .ZN(n4486) );
  INVX0 U4467 ( .INP(n4426), .ZN(n4487) );
  INVX0 U4468 ( .INP(n4426), .ZN(n4488) );
  INVX0 U4469 ( .INP(n4426), .ZN(n4489) );
  INVX0 U4470 ( .INP(n4426), .ZN(n4490) );
  INVX0 U4471 ( .INP(n4427), .ZN(n4491) );
  INVX0 U4472 ( .INP(n4427), .ZN(n4492) );
  INVX0 U4473 ( .INP(n4427), .ZN(n4493) );
  INVX0 U4474 ( .INP(n4427), .ZN(n4494) );
  INVX0 U4475 ( .INP(n4427), .ZN(n4495) );
  INVX0 U4476 ( .INP(n4427), .ZN(n4496) );
  INVX0 U4477 ( .INP(n4427), .ZN(n4497) );
  INVX0 U4478 ( .INP(n4427), .ZN(n4498) );
  INVX0 U4479 ( .INP(n4428), .ZN(n4499) );
  INVX0 U4480 ( .INP(n4428), .ZN(n4500) );
  INVX0 U4481 ( .INP(n4428), .ZN(n4501) );
  INVX0 U4482 ( .INP(n4428), .ZN(n4502) );
  INVX0 U4483 ( .INP(n4428), .ZN(n4503) );
  INVX0 U4484 ( .INP(n4428), .ZN(n4504) );
  INVX0 U4485 ( .INP(n4428), .ZN(n4505) );
  INVX0 U4486 ( .INP(n4428), .ZN(n4506) );
  INVX0 U4487 ( .INP(n4429), .ZN(n4507) );
  INVX0 U4488 ( .INP(n4429), .ZN(n4508) );
  INVX0 U4489 ( .INP(n4429), .ZN(n4509) );
  INVX0 U4490 ( .INP(n4429), .ZN(n4510) );
  INVX0 U4491 ( .INP(n4429), .ZN(n4511) );
  INVX0 U4492 ( .INP(n4429), .ZN(n4512) );
  INVX0 U4493 ( .INP(n4429), .ZN(n4513) );
  INVX0 U4494 ( .INP(n4429), .ZN(n4514) );
  INVX0 U4495 ( .INP(n4430), .ZN(n4515) );
  INVX0 U4496 ( .INP(n4430), .ZN(n4516) );
  INVX0 U4497 ( .INP(n4430), .ZN(n4517) );
  INVX0 U4498 ( .INP(n4430), .ZN(n4518) );
  INVX0 U4499 ( .INP(n4430), .ZN(n4519) );
  INVX0 U4500 ( .INP(n4430), .ZN(n4520) );
  INVX0 U4501 ( .INP(n4430), .ZN(n4521) );
  INVX0 U4502 ( .INP(n4430), .ZN(n4522) );
  INVX0 U4503 ( .INP(n4431), .ZN(n4523) );
  INVX0 U4504 ( .INP(n4431), .ZN(n4524) );
  INVX0 U4505 ( .INP(n4431), .ZN(n4525) );
  INVX0 U4506 ( .INP(n4431), .ZN(n4526) );
  INVX0 U4507 ( .INP(n4431), .ZN(n4527) );
  INVX0 U4508 ( .INP(n4431), .ZN(n4528) );
  INVX0 U4509 ( .INP(n4431), .ZN(n4529) );
  INVX0 U4510 ( .INP(n4432), .ZN(n4530) );
  INVX0 U4511 ( .INP(n4432), .ZN(n4531) );
  INVX0 U4512 ( .INP(n4432), .ZN(n4532) );
  INVX0 U4513 ( .INP(n4432), .ZN(n4533) );
  INVX0 U4514 ( .INP(n4432), .ZN(n4534) );
  INVX0 U4515 ( .INP(n4432), .ZN(n4535) );
  INVX0 U4516 ( .INP(n4432), .ZN(n4536) );
  INVX0 U4517 ( .INP(n4432), .ZN(n4537) );
  INVX0 U4518 ( .INP(n4433), .ZN(n4538) );
  INVX0 U4519 ( .INP(n4433), .ZN(n4539) );
  INVX0 U4520 ( .INP(n4433), .ZN(n4540) );
  INVX0 U4521 ( .INP(n4433), .ZN(n4541) );
  INVX0 U4522 ( .INP(n4433), .ZN(n4542) );
  INVX0 U4523 ( .INP(n4433), .ZN(n4543) );
  INVX0 U4524 ( .INP(n4433), .ZN(n4544) );
  INVX0 U4525 ( .INP(n4433), .ZN(n4545) );
  INVX0 U4526 ( .INP(n4434), .ZN(n4546) );
  INVX0 U4527 ( .INP(n4434), .ZN(n4547) );
  INVX0 U4528 ( .INP(n4434), .ZN(n4548) );
  INVX0 U4529 ( .INP(n4434), .ZN(n4549) );
  INVX0 U4530 ( .INP(n4434), .ZN(n4550) );
  INVX0 U4531 ( .INP(n4434), .ZN(n4551) );
  INVX0 U4532 ( .INP(n4434), .ZN(n4552) );
  INVX0 U4533 ( .INP(n4434), .ZN(n4553) );
  INVX0 U4534 ( .INP(n4435), .ZN(n4554) );
  INVX0 U4535 ( .INP(n4435), .ZN(n4555) );
  INVX0 U4536 ( .INP(n4435), .ZN(n4556) );
  INVX0 U4537 ( .INP(n4435), .ZN(n4557) );
  INVX0 U4538 ( .INP(n4435), .ZN(n4558) );
  INVX0 U4539 ( .INP(n4435), .ZN(n4559) );
  INVX0 U4540 ( .INP(n4435), .ZN(n4560) );
  INVX0 U4541 ( .INP(n4435), .ZN(n4561) );
  INVX0 U4542 ( .INP(n4436), .ZN(n4562) );
  INVX0 U4543 ( .INP(n4436), .ZN(n4563) );
  INVX0 U4544 ( .INP(n4436), .ZN(n4564) );
  INVX0 U4545 ( .INP(n4436), .ZN(n4565) );
  INVX0 U4546 ( .INP(n4436), .ZN(n4566) );
  INVX0 U4547 ( .INP(n4436), .ZN(n4567) );
  INVX0 U4548 ( .INP(n4431), .ZN(n4568) );
  NBUFFX2 U4549 ( .INP(n4751), .Z(n4713) );
  NBUFFX2 U4550 ( .INP(n4751), .Z(n4714) );
  NBUFFX2 U4551 ( .INP(n4750), .Z(n4715) );
  NBUFFX2 U4552 ( .INP(n4750), .Z(n4716) );
  NBUFFX2 U4553 ( .INP(n4750), .Z(n4717) );
  NBUFFX2 U4554 ( .INP(n4749), .Z(n4718) );
  NBUFFX2 U4555 ( .INP(n4749), .Z(n4719) );
  NBUFFX2 U4556 ( .INP(n4749), .Z(n4720) );
  NBUFFX2 U4557 ( .INP(n4748), .Z(n4721) );
  NBUFFX2 U4558 ( .INP(n4748), .Z(n4722) );
  NBUFFX2 U4559 ( .INP(n4748), .Z(n4723) );
  NBUFFX2 U4560 ( .INP(n4747), .Z(n4724) );
  NBUFFX2 U4561 ( .INP(n4747), .Z(n4725) );
  NBUFFX2 U4562 ( .INP(n4747), .Z(n4726) );
  NBUFFX2 U4563 ( .INP(n4746), .Z(n4727) );
  NBUFFX2 U4564 ( .INP(n4746), .Z(n4728) );
  NBUFFX2 U4565 ( .INP(n4746), .Z(n4729) );
  NBUFFX2 U4566 ( .INP(n4745), .Z(n4730) );
  NBUFFX2 U4567 ( .INP(n4745), .Z(n4731) );
  NBUFFX2 U4568 ( .INP(n4745), .Z(n4732) );
  NBUFFX2 U4569 ( .INP(n4744), .Z(n4733) );
  NBUFFX2 U4570 ( .INP(n4744), .Z(n4734) );
  NBUFFX2 U4571 ( .INP(n4744), .Z(n4735) );
  NBUFFX2 U4572 ( .INP(n4743), .Z(n4736) );
  NBUFFX2 U4573 ( .INP(n4743), .Z(n4737) );
  NBUFFX2 U4574 ( .INP(n4743), .Z(n4738) );
  NBUFFX2 U4575 ( .INP(n4742), .Z(n4739) );
  NBUFFX2 U4576 ( .INP(n4742), .Z(n4740) );
  NBUFFX2 U4577 ( .INP(n4742), .Z(n4741) );
  NBUFFX2 U4578 ( .INP(CK), .Z(n4742) );
  NBUFFX2 U4579 ( .INP(CK), .Z(n4743) );
  NBUFFX2 U4580 ( .INP(n4751), .Z(n4744) );
  NBUFFX2 U4581 ( .INP(CK), .Z(n4745) );
  NBUFFX2 U4582 ( .INP(n4747), .Z(n4746) );
  NBUFFX2 U4583 ( .INP(CK), .Z(n4747) );
  NBUFFX2 U4584 ( .INP(n4742), .Z(n4748) );
  NBUFFX2 U4585 ( .INP(n4743), .Z(n4749) );
  NBUFFX2 U4586 ( .INP(n4745), .Z(n4750) );
  NBUFFX2 U4587 ( .INP(n4582), .Z(n4751) );
  NOR2X0 U4588 ( .IN1(n7224), .IN2(n4483), .QN(n77) );
  NOR2X0 U4589 ( .IN1(n7236), .IN2(n4483), .QN(n67) );
  NOR2X0 U4590 ( .IN1(n7252), .IN2(n4483), .QN(n623) );
  NOR2X0 U4591 ( .IN1(n7253), .IN2(n4483), .QN(n621) );
  NOR2X0 U4592 ( .IN1(n7254), .IN2(n4483), .QN(n619) );
  NOR2X0 U4593 ( .IN1(n7094), .IN2(n4483), .QN(n548) );
  NOR2X0 U4594 ( .IN1(n7095), .IN2(n4483), .QN(n547) );
  NOR2X0 U4595 ( .IN1(n7096), .IN2(n4483), .QN(n546) );
  NOR2X0 U4596 ( .IN1(n7097), .IN2(n4483), .QN(n545) );
  INVX0 U4597 ( .INP(n4752), .ZN(n544) );
  NAND2X0 U4598 ( .IN1(n4445), .IN2(test_so80), .QN(n4752) );
  NOR2X0 U4599 ( .IN1(n7099), .IN2(n4483), .QN(n543) );
  NOR2X0 U4600 ( .IN1(n7100), .IN2(n4483), .QN(n542) );
  NOR2X0 U4601 ( .IN1(n7101), .IN2(n4483), .QN(n541) );
  NOR2X0 U4602 ( .IN1(n7102), .IN2(n4483), .QN(n540) );
  NOR2X0 U4603 ( .IN1(n7103), .IN2(n4484), .QN(n539) );
  NOR2X0 U4604 ( .IN1(n7104), .IN2(n4484), .QN(n538) );
  NOR2X0 U4605 ( .IN1(n7105), .IN2(n4484), .QN(n537) );
  NOR2X0 U4606 ( .IN1(n7106), .IN2(n4484), .QN(n536) );
  NOR2X0 U4607 ( .IN1(n7107), .IN2(n4484), .QN(n535) );
  NOR2X0 U4608 ( .IN1(n7108), .IN2(n4484), .QN(n534) );
  NOR2X0 U4609 ( .IN1(n7109), .IN2(n4484), .QN(n533) );
  NOR2X0 U4610 ( .IN1(n7122), .IN2(n4484), .QN(n470) );
  NOR2X0 U4611 ( .IN1(n7123), .IN2(n4484), .QN(n469) );
  NOR2X0 U4612 ( .IN1(n7124), .IN2(n4484), .QN(n468) );
  NOR2X0 U4613 ( .IN1(n7125), .IN2(n4484), .QN(n467) );
  NOR2X0 U4614 ( .IN1(n7126), .IN2(n4484), .QN(n466) );
  NOR2X0 U4615 ( .IN1(n7127), .IN2(n4484), .QN(n465) );
  NOR2X0 U4616 ( .IN1(n7128), .IN2(n4484), .QN(n464) );
  NOR2X0 U4617 ( .IN1(n7129), .IN2(n4484), .QN(n463) );
  NOR2X0 U4618 ( .IN1(n7130), .IN2(n4485), .QN(n462) );
  NOR2X0 U4619 ( .IN1(n7131), .IN2(n4485), .QN(n461) );
  NOR2X0 U4620 ( .IN1(n7132), .IN2(n4485), .QN(n460) );
  NOR2X0 U4621 ( .IN1(n7133), .IN2(n4485), .QN(n459) );
  NOR2X0 U4622 ( .IN1(n7134), .IN2(n4485), .QN(n458) );
  NOR2X0 U4623 ( .IN1(n7135), .IN2(n4485), .QN(n457) );
  NOR2X0 U4624 ( .IN1(n7136), .IN2(n4485), .QN(n456) );
  NOR2X0 U4625 ( .IN1(n7137), .IN2(n4485), .QN(n455) );
  NOR2X0 U4626 ( .IN1(n7150), .IN2(n4485), .QN(n392) );
  NOR2X0 U4627 ( .IN1(n7151), .IN2(n4485), .QN(n391) );
  NOR2X0 U4628 ( .IN1(n7152), .IN2(n4485), .QN(n390) );
  NOR2X0 U4629 ( .IN1(n7153), .IN2(n4485), .QN(n389) );
  NOR2X0 U4630 ( .IN1(n7154), .IN2(n4485), .QN(n388) );
  NOR2X0 U4631 ( .IN1(n7155), .IN2(n4485), .QN(n387) );
  NOR2X0 U4632 ( .IN1(n7156), .IN2(n4485), .QN(n386) );
  NOR2X0 U4633 ( .IN1(n7157), .IN2(n4486), .QN(n385) );
  NOR2X0 U4634 ( .IN1(n7158), .IN2(n4486), .QN(n384) );
  NOR2X0 U4635 ( .IN1(n7159), .IN2(n4486), .QN(n383) );
  NOR2X0 U4636 ( .IN1(n7160), .IN2(n4486), .QN(n382) );
  INVX0 U4637 ( .INP(n4753), .ZN(n381) );
  NAND2X0 U4638 ( .IN1(n4445), .IN2(test_so57), .QN(n4753) );
  NOR2X0 U4639 ( .IN1(n7162), .IN2(n4486), .QN(n380) );
  NOR2X0 U4640 ( .IN1(n7163), .IN2(n4486), .QN(n379) );
  NOR2X0 U4641 ( .IN1(n7164), .IN2(n4486), .QN(n378) );
  NOR2X0 U4642 ( .IN1(n7165), .IN2(n4486), .QN(n377) );
  NOR2X0 U4643 ( .IN1(TM1), .IN2(n4486), .QN(n3278) );
  NOR2X0 U4644 ( .IN1(n7178), .IN2(n4486), .QN(n314) );
  NOR2X0 U4645 ( .IN1(n7179), .IN2(n4486), .QN(n313) );
  NOR2X0 U4646 ( .IN1(n7180), .IN2(n4486), .QN(n312) );
  NOR2X0 U4647 ( .IN1(n7181), .IN2(n4486), .QN(n311) );
  NOR2X0 U4648 ( .IN1(n7182), .IN2(n4486), .QN(n310) );
  NOR2X0 U4649 ( .IN1(n7183), .IN2(n4486), .QN(n309) );
  INVX0 U4650 ( .INP(n4754), .ZN(n308) );
  NAND2X0 U4651 ( .IN1(n4445), .IN2(test_so46), .QN(n4754) );
  NOR2X0 U4652 ( .IN1(n7185), .IN2(n4487), .QN(n307) );
  NOR2X0 U4653 ( .IN1(n7186), .IN2(n4487), .QN(n306) );
  NOR2X0 U4654 ( .IN1(n7187), .IN2(n4491), .QN(n305) );
  NOR2X0 U4655 ( .IN1(n7188), .IN2(n4491), .QN(n304) );
  NOR2X0 U4656 ( .IN1(n7189), .IN2(n4490), .QN(n303) );
  NOR2X0 U4657 ( .IN1(n7190), .IN2(n4491), .QN(n302) );
  NOR2X0 U4658 ( .IN1(n7191), .IN2(n4490), .QN(n301) );
  NOR2X0 U4659 ( .IN1(n7192), .IN2(n4490), .QN(n300) );
  NOR2X0 U4660 ( .IN1(n7193), .IN2(n4490), .QN(n299) );
  NOR2X0 U4661 ( .IN1(n7199), .IN2(n4490), .QN(n236) );
  INVX0 U4662 ( .INP(n4755), .ZN(n235) );
  NAND2X0 U4663 ( .IN1(n4445), .IN2(test_so35), .QN(n4755) );
  NOR2X0 U4664 ( .IN1(n7201), .IN2(n4490), .QN(n234) );
  NOR2X0 U4665 ( .IN1(n7202), .IN2(n4490), .QN(n233) );
  NOR2X0 U4666 ( .IN1(n7203), .IN2(n4490), .QN(n232) );
  NOR2X0 U4667 ( .IN1(n7204), .IN2(n4490), .QN(n231) );
  NOR2X0 U4668 ( .IN1(n7205), .IN2(n4489), .QN(n230) );
  NOR2X0 U4669 ( .IN1(n7206), .IN2(n4490), .QN(n229) );
  NOR2X0 U4670 ( .IN1(n7207), .IN2(n4490), .QN(n228) );
  NOR2X0 U4671 ( .IN1(n7208), .IN2(n4490), .QN(n227) );
  NOR2X0 U4672 ( .IN1(n7209), .IN2(n4490), .QN(n226) );
  NOR2X0 U4673 ( .IN1(n7210), .IN2(n4490), .QN(n225) );
  NOR2X0 U4674 ( .IN1(n7211), .IN2(n4490), .QN(n224) );
  NOR2X0 U4675 ( .IN1(n7212), .IN2(n4489), .QN(n223) );
  NOR2X0 U4676 ( .IN1(n7213), .IN2(n4489), .QN(n222) );
  NOR2X0 U4677 ( .IN1(n7214), .IN2(n4489), .QN(n221) );
  INVX0 U4678 ( .INP(n4756), .ZN(n158) );
  NAND2X0 U4679 ( .IN1(n4445), .IN2(test_so24), .QN(n4756) );
  NOR2X0 U4680 ( .IN1(n7222), .IN2(n4489), .QN(n157) );
  NOR2X0 U4681 ( .IN1(n7223), .IN2(n4489), .QN(n156) );
  NOR2X0 U4682 ( .IN1(n7225), .IN2(n4489), .QN(n155) );
  NOR2X0 U4683 ( .IN1(n7226), .IN2(n4489), .QN(n154) );
  NOR2X0 U4684 ( .IN1(n7227), .IN2(n4489), .QN(n153) );
  NOR2X0 U4685 ( .IN1(n7228), .IN2(n4489), .QN(n152) );
  NOR2X0 U4686 ( .IN1(n7230), .IN2(n4489), .QN(n151) );
  NOR2X0 U4687 ( .IN1(n7231), .IN2(n4489), .QN(n150) );
  NOR2X0 U4688 ( .IN1(n7232), .IN2(n4489), .QN(n149) );
  NOR2X0 U4689 ( .IN1(n7233), .IN2(n4489), .QN(n148) );
  NOR2X0 U4690 ( .IN1(n7234), .IN2(n4489), .QN(n147) );
  NOR2X0 U4691 ( .IN1(n7235), .IN2(n4488), .QN(n146) );
  NOR2X0 U4692 ( .IN1(n7237), .IN2(n4488), .QN(n145) );
  NOR2X0 U4693 ( .IN1(n7238), .IN2(n4488), .QN(n144) );
  NOR2X0 U4694 ( .IN1(n7239), .IN2(n4488), .QN(n143) );
  NAND4X0 U4695 ( .IN1(n4757), .IN2(n4758), .IN3(n4759), .IN4(n4760), .QN(
        WX9757) );
  NAND2X0 U4696 ( .IN1(n3886), .IN2(n4762), .QN(n4760) );
  NAND2X0 U4697 ( .IN1(n3965), .IN2(n4763), .QN(n4759) );
  NAND2X0 U4698 ( .IN1(n532), .IN2(n3915), .QN(n4758) );
  INVX0 U4699 ( .INP(n4764), .ZN(n532) );
  NAND2X0 U4700 ( .IN1(n4445), .IN2(n8321), .QN(n4764) );
  NAND2X0 U4701 ( .IN1(n3934), .IN2(CRC_OUT_2_0), .QN(n4757) );
  NAND4X0 U4702 ( .IN1(n4765), .IN2(n4766), .IN3(n4767), .IN4(n4768), .QN(
        WX9755) );
  NAND2X0 U4703 ( .IN1(n4769), .IN2(n3901), .QN(n4768) );
  NAND2X0 U4704 ( .IN1(n3977), .IN2(n4770), .QN(n4767) );
  NAND2X0 U4705 ( .IN1(n531), .IN2(n3915), .QN(n4766) );
  INVX0 U4706 ( .INP(n4771), .ZN(n531) );
  NAND2X0 U4707 ( .IN1(n4444), .IN2(n8322), .QN(n4771) );
  NAND2X0 U4708 ( .IN1(n3951), .IN2(CRC_OUT_2_1), .QN(n4765) );
  NAND4X0 U4709 ( .IN1(n4772), .IN2(n4773), .IN3(n4774), .IN4(n4775), .QN(
        WX9753) );
  NAND2X0 U4710 ( .IN1(n3888), .IN2(n4776), .QN(n4775) );
  NAND2X0 U4711 ( .IN1(n4777), .IN2(n3983), .QN(n4774) );
  NAND2X0 U4712 ( .IN1(n530), .IN2(n3915), .QN(n4773) );
  INVX0 U4713 ( .INP(n4778), .ZN(n530) );
  NAND2X0 U4714 ( .IN1(n4444), .IN2(n8323), .QN(n4778) );
  NAND2X0 U4715 ( .IN1(test_so87), .IN2(n3957), .QN(n4772) );
  NAND4X0 U4716 ( .IN1(n4779), .IN2(n4780), .IN3(n4781), .IN4(n4782), .QN(
        WX9751) );
  NAND2X0 U4717 ( .IN1(n4783), .IN2(n3900), .QN(n4782) );
  NAND2X0 U4718 ( .IN1(n3974), .IN2(n4784), .QN(n4781) );
  NAND2X0 U4719 ( .IN1(n529), .IN2(n3915), .QN(n4780) );
  INVX0 U4720 ( .INP(n4785), .ZN(n529) );
  NAND2X0 U4721 ( .IN1(n4444), .IN2(n8324), .QN(n4785) );
  NAND2X0 U4722 ( .IN1(n3945), .IN2(CRC_OUT_2_3), .QN(n4779) );
  NAND4X0 U4723 ( .IN1(n4786), .IN2(n4787), .IN3(n4788), .IN4(n4789), .QN(
        WX9749) );
  NAND2X0 U4724 ( .IN1(n3888), .IN2(n4790), .QN(n4789) );
  NAND2X0 U4725 ( .IN1(n4791), .IN2(n3984), .QN(n4788) );
  NAND2X0 U4726 ( .IN1(n528), .IN2(n3915), .QN(n4787) );
  INVX0 U4727 ( .INP(n4792), .ZN(n528) );
  NAND2X0 U4728 ( .IN1(n4444), .IN2(n8325), .QN(n4792) );
  NAND2X0 U4729 ( .IN1(n3945), .IN2(CRC_OUT_2_4), .QN(n4786) );
  NAND4X0 U4730 ( .IN1(n4793), .IN2(n4794), .IN3(n4795), .IN4(n4796), .QN(
        WX9747) );
  NAND2X0 U4731 ( .IN1(n3888), .IN2(n4797), .QN(n4796) );
  NAND2X0 U4732 ( .IN1(n3974), .IN2(n4798), .QN(n4795) );
  NAND2X0 U4733 ( .IN1(n527), .IN2(n3915), .QN(n4794) );
  INVX0 U4734 ( .INP(n4799), .ZN(n527) );
  NAND2X0 U4735 ( .IN1(test_so79), .IN2(n4463), .QN(n4799) );
  NAND2X0 U4736 ( .IN1(n3945), .IN2(CRC_OUT_2_5), .QN(n4793) );
  NAND4X0 U4737 ( .IN1(n4800), .IN2(n4801), .IN3(n4802), .IN4(n4803), .QN(
        WX9745) );
  NAND2X0 U4738 ( .IN1(n3888), .IN2(n4804), .QN(n4803) );
  NAND2X0 U4739 ( .IN1(n4805), .IN2(n3984), .QN(n4802) );
  NAND2X0 U4740 ( .IN1(n526), .IN2(n3915), .QN(n4801) );
  INVX0 U4741 ( .INP(n4806), .ZN(n526) );
  NAND2X0 U4742 ( .IN1(n4444), .IN2(n8328), .QN(n4806) );
  NAND2X0 U4743 ( .IN1(n3945), .IN2(CRC_OUT_2_6), .QN(n4800) );
  NAND4X0 U4744 ( .IN1(n4807), .IN2(n4808), .IN3(n4809), .IN4(n4810), .QN(
        WX9743) );
  NAND2X0 U4745 ( .IN1(n3888), .IN2(n4811), .QN(n4810) );
  NAND2X0 U4746 ( .IN1(n3974), .IN2(n4812), .QN(n4809) );
  NAND2X0 U4747 ( .IN1(n525), .IN2(n3915), .QN(n4808) );
  INVX0 U4748 ( .INP(n4813), .ZN(n525) );
  NAND2X0 U4749 ( .IN1(n4444), .IN2(n8329), .QN(n4813) );
  NAND2X0 U4750 ( .IN1(n3946), .IN2(CRC_OUT_2_7), .QN(n4807) );
  NAND4X0 U4751 ( .IN1(n4814), .IN2(n4815), .IN3(n4816), .IN4(n4817), .QN(
        WX9741) );
  NAND2X0 U4752 ( .IN1(n3887), .IN2(n4818), .QN(n4817) );
  NAND2X0 U4753 ( .IN1(n4819), .IN2(n3983), .QN(n4816) );
  NAND2X0 U4754 ( .IN1(n524), .IN2(n3915), .QN(n4815) );
  INVX0 U4755 ( .INP(n4820), .ZN(n524) );
  NAND2X0 U4756 ( .IN1(n4444), .IN2(n8330), .QN(n4820) );
  NAND2X0 U4757 ( .IN1(n3946), .IN2(CRC_OUT_2_8), .QN(n4814) );
  NAND4X0 U4758 ( .IN1(n4821), .IN2(n4822), .IN3(n4823), .IN4(n4824), .QN(
        WX9739) );
  NAND2X0 U4759 ( .IN1(n3887), .IN2(n4825), .QN(n4824) );
  NAND2X0 U4760 ( .IN1(n3974), .IN2(n4826), .QN(n4823) );
  NAND2X0 U4761 ( .IN1(n523), .IN2(n3915), .QN(n4822) );
  INVX0 U4762 ( .INP(n4827), .ZN(n523) );
  NAND2X0 U4763 ( .IN1(n4444), .IN2(n8331), .QN(n4827) );
  NAND2X0 U4764 ( .IN1(n3946), .IN2(CRC_OUT_2_9), .QN(n4821) );
  NAND4X0 U4765 ( .IN1(n4828), .IN2(n4829), .IN3(n4830), .IN4(n4831), .QN(
        WX9737) );
  NAND2X0 U4766 ( .IN1(n3887), .IN2(n4832), .QN(n4831) );
  NAND2X0 U4767 ( .IN1(n3974), .IN2(n4833), .QN(n4830) );
  NAND2X0 U4768 ( .IN1(n522), .IN2(n3915), .QN(n4829) );
  INVX0 U4769 ( .INP(n4834), .ZN(n522) );
  NAND2X0 U4770 ( .IN1(n4444), .IN2(n8332), .QN(n4834) );
  NAND2X0 U4771 ( .IN1(n3946), .IN2(CRC_OUT_2_10), .QN(n4828) );
  NAND4X0 U4772 ( .IN1(n4835), .IN2(n4836), .IN3(n4837), .IN4(n4838), .QN(
        WX9735) );
  NAND2X0 U4773 ( .IN1(n3887), .IN2(n4839), .QN(n4838) );
  NAND2X0 U4774 ( .IN1(n3974), .IN2(n4840), .QN(n4837) );
  NAND2X0 U4775 ( .IN1(n521), .IN2(n3915), .QN(n4836) );
  INVX0 U4776 ( .INP(n4841), .ZN(n521) );
  NAND2X0 U4777 ( .IN1(n4443), .IN2(n8333), .QN(n4841) );
  NAND2X0 U4778 ( .IN1(n3946), .IN2(CRC_OUT_2_11), .QN(n4835) );
  NAND4X0 U4779 ( .IN1(n4842), .IN2(n4843), .IN3(n4844), .IN4(n4845), .QN(
        WX9733) );
  NAND2X0 U4780 ( .IN1(n3887), .IN2(n4846), .QN(n4845) );
  NAND2X0 U4781 ( .IN1(n3974), .IN2(n4847), .QN(n4844) );
  NAND2X0 U4782 ( .IN1(n520), .IN2(n3915), .QN(n4843) );
  INVX0 U4783 ( .INP(n4848), .ZN(n520) );
  NAND2X0 U4784 ( .IN1(n4443), .IN2(n8334), .QN(n4848) );
  NAND2X0 U4785 ( .IN1(n3946), .IN2(CRC_OUT_2_12), .QN(n4842) );
  NAND4X0 U4786 ( .IN1(n4849), .IN2(n4850), .IN3(n4851), .IN4(n4852), .QN(
        WX9731) );
  NAND2X0 U4787 ( .IN1(n3887), .IN2(n4853), .QN(n4852) );
  NAND2X0 U4788 ( .IN1(n3975), .IN2(n4854), .QN(n4851) );
  NAND2X0 U4789 ( .IN1(n519), .IN2(n3915), .QN(n4850) );
  INVX0 U4790 ( .INP(n4855), .ZN(n519) );
  NAND2X0 U4791 ( .IN1(n4443), .IN2(n8335), .QN(n4855) );
  NAND2X0 U4792 ( .IN1(n3946), .IN2(CRC_OUT_2_13), .QN(n4849) );
  NAND4X0 U4793 ( .IN1(n4856), .IN2(n4857), .IN3(n4858), .IN4(n4859), .QN(
        WX9729) );
  NAND2X0 U4794 ( .IN1(n4860), .IN2(n3900), .QN(n4859) );
  NAND2X0 U4795 ( .IN1(n3975), .IN2(n4861), .QN(n4858) );
  NAND2X0 U4796 ( .IN1(n518), .IN2(n3915), .QN(n4857) );
  INVX0 U4797 ( .INP(n4862), .ZN(n518) );
  NAND2X0 U4798 ( .IN1(n4443), .IN2(n8336), .QN(n4862) );
  NAND2X0 U4799 ( .IN1(n3946), .IN2(CRC_OUT_2_14), .QN(n4856) );
  NAND4X0 U4800 ( .IN1(n4863), .IN2(n4864), .IN3(n4865), .IN4(n4866), .QN(
        WX9727) );
  NAND2X0 U4801 ( .IN1(n3887), .IN2(n4867), .QN(n4866) );
  NAND2X0 U4802 ( .IN1(n3975), .IN2(n4868), .QN(n4865) );
  NAND2X0 U4803 ( .IN1(n517), .IN2(n3915), .QN(n4864) );
  INVX0 U4804 ( .INP(n4869), .ZN(n517) );
  NAND2X0 U4805 ( .IN1(n4443), .IN2(n8337), .QN(n4869) );
  NAND2X0 U4806 ( .IN1(n3946), .IN2(CRC_OUT_2_15), .QN(n4863) );
  NAND4X0 U4807 ( .IN1(n4870), .IN2(n4871), .IN3(n4872), .IN4(n4873), .QN(
        WX9725) );
  NAND2X0 U4808 ( .IN1(n4874), .IN2(n3900), .QN(n4873) );
  NAND2X0 U4809 ( .IN1(n3975), .IN2(n4875), .QN(n4872) );
  NAND2X0 U4810 ( .IN1(n516), .IN2(n3916), .QN(n4871) );
  INVX0 U4811 ( .INP(n4876), .ZN(n516) );
  NAND2X0 U4812 ( .IN1(n4443), .IN2(n8338), .QN(n4876) );
  NAND2X0 U4813 ( .IN1(n3946), .IN2(CRC_OUT_2_16), .QN(n4870) );
  NAND4X0 U4814 ( .IN1(n4877), .IN2(n4878), .IN3(n4879), .IN4(n4880), .QN(
        WX9723) );
  NAND2X0 U4815 ( .IN1(n3887), .IN2(n4881), .QN(n4880) );
  NAND2X0 U4816 ( .IN1(n3975), .IN2(n4882), .QN(n4879) );
  NAND2X0 U4817 ( .IN1(n515), .IN2(n3916), .QN(n4878) );
  INVX0 U4818 ( .INP(n4883), .ZN(n515) );
  NAND2X0 U4819 ( .IN1(n4443), .IN2(n8339), .QN(n4883) );
  NAND2X0 U4820 ( .IN1(n3946), .IN2(CRC_OUT_2_17), .QN(n4877) );
  NAND4X0 U4821 ( .IN1(n4884), .IN2(n4885), .IN3(n4886), .IN4(n4887), .QN(
        WX9721) );
  NAND2X0 U4822 ( .IN1(n4888), .IN2(n3900), .QN(n4887) );
  NAND2X0 U4823 ( .IN1(n3975), .IN2(n4889), .QN(n4886) );
  NAND2X0 U4824 ( .IN1(n514), .IN2(n3916), .QN(n4885) );
  INVX0 U4825 ( .INP(n4890), .ZN(n514) );
  NAND2X0 U4826 ( .IN1(n4443), .IN2(n8340), .QN(n4890) );
  NAND2X0 U4827 ( .IN1(n3946), .IN2(CRC_OUT_2_18), .QN(n4884) );
  NAND4X0 U4828 ( .IN1(n4891), .IN2(n4892), .IN3(n4893), .IN4(n4894), .QN(
        WX9719) );
  NAND2X0 U4829 ( .IN1(n3887), .IN2(n4895), .QN(n4894) );
  NAND2X0 U4830 ( .IN1(n4896), .IN2(n3984), .QN(n4893) );
  NAND2X0 U4831 ( .IN1(n513), .IN2(n3916), .QN(n4892) );
  INVX0 U4832 ( .INP(n4897), .ZN(n513) );
  NAND2X0 U4833 ( .IN1(n4443), .IN2(n8341), .QN(n4897) );
  NAND2X0 U4834 ( .IN1(test_so88), .IN2(n3956), .QN(n4891) );
  NAND4X0 U4835 ( .IN1(n4898), .IN2(n4899), .IN3(n4900), .IN4(n4901), .QN(
        WX9717) );
  NAND2X0 U4836 ( .IN1(n4902), .IN2(n3900), .QN(n4901) );
  NAND2X0 U4837 ( .IN1(n3975), .IN2(n4903), .QN(n4900) );
  NAND2X0 U4838 ( .IN1(n512), .IN2(n3916), .QN(n4899) );
  INVX0 U4839 ( .INP(n4904), .ZN(n512) );
  NAND2X0 U4840 ( .IN1(n4442), .IN2(n8342), .QN(n4904) );
  NAND2X0 U4841 ( .IN1(n3947), .IN2(CRC_OUT_2_20), .QN(n4898) );
  NAND4X0 U4842 ( .IN1(n4905), .IN2(n4906), .IN3(n4907), .IN4(n4908), .QN(
        WX9715) );
  NAND2X0 U4843 ( .IN1(n3887), .IN2(n4909), .QN(n4908) );
  NAND2X0 U4844 ( .IN1(n4910), .IN2(n3985), .QN(n4907) );
  NAND2X0 U4845 ( .IN1(n511), .IN2(n3916), .QN(n4906) );
  INVX0 U4846 ( .INP(n4911), .ZN(n511) );
  NAND2X0 U4847 ( .IN1(n4442), .IN2(n8343), .QN(n4911) );
  NAND2X0 U4848 ( .IN1(n3947), .IN2(CRC_OUT_2_21), .QN(n4905) );
  NAND4X0 U4849 ( .IN1(n4912), .IN2(n4913), .IN3(n4914), .IN4(n4915), .QN(
        WX9713) );
  NAND2X0 U4850 ( .IN1(n3887), .IN2(n4916), .QN(n4915) );
  NAND2X0 U4851 ( .IN1(n3975), .IN2(n4917), .QN(n4914) );
  NAND2X0 U4852 ( .IN1(n510), .IN2(n3916), .QN(n4913) );
  INVX0 U4853 ( .INP(n4918), .ZN(n510) );
  NAND2X0 U4854 ( .IN1(test_so78), .IN2(n4463), .QN(n4918) );
  NAND2X0 U4855 ( .IN1(n3947), .IN2(CRC_OUT_2_22), .QN(n4912) );
  NAND4X0 U4856 ( .IN1(n4919), .IN2(n4920), .IN3(n4921), .IN4(n4922), .QN(
        WX9711) );
  NAND2X0 U4857 ( .IN1(n3887), .IN2(n4923), .QN(n4922) );
  NAND2X0 U4858 ( .IN1(n4924), .IN2(n3985), .QN(n4921) );
  NAND2X0 U4859 ( .IN1(n509), .IN2(n3916), .QN(n4920) );
  INVX0 U4860 ( .INP(n4925), .ZN(n509) );
  NAND2X0 U4861 ( .IN1(n4442), .IN2(n8346), .QN(n4925) );
  NAND2X0 U4862 ( .IN1(n3947), .IN2(CRC_OUT_2_23), .QN(n4919) );
  NAND4X0 U4863 ( .IN1(n4926), .IN2(n4927), .IN3(n4928), .IN4(n4929), .QN(
        WX9709) );
  NAND2X0 U4864 ( .IN1(n3886), .IN2(n4930), .QN(n4929) );
  NAND2X0 U4865 ( .IN1(n3975), .IN2(n4931), .QN(n4928) );
  NAND2X0 U4866 ( .IN1(n508), .IN2(n3916), .QN(n4927) );
  INVX0 U4867 ( .INP(n4932), .ZN(n508) );
  NAND2X0 U4868 ( .IN1(n4442), .IN2(n8347), .QN(n4932) );
  NAND2X0 U4869 ( .IN1(n3947), .IN2(CRC_OUT_2_24), .QN(n4926) );
  NAND4X0 U4870 ( .IN1(n4933), .IN2(n4934), .IN3(n4935), .IN4(n4936), .QN(
        WX9707) );
  NAND2X0 U4871 ( .IN1(n3886), .IN2(n4937), .QN(n4936) );
  NAND2X0 U4872 ( .IN1(n4938), .IN2(n3985), .QN(n4935) );
  NAND2X0 U4873 ( .IN1(n507), .IN2(n3916), .QN(n4934) );
  INVX0 U4874 ( .INP(n4939), .ZN(n507) );
  NAND2X0 U4875 ( .IN1(n4442), .IN2(n8348), .QN(n4939) );
  NAND2X0 U4876 ( .IN1(n3947), .IN2(CRC_OUT_2_25), .QN(n4933) );
  NAND4X0 U4877 ( .IN1(n4940), .IN2(n4941), .IN3(n4942), .IN4(n4943), .QN(
        WX9705) );
  NAND2X0 U4878 ( .IN1(n3886), .IN2(n4944), .QN(n4943) );
  NAND2X0 U4879 ( .IN1(n3975), .IN2(n4945), .QN(n4942) );
  NAND2X0 U4880 ( .IN1(n506), .IN2(n3916), .QN(n4941) );
  INVX0 U4881 ( .INP(n4946), .ZN(n506) );
  NAND2X0 U4882 ( .IN1(n4442), .IN2(n8349), .QN(n4946) );
  NAND2X0 U4883 ( .IN1(n3947), .IN2(CRC_OUT_2_26), .QN(n4940) );
  NAND4X0 U4884 ( .IN1(n4947), .IN2(n4948), .IN3(n4949), .IN4(n4950), .QN(
        WX9703) );
  NAND2X0 U4885 ( .IN1(n3886), .IN2(n4951), .QN(n4950) );
  NAND2X0 U4886 ( .IN1(n3975), .IN2(n4952), .QN(n4949) );
  NAND2X0 U4887 ( .IN1(n505), .IN2(n3916), .QN(n4948) );
  INVX0 U4888 ( .INP(n4953), .ZN(n505) );
  NAND2X0 U4889 ( .IN1(n4442), .IN2(n8350), .QN(n4953) );
  NAND2X0 U4890 ( .IN1(n3947), .IN2(CRC_OUT_2_27), .QN(n4947) );
  NAND4X0 U4891 ( .IN1(n4954), .IN2(n4955), .IN3(n4956), .IN4(n4957), .QN(
        WX9701) );
  NAND2X0 U4892 ( .IN1(n3886), .IN2(n4958), .QN(n4957) );
  NAND2X0 U4893 ( .IN1(n3975), .IN2(n4959), .QN(n4956) );
  NAND2X0 U4894 ( .IN1(n504), .IN2(n3916), .QN(n4955) );
  INVX0 U4895 ( .INP(n4960), .ZN(n504) );
  NAND2X0 U4896 ( .IN1(n4442), .IN2(n8351), .QN(n4960) );
  NAND2X0 U4897 ( .IN1(n3947), .IN2(CRC_OUT_2_28), .QN(n4954) );
  NAND4X0 U4898 ( .IN1(n4961), .IN2(n4962), .IN3(n4963), .IN4(n4964), .QN(
        WX9699) );
  NAND2X0 U4899 ( .IN1(n3886), .IN2(n4965), .QN(n4964) );
  NAND2X0 U4900 ( .IN1(n3976), .IN2(n4966), .QN(n4963) );
  NAND2X0 U4901 ( .IN1(n503), .IN2(n3916), .QN(n4962) );
  INVX0 U4902 ( .INP(n4967), .ZN(n503) );
  NAND2X0 U4903 ( .IN1(n4442), .IN2(n8352), .QN(n4967) );
  NAND2X0 U4904 ( .IN1(n3947), .IN2(CRC_OUT_2_29), .QN(n4961) );
  NAND4X0 U4905 ( .IN1(n4968), .IN2(n4969), .IN3(n4970), .IN4(n4971), .QN(
        WX9697) );
  NAND2X0 U4906 ( .IN1(n3886), .IN2(n4972), .QN(n4971) );
  NAND2X0 U4907 ( .IN1(n3976), .IN2(n4973), .QN(n4970) );
  NAND2X0 U4908 ( .IN1(n502), .IN2(n3916), .QN(n4969) );
  INVX0 U4909 ( .INP(n4974), .ZN(n502) );
  NAND2X0 U4910 ( .IN1(n4441), .IN2(n8353), .QN(n4974) );
  NAND2X0 U4911 ( .IN1(n3947), .IN2(CRC_OUT_2_30), .QN(n4968) );
  NAND4X0 U4912 ( .IN1(n4975), .IN2(n4976), .IN3(n4977), .IN4(n4978), .QN(
        WX9695) );
  NAND2X0 U4913 ( .IN1(n4979), .IN2(n3899), .QN(n4978) );
  NAND2X0 U4914 ( .IN1(n3976), .IN2(n4980), .QN(n4977) );
  NAND2X0 U4915 ( .IN1(n3947), .IN2(CRC_OUT_2_31), .QN(n4976) );
  NAND2X0 U4916 ( .IN1(n2245), .IN2(WX9536), .QN(n4975) );
  NOR2X0 U4917 ( .IN1(n4550), .IN2(WX9536), .QN(WX9597) );
  NOR2X0 U4918 ( .IN1(n4563), .IN2(n4981), .QN(WX9084) );
  XOR2X1 U4919 ( .IN1(n3518), .IN2(DFF_1342_n1), .Q(n4981) );
  NOR2X0 U4920 ( .IN1(n4558), .IN2(n4982), .QN(WX9082) );
  XOR2X1 U4921 ( .IN1(n3520), .IN2(DFF_1341_n1), .Q(n4982) );
  NOR2X0 U4922 ( .IN1(n4558), .IN2(n4983), .QN(WX9080) );
  XOR2X1 U4923 ( .IN1(n3522), .IN2(DFF_1340_n1), .Q(n4983) );
  NOR2X0 U4924 ( .IN1(n4558), .IN2(n4984), .QN(WX9078) );
  XOR2X1 U4925 ( .IN1(n3523), .IN2(DFF_1339_n1), .Q(n4984) );
  NOR2X0 U4926 ( .IN1(n4558), .IN2(n4985), .QN(WX9076) );
  XOR2X1 U4927 ( .IN1(n3524), .IN2(DFF_1338_n1), .Q(n4985) );
  NOR2X0 U4928 ( .IN1(n4559), .IN2(n4986), .QN(WX9074) );
  XOR2X1 U4929 ( .IN1(CRC_OUT_3_25), .IN2(test_so74), .Q(n4986) );
  NOR2X0 U4930 ( .IN1(n4559), .IN2(n4987), .QN(WX9072) );
  XNOR2X1 U4931 ( .IN1(n3526), .IN2(test_so77), .Q(n4987) );
  NOR2X0 U4932 ( .IN1(n4559), .IN2(n4988), .QN(WX9070) );
  XOR2X1 U4933 ( .IN1(n3528), .IN2(DFF_1335_n1), .Q(n4988) );
  NOR2X0 U4934 ( .IN1(n4559), .IN2(n4989), .QN(WX9068) );
  XOR2X1 U4935 ( .IN1(n3530), .IN2(DFF_1334_n1), .Q(n4989) );
  NOR2X0 U4936 ( .IN1(n4559), .IN2(n4990), .QN(WX9066) );
  XOR2X1 U4937 ( .IN1(n3532), .IN2(DFF_1333_n1), .Q(n4990) );
  NOR2X0 U4938 ( .IN1(n4559), .IN2(n4991), .QN(WX9064) );
  XOR2X1 U4939 ( .IN1(n3534), .IN2(DFF_1332_n1), .Q(n4991) );
  NOR2X0 U4940 ( .IN1(n4559), .IN2(n4992), .QN(WX9062) );
  XOR2X1 U4941 ( .IN1(n3536), .IN2(DFF_1331_n1), .Q(n4992) );
  NOR2X0 U4942 ( .IN1(n4559), .IN2(n4993), .QN(WX9060) );
  XOR2X1 U4943 ( .IN1(n3538), .IN2(DFF_1330_n1), .Q(n4993) );
  NOR2X0 U4944 ( .IN1(n4559), .IN2(n4994), .QN(WX9058) );
  XOR2X1 U4945 ( .IN1(n3540), .IN2(DFF_1329_n1), .Q(n4994) );
  NOR2X0 U4946 ( .IN1(n4559), .IN2(n4995), .QN(WX9056) );
  XOR2X1 U4947 ( .IN1(n3542), .IN2(DFF_1328_n1), .Q(n4995) );
  NOR2X0 U4948 ( .IN1(n4559), .IN2(n4996), .QN(WX9054) );
  XOR3X1 U4949 ( .IN1(n3418), .IN2(DFF_1343_n1), .IN3(CRC_OUT_3_15), .Q(n4996)
         );
  NOR2X0 U4950 ( .IN1(n4559), .IN2(n4997), .QN(WX9052) );
  XOR2X1 U4951 ( .IN1(n3543), .IN2(DFF_1326_n1), .Q(n4997) );
  NOR2X0 U4952 ( .IN1(n4559), .IN2(n4998), .QN(WX9050) );
  XOR2X1 U4953 ( .IN1(n3544), .IN2(DFF_1325_n1), .Q(n4998) );
  NOR2X0 U4954 ( .IN1(n4559), .IN2(n4999), .QN(WX9048) );
  XOR2X1 U4955 ( .IN1(n3546), .IN2(DFF_1324_n1), .Q(n4999) );
  NOR2X0 U4956 ( .IN1(n4559), .IN2(n5000), .QN(WX9046) );
  XOR2X1 U4957 ( .IN1(n3548), .IN2(DFF_1323_n1), .Q(n5000) );
  NOR2X0 U4958 ( .IN1(n4559), .IN2(n5001), .QN(WX9044) );
  XOR3X1 U4959 ( .IN1(n3419), .IN2(DFF_1343_n1), .IN3(CRC_OUT_3_10), .Q(n5001)
         );
  NOR2X0 U4960 ( .IN1(n4560), .IN2(n5002), .QN(WX9042) );
  XOR2X1 U4961 ( .IN1(n3550), .IN2(DFF_1321_n1), .Q(n5002) );
  NOR2X0 U4962 ( .IN1(n4560), .IN2(n5003), .QN(WX9040) );
  XOR2X1 U4963 ( .IN1(CRC_OUT_3_8), .IN2(test_so75), .Q(n5003) );
  NOR2X0 U4964 ( .IN1(n4560), .IN2(n5004), .QN(WX9038) );
  XNOR2X1 U4965 ( .IN1(n3552), .IN2(test_so76), .Q(n5004) );
  NOR2X0 U4966 ( .IN1(n4560), .IN2(n5005), .QN(WX9036) );
  XOR2X1 U4967 ( .IN1(n3554), .IN2(DFF_1318_n1), .Q(n5005) );
  NOR2X0 U4968 ( .IN1(n4560), .IN2(n5006), .QN(WX9034) );
  XOR2X1 U4969 ( .IN1(n3556), .IN2(DFF_1317_n1), .Q(n5006) );
  NOR2X0 U4970 ( .IN1(n4560), .IN2(n5007), .QN(WX9032) );
  XOR2X1 U4971 ( .IN1(n3558), .IN2(DFF_1316_n1), .Q(n5007) );
  NOR2X0 U4972 ( .IN1(n4560), .IN2(n5008), .QN(WX9030) );
  XOR3X1 U4973 ( .IN1(n3420), .IN2(DFF_1343_n1), .IN3(CRC_OUT_3_3), .Q(n5008)
         );
  NOR2X0 U4974 ( .IN1(n4560), .IN2(n5009), .QN(WX9028) );
  XOR2X1 U4975 ( .IN1(n3560), .IN2(DFF_1314_n1), .Q(n5009) );
  NOR2X0 U4976 ( .IN1(n4560), .IN2(n5010), .QN(WX9026) );
  XOR2X1 U4977 ( .IN1(n3562), .IN2(DFF_1313_n1), .Q(n5010) );
  NOR2X0 U4978 ( .IN1(n4560), .IN2(n5011), .QN(WX9024) );
  XOR2X1 U4979 ( .IN1(n3564), .IN2(DFF_1312_n1), .Q(n5011) );
  NOR2X0 U4980 ( .IN1(n4560), .IN2(n5012), .QN(WX9022) );
  XOR2X1 U4981 ( .IN1(n3435), .IN2(DFF_1343_n1), .Q(n5012) );
  NAND4X0 U4982 ( .IN1(n5013), .IN2(n5014), .IN3(n5015), .IN4(n5016), .QN(
        WX8464) );
  NAND2X0 U4983 ( .IN1(n3976), .IN2(n4762), .QN(n5016) );
  XNOR3X1 U4984 ( .IN1(n3434), .IN2(n3303), .IN3(n5017), .Q(n4762) );
  XOR2X1 U4985 ( .IN1(WX9822), .IN2(n7081), .Q(n5017) );
  NAND2X0 U4986 ( .IN1(n3886), .IN2(n5018), .QN(n5015) );
  NAND2X0 U4987 ( .IN1(n454), .IN2(n3916), .QN(n5014) );
  INVX0 U4988 ( .INP(n5019), .ZN(n454) );
  NAND2X0 U4989 ( .IN1(test_so68), .IN2(n4463), .QN(n5019) );
  NAND2X0 U4990 ( .IN1(n3948), .IN2(CRC_OUT_3_0), .QN(n5013) );
  NAND4X0 U4991 ( .IN1(n5020), .IN2(n5021), .IN3(n5022), .IN4(n5023), .QN(
        WX8462) );
  NAND2X0 U4992 ( .IN1(n4769), .IN2(n3985), .QN(n5023) );
  XOR3X1 U4993 ( .IN1(n3516), .IN2(n3304), .IN3(n5024), .Q(n4769) );
  XOR2X1 U4994 ( .IN1(WX9756), .IN2(test_so83), .Q(n5024) );
  NAND2X0 U4995 ( .IN1(n3886), .IN2(n5025), .QN(n5022) );
  NAND2X0 U4996 ( .IN1(n453), .IN2(n3916), .QN(n5021) );
  INVX0 U4997 ( .INP(n5026), .ZN(n453) );
  NAND2X0 U4998 ( .IN1(n4441), .IN2(n8381), .QN(n5026) );
  NAND2X0 U4999 ( .IN1(n3948), .IN2(CRC_OUT_3_1), .QN(n5020) );
  NAND4X0 U5000 ( .IN1(n5027), .IN2(n5028), .IN3(n5029), .IN4(n5030), .QN(
        WX8460) );
  NAND2X0 U5001 ( .IN1(n3976), .IN2(n4776), .QN(n5030) );
  XNOR3X1 U5002 ( .IN1(n3514), .IN2(n3305), .IN3(n5031), .Q(n4776) );
  XOR2X1 U5003 ( .IN1(WX9818), .IN2(n7082), .Q(n5031) );
  NAND2X0 U5004 ( .IN1(n3886), .IN2(n5032), .QN(n5029) );
  NAND2X0 U5005 ( .IN1(n452), .IN2(n3917), .QN(n5028) );
  INVX0 U5006 ( .INP(n5033), .ZN(n452) );
  NAND2X0 U5007 ( .IN1(n4441), .IN2(n8382), .QN(n5033) );
  NAND2X0 U5008 ( .IN1(n3948), .IN2(CRC_OUT_3_2), .QN(n5027) );
  NAND4X0 U5009 ( .IN1(n5034), .IN2(n5035), .IN3(n5036), .IN4(n5037), .QN(
        WX8458) );
  NAND2X0 U5010 ( .IN1(n4783), .IN2(n3985), .QN(n5037) );
  XOR3X1 U5011 ( .IN1(n3569), .IN2(n3512), .IN3(n5038), .Q(n4783) );
  XOR2X1 U5012 ( .IN1(WX9880), .IN2(test_so81), .Q(n5038) );
  NAND2X0 U5013 ( .IN1(n3886), .IN2(n5039), .QN(n5036) );
  NAND2X0 U5014 ( .IN1(n451), .IN2(n3917), .QN(n5035) );
  INVX0 U5015 ( .INP(n5040), .ZN(n451) );
  NAND2X0 U5016 ( .IN1(n4441), .IN2(n8383), .QN(n5040) );
  NAND2X0 U5017 ( .IN1(n3948), .IN2(CRC_OUT_3_3), .QN(n5034) );
  NAND4X0 U5018 ( .IN1(n5041), .IN2(n5042), .IN3(n5043), .IN4(n5044), .QN(
        WX8456) );
  NAND2X0 U5019 ( .IN1(n3976), .IN2(n4790), .QN(n5044) );
  XNOR3X1 U5020 ( .IN1(n3417), .IN2(n3306), .IN3(n5045), .Q(n4790) );
  XOR2X1 U5021 ( .IN1(WX9814), .IN2(n7083), .Q(n5045) );
  NAND2X0 U5022 ( .IN1(n3888), .IN2(n5046), .QN(n5043) );
  NAND2X0 U5023 ( .IN1(n450), .IN2(n3917), .QN(n5042) );
  INVX0 U5024 ( .INP(n5047), .ZN(n450) );
  NAND2X0 U5025 ( .IN1(n4441), .IN2(n8384), .QN(n5047) );
  NAND2X0 U5026 ( .IN1(n3948), .IN2(CRC_OUT_3_4), .QN(n5041) );
  NAND4X0 U5027 ( .IN1(n5048), .IN2(n5049), .IN3(n5050), .IN4(n5051), .QN(
        WX8454) );
  NAND2X0 U5028 ( .IN1(n3976), .IN2(n4797), .QN(n5051) );
  XNOR3X1 U5029 ( .IN1(n3510), .IN2(n3307), .IN3(n5052), .Q(n4797) );
  XOR2X1 U5030 ( .IN1(WX9812), .IN2(n7084), .Q(n5052) );
  NAND2X0 U5031 ( .IN1(n3885), .IN2(n5053), .QN(n5050) );
  NAND2X0 U5032 ( .IN1(n449), .IN2(n3917), .QN(n5049) );
  INVX0 U5033 ( .INP(n5054), .ZN(n449) );
  NAND2X0 U5034 ( .IN1(n4441), .IN2(n8385), .QN(n5054) );
  NAND2X0 U5035 ( .IN1(n3948), .IN2(CRC_OUT_3_5), .QN(n5048) );
  NAND4X0 U5036 ( .IN1(n5055), .IN2(n5056), .IN3(n5057), .IN4(n5058), .QN(
        WX8452) );
  NAND2X0 U5037 ( .IN1(n3976), .IN2(n4804), .QN(n5058) );
  XNOR3X1 U5038 ( .IN1(n3508), .IN2(n3308), .IN3(n5059), .Q(n4804) );
  XOR2X1 U5039 ( .IN1(WX9810), .IN2(n7085), .Q(n5059) );
  NAND2X0 U5040 ( .IN1(n3885), .IN2(n5060), .QN(n5057) );
  NAND2X0 U5041 ( .IN1(n448), .IN2(n3917), .QN(n5056) );
  INVX0 U5042 ( .INP(n5061), .ZN(n448) );
  NAND2X0 U5043 ( .IN1(n4441), .IN2(n8386), .QN(n5061) );
  NAND2X0 U5044 ( .IN1(n3948), .IN2(CRC_OUT_3_6), .QN(n5055) );
  NAND4X0 U5045 ( .IN1(n5062), .IN2(n5063), .IN3(n5064), .IN4(n5065), .QN(
        WX8450) );
  NAND2X0 U5046 ( .IN1(n3976), .IN2(n4811), .QN(n5065) );
  XNOR3X1 U5047 ( .IN1(n3506), .IN2(n3309), .IN3(n5066), .Q(n4811) );
  XOR2X1 U5048 ( .IN1(WX9808), .IN2(n7086), .Q(n5066) );
  NAND2X0 U5049 ( .IN1(n3885), .IN2(n5067), .QN(n5064) );
  NAND2X0 U5050 ( .IN1(n447), .IN2(n3917), .QN(n5063) );
  INVX0 U5051 ( .INP(n5068), .ZN(n447) );
  NAND2X0 U5052 ( .IN1(n4441), .IN2(n8387), .QN(n5068) );
  NAND2X0 U5053 ( .IN1(test_so76), .IN2(n3957), .QN(n5062) );
  NAND4X0 U5054 ( .IN1(n5069), .IN2(n5070), .IN3(n5071), .IN4(n5072), .QN(
        WX8448) );
  NAND2X0 U5055 ( .IN1(n3976), .IN2(n4818), .QN(n5072) );
  XNOR3X1 U5056 ( .IN1(n3504), .IN2(n3310), .IN3(n5073), .Q(n4818) );
  XOR2X1 U5057 ( .IN1(WX9806), .IN2(n7087), .Q(n5073) );
  NAND2X0 U5058 ( .IN1(n3885), .IN2(n5074), .QN(n5071) );
  NAND2X0 U5059 ( .IN1(n446), .IN2(n3917), .QN(n5070) );
  INVX0 U5060 ( .INP(n5075), .ZN(n446) );
  NAND2X0 U5061 ( .IN1(n4440), .IN2(n8388), .QN(n5075) );
  NAND2X0 U5062 ( .IN1(n3948), .IN2(CRC_OUT_3_8), .QN(n5069) );
  NAND4X0 U5063 ( .IN1(n5076), .IN2(n5077), .IN3(n5078), .IN4(n5079), .QN(
        WX8446) );
  NAND2X0 U5064 ( .IN1(n3976), .IN2(n4825), .QN(n5079) );
  XNOR3X1 U5065 ( .IN1(n3502), .IN2(n3311), .IN3(n5080), .Q(n4825) );
  XOR2X1 U5066 ( .IN1(WX9804), .IN2(n7088), .Q(n5080) );
  NAND2X0 U5067 ( .IN1(n5081), .IN2(n3898), .QN(n5078) );
  NAND2X0 U5068 ( .IN1(n445), .IN2(n3917), .QN(n5077) );
  INVX0 U5069 ( .INP(n5082), .ZN(n445) );
  NAND2X0 U5070 ( .IN1(n4440), .IN2(n8389), .QN(n5082) );
  NAND2X0 U5071 ( .IN1(n3948), .IN2(CRC_OUT_3_9), .QN(n5076) );
  NAND4X0 U5072 ( .IN1(n5083), .IN2(n5084), .IN3(n5085), .IN4(n5086), .QN(
        WX8444) );
  NAND2X0 U5073 ( .IN1(n3976), .IN2(n4832), .QN(n5086) );
  XNOR3X1 U5074 ( .IN1(n3500), .IN2(n3312), .IN3(n5087), .Q(n4832) );
  XOR2X1 U5075 ( .IN1(WX9802), .IN2(n7089), .Q(n5087) );
  NAND2X0 U5076 ( .IN1(n3885), .IN2(n5088), .QN(n5085) );
  NAND2X0 U5077 ( .IN1(n444), .IN2(n3917), .QN(n5084) );
  INVX0 U5078 ( .INP(n5089), .ZN(n444) );
  NAND2X0 U5079 ( .IN1(n4440), .IN2(n8390), .QN(n5089) );
  NAND2X0 U5080 ( .IN1(n3948), .IN2(CRC_OUT_3_10), .QN(n5083) );
  NAND4X0 U5081 ( .IN1(n5090), .IN2(n5091), .IN3(n5092), .IN4(n5093), .QN(
        WX8442) );
  NAND2X0 U5082 ( .IN1(n3977), .IN2(n4839), .QN(n5093) );
  XNOR3X1 U5083 ( .IN1(n3416), .IN2(n3313), .IN3(n5094), .Q(n4839) );
  XOR2X1 U5084 ( .IN1(WX9800), .IN2(n7090), .Q(n5094) );
  NAND2X0 U5085 ( .IN1(n5095), .IN2(n3898), .QN(n5092) );
  NAND2X0 U5086 ( .IN1(n443), .IN2(n3917), .QN(n5091) );
  INVX0 U5087 ( .INP(n5096), .ZN(n443) );
  NAND2X0 U5088 ( .IN1(n4440), .IN2(n8391), .QN(n5096) );
  NAND2X0 U5089 ( .IN1(n3948), .IN2(CRC_OUT_3_11), .QN(n5090) );
  NAND4X0 U5090 ( .IN1(n5097), .IN2(n5098), .IN3(n5099), .IN4(n5100), .QN(
        WX8440) );
  NAND2X0 U5091 ( .IN1(n3978), .IN2(n4846), .QN(n5100) );
  XNOR3X1 U5092 ( .IN1(n3498), .IN2(n3314), .IN3(n5101), .Q(n4846) );
  XOR2X1 U5093 ( .IN1(WX9798), .IN2(n7091), .Q(n5101) );
  NAND2X0 U5094 ( .IN1(n3885), .IN2(n5102), .QN(n5099) );
  NAND2X0 U5095 ( .IN1(n442), .IN2(n3917), .QN(n5098) );
  INVX0 U5096 ( .INP(n5103), .ZN(n442) );
  NAND2X0 U5097 ( .IN1(n4440), .IN2(n8392), .QN(n5103) );
  NAND2X0 U5098 ( .IN1(n3948), .IN2(CRC_OUT_3_12), .QN(n5097) );
  NAND4X0 U5099 ( .IN1(n5104), .IN2(n5105), .IN3(n5106), .IN4(n5107), .QN(
        WX8438) );
  NAND2X0 U5100 ( .IN1(n3977), .IN2(n4853), .QN(n5107) );
  XNOR3X1 U5101 ( .IN1(n3496), .IN2(n3315), .IN3(n5108), .Q(n4853) );
  XOR2X1 U5102 ( .IN1(WX9796), .IN2(n7092), .Q(n5108) );
  NAND2X0 U5103 ( .IN1(n5109), .IN2(n3898), .QN(n5106) );
  NAND2X0 U5104 ( .IN1(n441), .IN2(n3917), .QN(n5105) );
  INVX0 U5105 ( .INP(n5110), .ZN(n441) );
  NAND2X0 U5106 ( .IN1(n4440), .IN2(n8393), .QN(n5110) );
  NAND2X0 U5107 ( .IN1(n3949), .IN2(CRC_OUT_3_13), .QN(n5104) );
  NAND4X0 U5108 ( .IN1(n5111), .IN2(n5112), .IN3(n5113), .IN4(n5114), .QN(
        WX8436) );
  NAND2X0 U5109 ( .IN1(n4860), .IN2(n3986), .QN(n5114) );
  XOR3X1 U5110 ( .IN1(n3591), .IN2(n3316), .IN3(n5115), .Q(n4860) );
  XOR2X1 U5111 ( .IN1(WX9730), .IN2(test_so86), .Q(n5115) );
  NAND2X0 U5112 ( .IN1(n3885), .IN2(n5116), .QN(n5113) );
  NAND2X0 U5113 ( .IN1(n440), .IN2(n3917), .QN(n5112) );
  INVX0 U5114 ( .INP(n5117), .ZN(n440) );
  NAND2X0 U5115 ( .IN1(n4440), .IN2(n8394), .QN(n5117) );
  NAND2X0 U5116 ( .IN1(n3949), .IN2(CRC_OUT_3_14), .QN(n5111) );
  NAND4X0 U5117 ( .IN1(n5118), .IN2(n5119), .IN3(n5120), .IN4(n5121), .QN(
        WX8434) );
  NAND2X0 U5118 ( .IN1(n3977), .IN2(n4867), .QN(n5121) );
  XNOR3X1 U5119 ( .IN1(n3494), .IN2(n3317), .IN3(n5122), .Q(n4867) );
  XOR2X1 U5120 ( .IN1(WX9792), .IN2(n7093), .Q(n5122) );
  NAND2X0 U5121 ( .IN1(n5123), .IN2(n3897), .QN(n5120) );
  NAND2X0 U5122 ( .IN1(n439), .IN2(n3917), .QN(n5119) );
  INVX0 U5123 ( .INP(n5124), .ZN(n439) );
  NAND2X0 U5124 ( .IN1(n4440), .IN2(n8395), .QN(n5124) );
  NAND2X0 U5125 ( .IN1(n3949), .IN2(CRC_OUT_3_15), .QN(n5118) );
  NAND4X0 U5126 ( .IN1(n5125), .IN2(n5126), .IN3(n5127), .IN4(n5128), .QN(
        WX8432) );
  NAND2X0 U5127 ( .IN1(n4874), .IN2(n3986), .QN(n5128) );
  XOR3X1 U5128 ( .IN1(n3102), .IN2(TM1), .IN3(n5129), .Q(n4874) );
  XNOR3X1 U5129 ( .IN1(test_so84), .IN2(n7094), .IN3(n3415), .Q(n5129) );
  NAND2X0 U5130 ( .IN1(n3885), .IN2(n5130), .QN(n5127) );
  NAND2X0 U5131 ( .IN1(n438), .IN2(n3917), .QN(n5126) );
  INVX0 U5132 ( .INP(n5131), .ZN(n438) );
  NAND2X0 U5133 ( .IN1(n4440), .IN2(n8396), .QN(n5131) );
  NAND2X0 U5134 ( .IN1(n3949), .IN2(CRC_OUT_3_16), .QN(n5125) );
  NAND4X0 U5135 ( .IN1(n5132), .IN2(n5133), .IN3(n5134), .IN4(n5135), .QN(
        WX8430) );
  NAND2X0 U5136 ( .IN1(n3977), .IN2(n4881), .QN(n5135) );
  XOR3X1 U5137 ( .IN1(n3103), .IN2(n3874), .IN3(n5136), .Q(n4881) );
  XOR3X1 U5138 ( .IN1(n7095), .IN2(n3492), .IN3(WX9852), .Q(n5136) );
  NAND2X0 U5139 ( .IN1(n3885), .IN2(n5137), .QN(n5134) );
  NAND2X0 U5140 ( .IN1(n437), .IN2(n3917), .QN(n5133) );
  INVX0 U5141 ( .INP(n5138), .ZN(n437) );
  NAND2X0 U5142 ( .IN1(test_so67), .IN2(n4464), .QN(n5138) );
  NAND2X0 U5143 ( .IN1(n3949), .IN2(CRC_OUT_3_17), .QN(n5132) );
  NAND4X0 U5144 ( .IN1(n5139), .IN2(n5140), .IN3(n5141), .IN4(n5142), .QN(
        WX8428) );
  NAND2X0 U5145 ( .IN1(n4888), .IN2(n3986), .QN(n5142) );
  XOR3X1 U5146 ( .IN1(n3105), .IN2(TM1), .IN3(n5143), .Q(n4888) );
  XNOR3X1 U5147 ( .IN1(test_so82), .IN2(n7096), .IN3(n3490), .Q(n5143) );
  NAND2X0 U5148 ( .IN1(n3885), .IN2(n5144), .QN(n5141) );
  NAND2X0 U5149 ( .IN1(WX8266), .IN2(n3917), .QN(n5140) );
  NAND2X0 U5150 ( .IN1(n3949), .IN2(CRC_OUT_3_18), .QN(n5139) );
  NAND4X0 U5151 ( .IN1(n5145), .IN2(n5146), .IN3(n5147), .IN4(n5148), .QN(
        WX8426) );
  NAND2X0 U5152 ( .IN1(n3977), .IN2(n4895), .QN(n5148) );
  XOR3X1 U5153 ( .IN1(n3106), .IN2(n3873), .IN3(n5149), .Q(n4895) );
  XOR3X1 U5154 ( .IN1(n7097), .IN2(n3488), .IN3(WX9848), .Q(n5149) );
  NAND2X0 U5155 ( .IN1(n3885), .IN2(n5150), .QN(n5147) );
  NAND2X0 U5156 ( .IN1(n435), .IN2(n3918), .QN(n5146) );
  INVX0 U5157 ( .INP(n5151), .ZN(n435) );
  NAND2X0 U5158 ( .IN1(n4439), .IN2(n8400), .QN(n5151) );
  NAND2X0 U5159 ( .IN1(n3949), .IN2(CRC_OUT_3_19), .QN(n5145) );
  NAND4X0 U5160 ( .IN1(n5152), .IN2(n5153), .IN3(n5154), .IN4(n5155), .QN(
        WX8424) );
  NAND2X0 U5161 ( .IN1(n4902), .IN2(n3986), .QN(n5155) );
  XOR3X1 U5162 ( .IN1(n3108), .IN2(TM1), .IN3(n5156), .Q(n4902) );
  XNOR3X1 U5163 ( .IN1(test_so80), .IN2(n7098), .IN3(n3487), .Q(n5156) );
  NAND2X0 U5164 ( .IN1(n3885), .IN2(n5157), .QN(n5154) );
  NAND2X0 U5165 ( .IN1(n434), .IN2(n3918), .QN(n5153) );
  INVX0 U5166 ( .INP(n5158), .ZN(n434) );
  NAND2X0 U5167 ( .IN1(n4439), .IN2(n8401), .QN(n5158) );
  NAND2X0 U5168 ( .IN1(n3949), .IN2(CRC_OUT_3_20), .QN(n5152) );
  NAND4X0 U5169 ( .IN1(n5159), .IN2(n5160), .IN3(n5161), .IN4(n5162), .QN(
        WX8422) );
  NAND2X0 U5170 ( .IN1(n3977), .IN2(n4909), .QN(n5162) );
  XOR3X1 U5171 ( .IN1(n3109), .IN2(n3872), .IN3(n5163), .Q(n4909) );
  XOR3X1 U5172 ( .IN1(n7099), .IN2(n3486), .IN3(WX9844), .Q(n5163) );
  NAND2X0 U5173 ( .IN1(n3884), .IN2(n5164), .QN(n5161) );
  NAND2X0 U5174 ( .IN1(n433), .IN2(n3918), .QN(n5160) );
  INVX0 U5175 ( .INP(n5165), .ZN(n433) );
  NAND2X0 U5176 ( .IN1(n4439), .IN2(n8402), .QN(n5165) );
  NAND2X0 U5177 ( .IN1(n3949), .IN2(CRC_OUT_3_21), .QN(n5159) );
  NAND4X0 U5178 ( .IN1(n5166), .IN2(n5167), .IN3(n5168), .IN4(n5169), .QN(
        WX8420) );
  NAND2X0 U5179 ( .IN1(n3977), .IN2(n4916), .QN(n5169) );
  XOR3X1 U5180 ( .IN1(n3111), .IN2(n3875), .IN3(n5170), .Q(n4916) );
  XOR3X1 U5181 ( .IN1(n7100), .IN2(n3484), .IN3(WX9842), .Q(n5170) );
  NAND2X0 U5182 ( .IN1(n3884), .IN2(n5171), .QN(n5168) );
  NAND2X0 U5183 ( .IN1(n432), .IN2(n3918), .QN(n5167) );
  INVX0 U5184 ( .INP(n5172), .ZN(n432) );
  NAND2X0 U5185 ( .IN1(n4439), .IN2(n8403), .QN(n5172) );
  NAND2X0 U5186 ( .IN1(n3949), .IN2(CRC_OUT_3_22), .QN(n5166) );
  NAND4X0 U5187 ( .IN1(n5173), .IN2(n5174), .IN3(n5175), .IN4(n5176), .QN(
        WX8418) );
  NAND2X0 U5188 ( .IN1(n3977), .IN2(n4923), .QN(n5176) );
  XOR3X1 U5189 ( .IN1(n3113), .IN2(n3874), .IN3(n5177), .Q(n4923) );
  XOR3X1 U5190 ( .IN1(n7101), .IN2(n3482), .IN3(WX9840), .Q(n5177) );
  NAND2X0 U5191 ( .IN1(n3884), .IN2(n5178), .QN(n5175) );
  NAND2X0 U5192 ( .IN1(n431), .IN2(n3918), .QN(n5174) );
  INVX0 U5193 ( .INP(n5179), .ZN(n431) );
  NAND2X0 U5194 ( .IN1(n4439), .IN2(n8404), .QN(n5179) );
  NAND2X0 U5195 ( .IN1(n3949), .IN2(CRC_OUT_3_23), .QN(n5173) );
  NAND4X0 U5196 ( .IN1(n5180), .IN2(n5181), .IN3(n5182), .IN4(n5183), .QN(
        WX8416) );
  NAND2X0 U5197 ( .IN1(n3977), .IN2(n4930), .QN(n5183) );
  XOR3X1 U5198 ( .IN1(n3115), .IN2(n3873), .IN3(n5184), .Q(n4930) );
  XOR3X1 U5199 ( .IN1(n7102), .IN2(n3480), .IN3(WX9838), .Q(n5184) );
  NAND2X0 U5200 ( .IN1(n3884), .IN2(n5185), .QN(n5182) );
  NAND2X0 U5201 ( .IN1(n430), .IN2(n3918), .QN(n5181) );
  INVX0 U5202 ( .INP(n5186), .ZN(n430) );
  NAND2X0 U5203 ( .IN1(n4439), .IN2(n8405), .QN(n5186) );
  NAND2X0 U5204 ( .IN1(test_so77), .IN2(n3956), .QN(n5180) );
  NAND4X0 U5205 ( .IN1(n5187), .IN2(n5188), .IN3(n5189), .IN4(n5190), .QN(
        WX8414) );
  NAND2X0 U5206 ( .IN1(n3977), .IN2(n4937), .QN(n5190) );
  XOR3X1 U5207 ( .IN1(n3117), .IN2(n3872), .IN3(n5191), .Q(n4937) );
  XOR3X1 U5208 ( .IN1(n7103), .IN2(n3478), .IN3(WX9836), .Q(n5191) );
  NAND2X0 U5209 ( .IN1(n3884), .IN2(n5192), .QN(n5189) );
  NAND2X0 U5210 ( .IN1(n429), .IN2(n3918), .QN(n5188) );
  INVX0 U5211 ( .INP(n5193), .ZN(n429) );
  NAND2X0 U5212 ( .IN1(n4439), .IN2(n8406), .QN(n5193) );
  NAND2X0 U5213 ( .IN1(n3949), .IN2(CRC_OUT_3_25), .QN(n5187) );
  NAND4X0 U5214 ( .IN1(n5194), .IN2(n5195), .IN3(n5196), .IN4(n5197), .QN(
        WX8412) );
  NAND2X0 U5215 ( .IN1(n3977), .IN2(n4944), .QN(n5197) );
  XOR3X1 U5216 ( .IN1(n3119), .IN2(n3875), .IN3(n5198), .Q(n4944) );
  XOR3X1 U5217 ( .IN1(n7104), .IN2(n3476), .IN3(WX9834), .Q(n5198) );
  NAND2X0 U5218 ( .IN1(n5199), .IN2(n3897), .QN(n5196) );
  NAND2X0 U5219 ( .IN1(n428), .IN2(n3918), .QN(n5195) );
  INVX0 U5220 ( .INP(n5200), .ZN(n428) );
  NAND2X0 U5221 ( .IN1(n4439), .IN2(n8407), .QN(n5200) );
  NAND2X0 U5222 ( .IN1(n3950), .IN2(CRC_OUT_3_26), .QN(n5194) );
  NAND4X0 U5223 ( .IN1(n5201), .IN2(n5202), .IN3(n5203), .IN4(n5204), .QN(
        WX8410) );
  NAND2X0 U5224 ( .IN1(n3978), .IN2(n4951), .QN(n5204) );
  XOR3X1 U5225 ( .IN1(n3121), .IN2(n3874), .IN3(n5205), .Q(n4951) );
  XOR3X1 U5226 ( .IN1(n7105), .IN2(n3474), .IN3(WX9832), .Q(n5205) );
  NAND2X0 U5227 ( .IN1(n3884), .IN2(n5206), .QN(n5203) );
  NAND2X0 U5228 ( .IN1(n427), .IN2(n3918), .QN(n5202) );
  INVX0 U5229 ( .INP(n5207), .ZN(n427) );
  NAND2X0 U5230 ( .IN1(n4439), .IN2(n8408), .QN(n5207) );
  NAND2X0 U5231 ( .IN1(n3950), .IN2(CRC_OUT_3_27), .QN(n5201) );
  NAND4X0 U5232 ( .IN1(n5208), .IN2(n5209), .IN3(n5210), .IN4(n5211), .QN(
        WX8408) );
  NAND2X0 U5233 ( .IN1(n3978), .IN2(n4958), .QN(n5211) );
  XOR3X1 U5234 ( .IN1(n3123), .IN2(n3873), .IN3(n5212), .Q(n4958) );
  XOR3X1 U5235 ( .IN1(n7106), .IN2(n3472), .IN3(WX9830), .Q(n5212) );
  NAND2X0 U5236 ( .IN1(n5213), .IN2(n3897), .QN(n5210) );
  NAND2X0 U5237 ( .IN1(n426), .IN2(n3918), .QN(n5209) );
  INVX0 U5238 ( .INP(n5214), .ZN(n426) );
  NAND2X0 U5239 ( .IN1(n4438), .IN2(n8409), .QN(n5214) );
  NAND2X0 U5240 ( .IN1(n3950), .IN2(CRC_OUT_3_28), .QN(n5208) );
  NAND4X0 U5241 ( .IN1(n5215), .IN2(n5216), .IN3(n5217), .IN4(n5218), .QN(
        WX8406) );
  NAND2X0 U5242 ( .IN1(n3978), .IN2(n4965), .QN(n5218) );
  XOR3X1 U5243 ( .IN1(n3125), .IN2(n3872), .IN3(n5219), .Q(n4965) );
  XOR3X1 U5244 ( .IN1(n7107), .IN2(n3470), .IN3(WX9828), .Q(n5219) );
  NAND2X0 U5245 ( .IN1(n3884), .IN2(n5220), .QN(n5217) );
  NAND2X0 U5246 ( .IN1(n425), .IN2(n3918), .QN(n5216) );
  INVX0 U5247 ( .INP(n5221), .ZN(n425) );
  NAND2X0 U5248 ( .IN1(n4438), .IN2(n8410), .QN(n5221) );
  NAND2X0 U5249 ( .IN1(n3950), .IN2(CRC_OUT_3_29), .QN(n5215) );
  NAND4X0 U5250 ( .IN1(n5222), .IN2(n5223), .IN3(n5224), .IN4(n5225), .QN(
        WX8404) );
  NAND2X0 U5251 ( .IN1(n3978), .IN2(n4972), .QN(n5225) );
  XOR3X1 U5252 ( .IN1(n3127), .IN2(n3875), .IN3(n5226), .Q(n4972) );
  XOR3X1 U5253 ( .IN1(n7108), .IN2(n3468), .IN3(WX9826), .Q(n5226) );
  NAND2X0 U5254 ( .IN1(n5227), .IN2(n3897), .QN(n5224) );
  NAND2X0 U5255 ( .IN1(n424), .IN2(n3918), .QN(n5223) );
  INVX0 U5256 ( .INP(n5228), .ZN(n424) );
  NAND2X0 U5257 ( .IN1(n4438), .IN2(n8411), .QN(n5228) );
  NAND2X0 U5258 ( .IN1(n3950), .IN2(CRC_OUT_3_30), .QN(n5222) );
  NAND4X0 U5259 ( .IN1(n5229), .IN2(n5230), .IN3(n5231), .IN4(n5232), .QN(
        WX8402) );
  NAND2X0 U5260 ( .IN1(n4979), .IN2(n3987), .QN(n5232) );
  XOR3X1 U5261 ( .IN1(n3063), .IN2(TM1), .IN3(n5233), .Q(n4979) );
  XOR3X1 U5262 ( .IN1(test_so85), .IN2(n7109), .IN3(WX9824), .Q(n5233) );
  NAND2X0 U5263 ( .IN1(n3884), .IN2(n5234), .QN(n5231) );
  NAND2X0 U5264 ( .IN1(n3950), .IN2(CRC_OUT_3_31), .QN(n5230) );
  NAND2X0 U5265 ( .IN1(n2245), .IN2(WX8243), .QN(n5229) );
  NOR2X0 U5266 ( .IN1(n4560), .IN2(WX8243), .QN(WX8304) );
  NOR2X0 U5267 ( .IN1(n5235), .IN2(n3870), .QN(WX8266) );
  NOR2X0 U5268 ( .IN1(n4560), .IN2(n5236), .QN(WX7791) );
  XOR2X1 U5269 ( .IN1(n3565), .IN2(DFF_1150_n1), .Q(n5236) );
  NOR2X0 U5270 ( .IN1(n4560), .IN2(n5237), .QN(WX7789) );
  XNOR2X1 U5271 ( .IN1(n3566), .IN2(test_so66), .Q(n5237) );
  NOR2X0 U5272 ( .IN1(n4560), .IN2(n5238), .QN(WX7787) );
  XOR2X1 U5273 ( .IN1(n3568), .IN2(DFF_1148_n1), .Q(n5238) );
  NOR2X0 U5274 ( .IN1(n4560), .IN2(n5239), .QN(WX7785) );
  XOR2X1 U5275 ( .IN1(n3570), .IN2(DFF_1147_n1), .Q(n5239) );
  NOR2X0 U5276 ( .IN1(n5235), .IN2(n5240), .QN(WX7783) );
  XOR2X1 U5277 ( .IN1(n3572), .IN2(DFF_1146_n1), .Q(n5240) );
  NOR2X0 U5278 ( .IN1(n4561), .IN2(n5241), .QN(WX7781) );
  XOR2X1 U5279 ( .IN1(n3574), .IN2(DFF_1145_n1), .Q(n5241) );
  NOR2X0 U5280 ( .IN1(n4561), .IN2(n5242), .QN(WX7779) );
  XOR2X1 U5281 ( .IN1(n3576), .IN2(DFF_1144_n1), .Q(n5242) );
  NOR2X0 U5282 ( .IN1(n4561), .IN2(n5243), .QN(WX7777) );
  XOR2X1 U5283 ( .IN1(n3578), .IN2(DFF_1143_n1), .Q(n5243) );
  NOR2X0 U5284 ( .IN1(n4561), .IN2(n5244), .QN(WX7775) );
  XOR2X1 U5285 ( .IN1(n3580), .IN2(DFF_1142_n1), .Q(n5244) );
  NOR2X0 U5286 ( .IN1(n4561), .IN2(n5245), .QN(WX7773) );
  XOR2X1 U5287 ( .IN1(n3582), .IN2(DFF_1141_n1), .Q(n5245) );
  NOR2X0 U5288 ( .IN1(n4561), .IN2(n5246), .QN(WX7771) );
  XOR2X1 U5289 ( .IN1(CRC_OUT_4_20), .IN2(test_so63), .Q(n5246) );
  NOR2X0 U5290 ( .IN1(n4561), .IN2(n5247), .QN(WX7769) );
  XOR2X1 U5291 ( .IN1(n3584), .IN2(DFF_1139_n1), .Q(n5247) );
  NOR2X0 U5292 ( .IN1(n4561), .IN2(n5248), .QN(WX7767) );
  XOR2X1 U5293 ( .IN1(n3586), .IN2(DFF_1138_n1), .Q(n5248) );
  NOR2X0 U5294 ( .IN1(n4561), .IN2(n5249), .QN(WX7765) );
  XOR2X1 U5295 ( .IN1(n3588), .IN2(DFF_1137_n1), .Q(n5249) );
  NOR2X0 U5296 ( .IN1(n4561), .IN2(n5250), .QN(WX7763) );
  XOR2X1 U5297 ( .IN1(n3590), .IN2(DFF_1136_n1), .Q(n5250) );
  NOR2X0 U5298 ( .IN1(n4561), .IN2(n5251), .QN(WX7761) );
  XOR3X1 U5299 ( .IN1(n3421), .IN2(DFF_1151_n1), .IN3(CRC_OUT_4_15), .Q(n5251)
         );
  NOR2X0 U5300 ( .IN1(n4561), .IN2(n5252), .QN(WX7759) );
  XOR2X1 U5301 ( .IN1(n3592), .IN2(DFF_1134_n1), .Q(n5252) );
  NOR2X0 U5302 ( .IN1(n4561), .IN2(n5253), .QN(WX7757) );
  XOR2X1 U5303 ( .IN1(n3594), .IN2(DFF_1133_n1), .Q(n5253) );
  NOR2X0 U5304 ( .IN1(n4561), .IN2(n5254), .QN(WX7755) );
  XNOR2X1 U5305 ( .IN1(n3596), .IN2(test_so65), .Q(n5254) );
  NOR2X0 U5306 ( .IN1(n4561), .IN2(n5255), .QN(WX7753) );
  XOR2X1 U5307 ( .IN1(n3598), .IN2(DFF_1131_n1), .Q(n5255) );
  NOR2X0 U5308 ( .IN1(n4561), .IN2(n5256), .QN(WX7751) );
  XOR3X1 U5309 ( .IN1(n3422), .IN2(DFF_1151_n1), .IN3(CRC_OUT_4_10), .Q(n5256)
         );
  NOR2X0 U5310 ( .IN1(n4562), .IN2(n5257), .QN(WX7749) );
  XOR2X1 U5311 ( .IN1(n3600), .IN2(DFF_1129_n1), .Q(n5257) );
  NOR2X0 U5312 ( .IN1(n4562), .IN2(n5258), .QN(WX7747) );
  XOR2X1 U5313 ( .IN1(n3602), .IN2(DFF_1128_n1), .Q(n5258) );
  NOR2X0 U5314 ( .IN1(n4562), .IN2(n5259), .QN(WX7745) );
  XOR2X1 U5315 ( .IN1(n3604), .IN2(DFF_1127_n1), .Q(n5259) );
  NOR2X0 U5316 ( .IN1(n4562), .IN2(n5260), .QN(WX7743) );
  XOR2X1 U5317 ( .IN1(n3606), .IN2(DFF_1126_n1), .Q(n5260) );
  NOR2X0 U5318 ( .IN1(n4562), .IN2(n5261), .QN(WX7741) );
  XOR2X1 U5319 ( .IN1(n3608), .IN2(DFF_1125_n1), .Q(n5261) );
  NOR2X0 U5320 ( .IN1(n4562), .IN2(n5262), .QN(WX7739) );
  XOR2X1 U5321 ( .IN1(n3610), .IN2(DFF_1124_n1), .Q(n5262) );
  NOR2X0 U5322 ( .IN1(n4562), .IN2(n5263), .QN(WX7737) );
  XOR3X1 U5323 ( .IN1(test_so64), .IN2(DFF_1151_n1), .IN3(DFF_1123_n1), .Q(
        n5263) );
  NOR2X0 U5324 ( .IN1(n4562), .IN2(n5264), .QN(WX7735) );
  XOR2X1 U5325 ( .IN1(n3612), .IN2(DFF_1122_n1), .Q(n5264) );
  NOR2X0 U5326 ( .IN1(n4562), .IN2(n5265), .QN(WX7733) );
  XOR2X1 U5327 ( .IN1(n3614), .IN2(DFF_1121_n1), .Q(n5265) );
  NOR2X0 U5328 ( .IN1(n4562), .IN2(n5266), .QN(WX7731) );
  XOR2X1 U5329 ( .IN1(n3616), .IN2(DFF_1120_n1), .Q(n5266) );
  NOR2X0 U5330 ( .IN1(n4562), .IN2(n5267), .QN(WX7729) );
  XOR2X1 U5331 ( .IN1(n3436), .IN2(DFF_1151_n1), .Q(n5267) );
  NAND4X0 U5332 ( .IN1(n5268), .IN2(n5269), .IN3(n5270), .IN4(n5271), .QN(
        WX7171) );
  NAND2X0 U5333 ( .IN1(n3978), .IN2(n5018), .QN(n5271) );
  XNOR3X1 U5334 ( .IN1(n3435), .IN2(n3318), .IN3(n5272), .Q(n5018) );
  XOR2X1 U5335 ( .IN1(WX8529), .IN2(n7110), .Q(n5272) );
  NAND2X0 U5336 ( .IN1(n3884), .IN2(n5273), .QN(n5270) );
  NAND2X0 U5337 ( .IN1(n376), .IN2(n3918), .QN(n5269) );
  INVX0 U5338 ( .INP(n5274), .ZN(n376) );
  NAND2X0 U5339 ( .IN1(n4438), .IN2(n8438), .QN(n5274) );
  NAND2X0 U5340 ( .IN1(n3950), .IN2(CRC_OUT_4_0), .QN(n5268) );
  NAND4X0 U5341 ( .IN1(n5275), .IN2(n5276), .IN3(n5277), .IN4(n5278), .QN(
        WX7169) );
  NAND2X0 U5342 ( .IN1(n3978), .IN2(n5025), .QN(n5278) );
  XNOR3X1 U5343 ( .IN1(n3564), .IN2(n3319), .IN3(n5279), .Q(n5025) );
  XOR2X1 U5344 ( .IN1(WX8527), .IN2(n7111), .Q(n5279) );
  NAND2X0 U5345 ( .IN1(n3884), .IN2(n5280), .QN(n5277) );
  NAND2X0 U5346 ( .IN1(n375), .IN2(n3918), .QN(n5276) );
  INVX0 U5347 ( .INP(n5281), .ZN(n375) );
  NAND2X0 U5348 ( .IN1(n4438), .IN2(n8439), .QN(n5281) );
  NAND2X0 U5349 ( .IN1(n3950), .IN2(CRC_OUT_4_1), .QN(n5275) );
  NAND4X0 U5350 ( .IN1(n5282), .IN2(n5283), .IN3(n5284), .IN4(n5285), .QN(
        WX7167) );
  NAND2X0 U5351 ( .IN1(n3978), .IN2(n5032), .QN(n5285) );
  XNOR3X1 U5352 ( .IN1(n3562), .IN2(n3320), .IN3(n5286), .Q(n5032) );
  XOR2X1 U5353 ( .IN1(WX8525), .IN2(n7112), .Q(n5286) );
  NAND2X0 U5354 ( .IN1(n3884), .IN2(n5287), .QN(n5284) );
  NAND2X0 U5355 ( .IN1(n374), .IN2(n3918), .QN(n5283) );
  INVX0 U5356 ( .INP(n5288), .ZN(n374) );
  NAND2X0 U5357 ( .IN1(n4438), .IN2(n8440), .QN(n5288) );
  NAND2X0 U5358 ( .IN1(n3950), .IN2(CRC_OUT_4_2), .QN(n5282) );
  NAND4X0 U5359 ( .IN1(n5289), .IN2(n5290), .IN3(n5291), .IN4(n5292), .QN(
        WX7165) );
  NAND2X0 U5360 ( .IN1(n3978), .IN2(n5039), .QN(n5292) );
  XNOR3X1 U5361 ( .IN1(n3560), .IN2(n3321), .IN3(n5293), .Q(n5039) );
  XOR2X1 U5362 ( .IN1(WX8523), .IN2(n7113), .Q(n5293) );
  NAND2X0 U5363 ( .IN1(n3884), .IN2(n5294), .QN(n5291) );
  NAND2X0 U5364 ( .IN1(n373), .IN2(n3918), .QN(n5290) );
  INVX0 U5365 ( .INP(n5295), .ZN(n373) );
  NAND2X0 U5366 ( .IN1(n4438), .IN2(n8441), .QN(n5295) );
  NAND2X0 U5367 ( .IN1(n3950), .IN2(CRC_OUT_4_3), .QN(n5289) );
  NAND4X0 U5368 ( .IN1(n5296), .IN2(n5297), .IN3(n5298), .IN4(n5299), .QN(
        WX7163) );
  NAND2X0 U5369 ( .IN1(n3978), .IN2(n5046), .QN(n5299) );
  XNOR3X1 U5370 ( .IN1(n3420), .IN2(n3322), .IN3(n5300), .Q(n5046) );
  XOR2X1 U5371 ( .IN1(WX8521), .IN2(n7114), .Q(n5300) );
  NAND2X0 U5372 ( .IN1(n5301), .IN2(n3897), .QN(n5298) );
  NAND2X0 U5373 ( .IN1(n372), .IN2(n3918), .QN(n5297) );
  INVX0 U5374 ( .INP(n5302), .ZN(n372) );
  NAND2X0 U5375 ( .IN1(n4438), .IN2(n8442), .QN(n5302) );
  NAND2X0 U5376 ( .IN1(n3950), .IN2(CRC_OUT_4_4), .QN(n5296) );
  NAND4X0 U5377 ( .IN1(n5303), .IN2(n5304), .IN3(n5305), .IN4(n5306), .QN(
        WX7161) );
  NAND2X0 U5378 ( .IN1(n3978), .IN2(n5053), .QN(n5306) );
  XNOR3X1 U5379 ( .IN1(n3558), .IN2(n3323), .IN3(n5307), .Q(n5053) );
  XOR2X1 U5380 ( .IN1(WX8519), .IN2(n7115), .Q(n5307) );
  NAND2X0 U5381 ( .IN1(n3883), .IN2(n5308), .QN(n5305) );
  NAND2X0 U5382 ( .IN1(WX6999), .IN2(n3919), .QN(n5304) );
  NAND2X0 U5383 ( .IN1(n3950), .IN2(CRC_OUT_4_5), .QN(n5303) );
  NAND4X0 U5384 ( .IN1(n5309), .IN2(n5310), .IN3(n5311), .IN4(n5312), .QN(
        WX7159) );
  NAND2X0 U5385 ( .IN1(n3978), .IN2(n5060), .QN(n5312) );
  XNOR3X1 U5386 ( .IN1(n3556), .IN2(n3324), .IN3(n5313), .Q(n5060) );
  XOR2X1 U5387 ( .IN1(WX8517), .IN2(n7116), .Q(n5313) );
  NAND2X0 U5388 ( .IN1(n5314), .IN2(n3897), .QN(n5311) );
  NAND2X0 U5389 ( .IN1(n370), .IN2(n3919), .QN(n5310) );
  INVX0 U5390 ( .INP(n5315), .ZN(n370) );
  NAND2X0 U5391 ( .IN1(n4438), .IN2(n8444), .QN(n5315) );
  NAND2X0 U5392 ( .IN1(n3951), .IN2(CRC_OUT_4_6), .QN(n5309) );
  NAND4X0 U5393 ( .IN1(n5316), .IN2(n5317), .IN3(n5318), .IN4(n5319), .QN(
        WX7157) );
  NAND2X0 U5394 ( .IN1(n3979), .IN2(n5067), .QN(n5319) );
  XNOR3X1 U5395 ( .IN1(n3554), .IN2(n3325), .IN3(n5320), .Q(n5067) );
  XOR2X1 U5396 ( .IN1(WX8515), .IN2(n7117), .Q(n5320) );
  NAND2X0 U5397 ( .IN1(n3883), .IN2(n5321), .QN(n5318) );
  NAND2X0 U5398 ( .IN1(n369), .IN2(n3919), .QN(n5317) );
  INVX0 U5399 ( .INP(n5322), .ZN(n369) );
  NAND2X0 U5400 ( .IN1(n4437), .IN2(n8445), .QN(n5322) );
  NAND2X0 U5401 ( .IN1(n3951), .IN2(CRC_OUT_4_7), .QN(n5316) );
  NAND4X0 U5402 ( .IN1(n5323), .IN2(n5324), .IN3(n5325), .IN4(n5326), .QN(
        WX7155) );
  NAND2X0 U5403 ( .IN1(n3979), .IN2(n5074), .QN(n5326) );
  XNOR3X1 U5404 ( .IN1(n3552), .IN2(n3326), .IN3(n5327), .Q(n5074) );
  XOR2X1 U5405 ( .IN1(WX8513), .IN2(n7118), .Q(n5327) );
  NAND2X0 U5406 ( .IN1(n5328), .IN2(n3897), .QN(n5325) );
  NAND2X0 U5407 ( .IN1(n368), .IN2(n3919), .QN(n5324) );
  INVX0 U5408 ( .INP(n5329), .ZN(n368) );
  NAND2X0 U5409 ( .IN1(n4437), .IN2(n8446), .QN(n5329) );
  NAND2X0 U5410 ( .IN1(n3951), .IN2(CRC_OUT_4_8), .QN(n5323) );
  NAND4X0 U5411 ( .IN1(n5330), .IN2(n5331), .IN3(n5332), .IN4(n5333), .QN(
        WX7153) );
  NAND2X0 U5412 ( .IN1(n5081), .IN2(n3987), .QN(n5333) );
  XOR3X1 U5413 ( .IN1(n3613), .IN2(n3327), .IN3(n5334), .Q(n5081) );
  XOR2X1 U5414 ( .IN1(WX8447), .IN2(test_so75), .Q(n5334) );
  NAND2X0 U5415 ( .IN1(n3883), .IN2(n5335), .QN(n5332) );
  NAND2X0 U5416 ( .IN1(n367), .IN2(n3919), .QN(n5331) );
  INVX0 U5417 ( .INP(n5336), .ZN(n367) );
  NAND2X0 U5418 ( .IN1(n4437), .IN2(n8447), .QN(n5336) );
  NAND2X0 U5419 ( .IN1(n3951), .IN2(CRC_OUT_4_9), .QN(n5330) );
  NAND4X0 U5420 ( .IN1(n5337), .IN2(n5338), .IN3(n5339), .IN4(n5340), .QN(
        WX7151) );
  NAND2X0 U5421 ( .IN1(n3979), .IN2(n5088), .QN(n5340) );
  XNOR3X1 U5422 ( .IN1(n3550), .IN2(n3328), .IN3(n5341), .Q(n5088) );
  XOR2X1 U5423 ( .IN1(WX8509), .IN2(n7119), .Q(n5341) );
  NAND2X0 U5424 ( .IN1(n5342), .IN2(n3896), .QN(n5339) );
  NAND2X0 U5425 ( .IN1(n366), .IN2(n3919), .QN(n5338) );
  INVX0 U5426 ( .INP(n5343), .ZN(n366) );
  NAND2X0 U5427 ( .IN1(n4437), .IN2(n8448), .QN(n5343) );
  NAND2X0 U5428 ( .IN1(n3951), .IN2(CRC_OUT_4_10), .QN(n5337) );
  NAND4X0 U5429 ( .IN1(n5344), .IN2(n5345), .IN3(n5346), .IN4(n5347), .QN(
        WX7149) );
  NAND2X0 U5430 ( .IN1(n5095), .IN2(n3987), .QN(n5347) );
  XOR3X1 U5431 ( .IN1(n3617), .IN2(n3419), .IN3(n5348), .Q(n5095) );
  XOR2X1 U5432 ( .IN1(WX8443), .IN2(test_so73), .Q(n5348) );
  NAND2X0 U5433 ( .IN1(n3883), .IN2(n5349), .QN(n5346) );
  NAND2X0 U5434 ( .IN1(n365), .IN2(n3919), .QN(n5345) );
  INVX0 U5435 ( .INP(n5350), .ZN(n365) );
  NAND2X0 U5436 ( .IN1(n4437), .IN2(n8449), .QN(n5350) );
  NAND2X0 U5437 ( .IN1(n3951), .IN2(CRC_OUT_4_11), .QN(n5344) );
  NAND4X0 U5438 ( .IN1(n5351), .IN2(n5352), .IN3(n5353), .IN4(n5354), .QN(
        WX7147) );
  NAND2X0 U5439 ( .IN1(n3979), .IN2(n5102), .QN(n5354) );
  XNOR3X1 U5440 ( .IN1(n3548), .IN2(n3329), .IN3(n5355), .Q(n5102) );
  XOR2X1 U5441 ( .IN1(WX8505), .IN2(n7120), .Q(n5355) );
  NAND2X0 U5442 ( .IN1(n3883), .IN2(n5356), .QN(n5353) );
  NAND2X0 U5443 ( .IN1(n364), .IN2(n3919), .QN(n5352) );
  INVX0 U5444 ( .INP(n5357), .ZN(n364) );
  NAND2X0 U5445 ( .IN1(test_so56), .IN2(n4464), .QN(n5357) );
  NAND2X0 U5446 ( .IN1(test_so65), .IN2(n3956), .QN(n5351) );
  NAND4X0 U5447 ( .IN1(n5358), .IN2(n5359), .IN3(n5360), .IN4(n5361), .QN(
        WX7145) );
  NAND2X0 U5448 ( .IN1(n5109), .IN2(n3987), .QN(n5361) );
  XOR3X1 U5449 ( .IN1(n3546), .IN2(n3330), .IN3(n5362), .Q(n5109) );
  XOR2X1 U5450 ( .IN1(WX8439), .IN2(test_so71), .Q(n5362) );
  NAND2X0 U5451 ( .IN1(n3883), .IN2(n5363), .QN(n5360) );
  NAND2X0 U5452 ( .IN1(n363), .IN2(n3919), .QN(n5359) );
  INVX0 U5453 ( .INP(n5364), .ZN(n363) );
  NAND2X0 U5454 ( .IN1(n4437), .IN2(n8452), .QN(n5364) );
  NAND2X0 U5455 ( .IN1(n3951), .IN2(CRC_OUT_4_13), .QN(n5358) );
  NAND4X0 U5456 ( .IN1(n5365), .IN2(n5366), .IN3(n5367), .IN4(n5368), .QN(
        WX7143) );
  NAND2X0 U5457 ( .IN1(n3979), .IN2(n5116), .QN(n5368) );
  XNOR3X1 U5458 ( .IN1(n3544), .IN2(n3331), .IN3(n5369), .Q(n5116) );
  XOR2X1 U5459 ( .IN1(WX8501), .IN2(n7121), .Q(n5369) );
  NAND2X0 U5460 ( .IN1(n3883), .IN2(n5370), .QN(n5367) );
  NAND2X0 U5461 ( .IN1(n362), .IN2(n3919), .QN(n5366) );
  INVX0 U5462 ( .INP(n5371), .ZN(n362) );
  NAND2X0 U5463 ( .IN1(n4437), .IN2(n8453), .QN(n5371) );
  NAND2X0 U5464 ( .IN1(n3951), .IN2(CRC_OUT_4_14), .QN(n5365) );
  NAND4X0 U5465 ( .IN1(n5372), .IN2(n5373), .IN3(n5374), .IN4(n5375), .QN(
        WX7141) );
  NAND2X0 U5466 ( .IN1(n5123), .IN2(n3987), .QN(n5375) );
  XOR3X1 U5467 ( .IN1(n3625), .IN2(n3543), .IN3(n5376), .Q(n5123) );
  XOR2X1 U5468 ( .IN1(WX8563), .IN2(test_so69), .Q(n5376) );
  NAND2X0 U5469 ( .IN1(n3883), .IN2(n5377), .QN(n5374) );
  NAND2X0 U5470 ( .IN1(n361), .IN2(n3919), .QN(n5373) );
  INVX0 U5471 ( .INP(n5378), .ZN(n361) );
  NAND2X0 U5472 ( .IN1(n4437), .IN2(n8454), .QN(n5378) );
  NAND2X0 U5473 ( .IN1(n3951), .IN2(CRC_OUT_4_15), .QN(n5372) );
  NAND4X0 U5474 ( .IN1(n5379), .IN2(n5380), .IN3(n5381), .IN4(n5382), .QN(
        WX7139) );
  NAND2X0 U5475 ( .IN1(n3979), .IN2(n5130), .QN(n5382) );
  XOR3X1 U5476 ( .IN1(n3129), .IN2(n3874), .IN3(n5383), .Q(n5130) );
  XOR3X1 U5477 ( .IN1(n7122), .IN2(n3418), .IN3(WX8561), .Q(n5383) );
  NAND2X0 U5478 ( .IN1(n3883), .IN2(n5384), .QN(n5381) );
  NAND2X0 U5479 ( .IN1(n360), .IN2(n3919), .QN(n5380) );
  INVX0 U5480 ( .INP(n5385), .ZN(n360) );
  NAND2X0 U5481 ( .IN1(n4437), .IN2(n8455), .QN(n5385) );
  NAND2X0 U5482 ( .IN1(n3952), .IN2(CRC_OUT_4_16), .QN(n5379) );
  NAND4X0 U5483 ( .IN1(n5386), .IN2(n5387), .IN3(n5388), .IN4(n5389), .QN(
        WX7137) );
  NAND2X0 U5484 ( .IN1(n3980), .IN2(n5137), .QN(n5389) );
  XOR3X1 U5485 ( .IN1(n3131), .IN2(n3873), .IN3(n5390), .Q(n5137) );
  XOR3X1 U5486 ( .IN1(n7123), .IN2(n3542), .IN3(WX8559), .Q(n5390) );
  NAND2X0 U5487 ( .IN1(n3883), .IN2(n5391), .QN(n5388) );
  NAND2X0 U5488 ( .IN1(n359), .IN2(n3919), .QN(n5387) );
  INVX0 U5489 ( .INP(n5392), .ZN(n359) );
  NAND2X0 U5490 ( .IN1(n4436), .IN2(n8456), .QN(n5392) );
  NAND2X0 U5491 ( .IN1(n3952), .IN2(CRC_OUT_4_17), .QN(n5386) );
  NAND4X0 U5492 ( .IN1(n5393), .IN2(n5394), .IN3(n5395), .IN4(n5396), .QN(
        WX7135) );
  NAND2X0 U5493 ( .IN1(n3979), .IN2(n5144), .QN(n5396) );
  XOR3X1 U5494 ( .IN1(n3133), .IN2(n3872), .IN3(n5397), .Q(n5144) );
  XOR3X1 U5495 ( .IN1(n7124), .IN2(n3540), .IN3(WX8557), .Q(n5397) );
  NAND2X0 U5496 ( .IN1(n3883), .IN2(n5398), .QN(n5395) );
  NAND2X0 U5497 ( .IN1(n358), .IN2(n3919), .QN(n5394) );
  INVX0 U5498 ( .INP(n5399), .ZN(n358) );
  NAND2X0 U5499 ( .IN1(n4436), .IN2(n8457), .QN(n5399) );
  NAND2X0 U5500 ( .IN1(n3952), .IN2(CRC_OUT_4_18), .QN(n5393) );
  NAND4X0 U5501 ( .IN1(n5400), .IN2(n5401), .IN3(n5402), .IN4(n5403), .QN(
        WX7133) );
  NAND2X0 U5502 ( .IN1(n3980), .IN2(n5150), .QN(n5403) );
  XOR3X1 U5503 ( .IN1(n3135), .IN2(n3875), .IN3(n5404), .Q(n5150) );
  XOR3X1 U5504 ( .IN1(n7125), .IN2(n3538), .IN3(WX8555), .Q(n5404) );
  NAND2X0 U5505 ( .IN1(n3882), .IN2(n5405), .QN(n5402) );
  NAND2X0 U5506 ( .IN1(n357), .IN2(n3919), .QN(n5401) );
  INVX0 U5507 ( .INP(n5406), .ZN(n357) );
  NAND2X0 U5508 ( .IN1(n4441), .IN2(n8458), .QN(n5406) );
  NAND2X0 U5509 ( .IN1(n3951), .IN2(CRC_OUT_4_19), .QN(n5400) );
  NAND4X0 U5510 ( .IN1(n5407), .IN2(n5408), .IN3(n5409), .IN4(n5410), .QN(
        WX7131) );
  NAND2X0 U5511 ( .IN1(n3980), .IN2(n5157), .QN(n5410) );
  XOR3X1 U5512 ( .IN1(n3137), .IN2(n3874), .IN3(n5411), .Q(n5157) );
  XOR3X1 U5513 ( .IN1(n7126), .IN2(n3536), .IN3(WX8553), .Q(n5411) );
  NAND2X0 U5514 ( .IN1(n3882), .IN2(n5412), .QN(n5409) );
  NAND2X0 U5515 ( .IN1(n356), .IN2(n3919), .QN(n5408) );
  INVX0 U5516 ( .INP(n5413), .ZN(n356) );
  NAND2X0 U5517 ( .IN1(n4459), .IN2(n8459), .QN(n5413) );
  NAND2X0 U5518 ( .IN1(n3952), .IN2(CRC_OUT_4_20), .QN(n5407) );
  NAND4X0 U5519 ( .IN1(n5414), .IN2(n5415), .IN3(n5416), .IN4(n5417), .QN(
        WX7129) );
  NAND2X0 U5520 ( .IN1(n3979), .IN2(n5164), .QN(n5417) );
  XOR3X1 U5521 ( .IN1(n3139), .IN2(n3873), .IN3(n5418), .Q(n5164) );
  XOR3X1 U5522 ( .IN1(n7127), .IN2(n3534), .IN3(WX8551), .Q(n5418) );
  NAND2X0 U5523 ( .IN1(n5419), .IN2(n3898), .QN(n5416) );
  NAND2X0 U5524 ( .IN1(n355), .IN2(n3919), .QN(n5415) );
  INVX0 U5525 ( .INP(n5420), .ZN(n355) );
  NAND2X0 U5526 ( .IN1(n4462), .IN2(n8460), .QN(n5420) );
  NAND2X0 U5527 ( .IN1(n3952), .IN2(CRC_OUT_4_21), .QN(n5414) );
  NAND4X0 U5528 ( .IN1(n5421), .IN2(n5422), .IN3(n5423), .IN4(n5424), .QN(
        WX7127) );
  NAND2X0 U5529 ( .IN1(n3980), .IN2(n5171), .QN(n5424) );
  XOR3X1 U5530 ( .IN1(n3141), .IN2(n3872), .IN3(n5425), .Q(n5171) );
  XOR3X1 U5531 ( .IN1(n7128), .IN2(n3532), .IN3(WX8549), .Q(n5425) );
  NAND2X0 U5532 ( .IN1(n3882), .IN2(n5426), .QN(n5423) );
  NAND2X0 U5533 ( .IN1(n354), .IN2(n3920), .QN(n5422) );
  INVX0 U5534 ( .INP(n5427), .ZN(n354) );
  NAND2X0 U5535 ( .IN1(n4461), .IN2(n8461), .QN(n5427) );
  NAND2X0 U5536 ( .IN1(n3952), .IN2(CRC_OUT_4_22), .QN(n5421) );
  NAND4X0 U5537 ( .IN1(n5428), .IN2(n5429), .IN3(n5430), .IN4(n5431), .QN(
        WX7125) );
  NAND2X0 U5538 ( .IN1(n3979), .IN2(n5178), .QN(n5431) );
  XOR3X1 U5539 ( .IN1(n3143), .IN2(n3875), .IN3(n5432), .Q(n5178) );
  XOR3X1 U5540 ( .IN1(n7129), .IN2(n3530), .IN3(WX8547), .Q(n5432) );
  NAND2X0 U5541 ( .IN1(n5433), .IN2(n3899), .QN(n5430) );
  NAND2X0 U5542 ( .IN1(n353), .IN2(n3920), .QN(n5429) );
  INVX0 U5543 ( .INP(n5434), .ZN(n353) );
  NAND2X0 U5544 ( .IN1(n4462), .IN2(n8462), .QN(n5434) );
  NAND2X0 U5545 ( .IN1(n3952), .IN2(CRC_OUT_4_23), .QN(n5428) );
  NAND4X0 U5546 ( .IN1(n5435), .IN2(n5436), .IN3(n5437), .IN4(n5438), .QN(
        WX7123) );
  NAND2X0 U5547 ( .IN1(n3980), .IN2(n5185), .QN(n5438) );
  XOR3X1 U5548 ( .IN1(n3145), .IN2(n3874), .IN3(n5439), .Q(n5185) );
  XOR3X1 U5549 ( .IN1(n7130), .IN2(n3528), .IN3(WX8545), .Q(n5439) );
  NAND2X0 U5550 ( .IN1(n3882), .IN2(n5440), .QN(n5437) );
  NAND2X0 U5551 ( .IN1(n352), .IN2(n3920), .QN(n5436) );
  INVX0 U5552 ( .INP(n5441), .ZN(n352) );
  NAND2X0 U5553 ( .IN1(n4462), .IN2(n8463), .QN(n5441) );
  NAND2X0 U5554 ( .IN1(n3952), .IN2(CRC_OUT_4_24), .QN(n5435) );
  NAND4X0 U5555 ( .IN1(n5442), .IN2(n5443), .IN3(n5444), .IN4(n5445), .QN(
        WX7121) );
  NAND2X0 U5556 ( .IN1(n3980), .IN2(n5192), .QN(n5445) );
  XOR3X1 U5557 ( .IN1(n3147), .IN2(n3873), .IN3(n5446), .Q(n5192) );
  XOR3X1 U5558 ( .IN1(n7131), .IN2(n3526), .IN3(WX8543), .Q(n5446) );
  NAND2X0 U5559 ( .IN1(n5447), .IN2(n3899), .QN(n5444) );
  NAND2X0 U5560 ( .IN1(n351), .IN2(n3920), .QN(n5443) );
  INVX0 U5561 ( .INP(n5448), .ZN(n351) );
  NAND2X0 U5562 ( .IN1(n4461), .IN2(n8464), .QN(n5448) );
  NAND2X0 U5563 ( .IN1(n3952), .IN2(CRC_OUT_4_25), .QN(n5442) );
  NAND4X0 U5564 ( .IN1(n5449), .IN2(n5450), .IN3(n5451), .IN4(n5452), .QN(
        WX7119) );
  NAND2X0 U5565 ( .IN1(n5199), .IN2(n3986), .QN(n5452) );
  XOR3X1 U5566 ( .IN1(n3149), .IN2(TM1), .IN3(n5453), .Q(n5199) );
  XOR3X1 U5567 ( .IN1(test_so74), .IN2(n7132), .IN3(WX8541), .Q(n5453) );
  NAND2X0 U5568 ( .IN1(n3882), .IN2(n5454), .QN(n5451) );
  NAND2X0 U5569 ( .IN1(n350), .IN2(n3920), .QN(n5450) );
  INVX0 U5570 ( .INP(n5455), .ZN(n350) );
  NAND2X0 U5571 ( .IN1(n4462), .IN2(n8465), .QN(n5455) );
  NAND2X0 U5572 ( .IN1(n3953), .IN2(CRC_OUT_4_26), .QN(n5449) );
  NAND4X0 U5573 ( .IN1(n5456), .IN2(n5457), .IN3(n5458), .IN4(n5459), .QN(
        WX7117) );
  NAND2X0 U5574 ( .IN1(n3981), .IN2(n5206), .QN(n5459) );
  XOR3X1 U5575 ( .IN1(n3150), .IN2(n3872), .IN3(n5460), .Q(n5206) );
  XOR3X1 U5576 ( .IN1(n7133), .IN2(n3524), .IN3(WX8539), .Q(n5460) );
  NAND2X0 U5577 ( .IN1(n5461), .IN2(n3899), .QN(n5458) );
  NAND2X0 U5578 ( .IN1(n349), .IN2(n3920), .QN(n5457) );
  INVX0 U5579 ( .INP(n5462), .ZN(n349) );
  NAND2X0 U5580 ( .IN1(n4461), .IN2(n8466), .QN(n5462) );
  NAND2X0 U5581 ( .IN1(n3953), .IN2(CRC_OUT_4_27), .QN(n5456) );
  NAND4X0 U5582 ( .IN1(n5463), .IN2(n5464), .IN3(n5465), .IN4(n5466), .QN(
        WX7115) );
  NAND2X0 U5583 ( .IN1(n5213), .IN2(n3986), .QN(n5466) );
  XOR3X1 U5584 ( .IN1(n3152), .IN2(TM1), .IN3(n5467), .Q(n5213) );
  XNOR3X1 U5585 ( .IN1(test_so72), .IN2(n7134), .IN3(n3523), .Q(n5467) );
  NAND2X0 U5586 ( .IN1(n3882), .IN2(n5468), .QN(n5465) );
  NAND2X0 U5587 ( .IN1(n348), .IN2(n3920), .QN(n5464) );
  INVX0 U5588 ( .INP(n5469), .ZN(n348) );
  NAND2X0 U5589 ( .IN1(n4462), .IN2(n8467), .QN(n5469) );
  NAND2X0 U5590 ( .IN1(n3953), .IN2(CRC_OUT_4_28), .QN(n5463) );
  NAND4X0 U5591 ( .IN1(n5470), .IN2(n5471), .IN3(n5472), .IN4(n5473), .QN(
        WX7113) );
  NAND2X0 U5592 ( .IN1(n3980), .IN2(n5220), .QN(n5473) );
  XOR3X1 U5593 ( .IN1(n3153), .IN2(n3875), .IN3(n5474), .Q(n5220) );
  XOR3X1 U5594 ( .IN1(n7135), .IN2(n3522), .IN3(WX8535), .Q(n5474) );
  NAND2X0 U5595 ( .IN1(n3882), .IN2(n5475), .QN(n5472) );
  NAND2X0 U5596 ( .IN1(n347), .IN2(n3920), .QN(n5471) );
  INVX0 U5597 ( .INP(n5476), .ZN(n347) );
  NAND2X0 U5598 ( .IN1(test_so55), .IN2(n4463), .QN(n5476) );
  NAND2X0 U5599 ( .IN1(test_so66), .IN2(n3957), .QN(n5470) );
  NAND4X0 U5600 ( .IN1(n5477), .IN2(n5478), .IN3(n5479), .IN4(n5480), .QN(
        WX7111) );
  NAND2X0 U5601 ( .IN1(n5227), .IN2(n3985), .QN(n5480) );
  XOR3X1 U5602 ( .IN1(n3155), .IN2(TM1), .IN3(n5481), .Q(n5227) );
  XNOR3X1 U5603 ( .IN1(test_so70), .IN2(n7136), .IN3(n3520), .Q(n5481) );
  NAND2X0 U5604 ( .IN1(n3882), .IN2(n5482), .QN(n5479) );
  NAND2X0 U5605 ( .IN1(n346), .IN2(n3920), .QN(n5478) );
  INVX0 U5606 ( .INP(n5483), .ZN(n346) );
  NAND2X0 U5607 ( .IN1(n4460), .IN2(n8470), .QN(n5483) );
  NAND2X0 U5608 ( .IN1(n3953), .IN2(CRC_OUT_4_30), .QN(n5477) );
  NAND4X0 U5609 ( .IN1(n5484), .IN2(n5485), .IN3(n5486), .IN4(n5487), .QN(
        WX7109) );
  NAND2X0 U5610 ( .IN1(n3980), .IN2(n5234), .QN(n5487) );
  XOR3X1 U5611 ( .IN1(n3064), .IN2(n3874), .IN3(n5488), .Q(n5234) );
  XOR3X1 U5612 ( .IN1(n7137), .IN2(n3518), .IN3(WX8531), .Q(n5488) );
  NAND2X0 U5613 ( .IN1(n3882), .IN2(n5489), .QN(n5486) );
  NAND2X0 U5614 ( .IN1(n3952), .IN2(CRC_OUT_4_31), .QN(n5485) );
  NAND2X0 U5615 ( .IN1(n2245), .IN2(WX6950), .QN(n5484) );
  NAND4X0 U5616 ( .IN1(n5490), .IN2(n5491), .IN3(n5492), .IN4(n5493), .QN(
        WX706) );
  NAND2X0 U5617 ( .IN1(n5494), .IN2(n3985), .QN(n5493) );
  NAND2X0 U5618 ( .IN1(n3882), .IN2(n5495), .QN(n5492) );
  NAND2X0 U5619 ( .IN1(WX544), .IN2(n3920), .QN(n5491) );
  NAND2X0 U5620 ( .IN1(n3953), .IN2(CRC_OUT_9_0), .QN(n5490) );
  NAND4X0 U5621 ( .IN1(n5496), .IN2(n5497), .IN3(n5498), .IN4(n5499), .QN(
        WX704) );
  NAND2X0 U5622 ( .IN1(n3981), .IN2(n5500), .QN(n5499) );
  NAND2X0 U5623 ( .IN1(n3882), .IN2(n5501), .QN(n5498) );
  NAND2X0 U5624 ( .IN1(WX542), .IN2(n3920), .QN(n5497) );
  NAND2X0 U5625 ( .IN1(test_so9), .IN2(n3957), .QN(n5496) );
  NAND4X0 U5626 ( .IN1(n5502), .IN2(n5503), .IN3(n5504), .IN4(n5505), .QN(
        WX702) );
  NAND2X0 U5627 ( .IN1(n3981), .IN2(n5506), .QN(n5505) );
  NAND2X0 U5628 ( .IN1(n5507), .IN2(n3900), .QN(n5504) );
  NAND2X0 U5629 ( .IN1(WX540), .IN2(n3920), .QN(n5503) );
  NAND2X0 U5630 ( .IN1(n3953), .IN2(CRC_OUT_9_2), .QN(n5502) );
  NOR2X0 U5631 ( .IN1(n4562), .IN2(WX6950), .QN(WX7011) );
  NAND4X0 U5632 ( .IN1(n5508), .IN2(n5509), .IN3(n5510), .IN4(n5511), .QN(
        WX700) );
  NAND2X0 U5633 ( .IN1(n3981), .IN2(n5512), .QN(n5511) );
  NAND2X0 U5634 ( .IN1(n3882), .IN2(n5513), .QN(n5510) );
  NAND2X0 U5635 ( .IN1(WX538), .IN2(n3920), .QN(n5509) );
  NAND2X0 U5636 ( .IN1(n3952), .IN2(CRC_OUT_9_3), .QN(n5508) );
  NOR2X0 U5637 ( .IN1(n5235), .IN2(n3871), .QN(WX6999) );
  NAND4X0 U5638 ( .IN1(n5514), .IN2(n5515), .IN3(n5516), .IN4(n5517), .QN(
        WX698) );
  NAND2X0 U5639 ( .IN1(n5518), .IN2(n3984), .QN(n5517) );
  NAND2X0 U5640 ( .IN1(n3881), .IN2(n5519), .QN(n5516) );
  NAND2X0 U5641 ( .IN1(WX536), .IN2(n3920), .QN(n5515) );
  NAND2X0 U5642 ( .IN1(n3953), .IN2(CRC_OUT_9_4), .QN(n5514) );
  NAND4X0 U5643 ( .IN1(n5520), .IN2(n5521), .IN3(n5522), .IN4(n5523), .QN(
        WX696) );
  NAND2X0 U5644 ( .IN1(n3981), .IN2(n5524), .QN(n5523) );
  NAND2X0 U5645 ( .IN1(n3881), .IN2(n5525), .QN(n5522) );
  NAND2X0 U5646 ( .IN1(WX534), .IN2(n3920), .QN(n5521) );
  NAND2X0 U5647 ( .IN1(n3954), .IN2(CRC_OUT_9_5), .QN(n5520) );
  NAND4X0 U5648 ( .IN1(n5526), .IN2(n5527), .IN3(n5528), .IN4(n5529), .QN(
        WX694) );
  NAND2X0 U5649 ( .IN1(n3980), .IN2(n5530), .QN(n5529) );
  NAND2X0 U5650 ( .IN1(n5531), .IN2(n3900), .QN(n5528) );
  NAND2X0 U5651 ( .IN1(WX532), .IN2(n3920), .QN(n5527) );
  NAND2X0 U5652 ( .IN1(n3953), .IN2(CRC_OUT_9_6), .QN(n5526) );
  NAND4X0 U5653 ( .IN1(n5532), .IN2(n5533), .IN3(n5534), .IN4(n5535), .QN(
        WX692) );
  NAND2X0 U5654 ( .IN1(n3981), .IN2(n5536), .QN(n5535) );
  NAND2X0 U5655 ( .IN1(n3881), .IN2(n5537), .QN(n5534) );
  NAND2X0 U5656 ( .IN1(WX530), .IN2(n3920), .QN(n5533) );
  NAND2X0 U5657 ( .IN1(n3954), .IN2(CRC_OUT_9_7), .QN(n5532) );
  NAND4X0 U5658 ( .IN1(n5538), .IN2(n5539), .IN3(n5540), .IN4(n5541), .QN(
        WX690) );
  NAND2X0 U5659 ( .IN1(n3979), .IN2(n5542), .QN(n5541) );
  NAND2X0 U5660 ( .IN1(n3881), .IN2(n5543), .QN(n5540) );
  NAND2X0 U5661 ( .IN1(WX528), .IN2(n3921), .QN(n5539) );
  NAND2X0 U5662 ( .IN1(n3952), .IN2(CRC_OUT_9_8), .QN(n5538) );
  NAND4X0 U5663 ( .IN1(n5544), .IN2(n5545), .IN3(n5546), .IN4(n5547), .QN(
        WX688) );
  NAND2X0 U5664 ( .IN1(n3980), .IN2(n5548), .QN(n5547) );
  NAND2X0 U5665 ( .IN1(n3881), .IN2(n5549), .QN(n5546) );
  NAND2X0 U5666 ( .IN1(WX526), .IN2(n3921), .QN(n5545) );
  NAND2X0 U5667 ( .IN1(n3954), .IN2(CRC_OUT_9_9), .QN(n5544) );
  NAND4X0 U5668 ( .IN1(n5550), .IN2(n5551), .IN3(n5552), .IN4(n5553), .QN(
        WX686) );
  NAND2X0 U5669 ( .IN1(n5554), .IN2(n3984), .QN(n5553) );
  NAND2X0 U5670 ( .IN1(n5555), .IN2(n3900), .QN(n5552) );
  NAND2X0 U5671 ( .IN1(WX524), .IN2(n3921), .QN(n5551) );
  NAND2X0 U5672 ( .IN1(n3954), .IN2(CRC_OUT_9_10), .QN(n5550) );
  NAND4X0 U5673 ( .IN1(n5556), .IN2(n5557), .IN3(n5558), .IN4(n5559), .QN(
        WX684) );
  NAND2X0 U5674 ( .IN1(n3980), .IN2(n5560), .QN(n5559) );
  NAND2X0 U5675 ( .IN1(n3881), .IN2(n5561), .QN(n5558) );
  NAND2X0 U5676 ( .IN1(WX522), .IN2(n3921), .QN(n5557) );
  NAND2X0 U5677 ( .IN1(n3954), .IN2(CRC_OUT_9_11), .QN(n5556) );
  NAND4X0 U5678 ( .IN1(n5562), .IN2(n5563), .IN3(n5564), .IN4(n5565), .QN(
        WX682) );
  NAND2X0 U5679 ( .IN1(n3980), .IN2(n5566), .QN(n5565) );
  NAND2X0 U5680 ( .IN1(n3881), .IN2(n5567), .QN(n5564) );
  NAND2X0 U5681 ( .IN1(WX520), .IN2(n3921), .QN(n5563) );
  NAND2X0 U5682 ( .IN1(n3953), .IN2(CRC_OUT_9_12), .QN(n5562) );
  NAND4X0 U5683 ( .IN1(n5568), .IN2(n5569), .IN3(n5570), .IN4(n5571), .QN(
        WX680) );
  NAND2X0 U5684 ( .IN1(n3979), .IN2(n5572), .QN(n5571) );
  NAND2X0 U5685 ( .IN1(n3881), .IN2(n5573), .QN(n5570) );
  NAND2X0 U5686 ( .IN1(WX518), .IN2(n3921), .QN(n5569) );
  NAND2X0 U5687 ( .IN1(n3951), .IN2(CRC_OUT_9_13), .QN(n5568) );
  NAND4X0 U5688 ( .IN1(n5574), .IN2(n5575), .IN3(n5576), .IN4(n5577), .QN(
        WX678) );
  NAND2X0 U5689 ( .IN1(n5578), .IN2(n3983), .QN(n5577) );
  NAND2X0 U5690 ( .IN1(n3881), .IN2(n5579), .QN(n5576) );
  NAND2X0 U5691 ( .IN1(WX516), .IN2(n3921), .QN(n5575) );
  NAND2X0 U5692 ( .IN1(n3953), .IN2(CRC_OUT_9_14), .QN(n5574) );
  NAND4X0 U5693 ( .IN1(n5580), .IN2(n5581), .IN3(n5582), .IN4(n5583), .QN(
        WX676) );
  NAND2X0 U5694 ( .IN1(n3979), .IN2(n5584), .QN(n5583) );
  NAND2X0 U5695 ( .IN1(n3881), .IN2(n5585), .QN(n5582) );
  NAND2X0 U5696 ( .IN1(WX514), .IN2(n3921), .QN(n5581) );
  NAND2X0 U5697 ( .IN1(n3955), .IN2(CRC_OUT_9_15), .QN(n5580) );
  NAND4X0 U5698 ( .IN1(n5586), .IN2(n5587), .IN3(n5588), .IN4(n5589), .QN(
        WX674) );
  NAND2X0 U5699 ( .IN1(n3969), .IN2(n5590), .QN(n5589) );
  NAND2X0 U5700 ( .IN1(n5591), .IN2(n3898), .QN(n5588) );
  NAND2X0 U5701 ( .IN1(WX512), .IN2(n3921), .QN(n5587) );
  NAND2X0 U5702 ( .IN1(n3954), .IN2(CRC_OUT_9_16), .QN(n5586) );
  NAND4X0 U5703 ( .IN1(n5592), .IN2(n5593), .IN3(n5594), .IN4(n5595), .QN(
        WX672) );
  NAND2X0 U5704 ( .IN1(n3965), .IN2(n5596), .QN(n5595) );
  NAND2X0 U5705 ( .IN1(n3881), .IN2(n5597), .QN(n5594) );
  NAND2X0 U5706 ( .IN1(WX510), .IN2(n3921), .QN(n5593) );
  NAND2X0 U5707 ( .IN1(n3955), .IN2(CRC_OUT_9_17), .QN(n5592) );
  NAND4X0 U5708 ( .IN1(n5598), .IN2(n5599), .IN3(n5600), .IN4(n5601), .QN(
        WX670) );
  NAND2X0 U5709 ( .IN1(n5602), .IN2(n3983), .QN(n5601) );
  NAND2X0 U5710 ( .IN1(n3881), .IN2(n5603), .QN(n5600) );
  NAND2X0 U5711 ( .IN1(WX508), .IN2(n3921), .QN(n5599) );
  NAND2X0 U5712 ( .IN1(n3953), .IN2(CRC_OUT_9_18), .QN(n5598) );
  NAND4X0 U5713 ( .IN1(n5604), .IN2(n5605), .IN3(n5606), .IN4(n5607), .QN(
        WX668) );
  NAND2X0 U5714 ( .IN1(n3965), .IN2(n5608), .QN(n5607) );
  NAND2X0 U5715 ( .IN1(n3880), .IN2(n5609), .QN(n5606) );
  NAND2X0 U6483 ( .IN1(WX506), .IN2(n3921), .QN(n5605) );
  NAND2X0 U6484 ( .IN1(test_so10), .IN2(n3956), .QN(n5604) );
  NAND4X0 U6485 ( .IN1(n5610), .IN2(n5611), .IN3(n5612), .IN4(n5613), .QN(
        WX666) );
  NAND2X0 U6486 ( .IN1(n3965), .IN2(n5614), .QN(n5613) );
  NAND2X0 U6487 ( .IN1(n5615), .IN2(n3896), .QN(n5612) );
  NAND2X0 U6488 ( .IN1(WX504), .IN2(n3921), .QN(n5611) );
  NAND2X0 U6489 ( .IN1(n3955), .IN2(CRC_OUT_9_20), .QN(n5610) );
  NAND4X0 U6490 ( .IN1(n5616), .IN2(n5617), .IN3(n5618), .IN4(n5619), .QN(
        WX664) );
  NAND2X0 U6491 ( .IN1(n3965), .IN2(n5620), .QN(n5619) );
  NAND2X0 U6492 ( .IN1(n3880), .IN2(n5621), .QN(n5618) );
  NAND2X0 U6493 ( .IN1(WX502), .IN2(n3921), .QN(n5617) );
  NAND2X0 U6494 ( .IN1(n3954), .IN2(CRC_OUT_9_21), .QN(n5616) );
  NAND4X0 U6495 ( .IN1(n5622), .IN2(n5623), .IN3(n5624), .IN4(n5625), .QN(
        WX662) );
  NAND2X0 U6496 ( .IN1(n5626), .IN2(n3984), .QN(n5625) );
  NAND2X0 U6497 ( .IN1(n3880), .IN2(n5627), .QN(n5624) );
  NAND2X0 U6498 ( .IN1(WX500), .IN2(n3921), .QN(n5623) );
  NAND2X0 U6499 ( .IN1(n3955), .IN2(CRC_OUT_9_22), .QN(n5622) );
  NAND4X0 U6500 ( .IN1(n5628), .IN2(n5629), .IN3(n5630), .IN4(n5631), .QN(
        WX660) );
  NAND2X0 U6501 ( .IN1(n3965), .IN2(n5632), .QN(n5631) );
  NAND2X0 U6502 ( .IN1(n3880), .IN2(n5633), .QN(n5630) );
  NAND2X0 U6503 ( .IN1(WX498), .IN2(n3921), .QN(n5629) );
  NAND2X0 U6504 ( .IN1(n3953), .IN2(CRC_OUT_9_23), .QN(n5628) );
  NAND4X0 U6505 ( .IN1(n5634), .IN2(n5635), .IN3(n5636), .IN4(n5637), .QN(
        WX658) );
  NAND2X0 U6506 ( .IN1(n3965), .IN2(n5638), .QN(n5637) );
  NAND2X0 U6507 ( .IN1(n5639), .IN2(n3896), .QN(n5636) );
  NAND2X0 U6508 ( .IN1(WX496), .IN2(n3921), .QN(n5635) );
  NAND2X0 U6509 ( .IN1(n3955), .IN2(CRC_OUT_9_24), .QN(n5634) );
  NAND4X0 U6510 ( .IN1(n5640), .IN2(n5641), .IN3(n5642), .IN4(n5643), .QN(
        WX656) );
  NAND2X0 U6511 ( .IN1(n3965), .IN2(n5644), .QN(n5643) );
  NAND2X0 U6512 ( .IN1(n3880), .IN2(n5645), .QN(n5642) );
  NAND2X0 U6513 ( .IN1(WX494), .IN2(n3922), .QN(n5641) );
  NAND2X0 U6514 ( .IN1(n3954), .IN2(CRC_OUT_9_25), .QN(n5640) );
  NAND4X0 U6515 ( .IN1(n5646), .IN2(n5647), .IN3(n5648), .IN4(n5649), .QN(
        WX654) );
  NAND2X0 U6516 ( .IN1(n3965), .IN2(n5650), .QN(n5649) );
  NAND2X0 U6517 ( .IN1(n3880), .IN2(n5651), .QN(n5648) );
  NAND2X0 U6518 ( .IN1(WX492), .IN2(n3922), .QN(n5647) );
  NAND2X0 U6519 ( .IN1(n3955), .IN2(CRC_OUT_9_26), .QN(n5646) );
  NAND4X0 U6520 ( .IN1(n5652), .IN2(n5653), .IN3(n5654), .IN4(n5655), .QN(
        WX652) );
  NAND2X0 U6521 ( .IN1(n3965), .IN2(n5656), .QN(n5655) );
  NAND2X0 U6522 ( .IN1(n3880), .IN2(n5657), .QN(n5654) );
  NAND2X0 U6523 ( .IN1(WX490), .IN2(n3922), .QN(n5653) );
  NAND2X0 U6524 ( .IN1(n3954), .IN2(CRC_OUT_9_27), .QN(n5652) );
  NAND4X0 U6525 ( .IN1(n5658), .IN2(n5659), .IN3(n5660), .IN4(n5661), .QN(
        WX650) );
  NAND2X0 U6526 ( .IN1(n5662), .IN2(n3984), .QN(n5661) );
  NAND2X0 U6527 ( .IN1(n5663), .IN2(n3896), .QN(n5660) );
  NAND2X0 U6528 ( .IN1(WX488), .IN2(n3922), .QN(n5659) );
  NAND2X0 U6529 ( .IN1(n3954), .IN2(CRC_OUT_9_28), .QN(n5658) );
  NOR2X0 U6530 ( .IN1(n4562), .IN2(n5664), .QN(WX6498) );
  XOR2X1 U6531 ( .IN1(n3618), .IN2(DFF_958_n1), .Q(n5664) );
  NOR2X0 U6532 ( .IN1(n4562), .IN2(n5665), .QN(WX6496) );
  XOR2X1 U6533 ( .IN1(n3620), .IN2(DFF_957_n1), .Q(n5665) );
  NOR2X0 U6534 ( .IN1(n4562), .IN2(n5666), .QN(WX6494) );
  XOR2X1 U6535 ( .IN1(n3621), .IN2(DFF_956_n1), .Q(n5666) );
  NOR2X0 U6536 ( .IN1(n4562), .IN2(n5667), .QN(WX6492) );
  XOR2X1 U6537 ( .IN1(n3622), .IN2(DFF_955_n1), .Q(n5667) );
  NOR2X0 U6538 ( .IN1(n4563), .IN2(n5668), .QN(WX6490) );
  XOR2X1 U6539 ( .IN1(n3624), .IN2(DFF_954_n1), .Q(n5668) );
  NOR2X0 U6540 ( .IN1(n4563), .IN2(n5669), .QN(WX6488) );
  XOR2X1 U6541 ( .IN1(n3626), .IN2(DFF_953_n1), .Q(n5669) );
  NOR2X0 U6542 ( .IN1(n4563), .IN2(n5670), .QN(WX6486) );
  XOR2X1 U6543 ( .IN1(n3628), .IN2(DFF_952_n1), .Q(n5670) );
  NOR2X0 U6544 ( .IN1(n5235), .IN2(n5671), .QN(WX6484) );
  XOR2X1 U6545 ( .IN1(n3630), .IN2(DFF_951_n1), .Q(n5671) );
  INVX0 U6546 ( .INP(n5672), .ZN(n5235) );
  NOR2X0 U6547 ( .IN1(n4563), .IN2(Tj_Trigger), .QN(n5672) );
  NOR2X0 U6548 ( .IN1(n4563), .IN2(n5673), .QN(WX6482) );
  XOR2X1 U6549 ( .IN1(n3632), .IN2(DFF_950_n1), .Q(n5673) );
  NOR2X0 U6550 ( .IN1(n4563), .IN2(n5674), .QN(WX6480) );
  XOR2X1 U6551 ( .IN1(n3634), .IN2(DFF_949_n1), .Q(n5674) );
  NAND4X0 U6552 ( .IN1(n5675), .IN2(n5676), .IN3(n5677), .IN4(n5678), .QN(
        WX648) );
  NAND2X0 U6553 ( .IN1(n3965), .IN2(n5679), .QN(n5678) );
  NAND2X0 U6554 ( .IN1(n3880), .IN2(n5680), .QN(n5677) );
  NAND2X0 U6555 ( .IN1(WX486), .IN2(n3922), .QN(n5676) );
  NAND2X0 U6556 ( .IN1(n3955), .IN2(CRC_OUT_9_29), .QN(n5675) );
  NOR2X0 U6557 ( .IN1(n4563), .IN2(n5681), .QN(WX6478) );
  XOR2X1 U6558 ( .IN1(n3636), .IN2(DFF_948_n1), .Q(n5681) );
  NOR2X0 U6559 ( .IN1(n4563), .IN2(n5682), .QN(WX6476) );
  XOR2X1 U6560 ( .IN1(n3638), .IN2(DFF_947_n1), .Q(n5682) );
  NOR2X0 U6561 ( .IN1(n4563), .IN2(n5683), .QN(WX6474) );
  XOR2X1 U6562 ( .IN1(n3640), .IN2(DFF_946_n1), .Q(n5683) );
  NOR2X0 U6563 ( .IN1(n4563), .IN2(n5684), .QN(WX6472) );
  XNOR2X1 U6564 ( .IN1(n3642), .IN2(test_so54), .Q(n5684) );
  NOR2X0 U6565 ( .IN1(n4563), .IN2(n5685), .QN(WX6470) );
  XOR2X1 U6566 ( .IN1(n3643), .IN2(DFF_944_n1), .Q(n5685) );
  NOR2X0 U6567 ( .IN1(n4563), .IN2(n5686), .QN(WX6468) );
  XOR3X1 U6568 ( .IN1(test_so52), .IN2(DFF_959_n1), .IN3(DFF_943_n1), .Q(n5686) );
  NOR2X0 U6569 ( .IN1(n4563), .IN2(n5687), .QN(WX6466) );
  XOR2X1 U6570 ( .IN1(n3644), .IN2(DFF_942_n1), .Q(n5687) );
  NOR2X0 U6571 ( .IN1(n4563), .IN2(n5688), .QN(WX6464) );
  XOR2X1 U6572 ( .IN1(n3646), .IN2(DFF_941_n1), .Q(n5688) );
  NOR2X0 U6573 ( .IN1(n4563), .IN2(n5689), .QN(WX6462) );
  XOR2X1 U6574 ( .IN1(n3648), .IN2(DFF_940_n1), .Q(n5689) );
  NOR2X0 U6575 ( .IN1(n4564), .IN2(n5690), .QN(WX6460) );
  XOR2X1 U6576 ( .IN1(n3650), .IN2(DFF_939_n1), .Q(n5690) );
  NAND4X0 U6577 ( .IN1(n5691), .IN2(n5692), .IN3(n5693), .IN4(n5694), .QN(
        WX646) );
  NAND2X0 U6578 ( .IN1(n3965), .IN2(n5695), .QN(n5694) );
  NAND2X0 U6579 ( .IN1(n3880), .IN2(n5696), .QN(n5693) );
  NAND2X0 U6580 ( .IN1(WX484), .IN2(n3922), .QN(n5692) );
  NAND2X0 U6581 ( .IN1(n3956), .IN2(CRC_OUT_9_30), .QN(n5691) );
  NOR2X0 U6582 ( .IN1(n4564), .IN2(n5697), .QN(WX6458) );
  XOR3X1 U6583 ( .IN1(n3423), .IN2(DFF_959_n1), .IN3(CRC_OUT_5_10), .Q(n5697)
         );
  NOR2X0 U6584 ( .IN1(n4564), .IN2(n5698), .QN(WX6456) );
  XOR2X1 U6585 ( .IN1(n3652), .IN2(DFF_937_n1), .Q(n5698) );
  NOR2X0 U6586 ( .IN1(n4564), .IN2(n5699), .QN(WX6454) );
  XOR2X1 U6587 ( .IN1(n3654), .IN2(DFF_936_n1), .Q(n5699) );
  NOR2X0 U6588 ( .IN1(n4564), .IN2(n5700), .QN(WX6452) );
  XOR2X1 U6589 ( .IN1(n3656), .IN2(DFF_935_n1), .Q(n5700) );
  NOR2X0 U6590 ( .IN1(n4564), .IN2(n5701), .QN(WX6450) );
  XOR2X1 U6591 ( .IN1(n3658), .IN2(DFF_934_n1), .Q(n5701) );
  NOR2X0 U6592 ( .IN1(n4564), .IN2(n5702), .QN(WX6448) );
  XOR2X1 U6593 ( .IN1(n3660), .IN2(DFF_933_n1), .Q(n5702) );
  NOR2X0 U6594 ( .IN1(n4564), .IN2(n5703), .QN(WX6446) );
  XOR2X1 U6595 ( .IN1(n3662), .IN2(DFF_932_n1), .Q(n5703) );
  NOR2X0 U6596 ( .IN1(n4564), .IN2(n5704), .QN(WX6444) );
  XOR3X1 U6597 ( .IN1(n3424), .IN2(DFF_959_n1), .IN3(CRC_OUT_5_3), .Q(n5704)
         );
  NOR2X0 U6598 ( .IN1(n4564), .IN2(n5705), .QN(WX6442) );
  XOR2X1 U6599 ( .IN1(n3664), .IN2(DFF_930_n1), .Q(n5705) );
  NOR2X0 U6600 ( .IN1(n4564), .IN2(n5706), .QN(WX6440) );
  XOR2X1 U6601 ( .IN1(n3665), .IN2(DFF_929_n1), .Q(n5706) );
  NAND4X0 U6602 ( .IN1(n5707), .IN2(n5708), .IN3(n5709), .IN4(n5710), .QN(
        WX644) );
  NAND2X0 U6603 ( .IN1(n3966), .IN2(n5711), .QN(n5710) );
  NAND2X0 U6604 ( .IN1(n3880), .IN2(n5712), .QN(n5709) );
  NAND2X0 U6605 ( .IN1(n3955), .IN2(CRC_OUT_9_31), .QN(n5708) );
  NAND2X0 U6606 ( .IN1(n2245), .IN2(WX485), .QN(n5707) );
  NOR2X0 U6607 ( .IN1(n4564), .IN2(n5713), .QN(WX6438) );
  XNOR2X1 U6608 ( .IN1(n3666), .IN2(test_so53), .Q(n5713) );
  NOR2X0 U6609 ( .IN1(n4564), .IN2(n5714), .QN(WX6436) );
  XOR2X1 U6610 ( .IN1(n3437), .IN2(DFF_959_n1), .Q(n5714) );
  NAND4X0 U6611 ( .IN1(n5715), .IN2(n5716), .IN3(n5717), .IN4(n5718), .QN(
        WX5878) );
  NAND2X0 U6612 ( .IN1(n3966), .IN2(n5273), .QN(n5718) );
  XNOR3X1 U6613 ( .IN1(n3436), .IN2(n3332), .IN3(n5719), .Q(n5273) );
  XOR2X1 U6614 ( .IN1(WX7236), .IN2(n7138), .Q(n5719) );
  NAND2X0 U6615 ( .IN1(n3880), .IN2(n5720), .QN(n5717) );
  NAND2X0 U6616 ( .IN1(n298), .IN2(n3922), .QN(n5716) );
  INVX0 U6617 ( .INP(n5721), .ZN(n298) );
  NAND2X0 U6618 ( .IN1(n4462), .IN2(n8496), .QN(n5721) );
  NAND2X0 U6619 ( .IN1(test_so53), .IN2(n3957), .QN(n5715) );
  NAND4X0 U6620 ( .IN1(n5722), .IN2(n5723), .IN3(n5724), .IN4(n5725), .QN(
        WX5876) );
  NAND2X0 U6621 ( .IN1(n3966), .IN2(n5280), .QN(n5725) );
  XNOR3X1 U6622 ( .IN1(n3616), .IN2(n3333), .IN3(n5726), .Q(n5280) );
  XOR2X1 U6623 ( .IN1(WX7234), .IN2(n7139), .Q(n5726) );
  NAND2X0 U6624 ( .IN1(n5727), .IN2(n3897), .QN(n5724) );
  NAND2X0 U6625 ( .IN1(n297), .IN2(n3922), .QN(n5723) );
  INVX0 U6626 ( .INP(n5728), .ZN(n297) );
  NAND2X0 U6627 ( .IN1(n4462), .IN2(n8497), .QN(n5728) );
  NAND2X0 U6628 ( .IN1(n3954), .IN2(CRC_OUT_5_1), .QN(n5722) );
  NAND4X0 U6629 ( .IN1(n5729), .IN2(n5730), .IN3(n5731), .IN4(n5732), .QN(
        WX5874) );
  NAND2X0 U6630 ( .IN1(n3966), .IN2(n5287), .QN(n5732) );
  XNOR3X1 U6631 ( .IN1(n3614), .IN2(n3334), .IN3(n5733), .Q(n5287) );
  XOR2X1 U6632 ( .IN1(WX7232), .IN2(n7140), .Q(n5733) );
  NAND2X0 U6633 ( .IN1(n3880), .IN2(n5734), .QN(n5731) );
  NAND2X0 U6634 ( .IN1(n296), .IN2(n3922), .QN(n5730) );
  INVX0 U6635 ( .INP(n5735), .ZN(n296) );
  NAND2X0 U6636 ( .IN1(n4460), .IN2(n8498), .QN(n5735) );
  NAND2X0 U6637 ( .IN1(n3956), .IN2(CRC_OUT_5_2), .QN(n5729) );
  NAND4X0 U6638 ( .IN1(n5736), .IN2(n5737), .IN3(n5738), .IN4(n5739), .QN(
        WX5872) );
  NAND2X0 U6639 ( .IN1(n3966), .IN2(n5294), .QN(n5739) );
  XNOR3X1 U6640 ( .IN1(n3612), .IN2(n3335), .IN3(n5740), .Q(n5294) );
  XOR2X1 U6641 ( .IN1(WX7230), .IN2(n7141), .Q(n5740) );
  NAND2X0 U6642 ( .IN1(n5741), .IN2(n3898), .QN(n5738) );
  NAND2X0 U6643 ( .IN1(n295), .IN2(n3922), .QN(n5737) );
  INVX0 U6644 ( .INP(n5742), .ZN(n295) );
  NAND2X0 U6645 ( .IN1(n4462), .IN2(n8499), .QN(n5742) );
  NAND2X0 U6646 ( .IN1(n3955), .IN2(CRC_OUT_5_3), .QN(n5736) );
  NAND4X0 U6647 ( .IN1(n5743), .IN2(n5744), .IN3(n5745), .IN4(n5746), .QN(
        WX5870) );
  NAND2X0 U6648 ( .IN1(n5301), .IN2(n3985), .QN(n5746) );
  XOR3X1 U6649 ( .IN1(n3635), .IN2(n3336), .IN3(n5747), .Q(n5301) );
  XOR2X1 U6650 ( .IN1(WX7164), .IN2(test_so64), .Q(n5747) );
  NAND2X0 U6651 ( .IN1(n3879), .IN2(n5748), .QN(n5745) );
  NAND2X0 U6652 ( .IN1(n294), .IN2(n3922), .QN(n5744) );
  INVX0 U6653 ( .INP(n5749), .ZN(n294) );
  NAND2X0 U6654 ( .IN1(n4462), .IN2(n8500), .QN(n5749) );
  NAND2X0 U6655 ( .IN1(n3956), .IN2(CRC_OUT_5_4), .QN(n5743) );
  NAND4X0 U6656 ( .IN1(n5750), .IN2(n5751), .IN3(n5752), .IN4(n5753), .QN(
        WX5868) );
  NAND2X0 U6657 ( .IN1(n3966), .IN2(n5308), .QN(n5753) );
  XNOR3X1 U6658 ( .IN1(n3610), .IN2(n3337), .IN3(n5754), .Q(n5308) );
  XOR2X1 U6659 ( .IN1(WX7226), .IN2(n7142), .Q(n5754) );
  NAND2X0 U6660 ( .IN1(n5755), .IN2(n3898), .QN(n5752) );
  NAND2X0 U6661 ( .IN1(n293), .IN2(n3922), .QN(n5751) );
  INVX0 U6662 ( .INP(n5756), .ZN(n293) );
  NAND2X0 U6663 ( .IN1(n4461), .IN2(n8501), .QN(n5756) );
  NAND2X0 U6664 ( .IN1(n3955), .IN2(CRC_OUT_5_5), .QN(n5750) );
  NAND4X0 U6665 ( .IN1(n5757), .IN2(n5758), .IN3(n5759), .IN4(n5760), .QN(
        WX5866) );
  NAND2X0 U6666 ( .IN1(n5314), .IN2(n3985), .QN(n5760) );
  XOR3X1 U6667 ( .IN1(n3639), .IN2(n3608), .IN3(n5761), .Q(n5314) );
  XOR2X1 U6668 ( .IN1(WX7160), .IN2(test_so62), .Q(n5761) );
  NAND2X0 U6669 ( .IN1(n3879), .IN2(n5762), .QN(n5759) );
  NAND2X0 U6670 ( .IN1(n292), .IN2(n3922), .QN(n5758) );
  INVX0 U6671 ( .INP(n5763), .ZN(n292) );
  NAND2X0 U6672 ( .IN1(n4461), .IN2(n8502), .QN(n5763) );
  NAND2X0 U6673 ( .IN1(n3956), .IN2(CRC_OUT_5_6), .QN(n5757) );
  NAND4X0 U6674 ( .IN1(n5764), .IN2(n5765), .IN3(n5766), .IN4(n5767), .QN(
        WX5864) );
  NAND2X0 U6675 ( .IN1(n3966), .IN2(n5321), .QN(n5767) );
  XNOR3X1 U6676 ( .IN1(n3606), .IN2(n3338), .IN3(n5768), .Q(n5321) );
  XOR2X1 U6677 ( .IN1(WX7222), .IN2(n7143), .Q(n5768) );
  NAND2X0 U6678 ( .IN1(n3879), .IN2(n5769), .QN(n5766) );
  NAND2X0 U6679 ( .IN1(n291), .IN2(n3922), .QN(n5765) );
  INVX0 U6680 ( .INP(n5770), .ZN(n291) );
  NAND2X0 U6681 ( .IN1(test_so45), .IN2(n4464), .QN(n5770) );
  NAND2X0 U6682 ( .IN1(n3956), .IN2(CRC_OUT_5_7), .QN(n5764) );
  NAND4X0 U6683 ( .IN1(n5771), .IN2(n5772), .IN3(n5773), .IN4(n5774), .QN(
        WX5862) );
  NAND2X0 U6684 ( .IN1(n5328), .IN2(n3985), .QN(n5774) );
  XOR3X1 U6685 ( .IN1(n3604), .IN2(n3339), .IN3(n5775), .Q(n5328) );
  XOR2X1 U6686 ( .IN1(WX7156), .IN2(test_so60), .Q(n5775) );
  NAND2X0 U6687 ( .IN1(n3879), .IN2(n5776), .QN(n5773) );
  NAND2X0 U6688 ( .IN1(n290), .IN2(n3922), .QN(n5772) );
  INVX0 U6689 ( .INP(n5777), .ZN(n290) );
  NAND2X0 U6690 ( .IN1(n4461), .IN2(n8505), .QN(n5777) );
  NAND2X0 U6691 ( .IN1(n3955), .IN2(CRC_OUT_5_8), .QN(n5771) );
  NAND4X0 U6692 ( .IN1(n5778), .IN2(n5779), .IN3(n5780), .IN4(n5781), .QN(
        WX5860) );
  NAND2X0 U6693 ( .IN1(n3966), .IN2(n5335), .QN(n5781) );
  XNOR3X1 U6694 ( .IN1(n3602), .IN2(n3340), .IN3(n5782), .Q(n5335) );
  XOR2X1 U6695 ( .IN1(WX7218), .IN2(n7144), .Q(n5782) );
  NAND2X0 U6696 ( .IN1(n3879), .IN2(n5783), .QN(n5780) );
  NAND2X0 U6697 ( .IN1(n289), .IN2(n3922), .QN(n5779) );
  INVX0 U6698 ( .INP(n5784), .ZN(n289) );
  NAND2X0 U6699 ( .IN1(n4461), .IN2(n8506), .QN(n5784) );
  NAND2X0 U6700 ( .IN1(n3956), .IN2(CRC_OUT_5_9), .QN(n5778) );
  NAND4X0 U6701 ( .IN1(n5785), .IN2(n5786), .IN3(n5787), .IN4(n5788), .QN(
        WX5858) );
  NAND2X0 U6702 ( .IN1(n5342), .IN2(n3986), .QN(n5788) );
  XOR3X1 U6703 ( .IN1(n3647), .IN2(n3600), .IN3(n5789), .Q(n5342) );
  XOR2X1 U6704 ( .IN1(WX7280), .IN2(test_so58), .Q(n5789) );
  NAND2X0 U6705 ( .IN1(n3879), .IN2(n5790), .QN(n5787) );
  NAND2X0 U6706 ( .IN1(n288), .IN2(n3922), .QN(n5786) );
  INVX0 U6707 ( .INP(n5791), .ZN(n288) );
  NAND2X0 U6708 ( .IN1(n4460), .IN2(n8507), .QN(n5791) );
  NAND2X0 U6709 ( .IN1(n3955), .IN2(CRC_OUT_5_10), .QN(n5785) );
  NAND4X0 U6710 ( .IN1(n5792), .IN2(n5793), .IN3(n5794), .IN4(n5795), .QN(
        WX5856) );
  NAND2X0 U6711 ( .IN1(n3966), .IN2(n5349), .QN(n5795) );
  XNOR3X1 U6712 ( .IN1(n3422), .IN2(n3341), .IN3(n5796), .Q(n5349) );
  XOR2X1 U6713 ( .IN1(WX7214), .IN2(n7145), .Q(n5796) );
  NAND2X0 U6714 ( .IN1(n3879), .IN2(n5797), .QN(n5794) );
  NAND2X0 U6715 ( .IN1(n287), .IN2(n3923), .QN(n5793) );
  INVX0 U6716 ( .INP(n5798), .ZN(n287) );
  NAND2X0 U6717 ( .IN1(n4461), .IN2(n8508), .QN(n5798) );
  NAND2X0 U6718 ( .IN1(n3954), .IN2(CRC_OUT_5_11), .QN(n5792) );
  NAND4X0 U6719 ( .IN1(n5799), .IN2(n5800), .IN3(n5801), .IN4(n5802), .QN(
        WX5854) );
  NAND2X0 U6720 ( .IN1(n3966), .IN2(n5356), .QN(n5802) );
  XNOR3X1 U6721 ( .IN1(n3598), .IN2(n3342), .IN3(n5803), .Q(n5356) );
  XOR2X1 U6722 ( .IN1(WX7212), .IN2(n7146), .Q(n5803) );
  NAND2X0 U6723 ( .IN1(n3879), .IN2(n5804), .QN(n5801) );
  NAND2X0 U6724 ( .IN1(n286), .IN2(n3923), .QN(n5800) );
  INVX0 U6725 ( .INP(n5805), .ZN(n286) );
  NAND2X0 U6726 ( .IN1(n4461), .IN2(n8509), .QN(n5805) );
  NAND2X0 U6727 ( .IN1(n3939), .IN2(CRC_OUT_5_12), .QN(n5799) );
  NAND4X0 U6728 ( .IN1(n5806), .IN2(n5807), .IN3(n5808), .IN4(n5809), .QN(
        WX5852) );
  NAND2X0 U6729 ( .IN1(n3966), .IN2(n5363), .QN(n5809) );
  XNOR3X1 U6730 ( .IN1(n3596), .IN2(n3343), .IN3(n5810), .Q(n5363) );
  XOR2X1 U6731 ( .IN1(WX7210), .IN2(n7147), .Q(n5810) );
  NAND2X0 U6732 ( .IN1(n3879), .IN2(n5811), .QN(n5808) );
  NAND2X0 U6733 ( .IN1(n285), .IN2(n3923), .QN(n5807) );
  INVX0 U6734 ( .INP(n5812), .ZN(n285) );
  NAND2X0 U6735 ( .IN1(n4459), .IN2(n8510), .QN(n5812) );
  NAND2X0 U6736 ( .IN1(n3934), .IN2(CRC_OUT_5_13), .QN(n5806) );
  NAND4X0 U6737 ( .IN1(n5813), .IN2(n5814), .IN3(n5815), .IN4(n5816), .QN(
        WX5850) );
  NAND2X0 U6738 ( .IN1(n3966), .IN2(n5370), .QN(n5816) );
  XNOR3X1 U6739 ( .IN1(n3594), .IN2(n3344), .IN3(n5817), .Q(n5370) );
  XOR2X1 U6740 ( .IN1(WX7208), .IN2(n7148), .Q(n5817) );
  NAND2X0 U6741 ( .IN1(n3879), .IN2(n5818), .QN(n5815) );
  NAND2X0 U6742 ( .IN1(n284), .IN2(n3923), .QN(n5814) );
  INVX0 U6743 ( .INP(n5819), .ZN(n284) );
  NAND2X0 U6744 ( .IN1(n4460), .IN2(n8511), .QN(n5819) );
  NAND2X0 U6745 ( .IN1(n3934), .IN2(CRC_OUT_5_14), .QN(n5813) );
  NAND4X0 U6746 ( .IN1(n5820), .IN2(n5821), .IN3(n5822), .IN4(n5823), .QN(
        WX5848) );
  NAND2X0 U6747 ( .IN1(n3967), .IN2(n5377), .QN(n5823) );
  XNOR3X1 U6748 ( .IN1(n3592), .IN2(n3345), .IN3(n5824), .Q(n5377) );
  XOR2X1 U6749 ( .IN1(WX7206), .IN2(n7149), .Q(n5824) );
  NAND2X0 U6750 ( .IN1(n3879), .IN2(n5825), .QN(n5822) );
  NAND2X0 U6751 ( .IN1(n283), .IN2(n3923), .QN(n5821) );
  INVX0 U6752 ( .INP(n5826), .ZN(n283) );
  NAND2X0 U6753 ( .IN1(n4460), .IN2(n8512), .QN(n5826) );
  NAND2X0 U6754 ( .IN1(n3934), .IN2(CRC_OUT_5_15), .QN(n5820) );
  NAND4X0 U6755 ( .IN1(n5827), .IN2(n5828), .IN3(n5829), .IN4(n5830), .QN(
        WX5846) );
  NAND2X0 U6756 ( .IN1(n3967), .IN2(n5384), .QN(n5830) );
  XOR3X1 U6757 ( .IN1(n3156), .IN2(n3873), .IN3(n5831), .Q(n5384) );
  XOR3X1 U6758 ( .IN1(n7150), .IN2(n3421), .IN3(WX7268), .Q(n5831) );
  NAND2X0 U6759 ( .IN1(n5832), .IN2(n3899), .QN(n5829) );
  NAND2X0 U6760 ( .IN1(n282), .IN2(n3923), .QN(n5828) );
  INVX0 U6761 ( .INP(n5833), .ZN(n282) );
  NAND2X0 U6762 ( .IN1(n4459), .IN2(n8513), .QN(n5833) );
  NAND2X0 U6763 ( .IN1(n3934), .IN2(CRC_OUT_5_16), .QN(n5827) );
  NAND4X0 U6764 ( .IN1(n5834), .IN2(n5835), .IN3(n5836), .IN4(n5837), .QN(
        WX5844) );
  NAND2X0 U6765 ( .IN1(n3967), .IN2(n5391), .QN(n5837) );
  XOR3X1 U6766 ( .IN1(n3158), .IN2(n3872), .IN3(n5838), .Q(n5391) );
  XOR3X1 U6767 ( .IN1(n7151), .IN2(n3590), .IN3(WX7266), .Q(n5838) );
  NAND2X0 U6768 ( .IN1(n3879), .IN2(n5839), .QN(n5836) );
  NAND2X0 U6769 ( .IN1(n281), .IN2(n3923), .QN(n5835) );
  INVX0 U6770 ( .INP(n5840), .ZN(n281) );
  NAND2X0 U6771 ( .IN1(n4460), .IN2(n8514), .QN(n5840) );
  NAND2X0 U6772 ( .IN1(test_so54), .IN2(n3957), .QN(n5834) );
  NAND4X0 U6773 ( .IN1(n5841), .IN2(n5842), .IN3(n5843), .IN4(n5844), .QN(
        WX5842) );
  NAND2X0 U6774 ( .IN1(n3967), .IN2(n5398), .QN(n5844) );
  XOR3X1 U6775 ( .IN1(n3160), .IN2(n3875), .IN3(n5845), .Q(n5398) );
  XOR3X1 U6776 ( .IN1(n7152), .IN2(n3588), .IN3(WX7264), .Q(n5845) );
  NAND2X0 U6777 ( .IN1(n5846), .IN2(n3899), .QN(n5843) );
  NAND2X0 U6778 ( .IN1(n280), .IN2(n3923), .QN(n5842) );
  INVX0 U6779 ( .INP(n5847), .ZN(n280) );
  NAND2X0 U6780 ( .IN1(n4460), .IN2(n8515), .QN(n5847) );
  NAND2X0 U6781 ( .IN1(n3934), .IN2(CRC_OUT_5_18), .QN(n5841) );
  NAND4X0 U6782 ( .IN1(n5848), .IN2(n5849), .IN3(n5850), .IN4(n5851), .QN(
        WX5840) );
  NAND2X0 U6783 ( .IN1(n3967), .IN2(n5405), .QN(n5851) );
  XOR3X1 U6784 ( .IN1(n3162), .IN2(n3874), .IN3(n5852), .Q(n5405) );
  XOR3X1 U6785 ( .IN1(n7153), .IN2(n3586), .IN3(WX7262), .Q(n5852) );
  NAND2X0 U6786 ( .IN1(n3878), .IN2(n5853), .QN(n5850) );
  NAND2X0 U6787 ( .IN1(n279), .IN2(n3923), .QN(n5849) );
  INVX0 U6788 ( .INP(n5854), .ZN(n279) );
  NAND2X0 U6789 ( .IN1(n4460), .IN2(n8516), .QN(n5854) );
  NAND2X0 U6790 ( .IN1(n3934), .IN2(CRC_OUT_5_19), .QN(n5848) );
  NAND4X0 U6791 ( .IN1(n5855), .IN2(n5856), .IN3(n5857), .IN4(n5858), .QN(
        WX5838) );
  NAND2X0 U6792 ( .IN1(n3967), .IN2(n5412), .QN(n5858) );
  XOR3X1 U6793 ( .IN1(n3164), .IN2(n3873), .IN3(n5859), .Q(n5412) );
  XOR3X1 U6794 ( .IN1(n7154), .IN2(n3584), .IN3(WX7260), .Q(n5859) );
  NAND2X0 U6795 ( .IN1(n5860), .IN2(n3899), .QN(n5857) );
  NAND2X0 U6796 ( .IN1(n278), .IN2(n3923), .QN(n5856) );
  INVX0 U6797 ( .INP(n5861), .ZN(n278) );
  NAND2X0 U6798 ( .IN1(n4458), .IN2(n8517), .QN(n5861) );
  NAND2X0 U6799 ( .IN1(n3934), .IN2(CRC_OUT_5_20), .QN(n5855) );
  NAND4X0 U6800 ( .IN1(n5862), .IN2(n5863), .IN3(n5864), .IN4(n5865), .QN(
        WX5836) );
  NAND2X0 U6801 ( .IN1(n5419), .IN2(n3986), .QN(n5865) );
  XOR3X1 U6802 ( .IN1(n3166), .IN2(TM1), .IN3(n5866), .Q(n5419) );
  XOR3X1 U6803 ( .IN1(test_so63), .IN2(n7155), .IN3(WX7258), .Q(n5866) );
  NAND2X0 U6804 ( .IN1(n3878), .IN2(n5867), .QN(n5864) );
  NAND2X0 U6805 ( .IN1(n277), .IN2(n3923), .QN(n5863) );
  INVX0 U6806 ( .INP(n5868), .ZN(n277) );
  NAND2X0 U6807 ( .IN1(n4460), .IN2(n8518), .QN(n5868) );
  NAND2X0 U6808 ( .IN1(n3934), .IN2(CRC_OUT_5_21), .QN(n5862) );
  NAND4X0 U6809 ( .IN1(n5869), .IN2(n5870), .IN3(n5871), .IN4(n5872), .QN(
        WX5834) );
  NAND2X0 U6810 ( .IN1(n3967), .IN2(n5426), .QN(n5872) );
  XOR3X1 U6811 ( .IN1(n3167), .IN2(n3872), .IN3(n5873), .Q(n5426) );
  XOR3X1 U6812 ( .IN1(n7156), .IN2(n3582), .IN3(WX7256), .Q(n5873) );
  NAND2X0 U6813 ( .IN1(n5874), .IN2(n3899), .QN(n5871) );
  NAND2X0 U6814 ( .IN1(n276), .IN2(n3923), .QN(n5870) );
  INVX0 U6815 ( .INP(n5875), .ZN(n276) );
  NAND2X0 U6816 ( .IN1(n4459), .IN2(n8519), .QN(n5875) );
  NAND2X0 U6817 ( .IN1(n3934), .IN2(CRC_OUT_5_22), .QN(n5869) );
  NAND4X0 U6818 ( .IN1(n5876), .IN2(n5877), .IN3(n5878), .IN4(n5879), .QN(
        WX5832) );
  NAND2X0 U6819 ( .IN1(n5433), .IN2(n3986), .QN(n5879) );
  XOR3X1 U6820 ( .IN1(n3169), .IN2(TM1), .IN3(n5880), .Q(n5433) );
  XNOR3X1 U6821 ( .IN1(test_so61), .IN2(n7157), .IN3(n3580), .Q(n5880) );
  NAND2X0 U6822 ( .IN1(n3878), .IN2(n5881), .QN(n5878) );
  NAND2X0 U6823 ( .IN1(n275), .IN2(n3923), .QN(n5877) );
  INVX0 U6824 ( .INP(n5882), .ZN(n275) );
  NAND2X0 U6825 ( .IN1(n4459), .IN2(n8520), .QN(n5882) );
  NAND2X0 U6826 ( .IN1(n3934), .IN2(CRC_OUT_5_23), .QN(n5876) );
  NAND4X0 U6827 ( .IN1(n5883), .IN2(n5884), .IN3(n5885), .IN4(n5886), .QN(
        WX5830) );
  NAND2X0 U6828 ( .IN1(n3967), .IN2(n5440), .QN(n5886) );
  XOR3X1 U6829 ( .IN1(n3170), .IN2(n3875), .IN3(n5887), .Q(n5440) );
  XOR3X1 U6830 ( .IN1(n7158), .IN2(n3578), .IN3(WX7252), .Q(n5887) );
  NAND2X0 U6831 ( .IN1(n3878), .IN2(n5888), .QN(n5885) );
  NAND2X0 U6832 ( .IN1(n274), .IN2(n3923), .QN(n5884) );
  INVX0 U6833 ( .INP(n5889), .ZN(n274) );
  NAND2X0 U6834 ( .IN1(test_so44), .IN2(n4464), .QN(n5889) );
  NAND2X0 U6835 ( .IN1(n3934), .IN2(CRC_OUT_5_24), .QN(n5883) );
  NAND4X0 U6836 ( .IN1(n5890), .IN2(n5891), .IN3(n5892), .IN4(n5893), .QN(
        WX5828) );
  NAND2X0 U6837 ( .IN1(n5447), .IN2(n3987), .QN(n5893) );
  XOR3X1 U6838 ( .IN1(n3172), .IN2(TM1), .IN3(n5894), .Q(n5447) );
  XNOR3X1 U6839 ( .IN1(test_so59), .IN2(n7159), .IN3(n3576), .Q(n5894) );
  NAND2X0 U6840 ( .IN1(n3878), .IN2(n5895), .QN(n5892) );
  NAND2X0 U6841 ( .IN1(n273), .IN2(n3923), .QN(n5891) );
  INVX0 U6842 ( .INP(n5896), .ZN(n273) );
  NAND2X0 U6843 ( .IN1(n4459), .IN2(n8523), .QN(n5896) );
  NAND2X0 U6844 ( .IN1(n3935), .IN2(CRC_OUT_5_25), .QN(n5890) );
  NAND4X0 U6845 ( .IN1(n5897), .IN2(n5898), .IN3(n5899), .IN4(n5900), .QN(
        WX5826) );
  NAND2X0 U6846 ( .IN1(n3967), .IN2(n5454), .QN(n5900) );
  XOR3X1 U6847 ( .IN1(n3173), .IN2(n3874), .IN3(n5901), .Q(n5454) );
  XOR3X1 U6848 ( .IN1(n7160), .IN2(n3574), .IN3(WX7248), .Q(n5901) );
  NAND2X0 U6849 ( .IN1(n3878), .IN2(n5902), .QN(n5899) );
  NAND2X0 U6850 ( .IN1(n272), .IN2(n3923), .QN(n5898) );
  INVX0 U6851 ( .INP(n5903), .ZN(n272) );
  NAND2X0 U6852 ( .IN1(n4458), .IN2(n8524), .QN(n5903) );
  NAND2X0 U6853 ( .IN1(n3935), .IN2(CRC_OUT_5_26), .QN(n5897) );
  NAND4X0 U6854 ( .IN1(n5904), .IN2(n5905), .IN3(n5906), .IN4(n5907), .QN(
        WX5824) );
  NAND2X0 U6855 ( .IN1(n5461), .IN2(n3987), .QN(n5907) );
  XOR3X1 U6856 ( .IN1(n3175), .IN2(TM1), .IN3(n5908), .Q(n5461) );
  XNOR3X1 U6857 ( .IN1(test_so57), .IN2(n7161), .IN3(n3572), .Q(n5908) );
  NAND2X0 U6858 ( .IN1(n3878), .IN2(n5909), .QN(n5906) );
  NAND2X0 U6859 ( .IN1(n271), .IN2(n3923), .QN(n5905) );
  INVX0 U6860 ( .INP(n5910), .ZN(n271) );
  NAND2X0 U6861 ( .IN1(n4459), .IN2(n8525), .QN(n5910) );
  NAND2X0 U6862 ( .IN1(n3935), .IN2(CRC_OUT_5_27), .QN(n5904) );
  NAND4X0 U6863 ( .IN1(n5911), .IN2(n5912), .IN3(n5913), .IN4(n5914), .QN(
        WX5822) );
  NAND2X0 U6864 ( .IN1(n3967), .IN2(n5468), .QN(n5914) );
  XOR3X1 U6865 ( .IN1(n3176), .IN2(n3873), .IN3(n5915), .Q(n5468) );
  XOR3X1 U6866 ( .IN1(n7162), .IN2(n3570), .IN3(WX7244), .Q(n5915) );
  NAND2X0 U6867 ( .IN1(n3878), .IN2(n5916), .QN(n5913) );
  NAND2X0 U6868 ( .IN1(n270), .IN2(n3924), .QN(n5912) );
  INVX0 U6869 ( .INP(n5917), .ZN(n270) );
  NAND2X0 U6870 ( .IN1(n4459), .IN2(n8526), .QN(n5917) );
  NAND2X0 U6871 ( .IN1(n3935), .IN2(CRC_OUT_5_28), .QN(n5911) );
  NAND4X0 U6872 ( .IN1(n5918), .IN2(n5919), .IN3(n5920), .IN4(n5921), .QN(
        WX5820) );
  NAND2X0 U6873 ( .IN1(n3967), .IN2(n5475), .QN(n5921) );
  XOR3X1 U6874 ( .IN1(n3178), .IN2(n3872), .IN3(n5922), .Q(n5475) );
  XOR3X1 U6875 ( .IN1(n7163), .IN2(n3568), .IN3(WX7242), .Q(n5922) );
  NAND2X0 U6876 ( .IN1(n3878), .IN2(n5923), .QN(n5920) );
  NAND2X0 U6877 ( .IN1(n269), .IN2(n3924), .QN(n5919) );
  INVX0 U6878 ( .INP(n5924), .ZN(n269) );
  NAND2X0 U6879 ( .IN1(n4458), .IN2(n8527), .QN(n5924) );
  NAND2X0 U6880 ( .IN1(n3935), .IN2(CRC_OUT_5_29), .QN(n5918) );
  NAND4X0 U6881 ( .IN1(n5925), .IN2(n5926), .IN3(n5927), .IN4(n5928), .QN(
        WX5818) );
  NAND2X0 U6882 ( .IN1(n3967), .IN2(n5482), .QN(n5928) );
  XOR3X1 U6883 ( .IN1(n3180), .IN2(n3875), .IN3(n5929), .Q(n5482) );
  XOR3X1 U6884 ( .IN1(n7164), .IN2(n3566), .IN3(WX7240), .Q(n5929) );
  NAND2X0 U6885 ( .IN1(n3878), .IN2(n5930), .QN(n5927) );
  NAND2X0 U6886 ( .IN1(n268), .IN2(n3924), .QN(n5926) );
  INVX0 U6887 ( .INP(n5931), .ZN(n268) );
  NAND2X0 U6888 ( .IN1(n4459), .IN2(n8528), .QN(n5931) );
  NAND2X0 U6889 ( .IN1(n3935), .IN2(CRC_OUT_5_30), .QN(n5925) );
  NAND4X0 U6890 ( .IN1(n5932), .IN2(n5933), .IN3(n5934), .IN4(n5935), .QN(
        WX5816) );
  NAND2X0 U6891 ( .IN1(n3968), .IN2(n5489), .QN(n5935) );
  XOR3X1 U6892 ( .IN1(n3066), .IN2(n3874), .IN3(n5936), .Q(n5489) );
  XOR3X1 U6893 ( .IN1(n7165), .IN2(n3565), .IN3(WX7238), .Q(n5936) );
  NAND2X0 U6894 ( .IN1(n3878), .IN2(n5937), .QN(n5934) );
  NAND2X0 U6895 ( .IN1(n3935), .IN2(CRC_OUT_5_31), .QN(n5933) );
  NAND2X0 U6896 ( .IN1(n2245), .IN2(WX5657), .QN(n5932) );
  NOR2X0 U6897 ( .IN1(n4564), .IN2(WX5657), .QN(WX5718) );
  NOR2X0 U6898 ( .IN1(n4564), .IN2(WX485), .QN(WX546) );
  NOR2X0 U6899 ( .IN1(n4564), .IN2(n5938), .QN(WX5205) );
  XOR2X1 U6900 ( .IN1(n3668), .IN2(DFF_766_n1), .Q(n5938) );
  NOR2X0 U6901 ( .IN1(n4565), .IN2(n5939), .QN(WX5203) );
  XOR2X1 U6902 ( .IN1(n3670), .IN2(DFF_765_n1), .Q(n5939) );
  NOR2X0 U6903 ( .IN1(n4565), .IN2(n5940), .QN(WX5201) );
  XOR2X1 U6904 ( .IN1(n3672), .IN2(DFF_764_n1), .Q(n5940) );
  NOR2X0 U6905 ( .IN1(n4565), .IN2(n5941), .QN(WX5199) );
  XOR2X1 U6906 ( .IN1(CRC_OUT_6_27), .IN2(test_so40), .Q(n5941) );
  NOR2X0 U6907 ( .IN1(n4565), .IN2(n5942), .QN(WX5197) );
  XOR2X1 U6908 ( .IN1(n3674), .IN2(DFF_762_n1), .Q(n5942) );
  NOR2X0 U6909 ( .IN1(n4565), .IN2(n5943), .QN(WX5195) );
  XOR2X1 U6910 ( .IN1(n3676), .IN2(DFF_761_n1), .Q(n5943) );
  NOR2X0 U6911 ( .IN1(n4565), .IN2(n5944), .QN(WX5193) );
  XOR2X1 U6912 ( .IN1(n3678), .IN2(DFF_760_n1), .Q(n5944) );
  NOR2X0 U6913 ( .IN1(n4565), .IN2(n5945), .QN(WX5191) );
  XOR2X1 U6914 ( .IN1(n3680), .IN2(DFF_759_n1), .Q(n5945) );
  NOR2X0 U6915 ( .IN1(n4565), .IN2(n5946), .QN(WX5189) );
  XNOR2X1 U6916 ( .IN1(n3682), .IN2(test_so43), .Q(n5946) );
  NOR2X0 U6917 ( .IN1(n4565), .IN2(n5947), .QN(WX5187) );
  XOR2X1 U6918 ( .IN1(n3684), .IN2(DFF_757_n1), .Q(n5947) );
  NOR2X0 U6919 ( .IN1(n4565), .IN2(n5948), .QN(WX5185) );
  XOR2X1 U6920 ( .IN1(n3686), .IN2(DFF_756_n1), .Q(n5948) );
  NOR2X0 U6921 ( .IN1(n4565), .IN2(n5949), .QN(WX5183) );
  XOR2X1 U6922 ( .IN1(n3688), .IN2(DFF_755_n1), .Q(n5949) );
  NOR2X0 U6923 ( .IN1(n4565), .IN2(n5950), .QN(WX5181) );
  XOR2X1 U6924 ( .IN1(n3690), .IN2(DFF_754_n1), .Q(n5950) );
  NOR2X0 U6925 ( .IN1(n4565), .IN2(n5951), .QN(WX5179) );
  XOR2X1 U6926 ( .IN1(n3692), .IN2(DFF_753_n1), .Q(n5951) );
  NOR2X0 U6927 ( .IN1(n4565), .IN2(n5952), .QN(WX5177) );
  XOR2X1 U6928 ( .IN1(n3694), .IN2(DFF_752_n1), .Q(n5952) );
  NOR2X0 U6929 ( .IN1(n4565), .IN2(n5953), .QN(WX5175) );
  XOR3X1 U6930 ( .IN1(n3425), .IN2(DFF_767_n1), .IN3(CRC_OUT_6_15), .Q(n5953)
         );
  NOR2X0 U6931 ( .IN1(n4565), .IN2(n5954), .QN(WX5173) );
  XOR2X1 U6932 ( .IN1(n3696), .IN2(DFF_750_n1), .Q(n5954) );
  NOR2X0 U6933 ( .IN1(n4566), .IN2(n5955), .QN(WX5171) );
  XOR2X1 U6934 ( .IN1(n3698), .IN2(DFF_749_n1), .Q(n5955) );
  NOR2X0 U6935 ( .IN1(n4566), .IN2(n5956), .QN(WX5169) );
  XOR2X1 U6936 ( .IN1(n3700), .IN2(DFF_748_n1), .Q(n5956) );
  NOR2X0 U6937 ( .IN1(n4566), .IN2(n5957), .QN(WX5167) );
  XOR2X1 U6938 ( .IN1(n3702), .IN2(DFF_747_n1), .Q(n5957) );
  NOR2X0 U6939 ( .IN1(n4566), .IN2(n5958), .QN(WX5165) );
  XOR3X1 U6940 ( .IN1(test_so41), .IN2(DFF_767_n1), .IN3(DFF_746_n1), .Q(n5958) );
  NOR2X0 U6941 ( .IN1(n4566), .IN2(n5959), .QN(WX5163) );
  XOR2X1 U6942 ( .IN1(n3704), .IN2(DFF_745_n1), .Q(n5959) );
  NOR2X0 U6943 ( .IN1(n4566), .IN2(n5960), .QN(WX5161) );
  XOR2X1 U6944 ( .IN1(n3706), .IN2(DFF_744_n1), .Q(n5960) );
  NOR2X0 U6945 ( .IN1(n4566), .IN2(n5961), .QN(WX5159) );
  XOR2X1 U6946 ( .IN1(n3708), .IN2(DFF_743_n1), .Q(n5961) );
  NOR2X0 U6947 ( .IN1(n4566), .IN2(n5962), .QN(WX5157) );
  XOR2X1 U6948 ( .IN1(n3710), .IN2(DFF_742_n1), .Q(n5962) );
  NOR2X0 U6949 ( .IN1(n4566), .IN2(n5963), .QN(WX5155) );
  XNOR2X1 U6950 ( .IN1(n3712), .IN2(test_so42), .Q(n5963) );
  NOR2X0 U6951 ( .IN1(n4566), .IN2(n5964), .QN(WX5153) );
  XOR2X1 U6952 ( .IN1(n3714), .IN2(DFF_740_n1), .Q(n5964) );
  NOR2X0 U6953 ( .IN1(n4566), .IN2(n5965), .QN(WX5151) );
  XOR3X1 U6954 ( .IN1(n3426), .IN2(DFF_767_n1), .IN3(CRC_OUT_6_3), .Q(n5965)
         );
  NOR2X0 U6955 ( .IN1(n4566), .IN2(n5966), .QN(WX5149) );
  XOR2X1 U6956 ( .IN1(n3716), .IN2(DFF_738_n1), .Q(n5966) );
  NOR2X0 U6957 ( .IN1(n4566), .IN2(n5967), .QN(WX5147) );
  XOR2X1 U6958 ( .IN1(n3718), .IN2(DFF_737_n1), .Q(n5967) );
  NOR2X0 U6959 ( .IN1(n4566), .IN2(n5968), .QN(WX5145) );
  XOR2X1 U6960 ( .IN1(n3720), .IN2(DFF_736_n1), .Q(n5968) );
  NOR2X0 U6961 ( .IN1(n4566), .IN2(n5969), .QN(WX5143) );
  XOR2X1 U6962 ( .IN1(n3438), .IN2(DFF_767_n1), .Q(n5969) );
  NAND4X0 U6963 ( .IN1(n5970), .IN2(n5971), .IN3(n5972), .IN4(n5973), .QN(
        WX4585) );
  NAND2X0 U6964 ( .IN1(n3968), .IN2(n5720), .QN(n5973) );
  XNOR3X1 U6965 ( .IN1(n3437), .IN2(n3346), .IN3(n5974), .Q(n5720) );
  XOR2X1 U6966 ( .IN1(WX5943), .IN2(n7166), .Q(n5974) );
  NAND2X0 U6967 ( .IN1(n5975), .IN2(n3901), .QN(n5972) );
  NAND2X0 U6968 ( .IN1(n220), .IN2(n3924), .QN(n5971) );
  INVX0 U6969 ( .INP(n5976), .ZN(n220) );
  NAND2X0 U6970 ( .IN1(n4458), .IN2(n8554), .QN(n5976) );
  NAND2X0 U6971 ( .IN1(n3935), .IN2(CRC_OUT_6_0), .QN(n5970) );
  NAND4X0 U6972 ( .IN1(n5977), .IN2(n5978), .IN3(n5979), .IN4(n5980), .QN(
        WX4583) );
  NAND2X0 U6973 ( .IN1(n5727), .IN2(n3987), .QN(n5980) );
  XOR3X1 U6974 ( .IN1(n3666), .IN2(n3661), .IN3(n5981), .Q(n5727) );
  XOR2X1 U6975 ( .IN1(WX5877), .IN2(test_so51), .Q(n5981) );
  NAND2X0 U6976 ( .IN1(n3883), .IN2(n5982), .QN(n5979) );
  NAND2X0 U6977 ( .IN1(n219), .IN2(n3924), .QN(n5978) );
  INVX0 U6978 ( .INP(n5983), .ZN(n219) );
  NAND2X0 U6979 ( .IN1(n4458), .IN2(n8555), .QN(n5983) );
  NAND2X0 U6980 ( .IN1(n3935), .IN2(CRC_OUT_6_1), .QN(n5977) );
  NAND4X0 U6981 ( .IN1(n5984), .IN2(n5985), .IN3(n5986), .IN4(n5987), .QN(
        WX4581) );
  NAND2X0 U6982 ( .IN1(n3968), .IN2(n5734), .QN(n5987) );
  XNOR3X1 U6983 ( .IN1(n3663), .IN2(n3347), .IN3(n5988), .Q(n5734) );
  XOR2X1 U6984 ( .IN1(WX6003), .IN2(n3665), .Q(n5988) );
  NAND2X0 U6985 ( .IN1(n3893), .IN2(n5989), .QN(n5986) );
  NAND2X0 U6986 ( .IN1(n218), .IN2(n3924), .QN(n5985) );
  INVX0 U6987 ( .INP(n5990), .ZN(n218) );
  NAND2X0 U6988 ( .IN1(test_so34), .IN2(n4463), .QN(n5990) );
  NAND2X0 U6989 ( .IN1(n3935), .IN2(CRC_OUT_6_2), .QN(n5984) );
  NAND4X0 U6990 ( .IN1(n5991), .IN2(n5992), .IN3(n5993), .IN4(n5994), .QN(
        WX4579) );
  NAND2X0 U6991 ( .IN1(n5741), .IN2(n3987), .QN(n5994) );
  XOR3X1 U6992 ( .IN1(n3664), .IN2(n3348), .IN3(n5995), .Q(n5741) );
  XOR2X1 U6993 ( .IN1(WX5873), .IN2(test_so49), .Q(n5995) );
  NAND2X0 U6994 ( .IN1(n3893), .IN2(n5996), .QN(n5993) );
  NAND2X0 U6995 ( .IN1(n217), .IN2(n3924), .QN(n5992) );
  INVX0 U6996 ( .INP(n5997), .ZN(n217) );
  NAND2X0 U6997 ( .IN1(n4458), .IN2(n8558), .QN(n5997) );
  NAND2X0 U6998 ( .IN1(n3935), .IN2(CRC_OUT_6_3), .QN(n5991) );
  NAND4X0 U6999 ( .IN1(n5998), .IN2(n5999), .IN3(n6000), .IN4(n6001), .QN(
        WX4577) );
  NAND2X0 U7000 ( .IN1(n3968), .IN2(n5748), .QN(n6001) );
  XNOR3X1 U7001 ( .IN1(n3424), .IN2(n3349), .IN3(n6002), .Q(n5748) );
  XOR2X1 U7002 ( .IN1(WX5935), .IN2(n7167), .Q(n6002) );
  NAND2X0 U7003 ( .IN1(n3893), .IN2(n6003), .QN(n6000) );
  NAND2X0 U7004 ( .IN1(n216), .IN2(n3924), .QN(n5999) );
  INVX0 U7005 ( .INP(n6004), .ZN(n216) );
  NAND2X0 U7006 ( .IN1(n4458), .IN2(n8559), .QN(n6004) );
  NAND2X0 U7007 ( .IN1(n3935), .IN2(CRC_OUT_6_4), .QN(n5998) );
  NAND4X0 U7008 ( .IN1(n6005), .IN2(n6006), .IN3(n6007), .IN4(n6008), .QN(
        WX4575) );
  NAND2X0 U7009 ( .IN1(n5755), .IN2(n3981), .QN(n6008) );
  XOR3X1 U7010 ( .IN1(n3669), .IN2(n3662), .IN3(n6009), .Q(n5755) );
  XOR2X1 U7011 ( .IN1(WX5997), .IN2(test_so47), .Q(n6009) );
  NAND2X0 U7012 ( .IN1(n3893), .IN2(n6010), .QN(n6007) );
  NAND2X0 U7013 ( .IN1(n215), .IN2(n3924), .QN(n6006) );
  INVX0 U7014 ( .INP(n6011), .ZN(n215) );
  NAND2X0 U7015 ( .IN1(n4456), .IN2(n8560), .QN(n6011) );
  NAND2X0 U7016 ( .IN1(test_so42), .IN2(n3957), .QN(n6005) );
  NAND4X0 U7017 ( .IN1(n6012), .IN2(n6013), .IN3(n6014), .IN4(n6015), .QN(
        WX4573) );
  NAND2X0 U7018 ( .IN1(n3968), .IN2(n5762), .QN(n6015) );
  XNOR3X1 U7019 ( .IN1(n3660), .IN2(n3350), .IN3(n6016), .Q(n5762) );
  XOR2X1 U7020 ( .IN1(WX5931), .IN2(n7168), .Q(n6016) );
  NAND2X0 U7021 ( .IN1(n3893), .IN2(n6017), .QN(n6014) );
  NAND2X0 U7022 ( .IN1(n214), .IN2(n3924), .QN(n6013) );
  INVX0 U7023 ( .INP(n6018), .ZN(n214) );
  NAND2X0 U7024 ( .IN1(n4458), .IN2(n8561), .QN(n6018) );
  NAND2X0 U7025 ( .IN1(n3936), .IN2(CRC_OUT_6_6), .QN(n6012) );
  NAND4X0 U7026 ( .IN1(n6019), .IN2(n6020), .IN3(n6021), .IN4(n6022), .QN(
        WX4571) );
  NAND2X0 U7027 ( .IN1(n3968), .IN2(n5769), .QN(n6022) );
  XNOR3X1 U7028 ( .IN1(n3658), .IN2(n3351), .IN3(n6023), .Q(n5769) );
  XOR2X1 U7029 ( .IN1(WX5929), .IN2(n7169), .Q(n6023) );
  NAND2X0 U7030 ( .IN1(n3893), .IN2(n6024), .QN(n6021) );
  NAND2X0 U7031 ( .IN1(n213), .IN2(n3924), .QN(n6020) );
  INVX0 U7032 ( .INP(n6025), .ZN(n213) );
  NAND2X0 U7033 ( .IN1(n4458), .IN2(n8562), .QN(n6025) );
  NAND2X0 U7034 ( .IN1(n3936), .IN2(CRC_OUT_6_7), .QN(n6019) );
  NAND4X0 U7035 ( .IN1(n6026), .IN2(n6027), .IN3(n6028), .IN4(n6029), .QN(
        WX4569) );
  NAND2X0 U7036 ( .IN1(n3968), .IN2(n5776), .QN(n6029) );
  XNOR3X1 U7037 ( .IN1(n3656), .IN2(n3352), .IN3(n6030), .Q(n5776) );
  XOR2X1 U7038 ( .IN1(WX5927), .IN2(n7170), .Q(n6030) );
  NAND2X0 U7039 ( .IN1(n3895), .IN2(n6031), .QN(n6028) );
  NAND2X0 U7040 ( .IN1(n212), .IN2(n3924), .QN(n6027) );
  INVX0 U7041 ( .INP(n6032), .ZN(n212) );
  NAND2X0 U7042 ( .IN1(n4457), .IN2(n8563), .QN(n6032) );
  NAND2X0 U7043 ( .IN1(n3936), .IN2(CRC_OUT_6_8), .QN(n6026) );
  NAND4X0 U7044 ( .IN1(n6033), .IN2(n6034), .IN3(n6035), .IN4(n6036), .QN(
        WX4567) );
  NAND2X0 U7045 ( .IN1(n3968), .IN2(n5783), .QN(n6036) );
  XNOR3X1 U7046 ( .IN1(n3654), .IN2(n3353), .IN3(n6037), .Q(n5783) );
  XOR2X1 U7047 ( .IN1(WX5925), .IN2(n7171), .Q(n6037) );
  NAND2X0 U7048 ( .IN1(n3894), .IN2(n6038), .QN(n6035) );
  NAND2X0 U7049 ( .IN1(n211), .IN2(n3924), .QN(n6034) );
  INVX0 U7050 ( .INP(n6039), .ZN(n211) );
  NAND2X0 U7051 ( .IN1(n4457), .IN2(n8564), .QN(n6039) );
  NAND2X0 U7052 ( .IN1(n3936), .IN2(CRC_OUT_6_9), .QN(n6033) );
  NAND4X0 U7053 ( .IN1(n6040), .IN2(n6041), .IN3(n6042), .IN4(n6043), .QN(
        WX4565) );
  NAND2X0 U7054 ( .IN1(n3968), .IN2(n5790), .QN(n6043) );
  XNOR3X1 U7055 ( .IN1(n3652), .IN2(n3354), .IN3(n6044), .Q(n5790) );
  XOR2X1 U7056 ( .IN1(WX5923), .IN2(n7172), .Q(n6044) );
  NAND2X0 U7057 ( .IN1(n3894), .IN2(n6045), .QN(n6042) );
  NAND2X0 U7058 ( .IN1(n210), .IN2(n3924), .QN(n6041) );
  INVX0 U7059 ( .INP(n6046), .ZN(n210) );
  NAND2X0 U7060 ( .IN1(n4457), .IN2(n8565), .QN(n6046) );
  NAND2X0 U7061 ( .IN1(n3936), .IN2(CRC_OUT_6_10), .QN(n6040) );
  NAND4X0 U7062 ( .IN1(n6047), .IN2(n6048), .IN3(n6049), .IN4(n6050), .QN(
        WX4563) );
  NAND2X0 U7063 ( .IN1(n3968), .IN2(n5797), .QN(n6050) );
  XNOR3X1 U7064 ( .IN1(n3423), .IN2(n3355), .IN3(n6051), .Q(n5797) );
  XOR2X1 U7065 ( .IN1(WX5921), .IN2(n7173), .Q(n6051) );
  NAND2X0 U7066 ( .IN1(n6052), .IN2(n3899), .QN(n6049) );
  NAND2X0 U7067 ( .IN1(n209), .IN2(n3924), .QN(n6048) );
  INVX0 U7068 ( .INP(n6053), .ZN(n209) );
  NAND2X0 U7069 ( .IN1(n4457), .IN2(n8566), .QN(n6053) );
  NAND2X0 U7070 ( .IN1(n3936), .IN2(CRC_OUT_6_11), .QN(n6047) );
  NAND4X0 U7071 ( .IN1(n6054), .IN2(n6055), .IN3(n6056), .IN4(n6057), .QN(
        WX4561) );
  NAND2X0 U7072 ( .IN1(n3968), .IN2(n5804), .QN(n6057) );
  XNOR3X1 U7073 ( .IN1(n3650), .IN2(n3356), .IN3(n6058), .Q(n5804) );
  XOR2X1 U7074 ( .IN1(WX5919), .IN2(n7174), .Q(n6058) );
  NAND2X0 U7075 ( .IN1(n3894), .IN2(n6059), .QN(n6056) );
  NAND2X0 U7076 ( .IN1(n208), .IN2(n3924), .QN(n6055) );
  INVX0 U7077 ( .INP(n6060), .ZN(n208) );
  NAND2X0 U7078 ( .IN1(n4457), .IN2(n8567), .QN(n6060) );
  NAND2X0 U7079 ( .IN1(n3936), .IN2(CRC_OUT_6_12), .QN(n6054) );
  NAND4X0 U7080 ( .IN1(n6061), .IN2(n6062), .IN3(n6063), .IN4(n6064), .QN(
        WX4559) );
  NAND2X0 U7081 ( .IN1(n3968), .IN2(n5811), .QN(n6064) );
  XNOR3X1 U7082 ( .IN1(n3648), .IN2(n3357), .IN3(n6065), .Q(n5811) );
  XOR2X1 U7083 ( .IN1(WX5917), .IN2(n7175), .Q(n6065) );
  NAND2X0 U7084 ( .IN1(n6066), .IN2(n3899), .QN(n6063) );
  NAND2X0 U7085 ( .IN1(n207), .IN2(n3924), .QN(n6062) );
  INVX0 U7086 ( .INP(n6067), .ZN(n207) );
  NAND2X0 U7087 ( .IN1(n4457), .IN2(n8568), .QN(n6067) );
  NAND2X0 U7088 ( .IN1(n3936), .IN2(CRC_OUT_6_13), .QN(n6061) );
  NAND4X0 U7089 ( .IN1(n6068), .IN2(n6069), .IN3(n6070), .IN4(n6071), .QN(
        WX4557) );
  NAND2X0 U7090 ( .IN1(n3969), .IN2(n5818), .QN(n6071) );
  XNOR3X1 U7091 ( .IN1(n3646), .IN2(n3358), .IN3(n6072), .Q(n5818) );
  XOR2X1 U7092 ( .IN1(WX5915), .IN2(n7176), .Q(n6072) );
  NAND2X0 U7093 ( .IN1(n3894), .IN2(n6073), .QN(n6070) );
  NAND2X0 U7094 ( .IN1(n206), .IN2(n3925), .QN(n6069) );
  INVX0 U7095 ( .INP(n6074), .ZN(n206) );
  NAND2X0 U7096 ( .IN1(n4457), .IN2(n8569), .QN(n6074) );
  NAND2X0 U7097 ( .IN1(n3936), .IN2(CRC_OUT_6_14), .QN(n6068) );
  NAND4X0 U7098 ( .IN1(n6075), .IN2(n6076), .IN3(n6077), .IN4(n6078), .QN(
        WX4555) );
  NAND2X0 U7099 ( .IN1(n3969), .IN2(n5825), .QN(n6078) );
  XNOR3X1 U7100 ( .IN1(n3644), .IN2(n3359), .IN3(n6079), .Q(n5825) );
  XOR2X1 U7101 ( .IN1(WX5913), .IN2(n7177), .Q(n6079) );
  NAND2X0 U7102 ( .IN1(n6080), .IN2(n3899), .QN(n6077) );
  NAND2X0 U7103 ( .IN1(n205), .IN2(n3925), .QN(n6076) );
  INVX0 U7104 ( .INP(n6081), .ZN(n205) );
  NAND2X0 U7105 ( .IN1(n4457), .IN2(n8570), .QN(n6081) );
  NAND2X0 U7106 ( .IN1(n3936), .IN2(CRC_OUT_6_15), .QN(n6075) );
  NAND4X0 U7107 ( .IN1(n6082), .IN2(n6083), .IN3(n6084), .IN4(n6085), .QN(
        WX4553) );
  NAND2X0 U7108 ( .IN1(n5832), .IN2(n3987), .QN(n6085) );
  XOR3X1 U7109 ( .IN1(n3182), .IN2(TM1), .IN3(n6086), .Q(n5832) );
  XOR3X1 U7110 ( .IN1(test_so52), .IN2(n7178), .IN3(WX5975), .Q(n6086) );
  NAND2X0 U7111 ( .IN1(n3894), .IN2(n6087), .QN(n6084) );
  NAND2X0 U7112 ( .IN1(n204), .IN2(n3925), .QN(n6083) );
  INVX0 U7113 ( .INP(n6088), .ZN(n204) );
  NAND2X0 U7114 ( .IN1(n4456), .IN2(n8571), .QN(n6088) );
  NAND2X0 U7115 ( .IN1(n3936), .IN2(CRC_OUT_6_16), .QN(n6082) );
  NAND4X0 U7116 ( .IN1(n6089), .IN2(n6090), .IN3(n6091), .IN4(n6092), .QN(
        WX4551) );
  NAND2X0 U7117 ( .IN1(n3969), .IN2(n5839), .QN(n6092) );
  XOR3X1 U7118 ( .IN1(n3183), .IN2(n3873), .IN3(n6093), .Q(n5839) );
  XOR3X1 U7119 ( .IN1(n7179), .IN2(n3643), .IN3(WX5973), .Q(n6093) );
  NAND2X0 U7120 ( .IN1(n6094), .IN2(n3899), .QN(n6091) );
  NAND2X0 U7121 ( .IN1(n203), .IN2(n3925), .QN(n6090) );
  INVX0 U7122 ( .INP(n6095), .ZN(n203) );
  NAND2X0 U7123 ( .IN1(n4457), .IN2(n8572), .QN(n6095) );
  NAND2X0 U7124 ( .IN1(n3936), .IN2(CRC_OUT_6_17), .QN(n6089) );
  NAND4X0 U7125 ( .IN1(n6096), .IN2(n6097), .IN3(n6098), .IN4(n6099), .QN(
        WX4549) );
  NAND2X0 U7126 ( .IN1(n5846), .IN2(n3987), .QN(n6099) );
  XOR3X1 U7127 ( .IN1(n3185), .IN2(TM1), .IN3(n6100), .Q(n5846) );
  XNOR3X1 U7128 ( .IN1(test_so50), .IN2(n7180), .IN3(n3642), .Q(n6100) );
  NAND2X0 U7129 ( .IN1(n3894), .IN2(n6101), .QN(n6098) );
  NAND2X0 U7130 ( .IN1(n202), .IN2(n3925), .QN(n6097) );
  INVX0 U7131 ( .INP(n6102), .ZN(n202) );
  NAND2X0 U7132 ( .IN1(n4456), .IN2(n8573), .QN(n6102) );
  NAND2X0 U7133 ( .IN1(n3937), .IN2(CRC_OUT_6_18), .QN(n6096) );
  NAND4X0 U7134 ( .IN1(n6103), .IN2(n6104), .IN3(n6105), .IN4(n6106), .QN(
        WX4547) );
  NAND2X0 U7135 ( .IN1(n3969), .IN2(n5853), .QN(n6106) );
  XOR3X1 U7136 ( .IN1(n3186), .IN2(n3872), .IN3(n6107), .Q(n5853) );
  XOR3X1 U7137 ( .IN1(n7181), .IN2(n3640), .IN3(WX5969), .Q(n6107) );
  NAND2X0 U7138 ( .IN1(n3894), .IN2(n6108), .QN(n6105) );
  NAND2X0 U7139 ( .IN1(n201), .IN2(n3925), .QN(n6104) );
  INVX0 U7140 ( .INP(n6109), .ZN(n201) );
  NAND2X0 U7141 ( .IN1(test_so33), .IN2(n4463), .QN(n6109) );
  NAND2X0 U7142 ( .IN1(n3937), .IN2(CRC_OUT_6_19), .QN(n6103) );
  NAND4X0 U7143 ( .IN1(n6110), .IN2(n6111), .IN3(n6112), .IN4(n6113), .QN(
        WX4545) );
  NAND2X0 U7144 ( .IN1(n5860), .IN2(n3987), .QN(n6113) );
  XOR3X1 U7145 ( .IN1(n3188), .IN2(TM1), .IN3(n6114), .Q(n5860) );
  XNOR3X1 U7146 ( .IN1(test_so48), .IN2(n7182), .IN3(n3638), .Q(n6114) );
  NAND2X0 U7147 ( .IN1(n3894), .IN2(n6115), .QN(n6112) );
  NAND2X0 U7148 ( .IN1(n200), .IN2(n3925), .QN(n6111) );
  INVX0 U7149 ( .INP(n6116), .ZN(n200) );
  NAND2X0 U7150 ( .IN1(n4456), .IN2(n8576), .QN(n6116) );
  NAND2X0 U7151 ( .IN1(n3937), .IN2(CRC_OUT_6_20), .QN(n6110) );
  NAND4X0 U7152 ( .IN1(n6117), .IN2(n6118), .IN3(n6119), .IN4(n6120), .QN(
        WX4543) );
  NAND2X0 U7153 ( .IN1(n3969), .IN2(n5867), .QN(n6120) );
  XOR3X1 U7154 ( .IN1(n3189), .IN2(n3875), .IN3(n6121), .Q(n5867) );
  XOR3X1 U7155 ( .IN1(n7183), .IN2(n3636), .IN3(WX5965), .Q(n6121) );
  NAND2X0 U7156 ( .IN1(n3894), .IN2(n6122), .QN(n6119) );
  NAND2X0 U7157 ( .IN1(n199), .IN2(n3925), .QN(n6118) );
  INVX0 U7158 ( .INP(n6123), .ZN(n199) );
  NAND2X0 U7159 ( .IN1(n4456), .IN2(n8577), .QN(n6123) );
  NAND2X0 U7160 ( .IN1(n3937), .IN2(CRC_OUT_6_21), .QN(n6117) );
  NAND4X0 U7161 ( .IN1(n6124), .IN2(n6125), .IN3(n6126), .IN4(n6127), .QN(
        WX4541) );
  NAND2X0 U7162 ( .IN1(n5874), .IN2(n3987), .QN(n6127) );
  XOR3X1 U7163 ( .IN1(n3191), .IN2(TM1), .IN3(n6128), .Q(n5874) );
  XNOR3X1 U7164 ( .IN1(test_so46), .IN2(n7184), .IN3(n3634), .Q(n6128) );
  NAND2X0 U7165 ( .IN1(n3894), .IN2(n6129), .QN(n6126) );
  NAND2X0 U7166 ( .IN1(n198), .IN2(n3925), .QN(n6125) );
  INVX0 U7167 ( .INP(n6130), .ZN(n198) );
  NAND2X0 U7168 ( .IN1(n4456), .IN2(n8578), .QN(n6130) );
  NAND2X0 U7169 ( .IN1(test_so43), .IN2(n3956), .QN(n6124) );
  NAND4X0 U7170 ( .IN1(n6131), .IN2(n6132), .IN3(n6133), .IN4(n6134), .QN(
        WX4539) );
  NAND2X0 U7171 ( .IN1(n3969), .IN2(n5881), .QN(n6134) );
  XOR3X1 U7172 ( .IN1(n3192), .IN2(n3874), .IN3(n6135), .Q(n5881) );
  XOR3X1 U7173 ( .IN1(n7185), .IN2(n3632), .IN3(WX5961), .Q(n6135) );
  NAND2X0 U7174 ( .IN1(n3894), .IN2(n6136), .QN(n6133) );
  NAND2X0 U7175 ( .IN1(n197), .IN2(n3925), .QN(n6132) );
  INVX0 U7176 ( .INP(n6137), .ZN(n197) );
  NAND2X0 U7177 ( .IN1(n4456), .IN2(n8579), .QN(n6137) );
  NAND2X0 U7178 ( .IN1(n3937), .IN2(CRC_OUT_6_23), .QN(n6131) );
  NAND4X0 U7179 ( .IN1(n6138), .IN2(n6139), .IN3(n6140), .IN4(n6141), .QN(
        WX4537) );
  NAND2X0 U7180 ( .IN1(n3969), .IN2(n5888), .QN(n6141) );
  XOR3X1 U7181 ( .IN1(n3194), .IN2(n3873), .IN3(n6142), .Q(n5888) );
  XOR3X1 U7182 ( .IN1(n7186), .IN2(n3630), .IN3(WX5959), .Q(n6142) );
  NAND2X0 U7183 ( .IN1(n3894), .IN2(n6143), .QN(n6140) );
  NAND2X0 U7184 ( .IN1(n196), .IN2(n3925), .QN(n6139) );
  INVX0 U7185 ( .INP(n6144), .ZN(n196) );
  NAND2X0 U7186 ( .IN1(n4456), .IN2(n8580), .QN(n6144) );
  NAND2X0 U7187 ( .IN1(n3937), .IN2(CRC_OUT_6_24), .QN(n6138) );
  NAND4X0 U7188 ( .IN1(n6145), .IN2(n6146), .IN3(n6147), .IN4(n6148), .QN(
        WX4535) );
  NAND2X0 U7189 ( .IN1(n3969), .IN2(n5895), .QN(n6148) );
  XOR3X1 U7190 ( .IN1(n3196), .IN2(n3872), .IN3(n6149), .Q(n5895) );
  XOR3X1 U7191 ( .IN1(n7187), .IN2(n3628), .IN3(WX5957), .Q(n6149) );
  NAND2X0 U7192 ( .IN1(n3895), .IN2(n6150), .QN(n6147) );
  NAND2X0 U7193 ( .IN1(n195), .IN2(n3925), .QN(n6146) );
  INVX0 U7194 ( .INP(n6151), .ZN(n195) );
  NAND2X0 U7195 ( .IN1(n4456), .IN2(n8581), .QN(n6151) );
  NAND2X0 U7196 ( .IN1(n3937), .IN2(CRC_OUT_6_25), .QN(n6145) );
  NAND4X0 U7197 ( .IN1(n6152), .IN2(n6153), .IN3(n6154), .IN4(n6155), .QN(
        WX4533) );
  NAND2X0 U7198 ( .IN1(n3969), .IN2(n5902), .QN(n6155) );
  XOR3X1 U7199 ( .IN1(n3198), .IN2(n3875), .IN3(n6156), .Q(n5902) );
  XOR3X1 U7200 ( .IN1(n7188), .IN2(n3626), .IN3(WX5955), .Q(n6156) );
  NAND2X0 U7201 ( .IN1(n3895), .IN2(n6157), .QN(n6154) );
  NAND2X0 U7202 ( .IN1(n194), .IN2(n3925), .QN(n6153) );
  INVX0 U7203 ( .INP(n6158), .ZN(n194) );
  NAND2X0 U7204 ( .IN1(n4455), .IN2(n8582), .QN(n6158) );
  NAND2X0 U7205 ( .IN1(n3937), .IN2(CRC_OUT_6_26), .QN(n6152) );
  NAND4X0 U7206 ( .IN1(n6159), .IN2(n6160), .IN3(n6161), .IN4(n6162), .QN(
        WX4531) );
  NAND2X0 U7207 ( .IN1(n3969), .IN2(n5909), .QN(n6162) );
  XOR3X1 U7208 ( .IN1(n3200), .IN2(n3874), .IN3(n6163), .Q(n5909) );
  XOR3X1 U7209 ( .IN1(n7189), .IN2(n3624), .IN3(WX5953), .Q(n6163) );
  NAND2X0 U7210 ( .IN1(n3895), .IN2(n6164), .QN(n6161) );
  NAND2X0 U7211 ( .IN1(n193), .IN2(n3925), .QN(n6160) );
  INVX0 U7212 ( .INP(n6165), .ZN(n193) );
  NAND2X0 U7213 ( .IN1(n4455), .IN2(n8583), .QN(n6165) );
  NAND2X0 U7214 ( .IN1(n3937), .IN2(CRC_OUT_6_27), .QN(n6159) );
  NAND4X0 U7215 ( .IN1(n6166), .IN2(n6167), .IN3(n6168), .IN4(n6169), .QN(
        WX4529) );
  NAND2X0 U7216 ( .IN1(n3969), .IN2(n5916), .QN(n6169) );
  XOR3X1 U7217 ( .IN1(n3202), .IN2(n3873), .IN3(n6170), .Q(n5916) );
  XOR3X1 U7218 ( .IN1(n7190), .IN2(n3622), .IN3(WX5951), .Q(n6170) );
  NAND2X0 U7219 ( .IN1(n6171), .IN2(n3898), .QN(n6168) );
  NAND2X0 U7220 ( .IN1(n192), .IN2(n3925), .QN(n6167) );
  INVX0 U7221 ( .INP(n6172), .ZN(n192) );
  NAND2X0 U7222 ( .IN1(n4455), .IN2(n8584), .QN(n6172) );
  NAND2X0 U7223 ( .IN1(n3937), .IN2(CRC_OUT_6_28), .QN(n6166) );
  NAND4X0 U7224 ( .IN1(n6173), .IN2(n6174), .IN3(n6175), .IN4(n6176), .QN(
        WX4527) );
  NAND2X0 U7225 ( .IN1(n3970), .IN2(n5923), .QN(n6176) );
  XOR3X1 U7226 ( .IN1(n3204), .IN2(n3872), .IN3(n6177), .Q(n5923) );
  XOR3X1 U7227 ( .IN1(n7191), .IN2(n3621), .IN3(WX5949), .Q(n6177) );
  NAND2X0 U7228 ( .IN1(n3895), .IN2(n6178), .QN(n6175) );
  NAND2X0 U7229 ( .IN1(n191), .IN2(n3925), .QN(n6174) );
  INVX0 U7230 ( .INP(n6179), .ZN(n191) );
  NAND2X0 U7231 ( .IN1(n4455), .IN2(n8585), .QN(n6179) );
  NAND2X0 U7232 ( .IN1(n3937), .IN2(CRC_OUT_6_29), .QN(n6173) );
  NAND4X0 U7233 ( .IN1(n6180), .IN2(n6181), .IN3(n6182), .IN4(n6183), .QN(
        WX4525) );
  NAND2X0 U7234 ( .IN1(n3970), .IN2(n5930), .QN(n6183) );
  XOR3X1 U7235 ( .IN1(n3206), .IN2(n3875), .IN3(n6184), .Q(n5930) );
  XOR3X1 U7236 ( .IN1(n7192), .IN2(n3620), .IN3(WX5947), .Q(n6184) );
  NAND2X0 U7237 ( .IN1(n6185), .IN2(n3897), .QN(n6182) );
  NAND2X0 U7238 ( .IN1(n190), .IN2(n3925), .QN(n6181) );
  INVX0 U7239 ( .INP(n6186), .ZN(n190) );
  NAND2X0 U7240 ( .IN1(n4455), .IN2(n8586), .QN(n6186) );
  NAND2X0 U7241 ( .IN1(n3937), .IN2(CRC_OUT_6_30), .QN(n6180) );
  NAND4X0 U7242 ( .IN1(n6187), .IN2(n6188), .IN3(n6189), .IN4(n6190), .QN(
        WX4523) );
  NAND2X0 U7243 ( .IN1(n3970), .IN2(n5937), .QN(n6190) );
  XOR3X1 U7244 ( .IN1(n3068), .IN2(n3874), .IN3(n6191), .Q(n5937) );
  XOR3X1 U7245 ( .IN1(n7193), .IN2(n3618), .IN3(WX5945), .Q(n6191) );
  NAND2X0 U7246 ( .IN1(n3895), .IN2(n6192), .QN(n6189) );
  NAND2X0 U7247 ( .IN1(n3938), .IN2(CRC_OUT_6_31), .QN(n6188) );
  NAND2X0 U7248 ( .IN1(n2245), .IN2(WX4364), .QN(n6187) );
  NOR2X0 U7249 ( .IN1(n4566), .IN2(WX4364), .QN(WX4425) );
  NOR2X0 U7250 ( .IN1(n4567), .IN2(n6193), .QN(WX3912) );
  XOR2X1 U7251 ( .IN1(n3721), .IN2(DFF_574_n1), .Q(n6193) );
  NOR2X0 U7252 ( .IN1(n4567), .IN2(n6194), .QN(WX3910) );
  XOR2X1 U7253 ( .IN1(n3722), .IN2(DFF_573_n1), .Q(n6194) );
  NOR2X0 U7254 ( .IN1(n4567), .IN2(n6195), .QN(WX3908) );
  XOR2X1 U7255 ( .IN1(n3724), .IN2(DFF_572_n1), .Q(n6195) );
  NOR2X0 U7256 ( .IN1(n4567), .IN2(n6196), .QN(WX3906) );
  XNOR2X1 U7257 ( .IN1(n3726), .IN2(test_so32), .Q(n6196) );
  NOR2X0 U7258 ( .IN1(n4567), .IN2(n6197), .QN(WX3904) );
  XOR2X1 U7259 ( .IN1(n3728), .IN2(DFF_570_n1), .Q(n6197) );
  NOR2X0 U7260 ( .IN1(n4567), .IN2(n6198), .QN(WX3902) );
  XOR2X1 U7261 ( .IN1(n3730), .IN2(DFF_569_n1), .Q(n6198) );
  NOR2X0 U7262 ( .IN1(n4567), .IN2(n6199), .QN(WX3900) );
  XOR2X1 U7263 ( .IN1(n3732), .IN2(DFF_568_n1), .Q(n6199) );
  NOR2X0 U7264 ( .IN1(n4567), .IN2(n6200), .QN(WX3898) );
  XOR2X1 U7265 ( .IN1(n3734), .IN2(DFF_567_n1), .Q(n6200) );
  NOR2X0 U7266 ( .IN1(n4567), .IN2(n6201), .QN(WX3896) );
  XOR2X1 U7267 ( .IN1(CRC_OUT_7_22), .IN2(test_so29), .Q(n6201) );
  NOR2X0 U7268 ( .IN1(n4567), .IN2(n6202), .QN(WX3894) );
  XOR2X1 U7269 ( .IN1(n3736), .IN2(DFF_565_n1), .Q(n6202) );
  NOR2X0 U7270 ( .IN1(n4567), .IN2(n6203), .QN(WX3892) );
  XOR2X1 U7271 ( .IN1(n3738), .IN2(DFF_564_n1), .Q(n6203) );
  NOR2X0 U7272 ( .IN1(n4567), .IN2(n6204), .QN(WX3890) );
  XOR2X1 U7273 ( .IN1(n3740), .IN2(DFF_563_n1), .Q(n6204) );
  NOR2X0 U7274 ( .IN1(n4567), .IN2(n6205), .QN(WX3888) );
  XOR2X1 U7275 ( .IN1(n3742), .IN2(DFF_562_n1), .Q(n6205) );
  NOR2X0 U7276 ( .IN1(n4567), .IN2(n6206), .QN(WX3886) );
  XOR2X1 U7277 ( .IN1(n3744), .IN2(DFF_561_n1), .Q(n6206) );
  NOR2X0 U7278 ( .IN1(n4567), .IN2(n6207), .QN(WX3884) );
  XOR2X1 U7279 ( .IN1(n3746), .IN2(DFF_560_n1), .Q(n6207) );
  NOR2X0 U7280 ( .IN1(n4567), .IN2(n6208), .QN(WX3882) );
  XOR3X1 U7281 ( .IN1(n3427), .IN2(DFF_575_n1), .IN3(CRC_OUT_7_15), .Q(n6208)
         );
  NOR2X0 U7282 ( .IN1(n4568), .IN2(n6209), .QN(WX3880) );
  XOR2X1 U7283 ( .IN1(n3747), .IN2(DFF_558_n1), .Q(n6209) );
  NOR2X0 U7284 ( .IN1(n4568), .IN2(n6210), .QN(WX3878) );
  XOR2X1 U7285 ( .IN1(n3748), .IN2(DFF_557_n1), .Q(n6210) );
  NOR2X0 U7286 ( .IN1(n4568), .IN2(n6211), .QN(WX3876) );
  XOR2X1 U7287 ( .IN1(n3750), .IN2(DFF_556_n1), .Q(n6211) );
  NOR2X0 U7288 ( .IN1(n4568), .IN2(n6212), .QN(WX3874) );
  XOR2X1 U7289 ( .IN1(n3752), .IN2(DFF_555_n1), .Q(n6212) );
  NOR2X0 U7290 ( .IN1(n4568), .IN2(n6213), .QN(WX3872) );
  XOR3X1 U7291 ( .IN1(test_so31), .IN2(n3428), .IN3(DFF_575_n1), .Q(n6213) );
  NOR2X0 U7292 ( .IN1(n4568), .IN2(n6214), .QN(WX3870) );
  XOR2X1 U7293 ( .IN1(n3754), .IN2(DFF_553_n1), .Q(n6214) );
  NOR2X0 U7294 ( .IN1(n4568), .IN2(n6215), .QN(WX3868) );
  XOR2X1 U7295 ( .IN1(n3755), .IN2(DFF_552_n1), .Q(n6215) );
  NOR2X0 U7296 ( .IN1(n4568), .IN2(n6216), .QN(WX3866) );
  XOR2X1 U7297 ( .IN1(n3756), .IN2(DFF_551_n1), .Q(n6216) );
  NOR2X0 U7298 ( .IN1(n4568), .IN2(n6217), .QN(WX3864) );
  XOR2X1 U7299 ( .IN1(n3758), .IN2(DFF_550_n1), .Q(n6217) );
  NOR2X0 U7300 ( .IN1(n4568), .IN2(n6218), .QN(WX3862) );
  XOR2X1 U7301 ( .IN1(CRC_OUT_7_5), .IN2(test_so30), .Q(n6218) );
  NOR2X0 U7302 ( .IN1(n4568), .IN2(n6219), .QN(WX3860) );
  XOR2X1 U7303 ( .IN1(n3760), .IN2(DFF_548_n1), .Q(n6219) );
  NOR2X0 U7304 ( .IN1(n4568), .IN2(n6220), .QN(WX3858) );
  XOR3X1 U7305 ( .IN1(n3429), .IN2(DFF_575_n1), .IN3(CRC_OUT_7_3), .Q(n6220)
         );
  NOR2X0 U7306 ( .IN1(n4554), .IN2(n6221), .QN(WX3856) );
  XOR2X1 U7307 ( .IN1(n3762), .IN2(DFF_546_n1), .Q(n6221) );
  NOR2X0 U7308 ( .IN1(n4554), .IN2(n6222), .QN(WX3854) );
  XOR2X1 U7309 ( .IN1(n3764), .IN2(DFF_545_n1), .Q(n6222) );
  NOR2X0 U7310 ( .IN1(n4553), .IN2(n6223), .QN(WX3852) );
  XOR2X1 U7311 ( .IN1(n3766), .IN2(DFF_544_n1), .Q(n6223) );
  NOR2X0 U7312 ( .IN1(n4553), .IN2(n6224), .QN(WX3850) );
  XOR2X1 U7313 ( .IN1(n3439), .IN2(DFF_575_n1), .Q(n6224) );
  NAND4X0 U7314 ( .IN1(n6225), .IN2(n6226), .IN3(n6227), .IN4(n6228), .QN(
        WX3292) );
  NAND2X0 U7315 ( .IN1(n5975), .IN2(n3986), .QN(n6228) );
  XOR3X1 U7316 ( .IN1(n3691), .IN2(n3438), .IN3(n6229), .Q(n5975) );
  XOR2X1 U7317 ( .IN1(WX4714), .IN2(test_so36), .Q(n6229) );
  NAND2X0 U7318 ( .IN1(n3895), .IN2(n6230), .QN(n6227) );
  NAND2X0 U7319 ( .IN1(n142), .IN2(n3926), .QN(n6226) );
  INVX0 U7320 ( .INP(n6231), .ZN(n142) );
  NAND2X0 U7321 ( .IN1(n4455), .IN2(n8612), .QN(n6231) );
  NAND2X0 U7322 ( .IN1(n3938), .IN2(CRC_OUT_7_0), .QN(n6225) );
  NAND4X0 U7323 ( .IN1(n6232), .IN2(n6233), .IN3(n6234), .IN4(n6235), .QN(
        WX3290) );
  NAND2X0 U7324 ( .IN1(n3970), .IN2(n5982), .QN(n6235) );
  XNOR3X1 U7325 ( .IN1(n3693), .IN2(n3360), .IN3(n6236), .Q(n5982) );
  XOR2X1 U7326 ( .IN1(WX4712), .IN2(n3720), .Q(n6236) );
  NAND2X0 U7327 ( .IN1(n3895), .IN2(n6237), .QN(n6234) );
  NAND2X0 U7328 ( .IN1(n141), .IN2(n3926), .QN(n6233) );
  INVX0 U7329 ( .INP(n6238), .ZN(n141) );
  NAND2X0 U7330 ( .IN1(n4455), .IN2(n8613), .QN(n6238) );
  NAND2X0 U7331 ( .IN1(n3938), .IN2(CRC_OUT_7_1), .QN(n6232) );
  NAND4X0 U7332 ( .IN1(n6239), .IN2(n6240), .IN3(n6241), .IN4(n6242), .QN(
        WX3288) );
  NAND2X0 U7333 ( .IN1(n3970), .IN2(n5989), .QN(n6242) );
  XNOR3X1 U7334 ( .IN1(n3695), .IN2(n3361), .IN3(n6243), .Q(n5989) );
  XOR2X1 U7335 ( .IN1(WX4710), .IN2(n3718), .Q(n6243) );
  NAND2X0 U7336 ( .IN1(n3895), .IN2(n6244), .QN(n6241) );
  NAND2X0 U7337 ( .IN1(n140), .IN2(n3926), .QN(n6240) );
  INVX0 U7338 ( .INP(n6245), .ZN(n140) );
  NAND2X0 U7339 ( .IN1(test_so23), .IN2(n4463), .QN(n6245) );
  NAND2X0 U7340 ( .IN1(n3938), .IN2(CRC_OUT_7_2), .QN(n6239) );
  NAND4X0 U7341 ( .IN1(n6246), .IN2(n6247), .IN3(n6248), .IN4(n6249), .QN(
        WX3286) );
  NAND2X0 U7342 ( .IN1(n3970), .IN2(n5996), .QN(n6249) );
  XNOR3X1 U7343 ( .IN1(n3697), .IN2(n3362), .IN3(n6250), .Q(n5996) );
  XOR2X1 U7344 ( .IN1(WX4708), .IN2(n3716), .Q(n6250) );
  NAND2X0 U7345 ( .IN1(n3895), .IN2(n6251), .QN(n6248) );
  NAND2X0 U7346 ( .IN1(n139), .IN2(n3926), .QN(n6247) );
  INVX0 U7347 ( .INP(n6252), .ZN(n139) );
  NAND2X0 U7348 ( .IN1(n4455), .IN2(n8616), .QN(n6252) );
  NAND2X0 U7349 ( .IN1(n3938), .IN2(CRC_OUT_7_3), .QN(n6246) );
  NAND4X0 U7350 ( .IN1(n6253), .IN2(n6254), .IN3(n6255), .IN4(n6256), .QN(
        WX3284) );
  NAND2X0 U7351 ( .IN1(n3970), .IN2(n6003), .QN(n6256) );
  XNOR3X1 U7352 ( .IN1(n3426), .IN2(n3363), .IN3(n6257), .Q(n6003) );
  XOR2X1 U7353 ( .IN1(WX4642), .IN2(n7194), .Q(n6257) );
  NAND2X0 U7354 ( .IN1(n3895), .IN2(n6258), .QN(n6255) );
  NAND2X0 U7355 ( .IN1(n138), .IN2(n3926), .QN(n6254) );
  INVX0 U7356 ( .INP(n6259), .ZN(n138) );
  NAND2X0 U7357 ( .IN1(n4455), .IN2(n8617), .QN(n6259) );
  NAND2X0 U7358 ( .IN1(n3938), .IN2(CRC_OUT_7_4), .QN(n6253) );
  NAND4X0 U7359 ( .IN1(n6260), .IN2(n6261), .IN3(n6262), .IN4(n6263), .QN(
        WX3282) );
  NAND2X0 U7360 ( .IN1(n3970), .IN2(n6010), .QN(n6263) );
  XNOR3X1 U7361 ( .IN1(n3701), .IN2(n3364), .IN3(n6264), .Q(n6010) );
  XOR2X1 U7362 ( .IN1(WX4704), .IN2(n3714), .Q(n6264) );
  NAND2X0 U7363 ( .IN1(n3895), .IN2(n6265), .QN(n6262) );
  NAND2X0 U7364 ( .IN1(n137), .IN2(n3926), .QN(n6261) );
  INVX0 U7365 ( .INP(n6266), .ZN(n137) );
  NAND2X0 U7366 ( .IN1(n4454), .IN2(n8618), .QN(n6266) );
  NAND2X0 U7367 ( .IN1(n3938), .IN2(CRC_OUT_7_5), .QN(n6260) );
  NAND4X0 U7368 ( .IN1(n6267), .IN2(n6268), .IN3(n6269), .IN4(n6270), .QN(
        WX3280) );
  NAND2X0 U7369 ( .IN1(n3970), .IN2(n6017), .QN(n6270) );
  XNOR3X1 U7370 ( .IN1(n3703), .IN2(n3365), .IN3(n6271), .Q(n6017) );
  XOR2X1 U7371 ( .IN1(WX4702), .IN2(n3712), .Q(n6271) );
  NAND2X0 U7372 ( .IN1(n6272), .IN2(n3897), .QN(n6269) );
  NAND2X0 U7373 ( .IN1(n136), .IN2(n3926), .QN(n6268) );
  INVX0 U7374 ( .INP(n6273), .ZN(n136) );
  NAND2X0 U7375 ( .IN1(n4454), .IN2(n8619), .QN(n6273) );
  NAND2X0 U7376 ( .IN1(n3938), .IN2(CRC_OUT_7_6), .QN(n6267) );
  NAND4X0 U7377 ( .IN1(n6274), .IN2(n6275), .IN3(n6276), .IN4(n6277), .QN(
        WX3278) );
  NAND2X0 U7378 ( .IN1(n3970), .IN2(n6024), .QN(n6277) );
  XNOR3X1 U7379 ( .IN1(n3705), .IN2(n3366), .IN3(n6278), .Q(n6024) );
  XOR2X1 U7380 ( .IN1(WX4700), .IN2(n3710), .Q(n6278) );
  NAND2X0 U7381 ( .IN1(n3896), .IN2(n6279), .QN(n6276) );
  NAND2X0 U7382 ( .IN1(n135), .IN2(n3926), .QN(n6275) );
  INVX0 U7383 ( .INP(n6280), .ZN(n135) );
  NAND2X0 U7384 ( .IN1(n4454), .IN2(n8620), .QN(n6280) );
  NAND2X0 U7385 ( .IN1(n3938), .IN2(CRC_OUT_7_7), .QN(n6274) );
  NAND4X0 U7386 ( .IN1(n6281), .IN2(n6282), .IN3(n6283), .IN4(n6284), .QN(
        WX3276) );
  NAND2X0 U7387 ( .IN1(n3970), .IN2(n6031), .QN(n6284) );
  XNOR3X1 U7388 ( .IN1(n3707), .IN2(n3367), .IN3(n6285), .Q(n6031) );
  XOR2X1 U7389 ( .IN1(WX4698), .IN2(n3708), .Q(n6285) );
  NAND2X0 U7390 ( .IN1(n6286), .IN2(n3898), .QN(n6283) );
  NAND2X0 U7391 ( .IN1(n134), .IN2(n3926), .QN(n6282) );
  INVX0 U7392 ( .INP(n6287), .ZN(n134) );
  NAND2X0 U7393 ( .IN1(n4454), .IN2(n8621), .QN(n6287) );
  NAND2X0 U7394 ( .IN1(n3938), .IN2(CRC_OUT_7_8), .QN(n6281) );
  NAND4X0 U7395 ( .IN1(n6288), .IN2(n6289), .IN3(n6290), .IN4(n6291), .QN(
        WX3274) );
  NAND2X0 U7396 ( .IN1(n3970), .IN2(n6038), .QN(n6291) );
  XNOR3X1 U7397 ( .IN1(n3706), .IN2(n3368), .IN3(n6292), .Q(n6038) );
  XOR2X1 U7398 ( .IN1(WX4632), .IN2(n7195), .Q(n6292) );
  NAND2X0 U7399 ( .IN1(n3896), .IN2(n6293), .QN(n6290) );
  NAND2X0 U7400 ( .IN1(n133), .IN2(n3926), .QN(n6289) );
  INVX0 U7401 ( .INP(n6294), .ZN(n133) );
  NAND2X0 U7402 ( .IN1(n4454), .IN2(n8622), .QN(n6294) );
  NAND2X0 U7403 ( .IN1(n3938), .IN2(CRC_OUT_7_9), .QN(n6288) );
  NAND4X0 U7404 ( .IN1(n6295), .IN2(n6296), .IN3(n6297), .IN4(n6298), .QN(
        WX3272) );
  NAND2X0 U7405 ( .IN1(n3971), .IN2(n6045), .QN(n6298) );
  XNOR3X1 U7406 ( .IN1(n3704), .IN2(n3369), .IN3(n6299), .Q(n6045) );
  XOR2X1 U7407 ( .IN1(WX4630), .IN2(n7196), .Q(n6299) );
  NAND2X0 U7408 ( .IN1(n3896), .IN2(n6300), .QN(n6297) );
  NAND2X0 U7409 ( .IN1(n132), .IN2(n3926), .QN(n6296) );
  INVX0 U7410 ( .INP(n6301), .ZN(n132) );
  NAND2X0 U7411 ( .IN1(n4454), .IN2(n8623), .QN(n6301) );
  NAND2X0 U7412 ( .IN1(test_so31), .IN2(n3957), .QN(n6295) );
  NAND4X0 U7413 ( .IN1(n6302), .IN2(n6303), .IN3(n6304), .IN4(n6305), .QN(
        WX3270) );
  NAND2X0 U7414 ( .IN1(n6052), .IN2(n3986), .QN(n6305) );
  XOR3X1 U7415 ( .IN1(n3713), .IN2(n3370), .IN3(n6306), .Q(n6052) );
  XOR2X1 U7416 ( .IN1(WX4564), .IN2(test_so41), .Q(n6306) );
  NAND2X0 U7417 ( .IN1(n3896), .IN2(n6307), .QN(n6304) );
  NAND2X0 U7418 ( .IN1(n131), .IN2(n3926), .QN(n6303) );
  INVX0 U7419 ( .INP(n6308), .ZN(n131) );
  NAND2X0 U7420 ( .IN1(n4454), .IN2(n8624), .QN(n6308) );
  NAND2X0 U7421 ( .IN1(n3938), .IN2(CRC_OUT_7_11), .QN(n6302) );
  NAND4X0 U7422 ( .IN1(n6309), .IN2(n6310), .IN3(n6311), .IN4(n6312), .QN(
        WX3268) );
  NAND2X0 U7423 ( .IN1(n3971), .IN2(n6059), .QN(n6312) );
  XNOR3X1 U7424 ( .IN1(n3702), .IN2(n3371), .IN3(n6313), .Q(n6059) );
  XOR2X1 U7425 ( .IN1(WX4626), .IN2(n7197), .Q(n6313) );
  NAND2X0 U7426 ( .IN1(n6314), .IN2(n3900), .QN(n6311) );
  NAND2X0 U7427 ( .IN1(n130), .IN2(n3926), .QN(n6310) );
  INVX0 U7428 ( .INP(n6315), .ZN(n130) );
  NAND2X0 U7429 ( .IN1(n4454), .IN2(n8625), .QN(n6315) );
  NAND2X0 U7430 ( .IN1(n3939), .IN2(CRC_OUT_7_12), .QN(n6309) );
  NAND4X0 U7431 ( .IN1(n6316), .IN2(n6317), .IN3(n6318), .IN4(n6319), .QN(
        WX3266) );
  NAND2X0 U7432 ( .IN1(n6066), .IN2(n3986), .QN(n6319) );
  XOR3X1 U7433 ( .IN1(n3717), .IN2(n3700), .IN3(n6320), .Q(n6066) );
  XOR2X1 U7434 ( .IN1(WX4560), .IN2(test_so39), .Q(n6320) );
  NAND2X0 U7435 ( .IN1(n3896), .IN2(n6321), .QN(n6318) );
  NAND2X0 U7436 ( .IN1(n129), .IN2(n3926), .QN(n6317) );
  INVX0 U7437 ( .INP(n6322), .ZN(n129) );
  NAND2X0 U7438 ( .IN1(n4453), .IN2(n8626), .QN(n6322) );
  NAND2X0 U7439 ( .IN1(n3939), .IN2(CRC_OUT_7_13), .QN(n6316) );
  NAND4X0 U7440 ( .IN1(n6323), .IN2(n6324), .IN3(n6325), .IN4(n6326), .QN(
        WX3264) );
  NAND2X0 U7441 ( .IN1(n3971), .IN2(n6073), .QN(n6326) );
  XNOR3X1 U7442 ( .IN1(n3698), .IN2(n3372), .IN3(n6327), .Q(n6073) );
  XOR2X1 U7443 ( .IN1(WX4622), .IN2(n7198), .Q(n6327) );
  NAND2X0 U7444 ( .IN1(n3896), .IN2(n6328), .QN(n6325) );
  NAND2X0 U7445 ( .IN1(n128), .IN2(n3926), .QN(n6324) );
  INVX0 U7446 ( .INP(n6329), .ZN(n128) );
  NAND2X0 U7447 ( .IN1(n4453), .IN2(n8627), .QN(n6329) );
  NAND2X0 U7448 ( .IN1(n3939), .IN2(CRC_OUT_7_14), .QN(n6323) );
  NAND4X0 U7449 ( .IN1(n6330), .IN2(n6331), .IN3(n6332), .IN4(n6333), .QN(
        WX3262) );
  NAND2X0 U7450 ( .IN1(n6080), .IN2(n3986), .QN(n6333) );
  XOR3X1 U7451 ( .IN1(n3696), .IN2(n3373), .IN3(n6334), .Q(n6080) );
  XOR2X1 U7452 ( .IN1(WX4556), .IN2(test_so37), .Q(n6334) );
  NAND2X0 U7453 ( .IN1(n3896), .IN2(n6335), .QN(n6332) );
  NAND2X0 U7454 ( .IN1(n126), .IN2(n3926), .QN(n6331) );
  INVX0 U7455 ( .INP(n6336), .ZN(n126) );
  NAND2X0 U7456 ( .IN1(n4453), .IN2(n8628), .QN(n6336) );
  NAND2X0 U7457 ( .IN1(n3939), .IN2(CRC_OUT_7_15), .QN(n6330) );
  NAND4X0 U7458 ( .IN1(n6337), .IN2(n6338), .IN3(n6339), .IN4(n6340), .QN(
        WX3260) );
  NAND2X0 U7459 ( .IN1(n3971), .IN2(n6087), .QN(n6340) );
  XOR3X1 U7460 ( .IN1(n3208), .IN2(n3873), .IN3(n6341), .Q(n6087) );
  XOR3X1 U7461 ( .IN1(n7199), .IN2(n3425), .IN3(WX4682), .Q(n6341) );
  NAND2X0 U7462 ( .IN1(n6342), .IN2(n3901), .QN(n6339) );
  NAND2X0 U7463 ( .IN1(n125), .IN2(n3926), .QN(n6338) );
  INVX0 U7464 ( .INP(n6343), .ZN(n125) );
  NAND2X0 U7465 ( .IN1(n4453), .IN2(n8629), .QN(n6343) );
  NAND2X0 U7466 ( .IN1(n3939), .IN2(CRC_OUT_7_16), .QN(n6337) );
  NAND4X0 U7467 ( .IN1(n6344), .IN2(n6345), .IN3(n6346), .IN4(n6347), .QN(
        WX3258) );
  NAND2X0 U7468 ( .IN1(n6094), .IN2(n3986), .QN(n6347) );
  XOR3X1 U7469 ( .IN1(n3210), .IN2(TM1), .IN3(n6348), .Q(n6094) );
  XNOR3X1 U7470 ( .IN1(test_so35), .IN2(n7200), .IN3(n3694), .Q(n6348) );
  NAND2X0 U7471 ( .IN1(n3893), .IN2(n6349), .QN(n6346) );
  NAND2X0 U7472 ( .IN1(n124), .IN2(n3927), .QN(n6345) );
  INVX0 U7473 ( .INP(n6350), .ZN(n124) );
  NAND2X0 U7474 ( .IN1(n4453), .IN2(n8630), .QN(n6350) );
  NAND2X0 U7475 ( .IN1(n3939), .IN2(CRC_OUT_7_17), .QN(n6344) );
  NAND4X0 U7476 ( .IN1(n6351), .IN2(n6352), .IN3(n6353), .IN4(n6354), .QN(
        WX3256) );
  NAND2X0 U7477 ( .IN1(n3971), .IN2(n6101), .QN(n6354) );
  XOR3X1 U7478 ( .IN1(n3211), .IN2(n3872), .IN3(n6355), .Q(n6101) );
  XOR3X1 U7479 ( .IN1(n7201), .IN2(n3692), .IN3(WX4678), .Q(n6355) );
  NAND2X0 U7480 ( .IN1(n3893), .IN2(n6356), .QN(n6353) );
  NAND2X0 U7481 ( .IN1(n123), .IN2(n3927), .QN(n6352) );
  INVX0 U7482 ( .INP(n6357), .ZN(n123) );
  NAND2X0 U7483 ( .IN1(n4453), .IN2(n8631), .QN(n6357) );
  NAND2X0 U7484 ( .IN1(n3939), .IN2(CRC_OUT_7_18), .QN(n6351) );
  NAND4X0 U7485 ( .IN1(n6358), .IN2(n6359), .IN3(n6360), .IN4(n6361), .QN(
        WX3254) );
  NAND2X0 U7486 ( .IN1(n3971), .IN2(n6108), .QN(n6361) );
  XOR3X1 U7487 ( .IN1(n3213), .IN2(n3875), .IN3(n6362), .Q(n6108) );
  XOR3X1 U7488 ( .IN1(n7202), .IN2(n3690), .IN3(WX4676), .Q(n6362) );
  NAND2X0 U7489 ( .IN1(n3893), .IN2(n6363), .QN(n6360) );
  NAND2X0 U7490 ( .IN1(n122), .IN2(n3927), .QN(n6359) );
  INVX0 U7491 ( .INP(n6364), .ZN(n122) );
  NAND2X0 U7492 ( .IN1(n4453), .IN2(n8632), .QN(n6364) );
  NAND2X0 U7493 ( .IN1(n3939), .IN2(CRC_OUT_7_19), .QN(n6358) );
  NAND4X0 U7494 ( .IN1(n6365), .IN2(n6366), .IN3(n6367), .IN4(n6368), .QN(
        WX3252) );
  NAND2X0 U7495 ( .IN1(n3971), .IN2(n6115), .QN(n6368) );
  XOR3X1 U7496 ( .IN1(n3215), .IN2(n3874), .IN3(n6369), .Q(n6115) );
  XOR3X1 U7497 ( .IN1(n7203), .IN2(n3688), .IN3(WX4674), .Q(n6369) );
  NAND2X0 U7498 ( .IN1(n3893), .IN2(n6370), .QN(n6367) );
  NAND2X0 U7499 ( .IN1(n121), .IN2(n3927), .QN(n6366) );
  INVX0 U7500 ( .INP(n6371), .ZN(n121) );
  NAND2X0 U7501 ( .IN1(test_so22), .IN2(n4463), .QN(n6371) );
  NAND2X0 U7502 ( .IN1(n3939), .IN2(CRC_OUT_7_20), .QN(n6365) );
  NAND4X0 U7503 ( .IN1(n6372), .IN2(n6373), .IN3(n6374), .IN4(n6375), .QN(
        WX3250) );
  NAND2X0 U7504 ( .IN1(n3971), .IN2(n6122), .QN(n6375) );
  XOR3X1 U7505 ( .IN1(n3217), .IN2(n3873), .IN3(n6376), .Q(n6122) );
  XOR3X1 U7506 ( .IN1(n7204), .IN2(n3686), .IN3(WX4672), .Q(n6376) );
  NAND2X0 U7507 ( .IN1(n3893), .IN2(n6377), .QN(n6374) );
  NAND2X0 U7508 ( .IN1(n120), .IN2(n3927), .QN(n6373) );
  INVX0 U7509 ( .INP(n6378), .ZN(n120) );
  NAND2X0 U7510 ( .IN1(n4453), .IN2(n8635), .QN(n6378) );
  NAND2X0 U7511 ( .IN1(n3939), .IN2(CRC_OUT_7_21), .QN(n6372) );
  NAND4X0 U7512 ( .IN1(n6379), .IN2(n6380), .IN3(n6381), .IN4(n6382), .QN(
        WX3248) );
  NAND2X0 U7513 ( .IN1(n3971), .IN2(n6129), .QN(n6382) );
  XOR3X1 U7514 ( .IN1(n3219), .IN2(n3872), .IN3(n6383), .Q(n6129) );
  XOR3X1 U7515 ( .IN1(n7205), .IN2(n3684), .IN3(WX4670), .Q(n6383) );
  NAND2X0 U7516 ( .IN1(n3892), .IN2(n6384), .QN(n6381) );
  NAND2X0 U7517 ( .IN1(n119), .IN2(n3927), .QN(n6380) );
  INVX0 U7518 ( .INP(n6385), .ZN(n119) );
  NAND2X0 U7519 ( .IN1(n4453), .IN2(n8636), .QN(n6385) );
  NAND2X0 U7520 ( .IN1(n3939), .IN2(CRC_OUT_7_22), .QN(n6379) );
  NAND4X0 U7521 ( .IN1(n6386), .IN2(n6387), .IN3(n6388), .IN4(n6389), .QN(
        WX3246) );
  NAND2X0 U7522 ( .IN1(n3974), .IN2(n6136), .QN(n6389) );
  XOR3X1 U7523 ( .IN1(n3221), .IN2(n3875), .IN3(n6390), .Q(n6136) );
  XOR3X1 U7524 ( .IN1(n7206), .IN2(n3682), .IN3(WX4668), .Q(n6390) );
  NAND2X0 U7525 ( .IN1(n6391), .IN2(n3900), .QN(n6388) );
  NAND2X0 U7526 ( .IN1(n118), .IN2(n3927), .QN(n6387) );
  INVX0 U7527 ( .INP(n6392), .ZN(n118) );
  NAND2X0 U7528 ( .IN1(n4452), .IN2(n8637), .QN(n6392) );
  NAND2X0 U7529 ( .IN1(n3945), .IN2(CRC_OUT_7_23), .QN(n6386) );
  NAND4X0 U7530 ( .IN1(n6393), .IN2(n6394), .IN3(n6395), .IN4(n6396), .QN(
        WX3244) );
  NAND2X0 U7531 ( .IN1(n3971), .IN2(n6143), .QN(n6396) );
  XOR3X1 U7532 ( .IN1(n3223), .IN2(n3874), .IN3(n6397), .Q(n6143) );
  XOR3X1 U7533 ( .IN1(n7207), .IN2(n3680), .IN3(WX4666), .Q(n6397) );
  NAND2X0 U7534 ( .IN1(n3892), .IN2(n6398), .QN(n6395) );
  NAND2X0 U7535 ( .IN1(n117), .IN2(n3927), .QN(n6394) );
  INVX0 U7536 ( .INP(n6399), .ZN(n117) );
  NAND2X0 U7537 ( .IN1(n4452), .IN2(n8638), .QN(n6399) );
  NAND2X0 U7538 ( .IN1(n3940), .IN2(CRC_OUT_7_24), .QN(n6393) );
  NAND4X0 U7539 ( .IN1(n6400), .IN2(n6401), .IN3(n6402), .IN4(n6403), .QN(
        WX3242) );
  NAND2X0 U7540 ( .IN1(n3971), .IN2(n6150), .QN(n6403) );
  XOR3X1 U7541 ( .IN1(n3225), .IN2(n3873), .IN3(n6404), .Q(n6150) );
  XOR3X1 U7542 ( .IN1(n7208), .IN2(n3678), .IN3(WX4664), .Q(n6404) );
  NAND2X0 U7543 ( .IN1(n3892), .IN2(n6405), .QN(n6402) );
  NAND2X0 U7544 ( .IN1(n116), .IN2(n3927), .QN(n6401) );
  INVX0 U7545 ( .INP(n6406), .ZN(n116) );
  NAND2X0 U7546 ( .IN1(n4452), .IN2(n8639), .QN(n6406) );
  NAND2X0 U7547 ( .IN1(n3940), .IN2(CRC_OUT_7_25), .QN(n6400) );
  NAND4X0 U7548 ( .IN1(n6407), .IN2(n6408), .IN3(n6409), .IN4(n6410), .QN(
        WX3240) );
  NAND2X0 U7549 ( .IN1(n3971), .IN2(n6157), .QN(n6410) );
  XOR3X1 U7550 ( .IN1(n3227), .IN2(n3872), .IN3(n6411), .Q(n6157) );
  XOR3X1 U7551 ( .IN1(n7209), .IN2(n3676), .IN3(WX4662), .Q(n6411) );
  NAND2X0 U7552 ( .IN1(n6412), .IN2(n3898), .QN(n6409) );
  NAND2X0 U7553 ( .IN1(n115), .IN2(n3927), .QN(n6408) );
  INVX0 U7554 ( .INP(n6413), .ZN(n115) );
  NAND2X0 U7555 ( .IN1(n4452), .IN2(n8640), .QN(n6413) );
  NAND2X0 U7556 ( .IN1(n3940), .IN2(CRC_OUT_7_26), .QN(n6407) );
  NAND4X0 U7557 ( .IN1(n6414), .IN2(n6415), .IN3(n6416), .IN4(n6417), .QN(
        WX3238) );
  NAND2X0 U7558 ( .IN1(n3972), .IN2(n6164), .QN(n6417) );
  XOR3X1 U7559 ( .IN1(n3229), .IN2(n3875), .IN3(n6418), .Q(n6164) );
  XOR3X1 U7560 ( .IN1(n7210), .IN2(n3674), .IN3(WX4660), .Q(n6418) );
  NAND2X0 U7561 ( .IN1(n3892), .IN2(n6419), .QN(n6416) );
  NAND2X0 U7562 ( .IN1(n114), .IN2(n3927), .QN(n6415) );
  INVX0 U7563 ( .INP(n6420), .ZN(n114) );
  NAND2X0 U7564 ( .IN1(n4452), .IN2(n8641), .QN(n6420) );
  NAND2X0 U7565 ( .IN1(test_so32), .IN2(n3956), .QN(n6414) );
  NAND4X0 U7566 ( .IN1(n6421), .IN2(n6422), .IN3(n6423), .IN4(n6424), .QN(
        WX3236) );
  NAND2X0 U7567 ( .IN1(n6171), .IN2(n3985), .QN(n6424) );
  XOR3X1 U7568 ( .IN1(n3231), .IN2(TM1), .IN3(n6425), .Q(n6171) );
  XOR3X1 U7569 ( .IN1(test_so40), .IN2(n7211), .IN3(WX4658), .Q(n6425) );
  NAND2X0 U7570 ( .IN1(n3892), .IN2(n6426), .QN(n6423) );
  NAND2X0 U7571 ( .IN1(n113), .IN2(n3927), .QN(n6422) );
  INVX0 U7572 ( .INP(n6427), .ZN(n113) );
  NAND2X0 U7573 ( .IN1(n4452), .IN2(n8642), .QN(n6427) );
  NAND2X0 U7574 ( .IN1(n3940), .IN2(CRC_OUT_7_28), .QN(n6421) );
  NAND4X0 U7575 ( .IN1(n6428), .IN2(n6429), .IN3(n6430), .IN4(n6431), .QN(
        WX3234) );
  NAND2X0 U7576 ( .IN1(n3972), .IN2(n6178), .QN(n6431) );
  XOR3X1 U7577 ( .IN1(n3232), .IN2(n3874), .IN3(n6432), .Q(n6178) );
  XOR3X1 U7578 ( .IN1(n7212), .IN2(n3672), .IN3(WX4656), .Q(n6432) );
  NAND2X0 U7579 ( .IN1(n3892), .IN2(n6433), .QN(n6430) );
  NAND2X0 U7580 ( .IN1(n112), .IN2(n3927), .QN(n6429) );
  INVX0 U7581 ( .INP(n6434), .ZN(n112) );
  NAND2X0 U7582 ( .IN1(n4452), .IN2(n8643), .QN(n6434) );
  NAND2X0 U7583 ( .IN1(n3940), .IN2(CRC_OUT_7_29), .QN(n6428) );
  NAND4X0 U7584 ( .IN1(n6435), .IN2(n6436), .IN3(n6437), .IN4(n6438), .QN(
        WX3232) );
  NAND2X0 U7585 ( .IN1(n6185), .IN2(n3985), .QN(n6438) );
  XOR3X1 U7586 ( .IN1(n3234), .IN2(TM1), .IN3(n6439), .Q(n6185) );
  XNOR3X1 U7587 ( .IN1(test_so38), .IN2(n7213), .IN3(n3670), .Q(n6439) );
  NAND2X0 U7588 ( .IN1(n6440), .IN2(n3897), .QN(n6437) );
  NAND2X0 U7589 ( .IN1(n111), .IN2(n3927), .QN(n6436) );
  INVX0 U7590 ( .INP(n6441), .ZN(n111) );
  NAND2X0 U7591 ( .IN1(n4452), .IN2(n8644), .QN(n6441) );
  NAND2X0 U7592 ( .IN1(n3940), .IN2(CRC_OUT_7_30), .QN(n6435) );
  NAND4X0 U7593 ( .IN1(n6442), .IN2(n6443), .IN3(n6444), .IN4(n6445), .QN(
        WX3230) );
  NAND2X0 U7594 ( .IN1(n3972), .IN2(n6192), .QN(n6445) );
  XOR3X1 U7595 ( .IN1(n3070), .IN2(n3873), .IN3(n6446), .Q(n6192) );
  XOR3X1 U7596 ( .IN1(n7214), .IN2(n3668), .IN3(WX4652), .Q(n6446) );
  NAND2X0 U7597 ( .IN1(n3892), .IN2(n6447), .QN(n6444) );
  NAND2X0 U7598 ( .IN1(n3940), .IN2(CRC_OUT_7_31), .QN(n6443) );
  NAND2X0 U7599 ( .IN1(n2245), .IN2(WX3071), .QN(n6442) );
  NOR2X0 U7600 ( .IN1(n4553), .IN2(WX3071), .QN(WX3132) );
  NOR2X0 U7601 ( .IN1(n4553), .IN2(n6448), .QN(WX2619) );
  XOR2X1 U7602 ( .IN1(n3768), .IN2(DFF_382_n1), .Q(n6448) );
  NOR2X0 U7603 ( .IN1(n4553), .IN2(n6449), .QN(WX2617) );
  XOR2X1 U7604 ( .IN1(n3770), .IN2(DFF_381_n1), .Q(n6449) );
  NOR2X0 U7605 ( .IN1(n4553), .IN2(n6450), .QN(WX2615) );
  XOR2X1 U7606 ( .IN1(n3772), .IN2(DFF_380_n1), .Q(n6450) );
  NOR2X0 U7607 ( .IN1(n4553), .IN2(n6451), .QN(WX2613) );
  XOR2X1 U7608 ( .IN1(CRC_OUT_8_27), .IN2(test_so18), .Q(n6451) );
  NOR2X0 U7609 ( .IN1(n4553), .IN2(n6452), .QN(WX2611) );
  XOR2X1 U7610 ( .IN1(n3774), .IN2(DFF_378_n1), .Q(n6452) );
  NOR2X0 U7611 ( .IN1(n4553), .IN2(n6453), .QN(WX2609) );
  XNOR2X1 U7612 ( .IN1(n3776), .IN2(test_so21), .Q(n6453) );
  NOR2X0 U7613 ( .IN1(n4553), .IN2(n6454), .QN(WX2607) );
  XOR2X1 U7614 ( .IN1(n3778), .IN2(DFF_376_n1), .Q(n6454) );
  NOR2X0 U7615 ( .IN1(n4553), .IN2(n6455), .QN(WX2605) );
  XOR2X1 U7616 ( .IN1(n3780), .IN2(DFF_375_n1), .Q(n6455) );
  NOR2X0 U7617 ( .IN1(n4553), .IN2(n6456), .QN(WX2603) );
  XOR2X1 U7618 ( .IN1(n3782), .IN2(DFF_374_n1), .Q(n6456) );
  NOR2X0 U7619 ( .IN1(n4553), .IN2(n6457), .QN(WX2601) );
  XOR2X1 U7620 ( .IN1(n3784), .IN2(DFF_373_n1), .Q(n6457) );
  NOR2X0 U7621 ( .IN1(n4553), .IN2(n6458), .QN(WX2599) );
  XOR2X1 U7622 ( .IN1(n3786), .IN2(DFF_372_n1), .Q(n6458) );
  NOR2X0 U7623 ( .IN1(n4553), .IN2(n6459), .QN(WX2597) );
  XOR2X1 U7624 ( .IN1(n3787), .IN2(DFF_371_n1), .Q(n6459) );
  NOR2X0 U7625 ( .IN1(n4553), .IN2(n6460), .QN(WX2595) );
  XOR2X1 U7626 ( .IN1(n3788), .IN2(DFF_370_n1), .Q(n6460) );
  NOR2X0 U7627 ( .IN1(n4552), .IN2(n6461), .QN(WX2593) );
  XOR2X1 U7628 ( .IN1(n3789), .IN2(DFF_369_n1), .Q(n6461) );
  NOR2X0 U7629 ( .IN1(n4552), .IN2(n6462), .QN(WX2591) );
  XOR2X1 U7630 ( .IN1(n3790), .IN2(DFF_368_n1), .Q(n6462) );
  NOR2X0 U7631 ( .IN1(n4552), .IN2(n6463), .QN(WX2589) );
  XOR3X1 U7632 ( .IN1(n3430), .IN2(DFF_383_n1), .IN3(CRC_OUT_8_15), .Q(n6463)
         );
  NOR2X0 U7633 ( .IN1(n4552), .IN2(n6464), .QN(WX2587) );
  XOR2X1 U7634 ( .IN1(n3791), .IN2(DFF_366_n1), .Q(n6464) );
  NOR2X0 U7635 ( .IN1(n4552), .IN2(n6465), .QN(WX2585) );
  XOR2X1 U7636 ( .IN1(n3792), .IN2(DFF_365_n1), .Q(n6465) );
  NOR2X0 U7637 ( .IN1(n4552), .IN2(n6466), .QN(WX2583) );
  XOR2X1 U7638 ( .IN1(n3793), .IN2(DFF_364_n1), .Q(n6466) );
  NOR2X0 U7639 ( .IN1(n4552), .IN2(n6467), .QN(WX2581) );
  XOR2X1 U7640 ( .IN1(n3794), .IN2(DFF_363_n1), .Q(n6467) );
  NOR2X0 U7641 ( .IN1(n4552), .IN2(n6468), .QN(WX2579) );
  XOR3X1 U7642 ( .IN1(n3431), .IN2(DFF_383_n1), .IN3(CRC_OUT_8_10), .Q(n6468)
         );
  NOR2X0 U7643 ( .IN1(n4552), .IN2(n6469), .QN(WX2577) );
  XOR2X1 U7644 ( .IN1(CRC_OUT_8_9), .IN2(test_so19), .Q(n6469) );
  NOR2X0 U7645 ( .IN1(n4552), .IN2(n6470), .QN(WX2575) );
  XOR2X1 U7646 ( .IN1(n3795), .IN2(DFF_360_n1), .Q(n6470) );
  NOR2X0 U7647 ( .IN1(n4552), .IN2(n6471), .QN(WX2573) );
  XNOR2X1 U7648 ( .IN1(n3796), .IN2(test_so20), .Q(n6471) );
  NOR2X0 U7649 ( .IN1(n4552), .IN2(n6472), .QN(WX2571) );
  XOR2X1 U7650 ( .IN1(n3797), .IN2(DFF_358_n1), .Q(n6472) );
  NOR2X0 U7651 ( .IN1(n4552), .IN2(n6473), .QN(WX2569) );
  XOR2X1 U7652 ( .IN1(n3798), .IN2(DFF_357_n1), .Q(n6473) );
  NOR2X0 U7653 ( .IN1(n4552), .IN2(n6474), .QN(WX2567) );
  XOR2X1 U7654 ( .IN1(n3799), .IN2(DFF_356_n1), .Q(n6474) );
  NOR2X0 U7655 ( .IN1(n4552), .IN2(n6475), .QN(WX2565) );
  XOR3X1 U7656 ( .IN1(n3432), .IN2(DFF_383_n1), .IN3(CRC_OUT_8_3), .Q(n6475)
         );
  NOR2X0 U7657 ( .IN1(n4552), .IN2(n6476), .QN(WX2563) );
  XOR2X1 U7658 ( .IN1(n3800), .IN2(DFF_354_n1), .Q(n6476) );
  NOR2X0 U7659 ( .IN1(n4551), .IN2(n6477), .QN(WX2561) );
  XOR2X1 U7660 ( .IN1(n3801), .IN2(DFF_353_n1), .Q(n6477) );
  NOR2X0 U7661 ( .IN1(n4551), .IN2(n6478), .QN(WX2559) );
  XOR2X1 U7662 ( .IN1(n3802), .IN2(DFF_352_n1), .Q(n6478) );
  NOR2X0 U7663 ( .IN1(n4551), .IN2(n6479), .QN(WX2557) );
  XOR2X1 U7664 ( .IN1(n3440), .IN2(DFF_383_n1), .Q(n6479) );
  NOR2X0 U7665 ( .IN1(n7068), .IN2(n4488), .QN(WX2031) );
  NOR2X0 U7666 ( .IN1(n7067), .IN2(n4488), .QN(WX2029) );
  NOR2X0 U7667 ( .IN1(n7066), .IN2(n4488), .QN(WX2025) );
  NOR2X0 U7668 ( .IN1(n7065), .IN2(n4488), .QN(WX2023) );
  NOR2X0 U7669 ( .IN1(n7064), .IN2(n4488), .QN(WX2021) );
  INVX0 U7670 ( .INP(n6480), .ZN(WX2019) );
  NAND2X0 U7671 ( .IN1(n4452), .IN2(test_so13), .QN(n6480) );
  NOR2X0 U7672 ( .IN1(n7063), .IN2(n4488), .QN(WX2017) );
  NOR2X0 U7673 ( .IN1(n7062), .IN2(n4488), .QN(WX2015) );
  NOR2X0 U7674 ( .IN1(n7061), .IN2(n4488), .QN(WX2013) );
  NOR2X0 U7675 ( .IN1(n7060), .IN2(n4488), .QN(WX2011) );
  NOR2X0 U7676 ( .IN1(n7059), .IN2(n4488), .QN(WX2009) );
  NOR2X0 U7677 ( .IN1(n7058), .IN2(n4488), .QN(WX2005) );
  NOR2X0 U7678 ( .IN1(n7057), .IN2(n4487), .QN(WX2003) );
  NOR2X0 U7679 ( .IN1(n7056), .IN2(n4487), .QN(WX2001) );
  NAND4X0 U7680 ( .IN1(n6481), .IN2(n6482), .IN3(n6483), .IN4(n6484), .QN(
        WX1999) );
  NAND2X0 U7681 ( .IN1(n3972), .IN2(n6230), .QN(n6484) );
  XNOR3X1 U7682 ( .IN1(n3439), .IN2(n3374), .IN3(n6485), .Q(n6230) );
  XOR2X1 U7683 ( .IN1(WX3357), .IN2(n7215), .Q(n6485) );
  NAND2X0 U7684 ( .IN1(n5494), .IN2(n3898), .QN(n6483) );
  XOR3X1 U7685 ( .IN1(n3440), .IN2(n3389), .IN3(n6486), .Q(n5494) );
  XOR2X1 U7686 ( .IN1(WX2000), .IN2(test_so16), .Q(n6486) );
  NAND2X0 U7687 ( .IN1(n63), .IN2(n3927), .QN(n6482) );
  INVX0 U7688 ( .INP(n6487), .ZN(n63) );
  NAND2X0 U7689 ( .IN1(n4451), .IN2(n8670), .QN(n6487) );
  NAND2X0 U7690 ( .IN1(n3940), .IN2(CRC_OUT_8_0), .QN(n6481) );
  NAND4X0 U7691 ( .IN1(n6488), .IN2(n6489), .IN3(n6490), .IN4(n6491), .QN(
        WX1997) );
  NAND2X0 U7692 ( .IN1(n3972), .IN2(n6237), .QN(n6491) );
  XNOR3X1 U7693 ( .IN1(n3725), .IN2(n3375), .IN3(n6492), .Q(n6237) );
  XOR2X1 U7694 ( .IN1(WX3419), .IN2(n3766), .Q(n6492) );
  NAND2X0 U7695 ( .IN1(n3892), .IN2(n5500), .QN(n6490) );
  XNOR3X1 U7696 ( .IN1(n3757), .IN2(n3390), .IN3(n6493), .Q(n5500) );
  XOR2X1 U7697 ( .IN1(WX2126), .IN2(n3802), .Q(n6493) );
  NAND2X0 U7698 ( .IN1(n62), .IN2(n3927), .QN(n6489) );
  INVX0 U7699 ( .INP(n6494), .ZN(n62) );
  NAND2X0 U7700 ( .IN1(n4451), .IN2(n8671), .QN(n6494) );
  NAND2X0 U7701 ( .IN1(n3940), .IN2(CRC_OUT_8_1), .QN(n6488) );
  NAND4X0 U7702 ( .IN1(n6495), .IN2(n6496), .IN3(n6497), .IN4(n6498), .QN(
        WX1995) );
  NAND2X0 U7703 ( .IN1(n3972), .IN2(n6244), .QN(n6498) );
  XNOR3X1 U7704 ( .IN1(n3727), .IN2(n3376), .IN3(n6499), .Q(n6244) );
  XOR2X1 U7705 ( .IN1(WX3417), .IN2(n3764), .Q(n6499) );
  NAND2X0 U7706 ( .IN1(n3892), .IN2(n5506), .QN(n6497) );
  XNOR3X1 U7707 ( .IN1(n3759), .IN2(n3391), .IN3(n6500), .Q(n5506) );
  XOR2X1 U7708 ( .IN1(WX2124), .IN2(n3801), .Q(n6500) );
  NAND2X0 U7709 ( .IN1(n61), .IN2(n3927), .QN(n6496) );
  INVX0 U7710 ( .INP(n6501), .ZN(n61) );
  NAND2X0 U7711 ( .IN1(n4451), .IN2(n8672), .QN(n6501) );
  NAND2X0 U7712 ( .IN1(n3940), .IN2(CRC_OUT_8_2), .QN(n6495) );
  NAND4X0 U7713 ( .IN1(n6502), .IN2(n6503), .IN3(n6504), .IN4(n6505), .QN(
        WX1993) );
  NAND2X0 U7714 ( .IN1(n3972), .IN2(n6251), .QN(n6505) );
  XNOR3X1 U7715 ( .IN1(n3729), .IN2(n3377), .IN3(n6506), .Q(n6251) );
  XOR2X1 U7716 ( .IN1(WX3415), .IN2(n3762), .Q(n6506) );
  NAND2X0 U7717 ( .IN1(n3892), .IN2(n5512), .QN(n6504) );
  XNOR3X1 U7718 ( .IN1(n3761), .IN2(n3392), .IN3(n6507), .Q(n5512) );
  XOR2X1 U7719 ( .IN1(WX2122), .IN2(n3800), .Q(n6507) );
  NAND2X0 U7720 ( .IN1(n60), .IN2(n3928), .QN(n6503) );
  INVX0 U7721 ( .INP(n6508), .ZN(n60) );
  NAND2X0 U7722 ( .IN1(n4451), .IN2(n8673), .QN(n6508) );
  NAND2X0 U7723 ( .IN1(n3940), .IN2(CRC_OUT_8_3), .QN(n6502) );
  NAND4X0 U7724 ( .IN1(n6509), .IN2(n6510), .IN3(n6511), .IN4(n6512), .QN(
        WX1991) );
  NAND2X0 U7725 ( .IN1(n3972), .IN2(n6258), .QN(n6512) );
  XNOR3X1 U7726 ( .IN1(n3429), .IN2(n3378), .IN3(n6513), .Q(n6258) );
  XOR2X1 U7727 ( .IN1(WX3349), .IN2(n7216), .Q(n6513) );
  NAND2X0 U7728 ( .IN1(n5518), .IN2(n3896), .QN(n6511) );
  XOR3X1 U7729 ( .IN1(n3763), .IN2(n3432), .IN3(n6514), .Q(n5518) );
  XOR2X1 U7730 ( .IN1(WX2120), .IN2(test_so14), .Q(n6514) );
  NAND2X0 U7731 ( .IN1(n59), .IN2(n3928), .QN(n6510) );
  INVX0 U7732 ( .INP(n6515), .ZN(n59) );
  NAND2X0 U7733 ( .IN1(n4451), .IN2(n8674), .QN(n6515) );
  NAND2X0 U7734 ( .IN1(n3940), .IN2(CRC_OUT_8_4), .QN(n6509) );
  NAND4X0 U7735 ( .IN1(n6516), .IN2(n6517), .IN3(n6518), .IN4(n6519), .QN(
        WX1989) );
  NAND2X0 U7736 ( .IN1(n3972), .IN2(n6265), .QN(n6519) );
  XNOR3X1 U7737 ( .IN1(n3733), .IN2(n3379), .IN3(n6520), .Q(n6265) );
  XOR2X1 U7738 ( .IN1(WX3411), .IN2(n3760), .Q(n6520) );
  NAND2X0 U7739 ( .IN1(n3892), .IN2(n5524), .QN(n6518) );
  XNOR3X1 U7740 ( .IN1(n3765), .IN2(n3393), .IN3(n6521), .Q(n5524) );
  XOR2X1 U7741 ( .IN1(WX2118), .IN2(n3799), .Q(n6521) );
  NAND2X0 U7742 ( .IN1(n58), .IN2(n3928), .QN(n6517) );
  INVX0 U7743 ( .INP(n6522), .ZN(n58) );
  NAND2X0 U7744 ( .IN1(n4451), .IN2(n8675), .QN(n6522) );
  NAND2X0 U7745 ( .IN1(n3941), .IN2(CRC_OUT_8_5), .QN(n6516) );
  NAND4X0 U7746 ( .IN1(n6523), .IN2(n6524), .IN3(n6525), .IN4(n6526), .QN(
        WX1987) );
  NAND2X0 U7747 ( .IN1(n6272), .IN2(n3985), .QN(n6526) );
  XOR3X1 U7748 ( .IN1(n3735), .IN2(n3380), .IN3(n6527), .Q(n6272) );
  XOR2X1 U7749 ( .IN1(WX3281), .IN2(test_so30), .Q(n6527) );
  NAND2X0 U7750 ( .IN1(n3892), .IN2(n5530), .QN(n6525) );
  XNOR3X1 U7751 ( .IN1(n3767), .IN2(n3394), .IN3(n6528), .Q(n5530) );
  XOR2X1 U7752 ( .IN1(WX2116), .IN2(n3798), .Q(n6528) );
  NAND2X0 U7753 ( .IN1(n57), .IN2(n3928), .QN(n6524) );
  INVX0 U7754 ( .INP(n6529), .ZN(n57) );
  NAND2X0 U7755 ( .IN1(n4451), .IN2(n8676), .QN(n6529) );
  NAND2X0 U7756 ( .IN1(n3941), .IN2(CRC_OUT_8_6), .QN(n6523) );
  NAND4X0 U7757 ( .IN1(n6530), .IN2(n6531), .IN3(n6532), .IN4(n6533), .QN(
        WX1985) );
  NAND2X0 U7758 ( .IN1(n3972), .IN2(n6279), .QN(n6533) );
  XNOR3X1 U7759 ( .IN1(n3737), .IN2(n3381), .IN3(n6534), .Q(n6279) );
  XOR2X1 U7760 ( .IN1(WX3407), .IN2(n3758), .Q(n6534) );
  NAND2X0 U7761 ( .IN1(n3891), .IN2(n5536), .QN(n6532) );
  XNOR3X1 U7762 ( .IN1(n3769), .IN2(n3395), .IN3(n6535), .Q(n5536) );
  XOR2X1 U7763 ( .IN1(WX2114), .IN2(n3797), .Q(n6535) );
  NAND2X0 U7764 ( .IN1(n56), .IN2(n3928), .QN(n6531) );
  INVX0 U7765 ( .INP(n6536), .ZN(n56) );
  NAND2X0 U7766 ( .IN1(n4451), .IN2(n8677), .QN(n6536) );
  NAND2X0 U7767 ( .IN1(test_so20), .IN2(n3957), .QN(n6530) );
  NAND4X0 U7768 ( .IN1(n6537), .IN2(n6538), .IN3(n6539), .IN4(n6540), .QN(
        WX1983) );
  NAND2X0 U7769 ( .IN1(n6286), .IN2(n3984), .QN(n6540) );
  XOR3X1 U7770 ( .IN1(n3756), .IN2(n3739), .IN3(n6541), .Q(n6286) );
  XOR2X1 U7771 ( .IN1(WX3277), .IN2(test_so28), .Q(n6541) );
  NAND2X0 U7772 ( .IN1(n3891), .IN2(n5542), .QN(n6539) );
  XNOR3X1 U7773 ( .IN1(n3771), .IN2(n3396), .IN3(n6542), .Q(n5542) );
  XOR2X1 U7774 ( .IN1(WX2112), .IN2(n3796), .Q(n6542) );
  NAND2X0 U7775 ( .IN1(n55), .IN2(n3928), .QN(n6538) );
  INVX0 U7776 ( .INP(n6543), .ZN(n55) );
  NAND2X0 U7777 ( .IN1(test_so12), .IN2(n4463), .QN(n6543) );
  NAND2X0 U7778 ( .IN1(n3941), .IN2(CRC_OUT_8_8), .QN(n6537) );
  NAND4X0 U7779 ( .IN1(n6544), .IN2(n6545), .IN3(n6546), .IN4(n6547), .QN(
        WX1981) );
  NAND2X0 U7780 ( .IN1(n3972), .IN2(n6293), .QN(n6547) );
  XNOR3X1 U7781 ( .IN1(n3741), .IN2(n3382), .IN3(n6548), .Q(n6293) );
  XOR2X1 U7782 ( .IN1(WX3403), .IN2(n3755), .Q(n6548) );
  NAND2X0 U7783 ( .IN1(n3891), .IN2(n5548), .QN(n6546) );
  XNOR3X1 U7784 ( .IN1(n3773), .IN2(n3397), .IN3(n6549), .Q(n5548) );
  XOR2X1 U7785 ( .IN1(WX2110), .IN2(n3795), .Q(n6549) );
  NAND2X0 U7786 ( .IN1(n54), .IN2(n3928), .QN(n6545) );
  INVX0 U7787 ( .INP(n6550), .ZN(n54) );
  NAND2X0 U7788 ( .IN1(n4451), .IN2(n8680), .QN(n6550) );
  NAND2X0 U7789 ( .IN1(n3941), .IN2(CRC_OUT_8_9), .QN(n6544) );
  NAND4X0 U7790 ( .IN1(n6551), .IN2(n6552), .IN3(n6553), .IN4(n6554), .QN(
        WX1979) );
  NAND2X0 U7791 ( .IN1(n3972), .IN2(n6300), .QN(n6554) );
  XNOR3X1 U7792 ( .IN1(n3743), .IN2(n3383), .IN3(n6555), .Q(n6300) );
  XOR2X1 U7793 ( .IN1(WX3401), .IN2(n3754), .Q(n6555) );
  NAND2X0 U7794 ( .IN1(n5554), .IN2(n3897), .QN(n6553) );
  XOR3X1 U7795 ( .IN1(n3775), .IN2(n3398), .IN3(n6556), .Q(n5554) );
  XOR2X1 U7796 ( .IN1(WX1980), .IN2(test_so19), .Q(n6556) );
  NAND2X0 U7797 ( .IN1(n53), .IN2(n3928), .QN(n6552) );
  INVX0 U7798 ( .INP(n6557), .ZN(n53) );
  NAND2X0 U7799 ( .IN1(n4450), .IN2(n8681), .QN(n6557) );
  NAND2X0 U7800 ( .IN1(n3941), .IN2(CRC_OUT_8_10), .QN(n6551) );
  NAND4X0 U7801 ( .IN1(n6558), .IN2(n6559), .IN3(n6560), .IN4(n6561), .QN(
        WX1977) );
  NAND2X0 U7802 ( .IN1(n3973), .IN2(n6307), .QN(n6561) );
  XNOR3X1 U7803 ( .IN1(n3428), .IN2(n3384), .IN3(n6562), .Q(n6307) );
  XOR2X1 U7804 ( .IN1(WX3335), .IN2(n7217), .Q(n6562) );
  NAND2X0 U7805 ( .IN1(n3891), .IN2(n5560), .QN(n6560) );
  XNOR3X1 U7806 ( .IN1(n3431), .IN2(n3399), .IN3(n6563), .Q(n5560) );
  XOR2X1 U7807 ( .IN1(WX2042), .IN2(n7218), .Q(n6563) );
  NAND2X0 U7808 ( .IN1(n52), .IN2(n3928), .QN(n6559) );
  INVX0 U7809 ( .INP(n6564), .ZN(n52) );
  NAND2X0 U7810 ( .IN1(n4450), .IN2(n8682), .QN(n6564) );
  NAND2X0 U7811 ( .IN1(n3941), .IN2(CRC_OUT_8_11), .QN(n6558) );
  NAND4X0 U7812 ( .IN1(n6565), .IN2(n6566), .IN3(n6567), .IN4(n6568), .QN(
        WX1975) );
  NAND2X0 U7813 ( .IN1(n6314), .IN2(n3984), .QN(n6568) );
  XOR3X1 U7814 ( .IN1(n3752), .IN2(n3385), .IN3(n6569), .Q(n6314) );
  XOR2X1 U7815 ( .IN1(WX3269), .IN2(test_so26), .Q(n6569) );
  NAND2X0 U7816 ( .IN1(n3891), .IN2(n5566), .QN(n6567) );
  XNOR3X1 U7817 ( .IN1(n3779), .IN2(n3400), .IN3(n6570), .Q(n5566) );
  XOR2X1 U7818 ( .IN1(WX2104), .IN2(n3794), .Q(n6570) );
  NAND2X0 U7819 ( .IN1(n51), .IN2(n3928), .QN(n6566) );
  INVX0 U7820 ( .INP(n6571), .ZN(n51) );
  NAND2X0 U7821 ( .IN1(n4450), .IN2(n8683), .QN(n6571) );
  NAND2X0 U7822 ( .IN1(n3941), .IN2(CRC_OUT_8_12), .QN(n6565) );
  NAND4X0 U7823 ( .IN1(n6572), .IN2(n6573), .IN3(n6574), .IN4(n6575), .QN(
        WX1973) );
  NAND2X0 U7824 ( .IN1(n3973), .IN2(n6321), .QN(n6575) );
  XNOR3X1 U7825 ( .IN1(n3749), .IN2(n3386), .IN3(n6576), .Q(n6321) );
  XOR2X1 U7826 ( .IN1(WX3395), .IN2(n3750), .Q(n6576) );
  NAND2X0 U7827 ( .IN1(n3891), .IN2(n5572), .QN(n6574) );
  XNOR3X1 U7828 ( .IN1(n3781), .IN2(n3401), .IN3(n6577), .Q(n5572) );
  XOR2X1 U7829 ( .IN1(WX2102), .IN2(n3793), .Q(n6577) );
  NAND2X0 U7830 ( .IN1(n50), .IN2(n3928), .QN(n6573) );
  INVX0 U7831 ( .INP(n6578), .ZN(n50) );
  NAND2X0 U7832 ( .IN1(n4450), .IN2(n8684), .QN(n6578) );
  NAND2X0 U7833 ( .IN1(n3941), .IN2(CRC_OUT_8_13), .QN(n6572) );
  NAND4X0 U7834 ( .IN1(n6579), .IN2(n6580), .IN3(n6581), .IN4(n6582), .QN(
        WX1971) );
  NAND2X0 U7835 ( .IN1(n3973), .IN2(n6328), .QN(n6582) );
  XNOR3X1 U7836 ( .IN1(n3748), .IN2(n3387), .IN3(n6583), .Q(n6328) );
  XOR2X1 U7837 ( .IN1(WX3329), .IN2(n7219), .Q(n6583) );
  NAND2X0 U7838 ( .IN1(n5578), .IN2(n3896), .QN(n6581) );
  XOR3X1 U7839 ( .IN1(n3792), .IN2(n3783), .IN3(n6584), .Q(n5578) );
  XOR2X1 U7840 ( .IN1(WX1972), .IN2(test_so17), .Q(n6584) );
  NAND2X0 U7841 ( .IN1(n49), .IN2(n3928), .QN(n6580) );
  INVX0 U7842 ( .INP(n6585), .ZN(n49) );
  NAND2X0 U7843 ( .IN1(n4450), .IN2(n8685), .QN(n6585) );
  NAND2X0 U7844 ( .IN1(n3941), .IN2(CRC_OUT_8_14), .QN(n6579) );
  NAND4X0 U7845 ( .IN1(n6586), .IN2(n6587), .IN3(n6588), .IN4(n6589), .QN(
        WX1969) );
  NAND2X0 U7846 ( .IN1(n3973), .IN2(n6335), .QN(n6589) );
  XNOR3X1 U7847 ( .IN1(n3747), .IN2(n3388), .IN3(n6590), .Q(n6335) );
  XOR2X1 U7848 ( .IN1(WX3327), .IN2(n7220), .Q(n6590) );
  NAND2X0 U7849 ( .IN1(n3891), .IN2(n5584), .QN(n6588) );
  XNOR3X1 U7850 ( .IN1(n3785), .IN2(n3402), .IN3(n6591), .Q(n5584) );
  XOR2X1 U7851 ( .IN1(WX2098), .IN2(n3791), .Q(n6591) );
  NAND2X0 U7852 ( .IN1(n48), .IN2(n3928), .QN(n6587) );
  INVX0 U7853 ( .INP(n6592), .ZN(n48) );
  NAND2X0 U7854 ( .IN1(n4450), .IN2(n8686), .QN(n6592) );
  NAND2X0 U7855 ( .IN1(n3941), .IN2(CRC_OUT_8_15), .QN(n6586) );
  NAND4X0 U7856 ( .IN1(n6593), .IN2(n6594), .IN3(n6595), .IN4(n6596), .QN(
        WX1967) );
  NAND2X0 U7857 ( .IN1(n6342), .IN2(n3984), .QN(n6596) );
  XOR3X1 U7858 ( .IN1(n3235), .IN2(TM1), .IN3(n6597), .Q(n6342) );
  XNOR3X1 U7859 ( .IN1(test_so24), .IN2(n7221), .IN3(n3427), .Q(n6597) );
  NAND2X0 U7860 ( .IN1(n3891), .IN2(n5590), .QN(n6595) );
  XOR3X1 U7861 ( .IN1(n3261), .IN2(n3872), .IN3(n6598), .Q(n5590) );
  XOR3X1 U7862 ( .IN1(n7068), .IN2(n3430), .IN3(WX2096), .Q(n6598) );
  NAND2X0 U7863 ( .IN1(n47), .IN2(n3928), .QN(n6594) );
  INVX0 U7864 ( .INP(n6599), .ZN(n47) );
  NAND2X0 U7865 ( .IN1(n4450), .IN2(n8687), .QN(n6599) );
  NAND2X0 U7866 ( .IN1(n3941), .IN2(CRC_OUT_8_16), .QN(n6593) );
  NAND4X0 U7867 ( .IN1(n6600), .IN2(n6601), .IN3(n6602), .IN4(n6603), .QN(
        WX1965) );
  NAND2X0 U7868 ( .IN1(n3973), .IN2(n6349), .QN(n6603) );
  XOR3X1 U7869 ( .IN1(n3236), .IN2(n3875), .IN3(n6604), .Q(n6349) );
  XOR3X1 U7870 ( .IN1(n7222), .IN2(n3746), .IN3(WX3387), .Q(n6604) );
  NAND2X0 U7871 ( .IN1(n3891), .IN2(n5596), .QN(n6602) );
  XOR3X1 U7872 ( .IN1(n3263), .IN2(n3874), .IN3(n6605), .Q(n5596) );
  XOR3X1 U7873 ( .IN1(n7067), .IN2(n3790), .IN3(WX2094), .Q(n6605) );
  NAND2X0 U7874 ( .IN1(n46), .IN2(n3928), .QN(n6601) );
  INVX0 U7875 ( .INP(n6606), .ZN(n46) );
  NAND2X0 U7876 ( .IN1(n4450), .IN2(n8688), .QN(n6606) );
  NAND2X0 U7877 ( .IN1(n3941), .IN2(CRC_OUT_8_17), .QN(n6600) );
  NAND4X0 U7878 ( .IN1(n6607), .IN2(n6608), .IN3(n6609), .IN4(n6610), .QN(
        WX1963) );
  NAND2X0 U7879 ( .IN1(n3973), .IN2(n6356), .QN(n6610) );
  XOR3X1 U7880 ( .IN1(n3238), .IN2(n3873), .IN3(n6611), .Q(n6356) );
  XOR3X1 U7881 ( .IN1(n7223), .IN2(n3744), .IN3(WX3385), .Q(n6611) );
  NAND2X0 U7882 ( .IN1(n5602), .IN2(n3897), .QN(n6609) );
  XOR3X1 U7883 ( .IN1(n3265), .IN2(TM1), .IN3(n6612), .Q(n5602) );
  XNOR3X1 U7884 ( .IN1(test_so15), .IN2(n7224), .IN3(n3789), .Q(n6612) );
  NAND2X0 U7885 ( .IN1(n45), .IN2(n3928), .QN(n6608) );
  INVX0 U7886 ( .INP(n6613), .ZN(n45) );
  NAND2X0 U7887 ( .IN1(n4450), .IN2(n8689), .QN(n6613) );
  NAND2X0 U7888 ( .IN1(n3942), .IN2(CRC_OUT_8_18), .QN(n6607) );
  NAND4X0 U7889 ( .IN1(n6614), .IN2(n6615), .IN3(n6616), .IN4(n6617), .QN(
        WX1961) );
  NAND2X0 U7890 ( .IN1(n3973), .IN2(n6363), .QN(n6617) );
  XOR3X1 U7891 ( .IN1(n3240), .IN2(n3872), .IN3(n6618), .Q(n6363) );
  XOR3X1 U7892 ( .IN1(n7225), .IN2(n3742), .IN3(WX3383), .Q(n6618) );
  NAND2X0 U7893 ( .IN1(n3891), .IN2(n5608), .QN(n6616) );
  XOR3X1 U7894 ( .IN1(n3266), .IN2(n3875), .IN3(n6619), .Q(n5608) );
  XOR3X1 U7895 ( .IN1(n7066), .IN2(n3788), .IN3(WX2090), .Q(n6619) );
  NAND2X0 U7896 ( .IN1(n44), .IN2(n3928), .QN(n6615) );
  INVX0 U7897 ( .INP(n6620), .ZN(n44) );
  NAND2X0 U7898 ( .IN1(n4449), .IN2(n8690), .QN(n6620) );
  NAND2X0 U7899 ( .IN1(n3942), .IN2(CRC_OUT_8_19), .QN(n6614) );
  NAND4X0 U7900 ( .IN1(n6621), .IN2(n6622), .IN3(n6623), .IN4(n6624), .QN(
        WX1959) );
  NAND2X0 U7901 ( .IN1(n3973), .IN2(n6370), .QN(n6624) );
  XOR3X1 U7902 ( .IN1(n3242), .IN2(n3874), .IN3(n6625), .Q(n6370) );
  XOR3X1 U7903 ( .IN1(n7226), .IN2(n3740), .IN3(WX3381), .Q(n6625) );
  NAND2X0 U7904 ( .IN1(n3891), .IN2(n5614), .QN(n6623) );
  XOR3X1 U7905 ( .IN1(n3268), .IN2(n3873), .IN3(n6626), .Q(n5614) );
  XOR3X1 U7906 ( .IN1(n7065), .IN2(n3787), .IN3(WX2088), .Q(n6626) );
  NAND2X0 U7907 ( .IN1(n43), .IN2(n3929), .QN(n6622) );
  INVX0 U7908 ( .INP(n6627), .ZN(n43) );
  NAND2X0 U7909 ( .IN1(n4449), .IN2(n8691), .QN(n6627) );
  NAND2X0 U7910 ( .IN1(n3942), .IN2(CRC_OUT_8_20), .QN(n6621) );
  NAND4X0 U7911 ( .IN1(n6628), .IN2(n6629), .IN3(n6630), .IN4(n6631), .QN(
        WX1957) );
  NAND2X0 U7912 ( .IN1(n3973), .IN2(n6377), .QN(n6631) );
  XOR3X1 U7913 ( .IN1(n3244), .IN2(n3872), .IN3(n6632), .Q(n6377) );
  XOR3X1 U7914 ( .IN1(n7227), .IN2(n3738), .IN3(WX3379), .Q(n6632) );
  NAND2X0 U7915 ( .IN1(n3891), .IN2(n5620), .QN(n6630) );
  XOR3X1 U7916 ( .IN1(n3270), .IN2(n3875), .IN3(n6633), .Q(n5620) );
  XOR3X1 U7917 ( .IN1(n7064), .IN2(n3786), .IN3(WX2086), .Q(n6633) );
  NAND2X0 U7918 ( .IN1(n42), .IN2(n3929), .QN(n6629) );
  INVX0 U7919 ( .INP(n6634), .ZN(n42) );
  NAND2X0 U7920 ( .IN1(n4449), .IN2(n8692), .QN(n6634) );
  NAND2X0 U7921 ( .IN1(n3942), .IN2(CRC_OUT_8_21), .QN(n6628) );
  NAND4X0 U7922 ( .IN1(n6635), .IN2(n6636), .IN3(n6637), .IN4(n6638), .QN(
        WX1955) );
  NAND2X0 U7923 ( .IN1(n3973), .IN2(n6384), .QN(n6638) );
  XOR3X1 U7924 ( .IN1(n3246), .IN2(n3874), .IN3(n6639), .Q(n6384) );
  XOR3X1 U7925 ( .IN1(n7228), .IN2(n3736), .IN3(WX3377), .Q(n6639) );
  NAND2X0 U7926 ( .IN1(n5626), .IN2(n3897), .QN(n6637) );
  XOR3X1 U7927 ( .IN1(n3272), .IN2(TM1), .IN3(n6640), .Q(n5626) );
  XNOR3X1 U7928 ( .IN1(test_so13), .IN2(n7229), .IN3(n3784), .Q(n6640) );
  NAND2X0 U7929 ( .IN1(n41), .IN2(n3929), .QN(n6636) );
  INVX0 U7930 ( .INP(n6641), .ZN(n41) );
  NAND2X0 U7931 ( .IN1(n4449), .IN2(n8693), .QN(n6641) );
  NAND2X0 U7932 ( .IN1(n3942), .IN2(CRC_OUT_8_22), .QN(n6635) );
  NAND4X0 U7933 ( .IN1(n6642), .IN2(n6643), .IN3(n6644), .IN4(n6645), .QN(
        WX1953) );
  NAND2X0 U7934 ( .IN1(n6391), .IN2(n3984), .QN(n6645) );
  XOR3X1 U7935 ( .IN1(n3248), .IN2(TM1), .IN3(n6646), .Q(n6391) );
  XOR3X1 U7936 ( .IN1(test_so29), .IN2(n7230), .IN3(WX3375), .Q(n6646) );
  NAND2X0 U7937 ( .IN1(n3890), .IN2(n5632), .QN(n6644) );
  XOR3X1 U7938 ( .IN1(n3273), .IN2(n3873), .IN3(n6647), .Q(n5632) );
  XOR3X1 U7939 ( .IN1(n7063), .IN2(n3782), .IN3(WX2082), .Q(n6647) );
  NAND2X0 U7940 ( .IN1(n40), .IN2(n3929), .QN(n6643) );
  INVX0 U7941 ( .INP(n6648), .ZN(n40) );
  NAND2X0 U7942 ( .IN1(n4449), .IN2(n8694), .QN(n6648) );
  NAND2X0 U7943 ( .IN1(n3942), .IN2(CRC_OUT_8_23), .QN(n6642) );
  NAND4X0 U7944 ( .IN1(n6649), .IN2(n6650), .IN3(n6651), .IN4(n6652), .QN(
        WX1951) );
  NAND2X0 U7945 ( .IN1(n3973), .IN2(n6398), .QN(n6652) );
  XOR3X1 U7946 ( .IN1(n3249), .IN2(n3872), .IN3(n6653), .Q(n6398) );
  XOR3X1 U7947 ( .IN1(n7231), .IN2(n3734), .IN3(WX3373), .Q(n6653) );
  NAND2X0 U7948 ( .IN1(n3890), .IN2(n5638), .QN(n6651) );
  XOR3X1 U7949 ( .IN1(n3275), .IN2(n3875), .IN3(n6654), .Q(n5638) );
  XOR3X1 U7950 ( .IN1(n7062), .IN2(n3780), .IN3(WX2080), .Q(n6654) );
  NAND2X0 U7951 ( .IN1(n39), .IN2(n3929), .QN(n6650) );
  INVX0 U7952 ( .INP(n6655), .ZN(n39) );
  NAND2X0 U7953 ( .IN1(n4449), .IN2(n8695), .QN(n6655) );
  NAND2X0 U7954 ( .IN1(n3942), .IN2(CRC_OUT_8_24), .QN(n6649) );
  NAND4X0 U7955 ( .IN1(n6656), .IN2(n6657), .IN3(n6658), .IN4(n6659), .QN(
        WX1949) );
  NAND2X0 U7956 ( .IN1(n3973), .IN2(n6405), .QN(n6659) );
  XOR3X1 U7957 ( .IN1(n3251), .IN2(n3874), .IN3(n6660), .Q(n6405) );
  XOR3X1 U7958 ( .IN1(n7232), .IN2(n3732), .IN3(WX3371), .Q(n6660) );
  NAND2X0 U7959 ( .IN1(n3890), .IN2(n5644), .QN(n6658) );
  XOR3X1 U7960 ( .IN1(n3277), .IN2(n3873), .IN3(n6661), .Q(n5644) );
  XOR3X1 U7961 ( .IN1(n7061), .IN2(n3778), .IN3(WX2078), .Q(n6661) );
  NAND2X0 U7962 ( .IN1(n38), .IN2(n3929), .QN(n6657) );
  INVX0 U7963 ( .INP(n6662), .ZN(n38) );
  NAND2X0 U7964 ( .IN1(n4449), .IN2(n8696), .QN(n6662) );
  NAND2X0 U7965 ( .IN1(test_so21), .IN2(n3957), .QN(n6656) );
  NAND4X0 U7966 ( .IN1(n6663), .IN2(n6664), .IN3(n6665), .IN4(n6666), .QN(
        WX1947) );
  NAND2X0 U7967 ( .IN1(n6412), .IN2(n3983), .QN(n6666) );
  XOR3X1 U7968 ( .IN1(n3253), .IN2(TM1), .IN3(n6667), .Q(n6412) );
  XNOR3X1 U7969 ( .IN1(test_so27), .IN2(n7233), .IN3(n3730), .Q(n6667) );
  NAND2X0 U7970 ( .IN1(n3890), .IN2(n5650), .QN(n6665) );
  XOR3X1 U7971 ( .IN1(n3280), .IN2(n3872), .IN3(n6668), .Q(n5650) );
  XOR3X1 U7972 ( .IN1(n7060), .IN2(n3776), .IN3(WX2076), .Q(n6668) );
  NAND2X0 U7973 ( .IN1(n37), .IN2(n3929), .QN(n6664) );
  INVX0 U7974 ( .INP(n6669), .ZN(n37) );
  NAND2X0 U7975 ( .IN1(test_so11), .IN2(n4463), .QN(n6669) );
  NAND2X0 U7976 ( .IN1(n3942), .IN2(CRC_OUT_8_26), .QN(n6663) );
  NAND4X0 U7977 ( .IN1(n6670), .IN2(n6671), .IN3(n6672), .IN4(n6673), .QN(
        WX1945) );
  NAND2X0 U7978 ( .IN1(n3974), .IN2(n6419), .QN(n6673) );
  XOR3X1 U7979 ( .IN1(n3254), .IN2(n3875), .IN3(n6674), .Q(n6419) );
  XOR3X1 U7980 ( .IN1(n7234), .IN2(n3728), .IN3(WX3367), .Q(n6674) );
  NAND2X0 U7981 ( .IN1(n3890), .IN2(n5656), .QN(n6672) );
  XOR3X1 U7982 ( .IN1(n3282), .IN2(n3874), .IN3(n6675), .Q(n5656) );
  XOR3X1 U7983 ( .IN1(n7059), .IN2(n3774), .IN3(WX2074), .Q(n6675) );
  NAND2X0 U7984 ( .IN1(n36), .IN2(n3929), .QN(n6671) );
  INVX0 U7985 ( .INP(n6676), .ZN(n36) );
  NAND2X0 U7986 ( .IN1(n4449), .IN2(n8699), .QN(n6676) );
  NAND2X0 U7987 ( .IN1(n3942), .IN2(CRC_OUT_8_27), .QN(n6670) );
  NAND4X0 U7988 ( .IN1(n6677), .IN2(n6678), .IN3(n6679), .IN4(n6680), .QN(
        WX1943) );
  NAND2X0 U7989 ( .IN1(n3974), .IN2(n6426), .QN(n6680) );
  XOR3X1 U7990 ( .IN1(n3256), .IN2(n3873), .IN3(n6681), .Q(n6426) );
  XOR3X1 U7991 ( .IN1(n7235), .IN2(n3726), .IN3(WX3365), .Q(n6681) );
  NAND2X0 U7992 ( .IN1(n5662), .IN2(n3898), .QN(n6679) );
  XOR3X1 U7993 ( .IN1(n3284), .IN2(TM1), .IN3(n6682), .Q(n5662) );
  XOR3X1 U7994 ( .IN1(test_so18), .IN2(n7236), .IN3(WX2072), .Q(n6682) );
  NAND2X0 U7995 ( .IN1(n35), .IN2(n3929), .QN(n6678) );
  INVX0 U7996 ( .INP(n6683), .ZN(n35) );
  NAND2X0 U7997 ( .IN1(n4449), .IN2(n8700), .QN(n6683) );
  NAND2X0 U7998 ( .IN1(n3942), .IN2(CRC_OUT_8_28), .QN(n6677) );
  NAND4X0 U7999 ( .IN1(n6684), .IN2(n6685), .IN3(n6686), .IN4(n6687), .QN(
        WX1941) );
  NAND2X0 U8000 ( .IN1(n3974), .IN2(n6433), .QN(n6687) );
  XOR3X1 U8001 ( .IN1(n3258), .IN2(n3872), .IN3(n6688), .Q(n6433) );
  XOR3X1 U8002 ( .IN1(n7237), .IN2(n3724), .IN3(WX3363), .Q(n6688) );
  NAND2X0 U8003 ( .IN1(n3890), .IN2(n5679), .QN(n6686) );
  XOR3X1 U8004 ( .IN1(n3285), .IN2(n3875), .IN3(n6689), .Q(n5679) );
  XOR3X1 U8005 ( .IN1(n7058), .IN2(n3772), .IN3(WX2070), .Q(n6689) );
  NAND2X0 U8006 ( .IN1(n34), .IN2(n3929), .QN(n6685) );
  INVX0 U8007 ( .INP(n6690), .ZN(n34) );
  NAND2X0 U8008 ( .IN1(n4448), .IN2(n8701), .QN(n6690) );
  NAND2X0 U8009 ( .IN1(n3942), .IN2(CRC_OUT_8_29), .QN(n6684) );
  NAND4X0 U8010 ( .IN1(n6691), .IN2(n6692), .IN3(n6693), .IN4(n6694), .QN(
        WX1939) );
  NAND2X0 U8011 ( .IN1(n6440), .IN2(n3983), .QN(n6694) );
  XOR3X1 U8012 ( .IN1(n3260), .IN2(TM1), .IN3(n6695), .Q(n6440) );
  XNOR3X1 U8013 ( .IN1(test_so25), .IN2(n7238), .IN3(n3722), .Q(n6695) );
  NAND2X0 U8014 ( .IN1(n3890), .IN2(n5695), .QN(n6693) );
  XOR3X1 U8015 ( .IN1(n3287), .IN2(n3874), .IN3(n6696), .Q(n5695) );
  XOR3X1 U8016 ( .IN1(n7057), .IN2(n3770), .IN3(WX2068), .Q(n6696) );
  NAND2X0 U8017 ( .IN1(n33), .IN2(n3929), .QN(n6692) );
  INVX0 U8018 ( .INP(n6697), .ZN(n33) );
  NAND2X0 U8019 ( .IN1(n4448), .IN2(n8702), .QN(n6697) );
  NAND2X0 U8020 ( .IN1(n3942), .IN2(CRC_OUT_8_30), .QN(n6691) );
  NAND4X0 U8021 ( .IN1(n6698), .IN2(n6699), .IN3(n6700), .IN4(n6701), .QN(
        WX1937) );
  NAND2X0 U8022 ( .IN1(n3890), .IN2(n5711), .QN(n6701) );
  XOR3X1 U8023 ( .IN1(n3074), .IN2(n3873), .IN3(n6702), .Q(n5711) );
  XOR3X1 U8024 ( .IN1(n7056), .IN2(n3768), .IN3(WX2066), .Q(n6702) );
  NAND2X0 U8025 ( .IN1(n3974), .IN2(n6447), .QN(n6700) );
  XOR3X1 U8026 ( .IN1(n3072), .IN2(n3872), .IN3(n6703), .Q(n6447) );
  XOR3X1 U8027 ( .IN1(n7239), .IN2(n3721), .IN3(WX3359), .Q(n6703) );
  NAND2X0 U8028 ( .IN1(n3943), .IN2(CRC_OUT_8_31), .QN(n6699) );
  NAND2X0 U8029 ( .IN1(n2245), .IN2(WX1778), .QN(n6698) );
  NOR2X0 U8030 ( .IN1(n4551), .IN2(WX1778), .QN(WX1839) );
  NOR2X0 U8031 ( .IN1(n4550), .IN2(n6704), .QN(WX1326) );
  XOR2X1 U8032 ( .IN1(n3855), .IN2(DFF_190_n1), .Q(n6704) );
  NOR2X0 U8033 ( .IN1(n4551), .IN2(n6705), .QN(WX1324) );
  XOR2X1 U8034 ( .IN1(n3805), .IN2(DFF_189_n1), .Q(n6705) );
  NOR2X0 U8035 ( .IN1(n4550), .IN2(n6706), .QN(WX1322) );
  XOR2X1 U8036 ( .IN1(n3810), .IN2(DFF_188_n1), .Q(n6706) );
  NOR2X0 U8037 ( .IN1(n4551), .IN2(n6707), .QN(WX1320) );
  XOR2X1 U8038 ( .IN1(n3816), .IN2(DFF_187_n1), .Q(n6707) );
  NOR2X0 U8039 ( .IN1(n4550), .IN2(n6708), .QN(WX1318) );
  XOR2X1 U8040 ( .IN1(n3819), .IN2(DFF_186_n1), .Q(n6708) );
  NOR2X0 U8041 ( .IN1(n4551), .IN2(n6709), .QN(WX1316) );
  XOR2X1 U8042 ( .IN1(n3821), .IN2(DFF_185_n1), .Q(n6709) );
  NOR2X0 U8043 ( .IN1(n4550), .IN2(n6710), .QN(WX1314) );
  XOR2X1 U8044 ( .IN1(n3826), .IN2(DFF_184_n1), .Q(n6710) );
  NOR2X0 U8045 ( .IN1(n4551), .IN2(n6711), .QN(WX1312) );
  XOR2X1 U8046 ( .IN1(n3832), .IN2(DFF_183_n1), .Q(n6711) );
  NOR2X0 U8047 ( .IN1(n4551), .IN2(n6712), .QN(WX1310) );
  XOR2X1 U8048 ( .IN1(n3833), .IN2(DFF_182_n1), .Q(n6712) );
  NOR2X0 U8049 ( .IN1(n4551), .IN2(n6713), .QN(WX1308) );
  XOR2X1 U8050 ( .IN1(n3844), .IN2(DFF_181_n1), .Q(n6713) );
  NOR2X0 U8051 ( .IN1(n4550), .IN2(n6714), .QN(WX1306) );
  XOR2X1 U8052 ( .IN1(n3850), .IN2(DFF_180_n1), .Q(n6714) );
  NOR2X0 U8053 ( .IN1(n4551), .IN2(n6715), .QN(WX1304) );
  XNOR2X1 U8054 ( .IN1(n3853), .IN2(test_so10), .Q(n6715) );
  NOR2X0 U8055 ( .IN1(n4550), .IN2(n6716), .QN(WX1302) );
  XOR2X1 U8056 ( .IN1(n3808), .IN2(DFF_178_n1), .Q(n6716) );
  NOR2X0 U8057 ( .IN1(n4551), .IN2(n6717), .QN(WX1300) );
  XOR2X1 U8058 ( .IN1(n3817), .IN2(DFF_177_n1), .Q(n6717) );
  NOR2X0 U8059 ( .IN1(n4550), .IN2(n6718), .QN(WX1298) );
  XOR2X1 U8060 ( .IN1(n3824), .IN2(DFF_176_n1), .Q(n6718) );
  NOR2X0 U8061 ( .IN1(n4551), .IN2(n6719), .QN(WX1296) );
  XOR3X1 U8062 ( .IN1(test_so8), .IN2(DFF_191_n1), .IN3(DFF_175_n1), .Q(n6719)
         );
  NOR2X0 U8063 ( .IN1(n4550), .IN2(n6720), .QN(WX1294) );
  XOR2X1 U8064 ( .IN1(n3847), .IN2(DFF_174_n1), .Q(n6720) );
  NOR2X0 U8065 ( .IN1(n4550), .IN2(n6721), .QN(WX1292) );
  XOR2X1 U8066 ( .IN1(n3856), .IN2(DFF_173_n1), .Q(n6721) );
  NOR2X0 U8067 ( .IN1(n4551), .IN2(n6722), .QN(WX1290) );
  XOR2X1 U8068 ( .IN1(n3812), .IN2(DFF_172_n1), .Q(n6722) );
  NOR2X0 U8069 ( .IN1(n4550), .IN2(n6723), .QN(WX1288) );
  XOR2X1 U8070 ( .IN1(n3828), .IN2(DFF_171_n1), .Q(n6723) );
  NOR2X0 U8071 ( .IN1(n4550), .IN2(n6724), .QN(WX1286) );
  XOR3X1 U8072 ( .IN1(n3863), .IN2(DFF_191_n1), .IN3(CRC_OUT_9_10), .Q(n6724)
         );
  NOR2X0 U8073 ( .IN1(n4551), .IN2(n6725), .QN(WX1284) );
  XOR2X1 U8074 ( .IN1(n3823), .IN2(DFF_169_n1), .Q(n6725) );
  NOR2X0 U8075 ( .IN1(n4551), .IN2(n6726), .QN(WX1282) );
  XOR2X1 U8076 ( .IN1(n3831), .IN2(DFF_168_n1), .Q(n6726) );
  NOR2X0 U8077 ( .IN1(n4554), .IN2(n6727), .QN(WX1280) );
  XOR2X1 U8078 ( .IN1(n3836), .IN2(DFF_167_n1), .Q(n6727) );
  NOR2X0 U8079 ( .IN1(n4554), .IN2(n6728), .QN(WX1278) );
  XOR2X1 U8080 ( .IN1(n3862), .IN2(DFF_166_n1), .Q(n6728) );
  NOR2X0 U8081 ( .IN1(n4554), .IN2(n6729), .QN(WX1276) );
  XOR2X1 U8082 ( .IN1(n3852), .IN2(DFF_165_n1), .Q(n6729) );
  NOR2X0 U8083 ( .IN1(n4554), .IN2(n6730), .QN(WX1274) );
  XOR2X1 U8084 ( .IN1(n3838), .IN2(DFF_164_n1), .Q(n6730) );
  NOR2X0 U8085 ( .IN1(n4554), .IN2(n6731), .QN(WX1272) );
  XOR3X1 U8086 ( .IN1(n3840), .IN2(DFF_191_n1), .IN3(CRC_OUT_9_3), .Q(n6731)
         );
  NOR2X0 U8087 ( .IN1(n4554), .IN2(n6732), .QN(WX1270) );
  XOR2X1 U8088 ( .IN1(n3806), .IN2(DFF_162_n1), .Q(n6732) );
  NOR2X0 U8089 ( .IN1(n4554), .IN2(n6733), .QN(WX1268) );
  XNOR2X1 U8090 ( .IN1(n3859), .IN2(test_so9), .Q(n6733) );
  NOR2X0 U8091 ( .IN1(n4554), .IN2(n6734), .QN(WX1266) );
  XOR2X1 U8092 ( .IN1(n3814), .IN2(DFF_160_n1), .Q(n6734) );
  NOR2X0 U8093 ( .IN1(n4554), .IN2(n6735), .QN(WX1264) );
  XOR2X1 U8094 ( .IN1(n3867), .IN2(DFF_191_n1), .Q(n6735) );
  NOR2X0 U8095 ( .IN1(n4554), .IN2(n6736), .QN(WX11670) );
  XOR2X1 U8096 ( .IN1(n3441), .IN2(DFF_1726_n1), .Q(n6736) );
  NOR2X0 U8097 ( .IN1(n4554), .IN2(n6737), .QN(WX11668) );
  XOR2X1 U8098 ( .IN1(n3442), .IN2(DFF_1725_n1), .Q(n6737) );
  NOR2X0 U8099 ( .IN1(n4554), .IN2(n6738), .QN(WX11666) );
  XOR2X1 U8100 ( .IN1(n3443), .IN2(DFF_1724_n1), .Q(n6738) );
  NOR2X0 U8101 ( .IN1(n4554), .IN2(n6739), .QN(WX11664) );
  XOR2X1 U8102 ( .IN1(n3444), .IN2(DFF_1723_n1), .Q(n6739) );
  NOR2X0 U8103 ( .IN1(n4554), .IN2(n6740), .QN(WX11662) );
  XOR2X1 U8104 ( .IN1(n3445), .IN2(DFF_1722_n1), .Q(n6740) );
  NOR2X0 U8105 ( .IN1(n4555), .IN2(n6741), .QN(WX11660) );
  XOR2X1 U8106 ( .IN1(n3446), .IN2(DFF_1721_n1), .Q(n6741) );
  NOR2X0 U8107 ( .IN1(n4555), .IN2(n6742), .QN(WX11658) );
  XOR2X1 U8108 ( .IN1(n3447), .IN2(DFF_1720_n1), .Q(n6742) );
  NOR2X0 U8109 ( .IN1(n4555), .IN2(n6743), .QN(WX11656) );
  XOR2X1 U8110 ( .IN1(n3448), .IN2(DFF_1719_n1), .Q(n6743) );
  NOR2X0 U8111 ( .IN1(n4555), .IN2(n6744), .QN(WX11654) );
  XOR2X1 U8112 ( .IN1(n3449), .IN2(DFF_1718_n1), .Q(n6744) );
  NOR2X0 U8113 ( .IN1(n4555), .IN2(n6745), .QN(WX11652) );
  XOR2X1 U8114 ( .IN1(n3450), .IN2(DFF_1717_n1), .Q(n6745) );
  NOR2X0 U8115 ( .IN1(n4555), .IN2(n6746), .QN(WX11650) );
  XOR2X1 U8116 ( .IN1(n3451), .IN2(DFF_1716_n1), .Q(n6746) );
  NOR2X0 U8117 ( .IN1(n4555), .IN2(n6747), .QN(WX11648) );
  XOR2X1 U8118 ( .IN1(n3452), .IN2(DFF_1715_n1), .Q(n6747) );
  NOR2X0 U8119 ( .IN1(n4555), .IN2(n6748), .QN(WX11646) );
  XOR2X1 U8120 ( .IN1(CRC_OUT_1_18), .IN2(test_so97), .Q(n6748) );
  NOR2X0 U8121 ( .IN1(n4555), .IN2(n6749), .QN(WX11644) );
  XOR2X1 U8122 ( .IN1(n3453), .IN2(DFF_1713_n1), .Q(n6749) );
  NOR2X0 U8123 ( .IN1(n4555), .IN2(n6750), .QN(WX11642) );
  XOR2X1 U8124 ( .IN1(n3454), .IN2(DFF_1712_n1), .Q(n6750) );
  NOR2X0 U8125 ( .IN1(n4555), .IN2(n6751), .QN(WX11640) );
  XOR3X1 U8126 ( .IN1(test_so100), .IN2(n3412), .IN3(DFF_1711_n1), .Q(n6751)
         );
  NOR2X0 U8127 ( .IN1(n4555), .IN2(n6752), .QN(WX11638) );
  XNOR2X1 U8128 ( .IN1(n3455), .IN2(test_so99), .Q(n6752) );
  NOR2X0 U8129 ( .IN1(n4555), .IN2(n6753), .QN(WX11636) );
  XOR2X1 U8130 ( .IN1(n3456), .IN2(DFF_1709_n1), .Q(n6753) );
  NOR2X0 U8131 ( .IN1(n4555), .IN2(n6754), .QN(WX11634) );
  XOR2X1 U8132 ( .IN1(n3457), .IN2(DFF_1708_n1), .Q(n6754) );
  NOR2X0 U8133 ( .IN1(n4555), .IN2(n6755), .QN(WX11632) );
  XOR2X1 U8134 ( .IN1(n3458), .IN2(DFF_1707_n1), .Q(n6755) );
  NOR2X0 U8135 ( .IN1(n4555), .IN2(n6756), .QN(WX11630) );
  XOR3X1 U8136 ( .IN1(test_so100), .IN2(n3413), .IN3(DFF_1706_n1), .Q(n6756)
         );
  NOR2X0 U8137 ( .IN1(n4556), .IN2(n6757), .QN(WX11628) );
  XOR2X1 U8138 ( .IN1(n3459), .IN2(DFF_1705_n1), .Q(n6757) );
  NOR2X0 U8139 ( .IN1(n4556), .IN2(n6758), .QN(WX11626) );
  XOR2X1 U8140 ( .IN1(n3460), .IN2(DFF_1704_n1), .Q(n6758) );
  NOR2X0 U8141 ( .IN1(n4556), .IN2(n6759), .QN(WX11624) );
  XOR2X1 U8142 ( .IN1(n3461), .IN2(DFF_1703_n1), .Q(n6759) );
  NOR2X0 U8143 ( .IN1(n4556), .IN2(n6760), .QN(WX11622) );
  XOR2X1 U8144 ( .IN1(n3462), .IN2(DFF_1702_n1), .Q(n6760) );
  NOR2X0 U8145 ( .IN1(n4556), .IN2(n6761), .QN(WX11620) );
  XOR2X1 U8146 ( .IN1(n3463), .IN2(DFF_1701_n1), .Q(n6761) );
  NOR2X0 U8147 ( .IN1(n4556), .IN2(n6762), .QN(WX11618) );
  XOR2X1 U8148 ( .IN1(n3464), .IN2(DFF_1700_n1), .Q(n6762) );
  NOR2X0 U8149 ( .IN1(n4556), .IN2(n6763), .QN(WX11616) );
  XOR3X1 U8150 ( .IN1(test_so100), .IN2(n3414), .IN3(DFF_1699_n1), .Q(n6763)
         );
  NOR2X0 U8151 ( .IN1(n4556), .IN2(n6764), .QN(WX11614) );
  XOR2X1 U8152 ( .IN1(n3465), .IN2(DFF_1698_n1), .Q(n6764) );
  NOR2X0 U8153 ( .IN1(n4556), .IN2(n6765), .QN(WX11612) );
  XOR2X1 U8154 ( .IN1(CRC_OUT_1_1), .IN2(test_so98), .Q(n6765) );
  NOR2X0 U8155 ( .IN1(n4556), .IN2(n6766), .QN(WX11610) );
  XOR2X1 U8156 ( .IN1(n3466), .IN2(DFF_1696_n1), .Q(n6766) );
  NOR2X0 U8157 ( .IN1(n4556), .IN2(n6767), .QN(WX11608) );
  XNOR2X1 U8158 ( .IN1(n3433), .IN2(test_so100), .Q(n6767) );
  NOR2X0 U8159 ( .IN1(n7080), .IN2(n4487), .QN(WX11082) );
  NOR2X0 U8160 ( .IN1(n7079), .IN2(n4487), .QN(WX11080) );
  NOR2X0 U8161 ( .IN1(n7078), .IN2(n4487), .QN(WX11078) );
  NOR2X0 U8162 ( .IN1(n7077), .IN2(n4487), .QN(WX11074) );
  NOR2X0 U8163 ( .IN1(n7076), .IN2(n4487), .QN(WX11070) );
  NOR2X0 U8164 ( .IN1(n7075), .IN2(n4487), .QN(WX11066) );
  INVX0 U8165 ( .INP(n6768), .ZN(WX11064) );
  NAND2X0 U8166 ( .IN1(n4448), .IN2(test_so91), .QN(n6768) );
  NOR2X0 U8167 ( .IN1(n7074), .IN2(n4487), .QN(WX11062) );
  NOR2X0 U8168 ( .IN1(n7073), .IN2(n4487), .QN(WX11060) );
  NOR2X0 U8169 ( .IN1(n7072), .IN2(n4487), .QN(WX11058) );
  NOR2X0 U8170 ( .IN1(n7071), .IN2(n4487), .QN(WX11056) );
  NOR2X0 U8171 ( .IN1(n7070), .IN2(n4487), .QN(WX11054) );
  NOR2X0 U8172 ( .IN1(n7069), .IN2(n4483), .QN(WX11052) );
  NAND4X0 U8173 ( .IN1(n6769), .IN2(n6770), .IN3(n6771), .IN4(n6772), .QN(
        WX11050) );
  NAND2X0 U8174 ( .IN1(n3890), .IN2(n4763), .QN(n6772) );
  XNOR3X1 U8175 ( .IN1(n3433), .IN2(n3289), .IN3(n6773), .Q(n4763) );
  XOR2X1 U8176 ( .IN1(WX11115), .IN2(n7240), .Q(n6773) );
  NAND2X0 U8177 ( .IN1(n610), .IN2(n3929), .QN(n6771) );
  INVX0 U8178 ( .INP(n6774), .ZN(n610) );
  NAND2X0 U8179 ( .IN1(n4448), .IN2(n8263), .QN(n6774) );
  NAND2X0 U8180 ( .IN1(DATA_0_0), .IN2(n3983), .QN(n6770) );
  NAND2X0 U8181 ( .IN1(n3943), .IN2(CRC_OUT_1_0), .QN(n6769) );
  NAND4X0 U8182 ( .IN1(n6775), .IN2(n6776), .IN3(n6777), .IN4(n6778), .QN(
        WX11048) );
  NAND2X0 U8183 ( .IN1(n3890), .IN2(n4770), .QN(n6778) );
  XNOR3X1 U8184 ( .IN1(n3466), .IN2(n3290), .IN3(n6779), .Q(n4770) );
  XOR2X1 U8185 ( .IN1(WX11113), .IN2(n7241), .Q(n6779) );
  NAND2X0 U8186 ( .IN1(n609), .IN2(n3929), .QN(n6777) );
  INVX0 U8187 ( .INP(n6780), .ZN(n609) );
  NAND2X0 U8188 ( .IN1(n4448), .IN2(n8264), .QN(n6780) );
  NAND2X0 U8189 ( .IN1(DATA_0_1), .IN2(n3984), .QN(n6776) );
  NAND2X0 U8190 ( .IN1(n3943), .IN2(CRC_OUT_1_1), .QN(n6775) );
  NAND4X0 U8191 ( .IN1(n6781), .IN2(n6782), .IN3(n6783), .IN4(n6784), .QN(
        WX11046) );
  NAND2X0 U8192 ( .IN1(n4777), .IN2(n3898), .QN(n6784) );
  XOR3X1 U8193 ( .IN1(n3535), .IN2(n3291), .IN3(n6785), .Q(n4777) );
  XOR2X1 U8194 ( .IN1(WX11047), .IN2(test_so98), .Q(n6785) );
  NAND2X0 U8195 ( .IN1(n608), .IN2(n3929), .QN(n6783) );
  INVX0 U8196 ( .INP(n6786), .ZN(n608) );
  NAND2X0 U8197 ( .IN1(n4448), .IN2(n8265), .QN(n6786) );
  NAND2X0 U8198 ( .IN1(DATA_0_2), .IN2(n3983), .QN(n6782) );
  NAND2X0 U8199 ( .IN1(n3943), .IN2(CRC_OUT_1_2), .QN(n6781) );
  NAND4X0 U8200 ( .IN1(n6787), .IN2(n6788), .IN3(n6789), .IN4(n6790), .QN(
        WX11044) );
  NAND2X0 U8201 ( .IN1(n3890), .IN2(n4784), .QN(n6790) );
  XNOR3X1 U8202 ( .IN1(n3465), .IN2(n3292), .IN3(n6791), .Q(n4784) );
  XOR2X1 U8203 ( .IN1(WX11109), .IN2(n7242), .Q(n6791) );
  NAND2X0 U8204 ( .IN1(n607), .IN2(n3929), .QN(n6789) );
  INVX0 U8205 ( .INP(n6792), .ZN(n607) );
  NAND2X0 U8206 ( .IN1(n4448), .IN2(n8266), .QN(n6792) );
  NAND2X0 U8207 ( .IN1(DATA_0_3), .IN2(n3982), .QN(n6788) );
  NAND2X0 U8208 ( .IN1(n3943), .IN2(CRC_OUT_1_3), .QN(n6787) );
  NAND4X0 U8209 ( .IN1(n6793), .IN2(n6794), .IN3(n6795), .IN4(n6796), .QN(
        WX11042) );
  NAND2X0 U8210 ( .IN1(n4791), .IN2(n3898), .QN(n6796) );
  XOR3X1 U8211 ( .IN1(n3539), .IN2(n3414), .IN3(n6797), .Q(n4791) );
  XOR2X1 U8212 ( .IN1(WX11043), .IN2(test_so96), .Q(n6797) );
  NAND2X0 U8213 ( .IN1(n606), .IN2(n3929), .QN(n6795) );
  INVX0 U8214 ( .INP(n6798), .ZN(n606) );
  NAND2X0 U8215 ( .IN1(n4448), .IN2(n8267), .QN(n6798) );
  NAND2X0 U8216 ( .IN1(DATA_0_4), .IN2(n3983), .QN(n6794) );
  NAND2X0 U8217 ( .IN1(n3943), .IN2(CRC_OUT_1_4), .QN(n6793) );
  NAND4X0 U8218 ( .IN1(n6799), .IN2(n6800), .IN3(n6801), .IN4(n6802), .QN(
        WX11040) );
  NAND2X0 U8219 ( .IN1(n3890), .IN2(n4798), .QN(n6802) );
  XNOR3X1 U8220 ( .IN1(n3464), .IN2(n3293), .IN3(n6803), .Q(n4798) );
  XOR2X1 U8221 ( .IN1(WX11105), .IN2(n7243), .Q(n6803) );
  NAND2X0 U8222 ( .IN1(n605), .IN2(n3929), .QN(n6801) );
  INVX0 U8223 ( .INP(n6804), .ZN(n605) );
  NAND2X0 U8224 ( .IN1(n4448), .IN2(n8268), .QN(n6804) );
  NAND2X0 U8225 ( .IN1(DATA_0_5), .IN2(n3982), .QN(n6800) );
  NAND2X0 U8226 ( .IN1(n3943), .IN2(CRC_OUT_1_5), .QN(n6799) );
  NAND4X0 U8227 ( .IN1(n6805), .IN2(n6806), .IN3(n6807), .IN4(n6808), .QN(
        WX11038) );
  NAND2X0 U8228 ( .IN1(n4805), .IN2(n3899), .QN(n6808) );
  XOR3X1 U8229 ( .IN1(n3463), .IN2(n3294), .IN3(n6809), .Q(n4805) );
  XOR2X1 U8230 ( .IN1(WX11039), .IN2(test_so94), .Q(n6809) );
  NAND2X0 U8231 ( .IN1(n604), .IN2(n3930), .QN(n6807) );
  INVX0 U8232 ( .INP(n6810), .ZN(n604) );
  NAND2X0 U8233 ( .IN1(n4447), .IN2(n8269), .QN(n6810) );
  NAND2X0 U8234 ( .IN1(DATA_0_6), .IN2(n3984), .QN(n6806) );
  NAND2X0 U8235 ( .IN1(n3943), .IN2(CRC_OUT_1_6), .QN(n6805) );
  NAND4X0 U8236 ( .IN1(n6811), .IN2(n6812), .IN3(n6813), .IN4(n6814), .QN(
        WX11036) );
  NAND2X0 U8237 ( .IN1(n3889), .IN2(n4812), .QN(n6814) );
  XNOR3X1 U8238 ( .IN1(n3462), .IN2(n3295), .IN3(n6815), .Q(n4812) );
  XOR2X1 U8239 ( .IN1(WX11101), .IN2(n7244), .Q(n6815) );
  NAND2X0 U8240 ( .IN1(n603), .IN2(n3930), .QN(n6813) );
  INVX0 U8241 ( .INP(n6816), .ZN(n603) );
  NAND2X0 U8242 ( .IN1(n4447), .IN2(n8270), .QN(n6816) );
  NAND2X0 U8243 ( .IN1(DATA_0_7), .IN2(n3984), .QN(n6812) );
  NAND2X0 U8244 ( .IN1(n3943), .IN2(CRC_OUT_1_7), .QN(n6811) );
  NAND4X0 U8245 ( .IN1(n6817), .IN2(n6818), .IN3(n6819), .IN4(n6820), .QN(
        WX11034) );
  NAND2X0 U8246 ( .IN1(n4819), .IN2(n3899), .QN(n6820) );
  XOR3X1 U8247 ( .IN1(n3547), .IN2(n3461), .IN3(n6821), .Q(n4819) );
  XOR2X1 U8248 ( .IN1(WX11163), .IN2(test_so92), .Q(n6821) );
  NAND2X0 U8249 ( .IN1(n602), .IN2(n3930), .QN(n6819) );
  INVX0 U8250 ( .INP(n6822), .ZN(n602) );
  NAND2X0 U8251 ( .IN1(n4447), .IN2(n8271), .QN(n6822) );
  NAND2X0 U8252 ( .IN1(DATA_0_8), .IN2(n3982), .QN(n6818) );
  NAND2X0 U8253 ( .IN1(n3943), .IN2(CRC_OUT_1_8), .QN(n6817) );
  NAND4X0 U8254 ( .IN1(n6823), .IN2(n6824), .IN3(n6825), .IN4(n6826), .QN(
        WX11032) );
  NAND2X0 U8255 ( .IN1(n3889), .IN2(n4826), .QN(n6826) );
  XNOR3X1 U8256 ( .IN1(n3460), .IN2(n3296), .IN3(n6827), .Q(n4826) );
  XOR2X1 U8257 ( .IN1(WX11097), .IN2(n7245), .Q(n6827) );
  NAND2X0 U8258 ( .IN1(n601), .IN2(n3930), .QN(n6825) );
  INVX0 U8259 ( .INP(n6828), .ZN(n601) );
  NAND2X0 U8260 ( .IN1(n4447), .IN2(n8272), .QN(n6828) );
  NAND2X0 U8261 ( .IN1(DATA_0_9), .IN2(n3983), .QN(n6824) );
  NAND2X0 U8262 ( .IN1(n3943), .IN2(CRC_OUT_1_9), .QN(n6823) );
  NAND4X0 U8263 ( .IN1(n6829), .IN2(n6830), .IN3(n6831), .IN4(n6832), .QN(
        WX11030) );
  NAND2X0 U8264 ( .IN1(n3889), .IN2(n4833), .QN(n6832) );
  XNOR3X1 U8265 ( .IN1(n3459), .IN2(n3297), .IN3(n6833), .Q(n4833) );
  XOR2X1 U8266 ( .IN1(WX11095), .IN2(n7246), .Q(n6833) );
  NAND2X0 U8267 ( .IN1(n600), .IN2(n3930), .QN(n6831) );
  INVX0 U8268 ( .INP(n6834), .ZN(n600) );
  NAND2X0 U8269 ( .IN1(test_so90), .IN2(n4464), .QN(n6834) );
  NAND2X0 U8270 ( .IN1(DATA_0_10), .IN2(n3983), .QN(n6830) );
  NAND2X0 U8271 ( .IN1(n3943), .IN2(CRC_OUT_1_10), .QN(n6829) );
  NAND4X0 U8272 ( .IN1(n6835), .IN2(n6836), .IN3(n6837), .IN4(n6838), .QN(
        WX11028) );
  NAND2X0 U8273 ( .IN1(n3889), .IN2(n4840), .QN(n6838) );
  XNOR3X1 U8274 ( .IN1(n3413), .IN2(n3298), .IN3(n6839), .Q(n4840) );
  XOR2X1 U8275 ( .IN1(WX11093), .IN2(n7247), .Q(n6839) );
  NAND2X0 U8276 ( .IN1(n599), .IN2(n3930), .QN(n6837) );
  INVX0 U8277 ( .INP(n6840), .ZN(n599) );
  NAND2X0 U8278 ( .IN1(n4447), .IN2(n8275), .QN(n6840) );
  NAND2X0 U8279 ( .IN1(DATA_0_11), .IN2(n3983), .QN(n6836) );
  NAND2X0 U8280 ( .IN1(n3944), .IN2(CRC_OUT_1_11), .QN(n6835) );
  NAND4X0 U8281 ( .IN1(n6841), .IN2(n6842), .IN3(n6843), .IN4(n6844), .QN(
        WX11026) );
  NAND2X0 U8282 ( .IN1(n3889), .IN2(n4847), .QN(n6844) );
  XNOR3X1 U8283 ( .IN1(n3458), .IN2(n3299), .IN3(n6845), .Q(n4847) );
  XOR2X1 U8284 ( .IN1(WX11091), .IN2(n7248), .Q(n6845) );
  NAND2X0 U8285 ( .IN1(n598), .IN2(n3930), .QN(n6843) );
  INVX0 U8286 ( .INP(n6846), .ZN(n598) );
  NAND2X0 U8287 ( .IN1(n4447), .IN2(n8276), .QN(n6846) );
  NAND2X0 U8288 ( .IN1(DATA_0_12), .IN2(n3982), .QN(n6842) );
  NAND2X0 U8289 ( .IN1(n3944), .IN2(CRC_OUT_1_12), .QN(n6841) );
  NAND4X0 U8290 ( .IN1(n6847), .IN2(n6848), .IN3(n6849), .IN4(n6850), .QN(
        WX11024) );
  NAND2X0 U8291 ( .IN1(n3889), .IN2(n4854), .QN(n6850) );
  XNOR3X1 U8292 ( .IN1(n3457), .IN2(n3300), .IN3(n6851), .Q(n4854) );
  XOR2X1 U8293 ( .IN1(WX11089), .IN2(n7249), .Q(n6851) );
  NAND2X0 U8294 ( .IN1(n597), .IN2(n3930), .QN(n6849) );
  INVX0 U8295 ( .INP(n6852), .ZN(n597) );
  NAND2X0 U8296 ( .IN1(n4447), .IN2(n8277), .QN(n6852) );
  NAND2X0 U8297 ( .IN1(DATA_0_13), .IN2(n3982), .QN(n6848) );
  NAND2X0 U8298 ( .IN1(n3944), .IN2(CRC_OUT_1_13), .QN(n6847) );
  NAND4X0 U8299 ( .IN1(n6853), .IN2(n6854), .IN3(n6855), .IN4(n6856), .QN(
        WX11022) );
  NAND2X0 U8300 ( .IN1(n3889), .IN2(n4861), .QN(n6856) );
  XNOR3X1 U8301 ( .IN1(n3456), .IN2(n3301), .IN3(n6857), .Q(n4861) );
  XOR2X1 U8302 ( .IN1(WX11087), .IN2(n7250), .Q(n6857) );
  NAND2X0 U8303 ( .IN1(n596), .IN2(n3930), .QN(n6855) );
  INVX0 U8304 ( .INP(n6858), .ZN(n596) );
  NAND2X0 U8305 ( .IN1(n4447), .IN2(n8278), .QN(n6858) );
  NAND2X0 U8306 ( .IN1(DATA_0_14), .IN2(n3982), .QN(n6854) );
  NAND2X0 U8307 ( .IN1(test_so99), .IN2(n3956), .QN(n6853) );
  NAND4X0 U8308 ( .IN1(n6859), .IN2(n6860), .IN3(n6861), .IN4(n6862), .QN(
        WX11020) );
  NAND2X0 U8309 ( .IN1(n3889), .IN2(n4868), .QN(n6862) );
  XNOR3X1 U8310 ( .IN1(n3455), .IN2(n3302), .IN3(n6863), .Q(n4868) );
  XOR2X1 U8311 ( .IN1(WX11085), .IN2(n7251), .Q(n6863) );
  NAND2X0 U8312 ( .IN1(n595), .IN2(n3930), .QN(n6861) );
  INVX0 U8313 ( .INP(n6864), .ZN(n595) );
  NAND2X0 U8314 ( .IN1(n4447), .IN2(n8279), .QN(n6864) );
  NAND2X0 U8315 ( .IN1(DATA_0_15), .IN2(n3982), .QN(n6860) );
  NAND2X0 U8316 ( .IN1(n3944), .IN2(CRC_OUT_1_15), .QN(n6859) );
  NAND4X0 U8317 ( .IN1(n6865), .IN2(n6866), .IN3(n6867), .IN4(n6868), .QN(
        WX11018) );
  NAND2X0 U8318 ( .IN1(n3889), .IN2(n4875), .QN(n6868) );
  XOR3X1 U8319 ( .IN1(n3076), .IN2(n3875), .IN3(n6869), .Q(n4875) );
  XOR3X1 U8320 ( .IN1(n7080), .IN2(n3412), .IN3(WX11147), .Q(n6869) );
  NAND2X0 U8321 ( .IN1(n594), .IN2(n3930), .QN(n6867) );
  INVX0 U8322 ( .INP(n6870), .ZN(n594) );
  NAND2X0 U8323 ( .IN1(n4446), .IN2(n8280), .QN(n6870) );
  NAND2X0 U8324 ( .IN1(DATA_0_16), .IN2(n3982), .QN(n6866) );
  NAND2X0 U8325 ( .IN1(n3944), .IN2(CRC_OUT_1_16), .QN(n6865) );
  NAND4X0 U8326 ( .IN1(n6871), .IN2(n6872), .IN3(n6873), .IN4(n6874), .QN(
        WX11016) );
  NAND2X0 U8327 ( .IN1(n3889), .IN2(n4882), .QN(n6874) );
  XOR3X1 U8328 ( .IN1(n3078), .IN2(n3874), .IN3(n6875), .Q(n4882) );
  XOR3X1 U8329 ( .IN1(n7079), .IN2(n3454), .IN3(WX11145), .Q(n6875) );
  NAND2X0 U8330 ( .IN1(n593), .IN2(n3930), .QN(n6873) );
  INVX0 U8331 ( .INP(n6876), .ZN(n593) );
  NAND2X0 U8332 ( .IN1(n4446), .IN2(n8281), .QN(n6876) );
  NAND2X0 U8333 ( .IN1(DATA_0_17), .IN2(n3982), .QN(n6872) );
  NAND2X0 U8334 ( .IN1(n3944), .IN2(CRC_OUT_1_17), .QN(n6871) );
  NAND4X0 U8335 ( .IN1(n6877), .IN2(n6878), .IN3(n6879), .IN4(n6880), .QN(
        WX11014) );
  NAND2X0 U8336 ( .IN1(n3889), .IN2(n4889), .QN(n6880) );
  XOR3X1 U8337 ( .IN1(n3080), .IN2(n3873), .IN3(n6881), .Q(n4889) );
  XOR3X1 U8338 ( .IN1(n7078), .IN2(n3453), .IN3(WX11143), .Q(n6881) );
  NAND2X0 U8339 ( .IN1(n592), .IN2(n3930), .QN(n6879) );
  INVX0 U8340 ( .INP(n6882), .ZN(n592) );
  NAND2X0 U8341 ( .IN1(n4446), .IN2(n8282), .QN(n6882) );
  NAND2X0 U8342 ( .IN1(DATA_0_18), .IN2(n3982), .QN(n6878) );
  NAND2X0 U8343 ( .IN1(n3944), .IN2(CRC_OUT_1_18), .QN(n6877) );
  NAND4X0 U8344 ( .IN1(n6883), .IN2(n6884), .IN3(n6885), .IN4(n6886), .QN(
        WX11012) );
  NAND2X0 U8345 ( .IN1(n4896), .IN2(n3900), .QN(n6886) );
  XOR3X1 U8346 ( .IN1(n3082), .IN2(TM1), .IN3(n6887), .Q(n4896) );
  XOR3X1 U8347 ( .IN1(test_so97), .IN2(n7252), .IN3(WX11141), .Q(n6887) );
  NAND2X0 U8348 ( .IN1(n591), .IN2(n3930), .QN(n6885) );
  INVX0 U8349 ( .INP(n6888), .ZN(n591) );
  NAND2X0 U8350 ( .IN1(n4446), .IN2(n8283), .QN(n6888) );
  NAND2X0 U8351 ( .IN1(DATA_0_19), .IN2(n3983), .QN(n6884) );
  NAND2X0 U8352 ( .IN1(n3944), .IN2(CRC_OUT_1_19), .QN(n6883) );
  NAND4X0 U8353 ( .IN1(n6889), .IN2(n6890), .IN3(n6891), .IN4(n6892), .QN(
        WX11010) );
  NAND2X0 U8354 ( .IN1(n3889), .IN2(n4903), .QN(n6892) );
  XOR3X1 U8355 ( .IN1(n3083), .IN2(n3872), .IN3(n6893), .Q(n4903) );
  XOR3X1 U8356 ( .IN1(n7077), .IN2(n3452), .IN3(WX11139), .Q(n6893) );
  NAND2X0 U8357 ( .IN1(n590), .IN2(n3930), .QN(n6891) );
  INVX0 U8358 ( .INP(n6894), .ZN(n590) );
  NAND2X0 U8359 ( .IN1(n4446), .IN2(n8284), .QN(n6894) );
  NAND2X0 U8360 ( .IN1(DATA_0_20), .IN2(n3982), .QN(n6890) );
  NAND2X0 U8361 ( .IN1(n3944), .IN2(CRC_OUT_1_20), .QN(n6889) );
  NAND4X0 U8362 ( .IN1(n6895), .IN2(n6896), .IN3(n6897), .IN4(n6898), .QN(
        WX11008) );
  NAND2X0 U8363 ( .IN1(n4910), .IN2(n3900), .QN(n6898) );
  XOR3X1 U8364 ( .IN1(n3085), .IN2(TM1), .IN3(n6899), .Q(n4910) );
  XNOR3X1 U8365 ( .IN1(test_so95), .IN2(n7253), .IN3(n3451), .Q(n6899) );
  NAND2X0 U8366 ( .IN1(n589), .IN2(n3930), .QN(n6897) );
  INVX0 U8367 ( .INP(n6900), .ZN(n589) );
  NAND2X0 U8368 ( .IN1(n4446), .IN2(n8285), .QN(n6900) );
  NAND2X0 U8369 ( .IN1(DATA_0_21), .IN2(n3981), .QN(n6896) );
  NAND2X0 U8370 ( .IN1(n3944), .IN2(CRC_OUT_1_21), .QN(n6895) );
  NAND4X0 U8371 ( .IN1(n6901), .IN2(n6902), .IN3(n6903), .IN4(n6904), .QN(
        WX11006) );
  NAND2X0 U8372 ( .IN1(n3888), .IN2(n4917), .QN(n6904) );
  XOR3X1 U8373 ( .IN1(n3086), .IN2(n3875), .IN3(n6905), .Q(n4917) );
  XOR3X1 U8374 ( .IN1(n7076), .IN2(n3450), .IN3(WX11135), .Q(n6905) );
  NAND2X0 U8375 ( .IN1(n588), .IN2(n3930), .QN(n6903) );
  INVX0 U8376 ( .INP(n6906), .ZN(n588) );
  NAND2X0 U8377 ( .IN1(n4446), .IN2(n8286), .QN(n6906) );
  NAND2X0 U8378 ( .IN1(DATA_0_22), .IN2(n3982), .QN(n6902) );
  NAND2X0 U8379 ( .IN1(n3944), .IN2(CRC_OUT_1_22), .QN(n6901) );
  NAND4X0 U8380 ( .IN1(n6907), .IN2(n6908), .IN3(n6909), .IN4(n6910), .QN(
        WX11004) );
  NAND2X0 U8381 ( .IN1(n4924), .IN2(n3900), .QN(n6910) );
  XOR3X1 U8382 ( .IN1(n3088), .IN2(TM1), .IN3(n6911), .Q(n4924) );
  XNOR3X1 U8383 ( .IN1(test_so93), .IN2(n7254), .IN3(n3449), .Q(n6911) );
  NAND2X0 U8384 ( .IN1(n587), .IN2(n3931), .QN(n6909) );
  INVX0 U8385 ( .INP(n6912), .ZN(n587) );
  NAND2X0 U8386 ( .IN1(n4446), .IN2(n8287), .QN(n6912) );
  NAND2X0 U8387 ( .IN1(DATA_0_23), .IN2(n3981), .QN(n6908) );
  NAND2X0 U8388 ( .IN1(n3944), .IN2(CRC_OUT_1_23), .QN(n6907) );
  NAND4X0 U8389 ( .IN1(n6913), .IN2(n6914), .IN3(n6915), .IN4(n6916), .QN(
        WX11002) );
  NAND2X0 U8390 ( .IN1(n3888), .IN2(n4931), .QN(n6916) );
  XOR3X1 U8391 ( .IN1(n3089), .IN2(n3874), .IN3(n6917), .Q(n4931) );
  XOR3X1 U8392 ( .IN1(n7075), .IN2(n3448), .IN3(WX11131), .Q(n6917) );
  NAND2X0 U8393 ( .IN1(n586), .IN2(n3931), .QN(n6915) );
  INVX0 U8394 ( .INP(n6918), .ZN(n586) );
  NAND2X0 U8395 ( .IN1(n4446), .IN2(n8288), .QN(n6918) );
  NAND2X0 U8396 ( .IN1(DATA_0_24), .IN2(n3981), .QN(n6914) );
  NAND2X0 U8397 ( .IN1(n3945), .IN2(CRC_OUT_1_24), .QN(n6913) );
  NAND4X0 U8398 ( .IN1(n6919), .IN2(n6920), .IN3(n6921), .IN4(n6922), .QN(
        WX11000) );
  NAND2X0 U8399 ( .IN1(n4938), .IN2(n3900), .QN(n6922) );
  XOR3X1 U8400 ( .IN1(n3091), .IN2(TM1), .IN3(n6923), .Q(n4938) );
  XNOR3X1 U8401 ( .IN1(test_so91), .IN2(n7255), .IN3(n3447), .Q(n6923) );
  NAND2X0 U8402 ( .IN1(n585), .IN2(n3931), .QN(n6921) );
  INVX0 U8403 ( .INP(n6924), .ZN(n585) );
  NAND2X0 U8404 ( .IN1(n4445), .IN2(n8289), .QN(n6924) );
  NAND2X0 U8405 ( .IN1(DATA_0_25), .IN2(n3982), .QN(n6920) );
  NAND2X0 U8406 ( .IN1(n3945), .IN2(CRC_OUT_1_25), .QN(n6919) );
  NAND4X0 U8407 ( .IN1(n6925), .IN2(n6926), .IN3(n6927), .IN4(n6928), .QN(
        WX10998) );
  NAND2X0 U8408 ( .IN1(n3888), .IN2(n4945), .QN(n6928) );
  XOR3X1 U8409 ( .IN1(n3092), .IN2(n3873), .IN3(n6929), .Q(n4945) );
  XOR3X1 U8410 ( .IN1(n7074), .IN2(n3446), .IN3(WX11127), .Q(n6929) );
  NAND2X0 U8411 ( .IN1(n584), .IN2(n3931), .QN(n6927) );
  INVX0 U8412 ( .INP(n6930), .ZN(n584) );
  NAND2X0 U8413 ( .IN1(n4445), .IN2(n8290), .QN(n6930) );
  NAND2X0 U8414 ( .IN1(DATA_0_26), .IN2(n3981), .QN(n6926) );
  NAND2X0 U8415 ( .IN1(n3945), .IN2(CRC_OUT_1_26), .QN(n6925) );
  NAND4X0 U8416 ( .IN1(n6931), .IN2(n6932), .IN3(n6933), .IN4(n6934), .QN(
        WX10996) );
  NAND2X0 U8417 ( .IN1(n3888), .IN2(n4952), .QN(n6934) );
  XOR3X1 U8418 ( .IN1(n3094), .IN2(n3872), .IN3(n6935), .Q(n4952) );
  XOR3X1 U8419 ( .IN1(n7073), .IN2(n3445), .IN3(WX11125), .Q(n6935) );
  NAND2X0 U8420 ( .IN1(n583), .IN2(n3931), .QN(n6933) );
  INVX0 U8421 ( .INP(n6936), .ZN(n583) );
  NAND2X0 U8422 ( .IN1(test_so89), .IN2(n4464), .QN(n6936) );
  NAND2X0 U8423 ( .IN1(DATA_0_27), .IN2(n3983), .QN(n6932) );
  NAND2X0 U8424 ( .IN1(n3945), .IN2(CRC_OUT_1_27), .QN(n6931) );
  NAND4X0 U8425 ( .IN1(n6937), .IN2(n6938), .IN3(n6939), .IN4(n6940), .QN(
        WX10994) );
  NAND2X0 U8426 ( .IN1(n3888), .IN2(n4959), .QN(n6940) );
  XOR3X1 U8427 ( .IN1(n3096), .IN2(n3875), .IN3(n6941), .Q(n4959) );
  XOR3X1 U8428 ( .IN1(n7072), .IN2(n3444), .IN3(WX11123), .Q(n6941) );
  NAND2X0 U8429 ( .IN1(n582), .IN2(n3931), .QN(n6939) );
  INVX0 U8430 ( .INP(n6942), .ZN(n582) );
  NAND2X0 U8431 ( .IN1(n4454), .IN2(n8293), .QN(n6942) );
  NAND2X0 U8432 ( .IN1(DATA_0_28), .IN2(n3981), .QN(n6938) );
  NAND2X0 U8433 ( .IN1(n3945), .IN2(CRC_OUT_1_28), .QN(n6937) );
  NAND4X0 U8434 ( .IN1(n6943), .IN2(n6944), .IN3(n6945), .IN4(n6946), .QN(
        WX10992) );
  NAND2X0 U8435 ( .IN1(n3888), .IN2(n4966), .QN(n6946) );
  XOR3X1 U8436 ( .IN1(n3098), .IN2(n3874), .IN3(n6947), .Q(n4966) );
  XOR3X1 U8437 ( .IN1(n7071), .IN2(n3443), .IN3(WX11121), .Q(n6947) );
  NAND2X0 U8438 ( .IN1(n581), .IN2(n3931), .QN(n6945) );
  INVX0 U8439 ( .INP(n6948), .ZN(n581) );
  NAND2X0 U8440 ( .IN1(n4436), .IN2(n8294), .QN(n6948) );
  NAND2X0 U8441 ( .IN1(DATA_0_29), .IN2(n3981), .QN(n6944) );
  NAND2X0 U8442 ( .IN1(n3945), .IN2(CRC_OUT_1_29), .QN(n6943) );
  NAND4X0 U8443 ( .IN1(n6949), .IN2(n6950), .IN3(n6951), .IN4(n6952), .QN(
        WX10990) );
  NAND2X0 U8444 ( .IN1(n3893), .IN2(n4973), .QN(n6952) );
  XOR3X1 U8445 ( .IN1(n3100), .IN2(n3873), .IN3(n6953), .Q(n4973) );
  XOR3X1 U8446 ( .IN1(n7070), .IN2(n3442), .IN3(WX11119), .Q(n6953) );
  NAND2X0 U8447 ( .IN1(n580), .IN2(n3931), .QN(n6951) );
  NOR2X0 U8448 ( .IN1(n3875), .IN2(n658), .QN(n2148) );
  INVX0 U8449 ( .INP(n6954), .ZN(n580) );
  NAND2X0 U8450 ( .IN1(n4445), .IN2(n8295), .QN(n6954) );
  NAND2X0 U8451 ( .IN1(DATA_0_30), .IN2(n3982), .QN(n6950) );
  NAND2X0 U8452 ( .IN1(n3945), .IN2(CRC_OUT_1_30), .QN(n6949) );
  NAND4X0 U8453 ( .IN1(n6955), .IN2(n6956), .IN3(n6957), .IN4(n6958), .QN(
        WX10988) );
  NAND2X0 U8454 ( .IN1(n3878), .IN2(n4980), .QN(n6958) );
  XOR3X1 U8455 ( .IN1(n3061), .IN2(n3872), .IN3(n6959), .Q(n4980) );
  XOR3X1 U8456 ( .IN1(n7069), .IN2(n3441), .IN3(WX11117), .Q(n6959) );
  NOR3X0 U8457 ( .IN1(n4483), .IN2(TM0), .IN3(n3875), .QN(n4761) );
  NAND2X0 U8458 ( .IN1(DATA_0_31), .IN2(n3985), .QN(n6957) );
  NAND2X0 U8459 ( .IN1(test_so100), .IN2(n3957), .QN(n6956) );
  NAND2X0 U8460 ( .IN1(n2245), .IN2(WX10829), .QN(n6955) );
  NOR2X0 U8461 ( .IN1(n4556), .IN2(WX10829), .QN(WX10890) );
  NOR2X0 U8462 ( .IN1(n4556), .IN2(n6960), .QN(WX10377) );
  XOR2X1 U8463 ( .IN1(CRC_OUT_2_30), .IN2(test_so85), .Q(n6960) );
  NOR2X0 U8464 ( .IN1(n4556), .IN2(n6961), .QN(WX10375) );
  XOR2X1 U8465 ( .IN1(n3468), .IN2(DFF_1533_n1), .Q(n6961) );
  NOR2X0 U8466 ( .IN1(n4556), .IN2(n6962), .QN(WX10373) );
  XOR2X1 U8467 ( .IN1(n3470), .IN2(DFF_1532_n1), .Q(n6962) );
  NOR2X0 U8468 ( .IN1(n4556), .IN2(n6963), .QN(WX10371) );
  XOR2X1 U8469 ( .IN1(n3472), .IN2(DFF_1531_n1), .Q(n6963) );
  NOR2X0 U8470 ( .IN1(n4557), .IN2(n6964), .QN(WX10369) );
  XOR2X1 U8471 ( .IN1(n3474), .IN2(DFF_1530_n1), .Q(n6964) );
  NOR2X0 U8472 ( .IN1(n4557), .IN2(n6965), .QN(WX10367) );
  XOR2X1 U8473 ( .IN1(n3476), .IN2(DFF_1529_n1), .Q(n6965) );
  NOR2X0 U8474 ( .IN1(n4557), .IN2(n6966), .QN(WX10365) );
  XOR2X1 U8475 ( .IN1(n3478), .IN2(DFF_1528_n1), .Q(n6966) );
  NOR2X0 U8476 ( .IN1(n4557), .IN2(n6967), .QN(WX10363) );
  XOR2X1 U8477 ( .IN1(n3480), .IN2(DFF_1527_n1), .Q(n6967) );
  NOR2X0 U8478 ( .IN1(n4557), .IN2(n6968), .QN(WX10361) );
  XOR2X1 U8479 ( .IN1(n3482), .IN2(DFF_1526_n1), .Q(n6968) );
  NOR2X0 U8480 ( .IN1(n4557), .IN2(n6969), .QN(WX10359) );
  XOR2X1 U8481 ( .IN1(n3484), .IN2(DFF_1525_n1), .Q(n6969) );
  NOR2X0 U8482 ( .IN1(n4557), .IN2(n6970), .QN(WX10357) );
  XOR2X1 U8483 ( .IN1(n3486), .IN2(DFF_1524_n1), .Q(n6970) );
  NOR2X0 U8484 ( .IN1(n4557), .IN2(n6971), .QN(WX10355) );
  XNOR2X1 U8485 ( .IN1(n3487), .IN2(test_so88), .Q(n6971) );
  NOR2X0 U8486 ( .IN1(n4557), .IN2(n6972), .QN(WX10353) );
  XOR2X1 U8487 ( .IN1(n3488), .IN2(DFF_1522_n1), .Q(n6972) );
  NOR2X0 U8488 ( .IN1(n4557), .IN2(n6973), .QN(WX10351) );
  XOR2X1 U8489 ( .IN1(n3490), .IN2(DFF_1521_n1), .Q(n6973) );
  NOR2X0 U8490 ( .IN1(n4557), .IN2(n6974), .QN(WX10349) );
  XOR2X1 U8491 ( .IN1(n3492), .IN2(DFF_1520_n1), .Q(n6974) );
  NOR2X0 U8492 ( .IN1(n4557), .IN2(n6975), .QN(WX10347) );
  XOR3X1 U8493 ( .IN1(n3415), .IN2(DFF_1535_n1), .IN3(CRC_OUT_2_15), .Q(n6975)
         );
  NOR2X0 U8494 ( .IN1(n4557), .IN2(n6976), .QN(WX10345) );
  XOR2X1 U8495 ( .IN1(n3494), .IN2(DFF_1518_n1), .Q(n6976) );
  NOR2X0 U8496 ( .IN1(n4557), .IN2(n6977), .QN(WX10343) );
  XOR2X1 U8497 ( .IN1(CRC_OUT_2_13), .IN2(test_so86), .Q(n6977) );
  NOR2X0 U8498 ( .IN1(n4557), .IN2(n6978), .QN(WX10341) );
  XOR2X1 U8499 ( .IN1(n3496), .IN2(DFF_1516_n1), .Q(n6978) );
  NOR2X0 U8500 ( .IN1(n4557), .IN2(n6979), .QN(WX10339) );
  XOR2X1 U8501 ( .IN1(n3498), .IN2(DFF_1515_n1), .Q(n6979) );
  NOR2X0 U8502 ( .IN1(n4558), .IN2(n6980), .QN(WX10337) );
  XOR3X1 U8503 ( .IN1(n3416), .IN2(DFF_1535_n1), .IN3(CRC_OUT_2_10), .Q(n6980)
         );
  NOR2X0 U8504 ( .IN1(n4558), .IN2(n6981), .QN(WX10335) );
  XOR2X1 U8505 ( .IN1(n3500), .IN2(DFF_1513_n1), .Q(n6981) );
  NOR2X0 U8506 ( .IN1(n4558), .IN2(n6982), .QN(WX10333) );
  XOR2X1 U8507 ( .IN1(n3502), .IN2(DFF_1512_n1), .Q(n6982) );
  NOR2X0 U8508 ( .IN1(n4558), .IN2(n6983), .QN(WX10331) );
  XOR2X1 U8509 ( .IN1(n3504), .IN2(DFF_1511_n1), .Q(n6983) );
  NOR2X0 U8510 ( .IN1(n4558), .IN2(n6984), .QN(WX10329) );
  XOR2X1 U8511 ( .IN1(n3506), .IN2(DFF_1510_n1), .Q(n6984) );
  NOR2X0 U8512 ( .IN1(n4558), .IN2(n6985), .QN(WX10327) );
  XOR2X1 U8513 ( .IN1(n3508), .IN2(DFF_1509_n1), .Q(n6985) );
  NOR2X0 U8514 ( .IN1(n4558), .IN2(n6986), .QN(WX10325) );
  XOR2X1 U8515 ( .IN1(n3510), .IN2(DFF_1508_n1), .Q(n6986) );
  NOR2X0 U8516 ( .IN1(n4558), .IN2(n6987), .QN(WX10323) );
  XOR3X1 U8517 ( .IN1(n3417), .IN2(DFF_1535_n1), .IN3(CRC_OUT_2_3), .Q(n6987)
         );
  NOR2X0 U8518 ( .IN1(n4558), .IN2(n6988), .QN(WX10321) );
  XNOR2X1 U8519 ( .IN1(n3512), .IN2(test_so87), .Q(n6988) );
  NOR2X0 U8520 ( .IN1(n4558), .IN2(n6989), .QN(WX10319) );
  XOR2X1 U8521 ( .IN1(n3514), .IN2(DFF_1505_n1), .Q(n6989) );
  NOR2X0 U8522 ( .IN1(n4558), .IN2(n6990), .QN(WX10317) );
  XOR2X1 U8523 ( .IN1(n3516), .IN2(DFF_1504_n1), .Q(n6990) );
  NOR2X0 U8524 ( .IN1(n4558), .IN2(n6991), .QN(WX10315) );
  XOR2X1 U8525 ( .IN1(n3434), .IN2(DFF_1535_n1), .Q(n6991) );
  XNOR2X1 U8526 ( .IN1(n6992), .IN2(n5549), .Q(DATA_9_9) );
  XNOR3X1 U8527 ( .IN1(n3485), .IN2(TM0), .IN3(n6993), .Q(n5549) );
  XOR3X1 U8528 ( .IN1(n7256), .IN2(n3831), .IN3(WX817), .Q(n6993) );
  NAND2X0 U8529 ( .IN1(TM0), .IN2(WX529), .QN(n6992) );
  XNOR2X1 U8530 ( .IN1(n6994), .IN2(n5543), .Q(DATA_9_8) );
  XNOR3X1 U8531 ( .IN1(n3483), .IN2(TM0), .IN3(n6995), .Q(n5543) );
  XNOR3X1 U8532 ( .IN1(n7257), .IN2(n3837), .IN3(n3836), .Q(n6995) );
  NAND2X0 U8533 ( .IN1(TM0), .IN2(WX531), .QN(n6994) );
  XNOR2X1 U8534 ( .IN1(n6996), .IN2(n5537), .Q(DATA_9_7) );
  XNOR3X1 U8535 ( .IN1(n3481), .IN2(TM0), .IN3(n6997), .Q(n5537) );
  XOR3X1 U8536 ( .IN1(n3862), .IN2(n3861), .IN3(WX757), .Q(n6997) );
  NAND2X0 U8537 ( .IN1(TM0), .IN2(WX533), .QN(n6996) );
  XNOR2X1 U8538 ( .IN1(n6998), .IN2(n5531), .Q(DATA_9_6) );
  XNOR3X1 U8539 ( .IN1(n3479), .IN2(n658), .IN3(n6999), .Q(n5531) );
  XOR3X1 U8540 ( .IN1(test_so5), .IN2(n3852), .IN3(WX823), .Q(n6999) );
  NAND2X0 U8541 ( .IN1(TM0), .IN2(WX535), .QN(n6998) );
  XNOR2X1 U8542 ( .IN1(n7000), .IN2(n5525), .Q(DATA_9_5) );
  XNOR3X1 U8543 ( .IN1(n3477), .IN2(TM0), .IN3(n7001), .Q(n5525) );
  XNOR3X1 U8544 ( .IN1(n7258), .IN2(n3839), .IN3(n3838), .Q(n7001) );
  NAND2X0 U8545 ( .IN1(TM0), .IN2(WX537), .QN(n7000) );
  XNOR2X1 U8546 ( .IN1(n7002), .IN2(n5519), .Q(DATA_9_4) );
  XNOR3X1 U8547 ( .IN1(n3475), .IN2(TM0), .IN3(n7003), .Q(n5519) );
  XNOR3X1 U8548 ( .IN1(n7259), .IN2(n3841), .IN3(n3840), .Q(n7003) );
  NAND2X0 U8549 ( .IN1(TM0), .IN2(WX539), .QN(n7002) );
  XNOR2X1 U8550 ( .IN1(n7004), .IN2(n5712), .Q(DATA_9_31) );
  XNOR3X1 U8551 ( .IN1(n3529), .IN2(TM1), .IN3(n7005), .Q(n5712) );
  XOR3X1 U8552 ( .IN1(n7260), .IN2(n3855), .IN3(WX773), .Q(n7005) );
  NAND2X0 U8553 ( .IN1(TM0), .IN2(WX485), .QN(n7004) );
  XNOR2X1 U8554 ( .IN1(n7006), .IN2(n5696), .Q(DATA_9_30) );
  XNOR3X1 U8555 ( .IN1(n3527), .IN2(TM1), .IN3(n7007), .Q(n5696) );
  XOR3X1 U8556 ( .IN1(n3805), .IN2(n3804), .IN3(WX711), .Q(n7007) );
  NAND2X0 U8557 ( .IN1(TM0), .IN2(WX487), .QN(n7006) );
  XNOR2X1 U8558 ( .IN1(n7008), .IN2(n5513), .Q(DATA_9_3) );
  XNOR3X1 U8559 ( .IN1(n3473), .IN2(TM0), .IN3(n7009), .Q(n5513) );
  XNOR3X1 U8560 ( .IN1(n7261), .IN2(n3807), .IN3(n3806), .Q(n7009) );
  NAND2X0 U8561 ( .IN1(TM0), .IN2(WX541), .QN(n7008) );
  XNOR2X1 U8562 ( .IN1(n7010), .IN2(n5680), .Q(DATA_9_29) );
  XNOR3X1 U8563 ( .IN1(n3525), .IN2(TM1), .IN3(n7011), .Q(n5680) );
  XNOR3X1 U8564 ( .IN1(n7262), .IN2(n3811), .IN3(n3810), .Q(n7011) );
  NAND2X0 U8565 ( .IN1(TM0), .IN2(WX489), .QN(n7010) );
  XNOR2X1 U8566 ( .IN1(n7012), .IN2(n5663), .Q(DATA_9_28) );
  XNOR3X1 U8567 ( .IN1(n3816), .IN2(n3875), .IN3(n7013), .Q(n5663) );
  XOR3X1 U8568 ( .IN1(test_so2), .IN2(n7263), .IN3(WX779), .Q(n7013) );
  NAND2X0 U8569 ( .IN1(TM0), .IN2(WX491), .QN(n7012) );
  XNOR2X1 U8570 ( .IN1(n7014), .IN2(n5657), .Q(DATA_9_27) );
  XNOR3X1 U8571 ( .IN1(n3521), .IN2(TM1), .IN3(n7015), .Q(n5657) );
  XNOR3X1 U8572 ( .IN1(n7264), .IN2(n3820), .IN3(n3819), .Q(n7015) );
  NAND2X0 U8573 ( .IN1(TM0), .IN2(WX493), .QN(n7014) );
  XNOR2X1 U8574 ( .IN1(n7016), .IN2(n5651), .Q(DATA_9_26) );
  XNOR3X1 U8575 ( .IN1(n3519), .IN2(TM1), .IN3(n7017), .Q(n5651) );
  XNOR3X1 U8576 ( .IN1(n7265), .IN2(n3822), .IN3(n3821), .Q(n7017) );
  NAND2X0 U8577 ( .IN1(TM0), .IN2(WX495), .QN(n7016) );
  XNOR2X1 U8578 ( .IN1(n7018), .IN2(n5645), .Q(DATA_9_25) );
  XNOR3X1 U8579 ( .IN1(n3517), .IN2(TM1), .IN3(n7019), .Q(n5645) );
  XNOR3X1 U8580 ( .IN1(n7266), .IN2(n3827), .IN3(n3826), .Q(n7019) );
  NAND2X0 U8581 ( .IN1(TM0), .IN2(WX497), .QN(n7018) );
  XNOR2X1 U8582 ( .IN1(n7020), .IN2(n5639), .Q(DATA_9_24) );
  XNOR3X1 U8583 ( .IN1(n3515), .IN2(n3874), .IN3(n7021), .Q(n5639) );
  XNOR3X1 U8584 ( .IN1(test_so4), .IN2(n7267), .IN3(n3832), .Q(n7021) );
  NAND2X0 U8585 ( .IN1(TM0), .IN2(WX499), .QN(n7020) );
  XNOR2X1 U8586 ( .IN1(n7022), .IN2(n5633), .Q(DATA_9_23) );
  XNOR3X1 U8587 ( .IN1(n3513), .IN2(TM1), .IN3(n7023), .Q(n5633) );
  XNOR3X1 U8588 ( .IN1(n7268), .IN2(n3834), .IN3(n3833), .Q(n7023) );
  NAND2X0 U8589 ( .IN1(TM0), .IN2(WX501), .QN(n7022) );
  XNOR2X1 U8590 ( .IN1(n7024), .IN2(n5627), .Q(DATA_9_22) );
  XNOR3X1 U8591 ( .IN1(n3511), .IN2(TM1), .IN3(n7025), .Q(n5627) );
  XOR3X1 U8592 ( .IN1(n3844), .IN2(n3843), .IN3(WX727), .Q(n7025) );
  NAND2X0 U8593 ( .IN1(TM0), .IN2(WX503), .QN(n7024) );
  XNOR2X1 U8594 ( .IN1(n7026), .IN2(n5621), .Q(DATA_9_21) );
  XNOR3X1 U8595 ( .IN1(n3509), .IN2(TM1), .IN3(n7027), .Q(n5621) );
  XOR3X1 U8596 ( .IN1(n3850), .IN2(n3849), .IN3(WX729), .Q(n7027) );
  NAND2X0 U8597 ( .IN1(TM0), .IN2(WX505), .QN(n7026) );
  XNOR2X1 U8598 ( .IN1(n7028), .IN2(n5615), .Q(DATA_9_20) );
  XNOR3X1 U8599 ( .IN1(n3507), .IN2(n3873), .IN3(n7029), .Q(n5615) );
  XNOR3X1 U8600 ( .IN1(test_so6), .IN2(n7269), .IN3(n3853), .Q(n7029) );
  NAND2X0 U8601 ( .IN1(TM0), .IN2(WX507), .QN(n7028) );
  XNOR2X1 U8602 ( .IN1(n7030), .IN2(n5507), .Q(DATA_9_2) );
  XNOR3X1 U8603 ( .IN1(n3471), .IN2(n658), .IN3(n7031), .Q(n5507) );
  XOR3X1 U8604 ( .IN1(test_so7), .IN2(n3859), .IN3(WX767), .Q(n7031) );
  NAND2X0 U8605 ( .IN1(TM0), .IN2(WX543), .QN(n7030) );
  XNOR2X1 U8606 ( .IN1(n7032), .IN2(n5609), .Q(DATA_9_19) );
  XNOR3X1 U8607 ( .IN1(n3505), .IN2(TM1), .IN3(n7033), .Q(n5609) );
  XNOR3X1 U8608 ( .IN1(n7270), .IN2(n3809), .IN3(n3808), .Q(n7033) );
  NAND2X0 U8609 ( .IN1(TM0), .IN2(WX509), .QN(n7032) );
  XNOR2X1 U8610 ( .IN1(n7034), .IN2(n5603), .Q(DATA_9_18) );
  XNOR3X1 U8611 ( .IN1(n3503), .IN2(TM1), .IN3(n7035), .Q(n5603) );
  XNOR3X1 U8612 ( .IN1(n7271), .IN2(n3818), .IN3(n3817), .Q(n7035) );
  NAND2X0 U8613 ( .IN1(TM0), .IN2(WX511), .QN(n7034) );
  XNOR2X1 U8614 ( .IN1(n7036), .IN2(n5597), .Q(DATA_9_17) );
  XNOR3X1 U8615 ( .IN1(n3501), .IN2(TM1), .IN3(n7037), .Q(n5597) );
  XNOR3X1 U8616 ( .IN1(n7272), .IN2(n3825), .IN3(n3824), .Q(n7037) );
  NAND2X0 U8617 ( .IN1(TM0), .IN2(WX513), .QN(n7036) );
  XNOR2X1 U8618 ( .IN1(n7038), .IN2(n5591), .Q(DATA_9_16) );
  XNOR3X1 U8619 ( .IN1(n3499), .IN2(n3872), .IN3(n7039), .Q(n5591) );
  XOR3X1 U8620 ( .IN1(test_so8), .IN2(n7273), .IN3(WX739), .Q(n7039) );
  NAND2X0 U8621 ( .IN1(TM0), .IN2(WX515), .QN(n7038) );
  XNOR2X1 U8622 ( .IN1(n7040), .IN2(n5585), .Q(DATA_9_15) );
  XNOR3X1 U8623 ( .IN1(n3497), .IN2(TM0), .IN3(n7041), .Q(n5585) );
  XOR3X1 U8624 ( .IN1(n3847), .IN2(n3846), .IN3(WX741), .Q(n7041) );
  NAND2X0 U8625 ( .IN1(TM0), .IN2(WX517), .QN(n7040) );
  XNOR2X1 U8626 ( .IN1(n7042), .IN2(n5579), .Q(DATA_9_14) );
  XNOR3X1 U8627 ( .IN1(n3495), .IN2(TM0), .IN3(n7043), .Q(n5579) );
  XNOR3X1 U8628 ( .IN1(n7274), .IN2(n3857), .IN3(n3856), .Q(n7043) );
  NAND2X0 U8629 ( .IN1(test_so1), .IN2(TM0), .QN(n7042) );
  XNOR2X1 U8630 ( .IN1(n7044), .IN2(n5573), .Q(DATA_9_13) );
  XNOR3X1 U8631 ( .IN1(n3493), .IN2(TM0), .IN3(n7045), .Q(n5573) );
  XNOR3X1 U8632 ( .IN1(n7275), .IN2(n3813), .IN3(n3812), .Q(n7045) );
  NAND2X0 U8633 ( .IN1(TM0), .IN2(WX521), .QN(n7044) );
  XNOR2X1 U8634 ( .IN1(n7046), .IN2(n5567), .Q(DATA_9_12) );
  XNOR3X1 U8635 ( .IN1(n3491), .IN2(TM0), .IN3(n7047), .Q(n5567) );
  XNOR3X1 U8636 ( .IN1(n7276), .IN2(n3829), .IN3(n3828), .Q(n7047) );
  NAND2X0 U8637 ( .IN1(TM0), .IN2(WX523), .QN(n7046) );
  XNOR2X1 U8638 ( .IN1(n7048), .IN2(n5561), .Q(DATA_9_11) );
  XNOR3X1 U8639 ( .IN1(n3489), .IN2(TM0), .IN3(n7049), .Q(n5561) );
  XNOR3X1 U8640 ( .IN1(n7277), .IN2(n3864), .IN3(n3863), .Q(n7049) );
  NAND2X0 U8641 ( .IN1(TM0), .IN2(WX525), .QN(n7048) );
  XNOR2X1 U8642 ( .IN1(n7050), .IN2(n5555), .Q(DATA_9_10) );
  XNOR3X1 U8643 ( .IN1(n3823), .IN2(n658), .IN3(n7051), .Q(n5555) );
  XOR3X1 U8644 ( .IN1(test_so3), .IN2(n7278), .IN3(WX815), .Q(n7051) );
  INVX0 U8645 ( .INP(TM0), .ZN(n658) );
  NAND2X0 U8646 ( .IN1(TM0), .IN2(WX527), .QN(n7050) );
  XNOR2X1 U8647 ( .IN1(n7052), .IN2(n5501), .Q(DATA_9_1) );
  XNOR3X1 U8648 ( .IN1(n3469), .IN2(TM0), .IN3(n7053), .Q(n5501) );
  XNOR3X1 U8649 ( .IN1(n7279), .IN2(n3815), .IN3(n3814), .Q(n7053) );
  NAND2X0 U8650 ( .IN1(TM0), .IN2(WX545), .QN(n7052) );
  XNOR2X1 U8651 ( .IN1(n7054), .IN2(n5495), .Q(DATA_9_0) );
  XNOR3X1 U8652 ( .IN1(n3467), .IN2(TM0), .IN3(n7055), .Q(n5495) );
  XOR3X1 U8653 ( .IN1(n3867), .IN2(n3866), .IN3(WX771), .Q(n7055) );
  NAND2X0 U8654 ( .IN1(TM0), .IN2(WX547), .QN(n7054) );
  NOR2X0 U3558_U2 ( .IN1(n4497), .IN2(U3558_n1), .QN(n2245) );
  INVX0 U3558_U1 ( .INP(n3915), .ZN(U3558_n1) );
  INVX0 U3871_U2 ( .INP(n3278), .ZN(U3871_n1) );
  NOR2X0 U3871_U1 ( .IN1(TM0), .IN2(U3871_n1), .QN(n2153) );
  INVX0 U3991_U2 ( .INP(n3278), .ZN(U3991_n1) );
  NOR2X0 U3991_U1 ( .IN1(n658), .IN2(U3991_n1), .QN(n2152) );
  INVX0 U5716_U2 ( .INP(WX547), .ZN(U5716_n1) );
  NOR2X0 U5716_U1 ( .IN1(n4541), .IN2(U5716_n1), .QN(WX544) );
  INVX0 U5717_U2 ( .INP(WX545), .ZN(U5717_n1) );
  NOR2X0 U5717_U1 ( .IN1(n4516), .IN2(U5717_n1), .QN(WX542) );
  INVX0 U5718_U2 ( .INP(WX543), .ZN(U5718_n1) );
  NOR2X0 U5718_U1 ( .IN1(n4528), .IN2(U5718_n1), .QN(WX540) );
  INVX0 U5719_U2 ( .INP(WX541), .ZN(U5719_n1) );
  NOR2X0 U5719_U1 ( .IN1(n4524), .IN2(U5719_n1), .QN(WX538) );
  INVX0 U5720_U2 ( .INP(WX539), .ZN(U5720_n1) );
  NOR2X0 U5720_U1 ( .IN1(n4524), .IN2(U5720_n1), .QN(WX536) );
  INVX0 U5721_U2 ( .INP(WX537), .ZN(U5721_n1) );
  NOR2X0 U5721_U1 ( .IN1(n4524), .IN2(U5721_n1), .QN(WX534) );
  INVX0 U5722_U2 ( .INP(WX535), .ZN(U5722_n1) );
  NOR2X0 U5722_U1 ( .IN1(n4524), .IN2(U5722_n1), .QN(WX532) );
  INVX0 U5723_U2 ( .INP(WX533), .ZN(U5723_n1) );
  NOR2X0 U5723_U1 ( .IN1(n4524), .IN2(U5723_n1), .QN(WX530) );
  INVX0 U5724_U2 ( .INP(WX531), .ZN(U5724_n1) );
  NOR2X0 U5724_U1 ( .IN1(n4525), .IN2(U5724_n1), .QN(WX528) );
  INVX0 U5725_U2 ( .INP(WX529), .ZN(U5725_n1) );
  NOR2X0 U5725_U1 ( .IN1(n4525), .IN2(U5725_n1), .QN(WX526) );
  INVX0 U5726_U2 ( .INP(WX527), .ZN(U5726_n1) );
  NOR2X0 U5726_U1 ( .IN1(n4525), .IN2(U5726_n1), .QN(WX524) );
  INVX0 U5727_U2 ( .INP(WX525), .ZN(U5727_n1) );
  NOR2X0 U5727_U1 ( .IN1(n4525), .IN2(U5727_n1), .QN(WX522) );
  INVX0 U5728_U2 ( .INP(WX523), .ZN(U5728_n1) );
  NOR2X0 U5728_U1 ( .IN1(n4525), .IN2(U5728_n1), .QN(WX520) );
  INVX0 U5729_U2 ( .INP(WX521), .ZN(U5729_n1) );
  NOR2X0 U5729_U1 ( .IN1(n4525), .IN2(U5729_n1), .QN(WX518) );
  INVX0 U5730_U2 ( .INP(test_so1), .ZN(U5730_n1) );
  NOR2X0 U5730_U1 ( .IN1(n4525), .IN2(U5730_n1), .QN(WX516) );
  INVX0 U5731_U2 ( .INP(WX517), .ZN(U5731_n1) );
  NOR2X0 U5731_U1 ( .IN1(n4525), .IN2(U5731_n1), .QN(WX514) );
  INVX0 U5732_U2 ( .INP(WX515), .ZN(U5732_n1) );
  NOR2X0 U5732_U1 ( .IN1(n4525), .IN2(U5732_n1), .QN(WX512) );
  INVX0 U5733_U2 ( .INP(WX513), .ZN(U5733_n1) );
  NOR2X0 U5733_U1 ( .IN1(n4525), .IN2(U5733_n1), .QN(WX510) );
  INVX0 U5734_U2 ( .INP(WX511), .ZN(U5734_n1) );
  NOR2X0 U5734_U1 ( .IN1(n4525), .IN2(U5734_n1), .QN(WX508) );
  INVX0 U5735_U2 ( .INP(WX509), .ZN(U5735_n1) );
  NOR2X0 U5735_U1 ( .IN1(n4525), .IN2(U5735_n1), .QN(WX506) );
  INVX0 U5736_U2 ( .INP(WX507), .ZN(U5736_n1) );
  NOR2X0 U5736_U1 ( .IN1(n4525), .IN2(U5736_n1), .QN(WX504) );
  INVX0 U5737_U2 ( .INP(WX505), .ZN(U5737_n1) );
  NOR2X0 U5737_U1 ( .IN1(n4526), .IN2(U5737_n1), .QN(WX502) );
  INVX0 U5738_U2 ( .INP(WX503), .ZN(U5738_n1) );
  NOR2X0 U5738_U1 ( .IN1(n4526), .IN2(U5738_n1), .QN(WX500) );
  INVX0 U5739_U2 ( .INP(WX501), .ZN(U5739_n1) );
  NOR2X0 U5739_U1 ( .IN1(n4526), .IN2(U5739_n1), .QN(WX498) );
  INVX0 U5740_U2 ( .INP(WX499), .ZN(U5740_n1) );
  NOR2X0 U5740_U1 ( .IN1(n4526), .IN2(U5740_n1), .QN(WX496) );
  INVX0 U5741_U2 ( .INP(WX497), .ZN(U5741_n1) );
  NOR2X0 U5741_U1 ( .IN1(n4526), .IN2(U5741_n1), .QN(WX494) );
  INVX0 U5742_U2 ( .INP(WX495), .ZN(U5742_n1) );
  NOR2X0 U5742_U1 ( .IN1(n4526), .IN2(U5742_n1), .QN(WX492) );
  INVX0 U5743_U2 ( .INP(WX493), .ZN(U5743_n1) );
  NOR2X0 U5743_U1 ( .IN1(n4526), .IN2(U5743_n1), .QN(WX490) );
  INVX0 U5744_U2 ( .INP(WX491), .ZN(U5744_n1) );
  NOR2X0 U5744_U1 ( .IN1(n4526), .IN2(U5744_n1), .QN(WX488) );
  INVX0 U5745_U2 ( .INP(WX489), .ZN(U5745_n1) );
  NOR2X0 U5745_U1 ( .IN1(n4526), .IN2(U5745_n1), .QN(WX486) );
  INVX0 U5746_U2 ( .INP(WX487), .ZN(U5746_n1) );
  NOR2X0 U5746_U1 ( .IN1(n4526), .IN2(U5746_n1), .QN(WX484) );
  INVX0 U5747_U2 ( .INP(WX5939), .ZN(U5747_n1) );
  NOR2X0 U5747_U1 ( .IN1(n4526), .IN2(U5747_n1), .QN(WX6002) );
  INVX0 U5748_U2 ( .INP(test_so49), .ZN(U5748_n1) );
  NOR2X0 U5748_U1 ( .IN1(n4526), .IN2(U5748_n1), .QN(WX6000) );
  INVX0 U5749_U2 ( .INP(WX5935), .ZN(U5749_n1) );
  NOR2X0 U5749_U1 ( .IN1(n4526), .IN2(U5749_n1), .QN(WX5998) );
  INVX0 U5750_U2 ( .INP(WX5933), .ZN(U5750_n1) );
  NOR2X0 U5750_U1 ( .IN1(n4527), .IN2(U5750_n1), .QN(WX5996) );
  INVX0 U5751_U2 ( .INP(WX5931), .ZN(U5751_n1) );
  NOR2X0 U5751_U1 ( .IN1(n4527), .IN2(U5751_n1), .QN(WX5994) );
  INVX0 U5752_U2 ( .INP(WX3269), .ZN(U5752_n1) );
  NOR2X0 U5752_U1 ( .IN1(n4527), .IN2(U5752_n1), .QN(WX3332) );
  INVX0 U5753_U2 ( .INP(WX3265), .ZN(U5753_n1) );
  NOR2X0 U5753_U1 ( .IN1(n4527), .IN2(U5753_n1), .QN(WX3328) );
  INVX0 U5754_U2 ( .INP(WX3263), .ZN(U5754_n1) );
  NOR2X0 U5754_U1 ( .IN1(n4527), .IN2(U5754_n1), .QN(WX3326) );
  INVX0 U5755_U2 ( .INP(WX11179), .ZN(U5755_n1) );
  NOR2X0 U5755_U1 ( .IN1(n4527), .IN2(U5755_n1), .QN(WX11242) );
  INVX0 U5756_U2 ( .INP(WX11177), .ZN(U5756_n1) );
  NOR2X0 U5756_U1 ( .IN1(n4527), .IN2(U5756_n1), .QN(WX11240) );
  INVX0 U5757_U2 ( .INP(WX11175), .ZN(U5757_n1) );
  NOR2X0 U5757_U1 ( .IN1(n4527), .IN2(U5757_n1), .QN(WX11238) );
  INVX0 U5758_U2 ( .INP(WX11173), .ZN(U5758_n1) );
  NOR2X0 U5758_U1 ( .IN1(n4527), .IN2(U5758_n1), .QN(WX11236) );
  INVX0 U5759_U2 ( .INP(test_so96), .ZN(U5759_n1) );
  NOR2X0 U5759_U1 ( .IN1(n4527), .IN2(U5759_n1), .QN(WX11234) );
  INVX0 U5760_U2 ( .INP(WX11169), .ZN(U5760_n1) );
  NOR2X0 U5760_U1 ( .IN1(n4527), .IN2(U5760_n1), .QN(WX11232) );
  INVX0 U5761_U2 ( .INP(WX11167), .ZN(U5761_n1) );
  NOR2X0 U5761_U1 ( .IN1(n4527), .IN2(U5761_n1), .QN(WX11230) );
  INVX0 U5762_U2 ( .INP(WX11165), .ZN(U5762_n1) );
  NOR2X0 U5762_U1 ( .IN1(n4527), .IN2(U5762_n1), .QN(WX11228) );
  INVX0 U5763_U2 ( .INP(WX11163), .ZN(U5763_n1) );
  NOR2X0 U5763_U1 ( .IN1(n4528), .IN2(U5763_n1), .QN(WX11226) );
  INVX0 U5764_U2 ( .INP(WX11161), .ZN(U5764_n1) );
  NOR2X0 U5764_U1 ( .IN1(n4528), .IN2(U5764_n1), .QN(WX11224) );
  INVX0 U5765_U2 ( .INP(WX11159), .ZN(U5765_n1) );
  NOR2X0 U5765_U1 ( .IN1(n4528), .IN2(U5765_n1), .QN(WX11222) );
  INVX0 U5766_U2 ( .INP(WX11157), .ZN(U5766_n1) );
  NOR2X0 U5766_U1 ( .IN1(n4528), .IN2(U5766_n1), .QN(WX11220) );
  INVX0 U5767_U2 ( .INP(WX11155), .ZN(U5767_n1) );
  NOR2X0 U5767_U1 ( .IN1(n4528), .IN2(U5767_n1), .QN(WX11218) );
  INVX0 U5768_U2 ( .INP(WX11153), .ZN(U5768_n1) );
  NOR2X0 U5768_U1 ( .IN1(n4528), .IN2(U5768_n1), .QN(WX11216) );
  INVX0 U5769_U2 ( .INP(WX11151), .ZN(U5769_n1) );
  NOR2X0 U5769_U1 ( .IN1(n4528), .IN2(U5769_n1), .QN(WX11214) );
  INVX0 U5770_U2 ( .INP(WX11149), .ZN(U5770_n1) );
  NOR2X0 U5770_U1 ( .IN1(n4528), .IN2(U5770_n1), .QN(WX11212) );
  INVX0 U5771_U2 ( .INP(WX11147), .ZN(U5771_n1) );
  NOR2X0 U5771_U1 ( .IN1(n4528), .IN2(U5771_n1), .QN(WX11210) );
  INVX0 U5772_U2 ( .INP(WX11145), .ZN(U5772_n1) );
  NOR2X0 U5772_U1 ( .IN1(n4528), .IN2(U5772_n1), .QN(WX11208) );
  INVX0 U5773_U2 ( .INP(WX11143), .ZN(U5773_n1) );
  NOR2X0 U5773_U1 ( .IN1(n4528), .IN2(U5773_n1), .QN(WX11206) );
  INVX0 U5774_U2 ( .INP(WX11141), .ZN(U5774_n1) );
  NOR2X0 U5774_U1 ( .IN1(n4528), .IN2(U5774_n1), .QN(WX11204) );
  INVX0 U5775_U2 ( .INP(WX11139), .ZN(U5775_n1) );
  NOR2X0 U5775_U1 ( .IN1(n4529), .IN2(U5775_n1), .QN(WX11202) );
  INVX0 U5776_U2 ( .INP(test_so95), .ZN(U5776_n1) );
  NOR2X0 U5776_U1 ( .IN1(n4529), .IN2(U5776_n1), .QN(WX11200) );
  INVX0 U5777_U2 ( .INP(WX11135), .ZN(U5777_n1) );
  NOR2X0 U5777_U1 ( .IN1(n4529), .IN2(U5777_n1), .QN(WX11198) );
  INVX0 U5778_U2 ( .INP(WX11133), .ZN(U5778_n1) );
  NOR2X0 U5778_U1 ( .IN1(n4529), .IN2(U5778_n1), .QN(WX11196) );
  INVX0 U5779_U2 ( .INP(WX11131), .ZN(U5779_n1) );
  NOR2X0 U5779_U1 ( .IN1(n4529), .IN2(U5779_n1), .QN(WX11194) );
  INVX0 U5780_U2 ( .INP(WX11129), .ZN(U5780_n1) );
  NOR2X0 U5780_U1 ( .IN1(n4529), .IN2(U5780_n1), .QN(WX11192) );
  INVX0 U5781_U2 ( .INP(WX11127), .ZN(U5781_n1) );
  NOR2X0 U5781_U1 ( .IN1(n4529), .IN2(U5781_n1), .QN(WX11190) );
  INVX0 U5782_U2 ( .INP(WX11125), .ZN(U5782_n1) );
  NOR2X0 U5782_U1 ( .IN1(n4529), .IN2(U5782_n1), .QN(WX11188) );
  INVX0 U5783_U2 ( .INP(WX11123), .ZN(U5783_n1) );
  NOR2X0 U5783_U1 ( .IN1(n4529), .IN2(U5783_n1), .QN(WX11186) );
  INVX0 U5784_U2 ( .INP(WX11121), .ZN(U5784_n1) );
  NOR2X0 U5784_U1 ( .IN1(n4529), .IN2(U5784_n1), .QN(WX11184) );
  INVX0 U5785_U2 ( .INP(WX11119), .ZN(U5785_n1) );
  NOR2X0 U5785_U1 ( .IN1(n4529), .IN2(U5785_n1), .QN(WX11182) );
  INVX0 U5786_U2 ( .INP(WX11117), .ZN(U5786_n1) );
  NOR2X0 U5786_U1 ( .IN1(n4529), .IN2(U5786_n1), .QN(WX11180) );
  INVX0 U5787_U2 ( .INP(WX11115), .ZN(U5787_n1) );
  NOR2X0 U5787_U1 ( .IN1(n4529), .IN2(U5787_n1), .QN(WX11178) );
  INVX0 U5788_U2 ( .INP(WX11113), .ZN(U5788_n1) );
  NOR2X0 U5788_U1 ( .IN1(n4530), .IN2(U5788_n1), .QN(WX11176) );
  INVX0 U5789_U2 ( .INP(WX11111), .ZN(U5789_n1) );
  NOR2X0 U5789_U1 ( .IN1(n4530), .IN2(U5789_n1), .QN(WX11174) );
  INVX0 U5790_U2 ( .INP(WX11109), .ZN(U5790_n1) );
  NOR2X0 U5790_U1 ( .IN1(n4530), .IN2(U5790_n1), .QN(WX11172) );
  INVX0 U5791_U2 ( .INP(WX11107), .ZN(U5791_n1) );
  NOR2X0 U5791_U1 ( .IN1(n4530), .IN2(U5791_n1), .QN(WX11170) );
  INVX0 U5792_U2 ( .INP(WX11105), .ZN(U5792_n1) );
  NOR2X0 U5792_U1 ( .IN1(n4530), .IN2(U5792_n1), .QN(WX11168) );
  INVX0 U5793_U2 ( .INP(test_so94), .ZN(U5793_n1) );
  NOR2X0 U5793_U1 ( .IN1(n4530), .IN2(U5793_n1), .QN(WX11166) );
  INVX0 U5794_U2 ( .INP(WX11101), .ZN(U5794_n1) );
  NOR2X0 U5794_U1 ( .IN1(n4530), .IN2(U5794_n1), .QN(WX11164) );
  INVX0 U5795_U2 ( .INP(WX11099), .ZN(U5795_n1) );
  NOR2X0 U5795_U1 ( .IN1(n4530), .IN2(U5795_n1), .QN(WX11162) );
  INVX0 U5796_U2 ( .INP(WX11097), .ZN(U5796_n1) );
  NOR2X0 U5796_U1 ( .IN1(n4530), .IN2(U5796_n1), .QN(WX11160) );
  INVX0 U5797_U2 ( .INP(WX11095), .ZN(U5797_n1) );
  NOR2X0 U5797_U1 ( .IN1(n4530), .IN2(U5797_n1), .QN(WX11158) );
  INVX0 U5798_U2 ( .INP(WX11093), .ZN(U5798_n1) );
  NOR2X0 U5798_U1 ( .IN1(n4530), .IN2(U5798_n1), .QN(WX11156) );
  INVX0 U5799_U2 ( .INP(WX11091), .ZN(U5799_n1) );
  NOR2X0 U5799_U1 ( .IN1(n4530), .IN2(U5799_n1), .QN(WX11154) );
  INVX0 U5800_U2 ( .INP(WX11089), .ZN(U5800_n1) );
  NOR2X0 U5800_U1 ( .IN1(n4530), .IN2(U5800_n1), .QN(WX11152) );
  INVX0 U5801_U2 ( .INP(WX11087), .ZN(U5801_n1) );
  NOR2X0 U5801_U1 ( .IN1(n4531), .IN2(U5801_n1), .QN(WX11150) );
  INVX0 U5802_U2 ( .INP(WX11085), .ZN(U5802_n1) );
  NOR2X0 U5802_U1 ( .IN1(n4531), .IN2(U5802_n1), .QN(WX11148) );
  INVX0 U5803_U2 ( .INP(WX11083), .ZN(U5803_n1) );
  NOR2X0 U5803_U1 ( .IN1(n4531), .IN2(U5803_n1), .QN(WX11146) );
  INVX0 U5804_U2 ( .INP(WX11081), .ZN(U5804_n1) );
  NOR2X0 U5804_U1 ( .IN1(n4531), .IN2(U5804_n1), .QN(WX11144) );
  INVX0 U5805_U2 ( .INP(WX11079), .ZN(U5805_n1) );
  NOR2X0 U5805_U1 ( .IN1(n4531), .IN2(U5805_n1), .QN(WX11142) );
  INVX0 U5806_U2 ( .INP(WX11077), .ZN(U5806_n1) );
  NOR2X0 U5806_U1 ( .IN1(n4531), .IN2(U5806_n1), .QN(WX11140) );
  INVX0 U5807_U2 ( .INP(WX11075), .ZN(U5807_n1) );
  NOR2X0 U5807_U1 ( .IN1(n4531), .IN2(U5807_n1), .QN(WX11138) );
  INVX0 U5808_U2 ( .INP(WX11073), .ZN(U5808_n1) );
  NOR2X0 U5808_U1 ( .IN1(n4531), .IN2(U5808_n1), .QN(WX11136) );
  INVX0 U5809_U2 ( .INP(WX11071), .ZN(U5809_n1) );
  NOR2X0 U5809_U1 ( .IN1(n4531), .IN2(U5809_n1), .QN(WX11134) );
  INVX0 U5810_U2 ( .INP(test_so93), .ZN(U5810_n1) );
  NOR2X0 U5810_U1 ( .IN1(n4531), .IN2(U5810_n1), .QN(WX11132) );
  INVX0 U5811_U2 ( .INP(WX11067), .ZN(U5811_n1) );
  NOR2X0 U5811_U1 ( .IN1(n4531), .IN2(U5811_n1), .QN(WX11130) );
  INVX0 U5812_U2 ( .INP(WX11065), .ZN(U5812_n1) );
  NOR2X0 U5812_U1 ( .IN1(n4531), .IN2(U5812_n1), .QN(WX11128) );
  INVX0 U5813_U2 ( .INP(WX11063), .ZN(U5813_n1) );
  NOR2X0 U5813_U1 ( .IN1(n4531), .IN2(U5813_n1), .QN(WX11126) );
  INVX0 U5814_U2 ( .INP(WX11061), .ZN(U5814_n1) );
  NOR2X0 U5814_U1 ( .IN1(n4532), .IN2(U5814_n1), .QN(WX11124) );
  INVX0 U5815_U2 ( .INP(WX11059), .ZN(U5815_n1) );
  NOR2X0 U5815_U1 ( .IN1(n4532), .IN2(U5815_n1), .QN(WX11122) );
  INVX0 U5816_U2 ( .INP(WX11057), .ZN(U5816_n1) );
  NOR2X0 U5816_U1 ( .IN1(n4532), .IN2(U5816_n1), .QN(WX11120) );
  INVX0 U5817_U2 ( .INP(WX11055), .ZN(U5817_n1) );
  NOR2X0 U5817_U1 ( .IN1(n4532), .IN2(U5817_n1), .QN(WX11118) );
  INVX0 U5818_U2 ( .INP(WX11053), .ZN(U5818_n1) );
  NOR2X0 U5818_U1 ( .IN1(n4532), .IN2(U5818_n1), .QN(WX11116) );
  INVX0 U5819_U2 ( .INP(WX11051), .ZN(U5819_n1) );
  NOR2X0 U5819_U1 ( .IN1(n4532), .IN2(U5819_n1), .QN(WX11114) );
  INVX0 U5820_U2 ( .INP(WX11049), .ZN(U5820_n1) );
  NOR2X0 U5820_U1 ( .IN1(n4532), .IN2(U5820_n1), .QN(WX11112) );
  INVX0 U5821_U2 ( .INP(WX11047), .ZN(U5821_n1) );
  NOR2X0 U5821_U1 ( .IN1(n4532), .IN2(U5821_n1), .QN(WX11110) );
  INVX0 U5822_U2 ( .INP(WX11045), .ZN(U5822_n1) );
  NOR2X0 U5822_U1 ( .IN1(n4532), .IN2(U5822_n1), .QN(WX11108) );
  INVX0 U5823_U2 ( .INP(WX11043), .ZN(U5823_n1) );
  NOR2X0 U5823_U1 ( .IN1(n4532), .IN2(U5823_n1), .QN(WX11106) );
  INVX0 U5824_U2 ( .INP(WX11041), .ZN(U5824_n1) );
  NOR2X0 U5824_U1 ( .IN1(n4532), .IN2(U5824_n1), .QN(WX11104) );
  INVX0 U5825_U2 ( .INP(WX11039), .ZN(U5825_n1) );
  NOR2X0 U5825_U1 ( .IN1(n4532), .IN2(U5825_n1), .QN(WX11102) );
  INVX0 U5826_U2 ( .INP(WX11037), .ZN(U5826_n1) );
  NOR2X0 U5826_U1 ( .IN1(n4532), .IN2(U5826_n1), .QN(WX11100) );
  INVX0 U5827_U2 ( .INP(test_so92), .ZN(U5827_n1) );
  NOR2X0 U5827_U1 ( .IN1(n4533), .IN2(U5827_n1), .QN(WX11098) );
  INVX0 U5828_U2 ( .INP(WX11033), .ZN(U5828_n1) );
  NOR2X0 U5828_U1 ( .IN1(n4533), .IN2(U5828_n1), .QN(WX11096) );
  INVX0 U5829_U2 ( .INP(WX11031), .ZN(U5829_n1) );
  NOR2X0 U5829_U1 ( .IN1(n4520), .IN2(U5829_n1), .QN(WX11094) );
  INVX0 U5830_U2 ( .INP(WX11029), .ZN(U5830_n1) );
  NOR2X0 U5830_U1 ( .IN1(n4516), .IN2(U5830_n1), .QN(WX11092) );
  INVX0 U5831_U2 ( .INP(WX11027), .ZN(U5831_n1) );
  NOR2X0 U5831_U1 ( .IN1(n4516), .IN2(U5831_n1), .QN(WX11090) );
  INVX0 U5832_U2 ( .INP(WX11025), .ZN(U5832_n1) );
  NOR2X0 U5832_U1 ( .IN1(n4516), .IN2(U5832_n1), .QN(WX11088) );
  INVX0 U5833_U2 ( .INP(WX11023), .ZN(U5833_n1) );
  NOR2X0 U5833_U1 ( .IN1(n4516), .IN2(U5833_n1), .QN(WX11086) );
  INVX0 U5834_U2 ( .INP(WX11021), .ZN(U5834_n1) );
  NOR2X0 U5834_U1 ( .IN1(n4516), .IN2(U5834_n1), .QN(WX11084) );
  INVX0 U5835_U2 ( .INP(WX9886), .ZN(U5835_n1) );
  NOR2X0 U5835_U1 ( .IN1(n4516), .IN2(U5835_n1), .QN(WX9949) );
  INVX0 U5836_U2 ( .INP(WX9884), .ZN(U5836_n1) );
  NOR2X0 U5836_U1 ( .IN1(n4516), .IN2(U5836_n1), .QN(WX9947) );
  INVX0 U5837_U2 ( .INP(WX9882), .ZN(U5837_n1) );
  NOR2X0 U5837_U1 ( .IN1(n4516), .IN2(U5837_n1), .QN(WX9945) );
  INVX0 U5838_U2 ( .INP(WX9880), .ZN(U5838_n1) );
  NOR2X0 U5838_U1 ( .IN1(n4516), .IN2(U5838_n1), .QN(WX9943) );
  INVX0 U5839_U2 ( .INP(WX9878), .ZN(U5839_n1) );
  NOR2X0 U5839_U1 ( .IN1(n4516), .IN2(U5839_n1), .QN(WX9941) );
  INVX0 U5840_U2 ( .INP(WX9876), .ZN(U5840_n1) );
  NOR2X0 U5840_U1 ( .IN1(n4516), .IN2(U5840_n1), .QN(WX9939) );
  INVX0 U5841_U2 ( .INP(WX9874), .ZN(U5841_n1) );
  NOR2X0 U5841_U1 ( .IN1(n4516), .IN2(U5841_n1), .QN(WX9937) );
  INVX0 U5842_U2 ( .INP(WX9872), .ZN(U5842_n1) );
  NOR2X0 U5842_U1 ( .IN1(n4517), .IN2(U5842_n1), .QN(WX9935) );
  INVX0 U5843_U2 ( .INP(WX9870), .ZN(U5843_n1) );
  NOR2X0 U5843_U1 ( .IN1(n4517), .IN2(U5843_n1), .QN(WX9933) );
  INVX0 U5844_U2 ( .INP(WX9868), .ZN(U5844_n1) );
  NOR2X0 U5844_U1 ( .IN1(n4517), .IN2(U5844_n1), .QN(WX9931) );
  INVX0 U5845_U2 ( .INP(WX9866), .ZN(U5845_n1) );
  NOR2X0 U5845_U1 ( .IN1(n4517), .IN2(U5845_n1), .QN(WX9929) );
  INVX0 U5846_U2 ( .INP(WX9864), .ZN(U5846_n1) );
  NOR2X0 U5846_U1 ( .IN1(n4517), .IN2(U5846_n1), .QN(WX9927) );
  INVX0 U5847_U2 ( .INP(WX9862), .ZN(U5847_n1) );
  NOR2X0 U5847_U1 ( .IN1(n4517), .IN2(U5847_n1), .QN(WX9925) );
  INVX0 U5848_U2 ( .INP(WX9860), .ZN(U5848_n1) );
  NOR2X0 U5848_U1 ( .IN1(n4517), .IN2(U5848_n1), .QN(WX9923) );
  INVX0 U5849_U2 ( .INP(WX9858), .ZN(U5849_n1) );
  NOR2X0 U5849_U1 ( .IN1(n4517), .IN2(U5849_n1), .QN(WX9921) );
  INVX0 U5850_U2 ( .INP(WX9856), .ZN(U5850_n1) );
  NOR2X0 U5850_U1 ( .IN1(n4517), .IN2(U5850_n1), .QN(WX9919) );
  INVX0 U5851_U2 ( .INP(test_so84), .ZN(U5851_n1) );
  NOR2X0 U5851_U1 ( .IN1(n4517), .IN2(U5851_n1), .QN(WX9917) );
  INVX0 U5852_U2 ( .INP(WX9852), .ZN(U5852_n1) );
  NOR2X0 U5852_U1 ( .IN1(n4517), .IN2(U5852_n1), .QN(WX9915) );
  INVX0 U5853_U2 ( .INP(WX9850), .ZN(U5853_n1) );
  NOR2X0 U5853_U1 ( .IN1(n4517), .IN2(U5853_n1), .QN(WX9913) );
  INVX0 U5854_U2 ( .INP(WX9848), .ZN(U5854_n1) );
  NOR2X0 U5854_U1 ( .IN1(n4517), .IN2(U5854_n1), .QN(WX9911) );
  INVX0 U5855_U2 ( .INP(WX9846), .ZN(U5855_n1) );
  NOR2X0 U5855_U1 ( .IN1(n4518), .IN2(U5855_n1), .QN(WX9909) );
  INVX0 U5856_U2 ( .INP(WX9844), .ZN(U5856_n1) );
  NOR2X0 U5856_U1 ( .IN1(n4518), .IN2(U5856_n1), .QN(WX9907) );
  INVX0 U5857_U2 ( .INP(WX9842), .ZN(U5857_n1) );
  NOR2X0 U5857_U1 ( .IN1(n4518), .IN2(U5857_n1), .QN(WX9905) );
  INVX0 U5858_U2 ( .INP(WX9840), .ZN(U5858_n1) );
  NOR2X0 U5858_U1 ( .IN1(n4518), .IN2(U5858_n1), .QN(WX9903) );
  INVX0 U5859_U2 ( .INP(WX9838), .ZN(U5859_n1) );
  NOR2X0 U5859_U1 ( .IN1(n4518), .IN2(U5859_n1), .QN(WX9901) );
  INVX0 U5860_U2 ( .INP(WX9836), .ZN(U5860_n1) );
  NOR2X0 U5860_U1 ( .IN1(n4518), .IN2(U5860_n1), .QN(WX9899) );
  INVX0 U5861_U2 ( .INP(WX9834), .ZN(U5861_n1) );
  NOR2X0 U5861_U1 ( .IN1(n4518), .IN2(U5861_n1), .QN(WX9897) );
  INVX0 U5862_U2 ( .INP(WX9832), .ZN(U5862_n1) );
  NOR2X0 U5862_U1 ( .IN1(n4518), .IN2(U5862_n1), .QN(WX9895) );
  INVX0 U5863_U2 ( .INP(WX9830), .ZN(U5863_n1) );
  NOR2X0 U5863_U1 ( .IN1(n4518), .IN2(U5863_n1), .QN(WX9893) );
  INVX0 U5864_U2 ( .INP(WX9828), .ZN(U5864_n1) );
  NOR2X0 U5864_U1 ( .IN1(n4518), .IN2(U5864_n1), .QN(WX9891) );
  INVX0 U5865_U2 ( .INP(WX9826), .ZN(U5865_n1) );
  NOR2X0 U5865_U1 ( .IN1(n4518), .IN2(U5865_n1), .QN(WX9889) );
  INVX0 U5866_U2 ( .INP(WX9824), .ZN(U5866_n1) );
  NOR2X0 U5866_U1 ( .IN1(n4518), .IN2(U5866_n1), .QN(WX9887) );
  INVX0 U5867_U2 ( .INP(WX9822), .ZN(U5867_n1) );
  NOR2X0 U5867_U1 ( .IN1(n4518), .IN2(U5867_n1), .QN(WX9885) );
  INVX0 U5868_U2 ( .INP(test_so83), .ZN(U5868_n1) );
  NOR2X0 U5868_U1 ( .IN1(n4519), .IN2(U5868_n1), .QN(WX9883) );
  INVX0 U5869_U2 ( .INP(WX9818), .ZN(U5869_n1) );
  NOR2X0 U5869_U1 ( .IN1(n4519), .IN2(U5869_n1), .QN(WX9881) );
  INVX0 U5870_U2 ( .INP(WX9816), .ZN(U5870_n1) );
  NOR2X0 U5870_U1 ( .IN1(n4519), .IN2(U5870_n1), .QN(WX9879) );
  INVX0 U5871_U2 ( .INP(WX9814), .ZN(U5871_n1) );
  NOR2X0 U5871_U1 ( .IN1(n4519), .IN2(U5871_n1), .QN(WX9877) );
  INVX0 U5872_U2 ( .INP(WX9812), .ZN(U5872_n1) );
  NOR2X0 U5872_U1 ( .IN1(n4519), .IN2(U5872_n1), .QN(WX9875) );
  INVX0 U5873_U2 ( .INP(WX9810), .ZN(U5873_n1) );
  NOR2X0 U5873_U1 ( .IN1(n4519), .IN2(U5873_n1), .QN(WX9873) );
  INVX0 U5874_U2 ( .INP(WX9808), .ZN(U5874_n1) );
  NOR2X0 U5874_U1 ( .IN1(n4519), .IN2(U5874_n1), .QN(WX9871) );
  INVX0 U5875_U2 ( .INP(WX9806), .ZN(U5875_n1) );
  NOR2X0 U5875_U1 ( .IN1(n4519), .IN2(U5875_n1), .QN(WX9869) );
  INVX0 U5876_U2 ( .INP(WX9804), .ZN(U5876_n1) );
  NOR2X0 U5876_U1 ( .IN1(n4519), .IN2(U5876_n1), .QN(WX9867) );
  INVX0 U5877_U2 ( .INP(WX9802), .ZN(U5877_n1) );
  NOR2X0 U5877_U1 ( .IN1(n4519), .IN2(U5877_n1), .QN(WX9865) );
  INVX0 U5878_U2 ( .INP(WX9800), .ZN(U5878_n1) );
  NOR2X0 U5878_U1 ( .IN1(n4519), .IN2(U5878_n1), .QN(WX9863) );
  INVX0 U5879_U2 ( .INP(WX9798), .ZN(U5879_n1) );
  NOR2X0 U5879_U1 ( .IN1(n4519), .IN2(U5879_n1), .QN(WX9861) );
  INVX0 U5880_U2 ( .INP(WX9796), .ZN(U5880_n1) );
  NOR2X0 U5880_U1 ( .IN1(n4519), .IN2(U5880_n1), .QN(WX9859) );
  INVX0 U5881_U2 ( .INP(WX9794), .ZN(U5881_n1) );
  NOR2X0 U5881_U1 ( .IN1(n4520), .IN2(U5881_n1), .QN(WX9857) );
  INVX0 U5882_U2 ( .INP(WX9792), .ZN(U5882_n1) );
  NOR2X0 U5882_U1 ( .IN1(n4520), .IN2(U5882_n1), .QN(WX9855) );
  INVX0 U5883_U2 ( .INP(WX9790), .ZN(U5883_n1) );
  NOR2X0 U5883_U1 ( .IN1(n4520), .IN2(U5883_n1), .QN(WX9853) );
  INVX0 U5884_U2 ( .INP(WX9788), .ZN(U5884_n1) );
  NOR2X0 U5884_U1 ( .IN1(n4520), .IN2(U5884_n1), .QN(WX9851) );
  INVX0 U5885_U2 ( .INP(test_so82), .ZN(U5885_n1) );
  NOR2X0 U5885_U1 ( .IN1(n4520), .IN2(U5885_n1), .QN(WX9849) );
  INVX0 U5886_U2 ( .INP(WX9784), .ZN(U5886_n1) );
  NOR2X0 U5886_U1 ( .IN1(n4520), .IN2(U5886_n1), .QN(WX9847) );
  INVX0 U5887_U2 ( .INP(WX9782), .ZN(U5887_n1) );
  NOR2X0 U5887_U1 ( .IN1(n4520), .IN2(U5887_n1), .QN(WX9845) );
  INVX0 U5888_U2 ( .INP(WX9780), .ZN(U5888_n1) );
  NOR2X0 U5888_U1 ( .IN1(n4520), .IN2(U5888_n1), .QN(WX9843) );
  INVX0 U5889_U2 ( .INP(WX9778), .ZN(U5889_n1) );
  NOR2X0 U5889_U1 ( .IN1(n4520), .IN2(U5889_n1), .QN(WX9841) );
  INVX0 U5890_U2 ( .INP(WX9776), .ZN(U5890_n1) );
  NOR2X0 U5890_U1 ( .IN1(n4520), .IN2(U5890_n1), .QN(WX9839) );
  INVX0 U5891_U2 ( .INP(WX9774), .ZN(U5891_n1) );
  NOR2X0 U5891_U1 ( .IN1(n4520), .IN2(U5891_n1), .QN(WX9837) );
  INVX0 U5892_U2 ( .INP(WX9772), .ZN(U5892_n1) );
  NOR2X0 U5892_U1 ( .IN1(n4520), .IN2(U5892_n1), .QN(WX9835) );
  INVX0 U5893_U2 ( .INP(WX9770), .ZN(U5893_n1) );
  NOR2X0 U5893_U1 ( .IN1(n4521), .IN2(U5893_n1), .QN(WX9833) );
  INVX0 U5894_U2 ( .INP(WX9768), .ZN(U5894_n1) );
  NOR2X0 U5894_U1 ( .IN1(n4521), .IN2(U5894_n1), .QN(WX9831) );
  INVX0 U5895_U2 ( .INP(WX9766), .ZN(U5895_n1) );
  NOR2X0 U5895_U1 ( .IN1(n4521), .IN2(U5895_n1), .QN(WX9829) );
  INVX0 U5896_U2 ( .INP(WX9764), .ZN(U5896_n1) );
  NOR2X0 U5896_U1 ( .IN1(n4521), .IN2(U5896_n1), .QN(WX9827) );
  INVX0 U5897_U2 ( .INP(WX9762), .ZN(U5897_n1) );
  NOR2X0 U5897_U1 ( .IN1(n4521), .IN2(U5897_n1), .QN(WX9825) );
  INVX0 U5898_U2 ( .INP(WX9760), .ZN(U5898_n1) );
  NOR2X0 U5898_U1 ( .IN1(n4521), .IN2(U5898_n1), .QN(WX9823) );
  INVX0 U5899_U2 ( .INP(WX9758), .ZN(U5899_n1) );
  NOR2X0 U5899_U1 ( .IN1(n4521), .IN2(U5899_n1), .QN(WX9821) );
  INVX0 U5900_U2 ( .INP(WX9756), .ZN(U5900_n1) );
  NOR2X0 U5900_U1 ( .IN1(n4521), .IN2(U5900_n1), .QN(WX9819) );
  INVX0 U5901_U2 ( .INP(WX9754), .ZN(U5901_n1) );
  NOR2X0 U5901_U1 ( .IN1(n4521), .IN2(U5901_n1), .QN(WX9817) );
  INVX0 U5902_U2 ( .INP(test_so81), .ZN(U5902_n1) );
  NOR2X0 U5902_U1 ( .IN1(n4521), .IN2(U5902_n1), .QN(WX9815) );
  INVX0 U5903_U2 ( .INP(WX9750), .ZN(U5903_n1) );
  NOR2X0 U5903_U1 ( .IN1(n4521), .IN2(U5903_n1), .QN(WX9813) );
  INVX0 U5904_U2 ( .INP(WX9748), .ZN(U5904_n1) );
  NOR2X0 U5904_U1 ( .IN1(n4521), .IN2(U5904_n1), .QN(WX9811) );
  INVX0 U5905_U2 ( .INP(WX9746), .ZN(U5905_n1) );
  NOR2X0 U5905_U1 ( .IN1(n4521), .IN2(U5905_n1), .QN(WX9809) );
  INVX0 U5906_U2 ( .INP(WX9744), .ZN(U5906_n1) );
  NOR2X0 U5906_U1 ( .IN1(n4522), .IN2(U5906_n1), .QN(WX9807) );
  INVX0 U5907_U2 ( .INP(WX9742), .ZN(U5907_n1) );
  NOR2X0 U5907_U1 ( .IN1(n4522), .IN2(U5907_n1), .QN(WX9805) );
  INVX0 U5908_U2 ( .INP(WX9740), .ZN(U5908_n1) );
  NOR2X0 U5908_U1 ( .IN1(n4522), .IN2(U5908_n1), .QN(WX9803) );
  INVX0 U5909_U2 ( .INP(WX9738), .ZN(U5909_n1) );
  NOR2X0 U5909_U1 ( .IN1(n4522), .IN2(U5909_n1), .QN(WX9801) );
  INVX0 U5910_U2 ( .INP(WX9736), .ZN(U5910_n1) );
  NOR2X0 U5910_U1 ( .IN1(n4522), .IN2(U5910_n1), .QN(WX9799) );
  INVX0 U5911_U2 ( .INP(WX9734), .ZN(U5911_n1) );
  NOR2X0 U5911_U1 ( .IN1(n4522), .IN2(U5911_n1), .QN(WX9797) );
  INVX0 U5912_U2 ( .INP(WX9732), .ZN(U5912_n1) );
  NOR2X0 U5912_U1 ( .IN1(n4522), .IN2(U5912_n1), .QN(WX9795) );
  INVX0 U5913_U2 ( .INP(WX9730), .ZN(U5913_n1) );
  NOR2X0 U5913_U1 ( .IN1(n4522), .IN2(U5913_n1), .QN(WX9793) );
  INVX0 U5914_U2 ( .INP(WX9728), .ZN(U5914_n1) );
  NOR2X0 U5914_U1 ( .IN1(n4522), .IN2(U5914_n1), .QN(WX9791) );
  INVX0 U5915_U2 ( .INP(WX8593), .ZN(U5915_n1) );
  NOR2X0 U5915_U1 ( .IN1(n4522), .IN2(U5915_n1), .QN(WX8656) );
  INVX0 U5916_U2 ( .INP(WX8591), .ZN(U5916_n1) );
  NOR2X0 U5916_U1 ( .IN1(n4522), .IN2(U5916_n1), .QN(WX8654) );
  INVX0 U5917_U2 ( .INP(WX8589), .ZN(U5917_n1) );
  NOR2X0 U5917_U1 ( .IN1(n4522), .IN2(U5917_n1), .QN(WX8652) );
  INVX0 U5918_U2 ( .INP(WX8587), .ZN(U5918_n1) );
  NOR2X0 U5918_U1 ( .IN1(n4522), .IN2(U5918_n1), .QN(WX8650) );
  INVX0 U5919_U2 ( .INP(WX8585), .ZN(U5919_n1) );
  NOR2X0 U5919_U1 ( .IN1(n4523), .IN2(U5919_n1), .QN(WX8648) );
  INVX0 U5920_U2 ( .INP(WX8583), .ZN(U5920_n1) );
  NOR2X0 U5920_U1 ( .IN1(n4523), .IN2(U5920_n1), .QN(WX8646) );
  INVX0 U5921_U2 ( .INP(WX8581), .ZN(U5921_n1) );
  NOR2X0 U5921_U1 ( .IN1(n4523), .IN2(U5921_n1), .QN(WX8644) );
  INVX0 U5922_U2 ( .INP(WX8579), .ZN(U5922_n1) );
  NOR2X0 U5922_U1 ( .IN1(n4523), .IN2(U5922_n1), .QN(WX8642) );
  INVX0 U5923_U2 ( .INP(WX8577), .ZN(U5923_n1) );
  NOR2X0 U5923_U1 ( .IN1(n4523), .IN2(U5923_n1), .QN(WX8640) );
  INVX0 U5924_U2 ( .INP(WX8575), .ZN(U5924_n1) );
  NOR2X0 U5924_U1 ( .IN1(n4523), .IN2(U5924_n1), .QN(WX8638) );
  INVX0 U5925_U2 ( .INP(WX8573), .ZN(U5925_n1) );
  NOR2X0 U5925_U1 ( .IN1(n4523), .IN2(U5925_n1), .QN(WX8636) );
  INVX0 U5926_U2 ( .INP(test_so73), .ZN(U5926_n1) );
  NOR2X0 U5926_U1 ( .IN1(n4523), .IN2(U5926_n1), .QN(WX8634) );
  INVX0 U5927_U2 ( .INP(WX8569), .ZN(U5927_n1) );
  NOR2X0 U5927_U1 ( .IN1(n4523), .IN2(U5927_n1), .QN(WX8632) );
  INVX0 U5928_U2 ( .INP(WX8567), .ZN(U5928_n1) );
  NOR2X0 U5928_U1 ( .IN1(n4523), .IN2(U5928_n1), .QN(WX8630) );
  INVX0 U5929_U2 ( .INP(WX8565), .ZN(U5929_n1) );
  NOR2X0 U5929_U1 ( .IN1(n4523), .IN2(U5929_n1), .QN(WX8628) );
  INVX0 U5930_U2 ( .INP(WX8563), .ZN(U5930_n1) );
  NOR2X0 U5930_U1 ( .IN1(n4523), .IN2(U5930_n1), .QN(WX8626) );
  INVX0 U5931_U2 ( .INP(WX8561), .ZN(U5931_n1) );
  NOR2X0 U5931_U1 ( .IN1(n4523), .IN2(U5931_n1), .QN(WX8624) );
  INVX0 U5932_U2 ( .INP(WX8559), .ZN(U5932_n1) );
  NOR2X0 U5932_U1 ( .IN1(n4524), .IN2(U5932_n1), .QN(WX8622) );
  INVX0 U5933_U2 ( .INP(WX8557), .ZN(U5933_n1) );
  NOR2X0 U5933_U1 ( .IN1(n4524), .IN2(U5933_n1), .QN(WX8620) );
  INVX0 U5934_U2 ( .INP(WX8555), .ZN(U5934_n1) );
  NOR2X0 U5934_U1 ( .IN1(n4524), .IN2(U5934_n1), .QN(WX8618) );
  INVX0 U5935_U2 ( .INP(WX8553), .ZN(U5935_n1) );
  NOR2X0 U5935_U1 ( .IN1(n4524), .IN2(U5935_n1), .QN(WX8616) );
  INVX0 U5936_U2 ( .INP(WX8551), .ZN(U5936_n1) );
  NOR2X0 U5936_U1 ( .IN1(n4524), .IN2(U5936_n1), .QN(WX8614) );
  INVX0 U5937_U2 ( .INP(WX8549), .ZN(U5937_n1) );
  NOR2X0 U5937_U1 ( .IN1(n4524), .IN2(U5937_n1), .QN(WX8612) );
  INVX0 U5938_U2 ( .INP(WX8547), .ZN(U5938_n1) );
  NOR2X0 U5938_U1 ( .IN1(n4524), .IN2(U5938_n1), .QN(WX8610) );
  INVX0 U5939_U2 ( .INP(WX8545), .ZN(U5939_n1) );
  NOR2X0 U5939_U1 ( .IN1(n4524), .IN2(U5939_n1), .QN(WX8608) );
  INVX0 U5940_U2 ( .INP(WX8543), .ZN(U5940_n1) );
  NOR2X0 U5940_U1 ( .IN1(n4543), .IN2(U5940_n1), .QN(WX8606) );
  INVX0 U5941_U2 ( .INP(WX8541), .ZN(U5941_n1) );
  NOR2X0 U5941_U1 ( .IN1(n4541), .IN2(U5941_n1), .QN(WX8604) );
  INVX0 U5942_U2 ( .INP(WX8539), .ZN(U5942_n1) );
  NOR2X0 U5942_U1 ( .IN1(n4541), .IN2(U5942_n1), .QN(WX8602) );
  INVX0 U5943_U2 ( .INP(test_so72), .ZN(U5943_n1) );
  NOR2X0 U5943_U1 ( .IN1(n4541), .IN2(U5943_n1), .QN(WX8600) );
  INVX0 U5944_U2 ( .INP(WX8535), .ZN(U5944_n1) );
  NOR2X0 U5944_U1 ( .IN1(n4546), .IN2(U5944_n1), .QN(WX8598) );
  INVX0 U5945_U2 ( .INP(WX8533), .ZN(U5945_n1) );
  NOR2X0 U5945_U1 ( .IN1(n4543), .IN2(U5945_n1), .QN(WX8596) );
  INVX0 U5946_U2 ( .INP(WX8531), .ZN(U5946_n1) );
  NOR2X0 U5946_U1 ( .IN1(n4543), .IN2(U5946_n1), .QN(WX8594) );
  INVX0 U5947_U2 ( .INP(WX8529), .ZN(U5947_n1) );
  NOR2X0 U5947_U1 ( .IN1(n4543), .IN2(U5947_n1), .QN(WX8592) );
  INVX0 U5948_U2 ( .INP(WX8527), .ZN(U5948_n1) );
  NOR2X0 U5948_U1 ( .IN1(n4543), .IN2(U5948_n1), .QN(WX8590) );
  INVX0 U5949_U2 ( .INP(WX8525), .ZN(U5949_n1) );
  NOR2X0 U5949_U1 ( .IN1(n4543), .IN2(U5949_n1), .QN(WX8588) );
  INVX0 U5950_U2 ( .INP(WX8523), .ZN(U5950_n1) );
  NOR2X0 U5950_U1 ( .IN1(n4543), .IN2(U5950_n1), .QN(WX8586) );
  INVX0 U5951_U2 ( .INP(WX8521), .ZN(U5951_n1) );
  NOR2X0 U5951_U1 ( .IN1(n4543), .IN2(U5951_n1), .QN(WX8584) );
  INVX0 U5952_U2 ( .INP(WX8519), .ZN(U5952_n1) );
  NOR2X0 U5952_U1 ( .IN1(n4543), .IN2(U5952_n1), .QN(WX8582) );
  INVX0 U5953_U2 ( .INP(WX8517), .ZN(U5953_n1) );
  NOR2X0 U5953_U1 ( .IN1(n4542), .IN2(U5953_n1), .QN(WX8580) );
  INVX0 U5954_U2 ( .INP(WX8515), .ZN(U5954_n1) );
  NOR2X0 U5954_U1 ( .IN1(n4542), .IN2(U5954_n1), .QN(WX8578) );
  INVX0 U5955_U2 ( .INP(WX8513), .ZN(U5955_n1) );
  NOR2X0 U5955_U1 ( .IN1(n4542), .IN2(U5955_n1), .QN(WX8576) );
  INVX0 U5956_U2 ( .INP(WX8511), .ZN(U5956_n1) );
  NOR2X0 U5956_U1 ( .IN1(n4542), .IN2(U5956_n1), .QN(WX8574) );
  INVX0 U5957_U2 ( .INP(WX8509), .ZN(U5957_n1) );
  NOR2X0 U5957_U1 ( .IN1(n4542), .IN2(U5957_n1), .QN(WX8572) );
  INVX0 U5958_U2 ( .INP(WX8507), .ZN(U5958_n1) );
  NOR2X0 U5958_U1 ( .IN1(n4542), .IN2(U5958_n1), .QN(WX8570) );
  INVX0 U5959_U2 ( .INP(WX8505), .ZN(U5959_n1) );
  NOR2X0 U5959_U1 ( .IN1(n4542), .IN2(U5959_n1), .QN(WX8568) );
  INVX0 U5960_U2 ( .INP(test_so71), .ZN(U5960_n1) );
  NOR2X0 U5960_U1 ( .IN1(n4542), .IN2(U5960_n1), .QN(WX8566) );
  INVX0 U5961_U2 ( .INP(WX8501), .ZN(U5961_n1) );
  NOR2X0 U5961_U1 ( .IN1(n4542), .IN2(U5961_n1), .QN(WX8564) );
  INVX0 U5962_U2 ( .INP(WX8499), .ZN(U5962_n1) );
  NOR2X0 U5962_U1 ( .IN1(n4542), .IN2(U5962_n1), .QN(WX8562) );
  INVX0 U5963_U2 ( .INP(WX8497), .ZN(U5963_n1) );
  NOR2X0 U5963_U1 ( .IN1(n4542), .IN2(U5963_n1), .QN(WX8560) );
  INVX0 U5964_U2 ( .INP(WX8495), .ZN(U5964_n1) );
  NOR2X0 U5964_U1 ( .IN1(n4542), .IN2(U5964_n1), .QN(WX8558) );
  INVX0 U5965_U2 ( .INP(WX8493), .ZN(U5965_n1) );
  NOR2X0 U5965_U1 ( .IN1(n4542), .IN2(U5965_n1), .QN(WX8556) );
  INVX0 U5966_U2 ( .INP(WX8491), .ZN(U5966_n1) );
  NOR2X0 U5966_U1 ( .IN1(n4543), .IN2(U5966_n1), .QN(WX8554) );
  INVX0 U5967_U2 ( .INP(WX8489), .ZN(U5967_n1) );
  NOR2X0 U5967_U1 ( .IN1(n4543), .IN2(U5967_n1), .QN(WX8552) );
  INVX0 U5968_U2 ( .INP(WX8487), .ZN(U5968_n1) );
  NOR2X0 U5968_U1 ( .IN1(n4543), .IN2(U5968_n1), .QN(WX8550) );
  INVX0 U5969_U2 ( .INP(WX8485), .ZN(U5969_n1) );
  NOR2X0 U5969_U1 ( .IN1(n4543), .IN2(U5969_n1), .QN(WX8548) );
  INVX0 U5970_U2 ( .INP(WX8483), .ZN(U5970_n1) );
  NOR2X0 U5970_U1 ( .IN1(n4544), .IN2(U5970_n1), .QN(WX8546) );
  INVX0 U5971_U2 ( .INP(WX8481), .ZN(U5971_n1) );
  NOR2X0 U5971_U1 ( .IN1(n4544), .IN2(U5971_n1), .QN(WX8544) );
  INVX0 U5972_U2 ( .INP(WX8479), .ZN(U5972_n1) );
  NOR2X0 U5972_U1 ( .IN1(n4544), .IN2(U5972_n1), .QN(WX8542) );
  INVX0 U5973_U2 ( .INP(WX8477), .ZN(U5973_n1) );
  NOR2X0 U5973_U1 ( .IN1(n4544), .IN2(U5973_n1), .QN(WX8540) );
  INVX0 U5974_U2 ( .INP(WX8475), .ZN(U5974_n1) );
  NOR2X0 U5974_U1 ( .IN1(n4544), .IN2(U5974_n1), .QN(WX8538) );
  INVX0 U5975_U2 ( .INP(WX8473), .ZN(U5975_n1) );
  NOR2X0 U5975_U1 ( .IN1(n4544), .IN2(U5975_n1), .QN(WX8536) );
  INVX0 U5976_U2 ( .INP(WX8471), .ZN(U5976_n1) );
  NOR2X0 U5976_U1 ( .IN1(n4544), .IN2(U5976_n1), .QN(WX8534) );
  INVX0 U5977_U2 ( .INP(test_so70), .ZN(U5977_n1) );
  NOR2X0 U5977_U1 ( .IN1(n4544), .IN2(U5977_n1), .QN(WX8532) );
  INVX0 U5978_U2 ( .INP(WX8467), .ZN(U5978_n1) );
  NOR2X0 U5978_U1 ( .IN1(n4544), .IN2(U5978_n1), .QN(WX8530) );
  INVX0 U5979_U2 ( .INP(WX8465), .ZN(U5979_n1) );
  NOR2X0 U5979_U1 ( .IN1(n4544), .IN2(U5979_n1), .QN(WX8528) );
  INVX0 U5980_U2 ( .INP(WX8463), .ZN(U5980_n1) );
  NOR2X0 U5980_U1 ( .IN1(n4544), .IN2(U5980_n1), .QN(WX8526) );
  INVX0 U5981_U2 ( .INP(WX8461), .ZN(U5981_n1) );
  NOR2X0 U5981_U1 ( .IN1(n4544), .IN2(U5981_n1), .QN(WX8524) );
  INVX0 U5982_U2 ( .INP(WX8459), .ZN(U5982_n1) );
  NOR2X0 U5982_U1 ( .IN1(n4544), .IN2(U5982_n1), .QN(WX8522) );
  INVX0 U5983_U2 ( .INP(WX8457), .ZN(U5983_n1) );
  NOR2X0 U5983_U1 ( .IN1(n4545), .IN2(U5983_n1), .QN(WX8520) );
  INVX0 U5984_U2 ( .INP(WX8455), .ZN(U5984_n1) );
  NOR2X0 U5984_U1 ( .IN1(n4545), .IN2(U5984_n1), .QN(WX8518) );
  INVX0 U5985_U2 ( .INP(WX8453), .ZN(U5985_n1) );
  NOR2X0 U5985_U1 ( .IN1(n4545), .IN2(U5985_n1), .QN(WX8516) );
  INVX0 U5986_U2 ( .INP(WX8451), .ZN(U5986_n1) );
  NOR2X0 U5986_U1 ( .IN1(n4545), .IN2(U5986_n1), .QN(WX8514) );
  INVX0 U5987_U2 ( .INP(WX8449), .ZN(U5987_n1) );
  NOR2X0 U5987_U1 ( .IN1(n4545), .IN2(U5987_n1), .QN(WX8512) );
  INVX0 U5988_U2 ( .INP(WX8447), .ZN(U5988_n1) );
  NOR2X0 U5988_U1 ( .IN1(n4545), .IN2(U5988_n1), .QN(WX8510) );
  INVX0 U5989_U2 ( .INP(WX8445), .ZN(U5989_n1) );
  NOR2X0 U5989_U1 ( .IN1(n4545), .IN2(U5989_n1), .QN(WX8508) );
  INVX0 U5990_U2 ( .INP(WX8443), .ZN(U5990_n1) );
  NOR2X0 U5990_U1 ( .IN1(n4545), .IN2(U5990_n1), .QN(WX8506) );
  INVX0 U5991_U2 ( .INP(WX8441), .ZN(U5991_n1) );
  NOR2X0 U5991_U1 ( .IN1(n4545), .IN2(U5991_n1), .QN(WX8504) );
  INVX0 U5992_U2 ( .INP(WX8439), .ZN(U5992_n1) );
  NOR2X0 U5992_U1 ( .IN1(n4545), .IN2(U5992_n1), .QN(WX8502) );
  INVX0 U5993_U2 ( .INP(WX8437), .ZN(U5993_n1) );
  NOR2X0 U5993_U1 ( .IN1(n4545), .IN2(U5993_n1), .QN(WX8500) );
  INVX0 U5994_U2 ( .INP(test_so69), .ZN(U5994_n1) );
  NOR2X0 U5994_U1 ( .IN1(n4545), .IN2(U5994_n1), .QN(WX8498) );
  INVX0 U5995_U2 ( .INP(WX7300), .ZN(U5995_n1) );
  NOR2X0 U5995_U1 ( .IN1(n4545), .IN2(U5995_n1), .QN(WX7363) );
  INVX0 U5996_U2 ( .INP(WX7298), .ZN(U5996_n1) );
  NOR2X0 U5996_U1 ( .IN1(n4546), .IN2(U5996_n1), .QN(WX7361) );
  INVX0 U5997_U2 ( .INP(WX7296), .ZN(U5997_n1) );
  NOR2X0 U5997_U1 ( .IN1(n4546), .IN2(U5997_n1), .QN(WX7359) );
  INVX0 U5998_U2 ( .INP(WX7294), .ZN(U5998_n1) );
  NOR2X0 U5998_U1 ( .IN1(n4546), .IN2(U5998_n1), .QN(WX7357) );
  INVX0 U5999_U2 ( .INP(WX7292), .ZN(U5999_n1) );
  NOR2X0 U5999_U1 ( .IN1(n4546), .IN2(U5999_n1), .QN(WX7355) );
  INVX0 U6000_U2 ( .INP(WX7290), .ZN(U6000_n1) );
  NOR2X0 U6000_U1 ( .IN1(n4546), .IN2(U6000_n1), .QN(WX7353) );
  INVX0 U6001_U2 ( .INP(test_so62), .ZN(U6001_n1) );
  NOR2X0 U6001_U1 ( .IN1(n4546), .IN2(U6001_n1), .QN(WX7351) );
  INVX0 U6002_U2 ( .INP(WX7286), .ZN(U6002_n1) );
  NOR2X0 U6002_U1 ( .IN1(n4546), .IN2(U6002_n1), .QN(WX7349) );
  INVX0 U6003_U2 ( .INP(WX7284), .ZN(U6003_n1) );
  NOR2X0 U6003_U1 ( .IN1(n4546), .IN2(U6003_n1), .QN(WX7347) );
  INVX0 U6004_U2 ( .INP(WX7282), .ZN(U6004_n1) );
  NOR2X0 U6004_U1 ( .IN1(n4546), .IN2(U6004_n1), .QN(WX7345) );
  INVX0 U6005_U2 ( .INP(WX7280), .ZN(U6005_n1) );
  NOR2X0 U6005_U1 ( .IN1(n4546), .IN2(U6005_n1), .QN(WX7343) );
  INVX0 U6006_U2 ( .INP(WX7278), .ZN(U6006_n1) );
  NOR2X0 U6006_U1 ( .IN1(n4546), .IN2(U6006_n1), .QN(WX7341) );
  INVX0 U6007_U2 ( .INP(WX7276), .ZN(U6007_n1) );
  NOR2X0 U6007_U1 ( .IN1(n4546), .IN2(U6007_n1), .QN(WX7339) );
  INVX0 U6008_U2 ( .INP(WX7274), .ZN(U6008_n1) );
  NOR2X0 U6008_U1 ( .IN1(n4547), .IN2(U6008_n1), .QN(WX7337) );
  INVX0 U6009_U2 ( .INP(WX7272), .ZN(U6009_n1) );
  NOR2X0 U6009_U1 ( .IN1(n4547), .IN2(U6009_n1), .QN(WX7335) );
  INVX0 U6010_U2 ( .INP(WX7270), .ZN(U6010_n1) );
  NOR2X0 U6010_U1 ( .IN1(n4547), .IN2(U6010_n1), .QN(WX7333) );
  INVX0 U6011_U2 ( .INP(WX7268), .ZN(U6011_n1) );
  NOR2X0 U6011_U1 ( .IN1(n4547), .IN2(U6011_n1), .QN(WX7331) );
  INVX0 U6012_U2 ( .INP(WX7266), .ZN(U6012_n1) );
  NOR2X0 U6012_U1 ( .IN1(n4547), .IN2(U6012_n1), .QN(WX7329) );
  INVX0 U6013_U2 ( .INP(WX7264), .ZN(U6013_n1) );
  NOR2X0 U6013_U1 ( .IN1(n4547), .IN2(U6013_n1), .QN(WX7327) );
  INVX0 U6014_U2 ( .INP(WX7262), .ZN(U6014_n1) );
  NOR2X0 U6014_U1 ( .IN1(n4547), .IN2(U6014_n1), .QN(WX7325) );
  INVX0 U6015_U2 ( .INP(WX7260), .ZN(U6015_n1) );
  NOR2X0 U6015_U1 ( .IN1(n4547), .IN2(U6015_n1), .QN(WX7323) );
  INVX0 U6016_U2 ( .INP(WX7258), .ZN(U6016_n1) );
  NOR2X0 U6016_U1 ( .IN1(n4547), .IN2(U6016_n1), .QN(WX7321) );
  INVX0 U6017_U2 ( .INP(WX7256), .ZN(U6017_n1) );
  NOR2X0 U6017_U1 ( .IN1(n4547), .IN2(U6017_n1), .QN(WX7319) );
  INVX0 U6018_U2 ( .INP(test_so61), .ZN(U6018_n1) );
  NOR2X0 U6018_U1 ( .IN1(n4547), .IN2(U6018_n1), .QN(WX7317) );
  INVX0 U6019_U2 ( .INP(WX7252), .ZN(U6019_n1) );
  NOR2X0 U6019_U1 ( .IN1(n4547), .IN2(U6019_n1), .QN(WX7315) );
  INVX0 U6020_U2 ( .INP(WX7250), .ZN(U6020_n1) );
  NOR2X0 U6020_U1 ( .IN1(n4547), .IN2(U6020_n1), .QN(WX7313) );
  INVX0 U6021_U2 ( .INP(WX7248), .ZN(U6021_n1) );
  NOR2X0 U6021_U1 ( .IN1(n4548), .IN2(U6021_n1), .QN(WX7311) );
  INVX0 U6022_U2 ( .INP(WX7246), .ZN(U6022_n1) );
  NOR2X0 U6022_U1 ( .IN1(n4548), .IN2(U6022_n1), .QN(WX7309) );
  INVX0 U6023_U2 ( .INP(WX7244), .ZN(U6023_n1) );
  NOR2X0 U6023_U1 ( .IN1(n4548), .IN2(U6023_n1), .QN(WX7307) );
  INVX0 U6024_U2 ( .INP(WX7242), .ZN(U6024_n1) );
  NOR2X0 U6024_U1 ( .IN1(n4548), .IN2(U6024_n1), .QN(WX7305) );
  INVX0 U6025_U2 ( .INP(WX7240), .ZN(U6025_n1) );
  NOR2X0 U6025_U1 ( .IN1(n4549), .IN2(U6025_n1), .QN(WX7303) );
  INVX0 U6026_U2 ( .INP(WX7238), .ZN(U6026_n1) );
  NOR2X0 U6026_U1 ( .IN1(n4548), .IN2(U6026_n1), .QN(WX7301) );
  INVX0 U6027_U2 ( .INP(WX7236), .ZN(U6027_n1) );
  NOR2X0 U6027_U1 ( .IN1(n4549), .IN2(U6027_n1), .QN(WX7299) );
  INVX0 U6028_U2 ( .INP(WX7234), .ZN(U6028_n1) );
  NOR2X0 U6028_U1 ( .IN1(n4548), .IN2(U6028_n1), .QN(WX7297) );
  INVX0 U6029_U2 ( .INP(WX7232), .ZN(U6029_n1) );
  NOR2X0 U6029_U1 ( .IN1(n4549), .IN2(U6029_n1), .QN(WX7295) );
  INVX0 U6030_U2 ( .INP(WX7230), .ZN(U6030_n1) );
  NOR2X0 U6030_U1 ( .IN1(n4548), .IN2(U6030_n1), .QN(WX7293) );
  INVX0 U6031_U2 ( .INP(WX7228), .ZN(U6031_n1) );
  NOR2X0 U6031_U1 ( .IN1(n4549), .IN2(U6031_n1), .QN(WX7291) );
  INVX0 U6032_U2 ( .INP(WX7226), .ZN(U6032_n1) );
  NOR2X0 U6032_U1 ( .IN1(n4548), .IN2(U6032_n1), .QN(WX7289) );
  INVX0 U6033_U2 ( .INP(WX7224), .ZN(U6033_n1) );
  NOR2X0 U6033_U1 ( .IN1(n4549), .IN2(U6033_n1), .QN(WX7287) );
  INVX0 U6034_U2 ( .INP(WX7222), .ZN(U6034_n1) );
  NOR2X0 U6034_U1 ( .IN1(n4548), .IN2(U6034_n1), .QN(WX7285) );
  INVX0 U6035_U2 ( .INP(test_so60), .ZN(U6035_n1) );
  NOR2X0 U6035_U1 ( .IN1(n4548), .IN2(U6035_n1), .QN(WX7283) );
  INVX0 U6036_U2 ( .INP(WX7218), .ZN(U6036_n1) );
  NOR2X0 U6036_U1 ( .IN1(n4549), .IN2(U6036_n1), .QN(WX7281) );
  INVX0 U6037_U2 ( .INP(WX7216), .ZN(U6037_n1) );
  NOR2X0 U6037_U1 ( .IN1(n4549), .IN2(U6037_n1), .QN(WX7279) );
  INVX0 U6038_U2 ( .INP(WX7214), .ZN(U6038_n1) );
  NOR2X0 U6038_U1 ( .IN1(n4548), .IN2(U6038_n1), .QN(WX7277) );
  INVX0 U6039_U2 ( .INP(WX7212), .ZN(U6039_n1) );
  NOR2X0 U6039_U1 ( .IN1(n4549), .IN2(U6039_n1), .QN(WX7275) );
  INVX0 U6040_U2 ( .INP(WX7210), .ZN(U6040_n1) );
  NOR2X0 U6040_U1 ( .IN1(n4549), .IN2(U6040_n1), .QN(WX7273) );
  INVX0 U6041_U2 ( .INP(WX7208), .ZN(U6041_n1) );
  NOR2X0 U6041_U1 ( .IN1(n4549), .IN2(U6041_n1), .QN(WX7271) );
  INVX0 U6042_U2 ( .INP(WX7206), .ZN(U6042_n1) );
  NOR2X0 U6042_U1 ( .IN1(n4549), .IN2(U6042_n1), .QN(WX7269) );
  INVX0 U6043_U2 ( .INP(WX7204), .ZN(U6043_n1) );
  NOR2X0 U6043_U1 ( .IN1(n4550), .IN2(U6043_n1), .QN(WX7267) );
  INVX0 U6044_U2 ( .INP(WX7202), .ZN(U6044_n1) );
  NOR2X0 U6044_U1 ( .IN1(n4548), .IN2(U6044_n1), .QN(WX7265) );
  INVX0 U6045_U2 ( .INP(WX7200), .ZN(U6045_n1) );
  NOR2X0 U6045_U1 ( .IN1(n4550), .IN2(U6045_n1), .QN(WX7263) );
  INVX0 U6046_U2 ( .INP(WX7198), .ZN(U6046_n1) );
  NOR2X0 U6046_U1 ( .IN1(n4549), .IN2(U6046_n1), .QN(WX7261) );
  INVX0 U6047_U2 ( .INP(WX7196), .ZN(U6047_n1) );
  NOR2X0 U6047_U1 ( .IN1(n4550), .IN2(U6047_n1), .QN(WX7259) );
  INVX0 U6048_U2 ( .INP(WX7194), .ZN(U6048_n1) );
  NOR2X0 U6048_U1 ( .IN1(n4549), .IN2(U6048_n1), .QN(WX7257) );
  INVX0 U6049_U2 ( .INP(WX7192), .ZN(U6049_n1) );
  NOR2X0 U6049_U1 ( .IN1(n4550), .IN2(U6049_n1), .QN(WX7255) );
  INVX0 U6050_U2 ( .INP(WX7190), .ZN(U6050_n1) );
  NOR2X0 U6050_U1 ( .IN1(n4548), .IN2(U6050_n1), .QN(WX7253) );
  INVX0 U6051_U2 ( .INP(WX7188), .ZN(U6051_n1) );
  NOR2X0 U6051_U1 ( .IN1(n4537), .IN2(U6051_n1), .QN(WX7251) );
  INVX0 U6052_U2 ( .INP(test_so59), .ZN(U6052_n1) );
  NOR2X0 U6052_U1 ( .IN1(n4533), .IN2(U6052_n1), .QN(WX7249) );
  INVX0 U6053_U2 ( .INP(WX7184), .ZN(U6053_n1) );
  NOR2X0 U6053_U1 ( .IN1(n4533), .IN2(U6053_n1), .QN(WX7247) );
  INVX0 U6054_U2 ( .INP(WX7182), .ZN(U6054_n1) );
  NOR2X0 U6054_U1 ( .IN1(n4533), .IN2(U6054_n1), .QN(WX7245) );
  INVX0 U6055_U2 ( .INP(WX7180), .ZN(U6055_n1) );
  NOR2X0 U6055_U1 ( .IN1(n4533), .IN2(U6055_n1), .QN(WX7243) );
  INVX0 U6056_U2 ( .INP(WX7178), .ZN(U6056_n1) );
  NOR2X0 U6056_U1 ( .IN1(n4533), .IN2(U6056_n1), .QN(WX7241) );
  INVX0 U6057_U2 ( .INP(WX7176), .ZN(U6057_n1) );
  NOR2X0 U6057_U1 ( .IN1(n4533), .IN2(U6057_n1), .QN(WX7239) );
  INVX0 U6058_U2 ( .INP(WX7174), .ZN(U6058_n1) );
  NOR2X0 U6058_U1 ( .IN1(n4533), .IN2(U6058_n1), .QN(WX7237) );
  INVX0 U6059_U2 ( .INP(WX7172), .ZN(U6059_n1) );
  NOR2X0 U6059_U1 ( .IN1(n4533), .IN2(U6059_n1), .QN(WX7235) );
  INVX0 U6060_U2 ( .INP(WX7170), .ZN(U6060_n1) );
  NOR2X0 U6060_U1 ( .IN1(n4533), .IN2(U6060_n1), .QN(WX7233) );
  INVX0 U6061_U2 ( .INP(WX7168), .ZN(U6061_n1) );
  NOR2X0 U6061_U1 ( .IN1(n4533), .IN2(U6061_n1), .QN(WX7231) );
  INVX0 U6062_U2 ( .INP(WX7166), .ZN(U6062_n1) );
  NOR2X0 U6062_U1 ( .IN1(n4534), .IN2(U6062_n1), .QN(WX7229) );
  INVX0 U6063_U2 ( .INP(WX7164), .ZN(U6063_n1) );
  NOR2X0 U6063_U1 ( .IN1(n4534), .IN2(U6063_n1), .QN(WX7227) );
  INVX0 U6064_U2 ( .INP(WX7162), .ZN(U6064_n1) );
  NOR2X0 U6064_U1 ( .IN1(n4534), .IN2(U6064_n1), .QN(WX7225) );
  INVX0 U6065_U2 ( .INP(WX7160), .ZN(U6065_n1) );
  NOR2X0 U6065_U1 ( .IN1(n4534), .IN2(U6065_n1), .QN(WX7223) );
  INVX0 U6066_U2 ( .INP(WX7158), .ZN(U6066_n1) );
  NOR2X0 U6066_U1 ( .IN1(n4534), .IN2(U6066_n1), .QN(WX7221) );
  INVX0 U6067_U2 ( .INP(WX7156), .ZN(U6067_n1) );
  NOR2X0 U6067_U1 ( .IN1(n4534), .IN2(U6067_n1), .QN(WX7219) );
  INVX0 U6068_U2 ( .INP(WX7154), .ZN(U6068_n1) );
  NOR2X0 U6068_U1 ( .IN1(n4534), .IN2(U6068_n1), .QN(WX7217) );
  INVX0 U6069_U2 ( .INP(test_so58), .ZN(U6069_n1) );
  NOR2X0 U6069_U1 ( .IN1(n4534), .IN2(U6069_n1), .QN(WX7215) );
  INVX0 U6070_U2 ( .INP(WX7150), .ZN(U6070_n1) );
  NOR2X0 U6070_U1 ( .IN1(n4534), .IN2(U6070_n1), .QN(WX7213) );
  INVX0 U6071_U2 ( .INP(WX7148), .ZN(U6071_n1) );
  NOR2X0 U6071_U1 ( .IN1(n4534), .IN2(U6071_n1), .QN(WX7211) );
  INVX0 U6072_U2 ( .INP(WX7146), .ZN(U6072_n1) );
  NOR2X0 U6072_U1 ( .IN1(n4534), .IN2(U6072_n1), .QN(WX7209) );
  INVX0 U6073_U2 ( .INP(WX7144), .ZN(U6073_n1) );
  NOR2X0 U6073_U1 ( .IN1(n4534), .IN2(U6073_n1), .QN(WX7207) );
  INVX0 U6074_U2 ( .INP(WX7142), .ZN(U6074_n1) );
  NOR2X0 U6074_U1 ( .IN1(n4534), .IN2(U6074_n1), .QN(WX7205) );
  INVX0 U6075_U2 ( .INP(WX6007), .ZN(U6075_n1) );
  NOR2X0 U6075_U1 ( .IN1(n4535), .IN2(U6075_n1), .QN(WX6070) );
  INVX0 U6076_U2 ( .INP(test_so51), .ZN(U6076_n1) );
  NOR2X0 U6076_U1 ( .IN1(n4535), .IN2(U6076_n1), .QN(WX6068) );
  INVX0 U6077_U2 ( .INP(WX6003), .ZN(U6077_n1) );
  NOR2X0 U6077_U1 ( .IN1(n4535), .IN2(U6077_n1), .QN(WX6066) );
  INVX0 U6078_U2 ( .INP(WX6001), .ZN(U6078_n1) );
  NOR2X0 U6078_U1 ( .IN1(n4535), .IN2(U6078_n1), .QN(WX6064) );
  INVX0 U6079_U2 ( .INP(WX5999), .ZN(U6079_n1) );
  NOR2X0 U6079_U1 ( .IN1(n4535), .IN2(U6079_n1), .QN(WX6062) );
  INVX0 U6080_U2 ( .INP(WX5997), .ZN(U6080_n1) );
  NOR2X0 U6080_U1 ( .IN1(n4535), .IN2(U6080_n1), .QN(WX6060) );
  INVX0 U6081_U2 ( .INP(WX5995), .ZN(U6081_n1) );
  NOR2X0 U6081_U1 ( .IN1(n4535), .IN2(U6081_n1), .QN(WX6058) );
  INVX0 U6082_U2 ( .INP(WX5993), .ZN(U6082_n1) );
  NOR2X0 U6082_U1 ( .IN1(n4535), .IN2(U6082_n1), .QN(WX6056) );
  INVX0 U6083_U2 ( .INP(WX5991), .ZN(U6083_n1) );
  NOR2X0 U6083_U1 ( .IN1(n4535), .IN2(U6083_n1), .QN(WX6054) );
  INVX0 U6084_U2 ( .INP(WX5989), .ZN(U6084_n1) );
  NOR2X0 U6084_U1 ( .IN1(n4535), .IN2(U6084_n1), .QN(WX6052) );
  INVX0 U6085_U2 ( .INP(WX5987), .ZN(U6085_n1) );
  NOR2X0 U6085_U1 ( .IN1(n4535), .IN2(U6085_n1), .QN(WX6050) );
  INVX0 U6086_U2 ( .INP(WX5985), .ZN(U6086_n1) );
  NOR2X0 U6086_U1 ( .IN1(n4535), .IN2(U6086_n1), .QN(WX6048) );
  INVX0 U6087_U2 ( .INP(WX5983), .ZN(U6087_n1) );
  NOR2X0 U6087_U1 ( .IN1(n4535), .IN2(U6087_n1), .QN(WX6046) );
  INVX0 U6088_U2 ( .INP(WX5981), .ZN(U6088_n1) );
  NOR2X0 U6088_U1 ( .IN1(n4536), .IN2(U6088_n1), .QN(WX6044) );
  INVX0 U6089_U2 ( .INP(WX5979), .ZN(U6089_n1) );
  NOR2X0 U6089_U1 ( .IN1(n4536), .IN2(U6089_n1), .QN(WX6042) );
  INVX0 U6090_U2 ( .INP(WX5977), .ZN(U6090_n1) );
  NOR2X0 U6090_U1 ( .IN1(n4536), .IN2(U6090_n1), .QN(WX6040) );
  INVX0 U6091_U2 ( .INP(WX5975), .ZN(U6091_n1) );
  NOR2X0 U6091_U1 ( .IN1(n4536), .IN2(U6091_n1), .QN(WX6038) );
  INVX0 U6092_U2 ( .INP(WX5973), .ZN(U6092_n1) );
  NOR2X0 U6092_U1 ( .IN1(n4536), .IN2(U6092_n1), .QN(WX6036) );
  INVX0 U6093_U2 ( .INP(test_so50), .ZN(U6093_n1) );
  NOR2X0 U6093_U1 ( .IN1(n4536), .IN2(U6093_n1), .QN(WX6034) );
  INVX0 U6094_U2 ( .INP(WX5969), .ZN(U6094_n1) );
  NOR2X0 U6094_U1 ( .IN1(n4536), .IN2(U6094_n1), .QN(WX6032) );
  INVX0 U6095_U2 ( .INP(WX5967), .ZN(U6095_n1) );
  NOR2X0 U6095_U1 ( .IN1(n4536), .IN2(U6095_n1), .QN(WX6030) );
  INVX0 U6096_U2 ( .INP(WX5965), .ZN(U6096_n1) );
  NOR2X0 U6096_U1 ( .IN1(n4536), .IN2(U6096_n1), .QN(WX6028) );
  INVX0 U6097_U2 ( .INP(WX5963), .ZN(U6097_n1) );
  NOR2X0 U6097_U1 ( .IN1(n4536), .IN2(U6097_n1), .QN(WX6026) );
  INVX0 U6098_U2 ( .INP(WX5961), .ZN(U6098_n1) );
  NOR2X0 U6098_U1 ( .IN1(n4536), .IN2(U6098_n1), .QN(WX6024) );
  INVX0 U6099_U2 ( .INP(WX5959), .ZN(U6099_n1) );
  NOR2X0 U6099_U1 ( .IN1(n4536), .IN2(U6099_n1), .QN(WX6022) );
  INVX0 U6100_U2 ( .INP(WX5957), .ZN(U6100_n1) );
  NOR2X0 U6100_U1 ( .IN1(n4536), .IN2(U6100_n1), .QN(WX6020) );
  INVX0 U6101_U2 ( .INP(WX5955), .ZN(U6101_n1) );
  NOR2X0 U6101_U1 ( .IN1(n4537), .IN2(U6101_n1), .QN(WX6018) );
  INVX0 U6102_U2 ( .INP(WX5953), .ZN(U6102_n1) );
  NOR2X0 U6102_U1 ( .IN1(n4537), .IN2(U6102_n1), .QN(WX6016) );
  INVX0 U6103_U2 ( .INP(WX5951), .ZN(U6103_n1) );
  NOR2X0 U6103_U1 ( .IN1(n4537), .IN2(U6103_n1), .QN(WX6014) );
  INVX0 U6104_U2 ( .INP(WX5949), .ZN(U6104_n1) );
  NOR2X0 U6104_U1 ( .IN1(n4537), .IN2(U6104_n1), .QN(WX6012) );
  INVX0 U6105_U2 ( .INP(WX5947), .ZN(U6105_n1) );
  NOR2X0 U6105_U1 ( .IN1(n4537), .IN2(U6105_n1), .QN(WX6010) );
  INVX0 U6106_U2 ( .INP(WX5945), .ZN(U6106_n1) );
  NOR2X0 U6106_U1 ( .IN1(n4537), .IN2(U6106_n1), .QN(WX6008) );
  INVX0 U6107_U2 ( .INP(WX5943), .ZN(U6107_n1) );
  NOR2X0 U6107_U1 ( .IN1(n4537), .IN2(U6107_n1), .QN(WX6006) );
  INVX0 U6108_U2 ( .INP(WX5941), .ZN(U6108_n1) );
  NOR2X0 U6108_U1 ( .IN1(n4537), .IN2(U6108_n1), .QN(WX6004) );
  INVX0 U6109_U2 ( .INP(WX5929), .ZN(U6109_n1) );
  NOR2X0 U6109_U1 ( .IN1(n4537), .IN2(U6109_n1), .QN(WX5992) );
  INVX0 U6110_U2 ( .INP(WX5927), .ZN(U6110_n1) );
  NOR2X0 U6110_U1 ( .IN1(n4537), .IN2(U6110_n1), .QN(WX5990) );
  INVX0 U6111_U2 ( .INP(WX5925), .ZN(U6111_n1) );
  NOR2X0 U6111_U1 ( .IN1(n4537), .IN2(U6111_n1), .QN(WX5988) );
  INVX0 U6112_U2 ( .INP(WX5923), .ZN(U6112_n1) );
  NOR2X0 U6112_U1 ( .IN1(n4537), .IN2(U6112_n1), .QN(WX5986) );
  INVX0 U6113_U2 ( .INP(WX5921), .ZN(U6113_n1) );
  NOR2X0 U6113_U1 ( .IN1(n4538), .IN2(U6113_n1), .QN(WX5984) );
  INVX0 U6114_U2 ( .INP(WX5919), .ZN(U6114_n1) );
  NOR2X0 U6114_U1 ( .IN1(n4538), .IN2(U6114_n1), .QN(WX5982) );
  INVX0 U6115_U2 ( .INP(WX5917), .ZN(U6115_n1) );
  NOR2X0 U6115_U1 ( .IN1(n4538), .IN2(U6115_n1), .QN(WX5980) );
  INVX0 U6116_U2 ( .INP(WX5915), .ZN(U6116_n1) );
  NOR2X0 U6116_U1 ( .IN1(n4538), .IN2(U6116_n1), .QN(WX5978) );
  INVX0 U6117_U2 ( .INP(WX5913), .ZN(U6117_n1) );
  NOR2X0 U6117_U1 ( .IN1(n4538), .IN2(U6117_n1), .QN(WX5976) );
  INVX0 U6118_U2 ( .INP(WX5911), .ZN(U6118_n1) );
  NOR2X0 U6118_U1 ( .IN1(n4538), .IN2(U6118_n1), .QN(WX5974) );
  INVX0 U6119_U2 ( .INP(WX5909), .ZN(U6119_n1) );
  NOR2X0 U6119_U1 ( .IN1(n4538), .IN2(U6119_n1), .QN(WX5972) );
  INVX0 U6120_U2 ( .INP(WX5907), .ZN(U6120_n1) );
  NOR2X0 U6120_U1 ( .IN1(n4538), .IN2(U6120_n1), .QN(WX5970) );
  INVX0 U6121_U2 ( .INP(WX5905), .ZN(U6121_n1) );
  NOR2X0 U6121_U1 ( .IN1(n4538), .IN2(U6121_n1), .QN(WX5968) );
  INVX0 U6122_U2 ( .INP(test_so48), .ZN(U6122_n1) );
  NOR2X0 U6122_U1 ( .IN1(n4538), .IN2(U6122_n1), .QN(WX5966) );
  INVX0 U6123_U2 ( .INP(WX5901), .ZN(U6123_n1) );
  NOR2X0 U6123_U1 ( .IN1(n4538), .IN2(U6123_n1), .QN(WX5964) );
  INVX0 U6124_U2 ( .INP(WX5899), .ZN(U6124_n1) );
  NOR2X0 U6124_U1 ( .IN1(n4538), .IN2(U6124_n1), .QN(WX5962) );
  INVX0 U6125_U2 ( .INP(WX5897), .ZN(U6125_n1) );
  NOR2X0 U6125_U1 ( .IN1(n4538), .IN2(U6125_n1), .QN(WX5960) );
  INVX0 U6126_U2 ( .INP(WX5895), .ZN(U6126_n1) );
  NOR2X0 U6126_U1 ( .IN1(n4539), .IN2(U6126_n1), .QN(WX5958) );
  INVX0 U6127_U2 ( .INP(WX5893), .ZN(U6127_n1) );
  NOR2X0 U6127_U1 ( .IN1(n4539), .IN2(U6127_n1), .QN(WX5956) );
  INVX0 U6128_U2 ( .INP(WX5891), .ZN(U6128_n1) );
  NOR2X0 U6128_U1 ( .IN1(n4539), .IN2(U6128_n1), .QN(WX5954) );
  INVX0 U6129_U2 ( .INP(WX5889), .ZN(U6129_n1) );
  NOR2X0 U6129_U1 ( .IN1(n4539), .IN2(U6129_n1), .QN(WX5952) );
  INVX0 U6130_U2 ( .INP(WX5887), .ZN(U6130_n1) );
  NOR2X0 U6130_U1 ( .IN1(n4539), .IN2(U6130_n1), .QN(WX5950) );
  INVX0 U6131_U2 ( .INP(WX5885), .ZN(U6131_n1) );
  NOR2X0 U6131_U1 ( .IN1(n4539), .IN2(U6131_n1), .QN(WX5948) );
  INVX0 U6132_U2 ( .INP(WX5883), .ZN(U6132_n1) );
  NOR2X0 U6132_U1 ( .IN1(n4539), .IN2(U6132_n1), .QN(WX5946) );
  INVX0 U6133_U2 ( .INP(WX5881), .ZN(U6133_n1) );
  NOR2X0 U6133_U1 ( .IN1(n4539), .IN2(U6133_n1), .QN(WX5944) );
  INVX0 U6134_U2 ( .INP(WX5879), .ZN(U6134_n1) );
  NOR2X0 U6134_U1 ( .IN1(n4539), .IN2(U6134_n1), .QN(WX5942) );
  INVX0 U6135_U2 ( .INP(WX5877), .ZN(U6135_n1) );
  NOR2X0 U6135_U1 ( .IN1(n4539), .IN2(U6135_n1), .QN(WX5940) );
  INVX0 U6136_U2 ( .INP(WX5875), .ZN(U6136_n1) );
  NOR2X0 U6136_U1 ( .IN1(n4533), .IN2(U6136_n1), .QN(WX5938) );
  INVX0 U6137_U2 ( .INP(WX5873), .ZN(U6137_n1) );
  NOR2X0 U6137_U1 ( .IN1(n4541), .IN2(U6137_n1), .QN(WX5936) );
  INVX0 U6138_U2 ( .INP(WX5871), .ZN(U6138_n1) );
  NOR2X0 U6138_U1 ( .IN1(n4541), .IN2(U6138_n1), .QN(WX5934) );
  INVX0 U6139_U2 ( .INP(test_so47), .ZN(U6139_n1) );
  NOR2X0 U6139_U1 ( .IN1(n4541), .IN2(U6139_n1), .QN(WX5932) );
  INVX0 U6140_U2 ( .INP(WX5867), .ZN(U6140_n1) );
  NOR2X0 U6140_U1 ( .IN1(n4541), .IN2(U6140_n1), .QN(WX5930) );
  INVX0 U6141_U2 ( .INP(WX5865), .ZN(U6141_n1) );
  NOR2X0 U6141_U1 ( .IN1(n4541), .IN2(U6141_n1), .QN(WX5928) );
  INVX0 U6142_U2 ( .INP(WX5863), .ZN(U6142_n1) );
  NOR2X0 U6142_U1 ( .IN1(n4541), .IN2(U6142_n1), .QN(WX5926) );
  INVX0 U6143_U2 ( .INP(WX5861), .ZN(U6143_n1) );
  NOR2X0 U6143_U1 ( .IN1(n4541), .IN2(U6143_n1), .QN(WX5924) );
  INVX0 U6144_U2 ( .INP(WX5859), .ZN(U6144_n1) );
  NOR2X0 U6144_U1 ( .IN1(n4541), .IN2(U6144_n1), .QN(WX5922) );
  INVX0 U6145_U2 ( .INP(WX5857), .ZN(U6145_n1) );
  NOR2X0 U6145_U1 ( .IN1(n4541), .IN2(U6145_n1), .QN(WX5920) );
  INVX0 U6146_U2 ( .INP(WX5855), .ZN(U6146_n1) );
  NOR2X0 U6146_U1 ( .IN1(n4540), .IN2(U6146_n1), .QN(WX5918) );
  INVX0 U6147_U2 ( .INP(WX5853), .ZN(U6147_n1) );
  NOR2X0 U6147_U1 ( .IN1(n4540), .IN2(U6147_n1), .QN(WX5916) );
  INVX0 U6148_U2 ( .INP(WX5851), .ZN(U6148_n1) );
  NOR2X0 U6148_U1 ( .IN1(n4540), .IN2(U6148_n1), .QN(WX5914) );
  INVX0 U6149_U2 ( .INP(WX5849), .ZN(U6149_n1) );
  NOR2X0 U6149_U1 ( .IN1(n4540), .IN2(U6149_n1), .QN(WX5912) );
  INVX0 U6150_U2 ( .INP(WX4714), .ZN(U6150_n1) );
  NOR2X0 U6150_U1 ( .IN1(n4540), .IN2(U6150_n1), .QN(WX4777) );
  INVX0 U6151_U2 ( .INP(WX4712), .ZN(U6151_n1) );
  NOR2X0 U6151_U1 ( .IN1(n4540), .IN2(U6151_n1), .QN(WX4775) );
  INVX0 U6152_U2 ( .INP(WX4710), .ZN(U6152_n1) );
  NOR2X0 U6152_U1 ( .IN1(n4540), .IN2(U6152_n1), .QN(WX4773) );
  INVX0 U6153_U2 ( .INP(WX4708), .ZN(U6153_n1) );
  NOR2X0 U6153_U1 ( .IN1(n4540), .IN2(U6153_n1), .QN(WX4771) );
  INVX0 U6154_U2 ( .INP(WX4706), .ZN(U6154_n1) );
  NOR2X0 U6154_U1 ( .IN1(n4540), .IN2(U6154_n1), .QN(WX4769) );
  INVX0 U6155_U2 ( .INP(WX4704), .ZN(U6155_n1) );
  NOR2X0 U6155_U1 ( .IN1(n4540), .IN2(U6155_n1), .QN(WX4767) );
  INVX0 U6156_U2 ( .INP(WX4702), .ZN(U6156_n1) );
  NOR2X0 U6156_U1 ( .IN1(n4540), .IN2(U6156_n1), .QN(WX4765) );
  INVX0 U6157_U2 ( .INP(WX4700), .ZN(U6157_n1) );
  NOR2X0 U6157_U1 ( .IN1(n4540), .IN2(U6157_n1), .QN(WX4763) );
  INVX0 U6158_U2 ( .INP(WX4698), .ZN(U6158_n1) );
  NOR2X0 U6158_U1 ( .IN1(n4540), .IN2(U6158_n1), .QN(WX4761) );
  INVX0 U6159_U2 ( .INP(WX4696), .ZN(U6159_n1) );
  NOR2X0 U6159_U1 ( .IN1(n4539), .IN2(U6159_n1), .QN(WX4759) );
  INVX0 U6160_U2 ( .INP(WX4694), .ZN(U6160_n1) );
  NOR2X0 U6160_U1 ( .IN1(n4539), .IN2(U6160_n1), .QN(WX4757) );
  INVX0 U6161_U2 ( .INP(WX4692), .ZN(U6161_n1) );
  NOR2X0 U6161_U1 ( .IN1(n4539), .IN2(U6161_n1), .QN(WX4755) );
  INVX0 U6162_U2 ( .INP(WX4690), .ZN(U6162_n1) );
  NOR2X0 U6162_U1 ( .IN1(n4503), .IN2(U6162_n1), .QN(WX4753) );
  INVX0 U6163_U2 ( .INP(test_so39), .ZN(U6163_n1) );
  NOR2X0 U6163_U1 ( .IN1(n4503), .IN2(U6163_n1), .QN(WX4751) );
  INVX0 U6164_U2 ( .INP(WX4686), .ZN(U6164_n1) );
  NOR2X0 U6164_U1 ( .IN1(n4503), .IN2(U6164_n1), .QN(WX4749) );
  INVX0 U6165_U2 ( .INP(WX4684), .ZN(U6165_n1) );
  NOR2X0 U6165_U1 ( .IN1(n4503), .IN2(U6165_n1), .QN(WX4747) );
  INVX0 U6166_U2 ( .INP(WX4682), .ZN(U6166_n1) );
  NOR2X0 U6166_U1 ( .IN1(n4503), .IN2(U6166_n1), .QN(WX4745) );
  INVX0 U6167_U2 ( .INP(WX4680), .ZN(U6167_n1) );
  NOR2X0 U6167_U1 ( .IN1(n4503), .IN2(U6167_n1), .QN(WX4743) );
  INVX0 U6168_U2 ( .INP(WX4678), .ZN(U6168_n1) );
  NOR2X0 U6168_U1 ( .IN1(n4503), .IN2(U6168_n1), .QN(WX4741) );
  INVX0 U6169_U2 ( .INP(WX4676), .ZN(U6169_n1) );
  NOR2X0 U6169_U1 ( .IN1(n4503), .IN2(U6169_n1), .QN(WX4739) );
  INVX0 U6170_U2 ( .INP(WX4674), .ZN(U6170_n1) );
  NOR2X0 U6170_U1 ( .IN1(n4503), .IN2(U6170_n1), .QN(WX4737) );
  INVX0 U6171_U2 ( .INP(WX4672), .ZN(U6171_n1) );
  NOR2X0 U6171_U1 ( .IN1(n4502), .IN2(U6171_n1), .QN(WX4735) );
  INVX0 U6172_U2 ( .INP(WX4670), .ZN(U6172_n1) );
  NOR2X0 U6172_U1 ( .IN1(n4502), .IN2(U6172_n1), .QN(WX4733) );
  INVX0 U6173_U2 ( .INP(WX4668), .ZN(U6173_n1) );
  NOR2X0 U6173_U1 ( .IN1(n4502), .IN2(U6173_n1), .QN(WX4731) );
  INVX0 U6174_U2 ( .INP(WX4666), .ZN(U6174_n1) );
  NOR2X0 U6174_U1 ( .IN1(n4502), .IN2(U6174_n1), .QN(WX4729) );
  INVX0 U6175_U2 ( .INP(WX4664), .ZN(U6175_n1) );
  NOR2X0 U6175_U1 ( .IN1(n4502), .IN2(U6175_n1), .QN(WX4727) );
  INVX0 U6176_U2 ( .INP(WX4662), .ZN(U6176_n1) );
  NOR2X0 U6176_U1 ( .IN1(n4502), .IN2(U6176_n1), .QN(WX4725) );
  INVX0 U6177_U2 ( .INP(WX4660), .ZN(U6177_n1) );
  NOR2X0 U6177_U1 ( .IN1(n4502), .IN2(U6177_n1), .QN(WX4723) );
  INVX0 U6178_U2 ( .INP(WX4658), .ZN(U6178_n1) );
  NOR2X0 U6178_U1 ( .IN1(n4502), .IN2(U6178_n1), .QN(WX4721) );
  INVX0 U6179_U2 ( .INP(WX4656), .ZN(U6179_n1) );
  NOR2X0 U6179_U1 ( .IN1(n4502), .IN2(U6179_n1), .QN(WX4719) );
  INVX0 U6180_U2 ( .INP(test_so38), .ZN(U6180_n1) );
  NOR2X0 U6180_U1 ( .IN1(n4502), .IN2(U6180_n1), .QN(WX4717) );
  INVX0 U6181_U2 ( .INP(WX4652), .ZN(U6181_n1) );
  NOR2X0 U6181_U1 ( .IN1(n4502), .IN2(U6181_n1), .QN(WX4715) );
  INVX0 U6182_U2 ( .INP(WX4650), .ZN(U6182_n1) );
  NOR2X0 U6182_U1 ( .IN1(n4502), .IN2(U6182_n1), .QN(WX4713) );
  INVX0 U6183_U2 ( .INP(WX4648), .ZN(U6183_n1) );
  NOR2X0 U6183_U1 ( .IN1(n4502), .IN2(U6183_n1), .QN(WX4711) );
  INVX0 U6184_U2 ( .INP(WX4646), .ZN(U6184_n1) );
  NOR2X0 U6184_U1 ( .IN1(n4501), .IN2(U6184_n1), .QN(WX4709) );
  INVX0 U6185_U2 ( .INP(WX4644), .ZN(U6185_n1) );
  NOR2X0 U6185_U1 ( .IN1(n4501), .IN2(U6185_n1), .QN(WX4707) );
  INVX0 U6186_U2 ( .INP(WX4642), .ZN(U6186_n1) );
  NOR2X0 U6186_U1 ( .IN1(n4501), .IN2(U6186_n1), .QN(WX4705) );
  INVX0 U6187_U2 ( .INP(WX4640), .ZN(U6187_n1) );
  NOR2X0 U6187_U1 ( .IN1(n4501), .IN2(U6187_n1), .QN(WX4703) );
  INVX0 U6188_U2 ( .INP(WX4638), .ZN(U6188_n1) );
  NOR2X0 U6188_U1 ( .IN1(n4501), .IN2(U6188_n1), .QN(WX4701) );
  INVX0 U6189_U2 ( .INP(WX4636), .ZN(U6189_n1) );
  NOR2X0 U6189_U1 ( .IN1(n4501), .IN2(U6189_n1), .QN(WX4699) );
  INVX0 U6190_U2 ( .INP(WX4634), .ZN(U6190_n1) );
  NOR2X0 U6190_U1 ( .IN1(n4501), .IN2(U6190_n1), .QN(WX4697) );
  INVX0 U6191_U2 ( .INP(WX4632), .ZN(U6191_n1) );
  NOR2X0 U6191_U1 ( .IN1(n4501), .IN2(U6191_n1), .QN(WX4695) );
  INVX0 U6192_U2 ( .INP(WX4630), .ZN(U6192_n1) );
  NOR2X0 U6192_U1 ( .IN1(n4501), .IN2(U6192_n1), .QN(WX4693) );
  INVX0 U6193_U2 ( .INP(WX4628), .ZN(U6193_n1) );
  NOR2X0 U6193_U1 ( .IN1(n4501), .IN2(U6193_n1), .QN(WX4691) );
  INVX0 U6194_U2 ( .INP(WX4626), .ZN(U6194_n1) );
  NOR2X0 U6194_U1 ( .IN1(n4501), .IN2(U6194_n1), .QN(WX4689) );
  INVX0 U6195_U2 ( .INP(WX4624), .ZN(U6195_n1) );
  NOR2X0 U6195_U1 ( .IN1(n4501), .IN2(U6195_n1), .QN(WX4687) );
  INVX0 U6196_U2 ( .INP(WX4622), .ZN(U6196_n1) );
  NOR2X0 U6196_U1 ( .IN1(n4501), .IN2(U6196_n1), .QN(WX4685) );
  INVX0 U6197_U2 ( .INP(test_so37), .ZN(U6197_n1) );
  NOR2X0 U6197_U1 ( .IN1(n4500), .IN2(U6197_n1), .QN(WX4683) );
  INVX0 U6198_U2 ( .INP(WX4618), .ZN(U6198_n1) );
  NOR2X0 U6198_U1 ( .IN1(n4500), .IN2(U6198_n1), .QN(WX4681) );
  INVX0 U6199_U2 ( .INP(WX4616), .ZN(U6199_n1) );
  NOR2X0 U6199_U1 ( .IN1(n4500), .IN2(U6199_n1), .QN(WX4679) );
  INVX0 U6200_U2 ( .INP(WX4614), .ZN(U6200_n1) );
  NOR2X0 U6200_U1 ( .IN1(n4500), .IN2(U6200_n1), .QN(WX4677) );
  INVX0 U6201_U2 ( .INP(WX4612), .ZN(U6201_n1) );
  NOR2X0 U6201_U1 ( .IN1(n4500), .IN2(U6201_n1), .QN(WX4675) );
  INVX0 U6202_U2 ( .INP(WX4610), .ZN(U6202_n1) );
  NOR2X0 U6202_U1 ( .IN1(n4500), .IN2(U6202_n1), .QN(WX4673) );
  INVX0 U6203_U2 ( .INP(WX4608), .ZN(U6203_n1) );
  NOR2X0 U6203_U1 ( .IN1(n4500), .IN2(U6203_n1), .QN(WX4671) );
  INVX0 U6204_U2 ( .INP(WX4606), .ZN(U6204_n1) );
  NOR2X0 U6204_U1 ( .IN1(n4500), .IN2(U6204_n1), .QN(WX4669) );
  INVX0 U6205_U2 ( .INP(WX4604), .ZN(U6205_n1) );
  NOR2X0 U6205_U1 ( .IN1(n4500), .IN2(U6205_n1), .QN(WX4667) );
  INVX0 U6206_U2 ( .INP(WX4602), .ZN(U6206_n1) );
  NOR2X0 U6206_U1 ( .IN1(n4500), .IN2(U6206_n1), .QN(WX4665) );
  INVX0 U6207_U2 ( .INP(WX4600), .ZN(U6207_n1) );
  NOR2X0 U6207_U1 ( .IN1(n4500), .IN2(U6207_n1), .QN(WX4663) );
  INVX0 U6208_U2 ( .INP(WX4598), .ZN(U6208_n1) );
  NOR2X0 U6208_U1 ( .IN1(n4500), .IN2(U6208_n1), .QN(WX4661) );
  INVX0 U6209_U2 ( .INP(WX4596), .ZN(U6209_n1) );
  NOR2X0 U6209_U1 ( .IN1(n4500), .IN2(U6209_n1), .QN(WX4659) );
  INVX0 U6210_U2 ( .INP(WX4594), .ZN(U6210_n1) );
  NOR2X0 U6210_U1 ( .IN1(n4499), .IN2(U6210_n1), .QN(WX4657) );
  INVX0 U6211_U2 ( .INP(WX4592), .ZN(U6211_n1) );
  NOR2X0 U6211_U1 ( .IN1(n4499), .IN2(U6211_n1), .QN(WX4655) );
  INVX0 U6212_U2 ( .INP(WX4590), .ZN(U6212_n1) );
  NOR2X0 U6212_U1 ( .IN1(n4499), .IN2(U6212_n1), .QN(WX4653) );
  INVX0 U6213_U2 ( .INP(WX4588), .ZN(U6213_n1) );
  NOR2X0 U6213_U1 ( .IN1(n4499), .IN2(U6213_n1), .QN(WX4651) );
  INVX0 U6214_U2 ( .INP(test_so36), .ZN(U6214_n1) );
  NOR2X0 U6214_U1 ( .IN1(n4499), .IN2(U6214_n1), .QN(WX4649) );
  INVX0 U6215_U2 ( .INP(WX4584), .ZN(U6215_n1) );
  NOR2X0 U6215_U1 ( .IN1(n4499), .IN2(U6215_n1), .QN(WX4647) );
  INVX0 U6216_U2 ( .INP(WX4582), .ZN(U6216_n1) );
  NOR2X0 U6216_U1 ( .IN1(n4499), .IN2(U6216_n1), .QN(WX4645) );
  INVX0 U6217_U2 ( .INP(WX4580), .ZN(U6217_n1) );
  NOR2X0 U6217_U1 ( .IN1(n4499), .IN2(U6217_n1), .QN(WX4643) );
  INVX0 U6218_U2 ( .INP(WX4578), .ZN(U6218_n1) );
  NOR2X0 U6218_U1 ( .IN1(n4499), .IN2(U6218_n1), .QN(WX4641) );
  INVX0 U6219_U2 ( .INP(WX4576), .ZN(U6219_n1) );
  NOR2X0 U6219_U1 ( .IN1(n4499), .IN2(U6219_n1), .QN(WX4639) );
  INVX0 U6220_U2 ( .INP(WX4574), .ZN(U6220_n1) );
  NOR2X0 U6220_U1 ( .IN1(n4499), .IN2(U6220_n1), .QN(WX4637) );
  INVX0 U6221_U2 ( .INP(WX4572), .ZN(U6221_n1) );
  NOR2X0 U6221_U1 ( .IN1(n4499), .IN2(U6221_n1), .QN(WX4635) );
  INVX0 U6222_U2 ( .INP(WX4570), .ZN(U6222_n1) );
  NOR2X0 U6222_U1 ( .IN1(n4499), .IN2(U6222_n1), .QN(WX4633) );
  INVX0 U6223_U2 ( .INP(WX4568), .ZN(U6223_n1) );
  NOR2X0 U6223_U1 ( .IN1(n4498), .IN2(U6223_n1), .QN(WX4631) );
  INVX0 U6224_U2 ( .INP(WX4566), .ZN(U6224_n1) );
  NOR2X0 U6224_U1 ( .IN1(n4498), .IN2(U6224_n1), .QN(WX4629) );
  INVX0 U6225_U2 ( .INP(WX4564), .ZN(U6225_n1) );
  NOR2X0 U6225_U1 ( .IN1(n4498), .IN2(U6225_n1), .QN(WX4627) );
  INVX0 U6226_U2 ( .INP(WX4562), .ZN(U6226_n1) );
  NOR2X0 U6226_U1 ( .IN1(n4498), .IN2(U6226_n1), .QN(WX4625) );
  INVX0 U6227_U2 ( .INP(WX4560), .ZN(U6227_n1) );
  NOR2X0 U6227_U1 ( .IN1(n4498), .IN2(U6227_n1), .QN(WX4623) );
  INVX0 U6228_U2 ( .INP(WX4558), .ZN(U6228_n1) );
  NOR2X0 U6228_U1 ( .IN1(n4498), .IN2(U6228_n1), .QN(WX4621) );
  INVX0 U6229_U2 ( .INP(WX4556), .ZN(U6229_n1) );
  NOR2X0 U6229_U1 ( .IN1(n4498), .IN2(U6229_n1), .QN(WX4619) );
  INVX0 U6230_U2 ( .INP(WX3421), .ZN(U6230_n1) );
  NOR2X0 U6230_U1 ( .IN1(n4498), .IN2(U6230_n1), .QN(WX3484) );
  INVX0 U6231_U2 ( .INP(WX3419), .ZN(U6231_n1) );
  NOR2X0 U6231_U1 ( .IN1(n4498), .IN2(U6231_n1), .QN(WX3482) );
  INVX0 U6232_U2 ( .INP(WX3417), .ZN(U6232_n1) );
  NOR2X0 U6232_U1 ( .IN1(n4498), .IN2(U6232_n1), .QN(WX3480) );
  INVX0 U6233_U2 ( .INP(WX3415), .ZN(U6233_n1) );
  NOR2X0 U6233_U1 ( .IN1(n4498), .IN2(U6233_n1), .QN(WX3478) );
  INVX0 U6234_U2 ( .INP(WX3413), .ZN(U6234_n1) );
  NOR2X0 U6234_U1 ( .IN1(n4498), .IN2(U6234_n1), .QN(WX3476) );
  INVX0 U6235_U2 ( .INP(WX3411), .ZN(U6235_n1) );
  NOR2X0 U6235_U1 ( .IN1(n4498), .IN2(U6235_n1), .QN(WX3474) );
  INVX0 U6236_U2 ( .INP(WX3409), .ZN(U6236_n1) );
  NOR2X0 U6236_U1 ( .IN1(n4497), .IN2(U6236_n1), .QN(WX3472) );
  INVX0 U6237_U2 ( .INP(WX3407), .ZN(U6237_n1) );
  NOR2X0 U6237_U1 ( .IN1(n4497), .IN2(U6237_n1), .QN(WX3470) );
  INVX0 U6238_U2 ( .INP(test_so28), .ZN(U6238_n1) );
  NOR2X0 U6238_U1 ( .IN1(n4497), .IN2(U6238_n1), .QN(WX3468) );
  INVX0 U6239_U2 ( .INP(WX3403), .ZN(U6239_n1) );
  NOR2X0 U6239_U1 ( .IN1(n4497), .IN2(U6239_n1), .QN(WX3466) );
  INVX0 U6240_U2 ( .INP(WX3401), .ZN(U6240_n1) );
  NOR2X0 U6240_U1 ( .IN1(n4497), .IN2(U6240_n1), .QN(WX3464) );
  INVX0 U6241_U2 ( .INP(WX3399), .ZN(U6241_n1) );
  NOR2X0 U6241_U1 ( .IN1(n4497), .IN2(U6241_n1), .QN(WX3462) );
  INVX0 U6242_U2 ( .INP(WX3397), .ZN(U6242_n1) );
  NOR2X0 U6242_U1 ( .IN1(n4497), .IN2(U6242_n1), .QN(WX3460) );
  INVX0 U6243_U2 ( .INP(WX3395), .ZN(U6243_n1) );
  NOR2X0 U6243_U1 ( .IN1(n4491), .IN2(U6243_n1), .QN(WX3458) );
  INVX0 U6244_U2 ( .INP(WX3393), .ZN(U6244_n1) );
  NOR2X0 U6244_U1 ( .IN1(n4491), .IN2(U6244_n1), .QN(WX3456) );
  INVX0 U6245_U2 ( .INP(WX3391), .ZN(U6245_n1) );
  NOR2X0 U6245_U1 ( .IN1(n4491), .IN2(U6245_n1), .QN(WX3454) );
  INVX0 U6246_U2 ( .INP(WX3389), .ZN(U6246_n1) );
  NOR2X0 U6246_U1 ( .IN1(n4491), .IN2(U6246_n1), .QN(WX3452) );
  INVX0 U6247_U2 ( .INP(WX3387), .ZN(U6247_n1) );
  NOR2X0 U6247_U1 ( .IN1(n4491), .IN2(U6247_n1), .QN(WX3450) );
  INVX0 U6248_U2 ( .INP(WX3385), .ZN(U6248_n1) );
  NOR2X0 U6248_U1 ( .IN1(n4491), .IN2(U6248_n1), .QN(WX3448) );
  INVX0 U6249_U2 ( .INP(WX3383), .ZN(U6249_n1) );
  NOR2X0 U6249_U1 ( .IN1(n4491), .IN2(U6249_n1), .QN(WX3446) );
  INVX0 U6250_U2 ( .INP(WX3381), .ZN(U6250_n1) );
  NOR2X0 U6250_U1 ( .IN1(n4491), .IN2(U6250_n1), .QN(WX3444) );
  INVX0 U6251_U2 ( .INP(WX3379), .ZN(U6251_n1) );
  NOR2X0 U6251_U1 ( .IN1(n4491), .IN2(U6251_n1), .QN(WX3442) );
  INVX0 U6252_U2 ( .INP(WX3377), .ZN(U6252_n1) );
  NOR2X0 U6252_U1 ( .IN1(n4492), .IN2(U6252_n1), .QN(WX3440) );
  INVX0 U6253_U2 ( .INP(WX3375), .ZN(U6253_n1) );
  NOR2X0 U6253_U1 ( .IN1(n4491), .IN2(U6253_n1), .QN(WX3438) );
  INVX0 U6254_U2 ( .INP(WX3373), .ZN(U6254_n1) );
  NOR2X0 U6254_U1 ( .IN1(n4492), .IN2(U6254_n1), .QN(WX3436) );
  INVX0 U6255_U2 ( .INP(WX3371), .ZN(U6255_n1) );
  NOR2X0 U6255_U1 ( .IN1(n4492), .IN2(U6255_n1), .QN(WX3434) );
  INVX0 U6256_U2 ( .INP(test_so27), .ZN(U6256_n1) );
  NOR2X0 U6256_U1 ( .IN1(n4492), .IN2(U6256_n1), .QN(WX3432) );
  INVX0 U6257_U2 ( .INP(WX3367), .ZN(U6257_n1) );
  NOR2X0 U6257_U1 ( .IN1(n4492), .IN2(U6257_n1), .QN(WX3430) );
  INVX0 U6258_U2 ( .INP(WX3365), .ZN(U6258_n1) );
  NOR2X0 U6258_U1 ( .IN1(n4492), .IN2(U6258_n1), .QN(WX3428) );
  INVX0 U6259_U2 ( .INP(WX3363), .ZN(U6259_n1) );
  NOR2X0 U6259_U1 ( .IN1(n4492), .IN2(U6259_n1), .QN(WX3426) );
  INVX0 U6260_U2 ( .INP(WX3361), .ZN(U6260_n1) );
  NOR2X0 U6260_U1 ( .IN1(n4492), .IN2(U6260_n1), .QN(WX3424) );
  INVX0 U6261_U2 ( .INP(WX3359), .ZN(U6261_n1) );
  NOR2X0 U6261_U1 ( .IN1(n4492), .IN2(U6261_n1), .QN(WX3422) );
  INVX0 U6262_U2 ( .INP(WX3357), .ZN(U6262_n1) );
  NOR2X0 U6262_U1 ( .IN1(n4493), .IN2(U6262_n1), .QN(WX3420) );
  INVX0 U6263_U2 ( .INP(WX3355), .ZN(U6263_n1) );
  NOR2X0 U6263_U1 ( .IN1(n4492), .IN2(U6263_n1), .QN(WX3418) );
  INVX0 U6264_U2 ( .INP(WX3353), .ZN(U6264_n1) );
  NOR2X0 U6264_U1 ( .IN1(n4492), .IN2(U6264_n1), .QN(WX3416) );
  INVX0 U6265_U2 ( .INP(WX3351), .ZN(U6265_n1) );
  NOR2X0 U6265_U1 ( .IN1(n4492), .IN2(U6265_n1), .QN(WX3414) );
  INVX0 U6266_U2 ( .INP(WX3349), .ZN(U6266_n1) );
  NOR2X0 U6266_U1 ( .IN1(n4492), .IN2(U6266_n1), .QN(WX3412) );
  INVX0 U6267_U2 ( .INP(WX3347), .ZN(U6267_n1) );
  NOR2X0 U6267_U1 ( .IN1(n4493), .IN2(U6267_n1), .QN(WX3410) );
  INVX0 U6268_U2 ( .INP(WX3345), .ZN(U6268_n1) );
  NOR2X0 U6268_U1 ( .IN1(n4493), .IN2(U6268_n1), .QN(WX3408) );
  INVX0 U6269_U2 ( .INP(WX3343), .ZN(U6269_n1) );
  NOR2X0 U6269_U1 ( .IN1(n4493), .IN2(U6269_n1), .QN(WX3406) );
  INVX0 U6270_U2 ( .INP(WX3341), .ZN(U6270_n1) );
  NOR2X0 U6270_U1 ( .IN1(n4493), .IN2(U6270_n1), .QN(WX3404) );
  INVX0 U6271_U2 ( .INP(WX3339), .ZN(U6271_n1) );
  NOR2X0 U6271_U1 ( .IN1(n4493), .IN2(U6271_n1), .QN(WX3402) );
  INVX0 U6272_U2 ( .INP(WX3337), .ZN(U6272_n1) );
  NOR2X0 U6272_U1 ( .IN1(n4493), .IN2(U6272_n1), .QN(WX3400) );
  INVX0 U6273_U2 ( .INP(WX3335), .ZN(U6273_n1) );
  NOR2X0 U6273_U1 ( .IN1(n4493), .IN2(U6273_n1), .QN(WX3398) );
  INVX0 U6274_U2 ( .INP(test_so26), .ZN(U6274_n1) );
  NOR2X0 U6274_U1 ( .IN1(n4493), .IN2(U6274_n1), .QN(WX3396) );
  INVX0 U6275_U2 ( .INP(WX3331), .ZN(U6275_n1) );
  NOR2X0 U6275_U1 ( .IN1(n4493), .IN2(U6275_n1), .QN(WX3394) );
  INVX0 U6276_U2 ( .INP(WX3329), .ZN(U6276_n1) );
  NOR2X0 U6276_U1 ( .IN1(n4493), .IN2(U6276_n1), .QN(WX3392) );
  INVX0 U6277_U2 ( .INP(WX3327), .ZN(U6277_n1) );
  NOR2X0 U6277_U1 ( .IN1(n4494), .IN2(U6277_n1), .QN(WX3390) );
  INVX0 U6278_U2 ( .INP(WX3325), .ZN(U6278_n1) );
  NOR2X0 U6278_U1 ( .IN1(n4493), .IN2(U6278_n1), .QN(WX3388) );
  INVX0 U6279_U2 ( .INP(WX3323), .ZN(U6279_n1) );
  NOR2X0 U6279_U1 ( .IN1(n4493), .IN2(U6279_n1), .QN(WX3386) );
  INVX0 U6280_U2 ( .INP(WX3321), .ZN(U6280_n1) );
  NOR2X0 U6280_U1 ( .IN1(n4494), .IN2(U6280_n1), .QN(WX3384) );
  INVX0 U6281_U2 ( .INP(WX3319), .ZN(U6281_n1) );
  NOR2X0 U6281_U1 ( .IN1(n4494), .IN2(U6281_n1), .QN(WX3382) );
  INVX0 U6282_U2 ( .INP(WX3317), .ZN(U6282_n1) );
  NOR2X0 U6282_U1 ( .IN1(n4494), .IN2(U6282_n1), .QN(WX3380) );
  INVX0 U6283_U2 ( .INP(WX3315), .ZN(U6283_n1) );
  NOR2X0 U6283_U1 ( .IN1(n4494), .IN2(U6283_n1), .QN(WX3378) );
  INVX0 U6284_U2 ( .INP(WX3313), .ZN(U6284_n1) );
  NOR2X0 U6284_U1 ( .IN1(n4494), .IN2(U6284_n1), .QN(WX3376) );
  INVX0 U6285_U2 ( .INP(WX3311), .ZN(U6285_n1) );
  NOR2X0 U6285_U1 ( .IN1(n4494), .IN2(U6285_n1), .QN(WX3374) );
  INVX0 U6286_U2 ( .INP(WX3309), .ZN(U6286_n1) );
  NOR2X0 U6286_U1 ( .IN1(n4494), .IN2(U6286_n1), .QN(WX3372) );
  INVX0 U6287_U2 ( .INP(WX3307), .ZN(U6287_n1) );
  NOR2X0 U6287_U1 ( .IN1(n4494), .IN2(U6287_n1), .QN(WX3370) );
  INVX0 U6288_U2 ( .INP(WX3305), .ZN(U6288_n1) );
  NOR2X0 U6288_U1 ( .IN1(n4494), .IN2(U6288_n1), .QN(WX3368) );
  INVX0 U6289_U2 ( .INP(WX3303), .ZN(U6289_n1) );
  NOR2X0 U6289_U1 ( .IN1(n4494), .IN2(U6289_n1), .QN(WX3366) );
  INVX0 U6290_U2 ( .INP(WX3301), .ZN(U6290_n1) );
  NOR2X0 U6290_U1 ( .IN1(n4494), .IN2(U6290_n1), .QN(WX3364) );
  INVX0 U6291_U2 ( .INP(WX3299), .ZN(U6291_n1) );
  NOR2X0 U6291_U1 ( .IN1(n4494), .IN2(U6291_n1), .QN(WX3362) );
  INVX0 U6292_U2 ( .INP(test_so25), .ZN(U6292_n1) );
  NOR2X0 U6292_U1 ( .IN1(n4495), .IN2(U6292_n1), .QN(WX3360) );
  INVX0 U6293_U2 ( .INP(WX3295), .ZN(U6293_n1) );
  NOR2X0 U6293_U1 ( .IN1(n4495), .IN2(U6293_n1), .QN(WX3358) );
  INVX0 U6294_U2 ( .INP(WX3293), .ZN(U6294_n1) );
  NOR2X0 U6294_U1 ( .IN1(n4495), .IN2(U6294_n1), .QN(WX3356) );
  INVX0 U6295_U2 ( .INP(WX3291), .ZN(U6295_n1) );
  NOR2X0 U6295_U1 ( .IN1(n4495), .IN2(U6295_n1), .QN(WX3354) );
  INVX0 U6296_U2 ( .INP(WX3289), .ZN(U6296_n1) );
  NOR2X0 U6296_U1 ( .IN1(n4495), .IN2(U6296_n1), .QN(WX3352) );
  INVX0 U6297_U2 ( .INP(WX3287), .ZN(U6297_n1) );
  NOR2X0 U6297_U1 ( .IN1(n4495), .IN2(U6297_n1), .QN(WX3350) );
  INVX0 U6298_U2 ( .INP(WX3285), .ZN(U6298_n1) );
  NOR2X0 U6298_U1 ( .IN1(n4495), .IN2(U6298_n1), .QN(WX3348) );
  INVX0 U6299_U2 ( .INP(WX3283), .ZN(U6299_n1) );
  NOR2X0 U6299_U1 ( .IN1(n4495), .IN2(U6299_n1), .QN(WX3346) );
  INVX0 U6300_U2 ( .INP(WX3281), .ZN(U6300_n1) );
  NOR2X0 U6300_U1 ( .IN1(n4495), .IN2(U6300_n1), .QN(WX3344) );
  INVX0 U6301_U2 ( .INP(WX3279), .ZN(U6301_n1) );
  NOR2X0 U6301_U1 ( .IN1(n4495), .IN2(U6301_n1), .QN(WX3342) );
  INVX0 U6302_U2 ( .INP(WX3277), .ZN(U6302_n1) );
  NOR2X0 U6302_U1 ( .IN1(n4495), .IN2(U6302_n1), .QN(WX3340) );
  INVX0 U6303_U2 ( .INP(WX3275), .ZN(U6303_n1) );
  NOR2X0 U6303_U1 ( .IN1(n4495), .IN2(U6303_n1), .QN(WX3338) );
  INVX0 U6304_U2 ( .INP(WX3273), .ZN(U6304_n1) );
  NOR2X0 U6304_U1 ( .IN1(n4495), .IN2(U6304_n1), .QN(WX3336) );
  INVX0 U6305_U2 ( .INP(WX3271), .ZN(U6305_n1) );
  NOR2X0 U6305_U1 ( .IN1(n4496), .IN2(U6305_n1), .QN(WX3334) );
  INVX0 U6306_U2 ( .INP(WX3267), .ZN(U6306_n1) );
  NOR2X0 U6306_U1 ( .IN1(n4496), .IN2(U6306_n1), .QN(WX3330) );
  INVX0 U6307_U2 ( .INP(WX2128), .ZN(U6307_n1) );
  NOR2X0 U6307_U1 ( .IN1(n4496), .IN2(U6307_n1), .QN(WX2191) );
  INVX0 U6308_U2 ( .INP(WX2126), .ZN(U6308_n1) );
  NOR2X0 U6308_U1 ( .IN1(n4496), .IN2(U6308_n1), .QN(WX2189) );
  INVX0 U6309_U2 ( .INP(WX2124), .ZN(U6309_n1) );
  NOR2X0 U6309_U1 ( .IN1(n4496), .IN2(U6309_n1), .QN(WX2187) );
  INVX0 U6310_U2 ( .INP(WX2122), .ZN(U6310_n1) );
  NOR2X0 U6310_U1 ( .IN1(n4496), .IN2(U6310_n1), .QN(WX2185) );
  INVX0 U6311_U2 ( .INP(WX2120), .ZN(U6311_n1) );
  NOR2X0 U6311_U1 ( .IN1(n4496), .IN2(U6311_n1), .QN(WX2183) );
  INVX0 U6312_U2 ( .INP(WX2118), .ZN(U6312_n1) );
  NOR2X0 U6312_U1 ( .IN1(n4496), .IN2(U6312_n1), .QN(WX2181) );
  INVX0 U6313_U2 ( .INP(WX2116), .ZN(U6313_n1) );
  NOR2X0 U6313_U1 ( .IN1(n4496), .IN2(U6313_n1), .QN(WX2179) );
  INVX0 U6314_U2 ( .INP(WX2114), .ZN(U6314_n1) );
  NOR2X0 U6314_U1 ( .IN1(n4496), .IN2(U6314_n1), .QN(WX2177) );
  INVX0 U6315_U2 ( .INP(WX2112), .ZN(U6315_n1) );
  NOR2X0 U6315_U1 ( .IN1(n4496), .IN2(U6315_n1), .QN(WX2175) );
  INVX0 U6316_U2 ( .INP(WX2110), .ZN(U6316_n1) );
  NOR2X0 U6316_U1 ( .IN1(n4496), .IN2(U6316_n1), .QN(WX2173) );
  INVX0 U6317_U2 ( .INP(WX2108), .ZN(U6317_n1) );
  NOR2X0 U6317_U1 ( .IN1(n4496), .IN2(U6317_n1), .QN(WX2171) );
  INVX0 U6318_U2 ( .INP(WX2106), .ZN(U6318_n1) );
  NOR2X0 U6318_U1 ( .IN1(n4497), .IN2(U6318_n1), .QN(WX2169) );
  INVX0 U6319_U2 ( .INP(WX2104), .ZN(U6319_n1) );
  NOR2X0 U6319_U1 ( .IN1(n4497), .IN2(U6319_n1), .QN(WX2167) );
  INVX0 U6320_U2 ( .INP(WX2102), .ZN(U6320_n1) );
  NOR2X0 U6320_U1 ( .IN1(n4497), .IN2(U6320_n1), .QN(WX2165) );
  INVX0 U6321_U2 ( .INP(test_so17), .ZN(U6321_n1) );
  NOR2X0 U6321_U1 ( .IN1(n4497), .IN2(U6321_n1), .QN(WX2163) );
  INVX0 U6322_U2 ( .INP(WX2098), .ZN(U6322_n1) );
  NOR2X0 U6322_U1 ( .IN1(n4497), .IN2(U6322_n1), .QN(WX2161) );
  INVX0 U6323_U2 ( .INP(WX2096), .ZN(U6323_n1) );
  NOR2X0 U6323_U1 ( .IN1(n4515), .IN2(U6323_n1), .QN(WX2159) );
  INVX0 U6324_U2 ( .INP(WX2094), .ZN(U6324_n1) );
  NOR2X0 U6324_U1 ( .IN1(n4515), .IN2(U6324_n1), .QN(WX2157) );
  INVX0 U6325_U2 ( .INP(WX2092), .ZN(U6325_n1) );
  NOR2X0 U6325_U1 ( .IN1(n4515), .IN2(U6325_n1), .QN(WX2155) );
  INVX0 U6326_U2 ( .INP(WX2090), .ZN(U6326_n1) );
  NOR2X0 U6326_U1 ( .IN1(n4515), .IN2(U6326_n1), .QN(WX2153) );
  INVX0 U6327_U2 ( .INP(WX2088), .ZN(U6327_n1) );
  NOR2X0 U6327_U1 ( .IN1(n4515), .IN2(U6327_n1), .QN(WX2151) );
  INVX0 U6328_U2 ( .INP(WX2086), .ZN(U6328_n1) );
  NOR2X0 U6328_U1 ( .IN1(n4515), .IN2(U6328_n1), .QN(WX2149) );
  INVX0 U6329_U2 ( .INP(WX2084), .ZN(U6329_n1) );
  NOR2X0 U6329_U1 ( .IN1(n4515), .IN2(U6329_n1), .QN(WX2147) );
  INVX0 U6330_U2 ( .INP(WX2082), .ZN(U6330_n1) );
  NOR2X0 U6330_U1 ( .IN1(n4515), .IN2(U6330_n1), .QN(WX2145) );
  INVX0 U6331_U2 ( .INP(WX2080), .ZN(U6331_n1) );
  NOR2X0 U6331_U1 ( .IN1(n4515), .IN2(U6331_n1), .QN(WX2143) );
  INVX0 U6332_U2 ( .INP(WX2078), .ZN(U6332_n1) );
  NOR2X0 U6332_U1 ( .IN1(n4515), .IN2(U6332_n1), .QN(WX2141) );
  INVX0 U6333_U2 ( .INP(WX2076), .ZN(U6333_n1) );
  NOR2X0 U6333_U1 ( .IN1(n4515), .IN2(U6333_n1), .QN(WX2139) );
  INVX0 U6334_U2 ( .INP(WX2074), .ZN(U6334_n1) );
  NOR2X0 U6334_U1 ( .IN1(n4515), .IN2(U6334_n1), .QN(WX2137) );
  INVX0 U6335_U2 ( .INP(WX2072), .ZN(U6335_n1) );
  NOR2X0 U6335_U1 ( .IN1(n4515), .IN2(U6335_n1), .QN(WX2135) );
  INVX0 U6336_U2 ( .INP(WX2070), .ZN(U6336_n1) );
  NOR2X0 U6336_U1 ( .IN1(n4514), .IN2(U6336_n1), .QN(WX2133) );
  INVX0 U6337_U2 ( .INP(WX2068), .ZN(U6337_n1) );
  NOR2X0 U6337_U1 ( .IN1(n4514), .IN2(U6337_n1), .QN(WX2131) );
  INVX0 U6338_U2 ( .INP(WX2066), .ZN(U6338_n1) );
  NOR2X0 U6338_U1 ( .IN1(n4514), .IN2(U6338_n1), .QN(WX2129) );
  INVX0 U6339_U2 ( .INP(test_so16), .ZN(U6339_n1) );
  NOR2X0 U6339_U1 ( .IN1(n4514), .IN2(U6339_n1), .QN(WX2127) );
  INVX0 U6340_U2 ( .INP(WX2062), .ZN(U6340_n1) );
  NOR2X0 U6340_U1 ( .IN1(n4514), .IN2(U6340_n1), .QN(WX2125) );
  INVX0 U6341_U2 ( .INP(WX2060), .ZN(U6341_n1) );
  NOR2X0 U6341_U1 ( .IN1(n4514), .IN2(U6341_n1), .QN(WX2123) );
  INVX0 U6342_U2 ( .INP(WX2058), .ZN(U6342_n1) );
  NOR2X0 U6342_U1 ( .IN1(n4514), .IN2(U6342_n1), .QN(WX2121) );
  INVX0 U6343_U2 ( .INP(WX2056), .ZN(U6343_n1) );
  NOR2X0 U6343_U1 ( .IN1(n4514), .IN2(U6343_n1), .QN(WX2119) );
  INVX0 U6344_U2 ( .INP(WX2054), .ZN(U6344_n1) );
  NOR2X0 U6344_U1 ( .IN1(n4514), .IN2(U6344_n1), .QN(WX2117) );
  INVX0 U6345_U2 ( .INP(WX2052), .ZN(U6345_n1) );
  NOR2X0 U6345_U1 ( .IN1(n4514), .IN2(U6345_n1), .QN(WX2115) );
  INVX0 U6346_U2 ( .INP(WX2050), .ZN(U6346_n1) );
  NOR2X0 U6346_U1 ( .IN1(n4514), .IN2(U6346_n1), .QN(WX2113) );
  INVX0 U6347_U2 ( .INP(WX2048), .ZN(U6347_n1) );
  NOR2X0 U6347_U1 ( .IN1(n4514), .IN2(U6347_n1), .QN(WX2111) );
  INVX0 U6348_U2 ( .INP(WX2046), .ZN(U6348_n1) );
  NOR2X0 U6348_U1 ( .IN1(n4514), .IN2(U6348_n1), .QN(WX2109) );
  INVX0 U6349_U2 ( .INP(WX2044), .ZN(U6349_n1) );
  NOR2X0 U6349_U1 ( .IN1(n4513), .IN2(U6349_n1), .QN(WX2107) );
  INVX0 U6350_U2 ( .INP(WX2042), .ZN(U6350_n1) );
  NOR2X0 U6350_U1 ( .IN1(n4513), .IN2(U6350_n1), .QN(WX2105) );
  INVX0 U6351_U2 ( .INP(WX2040), .ZN(U6351_n1) );
  NOR2X0 U6351_U1 ( .IN1(n4513), .IN2(U6351_n1), .QN(WX2103) );
  INVX0 U6352_U2 ( .INP(WX2038), .ZN(U6352_n1) );
  NOR2X0 U6352_U1 ( .IN1(n4513), .IN2(U6352_n1), .QN(WX2101) );
  INVX0 U6353_U2 ( .INP(WX2036), .ZN(U6353_n1) );
  NOR2X0 U6353_U1 ( .IN1(n4513), .IN2(U6353_n1), .QN(WX2099) );
  INVX0 U6354_U2 ( .INP(WX2034), .ZN(U6354_n1) );
  NOR2X0 U6354_U1 ( .IN1(n4513), .IN2(U6354_n1), .QN(WX2097) );
  INVX0 U6355_U2 ( .INP(WX2032), .ZN(U6355_n1) );
  NOR2X0 U6355_U1 ( .IN1(n4513), .IN2(U6355_n1), .QN(WX2095) );
  INVX0 U6356_U2 ( .INP(WX2030), .ZN(U6356_n1) );
  NOR2X0 U6356_U1 ( .IN1(n4513), .IN2(U6356_n1), .QN(WX2093) );
  INVX0 U6357_U2 ( .INP(test_so15), .ZN(U6357_n1) );
  NOR2X0 U6357_U1 ( .IN1(n4513), .IN2(U6357_n1), .QN(WX2091) );
  INVX0 U6358_U2 ( .INP(WX2026), .ZN(U6358_n1) );
  NOR2X0 U6358_U1 ( .IN1(n4513), .IN2(U6358_n1), .QN(WX2089) );
  INVX0 U6359_U2 ( .INP(WX2024), .ZN(U6359_n1) );
  NOR2X0 U6359_U1 ( .IN1(n4513), .IN2(U6359_n1), .QN(WX2087) );
  INVX0 U6360_U2 ( .INP(WX2022), .ZN(U6360_n1) );
  NOR2X0 U6360_U1 ( .IN1(n4513), .IN2(U6360_n1), .QN(WX2085) );
  INVX0 U6361_U2 ( .INP(WX2020), .ZN(U6361_n1) );
  NOR2X0 U6361_U1 ( .IN1(n4513), .IN2(U6361_n1), .QN(WX2083) );
  INVX0 U6362_U2 ( .INP(WX2018), .ZN(U6362_n1) );
  NOR2X0 U6362_U1 ( .IN1(n4512), .IN2(U6362_n1), .QN(WX2081) );
  INVX0 U6363_U2 ( .INP(WX2016), .ZN(U6363_n1) );
  NOR2X0 U6363_U1 ( .IN1(n4512), .IN2(U6363_n1), .QN(WX2079) );
  INVX0 U6364_U2 ( .INP(WX2014), .ZN(U6364_n1) );
  NOR2X0 U6364_U1 ( .IN1(n4512), .IN2(U6364_n1), .QN(WX2077) );
  INVX0 U6365_U2 ( .INP(WX2012), .ZN(U6365_n1) );
  NOR2X0 U6365_U1 ( .IN1(n4512), .IN2(U6365_n1), .QN(WX2075) );
  INVX0 U6366_U2 ( .INP(WX2010), .ZN(U6366_n1) );
  NOR2X0 U6366_U1 ( .IN1(n4512), .IN2(U6366_n1), .QN(WX2073) );
  INVX0 U6367_U2 ( .INP(WX2008), .ZN(U6367_n1) );
  NOR2X0 U6367_U1 ( .IN1(n4512), .IN2(U6367_n1), .QN(WX2071) );
  INVX0 U6368_U2 ( .INP(WX2006), .ZN(U6368_n1) );
  NOR2X0 U6368_U1 ( .IN1(n4512), .IN2(U6368_n1), .QN(WX2069) );
  INVX0 U6369_U2 ( .INP(WX2004), .ZN(U6369_n1) );
  NOR2X0 U6369_U1 ( .IN1(n4512), .IN2(U6369_n1), .QN(WX2067) );
  INVX0 U6370_U2 ( .INP(WX2002), .ZN(U6370_n1) );
  NOR2X0 U6370_U1 ( .IN1(n4512), .IN2(U6370_n1), .QN(WX2065) );
  INVX0 U6371_U2 ( .INP(WX2000), .ZN(U6371_n1) );
  NOR2X0 U6371_U1 ( .IN1(n4512), .IN2(U6371_n1), .QN(WX2063) );
  INVX0 U6372_U2 ( .INP(WX1998), .ZN(U6372_n1) );
  NOR2X0 U6372_U1 ( .IN1(n4512), .IN2(U6372_n1), .QN(WX2061) );
  INVX0 U6373_U2 ( .INP(WX1996), .ZN(U6373_n1) );
  NOR2X0 U6373_U1 ( .IN1(n4512), .IN2(U6373_n1), .QN(WX2059) );
  INVX0 U6374_U2 ( .INP(WX1994), .ZN(U6374_n1) );
  NOR2X0 U6374_U1 ( .IN1(n4512), .IN2(U6374_n1), .QN(WX2057) );
  INVX0 U6375_U2 ( .INP(test_so14), .ZN(U6375_n1) );
  NOR2X0 U6375_U1 ( .IN1(n4511), .IN2(U6375_n1), .QN(WX2055) );
  INVX0 U6376_U2 ( .INP(WX1990), .ZN(U6376_n1) );
  NOR2X0 U6376_U1 ( .IN1(n4511), .IN2(U6376_n1), .QN(WX2053) );
  INVX0 U6377_U2 ( .INP(WX1988), .ZN(U6377_n1) );
  NOR2X0 U6377_U1 ( .IN1(n4511), .IN2(U6377_n1), .QN(WX2051) );
  INVX0 U6378_U2 ( .INP(WX1986), .ZN(U6378_n1) );
  NOR2X0 U6378_U1 ( .IN1(n4511), .IN2(U6378_n1), .QN(WX2049) );
  INVX0 U6379_U2 ( .INP(WX1984), .ZN(U6379_n1) );
  NOR2X0 U6379_U1 ( .IN1(n4511), .IN2(U6379_n1), .QN(WX2047) );
  INVX0 U6380_U2 ( .INP(WX1982), .ZN(U6380_n1) );
  NOR2X0 U6380_U1 ( .IN1(n4511), .IN2(U6380_n1), .QN(WX2045) );
  INVX0 U6381_U2 ( .INP(WX1980), .ZN(U6381_n1) );
  NOR2X0 U6381_U1 ( .IN1(n4511), .IN2(U6381_n1), .QN(WX2043) );
  INVX0 U6382_U2 ( .INP(WX1978), .ZN(U6382_n1) );
  NOR2X0 U6382_U1 ( .IN1(n4511), .IN2(U6382_n1), .QN(WX2041) );
  INVX0 U6383_U2 ( .INP(WX1976), .ZN(U6383_n1) );
  NOR2X0 U6383_U1 ( .IN1(n4511), .IN2(U6383_n1), .QN(WX2039) );
  INVX0 U6384_U2 ( .INP(WX1974), .ZN(U6384_n1) );
  NOR2X0 U6384_U1 ( .IN1(n4511), .IN2(U6384_n1), .QN(WX2037) );
  INVX0 U6385_U2 ( .INP(WX1972), .ZN(U6385_n1) );
  NOR2X0 U6385_U1 ( .IN1(n4511), .IN2(U6385_n1), .QN(WX2035) );
  INVX0 U6386_U2 ( .INP(WX1970), .ZN(U6386_n1) );
  NOR2X0 U6386_U1 ( .IN1(n4511), .IN2(U6386_n1), .QN(WX2033) );
  INVX0 U6387_U2 ( .INP(WX835), .ZN(U6387_n1) );
  NOR2X0 U6387_U1 ( .IN1(n4511), .IN2(U6387_n1), .QN(WX898) );
  INVX0 U6388_U2 ( .INP(WX833), .ZN(U6388_n1) );
  NOR2X0 U6388_U1 ( .IN1(n4510), .IN2(U6388_n1), .QN(WX896) );
  INVX0 U6389_U2 ( .INP(test_so7), .ZN(U6389_n1) );
  NOR2X0 U6389_U1 ( .IN1(n4510), .IN2(U6389_n1), .QN(WX894) );
  INVX0 U6390_U2 ( .INP(WX829), .ZN(U6390_n1) );
  NOR2X0 U6390_U1 ( .IN1(n4510), .IN2(U6390_n1), .QN(WX892) );
  INVX0 U6391_U2 ( .INP(WX827), .ZN(U6391_n1) );
  NOR2X0 U6391_U1 ( .IN1(n4510), .IN2(U6391_n1), .QN(WX890) );
  INVX0 U6392_U2 ( .INP(WX825), .ZN(U6392_n1) );
  NOR2X0 U6392_U1 ( .IN1(n4510), .IN2(U6392_n1), .QN(WX888) );
  INVX0 U6393_U2 ( .INP(WX823), .ZN(U6393_n1) );
  NOR2X0 U6393_U1 ( .IN1(n4510), .IN2(U6393_n1), .QN(WX886) );
  INVX0 U6394_U2 ( .INP(WX821), .ZN(U6394_n1) );
  NOR2X0 U6394_U1 ( .IN1(n4510), .IN2(U6394_n1), .QN(WX884) );
  INVX0 U6395_U2 ( .INP(WX819), .ZN(U6395_n1) );
  NOR2X0 U6395_U1 ( .IN1(n4510), .IN2(U6395_n1), .QN(WX882) );
  INVX0 U6396_U2 ( .INP(WX817), .ZN(U6396_n1) );
  NOR2X0 U6396_U1 ( .IN1(n4510), .IN2(U6396_n1), .QN(WX880) );
  INVX0 U6397_U2 ( .INP(WX815), .ZN(U6397_n1) );
  NOR2X0 U6397_U1 ( .IN1(n4510), .IN2(U6397_n1), .QN(WX878) );
  INVX0 U6398_U2 ( .INP(WX813), .ZN(U6398_n1) );
  NOR2X0 U6398_U1 ( .IN1(n4510), .IN2(U6398_n1), .QN(WX876) );
  INVX0 U6399_U2 ( .INP(WX811), .ZN(U6399_n1) );
  NOR2X0 U6399_U1 ( .IN1(n4510), .IN2(U6399_n1), .QN(WX874) );
  INVX0 U6400_U2 ( .INP(WX809), .ZN(U6400_n1) );
  NOR2X0 U6400_U1 ( .IN1(n4510), .IN2(U6400_n1), .QN(WX872) );
  INVX0 U6401_U2 ( .INP(WX807), .ZN(U6401_n1) );
  NOR2X0 U6401_U1 ( .IN1(n4509), .IN2(U6401_n1), .QN(WX870) );
  INVX0 U6402_U2 ( .INP(WX805), .ZN(U6402_n1) );
  NOR2X0 U6402_U1 ( .IN1(n4509), .IN2(U6402_n1), .QN(WX868) );
  INVX0 U6403_U2 ( .INP(WX803), .ZN(U6403_n1) );
  NOR2X0 U6403_U1 ( .IN1(n4509), .IN2(U6403_n1), .QN(WX866) );
  INVX0 U6404_U2 ( .INP(WX801), .ZN(U6404_n1) );
  NOR2X0 U6404_U1 ( .IN1(n4509), .IN2(U6404_n1), .QN(WX864) );
  INVX0 U6405_U2 ( .INP(WX799), .ZN(U6405_n1) );
  NOR2X0 U6405_U1 ( .IN1(n4509), .IN2(U6405_n1), .QN(WX862) );
  INVX0 U6406_U2 ( .INP(WX797), .ZN(U6406_n1) );
  NOR2X0 U6406_U1 ( .IN1(n4509), .IN2(U6406_n1), .QN(WX860) );
  INVX0 U6407_U2 ( .INP(test_so6), .ZN(U6407_n1) );
  NOR2X0 U6407_U1 ( .IN1(n4509), .IN2(U6407_n1), .QN(WX858) );
  INVX0 U6408_U2 ( .INP(WX793), .ZN(U6408_n1) );
  NOR2X0 U6408_U1 ( .IN1(n4509), .IN2(U6408_n1), .QN(WX856) );
  INVX0 U6409_U2 ( .INP(WX791), .ZN(U6409_n1) );
  NOR2X0 U6409_U1 ( .IN1(n4509), .IN2(U6409_n1), .QN(WX854) );
  INVX0 U6410_U2 ( .INP(WX789), .ZN(U6410_n1) );
  NOR2X0 U6410_U1 ( .IN1(n4509), .IN2(U6410_n1), .QN(WX852) );
  INVX0 U6411_U2 ( .INP(WX787), .ZN(U6411_n1) );
  NOR2X0 U6411_U1 ( .IN1(n4509), .IN2(U6411_n1), .QN(WX850) );
  INVX0 U6412_U2 ( .INP(WX785), .ZN(U6412_n1) );
  NOR2X0 U6412_U1 ( .IN1(n4509), .IN2(U6412_n1), .QN(WX848) );
  INVX0 U6413_U2 ( .INP(WX783), .ZN(U6413_n1) );
  NOR2X0 U6413_U1 ( .IN1(n4508), .IN2(U6413_n1), .QN(WX846) );
  INVX0 U6414_U2 ( .INP(WX781), .ZN(U6414_n1) );
  NOR2X0 U6414_U1 ( .IN1(n4508), .IN2(U6414_n1), .QN(WX844) );
  INVX0 U6415_U2 ( .INP(WX779), .ZN(U6415_n1) );
  NOR2X0 U6415_U1 ( .IN1(n4508), .IN2(U6415_n1), .QN(WX842) );
  INVX0 U6416_U2 ( .INP(WX777), .ZN(U6416_n1) );
  NOR2X0 U6416_U1 ( .IN1(n4508), .IN2(U6416_n1), .QN(WX840) );
  INVX0 U6417_U2 ( .INP(WX775), .ZN(U6417_n1) );
  NOR2X0 U6417_U1 ( .IN1(n4508), .IN2(U6417_n1), .QN(WX838) );
  INVX0 U6418_U2 ( .INP(WX773), .ZN(U6418_n1) );
  NOR2X0 U6418_U1 ( .IN1(n4508), .IN2(U6418_n1), .QN(WX836) );
  INVX0 U6419_U2 ( .INP(WX771), .ZN(U6419_n1) );
  NOR2X0 U6419_U1 ( .IN1(n4508), .IN2(U6419_n1), .QN(WX834) );
  INVX0 U6420_U2 ( .INP(WX769), .ZN(U6420_n1) );
  NOR2X0 U6420_U1 ( .IN1(n4508), .IN2(U6420_n1), .QN(WX832) );
  INVX0 U6421_U2 ( .INP(WX767), .ZN(U6421_n1) );
  NOR2X0 U6421_U1 ( .IN1(n4508), .IN2(U6421_n1), .QN(WX830) );
  INVX0 U6422_U2 ( .INP(WX765), .ZN(U6422_n1) );
  NOR2X0 U6422_U1 ( .IN1(n4508), .IN2(U6422_n1), .QN(WX828) );
  INVX0 U6423_U2 ( .INP(WX763), .ZN(U6423_n1) );
  NOR2X0 U6423_U1 ( .IN1(n4508), .IN2(U6423_n1), .QN(WX826) );
  INVX0 U6424_U2 ( .INP(WX761), .ZN(U6424_n1) );
  NOR2X0 U6424_U1 ( .IN1(n4508), .IN2(U6424_n1), .QN(WX824) );
  INVX0 U6425_U2 ( .INP(test_so5), .ZN(U6425_n1) );
  NOR2X0 U6425_U1 ( .IN1(n4508), .IN2(U6425_n1), .QN(WX822) );
  INVX0 U6426_U2 ( .INP(WX757), .ZN(U6426_n1) );
  NOR2X0 U6426_U1 ( .IN1(n4507), .IN2(U6426_n1), .QN(WX820) );
  INVX0 U6427_U2 ( .INP(WX755), .ZN(U6427_n1) );
  NOR2X0 U6427_U1 ( .IN1(n4507), .IN2(U6427_n1), .QN(WX818) );
  INVX0 U6428_U2 ( .INP(WX753), .ZN(U6428_n1) );
  NOR2X0 U6428_U1 ( .IN1(n4507), .IN2(U6428_n1), .QN(WX816) );
  INVX0 U6429_U2 ( .INP(WX751), .ZN(U6429_n1) );
  NOR2X0 U6429_U1 ( .IN1(n4507), .IN2(U6429_n1), .QN(WX814) );
  INVX0 U6430_U2 ( .INP(WX749), .ZN(U6430_n1) );
  NOR2X0 U6430_U1 ( .IN1(n4507), .IN2(U6430_n1), .QN(WX812) );
  INVX0 U6431_U2 ( .INP(WX747), .ZN(U6431_n1) );
  NOR2X0 U6431_U1 ( .IN1(n4507), .IN2(U6431_n1), .QN(WX810) );
  INVX0 U6432_U2 ( .INP(WX745), .ZN(U6432_n1) );
  NOR2X0 U6432_U1 ( .IN1(n4507), .IN2(U6432_n1), .QN(WX808) );
  INVX0 U6433_U2 ( .INP(WX743), .ZN(U6433_n1) );
  NOR2X0 U6433_U1 ( .IN1(n4507), .IN2(U6433_n1), .QN(WX806) );
  INVX0 U6434_U2 ( .INP(WX741), .ZN(U6434_n1) );
  NOR2X0 U6434_U1 ( .IN1(n4507), .IN2(U6434_n1), .QN(WX804) );
  INVX0 U6435_U2 ( .INP(WX739), .ZN(U6435_n1) );
  NOR2X0 U6435_U1 ( .IN1(n4507), .IN2(U6435_n1), .QN(WX802) );
  INVX0 U6436_U2 ( .INP(WX737), .ZN(U6436_n1) );
  NOR2X0 U6436_U1 ( .IN1(n4507), .IN2(U6436_n1), .QN(WX800) );
  INVX0 U6437_U2 ( .INP(WX735), .ZN(U6437_n1) );
  NOR2X0 U6437_U1 ( .IN1(n4507), .IN2(U6437_n1), .QN(WX798) );
  INVX0 U6438_U2 ( .INP(WX733), .ZN(U6438_n1) );
  NOR2X0 U6438_U1 ( .IN1(n4507), .IN2(U6438_n1), .QN(WX796) );
  INVX0 U6439_U2 ( .INP(WX731), .ZN(U6439_n1) );
  NOR2X0 U6439_U1 ( .IN1(n4506), .IN2(U6439_n1), .QN(WX794) );
  INVX0 U6440_U2 ( .INP(WX729), .ZN(U6440_n1) );
  NOR2X0 U6440_U1 ( .IN1(n4506), .IN2(U6440_n1), .QN(WX792) );
  INVX0 U6441_U2 ( .INP(WX727), .ZN(U6441_n1) );
  NOR2X0 U6441_U1 ( .IN1(n4506), .IN2(U6441_n1), .QN(WX790) );
  INVX0 U6442_U2 ( .INP(WX725), .ZN(U6442_n1) );
  NOR2X0 U6442_U1 ( .IN1(n4506), .IN2(U6442_n1), .QN(WX788) );
  INVX0 U6443_U2 ( .INP(test_so4), .ZN(U6443_n1) );
  NOR2X0 U6443_U1 ( .IN1(n4506), .IN2(U6443_n1), .QN(WX786) );
  INVX0 U6444_U2 ( .INP(WX721), .ZN(U6444_n1) );
  NOR2X0 U6444_U1 ( .IN1(n4506), .IN2(U6444_n1), .QN(WX784) );
  INVX0 U6445_U2 ( .INP(WX719), .ZN(U6445_n1) );
  NOR2X0 U6445_U1 ( .IN1(n4506), .IN2(U6445_n1), .QN(WX782) );
  INVX0 U6446_U2 ( .INP(WX717), .ZN(U6446_n1) );
  NOR2X0 U6446_U1 ( .IN1(n4506), .IN2(U6446_n1), .QN(WX780) );
  INVX0 U6447_U2 ( .INP(WX715), .ZN(U6447_n1) );
  NOR2X0 U6447_U1 ( .IN1(n4506), .IN2(U6447_n1), .QN(WX778) );
  INVX0 U6448_U2 ( .INP(WX713), .ZN(U6448_n1) );
  NOR2X0 U6448_U1 ( .IN1(n4506), .IN2(U6448_n1), .QN(WX776) );
  INVX0 U6449_U2 ( .INP(WX711), .ZN(U6449_n1) );
  NOR2X0 U6449_U1 ( .IN1(n4506), .IN2(U6449_n1), .QN(WX774) );
  INVX0 U6450_U2 ( .INP(WX709), .ZN(U6450_n1) );
  NOR2X0 U6450_U1 ( .IN1(n4506), .IN2(U6450_n1), .QN(WX772) );
  INVX0 U6451_U2 ( .INP(WX707), .ZN(U6451_n1) );
  NOR2X0 U6451_U1 ( .IN1(n4506), .IN2(U6451_n1), .QN(WX770) );
  INVX0 U6452_U2 ( .INP(WX705), .ZN(U6452_n1) );
  NOR2X0 U6452_U1 ( .IN1(n4505), .IN2(U6452_n1), .QN(WX768) );
  INVX0 U6453_U2 ( .INP(WX703), .ZN(U6453_n1) );
  NOR2X0 U6453_U1 ( .IN1(n4505), .IN2(U6453_n1), .QN(WX766) );
  INVX0 U6454_U2 ( .INP(WX701), .ZN(U6454_n1) );
  NOR2X0 U6454_U1 ( .IN1(n4505), .IN2(U6454_n1), .QN(WX764) );
  INVX0 U6455_U2 ( .INP(WX699), .ZN(U6455_n1) );
  NOR2X0 U6455_U1 ( .IN1(n4505), .IN2(U6455_n1), .QN(WX762) );
  INVX0 U6456_U2 ( .INP(WX697), .ZN(U6456_n1) );
  NOR2X0 U6456_U1 ( .IN1(n4505), .IN2(U6456_n1), .QN(WX760) );
  INVX0 U6457_U2 ( .INP(WX695), .ZN(U6457_n1) );
  NOR2X0 U6457_U1 ( .IN1(n4505), .IN2(U6457_n1), .QN(WX758) );
  INVX0 U6458_U2 ( .INP(WX693), .ZN(U6458_n1) );
  NOR2X0 U6458_U1 ( .IN1(n4505), .IN2(U6458_n1), .QN(WX756) );
  INVX0 U6459_U2 ( .INP(WX691), .ZN(U6459_n1) );
  NOR2X0 U6459_U1 ( .IN1(n4505), .IN2(U6459_n1), .QN(WX754) );
  INVX0 U6460_U2 ( .INP(WX689), .ZN(U6460_n1) );
  NOR2X0 U6460_U1 ( .IN1(n4505), .IN2(U6460_n1), .QN(WX752) );
  INVX0 U6461_U2 ( .INP(test_so3), .ZN(U6461_n1) );
  NOR2X0 U6461_U1 ( .IN1(n4505), .IN2(U6461_n1), .QN(WX750) );
  INVX0 U6462_U2 ( .INP(WX685), .ZN(U6462_n1) );
  NOR2X0 U6462_U1 ( .IN1(n4505), .IN2(U6462_n1), .QN(WX748) );
  INVX0 U6463_U2 ( .INP(WX683), .ZN(U6463_n1) );
  NOR2X0 U6463_U1 ( .IN1(n4505), .IN2(U6463_n1), .QN(WX746) );
  INVX0 U6464_U2 ( .INP(WX681), .ZN(U6464_n1) );
  NOR2X0 U6464_U1 ( .IN1(n4505), .IN2(U6464_n1), .QN(WX744) );
  INVX0 U6465_U2 ( .INP(WX679), .ZN(U6465_n1) );
  NOR2X0 U6465_U1 ( .IN1(n4504), .IN2(U6465_n1), .QN(WX742) );
  INVX0 U6466_U2 ( .INP(WX677), .ZN(U6466_n1) );
  NOR2X0 U6466_U1 ( .IN1(n4504), .IN2(U6466_n1), .QN(WX740) );
  INVX0 U6467_U2 ( .INP(WX675), .ZN(U6467_n1) );
  NOR2X0 U6467_U1 ( .IN1(n4504), .IN2(U6467_n1), .QN(WX738) );
  INVX0 U6468_U2 ( .INP(WX673), .ZN(U6468_n1) );
  NOR2X0 U6468_U1 ( .IN1(n4504), .IN2(U6468_n1), .QN(WX736) );
  INVX0 U6469_U2 ( .INP(WX671), .ZN(U6469_n1) );
  NOR2X0 U6469_U1 ( .IN1(n4504), .IN2(U6469_n1), .QN(WX734) );
  INVX0 U6470_U2 ( .INP(WX669), .ZN(U6470_n1) );
  NOR2X0 U6470_U1 ( .IN1(n4504), .IN2(U6470_n1), .QN(WX732) );
  INVX0 U6471_U2 ( .INP(WX667), .ZN(U6471_n1) );
  NOR2X0 U6471_U1 ( .IN1(n4504), .IN2(U6471_n1), .QN(WX730) );
  INVX0 U6472_U2 ( .INP(WX665), .ZN(U6472_n1) );
  NOR2X0 U6472_U1 ( .IN1(n4504), .IN2(U6472_n1), .QN(WX728) );
  INVX0 U6473_U2 ( .INP(WX663), .ZN(U6473_n1) );
  NOR2X0 U6473_U1 ( .IN1(n4504), .IN2(U6473_n1), .QN(WX726) );
  INVX0 U6474_U2 ( .INP(WX661), .ZN(U6474_n1) );
  NOR2X0 U6474_U1 ( .IN1(n4504), .IN2(U6474_n1), .QN(WX724) );
  INVX0 U6475_U2 ( .INP(WX659), .ZN(U6475_n1) );
  NOR2X0 U6475_U1 ( .IN1(n4504), .IN2(U6475_n1), .QN(WX722) );
  INVX0 U6476_U2 ( .INP(WX657), .ZN(U6476_n1) );
  NOR2X0 U6476_U1 ( .IN1(n4504), .IN2(U6476_n1), .QN(WX720) );
  INVX0 U6477_U2 ( .INP(WX655), .ZN(U6477_n1) );
  NOR2X0 U6477_U1 ( .IN1(n4504), .IN2(U6477_n1), .QN(WX718) );
  INVX0 U6478_U2 ( .INP(WX653), .ZN(U6478_n1) );
  NOR2X0 U6478_U1 ( .IN1(n4503), .IN2(U6478_n1), .QN(WX716) );
  INVX0 U6479_U2 ( .INP(test_so2), .ZN(U6479_n1) );
  NOR2X0 U6479_U1 ( .IN1(n4503), .IN2(U6479_n1), .QN(WX714) );
  INVX0 U6480_U2 ( .INP(WX649), .ZN(U6480_n1) );
  NOR2X0 U6480_U1 ( .IN1(n4503), .IN2(U6480_n1), .QN(WX712) );
  INVX0 U6481_U2 ( .INP(WX647), .ZN(U6481_n1) );
  NOR2X0 U6481_U1 ( .IN1(n4503), .IN2(U6481_n1), .QN(WX710) );
  INVX0 U6482_U2 ( .INP(WX645), .ZN(U6482_n1) );
  NOR2X0 U6482_U1 ( .IN1(n4509), .IN2(U6482_n1), .QN(WX708) );
endmodule

