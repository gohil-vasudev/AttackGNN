module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n155_, new_n384_, new_n410_, new_n236_, new_n238_, new_n92_, new_n79_, new_n250_, new_n113_, new_n288_, new_n371_, new_n97_, new_n421_, new_n202_, new_n296_, new_n308_, new_n368_, new_n232_, new_n258_, new_n76_, new_n176_, new_n283_, new_n223_, new_n390_, new_n156_, new_n306_, new_n366_, new_n291_, new_n261_, new_n241_, new_n309_, new_n186_, new_n339_, new_n365_, new_n197_, new_n386_, new_n82_, new_n401_, new_n389_, new_n323_, new_n259_, new_n362_, new_n227_, new_n222_, new_n170_, new_n246_, new_n400_, new_n328_, new_n266_, new_n367_, new_n173_, new_n220_, new_n130_, new_n268_, new_n374_, new_n376_, new_n380_, new_n214_, new_n424_, new_n138_, new_n310_, new_n144_, new_n275_, new_n114_, new_n188_, new_n240_, new_n413_, new_n352_, new_n211_, new_n123_, new_n127_, new_n342_, new_n126_, new_n177_, new_n264_, new_n379_, new_n273_, new_n224_, new_n270_, new_n317_, new_n344_, new_n143_, new_n287_, new_n125_, new_n145_, new_n253_, new_n403_, new_n90_, new_n237_, new_n427_, new_n234_, new_n149_, new_n393_, new_n260_, new_n418_, new_n251_, new_n189_, new_n300_, new_n292_, new_n106_, new_n411_, new_n215_, new_n152_, new_n157_, new_n107_, new_n93_, new_n182_, new_n153_, new_n407_, new_n81_, new_n133_, new_n257_, new_n212_, new_n151_, new_n364_, new_n219_, new_n231_, new_n313_, new_n78_, new_n239_, new_n382_, new_n272_, new_n282_, new_n201_, new_n428_, new_n192_, new_n414_, new_n199_, new_n146_, new_n88_, new_n360_, new_n98_, new_n110_, new_n315_, new_n302_, new_n191_, new_n124_, new_n95_, new_n225_, new_n164_, new_n230_, new_n281_, new_n87_, new_n387_, new_n103_, new_n112_, new_n248_, new_n350_, new_n117_, new_n121_, new_n415_, new_n167_, new_n221_, new_n385_, new_n243_, new_n345_, new_n298_, new_n184_, new_n154_, new_n131_, new_n255_, new_n174_, new_n297_, new_n361_, new_n150_, new_n354_, new_n392_, new_n108_, new_n137_, new_n183_, new_n303_, new_n105_, new_n340_, new_n147_, new_n285_, new_n80_, new_n351_, new_n209_, new_n337_, new_n203_, new_n316_, new_n325_, new_n417_, new_n180_, new_n332_, new_n318_, new_n163_, new_n148_, new_n321_, new_n122_, new_n324_, new_n111_, new_n158_, new_n252_, new_n262_, new_n160_, new_n312_, new_n271_, new_n274_, new_n372_, new_n100_, new_n242_, new_n218_, new_n115_, new_n307_, new_n190_, new_n305_, new_n420_, new_n408_, new_n423_, new_n205_, new_n134_, new_n141_, new_n206_, new_n109_, new_n254_, new_n429_, new_n355_, new_n353_, new_n85_, new_n265_, new_n370_, new_n256_, new_n278_, new_n304_, new_n381_, new_n388_, new_n217_, new_n101_, new_n269_, new_n194_, new_n394_, new_n116_, new_n299_, new_n129_, new_n142_, new_n139_, new_n314_, new_n118_, new_n363_, new_n165_, new_n327_, new_n216_, new_n77_, new_n196_, new_n280_, new_n426_, new_n319_, new_n235_, new_n398_, new_n301_, new_n169_, new_n395_, new_n338_, new_n383_, new_n343_, new_n210_, new_n207_, new_n267_, new_n336_, new_n140_, new_n377_, new_n247_, new_n330_, new_n375_, new_n294_, new_n187_, new_n311_, new_n86_, new_n84_, new_n195_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n357_, new_n320_, new_n349_, new_n244_, new_n172_, new_n277_, new_n245_, new_n402_, new_n89_, new_n286_, new_n404_, new_n335_, new_n347_, new_n193_, new_n91_, new_n346_, new_n396_, new_n198_, new_n128_, new_n358_, new_n208_, new_n348_, new_n159_, new_n83_, new_n322_, new_n228_, new_n289_, new_n179_, new_n425_, new_n175_, new_n226_, new_n397_, new_n104_, new_n185_, new_n399_, new_n373_, new_n171_, new_n200_, new_n422_, new_n99_, new_n329_, new_n249_, new_n233_, new_n136_, new_n284_, new_n119_, new_n293_, new_n391_, new_n96_, new_n178_, new_n168_, new_n279_, new_n295_, new_n359_, new_n132_, new_n120_, new_n166_, new_n162_, new_n409_, new_n161_, new_n406_, new_n356_, new_n333_, new_n229_, new_n290_, new_n94_, new_n204_, new_n369_, new_n181_, new_n135_, new_n276_, new_n405_;

not g000 ( new_n76_, N108 );
or g001 ( new_n77_, new_n76_, N102 );
and g002 ( new_n78_, new_n77_, keyIn_0_4 );
not g003 ( new_n79_, keyIn_0_4 );
not g004 ( new_n80_, N102 );
and g005 ( new_n81_, new_n79_, new_n80_, N108 );
or g006 ( new_n82_, new_n78_, new_n81_ );
not g007 ( new_n83_, N69 );
or g008 ( new_n84_, new_n83_, N63 );
not g009 ( new_n85_, N56 );
or g010 ( new_n86_, new_n85_, N50 );
not g011 ( new_n87_, N95 );
or g012 ( new_n88_, new_n87_, N89 );
not g013 ( new_n89_, N82 );
or g014 ( new_n90_, new_n89_, N76 );
and g015 ( new_n91_, new_n84_, new_n86_, new_n88_, new_n90_ );
not g016 ( new_n92_, N17 );
or g017 ( new_n93_, new_n92_, N11 );
not g018 ( new_n94_, N4 );
or g019 ( new_n95_, new_n94_, N1 );
not g020 ( new_n96_, N43 );
or g021 ( new_n97_, new_n96_, N37 );
not g022 ( new_n98_, N30 );
or g023 ( new_n99_, new_n98_, N24 );
and g024 ( new_n100_, new_n93_, new_n95_, new_n97_, new_n99_ );
and g025 ( new_n101_, new_n82_, new_n91_, new_n100_ );
not g026 ( N223, new_n101_ );
not g027 ( new_n103_, N34 );
not g028 ( new_n104_, keyIn_0_11 );
not g029 ( new_n105_, new_n99_ );
or g030 ( new_n106_, new_n101_, new_n105_ );
and g031 ( new_n107_, new_n106_, new_n104_ );
and g032 ( new_n108_, N223, keyIn_0_11, new_n99_ );
or g033 ( new_n109_, new_n107_, new_n108_ );
and g034 ( new_n110_, new_n109_, N30, new_n103_ );
or g035 ( new_n111_, new_n110_, keyIn_0_16 );
and g036 ( new_n112_, new_n109_, keyIn_0_16, N30, new_n103_ );
not g037 ( new_n113_, new_n112_ );
and g038 ( new_n114_, new_n111_, new_n113_ );
not g039 ( new_n115_, new_n95_ );
or g040 ( new_n116_, new_n101_, new_n115_ );
and g041 ( new_n117_, new_n91_, new_n100_ );
and g042 ( new_n118_, new_n117_, new_n82_, new_n115_ );
not g043 ( new_n119_, new_n118_ );
not g044 ( new_n120_, N8 );
and g045 ( new_n121_, keyIn_0_0, N4 );
not g046 ( new_n122_, new_n121_ );
or g047 ( new_n123_, keyIn_0_0, N4 );
and g048 ( new_n124_, new_n122_, new_n123_ );
and g049 ( new_n125_, new_n124_, new_n120_ );
and g050 ( new_n126_, new_n116_, new_n119_, new_n125_ );
not g051 ( new_n127_, N60 );
not g052 ( new_n128_, new_n86_ );
and g053 ( new_n129_, new_n117_, new_n82_, new_n128_ );
not g054 ( new_n130_, new_n129_ );
or g055 ( new_n131_, new_n101_, new_n128_ );
and g056 ( new_n132_, new_n131_, new_n130_, N56, new_n127_ );
not g057 ( new_n133_, N86 );
not g058 ( new_n134_, new_n90_ );
or g059 ( new_n135_, new_n101_, new_n134_ );
and g060 ( new_n136_, new_n135_, N82, new_n133_ );
or g061 ( new_n137_, new_n132_, new_n126_, new_n136_ );
not g062 ( new_n138_, N21 );
not g063 ( new_n139_, new_n93_ );
or g064 ( new_n140_, new_n101_, new_n139_ );
and g065 ( new_n141_, new_n140_, keyIn_0_10 );
not g066 ( new_n142_, keyIn_0_10 );
and g067 ( new_n143_, N223, new_n142_, new_n93_ );
or g068 ( new_n144_, new_n141_, new_n143_ );
and g069 ( new_n145_, keyIn_0_1, N17 );
not g070 ( new_n146_, new_n145_ );
or g071 ( new_n147_, keyIn_0_1, N17 );
and g072 ( new_n148_, new_n146_, new_n147_ );
not g073 ( new_n149_, new_n148_ );
and g074 ( new_n150_, new_n144_, new_n138_, new_n149_ );
not g075 ( new_n151_, N47 );
and g076 ( new_n152_, new_n151_, N43 );
or g077 ( new_n153_, new_n152_, keyIn_0_6 );
and g078 ( new_n154_, new_n152_, keyIn_0_6 );
not g079 ( new_n155_, new_n154_ );
and g080 ( new_n156_, new_n155_, new_n153_ );
not g081 ( new_n157_, new_n156_ );
not g082 ( new_n158_, keyIn_0_12 );
not g083 ( new_n159_, new_n97_ );
or g084 ( new_n160_, new_n101_, new_n159_ );
and g085 ( new_n161_, new_n160_, new_n158_ );
not g086 ( new_n162_, new_n161_ );
or g087 ( new_n163_, new_n160_, new_n158_ );
and g088 ( new_n164_, new_n162_, new_n157_, new_n163_ );
not g089 ( new_n165_, new_n88_ );
or g090 ( new_n166_, new_n101_, new_n165_ );
not g091 ( new_n167_, N99 );
and g092 ( new_n168_, keyIn_0_2, N95 );
not g093 ( new_n169_, new_n168_ );
or g094 ( new_n170_, keyIn_0_2, N95 );
and g095 ( new_n171_, new_n169_, new_n170_ );
and g096 ( new_n172_, new_n171_, new_n167_ );
and g097 ( new_n173_, new_n166_, new_n172_ );
or g098 ( new_n174_, new_n173_, keyIn_0_17 );
and g099 ( new_n175_, new_n166_, keyIn_0_17, new_n172_ );
not g100 ( new_n176_, new_n175_ );
and g101 ( new_n177_, new_n174_, new_n176_ );
or g102 ( new_n178_, new_n150_, new_n177_, new_n137_, new_n164_ );
not g103 ( new_n179_, keyIn_0_14 );
and g104 ( new_n180_, new_n80_, N108 );
or g105 ( new_n181_, new_n180_, new_n79_ );
not g106 ( new_n182_, new_n81_ );
and g107 ( new_n183_, new_n181_, new_n182_ );
or g108 ( new_n184_, new_n117_, new_n183_ );
and g109 ( new_n185_, new_n184_, new_n179_ );
not g110 ( new_n186_, new_n117_ );
and g111 ( new_n187_, new_n186_, keyIn_0_14, new_n82_ );
or g112 ( new_n188_, new_n185_, new_n187_ );
not g113 ( new_n189_, N112 );
and g114 ( new_n190_, new_n76_, keyIn_0_3 );
not g115 ( new_n191_, new_n190_ );
or g116 ( new_n192_, new_n76_, keyIn_0_3 );
and g117 ( new_n193_, new_n191_, new_n192_ );
and g118 ( new_n194_, new_n193_, new_n189_ );
and g119 ( new_n195_, new_n188_, new_n194_ );
or g120 ( new_n196_, new_n195_, keyIn_0_18 );
and g121 ( new_n197_, new_n195_, keyIn_0_18 );
not g122 ( new_n198_, new_n197_ );
and g123 ( new_n199_, new_n198_, new_n196_ );
not g124 ( new_n200_, N73 );
and g125 ( new_n201_, N223, new_n84_ );
not g126 ( new_n202_, new_n84_ );
and g127 ( new_n203_, new_n101_, new_n202_ );
or g128 ( new_n204_, new_n201_, new_n203_ );
and g129 ( new_n205_, new_n204_, keyIn_0_13 );
not g130 ( new_n206_, keyIn_0_13 );
or g131 ( new_n207_, new_n101_, new_n202_ );
not g132 ( new_n208_, new_n203_ );
and g133 ( new_n209_, new_n208_, new_n207_ );
and g134 ( new_n210_, new_n209_, new_n206_ );
or g135 ( new_n211_, new_n205_, new_n210_ );
and g136 ( new_n212_, new_n211_, N69, new_n200_ );
or g137 ( N329, new_n114_, new_n178_, new_n199_, new_n212_ );
and g138 ( new_n214_, N329, new_n126_ );
not g139 ( new_n215_, new_n214_ );
not g140 ( new_n216_, keyIn_0_16 );
not g141 ( new_n217_, new_n109_ );
or g142 ( new_n218_, new_n98_, N34 );
or g143 ( new_n219_, new_n217_, new_n218_ );
and g144 ( new_n220_, new_n219_, new_n216_ );
or g145 ( new_n221_, new_n220_, new_n112_ );
not g146 ( new_n222_, new_n199_ );
not g147 ( new_n223_, new_n212_ );
not g148 ( new_n224_, new_n126_ );
not g149 ( new_n225_, new_n137_ );
not g150 ( new_n226_, new_n150_ );
not g151 ( new_n227_, new_n164_ );
not g152 ( new_n228_, new_n177_ );
and g153 ( new_n229_, new_n226_, new_n228_, new_n225_, new_n227_ );
and g154 ( new_n230_, new_n229_, new_n224_ );
and g155 ( new_n231_, new_n230_, new_n221_, new_n222_, new_n223_ );
not g156 ( new_n232_, new_n231_ );
and g157 ( new_n233_, new_n215_, keyIn_0_22, new_n232_ );
not g158 ( new_n234_, keyIn_0_22 );
or g159 ( new_n235_, new_n214_, new_n231_ );
and g160 ( new_n236_, new_n235_, new_n234_ );
not g161 ( new_n237_, N14 );
and g162 ( new_n238_, new_n116_, new_n237_, new_n119_, new_n124_ );
not g163 ( new_n239_, new_n238_ );
or g164 ( new_n240_, new_n236_, new_n233_, new_n239_ );
not g165 ( new_n241_, keyIn_0_26 );
and g166 ( new_n242_, new_n221_, new_n229_, new_n222_, new_n223_ );
or g167 ( new_n243_, new_n242_, new_n150_ );
not g168 ( new_n244_, new_n243_ );
not g169 ( new_n245_, N27 );
and g170 ( new_n246_, new_n144_, new_n245_, new_n149_ );
not g171 ( new_n247_, new_n246_ );
or g172 ( new_n248_, new_n244_, new_n241_, new_n247_ );
not g173 ( new_n249_, new_n132_ );
or g174 ( new_n250_, new_n242_, new_n249_ );
or g175 ( new_n251_, new_n114_, new_n178_, new_n199_, new_n212_ );
and g176 ( new_n252_, new_n250_, new_n251_ );
or g177 ( new_n253_, new_n129_, new_n85_ );
not g178 ( new_n254_, new_n131_ );
or g179 ( new_n255_, new_n254_, new_n253_, N66 );
not g180 ( new_n256_, new_n255_ );
or g181 ( new_n257_, new_n256_, keyIn_0_21 );
not g182 ( new_n258_, keyIn_0_21 );
or g183 ( new_n259_, new_n255_, new_n258_ );
and g184 ( new_n260_, new_n257_, new_n259_ );
or g185 ( new_n261_, new_n252_, new_n260_ );
not g186 ( new_n262_, keyIn_0_23 );
and g187 ( new_n263_, new_n222_, new_n223_, new_n229_ );
not g188 ( new_n264_, new_n263_ );
and g189 ( new_n265_, new_n264_, new_n262_, new_n221_ );
not g190 ( new_n266_, keyIn_0_20 );
not g191 ( new_n267_, keyIn_0_5 );
not g192 ( new_n268_, N40 );
and g193 ( new_n269_, new_n267_, new_n268_, N30 );
or g194 ( new_n270_, new_n98_, N40 );
and g195 ( new_n271_, new_n270_, keyIn_0_5 );
or g196 ( new_n272_, new_n271_, new_n269_ );
and g197 ( new_n273_, new_n109_, new_n272_ );
or g198 ( new_n274_, new_n273_, new_n266_ );
and g199 ( new_n275_, new_n273_, new_n266_ );
not g200 ( new_n276_, new_n275_ );
and g201 ( new_n277_, new_n276_, new_n274_ );
or g202 ( new_n278_, new_n263_, new_n114_ );
and g203 ( new_n279_, new_n278_, keyIn_0_23 );
or g204 ( new_n280_, new_n279_, new_n265_, new_n277_ );
and g205 ( new_n281_, new_n261_, new_n248_, new_n280_ );
and g206 ( new_n282_, N329, N86 );
not g207 ( new_n283_, N92 );
and g208 ( new_n284_, new_n135_, N82, new_n283_ );
not g209 ( new_n285_, new_n284_ );
or g210 ( new_n286_, new_n282_, new_n285_ );
and g211 ( new_n287_, N329, new_n228_ );
not g212 ( new_n288_, new_n166_ );
not g213 ( new_n289_, keyIn_0_8 );
not g214 ( new_n290_, N105 );
and g215 ( new_n291_, new_n171_, new_n290_ );
not g216 ( new_n292_, new_n291_ );
or g217 ( new_n293_, new_n292_, new_n289_ );
or g218 ( new_n294_, new_n291_, keyIn_0_8 );
and g219 ( new_n295_, new_n293_, new_n294_ );
or g220 ( new_n296_, new_n288_, new_n295_ );
or g221 ( new_n297_, new_n287_, new_n296_ );
and g222 ( new_n298_, N329, N73 );
not g223 ( new_n299_, new_n211_ );
or g224 ( new_n300_, new_n299_, new_n83_, N79 );
or g225 ( new_n301_, new_n298_, new_n300_ );
and g226 ( new_n302_, new_n286_, new_n297_, new_n301_ );
and g227 ( new_n303_, new_n243_, new_n246_ );
or g228 ( new_n304_, new_n303_, keyIn_0_26 );
and g229 ( new_n305_, N329, new_n227_ );
not g230 ( new_n306_, new_n163_ );
not g231 ( new_n307_, N53 );
and g232 ( new_n308_, new_n307_, N43 );
or g233 ( new_n309_, new_n308_, keyIn_0_7 );
not g234 ( new_n310_, keyIn_0_7 );
or g235 ( new_n311_, new_n310_, new_n96_, N53 );
and g236 ( new_n312_, new_n309_, new_n311_ );
or g237 ( new_n313_, new_n306_, new_n161_, new_n312_ );
or g238 ( new_n314_, new_n305_, new_n313_ );
and g239 ( new_n315_, N329, new_n222_ );
not g240 ( new_n316_, N115 );
and g241 ( new_n317_, new_n188_, new_n316_, new_n193_ );
or g242 ( new_n318_, new_n317_, keyIn_0_19 );
and g243 ( new_n319_, new_n317_, keyIn_0_19 );
not g244 ( new_n320_, new_n319_ );
and g245 ( new_n321_, new_n320_, new_n318_ );
or g246 ( new_n322_, new_n315_, new_n321_ );
and g247 ( new_n323_, new_n314_, new_n322_ );
and g248 ( new_n324_, new_n302_, new_n304_, new_n323_ );
and g249 ( new_n325_, new_n324_, new_n240_, new_n281_ );
not g250 ( N370, new_n325_ );
not g251 ( new_n327_, keyIn_0_28 );
or g252 ( new_n328_, new_n325_, new_n268_ );
and g253 ( new_n329_, N329, N34 );
or g254 ( new_n330_, new_n101_, keyIn_0_9 );
and g255 ( new_n331_, new_n101_, keyIn_0_9 );
not g256 ( new_n332_, new_n331_ );
and g257 ( new_n333_, new_n332_, new_n330_ );
not g258 ( new_n334_, new_n333_ );
and g259 ( new_n335_, new_n334_, N24 );
or g260 ( new_n336_, new_n329_, new_n98_, new_n335_ );
not g261 ( new_n337_, new_n336_ );
and g262 ( new_n338_, new_n328_, new_n337_ );
not g263 ( new_n339_, new_n338_ );
and g264 ( new_n340_, new_n339_, new_n327_ );
and g265 ( new_n341_, new_n338_, keyIn_0_28 );
or g266 ( new_n342_, new_n340_, new_n341_ );
not g267 ( new_n343_, new_n342_ );
and g268 ( new_n344_, N370, N27 );
and g269 ( new_n345_, N329, N21 );
and g270 ( new_n346_, new_n334_, N11 );
or g271 ( new_n347_, new_n344_, new_n92_, new_n345_, new_n346_ );
not g272 ( new_n348_, new_n347_ );
or g273 ( new_n349_, new_n343_, new_n348_ );
and g274 ( new_n350_, N370, N53 );
not g275 ( new_n351_, new_n350_ );
and g276 ( new_n352_, N329, N47 );
not g277 ( new_n353_, new_n352_ );
and g278 ( new_n354_, new_n334_, N37 );
not g279 ( new_n355_, new_n354_ );
and g280 ( new_n356_, new_n351_, N43, new_n353_, new_n355_ );
not g281 ( new_n357_, new_n356_ );
and g282 ( new_n358_, N370, N66 );
and g283 ( new_n359_, N329, N60 );
and g284 ( new_n360_, new_n334_, N50 );
or g285 ( new_n361_, new_n358_, new_n85_, new_n359_, new_n360_ );
and g286 ( new_n362_, new_n357_, new_n361_ );
not g287 ( new_n363_, new_n362_ );
or g288 ( new_n364_, new_n349_, new_n363_ );
not g289 ( new_n365_, keyIn_0_27 );
not g290 ( new_n366_, N79 );
or g291 ( new_n367_, new_n325_, new_n366_ );
and g292 ( new_n368_, new_n367_, new_n365_ );
and g293 ( new_n369_, N370, keyIn_0_27, N79 );
or g294 ( new_n370_, new_n368_, new_n369_ );
not g295 ( new_n371_, new_n298_ );
and g296 ( new_n372_, new_n371_, keyIn_0_24 );
or g297 ( new_n373_, new_n371_, keyIn_0_24 );
not g298 ( new_n374_, new_n373_ );
and g299 ( new_n375_, new_n334_, N63 );
or g300 ( new_n376_, new_n374_, new_n372_, new_n83_, new_n375_ );
not g301 ( new_n377_, new_n376_ );
and g302 ( new_n378_, new_n370_, new_n377_ );
or g303 ( new_n379_, new_n378_, keyIn_0_29 );
and g304 ( new_n380_, new_n370_, keyIn_0_29, new_n377_ );
not g305 ( new_n381_, new_n380_ );
and g306 ( new_n382_, new_n379_, new_n381_ );
and g307 ( new_n383_, N370, N92 );
not g308 ( new_n384_, keyIn_0_15 );
and g309 ( new_n385_, new_n334_, N76 );
and g310 ( new_n386_, new_n385_, new_n384_ );
or g311 ( new_n387_, new_n385_, new_n384_ );
not g312 ( new_n388_, new_n387_ );
or g313 ( new_n389_, new_n282_, new_n89_, new_n386_, new_n388_ );
or g314 ( new_n390_, new_n383_, new_n389_ );
not g315 ( new_n391_, new_n390_ );
or g316 ( new_n392_, new_n325_, new_n290_ );
and g317 ( new_n393_, N329, N99 );
not g318 ( new_n394_, new_n393_ );
and g319 ( new_n395_, new_n394_, keyIn_0_25 );
or g320 ( new_n396_, new_n394_, keyIn_0_25 );
not g321 ( new_n397_, new_n396_ );
and g322 ( new_n398_, new_n334_, N89 );
or g323 ( new_n399_, new_n397_, new_n395_, new_n87_, new_n398_ );
not g324 ( new_n400_, new_n399_ );
and g325 ( new_n401_, new_n392_, new_n400_ );
or g326 ( new_n402_, new_n325_, new_n316_ );
or g327 ( new_n403_, new_n242_, new_n189_ );
or g328 ( new_n404_, new_n333_, new_n80_ );
and g329 ( new_n405_, new_n402_, N108, new_n403_, new_n404_ );
or g330 ( new_n406_, new_n391_, new_n401_, new_n405_ );
or g331 ( new_n407_, new_n364_, new_n382_, new_n406_ );
and g332 ( new_n408_, N370, N14 );
and g333 ( new_n409_, N329, N8 );
and g334 ( new_n410_, new_n334_, N1 );
or g335 ( new_n411_, new_n408_, new_n94_, new_n409_, new_n410_ );
and g336 ( N421, new_n407_, new_n411_ );
and g337 ( new_n413_, new_n364_, keyIn_0_30 );
not g338 ( new_n414_, keyIn_0_30 );
and g339 ( new_n415_, new_n362_, new_n342_, new_n414_, new_n347_ );
or g340 ( N430, new_n413_, new_n415_ );
and g341 ( new_n417_, new_n379_, new_n342_, new_n362_, new_n381_ );
and g342 ( new_n418_, new_n362_, new_n391_ );
or g343 ( N431, new_n417_, new_n349_, new_n418_ );
not g344 ( new_n420_, keyIn_0_31 );
and g345 ( new_n421_, new_n390_, new_n401_ );
or g346 ( new_n422_, new_n421_, new_n356_ );
and g347 ( new_n423_, new_n342_, new_n422_ );
or g348 ( new_n424_, new_n423_, new_n348_ );
or g349 ( new_n425_, new_n424_, new_n417_ );
and g350 ( new_n426_, new_n425_, new_n420_ );
not g351 ( new_n427_, new_n417_ );
not g352 ( new_n428_, new_n423_ );
and g353 ( new_n429_, new_n427_, keyIn_0_31, new_n347_, new_n428_ );
or g354 ( N432, new_n426_, new_n429_ );
endmodule