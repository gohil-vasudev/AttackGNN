module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n614_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n641_, new_n339_, new_n365_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n636_, new_n670_, new_n456_, new_n691_, new_n246_, new_n682_, new_n812_, new_n679_, new_n266_, new_n667_, new_n367_, new_n821_, new_n548_, new_n669_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n602_, new_n695_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n462_, new_n761_, new_n564_, new_n752_, new_n735_, new_n500_, new_n786_, new_n799_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n742_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n774_, new_n701_, new_n792_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n634_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n230_, new_n281_, new_n430_, new_n822_, new_n482_, new_n606_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n385_, new_n829_, new_n478_, new_n461_, new_n297_, new_n361_, new_n565_, new_n764_, new_n683_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n530_, new_n318_, new_n622_, new_n629_, new_n702_, new_n833_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n763_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n816_, new_n768_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n498_, new_n496_, new_n650_, new_n708_, new_n750_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n506_, new_n680_, new_n256_, new_n778_, new_n452_, new_n381_, new_n656_, new_n820_, new_n771_, new_n388_, new_n508_, new_n714_, new_n483_, new_n394_, new_n299_, new_n657_, new_n652_, new_n314_, new_n582_, new_n363_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n646_, new_n395_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n790_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n488_, new_n705_, new_n277_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n438_, new_n696_, new_n208_, new_n632_, new_n671_, new_n528_, new_n572_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n805_, new_n559_, new_n838_, new_n233_, new_n469_, new_n391_, new_n437_, new_n295_, new_n359_, new_n794_, new_n628_, new_n409_, new_n745_, new_n457_, new_n553_, new_n668_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n688_, new_n384_, new_n410_, new_n543_, new_n775_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n323_, new_n259_, new_n362_, new_n809_, new_n654_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n505_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n749_, new_n310_, new_n275_, new_n352_, new_n575_, new_n839_, new_n485_, new_n525_, new_n562_, new_n578_, new_n810_, new_n808_, new_n493_, new_n547_, new_n264_, new_n665_, new_n800_, new_n379_, new_n719_, new_n273_, new_n224_, new_n270_, new_n570_, new_n598_, new_n824_, new_n520_, new_n253_, new_n717_, new_n403_, new_n475_, new_n237_, new_n825_, new_n557_, new_n260_, new_n251_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n748_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n592_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n428_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n755_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n499_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n468_, new_n782_, new_n354_, new_n392_, new_n444_, new_n737_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n789_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n519_, new_n662_, new_n440_, new_n733_, new_n531_, new_n593_, new_n252_, new_n585_, new_n751_, new_n312_, new_n535_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n307_, new_n597_, new_n408_, new_n470_, new_n213_, new_n769_, new_n651_, new_n433_, new_n435_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n815_, new_n278_, new_n304_, new_n523_, new_n638_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n754_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n803_, new_n330_, new_n727_, new_n375_, new_n294_, new_n760_, new_n627_, new_n704_, new_n567_, new_n576_, new_n831_, new_n791_, new_n357_, new_n320_, new_n780_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n490_, new_n358_, new_n348_, new_n610_, new_n322_, new_n228_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n226_, new_n802_, new_n697_, new_n709_, new_n373_, new_n434_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n551_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n521_, new_n406_, new_n828_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n573_, new_n405_;

not g000 ( new_n202_, keyIn_0_78 );
not g001 ( new_n203_, keyIn_0_40 );
not g002 ( new_n204_, N93 );
nand g003 ( new_n205_, new_n204_, N89 );
not g004 ( new_n206_, N89 );
nand g005 ( new_n207_, new_n206_, N93 );
nand g006 ( new_n208_, new_n205_, new_n207_ );
nand g007 ( new_n209_, new_n208_, keyIn_0_6 );
not g008 ( new_n210_, keyIn_0_6 );
xnor g009 ( new_n211_, N89, N93 );
nand g010 ( new_n212_, new_n211_, new_n210_ );
nand g011 ( new_n213_, new_n209_, new_n212_ );
xnor g012 ( new_n214_, N81, N85 );
nand g013 ( new_n215_, new_n214_, keyIn_0_5 );
not g014 ( new_n216_, keyIn_0_5 );
and g015 ( new_n217_, N81, N85 );
nor g016 ( new_n218_, N81, N85 );
nor g017 ( new_n219_, new_n217_, new_n218_ );
nand g018 ( new_n220_, new_n219_, new_n216_ );
nand g019 ( new_n221_, new_n220_, new_n215_ );
nand g020 ( new_n222_, new_n213_, new_n221_ );
and g021 ( new_n223_, new_n209_, new_n212_ );
xnor g022 ( new_n224_, new_n214_, new_n216_ );
nand g023 ( new_n225_, new_n223_, new_n224_ );
nand g024 ( new_n226_, new_n225_, new_n222_ );
nand g025 ( new_n227_, new_n226_, keyIn_0_28 );
not g026 ( new_n228_, keyIn_0_28 );
and g027 ( new_n229_, new_n213_, new_n221_ );
nor g028 ( new_n230_, new_n213_, new_n221_ );
nor g029 ( new_n231_, new_n229_, new_n230_ );
nand g030 ( new_n232_, new_n231_, new_n228_ );
nand g031 ( new_n233_, new_n232_, new_n227_ );
xnor g032 ( new_n234_, N73, N77 );
xnor g033 ( new_n235_, N65, N69 );
xnor g034 ( new_n236_, new_n234_, new_n235_ );
not g035 ( new_n237_, new_n236_ );
nand g036 ( new_n238_, new_n233_, new_n237_ );
xnor g037 ( new_n239_, new_n226_, new_n228_ );
nand g038 ( new_n240_, new_n239_, new_n236_ );
nand g039 ( new_n241_, new_n240_, new_n238_ );
nand g040 ( new_n242_, new_n241_, keyIn_0_34 );
not g041 ( new_n243_, keyIn_0_34 );
xnor g042 ( new_n244_, new_n233_, new_n236_ );
nand g043 ( new_n245_, new_n244_, new_n243_ );
nand g044 ( new_n246_, new_n245_, new_n242_ );
nand g045 ( new_n247_, N129, N137 );
xnor g046 ( new_n248_, new_n247_, keyIn_0_9 );
not g047 ( new_n249_, new_n248_ );
nand g048 ( new_n250_, new_n246_, new_n249_ );
xnor g049 ( new_n251_, new_n241_, new_n243_ );
nand g050 ( new_n252_, new_n251_, new_n248_ );
nand g051 ( new_n253_, new_n252_, new_n250_ );
nand g052 ( new_n254_, new_n253_, keyIn_0_36 );
not g053 ( new_n255_, keyIn_0_36 );
xnor g054 ( new_n256_, new_n246_, new_n248_ );
nand g055 ( new_n257_, new_n256_, new_n255_ );
nand g056 ( new_n258_, new_n257_, new_n254_ );
xor g057 ( new_n259_, N33, N49 );
xnor g058 ( new_n260_, new_n259_, keyIn_0_16 );
xnor g059 ( new_n261_, N1, N17 );
xnor g060 ( new_n262_, new_n260_, new_n261_ );
not g061 ( new_n263_, new_n262_ );
nand g062 ( new_n264_, new_n258_, new_n263_ );
xnor g063 ( new_n265_, new_n253_, new_n255_ );
nand g064 ( new_n266_, new_n265_, new_n262_ );
nand g065 ( new_n267_, new_n266_, new_n264_ );
xnor g066 ( new_n268_, new_n267_, new_n203_ );
xnor g067 ( new_n269_, new_n268_, keyIn_0_49 );
xnor g068 ( new_n270_, N121, N125 );
xnor g069 ( new_n271_, new_n270_, keyIn_0_8 );
xnor g070 ( new_n272_, N113, N117 );
xnor g071 ( new_n273_, new_n271_, new_n272_ );
not g072 ( new_n274_, new_n273_ );
nand g073 ( new_n275_, new_n233_, new_n274_ );
nand g074 ( new_n276_, new_n239_, new_n273_ );
nand g075 ( new_n277_, new_n276_, new_n275_ );
nand g076 ( new_n278_, N132, N137 );
xnor g077 ( new_n279_, new_n278_, keyIn_0_12 );
not g078 ( new_n280_, new_n279_ );
nand g079 ( new_n281_, new_n277_, new_n280_ );
xnor g080 ( new_n282_, new_n233_, new_n273_ );
nand g081 ( new_n283_, new_n282_, new_n279_ );
nand g082 ( new_n284_, new_n283_, new_n281_ );
nand g083 ( new_n285_, new_n284_, keyIn_0_37 );
not g084 ( new_n286_, keyIn_0_37 );
xnor g085 ( new_n287_, new_n277_, new_n279_ );
nand g086 ( new_n288_, new_n287_, new_n286_ );
nand g087 ( new_n289_, new_n288_, new_n285_ );
xor g088 ( new_n290_, N13, N29 );
xnor g089 ( new_n291_, new_n290_, keyIn_0_20 );
xor g090 ( new_n292_, N45, N61 );
xnor g091 ( new_n293_, new_n291_, new_n292_ );
xor g092 ( new_n294_, new_n293_, keyIn_0_30 );
not g093 ( new_n295_, new_n294_ );
nand g094 ( new_n296_, new_n289_, new_n295_ );
xnor g095 ( new_n297_, new_n284_, new_n286_ );
nand g096 ( new_n298_, new_n297_, new_n294_ );
nand g097 ( new_n299_, new_n298_, new_n296_ );
nand g098 ( new_n300_, new_n299_, keyIn_0_41 );
not g099 ( new_n301_, keyIn_0_41 );
xnor g100 ( new_n302_, new_n289_, new_n294_ );
nand g101 ( new_n303_, new_n302_, new_n301_ );
nand g102 ( new_n304_, new_n303_, new_n300_ );
xnor g103 ( new_n305_, N105, N109 );
xnor g104 ( new_n306_, new_n305_, keyIn_0_7 );
xor g105 ( new_n307_, N97, N101 );
xnor g106 ( new_n308_, new_n306_, new_n307_ );
xnor g107 ( new_n309_, new_n308_, new_n236_ );
nand g108 ( new_n310_, N131, N137 );
xor g109 ( new_n311_, new_n310_, keyIn_0_11 );
xnor g110 ( new_n312_, new_n309_, new_n311_ );
xor g111 ( new_n313_, N41, N57 );
xnor g112 ( new_n314_, new_n313_, keyIn_0_19 );
xor g113 ( new_n315_, N9, N25 );
xnor g114 ( new_n316_, new_n314_, new_n315_ );
xor g115 ( new_n317_, new_n316_, keyIn_0_29 );
xnor g116 ( new_n318_, new_n312_, new_n317_ );
xnor g117 ( new_n319_, new_n308_, new_n273_ );
xnor g118 ( new_n320_, new_n319_, keyIn_0_35 );
nand g119 ( new_n321_, N130, N137 );
xor g120 ( new_n322_, new_n321_, keyIn_0_10 );
xnor g121 ( new_n323_, new_n320_, new_n322_ );
xor g122 ( new_n324_, N37, N53 );
xnor g123 ( new_n325_, new_n324_, keyIn_0_18 );
xor g124 ( new_n326_, N5, N21 );
xnor g125 ( new_n327_, new_n326_, keyIn_0_17 );
xnor g126 ( new_n328_, new_n327_, new_n325_ );
xnor g127 ( new_n329_, new_n323_, new_n328_ );
xnor g128 ( new_n330_, new_n329_, keyIn_0_50 );
nand g129 ( new_n331_, new_n330_, new_n318_ );
nor g130 ( new_n332_, new_n331_, new_n304_ );
nand g131 ( new_n333_, new_n269_, new_n332_ );
xnor g132 ( new_n334_, new_n333_, keyIn_0_73 );
nand g133 ( new_n335_, new_n267_, keyIn_0_40 );
xnor g134 ( new_n336_, new_n258_, new_n262_ );
nand g135 ( new_n337_, new_n336_, new_n203_ );
nand g136 ( new_n338_, new_n337_, new_n335_ );
xnor g137 ( new_n339_, new_n338_, keyIn_0_46 );
xnor g138 ( new_n340_, new_n299_, new_n301_ );
not g139 ( new_n341_, new_n329_ );
nand g140 ( new_n342_, new_n341_, keyIn_0_47 );
nor g141 ( new_n343_, new_n341_, keyIn_0_47 );
xnor g142 ( new_n344_, new_n318_, keyIn_0_48 );
nor g143 ( new_n345_, new_n343_, new_n344_ );
nand g144 ( new_n346_, new_n345_, new_n342_ );
nor g145 ( new_n347_, new_n346_, new_n340_ );
not g146 ( new_n348_, new_n347_ );
nor g147 ( new_n349_, new_n339_, new_n348_ );
nand g148 ( new_n350_, new_n349_, keyIn_0_72 );
not g149 ( new_n351_, keyIn_0_72 );
not g150 ( new_n352_, keyIn_0_46 );
nand g151 ( new_n353_, new_n338_, new_n352_ );
nand g152 ( new_n354_, new_n268_, keyIn_0_46 );
nand g153 ( new_n355_, new_n354_, new_n353_ );
nand g154 ( new_n356_, new_n355_, new_n347_ );
nand g155 ( new_n357_, new_n356_, new_n351_ );
nand g156 ( new_n358_, new_n350_, new_n357_ );
nor g157 ( new_n359_, new_n341_, new_n318_ );
nand g158 ( new_n360_, new_n340_, new_n359_ );
nor g159 ( new_n361_, new_n268_, new_n360_ );
xnor g160 ( new_n362_, new_n361_, keyIn_0_75 );
nor g161 ( new_n363_, new_n338_, new_n329_ );
nor g162 ( new_n364_, new_n340_, keyIn_0_52 );
nand g163 ( new_n365_, new_n340_, keyIn_0_52 );
xnor g164 ( new_n366_, new_n318_, keyIn_0_51 );
not g165 ( new_n367_, new_n366_ );
nand g166 ( new_n368_, new_n365_, new_n367_ );
nor g167 ( new_n369_, new_n368_, new_n364_ );
nand g168 ( new_n370_, new_n363_, new_n369_ );
nand g169 ( new_n371_, new_n370_, keyIn_0_74 );
not g170 ( new_n372_, keyIn_0_74 );
nand g171 ( new_n373_, new_n268_, new_n341_ );
not g172 ( new_n374_, new_n364_ );
not g173 ( new_n375_, keyIn_0_52 );
nor g174 ( new_n376_, new_n304_, new_n375_ );
nor g175 ( new_n377_, new_n376_, new_n366_ );
nand g176 ( new_n378_, new_n377_, new_n374_ );
nor g177 ( new_n379_, new_n373_, new_n378_ );
nand g178 ( new_n380_, new_n379_, new_n372_ );
nand g179 ( new_n381_, new_n380_, new_n371_ );
nor g180 ( new_n382_, new_n381_, new_n362_ );
nand g181 ( new_n383_, new_n382_, new_n358_ );
nor g182 ( new_n384_, new_n383_, new_n334_ );
nand g183 ( new_n385_, new_n384_, new_n202_ );
xor g184 ( new_n386_, new_n333_, keyIn_0_73 );
xnor g185 ( new_n387_, new_n356_, keyIn_0_72 );
not g186 ( new_n388_, new_n362_ );
xnor g187 ( new_n389_, new_n370_, new_n372_ );
nand g188 ( new_n390_, new_n389_, new_n388_ );
nor g189 ( new_n391_, new_n390_, new_n387_ );
nand g190 ( new_n392_, new_n391_, new_n386_ );
nand g191 ( new_n393_, new_n392_, keyIn_0_78 );
nand g192 ( new_n394_, new_n393_, new_n385_ );
not g193 ( new_n395_, keyIn_0_43 );
not g194 ( new_n396_, keyIn_0_39 );
xnor g195 ( new_n397_, N41, N45 );
xor g196 ( new_n398_, N33, N37 );
xnor g197 ( new_n399_, keyIn_0_1, keyIn_0_2 );
xnor g198 ( new_n400_, new_n398_, new_n399_ );
xnor g199 ( new_n401_, new_n400_, new_n397_ );
nand g200 ( new_n402_, new_n401_, keyIn_0_26 );
not g201 ( new_n403_, keyIn_0_26 );
not g202 ( new_n404_, new_n397_ );
xnor g203 ( new_n405_, new_n400_, new_n404_ );
nand g204 ( new_n406_, new_n405_, new_n403_ );
nand g205 ( new_n407_, new_n402_, new_n406_ );
xnor g206 ( new_n408_, N49, N53 );
xor g207 ( new_n409_, N57, N61 );
xnor g208 ( new_n410_, keyIn_0_3, keyIn_0_4 );
xnor g209 ( new_n411_, new_n409_, new_n410_ );
xnor g210 ( new_n412_, new_n411_, new_n408_ );
nand g211 ( new_n413_, new_n412_, keyIn_0_27 );
not g212 ( new_n414_, keyIn_0_27 );
not g213 ( new_n415_, new_n408_ );
xnor g214 ( new_n416_, new_n411_, new_n415_ );
nand g215 ( new_n417_, new_n416_, new_n414_ );
nand g216 ( new_n418_, new_n413_, new_n417_ );
xnor g217 ( new_n419_, new_n407_, new_n418_ );
nand g218 ( new_n420_, new_n419_, keyIn_0_33 );
not g219 ( new_n421_, keyIn_0_33 );
and g220 ( new_n422_, new_n407_, new_n418_ );
nor g221 ( new_n423_, new_n407_, new_n418_ );
nor g222 ( new_n424_, new_n422_, new_n423_ );
nand g223 ( new_n425_, new_n424_, new_n421_ );
nand g224 ( new_n426_, new_n425_, new_n420_ );
nand g225 ( new_n427_, N134, N137 );
xnor g226 ( new_n428_, new_n427_, keyIn_0_14 );
not g227 ( new_n429_, new_n428_ );
nand g228 ( new_n430_, new_n426_, new_n429_ );
and g229 ( new_n431_, new_n425_, new_n420_ );
nand g230 ( new_n432_, new_n431_, new_n428_ );
nand g231 ( new_n433_, new_n432_, new_n430_ );
nand g232 ( new_n434_, new_n433_, new_n396_ );
xnor g233 ( new_n435_, new_n426_, new_n428_ );
nand g234 ( new_n436_, new_n435_, keyIn_0_39 );
nand g235 ( new_n437_, new_n436_, new_n434_ );
xor g236 ( new_n438_, N69, N85 );
xnor g237 ( new_n439_, new_n438_, keyIn_0_23 );
xor g238 ( new_n440_, N101, N117 );
xnor g239 ( new_n441_, new_n440_, keyIn_0_24 );
xnor g240 ( new_n442_, new_n439_, new_n441_ );
nand g241 ( new_n443_, new_n437_, new_n442_ );
xnor g242 ( new_n444_, new_n433_, keyIn_0_39 );
not g243 ( new_n445_, new_n442_ );
nand g244 ( new_n446_, new_n444_, new_n445_ );
nand g245 ( new_n447_, new_n446_, new_n443_ );
nand g246 ( new_n448_, new_n447_, new_n395_ );
xnor g247 ( new_n449_, new_n437_, new_n445_ );
nand g248 ( new_n450_, new_n449_, keyIn_0_43 );
nand g249 ( new_n451_, new_n450_, new_n448_ );
xor g250 ( new_n452_, new_n451_, keyIn_0_53 );
xor g251 ( new_n453_, N17, N21 );
xnor g252 ( new_n454_, N25, N29 );
xnor g253 ( new_n455_, new_n454_, keyIn_0_0 );
xnor g254 ( new_n456_, new_n455_, new_n453_ );
xnor g255 ( new_n457_, new_n456_, keyIn_0_25 );
xnor g256 ( new_n458_, N9, N13 );
xnor g257 ( new_n459_, N1, N5 );
xnor g258 ( new_n460_, new_n458_, new_n459_ );
xnor g259 ( new_n461_, new_n457_, new_n460_ );
nand g260 ( new_n462_, N133, N137 );
xnor g261 ( new_n463_, new_n462_, keyIn_0_13 );
xnor g262 ( new_n464_, new_n461_, new_n463_ );
xnor g263 ( new_n465_, new_n464_, keyIn_0_38 );
xor g264 ( new_n466_, N97, N113 );
xnor g265 ( new_n467_, new_n466_, keyIn_0_22 );
xor g266 ( new_n468_, N65, N81 );
xnor g267 ( new_n469_, new_n468_, keyIn_0_21 );
xor g268 ( new_n470_, new_n467_, new_n469_ );
not g269 ( new_n471_, new_n470_ );
nand g270 ( new_n472_, new_n465_, new_n471_ );
not g271 ( new_n473_, keyIn_0_38 );
xnor g272 ( new_n474_, new_n464_, new_n473_ );
nand g273 ( new_n475_, new_n474_, new_n470_ );
nand g274 ( new_n476_, new_n472_, new_n475_ );
xnor g275 ( new_n477_, new_n476_, keyIn_0_42 );
not g276 ( new_n478_, keyIn_0_45 );
xor g277 ( new_n479_, new_n418_, new_n457_ );
nand g278 ( new_n480_, N136, N137 );
xor g279 ( new_n481_, new_n480_, keyIn_0_15 );
xnor g280 ( new_n482_, new_n479_, new_n481_ );
xor g281 ( new_n483_, N109, N125 );
xnor g282 ( new_n484_, N77, N93 );
xnor g283 ( new_n485_, new_n483_, new_n484_ );
xor g284 ( new_n486_, new_n485_, keyIn_0_32 );
xnor g285 ( new_n487_, new_n482_, new_n486_ );
xnor g286 ( new_n488_, new_n487_, new_n478_ );
nor g287 ( new_n489_, new_n488_, keyIn_0_54 );
not g288 ( new_n490_, keyIn_0_44 );
xnor g289 ( new_n491_, new_n407_, new_n460_ );
nand g290 ( new_n492_, N135, N137 );
xnor g291 ( new_n493_, new_n491_, new_n492_ );
xor g292 ( new_n494_, N105, N121 );
xnor g293 ( new_n495_, N73, N89 );
xnor g294 ( new_n496_, new_n494_, new_n495_ );
xor g295 ( new_n497_, new_n496_, keyIn_0_31 );
not g296 ( new_n498_, new_n497_ );
xnor g297 ( new_n499_, new_n493_, new_n498_ );
nand g298 ( new_n500_, new_n499_, new_n490_ );
xnor g299 ( new_n501_, new_n493_, new_n497_ );
nand g300 ( new_n502_, new_n501_, keyIn_0_44 );
nand g301 ( new_n503_, new_n500_, new_n502_ );
not g302 ( new_n504_, new_n503_ );
nand g303 ( new_n505_, new_n488_, keyIn_0_54 );
nand g304 ( new_n506_, new_n505_, new_n504_ );
nor g305 ( new_n507_, new_n506_, new_n489_ );
and g306 ( new_n508_, new_n507_, new_n477_ );
nand g307 ( new_n509_, new_n452_, new_n508_ );
nor g308 ( new_n510_, new_n509_, new_n268_ );
nand g309 ( new_n511_, new_n394_, new_n510_ );
xnor g310 ( new_n512_, new_n511_, N1 );
xor g311 ( N724, new_n512_, keyIn_0_107 );
nor g312 ( new_n514_, new_n509_, new_n329_ );
nand g313 ( new_n515_, new_n394_, new_n514_ );
xnor g314 ( new_n516_, new_n515_, keyIn_0_86 );
xnor g315 ( new_n517_, new_n516_, N5 );
xnor g316 ( N725, new_n517_, keyIn_0_108 );
not g317 ( new_n519_, new_n318_ );
nor g318 ( new_n520_, new_n509_, new_n519_ );
nand g319 ( new_n521_, new_n394_, new_n520_ );
xnor g320 ( new_n522_, new_n521_, keyIn_0_87 );
xnor g321 ( new_n523_, new_n522_, N9 );
xor g322 ( N726, new_n523_, keyIn_0_109 );
nor g323 ( new_n525_, new_n509_, new_n340_ );
nand g324 ( new_n526_, new_n394_, new_n525_ );
xnor g325 ( new_n527_, new_n526_, keyIn_0_88 );
xnor g326 ( new_n528_, new_n527_, N13 );
xor g327 ( N727, new_n528_, keyIn_0_110 );
xor g328 ( new_n530_, new_n451_, keyIn_0_55 );
nor g329 ( new_n531_, new_n488_, new_n504_ );
nand g330 ( new_n532_, new_n477_, new_n531_ );
nor g331 ( new_n533_, new_n530_, new_n532_ );
nand g332 ( new_n534_, new_n394_, new_n533_ );
xor g333 ( new_n535_, new_n534_, keyIn_0_80 );
not g334 ( new_n536_, new_n535_ );
nand g335 ( new_n537_, new_n536_, new_n338_ );
xnor g336 ( N728, new_n537_, N17 );
nand g337 ( new_n539_, new_n536_, new_n341_ );
xnor g338 ( N729, new_n539_, N21 );
nand g339 ( new_n541_, new_n536_, new_n318_ );
xnor g340 ( N730, new_n541_, N25 );
nand g341 ( new_n543_, new_n536_, new_n304_ );
xnor g342 ( new_n544_, new_n543_, N29 );
xnor g343 ( N731, new_n544_, keyIn_0_111 );
nand g344 ( new_n546_, new_n477_, keyIn_0_56 );
nor g345 ( new_n547_, new_n477_, keyIn_0_56 );
nand g346 ( new_n548_, new_n488_, new_n504_ );
nor g347 ( new_n549_, new_n547_, new_n548_ );
nand g348 ( new_n550_, new_n549_, new_n546_ );
nor g349 ( new_n551_, new_n550_, new_n451_ );
nand g350 ( new_n552_, new_n394_, new_n551_ );
nor g351 ( new_n553_, new_n552_, new_n268_ );
xnor g352 ( new_n554_, new_n553_, keyIn_0_89 );
xor g353 ( new_n555_, new_n554_, N33 );
xnor g354 ( N732, new_n555_, keyIn_0_112 );
nor g355 ( new_n557_, new_n552_, new_n329_ );
xnor g356 ( new_n558_, new_n557_, keyIn_0_90 );
xnor g357 ( new_n559_, new_n558_, N37 );
xnor g358 ( N733, new_n559_, keyIn_0_113 );
nor g359 ( new_n561_, new_n552_, new_n519_ );
xor g360 ( new_n562_, new_n561_, keyIn_0_91 );
xnor g361 ( N734, new_n562_, N41 );
nor g362 ( new_n564_, new_n552_, new_n340_ );
xnor g363 ( new_n565_, new_n564_, N45 );
xnor g364 ( N735, new_n565_, keyIn_0_114 );
not g365 ( new_n567_, keyIn_0_81 );
not g366 ( new_n568_, keyIn_0_57 );
not g367 ( new_n569_, keyIn_0_42 );
xnor g368 ( new_n570_, new_n476_, new_n569_ );
nand g369 ( new_n571_, new_n570_, new_n568_ );
nor g370 ( new_n572_, new_n570_, new_n568_ );
xnor g371 ( new_n573_, new_n487_, keyIn_0_45 );
xor g372 ( new_n574_, new_n503_, keyIn_0_58 );
nand g373 ( new_n575_, new_n574_, new_n573_ );
nor g374 ( new_n576_, new_n575_, new_n572_ );
nand g375 ( new_n577_, new_n576_, new_n571_ );
nor g376 ( new_n578_, new_n577_, new_n451_ );
nand g377 ( new_n579_, new_n394_, new_n578_ );
xnor g378 ( new_n580_, new_n579_, new_n567_ );
nand g379 ( new_n581_, new_n580_, new_n338_ );
xnor g380 ( new_n582_, new_n581_, keyIn_0_92 );
xnor g381 ( N736, new_n582_, N49 );
nand g382 ( new_n584_, new_n580_, new_n341_ );
xnor g383 ( new_n585_, new_n584_, keyIn_0_93 );
xnor g384 ( N737, new_n585_, N53 );
not g385 ( new_n587_, keyIn_0_115 );
xnor g386 ( new_n588_, new_n579_, keyIn_0_81 );
nor g387 ( new_n589_, new_n588_, new_n519_ );
nand g388 ( new_n590_, new_n589_, keyIn_0_94 );
not g389 ( new_n591_, keyIn_0_94 );
nand g390 ( new_n592_, new_n580_, new_n318_ );
nand g391 ( new_n593_, new_n592_, new_n591_ );
nand g392 ( new_n594_, new_n590_, new_n593_ );
nand g393 ( new_n595_, new_n594_, N57 );
not g394 ( new_n596_, N57 );
xnor g395 ( new_n597_, new_n592_, keyIn_0_94 );
nand g396 ( new_n598_, new_n597_, new_n596_ );
nand g397 ( new_n599_, new_n598_, new_n595_ );
nand g398 ( new_n600_, new_n599_, new_n587_ );
xnor g399 ( new_n601_, new_n594_, new_n596_ );
nand g400 ( new_n602_, new_n601_, keyIn_0_115 );
nand g401 ( N738, new_n602_, new_n600_ );
nor g402 ( new_n604_, new_n588_, new_n340_ );
nand g403 ( new_n605_, new_n604_, keyIn_0_95 );
not g404 ( new_n606_, keyIn_0_95 );
nand g405 ( new_n607_, new_n580_, new_n304_ );
nand g406 ( new_n608_, new_n607_, new_n606_ );
nand g407 ( new_n609_, new_n605_, new_n608_ );
nand g408 ( new_n610_, new_n609_, N61 );
not g409 ( new_n611_, N61 );
xnor g410 ( new_n612_, new_n607_, keyIn_0_95 );
nand g411 ( new_n613_, new_n612_, new_n611_ );
nand g412 ( new_n614_, new_n613_, new_n610_ );
nand g413 ( new_n615_, new_n614_, keyIn_0_116 );
not g414 ( new_n616_, keyIn_0_116 );
xnor g415 ( new_n617_, new_n609_, new_n611_ );
nand g416 ( new_n618_, new_n617_, new_n616_ );
nand g417 ( N739, new_n618_, new_n615_ );
not g418 ( new_n620_, keyIn_0_117 );
not g419 ( new_n621_, keyIn_0_96 );
not g420 ( new_n622_, keyIn_0_79 );
nor g421 ( new_n623_, new_n451_, keyIn_0_59 );
nand g422 ( new_n624_, new_n451_, keyIn_0_59 );
xnor g423 ( new_n625_, new_n503_, keyIn_0_60 );
nand g424 ( new_n626_, new_n570_, new_n573_ );
nor g425 ( new_n627_, new_n626_, new_n625_ );
nand g426 ( new_n628_, new_n624_, new_n627_ );
nor g427 ( new_n629_, new_n628_, new_n623_ );
xnor g428 ( new_n630_, new_n629_, keyIn_0_76 );
xnor g429 ( new_n631_, new_n477_, keyIn_0_62 );
not g430 ( new_n632_, new_n451_ );
xnor g431 ( new_n633_, new_n573_, keyIn_0_64 );
xor g432 ( new_n634_, new_n503_, keyIn_0_63 );
nor g433 ( new_n635_, new_n633_, new_n634_ );
nand g434 ( new_n636_, new_n632_, new_n635_ );
nor g435 ( new_n637_, new_n636_, new_n631_ );
nor g436 ( new_n638_, new_n573_, keyIn_0_61 );
nand g437 ( new_n639_, new_n573_, keyIn_0_61 );
nand g438 ( new_n640_, new_n639_, new_n504_ );
nor g439 ( new_n641_, new_n640_, new_n638_ );
nand g440 ( new_n642_, new_n641_, new_n570_ );
nor g441 ( new_n643_, new_n642_, new_n632_ );
nor g442 ( new_n644_, new_n637_, new_n643_ );
xnor g443 ( new_n645_, new_n488_, keyIn_0_66 );
not g444 ( new_n646_, keyIn_0_65 );
xnor g445 ( new_n647_, new_n503_, new_n646_ );
nand g446 ( new_n648_, new_n647_, new_n477_ );
nor g447 ( new_n649_, new_n645_, new_n648_ );
nand g448 ( new_n650_, new_n649_, new_n451_ );
xnor g449 ( new_n651_, new_n650_, keyIn_0_77 );
nand g450 ( new_n652_, new_n651_, new_n644_ );
nor g451 ( new_n653_, new_n630_, new_n652_ );
nand g452 ( new_n654_, new_n653_, new_n622_ );
not g453 ( new_n655_, keyIn_0_76 );
xnor g454 ( new_n656_, new_n629_, new_n655_ );
not g455 ( new_n657_, new_n631_ );
and g456 ( new_n658_, new_n632_, new_n635_ );
nand g457 ( new_n659_, new_n658_, new_n657_ );
not g458 ( new_n660_, new_n643_ );
nand g459 ( new_n661_, new_n659_, new_n660_ );
not g460 ( new_n662_, keyIn_0_77 );
xnor g461 ( new_n663_, new_n650_, new_n662_ );
nor g462 ( new_n664_, new_n663_, new_n661_ );
nand g463 ( new_n665_, new_n656_, new_n664_ );
nand g464 ( new_n666_, new_n665_, keyIn_0_79 );
nand g465 ( new_n667_, new_n654_, new_n666_ );
nand g466 ( new_n668_, new_n304_, keyIn_0_68 );
nor g467 ( new_n669_, new_n304_, keyIn_0_68 );
nor g468 ( new_n670_, new_n329_, keyIn_0_67 );
nand g469 ( new_n671_, new_n329_, keyIn_0_67 );
nand g470 ( new_n672_, new_n671_, new_n318_ );
or g471 ( new_n673_, new_n672_, new_n670_ );
nor g472 ( new_n674_, new_n669_, new_n673_ );
nand g473 ( new_n675_, new_n674_, new_n668_ );
nor g474 ( new_n676_, new_n675_, new_n268_ );
nand g475 ( new_n677_, new_n667_, new_n676_ );
xnor g476 ( new_n678_, new_n677_, keyIn_0_82 );
nor g477 ( new_n679_, new_n678_, new_n570_ );
nand g478 ( new_n680_, new_n679_, new_n621_ );
not g479 ( new_n681_, keyIn_0_82 );
xnor g480 ( new_n682_, new_n677_, new_n681_ );
nand g481 ( new_n683_, new_n682_, new_n477_ );
nand g482 ( new_n684_, new_n683_, keyIn_0_96 );
nand g483 ( new_n685_, new_n680_, new_n684_ );
nand g484 ( new_n686_, new_n685_, N65 );
not g485 ( new_n687_, N65 );
xnor g486 ( new_n688_, new_n683_, new_n621_ );
nand g487 ( new_n689_, new_n688_, new_n687_ );
nand g488 ( new_n690_, new_n689_, new_n686_ );
nand g489 ( new_n691_, new_n690_, new_n620_ );
xnor g490 ( new_n692_, new_n685_, new_n687_ );
nand g491 ( new_n693_, new_n692_, keyIn_0_117 );
nand g492 ( N740, new_n693_, new_n691_ );
not g493 ( new_n695_, keyIn_0_118 );
nor g494 ( new_n696_, new_n678_, new_n451_ );
nand g495 ( new_n697_, new_n696_, keyIn_0_97 );
not g496 ( new_n698_, keyIn_0_97 );
nand g497 ( new_n699_, new_n682_, new_n632_ );
nand g498 ( new_n700_, new_n699_, new_n698_ );
nand g499 ( new_n701_, new_n697_, new_n700_ );
nand g500 ( new_n702_, new_n701_, N69 );
not g501 ( new_n703_, N69 );
xnor g502 ( new_n704_, new_n699_, keyIn_0_97 );
nand g503 ( new_n705_, new_n704_, new_n703_ );
nand g504 ( new_n706_, new_n705_, new_n702_ );
nand g505 ( new_n707_, new_n706_, new_n695_ );
xnor g506 ( new_n708_, new_n701_, new_n703_ );
nand g507 ( new_n709_, new_n708_, keyIn_0_118 );
nand g508 ( N741, new_n709_, new_n707_ );
nand g509 ( new_n711_, new_n682_, new_n504_ );
xnor g510 ( new_n712_, new_n711_, keyIn_0_98 );
xor g511 ( N742, new_n712_, N73 );
nand g512 ( new_n714_, new_n682_, new_n573_ );
xnor g513 ( new_n715_, new_n714_, N77 );
xor g514 ( N743, new_n715_, keyIn_0_119 );
not g515 ( new_n717_, keyIn_0_83 );
not g516 ( new_n718_, keyIn_0_69 );
nor g517 ( new_n719_, new_n341_, new_n718_ );
nand g518 ( new_n720_, new_n341_, new_n718_ );
xnor g519 ( new_n721_, new_n318_, keyIn_0_70 );
nand g520 ( new_n722_, new_n720_, new_n721_ );
nor g521 ( new_n723_, new_n722_, new_n719_ );
nand g522 ( new_n724_, new_n723_, new_n304_ );
nor g523 ( new_n725_, new_n268_, new_n724_ );
nand g524 ( new_n726_, new_n667_, new_n725_ );
xnor g525 ( new_n727_, new_n726_, new_n717_ );
nor g526 ( new_n728_, new_n727_, new_n570_ );
nand g527 ( new_n729_, new_n728_, keyIn_0_99 );
not g528 ( new_n730_, keyIn_0_99 );
xnor g529 ( new_n731_, new_n726_, keyIn_0_83 );
nand g530 ( new_n732_, new_n731_, new_n477_ );
nand g531 ( new_n733_, new_n732_, new_n730_ );
nand g532 ( new_n734_, new_n729_, new_n733_ );
nand g533 ( new_n735_, new_n734_, N81 );
not g534 ( new_n736_, N81 );
xnor g535 ( new_n737_, new_n732_, keyIn_0_99 );
nand g536 ( new_n738_, new_n737_, new_n736_ );
nand g537 ( new_n739_, new_n738_, new_n735_ );
nand g538 ( new_n740_, new_n739_, keyIn_0_120 );
not g539 ( new_n741_, keyIn_0_120 );
xnor g540 ( new_n742_, new_n734_, new_n736_ );
nand g541 ( new_n743_, new_n742_, new_n741_ );
nand g542 ( N744, new_n743_, new_n740_ );
nand g543 ( new_n745_, new_n731_, new_n632_ );
xnor g544 ( new_n746_, new_n745_, N85 );
xnor g545 ( N745, new_n746_, keyIn_0_121 );
nor g546 ( new_n748_, new_n727_, new_n503_ );
nand g547 ( new_n749_, new_n748_, keyIn_0_100 );
not g548 ( new_n750_, keyIn_0_100 );
nand g549 ( new_n751_, new_n731_, new_n504_ );
nand g550 ( new_n752_, new_n751_, new_n750_ );
nand g551 ( new_n753_, new_n749_, new_n752_ );
nand g552 ( new_n754_, new_n753_, N89 );
xnor g553 ( new_n755_, new_n751_, keyIn_0_100 );
nand g554 ( new_n756_, new_n755_, new_n206_ );
nand g555 ( new_n757_, new_n756_, new_n754_ );
nand g556 ( new_n758_, new_n757_, keyIn_0_122 );
not g557 ( new_n759_, keyIn_0_122 );
xnor g558 ( new_n760_, new_n753_, new_n206_ );
nand g559 ( new_n761_, new_n760_, new_n759_ );
nand g560 ( N746, new_n761_, new_n758_ );
nand g561 ( new_n763_, new_n731_, new_n573_ );
xnor g562 ( new_n764_, new_n763_, keyIn_0_101 );
xnor g563 ( N747, new_n764_, new_n204_ );
not g564 ( new_n766_, keyIn_0_84 );
nand g565 ( new_n767_, new_n340_, new_n318_ );
nor g566 ( new_n768_, new_n373_, new_n767_ );
nand g567 ( new_n769_, new_n667_, new_n768_ );
xnor g568 ( new_n770_, new_n769_, new_n766_ );
nand g569 ( new_n771_, new_n770_, new_n477_ );
xnor g570 ( new_n772_, new_n771_, keyIn_0_102 );
xor g571 ( N748, new_n772_, N97 );
nand g572 ( new_n774_, new_n770_, new_n632_ );
xnor g573 ( new_n775_, new_n774_, keyIn_0_103 );
xor g574 ( N749, new_n775_, N101 );
xnor g575 ( new_n777_, new_n769_, keyIn_0_84 );
nor g576 ( new_n778_, new_n777_, new_n503_ );
nand g577 ( new_n779_, new_n778_, keyIn_0_104 );
not g578 ( new_n780_, keyIn_0_104 );
nand g579 ( new_n781_, new_n770_, new_n504_ );
nand g580 ( new_n782_, new_n781_, new_n780_ );
nand g581 ( new_n783_, new_n779_, new_n782_ );
nand g582 ( new_n784_, new_n783_, N105 );
not g583 ( new_n785_, N105 );
xnor g584 ( new_n786_, new_n781_, keyIn_0_104 );
nand g585 ( new_n787_, new_n786_, new_n785_ );
nand g586 ( new_n788_, new_n787_, new_n784_ );
nand g587 ( new_n789_, new_n788_, keyIn_0_123 );
not g588 ( new_n790_, keyIn_0_123 );
xnor g589 ( new_n791_, new_n783_, new_n785_ );
nand g590 ( new_n792_, new_n791_, new_n790_ );
nand g591 ( N750, new_n792_, new_n789_ );
nand g592 ( new_n794_, new_n770_, new_n573_ );
xnor g593 ( N751, new_n794_, N109 );
not g594 ( new_n796_, keyIn_0_124 );
not g595 ( new_n797_, keyIn_0_85 );
xor g596 ( new_n798_, new_n318_, keyIn_0_71 );
nand g597 ( new_n799_, new_n304_, new_n798_ );
nor g598 ( new_n800_, new_n373_, new_n799_ );
nand g599 ( new_n801_, new_n667_, new_n800_ );
xnor g600 ( new_n802_, new_n801_, new_n797_ );
nor g601 ( new_n803_, new_n802_, new_n570_ );
nand g602 ( new_n804_, new_n803_, keyIn_0_105 );
not g603 ( new_n805_, keyIn_0_105 );
xnor g604 ( new_n806_, new_n801_, keyIn_0_85 );
nand g605 ( new_n807_, new_n806_, new_n477_ );
nand g606 ( new_n808_, new_n807_, new_n805_ );
nand g607 ( new_n809_, new_n804_, new_n808_ );
nand g608 ( new_n810_, new_n809_, N113 );
not g609 ( new_n811_, N113 );
xnor g610 ( new_n812_, new_n807_, keyIn_0_105 );
nand g611 ( new_n813_, new_n812_, new_n811_ );
nand g612 ( new_n814_, new_n813_, new_n810_ );
nand g613 ( new_n815_, new_n814_, new_n796_ );
xnor g614 ( new_n816_, new_n809_, new_n811_ );
nand g615 ( new_n817_, new_n816_, keyIn_0_124 );
nand g616 ( N752, new_n817_, new_n815_ );
not g617 ( new_n819_, keyIn_0_125 );
nor g618 ( new_n820_, new_n802_, new_n451_ );
nand g619 ( new_n821_, new_n820_, keyIn_0_106 );
not g620 ( new_n822_, keyIn_0_106 );
nand g621 ( new_n823_, new_n806_, new_n632_ );
nand g622 ( new_n824_, new_n823_, new_n822_ );
nand g623 ( new_n825_, new_n821_, new_n824_ );
nand g624 ( new_n826_, new_n825_, N117 );
not g625 ( new_n827_, N117 );
xnor g626 ( new_n828_, new_n823_, keyIn_0_106 );
nand g627 ( new_n829_, new_n828_, new_n827_ );
nand g628 ( new_n830_, new_n829_, new_n826_ );
nand g629 ( new_n831_, new_n830_, new_n819_ );
xnor g630 ( new_n832_, new_n825_, new_n827_ );
nand g631 ( new_n833_, new_n832_, keyIn_0_125 );
nand g632 ( N753, new_n833_, new_n831_ );
nand g633 ( new_n835_, new_n806_, new_n504_ );
xnor g634 ( new_n836_, new_n835_, N121 );
xor g635 ( N754, new_n836_, keyIn_0_126 );
nand g636 ( new_n838_, new_n806_, new_n573_ );
xnor g637 ( new_n839_, new_n838_, N125 );
xor g638 ( N755, new_n839_, keyIn_0_127 );
endmodule