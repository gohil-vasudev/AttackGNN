module locked_c2670 (  G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,  G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397, G329, G231, G308, G225  );
  input  G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire new_n359_, new_n360_, new_n361_, new_n362_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n384_, new_n386_, new_n387_, new_n388_, new_n389_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n408_, new_n409_, new_n410_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n527_, new_n528_, new_n530_, new_n532_, new_n533_, new_n534_, new_n535_, new_n537_, new_n538_, new_n539_, new_n540_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n558_, new_n559_, new_n560_, new_n561_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n592_, new_n593_, new_n594_, new_n595_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_;
  INV_X1 g000 ( .A(G44), .ZN(new_n359_) );
  NOR2_X1 g001 ( .A1(new_n359_), .A2(KEYINPUT3), .ZN(new_n360_) );
  NAND2_X1 g002 ( .A1(new_n359_), .A2(KEYINPUT3), .ZN(new_n361_) );
  INV_X1 g003 ( .A(new_n361_), .ZN(new_n362_) );
  NOR2_X1 g004 ( .A1(new_n362_), .A2(new_n360_), .ZN(G218) );
  INV_X1 g005 ( .A(G132), .ZN(G219) );
  INV_X1 g006 ( .A(G82), .ZN(G220) );
  INV_X1 g007 ( .A(G96), .ZN(G221) );
  INV_X1 g008 ( .A(G69), .ZN(G235) );
  INV_X1 g009 ( .A(G120), .ZN(G236) );
  INV_X1 g010 ( .A(G57), .ZN(G237) );
  INV_X1 g011 ( .A(G108), .ZN(G238) );
  INV_X1 g012 ( .A(KEYINPUT20), .ZN(new_n371_) );
  NAND2_X1 g013 ( .A1(G2078), .A2(G2084), .ZN(new_n372_) );
  NAND2_X1 g014 ( .A1(new_n372_), .A2(new_n371_), .ZN(new_n373_) );
  INV_X1 g015 ( .A(new_n372_), .ZN(new_n374_) );
  NAND2_X1 g016 ( .A1(new_n374_), .A2(KEYINPUT20), .ZN(new_n375_) );
  NAND2_X1 g017 ( .A1(new_n375_), .A2(new_n373_), .ZN(new_n376_) );
  NAND2_X1 g018 ( .A1(new_n376_), .A2(G2090), .ZN(new_n377_) );
  NAND2_X1 g019 ( .A1(new_n377_), .A2(KEYINPUT21), .ZN(new_n378_) );
  INV_X1 g020 ( .A(KEYINPUT21), .ZN(new_n379_) );
  NAND3_X1 g021 ( .A1(new_n376_), .A2(G2090), .A3(new_n379_), .ZN(new_n380_) );
  NAND2_X1 g022 ( .A1(new_n378_), .A2(new_n380_), .ZN(new_n381_) );
  NAND2_X1 g023 ( .A1(new_n381_), .A2(G2072), .ZN(G158) );
  NAND3_X1 g024 ( .A1(G2), .A2(G15), .A3(G661), .ZN(G259) );
  NAND2_X1 g025 ( .A1(G94), .A2(G452), .ZN(new_n384_) );
  INV_X1 g026 ( .A(new_n384_), .ZN(G173) );
  NAND2_X1 g027 ( .A1(G7), .A2(G661), .ZN(new_n386_) );
  NAND2_X1 g028 ( .A1(new_n386_), .A2(KEYINPUT10), .ZN(new_n387_) );
  INV_X1 g029 ( .A(KEYINPUT10), .ZN(new_n388_) );
  NAND3_X1 g030 ( .A1(new_n388_), .A2(G7), .A3(G661), .ZN(new_n389_) );
  NAND2_X1 g031 ( .A1(new_n387_), .A2(new_n389_), .ZN(G223) );
  INV_X1 g032 ( .A(KEYINPUT11), .ZN(new_n391_) );
  INV_X1 g033 ( .A(G223), .ZN(new_n392_) );
  NAND2_X1 g034 ( .A1(new_n392_), .A2(G567), .ZN(new_n393_) );
  NAND2_X1 g035 ( .A1(new_n393_), .A2(new_n391_), .ZN(new_n394_) );
  NAND3_X1 g036 ( .A1(new_n392_), .A2(G567), .A3(KEYINPUT11), .ZN(new_n395_) );
  NAND2_X1 g037 ( .A1(new_n394_), .A2(new_n395_), .ZN(G234) );
  NAND2_X1 g038 ( .A1(new_n392_), .A2(G2106), .ZN(G217) );
  INV_X1 g039 ( .A(G218), .ZN(new_n398_) );
  NAND2_X1 g040 ( .A1(G82), .A2(G132), .ZN(new_n399_) );
  NAND2_X1 g041 ( .A1(new_n399_), .A2(KEYINPUT22), .ZN(new_n400_) );
  INV_X1 g042 ( .A(KEYINPUT22), .ZN(new_n401_) );
  NAND3_X1 g043 ( .A1(new_n401_), .A2(G82), .A3(G132), .ZN(new_n402_) );
  NAND4_X1 g044 ( .A1(new_n398_), .A2(G96), .A3(new_n400_), .A4(new_n402_), .ZN(new_n403_) );
  NOR4_X1 g045 ( .A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n404_) );
  INV_X1 g046 ( .A(new_n404_), .ZN(new_n405_) );
  NOR2_X1 g047 ( .A1(new_n403_), .A2(new_n405_), .ZN(G325) );
  INV_X1 g048 ( .A(G325), .ZN(G261) );
  NAND2_X1 g049 ( .A1(new_n403_), .A2(G2106), .ZN(new_n408_) );
  NAND2_X1 g050 ( .A1(new_n405_), .A2(G567), .ZN(new_n409_) );
  NAND2_X1 g051 ( .A1(new_n408_), .A2(new_n409_), .ZN(new_n410_) );
  INV_X1 g052 ( .A(new_n410_), .ZN(G319) );
  INV_X1 g053 ( .A(G2104), .ZN(new_n412_) );
  INV_X1 g054 ( .A(G2105), .ZN(new_n413_) );
  NAND3_X1 g055 ( .A1(new_n412_), .A2(new_n413_), .A3(KEYINPUT17), .ZN(new_n414_) );
  INV_X1 g056 ( .A(KEYINPUT17), .ZN(new_n415_) );
  NAND2_X1 g057 ( .A1(new_n412_), .A2(new_n413_), .ZN(new_n416_) );
  NAND2_X1 g058 ( .A1(new_n416_), .A2(new_n415_), .ZN(new_n417_) );
  NAND3_X1 g059 ( .A1(new_n417_), .A2(G137), .A3(new_n414_), .ZN(new_n418_) );
  NAND3_X1 g060 ( .A1(new_n413_), .A2(G101), .A3(G2104), .ZN(new_n419_) );
  NAND2_X1 g061 ( .A1(new_n419_), .A2(KEYINPUT23), .ZN(new_n420_) );
  NOR2_X1 g062 ( .A1(new_n419_), .A2(KEYINPUT23), .ZN(new_n421_) );
  NAND3_X1 g063 ( .A1(new_n412_), .A2(G125), .A3(G2105), .ZN(new_n422_) );
  NAND3_X1 g064 ( .A1(G113), .A2(G2104), .A3(G2105), .ZN(new_n423_) );
  NAND2_X1 g065 ( .A1(new_n422_), .A2(new_n423_), .ZN(new_n424_) );
  NOR2_X1 g066 ( .A1(new_n421_), .A2(new_n424_), .ZN(new_n425_) );
  NAND3_X1 g067 ( .A1(new_n425_), .A2(new_n418_), .A3(new_n420_), .ZN(new_n426_) );
  INV_X1 g068 ( .A(new_n426_), .ZN(G160) );
  NAND2_X1 g069 ( .A1(new_n417_), .A2(new_n414_), .ZN(new_n428_) );
  INV_X1 g070 ( .A(new_n428_), .ZN(new_n429_) );
  NAND2_X1 g071 ( .A1(new_n429_), .A2(G136), .ZN(new_n430_) );
  NOR2_X1 g072 ( .A1(new_n413_), .A2(G2104), .ZN(new_n431_) );
  NAND2_X1 g073 ( .A1(new_n431_), .A2(G124), .ZN(new_n432_) );
  NAND2_X1 g074 ( .A1(new_n432_), .A2(KEYINPUT44), .ZN(new_n433_) );
  INV_X1 g075 ( .A(KEYINPUT44), .ZN(new_n434_) );
  NAND3_X1 g076 ( .A1(new_n431_), .A2(G124), .A3(new_n434_), .ZN(new_n435_) );
  NAND2_X1 g077 ( .A1(new_n433_), .A2(new_n435_), .ZN(new_n436_) );
  NOR2_X1 g078 ( .A1(new_n412_), .A2(G2105), .ZN(new_n437_) );
  NAND2_X1 g079 ( .A1(new_n437_), .A2(G100), .ZN(new_n438_) );
  NAND2_X1 g080 ( .A1(G2104), .A2(G2105), .ZN(new_n439_) );
  INV_X1 g081 ( .A(new_n439_), .ZN(new_n440_) );
  NAND2_X1 g082 ( .A1(new_n440_), .A2(G112), .ZN(new_n441_) );
  NAND2_X1 g083 ( .A1(new_n438_), .A2(new_n441_), .ZN(new_n442_) );
  INV_X1 g084 ( .A(new_n442_), .ZN(new_n443_) );
  NAND3_X1 g085 ( .A1(new_n430_), .A2(new_n436_), .A3(new_n443_), .ZN(new_n444_) );
  INV_X1 g086 ( .A(new_n444_), .ZN(G162) );
  NAND3_X1 g087 ( .A1(new_n417_), .A2(G138), .A3(new_n414_), .ZN(new_n446_) );
  NAND3_X1 g088 ( .A1(G114), .A2(G2104), .A3(G2105), .ZN(new_n447_) );
  NAND3_X1 g089 ( .A1(new_n413_), .A2(G102), .A3(G2104), .ZN(new_n448_) );
  NAND3_X1 g090 ( .A1(new_n412_), .A2(G126), .A3(G2105), .ZN(new_n449_) );
  NAND3_X1 g091 ( .A1(new_n448_), .A2(new_n449_), .A3(new_n447_), .ZN(new_n450_) );
  INV_X1 g092 ( .A(new_n450_), .ZN(new_n451_) );
  NAND2_X1 g093 ( .A1(new_n451_), .A2(new_n446_), .ZN(new_n452_) );
  INV_X1 g094 ( .A(new_n452_), .ZN(G164) );
  INV_X1 g095 ( .A(G651), .ZN(new_n454_) );
  INV_X1 g096 ( .A(KEYINPUT0), .ZN(new_n455_) );
  NAND2_X1 g097 ( .A1(new_n455_), .A2(G543), .ZN(new_n456_) );
  INV_X1 g098 ( .A(G543), .ZN(new_n457_) );
  NAND2_X1 g099 ( .A1(new_n457_), .A2(KEYINPUT0), .ZN(new_n458_) );
  NAND3_X1 g100 ( .A1(new_n456_), .A2(new_n458_), .A3(new_n454_), .ZN(new_n459_) );
  INV_X1 g101 ( .A(new_n459_), .ZN(new_n460_) );
  NAND2_X1 g102 ( .A1(new_n460_), .A2(G50), .ZN(new_n461_) );
  NOR2_X1 g103 ( .A1(G543), .A2(G651), .ZN(new_n462_) );
  NAND2_X1 g104 ( .A1(new_n462_), .A2(G88), .ZN(new_n463_) );
  NAND3_X1 g105 ( .A1(new_n456_), .A2(new_n458_), .A3(G651), .ZN(new_n464_) );
  INV_X1 g106 ( .A(new_n464_), .ZN(new_n465_) );
  NAND2_X1 g107 ( .A1(new_n465_), .A2(G75), .ZN(new_n466_) );
  NAND2_X1 g108 ( .A1(new_n457_), .A2(G651), .ZN(new_n467_) );
  NAND2_X1 g109 ( .A1(new_n467_), .A2(KEYINPUT1), .ZN(new_n468_) );
  INV_X1 g110 ( .A(KEYINPUT1), .ZN(new_n469_) );
  NAND3_X1 g111 ( .A1(new_n457_), .A2(new_n469_), .A3(G651), .ZN(new_n470_) );
  NAND2_X1 g112 ( .A1(new_n468_), .A2(new_n470_), .ZN(new_n471_) );
  NAND2_X1 g113 ( .A1(new_n471_), .A2(G62), .ZN(new_n472_) );
  NAND4_X1 g114 ( .A1(new_n461_), .A2(new_n466_), .A3(new_n463_), .A4(new_n472_), .ZN(G303) );
  INV_X1 g115 ( .A(G303), .ZN(G166) );
  INV_X1 g116 ( .A(KEYINPUT6), .ZN(new_n475_) );
  NAND2_X1 g117 ( .A1(new_n460_), .A2(G51), .ZN(new_n476_) );
  NAND2_X1 g118 ( .A1(new_n471_), .A2(G63), .ZN(new_n477_) );
  NAND2_X1 g119 ( .A1(new_n476_), .A2(new_n477_), .ZN(new_n478_) );
  NAND2_X1 g120 ( .A1(new_n478_), .A2(new_n475_), .ZN(new_n479_) );
  NAND3_X1 g121 ( .A1(new_n476_), .A2(new_n477_), .A3(KEYINPUT6), .ZN(new_n480_) );
  NAND2_X1 g122 ( .A1(new_n479_), .A2(new_n480_), .ZN(new_n481_) );
  NAND2_X1 g123 ( .A1(new_n465_), .A2(G76), .ZN(new_n482_) );
  NAND2_X1 g124 ( .A1(new_n462_), .A2(G89), .ZN(new_n483_) );
  NAND2_X1 g125 ( .A1(new_n483_), .A2(KEYINPUT4), .ZN(new_n484_) );
  INV_X1 g126 ( .A(KEYINPUT4), .ZN(new_n485_) );
  NAND3_X1 g127 ( .A1(new_n462_), .A2(G89), .A3(new_n485_), .ZN(new_n486_) );
  NAND2_X1 g128 ( .A1(new_n484_), .A2(new_n486_), .ZN(new_n487_) );
  NAND2_X1 g129 ( .A1(new_n482_), .A2(new_n487_), .ZN(new_n488_) );
  NAND2_X1 g130 ( .A1(new_n488_), .A2(KEYINPUT5), .ZN(new_n489_) );
  INV_X1 g131 ( .A(KEYINPUT5), .ZN(new_n490_) );
  NAND3_X1 g132 ( .A1(new_n482_), .A2(new_n490_), .A3(new_n487_), .ZN(new_n491_) );
  NAND2_X1 g133 ( .A1(new_n489_), .A2(new_n491_), .ZN(new_n492_) );
  NAND2_X1 g134 ( .A1(new_n481_), .A2(new_n492_), .ZN(new_n493_) );
  NAND2_X1 g135 ( .A1(new_n493_), .A2(KEYINPUT7), .ZN(new_n494_) );
  INV_X1 g136 ( .A(KEYINPUT7), .ZN(new_n495_) );
  NAND3_X1 g137 ( .A1(new_n481_), .A2(new_n492_), .A3(new_n495_), .ZN(new_n496_) );
  NAND2_X1 g138 ( .A1(new_n494_), .A2(new_n496_), .ZN(G168) );
  NAND2_X1 g139 ( .A1(new_n465_), .A2(G77), .ZN(new_n498_) );
  NAND2_X1 g140 ( .A1(new_n462_), .A2(G90), .ZN(new_n499_) );
  NAND3_X1 g141 ( .A1(new_n498_), .A2(KEYINPUT9), .A3(new_n499_), .ZN(new_n500_) );
  INV_X1 g142 ( .A(KEYINPUT9), .ZN(new_n501_) );
  NAND2_X1 g143 ( .A1(new_n498_), .A2(new_n499_), .ZN(new_n502_) );
  NAND2_X1 g144 ( .A1(new_n502_), .A2(new_n501_), .ZN(new_n503_) );
  NAND2_X1 g145 ( .A1(new_n460_), .A2(G52), .ZN(new_n504_) );
  NAND2_X1 g146 ( .A1(new_n471_), .A2(G64), .ZN(new_n505_) );
  NAND4_X1 g147 ( .A1(new_n503_), .A2(new_n500_), .A3(new_n504_), .A4(new_n505_), .ZN(G301) );
  INV_X1 g148 ( .A(G301), .ZN(G171) );
  NAND4_X1 g149 ( .A1(new_n456_), .A2(new_n458_), .A3(G68), .A4(G651), .ZN(new_n508_) );
  NAND3_X1 g150 ( .A1(new_n457_), .A2(new_n454_), .A3(G81), .ZN(new_n509_) );
  NAND2_X1 g151 ( .A1(new_n509_), .A2(KEYINPUT12), .ZN(new_n510_) );
  INV_X1 g152 ( .A(KEYINPUT12), .ZN(new_n511_) );
  NAND3_X1 g153 ( .A1(new_n462_), .A2(G81), .A3(new_n511_), .ZN(new_n512_) );
  NAND2_X1 g154 ( .A1(new_n510_), .A2(new_n512_), .ZN(new_n513_) );
  NAND2_X1 g155 ( .A1(new_n513_), .A2(new_n508_), .ZN(new_n514_) );
  NAND2_X1 g156 ( .A1(new_n514_), .A2(KEYINPUT13), .ZN(new_n515_) );
  INV_X1 g157 ( .A(KEYINPUT13), .ZN(new_n516_) );
  NAND3_X1 g158 ( .A1(new_n513_), .A2(new_n516_), .A3(new_n508_), .ZN(new_n517_) );
  NAND2_X1 g159 ( .A1(new_n515_), .A2(new_n517_), .ZN(new_n518_) );
  NAND3_X1 g160 ( .A1(new_n471_), .A2(G56), .A3(KEYINPUT14), .ZN(new_n519_) );
  INV_X1 g161 ( .A(KEYINPUT14), .ZN(new_n520_) );
  NAND2_X1 g162 ( .A1(new_n471_), .A2(G56), .ZN(new_n521_) );
  NAND2_X1 g163 ( .A1(new_n521_), .A2(new_n520_), .ZN(new_n522_) );
  NAND2_X1 g164 ( .A1(new_n460_), .A2(G43), .ZN(new_n523_) );
  NAND4_X1 g165 ( .A1(new_n518_), .A2(new_n519_), .A3(new_n522_), .A4(new_n523_), .ZN(new_n524_) );
  INV_X1 g166 ( .A(new_n524_), .ZN(new_n525_) );
  NAND2_X1 g167 ( .A1(new_n525_), .A2(G860), .ZN(G153) );
  NAND3_X1 g168 ( .A1(G319), .A2(G483), .A3(G661), .ZN(new_n527_) );
  INV_X1 g169 ( .A(new_n527_), .ZN(new_n528_) );
  NAND2_X1 g170 ( .A1(new_n528_), .A2(G36), .ZN(G176) );
  NAND2_X1 g171 ( .A1(G1), .A2(G3), .ZN(new_n530_) );
  NAND2_X1 g172 ( .A1(new_n528_), .A2(new_n530_), .ZN(G188) );
  NAND2_X1 g173 ( .A1(new_n465_), .A2(G78), .ZN(new_n532_) );
  NAND2_X1 g174 ( .A1(new_n462_), .A2(G91), .ZN(new_n533_) );
  NAND2_X1 g175 ( .A1(new_n460_), .A2(G53), .ZN(new_n534_) );
  NAND2_X1 g176 ( .A1(new_n471_), .A2(G65), .ZN(new_n535_) );
  NAND4_X1 g177 ( .A1(new_n532_), .A2(new_n534_), .A3(new_n533_), .A4(new_n535_), .ZN(G299) );
  INV_X1 g178 ( .A(KEYINPUT8), .ZN(new_n537_) );
  NAND2_X1 g179 ( .A1(G168), .A2(new_n537_), .ZN(new_n538_) );
  INV_X1 g180 ( .A(G168), .ZN(new_n539_) );
  NAND2_X1 g181 ( .A1(new_n539_), .A2(KEYINPUT8), .ZN(new_n540_) );
  NAND2_X1 g182 ( .A1(new_n540_), .A2(new_n538_), .ZN(G286) );
  INV_X1 g183 ( .A(new_n471_), .ZN(new_n542_) );
  NAND2_X1 g184 ( .A1(new_n460_), .A2(G49), .ZN(new_n543_) );
  NAND2_X1 g185 ( .A1(new_n456_), .A2(new_n458_), .ZN(new_n544_) );
  NAND2_X1 g186 ( .A1(new_n544_), .A2(G87), .ZN(new_n545_) );
  NAND2_X1 g187 ( .A1(G74), .A2(G651), .ZN(new_n546_) );
  NAND4_X1 g188 ( .A1(new_n543_), .A2(new_n542_), .A3(new_n545_), .A4(new_n546_), .ZN(G288) );
  NAND2_X1 g189 ( .A1(new_n465_), .A2(G73), .ZN(new_n548_) );
  NAND2_X1 g190 ( .A1(new_n548_), .A2(KEYINPUT2), .ZN(new_n549_) );
  INV_X1 g191 ( .A(new_n549_), .ZN(new_n550_) );
  NOR2_X1 g192 ( .A1(new_n548_), .A2(KEYINPUT2), .ZN(new_n551_) );
  NOR2_X1 g193 ( .A1(new_n550_), .A2(new_n551_), .ZN(new_n552_) );
  INV_X1 g194 ( .A(new_n552_), .ZN(new_n553_) );
  NAND2_X1 g195 ( .A1(new_n471_), .A2(G61), .ZN(new_n554_) );
  NAND2_X1 g196 ( .A1(new_n460_), .A2(G48), .ZN(new_n555_) );
  NAND2_X1 g197 ( .A1(new_n462_), .A2(G86), .ZN(new_n556_) );
  NAND4_X1 g198 ( .A1(new_n553_), .A2(new_n554_), .A3(new_n555_), .A4(new_n556_), .ZN(G305) );
  NAND2_X1 g199 ( .A1(new_n465_), .A2(G72), .ZN(new_n558_) );
  NAND2_X1 g200 ( .A1(new_n462_), .A2(G85), .ZN(new_n559_) );
  NAND2_X1 g201 ( .A1(new_n460_), .A2(G47), .ZN(new_n560_) );
  NAND2_X1 g202 ( .A1(new_n471_), .A2(G60), .ZN(new_n561_) );
  NAND4_X1 g203 ( .A1(new_n558_), .A2(new_n560_), .A3(new_n559_), .A4(new_n561_), .ZN(G290) );
  NAND2_X1 g204 ( .A1(G301), .A2(G868), .ZN(new_n563_) );
  INV_X1 g205 ( .A(G868), .ZN(new_n564_) );
  INV_X1 g206 ( .A(KEYINPUT15), .ZN(new_n565_) );
  NAND2_X1 g207 ( .A1(new_n460_), .A2(G54), .ZN(new_n566_) );
  NAND2_X1 g208 ( .A1(new_n462_), .A2(G92), .ZN(new_n567_) );
  NAND2_X1 g209 ( .A1(new_n566_), .A2(new_n567_), .ZN(new_n568_) );
  INV_X1 g210 ( .A(new_n568_), .ZN(new_n569_) );
  NAND2_X1 g211 ( .A1(new_n465_), .A2(G79), .ZN(new_n570_) );
  NAND2_X1 g212 ( .A1(new_n471_), .A2(G66), .ZN(new_n571_) );
  NAND4_X1 g213 ( .A1(new_n569_), .A2(new_n565_), .A3(new_n570_), .A4(new_n571_), .ZN(new_n572_) );
  NAND4_X1 g214 ( .A1(new_n566_), .A2(new_n570_), .A3(new_n567_), .A4(new_n571_), .ZN(new_n573_) );
  NAND2_X1 g215 ( .A1(new_n573_), .A2(KEYINPUT15), .ZN(new_n574_) );
  NAND2_X1 g216 ( .A1(new_n572_), .A2(new_n574_), .ZN(new_n575_) );
  INV_X1 g217 ( .A(new_n575_), .ZN(new_n576_) );
  NAND2_X1 g218 ( .A1(new_n576_), .A2(new_n564_), .ZN(new_n577_) );
  NAND2_X1 g219 ( .A1(new_n577_), .A2(new_n563_), .ZN(G284) );
  INV_X1 g220 ( .A(G286), .ZN(new_n579_) );
  NAND2_X1 g221 ( .A1(new_n579_), .A2(G868), .ZN(new_n580_) );
  INV_X1 g222 ( .A(G299), .ZN(new_n581_) );
  NAND2_X1 g223 ( .A1(new_n581_), .A2(new_n564_), .ZN(new_n582_) );
  NAND2_X1 g224 ( .A1(new_n580_), .A2(new_n582_), .ZN(new_n583_) );
  INV_X1 g225 ( .A(new_n583_), .ZN(G297) );
  INV_X1 g226 ( .A(KEYINPUT16), .ZN(new_n585_) );
  INV_X1 g227 ( .A(G860), .ZN(new_n586_) );
  NAND2_X1 g228 ( .A1(new_n586_), .A2(G559), .ZN(new_n587_) );
  NAND3_X1 g229 ( .A1(new_n575_), .A2(new_n585_), .A3(new_n587_), .ZN(new_n588_) );
  NAND2_X1 g230 ( .A1(new_n575_), .A2(new_n587_), .ZN(new_n589_) );
  NAND2_X1 g231 ( .A1(new_n589_), .A2(KEYINPUT16), .ZN(new_n590_) );
  NAND2_X1 g232 ( .A1(new_n590_), .A2(new_n588_), .ZN(G148) );
  INV_X1 g233 ( .A(G559), .ZN(new_n592_) );
  NAND3_X1 g234 ( .A1(new_n575_), .A2(new_n592_), .A3(G868), .ZN(new_n593_) );
  NAND2_X1 g235 ( .A1(new_n525_), .A2(new_n564_), .ZN(new_n594_) );
  NAND2_X1 g236 ( .A1(new_n593_), .A2(new_n594_), .ZN(new_n595_) );
  INV_X1 g237 ( .A(new_n595_), .ZN(G282) );
  INV_X1 g238 ( .A(G2100), .ZN(new_n597_) );
  NAND2_X1 g239 ( .A1(new_n429_), .A2(G135), .ZN(new_n598_) );
  NAND3_X1 g240 ( .A1(new_n431_), .A2(G123), .A3(KEYINPUT18), .ZN(new_n599_) );
  INV_X1 g241 ( .A(KEYINPUT18), .ZN(new_n600_) );
  NAND2_X1 g242 ( .A1(new_n431_), .A2(G123), .ZN(new_n601_) );
  NAND2_X1 g243 ( .A1(new_n601_), .A2(new_n600_), .ZN(new_n602_) );
  NAND2_X1 g244 ( .A1(new_n437_), .A2(G99), .ZN(new_n603_) );
  NAND2_X1 g245 ( .A1(new_n440_), .A2(G111), .ZN(new_n604_) );
  NAND2_X1 g246 ( .A1(new_n603_), .A2(new_n604_), .ZN(new_n605_) );
  INV_X1 g247 ( .A(new_n605_), .ZN(new_n606_) );
  NAND4_X1 g248 ( .A1(new_n598_), .A2(new_n606_), .A3(new_n599_), .A4(new_n602_), .ZN(new_n607_) );
  NAND2_X1 g249 ( .A1(new_n607_), .A2(G2096), .ZN(new_n608_) );
  INV_X1 g250 ( .A(G2096), .ZN(new_n609_) );
  INV_X1 g251 ( .A(new_n607_), .ZN(new_n610_) );
  NAND2_X1 g252 ( .A1(new_n610_), .A2(new_n609_), .ZN(new_n611_) );
  NAND3_X1 g253 ( .A1(new_n611_), .A2(new_n597_), .A3(new_n608_), .ZN(G156) );
  INV_X1 g254 ( .A(G2454), .ZN(new_n613_) );
  NAND2_X1 g255 ( .A1(new_n613_), .A2(G2430), .ZN(new_n614_) );
  INV_X1 g256 ( .A(G2430), .ZN(new_n615_) );
  NAND2_X1 g257 ( .A1(new_n615_), .A2(G2454), .ZN(new_n616_) );
  NAND2_X1 g258 ( .A1(new_n614_), .A2(new_n616_), .ZN(new_n617_) );
  NAND2_X1 g259 ( .A1(G1341), .A2(G1348), .ZN(new_n618_) );
  INV_X1 g260 ( .A(G1341), .ZN(new_n619_) );
  INV_X1 g261 ( .A(G1348), .ZN(new_n620_) );
  NAND2_X1 g262 ( .A1(new_n619_), .A2(new_n620_), .ZN(new_n621_) );
  NAND2_X1 g263 ( .A1(new_n621_), .A2(new_n618_), .ZN(new_n622_) );
  NAND2_X1 g264 ( .A1(new_n617_), .A2(new_n622_), .ZN(new_n623_) );
  NAND4_X1 g265 ( .A1(new_n621_), .A2(new_n614_), .A3(new_n616_), .A4(new_n618_), .ZN(new_n624_) );
  NAND2_X1 g266 ( .A1(new_n623_), .A2(new_n624_), .ZN(new_n625_) );
  NAND2_X1 g267 ( .A1(G2435), .A2(G2438), .ZN(new_n626_) );
  INV_X1 g268 ( .A(new_n626_), .ZN(new_n627_) );
  NOR2_X1 g269 ( .A1(G2435), .A2(G2438), .ZN(new_n628_) );
  NOR2_X1 g270 ( .A1(new_n627_), .A2(new_n628_), .ZN(new_n629_) );
  INV_X1 g271 ( .A(new_n629_), .ZN(new_n630_) );
  NAND2_X1 g272 ( .A1(new_n625_), .A2(new_n630_), .ZN(new_n631_) );
  NAND3_X1 g273 ( .A1(new_n623_), .A2(new_n624_), .A3(new_n629_), .ZN(new_n632_) );
  NAND2_X1 g274 ( .A1(G2446), .A2(G2451), .ZN(new_n633_) );
  INV_X1 g275 ( .A(G2446), .ZN(new_n634_) );
  INV_X1 g276 ( .A(G2451), .ZN(new_n635_) );
  NAND2_X1 g277 ( .A1(new_n634_), .A2(new_n635_), .ZN(new_n636_) );
  NAND2_X1 g278 ( .A1(new_n636_), .A2(new_n633_), .ZN(new_n637_) );
  NAND2_X1 g279 ( .A1(G2427), .A2(G2443), .ZN(new_n638_) );
  INV_X1 g280 ( .A(G2427), .ZN(new_n639_) );
  INV_X1 g281 ( .A(G2443), .ZN(new_n640_) );
  NAND2_X1 g282 ( .A1(new_n639_), .A2(new_n640_), .ZN(new_n641_) );
  NAND2_X1 g283 ( .A1(new_n641_), .A2(new_n638_), .ZN(new_n642_) );
  NAND2_X1 g284 ( .A1(new_n637_), .A2(new_n642_), .ZN(new_n643_) );
  NAND4_X1 g285 ( .A1(new_n636_), .A2(new_n641_), .A3(new_n633_), .A4(new_n638_), .ZN(new_n644_) );
  NAND4_X1 g286 ( .A1(new_n631_), .A2(new_n632_), .A3(new_n643_), .A4(new_n644_), .ZN(new_n645_) );
  NAND2_X1 g287 ( .A1(new_n631_), .A2(new_n632_), .ZN(new_n646_) );
  NAND2_X1 g288 ( .A1(new_n643_), .A2(new_n644_), .ZN(new_n647_) );
  NAND2_X1 g289 ( .A1(new_n646_), .A2(new_n647_), .ZN(new_n648_) );
  NAND3_X1 g290 ( .A1(new_n648_), .A2(G14), .A3(new_n645_), .ZN(new_n649_) );
  INV_X1 g291 ( .A(new_n649_), .ZN(G401) );
  INV_X1 g292 ( .A(KEYINPUT42), .ZN(new_n651_) );
  NAND2_X1 g293 ( .A1(new_n651_), .A2(G2090), .ZN(new_n652_) );
  INV_X1 g294 ( .A(G2090), .ZN(new_n653_) );
  NAND2_X1 g295 ( .A1(new_n653_), .A2(KEYINPUT42), .ZN(new_n654_) );
  NAND2_X1 g296 ( .A1(new_n652_), .A2(new_n654_), .ZN(new_n655_) );
  NAND2_X1 g297 ( .A1(G2067), .A2(G2072), .ZN(new_n656_) );
  INV_X1 g298 ( .A(G2067), .ZN(new_n657_) );
  INV_X1 g299 ( .A(G2072), .ZN(new_n658_) );
  NAND2_X1 g300 ( .A1(new_n657_), .A2(new_n658_), .ZN(new_n659_) );
  NAND2_X1 g301 ( .A1(new_n659_), .A2(new_n656_), .ZN(new_n660_) );
  NAND2_X1 g302 ( .A1(new_n655_), .A2(new_n660_), .ZN(new_n661_) );
  NAND4_X1 g303 ( .A1(new_n659_), .A2(new_n652_), .A3(new_n654_), .A4(new_n656_), .ZN(new_n662_) );
  NAND2_X1 g304 ( .A1(new_n661_), .A2(new_n662_), .ZN(new_n663_) );
  NAND2_X1 g305 ( .A1(G2096), .A2(G2100), .ZN(new_n664_) );
  NAND2_X1 g306 ( .A1(new_n609_), .A2(new_n597_), .ZN(new_n665_) );
  NAND2_X1 g307 ( .A1(new_n665_), .A2(new_n664_), .ZN(new_n666_) );
  NAND2_X1 g308 ( .A1(G2678), .A2(KEYINPUT43), .ZN(new_n667_) );
  INV_X1 g309 ( .A(G2678), .ZN(new_n668_) );
  INV_X1 g310 ( .A(KEYINPUT43), .ZN(new_n669_) );
  NAND2_X1 g311 ( .A1(new_n668_), .A2(new_n669_), .ZN(new_n670_) );
  NAND2_X1 g312 ( .A1(new_n670_), .A2(new_n667_), .ZN(new_n671_) );
  NAND2_X1 g313 ( .A1(new_n666_), .A2(new_n671_), .ZN(new_n672_) );
  NAND4_X1 g314 ( .A1(new_n665_), .A2(new_n670_), .A3(new_n664_), .A4(new_n667_), .ZN(new_n673_) );
  NAND2_X1 g315 ( .A1(new_n672_), .A2(new_n673_), .ZN(new_n674_) );
  NAND2_X1 g316 ( .A1(new_n663_), .A2(new_n674_), .ZN(new_n675_) );
  NAND4_X1 g317 ( .A1(new_n661_), .A2(new_n672_), .A3(new_n662_), .A4(new_n673_), .ZN(new_n676_) );
  NAND2_X1 g318 ( .A1(new_n675_), .A2(new_n676_), .ZN(new_n677_) );
  NOR2_X1 g319 ( .A1(G2078), .A2(G2084), .ZN(new_n678_) );
  NOR2_X1 g320 ( .A1(new_n374_), .A2(new_n678_), .ZN(new_n679_) );
  INV_X1 g321 ( .A(new_n679_), .ZN(new_n680_) );
  NAND2_X1 g322 ( .A1(new_n677_), .A2(new_n680_), .ZN(new_n681_) );
  NAND3_X1 g323 ( .A1(new_n675_), .A2(new_n676_), .A3(new_n679_), .ZN(new_n682_) );
  NAND2_X1 g324 ( .A1(new_n681_), .A2(new_n682_), .ZN(G227) );
  INV_X1 g325 ( .A(G1981), .ZN(new_n684_) );
  NAND2_X1 g326 ( .A1(new_n684_), .A2(G1976), .ZN(new_n685_) );
  INV_X1 g327 ( .A(G1976), .ZN(new_n686_) );
  NAND2_X1 g328 ( .A1(new_n686_), .A2(G1981), .ZN(new_n687_) );
  NAND2_X1 g329 ( .A1(new_n685_), .A2(new_n687_), .ZN(new_n688_) );
  NAND2_X1 g330 ( .A1(G1956), .A2(G1966), .ZN(new_n689_) );
  INV_X1 g331 ( .A(G1956), .ZN(new_n690_) );
  INV_X1 g332 ( .A(G1966), .ZN(new_n691_) );
  NAND2_X1 g333 ( .A1(new_n690_), .A2(new_n691_), .ZN(new_n692_) );
  NAND2_X1 g334 ( .A1(new_n692_), .A2(new_n689_), .ZN(new_n693_) );
  NAND2_X1 g335 ( .A1(new_n688_), .A2(new_n693_), .ZN(new_n694_) );
  NAND4_X1 g336 ( .A1(new_n692_), .A2(new_n685_), .A3(new_n687_), .A4(new_n689_), .ZN(new_n695_) );
  NAND2_X1 g337 ( .A1(new_n694_), .A2(new_n695_), .ZN(new_n696_) );
  NAND2_X1 g338 ( .A1(new_n696_), .A2(G2474), .ZN(new_n697_) );
  INV_X1 g339 ( .A(G2474), .ZN(new_n698_) );
  NAND3_X1 g340 ( .A1(new_n694_), .A2(new_n698_), .A3(new_n695_), .ZN(new_n699_) );
  NAND2_X1 g341 ( .A1(new_n697_), .A2(new_n699_), .ZN(new_n700_) );
  INV_X1 g342 ( .A(G1991), .ZN(new_n701_) );
  NOR2_X1 g343 ( .A1(new_n701_), .A2(G1996), .ZN(new_n702_) );
  INV_X1 g344 ( .A(G1996), .ZN(new_n703_) );
  NOR2_X1 g345 ( .A1(new_n703_), .A2(G1991), .ZN(new_n704_) );
  NOR2_X1 g346 ( .A1(new_n702_), .A2(new_n704_), .ZN(new_n705_) );
  INV_X1 g347 ( .A(new_n705_), .ZN(new_n706_) );
  NAND2_X1 g348 ( .A1(new_n700_), .A2(new_n706_), .ZN(new_n707_) );
  NAND3_X1 g349 ( .A1(new_n697_), .A2(new_n699_), .A3(new_n705_), .ZN(new_n708_) );
  NAND2_X1 g350 ( .A1(new_n707_), .A2(new_n708_), .ZN(new_n709_) );
  NAND2_X1 g351 ( .A1(G1971), .A2(KEYINPUT41), .ZN(new_n710_) );
  INV_X1 g352 ( .A(G1971), .ZN(new_n711_) );
  INV_X1 g353 ( .A(KEYINPUT41), .ZN(new_n712_) );
  NAND2_X1 g354 ( .A1(new_n711_), .A2(new_n712_), .ZN(new_n713_) );
  NAND2_X1 g355 ( .A1(new_n713_), .A2(new_n710_), .ZN(new_n714_) );
  NAND2_X1 g356 ( .A1(G1961), .A2(G1986), .ZN(new_n715_) );
  INV_X1 g357 ( .A(G1961), .ZN(new_n716_) );
  INV_X1 g358 ( .A(G1986), .ZN(new_n717_) );
  NAND2_X1 g359 ( .A1(new_n716_), .A2(new_n717_), .ZN(new_n718_) );
  NAND2_X1 g360 ( .A1(new_n718_), .A2(new_n715_), .ZN(new_n719_) );
  NAND2_X1 g361 ( .A1(new_n714_), .A2(new_n719_), .ZN(new_n720_) );
  NAND4_X1 g362 ( .A1(new_n713_), .A2(new_n718_), .A3(new_n710_), .A4(new_n715_), .ZN(new_n721_) );
  NAND2_X1 g363 ( .A1(new_n720_), .A2(new_n721_), .ZN(new_n722_) );
  NAND2_X1 g364 ( .A1(new_n709_), .A2(new_n722_), .ZN(new_n723_) );
  NAND4_X1 g365 ( .A1(new_n707_), .A2(new_n708_), .A3(new_n720_), .A4(new_n721_), .ZN(new_n724_) );
  NAND2_X1 g366 ( .A1(new_n723_), .A2(new_n724_), .ZN(new_n725_) );
  INV_X1 g367 ( .A(new_n725_), .ZN(G229) );
  INV_X1 g368 ( .A(KEYINPUT55), .ZN(new_n727_) );
  INV_X1 g369 ( .A(KEYINPUT52), .ZN(new_n728_) );
  INV_X1 g370 ( .A(G139), .ZN(new_n729_) );
  NOR2_X1 g371 ( .A1(new_n428_), .A2(new_n729_), .ZN(new_n730_) );
  NAND2_X1 g372 ( .A1(new_n437_), .A2(G103), .ZN(new_n731_) );
  INV_X1 g373 ( .A(new_n731_), .ZN(new_n732_) );
  NOR2_X1 g374 ( .A1(new_n730_), .A2(new_n732_), .ZN(new_n733_) );
  INV_X1 g375 ( .A(KEYINPUT47), .ZN(new_n734_) );
  NAND2_X1 g376 ( .A1(new_n431_), .A2(G127), .ZN(new_n735_) );
  NAND2_X1 g377 ( .A1(new_n440_), .A2(G115), .ZN(new_n736_) );
  NAND2_X1 g378 ( .A1(new_n735_), .A2(new_n736_), .ZN(new_n737_) );
  NAND2_X1 g379 ( .A1(new_n737_), .A2(new_n734_), .ZN(new_n738_) );
  NAND3_X1 g380 ( .A1(new_n735_), .A2(new_n736_), .A3(KEYINPUT47), .ZN(new_n739_) );
  NAND2_X1 g381 ( .A1(new_n738_), .A2(new_n739_), .ZN(new_n740_) );
  INV_X1 g382 ( .A(new_n740_), .ZN(new_n741_) );
  NAND2_X1 g383 ( .A1(new_n741_), .A2(new_n733_), .ZN(new_n742_) );
  NAND2_X1 g384 ( .A1(new_n742_), .A2(G2072), .ZN(new_n743_) );
  INV_X1 g385 ( .A(G2078), .ZN(new_n744_) );
  NAND2_X1 g386 ( .A1(new_n452_), .A2(new_n744_), .ZN(new_n745_) );
  NAND2_X1 g387 ( .A1(G164), .A2(G2078), .ZN(new_n746_) );
  NAND2_X1 g388 ( .A1(new_n746_), .A2(new_n745_), .ZN(new_n747_) );
  NAND3_X1 g389 ( .A1(new_n741_), .A2(new_n658_), .A3(new_n733_), .ZN(new_n748_) );
  NAND3_X1 g390 ( .A1(new_n743_), .A2(new_n747_), .A3(new_n748_), .ZN(new_n749_) );
  NAND2_X1 g391 ( .A1(new_n749_), .A2(KEYINPUT50), .ZN(new_n750_) );
  INV_X1 g392 ( .A(new_n750_), .ZN(new_n751_) );
  INV_X1 g393 ( .A(KEYINPUT51), .ZN(new_n752_) );
  NAND2_X1 g394 ( .A1(new_n429_), .A2(G141), .ZN(new_n753_) );
  NAND3_X1 g395 ( .A1(new_n437_), .A2(G105), .A3(KEYINPUT38), .ZN(new_n754_) );
  INV_X1 g396 ( .A(KEYINPUT38), .ZN(new_n755_) );
  NAND2_X1 g397 ( .A1(new_n437_), .A2(G105), .ZN(new_n756_) );
  NAND2_X1 g398 ( .A1(new_n756_), .A2(new_n755_), .ZN(new_n757_) );
  NAND2_X1 g399 ( .A1(new_n431_), .A2(G129), .ZN(new_n758_) );
  NAND2_X1 g400 ( .A1(new_n440_), .A2(G117), .ZN(new_n759_) );
  NAND2_X1 g401 ( .A1(new_n758_), .A2(new_n759_), .ZN(new_n760_) );
  INV_X1 g402 ( .A(new_n760_), .ZN(new_n761_) );
  NAND4_X1 g403 ( .A1(new_n753_), .A2(new_n761_), .A3(new_n754_), .A4(new_n757_), .ZN(new_n762_) );
  INV_X1 g404 ( .A(new_n762_), .ZN(new_n763_) );
  NAND2_X1 g405 ( .A1(new_n763_), .A2(new_n703_), .ZN(new_n764_) );
  NAND2_X1 g406 ( .A1(G162), .A2(new_n653_), .ZN(new_n765_) );
  NAND2_X1 g407 ( .A1(new_n444_), .A2(G2090), .ZN(new_n766_) );
  NAND3_X1 g408 ( .A1(new_n764_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n767_) );
  NAND2_X1 g409 ( .A1(new_n767_), .A2(new_n752_), .ZN(new_n768_) );
  INV_X1 g410 ( .A(KEYINPUT50), .ZN(new_n769_) );
  NAND4_X1 g411 ( .A1(new_n743_), .A2(new_n769_), .A3(new_n747_), .A4(new_n748_), .ZN(new_n770_) );
  NAND2_X1 g412 ( .A1(new_n768_), .A2(new_n770_), .ZN(new_n771_) );
  NOR2_X1 g413 ( .A1(new_n751_), .A2(new_n771_), .ZN(new_n772_) );
  INV_X1 g414 ( .A(KEYINPUT34), .ZN(new_n773_) );
  NAND2_X1 g415 ( .A1(new_n429_), .A2(G140), .ZN(new_n774_) );
  NAND2_X1 g416 ( .A1(new_n437_), .A2(G104), .ZN(new_n775_) );
  NAND3_X1 g417 ( .A1(new_n774_), .A2(new_n773_), .A3(new_n775_), .ZN(new_n776_) );
  NAND2_X1 g418 ( .A1(new_n774_), .A2(new_n775_), .ZN(new_n777_) );
  NAND2_X1 g419 ( .A1(new_n777_), .A2(KEYINPUT34), .ZN(new_n778_) );
  NAND2_X1 g420 ( .A1(new_n431_), .A2(G128), .ZN(new_n779_) );
  NAND2_X1 g421 ( .A1(new_n440_), .A2(G116), .ZN(new_n780_) );
  NAND2_X1 g422 ( .A1(new_n779_), .A2(new_n780_), .ZN(new_n781_) );
  NAND2_X1 g423 ( .A1(new_n781_), .A2(KEYINPUT35), .ZN(new_n782_) );
  INV_X1 g424 ( .A(KEYINPUT35), .ZN(new_n783_) );
  NAND3_X1 g425 ( .A1(new_n779_), .A2(new_n780_), .A3(new_n783_), .ZN(new_n784_) );
  NAND2_X1 g426 ( .A1(new_n782_), .A2(new_n784_), .ZN(new_n785_) );
  NAND4_X1 g427 ( .A1(new_n778_), .A2(KEYINPUT36), .A3(new_n776_), .A4(new_n785_), .ZN(new_n786_) );
  INV_X1 g428 ( .A(KEYINPUT36), .ZN(new_n787_) );
  NAND3_X1 g429 ( .A1(new_n778_), .A2(new_n785_), .A3(new_n776_), .ZN(new_n788_) );
  NAND2_X1 g430 ( .A1(new_n788_), .A2(new_n787_), .ZN(new_n789_) );
  NAND2_X1 g431 ( .A1(new_n789_), .A2(new_n786_), .ZN(new_n790_) );
  NAND2_X1 g432 ( .A1(G2067), .A2(KEYINPUT37), .ZN(new_n791_) );
  INV_X1 g433 ( .A(new_n791_), .ZN(new_n792_) );
  NOR2_X1 g434 ( .A1(G2067), .A2(KEYINPUT37), .ZN(new_n793_) );
  NOR2_X1 g435 ( .A1(new_n792_), .A2(new_n793_), .ZN(new_n794_) );
  INV_X1 g436 ( .A(new_n794_), .ZN(new_n795_) );
  NAND2_X1 g437 ( .A1(new_n790_), .A2(new_n795_), .ZN(new_n796_) );
  INV_X1 g438 ( .A(new_n790_), .ZN(new_n797_) );
  NAND2_X1 g439 ( .A1(new_n797_), .A2(new_n794_), .ZN(new_n798_) );
  INV_X1 g440 ( .A(new_n798_), .ZN(new_n799_) );
  NAND4_X1 g441 ( .A1(new_n764_), .A2(new_n765_), .A3(KEYINPUT51), .A4(new_n766_), .ZN(new_n800_) );
  INV_X1 g442 ( .A(new_n800_), .ZN(new_n801_) );
  NOR2_X1 g443 ( .A1(new_n763_), .A2(new_n703_), .ZN(new_n802_) );
  NAND2_X1 g444 ( .A1(new_n429_), .A2(G131), .ZN(new_n803_) );
  INV_X1 g445 ( .A(new_n803_), .ZN(new_n804_) );
  NAND2_X1 g446 ( .A1(new_n431_), .A2(G119), .ZN(new_n805_) );
  NAND2_X1 g447 ( .A1(new_n437_), .A2(G95), .ZN(new_n806_) );
  NAND2_X1 g448 ( .A1(new_n440_), .A2(G107), .ZN(new_n807_) );
  NAND3_X1 g449 ( .A1(new_n805_), .A2(new_n806_), .A3(new_n807_), .ZN(new_n808_) );
  NOR2_X1 g450 ( .A1(new_n804_), .A2(new_n808_), .ZN(new_n809_) );
  NOR2_X1 g451 ( .A1(new_n809_), .A2(new_n701_), .ZN(new_n810_) );
  NOR2_X1 g452 ( .A1(new_n802_), .A2(new_n810_), .ZN(new_n811_) );
  INV_X1 g453 ( .A(new_n811_), .ZN(new_n812_) );
  NAND2_X1 g454 ( .A1(new_n426_), .A2(G2084), .ZN(new_n813_) );
  INV_X1 g455 ( .A(G2084), .ZN(new_n814_) );
  NAND2_X1 g456 ( .A1(G160), .A2(new_n814_), .ZN(new_n815_) );
  NAND2_X1 g457 ( .A1(new_n809_), .A2(new_n701_), .ZN(new_n816_) );
  NAND4_X1 g458 ( .A1(new_n816_), .A2(new_n607_), .A3(new_n813_), .A4(new_n815_), .ZN(new_n817_) );
  NOR4_X1 g459 ( .A1(new_n799_), .A2(new_n801_), .A3(new_n812_), .A4(new_n817_), .ZN(new_n818_) );
  NAND4_X1 g460 ( .A1(new_n818_), .A2(new_n728_), .A3(new_n772_), .A4(new_n796_), .ZN(new_n819_) );
  NAND3_X1 g461 ( .A1(new_n818_), .A2(new_n772_), .A3(new_n796_), .ZN(new_n820_) );
  NAND2_X1 g462 ( .A1(new_n820_), .A2(KEYINPUT52), .ZN(new_n821_) );
  NAND3_X1 g463 ( .A1(new_n821_), .A2(new_n727_), .A3(new_n819_), .ZN(new_n822_) );
  NAND2_X1 g464 ( .A1(new_n822_), .A2(G29), .ZN(new_n823_) );
  NAND2_X1 g465 ( .A1(G168), .A2(G1966), .ZN(new_n824_) );
  NAND2_X1 g466 ( .A1(new_n539_), .A2(new_n691_), .ZN(new_n825_) );
  NAND2_X1 g467 ( .A1(new_n825_), .A2(new_n824_), .ZN(new_n826_) );
  NOR2_X1 g468 ( .A1(G305), .A2(G1981), .ZN(new_n827_) );
  INV_X1 g469 ( .A(new_n827_), .ZN(new_n828_) );
  NAND2_X1 g470 ( .A1(G305), .A2(G1981), .ZN(new_n829_) );
  NAND2_X1 g471 ( .A1(new_n828_), .A2(new_n829_), .ZN(new_n830_) );
  INV_X1 g472 ( .A(new_n830_), .ZN(new_n831_) );
  NAND2_X1 g473 ( .A1(new_n831_), .A2(new_n826_), .ZN(new_n832_) );
  NAND2_X1 g474 ( .A1(new_n832_), .A2(KEYINPUT57), .ZN(new_n833_) );
  INV_X1 g475 ( .A(KEYINPUT57), .ZN(new_n834_) );
  NAND3_X1 g476 ( .A1(new_n831_), .A2(new_n826_), .A3(new_n834_), .ZN(new_n835_) );
  NAND2_X1 g477 ( .A1(new_n833_), .A2(new_n835_), .ZN(new_n836_) );
  NAND2_X1 g478 ( .A1(G171), .A2(new_n716_), .ZN(new_n837_) );
  NAND2_X1 g479 ( .A1(new_n525_), .A2(new_n619_), .ZN(new_n838_) );
  NAND2_X1 g480 ( .A1(G301), .A2(G1961), .ZN(new_n839_) );
  NAND2_X1 g481 ( .A1(new_n524_), .A2(G1341), .ZN(new_n840_) );
  NAND4_X1 g482 ( .A1(new_n838_), .A2(new_n837_), .A3(new_n839_), .A4(new_n840_), .ZN(new_n841_) );
  NAND2_X1 g483 ( .A1(new_n575_), .A2(G1348), .ZN(new_n842_) );
  NAND2_X1 g484 ( .A1(new_n576_), .A2(new_n620_), .ZN(new_n843_) );
  NAND2_X1 g485 ( .A1(new_n843_), .A2(new_n842_), .ZN(new_n844_) );
  NAND2_X1 g486 ( .A1(G166), .A2(new_n711_), .ZN(new_n845_) );
  INV_X1 g487 ( .A(G288), .ZN(new_n846_) );
  NAND2_X1 g488 ( .A1(new_n846_), .A2(new_n686_), .ZN(new_n847_) );
  NAND2_X1 g489 ( .A1(new_n845_), .A2(new_n847_), .ZN(new_n848_) );
  NOR2_X1 g490 ( .A1(new_n846_), .A2(new_n686_), .ZN(new_n849_) );
  NAND2_X1 g491 ( .A1(G303), .A2(G1971), .ZN(new_n850_) );
  INV_X1 g492 ( .A(new_n850_), .ZN(new_n851_) );
  NOR3_X1 g493 ( .A1(new_n848_), .A2(new_n851_), .A3(new_n849_), .ZN(new_n852_) );
  NAND2_X1 g494 ( .A1(new_n581_), .A2(G1956), .ZN(new_n853_) );
  NAND2_X1 g495 ( .A1(G299), .A2(new_n690_), .ZN(new_n854_) );
  NAND2_X1 g496 ( .A1(new_n853_), .A2(new_n854_), .ZN(new_n855_) );
  INV_X1 g497 ( .A(G290), .ZN(new_n856_) );
  NAND2_X1 g498 ( .A1(new_n856_), .A2(new_n717_), .ZN(new_n857_) );
  NAND2_X1 g499 ( .A1(G290), .A2(G1986), .ZN(new_n858_) );
  NAND2_X1 g500 ( .A1(new_n857_), .A2(new_n858_), .ZN(new_n859_) );
  INV_X1 g501 ( .A(new_n859_), .ZN(new_n860_) );
  NAND4_X1 g502 ( .A1(new_n844_), .A2(new_n852_), .A3(new_n855_), .A4(new_n860_), .ZN(new_n861_) );
  NOR2_X1 g503 ( .A1(new_n861_), .A2(new_n841_), .ZN(new_n862_) );
  NAND2_X1 g504 ( .A1(new_n836_), .A2(new_n862_), .ZN(new_n863_) );
  NAND2_X1 g505 ( .A1(G16), .A2(KEYINPUT56), .ZN(new_n864_) );
  INV_X1 g506 ( .A(G16), .ZN(new_n865_) );
  INV_X1 g507 ( .A(KEYINPUT56), .ZN(new_n866_) );
  NAND2_X1 g508 ( .A1(new_n865_), .A2(new_n866_), .ZN(new_n867_) );
  NAND2_X1 g509 ( .A1(new_n867_), .A2(new_n864_), .ZN(new_n868_) );
  NAND2_X1 g510 ( .A1(new_n863_), .A2(new_n868_), .ZN(new_n869_) );
  INV_X1 g511 ( .A(G29), .ZN(new_n870_) );
  NAND2_X1 g512 ( .A1(G33), .A2(G2072), .ZN(new_n871_) );
  NAND2_X1 g513 ( .A1(new_n871_), .A2(G28), .ZN(new_n872_) );
  NAND2_X1 g514 ( .A1(G25), .A2(G1991), .ZN(new_n873_) );
  INV_X1 g515 ( .A(G25), .ZN(new_n874_) );
  NAND2_X1 g516 ( .A1(new_n874_), .A2(new_n701_), .ZN(new_n875_) );
  NAND2_X1 g517 ( .A1(G32), .A2(G1996), .ZN(new_n876_) );
  INV_X1 g518 ( .A(G32), .ZN(new_n877_) );
  NAND2_X1 g519 ( .A1(new_n877_), .A2(new_n703_), .ZN(new_n878_) );
  NAND4_X1 g520 ( .A1(new_n875_), .A2(new_n878_), .A3(new_n873_), .A4(new_n876_), .ZN(new_n879_) );
  NAND2_X1 g521 ( .A1(G2078), .A2(KEYINPUT25), .ZN(new_n880_) );
  INV_X1 g522 ( .A(new_n880_), .ZN(new_n881_) );
  NOR2_X1 g523 ( .A1(G2078), .A2(KEYINPUT25), .ZN(new_n882_) );
  NOR2_X1 g524 ( .A1(new_n881_), .A2(new_n882_), .ZN(new_n883_) );
  NAND2_X1 g525 ( .A1(new_n883_), .A2(G27), .ZN(new_n884_) );
  NOR2_X1 g526 ( .A1(new_n883_), .A2(G27), .ZN(new_n885_) );
  NOR2_X1 g527 ( .A1(G26), .A2(G2067), .ZN(new_n886_) );
  NOR2_X1 g528 ( .A1(G33), .A2(G2072), .ZN(new_n887_) );
  NAND2_X1 g529 ( .A1(G26), .A2(G2067), .ZN(new_n888_) );
  INV_X1 g530 ( .A(new_n888_), .ZN(new_n889_) );
  NOR4_X1 g531 ( .A1(new_n885_), .A2(new_n886_), .A3(new_n887_), .A4(new_n889_), .ZN(new_n890_) );
  NAND2_X1 g532 ( .A1(new_n890_), .A2(new_n884_), .ZN(new_n891_) );
  NOR3_X1 g533 ( .A1(new_n891_), .A2(new_n872_), .A3(new_n879_), .ZN(new_n892_) );
  NOR2_X1 g534 ( .A1(new_n892_), .A2(KEYINPUT53), .ZN(new_n893_) );
  INV_X1 g535 ( .A(new_n893_), .ZN(new_n894_) );
  NAND2_X1 g536 ( .A1(new_n892_), .A2(KEYINPUT53), .ZN(new_n895_) );
  INV_X1 g537 ( .A(KEYINPUT54), .ZN(new_n896_) );
  NAND2_X1 g538 ( .A1(new_n896_), .A2(G2084), .ZN(new_n897_) );
  NAND2_X1 g539 ( .A1(new_n814_), .A2(KEYINPUT54), .ZN(new_n898_) );
  NAND2_X1 g540 ( .A1(new_n897_), .A2(new_n898_), .ZN(new_n899_) );
  NAND2_X1 g541 ( .A1(new_n899_), .A2(G34), .ZN(new_n900_) );
  INV_X1 g542 ( .A(G34), .ZN(new_n901_) );
  NAND3_X1 g543 ( .A1(new_n897_), .A2(new_n898_), .A3(new_n901_), .ZN(new_n902_) );
  NAND2_X1 g544 ( .A1(new_n900_), .A2(new_n902_), .ZN(new_n903_) );
  NAND2_X1 g545 ( .A1(new_n653_), .A2(G35), .ZN(new_n904_) );
  INV_X1 g546 ( .A(G35), .ZN(new_n905_) );
  NAND2_X1 g547 ( .A1(new_n905_), .A2(G2090), .ZN(new_n906_) );
  NAND2_X1 g548 ( .A1(new_n904_), .A2(new_n906_), .ZN(new_n907_) );
  NAND4_X1 g549 ( .A1(new_n894_), .A2(new_n895_), .A3(new_n903_), .A4(new_n907_), .ZN(new_n908_) );
  INV_X1 g550 ( .A(new_n908_), .ZN(new_n909_) );
  NAND2_X1 g551 ( .A1(new_n909_), .A2(new_n727_), .ZN(new_n910_) );
  NAND2_X1 g552 ( .A1(new_n908_), .A2(KEYINPUT55), .ZN(new_n911_) );
  NAND3_X1 g553 ( .A1(new_n910_), .A2(new_n870_), .A3(new_n911_), .ZN(new_n912_) );
  INV_X1 g554 ( .A(KEYINPUT61), .ZN(new_n913_) );
  NAND2_X1 g555 ( .A1(G20), .A2(G1956), .ZN(new_n914_) );
  NOR2_X1 g556 ( .A1(G20), .A2(G1956), .ZN(new_n915_) );
  INV_X1 g557 ( .A(new_n915_), .ZN(new_n916_) );
  NAND2_X1 g558 ( .A1(new_n916_), .A2(new_n914_), .ZN(new_n917_) );
  NAND2_X1 g559 ( .A1(G6), .A2(G1981), .ZN(new_n918_) );
  NAND2_X1 g560 ( .A1(G19), .A2(G1341), .ZN(new_n919_) );
  NOR2_X1 g561 ( .A1(G19), .A2(G1341), .ZN(new_n920_) );
  NOR2_X1 g562 ( .A1(G6), .A2(G1981), .ZN(new_n921_) );
  NOR2_X1 g563 ( .A1(new_n920_), .A2(new_n921_), .ZN(new_n922_) );
  NAND3_X1 g564 ( .A1(new_n922_), .A2(new_n918_), .A3(new_n919_), .ZN(new_n923_) );
  INV_X1 g565 ( .A(KEYINPUT59), .ZN(new_n924_) );
  NAND2_X1 g566 ( .A1(new_n924_), .A2(G1348), .ZN(new_n925_) );
  NAND2_X1 g567 ( .A1(new_n620_), .A2(KEYINPUT59), .ZN(new_n926_) );
  NAND2_X1 g568 ( .A1(new_n925_), .A2(new_n926_), .ZN(new_n927_) );
  NAND2_X1 g569 ( .A1(new_n927_), .A2(G4), .ZN(new_n928_) );
  INV_X1 g570 ( .A(G4), .ZN(new_n929_) );
  NAND3_X1 g571 ( .A1(new_n925_), .A2(new_n926_), .A3(new_n929_), .ZN(new_n930_) );
  NAND2_X1 g572 ( .A1(new_n928_), .A2(new_n930_), .ZN(new_n931_) );
  NOR3_X1 g573 ( .A1(new_n931_), .A2(new_n917_), .A3(new_n923_), .ZN(new_n932_) );
  NAND2_X1 g574 ( .A1(new_n932_), .A2(KEYINPUT60), .ZN(new_n933_) );
  INV_X1 g575 ( .A(KEYINPUT60), .ZN(new_n934_) );
  INV_X1 g576 ( .A(new_n932_), .ZN(new_n935_) );
  NAND2_X1 g577 ( .A1(new_n935_), .A2(new_n934_), .ZN(new_n936_) );
  NAND2_X1 g578 ( .A1(new_n936_), .A2(new_n933_), .ZN(new_n937_) );
  INV_X1 g579 ( .A(KEYINPUT58), .ZN(new_n938_) );
  INV_X1 g580 ( .A(G24), .ZN(new_n939_) );
  NOR2_X1 g581 ( .A1(new_n939_), .A2(G1986), .ZN(new_n940_) );
  NOR2_X1 g582 ( .A1(new_n717_), .A2(G24), .ZN(new_n941_) );
  NOR2_X1 g583 ( .A1(new_n940_), .A2(new_n941_), .ZN(new_n942_) );
  INV_X1 g584 ( .A(new_n942_), .ZN(new_n943_) );
  NAND2_X1 g585 ( .A1(G23), .A2(G1976), .ZN(new_n944_) );
  INV_X1 g586 ( .A(new_n944_), .ZN(new_n945_) );
  NOR2_X1 g587 ( .A1(G23), .A2(G1976), .ZN(new_n946_) );
  NOR2_X1 g588 ( .A1(new_n945_), .A2(new_n946_), .ZN(new_n947_) );
  NAND2_X1 g589 ( .A1(G22), .A2(G1971), .ZN(new_n948_) );
  INV_X1 g590 ( .A(new_n948_), .ZN(new_n949_) );
  NOR2_X1 g591 ( .A1(G22), .A2(G1971), .ZN(new_n950_) );
  NOR2_X1 g592 ( .A1(new_n949_), .A2(new_n950_), .ZN(new_n951_) );
  NAND4_X1 g593 ( .A1(new_n943_), .A2(new_n938_), .A3(new_n947_), .A4(new_n951_), .ZN(new_n952_) );
  NAND3_X1 g594 ( .A1(new_n943_), .A2(new_n947_), .A3(new_n951_), .ZN(new_n953_) );
  NAND2_X1 g595 ( .A1(new_n953_), .A2(KEYINPUT58), .ZN(new_n954_) );
  NAND2_X1 g596 ( .A1(G5), .A2(G1961), .ZN(new_n955_) );
  INV_X1 g597 ( .A(G5), .ZN(new_n956_) );
  NAND2_X1 g598 ( .A1(new_n956_), .A2(new_n716_), .ZN(new_n957_) );
  NAND2_X1 g599 ( .A1(G21), .A2(G1966), .ZN(new_n958_) );
  INV_X1 g600 ( .A(G21), .ZN(new_n959_) );
  NAND2_X1 g601 ( .A1(new_n959_), .A2(new_n691_), .ZN(new_n960_) );
  NAND4_X1 g602 ( .A1(new_n957_), .A2(new_n960_), .A3(new_n955_), .A4(new_n958_), .ZN(new_n961_) );
  INV_X1 g603 ( .A(new_n961_), .ZN(new_n962_) );
  NAND3_X1 g604 ( .A1(new_n954_), .A2(new_n952_), .A3(new_n962_), .ZN(new_n963_) );
  INV_X1 g605 ( .A(new_n963_), .ZN(new_n964_) );
  NAND3_X1 g606 ( .A1(new_n937_), .A2(new_n913_), .A3(new_n964_), .ZN(new_n965_) );
  NAND2_X1 g607 ( .A1(new_n937_), .A2(new_n964_), .ZN(new_n966_) );
  NAND2_X1 g608 ( .A1(new_n966_), .A2(KEYINPUT61), .ZN(new_n967_) );
  NAND3_X1 g609 ( .A1(new_n967_), .A2(new_n865_), .A3(new_n965_), .ZN(new_n968_) );
  NAND3_X1 g610 ( .A1(new_n912_), .A2(G11), .A3(new_n968_), .ZN(new_n969_) );
  INV_X1 g611 ( .A(new_n969_), .ZN(new_n970_) );
  NAND4_X1 g612 ( .A1(new_n823_), .A2(KEYINPUT62), .A3(new_n869_), .A4(new_n970_), .ZN(new_n971_) );
  INV_X1 g613 ( .A(KEYINPUT62), .ZN(new_n972_) );
  NAND3_X1 g614 ( .A1(new_n823_), .A2(new_n869_), .A3(new_n970_), .ZN(new_n973_) );
  NAND2_X1 g615 ( .A1(new_n973_), .A2(new_n972_), .ZN(new_n974_) );
  NAND2_X1 g616 ( .A1(new_n974_), .A2(new_n971_), .ZN(G311) );
  INV_X1 g617 ( .A(G311), .ZN(G150) );
  NAND2_X1 g618 ( .A1(new_n575_), .A2(G559), .ZN(new_n977_) );
  INV_X1 g619 ( .A(new_n977_), .ZN(new_n978_) );
  NAND2_X1 g620 ( .A1(new_n978_), .A2(new_n525_), .ZN(new_n979_) );
  NAND2_X1 g621 ( .A1(new_n977_), .A2(new_n524_), .ZN(new_n980_) );
  NAND3_X1 g622 ( .A1(new_n979_), .A2(new_n586_), .A3(new_n980_), .ZN(new_n981_) );
  NAND2_X1 g623 ( .A1(new_n465_), .A2(G80), .ZN(new_n982_) );
  NAND2_X1 g624 ( .A1(new_n462_), .A2(G93), .ZN(new_n983_) );
  NAND2_X1 g625 ( .A1(new_n460_), .A2(G55), .ZN(new_n984_) );
  NAND2_X1 g626 ( .A1(new_n471_), .A2(G67), .ZN(new_n985_) );
  NAND4_X1 g627 ( .A1(new_n982_), .A2(new_n984_), .A3(new_n983_), .A4(new_n985_), .ZN(new_n986_) );
  NAND2_X1 g628 ( .A1(new_n981_), .A2(new_n986_), .ZN(new_n987_) );
  INV_X1 g629 ( .A(new_n986_), .ZN(new_n988_) );
  NAND4_X1 g630 ( .A1(new_n979_), .A2(new_n586_), .A3(new_n980_), .A4(new_n988_), .ZN(new_n989_) );
  NAND2_X1 g631 ( .A1(new_n987_), .A2(new_n989_), .ZN(G145) );
  INV_X1 g632 ( .A(G37), .ZN(new_n991_) );
  NAND2_X1 g633 ( .A1(new_n429_), .A2(G142), .ZN(new_n992_) );
  NAND2_X1 g634 ( .A1(new_n437_), .A2(G106), .ZN(new_n993_) );
  NAND3_X1 g635 ( .A1(new_n992_), .A2(KEYINPUT45), .A3(new_n993_), .ZN(new_n994_) );
  INV_X1 g636 ( .A(KEYINPUT45), .ZN(new_n995_) );
  NAND2_X1 g637 ( .A1(new_n992_), .A2(new_n993_), .ZN(new_n996_) );
  NAND2_X1 g638 ( .A1(new_n996_), .A2(new_n995_), .ZN(new_n997_) );
  NAND2_X1 g639 ( .A1(new_n431_), .A2(G130), .ZN(new_n998_) );
  NAND2_X1 g640 ( .A1(new_n440_), .A2(G118), .ZN(new_n999_) );
  NAND4_X1 g641 ( .A1(new_n997_), .A2(new_n994_), .A3(new_n998_), .A4(new_n999_), .ZN(new_n1000_) );
  INV_X1 g642 ( .A(new_n1000_), .ZN(new_n1001_) );
  NAND2_X1 g643 ( .A1(new_n1001_), .A2(new_n762_), .ZN(new_n1002_) );
  NAND2_X1 g644 ( .A1(new_n1000_), .A2(new_n763_), .ZN(new_n1003_) );
  NAND2_X1 g645 ( .A1(new_n1002_), .A2(new_n1003_), .ZN(new_n1004_) );
  NAND2_X1 g646 ( .A1(new_n1004_), .A2(G162), .ZN(new_n1005_) );
  NAND3_X1 g647 ( .A1(new_n1002_), .A2(new_n444_), .A3(new_n1003_), .ZN(new_n1006_) );
  NAND2_X1 g648 ( .A1(new_n1005_), .A2(new_n1006_), .ZN(new_n1007_) );
  NOR2_X1 g649 ( .A1(new_n742_), .A2(new_n426_), .ZN(new_n1008_) );
  NAND2_X1 g650 ( .A1(new_n742_), .A2(new_n426_), .ZN(new_n1009_) );
  INV_X1 g651 ( .A(new_n1009_), .ZN(new_n1010_) );
  NOR2_X1 g652 ( .A1(new_n1010_), .A2(new_n1008_), .ZN(new_n1011_) );
  INV_X1 g653 ( .A(new_n1011_), .ZN(new_n1012_) );
  NAND2_X1 g654 ( .A1(new_n1012_), .A2(new_n790_), .ZN(new_n1013_) );
  NAND2_X1 g655 ( .A1(new_n797_), .A2(new_n1011_), .ZN(new_n1014_) );
  NAND2_X1 g656 ( .A1(new_n1014_), .A2(new_n1013_), .ZN(new_n1015_) );
  NAND2_X1 g657 ( .A1(new_n1007_), .A2(new_n1015_), .ZN(new_n1016_) );
  NAND4_X1 g658 ( .A1(new_n1005_), .A2(new_n1014_), .A3(new_n1006_), .A4(new_n1013_), .ZN(new_n1017_) );
  NAND2_X1 g659 ( .A1(new_n1016_), .A2(new_n1017_), .ZN(new_n1018_) );
  INV_X1 g660 ( .A(new_n809_), .ZN(new_n1019_) );
  NAND2_X1 g661 ( .A1(new_n1019_), .A2(new_n607_), .ZN(new_n1020_) );
  NAND2_X1 g662 ( .A1(new_n610_), .A2(new_n809_), .ZN(new_n1021_) );
  NAND2_X1 g663 ( .A1(new_n1020_), .A2(new_n1021_), .ZN(new_n1022_) );
  INV_X1 g664 ( .A(KEYINPUT48), .ZN(new_n1023_) );
  NOR2_X1 g665 ( .A1(new_n1023_), .A2(KEYINPUT46), .ZN(new_n1024_) );
  NAND2_X1 g666 ( .A1(new_n1023_), .A2(KEYINPUT46), .ZN(new_n1025_) );
  INV_X1 g667 ( .A(new_n1025_), .ZN(new_n1026_) );
  NOR2_X1 g668 ( .A1(new_n1026_), .A2(new_n1024_), .ZN(new_n1027_) );
  INV_X1 g669 ( .A(new_n1027_), .ZN(new_n1028_) );
  NAND2_X1 g670 ( .A1(new_n1022_), .A2(new_n1028_), .ZN(new_n1029_) );
  NAND3_X1 g671 ( .A1(new_n1020_), .A2(new_n1021_), .A3(new_n1027_), .ZN(new_n1030_) );
  NAND2_X1 g672 ( .A1(new_n1029_), .A2(new_n1030_), .ZN(new_n1031_) );
  NAND2_X1 g673 ( .A1(new_n1031_), .A2(G164), .ZN(new_n1032_) );
  NAND3_X1 g674 ( .A1(new_n1029_), .A2(new_n452_), .A3(new_n1030_), .ZN(new_n1033_) );
  NAND2_X1 g675 ( .A1(new_n1032_), .A2(new_n1033_), .ZN(new_n1034_) );
  NAND2_X1 g676 ( .A1(new_n1018_), .A2(new_n1034_), .ZN(new_n1035_) );
  NAND4_X1 g677 ( .A1(new_n1016_), .A2(new_n1017_), .A3(new_n1032_), .A4(new_n1033_), .ZN(new_n1036_) );
  NAND3_X1 g678 ( .A1(new_n1035_), .A2(new_n991_), .A3(new_n1036_), .ZN(new_n1037_) );
  INV_X1 g679 ( .A(new_n1037_), .ZN(G395) );
  NAND2_X1 g680 ( .A1(new_n524_), .A2(new_n856_), .ZN(new_n1039_) );
  NAND2_X1 g681 ( .A1(new_n525_), .A2(G290), .ZN(new_n1040_) );
  NAND2_X1 g682 ( .A1(new_n1040_), .A2(new_n1039_), .ZN(new_n1041_) );
  NAND2_X1 g683 ( .A1(new_n1041_), .A2(new_n846_), .ZN(new_n1042_) );
  NAND3_X1 g684 ( .A1(new_n1040_), .A2(G288), .A3(new_n1039_), .ZN(new_n1043_) );
  NAND2_X1 g685 ( .A1(new_n1042_), .A2(new_n1043_), .ZN(new_n1044_) );
  INV_X1 g686 ( .A(G305), .ZN(new_n1045_) );
  NAND2_X1 g687 ( .A1(new_n581_), .A2(KEYINPUT19), .ZN(new_n1046_) );
  INV_X1 g688 ( .A(KEYINPUT19), .ZN(new_n1047_) );
  NAND2_X1 g689 ( .A1(G299), .A2(new_n1047_), .ZN(new_n1048_) );
  NAND2_X1 g690 ( .A1(new_n1046_), .A2(new_n1048_), .ZN(new_n1049_) );
  NAND2_X1 g691 ( .A1(new_n1045_), .A2(new_n1049_), .ZN(new_n1050_) );
  NAND3_X1 g692 ( .A1(G305), .A2(new_n1046_), .A3(new_n1048_), .ZN(new_n1051_) );
  NAND2_X1 g693 ( .A1(new_n1050_), .A2(new_n1051_), .ZN(new_n1052_) );
  NAND2_X1 g694 ( .A1(new_n1044_), .A2(new_n1052_), .ZN(new_n1053_) );
  NAND4_X1 g695 ( .A1(new_n1042_), .A2(new_n1050_), .A3(new_n1043_), .A4(new_n1051_), .ZN(new_n1054_) );
  NAND2_X1 g696 ( .A1(new_n1053_), .A2(new_n1054_), .ZN(new_n1055_) );
  NOR2_X1 g697 ( .A1(G303), .A2(new_n986_), .ZN(new_n1056_) );
  NAND2_X1 g698 ( .A1(G303), .A2(new_n986_), .ZN(new_n1057_) );
  INV_X1 g699 ( .A(new_n1057_), .ZN(new_n1058_) );
  NOR2_X1 g700 ( .A1(new_n1058_), .A2(new_n1056_), .ZN(new_n1059_) );
  INV_X1 g701 ( .A(new_n1059_), .ZN(new_n1060_) );
  NAND2_X1 g702 ( .A1(new_n1055_), .A2(new_n1060_), .ZN(new_n1061_) );
  NAND3_X1 g703 ( .A1(new_n1053_), .A2(new_n1054_), .A3(new_n1059_), .ZN(new_n1062_) );
  NAND2_X1 g704 ( .A1(new_n1061_), .A2(new_n1062_), .ZN(new_n1063_) );
  NAND2_X1 g705 ( .A1(new_n1063_), .A2(new_n978_), .ZN(new_n1064_) );
  INV_X1 g706 ( .A(new_n1063_), .ZN(new_n1065_) );
  NAND2_X1 g707 ( .A1(new_n1065_), .A2(new_n977_), .ZN(new_n1066_) );
  NAND2_X1 g708 ( .A1(new_n1066_), .A2(new_n1064_), .ZN(new_n1067_) );
  NAND2_X1 g709 ( .A1(new_n1067_), .A2(G868), .ZN(new_n1068_) );
  NAND2_X1 g710 ( .A1(new_n986_), .A2(new_n564_), .ZN(new_n1069_) );
  NAND2_X1 g711 ( .A1(new_n1068_), .A2(new_n1069_), .ZN(G295) );
  NAND2_X1 g712 ( .A1(G286), .A2(new_n576_), .ZN(new_n1071_) );
  NAND2_X1 g713 ( .A1(new_n579_), .A2(new_n575_), .ZN(new_n1072_) );
  NAND2_X1 g714 ( .A1(new_n1072_), .A2(new_n1071_), .ZN(new_n1073_) );
  NAND2_X1 g715 ( .A1(new_n1063_), .A2(new_n1073_), .ZN(new_n1074_) );
  NAND3_X1 g716 ( .A1(new_n1065_), .A2(new_n1071_), .A3(new_n1072_), .ZN(new_n1075_) );
  NAND2_X1 g717 ( .A1(new_n1075_), .A2(new_n1074_), .ZN(new_n1076_) );
  NAND2_X1 g718 ( .A1(new_n1076_), .A2(G301), .ZN(new_n1077_) );
  NAND3_X1 g719 ( .A1(new_n1075_), .A2(G171), .A3(new_n1074_), .ZN(new_n1078_) );
  NAND3_X1 g720 ( .A1(new_n1077_), .A2(new_n991_), .A3(new_n1078_), .ZN(new_n1079_) );
  INV_X1 g721 ( .A(new_n1079_), .ZN(G397) );
  INV_X1 g722 ( .A(KEYINPUT33), .ZN(new_n1081_) );
  INV_X1 g723 ( .A(new_n848_), .ZN(new_n1082_) );
  INV_X1 g724 ( .A(KEYINPUT29), .ZN(new_n1083_) );
  NAND4_X1 g725 ( .A1(new_n425_), .A2(G40), .A3(new_n418_), .A4(new_n420_), .ZN(new_n1084_) );
  INV_X1 g726 ( .A(G1384), .ZN(new_n1085_) );
  NAND2_X1 g727 ( .A1(new_n452_), .A2(new_n1085_), .ZN(new_n1086_) );
  NOR2_X1 g728 ( .A1(new_n1086_), .A2(new_n1084_), .ZN(new_n1087_) );
  NAND3_X1 g729 ( .A1(new_n1087_), .A2(G1996), .A3(KEYINPUT26), .ZN(new_n1088_) );
  INV_X1 g730 ( .A(KEYINPUT26), .ZN(new_n1089_) );
  NAND2_X1 g731 ( .A1(new_n1087_), .A2(G1996), .ZN(new_n1090_) );
  NAND2_X1 g732 ( .A1(new_n1090_), .A2(new_n1089_), .ZN(new_n1091_) );
  NOR2_X1 g733 ( .A1(new_n1087_), .A2(new_n619_), .ZN(new_n1092_) );
  NOR2_X1 g734 ( .A1(new_n1092_), .A2(new_n524_), .ZN(new_n1093_) );
  NAND4_X1 g735 ( .A1(new_n1093_), .A2(new_n575_), .A3(new_n1088_), .A4(new_n1091_), .ZN(new_n1094_) );
  INV_X1 g736 ( .A(new_n1087_), .ZN(new_n1095_) );
  NAND2_X1 g737 ( .A1(new_n1095_), .A2(G1348), .ZN(new_n1096_) );
  NAND2_X1 g738 ( .A1(new_n1087_), .A2(G2067), .ZN(new_n1097_) );
  NAND2_X1 g739 ( .A1(new_n1096_), .A2(new_n1097_), .ZN(new_n1098_) );
  NAND2_X1 g740 ( .A1(new_n1094_), .A2(new_n1098_), .ZN(new_n1099_) );
  NAND3_X1 g741 ( .A1(new_n1093_), .A2(new_n1088_), .A3(new_n1091_), .ZN(new_n1100_) );
  NAND2_X1 g742 ( .A1(new_n1100_), .A2(new_n576_), .ZN(new_n1101_) );
  NAND2_X1 g743 ( .A1(new_n1099_), .A2(new_n1101_), .ZN(new_n1102_) );
  INV_X1 g744 ( .A(KEYINPUT27), .ZN(new_n1103_) );
  NAND3_X1 g745 ( .A1(new_n1087_), .A2(G2072), .A3(new_n1103_), .ZN(new_n1104_) );
  NAND2_X1 g746 ( .A1(new_n1087_), .A2(G2072), .ZN(new_n1105_) );
  NAND2_X1 g747 ( .A1(new_n1105_), .A2(KEYINPUT27), .ZN(new_n1106_) );
  NAND2_X1 g748 ( .A1(new_n1095_), .A2(G1956), .ZN(new_n1107_) );
  NAND4_X1 g749 ( .A1(new_n1106_), .A2(new_n1107_), .A3(new_n581_), .A4(new_n1104_), .ZN(new_n1108_) );
  NAND2_X1 g750 ( .A1(new_n1102_), .A2(new_n1108_), .ZN(new_n1109_) );
  INV_X1 g751 ( .A(KEYINPUT28), .ZN(new_n1110_) );
  NAND3_X1 g752 ( .A1(new_n1106_), .A2(new_n1104_), .A3(new_n1107_), .ZN(new_n1111_) );
  NAND3_X1 g753 ( .A1(new_n1111_), .A2(new_n1110_), .A3(G299), .ZN(new_n1112_) );
  NAND2_X1 g754 ( .A1(new_n1111_), .A2(G299), .ZN(new_n1113_) );
  NAND2_X1 g755 ( .A1(new_n1113_), .A2(KEYINPUT28), .ZN(new_n1114_) );
  NAND2_X1 g756 ( .A1(new_n1114_), .A2(new_n1112_), .ZN(new_n1115_) );
  NAND2_X1 g757 ( .A1(new_n1109_), .A2(new_n1115_), .ZN(new_n1116_) );
  NAND2_X1 g758 ( .A1(new_n1116_), .A2(new_n1083_), .ZN(new_n1117_) );
  NAND3_X1 g759 ( .A1(new_n1109_), .A2(KEYINPUT29), .A3(new_n1115_), .ZN(new_n1118_) );
  NAND2_X1 g760 ( .A1(new_n1117_), .A2(new_n1118_), .ZN(new_n1119_) );
  NAND2_X1 g761 ( .A1(new_n1095_), .A2(new_n716_), .ZN(new_n1120_) );
  INV_X1 g762 ( .A(new_n883_), .ZN(new_n1121_) );
  NAND2_X1 g763 ( .A1(new_n1087_), .A2(new_n1121_), .ZN(new_n1122_) );
  NAND2_X1 g764 ( .A1(new_n1120_), .A2(new_n1122_), .ZN(new_n1123_) );
  NAND2_X1 g765 ( .A1(new_n1123_), .A2(G171), .ZN(new_n1124_) );
  NAND2_X1 g766 ( .A1(new_n1119_), .A2(new_n1124_), .ZN(new_n1125_) );
  INV_X1 g767 ( .A(KEYINPUT31), .ZN(new_n1126_) );
  INV_X1 g768 ( .A(KEYINPUT30), .ZN(new_n1127_) );
  INV_X1 g769 ( .A(G8), .ZN(new_n1128_) );
  NOR2_X1 g770 ( .A1(new_n1087_), .A2(new_n1128_), .ZN(new_n1129_) );
  NAND2_X1 g771 ( .A1(new_n1129_), .A2(new_n691_), .ZN(new_n1130_) );
  NOR2_X1 g772 ( .A1(new_n1095_), .A2(G2084), .ZN(new_n1131_) );
  NOR2_X1 g773 ( .A1(new_n1131_), .A2(new_n1128_), .ZN(new_n1132_) );
  NAND3_X1 g774 ( .A1(new_n1132_), .A2(new_n1127_), .A3(new_n1130_), .ZN(new_n1133_) );
  NAND2_X1 g775 ( .A1(new_n1132_), .A2(new_n1130_), .ZN(new_n1134_) );
  NAND2_X1 g776 ( .A1(new_n1134_), .A2(KEYINPUT30), .ZN(new_n1135_) );
  NAND3_X1 g777 ( .A1(new_n1135_), .A2(new_n539_), .A3(new_n1133_), .ZN(new_n1136_) );
  NAND3_X1 g778 ( .A1(new_n1120_), .A2(G301), .A3(new_n1122_), .ZN(new_n1137_) );
  NAND3_X1 g779 ( .A1(new_n1136_), .A2(new_n1126_), .A3(new_n1137_), .ZN(new_n1138_) );
  NAND2_X1 g780 ( .A1(new_n1136_), .A2(new_n1137_), .ZN(new_n1139_) );
  NAND2_X1 g781 ( .A1(new_n1139_), .A2(KEYINPUT31), .ZN(new_n1140_) );
  NAND2_X1 g782 ( .A1(new_n1140_), .A2(new_n1138_), .ZN(new_n1141_) );
  NAND2_X1 g783 ( .A1(new_n1125_), .A2(new_n1141_), .ZN(new_n1142_) );
  NAND2_X1 g784 ( .A1(new_n1142_), .A2(G286), .ZN(new_n1143_) );
  NAND2_X1 g785 ( .A1(new_n1129_), .A2(new_n711_), .ZN(new_n1144_) );
  NAND2_X1 g786 ( .A1(new_n1087_), .A2(new_n653_), .ZN(new_n1145_) );
  NAND3_X1 g787 ( .A1(new_n1144_), .A2(G303), .A3(new_n1145_), .ZN(new_n1146_) );
  NAND2_X1 g788 ( .A1(new_n1143_), .A2(new_n1146_), .ZN(new_n1147_) );
  NAND2_X1 g789 ( .A1(new_n1147_), .A2(G8), .ZN(new_n1148_) );
  NAND2_X1 g790 ( .A1(new_n1148_), .A2(KEYINPUT32), .ZN(new_n1149_) );
  INV_X1 g791 ( .A(KEYINPUT32), .ZN(new_n1150_) );
  NAND3_X1 g792 ( .A1(new_n1147_), .A2(G8), .A3(new_n1150_), .ZN(new_n1151_) );
  NAND2_X1 g793 ( .A1(new_n1149_), .A2(new_n1151_), .ZN(new_n1152_) );
  NAND2_X1 g794 ( .A1(new_n1131_), .A2(G8), .ZN(new_n1153_) );
  NAND3_X1 g795 ( .A1(new_n1142_), .A2(new_n1130_), .A3(new_n1153_), .ZN(new_n1154_) );
  NAND2_X1 g796 ( .A1(new_n1152_), .A2(new_n1154_), .ZN(new_n1155_) );
  NAND2_X1 g797 ( .A1(new_n1155_), .A2(new_n1082_), .ZN(new_n1156_) );
  INV_X1 g798 ( .A(new_n849_), .ZN(new_n1157_) );
  NAND2_X1 g799 ( .A1(new_n1157_), .A2(new_n1129_), .ZN(new_n1158_) );
  INV_X1 g800 ( .A(new_n1158_), .ZN(new_n1159_) );
  NAND2_X1 g801 ( .A1(new_n1156_), .A2(new_n1159_), .ZN(new_n1160_) );
  NAND2_X1 g802 ( .A1(new_n1160_), .A2(new_n1081_), .ZN(new_n1161_) );
  INV_X1 g803 ( .A(new_n1129_), .ZN(new_n1162_) );
  NOR3_X1 g804 ( .A1(new_n1162_), .A2(new_n1081_), .A3(new_n847_), .ZN(new_n1163_) );
  NOR2_X1 g805 ( .A1(new_n830_), .A2(new_n1163_), .ZN(new_n1164_) );
  NAND2_X1 g806 ( .A1(new_n1161_), .A2(new_n1164_), .ZN(new_n1165_) );
  NAND3_X1 g807 ( .A1(G166), .A2(G8), .A3(new_n653_), .ZN(new_n1166_) );
  NAND2_X1 g808 ( .A1(new_n1155_), .A2(new_n1166_), .ZN(new_n1167_) );
  NAND2_X1 g809 ( .A1(new_n1167_), .A2(new_n1162_), .ZN(new_n1168_) );
  NAND2_X1 g810 ( .A1(new_n828_), .A2(KEYINPUT24), .ZN(new_n1169_) );
  INV_X1 g811 ( .A(KEYINPUT24), .ZN(new_n1170_) );
  NAND2_X1 g812 ( .A1(new_n827_), .A2(new_n1170_), .ZN(new_n1171_) );
  NAND3_X1 g813 ( .A1(new_n1169_), .A2(new_n1129_), .A3(new_n1171_), .ZN(new_n1172_) );
  NAND2_X1 g814 ( .A1(new_n1168_), .A2(new_n1172_), .ZN(new_n1173_) );
  INV_X1 g815 ( .A(new_n1173_), .ZN(new_n1174_) );
  NAND2_X1 g816 ( .A1(new_n1165_), .A2(new_n1174_), .ZN(new_n1175_) );
  INV_X1 g817 ( .A(new_n1086_), .ZN(new_n1176_) );
  NOR2_X1 g818 ( .A1(new_n1176_), .A2(new_n1084_), .ZN(new_n1177_) );
  NAND2_X1 g819 ( .A1(new_n799_), .A2(new_n1177_), .ZN(new_n1178_) );
  INV_X1 g820 ( .A(new_n1178_), .ZN(new_n1179_) );
  NAND2_X1 g821 ( .A1(new_n812_), .A2(new_n1177_), .ZN(new_n1180_) );
  NAND2_X1 g822 ( .A1(new_n859_), .A2(new_n1177_), .ZN(new_n1181_) );
  NAND2_X1 g823 ( .A1(new_n1180_), .A2(new_n1181_), .ZN(new_n1182_) );
  NOR2_X1 g824 ( .A1(new_n1179_), .A2(new_n1182_), .ZN(new_n1183_) );
  NAND2_X1 g825 ( .A1(new_n1175_), .A2(new_n1183_), .ZN(new_n1184_) );
  INV_X1 g826 ( .A(KEYINPUT39), .ZN(new_n1185_) );
  NAND2_X1 g827 ( .A1(new_n816_), .A2(new_n857_), .ZN(new_n1186_) );
  NAND2_X1 g828 ( .A1(new_n1180_), .A2(new_n1186_), .ZN(new_n1187_) );
  NAND2_X1 g829 ( .A1(new_n1187_), .A2(new_n764_), .ZN(new_n1188_) );
  NAND2_X1 g830 ( .A1(new_n1188_), .A2(new_n1185_), .ZN(new_n1189_) );
  NAND3_X1 g831 ( .A1(new_n1187_), .A2(KEYINPUT39), .A3(new_n764_), .ZN(new_n1190_) );
  NAND2_X1 g832 ( .A1(new_n1189_), .A2(new_n1190_), .ZN(new_n1191_) );
  NAND2_X1 g833 ( .A1(new_n1191_), .A2(new_n1178_), .ZN(new_n1192_) );
  NAND2_X1 g834 ( .A1(new_n1192_), .A2(new_n796_), .ZN(new_n1193_) );
  NAND2_X1 g835 ( .A1(new_n1193_), .A2(new_n1177_), .ZN(new_n1194_) );
  NAND2_X1 g836 ( .A1(new_n1184_), .A2(new_n1194_), .ZN(new_n1195_) );
  NAND2_X1 g837 ( .A1(new_n1195_), .A2(KEYINPUT40), .ZN(new_n1196_) );
  INV_X1 g838 ( .A(KEYINPUT40), .ZN(new_n1197_) );
  NAND3_X1 g839 ( .A1(new_n1184_), .A2(new_n1197_), .A3(new_n1194_), .ZN(new_n1198_) );
  NAND2_X1 g840 ( .A1(new_n1196_), .A2(new_n1198_), .ZN(G329) );
  INV_X1 g841 ( .A(KEYINPUT49), .ZN(new_n1201_) );
  INV_X1 g842 ( .A(G227), .ZN(new_n1202_) );
  NAND2_X1 g843 ( .A1(new_n725_), .A2(new_n1202_), .ZN(new_n1203_) );
  NAND2_X1 g844 ( .A1(new_n1203_), .A2(new_n1201_), .ZN(new_n1204_) );
  NAND3_X1 g845 ( .A1(new_n725_), .A2(KEYINPUT49), .A3(new_n1202_), .ZN(new_n1205_) );
  NAND3_X1 g846 ( .A1(new_n1205_), .A2(G319), .A3(new_n649_), .ZN(new_n1206_) );
  INV_X1 g847 ( .A(new_n1206_), .ZN(new_n1207_) );
  NAND3_X1 g848 ( .A1(new_n1037_), .A2(new_n1204_), .A3(new_n1207_), .ZN(new_n1208_) );
  INV_X1 g849 ( .A(new_n1208_), .ZN(new_n1209_) );
  NAND2_X1 g850 ( .A1(new_n1079_), .A2(new_n1209_), .ZN(G225) );
  INV_X1 g851 ( .A(G225), .ZN(G308) );
  assign   G231 = 1'b0;
  BUF_X1 g852 ( .A(G452), .Z(G350) );
  BUF_X1 g853 ( .A(G452), .Z(G335) );
  BUF_X1 g854 ( .A(G452), .Z(G409) );
  BUF_X1 g855 ( .A(G1083), .Z(G369) );
  BUF_X1 g856 ( .A(G1083), .Z(G367) );
  BUF_X1 g857 ( .A(G2066), .Z(G411) );
  BUF_X1 g858 ( .A(G2066), .Z(G337) );
  BUF_X1 g859 ( .A(G2066), .Z(G384) );
  BUF_X1 g860 ( .A(G452), .Z(G391) );
  NAND2_X1 g861 ( .A1(new_n577_), .A2(new_n563_), .ZN(G321) );
  INV_X1 g862 ( .A(new_n583_), .ZN(G280) );
  INV_X1 g863 ( .A(new_n595_), .ZN(G323) );
  NAND2_X1 g864 ( .A1(new_n1068_), .A2(new_n1069_), .ZN(G331) );
endmodule


