module add_mul_combine_8_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, Result_mul_0_, 
        Result_mul_1_, Result_mul_2_, Result_mul_3_, Result_mul_4_, 
        Result_mul_5_, Result_mul_6_, Result_mul_7_, Result_mul_8_, 
        Result_mul_9_, Result_mul_10_, Result_mul_11_, Result_mul_12_, 
        Result_mul_13_, Result_mul_14_, Result_mul_15_, Result_add_0_, 
        Result_add_1_, Result_add_2_, Result_add_3_, Result_add_4_, 
        Result_add_5_, Result_add_6_, Result_add_7_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_,
         b_4_, b_5_, b_6_, b_7_;
  output Result_mul_0_, Result_mul_1_, Result_mul_2_, Result_mul_3_,
         Result_mul_4_, Result_mul_5_, Result_mul_6_, Result_mul_7_,
         Result_mul_8_, Result_mul_9_, Result_mul_10_, Result_mul_11_,
         Result_mul_12_, Result_mul_13_, Result_mul_14_, Result_mul_15_,
         Result_add_0_, Result_add_1_, Result_add_2_, Result_add_3_,
         Result_add_4_, Result_add_5_, Result_add_6_, Result_add_7_;
  wire   n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941;

  XNOR2_X1 U485 ( .A(n462), .B(n463), .ZN(Result_mul_9_) );
  XNOR2_X1 U486 ( .A(n464), .B(n465), .ZN(n462) );
  NOR2_X1 U487 ( .A1(n466), .A2(n467), .ZN(n465) );
  XNOR2_X1 U488 ( .A(n468), .B(n469), .ZN(Result_mul_8_) );
  NAND2_X1 U489 ( .A1(n470), .A2(n471), .ZN(n468) );
  XNOR2_X1 U490 ( .A(n472), .B(n473), .ZN(Result_mul_7_) );
  NOR2_X1 U491 ( .A1(n474), .A2(n475), .ZN(Result_mul_6_) );
  NOR2_X1 U492 ( .A1(n476), .A2(n477), .ZN(n475) );
  XNOR2_X1 U493 ( .A(n474), .B(n478), .ZN(Result_mul_5_) );
  NAND2_X1 U494 ( .A1(n479), .A2(n480), .ZN(n478) );
  NAND2_X1 U495 ( .A1(n481), .A2(n482), .ZN(n480) );
  INV_X1 U496 ( .A(n483), .ZN(n479) );
  XNOR2_X1 U497 ( .A(n484), .B(n485), .ZN(Result_mul_4_) );
  XOR2_X1 U498 ( .A(n486), .B(n487), .Z(Result_mul_3_) );
  NOR2_X1 U499 ( .A1(n488), .A2(n485), .ZN(n487) );
  INV_X1 U500 ( .A(n484), .ZN(n488) );
  NOR2_X1 U501 ( .A1(n489), .A2(n490), .ZN(n486) );
  NOR2_X1 U502 ( .A1(n491), .A2(n492), .ZN(n490) );
  XOR2_X1 U503 ( .A(n493), .B(n494), .Z(Result_mul_2_) );
  XNOR2_X1 U504 ( .A(n495), .B(n496), .ZN(Result_mul_1_) );
  NOR2_X1 U505 ( .A1(n497), .A2(n498), .ZN(n496) );
  XNOR2_X1 U506 ( .A(n499), .B(n500), .ZN(Result_mul_14_) );
  NAND2_X1 U507 ( .A1(b_7_), .A2(a_6_), .ZN(n500) );
  XOR2_X1 U508 ( .A(n501), .B(n502), .Z(Result_mul_13_) );
  XNOR2_X1 U509 ( .A(n503), .B(n504), .ZN(n502) );
  XNOR2_X1 U510 ( .A(n505), .B(n506), .ZN(Result_mul_12_) );
  XNOR2_X1 U511 ( .A(n507), .B(n508), .ZN(n506) );
  XOR2_X1 U512 ( .A(n509), .B(n510), .Z(Result_mul_11_) );
  XOR2_X1 U513 ( .A(n511), .B(n512), .Z(n509) );
  NOR2_X1 U514 ( .A1(n513), .A2(n466), .ZN(n512) );
  XOR2_X1 U515 ( .A(n514), .B(n515), .Z(Result_mul_10_) );
  XNOR2_X1 U516 ( .A(n516), .B(n517), .ZN(n515) );
  NAND2_X1 U517 ( .A1(n518), .A2(n519), .ZN(Result_mul_0_) );
  NAND2_X1 U518 ( .A1(a_0_), .A2(n520), .ZN(n519) );
  NOR2_X1 U519 ( .A1(n497), .A2(n521), .ZN(n518) );
  NOR2_X1 U520 ( .A1(n498), .A2(n495), .ZN(n521) );
  NAND2_X1 U521 ( .A1(n493), .A2(n494), .ZN(n495) );
  NAND2_X1 U522 ( .A1(n522), .A2(n523), .ZN(n494) );
  NAND2_X1 U523 ( .A1(n524), .A2(n525), .ZN(n523) );
  NOR2_X1 U524 ( .A1(n489), .A2(n526), .ZN(n522) );
  NOR2_X1 U525 ( .A1(n485), .A2(n527), .ZN(n526) );
  NAND2_X1 U526 ( .A1(n492), .A2(n484), .ZN(n527) );
  NAND2_X1 U527 ( .A1(n528), .A2(n529), .ZN(n484) );
  NAND2_X1 U528 ( .A1(n474), .A2(n530), .ZN(n529) );
  INV_X1 U529 ( .A(n481), .ZN(n530) );
  INV_X1 U530 ( .A(n531), .ZN(n474) );
  NAND2_X1 U531 ( .A1(n476), .A2(n477), .ZN(n531) );
  XOR2_X1 U532 ( .A(n532), .B(n533), .Z(n477) );
  NOR2_X1 U533 ( .A1(n534), .A2(n473), .ZN(n476) );
  XNOR2_X1 U534 ( .A(n535), .B(n536), .ZN(n473) );
  XNOR2_X1 U535 ( .A(n537), .B(n538), .ZN(n536) );
  INV_X1 U536 ( .A(n472), .ZN(n534) );
  NAND2_X1 U537 ( .A1(n470), .A2(n539), .ZN(n472) );
  NAND2_X1 U538 ( .A1(n469), .A2(n471), .ZN(n539) );
  NAND2_X1 U539 ( .A1(n540), .A2(n541), .ZN(n471) );
  NAND2_X1 U540 ( .A1(a_0_), .A2(b_7_), .ZN(n541) );
  INV_X1 U541 ( .A(n542), .ZN(n540) );
  XOR2_X1 U542 ( .A(n543), .B(n544), .Z(n469) );
  XOR2_X1 U543 ( .A(n545), .B(n546), .Z(n543) );
  NOR2_X1 U544 ( .A1(n547), .A2(n467), .ZN(n546) );
  NAND2_X1 U545 ( .A1(a_0_), .A2(n542), .ZN(n470) );
  NAND2_X1 U546 ( .A1(n548), .A2(n549), .ZN(n542) );
  NAND2_X1 U547 ( .A1(n550), .A2(a_1_), .ZN(n549) );
  NOR2_X1 U548 ( .A1(n551), .A2(n466), .ZN(n550) );
  NOR2_X1 U549 ( .A1(n464), .A2(n463), .ZN(n551) );
  NAND2_X1 U550 ( .A1(n463), .A2(n464), .ZN(n548) );
  NOR2_X1 U551 ( .A1(n552), .A2(n553), .ZN(n464) );
  INV_X1 U552 ( .A(n554), .ZN(n553) );
  NAND2_X1 U553 ( .A1(n514), .A2(n555), .ZN(n554) );
  NAND2_X1 U554 ( .A1(n517), .A2(n516), .ZN(n555) );
  XNOR2_X1 U555 ( .A(n556), .B(n557), .ZN(n514) );
  XOR2_X1 U556 ( .A(n558), .B(n559), .Z(n556) );
  NOR2_X1 U557 ( .A1(n516), .A2(n517), .ZN(n552) );
  NOR2_X1 U558 ( .A1(n466), .A2(n560), .ZN(n517) );
  NAND2_X1 U559 ( .A1(n561), .A2(n562), .ZN(n516) );
  NAND2_X1 U560 ( .A1(n563), .A2(b_7_), .ZN(n562) );
  NOR2_X1 U561 ( .A1(n564), .A2(n513), .ZN(n563) );
  NOR2_X1 U562 ( .A1(n510), .A2(n511), .ZN(n564) );
  NAND2_X1 U563 ( .A1(n510), .A2(n511), .ZN(n561) );
  NAND2_X1 U564 ( .A1(n565), .A2(n566), .ZN(n511) );
  NAND2_X1 U565 ( .A1(n508), .A2(n567), .ZN(n566) );
  INV_X1 U566 ( .A(n568), .ZN(n567) );
  NOR2_X1 U567 ( .A1(n507), .A2(n505), .ZN(n568) );
  NOR2_X1 U568 ( .A1(n466), .A2(n569), .ZN(n508) );
  NAND2_X1 U569 ( .A1(n505), .A2(n507), .ZN(n565) );
  NAND2_X1 U570 ( .A1(n570), .A2(n571), .ZN(n507) );
  INV_X1 U571 ( .A(n572), .ZN(n571) );
  NOR2_X1 U572 ( .A1(n503), .A2(n573), .ZN(n572) );
  NOR2_X1 U573 ( .A1(n501), .A2(n504), .ZN(n573) );
  NAND2_X1 U574 ( .A1(n504), .A2(n501), .ZN(n570) );
  XOR2_X1 U575 ( .A(n574), .B(n575), .Z(n501) );
  NOR2_X1 U576 ( .A1(n576), .A2(n577), .ZN(n575) );
  NOR2_X1 U577 ( .A1(n466), .A2(n578), .ZN(n504) );
  XNOR2_X1 U578 ( .A(n579), .B(n580), .ZN(n505) );
  XOR2_X1 U579 ( .A(n581), .B(n582), .Z(n579) );
  XNOR2_X1 U580 ( .A(n583), .B(n584), .ZN(n510) );
  XNOR2_X1 U581 ( .A(n585), .B(n586), .ZN(n583) );
  XOR2_X1 U582 ( .A(n587), .B(n588), .Z(n463) );
  XOR2_X1 U583 ( .A(n589), .B(n590), .Z(n587) );
  NOR2_X1 U584 ( .A1(n483), .A2(n591), .ZN(n528) );
  NOR2_X1 U585 ( .A1(n592), .A2(n593), .ZN(n591) );
  NOR2_X1 U586 ( .A1(n482), .A2(n481), .ZN(n483) );
  XNOR2_X1 U587 ( .A(n593), .B(n592), .ZN(n481) );
  XNOR2_X1 U588 ( .A(n594), .B(n595), .ZN(n592) );
  XOR2_X1 U589 ( .A(n596), .B(n597), .Z(n594) );
  NAND2_X1 U590 ( .A1(n598), .A2(n599), .ZN(n593) );
  NAND2_X1 U591 ( .A1(n600), .A2(n601), .ZN(n599) );
  NAND2_X1 U592 ( .A1(n602), .A2(n603), .ZN(n601) );
  INV_X1 U593 ( .A(n604), .ZN(n598) );
  NOR2_X1 U594 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U595 ( .A1(n532), .A2(n533), .ZN(n482) );
  XOR2_X1 U596 ( .A(n600), .B(n605), .Z(n533) );
  XNOR2_X1 U597 ( .A(n603), .B(n602), .ZN(n605) );
  NOR2_X1 U598 ( .A1(n606), .A2(n577), .ZN(n602) );
  NAND2_X1 U599 ( .A1(n607), .A2(n608), .ZN(n603) );
  NAND2_X1 U600 ( .A1(n609), .A2(a_1_), .ZN(n608) );
  NOR2_X1 U601 ( .A1(n610), .A2(n577), .ZN(n609) );
  NOR2_X1 U602 ( .A1(n611), .A2(n612), .ZN(n610) );
  NAND2_X1 U603 ( .A1(n612), .A2(n611), .ZN(n607) );
  XOR2_X1 U604 ( .A(n613), .B(n614), .Z(n600) );
  XNOR2_X1 U605 ( .A(n615), .B(n616), .ZN(n614) );
  NOR2_X1 U606 ( .A1(n617), .A2(n618), .ZN(n532) );
  INV_X1 U607 ( .A(n619), .ZN(n618) );
  NAND2_X1 U608 ( .A1(n535), .A2(n620), .ZN(n619) );
  NAND2_X1 U609 ( .A1(n538), .A2(n537), .ZN(n620) );
  XNOR2_X1 U610 ( .A(n621), .B(n612), .ZN(n535) );
  XNOR2_X1 U611 ( .A(n622), .B(n623), .ZN(n612) );
  XNOR2_X1 U612 ( .A(n624), .B(n625), .ZN(n623) );
  XOR2_X1 U613 ( .A(n611), .B(n626), .Z(n621) );
  NOR2_X1 U614 ( .A1(n577), .A2(n467), .ZN(n626) );
  NAND2_X1 U615 ( .A1(n627), .A2(n628), .ZN(n611) );
  NAND2_X1 U616 ( .A1(n629), .A2(a_2_), .ZN(n628) );
  NOR2_X1 U617 ( .A1(n630), .A2(n577), .ZN(n629) );
  NOR2_X1 U618 ( .A1(n631), .A2(n632), .ZN(n630) );
  NAND2_X1 U619 ( .A1(n631), .A2(n632), .ZN(n627) );
  NOR2_X1 U620 ( .A1(n537), .A2(n538), .ZN(n617) );
  NOR2_X1 U621 ( .A1(n606), .A2(n547), .ZN(n538) );
  NAND2_X1 U622 ( .A1(n633), .A2(n634), .ZN(n537) );
  NAND2_X1 U623 ( .A1(n635), .A2(a_1_), .ZN(n634) );
  NOR2_X1 U624 ( .A1(n636), .A2(n547), .ZN(n635) );
  NOR2_X1 U625 ( .A1(n545), .A2(n544), .ZN(n636) );
  NAND2_X1 U626 ( .A1(n544), .A2(n545), .ZN(n633) );
  NAND2_X1 U627 ( .A1(n637), .A2(n638), .ZN(n545) );
  NAND2_X1 U628 ( .A1(n590), .A2(n639), .ZN(n638) );
  INV_X1 U629 ( .A(n640), .ZN(n639) );
  NOR2_X1 U630 ( .A1(n588), .A2(n589), .ZN(n640) );
  NOR2_X1 U631 ( .A1(n560), .A2(n547), .ZN(n590) );
  NAND2_X1 U632 ( .A1(n588), .A2(n589), .ZN(n637) );
  NAND2_X1 U633 ( .A1(n641), .A2(n642), .ZN(n589) );
  NAND2_X1 U634 ( .A1(n559), .A2(n643), .ZN(n642) );
  INV_X1 U635 ( .A(n644), .ZN(n643) );
  NOR2_X1 U636 ( .A1(n558), .A2(n557), .ZN(n644) );
  NOR2_X1 U637 ( .A1(n547), .A2(n513), .ZN(n559) );
  NAND2_X1 U638 ( .A1(n557), .A2(n558), .ZN(n641) );
  NAND2_X1 U639 ( .A1(n645), .A2(n646), .ZN(n558) );
  NAND2_X1 U640 ( .A1(n586), .A2(n647), .ZN(n646) );
  INV_X1 U641 ( .A(n648), .ZN(n647) );
  NOR2_X1 U642 ( .A1(n584), .A2(n585), .ZN(n648) );
  NOR2_X1 U643 ( .A1(n547), .A2(n569), .ZN(n586) );
  NAND2_X1 U644 ( .A1(n585), .A2(n584), .ZN(n645) );
  XNOR2_X1 U645 ( .A(n649), .B(n650), .ZN(n584) );
  XOR2_X1 U646 ( .A(n651), .B(n652), .Z(n650) );
  NOR2_X1 U647 ( .A1(n653), .A2(n654), .ZN(n585) );
  INV_X1 U648 ( .A(n655), .ZN(n654) );
  NAND2_X1 U649 ( .A1(n656), .A2(n582), .ZN(n655) );
  NAND2_X1 U650 ( .A1(n499), .A2(n657), .ZN(n582) );
  NOR2_X1 U651 ( .A1(n547), .A2(n576), .ZN(n499) );
  NAND2_X1 U652 ( .A1(n581), .A2(n580), .ZN(n656) );
  NOR2_X1 U653 ( .A1(n580), .A2(n581), .ZN(n653) );
  NOR2_X1 U654 ( .A1(n547), .A2(n578), .ZN(n581) );
  XOR2_X1 U655 ( .A(n657), .B(n658), .Z(n580) );
  XNOR2_X1 U656 ( .A(n659), .B(n660), .ZN(n557) );
  NAND2_X1 U657 ( .A1(n661), .A2(n662), .ZN(n659) );
  XNOR2_X1 U658 ( .A(n663), .B(n664), .ZN(n588) );
  XOR2_X1 U659 ( .A(n665), .B(n666), .Z(n664) );
  NAND2_X1 U660 ( .A1(a_3_), .A2(b_5_), .ZN(n666) );
  XNOR2_X1 U661 ( .A(n631), .B(n667), .ZN(n544) );
  XOR2_X1 U662 ( .A(n632), .B(n668), .Z(n667) );
  NAND2_X1 U663 ( .A1(a_2_), .A2(b_5_), .ZN(n668) );
  NAND2_X1 U664 ( .A1(n669), .A2(n670), .ZN(n632) );
  NAND2_X1 U665 ( .A1(n671), .A2(a_3_), .ZN(n670) );
  NOR2_X1 U666 ( .A1(n672), .A2(n577), .ZN(n671) );
  NOR2_X1 U667 ( .A1(n663), .A2(n665), .ZN(n672) );
  NAND2_X1 U668 ( .A1(n663), .A2(n665), .ZN(n669) );
  NAND2_X1 U669 ( .A1(n661), .A2(n673), .ZN(n665) );
  NAND2_X1 U670 ( .A1(n660), .A2(n662), .ZN(n673) );
  NAND2_X1 U671 ( .A1(n674), .A2(n675), .ZN(n662) );
  NAND2_X1 U672 ( .A1(b_5_), .A2(a_4_), .ZN(n675) );
  XOR2_X1 U673 ( .A(n676), .B(n677), .Z(n660) );
  XNOR2_X1 U674 ( .A(n678), .B(n679), .ZN(n677) );
  INV_X1 U675 ( .A(n680), .ZN(n661) );
  NOR2_X1 U676 ( .A1(n674), .A2(n569), .ZN(n680) );
  NAND2_X1 U677 ( .A1(n681), .A2(n682), .ZN(n674) );
  NAND2_X1 U678 ( .A1(n683), .A2(n651), .ZN(n682) );
  NAND2_X1 U679 ( .A1(n657), .A2(n658), .ZN(n651) );
  NOR2_X1 U680 ( .A1(n684), .A2(n576), .ZN(n658) );
  NOR2_X1 U681 ( .A1(n577), .A2(n685), .ZN(n657) );
  INV_X1 U682 ( .A(n686), .ZN(n683) );
  NOR2_X1 U683 ( .A1(n652), .A2(n649), .ZN(n686) );
  NAND2_X1 U684 ( .A1(n649), .A2(n652), .ZN(n681) );
  NAND2_X1 U685 ( .A1(n687), .A2(n688), .ZN(n652) );
  NAND2_X1 U686 ( .A1(n689), .A2(n690), .ZN(n688) );
  XNOR2_X1 U687 ( .A(n691), .B(n692), .ZN(n663) );
  XNOR2_X1 U688 ( .A(n693), .B(n694), .ZN(n691) );
  XNOR2_X1 U689 ( .A(n695), .B(n696), .ZN(n631) );
  XNOR2_X1 U690 ( .A(n697), .B(n698), .ZN(n695) );
  XNOR2_X1 U691 ( .A(n699), .B(n700), .ZN(n485) );
  INV_X1 U692 ( .A(n701), .ZN(n489) );
  NAND2_X1 U693 ( .A1(n491), .A2(n492), .ZN(n701) );
  XOR2_X1 U694 ( .A(n525), .B(n524), .Z(n492) );
  XNOR2_X1 U695 ( .A(n702), .B(n703), .ZN(n524) );
  XNOR2_X1 U696 ( .A(n704), .B(n705), .ZN(n703) );
  NAND2_X1 U697 ( .A1(n706), .A2(n707), .ZN(n525) );
  INV_X1 U698 ( .A(n708), .ZN(n707) );
  NOR2_X1 U699 ( .A1(n709), .A2(n710), .ZN(n708) );
  NOR2_X1 U700 ( .A1(n711), .A2(n712), .ZN(n710) );
  NAND2_X1 U701 ( .A1(n712), .A2(n711), .ZN(n706) );
  NOR2_X1 U702 ( .A1(n699), .A2(n700), .ZN(n491) );
  XNOR2_X1 U703 ( .A(n713), .B(n714), .ZN(n700) );
  INV_X1 U704 ( .A(n709), .ZN(n714) );
  XOR2_X1 U705 ( .A(n715), .B(n716), .Z(n709) );
  XNOR2_X1 U706 ( .A(n717), .B(n718), .ZN(n715) );
  XOR2_X1 U707 ( .A(n712), .B(n711), .Z(n713) );
  NAND2_X1 U708 ( .A1(n719), .A2(n720), .ZN(n711) );
  NAND2_X1 U709 ( .A1(n721), .A2(n722), .ZN(n720) );
  INV_X1 U710 ( .A(n723), .ZN(n722) );
  NOR2_X1 U711 ( .A1(n724), .A2(n725), .ZN(n723) );
  NAND2_X1 U712 ( .A1(n725), .A2(n724), .ZN(n719) );
  NOR2_X1 U713 ( .A1(n606), .A2(n726), .ZN(n712) );
  INV_X1 U714 ( .A(n727), .ZN(n699) );
  NAND2_X1 U715 ( .A1(n728), .A2(n729), .ZN(n727) );
  NAND2_X1 U716 ( .A1(n597), .A2(n730), .ZN(n729) );
  INV_X1 U717 ( .A(n731), .ZN(n730) );
  NOR2_X1 U718 ( .A1(n595), .A2(n596), .ZN(n731) );
  NOR2_X1 U719 ( .A1(n606), .A2(n684), .ZN(n597) );
  NAND2_X1 U720 ( .A1(n595), .A2(n596), .ZN(n728) );
  NAND2_X1 U721 ( .A1(n732), .A2(n733), .ZN(n596) );
  NAND2_X1 U722 ( .A1(n616), .A2(n734), .ZN(n733) );
  INV_X1 U723 ( .A(n735), .ZN(n734) );
  NOR2_X1 U724 ( .A1(n613), .A2(n615), .ZN(n735) );
  NOR2_X1 U725 ( .A1(n467), .A2(n684), .ZN(n616) );
  NAND2_X1 U726 ( .A1(n613), .A2(n615), .ZN(n732) );
  NAND2_X1 U727 ( .A1(n736), .A2(n737), .ZN(n615) );
  NAND2_X1 U728 ( .A1(n625), .A2(n738), .ZN(n737) );
  INV_X1 U729 ( .A(n739), .ZN(n738) );
  NOR2_X1 U730 ( .A1(n624), .A2(n622), .ZN(n739) );
  NOR2_X1 U731 ( .A1(n560), .A2(n684), .ZN(n625) );
  NAND2_X1 U732 ( .A1(n622), .A2(n624), .ZN(n736) );
  NAND2_X1 U733 ( .A1(n740), .A2(n741), .ZN(n624) );
  NAND2_X1 U734 ( .A1(n698), .A2(n742), .ZN(n741) );
  INV_X1 U735 ( .A(n743), .ZN(n742) );
  NOR2_X1 U736 ( .A1(n696), .A2(n697), .ZN(n743) );
  NOR2_X1 U737 ( .A1(n513), .A2(n684), .ZN(n698) );
  NAND2_X1 U738 ( .A1(n696), .A2(n697), .ZN(n740) );
  NOR2_X1 U739 ( .A1(n744), .A2(n745), .ZN(n697) );
  NOR2_X1 U740 ( .A1(n746), .A2(n694), .ZN(n745) );
  NOR2_X1 U741 ( .A1(n692), .A2(n693), .ZN(n746) );
  INV_X1 U742 ( .A(n747), .ZN(n744) );
  NAND2_X1 U743 ( .A1(n692), .A2(n693), .ZN(n747) );
  NOR2_X1 U744 ( .A1(n748), .A2(n749), .ZN(n693) );
  INV_X1 U745 ( .A(n750), .ZN(n749) );
  NAND2_X1 U746 ( .A1(n676), .A2(n751), .ZN(n750) );
  NAND2_X1 U747 ( .A1(n679), .A2(n687), .ZN(n751) );
  NOR2_X1 U748 ( .A1(n684), .A2(n578), .ZN(n676) );
  NOR2_X1 U749 ( .A1(n687), .A2(n679), .ZN(n748) );
  NAND2_X1 U750 ( .A1(n752), .A2(n753), .ZN(n679) );
  NAND2_X1 U751 ( .A1(n754), .A2(n755), .ZN(n753) );
  INV_X1 U752 ( .A(n756), .ZN(n752) );
  INV_X1 U753 ( .A(n678), .ZN(n687) );
  NOR2_X1 U754 ( .A1(n690), .A2(n689), .ZN(n678) );
  NAND2_X1 U755 ( .A1(b_4_), .A2(a_6_), .ZN(n689) );
  NAND2_X1 U756 ( .A1(a_7_), .A2(b_3_), .ZN(n690) );
  XOR2_X1 U757 ( .A(n757), .B(n758), .Z(n692) );
  XNOR2_X1 U758 ( .A(n759), .B(n756), .ZN(n758) );
  XOR2_X1 U759 ( .A(n760), .B(n761), .Z(n696) );
  XOR2_X1 U760 ( .A(n762), .B(n763), .Z(n760) );
  XNOR2_X1 U761 ( .A(n764), .B(n765), .ZN(n622) );
  XNOR2_X1 U762 ( .A(n766), .B(n767), .ZN(n764) );
  XNOR2_X1 U763 ( .A(n768), .B(n769), .ZN(n613) );
  XNOR2_X1 U764 ( .A(n770), .B(n771), .ZN(n768) );
  XNOR2_X1 U765 ( .A(n721), .B(n772), .ZN(n595) );
  XNOR2_X1 U766 ( .A(n724), .B(n725), .ZN(n772) );
  NOR2_X1 U767 ( .A1(n467), .A2(n726), .ZN(n725) );
  NAND2_X1 U768 ( .A1(n773), .A2(n774), .ZN(n724) );
  NAND2_X1 U769 ( .A1(n769), .A2(n775), .ZN(n774) );
  INV_X1 U770 ( .A(n776), .ZN(n775) );
  NOR2_X1 U771 ( .A1(n771), .A2(n770), .ZN(n776) );
  XNOR2_X1 U772 ( .A(n777), .B(n778), .ZN(n769) );
  XOR2_X1 U773 ( .A(n779), .B(n780), .Z(n778) );
  NAND2_X1 U774 ( .A1(n771), .A2(n770), .ZN(n773) );
  NOR2_X1 U775 ( .A1(n781), .A2(n782), .ZN(n770) );
  NOR2_X1 U776 ( .A1(n783), .A2(n767), .ZN(n782) );
  NOR2_X1 U777 ( .A1(n765), .A2(n766), .ZN(n783) );
  INV_X1 U778 ( .A(n784), .ZN(n781) );
  NAND2_X1 U779 ( .A1(n765), .A2(n766), .ZN(n784) );
  NOR2_X1 U780 ( .A1(n785), .A2(n786), .ZN(n766) );
  INV_X1 U781 ( .A(n787), .ZN(n786) );
  NAND2_X1 U782 ( .A1(n761), .A2(n788), .ZN(n787) );
  NAND2_X1 U783 ( .A1(n762), .A2(n763), .ZN(n788) );
  XNOR2_X1 U784 ( .A(n789), .B(n790), .ZN(n761) );
  NAND2_X1 U785 ( .A1(n791), .A2(n792), .ZN(n789) );
  NOR2_X1 U786 ( .A1(n763), .A2(n762), .ZN(n785) );
  NOR2_X1 U787 ( .A1(n793), .A2(n794), .ZN(n762) );
  INV_X1 U788 ( .A(n795), .ZN(n794) );
  NAND2_X1 U789 ( .A1(n756), .A2(n796), .ZN(n795) );
  NAND2_X1 U790 ( .A1(n759), .A2(n757), .ZN(n796) );
  NOR2_X1 U791 ( .A1(n754), .A2(n755), .ZN(n756) );
  NAND2_X1 U792 ( .A1(a_6_), .A2(b_3_), .ZN(n754) );
  NOR2_X1 U793 ( .A1(n757), .A2(n759), .ZN(n793) );
  NAND2_X1 U794 ( .A1(n797), .A2(n798), .ZN(n759) );
  NAND2_X1 U795 ( .A1(n799), .A2(n800), .ZN(n798) );
  NAND2_X1 U796 ( .A1(b_2_), .A2(a_6_), .ZN(n799) );
  NAND2_X1 U797 ( .A1(b_3_), .A2(a_5_), .ZN(n757) );
  NAND2_X1 U798 ( .A1(a_4_), .A2(b_3_), .ZN(n763) );
  XOR2_X1 U799 ( .A(n801), .B(n802), .Z(n765) );
  NAND2_X1 U800 ( .A1(n803), .A2(n804), .ZN(n801) );
  NOR2_X1 U801 ( .A1(n560), .A2(n726), .ZN(n771) );
  XNOR2_X1 U802 ( .A(n805), .B(n806), .ZN(n721) );
  XNOR2_X1 U803 ( .A(n807), .B(n808), .ZN(n806) );
  XOR2_X1 U804 ( .A(n809), .B(n810), .Z(n493) );
  INV_X1 U805 ( .A(n811), .ZN(n498) );
  NAND2_X1 U806 ( .A1(n812), .A2(n813), .ZN(n811) );
  XNOR2_X1 U807 ( .A(n814), .B(n520), .ZN(n812) );
  NOR2_X1 U808 ( .A1(n815), .A2(n813), .ZN(n497) );
  NAND2_X1 U809 ( .A1(n810), .A2(n809), .ZN(n813) );
  NAND2_X1 U810 ( .A1(n816), .A2(n817), .ZN(n809) );
  NAND2_X1 U811 ( .A1(n705), .A2(n818), .ZN(n817) );
  INV_X1 U812 ( .A(n819), .ZN(n818) );
  NOR2_X1 U813 ( .A1(n702), .A2(n704), .ZN(n819) );
  NOR2_X1 U814 ( .A1(n606), .A2(n820), .ZN(n705) );
  NAND2_X1 U815 ( .A1(n702), .A2(n704), .ZN(n816) );
  NAND2_X1 U816 ( .A1(n821), .A2(n822), .ZN(n704) );
  NAND2_X1 U817 ( .A1(n718), .A2(n823), .ZN(n822) );
  INV_X1 U818 ( .A(n824), .ZN(n823) );
  NOR2_X1 U819 ( .A1(n716), .A2(n717), .ZN(n824) );
  NOR2_X1 U820 ( .A1(n467), .A2(n820), .ZN(n718) );
  NAND2_X1 U821 ( .A1(n716), .A2(n717), .ZN(n821) );
  NOR2_X1 U822 ( .A1(n825), .A2(n826), .ZN(n717) );
  NOR2_X1 U823 ( .A1(n827), .A2(n807), .ZN(n826) );
  NOR2_X1 U824 ( .A1(n805), .A2(n808), .ZN(n827) );
  INV_X1 U825 ( .A(n828), .ZN(n825) );
  NAND2_X1 U826 ( .A1(n805), .A2(n808), .ZN(n828) );
  NAND2_X1 U827 ( .A1(n829), .A2(n830), .ZN(n808) );
  NAND2_X1 U828 ( .A1(n831), .A2(n779), .ZN(n830) );
  NAND2_X1 U829 ( .A1(a_3_), .A2(b_2_), .ZN(n779) );
  NAND2_X1 U830 ( .A1(n777), .A2(n780), .ZN(n831) );
  INV_X1 U831 ( .A(n832), .ZN(n829) );
  NOR2_X1 U832 ( .A1(n780), .A2(n777), .ZN(n832) );
  XOR2_X1 U833 ( .A(n833), .B(n834), .Z(n777) );
  XOR2_X1 U834 ( .A(n835), .B(n836), .Z(n833) );
  NAND2_X1 U835 ( .A1(n803), .A2(n837), .ZN(n780) );
  NAND2_X1 U836 ( .A1(n802), .A2(n804), .ZN(n837) );
  NAND2_X1 U837 ( .A1(n838), .A2(n839), .ZN(n804) );
  NAND2_X1 U838 ( .A1(a_4_), .A2(b_2_), .ZN(n839) );
  INV_X1 U839 ( .A(n840), .ZN(n838) );
  XNOR2_X1 U840 ( .A(n841), .B(n842), .ZN(n802) );
  NOR2_X1 U841 ( .A1(n843), .A2(n844), .ZN(n842) );
  NAND2_X1 U842 ( .A1(a_4_), .A2(n840), .ZN(n803) );
  NAND2_X1 U843 ( .A1(n791), .A2(n845), .ZN(n840) );
  NAND2_X1 U844 ( .A1(n790), .A2(n792), .ZN(n845) );
  NAND2_X1 U845 ( .A1(n797), .A2(n846), .ZN(n792) );
  NAND2_X1 U846 ( .A1(b_2_), .A2(a_5_), .ZN(n846) );
  INV_X1 U847 ( .A(n847), .ZN(n797) );
  XOR2_X1 U848 ( .A(n848), .B(n849), .Z(n790) );
  NAND2_X1 U849 ( .A1(a_7_), .A2(b_0_), .ZN(n849) );
  NAND2_X1 U850 ( .A1(n847), .A2(a_5_), .ZN(n791) );
  NOR2_X1 U851 ( .A1(n755), .A2(n848), .ZN(n847) );
  NAND2_X1 U852 ( .A1(a_6_), .A2(b_1_), .ZN(n848) );
  NAND2_X1 U853 ( .A1(b_2_), .A2(a_7_), .ZN(n755) );
  XOR2_X1 U854 ( .A(n850), .B(n851), .Z(n805) );
  XNOR2_X1 U855 ( .A(n852), .B(n853), .ZN(n851) );
  XNOR2_X1 U856 ( .A(n854), .B(n855), .ZN(n716) );
  XOR2_X1 U857 ( .A(n856), .B(n857), .Z(n854) );
  XOR2_X1 U858 ( .A(n858), .B(n859), .Z(n702) );
  XNOR2_X1 U859 ( .A(n860), .B(n861), .ZN(n859) );
  XOR2_X1 U860 ( .A(n862), .B(n863), .Z(n810) );
  XOR2_X1 U861 ( .A(n864), .B(n865), .Z(n862) );
  NAND2_X1 U862 ( .A1(n814), .A2(n866), .ZN(n815) );
  INV_X1 U863 ( .A(n520), .ZN(n866) );
  NAND2_X1 U864 ( .A1(n867), .A2(n868), .ZN(n520) );
  NAND2_X1 U865 ( .A1(n863), .A2(n869), .ZN(n868) );
  INV_X1 U866 ( .A(n870), .ZN(n869) );
  NOR2_X1 U867 ( .A1(n864), .A2(n865), .ZN(n870) );
  NOR2_X1 U868 ( .A1(n871), .A2(n467), .ZN(n863) );
  NAND2_X1 U869 ( .A1(n865), .A2(n864), .ZN(n867) );
  NAND2_X1 U870 ( .A1(n872), .A2(n873), .ZN(n864) );
  NAND2_X1 U871 ( .A1(n858), .A2(n874), .ZN(n873) );
  NAND2_X1 U872 ( .A1(n875), .A2(n860), .ZN(n874) );
  NOR2_X1 U873 ( .A1(n871), .A2(n560), .ZN(n858) );
  INV_X1 U874 ( .A(n876), .ZN(n872) );
  NOR2_X1 U875 ( .A1(n875), .A2(n860), .ZN(n876) );
  NAND2_X1 U876 ( .A1(n877), .A2(n878), .ZN(n860) );
  NAND2_X1 U877 ( .A1(n879), .A2(n856), .ZN(n878) );
  NAND2_X1 U878 ( .A1(b_0_), .A2(a_3_), .ZN(n856) );
  INV_X1 U879 ( .A(n880), .ZN(n879) );
  NOR2_X1 U880 ( .A1(n855), .A2(n857), .ZN(n880) );
  NAND2_X1 U881 ( .A1(n857), .A2(n855), .ZN(n877) );
  NAND2_X1 U882 ( .A1(a_2_), .A2(b_1_), .ZN(n855) );
  NOR2_X1 U883 ( .A1(n881), .A2(n882), .ZN(n857) );
  INV_X1 U884 ( .A(n883), .ZN(n882) );
  NAND2_X1 U885 ( .A1(n850), .A2(n884), .ZN(n883) );
  NAND2_X1 U886 ( .A1(n852), .A2(n853), .ZN(n884) );
  NOR2_X1 U887 ( .A1(n871), .A2(n569), .ZN(n850) );
  NOR2_X1 U888 ( .A1(n853), .A2(n852), .ZN(n881) );
  NOR2_X1 U889 ( .A1(n885), .A2(n886), .ZN(n852) );
  INV_X1 U890 ( .A(n887), .ZN(n886) );
  NAND2_X1 U891 ( .A1(n834), .A2(n888), .ZN(n887) );
  NAND2_X1 U892 ( .A1(n836), .A2(n835), .ZN(n888) );
  NOR2_X1 U893 ( .A1(n871), .A2(n578), .ZN(n834) );
  NOR2_X1 U894 ( .A1(n835), .A2(n836), .ZN(n885) );
  NOR2_X1 U895 ( .A1(n889), .A2(n843), .ZN(n836) );
  NOR2_X1 U896 ( .A1(n800), .A2(n844), .ZN(n843) );
  NAND2_X1 U897 ( .A1(b_1_), .A2(a_7_), .ZN(n800) );
  NOR2_X1 U898 ( .A1(n841), .A2(n844), .ZN(n889) );
  NAND2_X1 U899 ( .A1(b_0_), .A2(a_6_), .ZN(n844) );
  NAND2_X1 U900 ( .A1(b_1_), .A2(a_5_), .ZN(n841) );
  NAND2_X1 U901 ( .A1(a_4_), .A2(b_1_), .ZN(n835) );
  NAND2_X1 U902 ( .A1(a_3_), .A2(b_1_), .ZN(n853) );
  NOR2_X1 U903 ( .A1(n606), .A2(n890), .ZN(n865) );
  XNOR2_X1 U904 ( .A(n466), .B(a_7_), .ZN(Result_add_7_) );
  NAND2_X1 U905 ( .A1(n891), .A2(n503), .ZN(Result_add_6_) );
  NAND2_X1 U906 ( .A1(n574), .A2(Result_mul_15_), .ZN(n503) );
  NOR2_X1 U907 ( .A1(n892), .A2(n893), .ZN(n891) );
  NOR2_X1 U908 ( .A1(n547), .A2(n894), .ZN(n893) );
  NAND2_X1 U909 ( .A1(n895), .A2(n685), .ZN(n894) );
  INV_X1 U910 ( .A(Result_mul_15_), .ZN(n895) );
  NOR2_X1 U911 ( .A1(b_6_), .A2(n896), .ZN(n892) );
  XNOR2_X1 U912 ( .A(Result_mul_15_), .B(a_6_), .ZN(n896) );
  NAND2_X1 U913 ( .A1(n897), .A2(n898), .ZN(Result_add_5_) );
  INV_X1 U914 ( .A(n899), .ZN(n898) );
  NOR2_X1 U915 ( .A1(n649), .A2(n900), .ZN(n899) );
  NOR2_X1 U916 ( .A1(n901), .A2(n902), .ZN(n897) );
  NOR2_X1 U917 ( .A1(b_5_), .A2(n903), .ZN(n902) );
  XNOR2_X1 U918 ( .A(n578), .B(n900), .ZN(n903) );
  NOR2_X1 U919 ( .A1(n577), .A2(n904), .ZN(n901) );
  NAND2_X1 U920 ( .A1(n900), .A2(n578), .ZN(n904) );
  XNOR2_X1 U921 ( .A(n905), .B(n906), .ZN(Result_add_4_) );
  NAND2_X1 U922 ( .A1(n907), .A2(n908), .ZN(n905) );
  NAND2_X1 U923 ( .A1(n909), .A2(n910), .ZN(Result_add_3_) );
  NAND2_X1 U924 ( .A1(n767), .A2(n911), .ZN(n910) );
  NOR2_X1 U925 ( .A1(n912), .A2(n913), .ZN(n909) );
  NOR2_X1 U926 ( .A1(b_3_), .A2(n914), .ZN(n913) );
  XNOR2_X1 U927 ( .A(a_3_), .B(n911), .ZN(n914) );
  NOR2_X1 U928 ( .A1(n726), .A2(n915), .ZN(n912) );
  NAND2_X1 U929 ( .A1(n916), .A2(n513), .ZN(n915) );
  XNOR2_X1 U930 ( .A(n917), .B(n918), .ZN(Result_add_2_) );
  NOR2_X1 U931 ( .A1(n919), .A2(n807), .ZN(n918) );
  NAND2_X1 U932 ( .A1(n920), .A2(n921), .ZN(Result_add_1_) );
  NAND2_X1 U933 ( .A1(n922), .A2(n923), .ZN(n921) );
  NAND2_X1 U934 ( .A1(n875), .A2(n924), .ZN(n922) );
  INV_X1 U935 ( .A(n925), .ZN(n924) );
  INV_X1 U936 ( .A(n861), .ZN(n875) );
  NAND2_X1 U937 ( .A1(n926), .A2(n927), .ZN(n920) );
  XNOR2_X1 U938 ( .A(n890), .B(a_1_), .ZN(n926) );
  XOR2_X1 U939 ( .A(n928), .B(n929), .Z(Result_add_0_) );
  NOR2_X1 U940 ( .A1(n930), .A2(n814), .ZN(n929) );
  NOR2_X1 U941 ( .A1(n871), .A2(n606), .ZN(n814) );
  INV_X1 U942 ( .A(a_0_), .ZN(n606) );
  INV_X1 U943 ( .A(b_0_), .ZN(n871) );
  NOR2_X1 U944 ( .A1(b_0_), .A2(a_0_), .ZN(n930) );
  NOR2_X1 U945 ( .A1(n925), .A2(n931), .ZN(n928) );
  NOR2_X1 U946 ( .A1(n861), .A2(n923), .ZN(n931) );
  INV_X1 U947 ( .A(n927), .ZN(n923) );
  NOR2_X1 U948 ( .A1(n807), .A2(n932), .ZN(n927) );
  NOR2_X1 U949 ( .A1(n919), .A2(n917), .ZN(n932) );
  NOR2_X1 U950 ( .A1(n767), .A2(n933), .ZN(n917) );
  NOR2_X1 U951 ( .A1(n934), .A2(n916), .ZN(n933) );
  INV_X1 U952 ( .A(n911), .ZN(n916) );
  NAND2_X1 U953 ( .A1(n907), .A2(n935), .ZN(n911) );
  NAND2_X1 U954 ( .A1(n908), .A2(n906), .ZN(n935) );
  NAND2_X1 U955 ( .A1(n649), .A2(n936), .ZN(n906) );
  NAND2_X1 U956 ( .A1(n937), .A2(n938), .ZN(n936) );
  INV_X1 U957 ( .A(n900), .ZN(n938) );
  NOR2_X1 U958 ( .A1(n574), .A2(n939), .ZN(n900) );
  INV_X1 U959 ( .A(n940), .ZN(n939) );
  NAND2_X1 U960 ( .A1(Result_mul_15_), .A2(n941), .ZN(n940) );
  NAND2_X1 U961 ( .A1(n547), .A2(n685), .ZN(n941) );
  NOR2_X1 U962 ( .A1(n466), .A2(n576), .ZN(Result_mul_15_) );
  INV_X1 U963 ( .A(a_7_), .ZN(n576) );
  INV_X1 U964 ( .A(b_7_), .ZN(n466) );
  NOR2_X1 U965 ( .A1(n547), .A2(n685), .ZN(n574) );
  INV_X1 U966 ( .A(a_6_), .ZN(n685) );
  INV_X1 U967 ( .A(b_6_), .ZN(n547) );
  NAND2_X1 U968 ( .A1(n577), .A2(n578), .ZN(n937) );
  INV_X1 U969 ( .A(a_5_), .ZN(n578) );
  INV_X1 U970 ( .A(b_5_), .ZN(n577) );
  NAND2_X1 U971 ( .A1(b_5_), .A2(a_5_), .ZN(n649) );
  NAND2_X1 U972 ( .A1(n684), .A2(n569), .ZN(n908) );
  INV_X1 U973 ( .A(n694), .ZN(n907) );
  NOR2_X1 U974 ( .A1(n569), .A2(n684), .ZN(n694) );
  INV_X1 U975 ( .A(b_4_), .ZN(n684) );
  INV_X1 U976 ( .A(a_4_), .ZN(n569) );
  NOR2_X1 U977 ( .A1(b_3_), .A2(a_3_), .ZN(n934) );
  NOR2_X1 U978 ( .A1(n513), .A2(n726), .ZN(n767) );
  INV_X1 U979 ( .A(b_3_), .ZN(n726) );
  INV_X1 U980 ( .A(a_3_), .ZN(n513) );
  NOR2_X1 U981 ( .A1(b_2_), .A2(a_2_), .ZN(n919) );
  NOR2_X1 U982 ( .A1(n560), .A2(n820), .ZN(n807) );
  INV_X1 U983 ( .A(b_2_), .ZN(n820) );
  INV_X1 U984 ( .A(a_2_), .ZN(n560) );
  NOR2_X1 U985 ( .A1(n467), .A2(n890), .ZN(n861) );
  INV_X1 U986 ( .A(b_1_), .ZN(n890) );
  INV_X1 U987 ( .A(a_1_), .ZN(n467) );
  NOR2_X1 U988 ( .A1(b_1_), .A2(a_1_), .ZN(n925) );
endmodule

