module add_mul_mix_4_bit ( a_0_, a_1_, a_2_, a_3_, b_0_, b_1_, b_2_, b_3_, 
        c_0_, c_1_, c_2_, c_3_, d_0_, d_1_, d_2_, d_3_, Result_0_, Result_1_, 
        Result_2_, Result_3_, Result_4_, Result_5_, Result_6_, Result_7_ );
  input a_0_, a_1_, a_2_, a_3_, b_0_, b_1_, b_2_, b_3_, c_0_, c_1_, c_2_, c_3_,
         d_0_, d_1_, d_2_, d_3_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_;
  wire   n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215;

  INV_X1 U116 ( .A(n109), .ZN(Result_7_) );
  XOR2_X1 U117 ( .A(n110), .B(n111), .Z(Result_6_) );
  OR2_X1 U118 ( .A1(n112), .A2(n113), .ZN(n111) );
  OR2_X1 U119 ( .A1(n114), .A2(n115), .ZN(n110) );
  XNOR2_X1 U120 ( .A(n116), .B(n117), .ZN(Result_5_) );
  XOR2_X1 U121 ( .A(n118), .B(n119), .Z(n117) );
  XOR2_X1 U122 ( .A(n120), .B(n121), .Z(Result_4_) );
  XNOR2_X1 U123 ( .A(n122), .B(n123), .ZN(n121) );
  XOR2_X1 U124 ( .A(n124), .B(n125), .Z(Result_3_) );
  XOR2_X1 U125 ( .A(n126), .B(n127), .Z(Result_2_) );
  XOR2_X1 U126 ( .A(n128), .B(n129), .Z(Result_1_) );
  INV_X1 U127 ( .A(n130), .ZN(Result_0_) );
  AND2_X1 U128 ( .A1(n131), .A2(n132), .ZN(n130) );
  AND2_X1 U129 ( .A1(n133), .A2(n134), .ZN(n132) );
  OR2_X1 U130 ( .A1(n129), .A2(n128), .ZN(n134) );
  OR2_X1 U131 ( .A1(n135), .A2(n136), .ZN(n128) );
  INV_X1 U132 ( .A(n133), .ZN(n136) );
  AND2_X1 U133 ( .A1(n137), .A2(n138), .ZN(n135) );
  OR2_X1 U134 ( .A1(n139), .A2(n140), .ZN(n138) );
  OR2_X1 U135 ( .A1(n127), .A2(n126), .ZN(n129) );
  OR2_X1 U136 ( .A1(n125), .A2(n124), .ZN(n126) );
  OR2_X1 U137 ( .A1(n141), .A2(n142), .ZN(n124) );
  AND2_X1 U138 ( .A1(n123), .A2(n122), .ZN(n142) );
  AND2_X1 U139 ( .A1(n120), .A2(n143), .ZN(n141) );
  OR2_X1 U140 ( .A1(n122), .A2(n123), .ZN(n143) );
  OR2_X1 U141 ( .A1(n144), .A2(n112), .ZN(n123) );
  OR2_X1 U142 ( .A1(n145), .A2(n146), .ZN(n122) );
  AND2_X1 U143 ( .A1(n116), .A2(n119), .ZN(n146) );
  AND2_X1 U144 ( .A1(n147), .A2(n118), .ZN(n145) );
  OR2_X1 U145 ( .A1(n148), .A2(n149), .ZN(n118) );
  INV_X1 U146 ( .A(n150), .ZN(n149) );
  AND2_X1 U147 ( .A1(n151), .A2(n152), .ZN(n148) );
  OR2_X1 U148 ( .A1(n119), .A2(n116), .ZN(n147) );
  OR2_X1 U149 ( .A1(n152), .A2(n109), .ZN(n116) );
  OR2_X1 U150 ( .A1(n112), .A2(n114), .ZN(n109) );
  OR2_X1 U151 ( .A1(n112), .A2(n153), .ZN(n119) );
  OR2_X1 U152 ( .A1(n154), .A2(n155), .ZN(n112) );
  INV_X1 U153 ( .A(n156), .ZN(n154) );
  OR2_X1 U154 ( .A1(c_3_), .A2(d_3_), .ZN(n156) );
  XNOR2_X1 U155 ( .A(n157), .B(n158), .ZN(n120) );
  XNOR2_X1 U156 ( .A(n159), .B(n150), .ZN(n157) );
  XNOR2_X1 U157 ( .A(n160), .B(n161), .ZN(n125) );
  XNOR2_X1 U158 ( .A(n162), .B(n163), .ZN(n160) );
  XNOR2_X1 U159 ( .A(n139), .B(n140), .ZN(n127) );
  OR2_X1 U160 ( .A1(n140), .A2(n164), .ZN(n133) );
  OR2_X1 U161 ( .A1(n137), .A2(n139), .ZN(n164) );
  XOR2_X1 U162 ( .A(n165), .B(n166), .Z(n139) );
  XOR2_X1 U163 ( .A(n167), .B(n168), .Z(n165) );
  XNOR2_X1 U164 ( .A(n169), .B(n170), .ZN(n137) );
  OR2_X1 U165 ( .A1(n171), .A2(n144), .ZN(n169) );
  OR2_X1 U166 ( .A1(n172), .A2(n173), .ZN(n140) );
  AND2_X1 U167 ( .A1(n162), .A2(n163), .ZN(n173) );
  AND2_X1 U168 ( .A1(n161), .A2(n174), .ZN(n172) );
  OR2_X1 U169 ( .A1(n163), .A2(n162), .ZN(n174) );
  OR2_X1 U170 ( .A1(n175), .A2(n176), .ZN(n162) );
  AND2_X1 U171 ( .A1(n158), .A2(n150), .ZN(n176) );
  AND2_X1 U172 ( .A1(n177), .A2(n159), .ZN(n175) );
  OR2_X1 U173 ( .A1(n178), .A2(n179), .ZN(n159) );
  AND2_X1 U174 ( .A1(n180), .A2(n181), .ZN(n178) );
  OR2_X1 U175 ( .A1(n150), .A2(n158), .ZN(n177) );
  OR2_X1 U176 ( .A1(n115), .A2(n153), .ZN(n158) );
  OR2_X1 U177 ( .A1(n152), .A2(n151), .ZN(n150) );
  OR2_X1 U178 ( .A1(n114), .A2(n182), .ZN(n151) );
  OR2_X1 U179 ( .A1(n115), .A2(n113), .ZN(n152) );
  OR2_X1 U180 ( .A1(n115), .A2(n144), .ZN(n163) );
  XNOR2_X1 U181 ( .A(n155), .B(n183), .ZN(n115) );
  XOR2_X1 U182 ( .A(d_2_), .B(c_2_), .Z(n183) );
  XNOR2_X1 U183 ( .A(n184), .B(n185), .ZN(n161) );
  OR2_X1 U184 ( .A1(n179), .A2(n186), .ZN(n184) );
  INV_X1 U185 ( .A(n187), .ZN(n179) );
  OR2_X1 U186 ( .A1(n170), .A2(n144), .ZN(n131) );
  OR2_X1 U187 ( .A1(n188), .A2(n189), .ZN(n170) );
  AND2_X1 U188 ( .A1(n166), .A2(n168), .ZN(n189) );
  AND2_X1 U189 ( .A1(n167), .A2(n190), .ZN(n188) );
  OR2_X1 U190 ( .A1(n168), .A2(n166), .ZN(n190) );
  OR2_X1 U191 ( .A1(n171), .A2(n153), .ZN(n166) );
  OR2_X1 U192 ( .A1(n144), .A2(n182), .ZN(n168) );
  XOR2_X1 U193 ( .A(n191), .B(n192), .Z(n144) );
  AND2_X1 U194 ( .A1(n193), .A2(n194), .ZN(n192) );
  OR2_X1 U195 ( .A1(b_1_), .A2(n195), .ZN(n194) );
  AND2_X1 U196 ( .A1(a_1_), .A2(n196), .ZN(n195) );
  OR2_X1 U197 ( .A1(a_1_), .A2(n196), .ZN(n193) );
  XNOR2_X1 U198 ( .A(b_0_), .B(a_0_), .ZN(n191) );
  AND2_X1 U199 ( .A1(n187), .A2(n197), .ZN(n167) );
  OR2_X1 U200 ( .A1(n185), .A2(n186), .ZN(n197) );
  OR2_X1 U201 ( .A1(n113), .A2(n171), .ZN(n186) );
  OR2_X1 U202 ( .A1(n182), .A2(n153), .ZN(n185) );
  XNOR2_X1 U203 ( .A(n196), .B(n198), .ZN(n153) );
  XOR2_X1 U204 ( .A(b_1_), .B(a_1_), .Z(n198) );
  OR2_X1 U205 ( .A1(n199), .A2(n200), .ZN(n196) );
  AND2_X1 U206 ( .A1(n201), .A2(a_2_), .ZN(n200) );
  AND2_X1 U207 ( .A1(b_2_), .A2(n202), .ZN(n199) );
  OR2_X1 U208 ( .A1(n201), .A2(a_2_), .ZN(n202) );
  OR2_X1 U209 ( .A1(n180), .A2(n181), .ZN(n187) );
  OR2_X1 U210 ( .A1(n171), .A2(n114), .ZN(n181) );
  OR2_X1 U211 ( .A1(n203), .A2(n201), .ZN(n114) );
  INV_X1 U212 ( .A(n204), .ZN(n203) );
  OR2_X1 U213 ( .A1(a_3_), .A2(b_3_), .ZN(n204) );
  XOR2_X1 U214 ( .A(n205), .B(n206), .Z(n171) );
  AND2_X1 U215 ( .A1(n207), .A2(n208), .ZN(n206) );
  OR2_X1 U216 ( .A1(d_1_), .A2(n209), .ZN(n208) );
  AND2_X1 U217 ( .A1(c_1_), .A2(n210), .ZN(n209) );
  OR2_X1 U218 ( .A1(c_1_), .A2(n210), .ZN(n207) );
  XNOR2_X1 U219 ( .A(d_0_), .B(c_0_), .ZN(n205) );
  OR2_X1 U220 ( .A1(n113), .A2(n182), .ZN(n180) );
  XNOR2_X1 U221 ( .A(n210), .B(n211), .ZN(n182) );
  XOR2_X1 U222 ( .A(d_1_), .B(c_1_), .Z(n211) );
  OR2_X1 U223 ( .A1(n212), .A2(n213), .ZN(n210) );
  AND2_X1 U224 ( .A1(n155), .A2(c_2_), .ZN(n213) );
  AND2_X1 U225 ( .A1(d_2_), .A2(n214), .ZN(n212) );
  OR2_X1 U226 ( .A1(n155), .A2(c_2_), .ZN(n214) );
  AND2_X1 U227 ( .A1(c_3_), .A2(d_3_), .ZN(n155) );
  XNOR2_X1 U228 ( .A(n201), .B(n215), .ZN(n113) );
  XOR2_X1 U229 ( .A(b_2_), .B(a_2_), .Z(n215) );
  AND2_X1 U230 ( .A1(a_3_), .A2(b_3_), .ZN(n201) );
endmodule

