module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n236_, new_n976_, new_n238_, new_n479_, new_n1009_, new_n955_, new_n608_, new_n847_, new_n250_, new_n888_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n246_, new_n682_, new_n812_, new_n911_, new_n679_, new_n937_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n188_, new_n695_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n500_, new_n898_, new_n786_, new_n799_, new_n946_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n862_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n959_, new_n990_, new_n774_, new_n716_, new_n701_, new_n792_, new_n953_, new_n257_, new_n481_, new_n212_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n903_, new_n230_, new_n983_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n849_, new_n1018_, new_n855_, new_n606_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n385_, new_n829_, new_n988_, new_n478_, new_n694_, new_n461_, new_n710_, new_n971_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n683_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n966_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n961_, new_n530_, new_n890_, new_n318_, new_n1006_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n1005_, new_n999_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n956_, new_n763_, new_n960_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n970_, new_n995_, new_n271_, new_n674_, new_n274_, new_n991_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n650_, new_n708_, new_n750_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n734_, new_n912_, new_n925_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n256_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n820_, new_n771_, new_n388_, new_n979_, new_n508_, new_n714_, new_n194_, new_n483_, new_n1004_, new_n394_, new_n299_, new_n1007_, new_n935_, new_n882_, new_n657_, new_n929_, new_n652_, new_n314_, new_n582_, new_n986_, new_n1020_, new_n363_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n917_, new_n426_, new_n235_, new_n398_, new_n301_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n207_, new_n267_, new_n473_, new_n790_, new_n187_, new_n311_, new_n587_, new_n465_, new_n783_, new_n969_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n996_, new_n621_, new_n846_, new_n915_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n874_, new_n943_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n198_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n208_, new_n632_, new_n671_, new_n965_, new_n528_, new_n952_, new_n179_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n397_, new_n729_, new_n975_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n559_, new_n948_, new_n762_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n794_, new_n628_, new_n409_, new_n745_, new_n457_, new_n553_, new_n668_, new_n333_, new_n1002_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n276_, new_n688_, new_n384_, new_n900_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n1000_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n176_, new_n860_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n938_, new_n809_, new_n654_, new_n713_, new_n880_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n749_, new_n861_, new_n310_, new_n275_, new_n998_, new_n352_, new_n931_, new_n575_, new_n839_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n177_, new_n493_, new_n547_, new_n907_, new_n264_, new_n665_, new_n800_, new_n379_, new_n897_, new_n1012_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n963_, new_n270_, new_n570_, new_n598_, new_n893_, new_n993_, new_n824_, new_n520_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n557_, new_n260_, new_n936_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1016_, new_n748_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n879_, new_n513_, new_n592_, new_n726_, new_n558_, new_n231_, new_n219_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n199_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n302_, new_n191_, new_n755_, new_n225_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n977_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n972_, new_n891_, new_n631_, new_n453_, new_n516_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n252_, new_n585_, new_n751_, new_n312_, new_n535_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n190_, new_n597_, new_n978_, new_n408_, new_n470_, new_n213_, new_n769_, new_n651_, new_n433_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n992_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n815_, new_n933_, new_n304_, new_n638_, new_n523_, new_n909_, new_n857_, new_n712_, new_n1017_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n989_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n319_, new_n1008_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n957_, new_n754_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n330_, new_n727_, new_n375_, new_n962_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n357_, new_n320_, new_n780_, new_n984_, new_n245_, new_n643_, new_n474_, new_n467_, new_n1013_, new_n404_, new_n193_, new_n490_, new_n560_, new_n865_, new_n358_, new_n877_, new_n348_, new_n610_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n1011_, new_n425_, new_n175_, new_n226_, new_n896_, new_n802_, new_n697_, new_n185_, new_n951_, new_n709_, new_n373_, new_n866_, new_n540_, new_n434_, new_n200_, new_n994_, new_n982_, new_n422_, new_n964_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n551_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n521_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n181_, new_n573_, new_n765_, new_n405_;

not g000 ( new_n172_, keyIn_0_36 );
not g001 ( new_n173_, N69 );
and g002 ( new_n174_, keyIn_0_10, N63 );
or g003 ( new_n175_, keyIn_0_10, N63 );
not g004 ( new_n176_, new_n175_ );
or g005 ( new_n177_, new_n176_, new_n173_, new_n174_ );
and g006 ( new_n178_, new_n177_, keyIn_0_24 );
not g007 ( new_n179_, keyIn_0_24 );
not g008 ( new_n180_, new_n174_ );
and g009 ( new_n181_, new_n180_, new_n179_, N69, new_n175_ );
or g010 ( new_n182_, new_n178_, new_n181_ );
not g011 ( new_n183_, N95 );
not g012 ( new_n184_, N89 );
and g013 ( new_n185_, new_n184_, keyIn_0_14 );
not g014 ( new_n186_, keyIn_0_14 );
and g015 ( new_n187_, new_n186_, N89 );
or g016 ( new_n188_, new_n185_, new_n187_, new_n183_ );
and g017 ( new_n189_, new_n188_, keyIn_0_26 );
not g018 ( new_n190_, keyIn_0_26 );
not g019 ( new_n191_, new_n185_ );
not g020 ( new_n192_, new_n187_ );
and g021 ( new_n193_, new_n191_, new_n192_, new_n190_, N95 );
or g022 ( new_n194_, new_n189_, new_n193_ );
not g023 ( new_n195_, N56 );
or g024 ( new_n196_, keyIn_0_8, N50 );
and g025 ( new_n197_, keyIn_0_8, N50 );
not g026 ( new_n198_, new_n197_ );
and g027 ( new_n199_, new_n198_, new_n196_ );
or g028 ( new_n200_, new_n199_, new_n195_ );
and g029 ( new_n201_, new_n200_, keyIn_0_23 );
not g030 ( new_n202_, keyIn_0_23 );
not g031 ( new_n203_, new_n199_ );
and g032 ( new_n204_, new_n203_, new_n202_, N56 );
or g033 ( new_n205_, new_n201_, new_n204_ );
and g034 ( new_n206_, new_n205_, new_n182_, new_n194_ );
not g035 ( new_n207_, keyIn_0_22 );
not g036 ( new_n208_, N43 );
not g037 ( new_n209_, N37 );
and g038 ( new_n210_, new_n209_, keyIn_0_6 );
not g039 ( new_n211_, keyIn_0_6 );
and g040 ( new_n212_, new_n211_, N37 );
or g041 ( new_n213_, new_n210_, new_n212_, new_n208_ );
and g042 ( new_n214_, new_n213_, new_n207_ );
not g043 ( new_n215_, new_n210_ );
not g044 ( new_n216_, new_n212_ );
and g045 ( new_n217_, new_n215_, new_n216_, keyIn_0_22, N43 );
or g046 ( new_n218_, new_n214_, new_n217_ );
not g047 ( new_n219_, N30 );
or g048 ( new_n220_, keyIn_0_4, N24 );
and g049 ( new_n221_, keyIn_0_4, N24 );
not g050 ( new_n222_, new_n221_ );
and g051 ( new_n223_, new_n222_, new_n220_ );
or g052 ( new_n224_, new_n223_, new_n219_ );
and g053 ( new_n225_, new_n224_, keyIn_0_21 );
not g054 ( new_n226_, keyIn_0_21 );
not g055 ( new_n227_, new_n223_ );
and g056 ( new_n228_, new_n227_, new_n226_, N30 );
or g057 ( new_n229_, new_n225_, new_n228_ );
and g058 ( new_n230_, new_n229_, new_n218_ );
and g059 ( new_n231_, keyIn_0_0, N1 );
not g060 ( new_n232_, new_n231_ );
or g061 ( new_n233_, keyIn_0_0, N1 );
and g062 ( new_n234_, new_n232_, N4, new_n233_ );
and g063 ( new_n235_, new_n234_, keyIn_0_18 );
not g064 ( new_n236_, keyIn_0_18 );
not g065 ( new_n237_, new_n234_ );
and g066 ( new_n238_, new_n237_, new_n236_ );
or g067 ( new_n239_, new_n238_, new_n235_ );
not g068 ( new_n240_, keyIn_0_20 );
not g069 ( new_n241_, N17 );
or g070 ( new_n242_, keyIn_0_2, N11 );
and g071 ( new_n243_, keyIn_0_2, N11 );
not g072 ( new_n244_, new_n243_ );
and g073 ( new_n245_, new_n244_, new_n242_ );
or g074 ( new_n246_, new_n245_, new_n241_ );
and g075 ( new_n247_, new_n246_, new_n240_ );
not g076 ( new_n248_, new_n245_ );
and g077 ( new_n249_, new_n248_, keyIn_0_20, N17 );
or g078 ( new_n250_, new_n247_, new_n249_ );
and g079 ( new_n251_, new_n250_, new_n239_ );
not g080 ( new_n252_, keyIn_0_27 );
not g081 ( new_n253_, N108 );
or g082 ( new_n254_, keyIn_0_16, N102 );
and g083 ( new_n255_, keyIn_0_16, N102 );
not g084 ( new_n256_, new_n255_ );
and g085 ( new_n257_, new_n256_, new_n254_ );
or g086 ( new_n258_, new_n257_, new_n253_ );
and g087 ( new_n259_, new_n258_, new_n252_ );
not g088 ( new_n260_, new_n257_ );
and g089 ( new_n261_, new_n260_, keyIn_0_27, N108 );
or g090 ( new_n262_, new_n259_, new_n261_ );
and g091 ( new_n263_, keyIn_0_12, N76 );
not g092 ( new_n264_, new_n263_ );
or g093 ( new_n265_, keyIn_0_12, N76 );
and g094 ( new_n266_, new_n264_, N82, new_n265_ );
and g095 ( new_n267_, new_n266_, keyIn_0_25 );
not g096 ( new_n268_, keyIn_0_25 );
not g097 ( new_n269_, new_n266_ );
and g098 ( new_n270_, new_n269_, new_n268_ );
or g099 ( new_n271_, new_n270_, new_n267_ );
and g100 ( new_n272_, new_n262_, new_n271_ );
and g101 ( new_n273_, new_n206_, new_n230_, new_n251_, new_n272_ );
or g102 ( new_n274_, new_n273_, new_n172_ );
and g103 ( new_n275_, new_n250_, new_n262_, new_n239_, new_n271_ );
and g104 ( new_n276_, new_n275_, new_n172_, new_n206_, new_n230_ );
not g105 ( new_n277_, new_n276_ );
and g106 ( N223, new_n274_, new_n277_ );
not g107 ( new_n279_, keyIn_0_51 );
not g108 ( new_n280_, keyIn_0_30 );
not g109 ( new_n281_, N47 );
or g110 ( new_n282_, keyIn_0_7, N43 );
and g111 ( new_n283_, keyIn_0_7, N43 );
not g112 ( new_n284_, new_n283_ );
and g113 ( new_n285_, new_n284_, new_n282_ );
and g114 ( new_n286_, new_n285_, new_n281_ );
not g115 ( new_n287_, new_n286_ );
and g116 ( new_n288_, new_n287_, new_n280_ );
and g117 ( new_n289_, new_n286_, keyIn_0_30 );
or g118 ( new_n290_, new_n288_, new_n289_ );
not g119 ( new_n291_, keyIn_0_41 );
not g120 ( new_n292_, new_n218_ );
or g121 ( new_n293_, N223, keyIn_0_37 );
and g122 ( new_n294_, new_n274_, keyIn_0_37, new_n277_ );
not g123 ( new_n295_, new_n294_ );
and g124 ( new_n296_, new_n293_, new_n295_ );
and g125 ( new_n297_, new_n296_, new_n292_ );
not g126 ( new_n298_, new_n297_ );
or g127 ( new_n299_, new_n296_, new_n292_ );
and g128 ( new_n300_, new_n298_, new_n299_ );
and g129 ( new_n301_, new_n300_, new_n291_ );
not g130 ( new_n302_, new_n301_ );
or g131 ( new_n303_, new_n300_, new_n291_ );
and g132 ( new_n304_, new_n302_, new_n290_, new_n303_ );
or g133 ( new_n305_, new_n304_, new_n279_ );
and g134 ( new_n306_, new_n302_, new_n279_, new_n290_, new_n303_ );
not g135 ( new_n307_, new_n306_ );
and g136 ( new_n308_, new_n305_, new_n307_ );
not g137 ( new_n309_, keyIn_0_42 );
or g138 ( new_n310_, new_n296_, new_n205_ );
and g139 ( new_n311_, new_n293_, new_n205_, new_n295_ );
not g140 ( new_n312_, new_n311_ );
and g141 ( new_n313_, new_n310_, new_n309_, new_n312_ );
not g142 ( new_n314_, new_n313_ );
and g143 ( new_n315_, new_n310_, new_n312_ );
or g144 ( new_n316_, new_n315_, new_n309_ );
and g145 ( new_n317_, new_n316_, new_n314_ );
not g146 ( new_n318_, keyIn_0_31 );
and g147 ( new_n319_, new_n195_, keyIn_0_9 );
not g148 ( new_n320_, new_n319_ );
or g149 ( new_n321_, new_n195_, keyIn_0_9 );
and g150 ( new_n322_, new_n320_, new_n321_ );
or g151 ( new_n323_, new_n322_, N60 );
and g152 ( new_n324_, new_n323_, new_n318_ );
not g153 ( new_n325_, new_n324_ );
or g154 ( new_n326_, new_n323_, new_n318_ );
and g155 ( new_n327_, new_n325_, new_n326_ );
or g156 ( new_n328_, new_n317_, new_n327_ );
and g157 ( new_n329_, new_n328_, keyIn_0_52 );
not g158 ( new_n330_, keyIn_0_52 );
not g159 ( new_n331_, new_n317_ );
not g160 ( new_n332_, new_n327_ );
and g161 ( new_n333_, new_n331_, new_n330_, new_n332_ );
or g162 ( new_n334_, new_n329_, new_n333_ );
or g163 ( new_n335_, new_n296_, new_n229_ );
and g164 ( new_n336_, new_n296_, new_n229_ );
not g165 ( new_n337_, new_n336_ );
and g166 ( new_n338_, new_n337_, new_n335_ );
and g167 ( new_n339_, new_n338_, keyIn_0_40 );
or g168 ( new_n340_, new_n338_, keyIn_0_40 );
not g169 ( new_n341_, new_n340_ );
or g170 ( new_n342_, new_n341_, new_n339_ );
not g171 ( new_n343_, keyIn_0_29 );
and g172 ( new_n344_, new_n219_, keyIn_0_5 );
not g173 ( new_n345_, new_n344_ );
or g174 ( new_n346_, new_n219_, keyIn_0_5 );
and g175 ( new_n347_, new_n345_, new_n346_ );
not g176 ( new_n348_, new_n347_ );
or g177 ( new_n349_, new_n348_, N34 );
not g178 ( new_n350_, new_n349_ );
and g179 ( new_n351_, new_n350_, new_n343_ );
and g180 ( new_n352_, new_n349_, keyIn_0_29 );
or g181 ( new_n353_, new_n351_, new_n352_ );
not g182 ( new_n354_, new_n353_ );
and g183 ( new_n355_, new_n342_, new_n354_ );
or g184 ( new_n356_, new_n355_, keyIn_0_50 );
not g185 ( new_n357_, keyIn_0_50 );
not g186 ( new_n358_, new_n342_ );
or g187 ( new_n359_, new_n358_, new_n357_, new_n353_ );
and g188 ( new_n360_, new_n334_, new_n356_, new_n308_, new_n359_ );
or g189 ( new_n361_, new_n296_, new_n239_ );
and g190 ( new_n362_, new_n293_, new_n239_, new_n295_ );
not g191 ( new_n363_, new_n362_ );
and g192 ( new_n364_, new_n361_, keyIn_0_38, new_n363_ );
not g193 ( new_n365_, new_n364_ );
and g194 ( new_n366_, new_n361_, new_n363_ );
or g195 ( new_n367_, new_n366_, keyIn_0_38 );
and g196 ( new_n368_, new_n367_, new_n365_ );
not g197 ( new_n369_, keyIn_0_19 );
not g198 ( new_n370_, N4 );
and g199 ( new_n371_, new_n370_, keyIn_0_1 );
not g200 ( new_n372_, new_n371_ );
or g201 ( new_n373_, new_n370_, keyIn_0_1 );
and g202 ( new_n374_, new_n372_, new_n373_ );
not g203 ( new_n375_, new_n374_ );
or g204 ( new_n376_, new_n375_, N8 );
not g205 ( new_n377_, new_n376_ );
and g206 ( new_n378_, new_n377_, new_n369_ );
and g207 ( new_n379_, new_n376_, keyIn_0_19 );
or g208 ( new_n380_, new_n378_, new_n379_ );
not g209 ( new_n381_, new_n380_ );
or g210 ( new_n382_, new_n368_, new_n381_ );
and g211 ( new_n383_, new_n382_, keyIn_0_48 );
not g212 ( new_n384_, keyIn_0_48 );
not g213 ( new_n385_, new_n368_ );
and g214 ( new_n386_, new_n385_, new_n384_, new_n380_ );
or g215 ( new_n387_, new_n383_, new_n386_ );
not g216 ( new_n388_, keyIn_0_49 );
not g217 ( new_n389_, keyIn_0_28 );
or g218 ( new_n390_, keyIn_0_3, N17 );
and g219 ( new_n391_, keyIn_0_3, N17 );
not g220 ( new_n392_, new_n391_ );
and g221 ( new_n393_, new_n392_, new_n390_ );
or g222 ( new_n394_, new_n393_, N21 );
and g223 ( new_n395_, new_n394_, new_n389_ );
not g224 ( new_n396_, new_n394_ );
and g225 ( new_n397_, new_n396_, keyIn_0_28 );
or g226 ( new_n398_, new_n397_, new_n395_ );
not g227 ( new_n399_, new_n250_ );
and g228 ( new_n400_, new_n296_, new_n399_ );
not g229 ( new_n401_, new_n400_ );
or g230 ( new_n402_, new_n296_, new_n399_ );
and g231 ( new_n403_, new_n401_, new_n402_ );
or g232 ( new_n404_, new_n403_, keyIn_0_39 );
and g233 ( new_n405_, new_n401_, keyIn_0_39, new_n402_ );
not g234 ( new_n406_, new_n405_ );
and g235 ( new_n407_, new_n404_, new_n398_, new_n406_ );
not g236 ( new_n408_, new_n407_ );
and g237 ( new_n409_, new_n408_, new_n388_ );
and g238 ( new_n410_, new_n407_, keyIn_0_49 );
or g239 ( new_n411_, new_n409_, new_n410_ );
and g240 ( new_n412_, new_n387_, new_n411_ );
not g241 ( new_n413_, keyIn_0_33 );
or g242 ( new_n414_, keyIn_0_13, N82 );
and g243 ( new_n415_, keyIn_0_13, N82 );
not g244 ( new_n416_, new_n415_ );
and g245 ( new_n417_, new_n416_, new_n414_ );
or g246 ( new_n418_, new_n417_, N86 );
not g247 ( new_n419_, new_n418_ );
and g248 ( new_n420_, new_n419_, new_n413_ );
and g249 ( new_n421_, new_n418_, keyIn_0_33 );
or g250 ( new_n422_, new_n420_, new_n421_ );
not g251 ( new_n423_, keyIn_0_44 );
not g252 ( new_n424_, new_n271_ );
or g253 ( new_n425_, new_n296_, new_n424_ );
and g254 ( new_n426_, new_n293_, new_n424_, new_n295_ );
not g255 ( new_n427_, new_n426_ );
and g256 ( new_n428_, new_n425_, new_n427_ );
or g257 ( new_n429_, new_n428_, new_n423_ );
and g258 ( new_n430_, new_n425_, new_n423_, new_n427_ );
not g259 ( new_n431_, new_n430_ );
and g260 ( new_n432_, new_n429_, new_n422_, new_n431_ );
not g261 ( new_n433_, new_n432_ );
and g262 ( new_n434_, new_n433_, keyIn_0_54 );
not g263 ( new_n435_, keyIn_0_54 );
and g264 ( new_n436_, new_n432_, new_n435_ );
or g265 ( new_n437_, new_n434_, new_n436_ );
not g266 ( new_n438_, keyIn_0_46 );
or g267 ( new_n439_, new_n296_, new_n194_ );
and g268 ( new_n440_, new_n293_, new_n194_, new_n295_ );
not g269 ( new_n441_, new_n440_ );
and g270 ( new_n442_, new_n439_, new_n438_, new_n441_ );
not g271 ( new_n443_, new_n442_ );
and g272 ( new_n444_, new_n439_, new_n441_ );
or g273 ( new_n445_, new_n444_, new_n438_ );
and g274 ( new_n446_, new_n445_, new_n443_ );
not g275 ( new_n447_, keyIn_0_34 );
and g276 ( new_n448_, new_n183_, keyIn_0_15 );
not g277 ( new_n449_, new_n448_ );
or g278 ( new_n450_, new_n183_, keyIn_0_15 );
and g279 ( new_n451_, new_n449_, new_n450_ );
or g280 ( new_n452_, new_n451_, N99 );
not g281 ( new_n453_, new_n452_ );
and g282 ( new_n454_, new_n453_, new_n447_ );
and g283 ( new_n455_, new_n452_, keyIn_0_34 );
or g284 ( new_n456_, new_n454_, new_n455_ );
not g285 ( new_n457_, new_n456_ );
or g286 ( new_n458_, new_n446_, new_n457_ );
and g287 ( new_n459_, new_n458_, keyIn_0_55 );
not g288 ( new_n460_, keyIn_0_55 );
not g289 ( new_n461_, new_n446_ );
and g290 ( new_n462_, new_n461_, new_n460_, new_n456_ );
or g291 ( new_n463_, new_n459_, new_n462_ );
not g292 ( new_n464_, keyIn_0_35 );
or g293 ( new_n465_, keyIn_0_17, N108 );
and g294 ( new_n466_, keyIn_0_17, N108 );
not g295 ( new_n467_, new_n466_ );
and g296 ( new_n468_, new_n467_, new_n465_ );
or g297 ( new_n469_, new_n468_, N112 );
and g298 ( new_n470_, new_n469_, new_n464_ );
not g299 ( new_n471_, new_n469_ );
and g300 ( new_n472_, new_n471_, keyIn_0_35 );
or g301 ( new_n473_, new_n472_, new_n470_ );
not g302 ( new_n474_, keyIn_0_47 );
not g303 ( new_n475_, new_n262_ );
and g304 ( new_n476_, new_n293_, new_n475_, new_n295_ );
not g305 ( new_n477_, new_n476_ );
or g306 ( new_n478_, new_n296_, new_n475_ );
and g307 ( new_n479_, new_n478_, new_n477_ );
or g308 ( new_n480_, new_n479_, new_n474_ );
and g309 ( new_n481_, new_n478_, new_n474_, new_n477_ );
not g310 ( new_n482_, new_n481_ );
and g311 ( new_n483_, new_n480_, new_n473_, new_n482_ );
not g312 ( new_n484_, new_n483_ );
and g313 ( new_n485_, new_n484_, keyIn_0_56 );
not g314 ( new_n486_, keyIn_0_56 );
and g315 ( new_n487_, new_n483_, new_n486_ );
or g316 ( new_n488_, new_n485_, new_n487_ );
not g317 ( new_n489_, keyIn_0_53 );
not g318 ( new_n490_, keyIn_0_43 );
not g319 ( new_n491_, new_n182_ );
and g320 ( new_n492_, new_n293_, new_n491_, new_n295_ );
not g321 ( new_n493_, new_n492_ );
or g322 ( new_n494_, new_n296_, new_n491_ );
and g323 ( new_n495_, new_n494_, new_n490_, new_n493_ );
not g324 ( new_n496_, new_n495_ );
and g325 ( new_n497_, new_n494_, new_n493_ );
or g326 ( new_n498_, new_n497_, new_n490_ );
and g327 ( new_n499_, new_n498_, new_n496_ );
not g328 ( new_n500_, keyIn_0_32 );
and g329 ( new_n501_, new_n173_, keyIn_0_11 );
not g330 ( new_n502_, new_n501_ );
or g331 ( new_n503_, new_n173_, keyIn_0_11 );
and g332 ( new_n504_, new_n502_, new_n503_ );
or g333 ( new_n505_, new_n504_, N73 );
not g334 ( new_n506_, new_n505_ );
and g335 ( new_n507_, new_n506_, new_n500_ );
and g336 ( new_n508_, new_n505_, keyIn_0_32 );
or g337 ( new_n509_, new_n507_, new_n508_ );
not g338 ( new_n510_, new_n509_ );
or g339 ( new_n511_, new_n499_, new_n510_ );
and g340 ( new_n512_, new_n511_, new_n489_ );
not g341 ( new_n513_, new_n499_ );
and g342 ( new_n514_, new_n513_, keyIn_0_53, new_n509_ );
or g343 ( new_n515_, new_n512_, new_n514_ );
and g344 ( new_n516_, new_n463_, new_n515_, new_n437_, new_n488_ );
and g345 ( new_n517_, new_n516_, new_n360_, new_n412_ );
or g346 ( new_n518_, new_n517_, keyIn_0_60 );
and g347 ( new_n519_, new_n516_, new_n360_, keyIn_0_60, new_n412_ );
not g348 ( new_n520_, new_n519_ );
and g349 ( new_n521_, new_n518_, new_n520_ );
not g350 ( N329, new_n521_ );
not g351 ( new_n523_, keyIn_0_95 );
not g352 ( new_n524_, keyIn_0_93 );
not g353 ( new_n525_, keyIn_0_89 );
not g354 ( new_n526_, new_n515_ );
not g355 ( new_n527_, keyIn_0_64 );
and g356 ( new_n528_, new_n518_, new_n527_, new_n520_ );
not g357 ( new_n529_, new_n528_ );
or g358 ( new_n530_, new_n521_, new_n527_ );
and g359 ( new_n531_, new_n530_, new_n529_ );
and g360 ( new_n532_, new_n531_, new_n526_ );
not g361 ( new_n533_, new_n531_ );
and g362 ( new_n534_, new_n533_, new_n515_ );
or g363 ( new_n535_, new_n534_, new_n532_ );
and g364 ( new_n536_, new_n535_, keyIn_0_73 );
not g365 ( new_n537_, keyIn_0_73 );
not g366 ( new_n538_, new_n535_ );
and g367 ( new_n539_, new_n538_, new_n537_ );
not g368 ( new_n540_, keyIn_0_62 );
not g369 ( new_n541_, keyIn_0_58 );
or g370 ( new_n542_, new_n499_, N79, new_n504_ );
and g371 ( new_n543_, new_n542_, new_n541_ );
not g372 ( new_n544_, new_n543_ );
or g373 ( new_n545_, new_n542_, new_n541_ );
and g374 ( new_n546_, new_n544_, new_n545_ );
and g375 ( new_n547_, new_n546_, new_n540_ );
or g376 ( new_n548_, new_n546_, new_n540_ );
not g377 ( new_n549_, new_n548_ );
or g378 ( new_n550_, new_n549_, new_n547_ );
or g379 ( new_n551_, new_n539_, new_n536_, new_n525_, new_n550_ );
not g380 ( new_n552_, keyIn_0_88 );
not g381 ( new_n553_, keyIn_0_71 );
not g382 ( new_n554_, new_n334_ );
or g383 ( new_n555_, new_n531_, new_n554_ );
and g384 ( new_n556_, new_n531_, new_n554_ );
not g385 ( new_n557_, new_n556_ );
and g386 ( new_n558_, new_n557_, new_n553_, new_n555_ );
not g387 ( new_n559_, new_n558_ );
and g388 ( new_n560_, new_n557_, new_n555_ );
or g389 ( new_n561_, new_n560_, new_n553_ );
not g390 ( new_n562_, keyIn_0_57 );
or g391 ( new_n563_, new_n317_, N66, new_n322_ );
not g392 ( new_n564_, new_n563_ );
and g393 ( new_n565_, new_n564_, new_n562_ );
and g394 ( new_n566_, new_n563_, keyIn_0_57 );
or g395 ( new_n567_, new_n565_, new_n566_ );
or g396 ( new_n568_, new_n567_, keyIn_0_61 );
not g397 ( new_n569_, keyIn_0_61 );
not g398 ( new_n570_, new_n567_ );
or g399 ( new_n571_, new_n570_, new_n569_ );
and g400 ( new_n572_, new_n571_, new_n568_ );
and g401 ( new_n573_, new_n561_, new_n559_, new_n572_ );
or g402 ( new_n574_, new_n573_, new_n552_ );
and g403 ( new_n575_, new_n561_, new_n552_, new_n559_, new_n572_ );
not g404 ( new_n576_, new_n575_ );
and g405 ( new_n577_, new_n574_, new_n551_, new_n576_ );
not g406 ( new_n578_, keyIn_0_90 );
not g407 ( new_n579_, keyIn_0_75 );
not g408 ( new_n580_, new_n437_ );
and g409 ( new_n581_, new_n531_, new_n580_ );
and g410 ( new_n582_, new_n533_, new_n437_ );
or g411 ( new_n583_, new_n582_, new_n581_ );
and g412 ( new_n584_, new_n583_, new_n579_ );
not g413 ( new_n585_, new_n584_ );
not g414 ( new_n586_, new_n581_ );
not g415 ( new_n587_, new_n582_ );
and g416 ( new_n588_, new_n587_, keyIn_0_75, new_n586_ );
not g417 ( new_n589_, new_n588_ );
not g418 ( new_n590_, N92 );
not g419 ( new_n591_, new_n417_ );
and g420 ( new_n592_, new_n429_, new_n431_ );
and g421 ( new_n593_, new_n592_, new_n590_, new_n591_ );
and g422 ( new_n594_, new_n585_, new_n578_, new_n589_, new_n593_ );
not g423 ( new_n595_, new_n593_ );
or g424 ( new_n596_, new_n584_, new_n588_, new_n595_ );
and g425 ( new_n597_, new_n596_, keyIn_0_90 );
or g426 ( new_n598_, new_n597_, new_n594_ );
not g427 ( new_n599_, keyIn_0_79 );
not g428 ( new_n600_, new_n488_ );
and g429 ( new_n601_, new_n530_, new_n600_, new_n529_ );
not g430 ( new_n602_, new_n601_ );
or g431 ( new_n603_, new_n531_, new_n600_ );
and g432 ( new_n604_, new_n603_, new_n599_, new_n602_ );
not g433 ( new_n605_, new_n604_ );
and g434 ( new_n606_, new_n603_, new_n602_ );
or g435 ( new_n607_, new_n606_, new_n599_ );
and g436 ( new_n608_, new_n607_, new_n605_ );
not g437 ( new_n609_, N115 );
not g438 ( new_n610_, new_n468_ );
and g439 ( new_n611_, new_n480_, new_n482_ );
and g440 ( new_n612_, new_n611_, new_n609_, new_n610_ );
not g441 ( new_n613_, new_n612_ );
or g442 ( new_n614_, new_n608_, new_n613_ );
and g443 ( new_n615_, new_n614_, keyIn_0_92 );
not g444 ( new_n616_, keyIn_0_92 );
not g445 ( new_n617_, new_n608_ );
and g446 ( new_n618_, new_n617_, new_n616_, new_n612_ );
or g447 ( new_n619_, new_n615_, new_n618_ );
and g448 ( new_n620_, new_n619_, new_n577_, new_n598_ );
not g449 ( new_n621_, keyIn_0_91 );
not g450 ( new_n622_, keyIn_0_77 );
or g451 ( new_n623_, new_n531_, new_n463_ );
and g452 ( new_n624_, new_n530_, new_n463_, new_n529_ );
not g453 ( new_n625_, new_n624_ );
and g454 ( new_n626_, new_n623_, new_n622_, new_n625_ );
not g455 ( new_n627_, new_n626_ );
and g456 ( new_n628_, new_n623_, new_n625_ );
or g457 ( new_n629_, new_n628_, new_n622_ );
and g458 ( new_n630_, new_n629_, new_n627_ );
not g459 ( new_n631_, keyIn_0_63 );
not g460 ( new_n632_, keyIn_0_59 );
or g461 ( new_n633_, new_n446_, N105, new_n451_ );
and g462 ( new_n634_, new_n633_, new_n632_ );
not g463 ( new_n635_, new_n634_ );
or g464 ( new_n636_, new_n633_, new_n632_ );
and g465 ( new_n637_, new_n635_, new_n636_ );
and g466 ( new_n638_, new_n637_, new_n631_ );
not g467 ( new_n639_, new_n638_ );
or g468 ( new_n640_, new_n637_, new_n631_ );
and g469 ( new_n641_, new_n639_, new_n640_ );
or g470 ( new_n642_, new_n630_, new_n641_ );
and g471 ( new_n643_, new_n642_, new_n621_ );
not g472 ( new_n644_, new_n630_ );
not g473 ( new_n645_, new_n641_ );
and g474 ( new_n646_, new_n644_, keyIn_0_91, new_n645_ );
or g475 ( new_n647_, new_n643_, new_n646_ );
not g476 ( new_n648_, new_n536_ );
not g477 ( new_n649_, new_n539_ );
not g478 ( new_n650_, new_n547_ );
and g479 ( new_n651_, new_n649_, new_n648_, new_n650_, new_n548_ );
or g480 ( new_n652_, new_n651_, keyIn_0_89 );
and g481 ( new_n653_, new_n647_, new_n652_ );
not g482 ( new_n654_, keyIn_0_86 );
not g483 ( new_n655_, N40 );
and g484 ( new_n656_, new_n356_, new_n359_ );
or g485 ( new_n657_, new_n531_, new_n656_ );
and g486 ( new_n658_, new_n531_, new_n656_ );
not g487 ( new_n659_, new_n658_ );
and g488 ( new_n660_, new_n659_, keyIn_0_68, new_n657_ );
not g489 ( new_n661_, keyIn_0_68 );
not g490 ( new_n662_, new_n656_ );
and g491 ( new_n663_, new_n533_, new_n662_ );
or g492 ( new_n664_, new_n663_, new_n658_ );
and g493 ( new_n665_, new_n664_, new_n661_ );
or g494 ( new_n666_, new_n665_, new_n660_ );
and g495 ( new_n667_, new_n666_, new_n655_, new_n342_, new_n347_ );
or g496 ( new_n668_, new_n667_, new_n654_ );
or g497 ( new_n669_, new_n531_, new_n308_ );
and g498 ( new_n670_, new_n531_, new_n308_ );
not g499 ( new_n671_, new_n670_ );
and g500 ( new_n672_, new_n671_, new_n669_ );
and g501 ( new_n673_, new_n672_, keyIn_0_69 );
not g502 ( new_n674_, new_n673_ );
or g503 ( new_n675_, new_n672_, keyIn_0_69 );
not g504 ( new_n676_, N53 );
and g505 ( new_n677_, new_n302_, new_n676_, new_n285_, new_n303_ );
and g506 ( new_n678_, new_n674_, new_n675_, new_n677_ );
or g507 ( new_n679_, new_n678_, keyIn_0_87 );
and g508 ( new_n680_, new_n674_, keyIn_0_87, new_n675_, new_n677_ );
not g509 ( new_n681_, new_n680_ );
not g510 ( new_n682_, new_n660_ );
and g511 ( new_n683_, new_n659_, new_n657_ );
or g512 ( new_n684_, new_n683_, keyIn_0_68 );
and g513 ( new_n685_, new_n684_, new_n682_ );
or g514 ( new_n686_, new_n358_, N40, new_n348_ );
or g515 ( new_n687_, new_n685_, keyIn_0_86, new_n686_ );
and g516 ( new_n688_, new_n687_, new_n681_ );
and g517 ( new_n689_, new_n668_, new_n679_, new_n688_ );
not g518 ( new_n690_, keyIn_0_85 );
not g519 ( new_n691_, keyIn_0_67 );
not g520 ( new_n692_, new_n411_ );
or g521 ( new_n693_, new_n531_, new_n692_ );
and g522 ( new_n694_, new_n530_, new_n692_, new_n529_ );
not g523 ( new_n695_, new_n694_ );
and g524 ( new_n696_, new_n693_, new_n691_, new_n695_ );
not g525 ( new_n697_, new_n696_ );
and g526 ( new_n698_, new_n693_, new_n695_ );
or g527 ( new_n699_, new_n698_, new_n691_ );
not g528 ( new_n700_, N27 );
not g529 ( new_n701_, new_n393_ );
and g530 ( new_n702_, new_n404_, new_n700_, new_n701_, new_n406_ );
and g531 ( new_n703_, new_n699_, new_n697_, new_n702_ );
not g532 ( new_n704_, new_n703_ );
and g533 ( new_n705_, new_n704_, new_n690_ );
and g534 ( new_n706_, new_n703_, keyIn_0_85 );
or g535 ( new_n707_, new_n705_, new_n706_ );
not g536 ( new_n708_, keyIn_0_66 );
or g537 ( new_n709_, new_n531_, new_n387_ );
and g538 ( new_n710_, new_n530_, new_n387_, new_n529_ );
not g539 ( new_n711_, new_n710_ );
and g540 ( new_n712_, new_n709_, new_n708_, new_n711_ );
not g541 ( new_n713_, new_n712_ );
and g542 ( new_n714_, new_n709_, new_n711_ );
or g543 ( new_n715_, new_n714_, new_n708_ );
and g544 ( new_n716_, new_n715_, new_n713_ );
or g545 ( new_n717_, new_n375_, N14 );
or g546 ( new_n718_, new_n368_, new_n717_ );
or g547 ( new_n719_, new_n716_, new_n718_ );
and g548 ( new_n720_, new_n719_, keyIn_0_84 );
not g549 ( new_n721_, keyIn_0_84 );
not g550 ( new_n722_, new_n716_ );
not g551 ( new_n723_, new_n717_ );
and g552 ( new_n724_, new_n722_, new_n721_, new_n385_, new_n723_ );
or g553 ( new_n725_, new_n720_, new_n724_ );
and g554 ( new_n726_, new_n725_, new_n707_ );
and g555 ( new_n727_, new_n620_, new_n653_, new_n726_, new_n689_ );
or g556 ( new_n728_, new_n727_, new_n524_ );
and g557 ( new_n729_, new_n707_, new_n524_ );
and g558 ( new_n730_, new_n717_, keyIn_0_84 );
or g559 ( new_n731_, new_n720_, new_n724_, new_n730_ );
and g560 ( new_n732_, new_n731_, new_n647_, new_n652_ );
and g561 ( new_n733_, new_n732_, new_n620_, new_n689_, new_n729_ );
not g562 ( new_n734_, new_n733_ );
and g563 ( new_n735_, new_n728_, new_n734_ );
and g564 ( new_n736_, new_n735_, new_n523_ );
not g565 ( new_n737_, new_n735_ );
and g566 ( new_n738_, new_n737_, keyIn_0_95 );
or g567 ( N370, new_n738_, new_n736_ );
not g568 ( new_n740_, keyIn_0_115 );
and g569 ( new_n741_, new_n728_, keyIn_0_94, new_n734_ );
not g570 ( new_n742_, new_n741_ );
or g571 ( new_n743_, new_n735_, keyIn_0_94 );
and g572 ( new_n744_, new_n743_, keyIn_0_103, N105, new_n742_ );
not g573 ( new_n745_, new_n744_ );
and g574 ( new_n746_, new_n743_, N105, new_n742_ );
or g575 ( new_n747_, new_n746_, keyIn_0_103 );
not g576 ( new_n748_, keyIn_0_82 );
or g577 ( new_n749_, new_n521_, keyIn_0_65 );
and g578 ( new_n750_, new_n521_, keyIn_0_65 );
not g579 ( new_n751_, new_n750_ );
and g580 ( new_n752_, new_n751_, new_n749_ );
and g581 ( new_n753_, new_n752_, N99 );
and g582 ( new_n754_, new_n753_, new_n748_ );
not g583 ( new_n755_, new_n753_ );
and g584 ( new_n756_, new_n755_, keyIn_0_82 );
or g585 ( new_n757_, new_n756_, new_n754_ );
and g586 ( new_n758_, N223, N89 );
not g587 ( new_n759_, new_n758_ );
and g588 ( new_n760_, new_n757_, N95, new_n759_ );
and g589 ( new_n761_, new_n747_, new_n745_, new_n760_ );
or g590 ( new_n762_, new_n761_, keyIn_0_112 );
and g591 ( new_n763_, new_n747_, keyIn_0_112, new_n745_, new_n760_ );
not g592 ( new_n764_, new_n763_ );
and g593 ( new_n765_, new_n762_, new_n764_ );
not g594 ( new_n766_, new_n765_ );
and g595 ( new_n767_, new_n743_, keyIn_0_101, N79, new_n742_ );
not g596 ( new_n768_, new_n767_ );
and g597 ( new_n769_, new_n743_, N79, new_n742_ );
or g598 ( new_n770_, new_n769_, keyIn_0_101 );
not g599 ( new_n771_, keyIn_0_80 );
and g600 ( new_n772_, new_n752_, N73 );
and g601 ( new_n773_, new_n772_, new_n771_ );
not g602 ( new_n774_, new_n773_ );
or g603 ( new_n775_, new_n772_, new_n771_ );
and g604 ( new_n776_, N223, N63 );
not g605 ( new_n777_, new_n776_ );
and g606 ( new_n778_, new_n774_, N69, new_n775_, new_n777_ );
and g607 ( new_n779_, new_n770_, new_n768_, new_n778_ );
not g608 ( new_n780_, new_n779_ );
and g609 ( new_n781_, new_n780_, keyIn_0_110 );
not g610 ( new_n782_, keyIn_0_110 );
and g611 ( new_n783_, new_n779_, new_n782_ );
or g612 ( new_n784_, new_n781_, new_n783_ );
not g613 ( new_n785_, keyIn_0_113 );
not g614 ( new_n786_, keyIn_0_104 );
and g615 ( new_n787_, new_n743_, N115, new_n742_ );
and g616 ( new_n788_, new_n787_, new_n786_ );
not g617 ( new_n789_, new_n788_ );
or g618 ( new_n790_, new_n787_, new_n786_ );
and g619 ( new_n791_, new_n789_, new_n790_ );
not g620 ( new_n792_, keyIn_0_83 );
and g621 ( new_n793_, new_n752_, N112 );
and g622 ( new_n794_, new_n793_, new_n792_ );
not g623 ( new_n795_, new_n794_ );
or g624 ( new_n796_, new_n793_, new_n792_ );
and g625 ( new_n797_, N223, N102 );
not g626 ( new_n798_, new_n797_ );
and g627 ( new_n799_, new_n795_, N108, new_n796_, new_n798_ );
not g628 ( new_n800_, new_n799_ );
or g629 ( new_n801_, new_n791_, new_n800_ );
and g630 ( new_n802_, new_n801_, new_n785_ );
not g631 ( new_n803_, new_n791_ );
and g632 ( new_n804_, new_n803_, keyIn_0_113, new_n799_ );
or g633 ( new_n805_, new_n802_, new_n804_ );
not g634 ( new_n806_, keyIn_0_111 );
and g635 ( new_n807_, new_n743_, N92, new_n742_ );
or g636 ( new_n808_, new_n807_, keyIn_0_102 );
and g637 ( new_n809_, new_n743_, keyIn_0_102, N92, new_n742_ );
not g638 ( new_n810_, new_n809_ );
and g639 ( new_n811_, new_n808_, new_n810_ );
not g640 ( new_n812_, keyIn_0_81 );
and g641 ( new_n813_, new_n752_, N86 );
and g642 ( new_n814_, new_n813_, new_n812_ );
not g643 ( new_n815_, new_n814_ );
or g644 ( new_n816_, new_n813_, new_n812_ );
and g645 ( new_n817_, N223, N76 );
not g646 ( new_n818_, new_n817_ );
and g647 ( new_n819_, new_n815_, N82, new_n816_, new_n818_ );
not g648 ( new_n820_, new_n819_ );
or g649 ( new_n821_, new_n811_, new_n820_ );
and g650 ( new_n822_, new_n821_, new_n806_ );
not g651 ( new_n823_, new_n811_ );
and g652 ( new_n824_, new_n823_, keyIn_0_111, new_n819_ );
or g653 ( new_n825_, new_n822_, new_n824_ );
and g654 ( new_n826_, new_n805_, new_n766_, new_n784_, new_n825_ );
not g655 ( new_n827_, keyIn_0_108 );
not g656 ( new_n828_, keyIn_0_99 );
and g657 ( new_n829_, new_n743_, N53, new_n742_ );
or g658 ( new_n830_, new_n829_, new_n828_ );
and g659 ( new_n831_, new_n743_, new_n828_, N53, new_n742_ );
not g660 ( new_n832_, new_n831_ );
and g661 ( new_n833_, new_n830_, new_n832_ );
not g662 ( new_n834_, keyIn_0_76 );
and g663 ( new_n835_, new_n752_, N47 );
and g664 ( new_n836_, new_n835_, new_n834_ );
not g665 ( new_n837_, new_n836_ );
or g666 ( new_n838_, new_n835_, new_n834_ );
and g667 ( new_n839_, N223, N37 );
not g668 ( new_n840_, new_n839_ );
and g669 ( new_n841_, new_n837_, N43, new_n838_, new_n840_ );
not g670 ( new_n842_, new_n841_ );
or g671 ( new_n843_, new_n833_, new_n842_ );
and g672 ( new_n844_, new_n843_, new_n827_ );
not g673 ( new_n845_, new_n833_ );
and g674 ( new_n846_, new_n845_, keyIn_0_108, new_n841_ );
or g675 ( new_n847_, new_n844_, new_n846_ );
and g676 ( new_n848_, new_n743_, N66, new_n742_ );
or g677 ( new_n849_, new_n848_, keyIn_0_100 );
and g678 ( new_n850_, new_n848_, keyIn_0_100 );
not g679 ( new_n851_, new_n850_ );
and g680 ( new_n852_, new_n851_, new_n849_ );
and g681 ( new_n853_, new_n752_, N60 );
and g682 ( new_n854_, new_n853_, keyIn_0_78 );
not g683 ( new_n855_, new_n854_ );
or g684 ( new_n856_, new_n853_, keyIn_0_78 );
and g685 ( new_n857_, N223, N50 );
not g686 ( new_n858_, new_n857_ );
and g687 ( new_n859_, new_n855_, N56, new_n856_, new_n858_ );
not g688 ( new_n860_, new_n859_ );
or g689 ( new_n861_, new_n852_, new_n860_ );
and g690 ( new_n862_, new_n861_, keyIn_0_109 );
not g691 ( new_n863_, keyIn_0_109 );
not g692 ( new_n864_, new_n852_ );
and g693 ( new_n865_, new_n864_, new_n863_, new_n859_ );
or g694 ( new_n866_, new_n862_, new_n865_ );
and g695 ( new_n867_, new_n866_, new_n847_ );
not g696 ( new_n868_, keyIn_0_106 );
and g697 ( new_n869_, new_n743_, N27, new_n742_ );
or g698 ( new_n870_, new_n869_, keyIn_0_97 );
and g699 ( new_n871_, new_n869_, keyIn_0_97 );
not g700 ( new_n872_, new_n871_ );
not g701 ( new_n873_, keyIn_0_72 );
and g702 ( new_n874_, new_n752_, N21 );
and g703 ( new_n875_, new_n874_, new_n873_ );
not g704 ( new_n876_, new_n875_ );
or g705 ( new_n877_, new_n874_, new_n873_ );
and g706 ( new_n878_, N223, N11 );
and g707 ( new_n879_, new_n878_, keyIn_0_45 );
not g708 ( new_n880_, new_n879_ );
or g709 ( new_n881_, new_n878_, keyIn_0_45 );
and g710 ( new_n882_, new_n880_, N17, new_n881_ );
and g711 ( new_n883_, new_n876_, new_n877_, new_n882_ );
and g712 ( new_n884_, new_n872_, new_n870_, new_n883_ );
and g713 ( new_n885_, new_n884_, new_n868_ );
not g714 ( new_n886_, new_n884_ );
and g715 ( new_n887_, new_n886_, keyIn_0_106 );
or g716 ( new_n888_, new_n887_, new_n885_ );
not g717 ( new_n889_, keyIn_0_98 );
and g718 ( new_n890_, new_n743_, N40, new_n742_ );
or g719 ( new_n891_, new_n890_, new_n889_ );
and g720 ( new_n892_, new_n743_, new_n889_, N40, new_n742_ );
not g721 ( new_n893_, new_n892_ );
and g722 ( new_n894_, new_n891_, new_n893_ );
not g723 ( new_n895_, keyIn_0_74 );
and g724 ( new_n896_, new_n752_, N34 );
and g725 ( new_n897_, new_n896_, new_n895_ );
not g726 ( new_n898_, new_n897_ );
or g727 ( new_n899_, new_n896_, new_n895_ );
and g728 ( new_n900_, N223, N24 );
not g729 ( new_n901_, new_n900_ );
and g730 ( new_n902_, new_n898_, N30, new_n899_, new_n901_ );
not g731 ( new_n903_, new_n902_ );
or g732 ( new_n904_, new_n894_, new_n903_ );
and g733 ( new_n905_, new_n904_, keyIn_0_107 );
not g734 ( new_n906_, keyIn_0_107 );
not g735 ( new_n907_, new_n894_ );
and g736 ( new_n908_, new_n907_, new_n906_, new_n902_ );
or g737 ( new_n909_, new_n905_, new_n908_ );
and g738 ( new_n910_, new_n909_, new_n888_ );
and g739 ( new_n911_, new_n867_, new_n910_ );
and g740 ( new_n912_, new_n911_, new_n826_ );
or g741 ( new_n913_, new_n912_, new_n740_ );
not g742 ( new_n914_, new_n913_ );
not g743 ( new_n915_, keyIn_0_114 );
not g744 ( new_n916_, keyIn_0_96 );
and g745 ( new_n917_, new_n743_, N14, new_n742_ );
and g746 ( new_n918_, new_n917_, new_n916_ );
not g747 ( new_n919_, new_n918_ );
or g748 ( new_n920_, new_n917_, new_n916_ );
and g749 ( new_n921_, new_n919_, new_n920_ );
not g750 ( new_n922_, new_n921_ );
not g751 ( new_n923_, keyIn_0_70 );
and g752 ( new_n924_, new_n752_, N8 );
and g753 ( new_n925_, new_n924_, new_n923_ );
not g754 ( new_n926_, new_n925_ );
or g755 ( new_n927_, new_n924_, new_n923_ );
and g756 ( new_n928_, N223, N1 );
not g757 ( new_n929_, new_n928_ );
and g758 ( new_n930_, new_n926_, N4, new_n927_, new_n929_ );
and g759 ( new_n931_, new_n922_, new_n930_ );
or g760 ( new_n932_, new_n931_, keyIn_0_105 );
and g761 ( new_n933_, new_n931_, keyIn_0_105 );
not g762 ( new_n934_, new_n933_ );
and g763 ( new_n935_, new_n934_, new_n932_ );
and g764 ( new_n936_, new_n935_, new_n915_ );
not g765 ( new_n937_, new_n936_ );
or g766 ( new_n938_, new_n935_, new_n915_ );
and g767 ( new_n939_, new_n937_, new_n938_ );
and g768 ( new_n940_, new_n912_, new_n740_ );
or g769 ( new_n941_, new_n914_, new_n939_, new_n940_ );
and g770 ( new_n942_, new_n941_, keyIn_0_120 );
not g771 ( new_n943_, keyIn_0_120 );
not g772 ( new_n944_, new_n939_ );
not g773 ( new_n945_, new_n940_ );
and g774 ( new_n946_, new_n945_, new_n943_, new_n913_, new_n944_ );
or g775 ( N421, new_n942_, new_n946_ );
not g776 ( new_n948_, keyIn_0_125 );
not g777 ( new_n949_, keyIn_0_121 );
not g778 ( new_n950_, keyIn_0_116 );
not g779 ( new_n951_, new_n844_ );
not g780 ( new_n952_, new_n846_ );
and g781 ( new_n953_, new_n951_, new_n950_, new_n952_ );
and g782 ( new_n954_, new_n847_, keyIn_0_116 );
or g783 ( new_n955_, new_n954_, new_n953_ );
and g784 ( new_n956_, new_n955_, new_n909_ );
or g785 ( new_n957_, new_n956_, new_n949_ );
and g786 ( new_n958_, new_n955_, new_n949_, new_n909_ );
not g787 ( new_n959_, new_n958_ );
and g788 ( new_n960_, new_n957_, new_n959_ );
and g789 ( new_n961_, new_n910_, new_n866_ );
not g790 ( new_n962_, new_n961_ );
or g791 ( new_n963_, new_n960_, new_n962_ );
and g792 ( new_n964_, new_n963_, new_n948_ );
not g793 ( new_n965_, new_n960_ );
and g794 ( new_n966_, new_n965_, keyIn_0_125, new_n961_ );
or g795 ( N430, new_n964_, new_n966_ );
not g796 ( new_n968_, new_n910_ );
not g797 ( new_n969_, new_n822_ );
not g798 ( new_n970_, new_n824_ );
and g799 ( new_n971_, new_n969_, keyIn_0_118, new_n970_ );
not g800 ( new_n972_, keyIn_0_118 );
and g801 ( new_n973_, new_n825_, new_n972_ );
or g802 ( new_n974_, new_n973_, new_n971_ );
and g803 ( new_n975_, new_n974_, new_n867_ );
or g804 ( new_n976_, new_n975_, keyIn_0_123 );
and g805 ( new_n977_, new_n974_, keyIn_0_123, new_n867_ );
not g806 ( new_n978_, new_n977_ );
and g807 ( new_n979_, new_n976_, new_n978_ );
not g808 ( new_n980_, keyIn_0_122 );
not g809 ( new_n981_, keyIn_0_117 );
or g810 ( new_n982_, new_n779_, new_n782_ );
not g811 ( new_n983_, new_n783_ );
and g812 ( new_n984_, new_n983_, new_n982_ );
and g813 ( new_n985_, new_n984_, new_n981_ );
and g814 ( new_n986_, new_n784_, keyIn_0_117 );
or g815 ( new_n987_, new_n986_, new_n985_ );
and g816 ( new_n988_, new_n987_, new_n867_, new_n909_ );
or g817 ( new_n989_, new_n988_, new_n980_ );
not g818 ( new_n990_, new_n867_ );
not g819 ( new_n991_, new_n909_ );
not g820 ( new_n992_, new_n987_ );
or g821 ( new_n993_, new_n992_, new_n990_, keyIn_0_122, new_n991_ );
and g822 ( new_n994_, new_n989_, new_n993_ );
or g823 ( new_n995_, new_n979_, new_n994_, new_n968_ );
and g824 ( new_n996_, new_n995_, keyIn_0_126 );
not g825 ( new_n997_, keyIn_0_126 );
not g826 ( new_n998_, new_n979_ );
not g827 ( new_n999_, new_n994_ );
and g828 ( new_n1000_, new_n998_, new_n999_, new_n997_, new_n910_ );
or g829 ( N431, new_n996_, new_n1000_ );
not g830 ( new_n1002_, new_n825_ );
not g831 ( new_n1003_, new_n847_ );
not g832 ( new_n1004_, keyIn_0_119 );
and g833 ( new_n1005_, new_n762_, new_n1004_, new_n764_ );
not g834 ( new_n1006_, new_n1005_ );
or g835 ( new_n1007_, new_n765_, new_n1004_ );
and g836 ( new_n1008_, new_n1007_, new_n1006_ );
or g837 ( new_n1009_, new_n1008_, new_n1002_, new_n1003_, new_n991_ );
and g838 ( new_n1010_, new_n1009_, keyIn_0_124 );
not g839 ( new_n1011_, new_n888_ );
not g840 ( new_n1012_, keyIn_0_124 );
not g841 ( new_n1013_, new_n1008_ );
and g842 ( new_n1014_, new_n825_, new_n847_, new_n909_ );
and g843 ( new_n1015_, new_n1013_, new_n1012_, new_n1014_ );
or g844 ( new_n1016_, new_n1015_, new_n1011_ );
or g845 ( new_n1017_, new_n1016_, new_n1010_ );
or g846 ( new_n1018_, new_n960_, new_n1017_, new_n994_ );
and g847 ( new_n1019_, new_n1018_, keyIn_0_127 );
not g848 ( new_n1020_, keyIn_0_127 );
not g849 ( new_n1021_, new_n1017_ );
and g850 ( new_n1022_, new_n965_, new_n1020_, new_n1021_, new_n999_ );
or g851 ( N432, new_n1019_, new_n1022_ );
endmodule