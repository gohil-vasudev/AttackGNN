module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n445_, new_n236_, new_n238_, new_n479_, new_n250_, new_n501_, new_n288_, new_n421_, new_n368_, new_n439_, new_n283_, new_n223_, new_n366_, new_n241_, new_n365_, new_n339_, new_n401_, new_n389_, new_n514_, new_n456_, new_n246_, new_n266_, new_n367_, new_n542_, new_n548_, new_n220_, new_n214_, new_n451_, new_n489_, new_n240_, new_n413_, new_n526_, new_n442_, new_n211_, new_n552_, new_n342_, new_n462_, new_n564_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n427_, new_n234_, new_n532_, new_n393_, new_n418_, new_n292_, new_n215_, new_n257_, new_n212_, new_n364_, new_n449_, new_n484_, new_n272_, new_n282_, new_n414_, new_n315_, new_n326_, new_n554_, new_n230_, new_n281_, new_n430_, new_n482_, new_n248_, new_n350_, new_n385_, new_n478_, new_n461_, new_n297_, new_n361_, new_n565_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n530_, new_n318_, new_n321_, new_n443_, new_n324_, new_n486_, new_n491_, new_n549_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n305_, new_n420_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n506_, new_n256_, new_n452_, new_n381_, new_n388_, new_n508_, new_n483_, new_n394_, new_n299_, new_n314_, new_n363_, new_n441_, new_n216_, new_n280_, new_n235_, new_n398_, new_n301_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n311_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n349_, new_n244_, new_n488_, new_n524_, new_n277_, new_n402_, new_n286_, new_n335_, new_n347_, new_n346_, new_n438_, new_n208_, new_n436_, new_n397_, new_n399_, new_n559_, new_n233_, new_n469_, new_n391_, new_n437_, new_n295_, new_n359_, new_n409_, new_n457_, new_n553_, new_n333_, new_n290_, new_n448_, new_n276_, new_n384_, new_n410_, new_n543_, new_n509_, new_n454_, new_n202_, new_n296_, new_n308_, new_n232_, new_n258_, new_n306_, new_n494_, new_n291_, new_n261_, new_n309_, new_n529_, new_n323_, new_n259_, new_n362_, new_n227_, new_n416_, new_n222_, new_n400_, new_n328_, new_n460_, new_n505_, new_n471_, new_n268_, new_n374_, new_n376_, new_n380_, new_n310_, new_n275_, new_n352_, new_n485_, new_n525_, new_n562_, new_n547_, new_n264_, new_n379_, new_n273_, new_n224_, new_n270_, new_n520_, new_n253_, new_n403_, new_n475_, new_n237_, new_n557_, new_n260_, new_n251_, new_n300_, new_n480_, new_n513_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n522_, new_n487_, new_n360_, new_n546_, new_n302_, new_n225_, new_n387_, new_n544_, new_n476_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n499_, new_n255_, new_n533_, new_n459_, new_n555_, new_n468_, new_n354_, new_n444_, new_n518_, new_n340_, new_n285_, new_n209_, new_n337_, new_n446_, new_n203_, new_n316_, new_n417_, new_n515_, new_n332_, new_n453_, new_n516_, new_n563_, new_n440_, new_n531_, new_n252_, new_n312_, new_n535_, new_n372_, new_n242_, new_n503_, new_n527_, new_n307_, new_n408_, new_n470_, new_n213_, new_n433_, new_n435_, new_n265_, new_n370_, new_n278_, new_n304_, new_n550_, new_n217_, new_n269_, new_n512_, new_n412_, new_n327_, new_n495_, new_n431_, new_n319_, new_n338_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n294_, new_n357_, new_n320_, new_n245_, new_n474_, new_n404_, new_n490_, new_n560_, new_n358_, new_n348_, new_n322_, new_n228_, new_n545_, new_n289_, new_n425_, new_n226_, new_n540_, new_n434_, new_n329_, new_n249_, new_n284_, new_n293_, new_n279_, new_n455_, new_n521_, new_n406_, new_n356_, new_n229_, new_n536_, new_n464_, new_n204_, new_n405_;

xor g000 ( new_n202_, N89, N93 );
xor g001 ( new_n203_, new_n202_, keyIn_0_11 );
xor g002 ( new_n204_, N81, N85 );
xnor g003 ( new_n205_, new_n204_, keyIn_0_10 );
xnor g004 ( new_n206_, new_n203_, new_n205_ );
xnor g005 ( new_n207_, new_n206_, keyIn_0_33 );
xnor g006 ( new_n208_, N73, N77 );
xor g007 ( new_n209_, new_n208_, keyIn_0_9 );
xnor g008 ( new_n210_, N65, N69 );
xnor g009 ( new_n211_, new_n210_, keyIn_0_8 );
xnor g010 ( new_n212_, new_n209_, new_n211_ );
xnor g011 ( new_n213_, new_n212_, keyIn_0_32 );
xnor g012 ( new_n214_, new_n207_, new_n213_ );
xor g013 ( new_n215_, new_n214_, keyIn_0_43 );
and g014 ( new_n216_, N129, N137 );
xnor g015 ( new_n217_, new_n215_, new_n216_ );
xnor g016 ( new_n218_, new_n217_, keyIn_0_47 );
xor g017 ( new_n219_, N33, N49 );
xnor g018 ( new_n220_, N1, N17 );
xnor g019 ( new_n221_, new_n219_, new_n220_ );
xnor g020 ( new_n222_, new_n218_, new_n221_ );
xor g021 ( new_n223_, new_n222_, keyIn_0_55 );
not g022 ( new_n224_, new_n223_ );
xnor g023 ( new_n225_, N113, N117 );
xnor g024 ( new_n226_, new_n225_, keyIn_0_14 );
xor g025 ( new_n227_, N121, N125 );
xnor g026 ( new_n228_, new_n227_, keyIn_0_15 );
xnor g027 ( new_n229_, new_n228_, new_n226_ );
xor g028 ( new_n230_, new_n229_, keyIn_0_35 );
xnor g029 ( new_n231_, N105, N109 );
xnor g030 ( new_n232_, new_n231_, keyIn_0_13 );
xnor g031 ( new_n233_, N97, N101 );
xnor g032 ( new_n234_, new_n233_, keyIn_0_12 );
xnor g033 ( new_n235_, new_n232_, new_n234_ );
xnor g034 ( new_n236_, new_n235_, keyIn_0_34 );
xnor g035 ( new_n237_, new_n230_, new_n236_ );
xnor g036 ( new_n238_, new_n237_, keyIn_0_44 );
and g037 ( new_n239_, N130, N137 );
xnor g038 ( new_n240_, new_n238_, new_n239_ );
xnor g039 ( new_n241_, new_n240_, keyIn_0_48 );
xor g040 ( new_n242_, N37, N53 );
xnor g041 ( new_n243_, N5, N21 );
xnor g042 ( new_n244_, new_n242_, new_n243_ );
xnor g043 ( new_n245_, new_n241_, new_n244_ );
xnor g044 ( new_n246_, new_n245_, keyIn_0_56 );
not g045 ( new_n247_, new_n246_ );
xnor g046 ( new_n248_, N13, N29 );
xnor g047 ( new_n249_, new_n248_, keyIn_0_23 );
xnor g048 ( new_n250_, N45, N61 );
xnor g049 ( new_n251_, new_n249_, new_n250_ );
xnor g050 ( new_n252_, new_n207_, new_n230_ );
xnor g051 ( new_n253_, new_n252_, keyIn_0_46 );
and g052 ( new_n254_, N132, N137 );
xnor g053 ( new_n255_, new_n253_, new_n254_ );
xnor g054 ( new_n256_, new_n255_, keyIn_0_50 );
xnor g055 ( new_n257_, new_n256_, new_n251_ );
xor g056 ( new_n258_, new_n257_, keyIn_0_58 );
not g057 ( new_n259_, new_n258_ );
xnor g058 ( new_n260_, new_n213_, new_n236_ );
xnor g059 ( new_n261_, new_n260_, keyIn_0_45 );
and g060 ( new_n262_, N131, N137 );
xor g061 ( new_n263_, new_n262_, keyIn_0_16 );
xnor g062 ( new_n264_, new_n261_, new_n263_ );
xnor g063 ( new_n265_, new_n264_, keyIn_0_49 );
xor g064 ( new_n266_, N9, N25 );
xor g065 ( new_n267_, new_n266_, keyIn_0_21 );
xor g066 ( new_n268_, N41, N57 );
xnor g067 ( new_n269_, new_n268_, keyIn_0_22 );
xnor g068 ( new_n270_, new_n267_, new_n269_ );
xnor g069 ( new_n271_, new_n270_, keyIn_0_36 );
xnor g070 ( new_n272_, new_n265_, new_n271_ );
xor g071 ( new_n273_, new_n272_, keyIn_0_57 );
or g072 ( new_n274_, new_n259_, new_n247_, new_n273_ );
and g073 ( new_n275_, new_n258_, new_n246_ );
not g074 ( new_n276_, new_n273_ );
or g075 ( new_n277_, new_n275_, new_n276_ );
and g076 ( new_n278_, new_n259_, new_n247_ );
not g077 ( new_n279_, new_n278_ );
and g078 ( new_n280_, new_n277_, new_n279_, new_n223_, new_n274_ );
not g079 ( new_n281_, keyIn_0_63 );
or g080 ( new_n282_, new_n276_, new_n281_ );
and g081 ( new_n283_, new_n224_, new_n246_ );
or g082 ( new_n284_, new_n273_, keyIn_0_63 );
and g083 ( new_n285_, new_n283_, new_n258_, new_n282_, new_n284_ );
or g084 ( new_n286_, new_n280_, new_n285_ );
not g085 ( new_n287_, keyIn_0_60 );
xnor g086 ( new_n288_, N49, N53 );
xnor g087 ( new_n289_, new_n288_, keyIn_0_6 );
xnor g088 ( new_n290_, N57, N61 );
xnor g089 ( new_n291_, new_n290_, keyIn_0_7 );
xor g090 ( new_n292_, new_n289_, new_n291_ );
xnor g091 ( new_n293_, new_n292_, keyIn_0_31 );
not g092 ( new_n294_, keyIn_0_30 );
not g093 ( new_n295_, keyIn_0_4 );
xnor g094 ( new_n296_, N33, N37 );
xnor g095 ( new_n297_, new_n296_, new_n295_ );
xnor g096 ( new_n298_, N41, N45 );
xnor g097 ( new_n299_, new_n298_, keyIn_0_5 );
xnor g098 ( new_n300_, new_n297_, new_n299_ );
xnor g099 ( new_n301_, new_n300_, new_n294_ );
xnor g100 ( new_n302_, new_n293_, new_n301_ );
xnor g101 ( new_n303_, new_n302_, keyIn_0_40 );
and g102 ( new_n304_, N134, N137 );
xor g103 ( new_n305_, new_n304_, keyIn_0_18 );
xnor g104 ( new_n306_, new_n303_, new_n305_ );
xnor g105 ( new_n307_, new_n306_, keyIn_0_52 );
xor g106 ( new_n308_, N69, N85 );
xnor g107 ( new_n309_, new_n308_, keyIn_0_24 );
xnor g108 ( new_n310_, N101, N117 );
xnor g109 ( new_n311_, new_n310_, keyIn_0_25 );
xnor g110 ( new_n312_, new_n309_, new_n311_ );
xnor g111 ( new_n313_, new_n312_, keyIn_0_37 );
xnor g112 ( new_n314_, new_n307_, new_n313_ );
xnor g113 ( new_n315_, new_n314_, new_n287_ );
xnor g114 ( new_n316_, N25, N29 );
xnor g115 ( new_n317_, new_n316_, keyIn_0_3 );
xor g116 ( new_n318_, N17, N21 );
xnor g117 ( new_n319_, new_n318_, keyIn_0_2 );
xnor g118 ( new_n320_, new_n319_, new_n317_ );
xnor g119 ( new_n321_, new_n320_, keyIn_0_29 );
xnor g120 ( new_n322_, N1, N5 );
xnor g121 ( new_n323_, new_n322_, keyIn_0_0 );
xnor g122 ( new_n324_, N9, N13 );
xnor g123 ( new_n325_, new_n324_, keyIn_0_1 );
xnor g124 ( new_n326_, new_n323_, new_n325_ );
xnor g125 ( new_n327_, new_n326_, keyIn_0_28 );
xnor g126 ( new_n328_, new_n321_, new_n327_ );
xnor g127 ( new_n329_, new_n328_, keyIn_0_39 );
and g128 ( new_n330_, N133, N137 );
xor g129 ( new_n331_, new_n330_, keyIn_0_17 );
xnor g130 ( new_n332_, new_n329_, new_n331_ );
xnor g131 ( new_n333_, new_n332_, keyIn_0_51 );
xnor g132 ( new_n334_, N97, N113 );
xnor g133 ( new_n335_, N65, N81 );
xnor g134 ( new_n336_, new_n334_, new_n335_ );
xnor g135 ( new_n337_, new_n333_, new_n336_ );
xnor g136 ( new_n338_, new_n337_, keyIn_0_59 );
not g137 ( new_n339_, new_n338_ );
and g138 ( new_n340_, new_n339_, new_n315_ );
xnor g139 ( new_n341_, new_n301_, new_n327_ );
xnor g140 ( new_n342_, new_n341_, keyIn_0_41 );
and g141 ( new_n343_, N135, N137 );
xnor g142 ( new_n344_, new_n343_, keyIn_0_19 );
xnor g143 ( new_n345_, new_n342_, new_n344_ );
xnor g144 ( new_n346_, new_n345_, keyIn_0_53 );
xnor g145 ( new_n347_, N73, N89 );
xnor g146 ( new_n348_, new_n347_, keyIn_0_26 );
xor g147 ( new_n349_, N105, N121 );
xnor g148 ( new_n350_, new_n349_, keyIn_0_27 );
xnor g149 ( new_n351_, new_n350_, new_n348_ );
xnor g150 ( new_n352_, new_n351_, keyIn_0_38 );
xnor g151 ( new_n353_, new_n346_, new_n352_ );
xnor g152 ( new_n354_, new_n353_, keyIn_0_61 );
xnor g153 ( new_n355_, new_n293_, new_n321_ );
xnor g154 ( new_n356_, new_n355_, keyIn_0_42 );
and g155 ( new_n357_, N136, N137 );
xnor g156 ( new_n358_, new_n357_, keyIn_0_20 );
xnor g157 ( new_n359_, new_n356_, new_n358_ );
xnor g158 ( new_n360_, new_n359_, keyIn_0_54 );
xor g159 ( new_n361_, N109, N125 );
xnor g160 ( new_n362_, N77, N93 );
xnor g161 ( new_n363_, new_n361_, new_n362_ );
xnor g162 ( new_n364_, new_n360_, new_n363_ );
xnor g163 ( new_n365_, new_n364_, keyIn_0_62 );
and g164 ( new_n366_, new_n365_, new_n354_ );
and g165 ( new_n367_, new_n286_, new_n340_, new_n366_ );
and g166 ( new_n368_, new_n367_, new_n224_ );
xor g167 ( N724, new_n368_, N1 );
and g168 ( new_n370_, new_n367_, new_n247_ );
xor g169 ( N725, new_n370_, N5 );
and g170 ( new_n372_, new_n367_, new_n273_ );
xor g171 ( N726, new_n372_, N9 );
and g172 ( new_n374_, new_n367_, new_n259_ );
xor g173 ( N727, new_n374_, N13 );
not g174 ( new_n376_, keyIn_0_76 );
not g175 ( new_n377_, new_n354_ );
not g176 ( new_n378_, new_n365_ );
and g177 ( new_n379_, new_n286_, new_n340_, new_n377_, new_n378_ );
and g178 ( new_n380_, new_n379_, new_n376_ );
not g179 ( new_n381_, new_n380_ );
or g180 ( new_n382_, new_n379_, new_n376_ );
and g181 ( new_n383_, new_n381_, new_n224_, new_n382_ );
xnor g182 ( new_n384_, new_n383_, keyIn_0_82 );
xor g183 ( new_n385_, new_n384_, N17 );
xnor g184 ( N728, new_n385_, keyIn_0_105 );
and g185 ( new_n387_, new_n381_, new_n247_, new_n382_ );
xor g186 ( new_n388_, new_n387_, keyIn_0_83 );
xnor g187 ( new_n389_, new_n388_, N21 );
xor g188 ( N729, new_n389_, keyIn_0_106 );
and g189 ( new_n391_, new_n381_, new_n273_, new_n382_ );
xor g190 ( N730, new_n391_, N25 );
and g191 ( new_n393_, new_n381_, new_n259_, new_n382_ );
xnor g192 ( new_n394_, new_n393_, keyIn_0_84 );
xnor g193 ( new_n395_, new_n394_, N29 );
xor g194 ( N731, new_n395_, keyIn_0_107 );
not g195 ( new_n397_, keyIn_0_77 );
or g196 ( new_n398_, new_n339_, new_n315_ );
not g197 ( new_n399_, new_n398_ );
and g198 ( new_n400_, new_n286_, new_n366_, new_n399_ );
and g199 ( new_n401_, new_n400_, new_n397_ );
not g200 ( new_n402_, new_n401_ );
or g201 ( new_n403_, new_n400_, new_n397_ );
and g202 ( new_n404_, new_n402_, new_n224_, new_n403_ );
xor g203 ( new_n405_, new_n404_, keyIn_0_85 );
xnor g204 ( new_n406_, new_n405_, N33 );
xnor g205 ( N732, new_n406_, keyIn_0_108 );
and g206 ( new_n408_, new_n402_, new_n247_, new_n403_ );
xnor g207 ( new_n409_, new_n408_, keyIn_0_86 );
xnor g208 ( new_n410_, new_n409_, N37 );
xor g209 ( N733, new_n410_, keyIn_0_109 );
and g210 ( new_n412_, new_n402_, new_n273_, new_n403_ );
xnor g211 ( new_n413_, new_n412_, keyIn_0_87 );
xor g212 ( new_n414_, new_n413_, N41 );
xnor g213 ( N734, new_n414_, keyIn_0_110 );
and g214 ( new_n416_, new_n402_, new_n259_, new_n403_ );
xnor g215 ( new_n417_, new_n416_, keyIn_0_88 );
xor g216 ( new_n418_, new_n417_, N45 );
xnor g217 ( N735, new_n418_, keyIn_0_111 );
and g218 ( new_n420_, new_n286_, new_n377_, new_n378_, new_n399_ );
and g219 ( new_n421_, new_n420_, new_n224_ );
xor g220 ( N736, new_n421_, N49 );
and g221 ( new_n423_, new_n420_, new_n247_ );
xor g222 ( N737, new_n423_, N53 );
and g223 ( new_n425_, new_n420_, new_n273_ );
xor g224 ( N738, new_n425_, N57 );
and g225 ( new_n427_, new_n420_, new_n259_ );
xor g226 ( N739, new_n427_, N61 );
not g227 ( new_n429_, N65 );
not g228 ( new_n430_, keyIn_0_65 );
xnor g229 ( new_n431_, new_n354_, new_n430_ );
not g230 ( new_n432_, new_n431_ );
or g231 ( new_n433_, new_n432_, new_n398_, keyIn_0_73, new_n378_ );
and g232 ( new_n434_, new_n315_, new_n365_, new_n338_, new_n354_ );
xor g233 ( new_n435_, new_n434_, keyIn_0_72 );
not g234 ( new_n436_, keyIn_0_73 );
xnor g235 ( new_n437_, new_n314_, keyIn_0_60 );
and g236 ( new_n438_, new_n437_, new_n365_, new_n338_ );
and g237 ( new_n439_, new_n431_, new_n438_ );
or g238 ( new_n440_, new_n439_, new_n436_ );
and g239 ( new_n441_, new_n440_, new_n435_ );
not g240 ( new_n442_, keyIn_0_71 );
and g241 ( new_n443_, new_n315_, new_n338_ );
not g242 ( new_n444_, keyIn_0_64 );
or g243 ( new_n445_, new_n377_, new_n444_ );
or g244 ( new_n446_, new_n354_, keyIn_0_64 );
and g245 ( new_n447_, new_n445_, new_n446_, new_n443_, new_n378_ );
xnor g246 ( new_n448_, new_n447_, new_n442_ );
not g247 ( new_n449_, keyIn_0_74 );
not g248 ( new_n450_, keyIn_0_66 );
xnor g249 ( new_n451_, new_n354_, new_n450_ );
and g250 ( new_n452_, new_n451_, new_n340_, new_n365_ );
xnor g251 ( new_n453_, new_n452_, new_n449_ );
and g252 ( new_n454_, new_n441_, new_n433_, new_n448_, new_n453_ );
xnor g253 ( new_n455_, new_n454_, keyIn_0_75 );
not g254 ( new_n456_, new_n455_ );
xnor g255 ( new_n457_, new_n246_, keyIn_0_67 );
and g256 ( new_n458_, new_n457_, new_n224_, new_n258_, new_n273_ );
not g257 ( new_n459_, new_n458_ );
or g258 ( new_n460_, new_n456_, keyIn_0_78, new_n459_ );
not g259 ( new_n461_, keyIn_0_78 );
and g260 ( new_n462_, new_n455_, new_n458_ );
or g261 ( new_n463_, new_n462_, new_n461_ );
and g262 ( new_n464_, new_n463_, new_n339_, new_n460_ );
xnor g263 ( new_n465_, new_n464_, keyIn_0_89 );
xnor g264 ( new_n466_, new_n465_, new_n429_ );
xnor g265 ( N740, new_n466_, keyIn_0_112 );
not g266 ( new_n468_, keyIn_0_113 );
and g267 ( new_n469_, new_n463_, new_n437_, new_n460_ );
xnor g268 ( new_n470_, new_n469_, keyIn_0_90 );
xnor g269 ( new_n471_, new_n470_, N69 );
xnor g270 ( N741, new_n471_, new_n468_ );
not g271 ( new_n473_, keyIn_0_114 );
and g272 ( new_n474_, new_n463_, new_n354_, new_n460_ );
xnor g273 ( new_n475_, new_n474_, keyIn_0_91 );
xnor g274 ( new_n476_, new_n475_, N73 );
xnor g275 ( N742, new_n476_, new_n473_ );
and g276 ( new_n478_, new_n463_, new_n378_, new_n460_ );
xnor g277 ( new_n479_, new_n478_, keyIn_0_92 );
xnor g278 ( new_n480_, new_n479_, N77 );
xnor g279 ( N743, new_n480_, keyIn_0_115 );
not g280 ( new_n482_, keyIn_0_116 );
not g281 ( new_n483_, keyIn_0_79 );
xnor g282 ( new_n484_, new_n273_, keyIn_0_68 );
and g283 ( new_n485_, new_n283_, new_n259_, new_n484_ );
not g284 ( new_n486_, new_n485_ );
or g285 ( new_n487_, new_n456_, new_n483_, new_n486_ );
and g286 ( new_n488_, new_n455_, new_n485_ );
or g287 ( new_n489_, new_n488_, keyIn_0_79 );
and g288 ( new_n490_, new_n489_, new_n339_, new_n487_ );
xnor g289 ( new_n491_, new_n490_, keyIn_0_93 );
xnor g290 ( new_n492_, new_n491_, N81 );
xnor g291 ( N744, new_n492_, new_n482_ );
and g292 ( new_n494_, new_n489_, new_n437_, new_n487_ );
xnor g293 ( new_n495_, new_n494_, keyIn_0_94 );
xnor g294 ( new_n496_, new_n495_, N85 );
xnor g295 ( N745, new_n496_, keyIn_0_117 );
not g296 ( new_n498_, keyIn_0_118 );
and g297 ( new_n499_, new_n489_, new_n354_, new_n487_ );
xnor g298 ( new_n500_, new_n499_, keyIn_0_95 );
xnor g299 ( new_n501_, new_n500_, N89 );
xnor g300 ( N746, new_n501_, new_n498_ );
not g301 ( new_n503_, keyIn_0_119 );
and g302 ( new_n504_, new_n489_, new_n378_, new_n487_ );
xnor g303 ( new_n505_, new_n504_, keyIn_0_96 );
xnor g304 ( new_n506_, new_n505_, N93 );
xnor g305 ( N747, new_n506_, new_n503_ );
not g306 ( new_n508_, keyIn_0_120 );
not g307 ( new_n509_, keyIn_0_97 );
and g308 ( new_n510_, new_n223_, new_n247_, new_n258_, new_n273_ );
not g309 ( new_n511_, new_n510_ );
or g310 ( new_n512_, new_n456_, keyIn_0_80, new_n511_ );
not g311 ( new_n513_, keyIn_0_80 );
and g312 ( new_n514_, new_n455_, new_n510_ );
or g313 ( new_n515_, new_n514_, new_n513_ );
and g314 ( new_n516_, new_n515_, new_n339_, new_n512_ );
xnor g315 ( new_n517_, new_n516_, new_n509_ );
xnor g316 ( new_n518_, new_n517_, N97 );
xnor g317 ( N748, new_n518_, new_n508_ );
and g318 ( new_n520_, new_n515_, new_n437_, new_n512_ );
xnor g319 ( new_n521_, new_n520_, keyIn_0_98 );
xnor g320 ( new_n522_, new_n521_, N101 );
xnor g321 ( N749, new_n522_, keyIn_0_121 );
not g322 ( new_n524_, keyIn_0_99 );
and g323 ( new_n525_, new_n515_, new_n354_, new_n512_ );
xnor g324 ( new_n526_, new_n525_, new_n524_ );
xnor g325 ( new_n527_, new_n526_, N105 );
xnor g326 ( N750, new_n527_, keyIn_0_122 );
not g327 ( new_n529_, keyIn_0_123 );
not g328 ( new_n530_, keyIn_0_100 );
and g329 ( new_n531_, new_n515_, new_n378_, new_n512_ );
xnor g330 ( new_n532_, new_n531_, new_n530_ );
xnor g331 ( new_n533_, new_n532_, N109 );
xnor g332 ( N751, new_n533_, new_n529_ );
not g333 ( new_n535_, keyIn_0_81 );
and g334 ( new_n536_, new_n276_, keyIn_0_70 );
not g335 ( new_n537_, new_n536_ );
and g336 ( new_n538_, new_n224_, keyIn_0_69 );
not g337 ( new_n539_, new_n538_ );
or g338 ( new_n540_, new_n276_, keyIn_0_70 );
or g339 ( new_n541_, new_n224_, keyIn_0_69 );
and g340 ( new_n542_, new_n541_, new_n540_ );
and g341 ( new_n543_, new_n542_, new_n278_, new_n537_, new_n539_ );
and g342 ( new_n544_, new_n455_, new_n543_ );
or g343 ( new_n545_, new_n544_, new_n535_ );
not g344 ( new_n546_, new_n543_ );
or g345 ( new_n547_, new_n456_, keyIn_0_81, new_n546_ );
and g346 ( new_n548_, new_n545_, new_n339_, new_n547_ );
xnor g347 ( new_n549_, new_n548_, keyIn_0_101 );
xnor g348 ( new_n550_, new_n549_, N113 );
xnor g349 ( N752, new_n550_, keyIn_0_124 );
not g350 ( new_n552_, keyIn_0_125 );
and g351 ( new_n553_, new_n545_, new_n437_, new_n547_ );
xnor g352 ( new_n554_, new_n553_, keyIn_0_102 );
xnor g353 ( new_n555_, new_n554_, N117 );
xnor g354 ( N753, new_n555_, new_n552_ );
not g355 ( new_n557_, N121 );
and g356 ( new_n558_, new_n545_, new_n354_, new_n547_ );
xnor g357 ( new_n559_, new_n558_, keyIn_0_103 );
xnor g358 ( new_n560_, new_n559_, new_n557_ );
xnor g359 ( N754, new_n560_, keyIn_0_126 );
not g360 ( new_n562_, keyIn_0_127 );
and g361 ( new_n563_, new_n545_, new_n378_, new_n547_ );
xnor g362 ( new_n564_, new_n563_, keyIn_0_104 );
xnor g363 ( new_n565_, new_n564_, N125 );
xnor g364 ( N755, new_n565_, new_n562_ );
endmodule