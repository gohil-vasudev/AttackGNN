module add_mul_mix_32_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, 
        a_18_, a_19_, a_20_, a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, 
        a_28_, a_29_, a_30_, a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, 
        b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, 
        b_17_, b_18_, b_19_, b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, 
        b_27_, b_28_, b_29_, b_30_, b_31_, c_0_, c_1_, c_2_, c_3_, c_4_, c_5_, 
        c_6_, c_7_, c_8_, c_9_, c_10_, c_11_, c_12_, c_13_, c_14_, c_15_, 
        c_16_, c_17_, c_18_, c_19_, c_20_, c_21_, c_22_, c_23_, c_24_, c_25_, 
        c_26_, c_27_, c_28_, c_29_, c_30_, c_31_, d_0_, d_1_, d_2_, d_3_, d_4_, 
        d_5_, d_6_, d_7_, d_8_, d_9_, d_10_, d_11_, d_12_, d_13_, d_14_, d_15_, 
        d_16_, d_17_, d_18_, d_19_, d_20_, d_21_, d_22_, d_23_, d_24_, d_25_, 
        d_26_, d_27_, d_28_, d_29_, d_30_, d_31_, Result_0_, Result_1_, 
        Result_2_, Result_3_, Result_4_, Result_5_, Result_6_, Result_7_, 
        Result_8_, Result_9_, Result_10_, Result_11_, Result_12_, Result_13_, 
        Result_14_, Result_15_, Result_16_, Result_17_, Result_18_, Result_19_, 
        Result_20_, Result_21_, Result_22_, Result_23_, Result_24_, Result_25_, 
        Result_26_, Result_27_, Result_28_, Result_29_, Result_30_, Result_31_, 
        Result_32_, Result_33_, Result_34_, Result_35_, Result_36_, Result_37_, 
        Result_38_, Result_39_, Result_40_, Result_41_, Result_42_, Result_43_, 
        Result_44_, Result_45_, Result_46_, Result_47_, Result_48_, Result_49_, 
        Result_50_, Result_51_, Result_52_, Result_53_, Result_54_, Result_55_, 
        Result_56_, Result_57_, Result_58_, Result_59_, Result_60_, Result_61_, 
        Result_62_, Result_63_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, a_19_, a_20_,
         a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, a_29_, a_30_,
         a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_,
         b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, b_18_, b_19_,
         b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, b_28_, b_29_,
         b_30_, b_31_, c_0_, c_1_, c_2_, c_3_, c_4_, c_5_, c_6_, c_7_, c_8_,
         c_9_, c_10_, c_11_, c_12_, c_13_, c_14_, c_15_, c_16_, c_17_, c_18_,
         c_19_, c_20_, c_21_, c_22_, c_23_, c_24_, c_25_, c_26_, c_27_, c_28_,
         c_29_, c_30_, c_31_, d_0_, d_1_, d_2_, d_3_, d_4_, d_5_, d_6_, d_7_,
         d_8_, d_9_, d_10_, d_11_, d_12_, d_13_, d_14_, d_15_, d_16_, d_17_,
         d_18_, d_19_, d_20_, d_21_, d_22_, d_23_, d_24_, d_25_, d_26_, d_27_,
         d_28_, d_29_, d_30_, d_31_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_,
         Result_32_, Result_33_, Result_34_, Result_35_, Result_36_,
         Result_37_, Result_38_, Result_39_, Result_40_, Result_41_,
         Result_42_, Result_43_, Result_44_, Result_45_, Result_46_,
         Result_47_, Result_48_, Result_49_, Result_50_, Result_51_,
         Result_52_, Result_53_, Result_54_, Result_55_, Result_56_,
         Result_57_, Result_58_, Result_59_, Result_60_, Result_61_,
         Result_62_, Result_63_;
  wire   n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,
         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,
         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,
         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,
         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,
         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
         n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
         n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
         n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088,
         n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,
         n17097, n17098;

  NAND2_X1 U8576 ( .A1(n16923), .A2(n16924), .ZN(n12731) );
  NAND2_X1 U8577 ( .A1(n16927), .A2(n16928), .ZN(n12460) );
  NAND2_X1 U8578 ( .A1(n16919), .A2(n16920), .ZN(n12984) );
  NAND2_X1 U8579 ( .A1(n17051), .A2(n17052), .ZN(n16810) );
  NAND2_X1 U8580 ( .A1(n17047), .A2(n17048), .ZN(n16812) );
  NAND2_X1 U8581 ( .A1(n17031), .A2(n17032), .ZN(n16821) );
  NAND2_X1 U8582 ( .A1(n17027), .A2(n17028), .ZN(n16823) );
  NAND2_X1 U8583 ( .A1(n17015), .A2(n17016), .ZN(n16831) );
  NAND2_X1 U8584 ( .A1(n16963), .A2(n16964), .ZN(n10256) );
  NAND2_X1 U8585 ( .A1(n16947), .A2(n16948), .ZN(n11185) );
  NAND2_X1 U8586 ( .A1(n16935), .A2(n16936), .ZN(n11939) );
  NAND2_X1 U8587 ( .A1(n16863), .A2(n16864), .ZN(n16552) );
  NAND2_X1 U8588 ( .A1(n17087), .A2(n17088), .ZN(n16791) );
  NAND2_X1 U8589 ( .A1(n17075), .A2(n17076), .ZN(n16797) );
  NAND2_X1 U8590 ( .A1(n17059), .A2(n17060), .ZN(n16805) );
  NAND2_X1 U8591 ( .A1(n17055), .A2(n17056), .ZN(n16808) );
  NAND2_X1 U8592 ( .A1(n16983), .A2(n16984), .ZN(n16428) );
  XNOR2_X1 U8593 ( .A(b_30_), .B(n16784), .ZN(n16783) );
  XOR2_X1 U8594 ( .A(d_30_), .B(c_30_), .Z(n9397) );
  XOR2_X1 U8595 ( .A(n16795), .B(n16796), .Z(n8512) );
  XOR2_X1 U8596 ( .A(n16843), .B(n16844), .Z(n8513) );
  XOR2_X1 U8597 ( .A(n16856), .B(n16857), .Z(n8514) );
  XOR2_X1 U8598 ( .A(n16803), .B(n16804), .Z(n8515) );
  XOR2_X1 U8599 ( .A(n16799), .B(n16800), .Z(n8516) );
  XOR2_X1 U8600 ( .A(n16817), .B(n16818), .Z(n8517) );
  XOR2_X1 U8601 ( .A(n10505), .B(n10506), .Z(n8518) );
  XOR2_X1 U8602 ( .A(n15271), .B(n15272), .Z(n8519) );
  XOR2_X1 U8603 ( .A(n13742), .B(n13743), .Z(n8520) );
  XOR2_X1 U8604 ( .A(n15777), .B(n15778), .Z(n8521) );
  XOR2_X1 U8605 ( .A(n15050), .B(n15051), .Z(n8522) );
  XOR2_X1 U8606 ( .A(n14764), .B(n14765), .Z(n8523) );
  XOR2_X1 U8607 ( .A(n14546), .B(n14547), .Z(n8524) );
  NAND2_X2 U8608 ( .A1(n8585), .A2(n8538), .ZN(n8624) );
  NAND2_X2 U8609 ( .A1(n16551), .A2(n8539), .ZN(n8630) );
  INV_X2 U8610 ( .A(n8534), .ZN(n14761) );
  INV_X2 U8611 ( .A(n8525), .ZN(n14248) );
  INV_X2 U8612 ( .A(n8523), .ZN(n8525) );
  INV_X2 U8613 ( .A(n8529), .ZN(n15268) );
  INV_X2 U8614 ( .A(n8524), .ZN(n8526) );
  INV_X2 U8615 ( .A(n8514), .ZN(n8527) );
  INV_X2 U8616 ( .A(n8513), .ZN(n8528) );
  INV_X2 U8617 ( .A(n8521), .ZN(n8529) );
  INV_X2 U8618 ( .A(n8522), .ZN(n8530) );
  INV_X2 U8619 ( .A(n8520), .ZN(n8531) );
  INV_X1 U8620 ( .A(n15557), .ZN(n8532) );
  INV_X2 U8621 ( .A(n8532), .ZN(n8533) );
  INV_X2 U8622 ( .A(n8519), .ZN(n8534) );
  INV_X2 U8623 ( .A(n8512), .ZN(n8535) );
  INV_X1 U8624 ( .A(n9149), .ZN(n8536) );
  INV_X2 U8625 ( .A(n8536), .ZN(n8537) );
  INV_X1 U8626 ( .A(n8632), .ZN(n8538) );
  INV_X2 U8627 ( .A(n8538), .ZN(n8539) );
  INV_X1 U8628 ( .A(n10410), .ZN(n8540) );
  INV_X2 U8629 ( .A(n8540), .ZN(n8541) );
  INV_X2 U8630 ( .A(n8518), .ZN(n8542) );
  INV_X1 U8631 ( .A(n9005), .ZN(n8543) );
  INV_X2 U8632 ( .A(n8543), .ZN(n8544) );
  INV_X2 U8633 ( .A(n8517), .ZN(n8545) );
  INV_X1 U8634 ( .A(n10804), .ZN(n8546) );
  INV_X2 U8635 ( .A(n8546), .ZN(n8547) );
  INV_X2 U8636 ( .A(n8516), .ZN(n8548) );
  INV_X1 U8637 ( .A(n9393), .ZN(n8549) );
  INV_X2 U8638 ( .A(n8549), .ZN(n8550) );
  INV_X2 U8639 ( .A(n8515), .ZN(n8551) );
  INV_X1 U8640 ( .A(n9268), .ZN(n8552) );
  XNOR2_X1 U8641 ( .A(n16975), .B(n16976), .ZN(n8982) );
  INV_X1 U8642 ( .A(n13504), .ZN(n8553) );
  INV_X1 U8643 ( .A(n15047), .ZN(n8554) );
  INV_X2 U8644 ( .A(n8982), .ZN(n9268) );
  INV_X1 U8645 ( .A(n9286), .ZN(n8555) );
  INV_X1 U8646 ( .A(n9304), .ZN(n8556) );
  INV_X1 U8647 ( .A(n12728), .ZN(n8557) );
  XNOR2_X2 U8648 ( .A(n16848), .B(n16849), .ZN(n8874) );
  INV_X1 U8649 ( .A(n11686), .ZN(n8558) );
  INV_X1 U8650 ( .A(n11182), .ZN(n8559) );
  INV_X1 U8651 ( .A(n9295), .ZN(n8560) );
  INV_X1 U8652 ( .A(n13739), .ZN(n8561) );
  INV_X1 U8653 ( .A(n9322), .ZN(n8562) );
  INV_X1 U8654 ( .A(n9098), .ZN(n8563) );
  INV_X1 U8655 ( .A(n10307), .ZN(n8564) );
  INV_X1 U8656 ( .A(n9138), .ZN(n8565) );
  INV_X1 U8657 ( .A(n9146), .ZN(n8566) );
  INV_X1 U8658 ( .A(n8566), .ZN(n8567) );
  INV_X1 U8659 ( .A(n9373), .ZN(n8568) );
  INV_X1 U8660 ( .A(n9331), .ZN(n8569) );
  INV_X1 U8661 ( .A(n12981), .ZN(n8570) );
  INV_X1 U8662 ( .A(n10159), .ZN(n8571) );
  INV_X1 U8663 ( .A(n9209), .ZN(n8572) );
  INV_X1 U8664 ( .A(n9157), .ZN(n8573) );
  INV_X1 U8665 ( .A(n9132), .ZN(n8574) );
  INV_X1 U8666 ( .A(n11936), .ZN(n8575) );
  INV_X1 U8667 ( .A(n10667), .ZN(n8576) );
  INV_X1 U8668 ( .A(n16040), .ZN(n8577) );
  INV_X1 U8669 ( .A(n12196), .ZN(n8578) );
  INV_X1 U8670 ( .A(n15774), .ZN(n8579) );
  INV_X2 U8671 ( .A(n15773), .ZN(n15774) );
  INV_X1 U8672 ( .A(n9070), .ZN(n8580) );
  INV_X1 U8673 ( .A(n11432), .ZN(n8581) );
  INV_X1 U8674 ( .A(n9313), .ZN(n8582) );
  INV_X1 U8675 ( .A(n9340), .ZN(n8583) );
  INV_X1 U8676 ( .A(n9112), .ZN(n8584) );
  INV_X1 U8677 ( .A(n16551), .ZN(n8585) );
  INV_X1 U8678 ( .A(n9650), .ZN(n8586) );
  INV_X1 U8679 ( .A(n12457), .ZN(n8587) );
  INV_X1 U8680 ( .A(n9080), .ZN(n8588) );
  INV_X1 U8681 ( .A(n9263), .ZN(n8589) );
  INV_X1 U8682 ( .A(n16285), .ZN(n8590) );
  INV_X2 U8683 ( .A(n16284), .ZN(n16285) );
  INV_X1 U8684 ( .A(n9721), .ZN(n8591) );
  INV_X1 U8685 ( .A(n8972), .ZN(n8592) );
  INV_X2 U8686 ( .A(n10722), .ZN(n8593) );
  INV_X2 U8687 ( .A(n10846), .ZN(n8594) );
  XNOR2_X1 U8688 ( .A(n9396), .B(n9397), .ZN(n8626) );
  INV_X1 U8689 ( .A(n8626), .ZN(n8595) );
  INV_X1 U8690 ( .A(n8626), .ZN(n8596) );
  XOR2_X1 U8691 ( .A(n8597), .B(n8598), .Z(Result_9_) );
  NOR2_X1 U8692 ( .A1(n8599), .A2(n8600), .ZN(n8598) );
  NOR2_X1 U8693 ( .A1(n8601), .A2(n8602), .ZN(n8600) );
  INV_X1 U8694 ( .A(n8603), .ZN(n8602) );
  NOR2_X1 U8695 ( .A1(n8604), .A2(n8605), .ZN(n8601) );
  XOR2_X1 U8696 ( .A(n8606), .B(n8607), .Z(Result_8_) );
  XNOR2_X1 U8697 ( .A(n8608), .B(n8609), .ZN(Result_7_) );
  NOR2_X1 U8698 ( .A1(n8610), .A2(n8611), .ZN(n8609) );
  NOR2_X1 U8699 ( .A1(n8612), .A2(n8613), .ZN(n8611) );
  INV_X1 U8700 ( .A(n8614), .ZN(n8613) );
  NOR2_X1 U8701 ( .A1(n8615), .A2(n8616), .ZN(n8612) );
  XOR2_X1 U8702 ( .A(n8617), .B(n8618), .Z(Result_6_) );
  NOR2_X1 U8703 ( .A1(n8538), .A2(n8619), .ZN(Result_63_) );
  NAND2_X1 U8704 ( .A1(n8620), .A2(n8621), .ZN(Result_62_) );
  NAND2_X1 U8705 ( .A1(n8622), .A2(n8623), .ZN(n8621) );
  NAND2_X1 U8706 ( .A1(n8624), .A2(n8625), .ZN(n8623) );
  NAND2_X1 U8707 ( .A1(n8596), .A2(n8585), .ZN(n8625) );
  NAND2_X1 U8708 ( .A1(n8628), .A2(n8629), .ZN(n8620) );
  NAND2_X1 U8709 ( .A1(n8630), .A2(n8631), .ZN(n8629) );
  NAND2_X1 U8710 ( .A1(n8539), .A2(n8619), .ZN(n8631) );
  XOR2_X1 U8711 ( .A(n8633), .B(n8634), .Z(Result_61_) );
  XOR2_X1 U8712 ( .A(n8635), .B(n8636), .Z(n8634) );
  XNOR2_X1 U8713 ( .A(n8637), .B(n8638), .ZN(Result_60_) );
  NAND2_X1 U8714 ( .A1(n8639), .A2(n8640), .ZN(n8637) );
  XNOR2_X1 U8715 ( .A(n8641), .B(n8642), .ZN(Result_5_) );
  NOR2_X1 U8716 ( .A1(n8643), .A2(n8644), .ZN(n8642) );
  NOR2_X1 U8717 ( .A1(n8645), .A2(n8646), .ZN(n8644) );
  INV_X1 U8718 ( .A(n8647), .ZN(n8646) );
  NOR2_X1 U8719 ( .A1(n8648), .A2(n8649), .ZN(n8645) );
  XNOR2_X1 U8720 ( .A(n8650), .B(n8651), .ZN(Result_59_) );
  XOR2_X1 U8721 ( .A(n8652), .B(n8653), .Z(n8651) );
  XNOR2_X1 U8722 ( .A(n8654), .B(n8655), .ZN(Result_58_) );
  XNOR2_X1 U8723 ( .A(n8656), .B(n8657), .ZN(n8655) );
  XOR2_X1 U8724 ( .A(n8658), .B(n8659), .Z(Result_57_) );
  XNOR2_X1 U8725 ( .A(n8660), .B(n8661), .ZN(n8658) );
  XNOR2_X1 U8726 ( .A(n8662), .B(n8663), .ZN(Result_56_) );
  NAND2_X1 U8727 ( .A1(n8664), .A2(n8665), .ZN(n8662) );
  XNOR2_X1 U8728 ( .A(n8666), .B(n8667), .ZN(Result_55_) );
  XOR2_X1 U8729 ( .A(n8668), .B(n8669), .Z(n8667) );
  XNOR2_X1 U8730 ( .A(n8670), .B(n8671), .ZN(Result_54_) );
  NAND2_X1 U8731 ( .A1(n8672), .A2(n8673), .ZN(n8670) );
  XNOR2_X1 U8732 ( .A(n8674), .B(n8675), .ZN(Result_53_) );
  XOR2_X1 U8733 ( .A(n8676), .B(n8677), .Z(n8675) );
  XNOR2_X1 U8734 ( .A(n8678), .B(n8679), .ZN(Result_52_) );
  NAND2_X1 U8735 ( .A1(n8680), .A2(n8681), .ZN(n8678) );
  XNOR2_X1 U8736 ( .A(n8682), .B(n8683), .ZN(Result_51_) );
  XOR2_X1 U8737 ( .A(n8684), .B(n8685), .Z(n8683) );
  XOR2_X1 U8738 ( .A(n8686), .B(n8687), .Z(Result_50_) );
  XOR2_X1 U8739 ( .A(n8688), .B(n8689), .Z(n8686) );
  XOR2_X1 U8740 ( .A(n8690), .B(n8691), .Z(Result_4_) );
  XOR2_X1 U8741 ( .A(n8692), .B(n8693), .Z(Result_49_) );
  XOR2_X1 U8742 ( .A(n8694), .B(n8695), .Z(n8693) );
  XNOR2_X1 U8743 ( .A(n8696), .B(n8697), .ZN(Result_48_) );
  XNOR2_X1 U8744 ( .A(n8698), .B(n8699), .ZN(n8697) );
  XNOR2_X1 U8745 ( .A(n8700), .B(n8701), .ZN(Result_47_) );
  XNOR2_X1 U8746 ( .A(n8702), .B(n8703), .ZN(n8701) );
  XOR2_X1 U8747 ( .A(n8704), .B(n8705), .Z(Result_46_) );
  XOR2_X1 U8748 ( .A(n8706), .B(n8707), .Z(n8705) );
  XNOR2_X1 U8749 ( .A(n8708), .B(n8709), .ZN(Result_45_) );
  XNOR2_X1 U8750 ( .A(n8710), .B(n8711), .ZN(n8709) );
  XOR2_X1 U8751 ( .A(n8712), .B(n8713), .Z(Result_44_) );
  XNOR2_X1 U8752 ( .A(n8714), .B(n8715), .ZN(n8713) );
  XNOR2_X1 U8753 ( .A(n8716), .B(n8717), .ZN(Result_43_) );
  XNOR2_X1 U8754 ( .A(n8718), .B(n8719), .ZN(n8716) );
  XOR2_X1 U8755 ( .A(n8720), .B(n8721), .Z(Result_42_) );
  XOR2_X1 U8756 ( .A(n8722), .B(n8723), .Z(n8721) );
  XNOR2_X1 U8757 ( .A(n8724), .B(n8725), .ZN(Result_41_) );
  XNOR2_X1 U8758 ( .A(n8726), .B(n8727), .ZN(n8724) );
  XOR2_X1 U8759 ( .A(n8728), .B(n8729), .Z(Result_40_) );
  XOR2_X1 U8760 ( .A(n8730), .B(n8731), .Z(n8729) );
  XNOR2_X1 U8761 ( .A(n8732), .B(n8733), .ZN(Result_3_) );
  NOR2_X1 U8762 ( .A1(n8734), .A2(n8735), .ZN(n8733) );
  NOR2_X1 U8763 ( .A1(n8736), .A2(n8737), .ZN(n8735) );
  INV_X1 U8764 ( .A(n8738), .ZN(n8737) );
  NOR2_X1 U8765 ( .A1(n8739), .A2(n8740), .ZN(n8736) );
  XOR2_X1 U8766 ( .A(n8741), .B(n8742), .Z(Result_39_) );
  XOR2_X1 U8767 ( .A(n8743), .B(n8744), .Z(n8741) );
  XNOR2_X1 U8768 ( .A(n8745), .B(n8746), .ZN(Result_38_) );
  XNOR2_X1 U8769 ( .A(n8747), .B(n8748), .ZN(n8746) );
  XOR2_X1 U8770 ( .A(n8749), .B(n8750), .Z(Result_37_) );
  XOR2_X1 U8771 ( .A(n8751), .B(n8752), .Z(n8749) );
  XOR2_X1 U8772 ( .A(n8753), .B(n8754), .Z(Result_36_) );
  XOR2_X1 U8773 ( .A(n8755), .B(n8756), .Z(n8754) );
  XOR2_X1 U8774 ( .A(n8757), .B(n8758), .Z(Result_35_) );
  XOR2_X1 U8775 ( .A(n8759), .B(n8760), .Z(n8757) );
  XOR2_X1 U8776 ( .A(n8761), .B(n8762), .Z(Result_34_) );
  XOR2_X1 U8777 ( .A(n8763), .B(n8764), .Z(n8762) );
  XOR2_X1 U8778 ( .A(n8765), .B(n8766), .Z(Result_33_) );
  XOR2_X1 U8779 ( .A(n8767), .B(n8768), .Z(n8765) );
  XNOR2_X1 U8780 ( .A(n8769), .B(n8770), .ZN(Result_32_) );
  XNOR2_X1 U8781 ( .A(n8771), .B(n8772), .ZN(n8770) );
  XOR2_X1 U8782 ( .A(n8773), .B(n8774), .Z(Result_31_) );
  NOR2_X1 U8783 ( .A1(n8775), .A2(n8776), .ZN(Result_30_) );
  NOR2_X1 U8784 ( .A1(n8777), .A2(n8778), .ZN(n8776) );
  NOR2_X1 U8785 ( .A1(n8773), .A2(n8774), .ZN(n8777) );
  XOR2_X1 U8786 ( .A(n8779), .B(n8780), .Z(Result_2_) );
  XNOR2_X1 U8787 ( .A(n8775), .B(n8781), .ZN(Result_29_) );
  NAND2_X1 U8788 ( .A1(n8782), .A2(n8783), .ZN(n8781) );
  XNOR2_X1 U8789 ( .A(n8784), .B(n8785), .ZN(Result_28_) );
  NAND2_X1 U8790 ( .A1(n8786), .A2(n8787), .ZN(n8784) );
  XNOR2_X1 U8791 ( .A(n8788), .B(n8789), .ZN(Result_27_) );
  NAND2_X1 U8792 ( .A1(n8790), .A2(n8791), .ZN(n8788) );
  XNOR2_X1 U8793 ( .A(n8792), .B(n8793), .ZN(Result_26_) );
  NAND2_X1 U8794 ( .A1(n8794), .A2(n8795), .ZN(n8792) );
  NAND2_X1 U8795 ( .A1(n8796), .A2(n8797), .ZN(n8795) );
  INV_X1 U8796 ( .A(n8798), .ZN(n8796) );
  XNOR2_X1 U8797 ( .A(n8799), .B(n8800), .ZN(Result_25_) );
  NAND2_X1 U8798 ( .A1(n8801), .A2(n8802), .ZN(n8799) );
  XNOR2_X1 U8799 ( .A(n8803), .B(n8804), .ZN(Result_24_) );
  NAND2_X1 U8800 ( .A1(n8805), .A2(n8806), .ZN(n8803) );
  XNOR2_X1 U8801 ( .A(n8807), .B(n8808), .ZN(Result_23_) );
  NAND2_X1 U8802 ( .A1(n8809), .A2(n8810), .ZN(n8807) );
  XNOR2_X1 U8803 ( .A(n8811), .B(n8812), .ZN(Result_22_) );
  NAND2_X1 U8804 ( .A1(n8813), .A2(n8814), .ZN(n8811) );
  XNOR2_X1 U8805 ( .A(n8815), .B(n8816), .ZN(Result_21_) );
  NAND2_X1 U8806 ( .A1(n8817), .A2(n8818), .ZN(n8815) );
  XNOR2_X1 U8807 ( .A(n8819), .B(n8820), .ZN(Result_20_) );
  NAND2_X1 U8808 ( .A1(n8821), .A2(n8822), .ZN(n8819) );
  XNOR2_X1 U8809 ( .A(n8823), .B(n8824), .ZN(Result_1_) );
  NOR2_X1 U8810 ( .A1(n8825), .A2(n8826), .ZN(n8824) );
  INV_X1 U8811 ( .A(n8827), .ZN(n8826) );
  NOR2_X1 U8812 ( .A1(n8828), .A2(n8829), .ZN(n8825) );
  XNOR2_X1 U8813 ( .A(n8830), .B(n8831), .ZN(Result_19_) );
  NAND2_X1 U8814 ( .A1(n8832), .A2(n8833), .ZN(n8830) );
  XNOR2_X1 U8815 ( .A(n8834), .B(n8835), .ZN(Result_18_) );
  NAND2_X1 U8816 ( .A1(n8836), .A2(n8837), .ZN(n8835) );
  XOR2_X1 U8817 ( .A(n8838), .B(n8839), .Z(Result_17_) );
  XOR2_X1 U8818 ( .A(n8840), .B(n8841), .Z(n8839) );
  XNOR2_X1 U8819 ( .A(n8842), .B(n8843), .ZN(Result_16_) );
  NAND2_X1 U8820 ( .A1(n8844), .A2(n8845), .ZN(n8843) );
  XNOR2_X1 U8821 ( .A(n8846), .B(n8847), .ZN(Result_15_) );
  NAND2_X1 U8822 ( .A1(n8848), .A2(n8849), .ZN(n8847) );
  XOR2_X1 U8823 ( .A(n8850), .B(n8851), .Z(Result_14_) );
  XOR2_X1 U8824 ( .A(n8852), .B(n8853), .Z(Result_13_) );
  NOR2_X1 U8825 ( .A1(n8854), .A2(n8855), .ZN(n8853) );
  INV_X1 U8826 ( .A(n8856), .ZN(n8855) );
  NOR2_X1 U8827 ( .A1(n8857), .A2(n8858), .ZN(n8854) );
  XOR2_X1 U8828 ( .A(n8859), .B(n8860), .Z(Result_12_) );
  XOR2_X1 U8829 ( .A(n8861), .B(n8862), .Z(Result_11_) );
  NOR2_X1 U8830 ( .A1(n8863), .A2(n8864), .ZN(n8862) );
  INV_X1 U8831 ( .A(n8865), .ZN(n8864) );
  NOR2_X1 U8832 ( .A1(n8866), .A2(n8867), .ZN(n8863) );
  XOR2_X1 U8833 ( .A(n8868), .B(n8869), .Z(Result_10_) );
  NAND3_X1 U8834 ( .A1(n8870), .A2(n8829), .A3(n8871), .ZN(Result_0_) );
  NAND2_X1 U8835 ( .A1(n8592), .A2(n8828), .ZN(n8871) );
  NAND4_X1 U8836 ( .A1(n8873), .A2(n8592), .A3(n8874), .A4(n8875), .ZN(n8829)
         );
  NAND2_X1 U8837 ( .A1(n8876), .A2(n8827), .ZN(n8870) );
  NAND2_X1 U8838 ( .A1(n8877), .A2(n8878), .ZN(n8827) );
  NAND2_X1 U8839 ( .A1(n8873), .A2(n8875), .ZN(n8878) );
  XOR2_X1 U8840 ( .A(n8828), .B(n8879), .Z(n8877) );
  NAND2_X1 U8841 ( .A1(n8592), .A2(n8874), .ZN(n8879) );
  NAND2_X1 U8842 ( .A1(n8880), .A2(n8881), .ZN(n8828) );
  NAND2_X1 U8843 ( .A1(n8882), .A2(n8883), .ZN(n8881) );
  NAND2_X1 U8844 ( .A1(n8589), .A2(n8885), .ZN(n8882) );
  INV_X1 U8845 ( .A(n8886), .ZN(n8880) );
  INV_X1 U8846 ( .A(n8823), .ZN(n8876) );
  NAND2_X1 U8847 ( .A1(n8779), .A2(n8780), .ZN(n8823) );
  NAND2_X1 U8848 ( .A1(n8887), .A2(n8888), .ZN(n8780) );
  NOR2_X1 U8849 ( .A1(n8734), .A2(n8889), .ZN(n8887) );
  NOR2_X1 U8850 ( .A1(n8732), .A2(n8738), .ZN(n8889) );
  NAND2_X1 U8851 ( .A1(n8690), .A2(n8691), .ZN(n8732) );
  NAND2_X1 U8852 ( .A1(n8890), .A2(n8891), .ZN(n8691) );
  NOR2_X1 U8853 ( .A1(n8643), .A2(n8892), .ZN(n8890) );
  NOR2_X1 U8854 ( .A1(n8641), .A2(n8647), .ZN(n8892) );
  NAND2_X1 U8855 ( .A1(n8617), .A2(n8618), .ZN(n8641) );
  NAND2_X1 U8856 ( .A1(n8893), .A2(n8894), .ZN(n8618) );
  NOR2_X1 U8857 ( .A1(n8610), .A2(n8895), .ZN(n8893) );
  NOR2_X1 U8858 ( .A1(n8608), .A2(n8614), .ZN(n8895) );
  NAND2_X1 U8859 ( .A1(n8606), .A2(n8607), .ZN(n8608) );
  NAND2_X1 U8860 ( .A1(n8896), .A2(n8897), .ZN(n8607) );
  NOR2_X1 U8861 ( .A1(n8599), .A2(n8898), .ZN(n8896) );
  NOR2_X1 U8862 ( .A1(n8899), .A2(n8603), .ZN(n8898) );
  INV_X1 U8863 ( .A(n8597), .ZN(n8899) );
  NOR2_X1 U8864 ( .A1(n8868), .A2(n8869), .ZN(n8597) );
  NOR2_X1 U8865 ( .A1(n8900), .A2(n8901), .ZN(n8869) );
  NAND2_X1 U8866 ( .A1(n8865), .A2(n8902), .ZN(n8901) );
  NAND2_X1 U8867 ( .A1(n8866), .A2(n8861), .ZN(n8902) );
  NOR2_X1 U8868 ( .A1(n8859), .A2(n8860), .ZN(n8861) );
  NOR2_X1 U8869 ( .A1(n8903), .A2(n8904), .ZN(n8860) );
  NAND2_X1 U8870 ( .A1(n8856), .A2(n8905), .ZN(n8904) );
  NAND2_X1 U8871 ( .A1(n8857), .A2(n8852), .ZN(n8905) );
  NOR2_X1 U8872 ( .A1(n8851), .A2(n8850), .ZN(n8852) );
  NOR2_X1 U8873 ( .A1(n8906), .A2(n8907), .ZN(n8850) );
  NAND2_X1 U8874 ( .A1(n8849), .A2(n8908), .ZN(n8907) );
  NAND2_X1 U8875 ( .A1(n8848), .A2(n8846), .ZN(n8908) );
  NAND2_X1 U8876 ( .A1(n8845), .A2(n8909), .ZN(n8846) );
  NAND2_X1 U8877 ( .A1(n8842), .A2(n8844), .ZN(n8909) );
  NAND2_X1 U8878 ( .A1(n8910), .A2(n8911), .ZN(n8844) );
  NOR2_X1 U8879 ( .A1(n8841), .A2(n8912), .ZN(n8842) );
  NOR2_X1 U8880 ( .A1(n8838), .A2(n8913), .ZN(n8912) );
  NAND2_X1 U8881 ( .A1(n8837), .A2(n8914), .ZN(n8838) );
  NAND2_X1 U8882 ( .A1(n8834), .A2(n8836), .ZN(n8914) );
  NAND2_X1 U8883 ( .A1(n8915), .A2(n8916), .ZN(n8836) );
  XNOR2_X1 U8884 ( .A(n8917), .B(n8918), .ZN(n8915) );
  NAND2_X1 U8885 ( .A1(n8833), .A2(n8919), .ZN(n8834) );
  NAND2_X1 U8886 ( .A1(n8831), .A2(n8832), .ZN(n8919) );
  NAND2_X1 U8887 ( .A1(n8920), .A2(n8921), .ZN(n8832) );
  NAND2_X1 U8888 ( .A1(n8922), .A2(n8916), .ZN(n8921) );
  NAND2_X1 U8889 ( .A1(n8923), .A2(n8924), .ZN(n8920) );
  NAND2_X1 U8890 ( .A1(n8822), .A2(n8925), .ZN(n8831) );
  NAND2_X1 U8891 ( .A1(n8820), .A2(n8821), .ZN(n8925) );
  NAND2_X1 U8892 ( .A1(n8926), .A2(n8927), .ZN(n8821) );
  NAND2_X1 U8893 ( .A1(n8928), .A2(n8929), .ZN(n8927) );
  XNOR2_X1 U8894 ( .A(n8924), .B(n8923), .ZN(n8926) );
  NAND2_X1 U8895 ( .A1(n8818), .A2(n8930), .ZN(n8820) );
  NAND2_X1 U8896 ( .A1(n8817), .A2(n8816), .ZN(n8930) );
  NAND2_X1 U8897 ( .A1(n8931), .A2(n8814), .ZN(n8816) );
  NAND2_X1 U8898 ( .A1(n8932), .A2(n8933), .ZN(n8814) );
  INV_X1 U8899 ( .A(n8934), .ZN(n8933) );
  NAND2_X1 U8900 ( .A1(n8812), .A2(n8813), .ZN(n8931) );
  NAND2_X1 U8901 ( .A1(n8934), .A2(n8935), .ZN(n8813) );
  XNOR2_X1 U8902 ( .A(n8936), .B(n8937), .ZN(n8934) );
  NAND2_X1 U8903 ( .A1(n8810), .A2(n8938), .ZN(n8812) );
  NAND2_X1 U8904 ( .A1(n8808), .A2(n8809), .ZN(n8938) );
  NAND2_X1 U8905 ( .A1(n8939), .A2(n8940), .ZN(n8809) );
  NAND2_X1 U8906 ( .A1(n8806), .A2(n8941), .ZN(n8808) );
  NAND2_X1 U8907 ( .A1(n8804), .A2(n8805), .ZN(n8941) );
  NAND2_X1 U8908 ( .A1(n8942), .A2(n8943), .ZN(n8805) );
  XNOR2_X1 U8909 ( .A(n8944), .B(n8945), .ZN(n8942) );
  NAND2_X1 U8910 ( .A1(n8802), .A2(n8946), .ZN(n8804) );
  NAND2_X1 U8911 ( .A1(n8800), .A2(n8801), .ZN(n8946) );
  NAND2_X1 U8912 ( .A1(n8947), .A2(n8948), .ZN(n8801) );
  NAND2_X1 U8913 ( .A1(n8949), .A2(n8943), .ZN(n8948) );
  NAND2_X1 U8914 ( .A1(n8950), .A2(n8951), .ZN(n8947) );
  NAND2_X1 U8915 ( .A1(n8794), .A2(n8952), .ZN(n8800) );
  NAND2_X1 U8916 ( .A1(n8798), .A2(n8793), .ZN(n8952) );
  NAND2_X1 U8917 ( .A1(n8953), .A2(n8790), .ZN(n8793) );
  NAND4_X1 U8918 ( .A1(n8954), .A2(n8955), .A3(n8956), .A4(n8797), .ZN(n8790)
         );
  NAND2_X1 U8919 ( .A1(n8791), .A2(n8789), .ZN(n8953) );
  NAND2_X1 U8920 ( .A1(n8787), .A2(n8957), .ZN(n8789) );
  NAND2_X1 U8921 ( .A1(n8785), .A2(n8786), .ZN(n8957) );
  NAND2_X1 U8922 ( .A1(n8958), .A2(n8959), .ZN(n8786) );
  NAND2_X1 U8923 ( .A1(n8960), .A2(n8961), .ZN(n8959) );
  XNOR2_X1 U8924 ( .A(n8956), .B(n8954), .ZN(n8958) );
  NAND2_X1 U8925 ( .A1(n8783), .A2(n8962), .ZN(n8785) );
  NAND2_X1 U8926 ( .A1(n8775), .A2(n8782), .ZN(n8962) );
  NAND2_X1 U8927 ( .A1(n8963), .A2(n8964), .ZN(n8782) );
  NAND2_X1 U8928 ( .A1(n8965), .A2(n8966), .ZN(n8964) );
  XNOR2_X1 U8929 ( .A(n8961), .B(n8960), .ZN(n8963) );
  NOR3_X1 U8930 ( .A1(n8774), .A2(n8773), .A3(n8967), .ZN(n8775) );
  INV_X1 U8931 ( .A(n8778), .ZN(n8967) );
  XOR2_X1 U8932 ( .A(n8966), .B(n8965), .Z(n8778) );
  NOR2_X1 U8933 ( .A1(n8968), .A2(n8969), .ZN(n8773) );
  INV_X1 U8934 ( .A(n8970), .ZN(n8969) );
  NAND2_X1 U8935 ( .A1(n8771), .A2(n8971), .ZN(n8970) );
  NAND2_X1 U8936 ( .A1(n8772), .A2(n8769), .ZN(n8971) );
  NOR2_X1 U8937 ( .A1(n8619), .A2(n8972), .ZN(n8771) );
  NOR2_X1 U8938 ( .A1(n8769), .A2(n8772), .ZN(n8968) );
  INV_X1 U8939 ( .A(n8973), .ZN(n8772) );
  NAND2_X1 U8940 ( .A1(n8974), .A2(n8975), .ZN(n8973) );
  NAND2_X1 U8941 ( .A1(n8768), .A2(n8976), .ZN(n8975) );
  INV_X1 U8942 ( .A(n8977), .ZN(n8976) );
  NOR2_X1 U8943 ( .A1(n8767), .A2(n8766), .ZN(n8977) );
  NOR2_X1 U8944 ( .A1(n8619), .A2(n8589), .ZN(n8768) );
  NAND2_X1 U8945 ( .A1(n8766), .A2(n8767), .ZN(n8974) );
  NAND2_X1 U8946 ( .A1(n8978), .A2(n8979), .ZN(n8767) );
  NAND2_X1 U8947 ( .A1(n8763), .A2(n8980), .ZN(n8979) );
  INV_X1 U8948 ( .A(n8981), .ZN(n8980) );
  NOR2_X1 U8949 ( .A1(n8764), .A2(n8761), .ZN(n8981) );
  NOR2_X1 U8950 ( .A1(n8619), .A2(n8552), .ZN(n8763) );
  NAND2_X1 U8951 ( .A1(n8761), .A2(n8764), .ZN(n8978) );
  NAND2_X1 U8952 ( .A1(n8983), .A2(n8984), .ZN(n8764) );
  NAND2_X1 U8953 ( .A1(n8760), .A2(n8985), .ZN(n8984) );
  INV_X1 U8954 ( .A(n8986), .ZN(n8985) );
  NOR2_X1 U8955 ( .A1(n8759), .A2(n8758), .ZN(n8986) );
  NOR2_X1 U8956 ( .A1(n8619), .A2(n8527), .ZN(n8760) );
  NAND2_X1 U8957 ( .A1(n8758), .A2(n8759), .ZN(n8983) );
  NAND2_X1 U8958 ( .A1(n8987), .A2(n8988), .ZN(n8759) );
  NAND2_X1 U8959 ( .A1(n8755), .A2(n8989), .ZN(n8988) );
  INV_X1 U8960 ( .A(n8990), .ZN(n8989) );
  NOR2_X1 U8961 ( .A1(n8756), .A2(n8753), .ZN(n8990) );
  NOR2_X1 U8962 ( .A1(n8619), .A2(n8528), .ZN(n8755) );
  NAND2_X1 U8963 ( .A1(n8753), .A2(n8756), .ZN(n8987) );
  NAND2_X1 U8964 ( .A1(n8991), .A2(n8992), .ZN(n8756) );
  NAND2_X1 U8965 ( .A1(n8752), .A2(n8993), .ZN(n8992) );
  INV_X1 U8966 ( .A(n8994), .ZN(n8993) );
  NOR2_X1 U8967 ( .A1(n8751), .A2(n8750), .ZN(n8994) );
  NOR2_X1 U8968 ( .A1(n8619), .A2(n8564), .ZN(n8752) );
  NAND2_X1 U8969 ( .A1(n8750), .A2(n8751), .ZN(n8991) );
  NAND2_X1 U8970 ( .A1(n8996), .A2(n8997), .ZN(n8751) );
  NAND2_X1 U8971 ( .A1(n8748), .A2(n8998), .ZN(n8997) );
  INV_X1 U8972 ( .A(n8999), .ZN(n8998) );
  NOR2_X1 U8973 ( .A1(n8747), .A2(n8745), .ZN(n8999) );
  NOR2_X1 U8974 ( .A1(n8619), .A2(n8555), .ZN(n8748) );
  NAND2_X1 U8975 ( .A1(n8745), .A2(n8747), .ZN(n8996) );
  NAND2_X1 U8976 ( .A1(n9001), .A2(n9002), .ZN(n8747) );
  NAND2_X1 U8977 ( .A1(n8744), .A2(n9003), .ZN(n9002) );
  INV_X1 U8978 ( .A(n9004), .ZN(n9003) );
  NOR2_X1 U8979 ( .A1(n8743), .A2(n8742), .ZN(n9004) );
  NOR2_X1 U8980 ( .A1(n8619), .A2(n8544), .ZN(n8744) );
  NAND2_X1 U8981 ( .A1(n8742), .A2(n8743), .ZN(n9001) );
  NAND2_X1 U8982 ( .A1(n9006), .A2(n9007), .ZN(n8743) );
  NAND2_X1 U8983 ( .A1(n8730), .A2(n9008), .ZN(n9007) );
  INV_X1 U8984 ( .A(n9009), .ZN(n9008) );
  NOR2_X1 U8985 ( .A1(n8731), .A2(n8728), .ZN(n9009) );
  NOR2_X1 U8986 ( .A1(n8619), .A2(n8560), .ZN(n8730) );
  NAND2_X1 U8987 ( .A1(n8728), .A2(n8731), .ZN(n9006) );
  NAND2_X1 U8988 ( .A1(n9011), .A2(n9012), .ZN(n8731) );
  NAND2_X1 U8989 ( .A1(n8727), .A2(n9013), .ZN(n9012) );
  NAND2_X1 U8990 ( .A1(n8726), .A2(n8725), .ZN(n9013) );
  NOR2_X1 U8991 ( .A1(n8619), .A2(n8594), .ZN(n8727) );
  INV_X1 U8992 ( .A(n9015), .ZN(n9011) );
  NOR2_X1 U8993 ( .A1(n8725), .A2(n8726), .ZN(n9015) );
  NOR2_X1 U8994 ( .A1(n9016), .A2(n9017), .ZN(n8726) );
  INV_X1 U8995 ( .A(n9018), .ZN(n9017) );
  NAND2_X1 U8996 ( .A1(n8723), .A2(n9019), .ZN(n9018) );
  NAND2_X1 U8997 ( .A1(n8722), .A2(n8720), .ZN(n9019) );
  NOR2_X1 U8998 ( .A1(n8619), .A2(n8556), .ZN(n8723) );
  NOR2_X1 U8999 ( .A1(n8720), .A2(n8722), .ZN(n9016) );
  NOR2_X1 U9000 ( .A1(n9021), .A2(n9022), .ZN(n8722) );
  INV_X1 U9001 ( .A(n9023), .ZN(n9022) );
  NAND2_X1 U9002 ( .A1(n8718), .A2(n9024), .ZN(n9023) );
  NAND2_X1 U9003 ( .A1(n8719), .A2(n8717), .ZN(n9024) );
  NOR2_X1 U9004 ( .A1(n8619), .A2(n8572), .ZN(n8718) );
  NOR2_X1 U9005 ( .A1(n8717), .A2(n8719), .ZN(n9021) );
  NOR2_X1 U9006 ( .A1(n9026), .A2(n9027), .ZN(n8719) );
  INV_X1 U9007 ( .A(n9028), .ZN(n9027) );
  NAND2_X1 U9008 ( .A1(n8715), .A2(n9029), .ZN(n9028) );
  NAND2_X1 U9009 ( .A1(n9030), .A2(n8712), .ZN(n9029) );
  NOR2_X1 U9010 ( .A1(n8619), .A2(n8582), .ZN(n8715) );
  NOR2_X1 U9011 ( .A1(n8712), .A2(n9030), .ZN(n9026) );
  INV_X1 U9012 ( .A(n8714), .ZN(n9030) );
  NAND2_X1 U9013 ( .A1(n9032), .A2(n9033), .ZN(n8714) );
  NAND2_X1 U9014 ( .A1(n8711), .A2(n9034), .ZN(n9033) );
  INV_X1 U9015 ( .A(n9035), .ZN(n9034) );
  NOR2_X1 U9016 ( .A1(n8710), .A2(n8708), .ZN(n9035) );
  NOR2_X1 U9017 ( .A1(n8619), .A2(n8591), .ZN(n8711) );
  NAND2_X1 U9018 ( .A1(n8708), .A2(n8710), .ZN(n9032) );
  NAND2_X1 U9019 ( .A1(n9037), .A2(n9038), .ZN(n8710) );
  NAND2_X1 U9020 ( .A1(n8707), .A2(n9039), .ZN(n9038) );
  INV_X1 U9021 ( .A(n9040), .ZN(n9039) );
  NOR2_X1 U9022 ( .A1(n8706), .A2(n8704), .ZN(n9040) );
  NOR2_X1 U9023 ( .A1(n8619), .A2(n8562), .ZN(n8707) );
  NAND2_X1 U9024 ( .A1(n8704), .A2(n8706), .ZN(n9037) );
  NAND2_X1 U9025 ( .A1(n9042), .A2(n9043), .ZN(n8706) );
  NAND2_X1 U9026 ( .A1(n8703), .A2(n9044), .ZN(n9043) );
  NAND2_X1 U9027 ( .A1(n9045), .A2(n9046), .ZN(n9044) );
  INV_X1 U9028 ( .A(n8700), .ZN(n9046) );
  INV_X1 U9029 ( .A(n8702), .ZN(n9045) );
  NOR2_X1 U9030 ( .A1(n8619), .A2(n8545), .ZN(n8703) );
  NAND2_X1 U9031 ( .A1(n8700), .A2(n8702), .ZN(n9042) );
  NAND2_X1 U9032 ( .A1(n9047), .A2(n9048), .ZN(n8702) );
  NAND2_X1 U9033 ( .A1(n8699), .A2(n9049), .ZN(n9048) );
  NAND2_X1 U9034 ( .A1(n8698), .A2(n8696), .ZN(n9049) );
  NOR2_X1 U9035 ( .A1(n8619), .A2(n8569), .ZN(n8699) );
  INV_X1 U9036 ( .A(n9051), .ZN(n9047) );
  NOR2_X1 U9037 ( .A1(n8696), .A2(n8698), .ZN(n9051) );
  NOR2_X1 U9038 ( .A1(n9052), .A2(n9053), .ZN(n8698) );
  INV_X1 U9039 ( .A(n9054), .ZN(n9053) );
  NAND2_X1 U9040 ( .A1(n8695), .A2(n9055), .ZN(n9054) );
  NAND2_X1 U9041 ( .A1(n8694), .A2(n8692), .ZN(n9055) );
  NOR2_X1 U9042 ( .A1(n8619), .A2(n8593), .ZN(n8695) );
  NOR2_X1 U9043 ( .A1(n8692), .A2(n8694), .ZN(n9052) );
  NOR2_X1 U9044 ( .A1(n9057), .A2(n9058), .ZN(n8694) );
  INV_X1 U9045 ( .A(n9059), .ZN(n9058) );
  NAND2_X1 U9046 ( .A1(n8689), .A2(n9060), .ZN(n9059) );
  NAND2_X1 U9047 ( .A1(n8687), .A2(n8688), .ZN(n9060) );
  NOR2_X1 U9048 ( .A1(n8619), .A2(n8583), .ZN(n8689) );
  NOR2_X1 U9049 ( .A1(n8688), .A2(n8687), .ZN(n9057) );
  XOR2_X1 U9050 ( .A(n9062), .B(n9063), .Z(n8687) );
  XNOR2_X1 U9051 ( .A(n9064), .B(n9065), .ZN(n9062) );
  NOR2_X1 U9052 ( .A1(n8596), .A2(n8580), .ZN(n9065) );
  NAND2_X1 U9053 ( .A1(n9067), .A2(n9068), .ZN(n8688) );
  NAND2_X1 U9054 ( .A1(n9069), .A2(n8684), .ZN(n9068) );
  NAND2_X1 U9055 ( .A1(n8622), .A2(n9070), .ZN(n8684) );
  NAND2_X1 U9056 ( .A1(n8682), .A2(n8685), .ZN(n9069) );
  INV_X1 U9057 ( .A(n9071), .ZN(n9067) );
  NOR2_X1 U9058 ( .A1(n8685), .A2(n8682), .ZN(n9071) );
  XNOR2_X1 U9059 ( .A(n9072), .B(n9073), .ZN(n8682) );
  XNOR2_X1 U9060 ( .A(n9074), .B(n9075), .ZN(n9072) );
  NOR2_X1 U9061 ( .A1(n8596), .A2(n8588), .ZN(n9075) );
  NAND2_X1 U9062 ( .A1(n8680), .A2(n9077), .ZN(n8685) );
  NAND2_X1 U9063 ( .A1(n8679), .A2(n8681), .ZN(n9077) );
  NAND2_X1 U9064 ( .A1(n9078), .A2(n9079), .ZN(n8681) );
  NAND2_X1 U9065 ( .A1(n8622), .A2(n9080), .ZN(n9078) );
  XNOR2_X1 U9066 ( .A(n9081), .B(n9082), .ZN(n8679) );
  XNOR2_X1 U9067 ( .A(n9083), .B(n9084), .ZN(n9081) );
  NOR2_X1 U9068 ( .A1(n8596), .A2(n8551), .ZN(n9084) );
  INV_X1 U9069 ( .A(n9085), .ZN(n8680) );
  NOR2_X1 U9070 ( .A1(n9079), .A2(n8588), .ZN(n9085) );
  NAND2_X1 U9071 ( .A1(n9086), .A2(n9087), .ZN(n9079) );
  NAND2_X1 U9072 ( .A1(n9088), .A2(n8676), .ZN(n9087) );
  NAND2_X1 U9073 ( .A1(n8622), .A2(n8515), .ZN(n8676) );
  NAND2_X1 U9074 ( .A1(n8674), .A2(n8677), .ZN(n9088) );
  INV_X1 U9075 ( .A(n9089), .ZN(n9086) );
  NOR2_X1 U9076 ( .A1(n8677), .A2(n8674), .ZN(n9089) );
  XNOR2_X1 U9077 ( .A(n9090), .B(n9091), .ZN(n8674) );
  XNOR2_X1 U9078 ( .A(n9092), .B(n9093), .ZN(n9090) );
  NOR2_X1 U9079 ( .A1(n8596), .A2(n8563), .ZN(n9093) );
  NAND2_X1 U9080 ( .A1(n8672), .A2(n9095), .ZN(n8677) );
  NAND2_X1 U9081 ( .A1(n8671), .A2(n8673), .ZN(n9095) );
  NAND2_X1 U9082 ( .A1(n9096), .A2(n9097), .ZN(n8673) );
  NAND2_X1 U9083 ( .A1(n8622), .A2(n9098), .ZN(n9097) );
  XNOR2_X1 U9084 ( .A(n9099), .B(n9100), .ZN(n8671) );
  XNOR2_X1 U9085 ( .A(n9101), .B(n9102), .ZN(n9099) );
  NOR2_X1 U9086 ( .A1(n8596), .A2(n8548), .ZN(n9102) );
  NAND2_X1 U9087 ( .A1(n9098), .A2(n9103), .ZN(n8672) );
  INV_X1 U9088 ( .A(n9096), .ZN(n9103) );
  NOR2_X1 U9089 ( .A1(n9104), .A2(n9105), .ZN(n9096) );
  NOR2_X1 U9090 ( .A1(n8668), .A2(n9106), .ZN(n9105) );
  NOR2_X1 U9091 ( .A1(n8669), .A2(n8666), .ZN(n9106) );
  NAND2_X1 U9092 ( .A1(n8622), .A2(n9107), .ZN(n8668) );
  INV_X1 U9093 ( .A(n9108), .ZN(n9104) );
  NAND2_X1 U9094 ( .A1(n8666), .A2(n8669), .ZN(n9108) );
  NAND2_X1 U9095 ( .A1(n8664), .A2(n9109), .ZN(n8669) );
  NAND2_X1 U9096 ( .A1(n8663), .A2(n8665), .ZN(n9109) );
  NAND2_X1 U9097 ( .A1(n9110), .A2(n9111), .ZN(n8665) );
  NAND2_X1 U9098 ( .A1(n8622), .A2(n9112), .ZN(n9111) );
  XNOR2_X1 U9099 ( .A(n9113), .B(n9114), .ZN(n8663) );
  XNOR2_X1 U9100 ( .A(n9115), .B(n9116), .ZN(n9113) );
  NOR2_X1 U9101 ( .A1(n8596), .A2(n8535), .ZN(n9116) );
  NAND2_X1 U9102 ( .A1(n9112), .A2(n9117), .ZN(n8664) );
  INV_X1 U9103 ( .A(n9110), .ZN(n9117) );
  NOR2_X1 U9104 ( .A1(n9118), .A2(n9119), .ZN(n9110) );
  NOR2_X1 U9105 ( .A1(n8660), .A2(n9120), .ZN(n9119) );
  NOR2_X1 U9106 ( .A1(n8661), .A2(n8659), .ZN(n9120) );
  NAND2_X1 U9107 ( .A1(n8622), .A2(n9121), .ZN(n8660) );
  INV_X1 U9108 ( .A(n9122), .ZN(n9118) );
  NAND2_X1 U9109 ( .A1(n8659), .A2(n8661), .ZN(n9122) );
  NAND2_X1 U9110 ( .A1(n9123), .A2(n9124), .ZN(n8661) );
  NAND2_X1 U9111 ( .A1(n8657), .A2(n9125), .ZN(n9124) );
  NAND2_X1 U9112 ( .A1(n8656), .A2(n8654), .ZN(n9125) );
  NOR2_X1 U9113 ( .A1(n8619), .A2(n8568), .ZN(n8657) );
  NAND2_X1 U9114 ( .A1(n9127), .A2(n9128), .ZN(n9123) );
  INV_X1 U9115 ( .A(n8656), .ZN(n9128) );
  NOR2_X1 U9116 ( .A1(n9129), .A2(n9130), .ZN(n8656) );
  NOR2_X1 U9117 ( .A1(n8652), .A2(n9131), .ZN(n9130) );
  NOR2_X1 U9118 ( .A1(n8653), .A2(n8650), .ZN(n9131) );
  NAND2_X1 U9119 ( .A1(n8622), .A2(n9132), .ZN(n8652) );
  INV_X1 U9120 ( .A(n9133), .ZN(n9129) );
  NAND2_X1 U9121 ( .A1(n8650), .A2(n8653), .ZN(n9133) );
  NAND2_X1 U9122 ( .A1(n8639), .A2(n9134), .ZN(n8653) );
  NAND2_X1 U9123 ( .A1(n8638), .A2(n8640), .ZN(n9134) );
  NAND2_X1 U9124 ( .A1(n9135), .A2(n9136), .ZN(n8640) );
  INV_X1 U9125 ( .A(n9137), .ZN(n9136) );
  NAND2_X1 U9126 ( .A1(n8622), .A2(n9138), .ZN(n9135) );
  XNOR2_X1 U9127 ( .A(n9139), .B(n9140), .ZN(n8638) );
  XNOR2_X1 U9128 ( .A(n9141), .B(n9142), .ZN(n9140) );
  NAND2_X1 U9129 ( .A1(n9137), .A2(n9138), .ZN(n8639) );
  NOR2_X1 U9130 ( .A1(n9143), .A2(n9144), .ZN(n9137) );
  NOR2_X1 U9131 ( .A1(n9145), .A2(n8635), .ZN(n9144) );
  NOR2_X1 U9132 ( .A1(n8619), .A2(n8567), .ZN(n8635) );
  INV_X1 U9133 ( .A(n8622), .ZN(n8619) );
  NOR2_X1 U9134 ( .A1(n8633), .A2(n8636), .ZN(n9145) );
  INV_X1 U9135 ( .A(n9147), .ZN(n8636) );
  NOR2_X1 U9136 ( .A1(n9147), .A2(n9148), .ZN(n9143) );
  INV_X1 U9137 ( .A(n8633), .ZN(n9148) );
  NAND3_X1 U9138 ( .A1(n8537), .A2(n8628), .A3(n8622), .ZN(n8633) );
  NOR2_X1 U9139 ( .A1(n9150), .A2(n9151), .ZN(n8622) );
  NOR2_X1 U9140 ( .A1(d_31_), .A2(c_31_), .ZN(n9150) );
  NAND2_X1 U9141 ( .A1(n9152), .A2(n9153), .ZN(n9147) );
  NAND2_X1 U9142 ( .A1(n8628), .A2(n9154), .ZN(n9153) );
  NAND2_X1 U9143 ( .A1(n8624), .A2(n9155), .ZN(n9154) );
  NAND2_X1 U9144 ( .A1(n8573), .A2(n8585), .ZN(n9155) );
  NAND2_X1 U9145 ( .A1(n9157), .A2(n9158), .ZN(n9152) );
  NAND2_X1 U9146 ( .A1(n8630), .A2(n9159), .ZN(n9158) );
  NAND2_X1 U9147 ( .A1(n8596), .A2(n8539), .ZN(n9159) );
  XNOR2_X1 U9148 ( .A(n9160), .B(n9161), .ZN(n8650) );
  XNOR2_X1 U9149 ( .A(n9162), .B(n9163), .ZN(n9160) );
  INV_X1 U9150 ( .A(n8654), .ZN(n9127) );
  XOR2_X1 U9151 ( .A(n9164), .B(n9165), .Z(n8654) );
  XNOR2_X1 U9152 ( .A(n9166), .B(n9167), .ZN(n9164) );
  XNOR2_X1 U9153 ( .A(n9168), .B(n9169), .ZN(n8659) );
  XNOR2_X1 U9154 ( .A(n9170), .B(n9171), .ZN(n9168) );
  NOR2_X1 U9155 ( .A1(n8596), .A2(n8568), .ZN(n9171) );
  XNOR2_X1 U9156 ( .A(n9172), .B(n9173), .ZN(n8666) );
  XNOR2_X1 U9157 ( .A(n9174), .B(n9175), .ZN(n9172) );
  NOR2_X1 U9158 ( .A1(n8596), .A2(n8584), .ZN(n9175) );
  XOR2_X1 U9159 ( .A(n9177), .B(n9178), .Z(n8692) );
  XNOR2_X1 U9160 ( .A(n9179), .B(n9180), .ZN(n9177) );
  NOR2_X1 U9161 ( .A1(n8596), .A2(n8583), .ZN(n9180) );
  XOR2_X1 U9162 ( .A(n9181), .B(n9182), .Z(n8696) );
  XNOR2_X1 U9163 ( .A(n9183), .B(n9184), .ZN(n9181) );
  NOR2_X1 U9164 ( .A1(n8596), .A2(n8593), .ZN(n9184) );
  XNOR2_X1 U9165 ( .A(n9185), .B(n9186), .ZN(n8700) );
  XNOR2_X1 U9166 ( .A(n9187), .B(n9188), .ZN(n9185) );
  NOR2_X1 U9167 ( .A1(n8596), .A2(n8569), .ZN(n9188) );
  XNOR2_X1 U9168 ( .A(n9189), .B(n9190), .ZN(n8704) );
  XNOR2_X1 U9169 ( .A(n9191), .B(n9192), .ZN(n9189) );
  NOR2_X1 U9170 ( .A1(n8596), .A2(n8545), .ZN(n9192) );
  XNOR2_X1 U9171 ( .A(n9193), .B(n9194), .ZN(n8708) );
  XNOR2_X1 U9172 ( .A(n9195), .B(n9196), .ZN(n9193) );
  NOR2_X1 U9173 ( .A1(n8596), .A2(n8562), .ZN(n9196) );
  XOR2_X1 U9174 ( .A(n9197), .B(n9198), .Z(n8712) );
  XNOR2_X1 U9175 ( .A(n9199), .B(n9200), .ZN(n9197) );
  NOR2_X1 U9176 ( .A1(n8596), .A2(n8591), .ZN(n9200) );
  XOR2_X1 U9177 ( .A(n9201), .B(n9202), .Z(n8717) );
  XNOR2_X1 U9178 ( .A(n9203), .B(n9204), .ZN(n9201) );
  NOR2_X1 U9179 ( .A1(n8596), .A2(n8582), .ZN(n9204) );
  XNOR2_X1 U9180 ( .A(n9205), .B(n9206), .ZN(n8720) );
  XNOR2_X1 U9181 ( .A(n9207), .B(n9208), .ZN(n9206) );
  NAND2_X1 U9182 ( .A1(n9209), .A2(n8628), .ZN(n9208) );
  XOR2_X1 U9183 ( .A(n9210), .B(n9211), .Z(n8725) );
  XNOR2_X1 U9184 ( .A(n9212), .B(n9213), .ZN(n9210) );
  NOR2_X1 U9185 ( .A1(n8596), .A2(n8556), .ZN(n9213) );
  XNOR2_X1 U9186 ( .A(n9214), .B(n9215), .ZN(n8728) );
  XNOR2_X1 U9187 ( .A(n9216), .B(n9217), .ZN(n9214) );
  NOR2_X1 U9188 ( .A1(n8595), .A2(n8594), .ZN(n9217) );
  XNOR2_X1 U9189 ( .A(n9218), .B(n9219), .ZN(n8742) );
  XNOR2_X1 U9190 ( .A(n9220), .B(n9221), .ZN(n9218) );
  NOR2_X1 U9191 ( .A1(n8595), .A2(n8560), .ZN(n9221) );
  XNOR2_X1 U9192 ( .A(n9222), .B(n9223), .ZN(n8745) );
  XNOR2_X1 U9193 ( .A(n9224), .B(n9225), .ZN(n9222) );
  NOR2_X1 U9194 ( .A1(n8595), .A2(n8544), .ZN(n9225) );
  XNOR2_X1 U9195 ( .A(n9226), .B(n9227), .ZN(n8750) );
  XNOR2_X1 U9196 ( .A(n9228), .B(n9229), .ZN(n9226) );
  NOR2_X1 U9197 ( .A1(n8595), .A2(n8555), .ZN(n9229) );
  XNOR2_X1 U9198 ( .A(n9230), .B(n9231), .ZN(n8753) );
  XNOR2_X1 U9199 ( .A(n9232), .B(n9233), .ZN(n9230) );
  NOR2_X1 U9200 ( .A1(n8595), .A2(n8564), .ZN(n9233) );
  XNOR2_X1 U9201 ( .A(n9234), .B(n9235), .ZN(n8758) );
  XNOR2_X1 U9202 ( .A(n9236), .B(n9237), .ZN(n9234) );
  NOR2_X1 U9203 ( .A1(n8595), .A2(n8528), .ZN(n9237) );
  XNOR2_X1 U9204 ( .A(n9238), .B(n9239), .ZN(n8761) );
  XNOR2_X1 U9205 ( .A(n9240), .B(n9241), .ZN(n9238) );
  NOR2_X1 U9206 ( .A1(n8595), .A2(n8527), .ZN(n9241) );
  XNOR2_X1 U9207 ( .A(n9242), .B(n9243), .ZN(n8766) );
  XNOR2_X1 U9208 ( .A(n9244), .B(n9245), .ZN(n9242) );
  NOR2_X1 U9209 ( .A1(n8595), .A2(n8552), .ZN(n9245) );
  XOR2_X1 U9210 ( .A(n9246), .B(n9247), .Z(n8769) );
  XNOR2_X1 U9211 ( .A(n9248), .B(n9249), .ZN(n9246) );
  NOR2_X1 U9212 ( .A1(n8595), .A2(n8589), .ZN(n9249) );
  XNOR2_X1 U9213 ( .A(n9250), .B(n9251), .ZN(n8774) );
  XNOR2_X1 U9214 ( .A(n9252), .B(n9253), .ZN(n9251) );
  NAND2_X1 U9215 ( .A1(n8628), .A2(n8592), .ZN(n9253) );
  NAND3_X1 U9216 ( .A1(n8965), .A2(n8966), .A3(n9254), .ZN(n8783) );
  XOR2_X1 U9217 ( .A(n8961), .B(n8960), .Z(n9254) );
  NAND2_X1 U9218 ( .A1(n9255), .A2(n9256), .ZN(n8966) );
  NAND3_X1 U9219 ( .A1(n8592), .A2(n9257), .A3(n8628), .ZN(n9256) );
  NAND2_X1 U9220 ( .A1(n9252), .A2(n9250), .ZN(n9257) );
  INV_X1 U9221 ( .A(n9258), .ZN(n9255) );
  NOR2_X1 U9222 ( .A1(n9250), .A2(n9252), .ZN(n9258) );
  NOR2_X1 U9223 ( .A1(n9259), .A2(n9260), .ZN(n9252) );
  INV_X1 U9224 ( .A(n9261), .ZN(n9260) );
  NAND3_X1 U9225 ( .A1(n8628), .A2(n9262), .A3(n9263), .ZN(n9261) );
  NAND2_X1 U9226 ( .A1(n9247), .A2(n9248), .ZN(n9262) );
  NOR2_X1 U9227 ( .A1(n9247), .A2(n9248), .ZN(n9259) );
  NOR2_X1 U9228 ( .A1(n9264), .A2(n9265), .ZN(n9248) );
  INV_X1 U9229 ( .A(n9266), .ZN(n9265) );
  NAND3_X1 U9230 ( .A1(n8628), .A2(n9267), .A3(n9268), .ZN(n9266) );
  NAND2_X1 U9231 ( .A1(n9244), .A2(n9243), .ZN(n9267) );
  NOR2_X1 U9232 ( .A1(n9243), .A2(n9244), .ZN(n9264) );
  NOR2_X1 U9233 ( .A1(n9269), .A2(n9270), .ZN(n9244) );
  NOR3_X1 U9234 ( .A1(n8595), .A2(n9271), .A3(n8527), .ZN(n9270) );
  INV_X1 U9235 ( .A(n9272), .ZN(n9271) );
  NAND2_X1 U9236 ( .A1(n9239), .A2(n9240), .ZN(n9272) );
  NOR2_X1 U9237 ( .A1(n9239), .A2(n9240), .ZN(n9269) );
  NOR2_X1 U9238 ( .A1(n9273), .A2(n9274), .ZN(n9240) );
  INV_X1 U9239 ( .A(n9275), .ZN(n9274) );
  NAND3_X1 U9240 ( .A1(n8628), .A2(n9276), .A3(n9277), .ZN(n9275) );
  NAND2_X1 U9241 ( .A1(n9236), .A2(n9235), .ZN(n9276) );
  NOR2_X1 U9242 ( .A1(n9235), .A2(n9236), .ZN(n9273) );
  NOR2_X1 U9243 ( .A1(n9278), .A2(n9279), .ZN(n9236) );
  NOR3_X1 U9244 ( .A1(n8595), .A2(n9280), .A3(n8564), .ZN(n9279) );
  INV_X1 U9245 ( .A(n9281), .ZN(n9280) );
  NAND2_X1 U9246 ( .A1(n9231), .A2(n9232), .ZN(n9281) );
  NOR2_X1 U9247 ( .A1(n9231), .A2(n9232), .ZN(n9278) );
  NOR2_X1 U9248 ( .A1(n9282), .A2(n9283), .ZN(n9232) );
  INV_X1 U9249 ( .A(n9284), .ZN(n9283) );
  NAND3_X1 U9250 ( .A1(n8628), .A2(n9285), .A3(n9286), .ZN(n9284) );
  NAND2_X1 U9251 ( .A1(n9228), .A2(n9227), .ZN(n9285) );
  NOR2_X1 U9252 ( .A1(n9227), .A2(n9228), .ZN(n9282) );
  NOR2_X1 U9253 ( .A1(n9287), .A2(n9288), .ZN(n9228) );
  NOR3_X1 U9254 ( .A1(n8595), .A2(n9289), .A3(n8544), .ZN(n9288) );
  INV_X1 U9255 ( .A(n9290), .ZN(n9289) );
  NAND2_X1 U9256 ( .A1(n9223), .A2(n9224), .ZN(n9290) );
  NOR2_X1 U9257 ( .A1(n9223), .A2(n9224), .ZN(n9287) );
  NOR2_X1 U9258 ( .A1(n9291), .A2(n9292), .ZN(n9224) );
  INV_X1 U9259 ( .A(n9293), .ZN(n9292) );
  NAND3_X1 U9260 ( .A1(n8628), .A2(n9294), .A3(n9295), .ZN(n9293) );
  NAND2_X1 U9261 ( .A1(n9220), .A2(n9219), .ZN(n9294) );
  NOR2_X1 U9262 ( .A1(n9219), .A2(n9220), .ZN(n9291) );
  NOR2_X1 U9263 ( .A1(n9296), .A2(n9297), .ZN(n9220) );
  NOR3_X1 U9264 ( .A1(n8595), .A2(n9298), .A3(n8594), .ZN(n9297) );
  INV_X1 U9265 ( .A(n9299), .ZN(n9298) );
  NAND2_X1 U9266 ( .A1(n9215), .A2(n9216), .ZN(n9299) );
  NOR2_X1 U9267 ( .A1(n9215), .A2(n9216), .ZN(n9296) );
  NOR2_X1 U9268 ( .A1(n9300), .A2(n9301), .ZN(n9216) );
  INV_X1 U9269 ( .A(n9302), .ZN(n9301) );
  NAND3_X1 U9270 ( .A1(n8628), .A2(n9303), .A3(n9304), .ZN(n9302) );
  NAND2_X1 U9271 ( .A1(n9212), .A2(n9211), .ZN(n9303) );
  NOR2_X1 U9272 ( .A1(n9211), .A2(n9212), .ZN(n9300) );
  NOR2_X1 U9273 ( .A1(n9305), .A2(n9306), .ZN(n9212) );
  NOR3_X1 U9274 ( .A1(n8595), .A2(n9307), .A3(n8572), .ZN(n9306) );
  INV_X1 U9275 ( .A(n9308), .ZN(n9307) );
  NAND2_X1 U9276 ( .A1(n9205), .A2(n9207), .ZN(n9308) );
  NOR2_X1 U9277 ( .A1(n9205), .A2(n9207), .ZN(n9305) );
  NOR2_X1 U9278 ( .A1(n9309), .A2(n9310), .ZN(n9207) );
  INV_X1 U9279 ( .A(n9311), .ZN(n9310) );
  NAND3_X1 U9280 ( .A1(n8628), .A2(n9312), .A3(n9313), .ZN(n9311) );
  NAND2_X1 U9281 ( .A1(n9203), .A2(n9202), .ZN(n9312) );
  NOR2_X1 U9282 ( .A1(n9202), .A2(n9203), .ZN(n9309) );
  NOR2_X1 U9283 ( .A1(n9314), .A2(n9315), .ZN(n9203) );
  NOR3_X1 U9284 ( .A1(n8595), .A2(n9316), .A3(n8591), .ZN(n9315) );
  INV_X1 U9285 ( .A(n9317), .ZN(n9316) );
  NAND2_X1 U9286 ( .A1(n9198), .A2(n9199), .ZN(n9317) );
  NOR2_X1 U9287 ( .A1(n9198), .A2(n9199), .ZN(n9314) );
  NOR2_X1 U9288 ( .A1(n9318), .A2(n9319), .ZN(n9199) );
  INV_X1 U9289 ( .A(n9320), .ZN(n9319) );
  NAND3_X1 U9290 ( .A1(n8628), .A2(n9321), .A3(n9322), .ZN(n9320) );
  NAND2_X1 U9291 ( .A1(n9195), .A2(n9194), .ZN(n9321) );
  NOR2_X1 U9292 ( .A1(n9194), .A2(n9195), .ZN(n9318) );
  NOR2_X1 U9293 ( .A1(n9323), .A2(n9324), .ZN(n9195) );
  NOR3_X1 U9294 ( .A1(n8595), .A2(n9325), .A3(n8545), .ZN(n9324) );
  INV_X1 U9295 ( .A(n9326), .ZN(n9325) );
  NAND2_X1 U9296 ( .A1(n9190), .A2(n9191), .ZN(n9326) );
  NOR2_X1 U9297 ( .A1(n9190), .A2(n9191), .ZN(n9323) );
  NOR2_X1 U9298 ( .A1(n9327), .A2(n9328), .ZN(n9191) );
  INV_X1 U9299 ( .A(n9329), .ZN(n9328) );
  NAND3_X1 U9300 ( .A1(n8628), .A2(n9330), .A3(n9331), .ZN(n9329) );
  NAND2_X1 U9301 ( .A1(n9187), .A2(n9186), .ZN(n9330) );
  NOR2_X1 U9302 ( .A1(n9186), .A2(n9187), .ZN(n9327) );
  NOR2_X1 U9303 ( .A1(n9332), .A2(n9333), .ZN(n9187) );
  NOR3_X1 U9304 ( .A1(n8595), .A2(n9334), .A3(n8593), .ZN(n9333) );
  INV_X1 U9305 ( .A(n9335), .ZN(n9334) );
  NAND2_X1 U9306 ( .A1(n9182), .A2(n9183), .ZN(n9335) );
  NOR2_X1 U9307 ( .A1(n9182), .A2(n9183), .ZN(n9332) );
  NOR2_X1 U9308 ( .A1(n9336), .A2(n9337), .ZN(n9183) );
  INV_X1 U9309 ( .A(n9338), .ZN(n9337) );
  NAND3_X1 U9310 ( .A1(n8628), .A2(n9339), .A3(n9340), .ZN(n9338) );
  NAND2_X1 U9311 ( .A1(n9179), .A2(n9178), .ZN(n9339) );
  NOR2_X1 U9312 ( .A1(n9178), .A2(n9179), .ZN(n9336) );
  NOR2_X1 U9313 ( .A1(n9341), .A2(n9342), .ZN(n9179) );
  NOR3_X1 U9314 ( .A1(n8595), .A2(n9343), .A3(n8580), .ZN(n9342) );
  INV_X1 U9315 ( .A(n9344), .ZN(n9343) );
  NAND2_X1 U9316 ( .A1(n9063), .A2(n9064), .ZN(n9344) );
  NOR2_X1 U9317 ( .A1(n9063), .A2(n9064), .ZN(n9341) );
  NOR2_X1 U9318 ( .A1(n9345), .A2(n9346), .ZN(n9064) );
  INV_X1 U9319 ( .A(n9347), .ZN(n9346) );
  NAND3_X1 U9320 ( .A1(n8628), .A2(n9348), .A3(n9080), .ZN(n9347) );
  NAND2_X1 U9321 ( .A1(n9074), .A2(n9073), .ZN(n9348) );
  NOR2_X1 U9322 ( .A1(n9073), .A2(n9074), .ZN(n9345) );
  NOR2_X1 U9323 ( .A1(n9349), .A2(n9350), .ZN(n9074) );
  NOR3_X1 U9324 ( .A1(n8595), .A2(n9351), .A3(n8551), .ZN(n9350) );
  INV_X1 U9325 ( .A(n9352), .ZN(n9351) );
  NAND2_X1 U9326 ( .A1(n9082), .A2(n9083), .ZN(n9352) );
  NOR2_X1 U9327 ( .A1(n9082), .A2(n9083), .ZN(n9349) );
  NOR2_X1 U9328 ( .A1(n9353), .A2(n9354), .ZN(n9083) );
  INV_X1 U9329 ( .A(n9355), .ZN(n9354) );
  NAND3_X1 U9330 ( .A1(n8628), .A2(n9356), .A3(n9098), .ZN(n9355) );
  NAND2_X1 U9331 ( .A1(n9092), .A2(n9091), .ZN(n9356) );
  NOR2_X1 U9332 ( .A1(n9091), .A2(n9092), .ZN(n9353) );
  NOR2_X1 U9333 ( .A1(n9357), .A2(n9358), .ZN(n9092) );
  NOR3_X1 U9334 ( .A1(n8595), .A2(n9359), .A3(n8548), .ZN(n9358) );
  INV_X1 U9335 ( .A(n9360), .ZN(n9359) );
  NAND2_X1 U9336 ( .A1(n9100), .A2(n9101), .ZN(n9360) );
  NOR2_X1 U9337 ( .A1(n9100), .A2(n9101), .ZN(n9357) );
  NOR2_X1 U9338 ( .A1(n9361), .A2(n9362), .ZN(n9101) );
  INV_X1 U9339 ( .A(n9363), .ZN(n9362) );
  NAND3_X1 U9340 ( .A1(n8628), .A2(n9364), .A3(n9112), .ZN(n9363) );
  NAND2_X1 U9341 ( .A1(n9174), .A2(n9173), .ZN(n9364) );
  NOR2_X1 U9342 ( .A1(n9173), .A2(n9174), .ZN(n9361) );
  NOR2_X1 U9343 ( .A1(n9365), .A2(n9366), .ZN(n9174) );
  NOR3_X1 U9344 ( .A1(n8595), .A2(n9367), .A3(n8535), .ZN(n9366) );
  INV_X1 U9345 ( .A(n9368), .ZN(n9367) );
  NAND2_X1 U9346 ( .A1(n9114), .A2(n9115), .ZN(n9368) );
  NOR2_X1 U9347 ( .A1(n9114), .A2(n9115), .ZN(n9365) );
  NOR2_X1 U9348 ( .A1(n9369), .A2(n9370), .ZN(n9115) );
  INV_X1 U9349 ( .A(n9371), .ZN(n9370) );
  NAND3_X1 U9350 ( .A1(n8628), .A2(n9372), .A3(n9373), .ZN(n9371) );
  NAND2_X1 U9351 ( .A1(n9170), .A2(n9169), .ZN(n9372) );
  NOR2_X1 U9352 ( .A1(n9169), .A2(n9170), .ZN(n9369) );
  NOR2_X1 U9353 ( .A1(n9374), .A2(n9375), .ZN(n9170) );
  INV_X1 U9354 ( .A(n9376), .ZN(n9375) );
  NAND2_X1 U9355 ( .A1(n9166), .A2(n9377), .ZN(n9376) );
  NAND2_X1 U9356 ( .A1(n9165), .A2(n9167), .ZN(n9377) );
  NOR2_X1 U9357 ( .A1(n9378), .A2(n8596), .ZN(n9166) );
  NOR2_X1 U9358 ( .A1(n9165), .A2(n9167), .ZN(n9374) );
  NOR2_X1 U9359 ( .A1(n9379), .A2(n9380), .ZN(n9167) );
  INV_X1 U9360 ( .A(n9381), .ZN(n9380) );
  NAND2_X1 U9361 ( .A1(n9162), .A2(n9382), .ZN(n9381) );
  NAND2_X1 U9362 ( .A1(n9163), .A2(n9161), .ZN(n9382) );
  NOR2_X1 U9363 ( .A1(n9383), .A2(n8596), .ZN(n9162) );
  NOR2_X1 U9364 ( .A1(n9161), .A2(n9163), .ZN(n9379) );
  NOR2_X1 U9365 ( .A1(n9384), .A2(n9385), .ZN(n9163) );
  INV_X1 U9366 ( .A(n9386), .ZN(n9385) );
  NAND2_X1 U9367 ( .A1(n9139), .A2(n9387), .ZN(n9386) );
  NAND2_X1 U9368 ( .A1(n9142), .A2(n9141), .ZN(n9387) );
  NOR2_X1 U9369 ( .A1(n9146), .A2(n8596), .ZN(n9139) );
  NOR2_X1 U9370 ( .A1(n9141), .A2(n9142), .ZN(n9384) );
  INV_X1 U9371 ( .A(n9388), .ZN(n9142) );
  NAND2_X1 U9372 ( .A1(n9389), .A2(n9390), .ZN(n9388) );
  NAND2_X1 U9373 ( .A1(n9157), .A2(n9391), .ZN(n9390) );
  NAND2_X1 U9374 ( .A1(n8624), .A2(n9392), .ZN(n9391) );
  NAND2_X1 U9375 ( .A1(n8550), .A2(n8585), .ZN(n9392) );
  NAND2_X1 U9376 ( .A1(n8549), .A2(n9394), .ZN(n9389) );
  NAND2_X1 U9377 ( .A1(n8630), .A2(n9395), .ZN(n9394) );
  NAND2_X1 U9378 ( .A1(n8539), .A2(n8573), .ZN(n9395) );
  NAND3_X1 U9379 ( .A1(n8537), .A2(n8628), .A3(n9157), .ZN(n9141) );
  INV_X1 U9380 ( .A(n8596), .ZN(n8628) );
  XOR2_X1 U9381 ( .A(n9398), .B(n9399), .Z(n9161) );
  XNOR2_X1 U9382 ( .A(n9400), .B(n9401), .ZN(n9399) );
  XOR2_X1 U9383 ( .A(n9402), .B(n9403), .Z(n9165) );
  XNOR2_X1 U9384 ( .A(n9404), .B(n9405), .ZN(n9402) );
  XOR2_X1 U9385 ( .A(n9406), .B(n9407), .Z(n9169) );
  XNOR2_X1 U9386 ( .A(n9408), .B(n9409), .ZN(n9406) );
  XOR2_X1 U9387 ( .A(n9410), .B(n9411), .Z(n9114) );
  XNOR2_X1 U9388 ( .A(n9412), .B(n9413), .ZN(n9410) );
  XOR2_X1 U9389 ( .A(n9414), .B(n9415), .Z(n9173) );
  XNOR2_X1 U9390 ( .A(n9416), .B(n9417), .ZN(n9414) );
  XOR2_X1 U9391 ( .A(n9418), .B(n9419), .Z(n9100) );
  XNOR2_X1 U9392 ( .A(n9420), .B(n9421), .ZN(n9418) );
  XNOR2_X1 U9393 ( .A(n9422), .B(n9423), .ZN(n9091) );
  XOR2_X1 U9394 ( .A(n9424), .B(n9425), .Z(n9423) );
  XOR2_X1 U9395 ( .A(n9426), .B(n9427), .Z(n9082) );
  XNOR2_X1 U9396 ( .A(n9428), .B(n9429), .ZN(n9426) );
  XNOR2_X1 U9397 ( .A(n9430), .B(n9431), .ZN(n9073) );
  XOR2_X1 U9398 ( .A(n9432), .B(n9433), .Z(n9431) );
  XOR2_X1 U9399 ( .A(n9434), .B(n9435), .Z(n9063) );
  XNOR2_X1 U9400 ( .A(n9436), .B(n9437), .ZN(n9434) );
  XNOR2_X1 U9401 ( .A(n9438), .B(n9439), .ZN(n9178) );
  XOR2_X1 U9402 ( .A(n9440), .B(n9441), .Z(n9439) );
  XOR2_X1 U9403 ( .A(n9442), .B(n9443), .Z(n9182) );
  XNOR2_X1 U9404 ( .A(n9444), .B(n9445), .ZN(n9442) );
  XNOR2_X1 U9405 ( .A(n9446), .B(n9447), .ZN(n9186) );
  XOR2_X1 U9406 ( .A(n9448), .B(n9449), .Z(n9447) );
  XOR2_X1 U9407 ( .A(n9450), .B(n9451), .Z(n9190) );
  XNOR2_X1 U9408 ( .A(n9452), .B(n9453), .ZN(n9450) );
  XOR2_X1 U9409 ( .A(n9454), .B(n9455), .Z(n9194) );
  XNOR2_X1 U9410 ( .A(n9456), .B(n9457), .ZN(n9454) );
  XOR2_X1 U9411 ( .A(n9458), .B(n9459), .Z(n9198) );
  XNOR2_X1 U9412 ( .A(n9460), .B(n9461), .ZN(n9458) );
  XOR2_X1 U9413 ( .A(n9462), .B(n9463), .Z(n9202) );
  XNOR2_X1 U9414 ( .A(n9464), .B(n9465), .ZN(n9462) );
  XOR2_X1 U9415 ( .A(n9466), .B(n9467), .Z(n9205) );
  XNOR2_X1 U9416 ( .A(n9468), .B(n9469), .ZN(n9466) );
  XOR2_X1 U9417 ( .A(n9470), .B(n9471), .Z(n9211) );
  XNOR2_X1 U9418 ( .A(n9472), .B(n9473), .ZN(n9470) );
  XNOR2_X1 U9419 ( .A(n9474), .B(n9475), .ZN(n9215) );
  XOR2_X1 U9420 ( .A(n9476), .B(n9477), .Z(n9475) );
  XNOR2_X1 U9421 ( .A(n9478), .B(n9479), .ZN(n9219) );
  XOR2_X1 U9422 ( .A(n9480), .B(n9481), .Z(n9478) );
  XNOR2_X1 U9423 ( .A(n9482), .B(n9483), .ZN(n9223) );
  XOR2_X1 U9424 ( .A(n9484), .B(n9485), .Z(n9482) );
  XOR2_X1 U9425 ( .A(n9486), .B(n9487), .Z(n9227) );
  XNOR2_X1 U9426 ( .A(n9488), .B(n9489), .ZN(n9486) );
  XNOR2_X1 U9427 ( .A(n9490), .B(n9491), .ZN(n9231) );
  XOR2_X1 U9428 ( .A(n9492), .B(n9493), .Z(n9491) );
  XNOR2_X1 U9429 ( .A(n9494), .B(n9495), .ZN(n9235) );
  XOR2_X1 U9430 ( .A(n9496), .B(n9497), .Z(n9494) );
  XOR2_X1 U9431 ( .A(n9498), .B(n9499), .Z(n9239) );
  XNOR2_X1 U9432 ( .A(n9500), .B(n9501), .ZN(n9499) );
  XNOR2_X1 U9433 ( .A(n9502), .B(n9503), .ZN(n9243) );
  XOR2_X1 U9434 ( .A(n9504), .B(n9505), .Z(n9502) );
  NOR2_X1 U9435 ( .A1(n8527), .A2(n8573), .ZN(n9505) );
  XNOR2_X1 U9436 ( .A(n9506), .B(n9507), .ZN(n9247) );
  XOR2_X1 U9437 ( .A(n9508), .B(n9509), .Z(n9507) );
  XOR2_X1 U9438 ( .A(n9510), .B(n9511), .Z(n9250) );
  XNOR2_X1 U9439 ( .A(n9512), .B(n9513), .ZN(n9510) );
  XNOR2_X1 U9440 ( .A(n9514), .B(n9515), .ZN(n8965) );
  NAND2_X1 U9441 ( .A1(n9516), .A2(n9517), .ZN(n9514) );
  NAND3_X1 U9442 ( .A1(n8960), .A2(n8961), .A3(n9518), .ZN(n8787) );
  XOR2_X1 U9443 ( .A(n8956), .B(n8954), .Z(n9518) );
  NAND2_X1 U9444 ( .A1(n9516), .A2(n9519), .ZN(n8961) );
  NAND2_X1 U9445 ( .A1(n9515), .A2(n9517), .ZN(n9519) );
  NAND2_X1 U9446 ( .A1(n9520), .A2(n9521), .ZN(n9517) );
  NAND2_X1 U9447 ( .A1(n9157), .A2(n8592), .ZN(n9521) );
  XOR2_X1 U9448 ( .A(n9522), .B(n9523), .Z(n9515) );
  XOR2_X1 U9449 ( .A(n9524), .B(n9525), .Z(n9522) );
  NAND2_X1 U9450 ( .A1(n8592), .A2(n9526), .ZN(n9516) );
  INV_X1 U9451 ( .A(n9520), .ZN(n9526) );
  NOR2_X1 U9452 ( .A1(n9527), .A2(n9528), .ZN(n9520) );
  INV_X1 U9453 ( .A(n9529), .ZN(n9528) );
  NAND2_X1 U9454 ( .A1(n9513), .A2(n9530), .ZN(n9529) );
  NAND2_X1 U9455 ( .A1(n9512), .A2(n9511), .ZN(n9530) );
  NOR2_X1 U9456 ( .A1(n8573), .A2(n8589), .ZN(n9513) );
  NOR2_X1 U9457 ( .A1(n9511), .A2(n9512), .ZN(n9527) );
  NOR2_X1 U9458 ( .A1(n9531), .A2(n9532), .ZN(n9512) );
  INV_X1 U9459 ( .A(n9533), .ZN(n9532) );
  NAND2_X1 U9460 ( .A1(n9508), .A2(n9534), .ZN(n9533) );
  NAND2_X1 U9461 ( .A1(n9506), .A2(n9509), .ZN(n9534) );
  NAND2_X1 U9462 ( .A1(n9535), .A2(n9536), .ZN(n9508) );
  INV_X1 U9463 ( .A(n9537), .ZN(n9536) );
  NOR3_X1 U9464 ( .A1(n8527), .A2(n9538), .A3(n8573), .ZN(n9537) );
  NOR2_X1 U9465 ( .A1(n9504), .A2(n9503), .ZN(n9538) );
  NAND2_X1 U9466 ( .A1(n9503), .A2(n9504), .ZN(n9535) );
  NAND2_X1 U9467 ( .A1(n9539), .A2(n9540), .ZN(n9504) );
  NAND2_X1 U9468 ( .A1(n9501), .A2(n9541), .ZN(n9540) );
  INV_X1 U9469 ( .A(n9542), .ZN(n9541) );
  NOR2_X1 U9470 ( .A1(n9500), .A2(n9498), .ZN(n9542) );
  NOR2_X1 U9471 ( .A1(n8573), .A2(n8528), .ZN(n9501) );
  NAND2_X1 U9472 ( .A1(n9498), .A2(n9500), .ZN(n9539) );
  NAND2_X1 U9473 ( .A1(n9543), .A2(n9544), .ZN(n9500) );
  NAND2_X1 U9474 ( .A1(n9497), .A2(n9545), .ZN(n9544) );
  INV_X1 U9475 ( .A(n9546), .ZN(n9545) );
  NOR2_X1 U9476 ( .A1(n9496), .A2(n9495), .ZN(n9546) );
  NOR2_X1 U9477 ( .A1(n8573), .A2(n8564), .ZN(n9497) );
  NAND2_X1 U9478 ( .A1(n9495), .A2(n9496), .ZN(n9543) );
  NAND2_X1 U9479 ( .A1(n9547), .A2(n9548), .ZN(n9496) );
  NAND2_X1 U9480 ( .A1(n9493), .A2(n9549), .ZN(n9548) );
  NAND2_X1 U9481 ( .A1(n9492), .A2(n9490), .ZN(n9549) );
  NOR2_X1 U9482 ( .A1(n8573), .A2(n8555), .ZN(n9493) );
  INV_X1 U9483 ( .A(n9550), .ZN(n9547) );
  NOR2_X1 U9484 ( .A1(n9490), .A2(n9492), .ZN(n9550) );
  NOR2_X1 U9485 ( .A1(n9551), .A2(n9552), .ZN(n9492) );
  INV_X1 U9486 ( .A(n9553), .ZN(n9552) );
  NAND2_X1 U9487 ( .A1(n9489), .A2(n9554), .ZN(n9553) );
  NAND2_X1 U9488 ( .A1(n9488), .A2(n9487), .ZN(n9554) );
  NOR2_X1 U9489 ( .A1(n8573), .A2(n8544), .ZN(n9489) );
  NOR2_X1 U9490 ( .A1(n9487), .A2(n9488), .ZN(n9551) );
  INV_X1 U9491 ( .A(n9555), .ZN(n9488) );
  NAND2_X1 U9492 ( .A1(n9556), .A2(n9557), .ZN(n9555) );
  NAND2_X1 U9493 ( .A1(n9484), .A2(n9558), .ZN(n9557) );
  INV_X1 U9494 ( .A(n9559), .ZN(n9558) );
  NOR2_X1 U9495 ( .A1(n9485), .A2(n9483), .ZN(n9559) );
  NOR2_X1 U9496 ( .A1(n8573), .A2(n8560), .ZN(n9484) );
  NAND2_X1 U9497 ( .A1(n9483), .A2(n9485), .ZN(n9556) );
  NAND2_X1 U9498 ( .A1(n9560), .A2(n9561), .ZN(n9485) );
  NAND2_X1 U9499 ( .A1(n9481), .A2(n9562), .ZN(n9561) );
  INV_X1 U9500 ( .A(n9563), .ZN(n9562) );
  NOR2_X1 U9501 ( .A1(n9480), .A2(n9479), .ZN(n9563) );
  NOR2_X1 U9502 ( .A1(n8573), .A2(n8594), .ZN(n9481) );
  NAND2_X1 U9503 ( .A1(n9479), .A2(n9480), .ZN(n9560) );
  NAND2_X1 U9504 ( .A1(n9564), .A2(n9565), .ZN(n9480) );
  NAND2_X1 U9505 ( .A1(n9477), .A2(n9566), .ZN(n9565) );
  NAND2_X1 U9506 ( .A1(n9476), .A2(n9474), .ZN(n9566) );
  NOR2_X1 U9507 ( .A1(n8573), .A2(n8556), .ZN(n9477) );
  INV_X1 U9508 ( .A(n9567), .ZN(n9564) );
  NOR2_X1 U9509 ( .A1(n9474), .A2(n9476), .ZN(n9567) );
  NOR2_X1 U9510 ( .A1(n9568), .A2(n9569), .ZN(n9476) );
  INV_X1 U9511 ( .A(n9570), .ZN(n9569) );
  NAND2_X1 U9512 ( .A1(n9473), .A2(n9571), .ZN(n9570) );
  NAND2_X1 U9513 ( .A1(n9472), .A2(n9471), .ZN(n9571) );
  NOR2_X1 U9514 ( .A1(n8573), .A2(n8572), .ZN(n9473) );
  NOR2_X1 U9515 ( .A1(n9471), .A2(n9472), .ZN(n9568) );
  NOR2_X1 U9516 ( .A1(n9572), .A2(n9573), .ZN(n9472) );
  INV_X1 U9517 ( .A(n9574), .ZN(n9573) );
  NAND2_X1 U9518 ( .A1(n9469), .A2(n9575), .ZN(n9574) );
  NAND2_X1 U9519 ( .A1(n9468), .A2(n9467), .ZN(n9575) );
  NOR2_X1 U9520 ( .A1(n8573), .A2(n8582), .ZN(n9469) );
  NOR2_X1 U9521 ( .A1(n9467), .A2(n9468), .ZN(n9572) );
  NOR2_X1 U9522 ( .A1(n9576), .A2(n9577), .ZN(n9468) );
  INV_X1 U9523 ( .A(n9578), .ZN(n9577) );
  NAND2_X1 U9524 ( .A1(n9464), .A2(n9579), .ZN(n9578) );
  NAND2_X1 U9525 ( .A1(n9465), .A2(n9463), .ZN(n9579) );
  NOR2_X1 U9526 ( .A1(n8573), .A2(n8591), .ZN(n9464) );
  NOR2_X1 U9527 ( .A1(n9463), .A2(n9465), .ZN(n9576) );
  NOR2_X1 U9528 ( .A1(n9580), .A2(n9581), .ZN(n9465) );
  INV_X1 U9529 ( .A(n9582), .ZN(n9581) );
  NAND2_X1 U9530 ( .A1(n9461), .A2(n9583), .ZN(n9582) );
  NAND2_X1 U9531 ( .A1(n9460), .A2(n9459), .ZN(n9583) );
  NOR2_X1 U9532 ( .A1(n8573), .A2(n8562), .ZN(n9461) );
  NOR2_X1 U9533 ( .A1(n9459), .A2(n9460), .ZN(n9580) );
  NOR2_X1 U9534 ( .A1(n9584), .A2(n9585), .ZN(n9460) );
  INV_X1 U9535 ( .A(n9586), .ZN(n9585) );
  NAND2_X1 U9536 ( .A1(n9456), .A2(n9587), .ZN(n9586) );
  NAND2_X1 U9537 ( .A1(n9457), .A2(n9455), .ZN(n9587) );
  NOR2_X1 U9538 ( .A1(n8573), .A2(n8545), .ZN(n9456) );
  NOR2_X1 U9539 ( .A1(n9455), .A2(n9457), .ZN(n9584) );
  NOR2_X1 U9540 ( .A1(n9588), .A2(n9589), .ZN(n9457) );
  INV_X1 U9541 ( .A(n9590), .ZN(n9589) );
  NAND2_X1 U9542 ( .A1(n9453), .A2(n9591), .ZN(n9590) );
  NAND2_X1 U9543 ( .A1(n9452), .A2(n9451), .ZN(n9591) );
  NOR2_X1 U9544 ( .A1(n8573), .A2(n8569), .ZN(n9453) );
  NOR2_X1 U9545 ( .A1(n9451), .A2(n9452), .ZN(n9588) );
  NOR2_X1 U9546 ( .A1(n9592), .A2(n9593), .ZN(n9452) );
  INV_X1 U9547 ( .A(n9594), .ZN(n9593) );
  NAND2_X1 U9548 ( .A1(n9449), .A2(n9595), .ZN(n9594) );
  NAND2_X1 U9549 ( .A1(n9448), .A2(n9446), .ZN(n9595) );
  NOR2_X1 U9550 ( .A1(n8573), .A2(n8593), .ZN(n9449) );
  NOR2_X1 U9551 ( .A1(n9446), .A2(n9448), .ZN(n9592) );
  NOR2_X1 U9552 ( .A1(n9596), .A2(n9597), .ZN(n9448) );
  INV_X1 U9553 ( .A(n9598), .ZN(n9597) );
  NAND2_X1 U9554 ( .A1(n9445), .A2(n9599), .ZN(n9598) );
  NAND2_X1 U9555 ( .A1(n9444), .A2(n9443), .ZN(n9599) );
  NOR2_X1 U9556 ( .A1(n8573), .A2(n8583), .ZN(n9445) );
  NOR2_X1 U9557 ( .A1(n9443), .A2(n9444), .ZN(n9596) );
  NOR2_X1 U9558 ( .A1(n9600), .A2(n9601), .ZN(n9444) );
  INV_X1 U9559 ( .A(n9602), .ZN(n9601) );
  NAND2_X1 U9560 ( .A1(n9441), .A2(n9603), .ZN(n9602) );
  NAND2_X1 U9561 ( .A1(n9440), .A2(n9438), .ZN(n9603) );
  NOR2_X1 U9562 ( .A1(n8573), .A2(n8580), .ZN(n9441) );
  NOR2_X1 U9563 ( .A1(n9438), .A2(n9440), .ZN(n9600) );
  NOR2_X1 U9564 ( .A1(n9604), .A2(n9605), .ZN(n9440) );
  INV_X1 U9565 ( .A(n9606), .ZN(n9605) );
  NAND2_X1 U9566 ( .A1(n9437), .A2(n9607), .ZN(n9606) );
  NAND2_X1 U9567 ( .A1(n9436), .A2(n9435), .ZN(n9607) );
  NOR2_X1 U9568 ( .A1(n9156), .A2(n8588), .ZN(n9437) );
  NOR2_X1 U9569 ( .A1(n9435), .A2(n9436), .ZN(n9604) );
  NOR2_X1 U9570 ( .A1(n9608), .A2(n9609), .ZN(n9436) );
  INV_X1 U9571 ( .A(n9610), .ZN(n9609) );
  NAND2_X1 U9572 ( .A1(n9433), .A2(n9611), .ZN(n9610) );
  NAND2_X1 U9573 ( .A1(n9432), .A2(n9430), .ZN(n9611) );
  NOR2_X1 U9574 ( .A1(n9156), .A2(n8551), .ZN(n9433) );
  NOR2_X1 U9575 ( .A1(n9430), .A2(n9432), .ZN(n9608) );
  NOR2_X1 U9576 ( .A1(n9612), .A2(n9613), .ZN(n9432) );
  INV_X1 U9577 ( .A(n9614), .ZN(n9613) );
  NAND2_X1 U9578 ( .A1(n9429), .A2(n9615), .ZN(n9614) );
  NAND2_X1 U9579 ( .A1(n9428), .A2(n9427), .ZN(n9615) );
  NOR2_X1 U9580 ( .A1(n9156), .A2(n8563), .ZN(n9429) );
  NOR2_X1 U9581 ( .A1(n9427), .A2(n9428), .ZN(n9612) );
  NOR2_X1 U9582 ( .A1(n9616), .A2(n9617), .ZN(n9428) );
  INV_X1 U9583 ( .A(n9618), .ZN(n9617) );
  NAND2_X1 U9584 ( .A1(n9425), .A2(n9619), .ZN(n9618) );
  NAND2_X1 U9585 ( .A1(n9424), .A2(n9422), .ZN(n9619) );
  NOR2_X1 U9586 ( .A1(n9156), .A2(n8548), .ZN(n9425) );
  NOR2_X1 U9587 ( .A1(n9422), .A2(n9424), .ZN(n9616) );
  NOR2_X1 U9588 ( .A1(n9620), .A2(n9621), .ZN(n9424) );
  INV_X1 U9589 ( .A(n9622), .ZN(n9621) );
  NAND2_X1 U9590 ( .A1(n9421), .A2(n9623), .ZN(n9622) );
  NAND2_X1 U9591 ( .A1(n9420), .A2(n9419), .ZN(n9623) );
  NOR2_X1 U9592 ( .A1(n9156), .A2(n8584), .ZN(n9421) );
  NOR2_X1 U9593 ( .A1(n9419), .A2(n9420), .ZN(n9620) );
  NOR2_X1 U9594 ( .A1(n9624), .A2(n9625), .ZN(n9420) );
  INV_X1 U9595 ( .A(n9626), .ZN(n9625) );
  NAND2_X1 U9596 ( .A1(n9416), .A2(n9627), .ZN(n9626) );
  NAND2_X1 U9597 ( .A1(n9417), .A2(n9415), .ZN(n9627) );
  NOR2_X1 U9598 ( .A1(n9156), .A2(n8535), .ZN(n9416) );
  NOR2_X1 U9599 ( .A1(n9415), .A2(n9417), .ZN(n9624) );
  NOR2_X1 U9600 ( .A1(n9628), .A2(n9629), .ZN(n9417) );
  INV_X1 U9601 ( .A(n9630), .ZN(n9629) );
  NAND2_X1 U9602 ( .A1(n9413), .A2(n9631), .ZN(n9630) );
  NAND2_X1 U9603 ( .A1(n9412), .A2(n9411), .ZN(n9631) );
  NOR2_X1 U9604 ( .A1(n9156), .A2(n8568), .ZN(n9413) );
  NOR2_X1 U9605 ( .A1(n9411), .A2(n9412), .ZN(n9628) );
  NOR2_X1 U9606 ( .A1(n9632), .A2(n9633), .ZN(n9412) );
  INV_X1 U9607 ( .A(n9634), .ZN(n9633) );
  NAND2_X1 U9608 ( .A1(n9408), .A2(n9635), .ZN(n9634) );
  NAND2_X1 U9609 ( .A1(n9409), .A2(n9407), .ZN(n9635) );
  NOR2_X1 U9610 ( .A1(n9156), .A2(n8574), .ZN(n9408) );
  NOR2_X1 U9611 ( .A1(n9407), .A2(n9409), .ZN(n9632) );
  NOR2_X1 U9612 ( .A1(n9636), .A2(n9637), .ZN(n9409) );
  INV_X1 U9613 ( .A(n9638), .ZN(n9637) );
  NAND2_X1 U9614 ( .A1(n9404), .A2(n9639), .ZN(n9638) );
  NAND2_X1 U9615 ( .A1(n9405), .A2(n9403), .ZN(n9639) );
  NOR2_X1 U9616 ( .A1(n9156), .A2(n8565), .ZN(n9404) );
  NOR2_X1 U9617 ( .A1(n9403), .A2(n9405), .ZN(n9636) );
  NOR2_X1 U9618 ( .A1(n9640), .A2(n9641), .ZN(n9405) );
  INV_X1 U9619 ( .A(n9642), .ZN(n9641) );
  NAND2_X1 U9620 ( .A1(n9398), .A2(n9643), .ZN(n9642) );
  NAND2_X1 U9621 ( .A1(n9401), .A2(n9400), .ZN(n9643) );
  NOR2_X1 U9622 ( .A1(n9156), .A2(n8567), .ZN(n9398) );
  NOR2_X1 U9623 ( .A1(n9400), .A2(n9401), .ZN(n9640) );
  INV_X1 U9624 ( .A(n9644), .ZN(n9401) );
  NAND2_X1 U9625 ( .A1(n9645), .A2(n9646), .ZN(n9644) );
  NAND2_X1 U9626 ( .A1(n8549), .A2(n9647), .ZN(n9646) );
  NAND2_X1 U9627 ( .A1(n8624), .A2(n9648), .ZN(n9647) );
  NAND2_X1 U9628 ( .A1(n8586), .A2(n8585), .ZN(n9648) );
  NAND2_X1 U9629 ( .A1(n9650), .A2(n9651), .ZN(n9645) );
  NAND2_X1 U9630 ( .A1(n8630), .A2(n9652), .ZN(n9651) );
  NAND2_X1 U9631 ( .A1(n8539), .A2(n8550), .ZN(n9652) );
  NAND3_X1 U9632 ( .A1(n8549), .A2(n8537), .A3(n9157), .ZN(n9400) );
  XOR2_X1 U9633 ( .A(n9653), .B(n9654), .Z(n9403) );
  XNOR2_X1 U9634 ( .A(n9655), .B(n9656), .ZN(n9654) );
  XOR2_X1 U9635 ( .A(n9657), .B(n9658), .Z(n9407) );
  XNOR2_X1 U9636 ( .A(n9659), .B(n9660), .ZN(n9657) );
  XOR2_X1 U9637 ( .A(n9661), .B(n9662), .Z(n9411) );
  XNOR2_X1 U9638 ( .A(n9663), .B(n9664), .ZN(n9661) );
  XOR2_X1 U9639 ( .A(n9665), .B(n9666), .Z(n9415) );
  XNOR2_X1 U9640 ( .A(n9667), .B(n9668), .ZN(n9665) );
  XOR2_X1 U9641 ( .A(n9669), .B(n9670), .Z(n9419) );
  XNOR2_X1 U9642 ( .A(n9671), .B(n9672), .ZN(n9669) );
  NOR2_X1 U9643 ( .A1(n8535), .A2(n8550), .ZN(n9672) );
  XOR2_X1 U9644 ( .A(n9673), .B(n9674), .Z(n9422) );
  XNOR2_X1 U9645 ( .A(n9675), .B(n9676), .ZN(n9673) );
  NOR2_X1 U9646 ( .A1(n8584), .A2(n8550), .ZN(n9676) );
  XOR2_X1 U9647 ( .A(n9677), .B(n9678), .Z(n9427) );
  XNOR2_X1 U9648 ( .A(n9679), .B(n9680), .ZN(n9677) );
  NOR2_X1 U9649 ( .A1(n8548), .A2(n8550), .ZN(n9680) );
  XOR2_X1 U9650 ( .A(n9681), .B(n9682), .Z(n9430) );
  XNOR2_X1 U9651 ( .A(n9683), .B(n9684), .ZN(n9681) );
  NOR2_X1 U9652 ( .A1(n8563), .A2(n8550), .ZN(n9684) );
  XOR2_X1 U9653 ( .A(n9685), .B(n9686), .Z(n9435) );
  XNOR2_X1 U9654 ( .A(n9687), .B(n9688), .ZN(n9685) );
  NOR2_X1 U9655 ( .A1(n8551), .A2(n8550), .ZN(n9688) );
  XOR2_X1 U9656 ( .A(n9689), .B(n9690), .Z(n9438) );
  XNOR2_X1 U9657 ( .A(n9691), .B(n9692), .ZN(n9689) );
  NOR2_X1 U9658 ( .A1(n8588), .A2(n8550), .ZN(n9692) );
  XOR2_X1 U9659 ( .A(n9693), .B(n9694), .Z(n9443) );
  XNOR2_X1 U9660 ( .A(n9695), .B(n9696), .ZN(n9693) );
  NOR2_X1 U9661 ( .A1(n8580), .A2(n8550), .ZN(n9696) );
  XOR2_X1 U9662 ( .A(n9697), .B(n9698), .Z(n9446) );
  XNOR2_X1 U9663 ( .A(n9699), .B(n9700), .ZN(n9697) );
  NOR2_X1 U9664 ( .A1(n8583), .A2(n8550), .ZN(n9700) );
  XOR2_X1 U9665 ( .A(n9701), .B(n9702), .Z(n9451) );
  XNOR2_X1 U9666 ( .A(n9703), .B(n9704), .ZN(n9701) );
  NOR2_X1 U9667 ( .A1(n8593), .A2(n8550), .ZN(n9704) );
  XOR2_X1 U9668 ( .A(n9705), .B(n9706), .Z(n9455) );
  XNOR2_X1 U9669 ( .A(n9707), .B(n9708), .ZN(n9705) );
  NOR2_X1 U9670 ( .A1(n8569), .A2(n8550), .ZN(n9708) );
  XOR2_X1 U9671 ( .A(n9709), .B(n9710), .Z(n9459) );
  XNOR2_X1 U9672 ( .A(n9711), .B(n9712), .ZN(n9709) );
  NOR2_X1 U9673 ( .A1(n8545), .A2(n8550), .ZN(n9712) );
  XOR2_X1 U9674 ( .A(n9713), .B(n9714), .Z(n9463) );
  XNOR2_X1 U9675 ( .A(n9715), .B(n9716), .ZN(n9713) );
  NOR2_X1 U9676 ( .A1(n8562), .A2(n8550), .ZN(n9716) );
  XNOR2_X1 U9677 ( .A(n9717), .B(n9718), .ZN(n9467) );
  XNOR2_X1 U9678 ( .A(n9719), .B(n9720), .ZN(n9718) );
  NAND2_X1 U9679 ( .A1(n8549), .A2(n9721), .ZN(n9720) );
  XOR2_X1 U9680 ( .A(n9722), .B(n9723), .Z(n9471) );
  XNOR2_X1 U9681 ( .A(n9724), .B(n9725), .ZN(n9722) );
  NOR2_X1 U9682 ( .A1(n8582), .A2(n8550), .ZN(n9725) );
  XOR2_X1 U9683 ( .A(n9726), .B(n9727), .Z(n9474) );
  XNOR2_X1 U9684 ( .A(n9728), .B(n9729), .ZN(n9726) );
  NOR2_X1 U9685 ( .A1(n8572), .A2(n8550), .ZN(n9729) );
  XNOR2_X1 U9686 ( .A(n9730), .B(n9731), .ZN(n9479) );
  XNOR2_X1 U9687 ( .A(n9732), .B(n9733), .ZN(n9730) );
  NOR2_X1 U9688 ( .A1(n8556), .A2(n8550), .ZN(n9733) );
  XNOR2_X1 U9689 ( .A(n9734), .B(n9735), .ZN(n9483) );
  XNOR2_X1 U9690 ( .A(n9736), .B(n9737), .ZN(n9734) );
  NOR2_X1 U9691 ( .A1(n8594), .A2(n8550), .ZN(n9737) );
  XOR2_X1 U9692 ( .A(n9738), .B(n9739), .Z(n9487) );
  XNOR2_X1 U9693 ( .A(n9740), .B(n9741), .ZN(n9738) );
  NOR2_X1 U9694 ( .A1(n8560), .A2(n8550), .ZN(n9741) );
  XOR2_X1 U9695 ( .A(n9742), .B(n9743), .Z(n9490) );
  XNOR2_X1 U9696 ( .A(n9744), .B(n9745), .ZN(n9742) );
  NOR2_X1 U9697 ( .A1(n8544), .A2(n8550), .ZN(n9745) );
  XNOR2_X1 U9698 ( .A(n9746), .B(n9747), .ZN(n9495) );
  XNOR2_X1 U9699 ( .A(n9748), .B(n9749), .ZN(n9746) );
  NOR2_X1 U9700 ( .A1(n8555), .A2(n8550), .ZN(n9749) );
  XNOR2_X1 U9701 ( .A(n9750), .B(n9751), .ZN(n9498) );
  XNOR2_X1 U9702 ( .A(n9752), .B(n9753), .ZN(n9750) );
  NOR2_X1 U9703 ( .A1(n8564), .A2(n8550), .ZN(n9753) );
  XNOR2_X1 U9704 ( .A(n9754), .B(n9755), .ZN(n9503) );
  XNOR2_X1 U9705 ( .A(n9756), .B(n9757), .ZN(n9754) );
  NOR2_X1 U9706 ( .A1(n8528), .A2(n8550), .ZN(n9757) );
  NOR2_X1 U9707 ( .A1(n9509), .A2(n9506), .ZN(n9531) );
  XOR2_X1 U9708 ( .A(n9758), .B(n9759), .Z(n9506) );
  XNOR2_X1 U9709 ( .A(n9760), .B(n9761), .ZN(n9758) );
  NOR2_X1 U9710 ( .A1(n8527), .A2(n8550), .ZN(n9761) );
  NAND2_X1 U9711 ( .A1(n9157), .A2(n9268), .ZN(n9509) );
  INV_X1 U9712 ( .A(n9156), .ZN(n9157) );
  XNOR2_X1 U9713 ( .A(n9762), .B(n9763), .ZN(n9156) );
  XOR2_X1 U9714 ( .A(d_29_), .B(c_29_), .Z(n9763) );
  XOR2_X1 U9715 ( .A(n9764), .B(n9765), .Z(n9511) );
  XNOR2_X1 U9716 ( .A(n9766), .B(n9767), .ZN(n9764) );
  XNOR2_X1 U9717 ( .A(n9768), .B(n9769), .ZN(n8960) );
  XOR2_X1 U9718 ( .A(n9770), .B(n9771), .Z(n9769) );
  NAND2_X1 U9719 ( .A1(n8549), .A2(n8592), .ZN(n9771) );
  NAND2_X1 U9720 ( .A1(n9772), .A2(n9773), .ZN(n8791) );
  NAND2_X1 U9721 ( .A1(n8955), .A2(n8797), .ZN(n9773) );
  INV_X1 U9722 ( .A(n9774), .ZN(n8797) );
  NAND2_X1 U9723 ( .A1(n9775), .A2(n9776), .ZN(n8955) );
  NAND2_X1 U9724 ( .A1(n8954), .A2(n8956), .ZN(n9772) );
  NAND2_X1 U9725 ( .A1(n9777), .A2(n9778), .ZN(n8956) );
  INV_X1 U9726 ( .A(n9779), .ZN(n9778) );
  NOR3_X1 U9727 ( .A1(n8972), .A2(n9780), .A3(n8550), .ZN(n9779) );
  NOR2_X1 U9728 ( .A1(n9770), .A2(n9768), .ZN(n9780) );
  NAND2_X1 U9729 ( .A1(n9768), .A2(n9770), .ZN(n9777) );
  NAND2_X1 U9730 ( .A1(n9781), .A2(n9782), .ZN(n9770) );
  NAND2_X1 U9731 ( .A1(n9524), .A2(n9783), .ZN(n9782) );
  INV_X1 U9732 ( .A(n9784), .ZN(n9783) );
  NOR2_X1 U9733 ( .A1(n9525), .A2(n9523), .ZN(n9784) );
  NOR2_X1 U9734 ( .A1(n8550), .A2(n8589), .ZN(n9524) );
  NAND2_X1 U9735 ( .A1(n9523), .A2(n9525), .ZN(n9781) );
  NAND2_X1 U9736 ( .A1(n9785), .A2(n9786), .ZN(n9525) );
  NAND2_X1 U9737 ( .A1(n9767), .A2(n9787), .ZN(n9786) );
  NAND2_X1 U9738 ( .A1(n9766), .A2(n9765), .ZN(n9787) );
  NOR2_X1 U9739 ( .A1(n8550), .A2(n8552), .ZN(n9767) );
  INV_X1 U9740 ( .A(n9788), .ZN(n9785) );
  NOR2_X1 U9741 ( .A1(n9765), .A2(n9766), .ZN(n9788) );
  NOR2_X1 U9742 ( .A1(n9789), .A2(n9790), .ZN(n9766) );
  INV_X1 U9743 ( .A(n9791), .ZN(n9790) );
  NAND3_X1 U9744 ( .A1(n9792), .A2(n9793), .A3(n8549), .ZN(n9791) );
  NAND2_X1 U9745 ( .A1(n9760), .A2(n9759), .ZN(n9793) );
  NOR2_X1 U9746 ( .A1(n9759), .A2(n9760), .ZN(n9789) );
  NOR2_X1 U9747 ( .A1(n9794), .A2(n9795), .ZN(n9760) );
  INV_X1 U9748 ( .A(n9796), .ZN(n9795) );
  NAND3_X1 U9749 ( .A1(n9277), .A2(n9797), .A3(n8549), .ZN(n9796) );
  NAND2_X1 U9750 ( .A1(n9756), .A2(n9755), .ZN(n9797) );
  NOR2_X1 U9751 ( .A1(n9755), .A2(n9756), .ZN(n9794) );
  NOR2_X1 U9752 ( .A1(n9798), .A2(n9799), .ZN(n9756) );
  NOR3_X1 U9753 ( .A1(n8995), .A2(n9800), .A3(n8550), .ZN(n9799) );
  INV_X1 U9754 ( .A(n9801), .ZN(n9800) );
  NAND2_X1 U9755 ( .A1(n9752), .A2(n9751), .ZN(n9801) );
  NOR2_X1 U9756 ( .A1(n9751), .A2(n9752), .ZN(n9798) );
  NOR2_X1 U9757 ( .A1(n9802), .A2(n9803), .ZN(n9752) );
  INV_X1 U9758 ( .A(n9804), .ZN(n9803) );
  NAND3_X1 U9759 ( .A1(n9286), .A2(n9805), .A3(n8549), .ZN(n9804) );
  NAND2_X1 U9760 ( .A1(n9748), .A2(n9747), .ZN(n9805) );
  NOR2_X1 U9761 ( .A1(n9747), .A2(n9748), .ZN(n9802) );
  NOR2_X1 U9762 ( .A1(n9806), .A2(n9807), .ZN(n9748) );
  NOR3_X1 U9763 ( .A1(n8544), .A2(n9808), .A3(n8550), .ZN(n9807) );
  INV_X1 U9764 ( .A(n9809), .ZN(n9808) );
  NAND2_X1 U9765 ( .A1(n9744), .A2(n9743), .ZN(n9809) );
  NOR2_X1 U9766 ( .A1(n9743), .A2(n9744), .ZN(n9806) );
  NOR2_X1 U9767 ( .A1(n9810), .A2(n9811), .ZN(n9744) );
  INV_X1 U9768 ( .A(n9812), .ZN(n9811) );
  NAND3_X1 U9769 ( .A1(n9295), .A2(n9813), .A3(n8549), .ZN(n9812) );
  NAND2_X1 U9770 ( .A1(n9740), .A2(n9739), .ZN(n9813) );
  NOR2_X1 U9771 ( .A1(n9739), .A2(n9740), .ZN(n9810) );
  NOR2_X1 U9772 ( .A1(n9814), .A2(n9815), .ZN(n9740) );
  NOR3_X1 U9773 ( .A1(n9014), .A2(n9816), .A3(n8550), .ZN(n9815) );
  INV_X1 U9774 ( .A(n9817), .ZN(n9816) );
  NAND2_X1 U9775 ( .A1(n9736), .A2(n9735), .ZN(n9817) );
  NOR2_X1 U9776 ( .A1(n9735), .A2(n9736), .ZN(n9814) );
  NOR2_X1 U9777 ( .A1(n9818), .A2(n9819), .ZN(n9736) );
  INV_X1 U9778 ( .A(n9820), .ZN(n9819) );
  NAND3_X1 U9779 ( .A1(n9304), .A2(n9821), .A3(n8549), .ZN(n9820) );
  NAND2_X1 U9780 ( .A1(n9732), .A2(n9731), .ZN(n9821) );
  NOR2_X1 U9781 ( .A1(n9731), .A2(n9732), .ZN(n9818) );
  NOR2_X1 U9782 ( .A1(n9822), .A2(n9823), .ZN(n9732) );
  NOR3_X1 U9783 ( .A1(n9025), .A2(n9824), .A3(n8550), .ZN(n9823) );
  INV_X1 U9784 ( .A(n9825), .ZN(n9824) );
  NAND2_X1 U9785 ( .A1(n9728), .A2(n9727), .ZN(n9825) );
  NOR2_X1 U9786 ( .A1(n9727), .A2(n9728), .ZN(n9822) );
  NOR2_X1 U9787 ( .A1(n9826), .A2(n9827), .ZN(n9728) );
  INV_X1 U9788 ( .A(n9828), .ZN(n9827) );
  NAND3_X1 U9789 ( .A1(n9313), .A2(n9829), .A3(n8549), .ZN(n9828) );
  NAND2_X1 U9790 ( .A1(n9724), .A2(n9723), .ZN(n9829) );
  NOR2_X1 U9791 ( .A1(n9723), .A2(n9724), .ZN(n9826) );
  NOR2_X1 U9792 ( .A1(n9830), .A2(n9831), .ZN(n9724) );
  NOR3_X1 U9793 ( .A1(n9036), .A2(n9832), .A3(n8550), .ZN(n9831) );
  INV_X1 U9794 ( .A(n9833), .ZN(n9832) );
  NAND2_X1 U9795 ( .A1(n9719), .A2(n9717), .ZN(n9833) );
  NOR2_X1 U9796 ( .A1(n9717), .A2(n9719), .ZN(n9830) );
  NOR2_X1 U9797 ( .A1(n9834), .A2(n9835), .ZN(n9719) );
  INV_X1 U9798 ( .A(n9836), .ZN(n9835) );
  NAND3_X1 U9799 ( .A1(n9322), .A2(n9837), .A3(n8549), .ZN(n9836) );
  NAND2_X1 U9800 ( .A1(n9715), .A2(n9714), .ZN(n9837) );
  NOR2_X1 U9801 ( .A1(n9714), .A2(n9715), .ZN(n9834) );
  NOR2_X1 U9802 ( .A1(n9838), .A2(n9839), .ZN(n9715) );
  NOR3_X1 U9803 ( .A1(n8545), .A2(n9840), .A3(n8550), .ZN(n9839) );
  INV_X1 U9804 ( .A(n9841), .ZN(n9840) );
  NAND2_X1 U9805 ( .A1(n9711), .A2(n9710), .ZN(n9841) );
  NOR2_X1 U9806 ( .A1(n9710), .A2(n9711), .ZN(n9838) );
  NOR2_X1 U9807 ( .A1(n9842), .A2(n9843), .ZN(n9711) );
  INV_X1 U9808 ( .A(n9844), .ZN(n9843) );
  NAND3_X1 U9809 ( .A1(n9331), .A2(n9845), .A3(n8549), .ZN(n9844) );
  NAND2_X1 U9810 ( .A1(n9707), .A2(n9706), .ZN(n9845) );
  NOR2_X1 U9811 ( .A1(n9706), .A2(n9707), .ZN(n9842) );
  NOR2_X1 U9812 ( .A1(n9846), .A2(n9847), .ZN(n9707) );
  NOR3_X1 U9813 ( .A1(n9056), .A2(n9848), .A3(n8550), .ZN(n9847) );
  INV_X1 U9814 ( .A(n9849), .ZN(n9848) );
  NAND2_X1 U9815 ( .A1(n9703), .A2(n9702), .ZN(n9849) );
  NOR2_X1 U9816 ( .A1(n9702), .A2(n9703), .ZN(n9846) );
  NOR2_X1 U9817 ( .A1(n9850), .A2(n9851), .ZN(n9703) );
  INV_X1 U9818 ( .A(n9852), .ZN(n9851) );
  NAND3_X1 U9819 ( .A1(n9340), .A2(n9853), .A3(n8549), .ZN(n9852) );
  NAND2_X1 U9820 ( .A1(n9699), .A2(n9698), .ZN(n9853) );
  NOR2_X1 U9821 ( .A1(n9698), .A2(n9699), .ZN(n9850) );
  NOR2_X1 U9822 ( .A1(n9854), .A2(n9855), .ZN(n9699) );
  NOR3_X1 U9823 ( .A1(n8580), .A2(n9856), .A3(n8550), .ZN(n9855) );
  INV_X1 U9824 ( .A(n9857), .ZN(n9856) );
  NAND2_X1 U9825 ( .A1(n9695), .A2(n9694), .ZN(n9857) );
  NOR2_X1 U9826 ( .A1(n9694), .A2(n9695), .ZN(n9854) );
  NOR2_X1 U9827 ( .A1(n9858), .A2(n9859), .ZN(n9695) );
  INV_X1 U9828 ( .A(n9860), .ZN(n9859) );
  NAND3_X1 U9829 ( .A1(n9080), .A2(n9861), .A3(n8549), .ZN(n9860) );
  NAND2_X1 U9830 ( .A1(n9691), .A2(n9690), .ZN(n9861) );
  NOR2_X1 U9831 ( .A1(n9690), .A2(n9691), .ZN(n9858) );
  NOR2_X1 U9832 ( .A1(n9862), .A2(n9863), .ZN(n9691) );
  NOR3_X1 U9833 ( .A1(n8551), .A2(n9864), .A3(n8550), .ZN(n9863) );
  INV_X1 U9834 ( .A(n9865), .ZN(n9864) );
  NAND2_X1 U9835 ( .A1(n9687), .A2(n9686), .ZN(n9865) );
  NOR2_X1 U9836 ( .A1(n9686), .A2(n9687), .ZN(n9862) );
  NOR2_X1 U9837 ( .A1(n9866), .A2(n9867), .ZN(n9687) );
  INV_X1 U9838 ( .A(n9868), .ZN(n9867) );
  NAND3_X1 U9839 ( .A1(n9098), .A2(n9869), .A3(n8549), .ZN(n9868) );
  NAND2_X1 U9840 ( .A1(n9683), .A2(n9682), .ZN(n9869) );
  NOR2_X1 U9841 ( .A1(n9682), .A2(n9683), .ZN(n9866) );
  NOR2_X1 U9842 ( .A1(n9870), .A2(n9871), .ZN(n9683) );
  NOR3_X1 U9843 ( .A1(n8548), .A2(n9872), .A3(n8550), .ZN(n9871) );
  INV_X1 U9844 ( .A(n9873), .ZN(n9872) );
  NAND2_X1 U9845 ( .A1(n9679), .A2(n9678), .ZN(n9873) );
  NOR2_X1 U9846 ( .A1(n9678), .A2(n9679), .ZN(n9870) );
  NOR2_X1 U9847 ( .A1(n9874), .A2(n9875), .ZN(n9679) );
  INV_X1 U9848 ( .A(n9876), .ZN(n9875) );
  NAND3_X1 U9849 ( .A1(n9112), .A2(n9877), .A3(n8549), .ZN(n9876) );
  NAND2_X1 U9850 ( .A1(n9675), .A2(n9674), .ZN(n9877) );
  NOR2_X1 U9851 ( .A1(n9674), .A2(n9675), .ZN(n9874) );
  NOR2_X1 U9852 ( .A1(n9878), .A2(n9879), .ZN(n9675) );
  INV_X1 U9853 ( .A(n9880), .ZN(n9879) );
  NAND3_X1 U9854 ( .A1(n9121), .A2(n9881), .A3(n8549), .ZN(n9880) );
  NAND2_X1 U9855 ( .A1(n9671), .A2(n9670), .ZN(n9881) );
  NOR2_X1 U9856 ( .A1(n9670), .A2(n9671), .ZN(n9878) );
  NOR2_X1 U9857 ( .A1(n9882), .A2(n9883), .ZN(n9671) );
  INV_X1 U9858 ( .A(n9884), .ZN(n9883) );
  NAND2_X1 U9859 ( .A1(n9667), .A2(n9885), .ZN(n9884) );
  NAND2_X1 U9860 ( .A1(n9668), .A2(n9666), .ZN(n9885) );
  NOR2_X1 U9861 ( .A1(n8550), .A2(n8568), .ZN(n9667) );
  NOR2_X1 U9862 ( .A1(n9666), .A2(n9668), .ZN(n9882) );
  NOR2_X1 U9863 ( .A1(n9886), .A2(n9887), .ZN(n9668) );
  INV_X1 U9864 ( .A(n9888), .ZN(n9887) );
  NAND2_X1 U9865 ( .A1(n9663), .A2(n9889), .ZN(n9888) );
  NAND2_X1 U9866 ( .A1(n9664), .A2(n9662), .ZN(n9889) );
  NOR2_X1 U9867 ( .A1(n8550), .A2(n8574), .ZN(n9663) );
  NOR2_X1 U9868 ( .A1(n9662), .A2(n9664), .ZN(n9886) );
  NOR2_X1 U9869 ( .A1(n9890), .A2(n9891), .ZN(n9664) );
  INV_X1 U9870 ( .A(n9892), .ZN(n9891) );
  NAND2_X1 U9871 ( .A1(n9659), .A2(n9893), .ZN(n9892) );
  NAND2_X1 U9872 ( .A1(n9660), .A2(n9658), .ZN(n9893) );
  NOR2_X1 U9873 ( .A1(n8550), .A2(n8565), .ZN(n9659) );
  NOR2_X1 U9874 ( .A1(n9658), .A2(n9660), .ZN(n9890) );
  NOR2_X1 U9875 ( .A1(n9894), .A2(n9895), .ZN(n9660) );
  INV_X1 U9876 ( .A(n9896), .ZN(n9895) );
  NAND2_X1 U9877 ( .A1(n9653), .A2(n9897), .ZN(n9896) );
  NAND2_X1 U9878 ( .A1(n9656), .A2(n9655), .ZN(n9897) );
  NOR2_X1 U9879 ( .A1(n8550), .A2(n8567), .ZN(n9653) );
  NOR2_X1 U9880 ( .A1(n9655), .A2(n9656), .ZN(n9894) );
  INV_X1 U9881 ( .A(n9898), .ZN(n9656) );
  NAND2_X1 U9882 ( .A1(n9899), .A2(n9900), .ZN(n9898) );
  NAND2_X1 U9883 ( .A1(n9650), .A2(n9901), .ZN(n9900) );
  NAND2_X1 U9884 ( .A1(n8624), .A2(n9902), .ZN(n9901) );
  NAND2_X1 U9885 ( .A1(n8542), .A2(n8585), .ZN(n9902) );
  NAND2_X1 U9886 ( .A1(n9903), .A2(n9904), .ZN(n9899) );
  NAND2_X1 U9887 ( .A1(n8630), .A2(n9905), .ZN(n9904) );
  NAND2_X1 U9888 ( .A1(n8539), .A2(n8586), .ZN(n9905) );
  NAND3_X1 U9889 ( .A1(n9650), .A2(n8537), .A3(n8549), .ZN(n9655) );
  XOR2_X1 U9890 ( .A(n9906), .B(n9907), .Z(n9393) );
  XNOR2_X1 U9891 ( .A(c_28_), .B(d_28_), .ZN(n9906) );
  XOR2_X1 U9892 ( .A(n9908), .B(n9909), .Z(n9658) );
  XNOR2_X1 U9893 ( .A(n9910), .B(n9911), .ZN(n9909) );
  XOR2_X1 U9894 ( .A(n9912), .B(n9913), .Z(n9662) );
  XNOR2_X1 U9895 ( .A(n9914), .B(n9915), .ZN(n9912) );
  XOR2_X1 U9896 ( .A(n9916), .B(n9917), .Z(n9666) );
  XNOR2_X1 U9897 ( .A(n9918), .B(n9919), .ZN(n9916) );
  XOR2_X1 U9898 ( .A(n9920), .B(n9921), .Z(n9670) );
  XNOR2_X1 U9899 ( .A(n9922), .B(n9923), .ZN(n9920) );
  XOR2_X1 U9900 ( .A(n9924), .B(n9925), .Z(n9674) );
  XNOR2_X1 U9901 ( .A(n9926), .B(n9927), .ZN(n9924) );
  XOR2_X1 U9902 ( .A(n9928), .B(n9929), .Z(n9678) );
  XNOR2_X1 U9903 ( .A(n9930), .B(n9931), .ZN(n9928) );
  XNOR2_X1 U9904 ( .A(n9932), .B(n9933), .ZN(n9682) );
  XOR2_X1 U9905 ( .A(n9934), .B(n9935), .Z(n9933) );
  XOR2_X1 U9906 ( .A(n9936), .B(n9937), .Z(n9686) );
  XNOR2_X1 U9907 ( .A(n9938), .B(n9939), .ZN(n9936) );
  XNOR2_X1 U9908 ( .A(n9940), .B(n9941), .ZN(n9690) );
  XOR2_X1 U9909 ( .A(n9942), .B(n9943), .Z(n9941) );
  XOR2_X1 U9910 ( .A(n9944), .B(n9945), .Z(n9694) );
  XNOR2_X1 U9911 ( .A(n9946), .B(n9947), .ZN(n9944) );
  XNOR2_X1 U9912 ( .A(n9948), .B(n9949), .ZN(n9698) );
  XOR2_X1 U9913 ( .A(n9950), .B(n9951), .Z(n9949) );
  XOR2_X1 U9914 ( .A(n9952), .B(n9953), .Z(n9702) );
  XNOR2_X1 U9915 ( .A(n9954), .B(n9955), .ZN(n9952) );
  XOR2_X1 U9916 ( .A(n9956), .B(n9957), .Z(n9706) );
  XNOR2_X1 U9917 ( .A(n9958), .B(n9959), .ZN(n9956) );
  XOR2_X1 U9918 ( .A(n9960), .B(n9961), .Z(n9710) );
  XNOR2_X1 U9919 ( .A(n9962), .B(n9963), .ZN(n9960) );
  XOR2_X1 U9920 ( .A(n9964), .B(n9965), .Z(n9714) );
  XNOR2_X1 U9921 ( .A(n9966), .B(n9967), .ZN(n9964) );
  XOR2_X1 U9922 ( .A(n9968), .B(n9969), .Z(n9717) );
  XNOR2_X1 U9923 ( .A(n9970), .B(n9971), .ZN(n9968) );
  XOR2_X1 U9924 ( .A(n9972), .B(n9973), .Z(n9723) );
  XNOR2_X1 U9925 ( .A(n9974), .B(n9975), .ZN(n9972) );
  XNOR2_X1 U9926 ( .A(n9976), .B(n9977), .ZN(n9727) );
  XOR2_X1 U9927 ( .A(n9978), .B(n9979), .Z(n9977) );
  XNOR2_X1 U9928 ( .A(n9980), .B(n9981), .ZN(n9731) );
  XOR2_X1 U9929 ( .A(n9982), .B(n9983), .Z(n9980) );
  XNOR2_X1 U9930 ( .A(n9984), .B(n9985), .ZN(n9735) );
  XOR2_X1 U9931 ( .A(n9986), .B(n9987), .Z(n9984) );
  XOR2_X1 U9932 ( .A(n9988), .B(n9989), .Z(n9739) );
  XNOR2_X1 U9933 ( .A(n9990), .B(n9991), .ZN(n9988) );
  XNOR2_X1 U9934 ( .A(n9992), .B(n9993), .ZN(n9743) );
  XOR2_X1 U9935 ( .A(n9994), .B(n9995), .Z(n9993) );
  XNOR2_X1 U9936 ( .A(n9996), .B(n9997), .ZN(n9747) );
  XOR2_X1 U9937 ( .A(n9998), .B(n9999), .Z(n9996) );
  NOR2_X1 U9938 ( .A1(n8544), .A2(n8586), .ZN(n9999) );
  XNOR2_X1 U9939 ( .A(n10000), .B(n10001), .ZN(n9751) );
  XOR2_X1 U9940 ( .A(n10002), .B(n10003), .Z(n10001) );
  XNOR2_X1 U9941 ( .A(n10004), .B(n10005), .ZN(n9755) );
  XOR2_X1 U9942 ( .A(n10006), .B(n10007), .Z(n10004) );
  XOR2_X1 U9943 ( .A(n10008), .B(n10009), .Z(n9759) );
  XNOR2_X1 U9944 ( .A(n10010), .B(n10011), .ZN(n10008) );
  XOR2_X1 U9945 ( .A(n10012), .B(n10013), .Z(n9765) );
  XNOR2_X1 U9946 ( .A(n10014), .B(n10015), .ZN(n10012) );
  NOR2_X1 U9947 ( .A1(n8527), .A2(n8586), .ZN(n10015) );
  XNOR2_X1 U9948 ( .A(n10016), .B(n10017), .ZN(n9523) );
  NAND2_X1 U9949 ( .A1(n10018), .A2(n10019), .ZN(n10016) );
  XOR2_X1 U9950 ( .A(n10020), .B(n10021), .Z(n9768) );
  XOR2_X1 U9951 ( .A(n10022), .B(n10023), .Z(n10020) );
  NOR2_X1 U9952 ( .A1(n8589), .A2(n8586), .ZN(n10023) );
  XOR2_X1 U9953 ( .A(n10024), .B(n10025), .Z(n8954) );
  XNOR2_X1 U9954 ( .A(n10026), .B(n10027), .ZN(n10025) );
  NAND2_X1 U9955 ( .A1(n9650), .A2(n8592), .ZN(n10027) );
  NAND2_X1 U9956 ( .A1(n9774), .A2(n8798), .ZN(n8794) );
  XOR2_X1 U9957 ( .A(n8951), .B(n8950), .Z(n8798) );
  NOR2_X1 U9958 ( .A1(n9776), .A2(n9775), .ZN(n9774) );
  NOR2_X1 U9959 ( .A1(n10028), .A2(n10029), .ZN(n9775) );
  NOR3_X1 U9960 ( .A1(n8972), .A2(n10030), .A3(n8586), .ZN(n10029) );
  INV_X1 U9961 ( .A(n10031), .ZN(n10030) );
  NAND2_X1 U9962 ( .A1(n10026), .A2(n10024), .ZN(n10031) );
  NOR2_X1 U9963 ( .A1(n10024), .A2(n10026), .ZN(n10028) );
  NOR2_X1 U9964 ( .A1(n10032), .A2(n10033), .ZN(n10026) );
  NOR3_X1 U9965 ( .A1(n8884), .A2(n10034), .A3(n8586), .ZN(n10033) );
  NOR2_X1 U9966 ( .A1(n10022), .A2(n10021), .ZN(n10034) );
  INV_X1 U9967 ( .A(n10035), .ZN(n10032) );
  NAND2_X1 U9968 ( .A1(n10021), .A2(n10022), .ZN(n10035) );
  NAND2_X1 U9969 ( .A1(n10018), .A2(n10036), .ZN(n10022) );
  NAND2_X1 U9970 ( .A1(n10017), .A2(n10019), .ZN(n10036) );
  NAND2_X1 U9971 ( .A1(n10037), .A2(n10038), .ZN(n10019) );
  NAND2_X1 U9972 ( .A1(n9650), .A2(n9268), .ZN(n10038) );
  XNOR2_X1 U9973 ( .A(n10039), .B(n10040), .ZN(n10017) );
  XOR2_X1 U9974 ( .A(n10041), .B(n10042), .Z(n10040) );
  NAND2_X1 U9975 ( .A1(n9268), .A2(n10043), .ZN(n10018) );
  INV_X1 U9976 ( .A(n10037), .ZN(n10043) );
  NOR2_X1 U9977 ( .A1(n10044), .A2(n10045), .ZN(n10037) );
  NOR3_X1 U9978 ( .A1(n8527), .A2(n10046), .A3(n8586), .ZN(n10045) );
  INV_X1 U9979 ( .A(n10047), .ZN(n10046) );
  NAND2_X1 U9980 ( .A1(n10014), .A2(n10013), .ZN(n10047) );
  NOR2_X1 U9981 ( .A1(n10013), .A2(n10014), .ZN(n10044) );
  NOR2_X1 U9982 ( .A1(n10048), .A2(n10049), .ZN(n10014) );
  INV_X1 U9983 ( .A(n10050), .ZN(n10049) );
  NAND2_X1 U9984 ( .A1(n10010), .A2(n10051), .ZN(n10050) );
  NAND2_X1 U9985 ( .A1(n10011), .A2(n10009), .ZN(n10051) );
  NOR2_X1 U9986 ( .A1(n8586), .A2(n8528), .ZN(n10010) );
  NOR2_X1 U9987 ( .A1(n10009), .A2(n10011), .ZN(n10048) );
  INV_X1 U9988 ( .A(n10052), .ZN(n10011) );
  NAND2_X1 U9989 ( .A1(n10053), .A2(n10054), .ZN(n10052) );
  NAND2_X1 U9990 ( .A1(n10007), .A2(n10055), .ZN(n10054) );
  INV_X1 U9991 ( .A(n10056), .ZN(n10055) );
  NOR2_X1 U9992 ( .A1(n10006), .A2(n10005), .ZN(n10056) );
  NOR2_X1 U9993 ( .A1(n8586), .A2(n8564), .ZN(n10007) );
  NAND2_X1 U9994 ( .A1(n10005), .A2(n10006), .ZN(n10053) );
  NAND2_X1 U9995 ( .A1(n10057), .A2(n10058), .ZN(n10006) );
  NAND2_X1 U9996 ( .A1(n10002), .A2(n10059), .ZN(n10058) );
  NAND2_X1 U9997 ( .A1(n10000), .A2(n10003), .ZN(n10059) );
  NAND2_X1 U9998 ( .A1(n10060), .A2(n10061), .ZN(n10002) );
  INV_X1 U9999 ( .A(n10062), .ZN(n10061) );
  NOR3_X1 U10000 ( .A1(n8544), .A2(n10063), .A3(n8586), .ZN(n10062) );
  NOR2_X1 U10001 ( .A1(n9998), .A2(n9997), .ZN(n10063) );
  NAND2_X1 U10002 ( .A1(n9997), .A2(n9998), .ZN(n10060) );
  NAND2_X1 U10003 ( .A1(n10064), .A2(n10065), .ZN(n9998) );
  NAND2_X1 U10004 ( .A1(n9995), .A2(n10066), .ZN(n10065) );
  NAND2_X1 U10005 ( .A1(n9994), .A2(n9992), .ZN(n10066) );
  NOR2_X1 U10006 ( .A1(n8586), .A2(n8560), .ZN(n9995) );
  INV_X1 U10007 ( .A(n10067), .ZN(n10064) );
  NOR2_X1 U10008 ( .A1(n9992), .A2(n9994), .ZN(n10067) );
  NOR2_X1 U10009 ( .A1(n10068), .A2(n10069), .ZN(n9994) );
  INV_X1 U10010 ( .A(n10070), .ZN(n10069) );
  NAND2_X1 U10011 ( .A1(n9991), .A2(n10071), .ZN(n10070) );
  NAND2_X1 U10012 ( .A1(n9990), .A2(n9989), .ZN(n10071) );
  NOR2_X1 U10013 ( .A1(n8586), .A2(n8594), .ZN(n9991) );
  NOR2_X1 U10014 ( .A1(n9989), .A2(n9990), .ZN(n10068) );
  INV_X1 U10015 ( .A(n10072), .ZN(n9990) );
  NAND2_X1 U10016 ( .A1(n10073), .A2(n10074), .ZN(n10072) );
  NAND2_X1 U10017 ( .A1(n9986), .A2(n10075), .ZN(n10074) );
  INV_X1 U10018 ( .A(n10076), .ZN(n10075) );
  NOR2_X1 U10019 ( .A1(n9987), .A2(n9985), .ZN(n10076) );
  NOR2_X1 U10020 ( .A1(n8586), .A2(n8556), .ZN(n9986) );
  NAND2_X1 U10021 ( .A1(n9985), .A2(n9987), .ZN(n10073) );
  NAND2_X1 U10022 ( .A1(n10077), .A2(n10078), .ZN(n9987) );
  NAND2_X1 U10023 ( .A1(n9983), .A2(n10079), .ZN(n10078) );
  INV_X1 U10024 ( .A(n10080), .ZN(n10079) );
  NOR2_X1 U10025 ( .A1(n9982), .A2(n9981), .ZN(n10080) );
  NOR2_X1 U10026 ( .A1(n8586), .A2(n8572), .ZN(n9983) );
  NAND2_X1 U10027 ( .A1(n9981), .A2(n9982), .ZN(n10077) );
  NAND2_X1 U10028 ( .A1(n10081), .A2(n10082), .ZN(n9982) );
  NAND2_X1 U10029 ( .A1(n9979), .A2(n10083), .ZN(n10082) );
  NAND2_X1 U10030 ( .A1(n9978), .A2(n9976), .ZN(n10083) );
  NOR2_X1 U10031 ( .A1(n8586), .A2(n8582), .ZN(n9979) );
  INV_X1 U10032 ( .A(n10084), .ZN(n10081) );
  NOR2_X1 U10033 ( .A1(n9976), .A2(n9978), .ZN(n10084) );
  NOR2_X1 U10034 ( .A1(n10085), .A2(n10086), .ZN(n9978) );
  INV_X1 U10035 ( .A(n10087), .ZN(n10086) );
  NAND2_X1 U10036 ( .A1(n9975), .A2(n10088), .ZN(n10087) );
  NAND2_X1 U10037 ( .A1(n9974), .A2(n9973), .ZN(n10088) );
  NOR2_X1 U10038 ( .A1(n8586), .A2(n8591), .ZN(n9975) );
  NOR2_X1 U10039 ( .A1(n9973), .A2(n9974), .ZN(n10085) );
  NOR2_X1 U10040 ( .A1(n10089), .A2(n10090), .ZN(n9974) );
  INV_X1 U10041 ( .A(n10091), .ZN(n10090) );
  NAND2_X1 U10042 ( .A1(n9971), .A2(n10092), .ZN(n10091) );
  NAND2_X1 U10043 ( .A1(n9970), .A2(n9969), .ZN(n10092) );
  NOR2_X1 U10044 ( .A1(n8586), .A2(n8562), .ZN(n9971) );
  NOR2_X1 U10045 ( .A1(n9969), .A2(n9970), .ZN(n10089) );
  NOR2_X1 U10046 ( .A1(n10093), .A2(n10094), .ZN(n9970) );
  INV_X1 U10047 ( .A(n10095), .ZN(n10094) );
  NAND2_X1 U10048 ( .A1(n9966), .A2(n10096), .ZN(n10095) );
  NAND2_X1 U10049 ( .A1(n9967), .A2(n9965), .ZN(n10096) );
  NOR2_X1 U10050 ( .A1(n8586), .A2(n8545), .ZN(n9966) );
  NOR2_X1 U10051 ( .A1(n9965), .A2(n9967), .ZN(n10093) );
  NOR2_X1 U10052 ( .A1(n10097), .A2(n10098), .ZN(n9967) );
  INV_X1 U10053 ( .A(n10099), .ZN(n10098) );
  NAND2_X1 U10054 ( .A1(n9963), .A2(n10100), .ZN(n10099) );
  NAND2_X1 U10055 ( .A1(n9962), .A2(n9961), .ZN(n10100) );
  NOR2_X1 U10056 ( .A1(n8586), .A2(n8569), .ZN(n9963) );
  NOR2_X1 U10057 ( .A1(n9961), .A2(n9962), .ZN(n10097) );
  NOR2_X1 U10058 ( .A1(n10101), .A2(n10102), .ZN(n9962) );
  INV_X1 U10059 ( .A(n10103), .ZN(n10102) );
  NAND2_X1 U10060 ( .A1(n9958), .A2(n10104), .ZN(n10103) );
  NAND2_X1 U10061 ( .A1(n9959), .A2(n9957), .ZN(n10104) );
  NOR2_X1 U10062 ( .A1(n8586), .A2(n8593), .ZN(n9958) );
  NOR2_X1 U10063 ( .A1(n9957), .A2(n9959), .ZN(n10101) );
  NOR2_X1 U10064 ( .A1(n10105), .A2(n10106), .ZN(n9959) );
  INV_X1 U10065 ( .A(n10107), .ZN(n10106) );
  NAND2_X1 U10066 ( .A1(n9955), .A2(n10108), .ZN(n10107) );
  NAND2_X1 U10067 ( .A1(n9954), .A2(n9953), .ZN(n10108) );
  NOR2_X1 U10068 ( .A1(n8586), .A2(n8583), .ZN(n9955) );
  NOR2_X1 U10069 ( .A1(n9953), .A2(n9954), .ZN(n10105) );
  NOR2_X1 U10070 ( .A1(n10109), .A2(n10110), .ZN(n9954) );
  INV_X1 U10071 ( .A(n10111), .ZN(n10110) );
  NAND2_X1 U10072 ( .A1(n9951), .A2(n10112), .ZN(n10111) );
  NAND2_X1 U10073 ( .A1(n9950), .A2(n9948), .ZN(n10112) );
  NOR2_X1 U10074 ( .A1(n8586), .A2(n8580), .ZN(n9951) );
  NOR2_X1 U10075 ( .A1(n9948), .A2(n9950), .ZN(n10109) );
  NOR2_X1 U10076 ( .A1(n10113), .A2(n10114), .ZN(n9950) );
  INV_X1 U10077 ( .A(n10115), .ZN(n10114) );
  NAND2_X1 U10078 ( .A1(n9947), .A2(n10116), .ZN(n10115) );
  NAND2_X1 U10079 ( .A1(n9946), .A2(n9945), .ZN(n10116) );
  NOR2_X1 U10080 ( .A1(n8586), .A2(n8588), .ZN(n9947) );
  NOR2_X1 U10081 ( .A1(n9945), .A2(n9946), .ZN(n10113) );
  NOR2_X1 U10082 ( .A1(n10117), .A2(n10118), .ZN(n9946) );
  INV_X1 U10083 ( .A(n10119), .ZN(n10118) );
  NAND2_X1 U10084 ( .A1(n9943), .A2(n10120), .ZN(n10119) );
  NAND2_X1 U10085 ( .A1(n9942), .A2(n9940), .ZN(n10120) );
  NOR2_X1 U10086 ( .A1(n8586), .A2(n8551), .ZN(n9943) );
  NOR2_X1 U10087 ( .A1(n9940), .A2(n9942), .ZN(n10117) );
  NOR2_X1 U10088 ( .A1(n10121), .A2(n10122), .ZN(n9942) );
  INV_X1 U10089 ( .A(n10123), .ZN(n10122) );
  NAND2_X1 U10090 ( .A1(n9939), .A2(n10124), .ZN(n10123) );
  NAND2_X1 U10091 ( .A1(n9938), .A2(n9937), .ZN(n10124) );
  NOR2_X1 U10092 ( .A1(n9649), .A2(n8563), .ZN(n9939) );
  NOR2_X1 U10093 ( .A1(n9937), .A2(n9938), .ZN(n10121) );
  NOR2_X1 U10094 ( .A1(n10125), .A2(n10126), .ZN(n9938) );
  INV_X1 U10095 ( .A(n10127), .ZN(n10126) );
  NAND2_X1 U10096 ( .A1(n9935), .A2(n10128), .ZN(n10127) );
  NAND2_X1 U10097 ( .A1(n9934), .A2(n9932), .ZN(n10128) );
  NOR2_X1 U10098 ( .A1(n9649), .A2(n8548), .ZN(n9935) );
  NOR2_X1 U10099 ( .A1(n9932), .A2(n9934), .ZN(n10125) );
  NOR2_X1 U10100 ( .A1(n10129), .A2(n10130), .ZN(n9934) );
  INV_X1 U10101 ( .A(n10131), .ZN(n10130) );
  NAND2_X1 U10102 ( .A1(n9931), .A2(n10132), .ZN(n10131) );
  NAND2_X1 U10103 ( .A1(n9930), .A2(n9929), .ZN(n10132) );
  NOR2_X1 U10104 ( .A1(n9649), .A2(n8584), .ZN(n9931) );
  NOR2_X1 U10105 ( .A1(n9929), .A2(n9930), .ZN(n10129) );
  NOR2_X1 U10106 ( .A1(n10133), .A2(n10134), .ZN(n9930) );
  INV_X1 U10107 ( .A(n10135), .ZN(n10134) );
  NAND2_X1 U10108 ( .A1(n9926), .A2(n10136), .ZN(n10135) );
  NAND2_X1 U10109 ( .A1(n9927), .A2(n9925), .ZN(n10136) );
  NOR2_X1 U10110 ( .A1(n9649), .A2(n8535), .ZN(n9926) );
  NOR2_X1 U10111 ( .A1(n9925), .A2(n9927), .ZN(n10133) );
  NOR2_X1 U10112 ( .A1(n10137), .A2(n10138), .ZN(n9927) );
  INV_X1 U10113 ( .A(n10139), .ZN(n10138) );
  NAND2_X1 U10114 ( .A1(n9923), .A2(n10140), .ZN(n10139) );
  NAND2_X1 U10115 ( .A1(n9922), .A2(n9921), .ZN(n10140) );
  NOR2_X1 U10116 ( .A1(n9649), .A2(n8568), .ZN(n9923) );
  NOR2_X1 U10117 ( .A1(n9921), .A2(n9922), .ZN(n10137) );
  NOR2_X1 U10118 ( .A1(n10141), .A2(n10142), .ZN(n9922) );
  INV_X1 U10119 ( .A(n10143), .ZN(n10142) );
  NAND2_X1 U10120 ( .A1(n9918), .A2(n10144), .ZN(n10143) );
  NAND2_X1 U10121 ( .A1(n9919), .A2(n9917), .ZN(n10144) );
  NOR2_X1 U10122 ( .A1(n9649), .A2(n8574), .ZN(n9918) );
  NOR2_X1 U10123 ( .A1(n9917), .A2(n9919), .ZN(n10141) );
  NOR2_X1 U10124 ( .A1(n10145), .A2(n10146), .ZN(n9919) );
  INV_X1 U10125 ( .A(n10147), .ZN(n10146) );
  NAND2_X1 U10126 ( .A1(n9914), .A2(n10148), .ZN(n10147) );
  NAND2_X1 U10127 ( .A1(n9915), .A2(n9913), .ZN(n10148) );
  NOR2_X1 U10128 ( .A1(n9649), .A2(n8565), .ZN(n9914) );
  NOR2_X1 U10129 ( .A1(n9913), .A2(n9915), .ZN(n10145) );
  NOR2_X1 U10130 ( .A1(n10149), .A2(n10150), .ZN(n9915) );
  INV_X1 U10131 ( .A(n10151), .ZN(n10150) );
  NAND2_X1 U10132 ( .A1(n9908), .A2(n10152), .ZN(n10151) );
  NAND2_X1 U10133 ( .A1(n9911), .A2(n9910), .ZN(n10152) );
  NOR2_X1 U10134 ( .A1(n9649), .A2(n8567), .ZN(n9908) );
  NOR2_X1 U10135 ( .A1(n9910), .A2(n9911), .ZN(n10149) );
  INV_X1 U10136 ( .A(n10153), .ZN(n9911) );
  NAND2_X1 U10137 ( .A1(n10154), .A2(n10155), .ZN(n10153) );
  NAND2_X1 U10138 ( .A1(n9903), .A2(n10156), .ZN(n10155) );
  NAND2_X1 U10139 ( .A1(n8624), .A2(n10157), .ZN(n10156) );
  NAND2_X1 U10140 ( .A1(n8571), .A2(n8585), .ZN(n10157) );
  NAND2_X1 U10141 ( .A1(n10159), .A2(n10160), .ZN(n10154) );
  NAND2_X1 U10142 ( .A1(n8630), .A2(n10161), .ZN(n10160) );
  NAND2_X1 U10143 ( .A1(n8539), .A2(n8542), .ZN(n10161) );
  NAND3_X1 U10144 ( .A1(n9903), .A2(n8537), .A3(n9650), .ZN(n9910) );
  XOR2_X1 U10145 ( .A(n10162), .B(n10163), .Z(n9913) );
  XNOR2_X1 U10146 ( .A(n10164), .B(n10165), .ZN(n10163) );
  XOR2_X1 U10147 ( .A(n10166), .B(n10167), .Z(n9917) );
  XNOR2_X1 U10148 ( .A(n10168), .B(n10169), .ZN(n10166) );
  XOR2_X1 U10149 ( .A(n10170), .B(n10171), .Z(n9921) );
  XNOR2_X1 U10150 ( .A(n10172), .B(n10173), .ZN(n10170) );
  XOR2_X1 U10151 ( .A(n10174), .B(n10175), .Z(n9925) );
  XNOR2_X1 U10152 ( .A(n10176), .B(n10177), .ZN(n10174) );
  XOR2_X1 U10153 ( .A(n10178), .B(n10179), .Z(n9929) );
  XNOR2_X1 U10154 ( .A(n10180), .B(n10181), .ZN(n10178) );
  NOR2_X1 U10155 ( .A1(n8535), .A2(n8542), .ZN(n10181) );
  XOR2_X1 U10156 ( .A(n10182), .B(n10183), .Z(n9932) );
  XNOR2_X1 U10157 ( .A(n10184), .B(n10185), .ZN(n10182) );
  NOR2_X1 U10158 ( .A1(n8584), .A2(n8542), .ZN(n10185) );
  XOR2_X1 U10159 ( .A(n10186), .B(n10187), .Z(n9937) );
  XNOR2_X1 U10160 ( .A(n10188), .B(n10189), .ZN(n10186) );
  NOR2_X1 U10161 ( .A1(n8548), .A2(n8542), .ZN(n10189) );
  XOR2_X1 U10162 ( .A(n10190), .B(n10191), .Z(n9940) );
  XNOR2_X1 U10163 ( .A(n10192), .B(n10193), .ZN(n10190) );
  NOR2_X1 U10164 ( .A1(n8563), .A2(n8542), .ZN(n10193) );
  XOR2_X1 U10165 ( .A(n10194), .B(n10195), .Z(n9945) );
  XNOR2_X1 U10166 ( .A(n10196), .B(n10197), .ZN(n10194) );
  NOR2_X1 U10167 ( .A1(n8551), .A2(n8542), .ZN(n10197) );
  XOR2_X1 U10168 ( .A(n10198), .B(n10199), .Z(n9948) );
  XNOR2_X1 U10169 ( .A(n10200), .B(n10201), .ZN(n10198) );
  NOR2_X1 U10170 ( .A1(n8588), .A2(n8542), .ZN(n10201) );
  XOR2_X1 U10171 ( .A(n10202), .B(n10203), .Z(n9953) );
  XNOR2_X1 U10172 ( .A(n10204), .B(n10205), .ZN(n10202) );
  NOR2_X1 U10173 ( .A1(n8580), .A2(n8542), .ZN(n10205) );
  XOR2_X1 U10174 ( .A(n10206), .B(n10207), .Z(n9957) );
  XNOR2_X1 U10175 ( .A(n10208), .B(n10209), .ZN(n10206) );
  NOR2_X1 U10176 ( .A1(n8583), .A2(n8542), .ZN(n10209) );
  XOR2_X1 U10177 ( .A(n10210), .B(n10211), .Z(n9961) );
  XNOR2_X1 U10178 ( .A(n10212), .B(n10213), .ZN(n10210) );
  NOR2_X1 U10179 ( .A1(n8593), .A2(n8542), .ZN(n10213) );
  XOR2_X1 U10180 ( .A(n10214), .B(n10215), .Z(n9965) );
  XNOR2_X1 U10181 ( .A(n10216), .B(n10217), .ZN(n10214) );
  NOR2_X1 U10182 ( .A1(n8569), .A2(n8542), .ZN(n10217) );
  XNOR2_X1 U10183 ( .A(n10218), .B(n10219), .ZN(n9969) );
  XNOR2_X1 U10184 ( .A(n10220), .B(n10221), .ZN(n10219) );
  NAND2_X1 U10185 ( .A1(n9903), .A2(n10222), .ZN(n10221) );
  XOR2_X1 U10186 ( .A(n10223), .B(n10224), .Z(n9973) );
  XNOR2_X1 U10187 ( .A(n10225), .B(n10226), .ZN(n10223) );
  NOR2_X1 U10188 ( .A1(n8562), .A2(n8542), .ZN(n10226) );
  XOR2_X1 U10189 ( .A(n10227), .B(n10228), .Z(n9976) );
  XNOR2_X1 U10190 ( .A(n10229), .B(n10230), .ZN(n10227) );
  NOR2_X1 U10191 ( .A1(n8591), .A2(n8542), .ZN(n10230) );
  XNOR2_X1 U10192 ( .A(n10231), .B(n10232), .ZN(n9981) );
  XNOR2_X1 U10193 ( .A(n10233), .B(n10234), .ZN(n10231) );
  NOR2_X1 U10194 ( .A1(n8582), .A2(n8542), .ZN(n10234) );
  XNOR2_X1 U10195 ( .A(n10235), .B(n10236), .ZN(n9985) );
  XNOR2_X1 U10196 ( .A(n10237), .B(n10238), .ZN(n10235) );
  NOR2_X1 U10197 ( .A1(n8572), .A2(n8542), .ZN(n10238) );
  XOR2_X1 U10198 ( .A(n10239), .B(n10240), .Z(n9989) );
  XNOR2_X1 U10199 ( .A(n10241), .B(n10242), .ZN(n10239) );
  NOR2_X1 U10200 ( .A1(n8556), .A2(n8542), .ZN(n10242) );
  XOR2_X1 U10201 ( .A(n10243), .B(n10244), .Z(n9992) );
  XNOR2_X1 U10202 ( .A(n10245), .B(n10246), .ZN(n10243) );
  NOR2_X1 U10203 ( .A1(n8594), .A2(n8542), .ZN(n10246) );
  XNOR2_X1 U10204 ( .A(n10247), .B(n10248), .ZN(n9997) );
  XNOR2_X1 U10205 ( .A(n10249), .B(n10250), .ZN(n10247) );
  NOR2_X1 U10206 ( .A1(n8560), .A2(n8542), .ZN(n10250) );
  INV_X1 U10207 ( .A(n10251), .ZN(n10057) );
  NOR2_X1 U10208 ( .A1(n10003), .A2(n10000), .ZN(n10251) );
  XNOR2_X1 U10209 ( .A(n10252), .B(n10253), .ZN(n10000) );
  XOR2_X1 U10210 ( .A(n10254), .B(n10255), .Z(n10252) );
  NOR2_X1 U10211 ( .A1(n8544), .A2(n8542), .ZN(n10255) );
  NAND2_X1 U10212 ( .A1(n9650), .A2(n9286), .ZN(n10003) );
  INV_X1 U10213 ( .A(n9649), .ZN(n9650) );
  XNOR2_X1 U10214 ( .A(n10256), .B(n10257), .ZN(n9649) );
  XOR2_X1 U10215 ( .A(d_27_), .B(c_27_), .Z(n10257) );
  XNOR2_X1 U10216 ( .A(n10258), .B(n10259), .ZN(n10005) );
  XNOR2_X1 U10217 ( .A(n10260), .B(n10261), .ZN(n10258) );
  XNOR2_X1 U10218 ( .A(n10262), .B(n10263), .ZN(n10009) );
  XOR2_X1 U10219 ( .A(n10264), .B(n10265), .Z(n10263) );
  NOR2_X1 U10220 ( .A1(n8564), .A2(n8542), .ZN(n10265) );
  XNOR2_X1 U10221 ( .A(n10266), .B(n10267), .ZN(n10013) );
  XNOR2_X1 U10222 ( .A(n10268), .B(n10269), .ZN(n10267) );
  NAND2_X1 U10223 ( .A1(n9903), .A2(n9277), .ZN(n10269) );
  XOR2_X1 U10224 ( .A(n10270), .B(n10271), .Z(n10021) );
  XNOR2_X1 U10225 ( .A(n10272), .B(n10273), .ZN(n10270) );
  XNOR2_X1 U10226 ( .A(n10274), .B(n10275), .ZN(n10024) );
  XOR2_X1 U10227 ( .A(n10276), .B(n10277), .Z(n10274) );
  NOR2_X1 U10228 ( .A1(n8589), .A2(n8542), .ZN(n10277) );
  XNOR2_X1 U10229 ( .A(n10278), .B(n10279), .ZN(n9776) );
  XNOR2_X1 U10230 ( .A(n10280), .B(n10281), .ZN(n10279) );
  NAND2_X1 U10231 ( .A1(n9903), .A2(n8592), .ZN(n10281) );
  NAND4_X1 U10232 ( .A1(n8950), .A2(n8949), .A3(n8951), .A4(n8943), .ZN(n8802)
         );
  INV_X1 U10233 ( .A(n10282), .ZN(n8943) );
  NAND2_X1 U10234 ( .A1(n10283), .A2(n10284), .ZN(n8951) );
  NAND3_X1 U10235 ( .A1(n8592), .A2(n10285), .A3(n9903), .ZN(n10284) );
  NAND2_X1 U10236 ( .A1(n10280), .A2(n10278), .ZN(n10285) );
  INV_X1 U10237 ( .A(n10286), .ZN(n10283) );
  NOR2_X1 U10238 ( .A1(n10278), .A2(n10280), .ZN(n10286) );
  NOR2_X1 U10239 ( .A1(n10287), .A2(n10288), .ZN(n10280) );
  NOR3_X1 U10240 ( .A1(n8884), .A2(n10289), .A3(n8542), .ZN(n10288) );
  NOR2_X1 U10241 ( .A1(n10276), .A2(n10275), .ZN(n10289) );
  INV_X1 U10242 ( .A(n10290), .ZN(n10287) );
  NAND2_X1 U10243 ( .A1(n10275), .A2(n10276), .ZN(n10290) );
  NAND2_X1 U10244 ( .A1(n10291), .A2(n10292), .ZN(n10276) );
  NAND2_X1 U10245 ( .A1(n10273), .A2(n10293), .ZN(n10292) );
  NAND2_X1 U10246 ( .A1(n10272), .A2(n10294), .ZN(n10293) );
  INV_X1 U10247 ( .A(n10271), .ZN(n10294) );
  NOR2_X1 U10248 ( .A1(n8542), .A2(n8552), .ZN(n10273) );
  NAND2_X1 U10249 ( .A1(n10271), .A2(n10295), .ZN(n10291) );
  INV_X1 U10250 ( .A(n10272), .ZN(n10295) );
  NOR2_X1 U10251 ( .A1(n10296), .A2(n10297), .ZN(n10272) );
  NOR2_X1 U10252 ( .A1(n10042), .A2(n10298), .ZN(n10297) );
  NOR2_X1 U10253 ( .A1(n10041), .A2(n10039), .ZN(n10298) );
  NAND2_X1 U10254 ( .A1(n9903), .A2(n9792), .ZN(n10042) );
  INV_X1 U10255 ( .A(n10299), .ZN(n10296) );
  NAND2_X1 U10256 ( .A1(n10039), .A2(n10041), .ZN(n10299) );
  NAND2_X1 U10257 ( .A1(n10300), .A2(n10301), .ZN(n10041) );
  NAND3_X1 U10258 ( .A1(n9277), .A2(n10302), .A3(n9903), .ZN(n10301) );
  NAND2_X1 U10259 ( .A1(n10268), .A2(n10266), .ZN(n10302) );
  INV_X1 U10260 ( .A(n10303), .ZN(n10300) );
  NOR2_X1 U10261 ( .A1(n10266), .A2(n10268), .ZN(n10303) );
  NOR2_X1 U10262 ( .A1(n10304), .A2(n10305), .ZN(n10268) );
  INV_X1 U10263 ( .A(n10306), .ZN(n10305) );
  NAND3_X1 U10264 ( .A1(n10307), .A2(n10308), .A3(n9903), .ZN(n10306) );
  NAND2_X1 U10265 ( .A1(n10264), .A2(n10262), .ZN(n10308) );
  NOR2_X1 U10266 ( .A1(n10262), .A2(n10264), .ZN(n10304) );
  NOR2_X1 U10267 ( .A1(n10309), .A2(n10310), .ZN(n10264) );
  INV_X1 U10268 ( .A(n10311), .ZN(n10310) );
  NAND2_X1 U10269 ( .A1(n10260), .A2(n10312), .ZN(n10311) );
  NAND2_X1 U10270 ( .A1(n10259), .A2(n10261), .ZN(n10312) );
  NAND2_X1 U10271 ( .A1(n10313), .A2(n10314), .ZN(n10260) );
  INV_X1 U10272 ( .A(n10315), .ZN(n10314) );
  NOR3_X1 U10273 ( .A1(n8544), .A2(n10316), .A3(n8542), .ZN(n10315) );
  NOR2_X1 U10274 ( .A1(n10254), .A2(n10253), .ZN(n10316) );
  NAND2_X1 U10275 ( .A1(n10253), .A2(n10254), .ZN(n10313) );
  NAND2_X1 U10276 ( .A1(n10317), .A2(n10318), .ZN(n10254) );
  NAND3_X1 U10277 ( .A1(n9295), .A2(n10319), .A3(n9903), .ZN(n10318) );
  NAND2_X1 U10278 ( .A1(n10249), .A2(n10248), .ZN(n10319) );
  INV_X1 U10279 ( .A(n10320), .ZN(n10317) );
  NOR2_X1 U10280 ( .A1(n10248), .A2(n10249), .ZN(n10320) );
  NOR2_X1 U10281 ( .A1(n10321), .A2(n10322), .ZN(n10249) );
  NOR3_X1 U10282 ( .A1(n9014), .A2(n10323), .A3(n8542), .ZN(n10322) );
  INV_X1 U10283 ( .A(n10324), .ZN(n10323) );
  NAND2_X1 U10284 ( .A1(n10245), .A2(n10244), .ZN(n10324) );
  NOR2_X1 U10285 ( .A1(n10244), .A2(n10245), .ZN(n10321) );
  NOR2_X1 U10286 ( .A1(n10325), .A2(n10326), .ZN(n10245) );
  INV_X1 U10287 ( .A(n10327), .ZN(n10326) );
  NAND3_X1 U10288 ( .A1(n9304), .A2(n10328), .A3(n9903), .ZN(n10327) );
  NAND2_X1 U10289 ( .A1(n10241), .A2(n10240), .ZN(n10328) );
  NOR2_X1 U10290 ( .A1(n10240), .A2(n10241), .ZN(n10325) );
  NOR2_X1 U10291 ( .A1(n10329), .A2(n10330), .ZN(n10241) );
  NOR3_X1 U10292 ( .A1(n9025), .A2(n10331), .A3(n8542), .ZN(n10330) );
  INV_X1 U10293 ( .A(n10332), .ZN(n10331) );
  NAND2_X1 U10294 ( .A1(n10237), .A2(n10236), .ZN(n10332) );
  NOR2_X1 U10295 ( .A1(n10236), .A2(n10237), .ZN(n10329) );
  NOR2_X1 U10296 ( .A1(n10333), .A2(n10334), .ZN(n10237) );
  INV_X1 U10297 ( .A(n10335), .ZN(n10334) );
  NAND3_X1 U10298 ( .A1(n9313), .A2(n10336), .A3(n9903), .ZN(n10335) );
  NAND2_X1 U10299 ( .A1(n10233), .A2(n10232), .ZN(n10336) );
  NOR2_X1 U10300 ( .A1(n10232), .A2(n10233), .ZN(n10333) );
  NOR2_X1 U10301 ( .A1(n10337), .A2(n10338), .ZN(n10233) );
  NOR3_X1 U10302 ( .A1(n9036), .A2(n10339), .A3(n8542), .ZN(n10338) );
  INV_X1 U10303 ( .A(n10340), .ZN(n10339) );
  NAND2_X1 U10304 ( .A1(n10229), .A2(n10228), .ZN(n10340) );
  NOR2_X1 U10305 ( .A1(n10228), .A2(n10229), .ZN(n10337) );
  NOR2_X1 U10306 ( .A1(n10341), .A2(n10342), .ZN(n10229) );
  INV_X1 U10307 ( .A(n10343), .ZN(n10342) );
  NAND3_X1 U10308 ( .A1(n9322), .A2(n10344), .A3(n9903), .ZN(n10343) );
  NAND2_X1 U10309 ( .A1(n10225), .A2(n10224), .ZN(n10344) );
  NOR2_X1 U10310 ( .A1(n10224), .A2(n10225), .ZN(n10341) );
  NOR2_X1 U10311 ( .A1(n10345), .A2(n10346), .ZN(n10225) );
  NOR3_X1 U10312 ( .A1(n8545), .A2(n10347), .A3(n8542), .ZN(n10346) );
  INV_X1 U10313 ( .A(n10348), .ZN(n10347) );
  NAND2_X1 U10314 ( .A1(n10220), .A2(n10218), .ZN(n10348) );
  NOR2_X1 U10315 ( .A1(n10218), .A2(n10220), .ZN(n10345) );
  NOR2_X1 U10316 ( .A1(n10349), .A2(n10350), .ZN(n10220) );
  INV_X1 U10317 ( .A(n10351), .ZN(n10350) );
  NAND3_X1 U10318 ( .A1(n9331), .A2(n10352), .A3(n9903), .ZN(n10351) );
  NAND2_X1 U10319 ( .A1(n10216), .A2(n10215), .ZN(n10352) );
  NOR2_X1 U10320 ( .A1(n10215), .A2(n10216), .ZN(n10349) );
  NOR2_X1 U10321 ( .A1(n10353), .A2(n10354), .ZN(n10216) );
  NOR3_X1 U10322 ( .A1(n9056), .A2(n10355), .A3(n8542), .ZN(n10354) );
  INV_X1 U10323 ( .A(n10356), .ZN(n10355) );
  NAND2_X1 U10324 ( .A1(n10212), .A2(n10211), .ZN(n10356) );
  NOR2_X1 U10325 ( .A1(n10211), .A2(n10212), .ZN(n10353) );
  NOR2_X1 U10326 ( .A1(n10357), .A2(n10358), .ZN(n10212) );
  INV_X1 U10327 ( .A(n10359), .ZN(n10358) );
  NAND3_X1 U10328 ( .A1(n9340), .A2(n10360), .A3(n9903), .ZN(n10359) );
  NAND2_X1 U10329 ( .A1(n10208), .A2(n10207), .ZN(n10360) );
  NOR2_X1 U10330 ( .A1(n10207), .A2(n10208), .ZN(n10357) );
  NOR2_X1 U10331 ( .A1(n10361), .A2(n10362), .ZN(n10208) );
  NOR3_X1 U10332 ( .A1(n8580), .A2(n10363), .A3(n8542), .ZN(n10362) );
  INV_X1 U10333 ( .A(n10364), .ZN(n10363) );
  NAND2_X1 U10334 ( .A1(n10204), .A2(n10203), .ZN(n10364) );
  NOR2_X1 U10335 ( .A1(n10203), .A2(n10204), .ZN(n10361) );
  NOR2_X1 U10336 ( .A1(n10365), .A2(n10366), .ZN(n10204) );
  INV_X1 U10337 ( .A(n10367), .ZN(n10366) );
  NAND3_X1 U10338 ( .A1(n9080), .A2(n10368), .A3(n9903), .ZN(n10367) );
  NAND2_X1 U10339 ( .A1(n10200), .A2(n10199), .ZN(n10368) );
  NOR2_X1 U10340 ( .A1(n10199), .A2(n10200), .ZN(n10365) );
  NOR2_X1 U10341 ( .A1(n10369), .A2(n10370), .ZN(n10200) );
  NOR3_X1 U10342 ( .A1(n8551), .A2(n10371), .A3(n8542), .ZN(n10370) );
  INV_X1 U10343 ( .A(n10372), .ZN(n10371) );
  NAND2_X1 U10344 ( .A1(n10196), .A2(n10195), .ZN(n10372) );
  NOR2_X1 U10345 ( .A1(n10195), .A2(n10196), .ZN(n10369) );
  NOR2_X1 U10346 ( .A1(n10373), .A2(n10374), .ZN(n10196) );
  INV_X1 U10347 ( .A(n10375), .ZN(n10374) );
  NAND3_X1 U10348 ( .A1(n9098), .A2(n10376), .A3(n9903), .ZN(n10375) );
  NAND2_X1 U10349 ( .A1(n10192), .A2(n10191), .ZN(n10376) );
  NOR2_X1 U10350 ( .A1(n10191), .A2(n10192), .ZN(n10373) );
  NOR2_X1 U10351 ( .A1(n10377), .A2(n10378), .ZN(n10192) );
  NOR3_X1 U10352 ( .A1(n8548), .A2(n10379), .A3(n8542), .ZN(n10378) );
  INV_X1 U10353 ( .A(n10380), .ZN(n10379) );
  NAND2_X1 U10354 ( .A1(n10188), .A2(n10187), .ZN(n10380) );
  NOR2_X1 U10355 ( .A1(n10187), .A2(n10188), .ZN(n10377) );
  NOR2_X1 U10356 ( .A1(n10381), .A2(n10382), .ZN(n10188) );
  INV_X1 U10357 ( .A(n10383), .ZN(n10382) );
  NAND3_X1 U10358 ( .A1(n9112), .A2(n10384), .A3(n9903), .ZN(n10383) );
  NAND2_X1 U10359 ( .A1(n10184), .A2(n10183), .ZN(n10384) );
  NOR2_X1 U10360 ( .A1(n10183), .A2(n10184), .ZN(n10381) );
  NOR2_X1 U10361 ( .A1(n10385), .A2(n10386), .ZN(n10184) );
  INV_X1 U10362 ( .A(n10387), .ZN(n10386) );
  NAND3_X1 U10363 ( .A1(n9121), .A2(n10388), .A3(n9903), .ZN(n10387) );
  NAND2_X1 U10364 ( .A1(n10180), .A2(n10179), .ZN(n10388) );
  NOR2_X1 U10365 ( .A1(n10179), .A2(n10180), .ZN(n10385) );
  NOR2_X1 U10366 ( .A1(n10389), .A2(n10390), .ZN(n10180) );
  INV_X1 U10367 ( .A(n10391), .ZN(n10390) );
  NAND2_X1 U10368 ( .A1(n10176), .A2(n10392), .ZN(n10391) );
  NAND2_X1 U10369 ( .A1(n10177), .A2(n10175), .ZN(n10392) );
  NOR2_X1 U10370 ( .A1(n8542), .A2(n8568), .ZN(n10176) );
  NOR2_X1 U10371 ( .A1(n10175), .A2(n10177), .ZN(n10389) );
  NOR2_X1 U10372 ( .A1(n10393), .A2(n10394), .ZN(n10177) );
  INV_X1 U10373 ( .A(n10395), .ZN(n10394) );
  NAND2_X1 U10374 ( .A1(n10172), .A2(n10396), .ZN(n10395) );
  NAND2_X1 U10375 ( .A1(n10173), .A2(n10171), .ZN(n10396) );
  NOR2_X1 U10376 ( .A1(n8542), .A2(n8574), .ZN(n10172) );
  NOR2_X1 U10377 ( .A1(n10171), .A2(n10173), .ZN(n10393) );
  NOR2_X1 U10378 ( .A1(n10397), .A2(n10398), .ZN(n10173) );
  INV_X1 U10379 ( .A(n10399), .ZN(n10398) );
  NAND2_X1 U10380 ( .A1(n10168), .A2(n10400), .ZN(n10399) );
  NAND2_X1 U10381 ( .A1(n10169), .A2(n10167), .ZN(n10400) );
  NOR2_X1 U10382 ( .A1(n8542), .A2(n8565), .ZN(n10168) );
  NOR2_X1 U10383 ( .A1(n10167), .A2(n10169), .ZN(n10397) );
  NOR2_X1 U10384 ( .A1(n10401), .A2(n10402), .ZN(n10169) );
  INV_X1 U10385 ( .A(n10403), .ZN(n10402) );
  NAND2_X1 U10386 ( .A1(n10162), .A2(n10404), .ZN(n10403) );
  NAND2_X1 U10387 ( .A1(n10165), .A2(n10164), .ZN(n10404) );
  NOR2_X1 U10388 ( .A1(n8542), .A2(n8567), .ZN(n10162) );
  NOR2_X1 U10389 ( .A1(n10164), .A2(n10165), .ZN(n10401) );
  INV_X1 U10390 ( .A(n10405), .ZN(n10165) );
  NAND2_X1 U10391 ( .A1(n10406), .A2(n10407), .ZN(n10405) );
  NAND2_X1 U10392 ( .A1(n10159), .A2(n10408), .ZN(n10407) );
  NAND2_X1 U10393 ( .A1(n8624), .A2(n10409), .ZN(n10408) );
  NAND2_X1 U10394 ( .A1(n8541), .A2(n8585), .ZN(n10409) );
  NAND2_X1 U10395 ( .A1(n8540), .A2(n10411), .ZN(n10406) );
  NAND2_X1 U10396 ( .A1(n8630), .A2(n10412), .ZN(n10411) );
  NAND2_X1 U10397 ( .A1(n8539), .A2(n8571), .ZN(n10412) );
  NAND3_X1 U10398 ( .A1(n10159), .A2(n8537), .A3(n9903), .ZN(n10164) );
  XOR2_X1 U10399 ( .A(n10413), .B(n10414), .Z(n10167) );
  XNOR2_X1 U10400 ( .A(n10415), .B(n10416), .ZN(n10414) );
  XOR2_X1 U10401 ( .A(n10417), .B(n10418), .Z(n10171) );
  XNOR2_X1 U10402 ( .A(n10419), .B(n10420), .ZN(n10417) );
  XOR2_X1 U10403 ( .A(n10421), .B(n10422), .Z(n10175) );
  XNOR2_X1 U10404 ( .A(n10423), .B(n10424), .ZN(n10421) );
  XOR2_X1 U10405 ( .A(n10425), .B(n10426), .Z(n10179) );
  XNOR2_X1 U10406 ( .A(n10427), .B(n10428), .ZN(n10425) );
  XOR2_X1 U10407 ( .A(n10429), .B(n10430), .Z(n10183) );
  XNOR2_X1 U10408 ( .A(n10431), .B(n10432), .ZN(n10429) );
  XOR2_X1 U10409 ( .A(n10433), .B(n10434), .Z(n10187) );
  XNOR2_X1 U10410 ( .A(n10435), .B(n10436), .ZN(n10433) );
  XNOR2_X1 U10411 ( .A(n10437), .B(n10438), .ZN(n10191) );
  XOR2_X1 U10412 ( .A(n10439), .B(n10440), .Z(n10438) );
  XOR2_X1 U10413 ( .A(n10441), .B(n10442), .Z(n10195) );
  XNOR2_X1 U10414 ( .A(n10443), .B(n10444), .ZN(n10441) );
  XNOR2_X1 U10415 ( .A(n10445), .B(n10446), .ZN(n10199) );
  XOR2_X1 U10416 ( .A(n10447), .B(n10448), .Z(n10446) );
  XOR2_X1 U10417 ( .A(n10449), .B(n10450), .Z(n10203) );
  XNOR2_X1 U10418 ( .A(n10451), .B(n10452), .ZN(n10449) );
  XOR2_X1 U10419 ( .A(n10453), .B(n10454), .Z(n10207) );
  XNOR2_X1 U10420 ( .A(n10455), .B(n10456), .ZN(n10453) );
  XOR2_X1 U10421 ( .A(n10457), .B(n10458), .Z(n10211) );
  XNOR2_X1 U10422 ( .A(n10459), .B(n10460), .ZN(n10457) );
  XOR2_X1 U10423 ( .A(n10461), .B(n10462), .Z(n10215) );
  XNOR2_X1 U10424 ( .A(n10463), .B(n10464), .ZN(n10461) );
  XOR2_X1 U10425 ( .A(n10465), .B(n10466), .Z(n10218) );
  XNOR2_X1 U10426 ( .A(n10467), .B(n10468), .ZN(n10465) );
  XOR2_X1 U10427 ( .A(n10469), .B(n10470), .Z(n10224) );
  XNOR2_X1 U10428 ( .A(n10471), .B(n10472), .ZN(n10469) );
  XNOR2_X1 U10429 ( .A(n10473), .B(n10474), .ZN(n10228) );
  XOR2_X1 U10430 ( .A(n10475), .B(n10476), .Z(n10474) );
  XNOR2_X1 U10431 ( .A(n10477), .B(n10478), .ZN(n10232) );
  XOR2_X1 U10432 ( .A(n10479), .B(n10480), .Z(n10477) );
  XNOR2_X1 U10433 ( .A(n10481), .B(n10482), .ZN(n10236) );
  XOR2_X1 U10434 ( .A(n10483), .B(n10484), .Z(n10481) );
  XNOR2_X1 U10435 ( .A(n10485), .B(n10486), .ZN(n10240) );
  XOR2_X1 U10436 ( .A(n10487), .B(n10488), .Z(n10485) );
  NOR2_X1 U10437 ( .A1(n8572), .A2(n8571), .ZN(n10488) );
  XNOR2_X1 U10438 ( .A(n10489), .B(n10490), .ZN(n10244) );
  XOR2_X1 U10439 ( .A(n10491), .B(n10492), .Z(n10490) );
  XNOR2_X1 U10440 ( .A(n10493), .B(n10494), .ZN(n10248) );
  XOR2_X1 U10441 ( .A(n10495), .B(n10496), .Z(n10493) );
  XOR2_X1 U10442 ( .A(n10497), .B(n10498), .Z(n10253) );
  XOR2_X1 U10443 ( .A(n10499), .B(n10500), .Z(n10497) );
  NOR2_X1 U10444 ( .A1(n10261), .A2(n10259), .ZN(n10309) );
  XNOR2_X1 U10445 ( .A(n10501), .B(n10502), .ZN(n10259) );
  XOR2_X1 U10446 ( .A(n10503), .B(n10504), .Z(n10501) );
  NOR2_X1 U10447 ( .A1(n8544), .A2(n8571), .ZN(n10504) );
  NAND2_X1 U10448 ( .A1(n9903), .A2(n9286), .ZN(n10261) );
  INV_X1 U10449 ( .A(n8542), .ZN(n9903) );
  XOR2_X1 U10450 ( .A(d_26_), .B(c_26_), .Z(n10506) );
  XNOR2_X1 U10451 ( .A(n10507), .B(n10508), .ZN(n10262) );
  XOR2_X1 U10452 ( .A(n10509), .B(n10510), .Z(n10508) );
  XOR2_X1 U10453 ( .A(n10511), .B(n10512), .Z(n10266) );
  XNOR2_X1 U10454 ( .A(n10513), .B(n10514), .ZN(n10511) );
  XNOR2_X1 U10455 ( .A(n10515), .B(n10516), .ZN(n10039) );
  NAND2_X1 U10456 ( .A1(n10517), .A2(n10518), .ZN(n10515) );
  XOR2_X1 U10457 ( .A(n10519), .B(n10520), .Z(n10271) );
  XOR2_X1 U10458 ( .A(n10521), .B(n10522), .Z(n10519) );
  NOR2_X1 U10459 ( .A1(n8527), .A2(n8571), .ZN(n10522) );
  XNOR2_X1 U10460 ( .A(n10523), .B(n10524), .ZN(n10275) );
  XOR2_X1 U10461 ( .A(n10525), .B(n10526), .Z(n10524) );
  NAND2_X1 U10462 ( .A1(n10159), .A2(n9268), .ZN(n10526) );
  XNOR2_X1 U10463 ( .A(n10527), .B(n10528), .ZN(n10278) );
  XOR2_X1 U10464 ( .A(n10529), .B(n10530), .Z(n10527) );
  NOR2_X1 U10465 ( .A1(n8589), .A2(n8571), .ZN(n10530) );
  NAND2_X1 U10466 ( .A1(n10531), .A2(n10532), .ZN(n8949) );
  XOR2_X1 U10467 ( .A(n10533), .B(n10534), .Z(n8950) );
  XOR2_X1 U10468 ( .A(n10535), .B(n10536), .Z(n10533) );
  NOR2_X1 U10469 ( .A1(n8972), .A2(n8571), .ZN(n10536) );
  NAND3_X1 U10470 ( .A1(n10537), .A2(n8940), .A3(n10282), .ZN(n8806) );
  NOR2_X1 U10471 ( .A1(n10532), .A2(n10531), .ZN(n10282) );
  NOR2_X1 U10472 ( .A1(n10538), .A2(n10539), .ZN(n10531) );
  NOR3_X1 U10473 ( .A1(n8972), .A2(n10540), .A3(n8571), .ZN(n10539) );
  NOR2_X1 U10474 ( .A1(n10535), .A2(n10534), .ZN(n10540) );
  INV_X1 U10475 ( .A(n10541), .ZN(n10538) );
  NAND2_X1 U10476 ( .A1(n10534), .A2(n10535), .ZN(n10541) );
  NAND2_X1 U10477 ( .A1(n10542), .A2(n10543), .ZN(n10535) );
  NAND3_X1 U10478 ( .A1(n9263), .A2(n10544), .A3(n10159), .ZN(n10543) );
  INV_X1 U10479 ( .A(n10545), .ZN(n10544) );
  NOR2_X1 U10480 ( .A1(n10529), .A2(n10528), .ZN(n10545) );
  NAND2_X1 U10481 ( .A1(n10528), .A2(n10529), .ZN(n10542) );
  NAND2_X1 U10482 ( .A1(n10546), .A2(n10547), .ZN(n10529) );
  NAND3_X1 U10483 ( .A1(n9268), .A2(n10548), .A3(n10159), .ZN(n10547) );
  INV_X1 U10484 ( .A(n10549), .ZN(n10548) );
  NOR2_X1 U10485 ( .A1(n10525), .A2(n10523), .ZN(n10549) );
  NAND2_X1 U10486 ( .A1(n10523), .A2(n10525), .ZN(n10546) );
  NAND2_X1 U10487 ( .A1(n10550), .A2(n10551), .ZN(n10525) );
  NAND3_X1 U10488 ( .A1(n9792), .A2(n10552), .A3(n10159), .ZN(n10551) );
  INV_X1 U10489 ( .A(n10553), .ZN(n10552) );
  NOR2_X1 U10490 ( .A1(n10521), .A2(n10520), .ZN(n10553) );
  NAND2_X1 U10491 ( .A1(n10520), .A2(n10521), .ZN(n10550) );
  NAND2_X1 U10492 ( .A1(n10517), .A2(n10554), .ZN(n10521) );
  NAND2_X1 U10493 ( .A1(n10516), .A2(n10518), .ZN(n10554) );
  NAND2_X1 U10494 ( .A1(n10555), .A2(n10556), .ZN(n10518) );
  NAND2_X1 U10495 ( .A1(n10159), .A2(n9277), .ZN(n10556) );
  XNOR2_X1 U10496 ( .A(n10557), .B(n10558), .ZN(n10516) );
  XOR2_X1 U10497 ( .A(n10559), .B(n10560), .Z(n10557) );
  NAND2_X1 U10498 ( .A1(n8540), .A2(n10307), .ZN(n10559) );
  NAND2_X1 U10499 ( .A1(n9277), .A2(n10561), .ZN(n10517) );
  INV_X1 U10500 ( .A(n10555), .ZN(n10561) );
  NOR2_X1 U10501 ( .A1(n10562), .A2(n10563), .ZN(n10555) );
  INV_X1 U10502 ( .A(n10564), .ZN(n10563) );
  NAND2_X1 U10503 ( .A1(n10514), .A2(n10565), .ZN(n10564) );
  NAND2_X1 U10504 ( .A1(n10513), .A2(n10512), .ZN(n10565) );
  NOR2_X1 U10505 ( .A1(n8571), .A2(n8564), .ZN(n10514) );
  NOR2_X1 U10506 ( .A1(n10512), .A2(n10513), .ZN(n10562) );
  NOR2_X1 U10507 ( .A1(n10566), .A2(n10567), .ZN(n10513) );
  INV_X1 U10508 ( .A(n10568), .ZN(n10567) );
  NAND2_X1 U10509 ( .A1(n10509), .A2(n10569), .ZN(n10568) );
  NAND2_X1 U10510 ( .A1(n10507), .A2(n10510), .ZN(n10569) );
  NAND2_X1 U10511 ( .A1(n10570), .A2(n10571), .ZN(n10509) );
  INV_X1 U10512 ( .A(n10572), .ZN(n10571) );
  NOR3_X1 U10513 ( .A1(n8544), .A2(n10573), .A3(n8571), .ZN(n10572) );
  NOR2_X1 U10514 ( .A1(n10503), .A2(n10502), .ZN(n10573) );
  NAND2_X1 U10515 ( .A1(n10502), .A2(n10503), .ZN(n10570) );
  NAND2_X1 U10516 ( .A1(n10574), .A2(n10575), .ZN(n10503) );
  NAND2_X1 U10517 ( .A1(n10499), .A2(n10576), .ZN(n10575) );
  INV_X1 U10518 ( .A(n10577), .ZN(n10576) );
  NOR2_X1 U10519 ( .A1(n10500), .A2(n10498), .ZN(n10577) );
  NOR2_X1 U10520 ( .A1(n8571), .A2(n8560), .ZN(n10499) );
  NAND2_X1 U10521 ( .A1(n10498), .A2(n10500), .ZN(n10574) );
  NAND2_X1 U10522 ( .A1(n10578), .A2(n10579), .ZN(n10500) );
  NAND2_X1 U10523 ( .A1(n10496), .A2(n10580), .ZN(n10579) );
  INV_X1 U10524 ( .A(n10581), .ZN(n10580) );
  NOR2_X1 U10525 ( .A1(n10495), .A2(n10494), .ZN(n10581) );
  NOR2_X1 U10526 ( .A1(n8571), .A2(n8594), .ZN(n10496) );
  NAND2_X1 U10527 ( .A1(n10494), .A2(n10495), .ZN(n10578) );
  NAND2_X1 U10528 ( .A1(n10582), .A2(n10583), .ZN(n10495) );
  NAND2_X1 U10529 ( .A1(n10491), .A2(n10584), .ZN(n10583) );
  NAND2_X1 U10530 ( .A1(n10489), .A2(n10492), .ZN(n10584) );
  NAND2_X1 U10531 ( .A1(n10585), .A2(n10586), .ZN(n10491) );
  INV_X1 U10532 ( .A(n10587), .ZN(n10586) );
  NOR3_X1 U10533 ( .A1(n9025), .A2(n10588), .A3(n8571), .ZN(n10587) );
  NOR2_X1 U10534 ( .A1(n10487), .A2(n10486), .ZN(n10588) );
  NAND2_X1 U10535 ( .A1(n10486), .A2(n10487), .ZN(n10585) );
  NAND2_X1 U10536 ( .A1(n10589), .A2(n10590), .ZN(n10487) );
  NAND2_X1 U10537 ( .A1(n10483), .A2(n10591), .ZN(n10590) );
  INV_X1 U10538 ( .A(n10592), .ZN(n10591) );
  NOR2_X1 U10539 ( .A1(n10484), .A2(n10482), .ZN(n10592) );
  NOR2_X1 U10540 ( .A1(n8571), .A2(n8582), .ZN(n10483) );
  NAND2_X1 U10541 ( .A1(n10482), .A2(n10484), .ZN(n10589) );
  NAND2_X1 U10542 ( .A1(n10593), .A2(n10594), .ZN(n10484) );
  NAND2_X1 U10543 ( .A1(n10480), .A2(n10595), .ZN(n10594) );
  INV_X1 U10544 ( .A(n10596), .ZN(n10595) );
  NOR2_X1 U10545 ( .A1(n10479), .A2(n10478), .ZN(n10596) );
  NOR2_X1 U10546 ( .A1(n8571), .A2(n8591), .ZN(n10480) );
  NAND2_X1 U10547 ( .A1(n10478), .A2(n10479), .ZN(n10593) );
  NAND2_X1 U10548 ( .A1(n10597), .A2(n10598), .ZN(n10479) );
  NAND2_X1 U10549 ( .A1(n10476), .A2(n10599), .ZN(n10598) );
  NAND2_X1 U10550 ( .A1(n10475), .A2(n10473), .ZN(n10599) );
  NOR2_X1 U10551 ( .A1(n8571), .A2(n8562), .ZN(n10476) );
  INV_X1 U10552 ( .A(n10600), .ZN(n10597) );
  NOR2_X1 U10553 ( .A1(n10473), .A2(n10475), .ZN(n10600) );
  NOR2_X1 U10554 ( .A1(n10601), .A2(n10602), .ZN(n10475) );
  INV_X1 U10555 ( .A(n10603), .ZN(n10602) );
  NAND2_X1 U10556 ( .A1(n10472), .A2(n10604), .ZN(n10603) );
  NAND2_X1 U10557 ( .A1(n10471), .A2(n10470), .ZN(n10604) );
  NOR2_X1 U10558 ( .A1(n8571), .A2(n8545), .ZN(n10472) );
  NOR2_X1 U10559 ( .A1(n10470), .A2(n10471), .ZN(n10601) );
  NOR2_X1 U10560 ( .A1(n10605), .A2(n10606), .ZN(n10471) );
  INV_X1 U10561 ( .A(n10607), .ZN(n10606) );
  NAND2_X1 U10562 ( .A1(n10468), .A2(n10608), .ZN(n10607) );
  NAND2_X1 U10563 ( .A1(n10467), .A2(n10466), .ZN(n10608) );
  NOR2_X1 U10564 ( .A1(n8571), .A2(n8569), .ZN(n10468) );
  NOR2_X1 U10565 ( .A1(n10466), .A2(n10467), .ZN(n10605) );
  NOR2_X1 U10566 ( .A1(n10609), .A2(n10610), .ZN(n10467) );
  INV_X1 U10567 ( .A(n10611), .ZN(n10610) );
  NAND2_X1 U10568 ( .A1(n10463), .A2(n10612), .ZN(n10611) );
  NAND2_X1 U10569 ( .A1(n10464), .A2(n10462), .ZN(n10612) );
  NOR2_X1 U10570 ( .A1(n8571), .A2(n8593), .ZN(n10463) );
  NOR2_X1 U10571 ( .A1(n10462), .A2(n10464), .ZN(n10609) );
  NOR2_X1 U10572 ( .A1(n10613), .A2(n10614), .ZN(n10464) );
  INV_X1 U10573 ( .A(n10615), .ZN(n10614) );
  NAND2_X1 U10574 ( .A1(n10460), .A2(n10616), .ZN(n10615) );
  NAND2_X1 U10575 ( .A1(n10459), .A2(n10458), .ZN(n10616) );
  NOR2_X1 U10576 ( .A1(n8571), .A2(n8583), .ZN(n10460) );
  NOR2_X1 U10577 ( .A1(n10458), .A2(n10459), .ZN(n10613) );
  NOR2_X1 U10578 ( .A1(n10617), .A2(n10618), .ZN(n10459) );
  INV_X1 U10579 ( .A(n10619), .ZN(n10618) );
  NAND2_X1 U10580 ( .A1(n10455), .A2(n10620), .ZN(n10619) );
  NAND2_X1 U10581 ( .A1(n10456), .A2(n10454), .ZN(n10620) );
  NOR2_X1 U10582 ( .A1(n8571), .A2(n8580), .ZN(n10455) );
  NOR2_X1 U10583 ( .A1(n10454), .A2(n10456), .ZN(n10617) );
  NOR2_X1 U10584 ( .A1(n10621), .A2(n10622), .ZN(n10456) );
  INV_X1 U10585 ( .A(n10623), .ZN(n10622) );
  NAND2_X1 U10586 ( .A1(n10452), .A2(n10624), .ZN(n10623) );
  NAND2_X1 U10587 ( .A1(n10451), .A2(n10450), .ZN(n10624) );
  NOR2_X1 U10588 ( .A1(n10158), .A2(n8588), .ZN(n10452) );
  NOR2_X1 U10589 ( .A1(n10450), .A2(n10451), .ZN(n10621) );
  NOR2_X1 U10590 ( .A1(n10625), .A2(n10626), .ZN(n10451) );
  INV_X1 U10591 ( .A(n10627), .ZN(n10626) );
  NAND2_X1 U10592 ( .A1(n10448), .A2(n10628), .ZN(n10627) );
  NAND2_X1 U10593 ( .A1(n10447), .A2(n10445), .ZN(n10628) );
  NOR2_X1 U10594 ( .A1(n10158), .A2(n8551), .ZN(n10448) );
  NOR2_X1 U10595 ( .A1(n10445), .A2(n10447), .ZN(n10625) );
  NOR2_X1 U10596 ( .A1(n10629), .A2(n10630), .ZN(n10447) );
  INV_X1 U10597 ( .A(n10631), .ZN(n10630) );
  NAND2_X1 U10598 ( .A1(n10444), .A2(n10632), .ZN(n10631) );
  NAND2_X1 U10599 ( .A1(n10443), .A2(n10442), .ZN(n10632) );
  NOR2_X1 U10600 ( .A1(n10158), .A2(n8563), .ZN(n10444) );
  NOR2_X1 U10601 ( .A1(n10442), .A2(n10443), .ZN(n10629) );
  NOR2_X1 U10602 ( .A1(n10633), .A2(n10634), .ZN(n10443) );
  INV_X1 U10603 ( .A(n10635), .ZN(n10634) );
  NAND2_X1 U10604 ( .A1(n10440), .A2(n10636), .ZN(n10635) );
  NAND2_X1 U10605 ( .A1(n10439), .A2(n10437), .ZN(n10636) );
  NOR2_X1 U10606 ( .A1(n10158), .A2(n8548), .ZN(n10440) );
  NOR2_X1 U10607 ( .A1(n10437), .A2(n10439), .ZN(n10633) );
  NOR2_X1 U10608 ( .A1(n10637), .A2(n10638), .ZN(n10439) );
  INV_X1 U10609 ( .A(n10639), .ZN(n10638) );
  NAND2_X1 U10610 ( .A1(n10436), .A2(n10640), .ZN(n10639) );
  NAND2_X1 U10611 ( .A1(n10435), .A2(n10434), .ZN(n10640) );
  NOR2_X1 U10612 ( .A1(n10158), .A2(n8584), .ZN(n10436) );
  NOR2_X1 U10613 ( .A1(n10434), .A2(n10435), .ZN(n10637) );
  NOR2_X1 U10614 ( .A1(n10641), .A2(n10642), .ZN(n10435) );
  INV_X1 U10615 ( .A(n10643), .ZN(n10642) );
  NAND2_X1 U10616 ( .A1(n10431), .A2(n10644), .ZN(n10643) );
  NAND2_X1 U10617 ( .A1(n10432), .A2(n10430), .ZN(n10644) );
  NOR2_X1 U10618 ( .A1(n10158), .A2(n8535), .ZN(n10431) );
  NOR2_X1 U10619 ( .A1(n10430), .A2(n10432), .ZN(n10641) );
  NOR2_X1 U10620 ( .A1(n10645), .A2(n10646), .ZN(n10432) );
  INV_X1 U10621 ( .A(n10647), .ZN(n10646) );
  NAND2_X1 U10622 ( .A1(n10428), .A2(n10648), .ZN(n10647) );
  NAND2_X1 U10623 ( .A1(n10427), .A2(n10426), .ZN(n10648) );
  NOR2_X1 U10624 ( .A1(n10158), .A2(n8568), .ZN(n10428) );
  NOR2_X1 U10625 ( .A1(n10426), .A2(n10427), .ZN(n10645) );
  NOR2_X1 U10626 ( .A1(n10649), .A2(n10650), .ZN(n10427) );
  INV_X1 U10627 ( .A(n10651), .ZN(n10650) );
  NAND2_X1 U10628 ( .A1(n10423), .A2(n10652), .ZN(n10651) );
  NAND2_X1 U10629 ( .A1(n10424), .A2(n10422), .ZN(n10652) );
  NOR2_X1 U10630 ( .A1(n10158), .A2(n8574), .ZN(n10423) );
  NOR2_X1 U10631 ( .A1(n10422), .A2(n10424), .ZN(n10649) );
  NOR2_X1 U10632 ( .A1(n10653), .A2(n10654), .ZN(n10424) );
  INV_X1 U10633 ( .A(n10655), .ZN(n10654) );
  NAND2_X1 U10634 ( .A1(n10419), .A2(n10656), .ZN(n10655) );
  NAND2_X1 U10635 ( .A1(n10420), .A2(n10418), .ZN(n10656) );
  NOR2_X1 U10636 ( .A1(n10158), .A2(n8565), .ZN(n10419) );
  NOR2_X1 U10637 ( .A1(n10418), .A2(n10420), .ZN(n10653) );
  NOR2_X1 U10638 ( .A1(n10657), .A2(n10658), .ZN(n10420) );
  INV_X1 U10639 ( .A(n10659), .ZN(n10658) );
  NAND2_X1 U10640 ( .A1(n10413), .A2(n10660), .ZN(n10659) );
  NAND2_X1 U10641 ( .A1(n10416), .A2(n10415), .ZN(n10660) );
  NOR2_X1 U10642 ( .A1(n10158), .A2(n8567), .ZN(n10413) );
  NOR2_X1 U10643 ( .A1(n10415), .A2(n10416), .ZN(n10657) );
  INV_X1 U10644 ( .A(n10661), .ZN(n10416) );
  NAND2_X1 U10645 ( .A1(n10662), .A2(n10663), .ZN(n10661) );
  NAND2_X1 U10646 ( .A1(n8540), .A2(n10664), .ZN(n10663) );
  NAND2_X1 U10647 ( .A1(n8624), .A2(n10665), .ZN(n10664) );
  NAND2_X1 U10648 ( .A1(n8576), .A2(n8585), .ZN(n10665) );
  NAND2_X1 U10649 ( .A1(n10667), .A2(n10668), .ZN(n10662) );
  NAND2_X1 U10650 ( .A1(n8630), .A2(n10669), .ZN(n10668) );
  NAND2_X1 U10651 ( .A1(n8539), .A2(n8541), .ZN(n10669) );
  NAND3_X1 U10652 ( .A1(n8540), .A2(n8537), .A3(n10159), .ZN(n10415) );
  XOR2_X1 U10653 ( .A(n10670), .B(n10671), .Z(n10418) );
  XNOR2_X1 U10654 ( .A(n10672), .B(n10673), .ZN(n10671) );
  XOR2_X1 U10655 ( .A(n10674), .B(n10675), .Z(n10422) );
  XNOR2_X1 U10656 ( .A(n10676), .B(n10677), .ZN(n10674) );
  XOR2_X1 U10657 ( .A(n10678), .B(n10679), .Z(n10426) );
  XNOR2_X1 U10658 ( .A(n10680), .B(n10681), .ZN(n10678) );
  XOR2_X1 U10659 ( .A(n10682), .B(n10683), .Z(n10430) );
  XNOR2_X1 U10660 ( .A(n10684), .B(n10685), .ZN(n10682) );
  XOR2_X1 U10661 ( .A(n10686), .B(n10687), .Z(n10434) );
  XNOR2_X1 U10662 ( .A(n10688), .B(n10689), .ZN(n10686) );
  NOR2_X1 U10663 ( .A1(n8535), .A2(n8541), .ZN(n10689) );
  XOR2_X1 U10664 ( .A(n10690), .B(n10691), .Z(n10437) );
  XNOR2_X1 U10665 ( .A(n10692), .B(n10693), .ZN(n10690) );
  NOR2_X1 U10666 ( .A1(n8584), .A2(n8541), .ZN(n10693) );
  XOR2_X1 U10667 ( .A(n10694), .B(n10695), .Z(n10442) );
  XNOR2_X1 U10668 ( .A(n10696), .B(n10697), .ZN(n10694) );
  NOR2_X1 U10669 ( .A1(n8548), .A2(n8541), .ZN(n10697) );
  XOR2_X1 U10670 ( .A(n10698), .B(n10699), .Z(n10445) );
  XNOR2_X1 U10671 ( .A(n10700), .B(n10701), .ZN(n10698) );
  NOR2_X1 U10672 ( .A1(n8563), .A2(n8541), .ZN(n10701) );
  XOR2_X1 U10673 ( .A(n10702), .B(n10703), .Z(n10450) );
  XNOR2_X1 U10674 ( .A(n10704), .B(n10705), .ZN(n10702) );
  NOR2_X1 U10675 ( .A1(n8551), .A2(n8541), .ZN(n10705) );
  XOR2_X1 U10676 ( .A(n10706), .B(n10707), .Z(n10454) );
  XNOR2_X1 U10677 ( .A(n10708), .B(n10709), .ZN(n10706) );
  NOR2_X1 U10678 ( .A1(n8588), .A2(n8541), .ZN(n10709) );
  XOR2_X1 U10679 ( .A(n10710), .B(n10711), .Z(n10458) );
  XNOR2_X1 U10680 ( .A(n10712), .B(n10713), .ZN(n10710) );
  NOR2_X1 U10681 ( .A1(n8580), .A2(n8541), .ZN(n10713) );
  XOR2_X1 U10682 ( .A(n10714), .B(n10715), .Z(n10462) );
  XNOR2_X1 U10683 ( .A(n10716), .B(n10717), .ZN(n10714) );
  NOR2_X1 U10684 ( .A1(n8583), .A2(n8541), .ZN(n10717) );
  XNOR2_X1 U10685 ( .A(n10718), .B(n10719), .ZN(n10466) );
  XNOR2_X1 U10686 ( .A(n10720), .B(n10721), .ZN(n10719) );
  NAND2_X1 U10687 ( .A1(n8540), .A2(n10722), .ZN(n10721) );
  XOR2_X1 U10688 ( .A(n10723), .B(n10724), .Z(n10470) );
  XNOR2_X1 U10689 ( .A(n10725), .B(n10726), .ZN(n10723) );
  NOR2_X1 U10690 ( .A1(n9050), .A2(n8541), .ZN(n10726) );
  XOR2_X1 U10691 ( .A(n10727), .B(n10728), .Z(n10473) );
  XNOR2_X1 U10692 ( .A(n10729), .B(n10730), .ZN(n10727) );
  NOR2_X1 U10693 ( .A1(n8545), .A2(n8541), .ZN(n10730) );
  XNOR2_X1 U10694 ( .A(n10731), .B(n10732), .ZN(n10478) );
  XNOR2_X1 U10695 ( .A(n10733), .B(n10734), .ZN(n10731) );
  NOR2_X1 U10696 ( .A1(n9041), .A2(n8541), .ZN(n10734) );
  XNOR2_X1 U10697 ( .A(n10735), .B(n10736), .ZN(n10482) );
  XNOR2_X1 U10698 ( .A(n10737), .B(n10738), .ZN(n10735) );
  NOR2_X1 U10699 ( .A1(n8591), .A2(n8541), .ZN(n10738) );
  XNOR2_X1 U10700 ( .A(n10739), .B(n10740), .ZN(n10486) );
  XNOR2_X1 U10701 ( .A(n10741), .B(n10742), .ZN(n10739) );
  NOR2_X1 U10702 ( .A1(n8582), .A2(n8541), .ZN(n10742) );
  INV_X1 U10703 ( .A(n10743), .ZN(n10582) );
  NOR2_X1 U10704 ( .A1(n10492), .A2(n10489), .ZN(n10743) );
  XNOR2_X1 U10705 ( .A(n10744), .B(n10745), .ZN(n10489) );
  XOR2_X1 U10706 ( .A(n10746), .B(n10747), .Z(n10744) );
  NOR2_X1 U10707 ( .A1(n8572), .A2(n8541), .ZN(n10747) );
  NAND2_X1 U10708 ( .A1(n10159), .A2(n9304), .ZN(n10492) );
  XNOR2_X1 U10709 ( .A(n10748), .B(n10749), .ZN(n10494) );
  XNOR2_X1 U10710 ( .A(n10750), .B(n10751), .ZN(n10748) );
  XOR2_X1 U10711 ( .A(n10752), .B(n10753), .Z(n10498) );
  XOR2_X1 U10712 ( .A(n10754), .B(n10755), .Z(n10753) );
  NOR2_X1 U10713 ( .A1(n8594), .A2(n8541), .ZN(n10755) );
  XNOR2_X1 U10714 ( .A(n10756), .B(n10757), .ZN(n10502) );
  XNOR2_X1 U10715 ( .A(n10758), .B(n10759), .ZN(n10756) );
  NOR2_X1 U10716 ( .A1(n8560), .A2(n8541), .ZN(n10759) );
  NOR2_X1 U10717 ( .A1(n10510), .A2(n10507), .ZN(n10566) );
  XOR2_X1 U10718 ( .A(n10760), .B(n10761), .Z(n10507) );
  XNOR2_X1 U10719 ( .A(n10762), .B(n10763), .ZN(n10760) );
  NOR2_X1 U10720 ( .A1(n8544), .A2(n8541), .ZN(n10763) );
  NAND2_X1 U10721 ( .A1(n10159), .A2(n9286), .ZN(n10510) );
  INV_X1 U10722 ( .A(n10158), .ZN(n10159) );
  XNOR2_X1 U10723 ( .A(n10764), .B(n10765), .ZN(n10158) );
  XOR2_X1 U10724 ( .A(d_25_), .B(c_25_), .Z(n10765) );
  XNOR2_X1 U10725 ( .A(n10766), .B(n10767), .ZN(n10512) );
  XOR2_X1 U10726 ( .A(n10768), .B(n10769), .Z(n10767) );
  XOR2_X1 U10727 ( .A(n10770), .B(n10771), .Z(n10520) );
  XNOR2_X1 U10728 ( .A(n10772), .B(n10773), .ZN(n10771) );
  NAND2_X1 U10729 ( .A1(n8540), .A2(n9277), .ZN(n10773) );
  XOR2_X1 U10730 ( .A(n10774), .B(n10775), .Z(n10523) );
  XOR2_X1 U10731 ( .A(n10776), .B(n10777), .Z(n10774) );
  XNOR2_X1 U10732 ( .A(n10778), .B(n10779), .ZN(n10528) );
  XOR2_X1 U10733 ( .A(n10780), .B(n10781), .Z(n10779) );
  NAND2_X1 U10734 ( .A1(n8540), .A2(n9268), .ZN(n10781) );
  XOR2_X1 U10735 ( .A(n10782), .B(n10783), .Z(n10534) );
  XNOR2_X1 U10736 ( .A(n10784), .B(n10785), .ZN(n10783) );
  XOR2_X1 U10737 ( .A(n10786), .B(n10787), .Z(n10532) );
  XNOR2_X1 U10738 ( .A(n10788), .B(n10789), .ZN(n10786) );
  NAND2_X1 U10739 ( .A1(n8944), .A2(n8945), .ZN(n10537) );
  INV_X1 U10740 ( .A(n10790), .ZN(n8810) );
  NOR2_X1 U10741 ( .A1(n8940), .A2(n8939), .ZN(n10790) );
  NAND2_X1 U10742 ( .A1(n8935), .A2(n10791), .ZN(n8939) );
  NAND2_X1 U10743 ( .A1(n10792), .A2(n10793), .ZN(n10791) );
  INV_X1 U10744 ( .A(n8932), .ZN(n8935) );
  NOR2_X1 U10745 ( .A1(n10793), .A2(n10792), .ZN(n8932) );
  NOR2_X1 U10746 ( .A1(n10794), .A2(n10795), .ZN(n10792) );
  INV_X1 U10747 ( .A(n10796), .ZN(n10795) );
  NAND3_X1 U10748 ( .A1(n8592), .A2(n10797), .A3(n10667), .ZN(n10796) );
  NAND2_X1 U10749 ( .A1(n10798), .A2(n10799), .ZN(n10797) );
  NOR2_X1 U10750 ( .A1(n10799), .A2(n10798), .ZN(n10794) );
  XNOR2_X1 U10751 ( .A(n10800), .B(n10801), .ZN(n10793) );
  XOR2_X1 U10752 ( .A(n10802), .B(n10803), .Z(n10800) );
  NOR2_X1 U10753 ( .A1(n8972), .A2(n8547), .ZN(n10803) );
  INV_X1 U10754 ( .A(n10805), .ZN(n8940) );
  NOR2_X1 U10755 ( .A1(n8945), .A2(n8944), .ZN(n10805) );
  NOR2_X1 U10756 ( .A1(n10806), .A2(n10807), .ZN(n8944) );
  INV_X1 U10757 ( .A(n10808), .ZN(n10807) );
  NAND2_X1 U10758 ( .A1(n10789), .A2(n10809), .ZN(n10808) );
  NAND2_X1 U10759 ( .A1(n10788), .A2(n10787), .ZN(n10809) );
  NOR2_X1 U10760 ( .A1(n8541), .A2(n8972), .ZN(n10789) );
  NOR2_X1 U10761 ( .A1(n10787), .A2(n10788), .ZN(n10806) );
  INV_X1 U10762 ( .A(n10810), .ZN(n10788) );
  NAND2_X1 U10763 ( .A1(n10811), .A2(n10812), .ZN(n10810) );
  NAND2_X1 U10764 ( .A1(n10784), .A2(n10813), .ZN(n10812) );
  NAND2_X1 U10765 ( .A1(n10782), .A2(n10814), .ZN(n10813) );
  INV_X1 U10766 ( .A(n10785), .ZN(n10814) );
  NAND2_X1 U10767 ( .A1(n10815), .A2(n10816), .ZN(n10784) );
  INV_X1 U10768 ( .A(n10817), .ZN(n10816) );
  NOR3_X1 U10769 ( .A1(n8982), .A2(n10818), .A3(n8541), .ZN(n10817) );
  NOR2_X1 U10770 ( .A1(n10780), .A2(n10778), .ZN(n10818) );
  NAND2_X1 U10771 ( .A1(n10778), .A2(n10780), .ZN(n10815) );
  NAND2_X1 U10772 ( .A1(n10819), .A2(n10820), .ZN(n10780) );
  NAND2_X1 U10773 ( .A1(n10776), .A2(n10821), .ZN(n10820) );
  INV_X1 U10774 ( .A(n10822), .ZN(n10821) );
  NOR2_X1 U10775 ( .A1(n10775), .A2(n10777), .ZN(n10822) );
  NAND2_X1 U10776 ( .A1(n10823), .A2(n10824), .ZN(n10776) );
  NAND3_X1 U10777 ( .A1(n9277), .A2(n10825), .A3(n8540), .ZN(n10824) );
  NAND2_X1 U10778 ( .A1(n10772), .A2(n10770), .ZN(n10825) );
  INV_X1 U10779 ( .A(n10826), .ZN(n10823) );
  NOR2_X1 U10780 ( .A1(n10770), .A2(n10772), .ZN(n10826) );
  NOR2_X1 U10781 ( .A1(n10827), .A2(n10828), .ZN(n10772) );
  NOR3_X1 U10782 ( .A1(n8995), .A2(n10829), .A3(n8541), .ZN(n10828) );
  INV_X1 U10783 ( .A(n10830), .ZN(n10829) );
  NAND2_X1 U10784 ( .A1(n10560), .A2(n10558), .ZN(n10830) );
  NOR2_X1 U10785 ( .A1(n10558), .A2(n10560), .ZN(n10827) );
  NOR2_X1 U10786 ( .A1(n10831), .A2(n10832), .ZN(n10560) );
  INV_X1 U10787 ( .A(n10833), .ZN(n10832) );
  NAND2_X1 U10788 ( .A1(n10768), .A2(n10834), .ZN(n10833) );
  NAND2_X1 U10789 ( .A1(n10769), .A2(n10766), .ZN(n10834) );
  NOR2_X1 U10790 ( .A1(n8541), .A2(n8555), .ZN(n10768) );
  NOR2_X1 U10791 ( .A1(n10766), .A2(n10769), .ZN(n10831) );
  NOR2_X1 U10792 ( .A1(n10835), .A2(n10836), .ZN(n10769) );
  NOR3_X1 U10793 ( .A1(n8544), .A2(n10837), .A3(n8541), .ZN(n10836) );
  INV_X1 U10794 ( .A(n10838), .ZN(n10837) );
  NAND2_X1 U10795 ( .A1(n10762), .A2(n10761), .ZN(n10838) );
  NOR2_X1 U10796 ( .A1(n10761), .A2(n10762), .ZN(n10835) );
  NOR2_X1 U10797 ( .A1(n10839), .A2(n10840), .ZN(n10762) );
  INV_X1 U10798 ( .A(n10841), .ZN(n10840) );
  NAND3_X1 U10799 ( .A1(n9295), .A2(n10842), .A3(n8540), .ZN(n10841) );
  NAND2_X1 U10800 ( .A1(n10758), .A2(n10757), .ZN(n10842) );
  NOR2_X1 U10801 ( .A1(n10757), .A2(n10758), .ZN(n10839) );
  NOR2_X1 U10802 ( .A1(n10843), .A2(n10844), .ZN(n10758) );
  INV_X1 U10803 ( .A(n10845), .ZN(n10844) );
  NAND3_X1 U10804 ( .A1(n10846), .A2(n10847), .A3(n8540), .ZN(n10845) );
  NAND2_X1 U10805 ( .A1(n10754), .A2(n10752), .ZN(n10847) );
  NOR2_X1 U10806 ( .A1(n10752), .A2(n10754), .ZN(n10843) );
  NOR2_X1 U10807 ( .A1(n10848), .A2(n10849), .ZN(n10754) );
  INV_X1 U10808 ( .A(n10850), .ZN(n10849) );
  NAND2_X1 U10809 ( .A1(n10750), .A2(n10851), .ZN(n10850) );
  NAND2_X1 U10810 ( .A1(n10749), .A2(n10751), .ZN(n10851) );
  NAND2_X1 U10811 ( .A1(n10852), .A2(n10853), .ZN(n10750) );
  INV_X1 U10812 ( .A(n10854), .ZN(n10853) );
  NOR3_X1 U10813 ( .A1(n9025), .A2(n10855), .A3(n8541), .ZN(n10854) );
  NOR2_X1 U10814 ( .A1(n10746), .A2(n10745), .ZN(n10855) );
  NAND2_X1 U10815 ( .A1(n10745), .A2(n10746), .ZN(n10852) );
  NAND2_X1 U10816 ( .A1(n10856), .A2(n10857), .ZN(n10746) );
  NAND3_X1 U10817 ( .A1(n9313), .A2(n10858), .A3(n8540), .ZN(n10857) );
  NAND2_X1 U10818 ( .A1(n10741), .A2(n10740), .ZN(n10858) );
  INV_X1 U10819 ( .A(n10859), .ZN(n10856) );
  NOR2_X1 U10820 ( .A1(n10740), .A2(n10741), .ZN(n10859) );
  NOR2_X1 U10821 ( .A1(n10860), .A2(n10861), .ZN(n10741) );
  NOR3_X1 U10822 ( .A1(n9036), .A2(n10862), .A3(n8541), .ZN(n10861) );
  INV_X1 U10823 ( .A(n10863), .ZN(n10862) );
  NAND2_X1 U10824 ( .A1(n10737), .A2(n10736), .ZN(n10863) );
  NOR2_X1 U10825 ( .A1(n10736), .A2(n10737), .ZN(n10860) );
  NOR2_X1 U10826 ( .A1(n10864), .A2(n10865), .ZN(n10737) );
  INV_X1 U10827 ( .A(n10866), .ZN(n10865) );
  NAND3_X1 U10828 ( .A1(n9322), .A2(n10867), .A3(n8540), .ZN(n10866) );
  NAND2_X1 U10829 ( .A1(n10733), .A2(n10732), .ZN(n10867) );
  NOR2_X1 U10830 ( .A1(n10732), .A2(n10733), .ZN(n10864) );
  NOR2_X1 U10831 ( .A1(n10868), .A2(n10869), .ZN(n10733) );
  NOR3_X1 U10832 ( .A1(n8545), .A2(n10870), .A3(n8541), .ZN(n10869) );
  INV_X1 U10833 ( .A(n10871), .ZN(n10870) );
  NAND2_X1 U10834 ( .A1(n10729), .A2(n10728), .ZN(n10871) );
  NOR2_X1 U10835 ( .A1(n10728), .A2(n10729), .ZN(n10868) );
  NOR2_X1 U10836 ( .A1(n10872), .A2(n10873), .ZN(n10729) );
  INV_X1 U10837 ( .A(n10874), .ZN(n10873) );
  NAND3_X1 U10838 ( .A1(n9331), .A2(n10875), .A3(n8540), .ZN(n10874) );
  NAND2_X1 U10839 ( .A1(n10725), .A2(n10724), .ZN(n10875) );
  NOR2_X1 U10840 ( .A1(n10724), .A2(n10725), .ZN(n10872) );
  NOR2_X1 U10841 ( .A1(n10876), .A2(n10877), .ZN(n10725) );
  NOR3_X1 U10842 ( .A1(n9056), .A2(n10878), .A3(n8541), .ZN(n10877) );
  INV_X1 U10843 ( .A(n10879), .ZN(n10878) );
  NAND2_X1 U10844 ( .A1(n10720), .A2(n10718), .ZN(n10879) );
  NOR2_X1 U10845 ( .A1(n10718), .A2(n10720), .ZN(n10876) );
  NOR2_X1 U10846 ( .A1(n10880), .A2(n10881), .ZN(n10720) );
  INV_X1 U10847 ( .A(n10882), .ZN(n10881) );
  NAND3_X1 U10848 ( .A1(n9340), .A2(n10883), .A3(n8540), .ZN(n10882) );
  NAND2_X1 U10849 ( .A1(n10716), .A2(n10715), .ZN(n10883) );
  NOR2_X1 U10850 ( .A1(n10715), .A2(n10716), .ZN(n10880) );
  NOR2_X1 U10851 ( .A1(n10884), .A2(n10885), .ZN(n10716) );
  NOR3_X1 U10852 ( .A1(n9066), .A2(n10886), .A3(n8541), .ZN(n10885) );
  INV_X1 U10853 ( .A(n10887), .ZN(n10886) );
  NAND2_X1 U10854 ( .A1(n10712), .A2(n10711), .ZN(n10887) );
  NOR2_X1 U10855 ( .A1(n10711), .A2(n10712), .ZN(n10884) );
  NOR2_X1 U10856 ( .A1(n10888), .A2(n10889), .ZN(n10712) );
  INV_X1 U10857 ( .A(n10890), .ZN(n10889) );
  NAND3_X1 U10858 ( .A1(n9080), .A2(n10891), .A3(n8540), .ZN(n10890) );
  NAND2_X1 U10859 ( .A1(n10708), .A2(n10707), .ZN(n10891) );
  NOR2_X1 U10860 ( .A1(n10707), .A2(n10708), .ZN(n10888) );
  NOR2_X1 U10861 ( .A1(n10892), .A2(n10893), .ZN(n10708) );
  NOR3_X1 U10862 ( .A1(n8551), .A2(n10894), .A3(n8541), .ZN(n10893) );
  INV_X1 U10863 ( .A(n10895), .ZN(n10894) );
  NAND2_X1 U10864 ( .A1(n10704), .A2(n10703), .ZN(n10895) );
  NOR2_X1 U10865 ( .A1(n10703), .A2(n10704), .ZN(n10892) );
  NOR2_X1 U10866 ( .A1(n10896), .A2(n10897), .ZN(n10704) );
  INV_X1 U10867 ( .A(n10898), .ZN(n10897) );
  NAND3_X1 U10868 ( .A1(n9098), .A2(n10899), .A3(n8540), .ZN(n10898) );
  NAND2_X1 U10869 ( .A1(n10700), .A2(n10699), .ZN(n10899) );
  NOR2_X1 U10870 ( .A1(n10699), .A2(n10700), .ZN(n10896) );
  NOR2_X1 U10871 ( .A1(n10900), .A2(n10901), .ZN(n10700) );
  NOR3_X1 U10872 ( .A1(n8548), .A2(n10902), .A3(n8541), .ZN(n10901) );
  INV_X1 U10873 ( .A(n10903), .ZN(n10902) );
  NAND2_X1 U10874 ( .A1(n10696), .A2(n10695), .ZN(n10903) );
  NOR2_X1 U10875 ( .A1(n10695), .A2(n10696), .ZN(n10900) );
  NOR2_X1 U10876 ( .A1(n10904), .A2(n10905), .ZN(n10696) );
  INV_X1 U10877 ( .A(n10906), .ZN(n10905) );
  NAND3_X1 U10878 ( .A1(n9112), .A2(n10907), .A3(n8540), .ZN(n10906) );
  NAND2_X1 U10879 ( .A1(n10692), .A2(n10691), .ZN(n10907) );
  NOR2_X1 U10880 ( .A1(n10691), .A2(n10692), .ZN(n10904) );
  NOR2_X1 U10881 ( .A1(n10908), .A2(n10909), .ZN(n10692) );
  INV_X1 U10882 ( .A(n10910), .ZN(n10909) );
  NAND3_X1 U10883 ( .A1(n9121), .A2(n10911), .A3(n8540), .ZN(n10910) );
  NAND2_X1 U10884 ( .A1(n10688), .A2(n10687), .ZN(n10911) );
  NOR2_X1 U10885 ( .A1(n10687), .A2(n10688), .ZN(n10908) );
  NOR2_X1 U10886 ( .A1(n10912), .A2(n10913), .ZN(n10688) );
  INV_X1 U10887 ( .A(n10914), .ZN(n10913) );
  NAND2_X1 U10888 ( .A1(n10684), .A2(n10915), .ZN(n10914) );
  NAND2_X1 U10889 ( .A1(n10685), .A2(n10683), .ZN(n10915) );
  NOR2_X1 U10890 ( .A1(n8541), .A2(n8568), .ZN(n10684) );
  NOR2_X1 U10891 ( .A1(n10683), .A2(n10685), .ZN(n10912) );
  NOR2_X1 U10892 ( .A1(n10916), .A2(n10917), .ZN(n10685) );
  INV_X1 U10893 ( .A(n10918), .ZN(n10917) );
  NAND2_X1 U10894 ( .A1(n10680), .A2(n10919), .ZN(n10918) );
  NAND2_X1 U10895 ( .A1(n10681), .A2(n10679), .ZN(n10919) );
  NOR2_X1 U10896 ( .A1(n8541), .A2(n8574), .ZN(n10680) );
  NOR2_X1 U10897 ( .A1(n10679), .A2(n10681), .ZN(n10916) );
  NOR2_X1 U10898 ( .A1(n10920), .A2(n10921), .ZN(n10681) );
  INV_X1 U10899 ( .A(n10922), .ZN(n10921) );
  NAND2_X1 U10900 ( .A1(n10676), .A2(n10923), .ZN(n10922) );
  NAND2_X1 U10901 ( .A1(n10677), .A2(n10675), .ZN(n10923) );
  NOR2_X1 U10902 ( .A1(n8541), .A2(n8565), .ZN(n10676) );
  NOR2_X1 U10903 ( .A1(n10675), .A2(n10677), .ZN(n10920) );
  NOR2_X1 U10904 ( .A1(n10924), .A2(n10925), .ZN(n10677) );
  INV_X1 U10905 ( .A(n10926), .ZN(n10925) );
  NAND2_X1 U10906 ( .A1(n10670), .A2(n10927), .ZN(n10926) );
  NAND2_X1 U10907 ( .A1(n10673), .A2(n10672), .ZN(n10927) );
  NOR2_X1 U10908 ( .A1(n8541), .A2(n8567), .ZN(n10670) );
  NOR2_X1 U10909 ( .A1(n10672), .A2(n10673), .ZN(n10924) );
  INV_X1 U10910 ( .A(n10928), .ZN(n10673) );
  NAND2_X1 U10911 ( .A1(n10929), .A2(n10930), .ZN(n10928) );
  NAND2_X1 U10912 ( .A1(n10667), .A2(n10931), .ZN(n10930) );
  NAND2_X1 U10913 ( .A1(n8624), .A2(n10932), .ZN(n10931) );
  NAND2_X1 U10914 ( .A1(n8547), .A2(n8585), .ZN(n10932) );
  NAND2_X1 U10915 ( .A1(n8546), .A2(n10933), .ZN(n10929) );
  NAND2_X1 U10916 ( .A1(n8630), .A2(n10934), .ZN(n10933) );
  NAND2_X1 U10917 ( .A1(n8539), .A2(n8576), .ZN(n10934) );
  NAND3_X1 U10918 ( .A1(n10667), .A2(n8537), .A3(n8540), .ZN(n10672) );
  XOR2_X1 U10919 ( .A(n10935), .B(n10936), .Z(n10675) );
  XNOR2_X1 U10920 ( .A(n10937), .B(n10938), .ZN(n10936) );
  XOR2_X1 U10921 ( .A(n10939), .B(n10940), .Z(n10679) );
  XNOR2_X1 U10922 ( .A(n10941), .B(n10942), .ZN(n10939) );
  XOR2_X1 U10923 ( .A(n10943), .B(n10944), .Z(n10683) );
  XNOR2_X1 U10924 ( .A(n10945), .B(n10946), .ZN(n10943) );
  XOR2_X1 U10925 ( .A(n10947), .B(n10948), .Z(n10687) );
  XNOR2_X1 U10926 ( .A(n10949), .B(n10950), .ZN(n10947) );
  XOR2_X1 U10927 ( .A(n10951), .B(n10952), .Z(n10691) );
  XNOR2_X1 U10928 ( .A(n10953), .B(n10954), .ZN(n10951) );
  XOR2_X1 U10929 ( .A(n10955), .B(n10956), .Z(n10695) );
  XNOR2_X1 U10930 ( .A(n10957), .B(n10958), .ZN(n10955) );
  XNOR2_X1 U10931 ( .A(n10959), .B(n10960), .ZN(n10699) );
  XOR2_X1 U10932 ( .A(n10961), .B(n10962), .Z(n10960) );
  XOR2_X1 U10933 ( .A(n10963), .B(n10964), .Z(n10703) );
  XNOR2_X1 U10934 ( .A(n10965), .B(n10966), .ZN(n10963) );
  XOR2_X1 U10935 ( .A(n10967), .B(n10968), .Z(n10707) );
  XNOR2_X1 U10936 ( .A(n10969), .B(n10970), .ZN(n10967) );
  XOR2_X1 U10937 ( .A(n10971), .B(n10972), .Z(n10711) );
  XNOR2_X1 U10938 ( .A(n10973), .B(n10974), .ZN(n10971) );
  XOR2_X1 U10939 ( .A(n10975), .B(n10976), .Z(n10715) );
  XNOR2_X1 U10940 ( .A(n10977), .B(n10978), .ZN(n10975) );
  XOR2_X1 U10941 ( .A(n10979), .B(n10980), .Z(n10718) );
  XNOR2_X1 U10942 ( .A(n10981), .B(n10982), .ZN(n10979) );
  XOR2_X1 U10943 ( .A(n10983), .B(n10984), .Z(n10724) );
  XNOR2_X1 U10944 ( .A(n10985), .B(n10986), .ZN(n10983) );
  XNOR2_X1 U10945 ( .A(n10987), .B(n10988), .ZN(n10728) );
  XOR2_X1 U10946 ( .A(n10989), .B(n10990), .Z(n10988) );
  XNOR2_X1 U10947 ( .A(n10991), .B(n10992), .ZN(n10732) );
  XOR2_X1 U10948 ( .A(n10993), .B(n10994), .Z(n10991) );
  NOR2_X1 U10949 ( .A1(n8545), .A2(n8576), .ZN(n10994) );
  XOR2_X1 U10950 ( .A(n10995), .B(n10996), .Z(n10736) );
  XNOR2_X1 U10951 ( .A(n10997), .B(n10998), .ZN(n10995) );
  XOR2_X1 U10952 ( .A(n10999), .B(n11000), .Z(n10740) );
  XNOR2_X1 U10953 ( .A(n11001), .B(n11002), .ZN(n10999) );
  NOR2_X1 U10954 ( .A1(n8591), .A2(n8576), .ZN(n11002) );
  XOR2_X1 U10955 ( .A(n11003), .B(n11004), .Z(n10745) );
  XOR2_X1 U10956 ( .A(n11005), .B(n11006), .Z(n11004) );
  NOR2_X1 U10957 ( .A1(n10751), .A2(n10749), .ZN(n10848) );
  XNOR2_X1 U10958 ( .A(n11007), .B(n11008), .ZN(n10749) );
  XOR2_X1 U10959 ( .A(n11009), .B(n11010), .Z(n11007) );
  NOR2_X1 U10960 ( .A1(n8572), .A2(n8576), .ZN(n11010) );
  NAND2_X1 U10961 ( .A1(n8540), .A2(n9304), .ZN(n10751) );
  XOR2_X1 U10962 ( .A(n11011), .B(n11012), .Z(n10752) );
  XOR2_X1 U10963 ( .A(n11013), .B(n11014), .Z(n11012) );
  NAND2_X1 U10964 ( .A1(n10667), .A2(n9304), .ZN(n11014) );
  XNOR2_X1 U10965 ( .A(n11015), .B(n11016), .ZN(n10757) );
  XOR2_X1 U10966 ( .A(n11017), .B(n11018), .Z(n11015) );
  NOR2_X1 U10967 ( .A1(n8594), .A2(n8576), .ZN(n11018) );
  XOR2_X1 U10968 ( .A(n11019), .B(n11020), .Z(n10761) );
  XNOR2_X1 U10969 ( .A(n11021), .B(n11022), .ZN(n11019) );
  XOR2_X1 U10970 ( .A(n11023), .B(n11024), .Z(n10766) );
  XNOR2_X1 U10971 ( .A(n11025), .B(n11026), .ZN(n11023) );
  NOR2_X1 U10972 ( .A1(n8544), .A2(n8576), .ZN(n11026) );
  XOR2_X1 U10973 ( .A(n11027), .B(n11028), .Z(n10558) );
  NAND2_X1 U10974 ( .A1(n11029), .A2(n11030), .ZN(n11027) );
  XOR2_X1 U10975 ( .A(n11031), .B(n11032), .Z(n10770) );
  XOR2_X1 U10976 ( .A(n11033), .B(n11034), .Z(n11032) );
  NAND2_X1 U10977 ( .A1(n10667), .A2(n10307), .ZN(n11034) );
  NAND2_X1 U10978 ( .A1(n10777), .A2(n10775), .ZN(n10819) );
  XNOR2_X1 U10979 ( .A(n11035), .B(n11036), .ZN(n10775) );
  XOR2_X1 U10980 ( .A(n11037), .B(n11038), .Z(n11036) );
  NAND2_X1 U10981 ( .A1(n10667), .A2(n9277), .ZN(n11038) );
  NOR2_X1 U10982 ( .A1(n8541), .A2(n8527), .ZN(n10777) );
  XOR2_X1 U10983 ( .A(n11039), .B(n11040), .Z(n10778) );
  XOR2_X1 U10984 ( .A(n11041), .B(n11042), .Z(n11039) );
  NOR2_X1 U10985 ( .A1(n8527), .A2(n8576), .ZN(n11042) );
  NAND2_X1 U10986 ( .A1(n10785), .A2(n11043), .ZN(n10811) );
  INV_X1 U10987 ( .A(n10782), .ZN(n11043) );
  XOR2_X1 U10988 ( .A(n11044), .B(n11045), .Z(n10782) );
  XOR2_X1 U10989 ( .A(n11046), .B(n11047), .Z(n11045) );
  NAND2_X1 U10990 ( .A1(n10667), .A2(n9268), .ZN(n11047) );
  NOR2_X1 U10991 ( .A1(n8541), .A2(n8589), .ZN(n10785) );
  XNOR2_X1 U10992 ( .A(n11048), .B(n11049), .ZN(n10410) );
  XOR2_X1 U10993 ( .A(d_24_), .B(c_24_), .Z(n11049) );
  XNOR2_X1 U10994 ( .A(n11050), .B(n11051), .ZN(n10787) );
  XOR2_X1 U10995 ( .A(n11052), .B(n11053), .Z(n11050) );
  NOR2_X1 U10996 ( .A1(n8589), .A2(n8576), .ZN(n11053) );
  XNOR2_X1 U10997 ( .A(n10799), .B(n11054), .ZN(n8945) );
  XNOR2_X1 U10998 ( .A(n10798), .B(n11055), .ZN(n11054) );
  NAND2_X1 U10999 ( .A1(n10667), .A2(n8592), .ZN(n11055) );
  NOR2_X1 U11000 ( .A1(n11056), .A2(n11057), .ZN(n10798) );
  NOR3_X1 U11001 ( .A1(n8884), .A2(n11058), .A3(n8576), .ZN(n11057) );
  NOR2_X1 U11002 ( .A1(n11052), .A2(n11051), .ZN(n11058) );
  INV_X1 U11003 ( .A(n11059), .ZN(n11056) );
  NAND2_X1 U11004 ( .A1(n11051), .A2(n11052), .ZN(n11059) );
  NAND2_X1 U11005 ( .A1(n11060), .A2(n11061), .ZN(n11052) );
  INV_X1 U11006 ( .A(n11062), .ZN(n11061) );
  NOR3_X1 U11007 ( .A1(n8982), .A2(n11063), .A3(n8576), .ZN(n11062) );
  NOR2_X1 U11008 ( .A1(n11046), .A2(n11044), .ZN(n11063) );
  NAND2_X1 U11009 ( .A1(n11044), .A2(n11046), .ZN(n11060) );
  NAND2_X1 U11010 ( .A1(n11064), .A2(n11065), .ZN(n11046) );
  NAND3_X1 U11011 ( .A1(n9792), .A2(n11066), .A3(n10667), .ZN(n11065) );
  INV_X1 U11012 ( .A(n11067), .ZN(n11066) );
  NOR2_X1 U11013 ( .A1(n11041), .A2(n11040), .ZN(n11067) );
  NAND2_X1 U11014 ( .A1(n11040), .A2(n11041), .ZN(n11064) );
  NAND2_X1 U11015 ( .A1(n11068), .A2(n11069), .ZN(n11041) );
  NAND3_X1 U11016 ( .A1(n9277), .A2(n11070), .A3(n10667), .ZN(n11069) );
  INV_X1 U11017 ( .A(n11071), .ZN(n11070) );
  NOR2_X1 U11018 ( .A1(n11037), .A2(n11035), .ZN(n11071) );
  NAND2_X1 U11019 ( .A1(n11035), .A2(n11037), .ZN(n11068) );
  NAND2_X1 U11020 ( .A1(n11072), .A2(n11073), .ZN(n11037) );
  NAND3_X1 U11021 ( .A1(n10307), .A2(n11074), .A3(n10667), .ZN(n11073) );
  INV_X1 U11022 ( .A(n11075), .ZN(n11074) );
  NOR2_X1 U11023 ( .A1(n11033), .A2(n11031), .ZN(n11075) );
  NAND2_X1 U11024 ( .A1(n11031), .A2(n11033), .ZN(n11072) );
  NAND2_X1 U11025 ( .A1(n11029), .A2(n11076), .ZN(n11033) );
  NAND2_X1 U11026 ( .A1(n11028), .A2(n11030), .ZN(n11076) );
  NAND2_X1 U11027 ( .A1(n11077), .A2(n11078), .ZN(n11030) );
  NAND2_X1 U11028 ( .A1(n10667), .A2(n9286), .ZN(n11078) );
  XNOR2_X1 U11029 ( .A(n11079), .B(n11080), .ZN(n11028) );
  XNOR2_X1 U11030 ( .A(n11081), .B(n11082), .ZN(n11079) );
  NAND2_X1 U11031 ( .A1(n9286), .A2(n11083), .ZN(n11029) );
  INV_X1 U11032 ( .A(n11077), .ZN(n11083) );
  NOR2_X1 U11033 ( .A1(n11084), .A2(n11085), .ZN(n11077) );
  NOR3_X1 U11034 ( .A1(n8544), .A2(n11086), .A3(n8576), .ZN(n11085) );
  INV_X1 U11035 ( .A(n11087), .ZN(n11086) );
  NAND2_X1 U11036 ( .A1(n11025), .A2(n11024), .ZN(n11087) );
  NOR2_X1 U11037 ( .A1(n11024), .A2(n11025), .ZN(n11084) );
  NOR2_X1 U11038 ( .A1(n11088), .A2(n11089), .ZN(n11025) );
  INV_X1 U11039 ( .A(n11090), .ZN(n11089) );
  NAND2_X1 U11040 ( .A1(n11022), .A2(n11091), .ZN(n11090) );
  NAND2_X1 U11041 ( .A1(n11021), .A2(n11020), .ZN(n11091) );
  NOR2_X1 U11042 ( .A1(n8576), .A2(n8560), .ZN(n11022) );
  NOR2_X1 U11043 ( .A1(n11020), .A2(n11021), .ZN(n11088) );
  NOR2_X1 U11044 ( .A1(n11092), .A2(n11093), .ZN(n11021) );
  NOR3_X1 U11045 ( .A1(n9014), .A2(n11094), .A3(n8576), .ZN(n11093) );
  NOR2_X1 U11046 ( .A1(n11017), .A2(n11016), .ZN(n11094) );
  INV_X1 U11047 ( .A(n11095), .ZN(n11092) );
  NAND2_X1 U11048 ( .A1(n11016), .A2(n11017), .ZN(n11095) );
  NAND2_X1 U11049 ( .A1(n11096), .A2(n11097), .ZN(n11017) );
  INV_X1 U11050 ( .A(n11098), .ZN(n11097) );
  NOR3_X1 U11051 ( .A1(n9020), .A2(n11099), .A3(n8576), .ZN(n11098) );
  NOR2_X1 U11052 ( .A1(n11013), .A2(n11011), .ZN(n11099) );
  NAND2_X1 U11053 ( .A1(n11011), .A2(n11013), .ZN(n11096) );
  NAND2_X1 U11054 ( .A1(n11100), .A2(n11101), .ZN(n11013) );
  NAND3_X1 U11055 ( .A1(n9209), .A2(n11102), .A3(n10667), .ZN(n11101) );
  INV_X1 U11056 ( .A(n11103), .ZN(n11102) );
  NOR2_X1 U11057 ( .A1(n11009), .A2(n11008), .ZN(n11103) );
  NAND2_X1 U11058 ( .A1(n11008), .A2(n11009), .ZN(n11100) );
  NAND2_X1 U11059 ( .A1(n11104), .A2(n11105), .ZN(n11009) );
  NAND2_X1 U11060 ( .A1(n11006), .A2(n11106), .ZN(n11105) );
  NAND2_X1 U11061 ( .A1(n11005), .A2(n11003), .ZN(n11106) );
  NOR2_X1 U11062 ( .A1(n8576), .A2(n8582), .ZN(n11006) );
  INV_X1 U11063 ( .A(n11107), .ZN(n11104) );
  NOR2_X1 U11064 ( .A1(n11003), .A2(n11005), .ZN(n11107) );
  NOR2_X1 U11065 ( .A1(n11108), .A2(n11109), .ZN(n11005) );
  INV_X1 U11066 ( .A(n11110), .ZN(n11109) );
  NAND3_X1 U11067 ( .A1(n9721), .A2(n11111), .A3(n10667), .ZN(n11110) );
  NAND2_X1 U11068 ( .A1(n11001), .A2(n11000), .ZN(n11111) );
  NOR2_X1 U11069 ( .A1(n11000), .A2(n11001), .ZN(n11108) );
  NOR2_X1 U11070 ( .A1(n11112), .A2(n11113), .ZN(n11001) );
  INV_X1 U11071 ( .A(n11114), .ZN(n11113) );
  NAND2_X1 U11072 ( .A1(n10998), .A2(n11115), .ZN(n11114) );
  NAND2_X1 U11073 ( .A1(n10997), .A2(n10996), .ZN(n11115) );
  NOR2_X1 U11074 ( .A1(n8576), .A2(n8562), .ZN(n10998) );
  NOR2_X1 U11075 ( .A1(n10996), .A2(n10997), .ZN(n11112) );
  NOR2_X1 U11076 ( .A1(n11116), .A2(n11117), .ZN(n10997) );
  NOR3_X1 U11077 ( .A1(n8545), .A2(n11118), .A3(n8576), .ZN(n11117) );
  NOR2_X1 U11078 ( .A1(n10993), .A2(n10992), .ZN(n11118) );
  INV_X1 U11079 ( .A(n11119), .ZN(n11116) );
  NAND2_X1 U11080 ( .A1(n10992), .A2(n10993), .ZN(n11119) );
  NAND2_X1 U11081 ( .A1(n11120), .A2(n11121), .ZN(n10993) );
  NAND2_X1 U11082 ( .A1(n10990), .A2(n11122), .ZN(n11121) );
  NAND2_X1 U11083 ( .A1(n10989), .A2(n10987), .ZN(n11122) );
  NOR2_X1 U11084 ( .A1(n8576), .A2(n8569), .ZN(n10990) );
  INV_X1 U11085 ( .A(n11123), .ZN(n11120) );
  NOR2_X1 U11086 ( .A1(n10987), .A2(n10989), .ZN(n11123) );
  NOR2_X1 U11087 ( .A1(n11124), .A2(n11125), .ZN(n10989) );
  INV_X1 U11088 ( .A(n11126), .ZN(n11125) );
  NAND2_X1 U11089 ( .A1(n10986), .A2(n11127), .ZN(n11126) );
  NAND2_X1 U11090 ( .A1(n10985), .A2(n10984), .ZN(n11127) );
  NOR2_X1 U11091 ( .A1(n8576), .A2(n8593), .ZN(n10986) );
  NOR2_X1 U11092 ( .A1(n10984), .A2(n10985), .ZN(n11124) );
  NOR2_X1 U11093 ( .A1(n11128), .A2(n11129), .ZN(n10985) );
  INV_X1 U11094 ( .A(n11130), .ZN(n11129) );
  NAND2_X1 U11095 ( .A1(n10982), .A2(n11131), .ZN(n11130) );
  NAND2_X1 U11096 ( .A1(n10981), .A2(n10980), .ZN(n11131) );
  NOR2_X1 U11097 ( .A1(n8576), .A2(n8583), .ZN(n10982) );
  NOR2_X1 U11098 ( .A1(n10980), .A2(n10981), .ZN(n11128) );
  NOR2_X1 U11099 ( .A1(n11132), .A2(n11133), .ZN(n10981) );
  INV_X1 U11100 ( .A(n11134), .ZN(n11133) );
  NAND2_X1 U11101 ( .A1(n10977), .A2(n11135), .ZN(n11134) );
  NAND2_X1 U11102 ( .A1(n10978), .A2(n10976), .ZN(n11135) );
  NOR2_X1 U11103 ( .A1(n8576), .A2(n8580), .ZN(n10977) );
  NOR2_X1 U11104 ( .A1(n10976), .A2(n10978), .ZN(n11132) );
  NOR2_X1 U11105 ( .A1(n11136), .A2(n11137), .ZN(n10978) );
  INV_X1 U11106 ( .A(n11138), .ZN(n11137) );
  NAND2_X1 U11107 ( .A1(n10974), .A2(n11139), .ZN(n11138) );
  NAND2_X1 U11108 ( .A1(n10973), .A2(n10972), .ZN(n11139) );
  NOR2_X1 U11109 ( .A1(n8576), .A2(n8588), .ZN(n10974) );
  NOR2_X1 U11110 ( .A1(n10972), .A2(n10973), .ZN(n11136) );
  NOR2_X1 U11111 ( .A1(n11140), .A2(n11141), .ZN(n10973) );
  INV_X1 U11112 ( .A(n11142), .ZN(n11141) );
  NAND2_X1 U11113 ( .A1(n10969), .A2(n11143), .ZN(n11142) );
  NAND2_X1 U11114 ( .A1(n10970), .A2(n10968), .ZN(n11143) );
  NOR2_X1 U11115 ( .A1(n8576), .A2(n8551), .ZN(n10969) );
  NOR2_X1 U11116 ( .A1(n10968), .A2(n10970), .ZN(n11140) );
  NOR2_X1 U11117 ( .A1(n11144), .A2(n11145), .ZN(n10970) );
  INV_X1 U11118 ( .A(n11146), .ZN(n11145) );
  NAND2_X1 U11119 ( .A1(n10966), .A2(n11147), .ZN(n11146) );
  NAND2_X1 U11120 ( .A1(n10965), .A2(n10964), .ZN(n11147) );
  NOR2_X1 U11121 ( .A1(n8576), .A2(n8563), .ZN(n10966) );
  NOR2_X1 U11122 ( .A1(n10964), .A2(n10965), .ZN(n11144) );
  NOR2_X1 U11123 ( .A1(n11148), .A2(n11149), .ZN(n10965) );
  INV_X1 U11124 ( .A(n11150), .ZN(n11149) );
  NAND2_X1 U11125 ( .A1(n10962), .A2(n11151), .ZN(n11150) );
  NAND2_X1 U11126 ( .A1(n10961), .A2(n10959), .ZN(n11151) );
  NOR2_X1 U11127 ( .A1(n10666), .A2(n8548), .ZN(n10962) );
  NOR2_X1 U11128 ( .A1(n10959), .A2(n10961), .ZN(n11148) );
  NOR2_X1 U11129 ( .A1(n11152), .A2(n11153), .ZN(n10961) );
  INV_X1 U11130 ( .A(n11154), .ZN(n11153) );
  NAND2_X1 U11131 ( .A1(n10958), .A2(n11155), .ZN(n11154) );
  NAND2_X1 U11132 ( .A1(n10957), .A2(n10956), .ZN(n11155) );
  NOR2_X1 U11133 ( .A1(n10666), .A2(n8584), .ZN(n10958) );
  NOR2_X1 U11134 ( .A1(n10956), .A2(n10957), .ZN(n11152) );
  NOR2_X1 U11135 ( .A1(n11156), .A2(n11157), .ZN(n10957) );
  INV_X1 U11136 ( .A(n11158), .ZN(n11157) );
  NAND2_X1 U11137 ( .A1(n10953), .A2(n11159), .ZN(n11158) );
  NAND2_X1 U11138 ( .A1(n10954), .A2(n10952), .ZN(n11159) );
  NOR2_X1 U11139 ( .A1(n10666), .A2(n8535), .ZN(n10953) );
  NOR2_X1 U11140 ( .A1(n10952), .A2(n10954), .ZN(n11156) );
  NOR2_X1 U11141 ( .A1(n11160), .A2(n11161), .ZN(n10954) );
  INV_X1 U11142 ( .A(n11162), .ZN(n11161) );
  NAND2_X1 U11143 ( .A1(n10949), .A2(n11163), .ZN(n11162) );
  NAND2_X1 U11144 ( .A1(n10950), .A2(n10948), .ZN(n11163) );
  NOR2_X1 U11145 ( .A1(n10666), .A2(n8568), .ZN(n10949) );
  NOR2_X1 U11146 ( .A1(n10948), .A2(n10950), .ZN(n11160) );
  NOR2_X1 U11147 ( .A1(n11164), .A2(n11165), .ZN(n10950) );
  INV_X1 U11148 ( .A(n11166), .ZN(n11165) );
  NAND2_X1 U11149 ( .A1(n10945), .A2(n11167), .ZN(n11166) );
  NAND2_X1 U11150 ( .A1(n10946), .A2(n10944), .ZN(n11167) );
  NOR2_X1 U11151 ( .A1(n10666), .A2(n8574), .ZN(n10945) );
  NOR2_X1 U11152 ( .A1(n10944), .A2(n10946), .ZN(n11164) );
  NOR2_X1 U11153 ( .A1(n11168), .A2(n11169), .ZN(n10946) );
  INV_X1 U11154 ( .A(n11170), .ZN(n11169) );
  NAND2_X1 U11155 ( .A1(n10941), .A2(n11171), .ZN(n11170) );
  NAND2_X1 U11156 ( .A1(n10942), .A2(n10940), .ZN(n11171) );
  NOR2_X1 U11157 ( .A1(n10666), .A2(n8565), .ZN(n10941) );
  NOR2_X1 U11158 ( .A1(n10940), .A2(n10942), .ZN(n11168) );
  NOR2_X1 U11159 ( .A1(n11172), .A2(n11173), .ZN(n10942) );
  INV_X1 U11160 ( .A(n11174), .ZN(n11173) );
  NAND2_X1 U11161 ( .A1(n10935), .A2(n11175), .ZN(n11174) );
  NAND2_X1 U11162 ( .A1(n10938), .A2(n10937), .ZN(n11175) );
  NOR2_X1 U11163 ( .A1(n10666), .A2(n8567), .ZN(n10935) );
  NOR2_X1 U11164 ( .A1(n10937), .A2(n10938), .ZN(n11172) );
  INV_X1 U11165 ( .A(n11176), .ZN(n10938) );
  NAND2_X1 U11166 ( .A1(n11177), .A2(n11178), .ZN(n11176) );
  NAND2_X1 U11167 ( .A1(n8546), .A2(n11179), .ZN(n11178) );
  NAND2_X1 U11168 ( .A1(n8624), .A2(n11180), .ZN(n11179) );
  NAND2_X1 U11169 ( .A1(n8559), .A2(n8585), .ZN(n11180) );
  NAND2_X1 U11170 ( .A1(n11182), .A2(n11183), .ZN(n11177) );
  NAND2_X1 U11171 ( .A1(n8630), .A2(n11184), .ZN(n11183) );
  NAND2_X1 U11172 ( .A1(n8539), .A2(n8547), .ZN(n11184) );
  NAND3_X1 U11173 ( .A1(n10667), .A2(n8537), .A3(n8546), .ZN(n10937) );
  INV_X1 U11174 ( .A(n10666), .ZN(n10667) );
  XNOR2_X1 U11175 ( .A(n11185), .B(n11186), .ZN(n10666) );
  XOR2_X1 U11176 ( .A(d_23_), .B(c_23_), .Z(n11186) );
  XOR2_X1 U11177 ( .A(n11187), .B(n11188), .Z(n10940) );
  XNOR2_X1 U11178 ( .A(n11189), .B(n11190), .ZN(n11188) );
  XOR2_X1 U11179 ( .A(n11191), .B(n11192), .Z(n10944) );
  XNOR2_X1 U11180 ( .A(n11193), .B(n11194), .ZN(n11191) );
  XOR2_X1 U11181 ( .A(n11195), .B(n11196), .Z(n10948) );
  XNOR2_X1 U11182 ( .A(n11197), .B(n11198), .ZN(n11195) );
  XOR2_X1 U11183 ( .A(n11199), .B(n11200), .Z(n10952) );
  XNOR2_X1 U11184 ( .A(n11201), .B(n11202), .ZN(n11199) );
  XOR2_X1 U11185 ( .A(n11203), .B(n11204), .Z(n10956) );
  XNOR2_X1 U11186 ( .A(n11205), .B(n11206), .ZN(n11203) );
  NOR2_X1 U11187 ( .A1(n8535), .A2(n8547), .ZN(n11206) );
  XOR2_X1 U11188 ( .A(n11207), .B(n11208), .Z(n10959) );
  XNOR2_X1 U11189 ( .A(n11209), .B(n11210), .ZN(n11207) );
  NOR2_X1 U11190 ( .A1(n8584), .A2(n8547), .ZN(n11210) );
  XOR2_X1 U11191 ( .A(n11211), .B(n11212), .Z(n10964) );
  XNOR2_X1 U11192 ( .A(n11213), .B(n11214), .ZN(n11211) );
  NOR2_X1 U11193 ( .A1(n8548), .A2(n8547), .ZN(n11214) );
  XOR2_X1 U11194 ( .A(n11215), .B(n11216), .Z(n10968) );
  XNOR2_X1 U11195 ( .A(n11217), .B(n11218), .ZN(n11215) );
  NOR2_X1 U11196 ( .A1(n8563), .A2(n8547), .ZN(n11218) );
  XOR2_X1 U11197 ( .A(n11219), .B(n11220), .Z(n10972) );
  XNOR2_X1 U11198 ( .A(n11221), .B(n11222), .ZN(n11219) );
  NOR2_X1 U11199 ( .A1(n8551), .A2(n8547), .ZN(n11222) );
  XOR2_X1 U11200 ( .A(n11223), .B(n11224), .Z(n10976) );
  XNOR2_X1 U11201 ( .A(n11225), .B(n11226), .ZN(n11223) );
  NOR2_X1 U11202 ( .A1(n8588), .A2(n8547), .ZN(n11226) );
  XNOR2_X1 U11203 ( .A(n11227), .B(n11228), .ZN(n10980) );
  XNOR2_X1 U11204 ( .A(n11229), .B(n11230), .ZN(n11228) );
  NAND2_X1 U11205 ( .A1(n8546), .A2(n9070), .ZN(n11230) );
  XOR2_X1 U11206 ( .A(n11231), .B(n11232), .Z(n10984) );
  XNOR2_X1 U11207 ( .A(n11233), .B(n11234), .ZN(n11231) );
  NOR2_X1 U11208 ( .A1(n8583), .A2(n8547), .ZN(n11234) );
  XOR2_X1 U11209 ( .A(n11235), .B(n11236), .Z(n10987) );
  XNOR2_X1 U11210 ( .A(n11237), .B(n11238), .ZN(n11235) );
  NOR2_X1 U11211 ( .A1(n8593), .A2(n8547), .ZN(n11238) );
  XNOR2_X1 U11212 ( .A(n11239), .B(n11240), .ZN(n10992) );
  XNOR2_X1 U11213 ( .A(n11241), .B(n11242), .ZN(n11239) );
  NOR2_X1 U11214 ( .A1(n9050), .A2(n8547), .ZN(n11242) );
  XOR2_X1 U11215 ( .A(n11243), .B(n11244), .Z(n10996) );
  XNOR2_X1 U11216 ( .A(n11245), .B(n11246), .ZN(n11243) );
  NOR2_X1 U11217 ( .A1(n8545), .A2(n8547), .ZN(n11246) );
  XOR2_X1 U11218 ( .A(n11247), .B(n11248), .Z(n11000) );
  XNOR2_X1 U11219 ( .A(n11249), .B(n11250), .ZN(n11247) );
  NOR2_X1 U11220 ( .A1(n9041), .A2(n8547), .ZN(n11250) );
  XOR2_X1 U11221 ( .A(n11251), .B(n11252), .Z(n11003) );
  XNOR2_X1 U11222 ( .A(n11253), .B(n11254), .ZN(n11251) );
  NOR2_X1 U11223 ( .A1(n8591), .A2(n8547), .ZN(n11254) );
  XNOR2_X1 U11224 ( .A(n11255), .B(n11256), .ZN(n11008) );
  XNOR2_X1 U11225 ( .A(n11257), .B(n11258), .ZN(n11255) );
  NOR2_X1 U11226 ( .A1(n8582), .A2(n8547), .ZN(n11258) );
  XNOR2_X1 U11227 ( .A(n11259), .B(n11260), .ZN(n11011) );
  XNOR2_X1 U11228 ( .A(n11261), .B(n11262), .ZN(n11259) );
  NOR2_X1 U11229 ( .A1(n8572), .A2(n8547), .ZN(n11262) );
  XNOR2_X1 U11230 ( .A(n11263), .B(n11264), .ZN(n11016) );
  XNOR2_X1 U11231 ( .A(n11265), .B(n11266), .ZN(n11263) );
  NOR2_X1 U11232 ( .A1(n8556), .A2(n8547), .ZN(n11266) );
  XOR2_X1 U11233 ( .A(n11267), .B(n11268), .Z(n11020) );
  XNOR2_X1 U11234 ( .A(n11269), .B(n11270), .ZN(n11267) );
  NOR2_X1 U11235 ( .A1(n8594), .A2(n8547), .ZN(n11270) );
  XOR2_X1 U11236 ( .A(n11271), .B(n11272), .Z(n11024) );
  XNOR2_X1 U11237 ( .A(n11273), .B(n11274), .ZN(n11271) );
  NOR2_X1 U11238 ( .A1(n8560), .A2(n8547), .ZN(n11274) );
  XOR2_X1 U11239 ( .A(n11275), .B(n11276), .Z(n11031) );
  XOR2_X1 U11240 ( .A(n11277), .B(n11278), .Z(n11275) );
  XOR2_X1 U11241 ( .A(n11279), .B(n11280), .Z(n11035) );
  XOR2_X1 U11242 ( .A(n11281), .B(n11282), .Z(n11279) );
  XNOR2_X1 U11243 ( .A(n11283), .B(n11284), .ZN(n11040) );
  XOR2_X1 U11244 ( .A(n11285), .B(n11286), .Z(n11284) );
  XNOR2_X1 U11245 ( .A(n11287), .B(n11288), .ZN(n11044) );
  XNOR2_X1 U11246 ( .A(n11289), .B(n11290), .ZN(n11287) );
  XNOR2_X1 U11247 ( .A(n11291), .B(n11292), .ZN(n11051) );
  XNOR2_X1 U11248 ( .A(n11293), .B(n11294), .ZN(n11291) );
  XOR2_X1 U11249 ( .A(n11295), .B(n11296), .Z(n10799) );
  XNOR2_X1 U11250 ( .A(n11297), .B(n11298), .ZN(n11295) );
  NAND2_X1 U11251 ( .A1(n11299), .A2(n11300), .ZN(n8817) );
  NAND2_X1 U11252 ( .A1(n8937), .A2(n8936), .ZN(n11300) );
  XNOR2_X1 U11253 ( .A(n8928), .B(n8929), .ZN(n11299) );
  NAND3_X1 U11254 ( .A1(n11301), .A2(n8936), .A3(n8937), .ZN(n8818) );
  XOR2_X1 U11255 ( .A(n11302), .B(n11303), .Z(n8937) );
  XNOR2_X1 U11256 ( .A(n11304), .B(n11305), .ZN(n11303) );
  NAND2_X1 U11257 ( .A1(n11182), .A2(n8872), .ZN(n11305) );
  NAND2_X1 U11258 ( .A1(n11306), .A2(n11307), .ZN(n8936) );
  INV_X1 U11259 ( .A(n11308), .ZN(n11307) );
  NOR3_X1 U11260 ( .A1(n8972), .A2(n11309), .A3(n8547), .ZN(n11308) );
  NOR2_X1 U11261 ( .A1(n10801), .A2(n10802), .ZN(n11309) );
  NAND2_X1 U11262 ( .A1(n10801), .A2(n10802), .ZN(n11306) );
  NAND2_X1 U11263 ( .A1(n11310), .A2(n11311), .ZN(n10802) );
  NAND2_X1 U11264 ( .A1(n11298), .A2(n11312), .ZN(n11311) );
  NAND2_X1 U11265 ( .A1(n11296), .A2(n11297), .ZN(n11312) );
  NOR2_X1 U11266 ( .A1(n8547), .A2(n8589), .ZN(n11298) );
  INV_X1 U11267 ( .A(n11313), .ZN(n11310) );
  NOR2_X1 U11268 ( .A1(n11296), .A2(n11297), .ZN(n11313) );
  NOR2_X1 U11269 ( .A1(n11314), .A2(n11315), .ZN(n11297) );
  INV_X1 U11270 ( .A(n11316), .ZN(n11315) );
  NAND2_X1 U11271 ( .A1(n11293), .A2(n11317), .ZN(n11316) );
  NAND2_X1 U11272 ( .A1(n11294), .A2(n11292), .ZN(n11317) );
  NOR2_X1 U11273 ( .A1(n8547), .A2(n8552), .ZN(n11293) );
  NOR2_X1 U11274 ( .A1(n11292), .A2(n11294), .ZN(n11314) );
  NOR2_X1 U11275 ( .A1(n11318), .A2(n11319), .ZN(n11294) );
  INV_X1 U11276 ( .A(n11320), .ZN(n11319) );
  NAND2_X1 U11277 ( .A1(n11290), .A2(n11321), .ZN(n11320) );
  NAND2_X1 U11278 ( .A1(n11289), .A2(n11288), .ZN(n11321) );
  NOR2_X1 U11279 ( .A1(n8547), .A2(n8527), .ZN(n11290) );
  NOR2_X1 U11280 ( .A1(n11288), .A2(n11289), .ZN(n11318) );
  NOR2_X1 U11281 ( .A1(n11322), .A2(n11323), .ZN(n11289) );
  NOR2_X1 U11282 ( .A1(n11286), .A2(n11324), .ZN(n11323) );
  NOR2_X1 U11283 ( .A1(n11285), .A2(n11283), .ZN(n11324) );
  NAND2_X1 U11284 ( .A1(n8546), .A2(n9277), .ZN(n11286) );
  INV_X1 U11285 ( .A(n11325), .ZN(n11322) );
  NAND2_X1 U11286 ( .A1(n11283), .A2(n11285), .ZN(n11325) );
  NAND2_X1 U11287 ( .A1(n11326), .A2(n11327), .ZN(n11285) );
  NAND2_X1 U11288 ( .A1(n11282), .A2(n11328), .ZN(n11327) );
  INV_X1 U11289 ( .A(n11329), .ZN(n11328) );
  NOR2_X1 U11290 ( .A1(n11280), .A2(n11281), .ZN(n11329) );
  NOR2_X1 U11291 ( .A1(n8547), .A2(n8564), .ZN(n11282) );
  NAND2_X1 U11292 ( .A1(n11280), .A2(n11281), .ZN(n11326) );
  NAND2_X1 U11293 ( .A1(n11330), .A2(n11331), .ZN(n11281) );
  NAND2_X1 U11294 ( .A1(n11278), .A2(n11332), .ZN(n11331) );
  INV_X1 U11295 ( .A(n11333), .ZN(n11332) );
  NOR2_X1 U11296 ( .A1(n11276), .A2(n11277), .ZN(n11333) );
  NOR2_X1 U11297 ( .A1(n8547), .A2(n8555), .ZN(n11278) );
  NAND2_X1 U11298 ( .A1(n11276), .A2(n11277), .ZN(n11330) );
  NAND2_X1 U11299 ( .A1(n11334), .A2(n11335), .ZN(n11277) );
  NAND2_X1 U11300 ( .A1(n11082), .A2(n11336), .ZN(n11335) );
  NAND2_X1 U11301 ( .A1(n11080), .A2(n11081), .ZN(n11336) );
  NOR2_X1 U11302 ( .A1(n8547), .A2(n8544), .ZN(n11082) );
  INV_X1 U11303 ( .A(n11337), .ZN(n11334) );
  NOR2_X1 U11304 ( .A1(n11080), .A2(n11081), .ZN(n11337) );
  NOR2_X1 U11305 ( .A1(n11338), .A2(n11339), .ZN(n11081) );
  INV_X1 U11306 ( .A(n11340), .ZN(n11339) );
  NAND3_X1 U11307 ( .A1(n9295), .A2(n11341), .A3(n8546), .ZN(n11340) );
  NAND2_X1 U11308 ( .A1(n11272), .A2(n11273), .ZN(n11341) );
  NOR2_X1 U11309 ( .A1(n11272), .A2(n11273), .ZN(n11338) );
  NOR2_X1 U11310 ( .A1(n11342), .A2(n11343), .ZN(n11273) );
  INV_X1 U11311 ( .A(n11344), .ZN(n11343) );
  NAND3_X1 U11312 ( .A1(n10846), .A2(n11345), .A3(n8546), .ZN(n11344) );
  NAND2_X1 U11313 ( .A1(n11268), .A2(n11269), .ZN(n11345) );
  NOR2_X1 U11314 ( .A1(n11268), .A2(n11269), .ZN(n11342) );
  NOR2_X1 U11315 ( .A1(n11346), .A2(n11347), .ZN(n11269) );
  INV_X1 U11316 ( .A(n11348), .ZN(n11347) );
  NAND3_X1 U11317 ( .A1(n9304), .A2(n11349), .A3(n8546), .ZN(n11348) );
  NAND2_X1 U11318 ( .A1(n11265), .A2(n11264), .ZN(n11349) );
  NOR2_X1 U11319 ( .A1(n11264), .A2(n11265), .ZN(n11346) );
  NOR2_X1 U11320 ( .A1(n11350), .A2(n11351), .ZN(n11265) );
  NOR3_X1 U11321 ( .A1(n9025), .A2(n11352), .A3(n8547), .ZN(n11351) );
  INV_X1 U11322 ( .A(n11353), .ZN(n11352) );
  NAND2_X1 U11323 ( .A1(n11260), .A2(n11261), .ZN(n11353) );
  NOR2_X1 U11324 ( .A1(n11260), .A2(n11261), .ZN(n11350) );
  NOR2_X1 U11325 ( .A1(n11354), .A2(n11355), .ZN(n11261) );
  INV_X1 U11326 ( .A(n11356), .ZN(n11355) );
  NAND3_X1 U11327 ( .A1(n9313), .A2(n11357), .A3(n8546), .ZN(n11356) );
  NAND2_X1 U11328 ( .A1(n11257), .A2(n11256), .ZN(n11357) );
  NOR2_X1 U11329 ( .A1(n11256), .A2(n11257), .ZN(n11354) );
  NOR2_X1 U11330 ( .A1(n11358), .A2(n11359), .ZN(n11257) );
  NOR3_X1 U11331 ( .A1(n9036), .A2(n11360), .A3(n8547), .ZN(n11359) );
  INV_X1 U11332 ( .A(n11361), .ZN(n11360) );
  NAND2_X1 U11333 ( .A1(n11252), .A2(n11253), .ZN(n11361) );
  NOR2_X1 U11334 ( .A1(n11252), .A2(n11253), .ZN(n11358) );
  NOR2_X1 U11335 ( .A1(n11362), .A2(n11363), .ZN(n11253) );
  INV_X1 U11336 ( .A(n11364), .ZN(n11363) );
  NAND3_X1 U11337 ( .A1(n9322), .A2(n11365), .A3(n8546), .ZN(n11364) );
  NAND2_X1 U11338 ( .A1(n11249), .A2(n11248), .ZN(n11365) );
  NOR2_X1 U11339 ( .A1(n11248), .A2(n11249), .ZN(n11362) );
  NOR2_X1 U11340 ( .A1(n11366), .A2(n11367), .ZN(n11249) );
  NOR3_X1 U11341 ( .A1(n8545), .A2(n11368), .A3(n8547), .ZN(n11367) );
  INV_X1 U11342 ( .A(n11369), .ZN(n11368) );
  NAND2_X1 U11343 ( .A1(n11244), .A2(n11245), .ZN(n11369) );
  NOR2_X1 U11344 ( .A1(n11244), .A2(n11245), .ZN(n11366) );
  NOR2_X1 U11345 ( .A1(n11370), .A2(n11371), .ZN(n11245) );
  INV_X1 U11346 ( .A(n11372), .ZN(n11371) );
  NAND3_X1 U11347 ( .A1(n9331), .A2(n11373), .A3(n8546), .ZN(n11372) );
  NAND2_X1 U11348 ( .A1(n11241), .A2(n11240), .ZN(n11373) );
  NOR2_X1 U11349 ( .A1(n11240), .A2(n11241), .ZN(n11370) );
  NOR2_X1 U11350 ( .A1(n11374), .A2(n11375), .ZN(n11241) );
  NOR3_X1 U11351 ( .A1(n9056), .A2(n11376), .A3(n8547), .ZN(n11375) );
  INV_X1 U11352 ( .A(n11377), .ZN(n11376) );
  NAND2_X1 U11353 ( .A1(n11236), .A2(n11237), .ZN(n11377) );
  NOR2_X1 U11354 ( .A1(n11236), .A2(n11237), .ZN(n11374) );
  NOR2_X1 U11355 ( .A1(n11378), .A2(n11379), .ZN(n11237) );
  INV_X1 U11356 ( .A(n11380), .ZN(n11379) );
  NAND3_X1 U11357 ( .A1(n9340), .A2(n11381), .A3(n8546), .ZN(n11380) );
  NAND2_X1 U11358 ( .A1(n11233), .A2(n11232), .ZN(n11381) );
  NOR2_X1 U11359 ( .A1(n11232), .A2(n11233), .ZN(n11378) );
  NOR2_X1 U11360 ( .A1(n11382), .A2(n11383), .ZN(n11233) );
  NOR3_X1 U11361 ( .A1(n9066), .A2(n11384), .A3(n8547), .ZN(n11383) );
  INV_X1 U11362 ( .A(n11385), .ZN(n11384) );
  NAND2_X1 U11363 ( .A1(n11227), .A2(n11229), .ZN(n11385) );
  NOR2_X1 U11364 ( .A1(n11227), .A2(n11229), .ZN(n11382) );
  NOR2_X1 U11365 ( .A1(n11386), .A2(n11387), .ZN(n11229) );
  INV_X1 U11366 ( .A(n11388), .ZN(n11387) );
  NAND3_X1 U11367 ( .A1(n9080), .A2(n11389), .A3(n8546), .ZN(n11388) );
  NAND2_X1 U11368 ( .A1(n11225), .A2(n11224), .ZN(n11389) );
  NOR2_X1 U11369 ( .A1(n11224), .A2(n11225), .ZN(n11386) );
  NOR2_X1 U11370 ( .A1(n11390), .A2(n11391), .ZN(n11225) );
  NOR3_X1 U11371 ( .A1(n8551), .A2(n11392), .A3(n8547), .ZN(n11391) );
  INV_X1 U11372 ( .A(n11393), .ZN(n11392) );
  NAND2_X1 U11373 ( .A1(n11220), .A2(n11221), .ZN(n11393) );
  NOR2_X1 U11374 ( .A1(n11220), .A2(n11221), .ZN(n11390) );
  NOR2_X1 U11375 ( .A1(n11394), .A2(n11395), .ZN(n11221) );
  INV_X1 U11376 ( .A(n11396), .ZN(n11395) );
  NAND3_X1 U11377 ( .A1(n9098), .A2(n11397), .A3(n8546), .ZN(n11396) );
  NAND2_X1 U11378 ( .A1(n11217), .A2(n11216), .ZN(n11397) );
  NOR2_X1 U11379 ( .A1(n11216), .A2(n11217), .ZN(n11394) );
  NOR2_X1 U11380 ( .A1(n11398), .A2(n11399), .ZN(n11217) );
  NOR3_X1 U11381 ( .A1(n8548), .A2(n11400), .A3(n8547), .ZN(n11399) );
  INV_X1 U11382 ( .A(n11401), .ZN(n11400) );
  NAND2_X1 U11383 ( .A1(n11212), .A2(n11213), .ZN(n11401) );
  NOR2_X1 U11384 ( .A1(n11212), .A2(n11213), .ZN(n11398) );
  NOR2_X1 U11385 ( .A1(n11402), .A2(n11403), .ZN(n11213) );
  INV_X1 U11386 ( .A(n11404), .ZN(n11403) );
  NAND3_X1 U11387 ( .A1(n9112), .A2(n11405), .A3(n8546), .ZN(n11404) );
  NAND2_X1 U11388 ( .A1(n11209), .A2(n11208), .ZN(n11405) );
  NOR2_X1 U11389 ( .A1(n11208), .A2(n11209), .ZN(n11402) );
  NOR2_X1 U11390 ( .A1(n11406), .A2(n11407), .ZN(n11209) );
  INV_X1 U11391 ( .A(n11408), .ZN(n11407) );
  NAND3_X1 U11392 ( .A1(n9121), .A2(n11409), .A3(n8546), .ZN(n11408) );
  NAND2_X1 U11393 ( .A1(n11204), .A2(n11205), .ZN(n11409) );
  NOR2_X1 U11394 ( .A1(n11204), .A2(n11205), .ZN(n11406) );
  NOR2_X1 U11395 ( .A1(n11410), .A2(n11411), .ZN(n11205) );
  INV_X1 U11396 ( .A(n11412), .ZN(n11411) );
  NAND2_X1 U11397 ( .A1(n11202), .A2(n11413), .ZN(n11412) );
  NAND2_X1 U11398 ( .A1(n11201), .A2(n11200), .ZN(n11413) );
  NOR2_X1 U11399 ( .A1(n8547), .A2(n8568), .ZN(n11202) );
  NOR2_X1 U11400 ( .A1(n11200), .A2(n11201), .ZN(n11410) );
  NOR2_X1 U11401 ( .A1(n11414), .A2(n11415), .ZN(n11201) );
  INV_X1 U11402 ( .A(n11416), .ZN(n11415) );
  NAND2_X1 U11403 ( .A1(n11197), .A2(n11417), .ZN(n11416) );
  NAND2_X1 U11404 ( .A1(n11196), .A2(n11198), .ZN(n11417) );
  NOR2_X1 U11405 ( .A1(n8547), .A2(n8574), .ZN(n11197) );
  NOR2_X1 U11406 ( .A1(n11196), .A2(n11198), .ZN(n11414) );
  NOR2_X1 U11407 ( .A1(n11418), .A2(n11419), .ZN(n11198) );
  INV_X1 U11408 ( .A(n11420), .ZN(n11419) );
  NAND2_X1 U11409 ( .A1(n11193), .A2(n11421), .ZN(n11420) );
  NAND2_X1 U11410 ( .A1(n11194), .A2(n11192), .ZN(n11421) );
  NOR2_X1 U11411 ( .A1(n8547), .A2(n8565), .ZN(n11193) );
  NOR2_X1 U11412 ( .A1(n11192), .A2(n11194), .ZN(n11418) );
  NOR2_X1 U11413 ( .A1(n11422), .A2(n11423), .ZN(n11194) );
  INV_X1 U11414 ( .A(n11424), .ZN(n11423) );
  NAND2_X1 U11415 ( .A1(n11187), .A2(n11425), .ZN(n11424) );
  NAND2_X1 U11416 ( .A1(n11190), .A2(n11189), .ZN(n11425) );
  NOR2_X1 U11417 ( .A1(n8547), .A2(n8567), .ZN(n11187) );
  NOR2_X1 U11418 ( .A1(n11189), .A2(n11190), .ZN(n11422) );
  INV_X1 U11419 ( .A(n11426), .ZN(n11190) );
  NAND2_X1 U11420 ( .A1(n11427), .A2(n11428), .ZN(n11426) );
  NAND2_X1 U11421 ( .A1(n11182), .A2(n11429), .ZN(n11428) );
  NAND2_X1 U11422 ( .A1(n8624), .A2(n11430), .ZN(n11429) );
  NAND2_X1 U11423 ( .A1(n8581), .A2(n8585), .ZN(n11430) );
  NAND2_X1 U11424 ( .A1(n11432), .A2(n11433), .ZN(n11427) );
  NAND2_X1 U11425 ( .A1(n8630), .A2(n11434), .ZN(n11433) );
  NAND2_X1 U11426 ( .A1(n8539), .A2(n8559), .ZN(n11434) );
  NAND3_X1 U11427 ( .A1(n11182), .A2(n8537), .A3(n8546), .ZN(n11189) );
  XNOR2_X1 U11428 ( .A(n11435), .B(n11436), .ZN(n10804) );
  XOR2_X1 U11429 ( .A(d_22_), .B(c_22_), .Z(n11436) );
  XOR2_X1 U11430 ( .A(n11437), .B(n11438), .Z(n11192) );
  XNOR2_X1 U11431 ( .A(n11439), .B(n11440), .ZN(n11438) );
  XOR2_X1 U11432 ( .A(n11441), .B(n11442), .Z(n11196) );
  XNOR2_X1 U11433 ( .A(n11443), .B(n11444), .ZN(n11441) );
  XOR2_X1 U11434 ( .A(n11445), .B(n11446), .Z(n11200) );
  XNOR2_X1 U11435 ( .A(n11447), .B(n11448), .ZN(n11445) );
  XOR2_X1 U11436 ( .A(n11449), .B(n11450), .Z(n11204) );
  XNOR2_X1 U11437 ( .A(n11451), .B(n11452), .ZN(n11449) );
  XOR2_X1 U11438 ( .A(n11453), .B(n11454), .Z(n11208) );
  XNOR2_X1 U11439 ( .A(n11455), .B(n11456), .ZN(n11453) );
  XOR2_X1 U11440 ( .A(n11457), .B(n11458), .Z(n11212) );
  XNOR2_X1 U11441 ( .A(n11459), .B(n11460), .ZN(n11457) );
  XOR2_X1 U11442 ( .A(n11461), .B(n11462), .Z(n11216) );
  XNOR2_X1 U11443 ( .A(n11463), .B(n11464), .ZN(n11461) );
  XOR2_X1 U11444 ( .A(n11465), .B(n11466), .Z(n11220) );
  XNOR2_X1 U11445 ( .A(n11467), .B(n11468), .ZN(n11465) );
  XOR2_X1 U11446 ( .A(n11469), .B(n11470), .Z(n11224) );
  XNOR2_X1 U11447 ( .A(n11471), .B(n11472), .ZN(n11469) );
  XOR2_X1 U11448 ( .A(n11473), .B(n11474), .Z(n11227) );
  XNOR2_X1 U11449 ( .A(n11475), .B(n11476), .ZN(n11473) );
  XOR2_X1 U11450 ( .A(n11477), .B(n11478), .Z(n11232) );
  XNOR2_X1 U11451 ( .A(n11479), .B(n11480), .ZN(n11477) );
  XNOR2_X1 U11452 ( .A(n11481), .B(n11482), .ZN(n11236) );
  XOR2_X1 U11453 ( .A(n11483), .B(n11484), .Z(n11482) );
  XNOR2_X1 U11454 ( .A(n11485), .B(n11486), .ZN(n11240) );
  XOR2_X1 U11455 ( .A(n11487), .B(n11488), .Z(n11485) );
  XNOR2_X1 U11456 ( .A(n11489), .B(n11490), .ZN(n11244) );
  XOR2_X1 U11457 ( .A(n11491), .B(n11492), .Z(n11489) );
  XOR2_X1 U11458 ( .A(n11493), .B(n11494), .Z(n11248) );
  XNOR2_X1 U11459 ( .A(n11495), .B(n11496), .ZN(n11493) );
  XNOR2_X1 U11460 ( .A(n11497), .B(n11498), .ZN(n11252) );
  XOR2_X1 U11461 ( .A(n11499), .B(n11500), .Z(n11498) );
  XNOR2_X1 U11462 ( .A(n11501), .B(n11502), .ZN(n11256) );
  XOR2_X1 U11463 ( .A(n11503), .B(n11504), .Z(n11501) );
  XOR2_X1 U11464 ( .A(n11505), .B(n11506), .Z(n11260) );
  XNOR2_X1 U11465 ( .A(n11507), .B(n11508), .ZN(n11506) );
  XNOR2_X1 U11466 ( .A(n11509), .B(n11510), .ZN(n11264) );
  XOR2_X1 U11467 ( .A(n11511), .B(n11512), .Z(n11509) );
  XNOR2_X1 U11468 ( .A(n11513), .B(n11514), .ZN(n11268) );
  XNOR2_X1 U11469 ( .A(n11515), .B(n11516), .ZN(n11514) );
  XOR2_X1 U11470 ( .A(n11517), .B(n11518), .Z(n11272) );
  XNOR2_X1 U11471 ( .A(n11519), .B(n11520), .ZN(n11517) );
  XOR2_X1 U11472 ( .A(n11521), .B(n11522), .Z(n11080) );
  NAND2_X1 U11473 ( .A1(n11523), .A2(n11524), .ZN(n11521) );
  XNOR2_X1 U11474 ( .A(n11525), .B(n11526), .ZN(n11276) );
  XOR2_X1 U11475 ( .A(n11527), .B(n11528), .Z(n11526) );
  NAND2_X1 U11476 ( .A1(n11182), .A2(n8543), .ZN(n11528) );
  XNOR2_X1 U11477 ( .A(n11529), .B(n11530), .ZN(n11280) );
  XOR2_X1 U11478 ( .A(n11531), .B(n11532), .Z(n11530) );
  NAND2_X1 U11479 ( .A1(n11182), .A2(n9286), .ZN(n11532) );
  XOR2_X1 U11480 ( .A(n11533), .B(n11534), .Z(n11283) );
  XOR2_X1 U11481 ( .A(n11535), .B(n11536), .Z(n11533) );
  NOR2_X1 U11482 ( .A1(n8564), .A2(n8559), .ZN(n11536) );
  XOR2_X1 U11483 ( .A(n11537), .B(n11538), .Z(n11288) );
  XOR2_X1 U11484 ( .A(n11539), .B(n11540), .Z(n11538) );
  NAND2_X1 U11485 ( .A1(n11182), .A2(n9277), .ZN(n11540) );
  XOR2_X1 U11486 ( .A(n11541), .B(n11542), .Z(n11292) );
  XOR2_X1 U11487 ( .A(n11543), .B(n11544), .Z(n11542) );
  NAND2_X1 U11488 ( .A1(n11182), .A2(n9792), .ZN(n11544) );
  XOR2_X1 U11489 ( .A(n11545), .B(n11546), .Z(n11296) );
  XOR2_X1 U11490 ( .A(n11547), .B(n11548), .Z(n11546) );
  NAND2_X1 U11491 ( .A1(n11182), .A2(n9268), .ZN(n11548) );
  XOR2_X1 U11492 ( .A(n11549), .B(n11550), .Z(n10801) );
  XNOR2_X1 U11493 ( .A(n11551), .B(n11552), .ZN(n11550) );
  NAND2_X1 U11494 ( .A1(n11182), .A2(n9263), .ZN(n11552) );
  XOR2_X1 U11495 ( .A(n8929), .B(n8928), .Z(n11301) );
  NAND3_X1 U11496 ( .A1(n8928), .A2(n8929), .A3(n11553), .ZN(n8822) );
  XOR2_X1 U11497 ( .A(n8924), .B(n8923), .Z(n11553) );
  NAND2_X1 U11498 ( .A1(n11554), .A2(n11555), .ZN(n8929) );
  NAND3_X1 U11499 ( .A1(n8592), .A2(n11556), .A3(n11182), .ZN(n11555) );
  NAND2_X1 U11500 ( .A1(n11304), .A2(n11302), .ZN(n11556) );
  INV_X1 U11501 ( .A(n11557), .ZN(n11554) );
  NOR2_X1 U11502 ( .A1(n11302), .A2(n11304), .ZN(n11557) );
  NOR2_X1 U11503 ( .A1(n11558), .A2(n11559), .ZN(n11304) );
  INV_X1 U11504 ( .A(n11560), .ZN(n11559) );
  NAND3_X1 U11505 ( .A1(n9263), .A2(n11561), .A3(n11182), .ZN(n11560) );
  NAND2_X1 U11506 ( .A1(n11551), .A2(n11549), .ZN(n11561) );
  NOR2_X1 U11507 ( .A1(n11549), .A2(n11551), .ZN(n11558) );
  NOR2_X1 U11508 ( .A1(n11562), .A2(n11563), .ZN(n11551) );
  NOR3_X1 U11509 ( .A1(n8982), .A2(n11564), .A3(n8559), .ZN(n11563) );
  NOR2_X1 U11510 ( .A1(n11547), .A2(n11545), .ZN(n11564) );
  INV_X1 U11511 ( .A(n11565), .ZN(n11562) );
  NAND2_X1 U11512 ( .A1(n11545), .A2(n11547), .ZN(n11565) );
  NAND2_X1 U11513 ( .A1(n11566), .A2(n11567), .ZN(n11547) );
  NAND3_X1 U11514 ( .A1(n9792), .A2(n11568), .A3(n11182), .ZN(n11567) );
  INV_X1 U11515 ( .A(n11569), .ZN(n11568) );
  NOR2_X1 U11516 ( .A1(n11543), .A2(n11541), .ZN(n11569) );
  NAND2_X1 U11517 ( .A1(n11541), .A2(n11543), .ZN(n11566) );
  NAND2_X1 U11518 ( .A1(n11570), .A2(n11571), .ZN(n11543) );
  INV_X1 U11519 ( .A(n11572), .ZN(n11571) );
  NOR3_X1 U11520 ( .A1(n8528), .A2(n11573), .A3(n8559), .ZN(n11572) );
  NOR2_X1 U11521 ( .A1(n11539), .A2(n11537), .ZN(n11573) );
  NAND2_X1 U11522 ( .A1(n11537), .A2(n11539), .ZN(n11570) );
  NAND2_X1 U11523 ( .A1(n11574), .A2(n11575), .ZN(n11539) );
  NAND3_X1 U11524 ( .A1(n10307), .A2(n11576), .A3(n11182), .ZN(n11575) );
  INV_X1 U11525 ( .A(n11577), .ZN(n11576) );
  NOR2_X1 U11526 ( .A1(n11535), .A2(n11534), .ZN(n11577) );
  NAND2_X1 U11527 ( .A1(n11534), .A2(n11535), .ZN(n11574) );
  NAND2_X1 U11528 ( .A1(n11578), .A2(n11579), .ZN(n11535) );
  INV_X1 U11529 ( .A(n11580), .ZN(n11579) );
  NOR3_X1 U11530 ( .A1(n9000), .A2(n11581), .A3(n8559), .ZN(n11580) );
  NOR2_X1 U11531 ( .A1(n11531), .A2(n11529), .ZN(n11581) );
  NAND2_X1 U11532 ( .A1(n11529), .A2(n11531), .ZN(n11578) );
  NAND2_X1 U11533 ( .A1(n11582), .A2(n11583), .ZN(n11531) );
  NAND3_X1 U11534 ( .A1(n8543), .A2(n11584), .A3(n11182), .ZN(n11583) );
  INV_X1 U11535 ( .A(n11585), .ZN(n11584) );
  NOR2_X1 U11536 ( .A1(n11527), .A2(n11525), .ZN(n11585) );
  NAND2_X1 U11537 ( .A1(n11525), .A2(n11527), .ZN(n11582) );
  NAND2_X1 U11538 ( .A1(n11523), .A2(n11586), .ZN(n11527) );
  NAND2_X1 U11539 ( .A1(n11522), .A2(n11524), .ZN(n11586) );
  NAND2_X1 U11540 ( .A1(n11587), .A2(n11588), .ZN(n11524) );
  NAND2_X1 U11541 ( .A1(n11182), .A2(n9295), .ZN(n11588) );
  XNOR2_X1 U11542 ( .A(n11589), .B(n11590), .ZN(n11522) );
  XOR2_X1 U11543 ( .A(n11591), .B(n11592), .Z(n11590) );
  NAND2_X1 U11544 ( .A1(n9295), .A2(n11593), .ZN(n11523) );
  INV_X1 U11545 ( .A(n11587), .ZN(n11593) );
  NOR2_X1 U11546 ( .A1(n11594), .A2(n11595), .ZN(n11587) );
  INV_X1 U11547 ( .A(n11596), .ZN(n11595) );
  NAND2_X1 U11548 ( .A1(n11520), .A2(n11597), .ZN(n11596) );
  NAND2_X1 U11549 ( .A1(n11519), .A2(n11518), .ZN(n11597) );
  NOR2_X1 U11550 ( .A1(n8559), .A2(n8594), .ZN(n11520) );
  NOR2_X1 U11551 ( .A1(n11518), .A2(n11519), .ZN(n11594) );
  NOR2_X1 U11552 ( .A1(n11598), .A2(n11599), .ZN(n11519) );
  INV_X1 U11553 ( .A(n11600), .ZN(n11599) );
  NAND2_X1 U11554 ( .A1(n11516), .A2(n11601), .ZN(n11600) );
  NAND2_X1 U11555 ( .A1(n11602), .A2(n11513), .ZN(n11601) );
  NOR2_X1 U11556 ( .A1(n8559), .A2(n8556), .ZN(n11516) );
  NOR2_X1 U11557 ( .A1(n11513), .A2(n11602), .ZN(n11598) );
  INV_X1 U11558 ( .A(n11515), .ZN(n11602) );
  NAND2_X1 U11559 ( .A1(n11603), .A2(n11604), .ZN(n11515) );
  NAND2_X1 U11560 ( .A1(n11512), .A2(n11605), .ZN(n11604) );
  INV_X1 U11561 ( .A(n11606), .ZN(n11605) );
  NOR2_X1 U11562 ( .A1(n11511), .A2(n11510), .ZN(n11606) );
  NOR2_X1 U11563 ( .A1(n8559), .A2(n8572), .ZN(n11512) );
  NAND2_X1 U11564 ( .A1(n11510), .A2(n11511), .ZN(n11603) );
  NAND2_X1 U11565 ( .A1(n11607), .A2(n11608), .ZN(n11511) );
  NAND2_X1 U11566 ( .A1(n11508), .A2(n11609), .ZN(n11608) );
  INV_X1 U11567 ( .A(n11610), .ZN(n11609) );
  NOR2_X1 U11568 ( .A1(n11507), .A2(n11505), .ZN(n11610) );
  NOR2_X1 U11569 ( .A1(n8559), .A2(n8582), .ZN(n11508) );
  NAND2_X1 U11570 ( .A1(n11505), .A2(n11507), .ZN(n11607) );
  NAND2_X1 U11571 ( .A1(n11611), .A2(n11612), .ZN(n11507) );
  NAND2_X1 U11572 ( .A1(n11504), .A2(n11613), .ZN(n11612) );
  INV_X1 U11573 ( .A(n11614), .ZN(n11613) );
  NOR2_X1 U11574 ( .A1(n11503), .A2(n11502), .ZN(n11614) );
  NOR2_X1 U11575 ( .A1(n8559), .A2(n8591), .ZN(n11504) );
  NAND2_X1 U11576 ( .A1(n11502), .A2(n11503), .ZN(n11611) );
  NAND2_X1 U11577 ( .A1(n11615), .A2(n11616), .ZN(n11503) );
  NAND2_X1 U11578 ( .A1(n11500), .A2(n11617), .ZN(n11616) );
  NAND2_X1 U11579 ( .A1(n11499), .A2(n11497), .ZN(n11617) );
  NOR2_X1 U11580 ( .A1(n8559), .A2(n8562), .ZN(n11500) );
  INV_X1 U11581 ( .A(n11618), .ZN(n11615) );
  NOR2_X1 U11582 ( .A1(n11497), .A2(n11499), .ZN(n11618) );
  NOR2_X1 U11583 ( .A1(n11619), .A2(n11620), .ZN(n11499) );
  INV_X1 U11584 ( .A(n11621), .ZN(n11620) );
  NAND2_X1 U11585 ( .A1(n11496), .A2(n11622), .ZN(n11621) );
  NAND2_X1 U11586 ( .A1(n11495), .A2(n11494), .ZN(n11622) );
  NOR2_X1 U11587 ( .A1(n8559), .A2(n8545), .ZN(n11496) );
  NOR2_X1 U11588 ( .A1(n11494), .A2(n11495), .ZN(n11619) );
  INV_X1 U11589 ( .A(n11623), .ZN(n11495) );
  NAND2_X1 U11590 ( .A1(n11624), .A2(n11625), .ZN(n11623) );
  NAND2_X1 U11591 ( .A1(n11491), .A2(n11626), .ZN(n11625) );
  INV_X1 U11592 ( .A(n11627), .ZN(n11626) );
  NOR2_X1 U11593 ( .A1(n11492), .A2(n11490), .ZN(n11627) );
  NOR2_X1 U11594 ( .A1(n8559), .A2(n8569), .ZN(n11491) );
  NAND2_X1 U11595 ( .A1(n11490), .A2(n11492), .ZN(n11624) );
  NAND2_X1 U11596 ( .A1(n11628), .A2(n11629), .ZN(n11492) );
  NAND2_X1 U11597 ( .A1(n11488), .A2(n11630), .ZN(n11629) );
  INV_X1 U11598 ( .A(n11631), .ZN(n11630) );
  NOR2_X1 U11599 ( .A1(n11487), .A2(n11486), .ZN(n11631) );
  NOR2_X1 U11600 ( .A1(n8559), .A2(n8593), .ZN(n11488) );
  NAND2_X1 U11601 ( .A1(n11486), .A2(n11487), .ZN(n11628) );
  NAND2_X1 U11602 ( .A1(n11632), .A2(n11633), .ZN(n11487) );
  NAND2_X1 U11603 ( .A1(n11484), .A2(n11634), .ZN(n11633) );
  NAND2_X1 U11604 ( .A1(n11483), .A2(n11481), .ZN(n11634) );
  NOR2_X1 U11605 ( .A1(n8559), .A2(n8583), .ZN(n11484) );
  INV_X1 U11606 ( .A(n11635), .ZN(n11632) );
  NOR2_X1 U11607 ( .A1(n11481), .A2(n11483), .ZN(n11635) );
  NOR2_X1 U11608 ( .A1(n11636), .A2(n11637), .ZN(n11483) );
  INV_X1 U11609 ( .A(n11638), .ZN(n11637) );
  NAND2_X1 U11610 ( .A1(n11480), .A2(n11639), .ZN(n11638) );
  NAND2_X1 U11611 ( .A1(n11479), .A2(n11478), .ZN(n11639) );
  NOR2_X1 U11612 ( .A1(n8559), .A2(n8580), .ZN(n11480) );
  NOR2_X1 U11613 ( .A1(n11478), .A2(n11479), .ZN(n11636) );
  NOR2_X1 U11614 ( .A1(n11640), .A2(n11641), .ZN(n11479) );
  INV_X1 U11615 ( .A(n11642), .ZN(n11641) );
  NAND2_X1 U11616 ( .A1(n11476), .A2(n11643), .ZN(n11642) );
  NAND2_X1 U11617 ( .A1(n11475), .A2(n11474), .ZN(n11643) );
  NOR2_X1 U11618 ( .A1(n8559), .A2(n8588), .ZN(n11476) );
  NOR2_X1 U11619 ( .A1(n11474), .A2(n11475), .ZN(n11640) );
  NOR2_X1 U11620 ( .A1(n11644), .A2(n11645), .ZN(n11475) );
  INV_X1 U11621 ( .A(n11646), .ZN(n11645) );
  NAND2_X1 U11622 ( .A1(n11471), .A2(n11647), .ZN(n11646) );
  NAND2_X1 U11623 ( .A1(n11472), .A2(n11470), .ZN(n11647) );
  NOR2_X1 U11624 ( .A1(n11181), .A2(n8551), .ZN(n11471) );
  NOR2_X1 U11625 ( .A1(n11470), .A2(n11472), .ZN(n11644) );
  NOR2_X1 U11626 ( .A1(n11648), .A2(n11649), .ZN(n11472) );
  INV_X1 U11627 ( .A(n11650), .ZN(n11649) );
  NAND2_X1 U11628 ( .A1(n11468), .A2(n11651), .ZN(n11650) );
  NAND2_X1 U11629 ( .A1(n11467), .A2(n11466), .ZN(n11651) );
  NOR2_X1 U11630 ( .A1(n11181), .A2(n8563), .ZN(n11468) );
  NOR2_X1 U11631 ( .A1(n11466), .A2(n11467), .ZN(n11648) );
  NOR2_X1 U11632 ( .A1(n11652), .A2(n11653), .ZN(n11467) );
  INV_X1 U11633 ( .A(n11654), .ZN(n11653) );
  NAND2_X1 U11634 ( .A1(n11463), .A2(n11655), .ZN(n11654) );
  NAND2_X1 U11635 ( .A1(n11464), .A2(n11462), .ZN(n11655) );
  NOR2_X1 U11636 ( .A1(n11181), .A2(n8548), .ZN(n11463) );
  NOR2_X1 U11637 ( .A1(n11462), .A2(n11464), .ZN(n11652) );
  NOR2_X1 U11638 ( .A1(n11656), .A2(n11657), .ZN(n11464) );
  INV_X1 U11639 ( .A(n11658), .ZN(n11657) );
  NAND2_X1 U11640 ( .A1(n11460), .A2(n11659), .ZN(n11658) );
  NAND2_X1 U11641 ( .A1(n11459), .A2(n11458), .ZN(n11659) );
  NOR2_X1 U11642 ( .A1(n11181), .A2(n8584), .ZN(n11460) );
  NOR2_X1 U11643 ( .A1(n11458), .A2(n11459), .ZN(n11656) );
  NOR2_X1 U11644 ( .A1(n11660), .A2(n11661), .ZN(n11459) );
  INV_X1 U11645 ( .A(n11662), .ZN(n11661) );
  NAND2_X1 U11646 ( .A1(n11455), .A2(n11663), .ZN(n11662) );
  NAND2_X1 U11647 ( .A1(n11456), .A2(n11454), .ZN(n11663) );
  NOR2_X1 U11648 ( .A1(n11181), .A2(n8535), .ZN(n11455) );
  NOR2_X1 U11649 ( .A1(n11454), .A2(n11456), .ZN(n11660) );
  NOR2_X1 U11650 ( .A1(n11664), .A2(n11665), .ZN(n11456) );
  INV_X1 U11651 ( .A(n11666), .ZN(n11665) );
  NAND2_X1 U11652 ( .A1(n11451), .A2(n11667), .ZN(n11666) );
  NAND2_X1 U11653 ( .A1(n11452), .A2(n11450), .ZN(n11667) );
  NOR2_X1 U11654 ( .A1(n11181), .A2(n8568), .ZN(n11451) );
  NOR2_X1 U11655 ( .A1(n11450), .A2(n11452), .ZN(n11664) );
  NOR2_X1 U11656 ( .A1(n11668), .A2(n11669), .ZN(n11452) );
  INV_X1 U11657 ( .A(n11670), .ZN(n11669) );
  NAND2_X1 U11658 ( .A1(n11447), .A2(n11671), .ZN(n11670) );
  NAND2_X1 U11659 ( .A1(n11448), .A2(n11446), .ZN(n11671) );
  NOR2_X1 U11660 ( .A1(n11181), .A2(n8574), .ZN(n11447) );
  NOR2_X1 U11661 ( .A1(n11446), .A2(n11448), .ZN(n11668) );
  NOR2_X1 U11662 ( .A1(n11672), .A2(n11673), .ZN(n11448) );
  INV_X1 U11663 ( .A(n11674), .ZN(n11673) );
  NAND2_X1 U11664 ( .A1(n11443), .A2(n11675), .ZN(n11674) );
  NAND2_X1 U11665 ( .A1(n11444), .A2(n11442), .ZN(n11675) );
  NOR2_X1 U11666 ( .A1(n11181), .A2(n8565), .ZN(n11443) );
  NOR2_X1 U11667 ( .A1(n11442), .A2(n11444), .ZN(n11672) );
  NOR2_X1 U11668 ( .A1(n11676), .A2(n11677), .ZN(n11444) );
  INV_X1 U11669 ( .A(n11678), .ZN(n11677) );
  NAND2_X1 U11670 ( .A1(n11437), .A2(n11679), .ZN(n11678) );
  NAND2_X1 U11671 ( .A1(n11440), .A2(n11439), .ZN(n11679) );
  NOR2_X1 U11672 ( .A1(n11181), .A2(n8567), .ZN(n11437) );
  NOR2_X1 U11673 ( .A1(n11439), .A2(n11440), .ZN(n11676) );
  INV_X1 U11674 ( .A(n11680), .ZN(n11440) );
  NAND2_X1 U11675 ( .A1(n11681), .A2(n11682), .ZN(n11680) );
  NAND2_X1 U11676 ( .A1(n11432), .A2(n11683), .ZN(n11682) );
  NAND2_X1 U11677 ( .A1(n8624), .A2(n11684), .ZN(n11683) );
  NAND2_X1 U11678 ( .A1(n8558), .A2(n8585), .ZN(n11684) );
  NAND2_X1 U11679 ( .A1(n11686), .A2(n11687), .ZN(n11681) );
  NAND2_X1 U11680 ( .A1(n8630), .A2(n11688), .ZN(n11687) );
  NAND2_X1 U11681 ( .A1(n8539), .A2(n8581), .ZN(n11688) );
  NAND3_X1 U11682 ( .A1(n11432), .A2(n8537), .A3(n11182), .ZN(n11439) );
  INV_X1 U11683 ( .A(n11181), .ZN(n11182) );
  XNOR2_X1 U11684 ( .A(n11689), .B(n11690), .ZN(n11181) );
  XOR2_X1 U11685 ( .A(d_21_), .B(c_21_), .Z(n11690) );
  XOR2_X1 U11686 ( .A(n11691), .B(n11692), .Z(n11442) );
  XNOR2_X1 U11687 ( .A(n11693), .B(n11694), .ZN(n11692) );
  XOR2_X1 U11688 ( .A(n11695), .B(n11696), .Z(n11446) );
  XNOR2_X1 U11689 ( .A(n11697), .B(n11698), .ZN(n11695) );
  XOR2_X1 U11690 ( .A(n11699), .B(n11700), .Z(n11450) );
  XNOR2_X1 U11691 ( .A(n11701), .B(n11702), .ZN(n11699) );
  XOR2_X1 U11692 ( .A(n11703), .B(n11704), .Z(n11454) );
  XNOR2_X1 U11693 ( .A(n11705), .B(n11706), .ZN(n11703) );
  XOR2_X1 U11694 ( .A(n11707), .B(n11708), .Z(n11458) );
  XNOR2_X1 U11695 ( .A(n11709), .B(n11710), .ZN(n11707) );
  NOR2_X1 U11696 ( .A1(n8535), .A2(n8581), .ZN(n11710) );
  XOR2_X1 U11697 ( .A(n11711), .B(n11712), .Z(n11462) );
  XNOR2_X1 U11698 ( .A(n11713), .B(n11714), .ZN(n11711) );
  NOR2_X1 U11699 ( .A1(n8584), .A2(n8581), .ZN(n11714) );
  XOR2_X1 U11700 ( .A(n11715), .B(n11716), .Z(n11466) );
  XNOR2_X1 U11701 ( .A(n11717), .B(n11718), .ZN(n11715) );
  NOR2_X1 U11702 ( .A1(n8548), .A2(n8581), .ZN(n11718) );
  XOR2_X1 U11703 ( .A(n11719), .B(n11720), .Z(n11470) );
  XNOR2_X1 U11704 ( .A(n11721), .B(n11722), .ZN(n11719) );
  NOR2_X1 U11705 ( .A1(n8563), .A2(n8581), .ZN(n11722) );
  XNOR2_X1 U11706 ( .A(n11723), .B(n11724), .ZN(n11474) );
  XNOR2_X1 U11707 ( .A(n11725), .B(n11726), .ZN(n11724) );
  NAND2_X1 U11708 ( .A1(n11432), .A2(n8515), .ZN(n11726) );
  XOR2_X1 U11709 ( .A(n11727), .B(n11728), .Z(n11478) );
  XNOR2_X1 U11710 ( .A(n11729), .B(n11730), .ZN(n11727) );
  NOR2_X1 U11711 ( .A1(n8588), .A2(n8581), .ZN(n11730) );
  XOR2_X1 U11712 ( .A(n11731), .B(n11732), .Z(n11481) );
  XNOR2_X1 U11713 ( .A(n11733), .B(n11734), .ZN(n11731) );
  NOR2_X1 U11714 ( .A1(n8580), .A2(n8581), .ZN(n11734) );
  XNOR2_X1 U11715 ( .A(n11735), .B(n11736), .ZN(n11486) );
  XNOR2_X1 U11716 ( .A(n11737), .B(n11738), .ZN(n11735) );
  NOR2_X1 U11717 ( .A1(n8583), .A2(n8581), .ZN(n11738) );
  XNOR2_X1 U11718 ( .A(n11739), .B(n11740), .ZN(n11490) );
  XNOR2_X1 U11719 ( .A(n11741), .B(n11742), .ZN(n11739) );
  NOR2_X1 U11720 ( .A1(n8593), .A2(n8581), .ZN(n11742) );
  XOR2_X1 U11721 ( .A(n11743), .B(n11744), .Z(n11494) );
  XNOR2_X1 U11722 ( .A(n11745), .B(n11746), .ZN(n11743) );
  NOR2_X1 U11723 ( .A1(n9050), .A2(n8581), .ZN(n11746) );
  XOR2_X1 U11724 ( .A(n11747), .B(n11748), .Z(n11497) );
  XNOR2_X1 U11725 ( .A(n11749), .B(n11750), .ZN(n11747) );
  NOR2_X1 U11726 ( .A1(n8545), .A2(n8581), .ZN(n11750) );
  XNOR2_X1 U11727 ( .A(n11751), .B(n11752), .ZN(n11502) );
  XNOR2_X1 U11728 ( .A(n11753), .B(n11754), .ZN(n11751) );
  NOR2_X1 U11729 ( .A1(n9041), .A2(n8581), .ZN(n11754) );
  XNOR2_X1 U11730 ( .A(n11755), .B(n11756), .ZN(n11505) );
  XNOR2_X1 U11731 ( .A(n11757), .B(n11758), .ZN(n11755) );
  NOR2_X1 U11732 ( .A1(n8591), .A2(n8581), .ZN(n11758) );
  XNOR2_X1 U11733 ( .A(n11759), .B(n11760), .ZN(n11510) );
  XNOR2_X1 U11734 ( .A(n11761), .B(n11762), .ZN(n11759) );
  NOR2_X1 U11735 ( .A1(n9031), .A2(n8581), .ZN(n11762) );
  XOR2_X1 U11736 ( .A(n11763), .B(n11764), .Z(n11513) );
  XNOR2_X1 U11737 ( .A(n11765), .B(n11766), .ZN(n11763) );
  NOR2_X1 U11738 ( .A1(n8572), .A2(n8581), .ZN(n11766) );
  XNOR2_X1 U11739 ( .A(n11767), .B(n11768), .ZN(n11518) );
  XNOR2_X1 U11740 ( .A(n11769), .B(n11770), .ZN(n11768) );
  NAND2_X1 U11741 ( .A1(n11432), .A2(n9304), .ZN(n11770) );
  XOR2_X1 U11742 ( .A(n11771), .B(n11772), .Z(n11525) );
  XNOR2_X1 U11743 ( .A(n11773), .B(n11774), .ZN(n11771) );
  XOR2_X1 U11744 ( .A(n11775), .B(n11776), .Z(n11529) );
  XOR2_X1 U11745 ( .A(n11777), .B(n11778), .Z(n11775) );
  XNOR2_X1 U11746 ( .A(n11779), .B(n11780), .ZN(n11534) );
  XOR2_X1 U11747 ( .A(n11781), .B(n11782), .Z(n11780) );
  XNOR2_X1 U11748 ( .A(n11783), .B(n11784), .ZN(n11537) );
  XNOR2_X1 U11749 ( .A(n11785), .B(n11786), .ZN(n11783) );
  XNOR2_X1 U11750 ( .A(n11787), .B(n11788), .ZN(n11541) );
  XNOR2_X1 U11751 ( .A(n11789), .B(n11790), .ZN(n11787) );
  XOR2_X1 U11752 ( .A(n11791), .B(n11792), .Z(n11545) );
  XNOR2_X1 U11753 ( .A(n11793), .B(n11794), .ZN(n11791) );
  XOR2_X1 U11754 ( .A(n11795), .B(n11796), .Z(n11549) );
  XOR2_X1 U11755 ( .A(n11797), .B(n11798), .Z(n11796) );
  XOR2_X1 U11756 ( .A(n11799), .B(n11800), .Z(n11302) );
  XNOR2_X1 U11757 ( .A(n11801), .B(n11802), .ZN(n11799) );
  XNOR2_X1 U11758 ( .A(n11803), .B(n11804), .ZN(n8928) );
  XNOR2_X1 U11759 ( .A(n11805), .B(n11806), .ZN(n11803) );
  NOR2_X1 U11760 ( .A1(n8972), .A2(n8581), .ZN(n11806) );
  NAND4_X1 U11761 ( .A1(n8923), .A2(n8922), .A3(n8924), .A4(n8916), .ZN(n8833)
         );
  INV_X1 U11762 ( .A(n11807), .ZN(n8916) );
  NAND2_X1 U11763 ( .A1(n11808), .A2(n11809), .ZN(n8924) );
  NAND3_X1 U11764 ( .A1(n8592), .A2(n11810), .A3(n11432), .ZN(n11809) );
  NAND2_X1 U11765 ( .A1(n11805), .A2(n11804), .ZN(n11810) );
  INV_X1 U11766 ( .A(n11811), .ZN(n11808) );
  NOR2_X1 U11767 ( .A1(n11804), .A2(n11805), .ZN(n11811) );
  NOR2_X1 U11768 ( .A1(n11812), .A2(n11813), .ZN(n11805) );
  INV_X1 U11769 ( .A(n11814), .ZN(n11813) );
  NAND2_X1 U11770 ( .A1(n11802), .A2(n11815), .ZN(n11814) );
  NAND2_X1 U11771 ( .A1(n11801), .A2(n11800), .ZN(n11815) );
  NOR2_X1 U11772 ( .A1(n8581), .A2(n8589), .ZN(n11802) );
  NOR2_X1 U11773 ( .A1(n11800), .A2(n11801), .ZN(n11812) );
  NOR2_X1 U11774 ( .A1(n11816), .A2(n11817), .ZN(n11801) );
  NOR2_X1 U11775 ( .A1(n11798), .A2(n11818), .ZN(n11817) );
  NOR2_X1 U11776 ( .A1(n11797), .A2(n11795), .ZN(n11818) );
  NAND2_X1 U11777 ( .A1(n11432), .A2(n9268), .ZN(n11798) );
  INV_X1 U11778 ( .A(n11819), .ZN(n11816) );
  NAND2_X1 U11779 ( .A1(n11795), .A2(n11797), .ZN(n11819) );
  NAND2_X1 U11780 ( .A1(n11820), .A2(n11821), .ZN(n11797) );
  NAND2_X1 U11781 ( .A1(n11794), .A2(n11822), .ZN(n11821) );
  NAND2_X1 U11782 ( .A1(n11793), .A2(n11823), .ZN(n11822) );
  INV_X1 U11783 ( .A(n11792), .ZN(n11823) );
  NOR2_X1 U11784 ( .A1(n8581), .A2(n8527), .ZN(n11794) );
  NAND2_X1 U11785 ( .A1(n11792), .A2(n11824), .ZN(n11820) );
  INV_X1 U11786 ( .A(n11793), .ZN(n11824) );
  NOR2_X1 U11787 ( .A1(n11825), .A2(n11826), .ZN(n11793) );
  INV_X1 U11788 ( .A(n11827), .ZN(n11826) );
  NAND2_X1 U11789 ( .A1(n11790), .A2(n11828), .ZN(n11827) );
  NAND2_X1 U11790 ( .A1(n11789), .A2(n11788), .ZN(n11828) );
  NOR2_X1 U11791 ( .A1(n11431), .A2(n8528), .ZN(n11790) );
  NOR2_X1 U11792 ( .A1(n11788), .A2(n11789), .ZN(n11825) );
  NOR2_X1 U11793 ( .A1(n11829), .A2(n11830), .ZN(n11789) );
  INV_X1 U11794 ( .A(n11831), .ZN(n11830) );
  NAND2_X1 U11795 ( .A1(n11786), .A2(n11832), .ZN(n11831) );
  NAND2_X1 U11796 ( .A1(n11785), .A2(n11784), .ZN(n11832) );
  NOR2_X1 U11797 ( .A1(n11431), .A2(n8564), .ZN(n11786) );
  NOR2_X1 U11798 ( .A1(n11784), .A2(n11785), .ZN(n11829) );
  NOR2_X1 U11799 ( .A1(n11833), .A2(n11834), .ZN(n11785) );
  NOR2_X1 U11800 ( .A1(n11782), .A2(n11835), .ZN(n11834) );
  NOR2_X1 U11801 ( .A1(n11781), .A2(n11779), .ZN(n11835) );
  NAND2_X1 U11802 ( .A1(n11432), .A2(n9286), .ZN(n11782) );
  INV_X1 U11803 ( .A(n11836), .ZN(n11833) );
  NAND2_X1 U11804 ( .A1(n11779), .A2(n11781), .ZN(n11836) );
  NAND2_X1 U11805 ( .A1(n11837), .A2(n11838), .ZN(n11781) );
  NAND2_X1 U11806 ( .A1(n11778), .A2(n11839), .ZN(n11838) );
  INV_X1 U11807 ( .A(n11840), .ZN(n11839) );
  NOR2_X1 U11808 ( .A1(n11777), .A2(n11776), .ZN(n11840) );
  NOR2_X1 U11809 ( .A1(n11431), .A2(n8544), .ZN(n11778) );
  NAND2_X1 U11810 ( .A1(n11776), .A2(n11777), .ZN(n11837) );
  NAND2_X1 U11811 ( .A1(n11841), .A2(n11842), .ZN(n11777) );
  NAND2_X1 U11812 ( .A1(n11774), .A2(n11843), .ZN(n11842) );
  NAND2_X1 U11813 ( .A1(n11773), .A2(n11844), .ZN(n11843) );
  INV_X1 U11814 ( .A(n11772), .ZN(n11844) );
  NOR2_X1 U11815 ( .A1(n11431), .A2(n8560), .ZN(n11774) );
  NAND2_X1 U11816 ( .A1(n11772), .A2(n11845), .ZN(n11841) );
  INV_X1 U11817 ( .A(n11773), .ZN(n11845) );
  NOR2_X1 U11818 ( .A1(n11846), .A2(n11847), .ZN(n11773) );
  NOR2_X1 U11819 ( .A1(n11592), .A2(n11848), .ZN(n11847) );
  NOR2_X1 U11820 ( .A1(n11591), .A2(n11589), .ZN(n11848) );
  NAND2_X1 U11821 ( .A1(n11432), .A2(n10846), .ZN(n11592) );
  INV_X1 U11822 ( .A(n11849), .ZN(n11846) );
  NAND2_X1 U11823 ( .A1(n11589), .A2(n11591), .ZN(n11849) );
  NAND2_X1 U11824 ( .A1(n11850), .A2(n11851), .ZN(n11591) );
  NAND3_X1 U11825 ( .A1(n9304), .A2(n11852), .A3(n11432), .ZN(n11851) );
  NAND2_X1 U11826 ( .A1(n11769), .A2(n11767), .ZN(n11852) );
  INV_X1 U11827 ( .A(n11853), .ZN(n11850) );
  NOR2_X1 U11828 ( .A1(n11767), .A2(n11769), .ZN(n11853) );
  NOR2_X1 U11829 ( .A1(n11854), .A2(n11855), .ZN(n11769) );
  INV_X1 U11830 ( .A(n11856), .ZN(n11855) );
  NAND3_X1 U11831 ( .A1(n9209), .A2(n11857), .A3(n11432), .ZN(n11856) );
  NAND2_X1 U11832 ( .A1(n11765), .A2(n11764), .ZN(n11857) );
  NOR2_X1 U11833 ( .A1(n11764), .A2(n11765), .ZN(n11854) );
  NOR2_X1 U11834 ( .A1(n11858), .A2(n11859), .ZN(n11765) );
  INV_X1 U11835 ( .A(n11860), .ZN(n11859) );
  NAND3_X1 U11836 ( .A1(n9313), .A2(n11861), .A3(n11432), .ZN(n11860) );
  NAND2_X1 U11837 ( .A1(n11761), .A2(n11760), .ZN(n11861) );
  NOR2_X1 U11838 ( .A1(n11760), .A2(n11761), .ZN(n11858) );
  NOR2_X1 U11839 ( .A1(n11862), .A2(n11863), .ZN(n11761) );
  NOR3_X1 U11840 ( .A1(n9036), .A2(n11864), .A3(n8581), .ZN(n11863) );
  INV_X1 U11841 ( .A(n11865), .ZN(n11864) );
  NAND2_X1 U11842 ( .A1(n11757), .A2(n11756), .ZN(n11865) );
  NOR2_X1 U11843 ( .A1(n11756), .A2(n11757), .ZN(n11862) );
  NOR2_X1 U11844 ( .A1(n11866), .A2(n11867), .ZN(n11757) );
  INV_X1 U11845 ( .A(n11868), .ZN(n11867) );
  NAND3_X1 U11846 ( .A1(n9322), .A2(n11869), .A3(n11432), .ZN(n11868) );
  NAND2_X1 U11847 ( .A1(n11753), .A2(n11752), .ZN(n11869) );
  NOR2_X1 U11848 ( .A1(n11752), .A2(n11753), .ZN(n11866) );
  NOR2_X1 U11849 ( .A1(n11870), .A2(n11871), .ZN(n11753) );
  NOR3_X1 U11850 ( .A1(n8545), .A2(n11872), .A3(n8581), .ZN(n11871) );
  INV_X1 U11851 ( .A(n11873), .ZN(n11872) );
  NAND2_X1 U11852 ( .A1(n11749), .A2(n11748), .ZN(n11873) );
  NOR2_X1 U11853 ( .A1(n11748), .A2(n11749), .ZN(n11870) );
  NOR2_X1 U11854 ( .A1(n11874), .A2(n11875), .ZN(n11749) );
  INV_X1 U11855 ( .A(n11876), .ZN(n11875) );
  NAND3_X1 U11856 ( .A1(n9331), .A2(n11877), .A3(n11432), .ZN(n11876) );
  NAND2_X1 U11857 ( .A1(n11745), .A2(n11744), .ZN(n11877) );
  NOR2_X1 U11858 ( .A1(n11744), .A2(n11745), .ZN(n11874) );
  NOR2_X1 U11859 ( .A1(n11878), .A2(n11879), .ZN(n11745) );
  NOR3_X1 U11860 ( .A1(n9056), .A2(n11880), .A3(n8581), .ZN(n11879) );
  INV_X1 U11861 ( .A(n11881), .ZN(n11880) );
  NAND2_X1 U11862 ( .A1(n11741), .A2(n11740), .ZN(n11881) );
  NOR2_X1 U11863 ( .A1(n11740), .A2(n11741), .ZN(n11878) );
  NOR2_X1 U11864 ( .A1(n11882), .A2(n11883), .ZN(n11741) );
  INV_X1 U11865 ( .A(n11884), .ZN(n11883) );
  NAND3_X1 U11866 ( .A1(n9340), .A2(n11885), .A3(n11432), .ZN(n11884) );
  NAND2_X1 U11867 ( .A1(n11737), .A2(n11736), .ZN(n11885) );
  NOR2_X1 U11868 ( .A1(n11736), .A2(n11737), .ZN(n11882) );
  NOR2_X1 U11869 ( .A1(n11886), .A2(n11887), .ZN(n11737) );
  NOR3_X1 U11870 ( .A1(n9066), .A2(n11888), .A3(n8581), .ZN(n11887) );
  INV_X1 U11871 ( .A(n11889), .ZN(n11888) );
  NAND2_X1 U11872 ( .A1(n11733), .A2(n11732), .ZN(n11889) );
  NOR2_X1 U11873 ( .A1(n11732), .A2(n11733), .ZN(n11886) );
  NOR2_X1 U11874 ( .A1(n11890), .A2(n11891), .ZN(n11733) );
  INV_X1 U11875 ( .A(n11892), .ZN(n11891) );
  NAND3_X1 U11876 ( .A1(n9080), .A2(n11893), .A3(n11432), .ZN(n11892) );
  NAND2_X1 U11877 ( .A1(n11729), .A2(n11728), .ZN(n11893) );
  NOR2_X1 U11878 ( .A1(n11728), .A2(n11729), .ZN(n11890) );
  NOR2_X1 U11879 ( .A1(n11894), .A2(n11895), .ZN(n11729) );
  NOR3_X1 U11880 ( .A1(n8551), .A2(n11896), .A3(n8581), .ZN(n11895) );
  INV_X1 U11881 ( .A(n11897), .ZN(n11896) );
  NAND2_X1 U11882 ( .A1(n11725), .A2(n11723), .ZN(n11897) );
  NOR2_X1 U11883 ( .A1(n11723), .A2(n11725), .ZN(n11894) );
  NOR2_X1 U11884 ( .A1(n11898), .A2(n11899), .ZN(n11725) );
  INV_X1 U11885 ( .A(n11900), .ZN(n11899) );
  NAND3_X1 U11886 ( .A1(n9098), .A2(n11901), .A3(n11432), .ZN(n11900) );
  NAND2_X1 U11887 ( .A1(n11721), .A2(n11720), .ZN(n11901) );
  NOR2_X1 U11888 ( .A1(n11720), .A2(n11721), .ZN(n11898) );
  NOR2_X1 U11889 ( .A1(n11902), .A2(n11903), .ZN(n11721) );
  NOR3_X1 U11890 ( .A1(n8548), .A2(n11904), .A3(n8581), .ZN(n11903) );
  INV_X1 U11891 ( .A(n11905), .ZN(n11904) );
  NAND2_X1 U11892 ( .A1(n11717), .A2(n11716), .ZN(n11905) );
  NOR2_X1 U11893 ( .A1(n11716), .A2(n11717), .ZN(n11902) );
  NOR2_X1 U11894 ( .A1(n11906), .A2(n11907), .ZN(n11717) );
  INV_X1 U11895 ( .A(n11908), .ZN(n11907) );
  NAND3_X1 U11896 ( .A1(n9112), .A2(n11909), .A3(n11432), .ZN(n11908) );
  NAND2_X1 U11897 ( .A1(n11713), .A2(n11712), .ZN(n11909) );
  NOR2_X1 U11898 ( .A1(n11712), .A2(n11713), .ZN(n11906) );
  NOR2_X1 U11899 ( .A1(n11910), .A2(n11911), .ZN(n11713) );
  INV_X1 U11900 ( .A(n11912), .ZN(n11911) );
  NAND3_X1 U11901 ( .A1(n9121), .A2(n11913), .A3(n11432), .ZN(n11912) );
  NAND2_X1 U11902 ( .A1(n11709), .A2(n11708), .ZN(n11913) );
  NOR2_X1 U11903 ( .A1(n11708), .A2(n11709), .ZN(n11910) );
  NOR2_X1 U11904 ( .A1(n11914), .A2(n11915), .ZN(n11709) );
  INV_X1 U11905 ( .A(n11916), .ZN(n11915) );
  NAND2_X1 U11906 ( .A1(n11705), .A2(n11917), .ZN(n11916) );
  NAND2_X1 U11907 ( .A1(n11706), .A2(n11704), .ZN(n11917) );
  NOR2_X1 U11908 ( .A1(n11431), .A2(n8568), .ZN(n11705) );
  NOR2_X1 U11909 ( .A1(n11704), .A2(n11706), .ZN(n11914) );
  NOR2_X1 U11910 ( .A1(n11918), .A2(n11919), .ZN(n11706) );
  INV_X1 U11911 ( .A(n11920), .ZN(n11919) );
  NAND2_X1 U11912 ( .A1(n11701), .A2(n11921), .ZN(n11920) );
  NAND2_X1 U11913 ( .A1(n11702), .A2(n11700), .ZN(n11921) );
  NOR2_X1 U11914 ( .A1(n11431), .A2(n8574), .ZN(n11701) );
  NOR2_X1 U11915 ( .A1(n11700), .A2(n11702), .ZN(n11918) );
  NOR2_X1 U11916 ( .A1(n11922), .A2(n11923), .ZN(n11702) );
  INV_X1 U11917 ( .A(n11924), .ZN(n11923) );
  NAND2_X1 U11918 ( .A1(n11697), .A2(n11925), .ZN(n11924) );
  NAND2_X1 U11919 ( .A1(n11698), .A2(n11696), .ZN(n11925) );
  NOR2_X1 U11920 ( .A1(n11431), .A2(n8565), .ZN(n11697) );
  NOR2_X1 U11921 ( .A1(n11696), .A2(n11698), .ZN(n11922) );
  NOR2_X1 U11922 ( .A1(n11926), .A2(n11927), .ZN(n11698) );
  INV_X1 U11923 ( .A(n11928), .ZN(n11927) );
  NAND2_X1 U11924 ( .A1(n11691), .A2(n11929), .ZN(n11928) );
  NAND2_X1 U11925 ( .A1(n11694), .A2(n11693), .ZN(n11929) );
  NOR2_X1 U11926 ( .A1(n11431), .A2(n8567), .ZN(n11691) );
  NOR2_X1 U11927 ( .A1(n11693), .A2(n11694), .ZN(n11926) );
  INV_X1 U11928 ( .A(n11930), .ZN(n11694) );
  NAND2_X1 U11929 ( .A1(n11931), .A2(n11932), .ZN(n11930) );
  NAND2_X1 U11930 ( .A1(n11686), .A2(n11933), .ZN(n11932) );
  NAND2_X1 U11931 ( .A1(n8624), .A2(n11934), .ZN(n11933) );
  NAND2_X1 U11932 ( .A1(n8575), .A2(n8585), .ZN(n11934) );
  NAND2_X1 U11933 ( .A1(n11936), .A2(n11937), .ZN(n11931) );
  NAND2_X1 U11934 ( .A1(n8630), .A2(n11938), .ZN(n11937) );
  NAND2_X1 U11935 ( .A1(n8539), .A2(n8558), .ZN(n11938) );
  NAND3_X1 U11936 ( .A1(n11686), .A2(n8537), .A3(n11432), .ZN(n11693) );
  INV_X1 U11937 ( .A(n11431), .ZN(n11432) );
  XNOR2_X1 U11938 ( .A(n11939), .B(n11940), .ZN(n11431) );
  XOR2_X1 U11939 ( .A(d_20_), .B(c_20_), .Z(n11940) );
  XOR2_X1 U11940 ( .A(n11941), .B(n11942), .Z(n11696) );
  XNOR2_X1 U11941 ( .A(n11943), .B(n11944), .ZN(n11942) );
  XOR2_X1 U11942 ( .A(n11945), .B(n11946), .Z(n11700) );
  XNOR2_X1 U11943 ( .A(n11947), .B(n11948), .ZN(n11945) );
  XOR2_X1 U11944 ( .A(n11949), .B(n11950), .Z(n11704) );
  XNOR2_X1 U11945 ( .A(n11951), .B(n11952), .ZN(n11949) );
  XOR2_X1 U11946 ( .A(n11953), .B(n11954), .Z(n11708) );
  XNOR2_X1 U11947 ( .A(n11955), .B(n11956), .ZN(n11953) );
  XOR2_X1 U11948 ( .A(n11957), .B(n11958), .Z(n11712) );
  XNOR2_X1 U11949 ( .A(n11959), .B(n11960), .ZN(n11957) );
  XOR2_X1 U11950 ( .A(n11961), .B(n11962), .Z(n11716) );
  XNOR2_X1 U11951 ( .A(n11963), .B(n11964), .ZN(n11961) );
  XOR2_X1 U11952 ( .A(n11965), .B(n11966), .Z(n11720) );
  XNOR2_X1 U11953 ( .A(n11967), .B(n11968), .ZN(n11965) );
  XOR2_X1 U11954 ( .A(n11969), .B(n11970), .Z(n11723) );
  XNOR2_X1 U11955 ( .A(n11971), .B(n11972), .ZN(n11969) );
  XOR2_X1 U11956 ( .A(n11973), .B(n11974), .Z(n11728) );
  XNOR2_X1 U11957 ( .A(n11975), .B(n11976), .ZN(n11973) );
  XNOR2_X1 U11958 ( .A(n11977), .B(n11978), .ZN(n11732) );
  XOR2_X1 U11959 ( .A(n11979), .B(n11980), .Z(n11978) );
  XNOR2_X1 U11960 ( .A(n11981), .B(n11982), .ZN(n11736) );
  XOR2_X1 U11961 ( .A(n11983), .B(n11984), .Z(n11981) );
  XNOR2_X1 U11962 ( .A(n11985), .B(n11986), .ZN(n11740) );
  XOR2_X1 U11963 ( .A(n11987), .B(n11988), .Z(n11985) );
  XOR2_X1 U11964 ( .A(n11989), .B(n11990), .Z(n11744) );
  XNOR2_X1 U11965 ( .A(n11991), .B(n11992), .ZN(n11989) );
  XNOR2_X1 U11966 ( .A(n11993), .B(n11994), .ZN(n11748) );
  XOR2_X1 U11967 ( .A(n11995), .B(n11996), .Z(n11994) );
  XNOR2_X1 U11968 ( .A(n11997), .B(n11998), .ZN(n11752) );
  XOR2_X1 U11969 ( .A(n11999), .B(n12000), .Z(n11997) );
  XOR2_X1 U11970 ( .A(n12001), .B(n12002), .Z(n11756) );
  XNOR2_X1 U11971 ( .A(n12003), .B(n12004), .ZN(n12002) );
  XNOR2_X1 U11972 ( .A(n12005), .B(n12006), .ZN(n11760) );
  XOR2_X1 U11973 ( .A(n12007), .B(n12008), .Z(n12005) );
  XNOR2_X1 U11974 ( .A(n12009), .B(n12010), .ZN(n11764) );
  XNOR2_X1 U11975 ( .A(n12011), .B(n12012), .ZN(n12010) );
  XOR2_X1 U11976 ( .A(n12013), .B(n12014), .Z(n11767) );
  XNOR2_X1 U11977 ( .A(n12015), .B(n12016), .ZN(n12013) );
  XNOR2_X1 U11978 ( .A(n12017), .B(n12018), .ZN(n11589) );
  NAND2_X1 U11979 ( .A1(n12019), .A2(n12020), .ZN(n12017) );
  XOR2_X1 U11980 ( .A(n12021), .B(n12022), .Z(n11772) );
  XOR2_X1 U11981 ( .A(n12023), .B(n12024), .Z(n12021) );
  NOR2_X1 U11982 ( .A1(n8594), .A2(n8558), .ZN(n12024) );
  XNOR2_X1 U11983 ( .A(n12025), .B(n12026), .ZN(n11776) );
  XOR2_X1 U11984 ( .A(n12027), .B(n12028), .Z(n12026) );
  NAND2_X1 U11985 ( .A1(n11686), .A2(n9295), .ZN(n12028) );
  XOR2_X1 U11986 ( .A(n12029), .B(n12030), .Z(n11779) );
  XOR2_X1 U11987 ( .A(n12031), .B(n12032), .Z(n12029) );
  NOR2_X1 U11988 ( .A1(n8544), .A2(n8558), .ZN(n12032) );
  XOR2_X1 U11989 ( .A(n12033), .B(n12034), .Z(n11784) );
  XOR2_X1 U11990 ( .A(n12035), .B(n12036), .Z(n12034) );
  NAND2_X1 U11991 ( .A1(n11686), .A2(n9286), .ZN(n12036) );
  XOR2_X1 U11992 ( .A(n12037), .B(n12038), .Z(n11788) );
  XOR2_X1 U11993 ( .A(n12039), .B(n12040), .Z(n12038) );
  NAND2_X1 U11994 ( .A1(n11686), .A2(n10307), .ZN(n12040) );
  XNOR2_X1 U11995 ( .A(n12041), .B(n12042), .ZN(n11792) );
  XOR2_X1 U11996 ( .A(n12043), .B(n12044), .Z(n12042) );
  NAND2_X1 U11997 ( .A1(n11686), .A2(n9277), .ZN(n12044) );
  XOR2_X1 U11998 ( .A(n12045), .B(n12046), .Z(n11795) );
  XNOR2_X1 U11999 ( .A(n12047), .B(n12048), .ZN(n12046) );
  NAND2_X1 U12000 ( .A1(n11686), .A2(n9792), .ZN(n12048) );
  XNOR2_X1 U12001 ( .A(n12049), .B(n12050), .ZN(n11800) );
  XNOR2_X1 U12002 ( .A(n12051), .B(n12052), .ZN(n12050) );
  NAND2_X1 U12003 ( .A1(n11686), .A2(n9268), .ZN(n12052) );
  XNOR2_X1 U12004 ( .A(n12053), .B(n12054), .ZN(n11804) );
  XNOR2_X1 U12005 ( .A(n12055), .B(n12056), .ZN(n12054) );
  NAND2_X1 U12006 ( .A1(n11686), .A2(n9263), .ZN(n12056) );
  NAND2_X1 U12007 ( .A1(n12057), .A2(n12058), .ZN(n8922) );
  XNOR2_X1 U12008 ( .A(n12059), .B(n12060), .ZN(n8923) );
  XOR2_X1 U12009 ( .A(n12061), .B(n12062), .Z(n12060) );
  NAND2_X1 U12010 ( .A1(n11686), .A2(n8872), .ZN(n12062) );
  NAND3_X1 U12011 ( .A1(n12063), .A2(n8840), .A3(n11807), .ZN(n8837) );
  NOR2_X1 U12012 ( .A1(n12058), .A2(n12057), .ZN(n11807) );
  NOR2_X1 U12013 ( .A1(n12064), .A2(n12065), .ZN(n12057) );
  NOR3_X1 U12014 ( .A1(n8972), .A2(n12066), .A3(n8558), .ZN(n12065) );
  NOR2_X1 U12015 ( .A1(n12061), .A2(n12059), .ZN(n12066) );
  INV_X1 U12016 ( .A(n12067), .ZN(n12064) );
  NAND2_X1 U12017 ( .A1(n12059), .A2(n12061), .ZN(n12067) );
  NAND2_X1 U12018 ( .A1(n12068), .A2(n12069), .ZN(n12061) );
  NAND3_X1 U12019 ( .A1(n9263), .A2(n12070), .A3(n11686), .ZN(n12069) );
  NAND2_X1 U12020 ( .A1(n12055), .A2(n12053), .ZN(n12070) );
  INV_X1 U12021 ( .A(n12071), .ZN(n12068) );
  NOR2_X1 U12022 ( .A1(n12053), .A2(n12055), .ZN(n12071) );
  NOR2_X1 U12023 ( .A1(n12072), .A2(n12073), .ZN(n12055) );
  INV_X1 U12024 ( .A(n12074), .ZN(n12073) );
  NAND3_X1 U12025 ( .A1(n9268), .A2(n12075), .A3(n11686), .ZN(n12074) );
  NAND2_X1 U12026 ( .A1(n12051), .A2(n12049), .ZN(n12075) );
  NOR2_X1 U12027 ( .A1(n12049), .A2(n12051), .ZN(n12072) );
  NOR2_X1 U12028 ( .A1(n12076), .A2(n12077), .ZN(n12051) );
  INV_X1 U12029 ( .A(n12078), .ZN(n12077) );
  NAND3_X1 U12030 ( .A1(n9792), .A2(n12079), .A3(n11686), .ZN(n12078) );
  NAND2_X1 U12031 ( .A1(n12047), .A2(n12045), .ZN(n12079) );
  NOR2_X1 U12032 ( .A1(n12045), .A2(n12047), .ZN(n12076) );
  NOR2_X1 U12033 ( .A1(n12080), .A2(n12081), .ZN(n12047) );
  NOR3_X1 U12034 ( .A1(n8528), .A2(n12082), .A3(n8558), .ZN(n12081) );
  NOR2_X1 U12035 ( .A1(n12043), .A2(n12041), .ZN(n12082) );
  INV_X1 U12036 ( .A(n12083), .ZN(n12080) );
  NAND2_X1 U12037 ( .A1(n12041), .A2(n12043), .ZN(n12083) );
  NAND2_X1 U12038 ( .A1(n12084), .A2(n12085), .ZN(n12043) );
  INV_X1 U12039 ( .A(n12086), .ZN(n12085) );
  NOR3_X1 U12040 ( .A1(n8995), .A2(n12087), .A3(n8558), .ZN(n12086) );
  NOR2_X1 U12041 ( .A1(n12039), .A2(n12037), .ZN(n12087) );
  NAND2_X1 U12042 ( .A1(n12037), .A2(n12039), .ZN(n12084) );
  NAND2_X1 U12043 ( .A1(n12088), .A2(n12089), .ZN(n12039) );
  INV_X1 U12044 ( .A(n12090), .ZN(n12089) );
  NOR3_X1 U12045 ( .A1(n9000), .A2(n12091), .A3(n8558), .ZN(n12090) );
  NOR2_X1 U12046 ( .A1(n12035), .A2(n12033), .ZN(n12091) );
  NAND2_X1 U12047 ( .A1(n12033), .A2(n12035), .ZN(n12088) );
  NAND2_X1 U12048 ( .A1(n12092), .A2(n12093), .ZN(n12035) );
  NAND3_X1 U12049 ( .A1(n8543), .A2(n12094), .A3(n11686), .ZN(n12093) );
  INV_X1 U12050 ( .A(n12095), .ZN(n12094) );
  NOR2_X1 U12051 ( .A1(n12031), .A2(n12030), .ZN(n12095) );
  NAND2_X1 U12052 ( .A1(n12030), .A2(n12031), .ZN(n12092) );
  NAND2_X1 U12053 ( .A1(n12096), .A2(n12097), .ZN(n12031) );
  NAND3_X1 U12054 ( .A1(n9295), .A2(n12098), .A3(n11686), .ZN(n12097) );
  INV_X1 U12055 ( .A(n12099), .ZN(n12098) );
  NOR2_X1 U12056 ( .A1(n12027), .A2(n12025), .ZN(n12099) );
  NAND2_X1 U12057 ( .A1(n12025), .A2(n12027), .ZN(n12096) );
  NAND2_X1 U12058 ( .A1(n12100), .A2(n12101), .ZN(n12027) );
  NAND3_X1 U12059 ( .A1(n10846), .A2(n12102), .A3(n11686), .ZN(n12101) );
  INV_X1 U12060 ( .A(n12103), .ZN(n12102) );
  NOR2_X1 U12061 ( .A1(n12023), .A2(n12022), .ZN(n12103) );
  NAND2_X1 U12062 ( .A1(n12022), .A2(n12023), .ZN(n12100) );
  NAND2_X1 U12063 ( .A1(n12019), .A2(n12104), .ZN(n12023) );
  NAND2_X1 U12064 ( .A1(n12018), .A2(n12020), .ZN(n12104) );
  NAND2_X1 U12065 ( .A1(n12105), .A2(n12106), .ZN(n12020) );
  NAND2_X1 U12066 ( .A1(n11686), .A2(n9304), .ZN(n12106) );
  XNOR2_X1 U12067 ( .A(n12107), .B(n12108), .ZN(n12018) );
  XOR2_X1 U12068 ( .A(n12109), .B(n12110), .Z(n12108) );
  NAND2_X1 U12069 ( .A1(n9304), .A2(n12111), .ZN(n12019) );
  INV_X1 U12070 ( .A(n12105), .ZN(n12111) );
  NOR2_X1 U12071 ( .A1(n12112), .A2(n12113), .ZN(n12105) );
  INV_X1 U12072 ( .A(n12114), .ZN(n12113) );
  NAND2_X1 U12073 ( .A1(n12016), .A2(n12115), .ZN(n12114) );
  NAND2_X1 U12074 ( .A1(n12015), .A2(n12014), .ZN(n12115) );
  NOR2_X1 U12075 ( .A1(n8558), .A2(n8572), .ZN(n12016) );
  NOR2_X1 U12076 ( .A1(n12014), .A2(n12015), .ZN(n12112) );
  NOR2_X1 U12077 ( .A1(n12116), .A2(n12117), .ZN(n12015) );
  INV_X1 U12078 ( .A(n12118), .ZN(n12117) );
  NAND2_X1 U12079 ( .A1(n12012), .A2(n12119), .ZN(n12118) );
  NAND2_X1 U12080 ( .A1(n12120), .A2(n12009), .ZN(n12119) );
  NOR2_X1 U12081 ( .A1(n8558), .A2(n8582), .ZN(n12012) );
  NOR2_X1 U12082 ( .A1(n12009), .A2(n12120), .ZN(n12116) );
  INV_X1 U12083 ( .A(n12011), .ZN(n12120) );
  NAND2_X1 U12084 ( .A1(n12121), .A2(n12122), .ZN(n12011) );
  NAND2_X1 U12085 ( .A1(n12008), .A2(n12123), .ZN(n12122) );
  INV_X1 U12086 ( .A(n12124), .ZN(n12123) );
  NOR2_X1 U12087 ( .A1(n12007), .A2(n12006), .ZN(n12124) );
  NOR2_X1 U12088 ( .A1(n8558), .A2(n8591), .ZN(n12008) );
  NAND2_X1 U12089 ( .A1(n12006), .A2(n12007), .ZN(n12121) );
  NAND2_X1 U12090 ( .A1(n12125), .A2(n12126), .ZN(n12007) );
  NAND2_X1 U12091 ( .A1(n12004), .A2(n12127), .ZN(n12126) );
  INV_X1 U12092 ( .A(n12128), .ZN(n12127) );
  NOR2_X1 U12093 ( .A1(n12003), .A2(n12001), .ZN(n12128) );
  NOR2_X1 U12094 ( .A1(n8558), .A2(n8562), .ZN(n12004) );
  NAND2_X1 U12095 ( .A1(n12001), .A2(n12003), .ZN(n12125) );
  NAND2_X1 U12096 ( .A1(n12129), .A2(n12130), .ZN(n12003) );
  NAND2_X1 U12097 ( .A1(n12000), .A2(n12131), .ZN(n12130) );
  INV_X1 U12098 ( .A(n12132), .ZN(n12131) );
  NOR2_X1 U12099 ( .A1(n11999), .A2(n11998), .ZN(n12132) );
  NOR2_X1 U12100 ( .A1(n8558), .A2(n8545), .ZN(n12000) );
  NAND2_X1 U12101 ( .A1(n11998), .A2(n11999), .ZN(n12129) );
  NAND2_X1 U12102 ( .A1(n12133), .A2(n12134), .ZN(n11999) );
  NAND2_X1 U12103 ( .A1(n11996), .A2(n12135), .ZN(n12134) );
  NAND2_X1 U12104 ( .A1(n11995), .A2(n11993), .ZN(n12135) );
  NOR2_X1 U12105 ( .A1(n8558), .A2(n8569), .ZN(n11996) );
  INV_X1 U12106 ( .A(n12136), .ZN(n12133) );
  NOR2_X1 U12107 ( .A1(n11993), .A2(n11995), .ZN(n12136) );
  NOR2_X1 U12108 ( .A1(n12137), .A2(n12138), .ZN(n11995) );
  INV_X1 U12109 ( .A(n12139), .ZN(n12138) );
  NAND2_X1 U12110 ( .A1(n11992), .A2(n12140), .ZN(n12139) );
  NAND2_X1 U12111 ( .A1(n11991), .A2(n11990), .ZN(n12140) );
  NOR2_X1 U12112 ( .A1(n8558), .A2(n8593), .ZN(n11992) );
  NOR2_X1 U12113 ( .A1(n11990), .A2(n11991), .ZN(n12137) );
  INV_X1 U12114 ( .A(n12141), .ZN(n11991) );
  NAND2_X1 U12115 ( .A1(n12142), .A2(n12143), .ZN(n12141) );
  NAND2_X1 U12116 ( .A1(n11987), .A2(n12144), .ZN(n12143) );
  INV_X1 U12117 ( .A(n12145), .ZN(n12144) );
  NOR2_X1 U12118 ( .A1(n11988), .A2(n11986), .ZN(n12145) );
  NOR2_X1 U12119 ( .A1(n8558), .A2(n8583), .ZN(n11987) );
  NAND2_X1 U12120 ( .A1(n11986), .A2(n11988), .ZN(n12142) );
  NAND2_X1 U12121 ( .A1(n12146), .A2(n12147), .ZN(n11988) );
  NAND2_X1 U12122 ( .A1(n11984), .A2(n12148), .ZN(n12147) );
  INV_X1 U12123 ( .A(n12149), .ZN(n12148) );
  NOR2_X1 U12124 ( .A1(n11983), .A2(n11982), .ZN(n12149) );
  NOR2_X1 U12125 ( .A1(n8558), .A2(n8580), .ZN(n11984) );
  NAND2_X1 U12126 ( .A1(n11982), .A2(n11983), .ZN(n12146) );
  NAND2_X1 U12127 ( .A1(n12150), .A2(n12151), .ZN(n11983) );
  NAND2_X1 U12128 ( .A1(n11980), .A2(n12152), .ZN(n12151) );
  NAND2_X1 U12129 ( .A1(n11979), .A2(n11977), .ZN(n12152) );
  NOR2_X1 U12130 ( .A1(n8558), .A2(n8588), .ZN(n11980) );
  INV_X1 U12131 ( .A(n12153), .ZN(n12150) );
  NOR2_X1 U12132 ( .A1(n11977), .A2(n11979), .ZN(n12153) );
  NOR2_X1 U12133 ( .A1(n12154), .A2(n12155), .ZN(n11979) );
  INV_X1 U12134 ( .A(n12156), .ZN(n12155) );
  NAND2_X1 U12135 ( .A1(n11976), .A2(n12157), .ZN(n12156) );
  NAND2_X1 U12136 ( .A1(n11975), .A2(n11974), .ZN(n12157) );
  NOR2_X1 U12137 ( .A1(n11685), .A2(n8551), .ZN(n11976) );
  NOR2_X1 U12138 ( .A1(n11974), .A2(n11975), .ZN(n12154) );
  NOR2_X1 U12139 ( .A1(n12158), .A2(n12159), .ZN(n11975) );
  INV_X1 U12140 ( .A(n12160), .ZN(n12159) );
  NAND2_X1 U12141 ( .A1(n11972), .A2(n12161), .ZN(n12160) );
  NAND2_X1 U12142 ( .A1(n11971), .A2(n11970), .ZN(n12161) );
  NOR2_X1 U12143 ( .A1(n11685), .A2(n8563), .ZN(n11972) );
  NOR2_X1 U12144 ( .A1(n11970), .A2(n11971), .ZN(n12158) );
  NOR2_X1 U12145 ( .A1(n12162), .A2(n12163), .ZN(n11971) );
  INV_X1 U12146 ( .A(n12164), .ZN(n12163) );
  NAND2_X1 U12147 ( .A1(n11967), .A2(n12165), .ZN(n12164) );
  NAND2_X1 U12148 ( .A1(n11968), .A2(n11966), .ZN(n12165) );
  NOR2_X1 U12149 ( .A1(n11685), .A2(n8548), .ZN(n11967) );
  NOR2_X1 U12150 ( .A1(n11966), .A2(n11968), .ZN(n12162) );
  NOR2_X1 U12151 ( .A1(n12166), .A2(n12167), .ZN(n11968) );
  INV_X1 U12152 ( .A(n12168), .ZN(n12167) );
  NAND2_X1 U12153 ( .A1(n11964), .A2(n12169), .ZN(n12168) );
  NAND2_X1 U12154 ( .A1(n11963), .A2(n11962), .ZN(n12169) );
  NOR2_X1 U12155 ( .A1(n11685), .A2(n8584), .ZN(n11964) );
  NOR2_X1 U12156 ( .A1(n11962), .A2(n11963), .ZN(n12166) );
  NOR2_X1 U12157 ( .A1(n12170), .A2(n12171), .ZN(n11963) );
  INV_X1 U12158 ( .A(n12172), .ZN(n12171) );
  NAND2_X1 U12159 ( .A1(n11959), .A2(n12173), .ZN(n12172) );
  NAND2_X1 U12160 ( .A1(n11960), .A2(n11958), .ZN(n12173) );
  NOR2_X1 U12161 ( .A1(n11685), .A2(n8535), .ZN(n11959) );
  NOR2_X1 U12162 ( .A1(n11958), .A2(n11960), .ZN(n12170) );
  NOR2_X1 U12163 ( .A1(n12174), .A2(n12175), .ZN(n11960) );
  INV_X1 U12164 ( .A(n12176), .ZN(n12175) );
  NAND2_X1 U12165 ( .A1(n11955), .A2(n12177), .ZN(n12176) );
  NAND2_X1 U12166 ( .A1(n11956), .A2(n11954), .ZN(n12177) );
  NOR2_X1 U12167 ( .A1(n11685), .A2(n8568), .ZN(n11955) );
  NOR2_X1 U12168 ( .A1(n11954), .A2(n11956), .ZN(n12174) );
  NOR2_X1 U12169 ( .A1(n12178), .A2(n12179), .ZN(n11956) );
  INV_X1 U12170 ( .A(n12180), .ZN(n12179) );
  NAND2_X1 U12171 ( .A1(n11951), .A2(n12181), .ZN(n12180) );
  NAND2_X1 U12172 ( .A1(n11952), .A2(n11950), .ZN(n12181) );
  NOR2_X1 U12173 ( .A1(n11685), .A2(n8574), .ZN(n11951) );
  NOR2_X1 U12174 ( .A1(n11950), .A2(n11952), .ZN(n12178) );
  NOR2_X1 U12175 ( .A1(n12182), .A2(n12183), .ZN(n11952) );
  INV_X1 U12176 ( .A(n12184), .ZN(n12183) );
  NAND2_X1 U12177 ( .A1(n11947), .A2(n12185), .ZN(n12184) );
  NAND2_X1 U12178 ( .A1(n11948), .A2(n11946), .ZN(n12185) );
  NOR2_X1 U12179 ( .A1(n11685), .A2(n8565), .ZN(n11947) );
  NOR2_X1 U12180 ( .A1(n11946), .A2(n11948), .ZN(n12182) );
  NOR2_X1 U12181 ( .A1(n12186), .A2(n12187), .ZN(n11948) );
  INV_X1 U12182 ( .A(n12188), .ZN(n12187) );
  NAND2_X1 U12183 ( .A1(n11941), .A2(n12189), .ZN(n12188) );
  NAND2_X1 U12184 ( .A1(n11944), .A2(n11943), .ZN(n12189) );
  NOR2_X1 U12185 ( .A1(n11685), .A2(n8567), .ZN(n11941) );
  NOR2_X1 U12186 ( .A1(n11943), .A2(n11944), .ZN(n12186) );
  INV_X1 U12187 ( .A(n12190), .ZN(n11944) );
  NAND2_X1 U12188 ( .A1(n12191), .A2(n12192), .ZN(n12190) );
  NAND2_X1 U12189 ( .A1(n11936), .A2(n12193), .ZN(n12192) );
  NAND2_X1 U12190 ( .A1(n8624), .A2(n12194), .ZN(n12193) );
  NAND2_X1 U12191 ( .A1(n8578), .A2(n8585), .ZN(n12194) );
  NAND2_X1 U12192 ( .A1(n12196), .A2(n12197), .ZN(n12191) );
  NAND2_X1 U12193 ( .A1(n8630), .A2(n12198), .ZN(n12197) );
  NAND2_X1 U12194 ( .A1(n8539), .A2(n8575), .ZN(n12198) );
  NAND3_X1 U12195 ( .A1(n11936), .A2(n8537), .A3(n11686), .ZN(n11943) );
  INV_X1 U12196 ( .A(n11685), .ZN(n11686) );
  XNOR2_X1 U12197 ( .A(n12199), .B(n12200), .ZN(n11685) );
  XOR2_X1 U12198 ( .A(d_19_), .B(c_19_), .Z(n12200) );
  XOR2_X1 U12199 ( .A(n12201), .B(n12202), .Z(n11946) );
  XNOR2_X1 U12200 ( .A(n12203), .B(n12204), .ZN(n12202) );
  XOR2_X1 U12201 ( .A(n12205), .B(n12206), .Z(n11950) );
  XNOR2_X1 U12202 ( .A(n12207), .B(n12208), .ZN(n12205) );
  XOR2_X1 U12203 ( .A(n12209), .B(n12210), .Z(n11954) );
  XNOR2_X1 U12204 ( .A(n12211), .B(n12212), .ZN(n12209) );
  XOR2_X1 U12205 ( .A(n12213), .B(n12214), .Z(n11958) );
  XNOR2_X1 U12206 ( .A(n12215), .B(n12216), .ZN(n12213) );
  XOR2_X1 U12207 ( .A(n12217), .B(n12218), .Z(n11962) );
  XNOR2_X1 U12208 ( .A(n12219), .B(n12220), .ZN(n12217) );
  NOR2_X1 U12209 ( .A1(n8535), .A2(n8575), .ZN(n12220) );
  XOR2_X1 U12210 ( .A(n12221), .B(n12222), .Z(n11966) );
  XNOR2_X1 U12211 ( .A(n12223), .B(n12224), .ZN(n12221) );
  NOR2_X1 U12212 ( .A1(n8584), .A2(n8575), .ZN(n12224) );
  XNOR2_X1 U12213 ( .A(n12225), .B(n12226), .ZN(n11970) );
  XNOR2_X1 U12214 ( .A(n12227), .B(n12228), .ZN(n12226) );
  NAND2_X1 U12215 ( .A1(n11936), .A2(n9107), .ZN(n12228) );
  XOR2_X1 U12216 ( .A(n12229), .B(n12230), .Z(n11974) );
  XNOR2_X1 U12217 ( .A(n12231), .B(n12232), .ZN(n12229) );
  NOR2_X1 U12218 ( .A1(n8563), .A2(n8575), .ZN(n12232) );
  XOR2_X1 U12219 ( .A(n12233), .B(n12234), .Z(n11977) );
  XNOR2_X1 U12220 ( .A(n12235), .B(n12236), .ZN(n12233) );
  NOR2_X1 U12221 ( .A1(n8551), .A2(n8575), .ZN(n12236) );
  XNOR2_X1 U12222 ( .A(n12237), .B(n12238), .ZN(n11982) );
  XNOR2_X1 U12223 ( .A(n12239), .B(n12240), .ZN(n12237) );
  NOR2_X1 U12224 ( .A1(n8588), .A2(n8575), .ZN(n12240) );
  XNOR2_X1 U12225 ( .A(n12241), .B(n12242), .ZN(n11986) );
  XNOR2_X1 U12226 ( .A(n12243), .B(n12244), .ZN(n12241) );
  NOR2_X1 U12227 ( .A1(n8580), .A2(n8575), .ZN(n12244) );
  XOR2_X1 U12228 ( .A(n12245), .B(n12246), .Z(n11990) );
  XNOR2_X1 U12229 ( .A(n12247), .B(n12248), .ZN(n12245) );
  NOR2_X1 U12230 ( .A1(n8583), .A2(n8575), .ZN(n12248) );
  XOR2_X1 U12231 ( .A(n12249), .B(n12250), .Z(n11993) );
  XNOR2_X1 U12232 ( .A(n12251), .B(n12252), .ZN(n12249) );
  NOR2_X1 U12233 ( .A1(n8593), .A2(n8575), .ZN(n12252) );
  XNOR2_X1 U12234 ( .A(n12253), .B(n12254), .ZN(n11998) );
  XNOR2_X1 U12235 ( .A(n12255), .B(n12256), .ZN(n12253) );
  NOR2_X1 U12236 ( .A1(n9050), .A2(n8575), .ZN(n12256) );
  XNOR2_X1 U12237 ( .A(n12257), .B(n12258), .ZN(n12001) );
  XNOR2_X1 U12238 ( .A(n12259), .B(n12260), .ZN(n12257) );
  NOR2_X1 U12239 ( .A1(n8545), .A2(n8575), .ZN(n12260) );
  XNOR2_X1 U12240 ( .A(n12261), .B(n12262), .ZN(n12006) );
  XNOR2_X1 U12241 ( .A(n12263), .B(n12264), .ZN(n12261) );
  NOR2_X1 U12242 ( .A1(n9041), .A2(n8575), .ZN(n12264) );
  XOR2_X1 U12243 ( .A(n12265), .B(n12266), .Z(n12009) );
  XNOR2_X1 U12244 ( .A(n12267), .B(n12268), .ZN(n12265) );
  NOR2_X1 U12245 ( .A1(n8591), .A2(n8575), .ZN(n12268) );
  XNOR2_X1 U12246 ( .A(n12269), .B(n12270), .ZN(n12014) );
  XNOR2_X1 U12247 ( .A(n12271), .B(n12272), .ZN(n12270) );
  NAND2_X1 U12248 ( .A1(n11936), .A2(n9313), .ZN(n12272) );
  XOR2_X1 U12249 ( .A(n12273), .B(n12274), .Z(n12022) );
  XOR2_X1 U12250 ( .A(n12275), .B(n12276), .Z(n12274) );
  XOR2_X1 U12251 ( .A(n12277), .B(n12278), .Z(n12025) );
  XOR2_X1 U12252 ( .A(n12279), .B(n12280), .Z(n12277) );
  XOR2_X1 U12253 ( .A(n12281), .B(n12282), .Z(n12030) );
  XNOR2_X1 U12254 ( .A(n12283), .B(n12284), .ZN(n12282) );
  XNOR2_X1 U12255 ( .A(n12285), .B(n12286), .ZN(n12033) );
  XNOR2_X1 U12256 ( .A(n12287), .B(n12288), .ZN(n12285) );
  XNOR2_X1 U12257 ( .A(n12289), .B(n12290), .ZN(n12037) );
  XNOR2_X1 U12258 ( .A(n12291), .B(n12292), .ZN(n12290) );
  XOR2_X1 U12259 ( .A(n12293), .B(n12294), .Z(n12041) );
  XOR2_X1 U12260 ( .A(n12295), .B(n12296), .Z(n12293) );
  XNOR2_X1 U12261 ( .A(n12297), .B(n12298), .ZN(n12045) );
  XOR2_X1 U12262 ( .A(n12299), .B(n12300), .Z(n12297) );
  XNOR2_X1 U12263 ( .A(n12301), .B(n12302), .ZN(n12049) );
  XOR2_X1 U12264 ( .A(n12303), .B(n12304), .Z(n12301) );
  XNOR2_X1 U12265 ( .A(n12305), .B(n12306), .ZN(n12053) );
  XOR2_X1 U12266 ( .A(n12307), .B(n12308), .Z(n12305) );
  XNOR2_X1 U12267 ( .A(n12309), .B(n12310), .ZN(n12059) );
  NAND2_X1 U12268 ( .A1(n12311), .A2(n12312), .ZN(n12309) );
  XOR2_X1 U12269 ( .A(n12313), .B(n12314), .Z(n12058) );
  NAND2_X1 U12270 ( .A1(n12315), .A2(n12316), .ZN(n12313) );
  INV_X1 U12271 ( .A(n8913), .ZN(n8840) );
  NOR2_X1 U12272 ( .A1(n8917), .A2(n8918), .ZN(n8913) );
  NAND2_X1 U12273 ( .A1(n8918), .A2(n8917), .ZN(n12063) );
  XOR2_X1 U12274 ( .A(n12317), .B(n12318), .Z(n8917) );
  XNOR2_X1 U12275 ( .A(n12319), .B(n12320), .ZN(n12318) );
  INV_X1 U12276 ( .A(n12321), .ZN(n8918) );
  NAND2_X1 U12277 ( .A1(n12315), .A2(n12322), .ZN(n12321) );
  NAND2_X1 U12278 ( .A1(n12314), .A2(n12316), .ZN(n12322) );
  NAND2_X1 U12279 ( .A1(n12323), .A2(n12324), .ZN(n12316) );
  NAND2_X1 U12280 ( .A1(n11936), .A2(n8872), .ZN(n12324) );
  INV_X1 U12281 ( .A(n12325), .ZN(n12323) );
  XNOR2_X1 U12282 ( .A(n12326), .B(n12327), .ZN(n12314) );
  XOR2_X1 U12283 ( .A(n12328), .B(n12329), .Z(n12326) );
  NAND2_X1 U12284 ( .A1(n8592), .A2(n12325), .ZN(n12315) );
  NAND2_X1 U12285 ( .A1(n12311), .A2(n12330), .ZN(n12325) );
  NAND2_X1 U12286 ( .A1(n12310), .A2(n12312), .ZN(n12330) );
  NAND2_X1 U12287 ( .A1(n12331), .A2(n12332), .ZN(n12312) );
  NAND2_X1 U12288 ( .A1(n11936), .A2(n9263), .ZN(n12332) );
  INV_X1 U12289 ( .A(n12333), .ZN(n12331) );
  XOR2_X1 U12290 ( .A(n12334), .B(n12335), .Z(n12310) );
  XOR2_X1 U12291 ( .A(n12336), .B(n12337), .Z(n12334) );
  NOR2_X1 U12292 ( .A1(n8552), .A2(n8578), .ZN(n12337) );
  NAND2_X1 U12293 ( .A1(n9263), .A2(n12333), .ZN(n12311) );
  NAND2_X1 U12294 ( .A1(n12338), .A2(n12339), .ZN(n12333) );
  NAND2_X1 U12295 ( .A1(n12308), .A2(n12340), .ZN(n12339) );
  INV_X1 U12296 ( .A(n12341), .ZN(n12340) );
  NOR2_X1 U12297 ( .A1(n12307), .A2(n12306), .ZN(n12341) );
  NOR2_X1 U12298 ( .A1(n8575), .A2(n8552), .ZN(n12308) );
  NAND2_X1 U12299 ( .A1(n12306), .A2(n12307), .ZN(n12338) );
  NAND2_X1 U12300 ( .A1(n12342), .A2(n12343), .ZN(n12307) );
  NAND2_X1 U12301 ( .A1(n12304), .A2(n12344), .ZN(n12343) );
  INV_X1 U12302 ( .A(n12345), .ZN(n12344) );
  NOR2_X1 U12303 ( .A1(n12303), .A2(n12302), .ZN(n12345) );
  NOR2_X1 U12304 ( .A1(n8575), .A2(n8527), .ZN(n12304) );
  NAND2_X1 U12305 ( .A1(n12302), .A2(n12303), .ZN(n12342) );
  NAND2_X1 U12306 ( .A1(n12346), .A2(n12347), .ZN(n12303) );
  NAND2_X1 U12307 ( .A1(n12300), .A2(n12348), .ZN(n12347) );
  INV_X1 U12308 ( .A(n12349), .ZN(n12348) );
  NOR2_X1 U12309 ( .A1(n12299), .A2(n12298), .ZN(n12349) );
  NOR2_X1 U12310 ( .A1(n8575), .A2(n8528), .ZN(n12300) );
  NAND2_X1 U12311 ( .A1(n12298), .A2(n12299), .ZN(n12346) );
  NAND2_X1 U12312 ( .A1(n12350), .A2(n12351), .ZN(n12299) );
  NAND2_X1 U12313 ( .A1(n12296), .A2(n12352), .ZN(n12351) );
  INV_X1 U12314 ( .A(n12353), .ZN(n12352) );
  NOR2_X1 U12315 ( .A1(n12295), .A2(n12294), .ZN(n12353) );
  NOR2_X1 U12316 ( .A1(n8575), .A2(n8564), .ZN(n12296) );
  NAND2_X1 U12317 ( .A1(n12294), .A2(n12295), .ZN(n12350) );
  NAND2_X1 U12318 ( .A1(n12354), .A2(n12355), .ZN(n12295) );
  NAND2_X1 U12319 ( .A1(n12292), .A2(n12356), .ZN(n12355) );
  INV_X1 U12320 ( .A(n12357), .ZN(n12356) );
  NOR2_X1 U12321 ( .A1(n12291), .A2(n12289), .ZN(n12357) );
  NOR2_X1 U12322 ( .A1(n8575), .A2(n8555), .ZN(n12292) );
  NAND2_X1 U12323 ( .A1(n12289), .A2(n12291), .ZN(n12354) );
  NAND2_X1 U12324 ( .A1(n12358), .A2(n12359), .ZN(n12291) );
  NAND2_X1 U12325 ( .A1(n12288), .A2(n12360), .ZN(n12359) );
  NAND2_X1 U12326 ( .A1(n12287), .A2(n12286), .ZN(n12360) );
  NOR2_X1 U12327 ( .A1(n8575), .A2(n8544), .ZN(n12288) );
  INV_X1 U12328 ( .A(n12361), .ZN(n12358) );
  NOR2_X1 U12329 ( .A1(n12286), .A2(n12287), .ZN(n12361) );
  NOR2_X1 U12330 ( .A1(n12362), .A2(n12363), .ZN(n12287) );
  INV_X1 U12331 ( .A(n12364), .ZN(n12363) );
  NAND2_X1 U12332 ( .A1(n12284), .A2(n12365), .ZN(n12364) );
  NAND2_X1 U12333 ( .A1(n12366), .A2(n12281), .ZN(n12365) );
  NOR2_X1 U12334 ( .A1(n11935), .A2(n8560), .ZN(n12284) );
  NOR2_X1 U12335 ( .A1(n12281), .A2(n12366), .ZN(n12362) );
  INV_X1 U12336 ( .A(n12283), .ZN(n12366) );
  NAND2_X1 U12337 ( .A1(n12367), .A2(n12368), .ZN(n12283) );
  NAND2_X1 U12338 ( .A1(n12280), .A2(n12369), .ZN(n12368) );
  INV_X1 U12339 ( .A(n12370), .ZN(n12369) );
  NOR2_X1 U12340 ( .A1(n12279), .A2(n12278), .ZN(n12370) );
  NOR2_X1 U12341 ( .A1(n11935), .A2(n8594), .ZN(n12280) );
  NAND2_X1 U12342 ( .A1(n12278), .A2(n12279), .ZN(n12367) );
  NAND2_X1 U12343 ( .A1(n12371), .A2(n12372), .ZN(n12279) );
  NAND2_X1 U12344 ( .A1(n12276), .A2(n12373), .ZN(n12372) );
  NAND2_X1 U12345 ( .A1(n12275), .A2(n12273), .ZN(n12373) );
  NOR2_X1 U12346 ( .A1(n11935), .A2(n8556), .ZN(n12276) );
  INV_X1 U12347 ( .A(n12374), .ZN(n12371) );
  NOR2_X1 U12348 ( .A1(n12273), .A2(n12275), .ZN(n12374) );
  NOR2_X1 U12349 ( .A1(n12375), .A2(n12376), .ZN(n12275) );
  NOR2_X1 U12350 ( .A1(n12110), .A2(n12377), .ZN(n12376) );
  NOR2_X1 U12351 ( .A1(n12109), .A2(n12107), .ZN(n12377) );
  NAND2_X1 U12352 ( .A1(n11936), .A2(n9209), .ZN(n12110) );
  INV_X1 U12353 ( .A(n12378), .ZN(n12375) );
  NAND2_X1 U12354 ( .A1(n12107), .A2(n12109), .ZN(n12378) );
  NAND2_X1 U12355 ( .A1(n12379), .A2(n12380), .ZN(n12109) );
  NAND3_X1 U12356 ( .A1(n9313), .A2(n12381), .A3(n11936), .ZN(n12380) );
  NAND2_X1 U12357 ( .A1(n12271), .A2(n12269), .ZN(n12381) );
  INV_X1 U12358 ( .A(n12382), .ZN(n12379) );
  NOR2_X1 U12359 ( .A1(n12269), .A2(n12271), .ZN(n12382) );
  NOR2_X1 U12360 ( .A1(n12383), .A2(n12384), .ZN(n12271) );
  INV_X1 U12361 ( .A(n12385), .ZN(n12384) );
  NAND3_X1 U12362 ( .A1(n9721), .A2(n12386), .A3(n11936), .ZN(n12385) );
  NAND2_X1 U12363 ( .A1(n12267), .A2(n12266), .ZN(n12386) );
  NOR2_X1 U12364 ( .A1(n12266), .A2(n12267), .ZN(n12383) );
  NOR2_X1 U12365 ( .A1(n12387), .A2(n12388), .ZN(n12267) );
  INV_X1 U12366 ( .A(n12389), .ZN(n12388) );
  NAND3_X1 U12367 ( .A1(n9322), .A2(n12390), .A3(n11936), .ZN(n12389) );
  NAND2_X1 U12368 ( .A1(n12263), .A2(n12262), .ZN(n12390) );
  NOR2_X1 U12369 ( .A1(n12262), .A2(n12263), .ZN(n12387) );
  NOR2_X1 U12370 ( .A1(n12391), .A2(n12392), .ZN(n12263) );
  NOR3_X1 U12371 ( .A1(n8545), .A2(n12393), .A3(n8575), .ZN(n12392) );
  INV_X1 U12372 ( .A(n12394), .ZN(n12393) );
  NAND2_X1 U12373 ( .A1(n12259), .A2(n12258), .ZN(n12394) );
  NOR2_X1 U12374 ( .A1(n12258), .A2(n12259), .ZN(n12391) );
  NOR2_X1 U12375 ( .A1(n12395), .A2(n12396), .ZN(n12259) );
  INV_X1 U12376 ( .A(n12397), .ZN(n12396) );
  NAND3_X1 U12377 ( .A1(n9331), .A2(n12398), .A3(n11936), .ZN(n12397) );
  NAND2_X1 U12378 ( .A1(n12255), .A2(n12254), .ZN(n12398) );
  NOR2_X1 U12379 ( .A1(n12254), .A2(n12255), .ZN(n12395) );
  NOR2_X1 U12380 ( .A1(n12399), .A2(n12400), .ZN(n12255) );
  NOR3_X1 U12381 ( .A1(n9056), .A2(n12401), .A3(n8575), .ZN(n12400) );
  INV_X1 U12382 ( .A(n12402), .ZN(n12401) );
  NAND2_X1 U12383 ( .A1(n12251), .A2(n12250), .ZN(n12402) );
  NOR2_X1 U12384 ( .A1(n12250), .A2(n12251), .ZN(n12399) );
  NOR2_X1 U12385 ( .A1(n12403), .A2(n12404), .ZN(n12251) );
  INV_X1 U12386 ( .A(n12405), .ZN(n12404) );
  NAND3_X1 U12387 ( .A1(n9340), .A2(n12406), .A3(n11936), .ZN(n12405) );
  NAND2_X1 U12388 ( .A1(n12247), .A2(n12246), .ZN(n12406) );
  NOR2_X1 U12389 ( .A1(n12246), .A2(n12247), .ZN(n12403) );
  NOR2_X1 U12390 ( .A1(n12407), .A2(n12408), .ZN(n12247) );
  NOR3_X1 U12391 ( .A1(n9066), .A2(n12409), .A3(n8575), .ZN(n12408) );
  INV_X1 U12392 ( .A(n12410), .ZN(n12409) );
  NAND2_X1 U12393 ( .A1(n12243), .A2(n12242), .ZN(n12410) );
  NOR2_X1 U12394 ( .A1(n12242), .A2(n12243), .ZN(n12407) );
  NOR2_X1 U12395 ( .A1(n12411), .A2(n12412), .ZN(n12243) );
  INV_X1 U12396 ( .A(n12413), .ZN(n12412) );
  NAND3_X1 U12397 ( .A1(n9080), .A2(n12414), .A3(n11936), .ZN(n12413) );
  NAND2_X1 U12398 ( .A1(n12239), .A2(n12238), .ZN(n12414) );
  NOR2_X1 U12399 ( .A1(n12238), .A2(n12239), .ZN(n12411) );
  NOR2_X1 U12400 ( .A1(n12415), .A2(n12416), .ZN(n12239) );
  NOR3_X1 U12401 ( .A1(n8551), .A2(n12417), .A3(n8575), .ZN(n12416) );
  INV_X1 U12402 ( .A(n12418), .ZN(n12417) );
  NAND2_X1 U12403 ( .A1(n12235), .A2(n12234), .ZN(n12418) );
  NOR2_X1 U12404 ( .A1(n12234), .A2(n12235), .ZN(n12415) );
  NOR2_X1 U12405 ( .A1(n12419), .A2(n12420), .ZN(n12235) );
  INV_X1 U12406 ( .A(n12421), .ZN(n12420) );
  NAND3_X1 U12407 ( .A1(n9098), .A2(n12422), .A3(n11936), .ZN(n12421) );
  NAND2_X1 U12408 ( .A1(n12231), .A2(n12230), .ZN(n12422) );
  NOR2_X1 U12409 ( .A1(n12230), .A2(n12231), .ZN(n12419) );
  NOR2_X1 U12410 ( .A1(n12423), .A2(n12424), .ZN(n12231) );
  NOR3_X1 U12411 ( .A1(n8548), .A2(n12425), .A3(n8575), .ZN(n12424) );
  INV_X1 U12412 ( .A(n12426), .ZN(n12425) );
  NAND2_X1 U12413 ( .A1(n12227), .A2(n12225), .ZN(n12426) );
  NOR2_X1 U12414 ( .A1(n12225), .A2(n12227), .ZN(n12423) );
  NOR2_X1 U12415 ( .A1(n12427), .A2(n12428), .ZN(n12227) );
  INV_X1 U12416 ( .A(n12429), .ZN(n12428) );
  NAND3_X1 U12417 ( .A1(n9112), .A2(n12430), .A3(n11936), .ZN(n12429) );
  NAND2_X1 U12418 ( .A1(n12223), .A2(n12222), .ZN(n12430) );
  NOR2_X1 U12419 ( .A1(n12222), .A2(n12223), .ZN(n12427) );
  NOR2_X1 U12420 ( .A1(n12431), .A2(n12432), .ZN(n12223) );
  INV_X1 U12421 ( .A(n12433), .ZN(n12432) );
  NAND3_X1 U12422 ( .A1(n9121), .A2(n12434), .A3(n11936), .ZN(n12433) );
  NAND2_X1 U12423 ( .A1(n12219), .A2(n12218), .ZN(n12434) );
  NOR2_X1 U12424 ( .A1(n12218), .A2(n12219), .ZN(n12431) );
  NOR2_X1 U12425 ( .A1(n12435), .A2(n12436), .ZN(n12219) );
  INV_X1 U12426 ( .A(n12437), .ZN(n12436) );
  NAND2_X1 U12427 ( .A1(n12215), .A2(n12438), .ZN(n12437) );
  NAND2_X1 U12428 ( .A1(n12216), .A2(n12214), .ZN(n12438) );
  NOR2_X1 U12429 ( .A1(n11935), .A2(n8568), .ZN(n12215) );
  NOR2_X1 U12430 ( .A1(n12214), .A2(n12216), .ZN(n12435) );
  NOR2_X1 U12431 ( .A1(n12439), .A2(n12440), .ZN(n12216) );
  INV_X1 U12432 ( .A(n12441), .ZN(n12440) );
  NAND2_X1 U12433 ( .A1(n12211), .A2(n12442), .ZN(n12441) );
  NAND2_X1 U12434 ( .A1(n12212), .A2(n12210), .ZN(n12442) );
  NOR2_X1 U12435 ( .A1(n11935), .A2(n8574), .ZN(n12211) );
  NOR2_X1 U12436 ( .A1(n12210), .A2(n12212), .ZN(n12439) );
  NOR2_X1 U12437 ( .A1(n12443), .A2(n12444), .ZN(n12212) );
  INV_X1 U12438 ( .A(n12445), .ZN(n12444) );
  NAND2_X1 U12439 ( .A1(n12207), .A2(n12446), .ZN(n12445) );
  NAND2_X1 U12440 ( .A1(n12208), .A2(n12206), .ZN(n12446) );
  NOR2_X1 U12441 ( .A1(n11935), .A2(n8565), .ZN(n12207) );
  NOR2_X1 U12442 ( .A1(n12206), .A2(n12208), .ZN(n12443) );
  NOR2_X1 U12443 ( .A1(n12447), .A2(n12448), .ZN(n12208) );
  INV_X1 U12444 ( .A(n12449), .ZN(n12448) );
  NAND2_X1 U12445 ( .A1(n12201), .A2(n12450), .ZN(n12449) );
  NAND2_X1 U12446 ( .A1(n12204), .A2(n12203), .ZN(n12450) );
  NOR2_X1 U12447 ( .A1(n11935), .A2(n8567), .ZN(n12201) );
  NOR2_X1 U12448 ( .A1(n12203), .A2(n12204), .ZN(n12447) );
  INV_X1 U12449 ( .A(n12451), .ZN(n12204) );
  NAND2_X1 U12450 ( .A1(n12452), .A2(n12453), .ZN(n12451) );
  NAND2_X1 U12451 ( .A1(n12196), .A2(n12454), .ZN(n12453) );
  NAND2_X1 U12452 ( .A1(n8624), .A2(n12455), .ZN(n12454) );
  NAND2_X1 U12453 ( .A1(n8587), .A2(n8585), .ZN(n12455) );
  NAND2_X1 U12454 ( .A1(n12457), .A2(n12458), .ZN(n12452) );
  NAND2_X1 U12455 ( .A1(n8630), .A2(n12459), .ZN(n12458) );
  NAND2_X1 U12456 ( .A1(n8539), .A2(n8578), .ZN(n12459) );
  NAND3_X1 U12457 ( .A1(n12196), .A2(n8537), .A3(n11936), .ZN(n12203) );
  INV_X1 U12458 ( .A(n11935), .ZN(n11936) );
  XNOR2_X1 U12459 ( .A(n12460), .B(n12461), .ZN(n11935) );
  XOR2_X1 U12460 ( .A(d_18_), .B(c_18_), .Z(n12461) );
  XOR2_X1 U12461 ( .A(n12462), .B(n12463), .Z(n12206) );
  XNOR2_X1 U12462 ( .A(n12464), .B(n12465), .ZN(n12463) );
  XOR2_X1 U12463 ( .A(n12466), .B(n12467), .Z(n12210) );
  XNOR2_X1 U12464 ( .A(n12468), .B(n12469), .ZN(n12466) );
  XOR2_X1 U12465 ( .A(n12470), .B(n12471), .Z(n12214) );
  XNOR2_X1 U12466 ( .A(n12472), .B(n12473), .ZN(n12470) );
  XOR2_X1 U12467 ( .A(n12474), .B(n12475), .Z(n12218) );
  XNOR2_X1 U12468 ( .A(n12476), .B(n12477), .ZN(n12474) );
  XOR2_X1 U12469 ( .A(n12478), .B(n12479), .Z(n12222) );
  XNOR2_X1 U12470 ( .A(n12480), .B(n12481), .ZN(n12478) );
  XOR2_X1 U12471 ( .A(n12482), .B(n12483), .Z(n12225) );
  XNOR2_X1 U12472 ( .A(n12484), .B(n12485), .ZN(n12482) );
  XOR2_X1 U12473 ( .A(n12486), .B(n12487), .Z(n12230) );
  XNOR2_X1 U12474 ( .A(n12488), .B(n12489), .ZN(n12486) );
  XNOR2_X1 U12475 ( .A(n12490), .B(n12491), .ZN(n12234) );
  XOR2_X1 U12476 ( .A(n12492), .B(n12493), .Z(n12491) );
  XNOR2_X1 U12477 ( .A(n12494), .B(n12495), .ZN(n12238) );
  XOR2_X1 U12478 ( .A(n12496), .B(n12497), .Z(n12494) );
  XNOR2_X1 U12479 ( .A(n12498), .B(n12499), .ZN(n12242) );
  XOR2_X1 U12480 ( .A(n12500), .B(n12501), .Z(n12498) );
  XOR2_X1 U12481 ( .A(n12502), .B(n12503), .Z(n12246) );
  XNOR2_X1 U12482 ( .A(n12504), .B(n12505), .ZN(n12502) );
  XNOR2_X1 U12483 ( .A(n12506), .B(n12507), .ZN(n12250) );
  XOR2_X1 U12484 ( .A(n12508), .B(n12509), .Z(n12507) );
  XNOR2_X1 U12485 ( .A(n12510), .B(n12511), .ZN(n12254) );
  XOR2_X1 U12486 ( .A(n12512), .B(n12513), .Z(n12510) );
  XOR2_X1 U12487 ( .A(n12514), .B(n12515), .Z(n12258) );
  XNOR2_X1 U12488 ( .A(n12516), .B(n12517), .ZN(n12515) );
  XNOR2_X1 U12489 ( .A(n12518), .B(n12519), .ZN(n12262) );
  XOR2_X1 U12490 ( .A(n12520), .B(n12521), .Z(n12518) );
  XNOR2_X1 U12491 ( .A(n12522), .B(n12523), .ZN(n12266) );
  XNOR2_X1 U12492 ( .A(n12524), .B(n12525), .ZN(n12523) );
  XOR2_X1 U12493 ( .A(n12526), .B(n12527), .Z(n12269) );
  XNOR2_X1 U12494 ( .A(n12528), .B(n12529), .ZN(n12526) );
  XNOR2_X1 U12495 ( .A(n12530), .B(n12531), .ZN(n12107) );
  NAND2_X1 U12496 ( .A1(n12532), .A2(n12533), .ZN(n12530) );
  XNOR2_X1 U12497 ( .A(n12534), .B(n12535), .ZN(n12273) );
  XOR2_X1 U12498 ( .A(n12536), .B(n12537), .Z(n12534) );
  NOR2_X1 U12499 ( .A1(n8572), .A2(n8578), .ZN(n12537) );
  XNOR2_X1 U12500 ( .A(n12538), .B(n12539), .ZN(n12278) );
  XNOR2_X1 U12501 ( .A(n12540), .B(n12541), .ZN(n12538) );
  NOR2_X1 U12502 ( .A1(n8556), .A2(n8578), .ZN(n12541) );
  XOR2_X1 U12503 ( .A(n12542), .B(n12543), .Z(n12281) );
  XNOR2_X1 U12504 ( .A(n12544), .B(n12545), .ZN(n12542) );
  NOR2_X1 U12505 ( .A1(n8594), .A2(n8578), .ZN(n12545) );
  XNOR2_X1 U12506 ( .A(n12546), .B(n12547), .ZN(n12286) );
  XNOR2_X1 U12507 ( .A(n12548), .B(n12549), .ZN(n12547) );
  NAND2_X1 U12508 ( .A1(n12196), .A2(n9295), .ZN(n12549) );
  XOR2_X1 U12509 ( .A(n12550), .B(n12551), .Z(n12289) );
  XOR2_X1 U12510 ( .A(n12552), .B(n12553), .Z(n12550) );
  NOR2_X1 U12511 ( .A1(n8544), .A2(n8578), .ZN(n12553) );
  XOR2_X1 U12512 ( .A(n12554), .B(n12555), .Z(n12294) );
  XNOR2_X1 U12513 ( .A(n12556), .B(n12557), .ZN(n12555) );
  NAND2_X1 U12514 ( .A1(n12196), .A2(n9286), .ZN(n12557) );
  XNOR2_X1 U12515 ( .A(n12558), .B(n12559), .ZN(n12298) );
  XNOR2_X1 U12516 ( .A(n12560), .B(n12561), .ZN(n12558) );
  NOR2_X1 U12517 ( .A1(n8564), .A2(n8578), .ZN(n12561) );
  XNOR2_X1 U12518 ( .A(n12562), .B(n12563), .ZN(n12302) );
  XNOR2_X1 U12519 ( .A(n12564), .B(n12565), .ZN(n12562) );
  NOR2_X1 U12520 ( .A1(n8528), .A2(n8578), .ZN(n12565) );
  XOR2_X1 U12521 ( .A(n12566), .B(n12567), .Z(n12306) );
  XNOR2_X1 U12522 ( .A(n12568), .B(n12569), .ZN(n12567) );
  NAND2_X1 U12523 ( .A1(n8911), .A2(n12570), .ZN(n8841) );
  NAND2_X1 U12524 ( .A1(n12571), .A2(n12572), .ZN(n12570) );
  INV_X1 U12525 ( .A(n12573), .ZN(n12572) );
  XOR2_X1 U12526 ( .A(n12574), .B(n12575), .Z(n12571) );
  INV_X1 U12527 ( .A(n12576), .ZN(n8845) );
  NOR2_X1 U12528 ( .A1(n8911), .A2(n8910), .ZN(n12576) );
  XNOR2_X1 U12529 ( .A(n12577), .B(n12578), .ZN(n8910) );
  NAND2_X1 U12530 ( .A1(n12579), .A2(n12573), .ZN(n8911) );
  NAND2_X1 U12531 ( .A1(n12580), .A2(n12581), .ZN(n12573) );
  NAND2_X1 U12532 ( .A1(n12320), .A2(n12582), .ZN(n12581) );
  NAND2_X1 U12533 ( .A1(n12317), .A2(n12319), .ZN(n12582) );
  NOR2_X1 U12534 ( .A1(n8578), .A2(n8972), .ZN(n12320) );
  INV_X1 U12535 ( .A(n12583), .ZN(n12580) );
  NOR2_X1 U12536 ( .A1(n12319), .A2(n12317), .ZN(n12583) );
  XNOR2_X1 U12537 ( .A(n12584), .B(n12585), .ZN(n12317) );
  XOR2_X1 U12538 ( .A(n12586), .B(n12587), .Z(n12584) );
  NOR2_X1 U12539 ( .A1(n8589), .A2(n8587), .ZN(n12587) );
  NAND2_X1 U12540 ( .A1(n12588), .A2(n12589), .ZN(n12319) );
  NAND2_X1 U12541 ( .A1(n12327), .A2(n12590), .ZN(n12589) );
  NAND2_X1 U12542 ( .A1(n12329), .A2(n12328), .ZN(n12590) );
  XOR2_X1 U12543 ( .A(n12591), .B(n12592), .Z(n12327) );
  XOR2_X1 U12544 ( .A(n12593), .B(n12594), .Z(n12591) );
  INV_X1 U12545 ( .A(n12595), .ZN(n12588) );
  NOR2_X1 U12546 ( .A1(n12328), .A2(n12329), .ZN(n12595) );
  NOR2_X1 U12547 ( .A1(n8578), .A2(n8589), .ZN(n12329) );
  NAND2_X1 U12548 ( .A1(n12596), .A2(n12597), .ZN(n12328) );
  NAND3_X1 U12549 ( .A1(n9268), .A2(n12598), .A3(n12196), .ZN(n12597) );
  NAND2_X1 U12550 ( .A1(n12335), .A2(n12336), .ZN(n12598) );
  INV_X1 U12551 ( .A(n12599), .ZN(n12596) );
  NOR2_X1 U12552 ( .A1(n12336), .A2(n12335), .ZN(n12599) );
  XOR2_X1 U12553 ( .A(n12600), .B(n12601), .Z(n12335) );
  NAND2_X1 U12554 ( .A1(n12602), .A2(n12603), .ZN(n12600) );
  NAND2_X1 U12555 ( .A1(n12604), .A2(n12605), .ZN(n12336) );
  NAND2_X1 U12556 ( .A1(n12566), .A2(n12606), .ZN(n12605) );
  NAND2_X1 U12557 ( .A1(n12569), .A2(n12568), .ZN(n12606) );
  XOR2_X1 U12558 ( .A(n12607), .B(n12608), .Z(n12566) );
  XOR2_X1 U12559 ( .A(n12609), .B(n12610), .Z(n12608) );
  NAND2_X1 U12560 ( .A1(n12457), .A2(n9277), .ZN(n12610) );
  INV_X1 U12561 ( .A(n12611), .ZN(n12604) );
  NOR2_X1 U12562 ( .A1(n12568), .A2(n12569), .ZN(n12611) );
  NOR2_X1 U12563 ( .A1(n8578), .A2(n8527), .ZN(n12569) );
  NAND2_X1 U12564 ( .A1(n12612), .A2(n12613), .ZN(n12568) );
  NAND3_X1 U12565 ( .A1(n9277), .A2(n12614), .A3(n12196), .ZN(n12613) );
  NAND2_X1 U12566 ( .A1(n12564), .A2(n12563), .ZN(n12614) );
  INV_X1 U12567 ( .A(n12615), .ZN(n12612) );
  NOR2_X1 U12568 ( .A1(n12563), .A2(n12564), .ZN(n12615) );
  NOR2_X1 U12569 ( .A1(n12616), .A2(n12617), .ZN(n12564) );
  INV_X1 U12570 ( .A(n12618), .ZN(n12617) );
  NAND3_X1 U12571 ( .A1(n10307), .A2(n12619), .A3(n12196), .ZN(n12618) );
  NAND2_X1 U12572 ( .A1(n12560), .A2(n12559), .ZN(n12619) );
  NOR2_X1 U12573 ( .A1(n12559), .A2(n12560), .ZN(n12616) );
  NOR2_X1 U12574 ( .A1(n12620), .A2(n12621), .ZN(n12560) );
  NOR3_X1 U12575 ( .A1(n9000), .A2(n12622), .A3(n8578), .ZN(n12621) );
  INV_X1 U12576 ( .A(n12623), .ZN(n12622) );
  NAND2_X1 U12577 ( .A1(n12556), .A2(n12554), .ZN(n12623) );
  NOR2_X1 U12578 ( .A1(n12554), .A2(n12556), .ZN(n12620) );
  NOR2_X1 U12579 ( .A1(n12624), .A2(n12625), .ZN(n12556) );
  NOR3_X1 U12580 ( .A1(n8544), .A2(n12626), .A3(n8578), .ZN(n12625) );
  NOR2_X1 U12581 ( .A1(n12552), .A2(n12551), .ZN(n12626) );
  INV_X1 U12582 ( .A(n12627), .ZN(n12624) );
  NAND2_X1 U12583 ( .A1(n12551), .A2(n12552), .ZN(n12627) );
  NAND2_X1 U12584 ( .A1(n12628), .A2(n12629), .ZN(n12552) );
  NAND3_X1 U12585 ( .A1(n9295), .A2(n12630), .A3(n12196), .ZN(n12629) );
  NAND2_X1 U12586 ( .A1(n12548), .A2(n12546), .ZN(n12630) );
  INV_X1 U12587 ( .A(n12631), .ZN(n12628) );
  NOR2_X1 U12588 ( .A1(n12546), .A2(n12548), .ZN(n12631) );
  NOR2_X1 U12589 ( .A1(n12632), .A2(n12633), .ZN(n12548) );
  INV_X1 U12590 ( .A(n12634), .ZN(n12633) );
  NAND3_X1 U12591 ( .A1(n10846), .A2(n12635), .A3(n12196), .ZN(n12634) );
  NAND2_X1 U12592 ( .A1(n12544), .A2(n12543), .ZN(n12635) );
  NOR2_X1 U12593 ( .A1(n12543), .A2(n12544), .ZN(n12632) );
  NOR2_X1 U12594 ( .A1(n12636), .A2(n12637), .ZN(n12544) );
  INV_X1 U12595 ( .A(n12638), .ZN(n12637) );
  NAND3_X1 U12596 ( .A1(n9304), .A2(n12639), .A3(n12196), .ZN(n12638) );
  NAND2_X1 U12597 ( .A1(n12540), .A2(n12539), .ZN(n12639) );
  NOR2_X1 U12598 ( .A1(n12539), .A2(n12540), .ZN(n12636) );
  NOR2_X1 U12599 ( .A1(n12640), .A2(n12641), .ZN(n12540) );
  NOR3_X1 U12600 ( .A1(n9025), .A2(n12642), .A3(n8578), .ZN(n12641) );
  NOR2_X1 U12601 ( .A1(n12536), .A2(n12535), .ZN(n12642) );
  INV_X1 U12602 ( .A(n12643), .ZN(n12640) );
  NAND2_X1 U12603 ( .A1(n12535), .A2(n12536), .ZN(n12643) );
  NAND2_X1 U12604 ( .A1(n12532), .A2(n12644), .ZN(n12536) );
  NAND2_X1 U12605 ( .A1(n12531), .A2(n12533), .ZN(n12644) );
  NAND2_X1 U12606 ( .A1(n12645), .A2(n12646), .ZN(n12533) );
  NAND2_X1 U12607 ( .A1(n12196), .A2(n9313), .ZN(n12646) );
  XOR2_X1 U12608 ( .A(n12647), .B(n12648), .Z(n12531) );
  XNOR2_X1 U12609 ( .A(n12649), .B(n12650), .ZN(n12648) );
  NAND2_X1 U12610 ( .A1(n9313), .A2(n12651), .ZN(n12532) );
  INV_X1 U12611 ( .A(n12645), .ZN(n12651) );
  NOR2_X1 U12612 ( .A1(n12652), .A2(n12653), .ZN(n12645) );
  INV_X1 U12613 ( .A(n12654), .ZN(n12653) );
  NAND2_X1 U12614 ( .A1(n12529), .A2(n12655), .ZN(n12654) );
  NAND2_X1 U12615 ( .A1(n12528), .A2(n12527), .ZN(n12655) );
  NOR2_X1 U12616 ( .A1(n8578), .A2(n8591), .ZN(n12529) );
  NOR2_X1 U12617 ( .A1(n12527), .A2(n12528), .ZN(n12652) );
  NOR2_X1 U12618 ( .A1(n12656), .A2(n12657), .ZN(n12528) );
  INV_X1 U12619 ( .A(n12658), .ZN(n12657) );
  NAND2_X1 U12620 ( .A1(n12525), .A2(n12659), .ZN(n12658) );
  NAND2_X1 U12621 ( .A1(n12660), .A2(n12522), .ZN(n12659) );
  NOR2_X1 U12622 ( .A1(n8578), .A2(n8562), .ZN(n12525) );
  NOR2_X1 U12623 ( .A1(n12522), .A2(n12660), .ZN(n12656) );
  INV_X1 U12624 ( .A(n12524), .ZN(n12660) );
  NAND2_X1 U12625 ( .A1(n12661), .A2(n12662), .ZN(n12524) );
  NAND2_X1 U12626 ( .A1(n12521), .A2(n12663), .ZN(n12662) );
  INV_X1 U12627 ( .A(n12664), .ZN(n12663) );
  NOR2_X1 U12628 ( .A1(n12520), .A2(n12519), .ZN(n12664) );
  NOR2_X1 U12629 ( .A1(n8578), .A2(n8545), .ZN(n12521) );
  NAND2_X1 U12630 ( .A1(n12519), .A2(n12520), .ZN(n12661) );
  NAND2_X1 U12631 ( .A1(n12665), .A2(n12666), .ZN(n12520) );
  NAND2_X1 U12632 ( .A1(n12517), .A2(n12667), .ZN(n12666) );
  INV_X1 U12633 ( .A(n12668), .ZN(n12667) );
  NOR2_X1 U12634 ( .A1(n12516), .A2(n12514), .ZN(n12668) );
  NOR2_X1 U12635 ( .A1(n8578), .A2(n8569), .ZN(n12517) );
  NAND2_X1 U12636 ( .A1(n12514), .A2(n12516), .ZN(n12665) );
  NAND2_X1 U12637 ( .A1(n12669), .A2(n12670), .ZN(n12516) );
  NAND2_X1 U12638 ( .A1(n12513), .A2(n12671), .ZN(n12670) );
  INV_X1 U12639 ( .A(n12672), .ZN(n12671) );
  NOR2_X1 U12640 ( .A1(n12512), .A2(n12511), .ZN(n12672) );
  NOR2_X1 U12641 ( .A1(n8578), .A2(n8593), .ZN(n12513) );
  NAND2_X1 U12642 ( .A1(n12511), .A2(n12512), .ZN(n12669) );
  NAND2_X1 U12643 ( .A1(n12673), .A2(n12674), .ZN(n12512) );
  NAND2_X1 U12644 ( .A1(n12509), .A2(n12675), .ZN(n12674) );
  NAND2_X1 U12645 ( .A1(n12508), .A2(n12506), .ZN(n12675) );
  NOR2_X1 U12646 ( .A1(n8578), .A2(n8583), .ZN(n12509) );
  INV_X1 U12647 ( .A(n12676), .ZN(n12673) );
  NOR2_X1 U12648 ( .A1(n12506), .A2(n12508), .ZN(n12676) );
  NOR2_X1 U12649 ( .A1(n12677), .A2(n12678), .ZN(n12508) );
  INV_X1 U12650 ( .A(n12679), .ZN(n12678) );
  NAND2_X1 U12651 ( .A1(n12505), .A2(n12680), .ZN(n12679) );
  NAND2_X1 U12652 ( .A1(n12504), .A2(n12503), .ZN(n12680) );
  NOR2_X1 U12653 ( .A1(n8578), .A2(n8580), .ZN(n12505) );
  NOR2_X1 U12654 ( .A1(n12503), .A2(n12504), .ZN(n12677) );
  INV_X1 U12655 ( .A(n12681), .ZN(n12504) );
  NAND2_X1 U12656 ( .A1(n12682), .A2(n12683), .ZN(n12681) );
  NAND2_X1 U12657 ( .A1(n12500), .A2(n12684), .ZN(n12683) );
  INV_X1 U12658 ( .A(n12685), .ZN(n12684) );
  NOR2_X1 U12659 ( .A1(n12501), .A2(n12499), .ZN(n12685) );
  NOR2_X1 U12660 ( .A1(n8578), .A2(n8588), .ZN(n12500) );
  NAND2_X1 U12661 ( .A1(n12499), .A2(n12501), .ZN(n12682) );
  NAND2_X1 U12662 ( .A1(n12686), .A2(n12687), .ZN(n12501) );
  NAND2_X1 U12663 ( .A1(n12497), .A2(n12688), .ZN(n12687) );
  INV_X1 U12664 ( .A(n12689), .ZN(n12688) );
  NOR2_X1 U12665 ( .A1(n12496), .A2(n12495), .ZN(n12689) );
  NOR2_X1 U12666 ( .A1(n8578), .A2(n8551), .ZN(n12497) );
  NAND2_X1 U12667 ( .A1(n12495), .A2(n12496), .ZN(n12686) );
  NAND2_X1 U12668 ( .A1(n12690), .A2(n12691), .ZN(n12496) );
  NAND2_X1 U12669 ( .A1(n12493), .A2(n12692), .ZN(n12691) );
  NAND2_X1 U12670 ( .A1(n12492), .A2(n12490), .ZN(n12692) );
  NOR2_X1 U12671 ( .A1(n8578), .A2(n8563), .ZN(n12493) );
  INV_X1 U12672 ( .A(n12693), .ZN(n12690) );
  NOR2_X1 U12673 ( .A1(n12490), .A2(n12492), .ZN(n12693) );
  NOR2_X1 U12674 ( .A1(n12694), .A2(n12695), .ZN(n12492) );
  INV_X1 U12675 ( .A(n12696), .ZN(n12695) );
  NAND2_X1 U12676 ( .A1(n12489), .A2(n12697), .ZN(n12696) );
  NAND2_X1 U12677 ( .A1(n12488), .A2(n12487), .ZN(n12697) );
  NOR2_X1 U12678 ( .A1(n12195), .A2(n8548), .ZN(n12489) );
  NOR2_X1 U12679 ( .A1(n12487), .A2(n12488), .ZN(n12694) );
  NOR2_X1 U12680 ( .A1(n12698), .A2(n12699), .ZN(n12488) );
  INV_X1 U12681 ( .A(n12700), .ZN(n12699) );
  NAND2_X1 U12682 ( .A1(n12485), .A2(n12701), .ZN(n12700) );
  NAND2_X1 U12683 ( .A1(n12484), .A2(n12483), .ZN(n12701) );
  NOR2_X1 U12684 ( .A1(n12195), .A2(n8584), .ZN(n12485) );
  NOR2_X1 U12685 ( .A1(n12483), .A2(n12484), .ZN(n12698) );
  NOR2_X1 U12686 ( .A1(n12702), .A2(n12703), .ZN(n12484) );
  INV_X1 U12687 ( .A(n12704), .ZN(n12703) );
  NAND2_X1 U12688 ( .A1(n12480), .A2(n12705), .ZN(n12704) );
  NAND2_X1 U12689 ( .A1(n12481), .A2(n12479), .ZN(n12705) );
  NOR2_X1 U12690 ( .A1(n12195), .A2(n8535), .ZN(n12480) );
  NOR2_X1 U12691 ( .A1(n12479), .A2(n12481), .ZN(n12702) );
  NOR2_X1 U12692 ( .A1(n12706), .A2(n12707), .ZN(n12481) );
  INV_X1 U12693 ( .A(n12708), .ZN(n12707) );
  NAND2_X1 U12694 ( .A1(n12476), .A2(n12709), .ZN(n12708) );
  NAND2_X1 U12695 ( .A1(n12477), .A2(n12475), .ZN(n12709) );
  NOR2_X1 U12696 ( .A1(n12195), .A2(n8568), .ZN(n12476) );
  NOR2_X1 U12697 ( .A1(n12475), .A2(n12477), .ZN(n12706) );
  NOR2_X1 U12698 ( .A1(n12710), .A2(n12711), .ZN(n12477) );
  INV_X1 U12699 ( .A(n12712), .ZN(n12711) );
  NAND2_X1 U12700 ( .A1(n12472), .A2(n12713), .ZN(n12712) );
  NAND2_X1 U12701 ( .A1(n12473), .A2(n12471), .ZN(n12713) );
  NOR2_X1 U12702 ( .A1(n12195), .A2(n8574), .ZN(n12472) );
  NOR2_X1 U12703 ( .A1(n12471), .A2(n12473), .ZN(n12710) );
  NOR2_X1 U12704 ( .A1(n12714), .A2(n12715), .ZN(n12473) );
  INV_X1 U12705 ( .A(n12716), .ZN(n12715) );
  NAND2_X1 U12706 ( .A1(n12468), .A2(n12717), .ZN(n12716) );
  NAND2_X1 U12707 ( .A1(n12469), .A2(n12467), .ZN(n12717) );
  NOR2_X1 U12708 ( .A1(n12195), .A2(n8565), .ZN(n12468) );
  NOR2_X1 U12709 ( .A1(n12467), .A2(n12469), .ZN(n12714) );
  NOR2_X1 U12710 ( .A1(n12718), .A2(n12719), .ZN(n12469) );
  INV_X1 U12711 ( .A(n12720), .ZN(n12719) );
  NAND2_X1 U12712 ( .A1(n12462), .A2(n12721), .ZN(n12720) );
  NAND2_X1 U12713 ( .A1(n12465), .A2(n12464), .ZN(n12721) );
  NOR2_X1 U12714 ( .A1(n12195), .A2(n8567), .ZN(n12462) );
  NOR2_X1 U12715 ( .A1(n12464), .A2(n12465), .ZN(n12718) );
  INV_X1 U12716 ( .A(n12722), .ZN(n12465) );
  NAND2_X1 U12717 ( .A1(n12723), .A2(n12724), .ZN(n12722) );
  NAND2_X1 U12718 ( .A1(n12457), .A2(n12725), .ZN(n12724) );
  NAND2_X1 U12719 ( .A1(n8624), .A2(n12726), .ZN(n12725) );
  NAND2_X1 U12720 ( .A1(n8557), .A2(n8585), .ZN(n12726) );
  NAND2_X1 U12721 ( .A1(n12728), .A2(n12729), .ZN(n12723) );
  NAND2_X1 U12722 ( .A1(n8630), .A2(n12730), .ZN(n12729) );
  NAND2_X1 U12723 ( .A1(n8539), .A2(n8587), .ZN(n12730) );
  NAND3_X1 U12724 ( .A1(n12196), .A2(n8537), .A3(n12457), .ZN(n12464) );
  INV_X1 U12725 ( .A(n12195), .ZN(n12196) );
  XNOR2_X1 U12726 ( .A(n12731), .B(n12732), .ZN(n12195) );
  XOR2_X1 U12727 ( .A(d_17_), .B(c_17_), .Z(n12732) );
  XOR2_X1 U12728 ( .A(n12733), .B(n12734), .Z(n12467) );
  XNOR2_X1 U12729 ( .A(n12735), .B(n12736), .ZN(n12734) );
  XOR2_X1 U12730 ( .A(n12737), .B(n12738), .Z(n12471) );
  XNOR2_X1 U12731 ( .A(n12739), .B(n12740), .ZN(n12737) );
  XOR2_X1 U12732 ( .A(n12741), .B(n12742), .Z(n12475) );
  XNOR2_X1 U12733 ( .A(n12743), .B(n12744), .ZN(n12741) );
  XOR2_X1 U12734 ( .A(n12745), .B(n12746), .Z(n12479) );
  XNOR2_X1 U12735 ( .A(n12747), .B(n12748), .ZN(n12745) );
  XOR2_X1 U12736 ( .A(n12749), .B(n12750), .Z(n12483) );
  XNOR2_X1 U12737 ( .A(n12751), .B(n12752), .ZN(n12749) );
  NOR2_X1 U12738 ( .A1(n8535), .A2(n8587), .ZN(n12752) );
  XOR2_X1 U12739 ( .A(n12753), .B(n12754), .Z(n12487) );
  XNOR2_X1 U12740 ( .A(n12755), .B(n12756), .ZN(n12753) );
  NOR2_X1 U12741 ( .A1(n8584), .A2(n8587), .ZN(n12756) );
  XOR2_X1 U12742 ( .A(n12757), .B(n12758), .Z(n12490) );
  XNOR2_X1 U12743 ( .A(n12759), .B(n12760), .ZN(n12757) );
  NOR2_X1 U12744 ( .A1(n8548), .A2(n8587), .ZN(n12760) );
  XNOR2_X1 U12745 ( .A(n12761), .B(n12762), .ZN(n12495) );
  XNOR2_X1 U12746 ( .A(n12763), .B(n12764), .ZN(n12761) );
  NOR2_X1 U12747 ( .A1(n9094), .A2(n8587), .ZN(n12764) );
  XNOR2_X1 U12748 ( .A(n12765), .B(n12766), .ZN(n12499) );
  XNOR2_X1 U12749 ( .A(n12767), .B(n12768), .ZN(n12765) );
  NOR2_X1 U12750 ( .A1(n8551), .A2(n8587), .ZN(n12768) );
  XOR2_X1 U12751 ( .A(n12769), .B(n12770), .Z(n12503) );
  XNOR2_X1 U12752 ( .A(n12771), .B(n12772), .ZN(n12769) );
  NOR2_X1 U12753 ( .A1(n8588), .A2(n8587), .ZN(n12772) );
  XOR2_X1 U12754 ( .A(n12773), .B(n12774), .Z(n12506) );
  XNOR2_X1 U12755 ( .A(n12775), .B(n12776), .ZN(n12773) );
  NOR2_X1 U12756 ( .A1(n8580), .A2(n8587), .ZN(n12776) );
  XNOR2_X1 U12757 ( .A(n12777), .B(n12778), .ZN(n12511) );
  XNOR2_X1 U12758 ( .A(n12779), .B(n12780), .ZN(n12777) );
  NOR2_X1 U12759 ( .A1(n8583), .A2(n8587), .ZN(n12780) );
  XNOR2_X1 U12760 ( .A(n12781), .B(n12782), .ZN(n12514) );
  XNOR2_X1 U12761 ( .A(n12783), .B(n12784), .ZN(n12781) );
  NOR2_X1 U12762 ( .A1(n8593), .A2(n8587), .ZN(n12784) );
  XNOR2_X1 U12763 ( .A(n12785), .B(n12786), .ZN(n12519) );
  XNOR2_X1 U12764 ( .A(n12787), .B(n12788), .ZN(n12785) );
  NOR2_X1 U12765 ( .A1(n9050), .A2(n8587), .ZN(n12788) );
  XOR2_X1 U12766 ( .A(n12789), .B(n12790), .Z(n12522) );
  XNOR2_X1 U12767 ( .A(n12791), .B(n12792), .ZN(n12789) );
  NOR2_X1 U12768 ( .A1(n8545), .A2(n8587), .ZN(n12792) );
  XOR2_X1 U12769 ( .A(n12793), .B(n12794), .Z(n12527) );
  XNOR2_X1 U12770 ( .A(n12795), .B(n12796), .ZN(n12793) );
  NOR2_X1 U12771 ( .A1(n9041), .A2(n8587), .ZN(n12796) );
  XOR2_X1 U12772 ( .A(n12797), .B(n12798), .Z(n12535) );
  XOR2_X1 U12773 ( .A(n12799), .B(n12800), .Z(n12797) );
  XOR2_X1 U12774 ( .A(n12801), .B(n12802), .Z(n12539) );
  XNOR2_X1 U12775 ( .A(n12803), .B(n12804), .ZN(n12801) );
  XNOR2_X1 U12776 ( .A(n12805), .B(n12806), .ZN(n12543) );
  XOR2_X1 U12777 ( .A(n12807), .B(n12808), .Z(n12806) );
  XOR2_X1 U12778 ( .A(n12809), .B(n12810), .Z(n12546) );
  XNOR2_X1 U12779 ( .A(n12811), .B(n12812), .ZN(n12809) );
  XNOR2_X1 U12780 ( .A(n12813), .B(n12814), .ZN(n12551) );
  XNOR2_X1 U12781 ( .A(n12815), .B(n12816), .ZN(n12813) );
  XOR2_X1 U12782 ( .A(n12817), .B(n12818), .Z(n12554) );
  XNOR2_X1 U12783 ( .A(n12819), .B(n12820), .ZN(n12817) );
  XNOR2_X1 U12784 ( .A(n12821), .B(n12822), .ZN(n12559) );
  XOR2_X1 U12785 ( .A(n12823), .B(n12824), .Z(n12821) );
  NOR2_X1 U12786 ( .A1(n8555), .A2(n8587), .ZN(n12824) );
  XOR2_X1 U12787 ( .A(n12825), .B(n12826), .Z(n12563) );
  NAND2_X1 U12788 ( .A1(n12827), .A2(n12828), .ZN(n12825) );
  XNOR2_X1 U12789 ( .A(n12574), .B(n12575), .ZN(n12579) );
  NAND2_X1 U12790 ( .A1(n12829), .A2(n12830), .ZN(n12574) );
  NAND2_X1 U12791 ( .A1(n12831), .A2(n12832), .ZN(n8848) );
  NAND2_X1 U12792 ( .A1(n12833), .A2(n12834), .ZN(n12832) );
  NAND2_X1 U12793 ( .A1(n12577), .A2(n12578), .ZN(n12831) );
  NAND4_X1 U12794 ( .A1(n12577), .A2(n12833), .A3(n12578), .A4(n12834), .ZN(
        n8849) );
  INV_X1 U12795 ( .A(n8906), .ZN(n12834) );
  NAND2_X1 U12796 ( .A1(n12829), .A2(n12835), .ZN(n12578) );
  NAND2_X1 U12797 ( .A1(n12575), .A2(n12830), .ZN(n12835) );
  NAND2_X1 U12798 ( .A1(n12836), .A2(n12837), .ZN(n12830) );
  NAND2_X1 U12799 ( .A1(n12457), .A2(n8872), .ZN(n12837) );
  XOR2_X1 U12800 ( .A(n12838), .B(n12839), .Z(n12575) );
  XOR2_X1 U12801 ( .A(n12840), .B(n12841), .Z(n12838) );
  NOR2_X1 U12802 ( .A1(n8589), .A2(n8557), .ZN(n12841) );
  NAND2_X1 U12803 ( .A1(n8592), .A2(n12842), .ZN(n12829) );
  INV_X1 U12804 ( .A(n12836), .ZN(n12842) );
  NOR2_X1 U12805 ( .A1(n12843), .A2(n12844), .ZN(n12836) );
  NOR3_X1 U12806 ( .A1(n8884), .A2(n12845), .A3(n8587), .ZN(n12844) );
  INV_X1 U12807 ( .A(n12846), .ZN(n12845) );
  NAND2_X1 U12808 ( .A1(n12585), .A2(n12586), .ZN(n12846) );
  NOR2_X1 U12809 ( .A1(n12585), .A2(n12586), .ZN(n12843) );
  NAND2_X1 U12810 ( .A1(n12847), .A2(n12848), .ZN(n12586) );
  NAND2_X1 U12811 ( .A1(n12592), .A2(n12849), .ZN(n12848) );
  NAND2_X1 U12812 ( .A1(n12594), .A2(n12593), .ZN(n12849) );
  XNOR2_X1 U12813 ( .A(n12850), .B(n12851), .ZN(n12592) );
  XOR2_X1 U12814 ( .A(n12852), .B(n12853), .Z(n12850) );
  NOR2_X1 U12815 ( .A1(n8527), .A2(n8557), .ZN(n12853) );
  INV_X1 U12816 ( .A(n12854), .ZN(n12847) );
  NOR2_X1 U12817 ( .A1(n12593), .A2(n12594), .ZN(n12854) );
  NOR2_X1 U12818 ( .A1(n8587), .A2(n8552), .ZN(n12594) );
  NAND2_X1 U12819 ( .A1(n12602), .A2(n12855), .ZN(n12593) );
  NAND2_X1 U12820 ( .A1(n12601), .A2(n12603), .ZN(n12855) );
  NAND2_X1 U12821 ( .A1(n12856), .A2(n12857), .ZN(n12603) );
  NAND2_X1 U12822 ( .A1(n12457), .A2(n9792), .ZN(n12857) );
  INV_X1 U12823 ( .A(n12858), .ZN(n12856) );
  XNOR2_X1 U12824 ( .A(n12859), .B(n12860), .ZN(n12601) );
  XOR2_X1 U12825 ( .A(n12861), .B(n12862), .Z(n12860) );
  NAND2_X1 U12826 ( .A1(n12728), .A2(n9277), .ZN(n12862) );
  NAND2_X1 U12827 ( .A1(n9792), .A2(n12858), .ZN(n12602) );
  NAND2_X1 U12828 ( .A1(n12863), .A2(n12864), .ZN(n12858) );
  INV_X1 U12829 ( .A(n12865), .ZN(n12864) );
  NOR3_X1 U12830 ( .A1(n8528), .A2(n12866), .A3(n8587), .ZN(n12865) );
  NOR2_X1 U12831 ( .A1(n12607), .A2(n12609), .ZN(n12866) );
  NAND2_X1 U12832 ( .A1(n12607), .A2(n12609), .ZN(n12863) );
  NAND2_X1 U12833 ( .A1(n12827), .A2(n12867), .ZN(n12609) );
  NAND2_X1 U12834 ( .A1(n12826), .A2(n12828), .ZN(n12867) );
  NAND2_X1 U12835 ( .A1(n12868), .A2(n12869), .ZN(n12828) );
  NAND2_X1 U12836 ( .A1(n12457), .A2(n10307), .ZN(n12869) );
  INV_X1 U12837 ( .A(n12870), .ZN(n12868) );
  XOR2_X1 U12838 ( .A(n12871), .B(n12872), .Z(n12826) );
  XNOR2_X1 U12839 ( .A(n12873), .B(n12874), .ZN(n12872) );
  NAND2_X1 U12840 ( .A1(n12728), .A2(n9286), .ZN(n12874) );
  NAND2_X1 U12841 ( .A1(n10307), .A2(n12870), .ZN(n12827) );
  NAND2_X1 U12842 ( .A1(n12875), .A2(n12876), .ZN(n12870) );
  INV_X1 U12843 ( .A(n12877), .ZN(n12876) );
  NOR3_X1 U12844 ( .A1(n9000), .A2(n12878), .A3(n8587), .ZN(n12877) );
  NOR2_X1 U12845 ( .A1(n12822), .A2(n12823), .ZN(n12878) );
  NAND2_X1 U12846 ( .A1(n12822), .A2(n12823), .ZN(n12875) );
  NAND2_X1 U12847 ( .A1(n12879), .A2(n12880), .ZN(n12823) );
  NAND2_X1 U12848 ( .A1(n12820), .A2(n12881), .ZN(n12880) );
  NAND2_X1 U12849 ( .A1(n12818), .A2(n12819), .ZN(n12881) );
  NOR2_X1 U12850 ( .A1(n8587), .A2(n8544), .ZN(n12820) );
  INV_X1 U12851 ( .A(n12882), .ZN(n12879) );
  NOR2_X1 U12852 ( .A1(n12818), .A2(n12819), .ZN(n12882) );
  NOR2_X1 U12853 ( .A1(n12883), .A2(n12884), .ZN(n12819) );
  INV_X1 U12854 ( .A(n12885), .ZN(n12884) );
  NAND2_X1 U12855 ( .A1(n12815), .A2(n12886), .ZN(n12885) );
  NAND2_X1 U12856 ( .A1(n12816), .A2(n12814), .ZN(n12886) );
  NOR2_X1 U12857 ( .A1(n12456), .A2(n8560), .ZN(n12815) );
  NOR2_X1 U12858 ( .A1(n12814), .A2(n12816), .ZN(n12883) );
  NOR2_X1 U12859 ( .A1(n12887), .A2(n12888), .ZN(n12816) );
  INV_X1 U12860 ( .A(n12889), .ZN(n12888) );
  NAND2_X1 U12861 ( .A1(n12812), .A2(n12890), .ZN(n12889) );
  NAND2_X1 U12862 ( .A1(n12811), .A2(n12810), .ZN(n12890) );
  NOR2_X1 U12863 ( .A1(n12456), .A2(n8594), .ZN(n12812) );
  NOR2_X1 U12864 ( .A1(n12810), .A2(n12811), .ZN(n12887) );
  NOR2_X1 U12865 ( .A1(n12891), .A2(n12892), .ZN(n12811) );
  INV_X1 U12866 ( .A(n12893), .ZN(n12892) );
  NAND2_X1 U12867 ( .A1(n12808), .A2(n12894), .ZN(n12893) );
  NAND2_X1 U12868 ( .A1(n12807), .A2(n12805), .ZN(n12894) );
  NOR2_X1 U12869 ( .A1(n12456), .A2(n8556), .ZN(n12808) );
  NOR2_X1 U12870 ( .A1(n12805), .A2(n12807), .ZN(n12891) );
  NOR2_X1 U12871 ( .A1(n12895), .A2(n12896), .ZN(n12807) );
  INV_X1 U12872 ( .A(n12897), .ZN(n12896) );
  NAND2_X1 U12873 ( .A1(n12804), .A2(n12898), .ZN(n12897) );
  NAND2_X1 U12874 ( .A1(n12802), .A2(n12803), .ZN(n12898) );
  NOR2_X1 U12875 ( .A1(n12456), .A2(n8572), .ZN(n12804) );
  NOR2_X1 U12876 ( .A1(n12802), .A2(n12803), .ZN(n12895) );
  NOR2_X1 U12877 ( .A1(n12899), .A2(n12900), .ZN(n12803) );
  INV_X1 U12878 ( .A(n12901), .ZN(n12900) );
  NAND2_X1 U12879 ( .A1(n12800), .A2(n12902), .ZN(n12901) );
  NAND2_X1 U12880 ( .A1(n12798), .A2(n12799), .ZN(n12902) );
  NOR2_X1 U12881 ( .A1(n12456), .A2(n8582), .ZN(n12800) );
  NOR2_X1 U12882 ( .A1(n12798), .A2(n12799), .ZN(n12899) );
  NAND2_X1 U12883 ( .A1(n12903), .A2(n12904), .ZN(n12799) );
  NAND2_X1 U12884 ( .A1(n12647), .A2(n12905), .ZN(n12904) );
  INV_X1 U12885 ( .A(n12906), .ZN(n12905) );
  NOR2_X1 U12886 ( .A1(n12650), .A2(n12649), .ZN(n12906) );
  XOR2_X1 U12887 ( .A(n12907), .B(n12908), .Z(n12647) );
  NAND2_X1 U12888 ( .A1(n12909), .A2(n12910), .ZN(n12907) );
  NAND2_X1 U12889 ( .A1(n12649), .A2(n12650), .ZN(n12903) );
  NAND2_X1 U12890 ( .A1(n12457), .A2(n9721), .ZN(n12650) );
  NOR2_X1 U12891 ( .A1(n12911), .A2(n12912), .ZN(n12649) );
  INV_X1 U12892 ( .A(n12913), .ZN(n12912) );
  NAND3_X1 U12893 ( .A1(n9322), .A2(n12914), .A3(n12457), .ZN(n12913) );
  NAND2_X1 U12894 ( .A1(n12794), .A2(n12795), .ZN(n12914) );
  NOR2_X1 U12895 ( .A1(n12794), .A2(n12795), .ZN(n12911) );
  NOR2_X1 U12896 ( .A1(n12915), .A2(n12916), .ZN(n12795) );
  INV_X1 U12897 ( .A(n12917), .ZN(n12916) );
  NAND3_X1 U12898 ( .A1(n10222), .A2(n12918), .A3(n12457), .ZN(n12917) );
  NAND2_X1 U12899 ( .A1(n12790), .A2(n12791), .ZN(n12918) );
  NOR2_X1 U12900 ( .A1(n12790), .A2(n12791), .ZN(n12915) );
  NOR2_X1 U12901 ( .A1(n12919), .A2(n12920), .ZN(n12791) );
  INV_X1 U12902 ( .A(n12921), .ZN(n12920) );
  NAND3_X1 U12903 ( .A1(n9331), .A2(n12922), .A3(n12457), .ZN(n12921) );
  NAND2_X1 U12904 ( .A1(n12787), .A2(n12786), .ZN(n12922) );
  NOR2_X1 U12905 ( .A1(n12786), .A2(n12787), .ZN(n12919) );
  NOR2_X1 U12906 ( .A1(n12923), .A2(n12924), .ZN(n12787) );
  NOR3_X1 U12907 ( .A1(n9056), .A2(n12925), .A3(n8587), .ZN(n12924) );
  INV_X1 U12908 ( .A(n12926), .ZN(n12925) );
  NAND2_X1 U12909 ( .A1(n12782), .A2(n12783), .ZN(n12926) );
  NOR2_X1 U12910 ( .A1(n12782), .A2(n12783), .ZN(n12923) );
  NOR2_X1 U12911 ( .A1(n12927), .A2(n12928), .ZN(n12783) );
  INV_X1 U12912 ( .A(n12929), .ZN(n12928) );
  NAND3_X1 U12913 ( .A1(n9340), .A2(n12930), .A3(n12457), .ZN(n12929) );
  NAND2_X1 U12914 ( .A1(n12779), .A2(n12778), .ZN(n12930) );
  NOR2_X1 U12915 ( .A1(n12778), .A2(n12779), .ZN(n12927) );
  NOR2_X1 U12916 ( .A1(n12931), .A2(n12932), .ZN(n12779) );
  NOR3_X1 U12917 ( .A1(n9066), .A2(n12933), .A3(n8587), .ZN(n12932) );
  INV_X1 U12918 ( .A(n12934), .ZN(n12933) );
  NAND2_X1 U12919 ( .A1(n12774), .A2(n12775), .ZN(n12934) );
  NOR2_X1 U12920 ( .A1(n12774), .A2(n12775), .ZN(n12931) );
  NOR2_X1 U12921 ( .A1(n12935), .A2(n12936), .ZN(n12775) );
  INV_X1 U12922 ( .A(n12937), .ZN(n12936) );
  NAND3_X1 U12923 ( .A1(n9080), .A2(n12938), .A3(n12457), .ZN(n12937) );
  NAND2_X1 U12924 ( .A1(n12771), .A2(n12770), .ZN(n12938) );
  NOR2_X1 U12925 ( .A1(n12770), .A2(n12771), .ZN(n12935) );
  NOR2_X1 U12926 ( .A1(n12939), .A2(n12940), .ZN(n12771) );
  NOR3_X1 U12927 ( .A1(n8551), .A2(n12941), .A3(n8587), .ZN(n12940) );
  INV_X1 U12928 ( .A(n12942), .ZN(n12941) );
  NAND2_X1 U12929 ( .A1(n12766), .A2(n12767), .ZN(n12942) );
  NOR2_X1 U12930 ( .A1(n12766), .A2(n12767), .ZN(n12939) );
  NOR2_X1 U12931 ( .A1(n12943), .A2(n12944), .ZN(n12767) );
  INV_X1 U12932 ( .A(n12945), .ZN(n12944) );
  NAND3_X1 U12933 ( .A1(n9098), .A2(n12946), .A3(n12457), .ZN(n12945) );
  NAND2_X1 U12934 ( .A1(n12763), .A2(n12762), .ZN(n12946) );
  NOR2_X1 U12935 ( .A1(n12762), .A2(n12763), .ZN(n12943) );
  NOR2_X1 U12936 ( .A1(n12947), .A2(n12948), .ZN(n12763) );
  NOR3_X1 U12937 ( .A1(n8548), .A2(n12949), .A3(n8587), .ZN(n12948) );
  INV_X1 U12938 ( .A(n12950), .ZN(n12949) );
  NAND2_X1 U12939 ( .A1(n12758), .A2(n12759), .ZN(n12950) );
  NOR2_X1 U12940 ( .A1(n12758), .A2(n12759), .ZN(n12947) );
  NOR2_X1 U12941 ( .A1(n12951), .A2(n12952), .ZN(n12759) );
  INV_X1 U12942 ( .A(n12953), .ZN(n12952) );
  NAND3_X1 U12943 ( .A1(n9112), .A2(n12954), .A3(n12457), .ZN(n12953) );
  NAND2_X1 U12944 ( .A1(n12755), .A2(n12754), .ZN(n12954) );
  NOR2_X1 U12945 ( .A1(n12754), .A2(n12755), .ZN(n12951) );
  NOR2_X1 U12946 ( .A1(n12955), .A2(n12956), .ZN(n12755) );
  INV_X1 U12947 ( .A(n12957), .ZN(n12956) );
  NAND3_X1 U12948 ( .A1(n9121), .A2(n12958), .A3(n12457), .ZN(n12957) );
  NAND2_X1 U12949 ( .A1(n12750), .A2(n12751), .ZN(n12958) );
  NOR2_X1 U12950 ( .A1(n12750), .A2(n12751), .ZN(n12955) );
  NOR2_X1 U12951 ( .A1(n12959), .A2(n12960), .ZN(n12751) );
  INV_X1 U12952 ( .A(n12961), .ZN(n12960) );
  NAND2_X1 U12953 ( .A1(n12748), .A2(n12962), .ZN(n12961) );
  NAND2_X1 U12954 ( .A1(n12747), .A2(n12746), .ZN(n12962) );
  NOR2_X1 U12955 ( .A1(n12456), .A2(n8568), .ZN(n12748) );
  NOR2_X1 U12956 ( .A1(n12746), .A2(n12747), .ZN(n12959) );
  NOR2_X1 U12957 ( .A1(n12963), .A2(n12964), .ZN(n12747) );
  INV_X1 U12958 ( .A(n12965), .ZN(n12964) );
  NAND2_X1 U12959 ( .A1(n12743), .A2(n12966), .ZN(n12965) );
  NAND2_X1 U12960 ( .A1(n12742), .A2(n12744), .ZN(n12966) );
  NOR2_X1 U12961 ( .A1(n12456), .A2(n8574), .ZN(n12743) );
  NOR2_X1 U12962 ( .A1(n12742), .A2(n12744), .ZN(n12963) );
  NOR2_X1 U12963 ( .A1(n12967), .A2(n12968), .ZN(n12744) );
  INV_X1 U12964 ( .A(n12969), .ZN(n12968) );
  NAND2_X1 U12965 ( .A1(n12739), .A2(n12970), .ZN(n12969) );
  NAND2_X1 U12966 ( .A1(n12740), .A2(n12738), .ZN(n12970) );
  NOR2_X1 U12967 ( .A1(n12456), .A2(n8565), .ZN(n12739) );
  NOR2_X1 U12968 ( .A1(n12738), .A2(n12740), .ZN(n12967) );
  NOR2_X1 U12969 ( .A1(n12971), .A2(n12972), .ZN(n12740) );
  INV_X1 U12970 ( .A(n12973), .ZN(n12972) );
  NAND2_X1 U12971 ( .A1(n12733), .A2(n12974), .ZN(n12973) );
  NAND2_X1 U12972 ( .A1(n12736), .A2(n12735), .ZN(n12974) );
  NOR2_X1 U12973 ( .A1(n12456), .A2(n8567), .ZN(n12733) );
  NOR2_X1 U12974 ( .A1(n12735), .A2(n12736), .ZN(n12971) );
  INV_X1 U12975 ( .A(n12975), .ZN(n12736) );
  NAND2_X1 U12976 ( .A1(n12976), .A2(n12977), .ZN(n12975) );
  NAND2_X1 U12977 ( .A1(n12728), .A2(n12978), .ZN(n12977) );
  NAND2_X1 U12978 ( .A1(n8624), .A2(n12979), .ZN(n12978) );
  NAND2_X1 U12979 ( .A1(n8570), .A2(n8585), .ZN(n12979) );
  NAND2_X1 U12980 ( .A1(n12981), .A2(n12982), .ZN(n12976) );
  NAND2_X1 U12981 ( .A1(n8630), .A2(n12983), .ZN(n12982) );
  NAND2_X1 U12982 ( .A1(n8539), .A2(n8557), .ZN(n12983) );
  NAND3_X1 U12983 ( .A1(n12728), .A2(n8537), .A3(n12457), .ZN(n12735) );
  INV_X1 U12984 ( .A(n12456), .ZN(n12457) );
  XNOR2_X1 U12985 ( .A(n12984), .B(n12985), .ZN(n12456) );
  XOR2_X1 U12986 ( .A(d_16_), .B(c_16_), .Z(n12985) );
  XOR2_X1 U12987 ( .A(n12986), .B(n12987), .Z(n12738) );
  XNOR2_X1 U12988 ( .A(n12988), .B(n12989), .ZN(n12987) );
  XOR2_X1 U12989 ( .A(n12990), .B(n12991), .Z(n12742) );
  XNOR2_X1 U12990 ( .A(n12992), .B(n12993), .ZN(n12990) );
  XOR2_X1 U12991 ( .A(n12994), .B(n12995), .Z(n12746) );
  XNOR2_X1 U12992 ( .A(n12996), .B(n12997), .ZN(n12994) );
  XOR2_X1 U12993 ( .A(n12998), .B(n12999), .Z(n12750) );
  XNOR2_X1 U12994 ( .A(n13000), .B(n13001), .ZN(n12998) );
  XOR2_X1 U12995 ( .A(n13002), .B(n13003), .Z(n12754) );
  XNOR2_X1 U12996 ( .A(n13004), .B(n13005), .ZN(n13002) );
  XOR2_X1 U12997 ( .A(n13006), .B(n13007), .Z(n12758) );
  XNOR2_X1 U12998 ( .A(n13008), .B(n13009), .ZN(n13006) );
  XNOR2_X1 U12999 ( .A(n13010), .B(n13011), .ZN(n12762) );
  XOR2_X1 U13000 ( .A(n13012), .B(n13013), .Z(n13010) );
  XNOR2_X1 U13001 ( .A(n13014), .B(n13015), .ZN(n12766) );
  XOR2_X1 U13002 ( .A(n13016), .B(n13017), .Z(n13014) );
  XOR2_X1 U13003 ( .A(n13018), .B(n13019), .Z(n12770) );
  XNOR2_X1 U13004 ( .A(n13020), .B(n13021), .ZN(n13018) );
  XNOR2_X1 U13005 ( .A(n13022), .B(n13023), .ZN(n12774) );
  XOR2_X1 U13006 ( .A(n13024), .B(n13025), .Z(n13023) );
  XNOR2_X1 U13007 ( .A(n13026), .B(n13027), .ZN(n12778) );
  XOR2_X1 U13008 ( .A(n13028), .B(n13029), .Z(n13026) );
  XOR2_X1 U13009 ( .A(n13030), .B(n13031), .Z(n12782) );
  XNOR2_X1 U13010 ( .A(n13032), .B(n13033), .ZN(n13031) );
  XNOR2_X1 U13011 ( .A(n13034), .B(n13035), .ZN(n12786) );
  XOR2_X1 U13012 ( .A(n13036), .B(n13037), .Z(n13034) );
  XNOR2_X1 U13013 ( .A(n13038), .B(n13039), .ZN(n12790) );
  XNOR2_X1 U13014 ( .A(n13040), .B(n13041), .ZN(n13039) );
  XOR2_X1 U13015 ( .A(n13042), .B(n13043), .Z(n12794) );
  XNOR2_X1 U13016 ( .A(n13044), .B(n13045), .ZN(n13042) );
  XNOR2_X1 U13017 ( .A(n13046), .B(n13047), .ZN(n12798) );
  XOR2_X1 U13018 ( .A(n13048), .B(n13049), .Z(n13046) );
  NOR2_X1 U13019 ( .A1(n8591), .A2(n8557), .ZN(n13049) );
  XOR2_X1 U13020 ( .A(n13050), .B(n13051), .Z(n12802) );
  XNOR2_X1 U13021 ( .A(n13052), .B(n13053), .ZN(n13050) );
  NOR2_X1 U13022 ( .A1(n9031), .A2(n8557), .ZN(n13053) );
  XOR2_X1 U13023 ( .A(n13054), .B(n13055), .Z(n12805) );
  XNOR2_X1 U13024 ( .A(n13056), .B(n13057), .ZN(n13054) );
  NOR2_X1 U13025 ( .A1(n9025), .A2(n8557), .ZN(n13057) );
  XNOR2_X1 U13026 ( .A(n13058), .B(n13059), .ZN(n12810) );
  XNOR2_X1 U13027 ( .A(n13060), .B(n13061), .ZN(n13059) );
  NAND2_X1 U13028 ( .A1(n12728), .A2(n9304), .ZN(n13061) );
  XNOR2_X1 U13029 ( .A(n13062), .B(n13063), .ZN(n12814) );
  XOR2_X1 U13030 ( .A(n13064), .B(n13065), .Z(n13062) );
  NOR2_X1 U13031 ( .A1(n8594), .A2(n8557), .ZN(n13065) );
  XNOR2_X1 U13032 ( .A(n13066), .B(n13067), .ZN(n12818) );
  XNOR2_X1 U13033 ( .A(n13068), .B(n13069), .ZN(n13067) );
  NAND2_X1 U13034 ( .A1(n12728), .A2(n9295), .ZN(n13069) );
  XNOR2_X1 U13035 ( .A(n13070), .B(n13071), .ZN(n12822) );
  XNOR2_X1 U13036 ( .A(n13072), .B(n13073), .ZN(n13070) );
  NOR2_X1 U13037 ( .A1(n8544), .A2(n8557), .ZN(n13073) );
  XOR2_X1 U13038 ( .A(n13074), .B(n13075), .Z(n12607) );
  XNOR2_X1 U13039 ( .A(n13076), .B(n13077), .ZN(n13075) );
  NAND2_X1 U13040 ( .A1(n12728), .A2(n10307), .ZN(n13077) );
  XOR2_X1 U13041 ( .A(n13078), .B(n13079), .Z(n12585) );
  XOR2_X1 U13042 ( .A(n13080), .B(n13081), .Z(n13079) );
  NAND2_X1 U13043 ( .A1(n12728), .A2(n9268), .ZN(n13081) );
  NAND2_X1 U13044 ( .A1(n13082), .A2(n13083), .ZN(n12833) );
  XOR2_X1 U13045 ( .A(n13084), .B(n13085), .Z(n12577) );
  XNOR2_X1 U13046 ( .A(n13086), .B(n13087), .ZN(n13085) );
  NAND2_X1 U13047 ( .A1(n12728), .A2(n8872), .ZN(n13087) );
  NOR2_X1 U13048 ( .A1(n13083), .A2(n13082), .ZN(n8906) );
  NOR2_X1 U13049 ( .A1(n13088), .A2(n13089), .ZN(n13082) );
  INV_X1 U13050 ( .A(n13090), .ZN(n13089) );
  NAND3_X1 U13051 ( .A1(n8592), .A2(n13091), .A3(n12728), .ZN(n13090) );
  NAND2_X1 U13052 ( .A1(n13086), .A2(n13084), .ZN(n13091) );
  NOR2_X1 U13053 ( .A1(n13084), .A2(n13086), .ZN(n13088) );
  NOR2_X1 U13054 ( .A1(n13092), .A2(n13093), .ZN(n13086) );
  NOR3_X1 U13055 ( .A1(n8884), .A2(n13094), .A3(n8557), .ZN(n13093) );
  NOR2_X1 U13056 ( .A1(n12840), .A2(n12839), .ZN(n13094) );
  INV_X1 U13057 ( .A(n13095), .ZN(n13092) );
  NAND2_X1 U13058 ( .A1(n12839), .A2(n12840), .ZN(n13095) );
  NAND2_X1 U13059 ( .A1(n13096), .A2(n13097), .ZN(n12840) );
  NAND3_X1 U13060 ( .A1(n9268), .A2(n13098), .A3(n12728), .ZN(n13097) );
  INV_X1 U13061 ( .A(n13099), .ZN(n13098) );
  NOR2_X1 U13062 ( .A1(n13080), .A2(n13078), .ZN(n13099) );
  NAND2_X1 U13063 ( .A1(n13078), .A2(n13080), .ZN(n13096) );
  NAND2_X1 U13064 ( .A1(n13100), .A2(n13101), .ZN(n13080) );
  NAND3_X1 U13065 ( .A1(n9792), .A2(n13102), .A3(n12728), .ZN(n13101) );
  INV_X1 U13066 ( .A(n13103), .ZN(n13102) );
  NOR2_X1 U13067 ( .A1(n12852), .A2(n12851), .ZN(n13103) );
  NAND2_X1 U13068 ( .A1(n12851), .A2(n12852), .ZN(n13100) );
  NAND2_X1 U13069 ( .A1(n13104), .A2(n13105), .ZN(n12852) );
  INV_X1 U13070 ( .A(n13106), .ZN(n13105) );
  NOR3_X1 U13071 ( .A1(n8528), .A2(n13107), .A3(n8557), .ZN(n13106) );
  NOR2_X1 U13072 ( .A1(n12861), .A2(n12859), .ZN(n13107) );
  NAND2_X1 U13073 ( .A1(n12859), .A2(n12861), .ZN(n13104) );
  NAND2_X1 U13074 ( .A1(n13108), .A2(n13109), .ZN(n12861) );
  NAND3_X1 U13075 ( .A1(n10307), .A2(n13110), .A3(n12728), .ZN(n13109) );
  NAND2_X1 U13076 ( .A1(n13076), .A2(n13074), .ZN(n13110) );
  INV_X1 U13077 ( .A(n13111), .ZN(n13108) );
  NOR2_X1 U13078 ( .A1(n13074), .A2(n13076), .ZN(n13111) );
  NOR2_X1 U13079 ( .A1(n13112), .A2(n13113), .ZN(n13076) );
  INV_X1 U13080 ( .A(n13114), .ZN(n13113) );
  NAND3_X1 U13081 ( .A1(n9286), .A2(n13115), .A3(n12728), .ZN(n13114) );
  NAND2_X1 U13082 ( .A1(n12873), .A2(n12871), .ZN(n13115) );
  NOR2_X1 U13083 ( .A1(n12871), .A2(n12873), .ZN(n13112) );
  NOR2_X1 U13084 ( .A1(n13116), .A2(n13117), .ZN(n12873) );
  INV_X1 U13085 ( .A(n13118), .ZN(n13117) );
  NAND3_X1 U13086 ( .A1(n8543), .A2(n13119), .A3(n12728), .ZN(n13118) );
  NAND2_X1 U13087 ( .A1(n13072), .A2(n13071), .ZN(n13119) );
  NOR2_X1 U13088 ( .A1(n13071), .A2(n13072), .ZN(n13116) );
  NOR2_X1 U13089 ( .A1(n13120), .A2(n13121), .ZN(n13072) );
  NOR3_X1 U13090 ( .A1(n9010), .A2(n13122), .A3(n8557), .ZN(n13121) );
  INV_X1 U13091 ( .A(n13123), .ZN(n13122) );
  NAND2_X1 U13092 ( .A1(n13068), .A2(n13066), .ZN(n13123) );
  NOR2_X1 U13093 ( .A1(n13066), .A2(n13068), .ZN(n13120) );
  NOR2_X1 U13094 ( .A1(n13124), .A2(n13125), .ZN(n13068) );
  NOR3_X1 U13095 ( .A1(n9014), .A2(n13126), .A3(n8557), .ZN(n13125) );
  NOR2_X1 U13096 ( .A1(n13064), .A2(n13063), .ZN(n13126) );
  INV_X1 U13097 ( .A(n13127), .ZN(n13124) );
  NAND2_X1 U13098 ( .A1(n13063), .A2(n13064), .ZN(n13127) );
  NAND2_X1 U13099 ( .A1(n13128), .A2(n13129), .ZN(n13064) );
  NAND3_X1 U13100 ( .A1(n9304), .A2(n13130), .A3(n12728), .ZN(n13129) );
  NAND2_X1 U13101 ( .A1(n13060), .A2(n13058), .ZN(n13130) );
  INV_X1 U13102 ( .A(n13131), .ZN(n13128) );
  NOR2_X1 U13103 ( .A1(n13058), .A2(n13060), .ZN(n13131) );
  NOR2_X1 U13104 ( .A1(n13132), .A2(n13133), .ZN(n13060) );
  INV_X1 U13105 ( .A(n13134), .ZN(n13133) );
  NAND3_X1 U13106 ( .A1(n9209), .A2(n13135), .A3(n12728), .ZN(n13134) );
  NAND2_X1 U13107 ( .A1(n13056), .A2(n13055), .ZN(n13135) );
  NOR2_X1 U13108 ( .A1(n13055), .A2(n13056), .ZN(n13132) );
  NOR2_X1 U13109 ( .A1(n13136), .A2(n13137), .ZN(n13056) );
  INV_X1 U13110 ( .A(n13138), .ZN(n13137) );
  NAND3_X1 U13111 ( .A1(n9313), .A2(n13139), .A3(n12728), .ZN(n13138) );
  NAND2_X1 U13112 ( .A1(n13052), .A2(n13051), .ZN(n13139) );
  NOR2_X1 U13113 ( .A1(n13051), .A2(n13052), .ZN(n13136) );
  NOR2_X1 U13114 ( .A1(n13140), .A2(n13141), .ZN(n13052) );
  NOR3_X1 U13115 ( .A1(n9036), .A2(n13142), .A3(n8557), .ZN(n13141) );
  NOR2_X1 U13116 ( .A1(n13048), .A2(n13047), .ZN(n13142) );
  INV_X1 U13117 ( .A(n13143), .ZN(n13140) );
  NAND2_X1 U13118 ( .A1(n13047), .A2(n13048), .ZN(n13143) );
  NAND2_X1 U13119 ( .A1(n12909), .A2(n13144), .ZN(n13048) );
  NAND2_X1 U13120 ( .A1(n12908), .A2(n12910), .ZN(n13144) );
  NAND2_X1 U13121 ( .A1(n13145), .A2(n13146), .ZN(n12910) );
  NAND2_X1 U13122 ( .A1(n12728), .A2(n9322), .ZN(n13146) );
  XNOR2_X1 U13123 ( .A(n13147), .B(n13148), .ZN(n12908) );
  XNOR2_X1 U13124 ( .A(n13149), .B(n13150), .ZN(n13148) );
  NAND2_X1 U13125 ( .A1(n9322), .A2(n13151), .ZN(n12909) );
  INV_X1 U13126 ( .A(n13145), .ZN(n13151) );
  NOR2_X1 U13127 ( .A1(n13152), .A2(n13153), .ZN(n13145) );
  INV_X1 U13128 ( .A(n13154), .ZN(n13153) );
  NAND2_X1 U13129 ( .A1(n13045), .A2(n13155), .ZN(n13154) );
  NAND2_X1 U13130 ( .A1(n13044), .A2(n13043), .ZN(n13155) );
  NOR2_X1 U13131 ( .A1(n8557), .A2(n8545), .ZN(n13045) );
  NOR2_X1 U13132 ( .A1(n13043), .A2(n13044), .ZN(n13152) );
  NOR2_X1 U13133 ( .A1(n13156), .A2(n13157), .ZN(n13044) );
  INV_X1 U13134 ( .A(n13158), .ZN(n13157) );
  NAND2_X1 U13135 ( .A1(n13041), .A2(n13159), .ZN(n13158) );
  NAND2_X1 U13136 ( .A1(n13160), .A2(n13038), .ZN(n13159) );
  NOR2_X1 U13137 ( .A1(n8557), .A2(n8569), .ZN(n13041) );
  NOR2_X1 U13138 ( .A1(n13038), .A2(n13160), .ZN(n13156) );
  INV_X1 U13139 ( .A(n13040), .ZN(n13160) );
  NAND2_X1 U13140 ( .A1(n13161), .A2(n13162), .ZN(n13040) );
  NAND2_X1 U13141 ( .A1(n13037), .A2(n13163), .ZN(n13162) );
  INV_X1 U13142 ( .A(n13164), .ZN(n13163) );
  NOR2_X1 U13143 ( .A1(n13036), .A2(n13035), .ZN(n13164) );
  NOR2_X1 U13144 ( .A1(n8557), .A2(n8593), .ZN(n13037) );
  NAND2_X1 U13145 ( .A1(n13035), .A2(n13036), .ZN(n13161) );
  NAND2_X1 U13146 ( .A1(n13165), .A2(n13166), .ZN(n13036) );
  NAND2_X1 U13147 ( .A1(n13033), .A2(n13167), .ZN(n13166) );
  INV_X1 U13148 ( .A(n13168), .ZN(n13167) );
  NOR2_X1 U13149 ( .A1(n13032), .A2(n13030), .ZN(n13168) );
  NOR2_X1 U13150 ( .A1(n8557), .A2(n8583), .ZN(n13033) );
  NAND2_X1 U13151 ( .A1(n13030), .A2(n13032), .ZN(n13165) );
  NAND2_X1 U13152 ( .A1(n13169), .A2(n13170), .ZN(n13032) );
  NAND2_X1 U13153 ( .A1(n13029), .A2(n13171), .ZN(n13170) );
  INV_X1 U13154 ( .A(n13172), .ZN(n13171) );
  NOR2_X1 U13155 ( .A1(n13028), .A2(n13027), .ZN(n13172) );
  NOR2_X1 U13156 ( .A1(n8557), .A2(n8580), .ZN(n13029) );
  NAND2_X1 U13157 ( .A1(n13027), .A2(n13028), .ZN(n13169) );
  NAND2_X1 U13158 ( .A1(n13173), .A2(n13174), .ZN(n13028) );
  NAND2_X1 U13159 ( .A1(n13025), .A2(n13175), .ZN(n13174) );
  NAND2_X1 U13160 ( .A1(n13024), .A2(n13022), .ZN(n13175) );
  NOR2_X1 U13161 ( .A1(n8557), .A2(n8588), .ZN(n13025) );
  INV_X1 U13162 ( .A(n13176), .ZN(n13173) );
  NOR2_X1 U13163 ( .A1(n13022), .A2(n13024), .ZN(n13176) );
  NOR2_X1 U13164 ( .A1(n13177), .A2(n13178), .ZN(n13024) );
  INV_X1 U13165 ( .A(n13179), .ZN(n13178) );
  NAND2_X1 U13166 ( .A1(n13021), .A2(n13180), .ZN(n13179) );
  NAND2_X1 U13167 ( .A1(n13020), .A2(n13019), .ZN(n13180) );
  NOR2_X1 U13168 ( .A1(n8557), .A2(n8551), .ZN(n13021) );
  NOR2_X1 U13169 ( .A1(n13019), .A2(n13020), .ZN(n13177) );
  INV_X1 U13170 ( .A(n13181), .ZN(n13020) );
  NAND2_X1 U13171 ( .A1(n13182), .A2(n13183), .ZN(n13181) );
  NAND2_X1 U13172 ( .A1(n13016), .A2(n13184), .ZN(n13183) );
  INV_X1 U13173 ( .A(n13185), .ZN(n13184) );
  NOR2_X1 U13174 ( .A1(n13017), .A2(n13015), .ZN(n13185) );
  NOR2_X1 U13175 ( .A1(n12727), .A2(n8563), .ZN(n13016) );
  NAND2_X1 U13176 ( .A1(n13015), .A2(n13017), .ZN(n13182) );
  NAND2_X1 U13177 ( .A1(n13186), .A2(n13187), .ZN(n13017) );
  NAND2_X1 U13178 ( .A1(n13013), .A2(n13188), .ZN(n13187) );
  INV_X1 U13179 ( .A(n13189), .ZN(n13188) );
  NOR2_X1 U13180 ( .A1(n13012), .A2(n13011), .ZN(n13189) );
  NOR2_X1 U13181 ( .A1(n12727), .A2(n8548), .ZN(n13013) );
  NAND2_X1 U13182 ( .A1(n13011), .A2(n13012), .ZN(n13186) );
  NAND2_X1 U13183 ( .A1(n13190), .A2(n13191), .ZN(n13012) );
  NAND2_X1 U13184 ( .A1(n13008), .A2(n13192), .ZN(n13191) );
  NAND2_X1 U13185 ( .A1(n13009), .A2(n13007), .ZN(n13192) );
  NOR2_X1 U13186 ( .A1(n12727), .A2(n8584), .ZN(n13008) );
  NAND2_X1 U13187 ( .A1(n13193), .A2(n13194), .ZN(n13190) );
  INV_X1 U13188 ( .A(n13009), .ZN(n13194) );
  NOR2_X1 U13189 ( .A1(n13195), .A2(n13196), .ZN(n13009) );
  INV_X1 U13190 ( .A(n13197), .ZN(n13196) );
  NAND2_X1 U13191 ( .A1(n13005), .A2(n13198), .ZN(n13197) );
  NAND2_X1 U13192 ( .A1(n13004), .A2(n13003), .ZN(n13198) );
  NOR2_X1 U13193 ( .A1(n12727), .A2(n8535), .ZN(n13005) );
  NOR2_X1 U13194 ( .A1(n13003), .A2(n13004), .ZN(n13195) );
  NOR2_X1 U13195 ( .A1(n13199), .A2(n13200), .ZN(n13004) );
  INV_X1 U13196 ( .A(n13201), .ZN(n13200) );
  NAND2_X1 U13197 ( .A1(n13000), .A2(n13202), .ZN(n13201) );
  NAND2_X1 U13198 ( .A1(n13001), .A2(n12999), .ZN(n13202) );
  NOR2_X1 U13199 ( .A1(n12727), .A2(n8568), .ZN(n13000) );
  NOR2_X1 U13200 ( .A1(n12999), .A2(n13001), .ZN(n13199) );
  NOR2_X1 U13201 ( .A1(n13203), .A2(n13204), .ZN(n13001) );
  INV_X1 U13202 ( .A(n13205), .ZN(n13204) );
  NAND2_X1 U13203 ( .A1(n12996), .A2(n13206), .ZN(n13205) );
  NAND2_X1 U13204 ( .A1(n12997), .A2(n12995), .ZN(n13206) );
  NOR2_X1 U13205 ( .A1(n12727), .A2(n8574), .ZN(n12996) );
  NOR2_X1 U13206 ( .A1(n12995), .A2(n12997), .ZN(n13203) );
  NOR2_X1 U13207 ( .A1(n13207), .A2(n13208), .ZN(n12997) );
  INV_X1 U13208 ( .A(n13209), .ZN(n13208) );
  NAND2_X1 U13209 ( .A1(n12992), .A2(n13210), .ZN(n13209) );
  NAND2_X1 U13210 ( .A1(n12993), .A2(n12991), .ZN(n13210) );
  NOR2_X1 U13211 ( .A1(n12727), .A2(n8565), .ZN(n12992) );
  NOR2_X1 U13212 ( .A1(n12991), .A2(n12993), .ZN(n13207) );
  NOR2_X1 U13213 ( .A1(n13211), .A2(n13212), .ZN(n12993) );
  INV_X1 U13214 ( .A(n13213), .ZN(n13212) );
  NAND2_X1 U13215 ( .A1(n12986), .A2(n13214), .ZN(n13213) );
  NAND2_X1 U13216 ( .A1(n12989), .A2(n12988), .ZN(n13214) );
  NOR2_X1 U13217 ( .A1(n12727), .A2(n8567), .ZN(n12986) );
  NOR2_X1 U13218 ( .A1(n12988), .A2(n12989), .ZN(n13211) );
  INV_X1 U13219 ( .A(n13215), .ZN(n12989) );
  NAND2_X1 U13220 ( .A1(n13216), .A2(n13217), .ZN(n13215) );
  NAND2_X1 U13221 ( .A1(n12981), .A2(n13218), .ZN(n13217) );
  NAND2_X1 U13222 ( .A1(n8624), .A2(n13219), .ZN(n13218) );
  NAND2_X1 U13223 ( .A1(n8531), .A2(n8585), .ZN(n13219) );
  NAND2_X1 U13224 ( .A1(n13220), .A2(n13221), .ZN(n13216) );
  NAND2_X1 U13225 ( .A1(n8630), .A2(n13222), .ZN(n13221) );
  NAND2_X1 U13226 ( .A1(n8539), .A2(n8570), .ZN(n13222) );
  NAND3_X1 U13227 ( .A1(n12728), .A2(n8537), .A3(n12981), .ZN(n12988) );
  INV_X1 U13228 ( .A(n12727), .ZN(n12728) );
  XNOR2_X1 U13229 ( .A(n13223), .B(n13224), .ZN(n12727) );
  XOR2_X1 U13230 ( .A(d_15_), .B(c_15_), .Z(n13224) );
  XOR2_X1 U13231 ( .A(n13225), .B(n13226), .Z(n12991) );
  XNOR2_X1 U13232 ( .A(n13227), .B(n13228), .ZN(n13226) );
  XOR2_X1 U13233 ( .A(n13229), .B(n13230), .Z(n12995) );
  XNOR2_X1 U13234 ( .A(n13231), .B(n13232), .ZN(n13229) );
  XOR2_X1 U13235 ( .A(n13233), .B(n13234), .Z(n12999) );
  XNOR2_X1 U13236 ( .A(n13235), .B(n13236), .ZN(n13233) );
  XOR2_X1 U13237 ( .A(n13237), .B(n13238), .Z(n13003) );
  XNOR2_X1 U13238 ( .A(n13239), .B(n13240), .ZN(n13237) );
  INV_X1 U13239 ( .A(n13007), .ZN(n13193) );
  XOR2_X1 U13240 ( .A(n13241), .B(n13242), .Z(n13007) );
  XOR2_X1 U13241 ( .A(n13243), .B(n13244), .Z(n13241) );
  NAND2_X1 U13242 ( .A1(n12981), .A2(n9121), .ZN(n13243) );
  XNOR2_X1 U13243 ( .A(n13245), .B(n13246), .ZN(n13011) );
  XNOR2_X1 U13244 ( .A(n13247), .B(n13248), .ZN(n13245) );
  NOR2_X1 U13245 ( .A1(n8584), .A2(n8570), .ZN(n13248) );
  XNOR2_X1 U13246 ( .A(n13249), .B(n13250), .ZN(n13015) );
  XNOR2_X1 U13247 ( .A(n13251), .B(n13252), .ZN(n13249) );
  NOR2_X1 U13248 ( .A1(n8548), .A2(n8570), .ZN(n13252) );
  XOR2_X1 U13249 ( .A(n13253), .B(n13254), .Z(n13019) );
  XNOR2_X1 U13250 ( .A(n13255), .B(n13256), .ZN(n13253) );
  NOR2_X1 U13251 ( .A1(n9094), .A2(n8570), .ZN(n13256) );
  XOR2_X1 U13252 ( .A(n13257), .B(n13258), .Z(n13022) );
  XNOR2_X1 U13253 ( .A(n13259), .B(n13260), .ZN(n13257) );
  NOR2_X1 U13254 ( .A1(n8551), .A2(n8570), .ZN(n13260) );
  XNOR2_X1 U13255 ( .A(n13261), .B(n13262), .ZN(n13027) );
  XNOR2_X1 U13256 ( .A(n13263), .B(n13264), .ZN(n13261) );
  NOR2_X1 U13257 ( .A1(n8588), .A2(n8570), .ZN(n13264) );
  XNOR2_X1 U13258 ( .A(n13265), .B(n13266), .ZN(n13030) );
  XNOR2_X1 U13259 ( .A(n13267), .B(n13268), .ZN(n13265) );
  NOR2_X1 U13260 ( .A1(n8580), .A2(n8570), .ZN(n13268) );
  XNOR2_X1 U13261 ( .A(n13269), .B(n13270), .ZN(n13035) );
  XNOR2_X1 U13262 ( .A(n13271), .B(n13272), .ZN(n13269) );
  NOR2_X1 U13263 ( .A1(n9061), .A2(n8570), .ZN(n13272) );
  XOR2_X1 U13264 ( .A(n13273), .B(n13274), .Z(n13038) );
  XNOR2_X1 U13265 ( .A(n13275), .B(n13276), .ZN(n13273) );
  NOR2_X1 U13266 ( .A1(n8593), .A2(n8570), .ZN(n13276) );
  XOR2_X1 U13267 ( .A(n13277), .B(n13278), .Z(n13043) );
  XNOR2_X1 U13268 ( .A(n13279), .B(n13280), .ZN(n13277) );
  NOR2_X1 U13269 ( .A1(n9050), .A2(n8570), .ZN(n13280) );
  XOR2_X1 U13270 ( .A(n13281), .B(n13282), .Z(n13047) );
  XOR2_X1 U13271 ( .A(n13283), .B(n13284), .Z(n13281) );
  XOR2_X1 U13272 ( .A(n13285), .B(n13286), .Z(n13051) );
  XNOR2_X1 U13273 ( .A(n13287), .B(n13288), .ZN(n13285) );
  XOR2_X1 U13274 ( .A(n13289), .B(n13290), .Z(n13055) );
  XNOR2_X1 U13275 ( .A(n13291), .B(n13292), .ZN(n13289) );
  XOR2_X1 U13276 ( .A(n13293), .B(n13294), .Z(n13058) );
  XNOR2_X1 U13277 ( .A(n13295), .B(n13296), .ZN(n13293) );
  XNOR2_X1 U13278 ( .A(n13297), .B(n13298), .ZN(n13063) );
  XNOR2_X1 U13279 ( .A(n13299), .B(n13300), .ZN(n13297) );
  XNOR2_X1 U13280 ( .A(n13301), .B(n13302), .ZN(n13066) );
  XNOR2_X1 U13281 ( .A(n13303), .B(n13304), .ZN(n13301) );
  NOR2_X1 U13282 ( .A1(n8594), .A2(n8570), .ZN(n13304) );
  XOR2_X1 U13283 ( .A(n13305), .B(n13306), .Z(n13071) );
  NAND2_X1 U13284 ( .A1(n13307), .A2(n13308), .ZN(n13305) );
  XOR2_X1 U13285 ( .A(n13309), .B(n13310), .Z(n12871) );
  XOR2_X1 U13286 ( .A(n13311), .B(n13312), .Z(n13310) );
  XNOR2_X1 U13287 ( .A(n13313), .B(n13314), .ZN(n13074) );
  XNOR2_X1 U13288 ( .A(n13315), .B(n13316), .ZN(n13313) );
  NOR2_X1 U13289 ( .A1(n8555), .A2(n8570), .ZN(n13316) );
  XNOR2_X1 U13290 ( .A(n13317), .B(n13318), .ZN(n12859) );
  NAND2_X1 U13291 ( .A1(n13319), .A2(n13320), .ZN(n13317) );
  XNOR2_X1 U13292 ( .A(n13321), .B(n13322), .ZN(n12851) );
  XOR2_X1 U13293 ( .A(n13323), .B(n13324), .Z(n13321) );
  XOR2_X1 U13294 ( .A(n13325), .B(n13326), .Z(n13078) );
  XNOR2_X1 U13295 ( .A(n13327), .B(n13328), .ZN(n13326) );
  NAND2_X1 U13296 ( .A1(n12981), .A2(n9792), .ZN(n13328) );
  XNOR2_X1 U13297 ( .A(n13329), .B(n13330), .ZN(n12839) );
  NAND2_X1 U13298 ( .A1(n13331), .A2(n13332), .ZN(n13329) );
  XOR2_X1 U13299 ( .A(n13333), .B(n13334), .Z(n13084) );
  XOR2_X1 U13300 ( .A(n13335), .B(n13336), .Z(n13333) );
  XNOR2_X1 U13301 ( .A(n13337), .B(n13338), .ZN(n13083) );
  XOR2_X1 U13302 ( .A(n13339), .B(n13340), .Z(n13338) );
  XNOR2_X1 U13303 ( .A(n13341), .B(n13342), .ZN(n8851) );
  NAND2_X1 U13304 ( .A1(n8858), .A2(n8857), .ZN(n8856) );
  NOR2_X1 U13305 ( .A1(n13343), .A2(n8903), .ZN(n8857) );
  INV_X1 U13306 ( .A(n13344), .ZN(n13343) );
  NAND2_X1 U13307 ( .A1(n13345), .A2(n13346), .ZN(n13344) );
  XNOR2_X1 U13308 ( .A(n13347), .B(n13348), .ZN(n13345) );
  INV_X1 U13309 ( .A(n13349), .ZN(n8858) );
  NAND2_X1 U13310 ( .A1(n13342), .A2(n13341), .ZN(n13349) );
  NAND2_X1 U13311 ( .A1(n13350), .A2(n13351), .ZN(n13341) );
  NAND2_X1 U13312 ( .A1(n13340), .A2(n13352), .ZN(n13351) );
  INV_X1 U13313 ( .A(n13353), .ZN(n13352) );
  NOR2_X1 U13314 ( .A1(n13337), .A2(n13339), .ZN(n13353) );
  NOR2_X1 U13315 ( .A1(n8570), .A2(n8972), .ZN(n13340) );
  NAND2_X1 U13316 ( .A1(n13337), .A2(n13339), .ZN(n13350) );
  NOR2_X1 U13317 ( .A1(n13354), .A2(n13355), .ZN(n13339) );
  INV_X1 U13318 ( .A(n13356), .ZN(n13355) );
  NAND2_X1 U13319 ( .A1(n13334), .A2(n13357), .ZN(n13356) );
  NAND2_X1 U13320 ( .A1(n13336), .A2(n13335), .ZN(n13357) );
  XOR2_X1 U13321 ( .A(n13358), .B(n13359), .Z(n13334) );
  XOR2_X1 U13322 ( .A(n13360), .B(n13361), .Z(n13359) );
  NAND2_X1 U13323 ( .A1(n13220), .A2(n9268), .ZN(n13361) );
  NOR2_X1 U13324 ( .A1(n13335), .A2(n13336), .ZN(n13354) );
  NOR2_X1 U13325 ( .A1(n8570), .A2(n8589), .ZN(n13336) );
  NAND2_X1 U13326 ( .A1(n13331), .A2(n13362), .ZN(n13335) );
  NAND2_X1 U13327 ( .A1(n13330), .A2(n13332), .ZN(n13362) );
  NAND2_X1 U13328 ( .A1(n13363), .A2(n13364), .ZN(n13332) );
  NAND2_X1 U13329 ( .A1(n12981), .A2(n9268), .ZN(n13364) );
  INV_X1 U13330 ( .A(n13365), .ZN(n13363) );
  XNOR2_X1 U13331 ( .A(n13366), .B(n13367), .ZN(n13330) );
  XOR2_X1 U13332 ( .A(n13368), .B(n13369), .Z(n13367) );
  NAND2_X1 U13333 ( .A1(n13220), .A2(n9792), .ZN(n13369) );
  NAND2_X1 U13334 ( .A1(n9268), .A2(n13365), .ZN(n13331) );
  NAND2_X1 U13335 ( .A1(n13370), .A2(n13371), .ZN(n13365) );
  NAND3_X1 U13336 ( .A1(n9792), .A2(n13372), .A3(n12981), .ZN(n13371) );
  NAND2_X1 U13337 ( .A1(n13373), .A2(n13374), .ZN(n13372) );
  INV_X1 U13338 ( .A(n13327), .ZN(n13374) );
  INV_X1 U13339 ( .A(n13325), .ZN(n13373) );
  NAND2_X1 U13340 ( .A1(n13327), .A2(n13325), .ZN(n13370) );
  XNOR2_X1 U13341 ( .A(n13375), .B(n13376), .ZN(n13325) );
  XOR2_X1 U13342 ( .A(n13377), .B(n13378), .Z(n13376) );
  NAND2_X1 U13343 ( .A1(n13220), .A2(n9277), .ZN(n13378) );
  NOR2_X1 U13344 ( .A1(n13379), .A2(n13380), .ZN(n13327) );
  INV_X1 U13345 ( .A(n13381), .ZN(n13380) );
  NAND2_X1 U13346 ( .A1(n13322), .A2(n13382), .ZN(n13381) );
  NAND2_X1 U13347 ( .A1(n13324), .A2(n13323), .ZN(n13382) );
  XOR2_X1 U13348 ( .A(n13383), .B(n13384), .Z(n13322) );
  XOR2_X1 U13349 ( .A(n13385), .B(n13386), .Z(n13384) );
  NAND2_X1 U13350 ( .A1(n13220), .A2(n10307), .ZN(n13386) );
  NOR2_X1 U13351 ( .A1(n13323), .A2(n13324), .ZN(n13379) );
  NOR2_X1 U13352 ( .A1(n8570), .A2(n8528), .ZN(n13324) );
  NAND2_X1 U13353 ( .A1(n13319), .A2(n13387), .ZN(n13323) );
  NAND2_X1 U13354 ( .A1(n13318), .A2(n13320), .ZN(n13387) );
  NAND2_X1 U13355 ( .A1(n13388), .A2(n13389), .ZN(n13320) );
  NAND2_X1 U13356 ( .A1(n12981), .A2(n10307), .ZN(n13389) );
  XOR2_X1 U13357 ( .A(n13390), .B(n13391), .Z(n13318) );
  XNOR2_X1 U13358 ( .A(n13392), .B(n13393), .ZN(n13391) );
  NAND2_X1 U13359 ( .A1(n13220), .A2(n9286), .ZN(n13393) );
  INV_X1 U13360 ( .A(n13394), .ZN(n13319) );
  NOR2_X1 U13361 ( .A1(n8564), .A2(n13388), .ZN(n13394) );
  NOR2_X1 U13362 ( .A1(n13395), .A2(n13396), .ZN(n13388) );
  NOR3_X1 U13363 ( .A1(n9000), .A2(n13397), .A3(n8570), .ZN(n13396) );
  NOR2_X1 U13364 ( .A1(n13314), .A2(n13398), .ZN(n13397) );
  INV_X1 U13365 ( .A(n13315), .ZN(n13398) );
  NOR2_X1 U13366 ( .A1(n13399), .A2(n13315), .ZN(n13395) );
  NOR2_X1 U13367 ( .A1(n13400), .A2(n13401), .ZN(n13315) );
  NOR2_X1 U13368 ( .A1(n13312), .A2(n13402), .ZN(n13401) );
  NOR2_X1 U13369 ( .A1(n13309), .A2(n13311), .ZN(n13402) );
  NAND2_X1 U13370 ( .A1(n12981), .A2(n8543), .ZN(n13312) );
  INV_X1 U13371 ( .A(n13403), .ZN(n13400) );
  NAND2_X1 U13372 ( .A1(n13309), .A2(n13311), .ZN(n13403) );
  NAND2_X1 U13373 ( .A1(n13307), .A2(n13404), .ZN(n13311) );
  NAND2_X1 U13374 ( .A1(n13306), .A2(n13308), .ZN(n13404) );
  NAND2_X1 U13375 ( .A1(n13405), .A2(n13406), .ZN(n13308) );
  NAND2_X1 U13376 ( .A1(n12981), .A2(n9295), .ZN(n13406) );
  XNOR2_X1 U13377 ( .A(n13407), .B(n13408), .ZN(n13306) );
  XOR2_X1 U13378 ( .A(n13409), .B(n13410), .Z(n13408) );
  NAND2_X1 U13379 ( .A1(n13220), .A2(n10846), .ZN(n13410) );
  INV_X1 U13380 ( .A(n13411), .ZN(n13307) );
  NOR2_X1 U13381 ( .A1(n9010), .A2(n13405), .ZN(n13411) );
  NOR2_X1 U13382 ( .A1(n13412), .A2(n13413), .ZN(n13405) );
  NOR3_X1 U13383 ( .A1(n9014), .A2(n13414), .A3(n8570), .ZN(n13413) );
  NOR2_X1 U13384 ( .A1(n13302), .A2(n13415), .ZN(n13414) );
  INV_X1 U13385 ( .A(n13303), .ZN(n13415) );
  NOR2_X1 U13386 ( .A1(n13416), .A2(n13303), .ZN(n13412) );
  NOR2_X1 U13387 ( .A1(n13417), .A2(n13418), .ZN(n13303) );
  INV_X1 U13388 ( .A(n13419), .ZN(n13418) );
  NAND2_X1 U13389 ( .A1(n13299), .A2(n13420), .ZN(n13419) );
  NAND2_X1 U13390 ( .A1(n13300), .A2(n13298), .ZN(n13420) );
  NOR2_X1 U13391 ( .A1(n12980), .A2(n8556), .ZN(n13299) );
  NOR2_X1 U13392 ( .A1(n13298), .A2(n13300), .ZN(n13417) );
  NOR2_X1 U13393 ( .A1(n13421), .A2(n13422), .ZN(n13300) );
  INV_X1 U13394 ( .A(n13423), .ZN(n13422) );
  NAND2_X1 U13395 ( .A1(n13296), .A2(n13424), .ZN(n13423) );
  NAND2_X1 U13396 ( .A1(n13295), .A2(n13294), .ZN(n13424) );
  NOR2_X1 U13397 ( .A1(n12980), .A2(n8572), .ZN(n13296) );
  NOR2_X1 U13398 ( .A1(n13294), .A2(n13295), .ZN(n13421) );
  NOR2_X1 U13399 ( .A1(n13425), .A2(n13426), .ZN(n13295) );
  INV_X1 U13400 ( .A(n13427), .ZN(n13426) );
  NAND2_X1 U13401 ( .A1(n13292), .A2(n13428), .ZN(n13427) );
  NAND2_X1 U13402 ( .A1(n13291), .A2(n13290), .ZN(n13428) );
  NOR2_X1 U13403 ( .A1(n12980), .A2(n8582), .ZN(n13292) );
  NOR2_X1 U13404 ( .A1(n13290), .A2(n13291), .ZN(n13425) );
  NOR2_X1 U13405 ( .A1(n13429), .A2(n13430), .ZN(n13291) );
  INV_X1 U13406 ( .A(n13431), .ZN(n13430) );
  NAND2_X1 U13407 ( .A1(n13288), .A2(n13432), .ZN(n13431) );
  NAND2_X1 U13408 ( .A1(n13286), .A2(n13287), .ZN(n13432) );
  NOR2_X1 U13409 ( .A1(n12980), .A2(n8591), .ZN(n13288) );
  NOR2_X1 U13410 ( .A1(n13286), .A2(n13287), .ZN(n13429) );
  INV_X1 U13411 ( .A(n13433), .ZN(n13287) );
  NAND2_X1 U13412 ( .A1(n13434), .A2(n13435), .ZN(n13433) );
  NAND2_X1 U13413 ( .A1(n13284), .A2(n13436), .ZN(n13435) );
  INV_X1 U13414 ( .A(n13437), .ZN(n13436) );
  NOR2_X1 U13415 ( .A1(n13283), .A2(n13282), .ZN(n13437) );
  NOR2_X1 U13416 ( .A1(n12980), .A2(n8562), .ZN(n13284) );
  NAND2_X1 U13417 ( .A1(n13282), .A2(n13283), .ZN(n13434) );
  NAND2_X1 U13418 ( .A1(n13438), .A2(n13439), .ZN(n13283) );
  NAND2_X1 U13419 ( .A1(n13150), .A2(n13440), .ZN(n13439) );
  INV_X1 U13420 ( .A(n13441), .ZN(n13440) );
  NOR2_X1 U13421 ( .A1(n13147), .A2(n13149), .ZN(n13441) );
  NOR2_X1 U13422 ( .A1(n12980), .A2(n8545), .ZN(n13150) );
  NAND2_X1 U13423 ( .A1(n13147), .A2(n13149), .ZN(n13438) );
  NAND2_X1 U13424 ( .A1(n13442), .A2(n13443), .ZN(n13149) );
  NAND3_X1 U13425 ( .A1(n9331), .A2(n13444), .A3(n12981), .ZN(n13443) );
  NAND2_X1 U13426 ( .A1(n13278), .A2(n13279), .ZN(n13444) );
  INV_X1 U13427 ( .A(n13445), .ZN(n13442) );
  NOR2_X1 U13428 ( .A1(n13278), .A2(n13279), .ZN(n13445) );
  NOR2_X1 U13429 ( .A1(n13446), .A2(n13447), .ZN(n13279) );
  INV_X1 U13430 ( .A(n13448), .ZN(n13447) );
  NAND3_X1 U13431 ( .A1(n10722), .A2(n13449), .A3(n12981), .ZN(n13448) );
  NAND2_X1 U13432 ( .A1(n13274), .A2(n13275), .ZN(n13449) );
  NOR2_X1 U13433 ( .A1(n13274), .A2(n13275), .ZN(n13446) );
  NOR2_X1 U13434 ( .A1(n13450), .A2(n13451), .ZN(n13275) );
  INV_X1 U13435 ( .A(n13452), .ZN(n13451) );
  NAND3_X1 U13436 ( .A1(n9340), .A2(n13453), .A3(n12981), .ZN(n13452) );
  NAND2_X1 U13437 ( .A1(n13271), .A2(n13270), .ZN(n13453) );
  NOR2_X1 U13438 ( .A1(n13270), .A2(n13271), .ZN(n13450) );
  NOR2_X1 U13439 ( .A1(n13454), .A2(n13455), .ZN(n13271) );
  NOR3_X1 U13440 ( .A1(n9066), .A2(n13456), .A3(n8570), .ZN(n13455) );
  INV_X1 U13441 ( .A(n13457), .ZN(n13456) );
  NAND2_X1 U13442 ( .A1(n13266), .A2(n13267), .ZN(n13457) );
  NOR2_X1 U13443 ( .A1(n13266), .A2(n13267), .ZN(n13454) );
  NOR2_X1 U13444 ( .A1(n13458), .A2(n13459), .ZN(n13267) );
  INV_X1 U13445 ( .A(n13460), .ZN(n13459) );
  NAND3_X1 U13446 ( .A1(n9080), .A2(n13461), .A3(n12981), .ZN(n13460) );
  NAND2_X1 U13447 ( .A1(n13263), .A2(n13262), .ZN(n13461) );
  NOR2_X1 U13448 ( .A1(n13262), .A2(n13263), .ZN(n13458) );
  NOR2_X1 U13449 ( .A1(n13462), .A2(n13463), .ZN(n13263) );
  NOR3_X1 U13450 ( .A1(n8551), .A2(n13464), .A3(n8570), .ZN(n13463) );
  INV_X1 U13451 ( .A(n13465), .ZN(n13464) );
  NAND2_X1 U13452 ( .A1(n13258), .A2(n13259), .ZN(n13465) );
  NOR2_X1 U13453 ( .A1(n13258), .A2(n13259), .ZN(n13462) );
  NOR2_X1 U13454 ( .A1(n13466), .A2(n13467), .ZN(n13259) );
  INV_X1 U13455 ( .A(n13468), .ZN(n13467) );
  NAND3_X1 U13456 ( .A1(n9098), .A2(n13469), .A3(n12981), .ZN(n13468) );
  NAND2_X1 U13457 ( .A1(n13255), .A2(n13254), .ZN(n13469) );
  NOR2_X1 U13458 ( .A1(n13254), .A2(n13255), .ZN(n13466) );
  NOR2_X1 U13459 ( .A1(n13470), .A2(n13471), .ZN(n13255) );
  NOR3_X1 U13460 ( .A1(n8548), .A2(n13472), .A3(n8570), .ZN(n13471) );
  INV_X1 U13461 ( .A(n13473), .ZN(n13472) );
  NAND2_X1 U13462 ( .A1(n13250), .A2(n13251), .ZN(n13473) );
  NOR2_X1 U13463 ( .A1(n13250), .A2(n13251), .ZN(n13470) );
  NOR2_X1 U13464 ( .A1(n13474), .A2(n13475), .ZN(n13251) );
  INV_X1 U13465 ( .A(n13476), .ZN(n13475) );
  NAND3_X1 U13466 ( .A1(n9112), .A2(n13477), .A3(n12981), .ZN(n13476) );
  NAND2_X1 U13467 ( .A1(n13247), .A2(n13246), .ZN(n13477) );
  NOR2_X1 U13468 ( .A1(n13246), .A2(n13247), .ZN(n13474) );
  NOR2_X1 U13469 ( .A1(n13478), .A2(n13479), .ZN(n13247) );
  INV_X1 U13470 ( .A(n13480), .ZN(n13479) );
  NAND3_X1 U13471 ( .A1(n9121), .A2(n13481), .A3(n12981), .ZN(n13480) );
  NAND2_X1 U13472 ( .A1(n13242), .A2(n13244), .ZN(n13481) );
  NOR2_X1 U13473 ( .A1(n13242), .A2(n13244), .ZN(n13478) );
  NOR2_X1 U13474 ( .A1(n13482), .A2(n13483), .ZN(n13244) );
  INV_X1 U13475 ( .A(n13484), .ZN(n13483) );
  NAND2_X1 U13476 ( .A1(n13240), .A2(n13485), .ZN(n13484) );
  NAND2_X1 U13477 ( .A1(n13239), .A2(n13238), .ZN(n13485) );
  NOR2_X1 U13478 ( .A1(n12980), .A2(n8568), .ZN(n13240) );
  NOR2_X1 U13479 ( .A1(n13238), .A2(n13239), .ZN(n13482) );
  NOR2_X1 U13480 ( .A1(n13486), .A2(n13487), .ZN(n13239) );
  INV_X1 U13481 ( .A(n13488), .ZN(n13487) );
  NAND2_X1 U13482 ( .A1(n13235), .A2(n13489), .ZN(n13488) );
  NAND2_X1 U13483 ( .A1(n13234), .A2(n13236), .ZN(n13489) );
  NOR2_X1 U13484 ( .A1(n12980), .A2(n8574), .ZN(n13235) );
  NOR2_X1 U13485 ( .A1(n13234), .A2(n13236), .ZN(n13486) );
  NOR2_X1 U13486 ( .A1(n13490), .A2(n13491), .ZN(n13236) );
  INV_X1 U13487 ( .A(n13492), .ZN(n13491) );
  NAND2_X1 U13488 ( .A1(n13231), .A2(n13493), .ZN(n13492) );
  NAND2_X1 U13489 ( .A1(n13232), .A2(n13230), .ZN(n13493) );
  NOR2_X1 U13490 ( .A1(n12980), .A2(n8565), .ZN(n13231) );
  NOR2_X1 U13491 ( .A1(n13230), .A2(n13232), .ZN(n13490) );
  NOR2_X1 U13492 ( .A1(n13494), .A2(n13495), .ZN(n13232) );
  INV_X1 U13493 ( .A(n13496), .ZN(n13495) );
  NAND2_X1 U13494 ( .A1(n13225), .A2(n13497), .ZN(n13496) );
  NAND2_X1 U13495 ( .A1(n13228), .A2(n13227), .ZN(n13497) );
  NOR2_X1 U13496 ( .A1(n12980), .A2(n8567), .ZN(n13225) );
  NOR2_X1 U13497 ( .A1(n13227), .A2(n13228), .ZN(n13494) );
  INV_X1 U13498 ( .A(n13498), .ZN(n13228) );
  NAND2_X1 U13499 ( .A1(n13499), .A2(n13500), .ZN(n13498) );
  NAND2_X1 U13500 ( .A1(n13220), .A2(n13501), .ZN(n13500) );
  NAND2_X1 U13501 ( .A1(n8624), .A2(n13502), .ZN(n13501) );
  NAND2_X1 U13502 ( .A1(n8553), .A2(n8585), .ZN(n13502) );
  NAND2_X1 U13503 ( .A1(n13504), .A2(n13505), .ZN(n13499) );
  NAND2_X1 U13504 ( .A1(n8630), .A2(n13506), .ZN(n13505) );
  NAND2_X1 U13505 ( .A1(n8539), .A2(n8531), .ZN(n13506) );
  NAND3_X1 U13506 ( .A1(n13220), .A2(n8537), .A3(n12981), .ZN(n13227) );
  INV_X1 U13507 ( .A(n12980), .ZN(n12981) );
  XNOR2_X1 U13508 ( .A(n13507), .B(n13508), .ZN(n12980) );
  XOR2_X1 U13509 ( .A(d_14_), .B(c_14_), .Z(n13508) );
  XOR2_X1 U13510 ( .A(n13509), .B(n13510), .Z(n13230) );
  XNOR2_X1 U13511 ( .A(n13511), .B(n13512), .ZN(n13510) );
  XOR2_X1 U13512 ( .A(n13513), .B(n13514), .Z(n13234) );
  XNOR2_X1 U13513 ( .A(n13515), .B(n13516), .ZN(n13513) );
  XOR2_X1 U13514 ( .A(n13517), .B(n13518), .Z(n13238) );
  XNOR2_X1 U13515 ( .A(n13519), .B(n13520), .ZN(n13517) );
  XOR2_X1 U13516 ( .A(n13521), .B(n13522), .Z(n13242) );
  XNOR2_X1 U13517 ( .A(n13523), .B(n13524), .ZN(n13521) );
  XOR2_X1 U13518 ( .A(n13525), .B(n13526), .Z(n13246) );
  XNOR2_X1 U13519 ( .A(n13527), .B(n13528), .ZN(n13525) );
  XOR2_X1 U13520 ( .A(n13529), .B(n13530), .Z(n13250) );
  XNOR2_X1 U13521 ( .A(n13531), .B(n13532), .ZN(n13529) );
  XOR2_X1 U13522 ( .A(n13533), .B(n13534), .Z(n13254) );
  XNOR2_X1 U13523 ( .A(n13535), .B(n13536), .ZN(n13533) );
  XNOR2_X1 U13524 ( .A(n13537), .B(n13538), .ZN(n13258) );
  XOR2_X1 U13525 ( .A(n13539), .B(n13540), .Z(n13538) );
  XNOR2_X1 U13526 ( .A(n13541), .B(n13542), .ZN(n13262) );
  XOR2_X1 U13527 ( .A(n13543), .B(n13544), .Z(n13541) );
  XOR2_X1 U13528 ( .A(n13545), .B(n13546), .Z(n13266) );
  XNOR2_X1 U13529 ( .A(n13547), .B(n13548), .ZN(n13546) );
  XNOR2_X1 U13530 ( .A(n13549), .B(n13550), .ZN(n13270) );
  XOR2_X1 U13531 ( .A(n13551), .B(n13552), .Z(n13549) );
  XNOR2_X1 U13532 ( .A(n13553), .B(n13554), .ZN(n13274) );
  XNOR2_X1 U13533 ( .A(n13555), .B(n13556), .ZN(n13554) );
  XOR2_X1 U13534 ( .A(n13557), .B(n13558), .Z(n13278) );
  XNOR2_X1 U13535 ( .A(n13559), .B(n13560), .ZN(n13557) );
  XNOR2_X1 U13536 ( .A(n13561), .B(n13562), .ZN(n13147) );
  NAND2_X1 U13537 ( .A1(n13563), .A2(n13564), .ZN(n13561) );
  XOR2_X1 U13538 ( .A(n13565), .B(n13566), .Z(n13282) );
  XOR2_X1 U13539 ( .A(n13567), .B(n13568), .Z(n13565) );
  NOR2_X1 U13540 ( .A1(n8545), .A2(n8531), .ZN(n13568) );
  XOR2_X1 U13541 ( .A(n13569), .B(n13570), .Z(n13286) );
  XOR2_X1 U13542 ( .A(n13571), .B(n13572), .Z(n13570) );
  NAND2_X1 U13543 ( .A1(n13220), .A2(n9322), .ZN(n13572) );
  XNOR2_X1 U13544 ( .A(n13573), .B(n13574), .ZN(n13290) );
  XOR2_X1 U13545 ( .A(n13575), .B(n13576), .Z(n13573) );
  NOR2_X1 U13546 ( .A1(n8591), .A2(n8531), .ZN(n13576) );
  XOR2_X1 U13547 ( .A(n13577), .B(n13578), .Z(n13294) );
  XOR2_X1 U13548 ( .A(n13579), .B(n13580), .Z(n13578) );
  NAND2_X1 U13549 ( .A1(n13220), .A2(n9313), .ZN(n13580) );
  XNOR2_X1 U13550 ( .A(n13581), .B(n13582), .ZN(n13298) );
  XOR2_X1 U13551 ( .A(n13583), .B(n13584), .Z(n13581) );
  NOR2_X1 U13552 ( .A1(n9025), .A2(n8531), .ZN(n13584) );
  INV_X1 U13553 ( .A(n13302), .ZN(n13416) );
  XNOR2_X1 U13554 ( .A(n13585), .B(n13586), .ZN(n13302) );
  XOR2_X1 U13555 ( .A(n13587), .B(n13588), .Z(n13586) );
  NAND2_X1 U13556 ( .A1(n13220), .A2(n9304), .ZN(n13588) );
  XNOR2_X1 U13557 ( .A(n13589), .B(n13590), .ZN(n13309) );
  XOR2_X1 U13558 ( .A(n13591), .B(n13592), .Z(n13590) );
  NAND2_X1 U13559 ( .A1(n13220), .A2(n9295), .ZN(n13592) );
  INV_X1 U13560 ( .A(n13314), .ZN(n13399) );
  XOR2_X1 U13561 ( .A(n13593), .B(n13594), .Z(n13314) );
  XNOR2_X1 U13562 ( .A(n13595), .B(n13596), .ZN(n13594) );
  NAND2_X1 U13563 ( .A1(n13220), .A2(n8543), .ZN(n13596) );
  XNOR2_X1 U13564 ( .A(n13597), .B(n13598), .ZN(n13337) );
  XOR2_X1 U13565 ( .A(n13599), .B(n13600), .Z(n13598) );
  NAND2_X1 U13566 ( .A1(n13220), .A2(n9263), .ZN(n13600) );
  XOR2_X1 U13567 ( .A(n13601), .B(n13602), .Z(n13342) );
  XNOR2_X1 U13568 ( .A(n13603), .B(n13604), .ZN(n13602) );
  NAND2_X1 U13569 ( .A1(n13220), .A2(n8872), .ZN(n13604) );
  NOR2_X1 U13570 ( .A1(n13605), .A2(n13346), .ZN(n8903) );
  NOR2_X1 U13571 ( .A1(n13606), .A2(n13607), .ZN(n13346) );
  INV_X1 U13572 ( .A(n13608), .ZN(n13607) );
  NAND3_X1 U13573 ( .A1(n8592), .A2(n13609), .A3(n13220), .ZN(n13608) );
  NAND2_X1 U13574 ( .A1(n13603), .A2(n13601), .ZN(n13609) );
  NOR2_X1 U13575 ( .A1(n13601), .A2(n13603), .ZN(n13606) );
  NOR2_X1 U13576 ( .A1(n13610), .A2(n13611), .ZN(n13603) );
  NOR3_X1 U13577 ( .A1(n8884), .A2(n13612), .A3(n8531), .ZN(n13611) );
  NOR2_X1 U13578 ( .A1(n13599), .A2(n13597), .ZN(n13612) );
  INV_X1 U13579 ( .A(n13613), .ZN(n13610) );
  NAND2_X1 U13580 ( .A1(n13597), .A2(n13599), .ZN(n13613) );
  NAND2_X1 U13581 ( .A1(n13614), .A2(n13615), .ZN(n13599) );
  INV_X1 U13582 ( .A(n13616), .ZN(n13615) );
  NOR3_X1 U13583 ( .A1(n8982), .A2(n13617), .A3(n8531), .ZN(n13616) );
  NOR2_X1 U13584 ( .A1(n13360), .A2(n13358), .ZN(n13617) );
  NAND2_X1 U13585 ( .A1(n13358), .A2(n13360), .ZN(n13614) );
  NAND2_X1 U13586 ( .A1(n13618), .A2(n13619), .ZN(n13360) );
  NAND3_X1 U13587 ( .A1(n9792), .A2(n13620), .A3(n13220), .ZN(n13619) );
  INV_X1 U13588 ( .A(n13621), .ZN(n13620) );
  NOR2_X1 U13589 ( .A1(n13368), .A2(n13366), .ZN(n13621) );
  NAND2_X1 U13590 ( .A1(n13366), .A2(n13368), .ZN(n13618) );
  NAND2_X1 U13591 ( .A1(n13622), .A2(n13623), .ZN(n13368) );
  INV_X1 U13592 ( .A(n13624), .ZN(n13623) );
  NOR3_X1 U13593 ( .A1(n8528), .A2(n13625), .A3(n8531), .ZN(n13624) );
  NOR2_X1 U13594 ( .A1(n13377), .A2(n13375), .ZN(n13625) );
  NAND2_X1 U13595 ( .A1(n13375), .A2(n13377), .ZN(n13622) );
  NAND2_X1 U13596 ( .A1(n13626), .A2(n13627), .ZN(n13377) );
  NAND3_X1 U13597 ( .A1(n10307), .A2(n13628), .A3(n13220), .ZN(n13627) );
  INV_X1 U13598 ( .A(n13629), .ZN(n13628) );
  NOR2_X1 U13599 ( .A1(n13385), .A2(n13383), .ZN(n13629) );
  NAND2_X1 U13600 ( .A1(n13383), .A2(n13385), .ZN(n13626) );
  NAND2_X1 U13601 ( .A1(n13630), .A2(n13631), .ZN(n13385) );
  NAND3_X1 U13602 ( .A1(n9286), .A2(n13632), .A3(n13220), .ZN(n13631) );
  NAND2_X1 U13603 ( .A1(n13392), .A2(n13390), .ZN(n13632) );
  INV_X1 U13604 ( .A(n13633), .ZN(n13630) );
  NOR2_X1 U13605 ( .A1(n13390), .A2(n13392), .ZN(n13633) );
  NOR2_X1 U13606 ( .A1(n13634), .A2(n13635), .ZN(n13392) );
  INV_X1 U13607 ( .A(n13636), .ZN(n13635) );
  NAND3_X1 U13608 ( .A1(n8543), .A2(n13637), .A3(n13220), .ZN(n13636) );
  NAND2_X1 U13609 ( .A1(n13595), .A2(n13593), .ZN(n13637) );
  NOR2_X1 U13610 ( .A1(n13593), .A2(n13595), .ZN(n13634) );
  NOR2_X1 U13611 ( .A1(n13638), .A2(n13639), .ZN(n13595) );
  NOR3_X1 U13612 ( .A1(n9010), .A2(n13640), .A3(n8531), .ZN(n13639) );
  NOR2_X1 U13613 ( .A1(n13591), .A2(n13589), .ZN(n13640) );
  INV_X1 U13614 ( .A(n13641), .ZN(n13638) );
  NAND2_X1 U13615 ( .A1(n13589), .A2(n13591), .ZN(n13641) );
  NAND2_X1 U13616 ( .A1(n13642), .A2(n13643), .ZN(n13591) );
  INV_X1 U13617 ( .A(n13644), .ZN(n13643) );
  NOR3_X1 U13618 ( .A1(n9014), .A2(n13645), .A3(n8531), .ZN(n13644) );
  NOR2_X1 U13619 ( .A1(n13409), .A2(n13407), .ZN(n13645) );
  NAND2_X1 U13620 ( .A1(n13407), .A2(n13409), .ZN(n13642) );
  NAND2_X1 U13621 ( .A1(n13646), .A2(n13647), .ZN(n13409) );
  INV_X1 U13622 ( .A(n13648), .ZN(n13647) );
  NOR3_X1 U13623 ( .A1(n9020), .A2(n13649), .A3(n8531), .ZN(n13648) );
  NOR2_X1 U13624 ( .A1(n13587), .A2(n13585), .ZN(n13649) );
  NAND2_X1 U13625 ( .A1(n13585), .A2(n13587), .ZN(n13646) );
  NAND2_X1 U13626 ( .A1(n13650), .A2(n13651), .ZN(n13587) );
  NAND3_X1 U13627 ( .A1(n9209), .A2(n13652), .A3(n13220), .ZN(n13651) );
  INV_X1 U13628 ( .A(n13653), .ZN(n13652) );
  NOR2_X1 U13629 ( .A1(n13583), .A2(n13582), .ZN(n13653) );
  NAND2_X1 U13630 ( .A1(n13582), .A2(n13583), .ZN(n13650) );
  NAND2_X1 U13631 ( .A1(n13654), .A2(n13655), .ZN(n13583) );
  INV_X1 U13632 ( .A(n13656), .ZN(n13655) );
  NOR3_X1 U13633 ( .A1(n9031), .A2(n13657), .A3(n8531), .ZN(n13656) );
  NOR2_X1 U13634 ( .A1(n13579), .A2(n13577), .ZN(n13657) );
  NAND2_X1 U13635 ( .A1(n13577), .A2(n13579), .ZN(n13654) );
  NAND2_X1 U13636 ( .A1(n13658), .A2(n13659), .ZN(n13579) );
  NAND3_X1 U13637 ( .A1(n9721), .A2(n13660), .A3(n13220), .ZN(n13659) );
  INV_X1 U13638 ( .A(n13661), .ZN(n13660) );
  NOR2_X1 U13639 ( .A1(n13575), .A2(n13574), .ZN(n13661) );
  NAND2_X1 U13640 ( .A1(n13574), .A2(n13575), .ZN(n13658) );
  NAND2_X1 U13641 ( .A1(n13662), .A2(n13663), .ZN(n13575) );
  INV_X1 U13642 ( .A(n13664), .ZN(n13663) );
  NOR3_X1 U13643 ( .A1(n9041), .A2(n13665), .A3(n8531), .ZN(n13664) );
  NOR2_X1 U13644 ( .A1(n13571), .A2(n13569), .ZN(n13665) );
  NAND2_X1 U13645 ( .A1(n13569), .A2(n13571), .ZN(n13662) );
  NAND2_X1 U13646 ( .A1(n13666), .A2(n13667), .ZN(n13571) );
  NAND3_X1 U13647 ( .A1(n10222), .A2(n13668), .A3(n13220), .ZN(n13667) );
  INV_X1 U13648 ( .A(n13669), .ZN(n13668) );
  NOR2_X1 U13649 ( .A1(n13567), .A2(n13566), .ZN(n13669) );
  NAND2_X1 U13650 ( .A1(n13566), .A2(n13567), .ZN(n13666) );
  NAND2_X1 U13651 ( .A1(n13563), .A2(n13670), .ZN(n13567) );
  NAND2_X1 U13652 ( .A1(n13562), .A2(n13564), .ZN(n13670) );
  NAND2_X1 U13653 ( .A1(n13671), .A2(n13672), .ZN(n13564) );
  NAND2_X1 U13654 ( .A1(n13220), .A2(n9331), .ZN(n13672) );
  XOR2_X1 U13655 ( .A(n13673), .B(n13674), .Z(n13562) );
  XOR2_X1 U13656 ( .A(n13675), .B(n13676), .Z(n13674) );
  NAND2_X1 U13657 ( .A1(n9331), .A2(n13677), .ZN(n13563) );
  INV_X1 U13658 ( .A(n13671), .ZN(n13677) );
  NOR2_X1 U13659 ( .A1(n13678), .A2(n13679), .ZN(n13671) );
  INV_X1 U13660 ( .A(n13680), .ZN(n13679) );
  NAND2_X1 U13661 ( .A1(n13560), .A2(n13681), .ZN(n13680) );
  NAND2_X1 U13662 ( .A1(n13559), .A2(n13558), .ZN(n13681) );
  NOR2_X1 U13663 ( .A1(n8531), .A2(n8593), .ZN(n13560) );
  NOR2_X1 U13664 ( .A1(n13558), .A2(n13559), .ZN(n13678) );
  NOR2_X1 U13665 ( .A1(n13682), .A2(n13683), .ZN(n13559) );
  INV_X1 U13666 ( .A(n13684), .ZN(n13683) );
  NAND2_X1 U13667 ( .A1(n13556), .A2(n13685), .ZN(n13684) );
  NAND2_X1 U13668 ( .A1(n13686), .A2(n13553), .ZN(n13685) );
  NOR2_X1 U13669 ( .A1(n8531), .A2(n8583), .ZN(n13556) );
  NOR2_X1 U13670 ( .A1(n13553), .A2(n13686), .ZN(n13682) );
  INV_X1 U13671 ( .A(n13555), .ZN(n13686) );
  NAND2_X1 U13672 ( .A1(n13687), .A2(n13688), .ZN(n13555) );
  NAND2_X1 U13673 ( .A1(n13552), .A2(n13689), .ZN(n13688) );
  INV_X1 U13674 ( .A(n13690), .ZN(n13689) );
  NOR2_X1 U13675 ( .A1(n13551), .A2(n13550), .ZN(n13690) );
  NOR2_X1 U13676 ( .A1(n8531), .A2(n8580), .ZN(n13552) );
  NAND2_X1 U13677 ( .A1(n13550), .A2(n13551), .ZN(n13687) );
  NAND2_X1 U13678 ( .A1(n13691), .A2(n13692), .ZN(n13551) );
  NAND2_X1 U13679 ( .A1(n13548), .A2(n13693), .ZN(n13692) );
  INV_X1 U13680 ( .A(n13694), .ZN(n13693) );
  NOR2_X1 U13681 ( .A1(n13547), .A2(n13545), .ZN(n13694) );
  NOR2_X1 U13682 ( .A1(n8531), .A2(n8588), .ZN(n13548) );
  NAND2_X1 U13683 ( .A1(n13545), .A2(n13547), .ZN(n13691) );
  NAND2_X1 U13684 ( .A1(n13695), .A2(n13696), .ZN(n13547) );
  NAND2_X1 U13685 ( .A1(n13544), .A2(n13697), .ZN(n13696) );
  INV_X1 U13686 ( .A(n13698), .ZN(n13697) );
  NOR2_X1 U13687 ( .A1(n13543), .A2(n13542), .ZN(n13698) );
  NOR2_X1 U13688 ( .A1(n8531), .A2(n8551), .ZN(n13544) );
  NAND2_X1 U13689 ( .A1(n13542), .A2(n13543), .ZN(n13695) );
  NAND2_X1 U13690 ( .A1(n13699), .A2(n13700), .ZN(n13543) );
  NAND2_X1 U13691 ( .A1(n13540), .A2(n13701), .ZN(n13700) );
  NAND2_X1 U13692 ( .A1(n13539), .A2(n13537), .ZN(n13701) );
  NOR2_X1 U13693 ( .A1(n8531), .A2(n8563), .ZN(n13540) );
  INV_X1 U13694 ( .A(n13702), .ZN(n13699) );
  NOR2_X1 U13695 ( .A1(n13537), .A2(n13539), .ZN(n13702) );
  NOR2_X1 U13696 ( .A1(n13703), .A2(n13704), .ZN(n13539) );
  INV_X1 U13697 ( .A(n13705), .ZN(n13704) );
  NAND2_X1 U13698 ( .A1(n13536), .A2(n13706), .ZN(n13705) );
  NAND2_X1 U13699 ( .A1(n13535), .A2(n13534), .ZN(n13706) );
  NOR2_X1 U13700 ( .A1(n8531), .A2(n8548), .ZN(n13536) );
  NOR2_X1 U13701 ( .A1(n13534), .A2(n13535), .ZN(n13703) );
  INV_X1 U13702 ( .A(n13707), .ZN(n13535) );
  NAND2_X1 U13703 ( .A1(n13708), .A2(n13709), .ZN(n13707) );
  NAND2_X1 U13704 ( .A1(n13531), .A2(n13710), .ZN(n13709) );
  NAND2_X1 U13705 ( .A1(n13532), .A2(n13530), .ZN(n13710) );
  NOR2_X1 U13706 ( .A1(n8531), .A2(n8584), .ZN(n13531) );
  NAND2_X1 U13707 ( .A1(n13711), .A2(n13712), .ZN(n13708) );
  INV_X1 U13708 ( .A(n13532), .ZN(n13712) );
  NOR2_X1 U13709 ( .A1(n13713), .A2(n13714), .ZN(n13532) );
  INV_X1 U13710 ( .A(n13715), .ZN(n13714) );
  NAND2_X1 U13711 ( .A1(n13528), .A2(n13716), .ZN(n13715) );
  NAND2_X1 U13712 ( .A1(n13527), .A2(n13526), .ZN(n13716) );
  NOR2_X1 U13713 ( .A1(n8531), .A2(n8535), .ZN(n13528) );
  NOR2_X1 U13714 ( .A1(n13526), .A2(n13527), .ZN(n13713) );
  NOR2_X1 U13715 ( .A1(n13717), .A2(n13718), .ZN(n13527) );
  INV_X1 U13716 ( .A(n13719), .ZN(n13718) );
  NAND2_X1 U13717 ( .A1(n13523), .A2(n13720), .ZN(n13719) );
  NAND2_X1 U13718 ( .A1(n13524), .A2(n13522), .ZN(n13720) );
  NOR2_X1 U13719 ( .A1(n8531), .A2(n8568), .ZN(n13523) );
  NOR2_X1 U13720 ( .A1(n13522), .A2(n13524), .ZN(n13717) );
  NOR2_X1 U13721 ( .A1(n13721), .A2(n13722), .ZN(n13524) );
  INV_X1 U13722 ( .A(n13723), .ZN(n13722) );
  NAND2_X1 U13723 ( .A1(n13519), .A2(n13724), .ZN(n13723) );
  NAND2_X1 U13724 ( .A1(n13520), .A2(n13518), .ZN(n13724) );
  NOR2_X1 U13725 ( .A1(n8531), .A2(n8574), .ZN(n13519) );
  NOR2_X1 U13726 ( .A1(n13518), .A2(n13520), .ZN(n13721) );
  NOR2_X1 U13727 ( .A1(n13725), .A2(n13726), .ZN(n13520) );
  INV_X1 U13728 ( .A(n13727), .ZN(n13726) );
  NAND2_X1 U13729 ( .A1(n13515), .A2(n13728), .ZN(n13727) );
  NAND2_X1 U13730 ( .A1(n13516), .A2(n13514), .ZN(n13728) );
  NOR2_X1 U13731 ( .A1(n8531), .A2(n8565), .ZN(n13515) );
  NOR2_X1 U13732 ( .A1(n13514), .A2(n13516), .ZN(n13725) );
  NOR2_X1 U13733 ( .A1(n13729), .A2(n13730), .ZN(n13516) );
  INV_X1 U13734 ( .A(n13731), .ZN(n13730) );
  NAND2_X1 U13735 ( .A1(n13509), .A2(n13732), .ZN(n13731) );
  NAND2_X1 U13736 ( .A1(n13512), .A2(n13511), .ZN(n13732) );
  NOR2_X1 U13737 ( .A1(n8531), .A2(n8567), .ZN(n13509) );
  NOR2_X1 U13738 ( .A1(n13511), .A2(n13512), .ZN(n13729) );
  INV_X1 U13739 ( .A(n13733), .ZN(n13512) );
  NAND2_X1 U13740 ( .A1(n13734), .A2(n13735), .ZN(n13733) );
  NAND2_X1 U13741 ( .A1(n13504), .A2(n13736), .ZN(n13735) );
  NAND2_X1 U13742 ( .A1(n8624), .A2(n13737), .ZN(n13736) );
  NAND2_X1 U13743 ( .A1(n8561), .A2(n8585), .ZN(n13737) );
  NAND2_X1 U13744 ( .A1(n13739), .A2(n13740), .ZN(n13734) );
  NAND2_X1 U13745 ( .A1(n8630), .A2(n13741), .ZN(n13740) );
  NAND2_X1 U13746 ( .A1(n8539), .A2(n8553), .ZN(n13741) );
  NAND3_X1 U13747 ( .A1(n13220), .A2(n8537), .A3(n13504), .ZN(n13511) );
  INV_X1 U13748 ( .A(n8531), .ZN(n13220) );
  XOR2_X1 U13749 ( .A(d_13_), .B(c_13_), .Z(n13743) );
  XOR2_X1 U13750 ( .A(n13744), .B(n13745), .Z(n13514) );
  XNOR2_X1 U13751 ( .A(n13746), .B(n13747), .ZN(n13745) );
  XOR2_X1 U13752 ( .A(n13748), .B(n13749), .Z(n13518) );
  XNOR2_X1 U13753 ( .A(n13750), .B(n13751), .ZN(n13748) );
  XOR2_X1 U13754 ( .A(n13752), .B(n13753), .Z(n13522) );
  XNOR2_X1 U13755 ( .A(n13754), .B(n13755), .ZN(n13752) );
  XOR2_X1 U13756 ( .A(n13756), .B(n13757), .Z(n13526) );
  XNOR2_X1 U13757 ( .A(n13758), .B(n13759), .ZN(n13756) );
  INV_X1 U13758 ( .A(n13530), .ZN(n13711) );
  XOR2_X1 U13759 ( .A(n13760), .B(n13761), .Z(n13530) );
  XOR2_X1 U13760 ( .A(n13762), .B(n13763), .Z(n13760) );
  NAND2_X1 U13761 ( .A1(n13504), .A2(n9121), .ZN(n13762) );
  XOR2_X1 U13762 ( .A(n13764), .B(n13765), .Z(n13534) );
  XNOR2_X1 U13763 ( .A(n13766), .B(n13767), .ZN(n13764) );
  NOR2_X1 U13764 ( .A1(n8584), .A2(n8553), .ZN(n13767) );
  XOR2_X1 U13765 ( .A(n13768), .B(n13769), .Z(n13537) );
  XNOR2_X1 U13766 ( .A(n13770), .B(n13771), .ZN(n13768) );
  NOR2_X1 U13767 ( .A1(n8548), .A2(n8553), .ZN(n13771) );
  XNOR2_X1 U13768 ( .A(n13772), .B(n13773), .ZN(n13542) );
  XNOR2_X1 U13769 ( .A(n13774), .B(n13775), .ZN(n13772) );
  NOR2_X1 U13770 ( .A1(n9094), .A2(n8553), .ZN(n13775) );
  XNOR2_X1 U13771 ( .A(n13776), .B(n13777), .ZN(n13545) );
  XNOR2_X1 U13772 ( .A(n13778), .B(n13779), .ZN(n13776) );
  NOR2_X1 U13773 ( .A1(n8551), .A2(n8553), .ZN(n13779) );
  XNOR2_X1 U13774 ( .A(n13780), .B(n13781), .ZN(n13550) );
  XNOR2_X1 U13775 ( .A(n13782), .B(n13783), .ZN(n13780) );
  NOR2_X1 U13776 ( .A1(n8588), .A2(n8553), .ZN(n13783) );
  XOR2_X1 U13777 ( .A(n13784), .B(n13785), .Z(n13553) );
  XNOR2_X1 U13778 ( .A(n13786), .B(n13787), .ZN(n13784) );
  NOR2_X1 U13779 ( .A1(n8580), .A2(n8553), .ZN(n13787) );
  XOR2_X1 U13780 ( .A(n13788), .B(n13789), .Z(n13558) );
  XNOR2_X1 U13781 ( .A(n13790), .B(n13791), .ZN(n13788) );
  NOR2_X1 U13782 ( .A1(n9061), .A2(n8553), .ZN(n13791) );
  XNOR2_X1 U13783 ( .A(n13792), .B(n13793), .ZN(n13566) );
  XOR2_X1 U13784 ( .A(n13794), .B(n13795), .Z(n13793) );
  XNOR2_X1 U13785 ( .A(n13796), .B(n13797), .ZN(n13569) );
  XNOR2_X1 U13786 ( .A(n13798), .B(n13799), .ZN(n13796) );
  XNOR2_X1 U13787 ( .A(n13800), .B(n13801), .ZN(n13574) );
  XNOR2_X1 U13788 ( .A(n13802), .B(n13803), .ZN(n13800) );
  XNOR2_X1 U13789 ( .A(n13804), .B(n13805), .ZN(n13577) );
  XNOR2_X1 U13790 ( .A(n13806), .B(n13807), .ZN(n13804) );
  XNOR2_X1 U13791 ( .A(n13808), .B(n13809), .ZN(n13582) );
  XOR2_X1 U13792 ( .A(n13810), .B(n13811), .Z(n13808) );
  NAND2_X1 U13793 ( .A1(n13504), .A2(n9313), .ZN(n13810) );
  XNOR2_X1 U13794 ( .A(n13812), .B(n13813), .ZN(n13585) );
  NAND2_X1 U13795 ( .A1(n13814), .A2(n13815), .ZN(n13812) );
  XOR2_X1 U13796 ( .A(n13816), .B(n13817), .Z(n13407) );
  XNOR2_X1 U13797 ( .A(n13818), .B(n13819), .ZN(n13817) );
  XNOR2_X1 U13798 ( .A(n13820), .B(n13821), .ZN(n13589) );
  NAND2_X1 U13799 ( .A1(n13822), .A2(n13823), .ZN(n13820) );
  XNOR2_X1 U13800 ( .A(n13824), .B(n13825), .ZN(n13593) );
  XNOR2_X1 U13801 ( .A(n13826), .B(n13827), .ZN(n13825) );
  XOR2_X1 U13802 ( .A(n13828), .B(n13829), .Z(n13390) );
  NAND2_X1 U13803 ( .A1(n13830), .A2(n13831), .ZN(n13828) );
  XOR2_X1 U13804 ( .A(n13832), .B(n13833), .Z(n13383) );
  XNOR2_X1 U13805 ( .A(n13834), .B(n13835), .ZN(n13833) );
  XNOR2_X1 U13806 ( .A(n13836), .B(n13837), .ZN(n13375) );
  NAND2_X1 U13807 ( .A1(n13838), .A2(n13839), .ZN(n13836) );
  XOR2_X1 U13808 ( .A(n13840), .B(n13841), .Z(n13366) );
  XNOR2_X1 U13809 ( .A(n13842), .B(n13843), .ZN(n13841) );
  XNOR2_X1 U13810 ( .A(n13844), .B(n13845), .ZN(n13358) );
  NAND2_X1 U13811 ( .A1(n13846), .A2(n13847), .ZN(n13844) );
  XNOR2_X1 U13812 ( .A(n13848), .B(n13849), .ZN(n13597) );
  XOR2_X1 U13813 ( .A(n13850), .B(n13851), .Z(n13849) );
  NAND2_X1 U13814 ( .A1(n13504), .A2(n9268), .ZN(n13851) );
  XOR2_X1 U13815 ( .A(n13852), .B(n13853), .Z(n13601) );
  NAND2_X1 U13816 ( .A1(n13854), .A2(n13855), .ZN(n13852) );
  XOR2_X1 U13817 ( .A(n13856), .B(n13347), .Z(n13605) );
  XNOR2_X1 U13818 ( .A(n13857), .B(n13858), .ZN(n13347) );
  XNOR2_X1 U13819 ( .A(n13859), .B(n13860), .ZN(n8859) );
  NAND2_X1 U13820 ( .A1(n8867), .A2(n8866), .ZN(n8865) );
  NOR2_X1 U13821 ( .A1(n13861), .A2(n8900), .ZN(n8866) );
  INV_X1 U13822 ( .A(n13862), .ZN(n13861) );
  NAND2_X1 U13823 ( .A1(n13863), .A2(n13864), .ZN(n13862) );
  NOR2_X1 U13824 ( .A1(n13860), .A2(n13859), .ZN(n8867) );
  INV_X1 U13825 ( .A(n13865), .ZN(n13859) );
  NAND2_X1 U13826 ( .A1(n13866), .A2(n13867), .ZN(n13865) );
  NAND2_X1 U13827 ( .A1(n13858), .A2(n13868), .ZN(n13867) );
  NAND2_X1 U13828 ( .A1(n13869), .A2(n13348), .ZN(n13868) );
  INV_X1 U13829 ( .A(n13856), .ZN(n13348) );
  INV_X1 U13830 ( .A(n13857), .ZN(n13869) );
  NOR2_X1 U13831 ( .A1(n8553), .A2(n8972), .ZN(n13858) );
  NAND2_X1 U13832 ( .A1(n13856), .A2(n13857), .ZN(n13866) );
  NAND2_X1 U13833 ( .A1(n13854), .A2(n13870), .ZN(n13857) );
  NAND2_X1 U13834 ( .A1(n13853), .A2(n13855), .ZN(n13870) );
  NAND2_X1 U13835 ( .A1(n13871), .A2(n13872), .ZN(n13855) );
  NAND2_X1 U13836 ( .A1(n13504), .A2(n9263), .ZN(n13872) );
  XNOR2_X1 U13837 ( .A(n13873), .B(n13874), .ZN(n13853) );
  XOR2_X1 U13838 ( .A(n13875), .B(n13876), .Z(n13874) );
  NAND2_X1 U13839 ( .A1(n9268), .A2(n13739), .ZN(n13876) );
  INV_X1 U13840 ( .A(n13877), .ZN(n13854) );
  NOR2_X1 U13841 ( .A1(n8589), .A2(n13871), .ZN(n13877) );
  NOR2_X1 U13842 ( .A1(n13878), .A2(n13879), .ZN(n13871) );
  NOR3_X1 U13843 ( .A1(n8982), .A2(n13880), .A3(n8553), .ZN(n13879) );
  NOR2_X1 U13844 ( .A1(n13850), .A2(n13848), .ZN(n13880) );
  INV_X1 U13845 ( .A(n13881), .ZN(n13878) );
  NAND2_X1 U13846 ( .A1(n13848), .A2(n13850), .ZN(n13881) );
  NAND2_X1 U13847 ( .A1(n13846), .A2(n13882), .ZN(n13850) );
  NAND2_X1 U13848 ( .A1(n13845), .A2(n13847), .ZN(n13882) );
  NAND2_X1 U13849 ( .A1(n13883), .A2(n13884), .ZN(n13847) );
  NAND2_X1 U13850 ( .A1(n13504), .A2(n9792), .ZN(n13883) );
  XNOR2_X1 U13851 ( .A(n13885), .B(n13886), .ZN(n13845) );
  XOR2_X1 U13852 ( .A(n13887), .B(n13888), .Z(n13886) );
  NAND2_X1 U13853 ( .A1(n9277), .A2(n13739), .ZN(n13888) );
  INV_X1 U13854 ( .A(n13889), .ZN(n13846) );
  NOR2_X1 U13855 ( .A1(n13884), .A2(n8527), .ZN(n13889) );
  NAND2_X1 U13856 ( .A1(n13890), .A2(n13891), .ZN(n13884) );
  NAND2_X1 U13857 ( .A1(n13840), .A2(n13892), .ZN(n13891) );
  NAND2_X1 U13858 ( .A1(n13843), .A2(n13842), .ZN(n13892) );
  XNOR2_X1 U13859 ( .A(n13893), .B(n13894), .ZN(n13840) );
  XOR2_X1 U13860 ( .A(n13895), .B(n13896), .Z(n13893) );
  NOR2_X1 U13861 ( .A1(n8561), .A2(n8564), .ZN(n13896) );
  INV_X1 U13862 ( .A(n13897), .ZN(n13890) );
  NOR2_X1 U13863 ( .A1(n13842), .A2(n13843), .ZN(n13897) );
  NOR2_X1 U13864 ( .A1(n8553), .A2(n8528), .ZN(n13843) );
  NAND2_X1 U13865 ( .A1(n13838), .A2(n13898), .ZN(n13842) );
  NAND2_X1 U13866 ( .A1(n13837), .A2(n13839), .ZN(n13898) );
  NAND2_X1 U13867 ( .A1(n13899), .A2(n13900), .ZN(n13839) );
  NAND2_X1 U13868 ( .A1(n13504), .A2(n10307), .ZN(n13899) );
  XNOR2_X1 U13869 ( .A(n13901), .B(n13902), .ZN(n13837) );
  XOR2_X1 U13870 ( .A(n13903), .B(n13904), .Z(n13902) );
  NAND2_X1 U13871 ( .A1(n9286), .A2(n13739), .ZN(n13904) );
  INV_X1 U13872 ( .A(n13905), .ZN(n13838) );
  NOR2_X1 U13873 ( .A1(n13900), .A2(n8564), .ZN(n13905) );
  NAND2_X1 U13874 ( .A1(n13906), .A2(n13907), .ZN(n13900) );
  NAND2_X1 U13875 ( .A1(n13832), .A2(n13908), .ZN(n13907) );
  NAND2_X1 U13876 ( .A1(n13835), .A2(n13834), .ZN(n13908) );
  XNOR2_X1 U13877 ( .A(n13909), .B(n13910), .ZN(n13832) );
  XOR2_X1 U13878 ( .A(n13911), .B(n13912), .Z(n13909) );
  NOR2_X1 U13879 ( .A1(n8561), .A2(n8544), .ZN(n13912) );
  INV_X1 U13880 ( .A(n13913), .ZN(n13906) );
  NOR2_X1 U13881 ( .A1(n13834), .A2(n13835), .ZN(n13913) );
  NOR2_X1 U13882 ( .A1(n8553), .A2(n8555), .ZN(n13835) );
  NAND2_X1 U13883 ( .A1(n13830), .A2(n13914), .ZN(n13834) );
  NAND2_X1 U13884 ( .A1(n13829), .A2(n13831), .ZN(n13914) );
  NAND2_X1 U13885 ( .A1(n13915), .A2(n13916), .ZN(n13831) );
  NAND2_X1 U13886 ( .A1(n13504), .A2(n8543), .ZN(n13915) );
  XOR2_X1 U13887 ( .A(n13917), .B(n13918), .Z(n13829) );
  XNOR2_X1 U13888 ( .A(n13919), .B(n13920), .ZN(n13918) );
  NAND2_X1 U13889 ( .A1(n9295), .A2(n13739), .ZN(n13920) );
  INV_X1 U13890 ( .A(n13921), .ZN(n13830) );
  NOR2_X1 U13891 ( .A1(n13916), .A2(n8544), .ZN(n13921) );
  NAND2_X1 U13892 ( .A1(n13922), .A2(n13923), .ZN(n13916) );
  NAND2_X1 U13893 ( .A1(n13824), .A2(n13924), .ZN(n13923) );
  NAND2_X1 U13894 ( .A1(n13827), .A2(n13826), .ZN(n13924) );
  XOR2_X1 U13895 ( .A(n13925), .B(n13926), .Z(n13824) );
  XNOR2_X1 U13896 ( .A(n13927), .B(n13928), .ZN(n13925) );
  NOR2_X1 U13897 ( .A1(n8561), .A2(n8594), .ZN(n13928) );
  INV_X1 U13898 ( .A(n13929), .ZN(n13922) );
  NOR2_X1 U13899 ( .A1(n13826), .A2(n13827), .ZN(n13929) );
  NOR2_X1 U13900 ( .A1(n8553), .A2(n8560), .ZN(n13827) );
  NAND2_X1 U13901 ( .A1(n13822), .A2(n13930), .ZN(n13826) );
  NAND2_X1 U13902 ( .A1(n13821), .A2(n13823), .ZN(n13930) );
  NAND2_X1 U13903 ( .A1(n13931), .A2(n13932), .ZN(n13823) );
  NAND2_X1 U13904 ( .A1(n13504), .A2(n10846), .ZN(n13931) );
  XOR2_X1 U13905 ( .A(n13933), .B(n13934), .Z(n13821) );
  XOR2_X1 U13906 ( .A(n13935), .B(n13936), .Z(n13933) );
  NOR2_X1 U13907 ( .A1(n8561), .A2(n8556), .ZN(n13936) );
  INV_X1 U13908 ( .A(n13937), .ZN(n13822) );
  NOR2_X1 U13909 ( .A1(n13932), .A2(n8594), .ZN(n13937) );
  NAND2_X1 U13910 ( .A1(n13938), .A2(n13939), .ZN(n13932) );
  NAND2_X1 U13911 ( .A1(n13816), .A2(n13940), .ZN(n13939) );
  NAND2_X1 U13912 ( .A1(n13819), .A2(n13818), .ZN(n13940) );
  XNOR2_X1 U13913 ( .A(n13941), .B(n13942), .ZN(n13816) );
  XNOR2_X1 U13914 ( .A(n13943), .B(n13944), .ZN(n13942) );
  NAND2_X1 U13915 ( .A1(n9209), .A2(n13739), .ZN(n13944) );
  INV_X1 U13916 ( .A(n13945), .ZN(n13938) );
  NOR2_X1 U13917 ( .A1(n13818), .A2(n13819), .ZN(n13945) );
  NOR2_X1 U13918 ( .A1(n13503), .A2(n8556), .ZN(n13819) );
  NAND2_X1 U13919 ( .A1(n13814), .A2(n13946), .ZN(n13818) );
  NAND2_X1 U13920 ( .A1(n13813), .A2(n13815), .ZN(n13946) );
  NAND2_X1 U13921 ( .A1(n13947), .A2(n13948), .ZN(n13815) );
  NAND2_X1 U13922 ( .A1(n13504), .A2(n9209), .ZN(n13948) );
  XOR2_X1 U13923 ( .A(n13949), .B(n13950), .Z(n13813) );
  XOR2_X1 U13924 ( .A(n13951), .B(n13952), .Z(n13949) );
  NOR2_X1 U13925 ( .A1(n8561), .A2(n8582), .ZN(n13952) );
  NAND2_X1 U13926 ( .A1(n9209), .A2(n13953), .ZN(n13814) );
  INV_X1 U13927 ( .A(n13947), .ZN(n13953) );
  NOR2_X1 U13928 ( .A1(n13954), .A2(n13955), .ZN(n13947) );
  NOR3_X1 U13929 ( .A1(n9031), .A2(n13956), .A3(n8553), .ZN(n13955) );
  INV_X1 U13930 ( .A(n13957), .ZN(n13956) );
  NAND2_X1 U13931 ( .A1(n13811), .A2(n13809), .ZN(n13957) );
  NOR2_X1 U13932 ( .A1(n13809), .A2(n13811), .ZN(n13954) );
  NOR2_X1 U13933 ( .A1(n13958), .A2(n13959), .ZN(n13811) );
  INV_X1 U13934 ( .A(n13960), .ZN(n13959) );
  NAND2_X1 U13935 ( .A1(n13807), .A2(n13961), .ZN(n13960) );
  NAND2_X1 U13936 ( .A1(n13806), .A2(n13805), .ZN(n13961) );
  NOR2_X1 U13937 ( .A1(n13503), .A2(n8591), .ZN(n13807) );
  NOR2_X1 U13938 ( .A1(n13805), .A2(n13806), .ZN(n13958) );
  NOR2_X1 U13939 ( .A1(n13962), .A2(n13963), .ZN(n13806) );
  INV_X1 U13940 ( .A(n13964), .ZN(n13963) );
  NAND2_X1 U13941 ( .A1(n13803), .A2(n13965), .ZN(n13964) );
  NAND2_X1 U13942 ( .A1(n13802), .A2(n13801), .ZN(n13965) );
  NOR2_X1 U13943 ( .A1(n13503), .A2(n8562), .ZN(n13803) );
  NOR2_X1 U13944 ( .A1(n13801), .A2(n13802), .ZN(n13962) );
  NOR2_X1 U13945 ( .A1(n13966), .A2(n13967), .ZN(n13802) );
  INV_X1 U13946 ( .A(n13968), .ZN(n13967) );
  NAND2_X1 U13947 ( .A1(n13799), .A2(n13969), .ZN(n13968) );
  NAND2_X1 U13948 ( .A1(n13797), .A2(n13798), .ZN(n13969) );
  NOR2_X1 U13949 ( .A1(n13503), .A2(n8545), .ZN(n13799) );
  NOR2_X1 U13950 ( .A1(n13797), .A2(n13798), .ZN(n13966) );
  NOR2_X1 U13951 ( .A1(n13970), .A2(n13971), .ZN(n13798) );
  NOR2_X1 U13952 ( .A1(n13795), .A2(n13972), .ZN(n13971) );
  NOR2_X1 U13953 ( .A1(n13794), .A2(n13792), .ZN(n13972) );
  NAND2_X1 U13954 ( .A1(n13504), .A2(n9331), .ZN(n13795) );
  INV_X1 U13955 ( .A(n13973), .ZN(n13970) );
  NAND2_X1 U13956 ( .A1(n13792), .A2(n13794), .ZN(n13973) );
  NAND2_X1 U13957 ( .A1(n13974), .A2(n13975), .ZN(n13794) );
  NAND2_X1 U13958 ( .A1(n13676), .A2(n13976), .ZN(n13975) );
  NAND2_X1 U13959 ( .A1(n13675), .A2(n13673), .ZN(n13976) );
  NOR2_X1 U13960 ( .A1(n13503), .A2(n8593), .ZN(n13676) );
  INV_X1 U13961 ( .A(n13977), .ZN(n13974) );
  NOR2_X1 U13962 ( .A1(n13673), .A2(n13675), .ZN(n13977) );
  NOR2_X1 U13963 ( .A1(n13978), .A2(n13979), .ZN(n13675) );
  NOR3_X1 U13964 ( .A1(n9061), .A2(n13980), .A3(n8553), .ZN(n13979) );
  INV_X1 U13965 ( .A(n13981), .ZN(n13980) );
  NAND2_X1 U13966 ( .A1(n13789), .A2(n13790), .ZN(n13981) );
  NOR2_X1 U13967 ( .A1(n13789), .A2(n13790), .ZN(n13978) );
  NOR2_X1 U13968 ( .A1(n13982), .A2(n13983), .ZN(n13790) );
  INV_X1 U13969 ( .A(n13984), .ZN(n13983) );
  NAND3_X1 U13970 ( .A1(n9070), .A2(n13985), .A3(n13504), .ZN(n13984) );
  NAND2_X1 U13971 ( .A1(n13785), .A2(n13786), .ZN(n13985) );
  NOR2_X1 U13972 ( .A1(n13785), .A2(n13786), .ZN(n13982) );
  NOR2_X1 U13973 ( .A1(n13986), .A2(n13987), .ZN(n13786) );
  INV_X1 U13974 ( .A(n13988), .ZN(n13987) );
  NAND3_X1 U13975 ( .A1(n9080), .A2(n13989), .A3(n13504), .ZN(n13988) );
  NAND2_X1 U13976 ( .A1(n13782), .A2(n13781), .ZN(n13989) );
  NOR2_X1 U13977 ( .A1(n13781), .A2(n13782), .ZN(n13986) );
  NOR2_X1 U13978 ( .A1(n13990), .A2(n13991), .ZN(n13782) );
  NOR3_X1 U13979 ( .A1(n8551), .A2(n13992), .A3(n8553), .ZN(n13991) );
  INV_X1 U13980 ( .A(n13993), .ZN(n13992) );
  NAND2_X1 U13981 ( .A1(n13777), .A2(n13778), .ZN(n13993) );
  NOR2_X1 U13982 ( .A1(n13777), .A2(n13778), .ZN(n13990) );
  NOR2_X1 U13983 ( .A1(n13994), .A2(n13995), .ZN(n13778) );
  INV_X1 U13984 ( .A(n13996), .ZN(n13995) );
  NAND3_X1 U13985 ( .A1(n9098), .A2(n13997), .A3(n13504), .ZN(n13996) );
  NAND2_X1 U13986 ( .A1(n13774), .A2(n13773), .ZN(n13997) );
  NOR2_X1 U13987 ( .A1(n13773), .A2(n13774), .ZN(n13994) );
  NOR2_X1 U13988 ( .A1(n13998), .A2(n13999), .ZN(n13774) );
  NOR3_X1 U13989 ( .A1(n8548), .A2(n14000), .A3(n8553), .ZN(n13999) );
  INV_X1 U13990 ( .A(n14001), .ZN(n14000) );
  NAND2_X1 U13991 ( .A1(n13769), .A2(n13770), .ZN(n14001) );
  NOR2_X1 U13992 ( .A1(n13769), .A2(n13770), .ZN(n13998) );
  NOR2_X1 U13993 ( .A1(n14002), .A2(n14003), .ZN(n13770) );
  INV_X1 U13994 ( .A(n14004), .ZN(n14003) );
  NAND3_X1 U13995 ( .A1(n9112), .A2(n14005), .A3(n13504), .ZN(n14004) );
  NAND2_X1 U13996 ( .A1(n13766), .A2(n13765), .ZN(n14005) );
  NOR2_X1 U13997 ( .A1(n13765), .A2(n13766), .ZN(n14002) );
  NOR2_X1 U13998 ( .A1(n14006), .A2(n14007), .ZN(n13766) );
  INV_X1 U13999 ( .A(n14008), .ZN(n14007) );
  NAND3_X1 U14000 ( .A1(n9121), .A2(n14009), .A3(n13504), .ZN(n14008) );
  NAND2_X1 U14001 ( .A1(n13761), .A2(n13763), .ZN(n14009) );
  NOR2_X1 U14002 ( .A1(n13761), .A2(n13763), .ZN(n14006) );
  NOR2_X1 U14003 ( .A1(n14010), .A2(n14011), .ZN(n13763) );
  INV_X1 U14004 ( .A(n14012), .ZN(n14011) );
  NAND2_X1 U14005 ( .A1(n13759), .A2(n14013), .ZN(n14012) );
  NAND2_X1 U14006 ( .A1(n13758), .A2(n13757), .ZN(n14013) );
  NOR2_X1 U14007 ( .A1(n13503), .A2(n8568), .ZN(n13759) );
  NOR2_X1 U14008 ( .A1(n13757), .A2(n13758), .ZN(n14010) );
  NOR2_X1 U14009 ( .A1(n14014), .A2(n14015), .ZN(n13758) );
  INV_X1 U14010 ( .A(n14016), .ZN(n14015) );
  NAND2_X1 U14011 ( .A1(n13754), .A2(n14017), .ZN(n14016) );
  NAND2_X1 U14012 ( .A1(n13753), .A2(n13755), .ZN(n14017) );
  NOR2_X1 U14013 ( .A1(n13503), .A2(n8574), .ZN(n13754) );
  NOR2_X1 U14014 ( .A1(n13753), .A2(n13755), .ZN(n14014) );
  NOR2_X1 U14015 ( .A1(n14018), .A2(n14019), .ZN(n13755) );
  INV_X1 U14016 ( .A(n14020), .ZN(n14019) );
  NAND2_X1 U14017 ( .A1(n13750), .A2(n14021), .ZN(n14020) );
  NAND2_X1 U14018 ( .A1(n13751), .A2(n13749), .ZN(n14021) );
  NOR2_X1 U14019 ( .A1(n13503), .A2(n8565), .ZN(n13750) );
  NOR2_X1 U14020 ( .A1(n13749), .A2(n13751), .ZN(n14018) );
  NOR2_X1 U14021 ( .A1(n14022), .A2(n14023), .ZN(n13751) );
  INV_X1 U14022 ( .A(n14024), .ZN(n14023) );
  NAND2_X1 U14023 ( .A1(n13744), .A2(n14025), .ZN(n14024) );
  NAND2_X1 U14024 ( .A1(n13747), .A2(n13746), .ZN(n14025) );
  NOR2_X1 U14025 ( .A1(n13503), .A2(n8567), .ZN(n13744) );
  NOR2_X1 U14026 ( .A1(n13746), .A2(n13747), .ZN(n14022) );
  INV_X1 U14027 ( .A(n14026), .ZN(n13747) );
  NAND2_X1 U14028 ( .A1(n14027), .A2(n14028), .ZN(n14026) );
  NAND2_X1 U14029 ( .A1(n13739), .A2(n14029), .ZN(n14028) );
  NAND2_X1 U14030 ( .A1(n8624), .A2(n14030), .ZN(n14029) );
  NAND2_X1 U14031 ( .A1(n8526), .A2(n8585), .ZN(n14030) );
  NAND2_X1 U14032 ( .A1(n14031), .A2(n14032), .ZN(n14027) );
  NAND2_X1 U14033 ( .A1(n8630), .A2(n14033), .ZN(n14032) );
  NAND2_X1 U14034 ( .A1(n8539), .A2(n8561), .ZN(n14033) );
  NAND3_X1 U14035 ( .A1(n13739), .A2(n8537), .A3(n13504), .ZN(n13746) );
  INV_X1 U14036 ( .A(n13503), .ZN(n13504) );
  XNOR2_X1 U14037 ( .A(n14034), .B(n14035), .ZN(n13503) );
  XOR2_X1 U14038 ( .A(d_12_), .B(c_12_), .Z(n14035) );
  XOR2_X1 U14039 ( .A(n14036), .B(n14037), .Z(n13749) );
  XNOR2_X1 U14040 ( .A(n14038), .B(n14039), .ZN(n14037) );
  XOR2_X1 U14041 ( .A(n14040), .B(n14041), .Z(n13753) );
  XNOR2_X1 U14042 ( .A(n14042), .B(n14043), .ZN(n14040) );
  XOR2_X1 U14043 ( .A(n14044), .B(n14045), .Z(n13757) );
  XNOR2_X1 U14044 ( .A(n14046), .B(n14047), .ZN(n14044) );
  XOR2_X1 U14045 ( .A(n14048), .B(n14049), .Z(n13761) );
  XNOR2_X1 U14046 ( .A(n14050), .B(n14051), .ZN(n14048) );
  XOR2_X1 U14047 ( .A(n14052), .B(n14053), .Z(n13765) );
  XNOR2_X1 U14048 ( .A(n14054), .B(n14055), .ZN(n14052) );
  XOR2_X1 U14049 ( .A(n14056), .B(n14057), .Z(n13769) );
  XNOR2_X1 U14050 ( .A(n14058), .B(n14059), .ZN(n14056) );
  XOR2_X1 U14051 ( .A(n14060), .B(n14061), .Z(n13773) );
  XNOR2_X1 U14052 ( .A(n14062), .B(n14063), .ZN(n14060) );
  XNOR2_X1 U14053 ( .A(n14064), .B(n14065), .ZN(n13777) );
  XOR2_X1 U14054 ( .A(n14066), .B(n14067), .Z(n14065) );
  XNOR2_X1 U14055 ( .A(n14068), .B(n14069), .ZN(n13781) );
  XOR2_X1 U14056 ( .A(n14070), .B(n14071), .Z(n14068) );
  XNOR2_X1 U14057 ( .A(n14072), .B(n14073), .ZN(n13785) );
  XNOR2_X1 U14058 ( .A(n14074), .B(n14075), .ZN(n14073) );
  XOR2_X1 U14059 ( .A(n14076), .B(n14077), .Z(n13789) );
  XNOR2_X1 U14060 ( .A(n14078), .B(n14079), .ZN(n14076) );
  XOR2_X1 U14061 ( .A(n14080), .B(n14081), .Z(n13673) );
  NAND2_X1 U14062 ( .A1(n14082), .A2(n14083), .ZN(n14080) );
  XNOR2_X1 U14063 ( .A(n14084), .B(n14085), .ZN(n13792) );
  XOR2_X1 U14064 ( .A(n14086), .B(n14087), .Z(n14085) );
  NAND2_X1 U14065 ( .A1(n10722), .A2(n13739), .ZN(n14087) );
  XOR2_X1 U14066 ( .A(n14088), .B(n14089), .Z(n13797) );
  XOR2_X1 U14067 ( .A(n14090), .B(n14091), .Z(n14089) );
  NAND2_X1 U14068 ( .A1(n9331), .A2(n13739), .ZN(n14091) );
  XNOR2_X1 U14069 ( .A(n14092), .B(n14093), .ZN(n13801) );
  XOR2_X1 U14070 ( .A(n14094), .B(n14095), .Z(n14092) );
  NOR2_X1 U14071 ( .A1(n8561), .A2(n8545), .ZN(n14095) );
  XOR2_X1 U14072 ( .A(n14096), .B(n14097), .Z(n13805) );
  XOR2_X1 U14073 ( .A(n14098), .B(n14099), .Z(n14097) );
  NAND2_X1 U14074 ( .A1(n9322), .A2(n13739), .ZN(n14099) );
  XOR2_X1 U14075 ( .A(n14100), .B(n14101), .Z(n13809) );
  XOR2_X1 U14076 ( .A(n14102), .B(n14103), .Z(n14101) );
  NAND2_X1 U14077 ( .A1(n9721), .A2(n13739), .ZN(n14103) );
  XOR2_X1 U14078 ( .A(n14104), .B(n14105), .Z(n13848) );
  XOR2_X1 U14079 ( .A(n14106), .B(n14107), .Z(n14104) );
  NOR2_X1 U14080 ( .A1(n8561), .A2(n8527), .ZN(n14107) );
  XOR2_X1 U14081 ( .A(n14108), .B(n14109), .Z(n13856) );
  XOR2_X1 U14082 ( .A(n14110), .B(n14111), .Z(n14108) );
  NOR2_X1 U14083 ( .A1(n8561), .A2(n8589), .ZN(n14111) );
  XNOR2_X1 U14084 ( .A(n14112), .B(n14113), .ZN(n13860) );
  XNOR2_X1 U14085 ( .A(n14114), .B(n14115), .ZN(n14113) );
  NAND2_X1 U14086 ( .A1(n13739), .A2(n8872), .ZN(n14115) );
  NOR2_X1 U14087 ( .A1(n13863), .A2(n13864), .ZN(n8900) );
  NOR2_X1 U14088 ( .A1(n14116), .A2(n14117), .ZN(n13864) );
  INV_X1 U14089 ( .A(n14118), .ZN(n14117) );
  NAND3_X1 U14090 ( .A1(n8592), .A2(n14119), .A3(n13739), .ZN(n14118) );
  NAND2_X1 U14091 ( .A1(n14114), .A2(n14112), .ZN(n14119) );
  NOR2_X1 U14092 ( .A1(n14112), .A2(n14114), .ZN(n14116) );
  NOR2_X1 U14093 ( .A1(n14120), .A2(n14121), .ZN(n14114) );
  NOR3_X1 U14094 ( .A1(n13738), .A2(n14122), .A3(n8589), .ZN(n14121) );
  NOR2_X1 U14095 ( .A1(n14110), .A2(n14109), .ZN(n14122) );
  INV_X1 U14096 ( .A(n14123), .ZN(n14120) );
  NAND2_X1 U14097 ( .A1(n14109), .A2(n14110), .ZN(n14123) );
  NAND2_X1 U14098 ( .A1(n14124), .A2(n14125), .ZN(n14110) );
  INV_X1 U14099 ( .A(n14126), .ZN(n14125) );
  NOR3_X1 U14100 ( .A1(n13738), .A2(n14127), .A3(n8552), .ZN(n14126) );
  NOR2_X1 U14101 ( .A1(n13875), .A2(n13873), .ZN(n14127) );
  NAND2_X1 U14102 ( .A1(n13873), .A2(n13875), .ZN(n14124) );
  NAND2_X1 U14103 ( .A1(n14128), .A2(n14129), .ZN(n13875) );
  NAND3_X1 U14104 ( .A1(n13739), .A2(n14130), .A3(n9792), .ZN(n14129) );
  INV_X1 U14105 ( .A(n14131), .ZN(n14130) );
  NOR2_X1 U14106 ( .A1(n14106), .A2(n14105), .ZN(n14131) );
  NAND2_X1 U14107 ( .A1(n14105), .A2(n14106), .ZN(n14128) );
  NAND2_X1 U14108 ( .A1(n14132), .A2(n14133), .ZN(n14106) );
  NAND3_X1 U14109 ( .A1(n13739), .A2(n14134), .A3(n9277), .ZN(n14133) );
  INV_X1 U14110 ( .A(n14135), .ZN(n14134) );
  NOR2_X1 U14111 ( .A1(n13887), .A2(n13885), .ZN(n14135) );
  NAND2_X1 U14112 ( .A1(n13885), .A2(n13887), .ZN(n14132) );
  NAND2_X1 U14113 ( .A1(n14136), .A2(n14137), .ZN(n13887) );
  NAND3_X1 U14114 ( .A1(n13739), .A2(n14138), .A3(n10307), .ZN(n14137) );
  INV_X1 U14115 ( .A(n14139), .ZN(n14138) );
  NOR2_X1 U14116 ( .A1(n13895), .A2(n13894), .ZN(n14139) );
  NAND2_X1 U14117 ( .A1(n13894), .A2(n13895), .ZN(n14136) );
  NAND2_X1 U14118 ( .A1(n14140), .A2(n14141), .ZN(n13895) );
  INV_X1 U14119 ( .A(n14142), .ZN(n14141) );
  NOR3_X1 U14120 ( .A1(n13738), .A2(n14143), .A3(n8555), .ZN(n14142) );
  NOR2_X1 U14121 ( .A1(n13903), .A2(n13901), .ZN(n14143) );
  NAND2_X1 U14122 ( .A1(n13901), .A2(n13903), .ZN(n14140) );
  NAND2_X1 U14123 ( .A1(n14144), .A2(n14145), .ZN(n13903) );
  NAND3_X1 U14124 ( .A1(n13739), .A2(n14146), .A3(n8543), .ZN(n14145) );
  INV_X1 U14125 ( .A(n14147), .ZN(n14146) );
  NOR2_X1 U14126 ( .A1(n13911), .A2(n13910), .ZN(n14147) );
  NAND2_X1 U14127 ( .A1(n13910), .A2(n13911), .ZN(n14144) );
  NAND2_X1 U14128 ( .A1(n14148), .A2(n14149), .ZN(n13911) );
  NAND3_X1 U14129 ( .A1(n13739), .A2(n14150), .A3(n9295), .ZN(n14149) );
  NAND2_X1 U14130 ( .A1(n13919), .A2(n13917), .ZN(n14150) );
  INV_X1 U14131 ( .A(n14151), .ZN(n14148) );
  NOR2_X1 U14132 ( .A1(n13917), .A2(n13919), .ZN(n14151) );
  NOR2_X1 U14133 ( .A1(n14152), .A2(n14153), .ZN(n13919) );
  INV_X1 U14134 ( .A(n14154), .ZN(n14153) );
  NAND3_X1 U14135 ( .A1(n13739), .A2(n14155), .A3(n10846), .ZN(n14154) );
  NAND2_X1 U14136 ( .A1(n13927), .A2(n13926), .ZN(n14155) );
  NOR2_X1 U14137 ( .A1(n13926), .A2(n13927), .ZN(n14152) );
  NOR2_X1 U14138 ( .A1(n14156), .A2(n14157), .ZN(n13927) );
  NOR3_X1 U14139 ( .A1(n13738), .A2(n14158), .A3(n8556), .ZN(n14157) );
  NOR2_X1 U14140 ( .A1(n13935), .A2(n13934), .ZN(n14158) );
  INV_X1 U14141 ( .A(n14159), .ZN(n14156) );
  NAND2_X1 U14142 ( .A1(n13934), .A2(n13935), .ZN(n14159) );
  NAND2_X1 U14143 ( .A1(n14160), .A2(n14161), .ZN(n13935) );
  NAND3_X1 U14144 ( .A1(n13739), .A2(n14162), .A3(n9209), .ZN(n14161) );
  NAND2_X1 U14145 ( .A1(n13943), .A2(n13941), .ZN(n14162) );
  INV_X1 U14146 ( .A(n14163), .ZN(n14160) );
  NOR2_X1 U14147 ( .A1(n13941), .A2(n13943), .ZN(n14163) );
  NOR2_X1 U14148 ( .A1(n14164), .A2(n14165), .ZN(n13943) );
  NOR3_X1 U14149 ( .A1(n13738), .A2(n14166), .A3(n8582), .ZN(n14165) );
  NOR2_X1 U14150 ( .A1(n13951), .A2(n13950), .ZN(n14166) );
  INV_X1 U14151 ( .A(n14167), .ZN(n14164) );
  NAND2_X1 U14152 ( .A1(n13950), .A2(n13951), .ZN(n14167) );
  NAND2_X1 U14153 ( .A1(n14168), .A2(n14169), .ZN(n13951) );
  INV_X1 U14154 ( .A(n14170), .ZN(n14169) );
  NOR3_X1 U14155 ( .A1(n13738), .A2(n14171), .A3(n8591), .ZN(n14170) );
  NOR2_X1 U14156 ( .A1(n14102), .A2(n14100), .ZN(n14171) );
  NAND2_X1 U14157 ( .A1(n14100), .A2(n14102), .ZN(n14168) );
  NAND2_X1 U14158 ( .A1(n14172), .A2(n14173), .ZN(n14102) );
  INV_X1 U14159 ( .A(n14174), .ZN(n14173) );
  NOR3_X1 U14160 ( .A1(n13738), .A2(n14175), .A3(n8562), .ZN(n14174) );
  NOR2_X1 U14161 ( .A1(n14098), .A2(n14096), .ZN(n14175) );
  NAND2_X1 U14162 ( .A1(n14096), .A2(n14098), .ZN(n14172) );
  NAND2_X1 U14163 ( .A1(n14176), .A2(n14177), .ZN(n14098) );
  NAND3_X1 U14164 ( .A1(n13739), .A2(n14178), .A3(n10222), .ZN(n14177) );
  INV_X1 U14165 ( .A(n14179), .ZN(n14178) );
  NOR2_X1 U14166 ( .A1(n14094), .A2(n14093), .ZN(n14179) );
  NAND2_X1 U14167 ( .A1(n14093), .A2(n14094), .ZN(n14176) );
  NAND2_X1 U14168 ( .A1(n14180), .A2(n14181), .ZN(n14094) );
  INV_X1 U14169 ( .A(n14182), .ZN(n14181) );
  NOR3_X1 U14170 ( .A1(n13738), .A2(n14183), .A3(n8569), .ZN(n14182) );
  NOR2_X1 U14171 ( .A1(n14090), .A2(n14088), .ZN(n14183) );
  NAND2_X1 U14172 ( .A1(n14088), .A2(n14090), .ZN(n14180) );
  NAND2_X1 U14173 ( .A1(n14184), .A2(n14185), .ZN(n14090) );
  NAND3_X1 U14174 ( .A1(n13739), .A2(n14186), .A3(n10722), .ZN(n14185) );
  INV_X1 U14175 ( .A(n14187), .ZN(n14186) );
  NOR2_X1 U14176 ( .A1(n14086), .A2(n14084), .ZN(n14187) );
  NAND2_X1 U14177 ( .A1(n14084), .A2(n14086), .ZN(n14184) );
  NAND2_X1 U14178 ( .A1(n14082), .A2(n14188), .ZN(n14086) );
  NAND2_X1 U14179 ( .A1(n14081), .A2(n14083), .ZN(n14188) );
  NAND2_X1 U14180 ( .A1(n14189), .A2(n14190), .ZN(n14083) );
  NAND2_X1 U14181 ( .A1(n9340), .A2(n13739), .ZN(n14190) );
  XNOR2_X1 U14182 ( .A(n14191), .B(n14192), .ZN(n14081) );
  XOR2_X1 U14183 ( .A(n14193), .B(n14194), .Z(n14192) );
  NAND2_X1 U14184 ( .A1(n9340), .A2(n14195), .ZN(n14082) );
  INV_X1 U14185 ( .A(n14189), .ZN(n14195) );
  NOR2_X1 U14186 ( .A1(n14196), .A2(n14197), .ZN(n14189) );
  INV_X1 U14187 ( .A(n14198), .ZN(n14197) );
  NAND2_X1 U14188 ( .A1(n14079), .A2(n14199), .ZN(n14198) );
  NAND2_X1 U14189 ( .A1(n14078), .A2(n14077), .ZN(n14199) );
  NOR2_X1 U14190 ( .A1(n8580), .A2(n8561), .ZN(n14079) );
  NOR2_X1 U14191 ( .A1(n14077), .A2(n14078), .ZN(n14196) );
  NOR2_X1 U14192 ( .A1(n14200), .A2(n14201), .ZN(n14078) );
  INV_X1 U14193 ( .A(n14202), .ZN(n14201) );
  NAND2_X1 U14194 ( .A1(n14075), .A2(n14203), .ZN(n14202) );
  NAND2_X1 U14195 ( .A1(n14204), .A2(n14072), .ZN(n14203) );
  NOR2_X1 U14196 ( .A1(n9076), .A2(n8561), .ZN(n14075) );
  NOR2_X1 U14197 ( .A1(n14072), .A2(n14204), .ZN(n14200) );
  INV_X1 U14198 ( .A(n14074), .ZN(n14204) );
  NAND2_X1 U14199 ( .A1(n14205), .A2(n14206), .ZN(n14074) );
  NAND2_X1 U14200 ( .A1(n14071), .A2(n14207), .ZN(n14206) );
  INV_X1 U14201 ( .A(n14208), .ZN(n14207) );
  NOR2_X1 U14202 ( .A1(n14070), .A2(n14069), .ZN(n14208) );
  NOR2_X1 U14203 ( .A1(n8551), .A2(n8561), .ZN(n14071) );
  NAND2_X1 U14204 ( .A1(n14069), .A2(n14070), .ZN(n14205) );
  NAND2_X1 U14205 ( .A1(n14209), .A2(n14210), .ZN(n14070) );
  NAND2_X1 U14206 ( .A1(n14067), .A2(n14211), .ZN(n14210) );
  NAND2_X1 U14207 ( .A1(n14066), .A2(n14064), .ZN(n14211) );
  NOR2_X1 U14208 ( .A1(n9094), .A2(n8561), .ZN(n14067) );
  INV_X1 U14209 ( .A(n14212), .ZN(n14209) );
  NOR2_X1 U14210 ( .A1(n14064), .A2(n14066), .ZN(n14212) );
  NOR2_X1 U14211 ( .A1(n14213), .A2(n14214), .ZN(n14066) );
  INV_X1 U14212 ( .A(n14215), .ZN(n14214) );
  NAND2_X1 U14213 ( .A1(n14063), .A2(n14216), .ZN(n14215) );
  NAND2_X1 U14214 ( .A1(n14062), .A2(n14061), .ZN(n14216) );
  NOR2_X1 U14215 ( .A1(n8548), .A2(n8561), .ZN(n14063) );
  NOR2_X1 U14216 ( .A1(n14061), .A2(n14062), .ZN(n14213) );
  INV_X1 U14217 ( .A(n14217), .ZN(n14062) );
  NAND2_X1 U14218 ( .A1(n14218), .A2(n14219), .ZN(n14217) );
  NAND2_X1 U14219 ( .A1(n14058), .A2(n14220), .ZN(n14219) );
  NAND2_X1 U14220 ( .A1(n14059), .A2(n14057), .ZN(n14220) );
  NOR2_X1 U14221 ( .A1(n8584), .A2(n8561), .ZN(n14058) );
  NAND2_X1 U14222 ( .A1(n14221), .A2(n14222), .ZN(n14218) );
  INV_X1 U14223 ( .A(n14059), .ZN(n14222) );
  NOR2_X1 U14224 ( .A1(n14223), .A2(n14224), .ZN(n14059) );
  INV_X1 U14225 ( .A(n14225), .ZN(n14224) );
  NAND2_X1 U14226 ( .A1(n14055), .A2(n14226), .ZN(n14225) );
  NAND2_X1 U14227 ( .A1(n14054), .A2(n14053), .ZN(n14226) );
  NOR2_X1 U14228 ( .A1(n8535), .A2(n8561), .ZN(n14055) );
  NOR2_X1 U14229 ( .A1(n14053), .A2(n14054), .ZN(n14223) );
  NOR2_X1 U14230 ( .A1(n14227), .A2(n14228), .ZN(n14054) );
  INV_X1 U14231 ( .A(n14229), .ZN(n14228) );
  NAND2_X1 U14232 ( .A1(n14050), .A2(n14230), .ZN(n14229) );
  NAND2_X1 U14233 ( .A1(n14051), .A2(n14049), .ZN(n14230) );
  NOR2_X1 U14234 ( .A1(n9126), .A2(n8561), .ZN(n14050) );
  NOR2_X1 U14235 ( .A1(n14049), .A2(n14051), .ZN(n14227) );
  NOR2_X1 U14236 ( .A1(n14231), .A2(n14232), .ZN(n14051) );
  INV_X1 U14237 ( .A(n14233), .ZN(n14232) );
  NAND2_X1 U14238 ( .A1(n14046), .A2(n14234), .ZN(n14233) );
  NAND2_X1 U14239 ( .A1(n14047), .A2(n14045), .ZN(n14234) );
  NOR2_X1 U14240 ( .A1(n9378), .A2(n8561), .ZN(n14046) );
  NOR2_X1 U14241 ( .A1(n14045), .A2(n14047), .ZN(n14231) );
  NOR2_X1 U14242 ( .A1(n14235), .A2(n14236), .ZN(n14047) );
  INV_X1 U14243 ( .A(n14237), .ZN(n14236) );
  NAND2_X1 U14244 ( .A1(n14042), .A2(n14238), .ZN(n14237) );
  NAND2_X1 U14245 ( .A1(n14043), .A2(n14041), .ZN(n14238) );
  NOR2_X1 U14246 ( .A1(n9383), .A2(n8561), .ZN(n14042) );
  NOR2_X1 U14247 ( .A1(n14041), .A2(n14043), .ZN(n14235) );
  NOR2_X1 U14248 ( .A1(n14239), .A2(n14240), .ZN(n14043) );
  INV_X1 U14249 ( .A(n14241), .ZN(n14240) );
  NAND2_X1 U14250 ( .A1(n14036), .A2(n14242), .ZN(n14241) );
  NAND2_X1 U14251 ( .A1(n14039), .A2(n14038), .ZN(n14242) );
  NOR2_X1 U14252 ( .A1(n9146), .A2(n8561), .ZN(n14036) );
  NOR2_X1 U14253 ( .A1(n14038), .A2(n14039), .ZN(n14239) );
  INV_X1 U14254 ( .A(n14243), .ZN(n14039) );
  NAND2_X1 U14255 ( .A1(n14244), .A2(n14245), .ZN(n14243) );
  NAND2_X1 U14256 ( .A1(n14031), .A2(n14246), .ZN(n14245) );
  NAND2_X1 U14257 ( .A1(n8624), .A2(n14247), .ZN(n14246) );
  NAND2_X1 U14258 ( .A1(n8585), .A2(n8525), .ZN(n14247) );
  NAND2_X1 U14259 ( .A1(n14248), .A2(n14249), .ZN(n14244) );
  NAND2_X1 U14260 ( .A1(n8630), .A2(n14250), .ZN(n14249) );
  NAND2_X1 U14261 ( .A1(n8539), .A2(n8526), .ZN(n14250) );
  NAND3_X1 U14262 ( .A1(n13739), .A2(n14031), .A3(n8537), .ZN(n14038) );
  INV_X1 U14263 ( .A(n13738), .ZN(n13739) );
  XNOR2_X1 U14264 ( .A(n14251), .B(n14252), .ZN(n13738) );
  XOR2_X1 U14265 ( .A(d_11_), .B(c_11_), .Z(n14252) );
  XOR2_X1 U14266 ( .A(n14253), .B(n14254), .Z(n14041) );
  XNOR2_X1 U14267 ( .A(n14255), .B(n14256), .ZN(n14254) );
  XOR2_X1 U14268 ( .A(n14257), .B(n14258), .Z(n14045) );
  XNOR2_X1 U14269 ( .A(n14259), .B(n14260), .ZN(n14257) );
  XOR2_X1 U14270 ( .A(n14261), .B(n14262), .Z(n14049) );
  XNOR2_X1 U14271 ( .A(n14263), .B(n14264), .ZN(n14261) );
  XOR2_X1 U14272 ( .A(n14265), .B(n14266), .Z(n14053) );
  XNOR2_X1 U14273 ( .A(n14267), .B(n14268), .ZN(n14265) );
  INV_X1 U14274 ( .A(n14057), .ZN(n14221) );
  XOR2_X1 U14275 ( .A(n14269), .B(n14270), .Z(n14057) );
  XOR2_X1 U14276 ( .A(n14271), .B(n14272), .Z(n14269) );
  NAND2_X1 U14277 ( .A1(n14031), .A2(n9121), .ZN(n14271) );
  XOR2_X1 U14278 ( .A(n14273), .B(n14274), .Z(n14061) );
  XNOR2_X1 U14279 ( .A(n14275), .B(n14276), .ZN(n14273) );
  NOR2_X1 U14280 ( .A1(n9176), .A2(n8526), .ZN(n14276) );
  XOR2_X1 U14281 ( .A(n14277), .B(n14278), .Z(n14064) );
  XNOR2_X1 U14282 ( .A(n14279), .B(n14280), .ZN(n14277) );
  NOR2_X1 U14283 ( .A1(n8548), .A2(n8526), .ZN(n14280) );
  XNOR2_X1 U14284 ( .A(n14281), .B(n14282), .ZN(n14069) );
  XNOR2_X1 U14285 ( .A(n14283), .B(n14284), .ZN(n14281) );
  NOR2_X1 U14286 ( .A1(n9094), .A2(n8526), .ZN(n14284) );
  XOR2_X1 U14287 ( .A(n14285), .B(n14286), .Z(n14072) );
  XNOR2_X1 U14288 ( .A(n14287), .B(n14288), .ZN(n14285) );
  NOR2_X1 U14289 ( .A1(n8551), .A2(n8526), .ZN(n14288) );
  XNOR2_X1 U14290 ( .A(n14289), .B(n14290), .ZN(n14077) );
  XNOR2_X1 U14291 ( .A(n14291), .B(n14292), .ZN(n14290) );
  NAND2_X1 U14292 ( .A1(n14031), .A2(n9080), .ZN(n14292) );
  XNOR2_X1 U14293 ( .A(n14293), .B(n14294), .ZN(n14084) );
  XNOR2_X1 U14294 ( .A(n14295), .B(n14296), .ZN(n14293) );
  XNOR2_X1 U14295 ( .A(n14297), .B(n14298), .ZN(n14088) );
  XNOR2_X1 U14296 ( .A(n14299), .B(n14300), .ZN(n14297) );
  XNOR2_X1 U14297 ( .A(n14301), .B(n14302), .ZN(n14093) );
  XNOR2_X1 U14298 ( .A(n14303), .B(n14304), .ZN(n14301) );
  XNOR2_X1 U14299 ( .A(n14305), .B(n14306), .ZN(n14096) );
  XNOR2_X1 U14300 ( .A(n14307), .B(n14308), .ZN(n14305) );
  NOR2_X1 U14301 ( .A1(n8526), .A2(n8545), .ZN(n14308) );
  XNOR2_X1 U14302 ( .A(n14309), .B(n14310), .ZN(n14100) );
  NAND2_X1 U14303 ( .A1(n14311), .A2(n14312), .ZN(n14309) );
  XNOR2_X1 U14304 ( .A(n14313), .B(n14314), .ZN(n13950) );
  XOR2_X1 U14305 ( .A(n14315), .B(n14316), .Z(n14313) );
  XNOR2_X1 U14306 ( .A(n14317), .B(n14318), .ZN(n13941) );
  XNOR2_X1 U14307 ( .A(n14319), .B(n14320), .ZN(n14318) );
  NAND2_X1 U14308 ( .A1(n9313), .A2(n14031), .ZN(n14320) );
  XNOR2_X1 U14309 ( .A(n14321), .B(n14322), .ZN(n13934) );
  NAND2_X1 U14310 ( .A1(n14323), .A2(n14324), .ZN(n14321) );
  XOR2_X1 U14311 ( .A(n14325), .B(n14326), .Z(n13926) );
  XOR2_X1 U14312 ( .A(n14327), .B(n14328), .Z(n14325) );
  XOR2_X1 U14313 ( .A(n14329), .B(n14330), .Z(n13917) );
  NAND2_X1 U14314 ( .A1(n14331), .A2(n14332), .ZN(n14329) );
  XOR2_X1 U14315 ( .A(n14333), .B(n14334), .Z(n13910) );
  XNOR2_X1 U14316 ( .A(n14335), .B(n14336), .ZN(n14334) );
  XNOR2_X1 U14317 ( .A(n14337), .B(n14338), .ZN(n13901) );
  NAND2_X1 U14318 ( .A1(n14339), .A2(n14340), .ZN(n14337) );
  XNOR2_X1 U14319 ( .A(n14341), .B(n14342), .ZN(n13894) );
  XOR2_X1 U14320 ( .A(n14343), .B(n14344), .Z(n14342) );
  XNOR2_X1 U14321 ( .A(n14345), .B(n14346), .ZN(n13885) );
  XNOR2_X1 U14322 ( .A(n14347), .B(n14348), .ZN(n14346) );
  XOR2_X1 U14323 ( .A(n14349), .B(n14350), .Z(n14105) );
  XOR2_X1 U14324 ( .A(n14351), .B(n14352), .Z(n14349) );
  XNOR2_X1 U14325 ( .A(n14353), .B(n14354), .ZN(n13873) );
  XNOR2_X1 U14326 ( .A(n14355), .B(n14356), .ZN(n14354) );
  XOR2_X1 U14327 ( .A(n14357), .B(n14358), .Z(n14109) );
  XOR2_X1 U14328 ( .A(n14359), .B(n14360), .Z(n14357) );
  XOR2_X1 U14329 ( .A(n14361), .B(n14362), .Z(n14112) );
  XNOR2_X1 U14330 ( .A(n14363), .B(n14364), .ZN(n14362) );
  XNOR2_X1 U14331 ( .A(n14365), .B(n14366), .ZN(n13863) );
  XOR2_X1 U14332 ( .A(n14367), .B(n14368), .Z(n14366) );
  XNOR2_X1 U14333 ( .A(n8604), .B(n8605), .ZN(n8868) );
  NOR3_X1 U14334 ( .A1(n8605), .A2(n8604), .A3(n8603), .ZN(n8599) );
  NAND2_X1 U14335 ( .A1(n14369), .A2(n8897), .ZN(n8603) );
  INV_X1 U14336 ( .A(n14370), .ZN(n8897) );
  NOR2_X1 U14337 ( .A1(n14371), .A2(n14372), .ZN(n14370) );
  NAND2_X1 U14338 ( .A1(n14371), .A2(n14372), .ZN(n14369) );
  NOR2_X1 U14339 ( .A1(n14373), .A2(n14374), .ZN(n14372) );
  INV_X1 U14340 ( .A(n14375), .ZN(n14374) );
  NAND3_X1 U14341 ( .A1(n8592), .A2(n14376), .A3(n14248), .ZN(n14375) );
  NAND2_X1 U14342 ( .A1(n14377), .A2(n14378), .ZN(n14376) );
  NOR2_X1 U14343 ( .A1(n14377), .A2(n14378), .ZN(n14373) );
  XNOR2_X1 U14344 ( .A(n14379), .B(n14380), .ZN(n14371) );
  XOR2_X1 U14345 ( .A(n14381), .B(n14382), .Z(n14379) );
  NOR2_X1 U14346 ( .A1(n14383), .A2(n14384), .ZN(n8604) );
  INV_X1 U14347 ( .A(n14385), .ZN(n14384) );
  NAND2_X1 U14348 ( .A1(n14368), .A2(n14386), .ZN(n14385) );
  NAND2_X1 U14349 ( .A1(n14367), .A2(n14365), .ZN(n14386) );
  NOR2_X1 U14350 ( .A1(n8526), .A2(n8972), .ZN(n14368) );
  NOR2_X1 U14351 ( .A1(n14365), .A2(n14367), .ZN(n14383) );
  INV_X1 U14352 ( .A(n14387), .ZN(n14367) );
  NAND2_X1 U14353 ( .A1(n14388), .A2(n14389), .ZN(n14387) );
  NAND2_X1 U14354 ( .A1(n14364), .A2(n14390), .ZN(n14389) );
  INV_X1 U14355 ( .A(n14391), .ZN(n14390) );
  NOR2_X1 U14356 ( .A1(n14363), .A2(n14361), .ZN(n14391) );
  NOR2_X1 U14357 ( .A1(n8589), .A2(n8526), .ZN(n14364) );
  NAND2_X1 U14358 ( .A1(n14361), .A2(n14363), .ZN(n14388) );
  NAND2_X1 U14359 ( .A1(n14392), .A2(n14393), .ZN(n14363) );
  NAND2_X1 U14360 ( .A1(n14360), .A2(n14394), .ZN(n14393) );
  INV_X1 U14361 ( .A(n14395), .ZN(n14394) );
  NOR2_X1 U14362 ( .A1(n14359), .A2(n14358), .ZN(n14395) );
  NOR2_X1 U14363 ( .A1(n8552), .A2(n8526), .ZN(n14360) );
  NAND2_X1 U14364 ( .A1(n14358), .A2(n14359), .ZN(n14392) );
  NAND2_X1 U14365 ( .A1(n14396), .A2(n14397), .ZN(n14359) );
  NAND2_X1 U14366 ( .A1(n14356), .A2(n14398), .ZN(n14397) );
  INV_X1 U14367 ( .A(n14399), .ZN(n14398) );
  NOR2_X1 U14368 ( .A1(n14355), .A2(n14353), .ZN(n14399) );
  NOR2_X1 U14369 ( .A1(n8527), .A2(n8526), .ZN(n14356) );
  NAND2_X1 U14370 ( .A1(n14353), .A2(n14355), .ZN(n14396) );
  NAND2_X1 U14371 ( .A1(n14400), .A2(n14401), .ZN(n14355) );
  NAND2_X1 U14372 ( .A1(n14352), .A2(n14402), .ZN(n14401) );
  INV_X1 U14373 ( .A(n14403), .ZN(n14402) );
  NOR2_X1 U14374 ( .A1(n14351), .A2(n14350), .ZN(n14403) );
  NOR2_X1 U14375 ( .A1(n8528), .A2(n8526), .ZN(n14352) );
  NAND2_X1 U14376 ( .A1(n14350), .A2(n14351), .ZN(n14400) );
  NAND2_X1 U14377 ( .A1(n14404), .A2(n14405), .ZN(n14351) );
  NAND2_X1 U14378 ( .A1(n14348), .A2(n14406), .ZN(n14405) );
  NAND2_X1 U14379 ( .A1(n14407), .A2(n14408), .ZN(n14406) );
  INV_X1 U14380 ( .A(n14347), .ZN(n14408) );
  INV_X1 U14381 ( .A(n14345), .ZN(n14407) );
  NOR2_X1 U14382 ( .A1(n8995), .A2(n8526), .ZN(n14348) );
  NAND2_X1 U14383 ( .A1(n14345), .A2(n14347), .ZN(n14404) );
  NAND2_X1 U14384 ( .A1(n14409), .A2(n14410), .ZN(n14347) );
  INV_X1 U14385 ( .A(n14411), .ZN(n14410) );
  NOR2_X1 U14386 ( .A1(n14344), .A2(n14412), .ZN(n14411) );
  NOR2_X1 U14387 ( .A1(n14343), .A2(n14341), .ZN(n14412) );
  NAND2_X1 U14388 ( .A1(n9286), .A2(n14031), .ZN(n14344) );
  NAND2_X1 U14389 ( .A1(n14341), .A2(n14343), .ZN(n14409) );
  NAND2_X1 U14390 ( .A1(n14339), .A2(n14413), .ZN(n14343) );
  NAND2_X1 U14391 ( .A1(n14338), .A2(n14340), .ZN(n14413) );
  NAND2_X1 U14392 ( .A1(n14414), .A2(n14415), .ZN(n14340) );
  NAND2_X1 U14393 ( .A1(n8543), .A2(n14031), .ZN(n14414) );
  XNOR2_X1 U14394 ( .A(n14416), .B(n14417), .ZN(n14338) );
  XOR2_X1 U14395 ( .A(n14418), .B(n14419), .Z(n14417) );
  NAND2_X1 U14396 ( .A1(n9295), .A2(n14248), .ZN(n14419) );
  INV_X1 U14397 ( .A(n14420), .ZN(n14339) );
  NOR2_X1 U14398 ( .A1(n14415), .A2(n8544), .ZN(n14420) );
  NAND2_X1 U14399 ( .A1(n14421), .A2(n14422), .ZN(n14415) );
  NAND2_X1 U14400 ( .A1(n14333), .A2(n14423), .ZN(n14422) );
  NAND2_X1 U14401 ( .A1(n14336), .A2(n14335), .ZN(n14423) );
  XNOR2_X1 U14402 ( .A(n14424), .B(n14425), .ZN(n14333) );
  XOR2_X1 U14403 ( .A(n14426), .B(n14427), .Z(n14424) );
  NOR2_X1 U14404 ( .A1(n8525), .A2(n8594), .ZN(n14427) );
  INV_X1 U14405 ( .A(n14428), .ZN(n14421) );
  NOR2_X1 U14406 ( .A1(n14335), .A2(n14336), .ZN(n14428) );
  NOR2_X1 U14407 ( .A1(n9010), .A2(n8526), .ZN(n14336) );
  NAND2_X1 U14408 ( .A1(n14331), .A2(n14429), .ZN(n14335) );
  NAND2_X1 U14409 ( .A1(n14330), .A2(n14332), .ZN(n14429) );
  NAND2_X1 U14410 ( .A1(n14430), .A2(n14431), .ZN(n14332) );
  NAND2_X1 U14411 ( .A1(n10846), .A2(n14031), .ZN(n14430) );
  XOR2_X1 U14412 ( .A(n14432), .B(n14433), .Z(n14330) );
  XNOR2_X1 U14413 ( .A(n14434), .B(n14435), .ZN(n14433) );
  NAND2_X1 U14414 ( .A1(n9304), .A2(n14248), .ZN(n14435) );
  INV_X1 U14415 ( .A(n14436), .ZN(n14331) );
  NOR2_X1 U14416 ( .A1(n14431), .A2(n8594), .ZN(n14436) );
  NAND2_X1 U14417 ( .A1(n14437), .A2(n14438), .ZN(n14431) );
  NAND2_X1 U14418 ( .A1(n14326), .A2(n14439), .ZN(n14438) );
  NAND2_X1 U14419 ( .A1(n14328), .A2(n14327), .ZN(n14439) );
  XOR2_X1 U14420 ( .A(n14440), .B(n14441), .Z(n14326) );
  XNOR2_X1 U14421 ( .A(n14442), .B(n14443), .ZN(n14440) );
  NOR2_X1 U14422 ( .A1(n8525), .A2(n8572), .ZN(n14443) );
  INV_X1 U14423 ( .A(n14444), .ZN(n14437) );
  NOR2_X1 U14424 ( .A1(n14327), .A2(n14328), .ZN(n14444) );
  NOR2_X1 U14425 ( .A1(n9020), .A2(n8526), .ZN(n14328) );
  NAND2_X1 U14426 ( .A1(n14323), .A2(n14445), .ZN(n14327) );
  NAND2_X1 U14427 ( .A1(n14322), .A2(n14324), .ZN(n14445) );
  NAND2_X1 U14428 ( .A1(n14446), .A2(n14447), .ZN(n14324) );
  NAND2_X1 U14429 ( .A1(n9209), .A2(n14031), .ZN(n14447) );
  INV_X1 U14430 ( .A(n14448), .ZN(n14446) );
  XOR2_X1 U14431 ( .A(n14449), .B(n14450), .Z(n14322) );
  XNOR2_X1 U14432 ( .A(n14451), .B(n14452), .ZN(n14450) );
  NAND2_X1 U14433 ( .A1(n9313), .A2(n14248), .ZN(n14452) );
  NAND2_X1 U14434 ( .A1(n9209), .A2(n14448), .ZN(n14323) );
  NAND2_X1 U14435 ( .A1(n14453), .A2(n14454), .ZN(n14448) );
  NAND3_X1 U14436 ( .A1(n14031), .A2(n14455), .A3(n9313), .ZN(n14454) );
  NAND2_X1 U14437 ( .A1(n14456), .A2(n14457), .ZN(n14455) );
  INV_X1 U14438 ( .A(n14319), .ZN(n14457) );
  INV_X1 U14439 ( .A(n14317), .ZN(n14456) );
  NAND2_X1 U14440 ( .A1(n14319), .A2(n14317), .ZN(n14453) );
  XNOR2_X1 U14441 ( .A(n14458), .B(n14459), .ZN(n14317) );
  XNOR2_X1 U14442 ( .A(n14460), .B(n14461), .ZN(n14458) );
  NOR2_X1 U14443 ( .A1(n8525), .A2(n8591), .ZN(n14461) );
  NOR2_X1 U14444 ( .A1(n14462), .A2(n14463), .ZN(n14319) );
  INV_X1 U14445 ( .A(n14464), .ZN(n14463) );
  NAND2_X1 U14446 ( .A1(n14314), .A2(n14465), .ZN(n14464) );
  NAND2_X1 U14447 ( .A1(n14316), .A2(n14315), .ZN(n14465) );
  XNOR2_X1 U14448 ( .A(n14466), .B(n14467), .ZN(n14314) );
  XNOR2_X1 U14449 ( .A(n14468), .B(n14469), .ZN(n14467) );
  NAND2_X1 U14450 ( .A1(n9322), .A2(n14248), .ZN(n14469) );
  NOR2_X1 U14451 ( .A1(n14315), .A2(n14316), .ZN(n14462) );
  NOR2_X1 U14452 ( .A1(n9036), .A2(n8526), .ZN(n14316) );
  NAND2_X1 U14453 ( .A1(n14311), .A2(n14470), .ZN(n14315) );
  NAND2_X1 U14454 ( .A1(n14310), .A2(n14312), .ZN(n14470) );
  NAND2_X1 U14455 ( .A1(n14471), .A2(n14472), .ZN(n14312) );
  NAND2_X1 U14456 ( .A1(n9322), .A2(n14031), .ZN(n14472) );
  XNOR2_X1 U14457 ( .A(n14473), .B(n14474), .ZN(n14310) );
  XOR2_X1 U14458 ( .A(n14475), .B(n14476), .Z(n14474) );
  NAND2_X1 U14459 ( .A1(n10222), .A2(n14248), .ZN(n14476) );
  NAND2_X1 U14460 ( .A1(n9322), .A2(n14477), .ZN(n14311) );
  INV_X1 U14461 ( .A(n14471), .ZN(n14477) );
  NOR2_X1 U14462 ( .A1(n14478), .A2(n14479), .ZN(n14471) );
  NOR3_X1 U14463 ( .A1(n8526), .A2(n14480), .A3(n8545), .ZN(n14479) );
  INV_X1 U14464 ( .A(n14481), .ZN(n14480) );
  NAND2_X1 U14465 ( .A1(n14307), .A2(n14306), .ZN(n14481) );
  NOR2_X1 U14466 ( .A1(n14306), .A2(n14307), .ZN(n14478) );
  NOR2_X1 U14467 ( .A1(n14482), .A2(n14483), .ZN(n14307) );
  INV_X1 U14468 ( .A(n14484), .ZN(n14483) );
  NAND2_X1 U14469 ( .A1(n14304), .A2(n14485), .ZN(n14484) );
  NAND2_X1 U14470 ( .A1(n14303), .A2(n14302), .ZN(n14485) );
  NOR2_X1 U14471 ( .A1(n9050), .A2(n8526), .ZN(n14304) );
  NOR2_X1 U14472 ( .A1(n14302), .A2(n14303), .ZN(n14482) );
  NOR2_X1 U14473 ( .A1(n14486), .A2(n14487), .ZN(n14303) );
  INV_X1 U14474 ( .A(n14488), .ZN(n14487) );
  NAND2_X1 U14475 ( .A1(n14300), .A2(n14489), .ZN(n14488) );
  NAND2_X1 U14476 ( .A1(n14298), .A2(n14299), .ZN(n14489) );
  NOR2_X1 U14477 ( .A1(n8593), .A2(n8526), .ZN(n14300) );
  NOR2_X1 U14478 ( .A1(n14298), .A2(n14299), .ZN(n14486) );
  NOR2_X1 U14479 ( .A1(n14490), .A2(n14491), .ZN(n14299) );
  INV_X1 U14480 ( .A(n14492), .ZN(n14491) );
  NAND2_X1 U14481 ( .A1(n14296), .A2(n14493), .ZN(n14492) );
  NAND2_X1 U14482 ( .A1(n14295), .A2(n14294), .ZN(n14493) );
  NOR2_X1 U14483 ( .A1(n9061), .A2(n8526), .ZN(n14296) );
  NOR2_X1 U14484 ( .A1(n14294), .A2(n14295), .ZN(n14490) );
  NOR2_X1 U14485 ( .A1(n14494), .A2(n14495), .ZN(n14295) );
  NOR2_X1 U14486 ( .A1(n14194), .A2(n14496), .ZN(n14495) );
  NOR2_X1 U14487 ( .A1(n14191), .A2(n14193), .ZN(n14496) );
  NAND2_X1 U14488 ( .A1(n14031), .A2(n9070), .ZN(n14194) );
  INV_X1 U14489 ( .A(n14497), .ZN(n14494) );
  NAND2_X1 U14490 ( .A1(n14191), .A2(n14193), .ZN(n14497) );
  NAND2_X1 U14491 ( .A1(n14498), .A2(n14499), .ZN(n14193) );
  NAND3_X1 U14492 ( .A1(n9080), .A2(n14500), .A3(n14031), .ZN(n14499) );
  NAND2_X1 U14493 ( .A1(n14289), .A2(n14291), .ZN(n14500) );
  INV_X1 U14494 ( .A(n14501), .ZN(n14498) );
  NOR2_X1 U14495 ( .A1(n14289), .A2(n14291), .ZN(n14501) );
  NOR2_X1 U14496 ( .A1(n14502), .A2(n14503), .ZN(n14291) );
  INV_X1 U14497 ( .A(n14504), .ZN(n14503) );
  NAND3_X1 U14498 ( .A1(n8515), .A2(n14505), .A3(n14031), .ZN(n14504) );
  NAND2_X1 U14499 ( .A1(n14286), .A2(n14287), .ZN(n14505) );
  NOR2_X1 U14500 ( .A1(n14286), .A2(n14287), .ZN(n14502) );
  NOR2_X1 U14501 ( .A1(n14506), .A2(n14507), .ZN(n14287) );
  INV_X1 U14502 ( .A(n14508), .ZN(n14507) );
  NAND3_X1 U14503 ( .A1(n9098), .A2(n14509), .A3(n14031), .ZN(n14508) );
  NAND2_X1 U14504 ( .A1(n14283), .A2(n14282), .ZN(n14509) );
  NOR2_X1 U14505 ( .A1(n14282), .A2(n14283), .ZN(n14506) );
  NOR2_X1 U14506 ( .A1(n14510), .A2(n14511), .ZN(n14283) );
  NOR3_X1 U14507 ( .A1(n8548), .A2(n14512), .A3(n8526), .ZN(n14511) );
  INV_X1 U14508 ( .A(n14513), .ZN(n14512) );
  NAND2_X1 U14509 ( .A1(n14278), .A2(n14279), .ZN(n14513) );
  NOR2_X1 U14510 ( .A1(n14278), .A2(n14279), .ZN(n14510) );
  NOR2_X1 U14511 ( .A1(n14514), .A2(n14515), .ZN(n14279) );
  INV_X1 U14512 ( .A(n14516), .ZN(n14515) );
  NAND3_X1 U14513 ( .A1(n9112), .A2(n14517), .A3(n14031), .ZN(n14516) );
  NAND2_X1 U14514 ( .A1(n14275), .A2(n14274), .ZN(n14517) );
  NOR2_X1 U14515 ( .A1(n14274), .A2(n14275), .ZN(n14514) );
  NOR2_X1 U14516 ( .A1(n14518), .A2(n14519), .ZN(n14275) );
  INV_X1 U14517 ( .A(n14520), .ZN(n14519) );
  NAND3_X1 U14518 ( .A1(n9121), .A2(n14521), .A3(n14031), .ZN(n14520) );
  NAND2_X1 U14519 ( .A1(n14270), .A2(n14272), .ZN(n14521) );
  NOR2_X1 U14520 ( .A1(n14270), .A2(n14272), .ZN(n14518) );
  NOR2_X1 U14521 ( .A1(n14522), .A2(n14523), .ZN(n14272) );
  INV_X1 U14522 ( .A(n14524), .ZN(n14523) );
  NAND2_X1 U14523 ( .A1(n14268), .A2(n14525), .ZN(n14524) );
  NAND2_X1 U14524 ( .A1(n14267), .A2(n14266), .ZN(n14525) );
  NOR2_X1 U14525 ( .A1(n8526), .A2(n8568), .ZN(n14268) );
  NOR2_X1 U14526 ( .A1(n14266), .A2(n14267), .ZN(n14522) );
  NOR2_X1 U14527 ( .A1(n14526), .A2(n14527), .ZN(n14267) );
  INV_X1 U14528 ( .A(n14528), .ZN(n14527) );
  NAND2_X1 U14529 ( .A1(n14263), .A2(n14529), .ZN(n14528) );
  NAND2_X1 U14530 ( .A1(n14262), .A2(n14264), .ZN(n14529) );
  NOR2_X1 U14531 ( .A1(n8526), .A2(n8574), .ZN(n14263) );
  NOR2_X1 U14532 ( .A1(n14262), .A2(n14264), .ZN(n14526) );
  NOR2_X1 U14533 ( .A1(n14530), .A2(n14531), .ZN(n14264) );
  INV_X1 U14534 ( .A(n14532), .ZN(n14531) );
  NAND2_X1 U14535 ( .A1(n14259), .A2(n14533), .ZN(n14532) );
  NAND2_X1 U14536 ( .A1(n14260), .A2(n14258), .ZN(n14533) );
  NOR2_X1 U14537 ( .A1(n8526), .A2(n8565), .ZN(n14259) );
  NOR2_X1 U14538 ( .A1(n14258), .A2(n14260), .ZN(n14530) );
  NOR2_X1 U14539 ( .A1(n14534), .A2(n14535), .ZN(n14260) );
  INV_X1 U14540 ( .A(n14536), .ZN(n14535) );
  NAND2_X1 U14541 ( .A1(n14253), .A2(n14537), .ZN(n14536) );
  NAND2_X1 U14542 ( .A1(n14256), .A2(n14255), .ZN(n14537) );
  NOR2_X1 U14543 ( .A1(n8526), .A2(n8567), .ZN(n14253) );
  NOR2_X1 U14544 ( .A1(n14255), .A2(n14256), .ZN(n14534) );
  INV_X1 U14545 ( .A(n14538), .ZN(n14256) );
  NAND2_X1 U14546 ( .A1(n14539), .A2(n14540), .ZN(n14538) );
  NAND2_X1 U14547 ( .A1(n14248), .A2(n14541), .ZN(n14540) );
  NAND2_X1 U14548 ( .A1(n8624), .A2(n14542), .ZN(n14541) );
  NAND2_X1 U14549 ( .A1(n8530), .A2(n8585), .ZN(n14542) );
  NAND2_X1 U14550 ( .A1(n14543), .A2(n14544), .ZN(n14539) );
  NAND2_X1 U14551 ( .A1(n8630), .A2(n14545), .ZN(n14544) );
  NAND2_X1 U14552 ( .A1(n8539), .A2(n8525), .ZN(n14545) );
  NAND3_X1 U14553 ( .A1(n14031), .A2(n8537), .A3(n14248), .ZN(n14255) );
  INV_X1 U14554 ( .A(n8526), .ZN(n14031) );
  XOR2_X1 U14555 ( .A(d_10_), .B(c_10_), .Z(n14547) );
  XOR2_X1 U14556 ( .A(n14548), .B(n14549), .Z(n14258) );
  XNOR2_X1 U14557 ( .A(n14550), .B(n14551), .ZN(n14549) );
  XOR2_X1 U14558 ( .A(n14552), .B(n14553), .Z(n14262) );
  XNOR2_X1 U14559 ( .A(n14554), .B(n14555), .ZN(n14552) );
  XOR2_X1 U14560 ( .A(n14556), .B(n14557), .Z(n14266) );
  XNOR2_X1 U14561 ( .A(n14558), .B(n14559), .ZN(n14556) );
  XOR2_X1 U14562 ( .A(n14560), .B(n14561), .Z(n14270) );
  XNOR2_X1 U14563 ( .A(n14562), .B(n14563), .ZN(n14560) );
  XOR2_X1 U14564 ( .A(n14564), .B(n14565), .Z(n14274) );
  XNOR2_X1 U14565 ( .A(n14566), .B(n14567), .ZN(n14564) );
  XOR2_X1 U14566 ( .A(n14568), .B(n14569), .Z(n14278) );
  XNOR2_X1 U14567 ( .A(n14570), .B(n14571), .ZN(n14568) );
  XOR2_X1 U14568 ( .A(n14572), .B(n14573), .Z(n14282) );
  XNOR2_X1 U14569 ( .A(n14574), .B(n14575), .ZN(n14572) );
  XNOR2_X1 U14570 ( .A(n14576), .B(n14577), .ZN(n14286) );
  XOR2_X1 U14571 ( .A(n14578), .B(n14579), .Z(n14577) );
  XOR2_X1 U14572 ( .A(n14580), .B(n14581), .Z(n14289) );
  XNOR2_X1 U14573 ( .A(n14582), .B(n14583), .ZN(n14580) );
  XNOR2_X1 U14574 ( .A(n14584), .B(n14585), .ZN(n14191) );
  NAND2_X1 U14575 ( .A1(n14586), .A2(n14587), .ZN(n14584) );
  XOR2_X1 U14576 ( .A(n14588), .B(n14589), .Z(n14294) );
  XOR2_X1 U14577 ( .A(n14590), .B(n14591), .Z(n14589) );
  NAND2_X1 U14578 ( .A1(n14248), .A2(n9070), .ZN(n14591) );
  XOR2_X1 U14579 ( .A(n14592), .B(n14593), .Z(n14298) );
  XOR2_X1 U14580 ( .A(n14594), .B(n14595), .Z(n14593) );
  NAND2_X1 U14581 ( .A1(n9340), .A2(n14248), .ZN(n14595) );
  XOR2_X1 U14582 ( .A(n14596), .B(n14597), .Z(n14302) );
  XOR2_X1 U14583 ( .A(n14598), .B(n14599), .Z(n14597) );
  NAND2_X1 U14584 ( .A1(n10722), .A2(n14248), .ZN(n14599) );
  XOR2_X1 U14585 ( .A(n14600), .B(n14601), .Z(n14306) );
  XOR2_X1 U14586 ( .A(n14602), .B(n14603), .Z(n14601) );
  NAND2_X1 U14587 ( .A1(n9331), .A2(n14248), .ZN(n14603) );
  XOR2_X1 U14588 ( .A(n14604), .B(n14605), .Z(n14341) );
  XOR2_X1 U14589 ( .A(n14606), .B(n14607), .Z(n14604) );
  NOR2_X1 U14590 ( .A1(n8525), .A2(n8544), .ZN(n14607) );
  XNOR2_X1 U14591 ( .A(n14608), .B(n14609), .ZN(n14345) );
  XOR2_X1 U14592 ( .A(n14610), .B(n14611), .Z(n14609) );
  NAND2_X1 U14593 ( .A1(n9286), .A2(n14248), .ZN(n14611) );
  XOR2_X1 U14594 ( .A(n14612), .B(n14613), .Z(n14350) );
  XOR2_X1 U14595 ( .A(n14614), .B(n14615), .Z(n14612) );
  NOR2_X1 U14596 ( .A1(n8525), .A2(n8564), .ZN(n14615) );
  XNOR2_X1 U14597 ( .A(n14616), .B(n14617), .ZN(n14353) );
  XOR2_X1 U14598 ( .A(n14618), .B(n14619), .Z(n14617) );
  NAND2_X1 U14599 ( .A1(n9277), .A2(n14248), .ZN(n14619) );
  XOR2_X1 U14600 ( .A(n14620), .B(n14621), .Z(n14358) );
  XNOR2_X1 U14601 ( .A(n14622), .B(n14623), .ZN(n14620) );
  NAND2_X1 U14602 ( .A1(n9792), .A2(n14248), .ZN(n14622) );
  XNOR2_X1 U14603 ( .A(n14624), .B(n14625), .ZN(n14361) );
  XOR2_X1 U14604 ( .A(n14626), .B(n14627), .Z(n14625) );
  NAND2_X1 U14605 ( .A1(n9268), .A2(n14248), .ZN(n14627) );
  XOR2_X1 U14606 ( .A(n14628), .B(n14629), .Z(n14365) );
  XOR2_X1 U14607 ( .A(n14630), .B(n14631), .Z(n14628) );
  NAND2_X1 U14608 ( .A1(n9263), .A2(n14248), .ZN(n14630) );
  XNOR2_X1 U14609 ( .A(n14377), .B(n14632), .ZN(n8605) );
  XNOR2_X1 U14610 ( .A(n14378), .B(n14633), .ZN(n14632) );
  NAND2_X1 U14611 ( .A1(n14248), .A2(n8872), .ZN(n14633) );
  NOR2_X1 U14612 ( .A1(n14634), .A2(n14635), .ZN(n14378) );
  INV_X1 U14613 ( .A(n14636), .ZN(n14635) );
  NAND3_X1 U14614 ( .A1(n14248), .A2(n14637), .A3(n9263), .ZN(n14636) );
  NAND2_X1 U14615 ( .A1(n14629), .A2(n14631), .ZN(n14637) );
  NOR2_X1 U14616 ( .A1(n14629), .A2(n14631), .ZN(n14634) );
  NOR2_X1 U14617 ( .A1(n14638), .A2(n14639), .ZN(n14631) );
  NOR3_X1 U14618 ( .A1(n8525), .A2(n14640), .A3(n8552), .ZN(n14639) );
  NOR2_X1 U14619 ( .A1(n14624), .A2(n14626), .ZN(n14640) );
  INV_X1 U14620 ( .A(n14641), .ZN(n14638) );
  NAND2_X1 U14621 ( .A1(n14624), .A2(n14626), .ZN(n14641) );
  NAND2_X1 U14622 ( .A1(n14642), .A2(n14643), .ZN(n14626) );
  NAND3_X1 U14623 ( .A1(n14248), .A2(n14644), .A3(n9792), .ZN(n14643) );
  INV_X1 U14624 ( .A(n14645), .ZN(n14644) );
  NOR2_X1 U14625 ( .A1(n14621), .A2(n14623), .ZN(n14645) );
  NAND2_X1 U14626 ( .A1(n14621), .A2(n14623), .ZN(n14642) );
  NAND2_X1 U14627 ( .A1(n14646), .A2(n14647), .ZN(n14623) );
  INV_X1 U14628 ( .A(n14648), .ZN(n14647) );
  NOR3_X1 U14629 ( .A1(n8525), .A2(n14649), .A3(n8528), .ZN(n14648) );
  NOR2_X1 U14630 ( .A1(n14616), .A2(n14618), .ZN(n14649) );
  NAND2_X1 U14631 ( .A1(n14616), .A2(n14618), .ZN(n14646) );
  NAND2_X1 U14632 ( .A1(n14650), .A2(n14651), .ZN(n14618) );
  NAND3_X1 U14633 ( .A1(n14248), .A2(n14652), .A3(n10307), .ZN(n14651) );
  INV_X1 U14634 ( .A(n14653), .ZN(n14652) );
  NOR2_X1 U14635 ( .A1(n14613), .A2(n14614), .ZN(n14653) );
  NAND2_X1 U14636 ( .A1(n14613), .A2(n14614), .ZN(n14650) );
  NAND2_X1 U14637 ( .A1(n14654), .A2(n14655), .ZN(n14614) );
  INV_X1 U14638 ( .A(n14656), .ZN(n14655) );
  NOR3_X1 U14639 ( .A1(n8525), .A2(n14657), .A3(n8555), .ZN(n14656) );
  NOR2_X1 U14640 ( .A1(n14610), .A2(n14608), .ZN(n14657) );
  NAND2_X1 U14641 ( .A1(n14608), .A2(n14610), .ZN(n14654) );
  NAND2_X1 U14642 ( .A1(n14658), .A2(n14659), .ZN(n14610) );
  NAND3_X1 U14643 ( .A1(n14248), .A2(n14660), .A3(n8543), .ZN(n14659) );
  INV_X1 U14644 ( .A(n14661), .ZN(n14660) );
  NOR2_X1 U14645 ( .A1(n14605), .A2(n14606), .ZN(n14661) );
  NAND2_X1 U14646 ( .A1(n14605), .A2(n14606), .ZN(n14658) );
  NAND2_X1 U14647 ( .A1(n14662), .A2(n14663), .ZN(n14606) );
  NAND3_X1 U14648 ( .A1(n14248), .A2(n14664), .A3(n9295), .ZN(n14663) );
  INV_X1 U14649 ( .A(n14665), .ZN(n14664) );
  NOR2_X1 U14650 ( .A1(n14418), .A2(n14416), .ZN(n14665) );
  NAND2_X1 U14651 ( .A1(n14416), .A2(n14418), .ZN(n14662) );
  NAND2_X1 U14652 ( .A1(n14666), .A2(n14667), .ZN(n14418) );
  NAND3_X1 U14653 ( .A1(n14248), .A2(n14668), .A3(n10846), .ZN(n14667) );
  INV_X1 U14654 ( .A(n14669), .ZN(n14668) );
  NOR2_X1 U14655 ( .A1(n14425), .A2(n14426), .ZN(n14669) );
  NAND2_X1 U14656 ( .A1(n14425), .A2(n14426), .ZN(n14666) );
  NAND2_X1 U14657 ( .A1(n14670), .A2(n14671), .ZN(n14426) );
  NAND3_X1 U14658 ( .A1(n14248), .A2(n14672), .A3(n9304), .ZN(n14671) );
  NAND2_X1 U14659 ( .A1(n14434), .A2(n14432), .ZN(n14672) );
  INV_X1 U14660 ( .A(n14673), .ZN(n14670) );
  NOR2_X1 U14661 ( .A1(n14432), .A2(n14434), .ZN(n14673) );
  NOR2_X1 U14662 ( .A1(n14674), .A2(n14675), .ZN(n14434) );
  INV_X1 U14663 ( .A(n14676), .ZN(n14675) );
  NAND3_X1 U14664 ( .A1(n14248), .A2(n14677), .A3(n9209), .ZN(n14676) );
  NAND2_X1 U14665 ( .A1(n14442), .A2(n14441), .ZN(n14677) );
  NOR2_X1 U14666 ( .A1(n14441), .A2(n14442), .ZN(n14674) );
  NOR2_X1 U14667 ( .A1(n14678), .A2(n14679), .ZN(n14442) );
  NOR3_X1 U14668 ( .A1(n8525), .A2(n14680), .A3(n8582), .ZN(n14679) );
  INV_X1 U14669 ( .A(n14681), .ZN(n14680) );
  NAND2_X1 U14670 ( .A1(n14451), .A2(n14449), .ZN(n14681) );
  NOR2_X1 U14671 ( .A1(n14449), .A2(n14451), .ZN(n14678) );
  NOR2_X1 U14672 ( .A1(n14682), .A2(n14683), .ZN(n14451) );
  INV_X1 U14673 ( .A(n14684), .ZN(n14683) );
  NAND3_X1 U14674 ( .A1(n14248), .A2(n14685), .A3(n9721), .ZN(n14684) );
  NAND2_X1 U14675 ( .A1(n14460), .A2(n14459), .ZN(n14685) );
  NOR2_X1 U14676 ( .A1(n14459), .A2(n14460), .ZN(n14682) );
  NOR2_X1 U14677 ( .A1(n14686), .A2(n14687), .ZN(n14460) );
  NOR3_X1 U14678 ( .A1(n8525), .A2(n14688), .A3(n8562), .ZN(n14687) );
  INV_X1 U14679 ( .A(n14689), .ZN(n14688) );
  NAND2_X1 U14680 ( .A1(n14466), .A2(n14468), .ZN(n14689) );
  NOR2_X1 U14681 ( .A1(n14466), .A2(n14468), .ZN(n14686) );
  NOR2_X1 U14682 ( .A1(n14690), .A2(n14691), .ZN(n14468) );
  NOR3_X1 U14683 ( .A1(n8525), .A2(n14692), .A3(n8545), .ZN(n14691) );
  NOR2_X1 U14684 ( .A1(n14475), .A2(n14473), .ZN(n14692) );
  INV_X1 U14685 ( .A(n14693), .ZN(n14690) );
  NAND2_X1 U14686 ( .A1(n14473), .A2(n14475), .ZN(n14693) );
  NAND2_X1 U14687 ( .A1(n14694), .A2(n14695), .ZN(n14475) );
  INV_X1 U14688 ( .A(n14696), .ZN(n14695) );
  NOR3_X1 U14689 ( .A1(n8525), .A2(n14697), .A3(n8569), .ZN(n14696) );
  NOR2_X1 U14690 ( .A1(n14600), .A2(n14602), .ZN(n14697) );
  NAND2_X1 U14691 ( .A1(n14600), .A2(n14602), .ZN(n14694) );
  NAND2_X1 U14692 ( .A1(n14698), .A2(n14699), .ZN(n14602) );
  NAND3_X1 U14693 ( .A1(n14248), .A2(n14700), .A3(n10722), .ZN(n14699) );
  INV_X1 U14694 ( .A(n14701), .ZN(n14700) );
  NOR2_X1 U14695 ( .A1(n14596), .A2(n14598), .ZN(n14701) );
  NAND2_X1 U14696 ( .A1(n14596), .A2(n14598), .ZN(n14698) );
  NAND2_X1 U14697 ( .A1(n14702), .A2(n14703), .ZN(n14598) );
  INV_X1 U14698 ( .A(n14704), .ZN(n14703) );
  NOR3_X1 U14699 ( .A1(n8525), .A2(n14705), .A3(n8583), .ZN(n14704) );
  NOR2_X1 U14700 ( .A1(n14594), .A2(n14592), .ZN(n14705) );
  NAND2_X1 U14701 ( .A1(n14592), .A2(n14594), .ZN(n14702) );
  NAND2_X1 U14702 ( .A1(n14706), .A2(n14707), .ZN(n14594) );
  NAND3_X1 U14703 ( .A1(n9070), .A2(n14708), .A3(n14248), .ZN(n14707) );
  INV_X1 U14704 ( .A(n14709), .ZN(n14708) );
  NOR2_X1 U14705 ( .A1(n14588), .A2(n14590), .ZN(n14709) );
  NAND2_X1 U14706 ( .A1(n14588), .A2(n14590), .ZN(n14706) );
  NAND2_X1 U14707 ( .A1(n14586), .A2(n14710), .ZN(n14590) );
  NAND2_X1 U14708 ( .A1(n14585), .A2(n14587), .ZN(n14710) );
  NAND2_X1 U14709 ( .A1(n14711), .A2(n14712), .ZN(n14587) );
  NAND2_X1 U14710 ( .A1(n14248), .A2(n9080), .ZN(n14712) );
  XNOR2_X1 U14711 ( .A(n14713), .B(n14714), .ZN(n14585) );
  XOR2_X1 U14712 ( .A(n14715), .B(n14716), .Z(n14714) );
  NAND2_X1 U14713 ( .A1(n9080), .A2(n14717), .ZN(n14586) );
  INV_X1 U14714 ( .A(n14711), .ZN(n14717) );
  NOR2_X1 U14715 ( .A1(n14718), .A2(n14719), .ZN(n14711) );
  INV_X1 U14716 ( .A(n14720), .ZN(n14719) );
  NAND2_X1 U14717 ( .A1(n14583), .A2(n14721), .ZN(n14720) );
  NAND2_X1 U14718 ( .A1(n14582), .A2(n14581), .ZN(n14721) );
  NOR2_X1 U14719 ( .A1(n8525), .A2(n8551), .ZN(n14583) );
  NOR2_X1 U14720 ( .A1(n14581), .A2(n14582), .ZN(n14718) );
  NOR2_X1 U14721 ( .A1(n14722), .A2(n14723), .ZN(n14582) );
  INV_X1 U14722 ( .A(n14724), .ZN(n14723) );
  NAND2_X1 U14723 ( .A1(n14579), .A2(n14725), .ZN(n14724) );
  NAND2_X1 U14724 ( .A1(n14578), .A2(n14576), .ZN(n14725) );
  NOR2_X1 U14725 ( .A1(n8525), .A2(n8563), .ZN(n14579) );
  NOR2_X1 U14726 ( .A1(n14576), .A2(n14578), .ZN(n14722) );
  NOR2_X1 U14727 ( .A1(n14726), .A2(n14727), .ZN(n14578) );
  INV_X1 U14728 ( .A(n14728), .ZN(n14727) );
  NAND2_X1 U14729 ( .A1(n14575), .A2(n14729), .ZN(n14728) );
  NAND2_X1 U14730 ( .A1(n14573), .A2(n14574), .ZN(n14729) );
  NOR2_X1 U14731 ( .A1(n8525), .A2(n8548), .ZN(n14575) );
  NOR2_X1 U14732 ( .A1(n14573), .A2(n14574), .ZN(n14726) );
  INV_X1 U14733 ( .A(n14730), .ZN(n14574) );
  NAND2_X1 U14734 ( .A1(n14731), .A2(n14732), .ZN(n14730) );
  NAND2_X1 U14735 ( .A1(n14571), .A2(n14733), .ZN(n14732) );
  NAND2_X1 U14736 ( .A1(n14570), .A2(n14569), .ZN(n14733) );
  NOR2_X1 U14737 ( .A1(n8525), .A2(n8584), .ZN(n14571) );
  NAND2_X1 U14738 ( .A1(n14734), .A2(n14735), .ZN(n14731) );
  INV_X1 U14739 ( .A(n14570), .ZN(n14735) );
  NOR2_X1 U14740 ( .A1(n14736), .A2(n14737), .ZN(n14570) );
  INV_X1 U14741 ( .A(n14738), .ZN(n14737) );
  NAND2_X1 U14742 ( .A1(n14567), .A2(n14739), .ZN(n14738) );
  NAND2_X1 U14743 ( .A1(n14565), .A2(n14566), .ZN(n14739) );
  NOR2_X1 U14744 ( .A1(n8525), .A2(n8535), .ZN(n14567) );
  NOR2_X1 U14745 ( .A1(n14565), .A2(n14566), .ZN(n14736) );
  NOR2_X1 U14746 ( .A1(n14740), .A2(n14741), .ZN(n14566) );
  INV_X1 U14747 ( .A(n14742), .ZN(n14741) );
  NAND2_X1 U14748 ( .A1(n14563), .A2(n14743), .ZN(n14742) );
  NAND2_X1 U14749 ( .A1(n14562), .A2(n14561), .ZN(n14743) );
  NOR2_X1 U14750 ( .A1(n8525), .A2(n9126), .ZN(n14563) );
  NOR2_X1 U14751 ( .A1(n14561), .A2(n14562), .ZN(n14740) );
  NOR2_X1 U14752 ( .A1(n14744), .A2(n14745), .ZN(n14562) );
  INV_X1 U14753 ( .A(n14746), .ZN(n14745) );
  NAND2_X1 U14754 ( .A1(n14558), .A2(n14747), .ZN(n14746) );
  NAND2_X1 U14755 ( .A1(n14557), .A2(n14559), .ZN(n14747) );
  NOR2_X1 U14756 ( .A1(n8525), .A2(n8574), .ZN(n14558) );
  NOR2_X1 U14757 ( .A1(n14557), .A2(n14559), .ZN(n14744) );
  NOR2_X1 U14758 ( .A1(n14748), .A2(n14749), .ZN(n14559) );
  INV_X1 U14759 ( .A(n14750), .ZN(n14749) );
  NAND2_X1 U14760 ( .A1(n14554), .A2(n14751), .ZN(n14750) );
  NAND2_X1 U14761 ( .A1(n14555), .A2(n14553), .ZN(n14751) );
  NOR2_X1 U14762 ( .A1(n8525), .A2(n8565), .ZN(n14554) );
  NOR2_X1 U14763 ( .A1(n14553), .A2(n14555), .ZN(n14748) );
  NOR2_X1 U14764 ( .A1(n14752), .A2(n14753), .ZN(n14555) );
  INV_X1 U14765 ( .A(n14754), .ZN(n14753) );
  NAND2_X1 U14766 ( .A1(n14548), .A2(n14755), .ZN(n14754) );
  NAND2_X1 U14767 ( .A1(n14551), .A2(n14550), .ZN(n14755) );
  NOR2_X1 U14768 ( .A1(n8525), .A2(n8567), .ZN(n14548) );
  NOR2_X1 U14769 ( .A1(n14550), .A2(n14551), .ZN(n14752) );
  INV_X1 U14770 ( .A(n14756), .ZN(n14551) );
  NAND2_X1 U14771 ( .A1(n14757), .A2(n14758), .ZN(n14756) );
  NAND2_X1 U14772 ( .A1(n14543), .A2(n14759), .ZN(n14758) );
  NAND2_X1 U14773 ( .A1(n8624), .A2(n14760), .ZN(n14759) );
  NAND2_X1 U14774 ( .A1(n8534), .A2(n8627), .ZN(n14760) );
  NAND2_X1 U14775 ( .A1(n14761), .A2(n14762), .ZN(n14757) );
  NAND2_X1 U14776 ( .A1(n8630), .A2(n14763), .ZN(n14762) );
  NAND2_X1 U14777 ( .A1(n8539), .A2(n8530), .ZN(n14763) );
  NAND3_X1 U14778 ( .A1(n14248), .A2(n8537), .A3(n14543), .ZN(n14550) );
  XOR2_X1 U14779 ( .A(d_9_), .B(c_9_), .Z(n14765) );
  XOR2_X1 U14780 ( .A(n14766), .B(n14767), .Z(n14553) );
  XNOR2_X1 U14781 ( .A(n14768), .B(n14769), .ZN(n14767) );
  XOR2_X1 U14782 ( .A(n14770), .B(n14771), .Z(n14557) );
  XNOR2_X1 U14783 ( .A(n14772), .B(n14773), .ZN(n14770) );
  XOR2_X1 U14784 ( .A(n14774), .B(n14775), .Z(n14561) );
  XNOR2_X1 U14785 ( .A(n14776), .B(n14777), .ZN(n14774) );
  XOR2_X1 U14786 ( .A(n14778), .B(n14779), .Z(n14565) );
  XNOR2_X1 U14787 ( .A(n14780), .B(n14781), .ZN(n14778) );
  INV_X1 U14788 ( .A(n14569), .ZN(n14734) );
  XOR2_X1 U14789 ( .A(n14782), .B(n14783), .Z(n14569) );
  XOR2_X1 U14790 ( .A(n14784), .B(n14785), .Z(n14782) );
  NAND2_X1 U14791 ( .A1(n14543), .A2(n9121), .ZN(n14784) );
  XOR2_X1 U14792 ( .A(n14786), .B(n14787), .Z(n14573) );
  XNOR2_X1 U14793 ( .A(n14788), .B(n14789), .ZN(n14786) );
  NOR2_X1 U14794 ( .A1(n9176), .A2(n8530), .ZN(n14789) );
  XOR2_X1 U14795 ( .A(n14790), .B(n14791), .Z(n14576) );
  XNOR2_X1 U14796 ( .A(n14792), .B(n14793), .ZN(n14790) );
  NOR2_X1 U14797 ( .A1(n8548), .A2(n8530), .ZN(n14793) );
  XNOR2_X1 U14798 ( .A(n14794), .B(n14795), .ZN(n14581) );
  XNOR2_X1 U14799 ( .A(n14796), .B(n14797), .ZN(n14795) );
  NAND2_X1 U14800 ( .A1(n14543), .A2(n9098), .ZN(n14797) );
  XNOR2_X1 U14801 ( .A(n14798), .B(n14799), .ZN(n14588) );
  XNOR2_X1 U14802 ( .A(n14800), .B(n14801), .ZN(n14798) );
  NOR2_X1 U14803 ( .A1(n9076), .A2(n8530), .ZN(n14801) );
  XNOR2_X1 U14804 ( .A(n14802), .B(n14803), .ZN(n14592) );
  NAND2_X1 U14805 ( .A1(n14804), .A2(n14805), .ZN(n14802) );
  XNOR2_X1 U14806 ( .A(n14806), .B(n14807), .ZN(n14596) );
  XOR2_X1 U14807 ( .A(n14808), .B(n14809), .Z(n14806) );
  XNOR2_X1 U14808 ( .A(n14810), .B(n14811), .ZN(n14600) );
  XNOR2_X1 U14809 ( .A(n14812), .B(n14813), .ZN(n14810) );
  NOR2_X1 U14810 ( .A1(n8530), .A2(n8593), .ZN(n14813) );
  XNOR2_X1 U14811 ( .A(n14814), .B(n14815), .ZN(n14473) );
  NAND2_X1 U14812 ( .A1(n14816), .A2(n14817), .ZN(n14814) );
  XOR2_X1 U14813 ( .A(n14818), .B(n14819), .Z(n14466) );
  NAND2_X1 U14814 ( .A1(n14820), .A2(n14821), .ZN(n14818) );
  XOR2_X1 U14815 ( .A(n14822), .B(n14823), .Z(n14459) );
  NAND2_X1 U14816 ( .A1(n14824), .A2(n14825), .ZN(n14822) );
  XOR2_X1 U14817 ( .A(n14826), .B(n14827), .Z(n14449) );
  XOR2_X1 U14818 ( .A(n14828), .B(n14829), .Z(n14826) );
  XNOR2_X1 U14819 ( .A(n14830), .B(n14831), .ZN(n14441) );
  XOR2_X1 U14820 ( .A(n14832), .B(n14833), .Z(n14831) );
  XOR2_X1 U14821 ( .A(n14834), .B(n14835), .Z(n14432) );
  XOR2_X1 U14822 ( .A(n14836), .B(n14837), .Z(n14835) );
  XNOR2_X1 U14823 ( .A(n14838), .B(n14839), .ZN(n14425) );
  XNOR2_X1 U14824 ( .A(n14840), .B(n14841), .ZN(n14838) );
  XOR2_X1 U14825 ( .A(n14842), .B(n14843), .Z(n14416) );
  XOR2_X1 U14826 ( .A(n14844), .B(n14845), .Z(n14843) );
  XOR2_X1 U14827 ( .A(n14846), .B(n14847), .Z(n14605) );
  XOR2_X1 U14828 ( .A(n14848), .B(n14849), .Z(n14846) );
  XNOR2_X1 U14829 ( .A(n14850), .B(n14851), .ZN(n14608) );
  XNOR2_X1 U14830 ( .A(n14852), .B(n14853), .ZN(n14851) );
  XOR2_X1 U14831 ( .A(n14854), .B(n14855), .Z(n14613) );
  XOR2_X1 U14832 ( .A(n14856), .B(n14857), .Z(n14854) );
  XNOR2_X1 U14833 ( .A(n14858), .B(n14859), .ZN(n14616) );
  XNOR2_X1 U14834 ( .A(n14860), .B(n14861), .ZN(n14859) );
  XOR2_X1 U14835 ( .A(n14862), .B(n14863), .Z(n14621) );
  XOR2_X1 U14836 ( .A(n14864), .B(n14865), .Z(n14862) );
  XOR2_X1 U14837 ( .A(n14866), .B(n14867), .Z(n14624) );
  XNOR2_X1 U14838 ( .A(n14868), .B(n14869), .ZN(n14867) );
  XOR2_X1 U14839 ( .A(n14870), .B(n14871), .Z(n14629) );
  XNOR2_X1 U14840 ( .A(n14872), .B(n14873), .ZN(n14870) );
  XNOR2_X1 U14841 ( .A(n14874), .B(n14875), .ZN(n14377) );
  XOR2_X1 U14842 ( .A(n14876), .B(n14877), .Z(n14875) );
  XOR2_X1 U14843 ( .A(n8615), .B(n8616), .Z(n8606) );
  NOR3_X1 U14844 ( .A1(n8616), .A2(n8615), .A3(n8614), .ZN(n8610) );
  NAND2_X1 U14845 ( .A1(n14878), .A2(n8894), .ZN(n8614) );
  INV_X1 U14846 ( .A(n14879), .ZN(n8894) );
  NOR2_X1 U14847 ( .A1(n14880), .A2(n14881), .ZN(n14879) );
  NAND2_X1 U14848 ( .A1(n14880), .A2(n14881), .ZN(n14878) );
  NOR2_X1 U14849 ( .A1(n14882), .A2(n14883), .ZN(n14881) );
  INV_X1 U14850 ( .A(n14884), .ZN(n14883) );
  NAND3_X1 U14851 ( .A1(n8592), .A2(n14885), .A3(n14761), .ZN(n14884) );
  NAND2_X1 U14852 ( .A1(n14886), .A2(n14887), .ZN(n14885) );
  NOR2_X1 U14853 ( .A1(n14886), .A2(n14887), .ZN(n14882) );
  XNOR2_X1 U14854 ( .A(n14888), .B(n14889), .ZN(n14880) );
  XOR2_X1 U14855 ( .A(n14890), .B(n14891), .Z(n14888) );
  NOR2_X1 U14856 ( .A1(n14892), .A2(n14893), .ZN(n8615) );
  INV_X1 U14857 ( .A(n14894), .ZN(n14893) );
  NAND2_X1 U14858 ( .A1(n14382), .A2(n14895), .ZN(n14894) );
  NAND2_X1 U14859 ( .A1(n14381), .A2(n14380), .ZN(n14895) );
  NOR2_X1 U14860 ( .A1(n8530), .A2(n8972), .ZN(n14382) );
  NOR2_X1 U14861 ( .A1(n14380), .A2(n14381), .ZN(n14892) );
  NOR2_X1 U14862 ( .A1(n14896), .A2(n14897), .ZN(n14381) );
  INV_X1 U14863 ( .A(n14898), .ZN(n14897) );
  NAND2_X1 U14864 ( .A1(n14877), .A2(n14899), .ZN(n14898) );
  NAND2_X1 U14865 ( .A1(n14876), .A2(n14874), .ZN(n14899) );
  NOR2_X1 U14866 ( .A1(n8589), .A2(n8530), .ZN(n14877) );
  NOR2_X1 U14867 ( .A1(n14874), .A2(n14876), .ZN(n14896) );
  NOR2_X1 U14868 ( .A1(n14900), .A2(n14901), .ZN(n14876) );
  INV_X1 U14869 ( .A(n14902), .ZN(n14901) );
  NAND2_X1 U14870 ( .A1(n14872), .A2(n14903), .ZN(n14902) );
  NAND2_X1 U14871 ( .A1(n14873), .A2(n14871), .ZN(n14903) );
  NOR2_X1 U14872 ( .A1(n8982), .A2(n8530), .ZN(n14872) );
  NOR2_X1 U14873 ( .A1(n14871), .A2(n14873), .ZN(n14900) );
  NOR2_X1 U14874 ( .A1(n14904), .A2(n14905), .ZN(n14873) );
  INV_X1 U14875 ( .A(n14906), .ZN(n14905) );
  NAND2_X1 U14876 ( .A1(n14869), .A2(n14907), .ZN(n14906) );
  NAND2_X1 U14877 ( .A1(n14908), .A2(n14866), .ZN(n14907) );
  NOR2_X1 U14878 ( .A1(n8527), .A2(n8530), .ZN(n14869) );
  NOR2_X1 U14879 ( .A1(n14866), .A2(n14908), .ZN(n14904) );
  INV_X1 U14880 ( .A(n14868), .ZN(n14908) );
  NAND2_X1 U14881 ( .A1(n14909), .A2(n14910), .ZN(n14868) );
  NAND2_X1 U14882 ( .A1(n14864), .A2(n14911), .ZN(n14910) );
  INV_X1 U14883 ( .A(n14912), .ZN(n14911) );
  NOR2_X1 U14884 ( .A1(n14865), .A2(n14863), .ZN(n14912) );
  NOR2_X1 U14885 ( .A1(n8528), .A2(n8530), .ZN(n14864) );
  NAND2_X1 U14886 ( .A1(n14863), .A2(n14865), .ZN(n14909) );
  NAND2_X1 U14887 ( .A1(n14913), .A2(n14914), .ZN(n14865) );
  NAND2_X1 U14888 ( .A1(n14861), .A2(n14915), .ZN(n14914) );
  INV_X1 U14889 ( .A(n14916), .ZN(n14915) );
  NOR2_X1 U14890 ( .A1(n14860), .A2(n14858), .ZN(n14916) );
  NOR2_X1 U14891 ( .A1(n8995), .A2(n8530), .ZN(n14861) );
  NAND2_X1 U14892 ( .A1(n14858), .A2(n14860), .ZN(n14913) );
  NAND2_X1 U14893 ( .A1(n14917), .A2(n14918), .ZN(n14860) );
  NAND2_X1 U14894 ( .A1(n14857), .A2(n14919), .ZN(n14918) );
  INV_X1 U14895 ( .A(n14920), .ZN(n14919) );
  NOR2_X1 U14896 ( .A1(n14856), .A2(n14855), .ZN(n14920) );
  NOR2_X1 U14897 ( .A1(n8555), .A2(n8530), .ZN(n14857) );
  NAND2_X1 U14898 ( .A1(n14855), .A2(n14856), .ZN(n14917) );
  NAND2_X1 U14899 ( .A1(n14921), .A2(n14922), .ZN(n14856) );
  NAND2_X1 U14900 ( .A1(n14853), .A2(n14923), .ZN(n14922) );
  INV_X1 U14901 ( .A(n14924), .ZN(n14923) );
  NOR2_X1 U14902 ( .A1(n14850), .A2(n14852), .ZN(n14924) );
  NOR2_X1 U14903 ( .A1(n8544), .A2(n8530), .ZN(n14853) );
  NAND2_X1 U14904 ( .A1(n14850), .A2(n14852), .ZN(n14921) );
  NAND2_X1 U14905 ( .A1(n14925), .A2(n14926), .ZN(n14852) );
  NAND2_X1 U14906 ( .A1(n14849), .A2(n14927), .ZN(n14926) );
  INV_X1 U14907 ( .A(n14928), .ZN(n14927) );
  NOR2_X1 U14908 ( .A1(n14848), .A2(n14847), .ZN(n14928) );
  NOR2_X1 U14909 ( .A1(n9010), .A2(n8530), .ZN(n14849) );
  NAND2_X1 U14910 ( .A1(n14847), .A2(n14848), .ZN(n14925) );
  NAND2_X1 U14911 ( .A1(n14929), .A2(n14930), .ZN(n14848) );
  NAND2_X1 U14912 ( .A1(n14845), .A2(n14931), .ZN(n14930) );
  NAND2_X1 U14913 ( .A1(n14842), .A2(n14844), .ZN(n14931) );
  NOR2_X1 U14914 ( .A1(n8594), .A2(n8530), .ZN(n14845) );
  INV_X1 U14915 ( .A(n14932), .ZN(n14929) );
  NOR2_X1 U14916 ( .A1(n14842), .A2(n14844), .ZN(n14932) );
  NOR2_X1 U14917 ( .A1(n14933), .A2(n14934), .ZN(n14844) );
  INV_X1 U14918 ( .A(n14935), .ZN(n14934) );
  NAND2_X1 U14919 ( .A1(n14841), .A2(n14936), .ZN(n14935) );
  NAND2_X1 U14920 ( .A1(n14840), .A2(n14839), .ZN(n14936) );
  NOR2_X1 U14921 ( .A1(n9020), .A2(n8530), .ZN(n14841) );
  NOR2_X1 U14922 ( .A1(n14839), .A2(n14840), .ZN(n14933) );
  NOR2_X1 U14923 ( .A1(n14937), .A2(n14938), .ZN(n14840) );
  NOR2_X1 U14924 ( .A1(n14837), .A2(n14939), .ZN(n14938) );
  NOR2_X1 U14925 ( .A1(n14834), .A2(n14836), .ZN(n14939) );
  NAND2_X1 U14926 ( .A1(n9209), .A2(n14543), .ZN(n14837) );
  INV_X1 U14927 ( .A(n14940), .ZN(n14937) );
  NAND2_X1 U14928 ( .A1(n14834), .A2(n14836), .ZN(n14940) );
  NAND2_X1 U14929 ( .A1(n14941), .A2(n14942), .ZN(n14836) );
  NAND2_X1 U14930 ( .A1(n14833), .A2(n14943), .ZN(n14942) );
  INV_X1 U14931 ( .A(n14944), .ZN(n14943) );
  NOR2_X1 U14932 ( .A1(n14830), .A2(n14832), .ZN(n14944) );
  NOR2_X1 U14933 ( .A1(n9031), .A2(n8530), .ZN(n14833) );
  NAND2_X1 U14934 ( .A1(n14830), .A2(n14832), .ZN(n14941) );
  NOR2_X1 U14935 ( .A1(n14945), .A2(n14946), .ZN(n14832) );
  INV_X1 U14936 ( .A(n14947), .ZN(n14946) );
  NAND2_X1 U14937 ( .A1(n14827), .A2(n14948), .ZN(n14947) );
  NAND2_X1 U14938 ( .A1(n14829), .A2(n14828), .ZN(n14948) );
  XNOR2_X1 U14939 ( .A(n14949), .B(n14950), .ZN(n14827) );
  XNOR2_X1 U14940 ( .A(n14951), .B(n14952), .ZN(n14950) );
  NAND2_X1 U14941 ( .A1(n9322), .A2(n14761), .ZN(n14952) );
  NOR2_X1 U14942 ( .A1(n14828), .A2(n14829), .ZN(n14945) );
  NOR2_X1 U14943 ( .A1(n9036), .A2(n8530), .ZN(n14829) );
  NAND2_X1 U14944 ( .A1(n14824), .A2(n14953), .ZN(n14828) );
  NAND2_X1 U14945 ( .A1(n14823), .A2(n14825), .ZN(n14953) );
  NAND2_X1 U14946 ( .A1(n14954), .A2(n14955), .ZN(n14825) );
  NAND2_X1 U14947 ( .A1(n9322), .A2(n14543), .ZN(n14955) );
  INV_X1 U14948 ( .A(n14956), .ZN(n14954) );
  XOR2_X1 U14949 ( .A(n14957), .B(n14958), .Z(n14823) );
  XOR2_X1 U14950 ( .A(n14959), .B(n14960), .Z(n14957) );
  NOR2_X1 U14951 ( .A1(n8534), .A2(n8545), .ZN(n14960) );
  NAND2_X1 U14952 ( .A1(n9322), .A2(n14956), .ZN(n14824) );
  NAND2_X1 U14953 ( .A1(n14820), .A2(n14961), .ZN(n14956) );
  NAND2_X1 U14954 ( .A1(n14819), .A2(n14821), .ZN(n14961) );
  NAND2_X1 U14955 ( .A1(n14962), .A2(n14963), .ZN(n14821) );
  NAND2_X1 U14956 ( .A1(n10222), .A2(n14543), .ZN(n14963) );
  INV_X1 U14957 ( .A(n14964), .ZN(n14962) );
  XNOR2_X1 U14958 ( .A(n14965), .B(n14966), .ZN(n14819) );
  XOR2_X1 U14959 ( .A(n14967), .B(n14968), .Z(n14966) );
  NAND2_X1 U14960 ( .A1(n9331), .A2(n14761), .ZN(n14968) );
  NAND2_X1 U14961 ( .A1(n10222), .A2(n14964), .ZN(n14820) );
  NAND2_X1 U14962 ( .A1(n14816), .A2(n14969), .ZN(n14964) );
  NAND2_X1 U14963 ( .A1(n14815), .A2(n14817), .ZN(n14969) );
  NAND2_X1 U14964 ( .A1(n14970), .A2(n14971), .ZN(n14817) );
  NAND2_X1 U14965 ( .A1(n9331), .A2(n14543), .ZN(n14971) );
  INV_X1 U14966 ( .A(n14972), .ZN(n14970) );
  XNOR2_X1 U14967 ( .A(n14973), .B(n14974), .ZN(n14815) );
  XNOR2_X1 U14968 ( .A(n14975), .B(n14976), .ZN(n14973) );
  NOR2_X1 U14969 ( .A1(n8534), .A2(n8593), .ZN(n14976) );
  NAND2_X1 U14970 ( .A1(n9331), .A2(n14972), .ZN(n14816) );
  NAND2_X1 U14971 ( .A1(n14977), .A2(n14978), .ZN(n14972) );
  INV_X1 U14972 ( .A(n14979), .ZN(n14978) );
  NOR3_X1 U14973 ( .A1(n8530), .A2(n14980), .A3(n8593), .ZN(n14979) );
  NOR2_X1 U14974 ( .A1(n14811), .A2(n14812), .ZN(n14980) );
  NAND2_X1 U14975 ( .A1(n14812), .A2(n14811), .ZN(n14977) );
  XOR2_X1 U14976 ( .A(n14981), .B(n14982), .Z(n14811) );
  XNOR2_X1 U14977 ( .A(n14983), .B(n14984), .ZN(n14982) );
  NAND2_X1 U14978 ( .A1(n9340), .A2(n14761), .ZN(n14984) );
  NOR2_X1 U14979 ( .A1(n14985), .A2(n14986), .ZN(n14812) );
  INV_X1 U14980 ( .A(n14987), .ZN(n14986) );
  NAND2_X1 U14981 ( .A1(n14807), .A2(n14988), .ZN(n14987) );
  NAND2_X1 U14982 ( .A1(n14809), .A2(n14808), .ZN(n14988) );
  XNOR2_X1 U14983 ( .A(n14989), .B(n14990), .ZN(n14807) );
  XNOR2_X1 U14984 ( .A(n14991), .B(n14992), .ZN(n14990) );
  NAND2_X1 U14985 ( .A1(n14761), .A2(n9070), .ZN(n14992) );
  NOR2_X1 U14986 ( .A1(n14808), .A2(n14809), .ZN(n14985) );
  NOR2_X1 U14987 ( .A1(n9061), .A2(n8530), .ZN(n14809) );
  NAND2_X1 U14988 ( .A1(n14804), .A2(n14993), .ZN(n14808) );
  NAND2_X1 U14989 ( .A1(n14803), .A2(n14805), .ZN(n14993) );
  NAND2_X1 U14990 ( .A1(n14994), .A2(n14995), .ZN(n14805) );
  NAND2_X1 U14991 ( .A1(n14543), .A2(n9070), .ZN(n14995) );
  XOR2_X1 U14992 ( .A(n14996), .B(n14997), .Z(n14803) );
  XOR2_X1 U14993 ( .A(n14998), .B(n14999), .Z(n14996) );
  NOR2_X1 U14994 ( .A1(n9076), .A2(n8534), .ZN(n14999) );
  NAND2_X1 U14995 ( .A1(n9070), .A2(n15000), .ZN(n14804) );
  INV_X1 U14996 ( .A(n14994), .ZN(n15000) );
  NOR2_X1 U14997 ( .A1(n15001), .A2(n15002), .ZN(n14994) );
  NOR3_X1 U14998 ( .A1(n9076), .A2(n15003), .A3(n8530), .ZN(n15002) );
  INV_X1 U14999 ( .A(n15004), .ZN(n15003) );
  NAND2_X1 U15000 ( .A1(n14800), .A2(n14799), .ZN(n15004) );
  NOR2_X1 U15001 ( .A1(n14799), .A2(n14800), .ZN(n15001) );
  NOR2_X1 U15002 ( .A1(n15005), .A2(n15006), .ZN(n14800) );
  NOR2_X1 U15003 ( .A1(n14716), .A2(n15007), .ZN(n15006) );
  NOR2_X1 U15004 ( .A1(n14715), .A2(n14713), .ZN(n15007) );
  NAND2_X1 U15005 ( .A1(n14543), .A2(n8515), .ZN(n14716) );
  INV_X1 U15006 ( .A(n15008), .ZN(n15005) );
  NAND2_X1 U15007 ( .A1(n14713), .A2(n14715), .ZN(n15008) );
  NAND2_X1 U15008 ( .A1(n15009), .A2(n15010), .ZN(n14715) );
  NAND3_X1 U15009 ( .A1(n9098), .A2(n15011), .A3(n14543), .ZN(n15010) );
  NAND2_X1 U15010 ( .A1(n14794), .A2(n14796), .ZN(n15011) );
  INV_X1 U15011 ( .A(n15012), .ZN(n15009) );
  NOR2_X1 U15012 ( .A1(n14794), .A2(n14796), .ZN(n15012) );
  NOR2_X1 U15013 ( .A1(n15013), .A2(n15014), .ZN(n14796) );
  INV_X1 U15014 ( .A(n15015), .ZN(n15014) );
  NAND3_X1 U15015 ( .A1(n9107), .A2(n15016), .A3(n14543), .ZN(n15015) );
  NAND2_X1 U15016 ( .A1(n14791), .A2(n14792), .ZN(n15016) );
  NOR2_X1 U15017 ( .A1(n14791), .A2(n14792), .ZN(n15013) );
  NOR2_X1 U15018 ( .A1(n15017), .A2(n15018), .ZN(n14792) );
  INV_X1 U15019 ( .A(n15019), .ZN(n15018) );
  NAND3_X1 U15020 ( .A1(n9112), .A2(n15020), .A3(n14543), .ZN(n15019) );
  NAND2_X1 U15021 ( .A1(n14788), .A2(n14787), .ZN(n15020) );
  NOR2_X1 U15022 ( .A1(n14787), .A2(n14788), .ZN(n15017) );
  NOR2_X1 U15023 ( .A1(n15021), .A2(n15022), .ZN(n14788) );
  INV_X1 U15024 ( .A(n15023), .ZN(n15022) );
  NAND3_X1 U15025 ( .A1(n9121), .A2(n15024), .A3(n14543), .ZN(n15023) );
  NAND2_X1 U15026 ( .A1(n14783), .A2(n14785), .ZN(n15024) );
  NOR2_X1 U15027 ( .A1(n14783), .A2(n14785), .ZN(n15021) );
  NOR2_X1 U15028 ( .A1(n15025), .A2(n15026), .ZN(n14785) );
  INV_X1 U15029 ( .A(n15027), .ZN(n15026) );
  NAND2_X1 U15030 ( .A1(n14781), .A2(n15028), .ZN(n15027) );
  NAND2_X1 U15031 ( .A1(n14780), .A2(n14779), .ZN(n15028) );
  NOR2_X1 U15032 ( .A1(n8530), .A2(n9126), .ZN(n14781) );
  NOR2_X1 U15033 ( .A1(n14779), .A2(n14780), .ZN(n15025) );
  NOR2_X1 U15034 ( .A1(n15029), .A2(n15030), .ZN(n14780) );
  INV_X1 U15035 ( .A(n15031), .ZN(n15030) );
  NAND2_X1 U15036 ( .A1(n14776), .A2(n15032), .ZN(n15031) );
  NAND2_X1 U15037 ( .A1(n14775), .A2(n14777), .ZN(n15032) );
  NOR2_X1 U15038 ( .A1(n8530), .A2(n9378), .ZN(n14776) );
  NOR2_X1 U15039 ( .A1(n14775), .A2(n14777), .ZN(n15029) );
  NOR2_X1 U15040 ( .A1(n15033), .A2(n15034), .ZN(n14777) );
  INV_X1 U15041 ( .A(n15035), .ZN(n15034) );
  NAND2_X1 U15042 ( .A1(n14772), .A2(n15036), .ZN(n15035) );
  NAND2_X1 U15043 ( .A1(n14773), .A2(n14771), .ZN(n15036) );
  NOR2_X1 U15044 ( .A1(n8530), .A2(n8565), .ZN(n14772) );
  NOR2_X1 U15045 ( .A1(n14771), .A2(n14773), .ZN(n15033) );
  NOR2_X1 U15046 ( .A1(n15037), .A2(n15038), .ZN(n14773) );
  INV_X1 U15047 ( .A(n15039), .ZN(n15038) );
  NAND2_X1 U15048 ( .A1(n14766), .A2(n15040), .ZN(n15039) );
  NAND2_X1 U15049 ( .A1(n14769), .A2(n14768), .ZN(n15040) );
  NOR2_X1 U15050 ( .A1(n8530), .A2(n9146), .ZN(n14766) );
  NOR2_X1 U15051 ( .A1(n14768), .A2(n14769), .ZN(n15037) );
  INV_X1 U15052 ( .A(n15041), .ZN(n14769) );
  NAND2_X1 U15053 ( .A1(n15042), .A2(n15043), .ZN(n15041) );
  NAND2_X1 U15054 ( .A1(n14761), .A2(n15044), .ZN(n15043) );
  NAND2_X1 U15055 ( .A1(n8624), .A2(n15045), .ZN(n15044) );
  NAND2_X1 U15056 ( .A1(n8554), .A2(n8627), .ZN(n15045) );
  NAND2_X1 U15057 ( .A1(n15047), .A2(n15048), .ZN(n15042) );
  NAND2_X1 U15058 ( .A1(n8630), .A2(n15049), .ZN(n15048) );
  NAND2_X1 U15059 ( .A1(n8539), .A2(n8534), .ZN(n15049) );
  NAND3_X1 U15060 ( .A1(n14543), .A2(n8537), .A3(n14761), .ZN(n14768) );
  INV_X1 U15061 ( .A(n8530), .ZN(n14543) );
  XOR2_X1 U15062 ( .A(d_8_), .B(c_8_), .Z(n15051) );
  XOR2_X1 U15063 ( .A(n15052), .B(n15053), .Z(n14771) );
  XNOR2_X1 U15064 ( .A(n15054), .B(n15055), .ZN(n15053) );
  XOR2_X1 U15065 ( .A(n15056), .B(n15057), .Z(n14775) );
  XNOR2_X1 U15066 ( .A(n15058), .B(n15059), .ZN(n15056) );
  XOR2_X1 U15067 ( .A(n15060), .B(n15061), .Z(n14779) );
  XNOR2_X1 U15068 ( .A(n15062), .B(n15063), .ZN(n15060) );
  XNOR2_X1 U15069 ( .A(n15064), .B(n15065), .ZN(n14783) );
  XOR2_X1 U15070 ( .A(n15066), .B(n15067), .Z(n15064) );
  XOR2_X1 U15071 ( .A(n15068), .B(n15069), .Z(n14787) );
  XNOR2_X1 U15072 ( .A(n15070), .B(n15071), .ZN(n15068) );
  XOR2_X1 U15073 ( .A(n15072), .B(n15073), .Z(n14791) );
  XNOR2_X1 U15074 ( .A(n15074), .B(n15075), .ZN(n15072) );
  XOR2_X1 U15075 ( .A(n15076), .B(n15077), .Z(n14794) );
  XNOR2_X1 U15076 ( .A(n15078), .B(n15079), .ZN(n15076) );
  XNOR2_X1 U15077 ( .A(n15080), .B(n15081), .ZN(n14713) );
  NAND2_X1 U15078 ( .A1(n15082), .A2(n15083), .ZN(n15080) );
  XOR2_X1 U15079 ( .A(n15084), .B(n15085), .Z(n14799) );
  XOR2_X1 U15080 ( .A(n15086), .B(n15087), .Z(n15085) );
  NAND2_X1 U15081 ( .A1(n14761), .A2(n8515), .ZN(n15087) );
  XOR2_X1 U15082 ( .A(n15088), .B(n15089), .Z(n14830) );
  XOR2_X1 U15083 ( .A(n15090), .B(n15091), .Z(n15088) );
  NOR2_X1 U15084 ( .A1(n8534), .A2(n8591), .ZN(n15091) );
  XNOR2_X1 U15085 ( .A(n15092), .B(n15093), .ZN(n14834) );
  XOR2_X1 U15086 ( .A(n15094), .B(n15095), .Z(n15093) );
  NAND2_X1 U15087 ( .A1(n9313), .A2(n14761), .ZN(n15095) );
  XNOR2_X1 U15088 ( .A(n15096), .B(n15097), .ZN(n14839) );
  XOR2_X1 U15089 ( .A(n15098), .B(n15099), .Z(n15096) );
  NOR2_X1 U15090 ( .A1(n8534), .A2(n8572), .ZN(n15099) );
  XOR2_X1 U15091 ( .A(n15100), .B(n15101), .Z(n14842) );
  XOR2_X1 U15092 ( .A(n15102), .B(n15103), .Z(n15101) );
  NAND2_X1 U15093 ( .A1(n9304), .A2(n14761), .ZN(n15103) );
  XOR2_X1 U15094 ( .A(n15104), .B(n15105), .Z(n14847) );
  XOR2_X1 U15095 ( .A(n15106), .B(n15107), .Z(n15104) );
  NOR2_X1 U15096 ( .A1(n8534), .A2(n8594), .ZN(n15107) );
  XNOR2_X1 U15097 ( .A(n15108), .B(n15109), .ZN(n14850) );
  XOR2_X1 U15098 ( .A(n15110), .B(n15111), .Z(n15109) );
  NAND2_X1 U15099 ( .A1(n9295), .A2(n14761), .ZN(n15111) );
  XOR2_X1 U15100 ( .A(n15112), .B(n15113), .Z(n14855) );
  XOR2_X1 U15101 ( .A(n15114), .B(n15115), .Z(n15112) );
  NOR2_X1 U15102 ( .A1(n8534), .A2(n8544), .ZN(n15115) );
  XNOR2_X1 U15103 ( .A(n15116), .B(n15117), .ZN(n14858) );
  XOR2_X1 U15104 ( .A(n15118), .B(n15119), .Z(n15117) );
  NAND2_X1 U15105 ( .A1(n9286), .A2(n14761), .ZN(n15119) );
  XOR2_X1 U15106 ( .A(n15120), .B(n15121), .Z(n14863) );
  XOR2_X1 U15107 ( .A(n15122), .B(n15123), .Z(n15120) );
  NOR2_X1 U15108 ( .A1(n8534), .A2(n8564), .ZN(n15123) );
  XNOR2_X1 U15109 ( .A(n15124), .B(n15125), .ZN(n14866) );
  XNOR2_X1 U15110 ( .A(n15126), .B(n15127), .ZN(n15125) );
  NAND2_X1 U15111 ( .A1(n9277), .A2(n14761), .ZN(n15127) );
  XNOR2_X1 U15112 ( .A(n15128), .B(n15129), .ZN(n14871) );
  XNOR2_X1 U15113 ( .A(n15130), .B(n15131), .ZN(n15129) );
  NAND2_X1 U15114 ( .A1(n9792), .A2(n14761), .ZN(n15131) );
  XNOR2_X1 U15115 ( .A(n15132), .B(n15133), .ZN(n14874) );
  XNOR2_X1 U15116 ( .A(n15134), .B(n15135), .ZN(n15133) );
  NAND2_X1 U15117 ( .A1(n9268), .A2(n14761), .ZN(n15135) );
  XNOR2_X1 U15118 ( .A(n15136), .B(n15137), .ZN(n14380) );
  XNOR2_X1 U15119 ( .A(n15138), .B(n15139), .ZN(n15137) );
  NAND2_X1 U15120 ( .A1(n9263), .A2(n14761), .ZN(n15139) );
  XNOR2_X1 U15121 ( .A(n14886), .B(n15140), .ZN(n8616) );
  XNOR2_X1 U15122 ( .A(n14887), .B(n15141), .ZN(n15140) );
  NAND2_X1 U15123 ( .A1(n14761), .A2(n8872), .ZN(n15141) );
  NOR2_X1 U15124 ( .A1(n15142), .A2(n15143), .ZN(n14887) );
  INV_X1 U15125 ( .A(n15144), .ZN(n15143) );
  NAND3_X1 U15126 ( .A1(n14761), .A2(n15145), .A3(n9263), .ZN(n15144) );
  NAND2_X1 U15127 ( .A1(n15136), .A2(n15138), .ZN(n15145) );
  NOR2_X1 U15128 ( .A1(n15136), .A2(n15138), .ZN(n15142) );
  NOR2_X1 U15129 ( .A1(n15146), .A2(n15147), .ZN(n15138) );
  INV_X1 U15130 ( .A(n15148), .ZN(n15147) );
  NAND3_X1 U15131 ( .A1(n14761), .A2(n15149), .A3(n9268), .ZN(n15148) );
  NAND2_X1 U15132 ( .A1(n15132), .A2(n15134), .ZN(n15149) );
  NOR2_X1 U15133 ( .A1(n15132), .A2(n15134), .ZN(n15146) );
  NOR2_X1 U15134 ( .A1(n15150), .A2(n15151), .ZN(n15134) );
  INV_X1 U15135 ( .A(n15152), .ZN(n15151) );
  NAND3_X1 U15136 ( .A1(n14761), .A2(n15153), .A3(n9792), .ZN(n15152) );
  NAND2_X1 U15137 ( .A1(n15128), .A2(n15130), .ZN(n15153) );
  NOR2_X1 U15138 ( .A1(n15128), .A2(n15130), .ZN(n15150) );
  NOR2_X1 U15139 ( .A1(n15154), .A2(n15155), .ZN(n15130) );
  INV_X1 U15140 ( .A(n15156), .ZN(n15155) );
  NAND3_X1 U15141 ( .A1(n14761), .A2(n15157), .A3(n9277), .ZN(n15156) );
  NAND2_X1 U15142 ( .A1(n15124), .A2(n15126), .ZN(n15157) );
  NOR2_X1 U15143 ( .A1(n15124), .A2(n15126), .ZN(n15154) );
  NOR2_X1 U15144 ( .A1(n15158), .A2(n15159), .ZN(n15126) );
  NOR3_X1 U15145 ( .A1(n8534), .A2(n15160), .A3(n8564), .ZN(n15159) );
  NOR2_X1 U15146 ( .A1(n15121), .A2(n15122), .ZN(n15160) );
  INV_X1 U15147 ( .A(n15161), .ZN(n15158) );
  NAND2_X1 U15148 ( .A1(n15121), .A2(n15122), .ZN(n15161) );
  NAND2_X1 U15149 ( .A1(n15162), .A2(n15163), .ZN(n15122) );
  INV_X1 U15150 ( .A(n15164), .ZN(n15163) );
  NOR3_X1 U15151 ( .A1(n8534), .A2(n15165), .A3(n8555), .ZN(n15164) );
  NOR2_X1 U15152 ( .A1(n15116), .A2(n15118), .ZN(n15165) );
  NAND2_X1 U15153 ( .A1(n15116), .A2(n15118), .ZN(n15162) );
  NAND2_X1 U15154 ( .A1(n15166), .A2(n15167), .ZN(n15118) );
  NAND3_X1 U15155 ( .A1(n14761), .A2(n15168), .A3(n8543), .ZN(n15167) );
  INV_X1 U15156 ( .A(n15169), .ZN(n15168) );
  NOR2_X1 U15157 ( .A1(n15113), .A2(n15114), .ZN(n15169) );
  NAND2_X1 U15158 ( .A1(n15113), .A2(n15114), .ZN(n15166) );
  NAND2_X1 U15159 ( .A1(n15170), .A2(n15171), .ZN(n15114) );
  INV_X1 U15160 ( .A(n15172), .ZN(n15171) );
  NOR3_X1 U15161 ( .A1(n8534), .A2(n15173), .A3(n8560), .ZN(n15172) );
  NOR2_X1 U15162 ( .A1(n15110), .A2(n15108), .ZN(n15173) );
  NAND2_X1 U15163 ( .A1(n15108), .A2(n15110), .ZN(n15170) );
  NAND2_X1 U15164 ( .A1(n15174), .A2(n15175), .ZN(n15110) );
  NAND3_X1 U15165 ( .A1(n14761), .A2(n15176), .A3(n10846), .ZN(n15175) );
  INV_X1 U15166 ( .A(n15177), .ZN(n15176) );
  NOR2_X1 U15167 ( .A1(n15105), .A2(n15106), .ZN(n15177) );
  NAND2_X1 U15168 ( .A1(n15105), .A2(n15106), .ZN(n15174) );
  NAND2_X1 U15169 ( .A1(n15178), .A2(n15179), .ZN(n15106) );
  INV_X1 U15170 ( .A(n15180), .ZN(n15179) );
  NOR3_X1 U15171 ( .A1(n8534), .A2(n15181), .A3(n8556), .ZN(n15180) );
  NOR2_X1 U15172 ( .A1(n15102), .A2(n15100), .ZN(n15181) );
  NAND2_X1 U15173 ( .A1(n15100), .A2(n15102), .ZN(n15178) );
  NAND2_X1 U15174 ( .A1(n15182), .A2(n15183), .ZN(n15102) );
  NAND3_X1 U15175 ( .A1(n14761), .A2(n15184), .A3(n9209), .ZN(n15183) );
  INV_X1 U15176 ( .A(n15185), .ZN(n15184) );
  NOR2_X1 U15177 ( .A1(n15097), .A2(n15098), .ZN(n15185) );
  NAND2_X1 U15178 ( .A1(n15097), .A2(n15098), .ZN(n15182) );
  NAND2_X1 U15179 ( .A1(n15186), .A2(n15187), .ZN(n15098) );
  INV_X1 U15180 ( .A(n15188), .ZN(n15187) );
  NOR3_X1 U15181 ( .A1(n8534), .A2(n15189), .A3(n8582), .ZN(n15188) );
  NOR2_X1 U15182 ( .A1(n15094), .A2(n15092), .ZN(n15189) );
  NAND2_X1 U15183 ( .A1(n15092), .A2(n15094), .ZN(n15186) );
  NAND2_X1 U15184 ( .A1(n15190), .A2(n15191), .ZN(n15094) );
  NAND3_X1 U15185 ( .A1(n14761), .A2(n15192), .A3(n9721), .ZN(n15191) );
  INV_X1 U15186 ( .A(n15193), .ZN(n15192) );
  NOR2_X1 U15187 ( .A1(n15089), .A2(n15090), .ZN(n15193) );
  NAND2_X1 U15188 ( .A1(n15089), .A2(n15090), .ZN(n15190) );
  NAND2_X1 U15189 ( .A1(n15194), .A2(n15195), .ZN(n15090) );
  NAND3_X1 U15190 ( .A1(n14761), .A2(n15196), .A3(n9322), .ZN(n15195) );
  NAND2_X1 U15191 ( .A1(n14951), .A2(n14949), .ZN(n15196) );
  INV_X1 U15192 ( .A(n15197), .ZN(n15194) );
  NOR2_X1 U15193 ( .A1(n14949), .A2(n14951), .ZN(n15197) );
  NOR2_X1 U15194 ( .A1(n15198), .A2(n15199), .ZN(n14951) );
  NOR3_X1 U15195 ( .A1(n8534), .A2(n15200), .A3(n8545), .ZN(n15199) );
  NOR2_X1 U15196 ( .A1(n14958), .A2(n14959), .ZN(n15200) );
  INV_X1 U15197 ( .A(n15201), .ZN(n15198) );
  NAND2_X1 U15198 ( .A1(n14958), .A2(n14959), .ZN(n15201) );
  NAND2_X1 U15199 ( .A1(n15202), .A2(n15203), .ZN(n14959) );
  NAND3_X1 U15200 ( .A1(n14761), .A2(n15204), .A3(n9331), .ZN(n15203) );
  INV_X1 U15201 ( .A(n15205), .ZN(n15204) );
  NOR2_X1 U15202 ( .A1(n14967), .A2(n14965), .ZN(n15205) );
  NAND2_X1 U15203 ( .A1(n14965), .A2(n14967), .ZN(n15202) );
  NAND2_X1 U15204 ( .A1(n15206), .A2(n15207), .ZN(n14967) );
  NAND3_X1 U15205 ( .A1(n14761), .A2(n15208), .A3(n10722), .ZN(n15207) );
  NAND2_X1 U15206 ( .A1(n14974), .A2(n14975), .ZN(n15208) );
  INV_X1 U15207 ( .A(n15209), .ZN(n15206) );
  NOR2_X1 U15208 ( .A1(n14974), .A2(n14975), .ZN(n15209) );
  NOR2_X1 U15209 ( .A1(n15210), .A2(n15211), .ZN(n14975) );
  NOR3_X1 U15210 ( .A1(n8534), .A2(n15212), .A3(n8583), .ZN(n15211) );
  INV_X1 U15211 ( .A(n15213), .ZN(n15212) );
  NAND2_X1 U15212 ( .A1(n14983), .A2(n14981), .ZN(n15213) );
  NOR2_X1 U15213 ( .A1(n14981), .A2(n14983), .ZN(n15210) );
  NOR2_X1 U15214 ( .A1(n15214), .A2(n15215), .ZN(n14983) );
  INV_X1 U15215 ( .A(n15216), .ZN(n15215) );
  NAND3_X1 U15216 ( .A1(n9070), .A2(n15217), .A3(n14761), .ZN(n15216) );
  NAND2_X1 U15217 ( .A1(n14989), .A2(n14991), .ZN(n15217) );
  NOR2_X1 U15218 ( .A1(n14989), .A2(n14991), .ZN(n15214) );
  NOR2_X1 U15219 ( .A1(n15218), .A2(n15219), .ZN(n14991) );
  NOR3_X1 U15220 ( .A1(n9076), .A2(n15220), .A3(n8534), .ZN(n15219) );
  NOR2_X1 U15221 ( .A1(n14997), .A2(n14998), .ZN(n15220) );
  INV_X1 U15222 ( .A(n15221), .ZN(n15218) );
  NAND2_X1 U15223 ( .A1(n14997), .A2(n14998), .ZN(n15221) );
  NAND2_X1 U15224 ( .A1(n15222), .A2(n15223), .ZN(n14998) );
  INV_X1 U15225 ( .A(n15224), .ZN(n15223) );
  NOR3_X1 U15226 ( .A1(n8551), .A2(n15225), .A3(n8534), .ZN(n15224) );
  NOR2_X1 U15227 ( .A1(n15084), .A2(n15086), .ZN(n15225) );
  NAND2_X1 U15228 ( .A1(n15084), .A2(n15086), .ZN(n15222) );
  NAND2_X1 U15229 ( .A1(n15082), .A2(n15226), .ZN(n15086) );
  NAND2_X1 U15230 ( .A1(n15081), .A2(n15083), .ZN(n15226) );
  NAND2_X1 U15231 ( .A1(n15227), .A2(n15228), .ZN(n15083) );
  NAND2_X1 U15232 ( .A1(n14761), .A2(n9098), .ZN(n15228) );
  XNOR2_X1 U15233 ( .A(n15229), .B(n15230), .ZN(n15081) );
  XOR2_X1 U15234 ( .A(n15231), .B(n15232), .Z(n15230) );
  NAND2_X1 U15235 ( .A1(n9098), .A2(n15233), .ZN(n15082) );
  INV_X1 U15236 ( .A(n15227), .ZN(n15233) );
  NOR2_X1 U15237 ( .A1(n15234), .A2(n15235), .ZN(n15227) );
  INV_X1 U15238 ( .A(n15236), .ZN(n15235) );
  NAND2_X1 U15239 ( .A1(n15079), .A2(n15237), .ZN(n15236) );
  NAND2_X1 U15240 ( .A1(n15078), .A2(n15077), .ZN(n15237) );
  NOR2_X1 U15241 ( .A1(n8534), .A2(n8548), .ZN(n15079) );
  NOR2_X1 U15242 ( .A1(n15077), .A2(n15078), .ZN(n15234) );
  NOR2_X1 U15243 ( .A1(n15238), .A2(n15239), .ZN(n15078) );
  INV_X1 U15244 ( .A(n15240), .ZN(n15239) );
  NAND2_X1 U15245 ( .A1(n15075), .A2(n15241), .ZN(n15240) );
  NAND2_X1 U15246 ( .A1(n15074), .A2(n15073), .ZN(n15241) );
  NOR2_X1 U15247 ( .A1(n8534), .A2(n8584), .ZN(n15075) );
  NOR2_X1 U15248 ( .A1(n15073), .A2(n15074), .ZN(n15238) );
  NOR2_X1 U15249 ( .A1(n15242), .A2(n15243), .ZN(n15074) );
  INV_X1 U15250 ( .A(n15244), .ZN(n15243) );
  NAND2_X1 U15251 ( .A1(n15071), .A2(n15245), .ZN(n15244) );
  NAND2_X1 U15252 ( .A1(n15069), .A2(n15070), .ZN(n15245) );
  NOR2_X1 U15253 ( .A1(n8534), .A2(n8535), .ZN(n15071) );
  NOR2_X1 U15254 ( .A1(n15069), .A2(n15070), .ZN(n15242) );
  INV_X1 U15255 ( .A(n15246), .ZN(n15070) );
  NAND2_X1 U15256 ( .A1(n15247), .A2(n15248), .ZN(n15246) );
  NAND2_X1 U15257 ( .A1(n15067), .A2(n15249), .ZN(n15248) );
  INV_X1 U15258 ( .A(n15250), .ZN(n15249) );
  NOR2_X1 U15259 ( .A1(n15066), .A2(n15065), .ZN(n15250) );
  NOR2_X1 U15260 ( .A1(n8534), .A2(n9126), .ZN(n15067) );
  NAND2_X1 U15261 ( .A1(n15065), .A2(n15066), .ZN(n15247) );
  NAND2_X1 U15262 ( .A1(n15251), .A2(n15252), .ZN(n15066) );
  NAND2_X1 U15263 ( .A1(n15063), .A2(n15253), .ZN(n15252) );
  NAND2_X1 U15264 ( .A1(n15061), .A2(n15062), .ZN(n15253) );
  NOR2_X1 U15265 ( .A1(n8534), .A2(n9378), .ZN(n15063) );
  INV_X1 U15266 ( .A(n15254), .ZN(n15251) );
  NOR2_X1 U15267 ( .A1(n15061), .A2(n15062), .ZN(n15254) );
  NOR2_X1 U15268 ( .A1(n15255), .A2(n15256), .ZN(n15062) );
  INV_X1 U15269 ( .A(n15257), .ZN(n15256) );
  NAND2_X1 U15270 ( .A1(n15058), .A2(n15258), .ZN(n15257) );
  NAND2_X1 U15271 ( .A1(n15059), .A2(n15057), .ZN(n15258) );
  NOR2_X1 U15272 ( .A1(n8534), .A2(n9383), .ZN(n15058) );
  NOR2_X1 U15273 ( .A1(n15057), .A2(n15059), .ZN(n15255) );
  NOR2_X1 U15274 ( .A1(n15259), .A2(n15260), .ZN(n15059) );
  INV_X1 U15275 ( .A(n15261), .ZN(n15260) );
  NAND2_X1 U15276 ( .A1(n15052), .A2(n15262), .ZN(n15261) );
  NAND2_X1 U15277 ( .A1(n15055), .A2(n15054), .ZN(n15262) );
  NOR2_X1 U15278 ( .A1(n8534), .A2(n9146), .ZN(n15052) );
  NOR2_X1 U15279 ( .A1(n15054), .A2(n15055), .ZN(n15259) );
  INV_X1 U15280 ( .A(n15263), .ZN(n15055) );
  NAND2_X1 U15281 ( .A1(n15264), .A2(n15265), .ZN(n15263) );
  NAND2_X1 U15282 ( .A1(n15047), .A2(n15266), .ZN(n15265) );
  NAND2_X1 U15283 ( .A1(n8624), .A2(n15267), .ZN(n15266) );
  NAND2_X1 U15284 ( .A1(n8529), .A2(n8627), .ZN(n15267) );
  NAND2_X1 U15285 ( .A1(n15268), .A2(n15269), .ZN(n15264) );
  NAND2_X1 U15286 ( .A1(n8630), .A2(n15270), .ZN(n15269) );
  NAND2_X1 U15287 ( .A1(n8539), .A2(n8554), .ZN(n15270) );
  NAND3_X1 U15288 ( .A1(n14761), .A2(n8537), .A3(n15047), .ZN(n15054) );
  XOR2_X1 U15289 ( .A(d_7_), .B(c_7_), .Z(n15272) );
  XOR2_X1 U15290 ( .A(n15273), .B(n15274), .Z(n15057) );
  XNOR2_X1 U15291 ( .A(n15275), .B(n15276), .ZN(n15274) );
  XOR2_X1 U15292 ( .A(n15277), .B(n15278), .Z(n15061) );
  XNOR2_X1 U15293 ( .A(n15279), .B(n15280), .ZN(n15277) );
  XNOR2_X1 U15294 ( .A(n15281), .B(n15282), .ZN(n15065) );
  XNOR2_X1 U15295 ( .A(n15283), .B(n15284), .ZN(n15281) );
  XOR2_X1 U15296 ( .A(n15285), .B(n15286), .Z(n15069) );
  XNOR2_X1 U15297 ( .A(n15287), .B(n15288), .ZN(n15285) );
  XOR2_X1 U15298 ( .A(n15289), .B(n15290), .Z(n15073) );
  XOR2_X1 U15299 ( .A(n15291), .B(n15292), .Z(n15289) );
  NAND2_X1 U15300 ( .A1(n15047), .A2(n9121), .ZN(n15291) );
  XNOR2_X1 U15301 ( .A(n15293), .B(n15294), .ZN(n15077) );
  XNOR2_X1 U15302 ( .A(n15295), .B(n15296), .ZN(n15294) );
  NAND2_X1 U15303 ( .A1(n15047), .A2(n9112), .ZN(n15296) );
  XNOR2_X1 U15304 ( .A(n15297), .B(n15298), .ZN(n15084) );
  XOR2_X1 U15305 ( .A(n15299), .B(n15300), .Z(n15297) );
  NAND2_X1 U15306 ( .A1(n15047), .A2(n9098), .ZN(n15299) );
  XNOR2_X1 U15307 ( .A(n15301), .B(n15302), .ZN(n14997) );
  NAND2_X1 U15308 ( .A1(n15303), .A2(n15304), .ZN(n15301) );
  XOR2_X1 U15309 ( .A(n15305), .B(n15306), .Z(n14989) );
  XOR2_X1 U15310 ( .A(n15307), .B(n15308), .Z(n15305) );
  XOR2_X1 U15311 ( .A(n15309), .B(n15310), .Z(n14981) );
  NAND2_X1 U15312 ( .A1(n15311), .A2(n15312), .ZN(n15309) );
  XOR2_X1 U15313 ( .A(n15313), .B(n15314), .Z(n14974) );
  XOR2_X1 U15314 ( .A(n15315), .B(n15316), .Z(n15314) );
  NAND2_X1 U15315 ( .A1(n9340), .A2(n15047), .ZN(n15316) );
  XNOR2_X1 U15316 ( .A(n15317), .B(n15318), .ZN(n14965) );
  NAND2_X1 U15317 ( .A1(n15319), .A2(n15320), .ZN(n15317) );
  XOR2_X1 U15318 ( .A(n15321), .B(n15322), .Z(n14958) );
  XOR2_X1 U15319 ( .A(n15323), .B(n15324), .Z(n15321) );
  NOR2_X1 U15320 ( .A1(n8554), .A2(n8569), .ZN(n15324) );
  XOR2_X1 U15321 ( .A(n15325), .B(n15326), .Z(n14949) );
  NAND2_X1 U15322 ( .A1(n15327), .A2(n15328), .ZN(n15325) );
  XOR2_X1 U15323 ( .A(n15329), .B(n15330), .Z(n15089) );
  XOR2_X1 U15324 ( .A(n15331), .B(n15332), .Z(n15329) );
  NOR2_X1 U15325 ( .A1(n8554), .A2(n8562), .ZN(n15332) );
  XNOR2_X1 U15326 ( .A(n15333), .B(n15334), .ZN(n15092) );
  NAND2_X1 U15327 ( .A1(n15335), .A2(n15336), .ZN(n15333) );
  XOR2_X1 U15328 ( .A(n15337), .B(n15338), .Z(n15097) );
  XOR2_X1 U15329 ( .A(n15339), .B(n15340), .Z(n15337) );
  NOR2_X1 U15330 ( .A1(n8554), .A2(n8582), .ZN(n15340) );
  XNOR2_X1 U15331 ( .A(n15341), .B(n15342), .ZN(n15100) );
  NAND2_X1 U15332 ( .A1(n15343), .A2(n15344), .ZN(n15341) );
  XOR2_X1 U15333 ( .A(n15345), .B(n15346), .Z(n15105) );
  XOR2_X1 U15334 ( .A(n15347), .B(n15348), .Z(n15345) );
  NOR2_X1 U15335 ( .A1(n8554), .A2(n8556), .ZN(n15348) );
  XNOR2_X1 U15336 ( .A(n15349), .B(n15350), .ZN(n15108) );
  NAND2_X1 U15337 ( .A1(n15351), .A2(n15352), .ZN(n15349) );
  XOR2_X1 U15338 ( .A(n15353), .B(n15354), .Z(n15113) );
  XOR2_X1 U15339 ( .A(n15355), .B(n15356), .Z(n15353) );
  NOR2_X1 U15340 ( .A1(n8554), .A2(n8560), .ZN(n15356) );
  XOR2_X1 U15341 ( .A(n15357), .B(n15358), .Z(n15116) );
  XOR2_X1 U15342 ( .A(n15359), .B(n15360), .Z(n15358) );
  XOR2_X1 U15343 ( .A(n15361), .B(n15362), .Z(n15121) );
  XOR2_X1 U15344 ( .A(n15363), .B(n15364), .Z(n15361) );
  XNOR2_X1 U15345 ( .A(n15365), .B(n15366), .ZN(n15124) );
  XNOR2_X1 U15346 ( .A(n15367), .B(n15368), .ZN(n15366) );
  XOR2_X1 U15347 ( .A(n15369), .B(n15370), .Z(n15128) );
  XNOR2_X1 U15348 ( .A(n15371), .B(n15372), .ZN(n15369) );
  XNOR2_X1 U15349 ( .A(n15373), .B(n15374), .ZN(n15132) );
  XOR2_X1 U15350 ( .A(n15375), .B(n15376), .Z(n15374) );
  XOR2_X1 U15351 ( .A(n15377), .B(n15378), .Z(n15136) );
  XNOR2_X1 U15352 ( .A(n15379), .B(n15380), .ZN(n15377) );
  XNOR2_X1 U15353 ( .A(n15381), .B(n15382), .ZN(n14886) );
  XOR2_X1 U15354 ( .A(n15383), .B(n15384), .Z(n15382) );
  XOR2_X1 U15355 ( .A(n8648), .B(n8649), .Z(n8617) );
  NOR3_X1 U15356 ( .A1(n8649), .A2(n8648), .A3(n8647), .ZN(n8643) );
  NAND2_X1 U15357 ( .A1(n15385), .A2(n8891), .ZN(n8647) );
  INV_X1 U15358 ( .A(n15386), .ZN(n8891) );
  NOR2_X1 U15359 ( .A1(n15387), .A2(n15388), .ZN(n15386) );
  NAND2_X1 U15360 ( .A1(n15387), .A2(n15388), .ZN(n15385) );
  NOR2_X1 U15361 ( .A1(n15389), .A2(n15390), .ZN(n15388) );
  INV_X1 U15362 ( .A(n15391), .ZN(n15390) );
  NAND3_X1 U15363 ( .A1(n8592), .A2(n15392), .A3(n15268), .ZN(n15391) );
  NAND2_X1 U15364 ( .A1(n15393), .A2(n15394), .ZN(n15392) );
  NOR2_X1 U15365 ( .A1(n15393), .A2(n15394), .ZN(n15389) );
  XNOR2_X1 U15366 ( .A(n15395), .B(n15396), .ZN(n15387) );
  XOR2_X1 U15367 ( .A(n15397), .B(n15398), .Z(n15395) );
  NOR2_X1 U15368 ( .A1(n15399), .A2(n15400), .ZN(n8648) );
  INV_X1 U15369 ( .A(n15401), .ZN(n15400) );
  NAND2_X1 U15370 ( .A1(n14891), .A2(n15402), .ZN(n15401) );
  NAND2_X1 U15371 ( .A1(n14890), .A2(n14889), .ZN(n15402) );
  NOR2_X1 U15372 ( .A1(n8554), .A2(n8972), .ZN(n14891) );
  NOR2_X1 U15373 ( .A1(n14889), .A2(n14890), .ZN(n15399) );
  NOR2_X1 U15374 ( .A1(n15403), .A2(n15404), .ZN(n14890) );
  INV_X1 U15375 ( .A(n15405), .ZN(n15404) );
  NAND2_X1 U15376 ( .A1(n15384), .A2(n15406), .ZN(n15405) );
  NAND2_X1 U15377 ( .A1(n15383), .A2(n15381), .ZN(n15406) );
  NOR2_X1 U15378 ( .A1(n8589), .A2(n8554), .ZN(n15384) );
  NOR2_X1 U15379 ( .A1(n15381), .A2(n15383), .ZN(n15403) );
  NOR2_X1 U15380 ( .A1(n15407), .A2(n15408), .ZN(n15383) );
  INV_X1 U15381 ( .A(n15409), .ZN(n15408) );
  NAND2_X1 U15382 ( .A1(n15380), .A2(n15410), .ZN(n15409) );
  NAND2_X1 U15383 ( .A1(n15379), .A2(n15378), .ZN(n15410) );
  NOR2_X1 U15384 ( .A1(n8982), .A2(n8554), .ZN(n15380) );
  NOR2_X1 U15385 ( .A1(n15378), .A2(n15379), .ZN(n15407) );
  NOR2_X1 U15386 ( .A1(n15411), .A2(n15412), .ZN(n15379) );
  INV_X1 U15387 ( .A(n15413), .ZN(n15412) );
  NAND2_X1 U15388 ( .A1(n15376), .A2(n15414), .ZN(n15413) );
  NAND2_X1 U15389 ( .A1(n15375), .A2(n15373), .ZN(n15414) );
  NOR2_X1 U15390 ( .A1(n8527), .A2(n8554), .ZN(n15376) );
  NOR2_X1 U15391 ( .A1(n15373), .A2(n15375), .ZN(n15411) );
  NOR2_X1 U15392 ( .A1(n15415), .A2(n15416), .ZN(n15375) );
  INV_X1 U15393 ( .A(n15417), .ZN(n15416) );
  NAND2_X1 U15394 ( .A1(n15372), .A2(n15418), .ZN(n15417) );
  NAND2_X1 U15395 ( .A1(n15371), .A2(n15370), .ZN(n15418) );
  NOR2_X1 U15396 ( .A1(n8528), .A2(n8554), .ZN(n15372) );
  NOR2_X1 U15397 ( .A1(n15370), .A2(n15371), .ZN(n15415) );
  NOR2_X1 U15398 ( .A1(n15419), .A2(n15420), .ZN(n15371) );
  INV_X1 U15399 ( .A(n15421), .ZN(n15420) );
  NAND2_X1 U15400 ( .A1(n15368), .A2(n15422), .ZN(n15421) );
  NAND2_X1 U15401 ( .A1(n15423), .A2(n15365), .ZN(n15422) );
  NOR2_X1 U15402 ( .A1(n8995), .A2(n8554), .ZN(n15368) );
  NOR2_X1 U15403 ( .A1(n15365), .A2(n15423), .ZN(n15419) );
  INV_X1 U15404 ( .A(n15367), .ZN(n15423) );
  NAND2_X1 U15405 ( .A1(n15424), .A2(n15425), .ZN(n15367) );
  NAND2_X1 U15406 ( .A1(n15363), .A2(n15426), .ZN(n15425) );
  INV_X1 U15407 ( .A(n15427), .ZN(n15426) );
  NOR2_X1 U15408 ( .A1(n15364), .A2(n15362), .ZN(n15427) );
  NOR2_X1 U15409 ( .A1(n8555), .A2(n8554), .ZN(n15363) );
  NAND2_X1 U15410 ( .A1(n15362), .A2(n15364), .ZN(n15424) );
  NAND2_X1 U15411 ( .A1(n15428), .A2(n15429), .ZN(n15364) );
  NAND2_X1 U15412 ( .A1(n15360), .A2(n15430), .ZN(n15429) );
  NAND2_X1 U15413 ( .A1(n15359), .A2(n15357), .ZN(n15430) );
  NOR2_X1 U15414 ( .A1(n8544), .A2(n8554), .ZN(n15360) );
  INV_X1 U15415 ( .A(n15431), .ZN(n15428) );
  NOR2_X1 U15416 ( .A1(n15357), .A2(n15359), .ZN(n15431) );
  NOR2_X1 U15417 ( .A1(n15432), .A2(n15433), .ZN(n15359) );
  NOR3_X1 U15418 ( .A1(n15046), .A2(n15434), .A3(n8560), .ZN(n15433) );
  NOR2_X1 U15419 ( .A1(n15355), .A2(n15354), .ZN(n15434) );
  INV_X1 U15420 ( .A(n15435), .ZN(n15432) );
  NAND2_X1 U15421 ( .A1(n15354), .A2(n15355), .ZN(n15435) );
  NAND2_X1 U15422 ( .A1(n15351), .A2(n15436), .ZN(n15355) );
  NAND2_X1 U15423 ( .A1(n15350), .A2(n15352), .ZN(n15436) );
  NAND2_X1 U15424 ( .A1(n15437), .A2(n15438), .ZN(n15352) );
  NAND2_X1 U15425 ( .A1(n10846), .A2(n15047), .ZN(n15438) );
  XNOR2_X1 U15426 ( .A(n15439), .B(n15440), .ZN(n15350) );
  XOR2_X1 U15427 ( .A(n15441), .B(n15442), .Z(n15440) );
  NAND2_X1 U15428 ( .A1(n9304), .A2(n15268), .ZN(n15442) );
  INV_X1 U15429 ( .A(n15443), .ZN(n15351) );
  NOR2_X1 U15430 ( .A1(n8594), .A2(n15437), .ZN(n15443) );
  NOR2_X1 U15431 ( .A1(n15444), .A2(n15445), .ZN(n15437) );
  NOR3_X1 U15432 ( .A1(n15046), .A2(n15446), .A3(n8556), .ZN(n15445) );
  NOR2_X1 U15433 ( .A1(n15347), .A2(n15346), .ZN(n15446) );
  INV_X1 U15434 ( .A(n15447), .ZN(n15444) );
  NAND2_X1 U15435 ( .A1(n15346), .A2(n15347), .ZN(n15447) );
  NAND2_X1 U15436 ( .A1(n15343), .A2(n15448), .ZN(n15347) );
  NAND2_X1 U15437 ( .A1(n15342), .A2(n15344), .ZN(n15448) );
  NAND2_X1 U15438 ( .A1(n15449), .A2(n15450), .ZN(n15344) );
  NAND2_X1 U15439 ( .A1(n9209), .A2(n15047), .ZN(n15450) );
  XNOR2_X1 U15440 ( .A(n15451), .B(n15452), .ZN(n15342) );
  XOR2_X1 U15441 ( .A(n15453), .B(n15454), .Z(n15452) );
  NAND2_X1 U15442 ( .A1(n9313), .A2(n15268), .ZN(n15454) );
  INV_X1 U15443 ( .A(n15455), .ZN(n15343) );
  NOR2_X1 U15444 ( .A1(n9025), .A2(n15449), .ZN(n15455) );
  NOR2_X1 U15445 ( .A1(n15456), .A2(n15457), .ZN(n15449) );
  NOR3_X1 U15446 ( .A1(n15046), .A2(n15458), .A3(n8582), .ZN(n15457) );
  NOR2_X1 U15447 ( .A1(n15339), .A2(n15338), .ZN(n15458) );
  INV_X1 U15448 ( .A(n15459), .ZN(n15456) );
  NAND2_X1 U15449 ( .A1(n15338), .A2(n15339), .ZN(n15459) );
  NAND2_X1 U15450 ( .A1(n15335), .A2(n15460), .ZN(n15339) );
  NAND2_X1 U15451 ( .A1(n15334), .A2(n15336), .ZN(n15460) );
  NAND2_X1 U15452 ( .A1(n15461), .A2(n15462), .ZN(n15336) );
  NAND2_X1 U15453 ( .A1(n9721), .A2(n15047), .ZN(n15462) );
  XNOR2_X1 U15454 ( .A(n15463), .B(n15464), .ZN(n15334) );
  XOR2_X1 U15455 ( .A(n15465), .B(n15466), .Z(n15464) );
  NAND2_X1 U15456 ( .A1(n9322), .A2(n15268), .ZN(n15466) );
  INV_X1 U15457 ( .A(n15467), .ZN(n15335) );
  NOR2_X1 U15458 ( .A1(n9036), .A2(n15461), .ZN(n15467) );
  NOR2_X1 U15459 ( .A1(n15468), .A2(n15469), .ZN(n15461) );
  NOR3_X1 U15460 ( .A1(n15046), .A2(n15470), .A3(n8562), .ZN(n15469) );
  NOR2_X1 U15461 ( .A1(n15331), .A2(n15330), .ZN(n15470) );
  INV_X1 U15462 ( .A(n15471), .ZN(n15468) );
  NAND2_X1 U15463 ( .A1(n15330), .A2(n15331), .ZN(n15471) );
  NAND2_X1 U15464 ( .A1(n15327), .A2(n15472), .ZN(n15331) );
  NAND2_X1 U15465 ( .A1(n15326), .A2(n15328), .ZN(n15472) );
  NAND2_X1 U15466 ( .A1(n15473), .A2(n15474), .ZN(n15328) );
  NAND2_X1 U15467 ( .A1(n10222), .A2(n15047), .ZN(n15474) );
  XNOR2_X1 U15468 ( .A(n15475), .B(n15476), .ZN(n15326) );
  XOR2_X1 U15469 ( .A(n15477), .B(n15478), .Z(n15476) );
  NAND2_X1 U15470 ( .A1(n9331), .A2(n15268), .ZN(n15478) );
  INV_X1 U15471 ( .A(n15479), .ZN(n15327) );
  NOR2_X1 U15472 ( .A1(n8545), .A2(n15473), .ZN(n15479) );
  NOR2_X1 U15473 ( .A1(n15480), .A2(n15481), .ZN(n15473) );
  NOR3_X1 U15474 ( .A1(n15046), .A2(n15482), .A3(n8569), .ZN(n15481) );
  NOR2_X1 U15475 ( .A1(n15323), .A2(n15322), .ZN(n15482) );
  INV_X1 U15476 ( .A(n15483), .ZN(n15480) );
  NAND2_X1 U15477 ( .A1(n15322), .A2(n15323), .ZN(n15483) );
  NAND2_X1 U15478 ( .A1(n15319), .A2(n15484), .ZN(n15323) );
  NAND2_X1 U15479 ( .A1(n15318), .A2(n15320), .ZN(n15484) );
  NAND2_X1 U15480 ( .A1(n15485), .A2(n15486), .ZN(n15320) );
  NAND2_X1 U15481 ( .A1(n10722), .A2(n15047), .ZN(n15486) );
  XNOR2_X1 U15482 ( .A(n15487), .B(n15488), .ZN(n15318) );
  XOR2_X1 U15483 ( .A(n15489), .B(n15490), .Z(n15488) );
  NAND2_X1 U15484 ( .A1(n9340), .A2(n15268), .ZN(n15490) );
  INV_X1 U15485 ( .A(n15491), .ZN(n15319) );
  NOR2_X1 U15486 ( .A1(n8593), .A2(n15485), .ZN(n15491) );
  NOR2_X1 U15487 ( .A1(n15492), .A2(n15493), .ZN(n15485) );
  NOR3_X1 U15488 ( .A1(n15046), .A2(n15494), .A3(n8583), .ZN(n15493) );
  NOR2_X1 U15489 ( .A1(n15315), .A2(n15313), .ZN(n15494) );
  INV_X1 U15490 ( .A(n15495), .ZN(n15492) );
  NAND2_X1 U15491 ( .A1(n15313), .A2(n15315), .ZN(n15495) );
  NAND2_X1 U15492 ( .A1(n15311), .A2(n15496), .ZN(n15315) );
  NAND2_X1 U15493 ( .A1(n15310), .A2(n15312), .ZN(n15496) );
  NAND2_X1 U15494 ( .A1(n15497), .A2(n15498), .ZN(n15312) );
  NAND2_X1 U15495 ( .A1(n15047), .A2(n9070), .ZN(n15497) );
  XNOR2_X1 U15496 ( .A(n15499), .B(n15500), .ZN(n15310) );
  XOR2_X1 U15497 ( .A(n15501), .B(n15502), .Z(n15500) );
  NAND2_X1 U15498 ( .A1(n15268), .A2(n9080), .ZN(n15502) );
  INV_X1 U15499 ( .A(n15503), .ZN(n15311) );
  NOR2_X1 U15500 ( .A1(n15498), .A2(n8580), .ZN(n15503) );
  NAND2_X1 U15501 ( .A1(n15504), .A2(n15505), .ZN(n15498) );
  NAND2_X1 U15502 ( .A1(n15306), .A2(n15506), .ZN(n15505) );
  NAND2_X1 U15503 ( .A1(n15308), .A2(n15307), .ZN(n15506) );
  XNOR2_X1 U15504 ( .A(n15507), .B(n15508), .ZN(n15306) );
  XOR2_X1 U15505 ( .A(n15509), .B(n15510), .Z(n15507) );
  NOR2_X1 U15506 ( .A1(n8551), .A2(n8529), .ZN(n15510) );
  INV_X1 U15507 ( .A(n15511), .ZN(n15504) );
  NOR2_X1 U15508 ( .A1(n15307), .A2(n15308), .ZN(n15511) );
  NOR2_X1 U15509 ( .A1(n8554), .A2(n8588), .ZN(n15308) );
  NAND2_X1 U15510 ( .A1(n15303), .A2(n15512), .ZN(n15307) );
  NAND2_X1 U15511 ( .A1(n15302), .A2(n15304), .ZN(n15512) );
  NAND2_X1 U15512 ( .A1(n15513), .A2(n15514), .ZN(n15304) );
  NAND2_X1 U15513 ( .A1(n15047), .A2(n8515), .ZN(n15514) );
  XNOR2_X1 U15514 ( .A(n15515), .B(n15516), .ZN(n15302) );
  XOR2_X1 U15515 ( .A(n15517), .B(n15518), .Z(n15516) );
  NAND2_X1 U15516 ( .A1(n15268), .A2(n9098), .ZN(n15518) );
  NAND2_X1 U15517 ( .A1(n8515), .A2(n15519), .ZN(n15303) );
  INV_X1 U15518 ( .A(n15513), .ZN(n15519) );
  NOR2_X1 U15519 ( .A1(n15520), .A2(n15521), .ZN(n15513) );
  NOR3_X1 U15520 ( .A1(n9094), .A2(n15522), .A3(n8554), .ZN(n15521) );
  INV_X1 U15521 ( .A(n15523), .ZN(n15522) );
  NAND2_X1 U15522 ( .A1(n15300), .A2(n15298), .ZN(n15523) );
  NOR2_X1 U15523 ( .A1(n15298), .A2(n15300), .ZN(n15520) );
  NOR2_X1 U15524 ( .A1(n15524), .A2(n15525), .ZN(n15300) );
  NOR2_X1 U15525 ( .A1(n15232), .A2(n15526), .ZN(n15525) );
  NOR2_X1 U15526 ( .A1(n15229), .A2(n15231), .ZN(n15526) );
  NAND2_X1 U15527 ( .A1(n15047), .A2(n9107), .ZN(n15232) );
  INV_X1 U15528 ( .A(n15527), .ZN(n15524) );
  NAND2_X1 U15529 ( .A1(n15229), .A2(n15231), .ZN(n15527) );
  NAND2_X1 U15530 ( .A1(n15528), .A2(n15529), .ZN(n15231) );
  NAND3_X1 U15531 ( .A1(n9112), .A2(n15530), .A3(n15047), .ZN(n15529) );
  NAND2_X1 U15532 ( .A1(n15293), .A2(n15295), .ZN(n15530) );
  INV_X1 U15533 ( .A(n15531), .ZN(n15528) );
  NOR2_X1 U15534 ( .A1(n15293), .A2(n15295), .ZN(n15531) );
  NOR2_X1 U15535 ( .A1(n15532), .A2(n15533), .ZN(n15295) );
  INV_X1 U15536 ( .A(n15534), .ZN(n15533) );
  NAND3_X1 U15537 ( .A1(n9121), .A2(n15535), .A3(n15047), .ZN(n15534) );
  NAND2_X1 U15538 ( .A1(n15290), .A2(n15292), .ZN(n15535) );
  NOR2_X1 U15539 ( .A1(n15290), .A2(n15292), .ZN(n15532) );
  NOR2_X1 U15540 ( .A1(n15536), .A2(n15537), .ZN(n15292) );
  INV_X1 U15541 ( .A(n15538), .ZN(n15537) );
  NAND2_X1 U15542 ( .A1(n15288), .A2(n15539), .ZN(n15538) );
  NAND2_X1 U15543 ( .A1(n15287), .A2(n15286), .ZN(n15539) );
  NOR2_X1 U15544 ( .A1(n8554), .A2(n9126), .ZN(n15288) );
  NOR2_X1 U15545 ( .A1(n15286), .A2(n15287), .ZN(n15536) );
  NOR2_X1 U15546 ( .A1(n15540), .A2(n15541), .ZN(n15287) );
  INV_X1 U15547 ( .A(n15542), .ZN(n15541) );
  NAND2_X1 U15548 ( .A1(n15283), .A2(n15543), .ZN(n15542) );
  NAND2_X1 U15549 ( .A1(n15282), .A2(n15284), .ZN(n15543) );
  NOR2_X1 U15550 ( .A1(n15046), .A2(n9378), .ZN(n15283) );
  NOR2_X1 U15551 ( .A1(n15282), .A2(n15284), .ZN(n15540) );
  NOR2_X1 U15552 ( .A1(n15544), .A2(n15545), .ZN(n15284) );
  INV_X1 U15553 ( .A(n15546), .ZN(n15545) );
  NAND2_X1 U15554 ( .A1(n15279), .A2(n15547), .ZN(n15546) );
  NAND2_X1 U15555 ( .A1(n15280), .A2(n15278), .ZN(n15547) );
  NOR2_X1 U15556 ( .A1(n15046), .A2(n9383), .ZN(n15279) );
  NOR2_X1 U15557 ( .A1(n15278), .A2(n15280), .ZN(n15544) );
  NOR2_X1 U15558 ( .A1(n15548), .A2(n15549), .ZN(n15280) );
  INV_X1 U15559 ( .A(n15550), .ZN(n15549) );
  NAND2_X1 U15560 ( .A1(n15273), .A2(n15551), .ZN(n15550) );
  NAND2_X1 U15561 ( .A1(n15276), .A2(n15275), .ZN(n15551) );
  NOR2_X1 U15562 ( .A1(n15046), .A2(n9146), .ZN(n15273) );
  NOR2_X1 U15563 ( .A1(n15275), .A2(n15276), .ZN(n15548) );
  INV_X1 U15564 ( .A(n15552), .ZN(n15276) );
  NAND2_X1 U15565 ( .A1(n15553), .A2(n15554), .ZN(n15552) );
  NAND2_X1 U15566 ( .A1(n15268), .A2(n15555), .ZN(n15554) );
  NAND2_X1 U15567 ( .A1(n8624), .A2(n15556), .ZN(n15555) );
  NAND2_X1 U15568 ( .A1(n8533), .A2(n8627), .ZN(n15556) );
  NAND2_X1 U15569 ( .A1(n8532), .A2(n15558), .ZN(n15553) );
  NAND2_X1 U15570 ( .A1(n8630), .A2(n15559), .ZN(n15558) );
  NAND2_X1 U15571 ( .A1(n8539), .A2(n8529), .ZN(n15559) );
  NAND3_X1 U15572 ( .A1(n15047), .A2(n8537), .A3(n15268), .ZN(n15275) );
  INV_X1 U15573 ( .A(n15046), .ZN(n15047) );
  XNOR2_X1 U15574 ( .A(n15560), .B(n15561), .ZN(n15046) );
  XOR2_X1 U15575 ( .A(d_6_), .B(c_6_), .Z(n15561) );
  XOR2_X1 U15576 ( .A(n15562), .B(n15563), .Z(n15278) );
  XNOR2_X1 U15577 ( .A(n15564), .B(n15565), .ZN(n15563) );
  XOR2_X1 U15578 ( .A(n15566), .B(n15567), .Z(n15282) );
  XNOR2_X1 U15579 ( .A(n15568), .B(n15569), .ZN(n15566) );
  XOR2_X1 U15580 ( .A(n15570), .B(n15571), .Z(n15286) );
  XNOR2_X1 U15581 ( .A(n15572), .B(n15573), .ZN(n15570) );
  XOR2_X1 U15582 ( .A(n15574), .B(n15575), .Z(n15290) );
  XNOR2_X1 U15583 ( .A(n15576), .B(n15577), .ZN(n15574) );
  XNOR2_X1 U15584 ( .A(n15578), .B(n15579), .ZN(n15293) );
  XOR2_X1 U15585 ( .A(n15580), .B(n15581), .Z(n15579) );
  XNOR2_X1 U15586 ( .A(n15582), .B(n15583), .ZN(n15229) );
  NAND2_X1 U15587 ( .A1(n15584), .A2(n15585), .ZN(n15582) );
  XNOR2_X1 U15588 ( .A(n15586), .B(n15587), .ZN(n15298) );
  XOR2_X1 U15589 ( .A(n15588), .B(n15589), .Z(n15586) );
  NOR2_X1 U15590 ( .A1(n8548), .A2(n8529), .ZN(n15589) );
  XOR2_X1 U15591 ( .A(n15590), .B(n15591), .Z(n15313) );
  XOR2_X1 U15592 ( .A(n15592), .B(n15593), .Z(n15590) );
  NOR2_X1 U15593 ( .A1(n8580), .A2(n8529), .ZN(n15593) );
  XOR2_X1 U15594 ( .A(n15594), .B(n15595), .Z(n15322) );
  XOR2_X1 U15595 ( .A(n15596), .B(n15597), .Z(n15594) );
  NOR2_X1 U15596 ( .A1(n8529), .A2(n8593), .ZN(n15597) );
  XOR2_X1 U15597 ( .A(n15598), .B(n15599), .Z(n15330) );
  XOR2_X1 U15598 ( .A(n15600), .B(n15601), .Z(n15598) );
  NOR2_X1 U15599 ( .A1(n8529), .A2(n8545), .ZN(n15601) );
  XOR2_X1 U15600 ( .A(n15602), .B(n15603), .Z(n15338) );
  XOR2_X1 U15601 ( .A(n15604), .B(n15605), .Z(n15602) );
  NOR2_X1 U15602 ( .A1(n8529), .A2(n8591), .ZN(n15605) );
  XOR2_X1 U15603 ( .A(n15606), .B(n15607), .Z(n15346) );
  XOR2_X1 U15604 ( .A(n15608), .B(n15609), .Z(n15606) );
  NOR2_X1 U15605 ( .A1(n8529), .A2(n8572), .ZN(n15609) );
  XOR2_X1 U15606 ( .A(n15610), .B(n15611), .Z(n15354) );
  XOR2_X1 U15607 ( .A(n15612), .B(n15613), .Z(n15610) );
  NOR2_X1 U15608 ( .A1(n8529), .A2(n8594), .ZN(n15613) );
  XOR2_X1 U15609 ( .A(n15614), .B(n15615), .Z(n15357) );
  XOR2_X1 U15610 ( .A(n15616), .B(n15617), .Z(n15615) );
  NAND2_X1 U15611 ( .A1(n9295), .A2(n15268), .ZN(n15617) );
  XOR2_X1 U15612 ( .A(n15618), .B(n15619), .Z(n15362) );
  XOR2_X1 U15613 ( .A(n15620), .B(n15621), .Z(n15618) );
  NOR2_X1 U15614 ( .A1(n8529), .A2(n8544), .ZN(n15621) );
  XNOR2_X1 U15615 ( .A(n15622), .B(n15623), .ZN(n15365) );
  XNOR2_X1 U15616 ( .A(n15624), .B(n15625), .ZN(n15623) );
  NAND2_X1 U15617 ( .A1(n9286), .A2(n15268), .ZN(n15625) );
  XOR2_X1 U15618 ( .A(n15626), .B(n15627), .Z(n15370) );
  XNOR2_X1 U15619 ( .A(n15628), .B(n15629), .ZN(n15626) );
  NOR2_X1 U15620 ( .A1(n8529), .A2(n8564), .ZN(n15629) );
  XNOR2_X1 U15621 ( .A(n15630), .B(n15631), .ZN(n15373) );
  XNOR2_X1 U15622 ( .A(n15632), .B(n15633), .ZN(n15631) );
  NAND2_X1 U15623 ( .A1(n9277), .A2(n15268), .ZN(n15633) );
  XNOR2_X1 U15624 ( .A(n15634), .B(n15635), .ZN(n15378) );
  XNOR2_X1 U15625 ( .A(n15636), .B(n15637), .ZN(n15635) );
  NAND2_X1 U15626 ( .A1(n9792), .A2(n15268), .ZN(n15637) );
  XNOR2_X1 U15627 ( .A(n15638), .B(n15639), .ZN(n15381) );
  XNOR2_X1 U15628 ( .A(n15640), .B(n15641), .ZN(n15639) );
  NAND2_X1 U15629 ( .A1(n9268), .A2(n15268), .ZN(n15641) );
  XNOR2_X1 U15630 ( .A(n15642), .B(n15643), .ZN(n14889) );
  XNOR2_X1 U15631 ( .A(n15644), .B(n15645), .ZN(n15643) );
  NAND2_X1 U15632 ( .A1(n9263), .A2(n15268), .ZN(n15645) );
  XNOR2_X1 U15633 ( .A(n15393), .B(n15646), .ZN(n8649) );
  XNOR2_X1 U15634 ( .A(n15394), .B(n15647), .ZN(n15646) );
  NAND2_X1 U15635 ( .A1(n15268), .A2(n8872), .ZN(n15647) );
  NOR2_X1 U15636 ( .A1(n15648), .A2(n15649), .ZN(n15394) );
  INV_X1 U15637 ( .A(n15650), .ZN(n15649) );
  NAND3_X1 U15638 ( .A1(n15268), .A2(n15651), .A3(n9263), .ZN(n15650) );
  NAND2_X1 U15639 ( .A1(n15642), .A2(n15644), .ZN(n15651) );
  NOR2_X1 U15640 ( .A1(n15642), .A2(n15644), .ZN(n15648) );
  NOR2_X1 U15641 ( .A1(n15652), .A2(n15653), .ZN(n15644) );
  INV_X1 U15642 ( .A(n15654), .ZN(n15653) );
  NAND3_X1 U15643 ( .A1(n15268), .A2(n15655), .A3(n9268), .ZN(n15654) );
  NAND2_X1 U15644 ( .A1(n15638), .A2(n15640), .ZN(n15655) );
  NOR2_X1 U15645 ( .A1(n15638), .A2(n15640), .ZN(n15652) );
  NOR2_X1 U15646 ( .A1(n15656), .A2(n15657), .ZN(n15640) );
  INV_X1 U15647 ( .A(n15658), .ZN(n15657) );
  NAND3_X1 U15648 ( .A1(n15268), .A2(n15659), .A3(n9792), .ZN(n15658) );
  NAND2_X1 U15649 ( .A1(n15634), .A2(n15636), .ZN(n15659) );
  NOR2_X1 U15650 ( .A1(n15634), .A2(n15636), .ZN(n15656) );
  NOR2_X1 U15651 ( .A1(n15660), .A2(n15661), .ZN(n15636) );
  INV_X1 U15652 ( .A(n15662), .ZN(n15661) );
  NAND3_X1 U15653 ( .A1(n15268), .A2(n15663), .A3(n9277), .ZN(n15662) );
  NAND2_X1 U15654 ( .A1(n15630), .A2(n15632), .ZN(n15663) );
  NOR2_X1 U15655 ( .A1(n15630), .A2(n15632), .ZN(n15660) );
  NOR2_X1 U15656 ( .A1(n15664), .A2(n15665), .ZN(n15632) );
  INV_X1 U15657 ( .A(n15666), .ZN(n15665) );
  NAND3_X1 U15658 ( .A1(n15268), .A2(n15667), .A3(n10307), .ZN(n15666) );
  NAND2_X1 U15659 ( .A1(n15627), .A2(n15628), .ZN(n15667) );
  NOR2_X1 U15660 ( .A1(n15627), .A2(n15628), .ZN(n15664) );
  NOR2_X1 U15661 ( .A1(n15668), .A2(n15669), .ZN(n15628) );
  INV_X1 U15662 ( .A(n15670), .ZN(n15669) );
  NAND3_X1 U15663 ( .A1(n15268), .A2(n15671), .A3(n9286), .ZN(n15670) );
  NAND2_X1 U15664 ( .A1(n15622), .A2(n15624), .ZN(n15671) );
  NOR2_X1 U15665 ( .A1(n15622), .A2(n15624), .ZN(n15668) );
  NOR2_X1 U15666 ( .A1(n15672), .A2(n15673), .ZN(n15624) );
  NOR3_X1 U15667 ( .A1(n8529), .A2(n15674), .A3(n8544), .ZN(n15673) );
  NOR2_X1 U15668 ( .A1(n15619), .A2(n15620), .ZN(n15674) );
  INV_X1 U15669 ( .A(n15675), .ZN(n15672) );
  NAND2_X1 U15670 ( .A1(n15619), .A2(n15620), .ZN(n15675) );
  NAND2_X1 U15671 ( .A1(n15676), .A2(n15677), .ZN(n15620) );
  INV_X1 U15672 ( .A(n15678), .ZN(n15677) );
  NOR3_X1 U15673 ( .A1(n8529), .A2(n15679), .A3(n8560), .ZN(n15678) );
  NOR2_X1 U15674 ( .A1(n15614), .A2(n15616), .ZN(n15679) );
  NAND2_X1 U15675 ( .A1(n15614), .A2(n15616), .ZN(n15676) );
  NAND2_X1 U15676 ( .A1(n15680), .A2(n15681), .ZN(n15616) );
  NAND3_X1 U15677 ( .A1(n15268), .A2(n15682), .A3(n10846), .ZN(n15681) );
  INV_X1 U15678 ( .A(n15683), .ZN(n15682) );
  NOR2_X1 U15679 ( .A1(n15611), .A2(n15612), .ZN(n15683) );
  NAND2_X1 U15680 ( .A1(n15611), .A2(n15612), .ZN(n15680) );
  NAND2_X1 U15681 ( .A1(n15684), .A2(n15685), .ZN(n15612) );
  INV_X1 U15682 ( .A(n15686), .ZN(n15685) );
  NOR3_X1 U15683 ( .A1(n8529), .A2(n15687), .A3(n8556), .ZN(n15686) );
  NOR2_X1 U15684 ( .A1(n15439), .A2(n15441), .ZN(n15687) );
  NAND2_X1 U15685 ( .A1(n15439), .A2(n15441), .ZN(n15684) );
  NAND2_X1 U15686 ( .A1(n15688), .A2(n15689), .ZN(n15441) );
  NAND3_X1 U15687 ( .A1(n15268), .A2(n15690), .A3(n9209), .ZN(n15689) );
  INV_X1 U15688 ( .A(n15691), .ZN(n15690) );
  NOR2_X1 U15689 ( .A1(n15607), .A2(n15608), .ZN(n15691) );
  NAND2_X1 U15690 ( .A1(n15607), .A2(n15608), .ZN(n15688) );
  NAND2_X1 U15691 ( .A1(n15692), .A2(n15693), .ZN(n15608) );
  INV_X1 U15692 ( .A(n15694), .ZN(n15693) );
  NOR3_X1 U15693 ( .A1(n8529), .A2(n15695), .A3(n8582), .ZN(n15694) );
  NOR2_X1 U15694 ( .A1(n15451), .A2(n15453), .ZN(n15695) );
  NAND2_X1 U15695 ( .A1(n15451), .A2(n15453), .ZN(n15692) );
  NAND2_X1 U15696 ( .A1(n15696), .A2(n15697), .ZN(n15453) );
  NAND3_X1 U15697 ( .A1(n15268), .A2(n15698), .A3(n9721), .ZN(n15697) );
  INV_X1 U15698 ( .A(n15699), .ZN(n15698) );
  NOR2_X1 U15699 ( .A1(n15603), .A2(n15604), .ZN(n15699) );
  NAND2_X1 U15700 ( .A1(n15603), .A2(n15604), .ZN(n15696) );
  NAND2_X1 U15701 ( .A1(n15700), .A2(n15701), .ZN(n15604) );
  INV_X1 U15702 ( .A(n15702), .ZN(n15701) );
  NOR3_X1 U15703 ( .A1(n8529), .A2(n15703), .A3(n8562), .ZN(n15702) );
  NOR2_X1 U15704 ( .A1(n15463), .A2(n15465), .ZN(n15703) );
  NAND2_X1 U15705 ( .A1(n15463), .A2(n15465), .ZN(n15700) );
  NAND2_X1 U15706 ( .A1(n15704), .A2(n15705), .ZN(n15465) );
  NAND3_X1 U15707 ( .A1(n15268), .A2(n15706), .A3(n10222), .ZN(n15705) );
  INV_X1 U15708 ( .A(n15707), .ZN(n15706) );
  NOR2_X1 U15709 ( .A1(n15599), .A2(n15600), .ZN(n15707) );
  NAND2_X1 U15710 ( .A1(n15599), .A2(n15600), .ZN(n15704) );
  NAND2_X1 U15711 ( .A1(n15708), .A2(n15709), .ZN(n15600) );
  INV_X1 U15712 ( .A(n15710), .ZN(n15709) );
  NOR3_X1 U15713 ( .A1(n8529), .A2(n15711), .A3(n8569), .ZN(n15710) );
  NOR2_X1 U15714 ( .A1(n15475), .A2(n15477), .ZN(n15711) );
  NAND2_X1 U15715 ( .A1(n15475), .A2(n15477), .ZN(n15708) );
  NAND2_X1 U15716 ( .A1(n15712), .A2(n15713), .ZN(n15477) );
  NAND3_X1 U15717 ( .A1(n15268), .A2(n15714), .A3(n10722), .ZN(n15713) );
  INV_X1 U15718 ( .A(n15715), .ZN(n15714) );
  NOR2_X1 U15719 ( .A1(n15595), .A2(n15596), .ZN(n15715) );
  NAND2_X1 U15720 ( .A1(n15595), .A2(n15596), .ZN(n15712) );
  NAND2_X1 U15721 ( .A1(n15716), .A2(n15717), .ZN(n15596) );
  INV_X1 U15722 ( .A(n15718), .ZN(n15717) );
  NOR3_X1 U15723 ( .A1(n8529), .A2(n15719), .A3(n8583), .ZN(n15718) );
  NOR2_X1 U15724 ( .A1(n15487), .A2(n15489), .ZN(n15719) );
  NAND2_X1 U15725 ( .A1(n15487), .A2(n15489), .ZN(n15716) );
  NAND2_X1 U15726 ( .A1(n15720), .A2(n15721), .ZN(n15489) );
  NAND3_X1 U15727 ( .A1(n9070), .A2(n15722), .A3(n15268), .ZN(n15721) );
  INV_X1 U15728 ( .A(n15723), .ZN(n15722) );
  NOR2_X1 U15729 ( .A1(n15591), .A2(n15592), .ZN(n15723) );
  NAND2_X1 U15730 ( .A1(n15591), .A2(n15592), .ZN(n15720) );
  NAND2_X1 U15731 ( .A1(n15724), .A2(n15725), .ZN(n15592) );
  INV_X1 U15732 ( .A(n15726), .ZN(n15725) );
  NOR3_X1 U15733 ( .A1(n9076), .A2(n15727), .A3(n8529), .ZN(n15726) );
  NOR2_X1 U15734 ( .A1(n15499), .A2(n15501), .ZN(n15727) );
  NAND2_X1 U15735 ( .A1(n15499), .A2(n15501), .ZN(n15724) );
  NAND2_X1 U15736 ( .A1(n15728), .A2(n15729), .ZN(n15501) );
  NAND3_X1 U15737 ( .A1(n8515), .A2(n15730), .A3(n15268), .ZN(n15729) );
  INV_X1 U15738 ( .A(n15731), .ZN(n15730) );
  NOR2_X1 U15739 ( .A1(n15508), .A2(n15509), .ZN(n15731) );
  NAND2_X1 U15740 ( .A1(n15508), .A2(n15509), .ZN(n15728) );
  NAND2_X1 U15741 ( .A1(n15732), .A2(n15733), .ZN(n15509) );
  NAND3_X1 U15742 ( .A1(n9098), .A2(n15734), .A3(n15268), .ZN(n15733) );
  INV_X1 U15743 ( .A(n15735), .ZN(n15734) );
  NOR2_X1 U15744 ( .A1(n15517), .A2(n15515), .ZN(n15735) );
  NAND2_X1 U15745 ( .A1(n15515), .A2(n15517), .ZN(n15732) );
  NAND2_X1 U15746 ( .A1(n15736), .A2(n15737), .ZN(n15517) );
  NAND3_X1 U15747 ( .A1(n9107), .A2(n15738), .A3(n15268), .ZN(n15737) );
  INV_X1 U15748 ( .A(n15739), .ZN(n15738) );
  NOR2_X1 U15749 ( .A1(n15587), .A2(n15588), .ZN(n15739) );
  NAND2_X1 U15750 ( .A1(n15587), .A2(n15588), .ZN(n15736) );
  NAND2_X1 U15751 ( .A1(n15584), .A2(n15740), .ZN(n15588) );
  NAND2_X1 U15752 ( .A1(n15583), .A2(n15585), .ZN(n15740) );
  NAND2_X1 U15753 ( .A1(n15741), .A2(n15742), .ZN(n15585) );
  NAND2_X1 U15754 ( .A1(n15268), .A2(n9112), .ZN(n15742) );
  XNOR2_X1 U15755 ( .A(n15743), .B(n15744), .ZN(n15583) );
  XNOR2_X1 U15756 ( .A(n15745), .B(n15746), .ZN(n15743) );
  INV_X1 U15757 ( .A(n15747), .ZN(n15584) );
  NOR2_X1 U15758 ( .A1(n9176), .A2(n15741), .ZN(n15747) );
  NOR2_X1 U15759 ( .A1(n15748), .A2(n15749), .ZN(n15741) );
  INV_X1 U15760 ( .A(n15750), .ZN(n15749) );
  NAND2_X1 U15761 ( .A1(n15581), .A2(n15751), .ZN(n15750) );
  NAND2_X1 U15762 ( .A1(n15580), .A2(n15578), .ZN(n15751) );
  NOR2_X1 U15763 ( .A1(n8529), .A2(n8535), .ZN(n15581) );
  NOR2_X1 U15764 ( .A1(n15578), .A2(n15580), .ZN(n15748) );
  NOR2_X1 U15765 ( .A1(n15752), .A2(n15753), .ZN(n15580) );
  INV_X1 U15766 ( .A(n15754), .ZN(n15753) );
  NAND2_X1 U15767 ( .A1(n15577), .A2(n15755), .ZN(n15754) );
  NAND2_X1 U15768 ( .A1(n15576), .A2(n15575), .ZN(n15755) );
  NOR2_X1 U15769 ( .A1(n8529), .A2(n9126), .ZN(n15577) );
  NOR2_X1 U15770 ( .A1(n15575), .A2(n15576), .ZN(n15752) );
  NOR2_X1 U15771 ( .A1(n15756), .A2(n15757), .ZN(n15576) );
  INV_X1 U15772 ( .A(n15758), .ZN(n15757) );
  NAND2_X1 U15773 ( .A1(n15572), .A2(n15759), .ZN(n15758) );
  NAND2_X1 U15774 ( .A1(n15571), .A2(n15573), .ZN(n15759) );
  NOR2_X1 U15775 ( .A1(n8529), .A2(n9378), .ZN(n15572) );
  NOR2_X1 U15776 ( .A1(n15571), .A2(n15573), .ZN(n15756) );
  NOR2_X1 U15777 ( .A1(n15760), .A2(n15761), .ZN(n15573) );
  INV_X1 U15778 ( .A(n15762), .ZN(n15761) );
  NAND2_X1 U15779 ( .A1(n15568), .A2(n15763), .ZN(n15762) );
  NAND2_X1 U15780 ( .A1(n15569), .A2(n15567), .ZN(n15763) );
  NOR2_X1 U15781 ( .A1(n8529), .A2(n9383), .ZN(n15568) );
  NOR2_X1 U15782 ( .A1(n15567), .A2(n15569), .ZN(n15760) );
  NOR2_X1 U15783 ( .A1(n15764), .A2(n15765), .ZN(n15569) );
  INV_X1 U15784 ( .A(n15766), .ZN(n15765) );
  NAND2_X1 U15785 ( .A1(n15562), .A2(n15767), .ZN(n15766) );
  NAND2_X1 U15786 ( .A1(n15565), .A2(n15564), .ZN(n15767) );
  NOR2_X1 U15787 ( .A1(n8529), .A2(n9146), .ZN(n15562) );
  NOR2_X1 U15788 ( .A1(n15564), .A2(n15565), .ZN(n15764) );
  INV_X1 U15789 ( .A(n15768), .ZN(n15565) );
  NAND2_X1 U15790 ( .A1(n15769), .A2(n15770), .ZN(n15768) );
  NAND2_X1 U15791 ( .A1(n8532), .A2(n15771), .ZN(n15770) );
  NAND2_X1 U15792 ( .A1(n8624), .A2(n15772), .ZN(n15771) );
  NAND2_X1 U15793 ( .A1(n8579), .A2(n8627), .ZN(n15772) );
  NAND2_X1 U15794 ( .A1(n15774), .A2(n15775), .ZN(n15769) );
  NAND2_X1 U15795 ( .A1(n8630), .A2(n15776), .ZN(n15775) );
  NAND2_X1 U15796 ( .A1(n8539), .A2(n8533), .ZN(n15776) );
  NAND3_X1 U15797 ( .A1(n15268), .A2(n8537), .A3(n8532), .ZN(n15564) );
  XOR2_X1 U15798 ( .A(d_5_), .B(c_5_), .Z(n15778) );
  XOR2_X1 U15799 ( .A(n15779), .B(n15780), .Z(n15567) );
  XNOR2_X1 U15800 ( .A(n15781), .B(n15782), .ZN(n15780) );
  XOR2_X1 U15801 ( .A(n15783), .B(n15784), .Z(n15571) );
  XNOR2_X1 U15802 ( .A(n15785), .B(n15786), .ZN(n15783) );
  XOR2_X1 U15803 ( .A(n15787), .B(n15788), .Z(n15575) );
  XNOR2_X1 U15804 ( .A(n15789), .B(n15790), .ZN(n15787) );
  XOR2_X1 U15805 ( .A(n15791), .B(n15792), .Z(n15578) );
  XNOR2_X1 U15806 ( .A(n15793), .B(n15794), .ZN(n15791) );
  XNOR2_X1 U15807 ( .A(n15795), .B(n15796), .ZN(n15587) );
  XNOR2_X1 U15808 ( .A(n15797), .B(n15798), .ZN(n15795) );
  NOR2_X1 U15809 ( .A1(n9176), .A2(n8533), .ZN(n15798) );
  XNOR2_X1 U15810 ( .A(n15799), .B(n15800), .ZN(n15515) );
  NAND2_X1 U15811 ( .A1(n15801), .A2(n15802), .ZN(n15799) );
  XNOR2_X1 U15812 ( .A(n15803), .B(n15804), .ZN(n15508) );
  XNOR2_X1 U15813 ( .A(n15805), .B(n15806), .ZN(n15803) );
  XNOR2_X1 U15814 ( .A(n15807), .B(n15808), .ZN(n15499) );
  XNOR2_X1 U15815 ( .A(n15809), .B(n15810), .ZN(n15807) );
  XNOR2_X1 U15816 ( .A(n15811), .B(n15812), .ZN(n15591) );
  XNOR2_X1 U15817 ( .A(n15813), .B(n15814), .ZN(n15812) );
  XNOR2_X1 U15818 ( .A(n15815), .B(n15816), .ZN(n15487) );
  XOR2_X1 U15819 ( .A(n15817), .B(n15818), .Z(n15816) );
  XOR2_X1 U15820 ( .A(n15819), .B(n15820), .Z(n15595) );
  XNOR2_X1 U15821 ( .A(n15821), .B(n15822), .ZN(n15820) );
  XNOR2_X1 U15822 ( .A(n15823), .B(n15824), .ZN(n15475) );
  XOR2_X1 U15823 ( .A(n15825), .B(n15826), .Z(n15824) );
  XOR2_X1 U15824 ( .A(n15827), .B(n15828), .Z(n15599) );
  XNOR2_X1 U15825 ( .A(n15829), .B(n15830), .ZN(n15828) );
  XNOR2_X1 U15826 ( .A(n15831), .B(n15832), .ZN(n15463) );
  XOR2_X1 U15827 ( .A(n15833), .B(n15834), .Z(n15832) );
  XOR2_X1 U15828 ( .A(n15835), .B(n15836), .Z(n15603) );
  XNOR2_X1 U15829 ( .A(n15837), .B(n15838), .ZN(n15836) );
  XNOR2_X1 U15830 ( .A(n15839), .B(n15840), .ZN(n15451) );
  XOR2_X1 U15831 ( .A(n15841), .B(n15842), .Z(n15840) );
  XOR2_X1 U15832 ( .A(n15843), .B(n15844), .Z(n15607) );
  XNOR2_X1 U15833 ( .A(n15845), .B(n15846), .ZN(n15844) );
  XNOR2_X1 U15834 ( .A(n15847), .B(n15848), .ZN(n15439) );
  XOR2_X1 U15835 ( .A(n15849), .B(n15850), .Z(n15848) );
  XOR2_X1 U15836 ( .A(n15851), .B(n15852), .Z(n15611) );
  XOR2_X1 U15837 ( .A(n15853), .B(n15854), .Z(n15852) );
  XOR2_X1 U15838 ( .A(n15855), .B(n15856), .Z(n15614) );
  XOR2_X1 U15839 ( .A(n15857), .B(n15858), .Z(n15856) );
  XOR2_X1 U15840 ( .A(n15859), .B(n15860), .Z(n15619) );
  XOR2_X1 U15841 ( .A(n15861), .B(n15862), .Z(n15860) );
  XNOR2_X1 U15842 ( .A(n15863), .B(n15864), .ZN(n15622) );
  XOR2_X1 U15843 ( .A(n15865), .B(n15866), .Z(n15864) );
  XNOR2_X1 U15844 ( .A(n15867), .B(n15868), .ZN(n15627) );
  XOR2_X1 U15845 ( .A(n15869), .B(n15870), .Z(n15868) );
  XNOR2_X1 U15846 ( .A(n15871), .B(n15872), .ZN(n15630) );
  XOR2_X1 U15847 ( .A(n15873), .B(n15874), .Z(n15872) );
  XNOR2_X1 U15848 ( .A(n15875), .B(n15876), .ZN(n15634) );
  XOR2_X1 U15849 ( .A(n15877), .B(n15878), .Z(n15876) );
  XNOR2_X1 U15850 ( .A(n15879), .B(n15880), .ZN(n15638) );
  XOR2_X1 U15851 ( .A(n15881), .B(n15882), .Z(n15880) );
  XNOR2_X1 U15852 ( .A(n15883), .B(n15884), .ZN(n15642) );
  XOR2_X1 U15853 ( .A(n15885), .B(n15886), .Z(n15884) );
  XNOR2_X1 U15854 ( .A(n15887), .B(n15888), .ZN(n15393) );
  XOR2_X1 U15855 ( .A(n15889), .B(n15890), .Z(n15888) );
  XOR2_X1 U15856 ( .A(n8740), .B(n8739), .Z(n8690) );
  NOR3_X1 U15857 ( .A1(n8740), .A2(n8739), .A3(n8738), .ZN(n8734) );
  NAND2_X1 U15858 ( .A1(n15891), .A2(n8888), .ZN(n8738) );
  INV_X1 U15859 ( .A(n15892), .ZN(n8888) );
  NOR2_X1 U15860 ( .A1(n15893), .A2(n15894), .ZN(n15892) );
  NAND2_X1 U15861 ( .A1(n15894), .A2(n15893), .ZN(n15891) );
  XOR2_X1 U15862 ( .A(n15895), .B(n15896), .Z(n15893) );
  NAND2_X1 U15863 ( .A1(n15897), .A2(n15898), .ZN(n15895) );
  NOR2_X1 U15864 ( .A1(n15899), .A2(n15900), .ZN(n15894) );
  INV_X1 U15865 ( .A(n15901), .ZN(n15900) );
  NAND3_X1 U15866 ( .A1(n8592), .A2(n15902), .A3(n15774), .ZN(n15901) );
  NAND2_X1 U15867 ( .A1(n15903), .A2(n15904), .ZN(n15902) );
  NOR2_X1 U15868 ( .A1(n15903), .A2(n15904), .ZN(n15899) );
  NOR2_X1 U15869 ( .A1(n15905), .A2(n15906), .ZN(n8739) );
  INV_X1 U15870 ( .A(n15907), .ZN(n15906) );
  NAND2_X1 U15871 ( .A1(n15398), .A2(n15908), .ZN(n15907) );
  NAND2_X1 U15872 ( .A1(n15397), .A2(n15396), .ZN(n15908) );
  NOR2_X1 U15873 ( .A1(n8533), .A2(n8972), .ZN(n15398) );
  NOR2_X1 U15874 ( .A1(n15396), .A2(n15397), .ZN(n15905) );
  NOR2_X1 U15875 ( .A1(n15909), .A2(n15910), .ZN(n15397) );
  INV_X1 U15876 ( .A(n15911), .ZN(n15910) );
  NAND2_X1 U15877 ( .A1(n15890), .A2(n15912), .ZN(n15911) );
  NAND2_X1 U15878 ( .A1(n15889), .A2(n15887), .ZN(n15912) );
  NOR2_X1 U15879 ( .A1(n8884), .A2(n8533), .ZN(n15890) );
  NOR2_X1 U15880 ( .A1(n15887), .A2(n15889), .ZN(n15909) );
  NOR2_X1 U15881 ( .A1(n15913), .A2(n15914), .ZN(n15889) );
  INV_X1 U15882 ( .A(n15915), .ZN(n15914) );
  NAND2_X1 U15883 ( .A1(n15886), .A2(n15916), .ZN(n15915) );
  NAND2_X1 U15884 ( .A1(n15885), .A2(n15883), .ZN(n15916) );
  NOR2_X1 U15885 ( .A1(n8982), .A2(n8533), .ZN(n15886) );
  NOR2_X1 U15886 ( .A1(n15883), .A2(n15885), .ZN(n15913) );
  NOR2_X1 U15887 ( .A1(n15917), .A2(n15918), .ZN(n15885) );
  INV_X1 U15888 ( .A(n15919), .ZN(n15918) );
  NAND2_X1 U15889 ( .A1(n15882), .A2(n15920), .ZN(n15919) );
  NAND2_X1 U15890 ( .A1(n15881), .A2(n15879), .ZN(n15920) );
  NOR2_X1 U15891 ( .A1(n8527), .A2(n8533), .ZN(n15882) );
  NOR2_X1 U15892 ( .A1(n15879), .A2(n15881), .ZN(n15917) );
  NOR2_X1 U15893 ( .A1(n15921), .A2(n15922), .ZN(n15881) );
  INV_X1 U15894 ( .A(n15923), .ZN(n15922) );
  NAND2_X1 U15895 ( .A1(n15878), .A2(n15924), .ZN(n15923) );
  NAND2_X1 U15896 ( .A1(n15877), .A2(n15875), .ZN(n15924) );
  NOR2_X1 U15897 ( .A1(n8528), .A2(n8533), .ZN(n15878) );
  NOR2_X1 U15898 ( .A1(n15875), .A2(n15877), .ZN(n15921) );
  NOR2_X1 U15899 ( .A1(n15925), .A2(n15926), .ZN(n15877) );
  INV_X1 U15900 ( .A(n15927), .ZN(n15926) );
  NAND2_X1 U15901 ( .A1(n15874), .A2(n15928), .ZN(n15927) );
  NAND2_X1 U15902 ( .A1(n15873), .A2(n15871), .ZN(n15928) );
  NOR2_X1 U15903 ( .A1(n8995), .A2(n8533), .ZN(n15874) );
  NOR2_X1 U15904 ( .A1(n15871), .A2(n15873), .ZN(n15925) );
  NOR2_X1 U15905 ( .A1(n15929), .A2(n15930), .ZN(n15873) );
  INV_X1 U15906 ( .A(n15931), .ZN(n15930) );
  NAND2_X1 U15907 ( .A1(n15870), .A2(n15932), .ZN(n15931) );
  NAND2_X1 U15908 ( .A1(n15869), .A2(n15867), .ZN(n15932) );
  NOR2_X1 U15909 ( .A1(n8555), .A2(n8533), .ZN(n15870) );
  NOR2_X1 U15910 ( .A1(n15867), .A2(n15869), .ZN(n15929) );
  NOR2_X1 U15911 ( .A1(n15933), .A2(n15934), .ZN(n15869) );
  INV_X1 U15912 ( .A(n15935), .ZN(n15934) );
  NAND2_X1 U15913 ( .A1(n15866), .A2(n15936), .ZN(n15935) );
  NAND2_X1 U15914 ( .A1(n15865), .A2(n15863), .ZN(n15936) );
  NOR2_X1 U15915 ( .A1(n8544), .A2(n8533), .ZN(n15866) );
  NOR2_X1 U15916 ( .A1(n15863), .A2(n15865), .ZN(n15933) );
  NOR2_X1 U15917 ( .A1(n15937), .A2(n15938), .ZN(n15865) );
  INV_X1 U15918 ( .A(n15939), .ZN(n15938) );
  NAND2_X1 U15919 ( .A1(n15862), .A2(n15940), .ZN(n15939) );
  NAND2_X1 U15920 ( .A1(n15861), .A2(n15859), .ZN(n15940) );
  NOR2_X1 U15921 ( .A1(n9010), .A2(n8533), .ZN(n15862) );
  NOR2_X1 U15922 ( .A1(n15859), .A2(n15861), .ZN(n15937) );
  NOR2_X1 U15923 ( .A1(n15941), .A2(n15942), .ZN(n15861) );
  INV_X1 U15924 ( .A(n15943), .ZN(n15942) );
  NAND2_X1 U15925 ( .A1(n15858), .A2(n15944), .ZN(n15943) );
  NAND2_X1 U15926 ( .A1(n15857), .A2(n15855), .ZN(n15944) );
  NOR2_X1 U15927 ( .A1(n8594), .A2(n8533), .ZN(n15858) );
  NOR2_X1 U15928 ( .A1(n15855), .A2(n15857), .ZN(n15941) );
  NOR2_X1 U15929 ( .A1(n15945), .A2(n15946), .ZN(n15857) );
  INV_X1 U15930 ( .A(n15947), .ZN(n15946) );
  NAND2_X1 U15931 ( .A1(n15854), .A2(n15948), .ZN(n15947) );
  NAND2_X1 U15932 ( .A1(n15853), .A2(n15851), .ZN(n15948) );
  NOR2_X1 U15933 ( .A1(n9020), .A2(n8533), .ZN(n15854) );
  NOR2_X1 U15934 ( .A1(n15851), .A2(n15853), .ZN(n15945) );
  NOR2_X1 U15935 ( .A1(n15949), .A2(n15950), .ZN(n15853) );
  NOR2_X1 U15936 ( .A1(n15850), .A2(n15951), .ZN(n15950) );
  NOR2_X1 U15937 ( .A1(n15849), .A2(n15847), .ZN(n15951) );
  NAND2_X1 U15938 ( .A1(n9209), .A2(n8532), .ZN(n15850) );
  INV_X1 U15939 ( .A(n15952), .ZN(n15949) );
  NAND2_X1 U15940 ( .A1(n15847), .A2(n15849), .ZN(n15952) );
  NAND2_X1 U15941 ( .A1(n15953), .A2(n15954), .ZN(n15849) );
  NAND2_X1 U15942 ( .A1(n15846), .A2(n15955), .ZN(n15954) );
  NAND2_X1 U15943 ( .A1(n15956), .A2(n15843), .ZN(n15955) );
  INV_X1 U15944 ( .A(n15845), .ZN(n15956) );
  NOR2_X1 U15945 ( .A1(n9031), .A2(n8533), .ZN(n15846) );
  NAND2_X1 U15946 ( .A1(n15957), .A2(n15845), .ZN(n15953) );
  NAND2_X1 U15947 ( .A1(n15958), .A2(n15959), .ZN(n15845) );
  INV_X1 U15948 ( .A(n15960), .ZN(n15959) );
  NOR2_X1 U15949 ( .A1(n15842), .A2(n15961), .ZN(n15960) );
  NOR2_X1 U15950 ( .A1(n15841), .A2(n15839), .ZN(n15961) );
  NAND2_X1 U15951 ( .A1(n9721), .A2(n8532), .ZN(n15842) );
  NAND2_X1 U15952 ( .A1(n15839), .A2(n15841), .ZN(n15958) );
  NAND2_X1 U15953 ( .A1(n15962), .A2(n15963), .ZN(n15841) );
  NAND2_X1 U15954 ( .A1(n15838), .A2(n15964), .ZN(n15963) );
  NAND2_X1 U15955 ( .A1(n15965), .A2(n15835), .ZN(n15964) );
  INV_X1 U15956 ( .A(n15837), .ZN(n15965) );
  NOR2_X1 U15957 ( .A1(n9041), .A2(n8533), .ZN(n15838) );
  NAND2_X1 U15958 ( .A1(n15966), .A2(n15837), .ZN(n15962) );
  NAND2_X1 U15959 ( .A1(n15967), .A2(n15968), .ZN(n15837) );
  INV_X1 U15960 ( .A(n15969), .ZN(n15968) );
  NOR2_X1 U15961 ( .A1(n15834), .A2(n15970), .ZN(n15969) );
  NOR2_X1 U15962 ( .A1(n15833), .A2(n15831), .ZN(n15970) );
  NAND2_X1 U15963 ( .A1(n10222), .A2(n8532), .ZN(n15834) );
  NAND2_X1 U15964 ( .A1(n15831), .A2(n15833), .ZN(n15967) );
  NAND2_X1 U15965 ( .A1(n15971), .A2(n15972), .ZN(n15833) );
  NAND2_X1 U15966 ( .A1(n15830), .A2(n15973), .ZN(n15972) );
  NAND2_X1 U15967 ( .A1(n15974), .A2(n15827), .ZN(n15973) );
  INV_X1 U15968 ( .A(n15829), .ZN(n15974) );
  NOR2_X1 U15969 ( .A1(n9050), .A2(n8533), .ZN(n15830) );
  NAND2_X1 U15970 ( .A1(n15975), .A2(n15829), .ZN(n15971) );
  NAND2_X1 U15971 ( .A1(n15976), .A2(n15977), .ZN(n15829) );
  INV_X1 U15972 ( .A(n15978), .ZN(n15977) );
  NOR2_X1 U15973 ( .A1(n15826), .A2(n15979), .ZN(n15978) );
  NOR2_X1 U15974 ( .A1(n15825), .A2(n15823), .ZN(n15979) );
  NAND2_X1 U15975 ( .A1(n10722), .A2(n8532), .ZN(n15826) );
  NAND2_X1 U15976 ( .A1(n15823), .A2(n15825), .ZN(n15976) );
  NAND2_X1 U15977 ( .A1(n15980), .A2(n15981), .ZN(n15825) );
  NAND2_X1 U15978 ( .A1(n15822), .A2(n15982), .ZN(n15981) );
  NAND2_X1 U15979 ( .A1(n15983), .A2(n15819), .ZN(n15982) );
  INV_X1 U15980 ( .A(n15821), .ZN(n15983) );
  NOR2_X1 U15981 ( .A1(n9061), .A2(n8533), .ZN(n15822) );
  NAND2_X1 U15982 ( .A1(n15984), .A2(n15821), .ZN(n15980) );
  NAND2_X1 U15983 ( .A1(n15985), .A2(n15986), .ZN(n15821) );
  INV_X1 U15984 ( .A(n15987), .ZN(n15986) );
  NOR2_X1 U15985 ( .A1(n15818), .A2(n15988), .ZN(n15987) );
  NOR2_X1 U15986 ( .A1(n15817), .A2(n15815), .ZN(n15988) );
  NAND2_X1 U15987 ( .A1(n8532), .A2(n9070), .ZN(n15818) );
  NAND2_X1 U15988 ( .A1(n15815), .A2(n15817), .ZN(n15985) );
  NAND2_X1 U15989 ( .A1(n15989), .A2(n15990), .ZN(n15817) );
  NAND2_X1 U15990 ( .A1(n15814), .A2(n15991), .ZN(n15990) );
  INV_X1 U15991 ( .A(n15992), .ZN(n15991) );
  NOR2_X1 U15992 ( .A1(n15813), .A2(n15811), .ZN(n15992) );
  NOR2_X1 U15993 ( .A1(n8533), .A2(n8588), .ZN(n15814) );
  NAND2_X1 U15994 ( .A1(n15811), .A2(n15813), .ZN(n15989) );
  NAND2_X1 U15995 ( .A1(n15993), .A2(n15994), .ZN(n15813) );
  NAND2_X1 U15996 ( .A1(n15810), .A2(n15995), .ZN(n15994) );
  NAND2_X1 U15997 ( .A1(n15809), .A2(n15808), .ZN(n15995) );
  NOR2_X1 U15998 ( .A1(n8533), .A2(n8551), .ZN(n15810) );
  INV_X1 U15999 ( .A(n15996), .ZN(n15993) );
  NOR2_X1 U16000 ( .A1(n15808), .A2(n15809), .ZN(n15996) );
  NOR2_X1 U16001 ( .A1(n15997), .A2(n15998), .ZN(n15809) );
  INV_X1 U16002 ( .A(n15999), .ZN(n15998) );
  NAND2_X1 U16003 ( .A1(n15806), .A2(n16000), .ZN(n15999) );
  NAND2_X1 U16004 ( .A1(n15805), .A2(n15804), .ZN(n16000) );
  NOR2_X1 U16005 ( .A1(n8533), .A2(n8563), .ZN(n15806) );
  NOR2_X1 U16006 ( .A1(n15804), .A2(n15805), .ZN(n15997) );
  INV_X1 U16007 ( .A(n16001), .ZN(n15805) );
  NAND2_X1 U16008 ( .A1(n15801), .A2(n16002), .ZN(n16001) );
  NAND2_X1 U16009 ( .A1(n15800), .A2(n15802), .ZN(n16002) );
  NAND2_X1 U16010 ( .A1(n16003), .A2(n16004), .ZN(n15802) );
  NAND2_X1 U16011 ( .A1(n8532), .A2(n9107), .ZN(n16004) );
  XNOR2_X1 U16012 ( .A(n16005), .B(n16006), .ZN(n15800) );
  XNOR2_X1 U16013 ( .A(n16007), .B(n16008), .ZN(n16005) );
  NOR2_X1 U16014 ( .A1(n9176), .A2(n8579), .ZN(n16008) );
  INV_X1 U16015 ( .A(n16009), .ZN(n15801) );
  NOR2_X1 U16016 ( .A1(n8548), .A2(n16003), .ZN(n16009) );
  NOR2_X1 U16017 ( .A1(n16010), .A2(n16011), .ZN(n16003) );
  INV_X1 U16018 ( .A(n16012), .ZN(n16011) );
  NAND3_X1 U16019 ( .A1(n9112), .A2(n16013), .A3(n8532), .ZN(n16012) );
  NAND2_X1 U16020 ( .A1(n15797), .A2(n15796), .ZN(n16013) );
  INV_X1 U16021 ( .A(n9176), .ZN(n9112) );
  NOR2_X1 U16022 ( .A1(n15796), .A2(n15797), .ZN(n16010) );
  NOR2_X1 U16023 ( .A1(n16014), .A2(n16015), .ZN(n15797) );
  INV_X1 U16024 ( .A(n16016), .ZN(n16015) );
  NAND2_X1 U16025 ( .A1(n15746), .A2(n16017), .ZN(n16016) );
  NAND2_X1 U16026 ( .A1(n15745), .A2(n15744), .ZN(n16017) );
  NOR2_X1 U16027 ( .A1(n8533), .A2(n8535), .ZN(n15746) );
  NOR2_X1 U16028 ( .A1(n15744), .A2(n15745), .ZN(n16014) );
  NOR2_X1 U16029 ( .A1(n16018), .A2(n16019), .ZN(n15745) );
  INV_X1 U16030 ( .A(n16020), .ZN(n16019) );
  NAND2_X1 U16031 ( .A1(n15794), .A2(n16021), .ZN(n16020) );
  NAND2_X1 U16032 ( .A1(n15792), .A2(n15793), .ZN(n16021) );
  NOR2_X1 U16033 ( .A1(n8533), .A2(n9126), .ZN(n15794) );
  NOR2_X1 U16034 ( .A1(n15792), .A2(n15793), .ZN(n16018) );
  NOR2_X1 U16035 ( .A1(n16022), .A2(n16023), .ZN(n15793) );
  INV_X1 U16036 ( .A(n16024), .ZN(n16023) );
  NAND2_X1 U16037 ( .A1(n15789), .A2(n16025), .ZN(n16024) );
  NAND2_X1 U16038 ( .A1(n15788), .A2(n15790), .ZN(n16025) );
  NOR2_X1 U16039 ( .A1(n8533), .A2(n9378), .ZN(n15789) );
  NOR2_X1 U16040 ( .A1(n15788), .A2(n15790), .ZN(n16022) );
  NOR2_X1 U16041 ( .A1(n16026), .A2(n16027), .ZN(n15790) );
  INV_X1 U16042 ( .A(n16028), .ZN(n16027) );
  NAND2_X1 U16043 ( .A1(n15785), .A2(n16029), .ZN(n16028) );
  NAND2_X1 U16044 ( .A1(n15786), .A2(n15784), .ZN(n16029) );
  NOR2_X1 U16045 ( .A1(n8533), .A2(n9383), .ZN(n15785) );
  NOR2_X1 U16046 ( .A1(n15784), .A2(n15786), .ZN(n16026) );
  NOR2_X1 U16047 ( .A1(n16030), .A2(n16031), .ZN(n15786) );
  INV_X1 U16048 ( .A(n16032), .ZN(n16031) );
  NAND2_X1 U16049 ( .A1(n15779), .A2(n16033), .ZN(n16032) );
  NAND2_X1 U16050 ( .A1(n15782), .A2(n15781), .ZN(n16033) );
  NOR2_X1 U16051 ( .A1(n8533), .A2(n9146), .ZN(n15779) );
  NOR2_X1 U16052 ( .A1(n15781), .A2(n15782), .ZN(n16030) );
  INV_X1 U16053 ( .A(n16034), .ZN(n15782) );
  NAND2_X1 U16054 ( .A1(n16035), .A2(n16036), .ZN(n16034) );
  NAND2_X1 U16055 ( .A1(n15774), .A2(n16037), .ZN(n16036) );
  NAND2_X1 U16056 ( .A1(n8624), .A2(n16038), .ZN(n16037) );
  NAND2_X1 U16057 ( .A1(n8577), .A2(n8627), .ZN(n16038) );
  NAND2_X1 U16058 ( .A1(n16040), .A2(n16041), .ZN(n16035) );
  NAND2_X1 U16059 ( .A1(n8630), .A2(n16042), .ZN(n16041) );
  NAND2_X1 U16060 ( .A1(n8539), .A2(n8579), .ZN(n16042) );
  NAND3_X1 U16061 ( .A1(n8532), .A2(n8537), .A3(n15774), .ZN(n15781) );
  XNOR2_X1 U16062 ( .A(n16043), .B(n16044), .ZN(n15557) );
  XOR2_X1 U16063 ( .A(d_4_), .B(c_4_), .Z(n16044) );
  XOR2_X1 U16064 ( .A(n16045), .B(n16046), .Z(n15784) );
  XNOR2_X1 U16065 ( .A(n16047), .B(n16048), .ZN(n16046) );
  XOR2_X1 U16066 ( .A(n16049), .B(n16050), .Z(n15788) );
  XNOR2_X1 U16067 ( .A(n16051), .B(n16052), .ZN(n16049) );
  XOR2_X1 U16068 ( .A(n16053), .B(n16054), .Z(n15792) );
  XNOR2_X1 U16069 ( .A(n16055), .B(n16056), .ZN(n16053) );
  XOR2_X1 U16070 ( .A(n16057), .B(n16058), .Z(n15744) );
  XNOR2_X1 U16071 ( .A(n16059), .B(n16060), .ZN(n16057) );
  NOR2_X1 U16072 ( .A1(n9126), .A2(n8579), .ZN(n16060) );
  XOR2_X1 U16073 ( .A(n16061), .B(n16062), .Z(n15796) );
  XNOR2_X1 U16074 ( .A(n16063), .B(n16064), .ZN(n16061) );
  NOR2_X1 U16075 ( .A1(n8535), .A2(n8579), .ZN(n16064) );
  XNOR2_X1 U16076 ( .A(n16065), .B(n16066), .ZN(n15804) );
  XNOR2_X1 U16077 ( .A(n16067), .B(n16068), .ZN(n16066) );
  NAND2_X1 U16078 ( .A1(n15774), .A2(n9107), .ZN(n16068) );
  XNOR2_X1 U16079 ( .A(n16069), .B(n16070), .ZN(n15808) );
  XOR2_X1 U16080 ( .A(n16071), .B(n16072), .Z(n16069) );
  NOR2_X1 U16081 ( .A1(n9094), .A2(n8579), .ZN(n16072) );
  XNOR2_X1 U16082 ( .A(n16073), .B(n16074), .ZN(n15811) );
  XOR2_X1 U16083 ( .A(n16075), .B(n16076), .Z(n16074) );
  NAND2_X1 U16084 ( .A1(n15774), .A2(n8515), .ZN(n16076) );
  XOR2_X1 U16085 ( .A(n16077), .B(n16078), .Z(n15815) );
  XOR2_X1 U16086 ( .A(n16079), .B(n16080), .Z(n16077) );
  NOR2_X1 U16087 ( .A1(n9076), .A2(n8579), .ZN(n16080) );
  INV_X1 U16088 ( .A(n15819), .ZN(n15984) );
  XOR2_X1 U16089 ( .A(n16081), .B(n16082), .Z(n15819) );
  XOR2_X1 U16090 ( .A(n16083), .B(n16084), .Z(n16082) );
  NAND2_X1 U16091 ( .A1(n15774), .A2(n9070), .ZN(n16084) );
  XOR2_X1 U16092 ( .A(n16085), .B(n16086), .Z(n15823) );
  XOR2_X1 U16093 ( .A(n16087), .B(n16088), .Z(n16085) );
  NOR2_X1 U16094 ( .A1(n8579), .A2(n8583), .ZN(n16088) );
  INV_X1 U16095 ( .A(n15827), .ZN(n15975) );
  XOR2_X1 U16096 ( .A(n16089), .B(n16090), .Z(n15827) );
  XOR2_X1 U16097 ( .A(n16091), .B(n16092), .Z(n16090) );
  NAND2_X1 U16098 ( .A1(n10722), .A2(n15774), .ZN(n16092) );
  XOR2_X1 U16099 ( .A(n16093), .B(n16094), .Z(n15831) );
  XOR2_X1 U16100 ( .A(n16095), .B(n16096), .Z(n16093) );
  NOR2_X1 U16101 ( .A1(n8579), .A2(n8569), .ZN(n16096) );
  INV_X1 U16102 ( .A(n15835), .ZN(n15966) );
  XOR2_X1 U16103 ( .A(n16097), .B(n16098), .Z(n15835) );
  XOR2_X1 U16104 ( .A(n16099), .B(n16100), .Z(n16098) );
  NAND2_X1 U16105 ( .A1(n10222), .A2(n15774), .ZN(n16100) );
  XOR2_X1 U16106 ( .A(n16101), .B(n16102), .Z(n15839) );
  XOR2_X1 U16107 ( .A(n16103), .B(n16104), .Z(n16101) );
  NOR2_X1 U16108 ( .A1(n8579), .A2(n8562), .ZN(n16104) );
  INV_X1 U16109 ( .A(n15843), .ZN(n15957) );
  XOR2_X1 U16110 ( .A(n16105), .B(n16106), .Z(n15843) );
  XOR2_X1 U16111 ( .A(n16107), .B(n16108), .Z(n16106) );
  NAND2_X1 U16112 ( .A1(n9721), .A2(n15774), .ZN(n16108) );
  XOR2_X1 U16113 ( .A(n16109), .B(n16110), .Z(n15847) );
  XOR2_X1 U16114 ( .A(n16111), .B(n16112), .Z(n16109) );
  NOR2_X1 U16115 ( .A1(n8579), .A2(n8582), .ZN(n16112) );
  XNOR2_X1 U16116 ( .A(n16113), .B(n16114), .ZN(n15851) );
  XOR2_X1 U16117 ( .A(n16115), .B(n16116), .Z(n16113) );
  NOR2_X1 U16118 ( .A1(n8579), .A2(n8572), .ZN(n16116) );
  XOR2_X1 U16119 ( .A(n16117), .B(n16118), .Z(n15855) );
  XNOR2_X1 U16120 ( .A(n16119), .B(n16120), .ZN(n16117) );
  NOR2_X1 U16121 ( .A1(n8579), .A2(n8556), .ZN(n16120) );
  XOR2_X1 U16122 ( .A(n16121), .B(n16122), .Z(n15859) );
  XNOR2_X1 U16123 ( .A(n16123), .B(n16124), .ZN(n16121) );
  NOR2_X1 U16124 ( .A1(n8579), .A2(n8594), .ZN(n16124) );
  XOR2_X1 U16125 ( .A(n16125), .B(n16126), .Z(n15863) );
  XNOR2_X1 U16126 ( .A(n16127), .B(n16128), .ZN(n16125) );
  NOR2_X1 U16127 ( .A1(n8579), .A2(n8560), .ZN(n16128) );
  XOR2_X1 U16128 ( .A(n16129), .B(n16130), .Z(n15867) );
  XNOR2_X1 U16129 ( .A(n16131), .B(n16132), .ZN(n16129) );
  NOR2_X1 U16130 ( .A1(n8579), .A2(n8544), .ZN(n16132) );
  XOR2_X1 U16131 ( .A(n16133), .B(n16134), .Z(n15871) );
  XNOR2_X1 U16132 ( .A(n16135), .B(n16136), .ZN(n16133) );
  NOR2_X1 U16133 ( .A1(n8579), .A2(n8555), .ZN(n16136) );
  XOR2_X1 U16134 ( .A(n16137), .B(n16138), .Z(n15875) );
  XNOR2_X1 U16135 ( .A(n16139), .B(n16140), .ZN(n16137) );
  NOR2_X1 U16136 ( .A1(n8579), .A2(n8564), .ZN(n16140) );
  XOR2_X1 U16137 ( .A(n16141), .B(n16142), .Z(n15879) );
  XNOR2_X1 U16138 ( .A(n16143), .B(n16144), .ZN(n16141) );
  NOR2_X1 U16139 ( .A1(n8579), .A2(n8528), .ZN(n16144) );
  XOR2_X1 U16140 ( .A(n16145), .B(n16146), .Z(n15883) );
  XNOR2_X1 U16141 ( .A(n16147), .B(n16148), .ZN(n16145) );
  NOR2_X1 U16142 ( .A1(n8579), .A2(n8527), .ZN(n16148) );
  XOR2_X1 U16143 ( .A(n16149), .B(n16150), .Z(n15887) );
  XNOR2_X1 U16144 ( .A(n16151), .B(n16152), .ZN(n16149) );
  NOR2_X1 U16145 ( .A1(n8579), .A2(n8552), .ZN(n16152) );
  XNOR2_X1 U16146 ( .A(n16153), .B(n16154), .ZN(n15396) );
  XNOR2_X1 U16147 ( .A(n16155), .B(n16156), .ZN(n16154) );
  NAND2_X1 U16148 ( .A1(n9263), .A2(n15774), .ZN(n16156) );
  XOR2_X1 U16149 ( .A(n16157), .B(n15903), .Z(n8740) );
  XOR2_X1 U16150 ( .A(n16158), .B(n16159), .Z(n15903) );
  XNOR2_X1 U16151 ( .A(n16160), .B(n16161), .ZN(n16158) );
  NOR2_X1 U16152 ( .A1(n8577), .A2(n8589), .ZN(n16161) );
  XNOR2_X1 U16153 ( .A(n15904), .B(n16162), .ZN(n16157) );
  NOR2_X1 U16154 ( .A1(n8972), .A2(n8579), .ZN(n16162) );
  NOR2_X1 U16155 ( .A1(n16163), .A2(n16164), .ZN(n15904) );
  INV_X1 U16156 ( .A(n16165), .ZN(n16164) );
  NAND3_X1 U16157 ( .A1(n15774), .A2(n16166), .A3(n9263), .ZN(n16165) );
  INV_X1 U16158 ( .A(n8884), .ZN(n9263) );
  NAND2_X1 U16159 ( .A1(n16153), .A2(n16155), .ZN(n16166) );
  NOR2_X1 U16160 ( .A1(n16153), .A2(n16155), .ZN(n16163) );
  NOR2_X1 U16161 ( .A1(n16167), .A2(n16168), .ZN(n16155) );
  INV_X1 U16162 ( .A(n16169), .ZN(n16168) );
  NAND3_X1 U16163 ( .A1(n15774), .A2(n16170), .A3(n9268), .ZN(n16169) );
  NAND2_X1 U16164 ( .A1(n16150), .A2(n16151), .ZN(n16170) );
  NOR2_X1 U16165 ( .A1(n16150), .A2(n16151), .ZN(n16167) );
  NOR2_X1 U16166 ( .A1(n16171), .A2(n16172), .ZN(n16151) );
  INV_X1 U16167 ( .A(n16173), .ZN(n16172) );
  NAND3_X1 U16168 ( .A1(n15774), .A2(n16174), .A3(n9792), .ZN(n16173) );
  NAND2_X1 U16169 ( .A1(n16146), .A2(n16147), .ZN(n16174) );
  NOR2_X1 U16170 ( .A1(n16146), .A2(n16147), .ZN(n16171) );
  NOR2_X1 U16171 ( .A1(n16175), .A2(n16176), .ZN(n16147) );
  INV_X1 U16172 ( .A(n16177), .ZN(n16176) );
  NAND3_X1 U16173 ( .A1(n15774), .A2(n16178), .A3(n9277), .ZN(n16177) );
  NAND2_X1 U16174 ( .A1(n16142), .A2(n16143), .ZN(n16178) );
  NOR2_X1 U16175 ( .A1(n16142), .A2(n16143), .ZN(n16175) );
  NOR2_X1 U16176 ( .A1(n16179), .A2(n16180), .ZN(n16143) );
  INV_X1 U16177 ( .A(n16181), .ZN(n16180) );
  NAND3_X1 U16178 ( .A1(n15774), .A2(n16182), .A3(n10307), .ZN(n16181) );
  NAND2_X1 U16179 ( .A1(n16138), .A2(n16139), .ZN(n16182) );
  NOR2_X1 U16180 ( .A1(n16138), .A2(n16139), .ZN(n16179) );
  NOR2_X1 U16181 ( .A1(n16183), .A2(n16184), .ZN(n16139) );
  INV_X1 U16182 ( .A(n16185), .ZN(n16184) );
  NAND3_X1 U16183 ( .A1(n15774), .A2(n16186), .A3(n9286), .ZN(n16185) );
  NAND2_X1 U16184 ( .A1(n16134), .A2(n16135), .ZN(n16186) );
  NOR2_X1 U16185 ( .A1(n16134), .A2(n16135), .ZN(n16183) );
  NOR2_X1 U16186 ( .A1(n16187), .A2(n16188), .ZN(n16135) );
  INV_X1 U16187 ( .A(n16189), .ZN(n16188) );
  NAND3_X1 U16188 ( .A1(n15774), .A2(n16190), .A3(n8543), .ZN(n16189) );
  NAND2_X1 U16189 ( .A1(n16130), .A2(n16131), .ZN(n16190) );
  NOR2_X1 U16190 ( .A1(n16130), .A2(n16131), .ZN(n16187) );
  NOR2_X1 U16191 ( .A1(n16191), .A2(n16192), .ZN(n16131) );
  INV_X1 U16192 ( .A(n16193), .ZN(n16192) );
  NAND3_X1 U16193 ( .A1(n15774), .A2(n16194), .A3(n9295), .ZN(n16193) );
  NAND2_X1 U16194 ( .A1(n16126), .A2(n16127), .ZN(n16194) );
  NOR2_X1 U16195 ( .A1(n16126), .A2(n16127), .ZN(n16191) );
  NOR2_X1 U16196 ( .A1(n16195), .A2(n16196), .ZN(n16127) );
  INV_X1 U16197 ( .A(n16197), .ZN(n16196) );
  NAND3_X1 U16198 ( .A1(n15774), .A2(n16198), .A3(n10846), .ZN(n16197) );
  NAND2_X1 U16199 ( .A1(n16122), .A2(n16123), .ZN(n16198) );
  NOR2_X1 U16200 ( .A1(n16122), .A2(n16123), .ZN(n16195) );
  NOR2_X1 U16201 ( .A1(n16199), .A2(n16200), .ZN(n16123) );
  INV_X1 U16202 ( .A(n16201), .ZN(n16200) );
  NAND3_X1 U16203 ( .A1(n15774), .A2(n16202), .A3(n9304), .ZN(n16201) );
  NAND2_X1 U16204 ( .A1(n16118), .A2(n16119), .ZN(n16202) );
  NOR2_X1 U16205 ( .A1(n16118), .A2(n16119), .ZN(n16199) );
  NOR2_X1 U16206 ( .A1(n16203), .A2(n16204), .ZN(n16119) );
  NOR3_X1 U16207 ( .A1(n15773), .A2(n16205), .A3(n8572), .ZN(n16204) );
  NOR2_X1 U16208 ( .A1(n16114), .A2(n16115), .ZN(n16205) );
  INV_X1 U16209 ( .A(n16206), .ZN(n16203) );
  NAND2_X1 U16210 ( .A1(n16114), .A2(n16115), .ZN(n16206) );
  NAND2_X1 U16211 ( .A1(n16207), .A2(n16208), .ZN(n16115) );
  NAND3_X1 U16212 ( .A1(n15774), .A2(n16209), .A3(n9313), .ZN(n16208) );
  INV_X1 U16213 ( .A(n9031), .ZN(n9313) );
  INV_X1 U16214 ( .A(n16210), .ZN(n16209) );
  NOR2_X1 U16215 ( .A1(n16110), .A2(n16111), .ZN(n16210) );
  NAND2_X1 U16216 ( .A1(n16110), .A2(n16111), .ZN(n16207) );
  NAND2_X1 U16217 ( .A1(n16211), .A2(n16212), .ZN(n16111) );
  INV_X1 U16218 ( .A(n16213), .ZN(n16212) );
  NOR3_X1 U16219 ( .A1(n15773), .A2(n16214), .A3(n8591), .ZN(n16213) );
  NOR2_X1 U16220 ( .A1(n16105), .A2(n16107), .ZN(n16214) );
  NAND2_X1 U16221 ( .A1(n16105), .A2(n16107), .ZN(n16211) );
  NAND2_X1 U16222 ( .A1(n16215), .A2(n16216), .ZN(n16107) );
  NAND3_X1 U16223 ( .A1(n15774), .A2(n16217), .A3(n9322), .ZN(n16216) );
  INV_X1 U16224 ( .A(n16218), .ZN(n16217) );
  NOR2_X1 U16225 ( .A1(n16102), .A2(n16103), .ZN(n16218) );
  NAND2_X1 U16226 ( .A1(n16102), .A2(n16103), .ZN(n16215) );
  NAND2_X1 U16227 ( .A1(n16219), .A2(n16220), .ZN(n16103) );
  INV_X1 U16228 ( .A(n16221), .ZN(n16220) );
  NOR3_X1 U16229 ( .A1(n15773), .A2(n16222), .A3(n8545), .ZN(n16221) );
  NOR2_X1 U16230 ( .A1(n16097), .A2(n16099), .ZN(n16222) );
  NAND2_X1 U16231 ( .A1(n16097), .A2(n16099), .ZN(n16219) );
  NAND2_X1 U16232 ( .A1(n16223), .A2(n16224), .ZN(n16099) );
  NAND3_X1 U16233 ( .A1(n15774), .A2(n16225), .A3(n9331), .ZN(n16224) );
  INV_X1 U16234 ( .A(n9050), .ZN(n9331) );
  INV_X1 U16235 ( .A(n16226), .ZN(n16225) );
  NOR2_X1 U16236 ( .A1(n16094), .A2(n16095), .ZN(n16226) );
  NAND2_X1 U16237 ( .A1(n16094), .A2(n16095), .ZN(n16223) );
  NAND2_X1 U16238 ( .A1(n16227), .A2(n16228), .ZN(n16095) );
  INV_X1 U16239 ( .A(n16229), .ZN(n16228) );
  NOR3_X1 U16240 ( .A1(n15773), .A2(n16230), .A3(n8593), .ZN(n16229) );
  NOR2_X1 U16241 ( .A1(n16089), .A2(n16091), .ZN(n16230) );
  NAND2_X1 U16242 ( .A1(n16089), .A2(n16091), .ZN(n16227) );
  NAND2_X1 U16243 ( .A1(n16231), .A2(n16232), .ZN(n16091) );
  NAND3_X1 U16244 ( .A1(n15774), .A2(n16233), .A3(n9340), .ZN(n16232) );
  INV_X1 U16245 ( .A(n16234), .ZN(n16233) );
  NOR2_X1 U16246 ( .A1(n16086), .A2(n16087), .ZN(n16234) );
  NAND2_X1 U16247 ( .A1(n16086), .A2(n16087), .ZN(n16231) );
  NAND2_X1 U16248 ( .A1(n16235), .A2(n16236), .ZN(n16087) );
  INV_X1 U16249 ( .A(n16237), .ZN(n16236) );
  NOR3_X1 U16250 ( .A1(n9066), .A2(n16238), .A3(n8579), .ZN(n16237) );
  NOR2_X1 U16251 ( .A1(n16081), .A2(n16083), .ZN(n16238) );
  NAND2_X1 U16252 ( .A1(n16081), .A2(n16083), .ZN(n16235) );
  NAND2_X1 U16253 ( .A1(n16239), .A2(n16240), .ZN(n16083) );
  NAND3_X1 U16254 ( .A1(n9080), .A2(n16241), .A3(n15774), .ZN(n16240) );
  INV_X1 U16255 ( .A(n16242), .ZN(n16241) );
  NOR2_X1 U16256 ( .A1(n16078), .A2(n16079), .ZN(n16242) );
  INV_X1 U16257 ( .A(n9076), .ZN(n9080) );
  NAND2_X1 U16258 ( .A1(n16078), .A2(n16079), .ZN(n16239) );
  NAND2_X1 U16259 ( .A1(n16243), .A2(n16244), .ZN(n16079) );
  INV_X1 U16260 ( .A(n16245), .ZN(n16244) );
  NOR3_X1 U16261 ( .A1(n8551), .A2(n16246), .A3(n8579), .ZN(n16245) );
  NOR2_X1 U16262 ( .A1(n16073), .A2(n16075), .ZN(n16246) );
  NAND2_X1 U16263 ( .A1(n16073), .A2(n16075), .ZN(n16243) );
  NAND2_X1 U16264 ( .A1(n16247), .A2(n16248), .ZN(n16075) );
  NAND3_X1 U16265 ( .A1(n9098), .A2(n16249), .A3(n15774), .ZN(n16248) );
  INV_X1 U16266 ( .A(n16250), .ZN(n16249) );
  NOR2_X1 U16267 ( .A1(n16070), .A2(n16071), .ZN(n16250) );
  INV_X1 U16268 ( .A(n9094), .ZN(n9098) );
  NAND2_X1 U16269 ( .A1(n16070), .A2(n16071), .ZN(n16247) );
  NAND2_X1 U16270 ( .A1(n16251), .A2(n16252), .ZN(n16071) );
  NAND3_X1 U16271 ( .A1(n9107), .A2(n16253), .A3(n15774), .ZN(n16252) );
  NAND2_X1 U16272 ( .A1(n16065), .A2(n16067), .ZN(n16253) );
  INV_X1 U16273 ( .A(n16254), .ZN(n16251) );
  NOR2_X1 U16274 ( .A1(n16065), .A2(n16067), .ZN(n16254) );
  NOR2_X1 U16275 ( .A1(n16255), .A2(n16256), .ZN(n16067) );
  NOR3_X1 U16276 ( .A1(n9176), .A2(n16257), .A3(n8579), .ZN(n16256) );
  INV_X1 U16277 ( .A(n16258), .ZN(n16257) );
  NAND2_X1 U16278 ( .A1(n16006), .A2(n16007), .ZN(n16258) );
  NOR2_X1 U16279 ( .A1(n16006), .A2(n16007), .ZN(n16255) );
  NOR2_X1 U16280 ( .A1(n16259), .A2(n16260), .ZN(n16007) );
  INV_X1 U16281 ( .A(n16261), .ZN(n16260) );
  NAND3_X1 U16282 ( .A1(n9121), .A2(n16262), .A3(n15774), .ZN(n16261) );
  NAND2_X1 U16283 ( .A1(n16062), .A2(n16063), .ZN(n16262) );
  NOR2_X1 U16284 ( .A1(n16062), .A2(n16063), .ZN(n16259) );
  NOR2_X1 U16285 ( .A1(n16263), .A2(n16264), .ZN(n16063) );
  INV_X1 U16286 ( .A(n16265), .ZN(n16264) );
  NAND3_X1 U16287 ( .A1(n9373), .A2(n16266), .A3(n15774), .ZN(n16265) );
  NAND2_X1 U16288 ( .A1(n16058), .A2(n16059), .ZN(n16266) );
  NOR2_X1 U16289 ( .A1(n16058), .A2(n16059), .ZN(n16263) );
  NOR2_X1 U16290 ( .A1(n16267), .A2(n16268), .ZN(n16059) );
  INV_X1 U16291 ( .A(n16269), .ZN(n16268) );
  NAND2_X1 U16292 ( .A1(n16055), .A2(n16270), .ZN(n16269) );
  NAND2_X1 U16293 ( .A1(n16056), .A2(n16054), .ZN(n16270) );
  NOR2_X1 U16294 ( .A1(n15773), .A2(n9378), .ZN(n16055) );
  NOR2_X1 U16295 ( .A1(n16054), .A2(n16056), .ZN(n16267) );
  NOR2_X1 U16296 ( .A1(n16271), .A2(n16272), .ZN(n16056) );
  INV_X1 U16297 ( .A(n16273), .ZN(n16272) );
  NAND2_X1 U16298 ( .A1(n16051), .A2(n16274), .ZN(n16273) );
  NAND2_X1 U16299 ( .A1(n16052), .A2(n16050), .ZN(n16274) );
  NOR2_X1 U16300 ( .A1(n15773), .A2(n9383), .ZN(n16051) );
  NOR2_X1 U16301 ( .A1(n16050), .A2(n16052), .ZN(n16271) );
  NOR2_X1 U16302 ( .A1(n16275), .A2(n16276), .ZN(n16052) );
  INV_X1 U16303 ( .A(n16277), .ZN(n16276) );
  NAND2_X1 U16304 ( .A1(n16045), .A2(n16278), .ZN(n16277) );
  NAND2_X1 U16305 ( .A1(n16048), .A2(n16047), .ZN(n16278) );
  NOR2_X1 U16306 ( .A1(n15773), .A2(n9146), .ZN(n16045) );
  NOR2_X1 U16307 ( .A1(n16047), .A2(n16048), .ZN(n16275) );
  INV_X1 U16308 ( .A(n16279), .ZN(n16048) );
  NAND2_X1 U16309 ( .A1(n16280), .A2(n16281), .ZN(n16279) );
  NAND2_X1 U16310 ( .A1(n16040), .A2(n16282), .ZN(n16281) );
  NAND2_X1 U16311 ( .A1(n8624), .A2(n16283), .ZN(n16282) );
  NAND2_X1 U16312 ( .A1(n8590), .A2(n8627), .ZN(n16283) );
  NAND2_X1 U16313 ( .A1(n16285), .A2(n16286), .ZN(n16280) );
  NAND2_X1 U16314 ( .A1(n8630), .A2(n16287), .ZN(n16286) );
  NAND2_X1 U16315 ( .A1(n8539), .A2(n8577), .ZN(n16287) );
  NAND3_X1 U16316 ( .A1(n15774), .A2(n8537), .A3(n16040), .ZN(n16047) );
  XNOR2_X1 U16317 ( .A(n16288), .B(n16289), .ZN(n15773) );
  XOR2_X1 U16318 ( .A(d_3_), .B(c_3_), .Z(n16289) );
  XOR2_X1 U16319 ( .A(n16290), .B(n16291), .Z(n16050) );
  XNOR2_X1 U16320 ( .A(n16292), .B(n16293), .ZN(n16291) );
  XOR2_X1 U16321 ( .A(n16294), .B(n16295), .Z(n16054) );
  XNOR2_X1 U16322 ( .A(n16296), .B(n16297), .ZN(n16294) );
  XOR2_X1 U16323 ( .A(n16298), .B(n16299), .Z(n16058) );
  XNOR2_X1 U16324 ( .A(n16300), .B(n16301), .ZN(n16298) );
  XOR2_X1 U16325 ( .A(n16302), .B(n16303), .Z(n16062) );
  XNOR2_X1 U16326 ( .A(n16304), .B(n16305), .ZN(n16302) );
  XOR2_X1 U16327 ( .A(n16306), .B(n16307), .Z(n16006) );
  XNOR2_X1 U16328 ( .A(n16308), .B(n16309), .ZN(n16306) );
  XOR2_X1 U16329 ( .A(n16310), .B(n16311), .Z(n16065) );
  XNOR2_X1 U16330 ( .A(n16312), .B(n16313), .ZN(n16310) );
  XNOR2_X1 U16331 ( .A(n16314), .B(n16315), .ZN(n16070) );
  XNOR2_X1 U16332 ( .A(n16316), .B(n16317), .ZN(n16314) );
  XNOR2_X1 U16333 ( .A(n16318), .B(n16319), .ZN(n16073) );
  XNOR2_X1 U16334 ( .A(n16320), .B(n16321), .ZN(n16318) );
  XNOR2_X1 U16335 ( .A(n16322), .B(n16323), .ZN(n16078) );
  XNOR2_X1 U16336 ( .A(n16324), .B(n16325), .ZN(n16322) );
  XNOR2_X1 U16337 ( .A(n16326), .B(n16327), .ZN(n16081) );
  XNOR2_X1 U16338 ( .A(n16328), .B(n16329), .ZN(n16326) );
  XNOR2_X1 U16339 ( .A(n16330), .B(n16331), .ZN(n16086) );
  XNOR2_X1 U16340 ( .A(n16332), .B(n16333), .ZN(n16330) );
  XNOR2_X1 U16341 ( .A(n16334), .B(n16335), .ZN(n16089) );
  XNOR2_X1 U16342 ( .A(n16336), .B(n16337), .ZN(n16334) );
  XNOR2_X1 U16343 ( .A(n16338), .B(n16339), .ZN(n16094) );
  XNOR2_X1 U16344 ( .A(n16340), .B(n16341), .ZN(n16338) );
  XNOR2_X1 U16345 ( .A(n16342), .B(n16343), .ZN(n16097) );
  XNOR2_X1 U16346 ( .A(n16344), .B(n16345), .ZN(n16342) );
  XNOR2_X1 U16347 ( .A(n16346), .B(n16347), .ZN(n16102) );
  XNOR2_X1 U16348 ( .A(n16348), .B(n16349), .ZN(n16346) );
  XNOR2_X1 U16349 ( .A(n16350), .B(n16351), .ZN(n16105) );
  XNOR2_X1 U16350 ( .A(n16352), .B(n16353), .ZN(n16350) );
  XNOR2_X1 U16351 ( .A(n16354), .B(n16355), .ZN(n16110) );
  XNOR2_X1 U16352 ( .A(n16356), .B(n16357), .ZN(n16354) );
  XNOR2_X1 U16353 ( .A(n16358), .B(n16359), .ZN(n16114) );
  XNOR2_X1 U16354 ( .A(n16360), .B(n16361), .ZN(n16358) );
  XOR2_X1 U16355 ( .A(n16362), .B(n16363), .Z(n16118) );
  XNOR2_X1 U16356 ( .A(n16364), .B(n16365), .ZN(n16362) );
  XOR2_X1 U16357 ( .A(n16366), .B(n16367), .Z(n16122) );
  XNOR2_X1 U16358 ( .A(n16368), .B(n16369), .ZN(n16366) );
  XOR2_X1 U16359 ( .A(n16370), .B(n16371), .Z(n16126) );
  XNOR2_X1 U16360 ( .A(n16372), .B(n16373), .ZN(n16370) );
  XOR2_X1 U16361 ( .A(n16374), .B(n16375), .Z(n16130) );
  XNOR2_X1 U16362 ( .A(n16376), .B(n16377), .ZN(n16374) );
  XOR2_X1 U16363 ( .A(n16378), .B(n16379), .Z(n16134) );
  XNOR2_X1 U16364 ( .A(n16380), .B(n16381), .ZN(n16378) );
  XOR2_X1 U16365 ( .A(n16382), .B(n16383), .Z(n16138) );
  XNOR2_X1 U16366 ( .A(n16384), .B(n16385), .ZN(n16382) );
  XOR2_X1 U16367 ( .A(n16386), .B(n16387), .Z(n16142) );
  XNOR2_X1 U16368 ( .A(n16388), .B(n16389), .ZN(n16386) );
  XOR2_X1 U16369 ( .A(n16390), .B(n16391), .Z(n16146) );
  XNOR2_X1 U16370 ( .A(n16392), .B(n16393), .ZN(n16390) );
  XOR2_X1 U16371 ( .A(n16394), .B(n16395), .Z(n16150) );
  XNOR2_X1 U16372 ( .A(n16396), .B(n16397), .ZN(n16394) );
  XOR2_X1 U16373 ( .A(n16398), .B(n16399), .Z(n16153) );
  XNOR2_X1 U16374 ( .A(n16400), .B(n16401), .ZN(n16398) );
  XOR2_X1 U16375 ( .A(n8875), .B(n8873), .Z(n8779) );
  XOR2_X1 U16376 ( .A(n8883), .B(n16402), .Z(n8873) );
  NOR2_X1 U16377 ( .A1(n16403), .A2(n8886), .ZN(n16402) );
  NOR3_X1 U16378 ( .A1(n8884), .A2(n16404), .A3(n8885), .ZN(n8886) );
  INV_X1 U16379 ( .A(n16405), .ZN(n8885) );
  NOR2_X1 U16380 ( .A1(n16405), .A2(n16406), .ZN(n16403) );
  NOR2_X1 U16381 ( .A1(n16404), .A2(n8589), .ZN(n16406) );
  NOR2_X1 U16382 ( .A1(n8590), .A2(n8972), .ZN(n16405) );
  INV_X1 U16383 ( .A(n8872), .ZN(n8972) );
  NAND2_X1 U16384 ( .A1(n16407), .A2(n16408), .ZN(n8883) );
  NAND3_X1 U16385 ( .A1(n8874), .A2(n16409), .A3(n9268), .ZN(n16408) );
  NAND2_X1 U16386 ( .A1(n16410), .A2(n16411), .ZN(n16409) );
  NAND2_X1 U16387 ( .A1(n16412), .A2(n16413), .ZN(n16407) );
  NAND2_X1 U16388 ( .A1(n15897), .A2(n16414), .ZN(n8875) );
  NAND2_X1 U16389 ( .A1(n15896), .A2(n15898), .ZN(n16414) );
  NAND2_X1 U16390 ( .A1(n16415), .A2(n16416), .ZN(n15898) );
  NAND2_X1 U16391 ( .A1(n16040), .A2(n8872), .ZN(n16416) );
  XOR2_X1 U16392 ( .A(n16417), .B(n16418), .Z(n15896) );
  XNOR2_X1 U16393 ( .A(n16411), .B(n16410), .ZN(n16418) );
  INV_X1 U16394 ( .A(n16413), .ZN(n16410) );
  NAND2_X1 U16395 ( .A1(n16419), .A2(n16420), .ZN(n16413) );
  NAND2_X1 U16396 ( .A1(n16421), .A2(n16422), .ZN(n16420) );
  NAND2_X1 U16397 ( .A1(n8552), .A2(n16423), .ZN(n16421) );
  INV_X1 U16398 ( .A(n16412), .ZN(n16411) );
  NOR2_X1 U16399 ( .A1(n8884), .A2(n8590), .ZN(n16412) );
  NAND2_X1 U16400 ( .A1(n9268), .A2(n8874), .ZN(n16417) );
  NAND2_X1 U16401 ( .A1(n8592), .A2(n16424), .ZN(n15897) );
  INV_X1 U16402 ( .A(n16415), .ZN(n16424) );
  NOR2_X1 U16403 ( .A1(n16425), .A2(n16426), .ZN(n16415) );
  NOR3_X1 U16404 ( .A1(n16039), .A2(n16427), .A3(n8589), .ZN(n16426) );
  XNOR2_X1 U16405 ( .A(n16428), .B(n16429), .ZN(n8884) );
  XNOR2_X1 U16406 ( .A(n16430), .B(a_1_), .ZN(n16429) );
  INV_X1 U16407 ( .A(n16431), .ZN(n16427) );
  NAND2_X1 U16408 ( .A1(n16160), .A2(n16159), .ZN(n16431) );
  NOR2_X1 U16409 ( .A1(n16159), .A2(n16160), .ZN(n16425) );
  NOR2_X1 U16410 ( .A1(n16432), .A2(n16433), .ZN(n16160) );
  INV_X1 U16411 ( .A(n16434), .ZN(n16433) );
  NAND2_X1 U16412 ( .A1(n16400), .A2(n16435), .ZN(n16434) );
  NAND2_X1 U16413 ( .A1(n16401), .A2(n16399), .ZN(n16435) );
  NOR2_X1 U16414 ( .A1(n8982), .A2(n8577), .ZN(n16400) );
  NOR2_X1 U16415 ( .A1(n16399), .A2(n16401), .ZN(n16432) );
  NOR2_X1 U16416 ( .A1(n16436), .A2(n16437), .ZN(n16401) );
  INV_X1 U16417 ( .A(n16438), .ZN(n16437) );
  NAND2_X1 U16418 ( .A1(n16397), .A2(n16439), .ZN(n16438) );
  NAND2_X1 U16419 ( .A1(n16396), .A2(n16395), .ZN(n16439) );
  NOR2_X1 U16420 ( .A1(n8527), .A2(n8577), .ZN(n16397) );
  NOR2_X1 U16421 ( .A1(n16395), .A2(n16396), .ZN(n16436) );
  NOR2_X1 U16422 ( .A1(n16440), .A2(n16441), .ZN(n16396) );
  INV_X1 U16423 ( .A(n16442), .ZN(n16441) );
  NAND2_X1 U16424 ( .A1(n16392), .A2(n16443), .ZN(n16442) );
  NAND2_X1 U16425 ( .A1(n16393), .A2(n16391), .ZN(n16443) );
  NOR2_X1 U16426 ( .A1(n8528), .A2(n8577), .ZN(n16392) );
  NOR2_X1 U16427 ( .A1(n16391), .A2(n16393), .ZN(n16440) );
  NOR2_X1 U16428 ( .A1(n16444), .A2(n16445), .ZN(n16393) );
  INV_X1 U16429 ( .A(n16446), .ZN(n16445) );
  NAND2_X1 U16430 ( .A1(n16389), .A2(n16447), .ZN(n16446) );
  NAND2_X1 U16431 ( .A1(n16388), .A2(n16387), .ZN(n16447) );
  NOR2_X1 U16432 ( .A1(n8995), .A2(n8577), .ZN(n16389) );
  NOR2_X1 U16433 ( .A1(n16387), .A2(n16388), .ZN(n16444) );
  NOR2_X1 U16434 ( .A1(n16448), .A2(n16449), .ZN(n16388) );
  INV_X1 U16435 ( .A(n16450), .ZN(n16449) );
  NAND2_X1 U16436 ( .A1(n16384), .A2(n16451), .ZN(n16450) );
  NAND2_X1 U16437 ( .A1(n16385), .A2(n16383), .ZN(n16451) );
  NOR2_X1 U16438 ( .A1(n9000), .A2(n8577), .ZN(n16384) );
  NOR2_X1 U16439 ( .A1(n16383), .A2(n16385), .ZN(n16448) );
  NOR2_X1 U16440 ( .A1(n16452), .A2(n16453), .ZN(n16385) );
  INV_X1 U16441 ( .A(n16454), .ZN(n16453) );
  NAND2_X1 U16442 ( .A1(n16381), .A2(n16455), .ZN(n16454) );
  NAND2_X1 U16443 ( .A1(n16380), .A2(n16379), .ZN(n16455) );
  NOR2_X1 U16444 ( .A1(n8544), .A2(n8577), .ZN(n16381) );
  NOR2_X1 U16445 ( .A1(n16379), .A2(n16380), .ZN(n16452) );
  NOR2_X1 U16446 ( .A1(n16456), .A2(n16457), .ZN(n16380) );
  INV_X1 U16447 ( .A(n16458), .ZN(n16457) );
  NAND2_X1 U16448 ( .A1(n16376), .A2(n16459), .ZN(n16458) );
  NAND2_X1 U16449 ( .A1(n16377), .A2(n16375), .ZN(n16459) );
  NOR2_X1 U16450 ( .A1(n9010), .A2(n8577), .ZN(n16376) );
  NOR2_X1 U16451 ( .A1(n16375), .A2(n16377), .ZN(n16456) );
  NOR2_X1 U16452 ( .A1(n16460), .A2(n16461), .ZN(n16377) );
  INV_X1 U16453 ( .A(n16462), .ZN(n16461) );
  NAND2_X1 U16454 ( .A1(n16373), .A2(n16463), .ZN(n16462) );
  NAND2_X1 U16455 ( .A1(n16372), .A2(n16371), .ZN(n16463) );
  NOR2_X1 U16456 ( .A1(n8594), .A2(n8577), .ZN(n16373) );
  NOR2_X1 U16457 ( .A1(n16371), .A2(n16372), .ZN(n16460) );
  NOR2_X1 U16458 ( .A1(n16464), .A2(n16465), .ZN(n16372) );
  INV_X1 U16459 ( .A(n16466), .ZN(n16465) );
  NAND2_X1 U16460 ( .A1(n16368), .A2(n16467), .ZN(n16466) );
  NAND2_X1 U16461 ( .A1(n16369), .A2(n16367), .ZN(n16467) );
  NOR2_X1 U16462 ( .A1(n9020), .A2(n8577), .ZN(n16368) );
  NOR2_X1 U16463 ( .A1(n16367), .A2(n16369), .ZN(n16464) );
  NOR2_X1 U16464 ( .A1(n16468), .A2(n16469), .ZN(n16369) );
  INV_X1 U16465 ( .A(n16470), .ZN(n16469) );
  NAND2_X1 U16466 ( .A1(n16365), .A2(n16471), .ZN(n16470) );
  NAND2_X1 U16467 ( .A1(n16364), .A2(n16363), .ZN(n16471) );
  NOR2_X1 U16468 ( .A1(n9025), .A2(n8577), .ZN(n16365) );
  NOR2_X1 U16469 ( .A1(n16363), .A2(n16364), .ZN(n16468) );
  NOR2_X1 U16470 ( .A1(n16472), .A2(n16473), .ZN(n16364) );
  INV_X1 U16471 ( .A(n16474), .ZN(n16473) );
  NAND2_X1 U16472 ( .A1(n16360), .A2(n16475), .ZN(n16474) );
  NAND2_X1 U16473 ( .A1(n16361), .A2(n16359), .ZN(n16475) );
  NOR2_X1 U16474 ( .A1(n9031), .A2(n8577), .ZN(n16360) );
  NOR2_X1 U16475 ( .A1(n16359), .A2(n16361), .ZN(n16472) );
  NOR2_X1 U16476 ( .A1(n16476), .A2(n16477), .ZN(n16361) );
  INV_X1 U16477 ( .A(n16478), .ZN(n16477) );
  NAND2_X1 U16478 ( .A1(n16357), .A2(n16479), .ZN(n16478) );
  NAND2_X1 U16479 ( .A1(n16356), .A2(n16355), .ZN(n16479) );
  NOR2_X1 U16480 ( .A1(n9036), .A2(n8577), .ZN(n16357) );
  NOR2_X1 U16481 ( .A1(n16355), .A2(n16356), .ZN(n16476) );
  NOR2_X1 U16482 ( .A1(n16480), .A2(n16481), .ZN(n16356) );
  INV_X1 U16483 ( .A(n16482), .ZN(n16481) );
  NAND2_X1 U16484 ( .A1(n16352), .A2(n16483), .ZN(n16482) );
  NAND2_X1 U16485 ( .A1(n16353), .A2(n16351), .ZN(n16483) );
  NOR2_X1 U16486 ( .A1(n9041), .A2(n8577), .ZN(n16352) );
  NOR2_X1 U16487 ( .A1(n16351), .A2(n16353), .ZN(n16480) );
  NOR2_X1 U16488 ( .A1(n16484), .A2(n16485), .ZN(n16353) );
  INV_X1 U16489 ( .A(n16486), .ZN(n16485) );
  NAND2_X1 U16490 ( .A1(n16349), .A2(n16487), .ZN(n16486) );
  NAND2_X1 U16491 ( .A1(n16348), .A2(n16347), .ZN(n16487) );
  NOR2_X1 U16492 ( .A1(n8545), .A2(n8577), .ZN(n16349) );
  NOR2_X1 U16493 ( .A1(n16347), .A2(n16348), .ZN(n16484) );
  NOR2_X1 U16494 ( .A1(n16488), .A2(n16489), .ZN(n16348) );
  INV_X1 U16495 ( .A(n16490), .ZN(n16489) );
  NAND2_X1 U16496 ( .A1(n16344), .A2(n16491), .ZN(n16490) );
  NAND2_X1 U16497 ( .A1(n16345), .A2(n16343), .ZN(n16491) );
  NOR2_X1 U16498 ( .A1(n9050), .A2(n8577), .ZN(n16344) );
  NOR2_X1 U16499 ( .A1(n16343), .A2(n16345), .ZN(n16488) );
  NOR2_X1 U16500 ( .A1(n16492), .A2(n16493), .ZN(n16345) );
  INV_X1 U16501 ( .A(n16494), .ZN(n16493) );
  NAND2_X1 U16502 ( .A1(n16341), .A2(n16495), .ZN(n16494) );
  NAND2_X1 U16503 ( .A1(n16340), .A2(n16339), .ZN(n16495) );
  NOR2_X1 U16504 ( .A1(n8593), .A2(n8577), .ZN(n16341) );
  NOR2_X1 U16505 ( .A1(n16339), .A2(n16340), .ZN(n16492) );
  NOR2_X1 U16506 ( .A1(n16496), .A2(n16497), .ZN(n16340) );
  INV_X1 U16507 ( .A(n16498), .ZN(n16497) );
  NAND2_X1 U16508 ( .A1(n16336), .A2(n16499), .ZN(n16498) );
  NAND2_X1 U16509 ( .A1(n16337), .A2(n16335), .ZN(n16499) );
  NOR2_X1 U16510 ( .A1(n9061), .A2(n8577), .ZN(n16336) );
  NOR2_X1 U16511 ( .A1(n16335), .A2(n16337), .ZN(n16496) );
  NOR2_X1 U16512 ( .A1(n16500), .A2(n16501), .ZN(n16337) );
  INV_X1 U16513 ( .A(n16502), .ZN(n16501) );
  NAND2_X1 U16514 ( .A1(n16333), .A2(n16503), .ZN(n16502) );
  NAND2_X1 U16515 ( .A1(n16332), .A2(n16331), .ZN(n16503) );
  NOR2_X1 U16516 ( .A1(n8577), .A2(n8580), .ZN(n16333) );
  NOR2_X1 U16517 ( .A1(n16331), .A2(n16332), .ZN(n16500) );
  NOR2_X1 U16518 ( .A1(n16504), .A2(n16505), .ZN(n16332) );
  INV_X1 U16519 ( .A(n16506), .ZN(n16505) );
  NAND2_X1 U16520 ( .A1(n16328), .A2(n16507), .ZN(n16506) );
  NAND2_X1 U16521 ( .A1(n16329), .A2(n16327), .ZN(n16507) );
  NOR2_X1 U16522 ( .A1(n8577), .A2(n8588), .ZN(n16328) );
  NOR2_X1 U16523 ( .A1(n16327), .A2(n16329), .ZN(n16504) );
  NOR2_X1 U16524 ( .A1(n16508), .A2(n16509), .ZN(n16329) );
  INV_X1 U16525 ( .A(n16510), .ZN(n16509) );
  NAND2_X1 U16526 ( .A1(n16325), .A2(n16511), .ZN(n16510) );
  NAND2_X1 U16527 ( .A1(n16324), .A2(n16323), .ZN(n16511) );
  NOR2_X1 U16528 ( .A1(n8577), .A2(n8551), .ZN(n16325) );
  NOR2_X1 U16529 ( .A1(n16323), .A2(n16324), .ZN(n16508) );
  NOR2_X1 U16530 ( .A1(n16512), .A2(n16513), .ZN(n16324) );
  INV_X1 U16531 ( .A(n16514), .ZN(n16513) );
  NAND2_X1 U16532 ( .A1(n16320), .A2(n16515), .ZN(n16514) );
  NAND2_X1 U16533 ( .A1(n16321), .A2(n16319), .ZN(n16515) );
  NOR2_X1 U16534 ( .A1(n8577), .A2(n8563), .ZN(n16320) );
  NOR2_X1 U16535 ( .A1(n16319), .A2(n16321), .ZN(n16512) );
  NOR2_X1 U16536 ( .A1(n16516), .A2(n16517), .ZN(n16321) );
  INV_X1 U16537 ( .A(n16518), .ZN(n16517) );
  NAND2_X1 U16538 ( .A1(n16317), .A2(n16519), .ZN(n16518) );
  NAND2_X1 U16539 ( .A1(n16316), .A2(n16315), .ZN(n16519) );
  NOR2_X1 U16540 ( .A1(n8577), .A2(n8548), .ZN(n16317) );
  NOR2_X1 U16541 ( .A1(n16315), .A2(n16316), .ZN(n16516) );
  NOR2_X1 U16542 ( .A1(n16520), .A2(n16521), .ZN(n16316) );
  INV_X1 U16543 ( .A(n16522), .ZN(n16521) );
  NAND2_X1 U16544 ( .A1(n16312), .A2(n16523), .ZN(n16522) );
  NAND2_X1 U16545 ( .A1(n16313), .A2(n16311), .ZN(n16523) );
  NOR2_X1 U16546 ( .A1(n16039), .A2(n8584), .ZN(n16312) );
  NOR2_X1 U16547 ( .A1(n16311), .A2(n16313), .ZN(n16520) );
  NOR2_X1 U16548 ( .A1(n16524), .A2(n16525), .ZN(n16313) );
  INV_X1 U16549 ( .A(n16526), .ZN(n16525) );
  NAND2_X1 U16550 ( .A1(n16309), .A2(n16527), .ZN(n16526) );
  NAND2_X1 U16551 ( .A1(n16308), .A2(n16307), .ZN(n16527) );
  NOR2_X1 U16552 ( .A1(n16039), .A2(n8535), .ZN(n16309) );
  NOR2_X1 U16553 ( .A1(n16307), .A2(n16308), .ZN(n16524) );
  NOR2_X1 U16554 ( .A1(n16528), .A2(n16529), .ZN(n16308) );
  INV_X1 U16555 ( .A(n16530), .ZN(n16529) );
  NAND2_X1 U16556 ( .A1(n16304), .A2(n16531), .ZN(n16530) );
  NAND2_X1 U16557 ( .A1(n16305), .A2(n16303), .ZN(n16531) );
  NOR2_X1 U16558 ( .A1(n16039), .A2(n9126), .ZN(n16304) );
  NOR2_X1 U16559 ( .A1(n16303), .A2(n16305), .ZN(n16528) );
  NOR2_X1 U16560 ( .A1(n16532), .A2(n16533), .ZN(n16305) );
  INV_X1 U16561 ( .A(n16534), .ZN(n16533) );
  NAND2_X1 U16562 ( .A1(n16301), .A2(n16535), .ZN(n16534) );
  NAND2_X1 U16563 ( .A1(n16300), .A2(n16299), .ZN(n16535) );
  NOR2_X1 U16564 ( .A1(n16039), .A2(n9378), .ZN(n16301) );
  NOR2_X1 U16565 ( .A1(n16299), .A2(n16300), .ZN(n16532) );
  NOR2_X1 U16566 ( .A1(n16536), .A2(n16537), .ZN(n16300) );
  INV_X1 U16567 ( .A(n16538), .ZN(n16537) );
  NAND2_X1 U16568 ( .A1(n16296), .A2(n16539), .ZN(n16538) );
  NAND2_X1 U16569 ( .A1(n16295), .A2(n16297), .ZN(n16539) );
  NOR2_X1 U16570 ( .A1(n16039), .A2(n9383), .ZN(n16296) );
  NOR2_X1 U16571 ( .A1(n16295), .A2(n16297), .ZN(n16536) );
  NOR2_X1 U16572 ( .A1(n16540), .A2(n16541), .ZN(n16297) );
  INV_X1 U16573 ( .A(n16542), .ZN(n16541) );
  NAND2_X1 U16574 ( .A1(n16290), .A2(n16543), .ZN(n16542) );
  NAND2_X1 U16575 ( .A1(n16293), .A2(n16292), .ZN(n16543) );
  NOR2_X1 U16576 ( .A1(n16039), .A2(n9146), .ZN(n16290) );
  NOR2_X1 U16577 ( .A1(n16292), .A2(n16293), .ZN(n16540) );
  INV_X1 U16578 ( .A(n16544), .ZN(n16293) );
  NAND2_X1 U16579 ( .A1(n16545), .A2(n16546), .ZN(n16544) );
  NAND2_X1 U16580 ( .A1(n16285), .A2(n16547), .ZN(n16546) );
  NAND2_X1 U16581 ( .A1(n8624), .A2(n16548), .ZN(n16547) );
  NAND2_X1 U16582 ( .A1(n16404), .A2(n8627), .ZN(n16548) );
  NAND2_X1 U16583 ( .A1(n8874), .A2(n16549), .ZN(n16545) );
  NAND2_X1 U16584 ( .A1(n8630), .A2(n16550), .ZN(n16549) );
  NAND2_X1 U16585 ( .A1(n8539), .A2(n8590), .ZN(n16550) );
  NAND3_X1 U16586 ( .A1(n16040), .A2(n8537), .A3(n16285), .ZN(n16292) );
  INV_X1 U16587 ( .A(n16039), .ZN(n16040) );
  XNOR2_X1 U16588 ( .A(n16552), .B(n16553), .ZN(n16039) );
  XOR2_X1 U16589 ( .A(d_2_), .B(c_2_), .Z(n16553) );
  XOR2_X1 U16590 ( .A(n16554), .B(n16555), .Z(n16295) );
  NOR2_X1 U16591 ( .A1(n16551), .A2(n16404), .ZN(n16555) );
  XOR2_X1 U16592 ( .A(n16556), .B(n16557), .Z(n16554) );
  XNOR2_X1 U16593 ( .A(n16558), .B(n16559), .ZN(n16299) );
  NOR2_X1 U16594 ( .A1(n9383), .A2(n8590), .ZN(n16559) );
  XOR2_X1 U16595 ( .A(n16560), .B(n16561), .Z(n16558) );
  XOR2_X1 U16596 ( .A(n16562), .B(n16563), .Z(n16303) );
  NAND2_X1 U16597 ( .A1(n16564), .A2(n16565), .ZN(n16562) );
  NAND2_X1 U16598 ( .A1(n16566), .A2(n16567), .ZN(n16565) );
  NAND2_X1 U16599 ( .A1(n16285), .A2(n9132), .ZN(n16566) );
  INV_X1 U16600 ( .A(n9378), .ZN(n9132) );
  XNOR2_X1 U16601 ( .A(n16568), .B(n16569), .ZN(n16307) );
  XNOR2_X1 U16602 ( .A(n16570), .B(n16571), .ZN(n16569) );
  NAND2_X1 U16603 ( .A1(n16285), .A2(n9373), .ZN(n16568) );
  XNOR2_X1 U16604 ( .A(n16572), .B(n16573), .ZN(n16311) );
  NOR2_X1 U16605 ( .A1(n8535), .A2(n8590), .ZN(n16573) );
  XOR2_X1 U16606 ( .A(n16574), .B(n16575), .Z(n16572) );
  XNOR2_X1 U16607 ( .A(n16576), .B(n16577), .ZN(n16315) );
  NOR2_X1 U16608 ( .A1(n16578), .A2(n16579), .ZN(n16577) );
  NOR2_X1 U16609 ( .A1(n16580), .A2(n16581), .ZN(n16578) );
  NOR2_X1 U16610 ( .A1(n9176), .A2(n8590), .ZN(n16581) );
  INV_X1 U16611 ( .A(n16582), .ZN(n16580) );
  XNOR2_X1 U16612 ( .A(n16583), .B(n16584), .ZN(n16319) );
  XNOR2_X1 U16613 ( .A(n16585), .B(n16586), .ZN(n16584) );
  NAND2_X1 U16614 ( .A1(n16285), .A2(n9107), .ZN(n16583) );
  XNOR2_X1 U16615 ( .A(n16587), .B(n16588), .ZN(n16323) );
  NOR2_X1 U16616 ( .A1(n16589), .A2(n16590), .ZN(n16588) );
  NOR2_X1 U16617 ( .A1(n16591), .A2(n16592), .ZN(n16589) );
  NOR2_X1 U16618 ( .A1(n9094), .A2(n8590), .ZN(n16592) );
  INV_X1 U16619 ( .A(n16593), .ZN(n16591) );
  XNOR2_X1 U16620 ( .A(n16594), .B(n16595), .ZN(n16327) );
  NOR2_X1 U16621 ( .A1(n8551), .A2(n8590), .ZN(n16595) );
  XOR2_X1 U16622 ( .A(n16596), .B(n16597), .Z(n16594) );
  XNOR2_X1 U16623 ( .A(n16598), .B(n16599), .ZN(n16331) );
  NOR2_X1 U16624 ( .A1(n16600), .A2(n16601), .ZN(n16599) );
  NOR2_X1 U16625 ( .A1(n16602), .A2(n16603), .ZN(n16600) );
  NOR2_X1 U16626 ( .A1(n9076), .A2(n8590), .ZN(n16603) );
  INV_X1 U16627 ( .A(n16604), .ZN(n16602) );
  XNOR2_X1 U16628 ( .A(n16605), .B(n16606), .ZN(n16335) );
  XNOR2_X1 U16629 ( .A(n16607), .B(n16608), .ZN(n16606) );
  NAND2_X1 U16630 ( .A1(n16285), .A2(n9070), .ZN(n16605) );
  XOR2_X1 U16631 ( .A(n16609), .B(n16610), .Z(n16339) );
  NAND2_X1 U16632 ( .A1(n16611), .A2(n16612), .ZN(n16609) );
  NAND2_X1 U16633 ( .A1(n16613), .A2(n16614), .ZN(n16612) );
  NAND2_X1 U16634 ( .A1(n9340), .A2(n16285), .ZN(n16613) );
  INV_X1 U16635 ( .A(n9061), .ZN(n9340) );
  XNOR2_X1 U16636 ( .A(n16615), .B(n16616), .ZN(n16343) );
  XNOR2_X1 U16637 ( .A(n16617), .B(n16618), .ZN(n16616) );
  NAND2_X1 U16638 ( .A1(n10722), .A2(n16285), .ZN(n16615) );
  XNOR2_X1 U16639 ( .A(n16619), .B(n16620), .ZN(n16347) );
  NOR2_X1 U16640 ( .A1(n16621), .A2(n16622), .ZN(n16620) );
  NOR2_X1 U16641 ( .A1(n16623), .A2(n16624), .ZN(n16621) );
  NOR2_X1 U16642 ( .A1(n8590), .A2(n8569), .ZN(n16624) );
  INV_X1 U16643 ( .A(n16625), .ZN(n16623) );
  XNOR2_X1 U16644 ( .A(n16626), .B(n16627), .ZN(n16351) );
  XNOR2_X1 U16645 ( .A(n16628), .B(n16629), .ZN(n16627) );
  NAND2_X1 U16646 ( .A1(n10222), .A2(n16285), .ZN(n16626) );
  XOR2_X1 U16647 ( .A(n16630), .B(n16631), .Z(n16355) );
  NAND2_X1 U16648 ( .A1(n16632), .A2(n16633), .ZN(n16630) );
  NAND2_X1 U16649 ( .A1(n16634), .A2(n16635), .ZN(n16633) );
  NAND2_X1 U16650 ( .A1(n9322), .A2(n16285), .ZN(n16634) );
  INV_X1 U16651 ( .A(n9041), .ZN(n9322) );
  XNOR2_X1 U16652 ( .A(n16636), .B(n16637), .ZN(n16359) );
  XNOR2_X1 U16653 ( .A(n16638), .B(n16639), .ZN(n16637) );
  NAND2_X1 U16654 ( .A1(n9721), .A2(n16285), .ZN(n16636) );
  XNOR2_X1 U16655 ( .A(n16640), .B(n16641), .ZN(n16363) );
  NOR2_X1 U16656 ( .A1(n16642), .A2(n16643), .ZN(n16641) );
  NOR2_X1 U16657 ( .A1(n16644), .A2(n16645), .ZN(n16642) );
  NOR2_X1 U16658 ( .A1(n8590), .A2(n8582), .ZN(n16645) );
  INV_X1 U16659 ( .A(n16646), .ZN(n16644) );
  XNOR2_X1 U16660 ( .A(n16647), .B(n16648), .ZN(n16367) );
  XNOR2_X1 U16661 ( .A(n16649), .B(n16650), .ZN(n16648) );
  NAND2_X1 U16662 ( .A1(n9209), .A2(n16285), .ZN(n16647) );
  XOR2_X1 U16663 ( .A(n16651), .B(n16652), .Z(n16371) );
  NAND2_X1 U16664 ( .A1(n16653), .A2(n16654), .ZN(n16651) );
  NAND2_X1 U16665 ( .A1(n16655), .A2(n16656), .ZN(n16654) );
  NAND2_X1 U16666 ( .A1(n9304), .A2(n16285), .ZN(n16655) );
  INV_X1 U16667 ( .A(n9020), .ZN(n9304) );
  XNOR2_X1 U16668 ( .A(n16657), .B(n16658), .ZN(n16375) );
  XNOR2_X1 U16669 ( .A(n16659), .B(n16660), .ZN(n16658) );
  NAND2_X1 U16670 ( .A1(n10846), .A2(n16285), .ZN(n16657) );
  XNOR2_X1 U16671 ( .A(n16661), .B(n16662), .ZN(n16379) );
  NOR2_X1 U16672 ( .A1(n16663), .A2(n16664), .ZN(n16662) );
  NOR2_X1 U16673 ( .A1(n16665), .A2(n16666), .ZN(n16663) );
  NOR2_X1 U16674 ( .A1(n8590), .A2(n8560), .ZN(n16666) );
  XNOR2_X1 U16675 ( .A(n16667), .B(n16668), .ZN(n16383) );
  NOR2_X1 U16676 ( .A1(n8590), .A2(n8544), .ZN(n16668) );
  XOR2_X1 U16677 ( .A(n16669), .B(n16670), .Z(n16667) );
  XOR2_X1 U16678 ( .A(n16671), .B(n16672), .Z(n16387) );
  NAND2_X1 U16679 ( .A1(n16673), .A2(n16674), .ZN(n16671) );
  NAND2_X1 U16680 ( .A1(n16675), .A2(n16676), .ZN(n16674) );
  NAND2_X1 U16681 ( .A1(n9286), .A2(n16285), .ZN(n16675) );
  INV_X1 U16682 ( .A(n9000), .ZN(n9286) );
  XNOR2_X1 U16683 ( .A(n16677), .B(n16678), .ZN(n16391) );
  XNOR2_X1 U16684 ( .A(n16679), .B(n16680), .ZN(n16678) );
  NAND2_X1 U16685 ( .A1(n10307), .A2(n16285), .ZN(n16677) );
  XNOR2_X1 U16686 ( .A(n16681), .B(n16682), .ZN(n16395) );
  NOR2_X1 U16687 ( .A1(n16683), .A2(n16684), .ZN(n16682) );
  NOR2_X1 U16688 ( .A1(n16685), .A2(n16686), .ZN(n16683) );
  NOR2_X1 U16689 ( .A1(n8590), .A2(n8528), .ZN(n16686) );
  XNOR2_X1 U16690 ( .A(n16687), .B(n16688), .ZN(n16399) );
  NOR2_X1 U16691 ( .A1(n8590), .A2(n8527), .ZN(n16688) );
  XOR2_X1 U16692 ( .A(n16689), .B(n16690), .Z(n16687) );
  XOR2_X1 U16693 ( .A(n16691), .B(n16422), .Z(n16159) );
  NAND2_X1 U16694 ( .A1(n16692), .A2(n16693), .ZN(n16422) );
  NAND3_X1 U16695 ( .A1(n16285), .A2(n16694), .A3(n9792), .ZN(n16693) );
  NAND2_X1 U16696 ( .A1(n16689), .A2(n16690), .ZN(n16694) );
  INV_X1 U16697 ( .A(n16695), .ZN(n16692) );
  NOR2_X1 U16698 ( .A1(n16690), .A2(n16689), .ZN(n16695) );
  NOR2_X1 U16699 ( .A1(n16684), .A2(n16696), .ZN(n16689) );
  INV_X1 U16700 ( .A(n16697), .ZN(n16696) );
  NAND2_X1 U16701 ( .A1(n16698), .A2(n16681), .ZN(n16697) );
  NAND2_X1 U16702 ( .A1(n16699), .A2(n16700), .ZN(n16681) );
  NAND3_X1 U16703 ( .A1(n16285), .A2(n16701), .A3(n10307), .ZN(n16700) );
  INV_X1 U16704 ( .A(n8995), .ZN(n10307) );
  NAND2_X1 U16705 ( .A1(n16680), .A2(n16679), .ZN(n16701) );
  INV_X1 U16706 ( .A(n16702), .ZN(n16679) );
  INV_X1 U16707 ( .A(n16703), .ZN(n16680) );
  NAND2_X1 U16708 ( .A1(n16702), .A2(n16703), .ZN(n16699) );
  NAND2_X1 U16709 ( .A1(n16673), .A2(n16704), .ZN(n16703) );
  NAND2_X1 U16710 ( .A1(n16705), .A2(n16672), .ZN(n16704) );
  NAND2_X1 U16711 ( .A1(n16706), .A2(n16707), .ZN(n16672) );
  NAND3_X1 U16712 ( .A1(n16285), .A2(n16708), .A3(n8543), .ZN(n16707) );
  NAND2_X1 U16713 ( .A1(n16669), .A2(n16670), .ZN(n16708) );
  INV_X1 U16714 ( .A(n16709), .ZN(n16706) );
  NOR2_X1 U16715 ( .A1(n16670), .A2(n16669), .ZN(n16709) );
  NOR2_X1 U16716 ( .A1(n16664), .A2(n16710), .ZN(n16669) );
  INV_X1 U16717 ( .A(n16711), .ZN(n16710) );
  NAND2_X1 U16718 ( .A1(n16712), .A2(n16661), .ZN(n16711) );
  NAND2_X1 U16719 ( .A1(n16713), .A2(n16714), .ZN(n16661) );
  NAND3_X1 U16720 ( .A1(n16285), .A2(n16715), .A3(n10846), .ZN(n16714) );
  INV_X1 U16721 ( .A(n9014), .ZN(n10846) );
  NAND2_X1 U16722 ( .A1(n16660), .A2(n16659), .ZN(n16715) );
  INV_X1 U16723 ( .A(n16716), .ZN(n16659) );
  INV_X1 U16724 ( .A(n16717), .ZN(n16660) );
  NAND2_X1 U16725 ( .A1(n16716), .A2(n16717), .ZN(n16713) );
  NAND2_X1 U16726 ( .A1(n16653), .A2(n16718), .ZN(n16717) );
  NAND2_X1 U16727 ( .A1(n16719), .A2(n16652), .ZN(n16718) );
  NAND2_X1 U16728 ( .A1(n16720), .A2(n16721), .ZN(n16652) );
  NAND3_X1 U16729 ( .A1(n16285), .A2(n16722), .A3(n9209), .ZN(n16721) );
  INV_X1 U16730 ( .A(n16723), .ZN(n16722) );
  NOR2_X1 U16731 ( .A1(n16650), .A2(n16649), .ZN(n16723) );
  NAND2_X1 U16732 ( .A1(n16649), .A2(n16650), .ZN(n16720) );
  NAND2_X1 U16733 ( .A1(n16724), .A2(n16725), .ZN(n16650) );
  NAND2_X1 U16734 ( .A1(n16726), .A2(n16640), .ZN(n16725) );
  NAND2_X1 U16735 ( .A1(n16727), .A2(n16728), .ZN(n16640) );
  INV_X1 U16736 ( .A(n16729), .ZN(n16728) );
  NOR3_X1 U16737 ( .A1(n8590), .A2(n16730), .A3(n8591), .ZN(n16729) );
  NOR2_X1 U16738 ( .A1(n16639), .A2(n16638), .ZN(n16730) );
  NAND2_X1 U16739 ( .A1(n16638), .A2(n16639), .ZN(n16727) );
  NAND2_X1 U16740 ( .A1(n16632), .A2(n16731), .ZN(n16639) );
  NAND2_X1 U16741 ( .A1(n16732), .A2(n16631), .ZN(n16731) );
  NAND2_X1 U16742 ( .A1(n16733), .A2(n16734), .ZN(n16631) );
  NAND3_X1 U16743 ( .A1(n16285), .A2(n16735), .A3(n10222), .ZN(n16734) );
  INV_X1 U16744 ( .A(n16736), .ZN(n16735) );
  NOR2_X1 U16745 ( .A1(n16629), .A2(n16628), .ZN(n16736) );
  NAND2_X1 U16746 ( .A1(n16628), .A2(n16629), .ZN(n16733) );
  NAND2_X1 U16747 ( .A1(n16737), .A2(n16738), .ZN(n16629) );
  NAND2_X1 U16748 ( .A1(n16739), .A2(n16619), .ZN(n16738) );
  NAND2_X1 U16749 ( .A1(n16740), .A2(n16741), .ZN(n16619) );
  INV_X1 U16750 ( .A(n16742), .ZN(n16741) );
  NOR3_X1 U16751 ( .A1(n16284), .A2(n16743), .A3(n8593), .ZN(n16742) );
  NOR2_X1 U16752 ( .A1(n16618), .A2(n16617), .ZN(n16743) );
  NAND2_X1 U16753 ( .A1(n16617), .A2(n16618), .ZN(n16740) );
  NAND2_X1 U16754 ( .A1(n16611), .A2(n16744), .ZN(n16618) );
  NAND2_X1 U16755 ( .A1(n16745), .A2(n16610), .ZN(n16744) );
  NAND2_X1 U16756 ( .A1(n16746), .A2(n16747), .ZN(n16610) );
  NAND3_X1 U16757 ( .A1(n9070), .A2(n16748), .A3(n16285), .ZN(n16747) );
  INV_X1 U16758 ( .A(n16749), .ZN(n16748) );
  NOR2_X1 U16759 ( .A1(n16608), .A2(n16607), .ZN(n16749) );
  NAND2_X1 U16760 ( .A1(n16607), .A2(n16608), .ZN(n16746) );
  NAND2_X1 U16761 ( .A1(n16750), .A2(n16751), .ZN(n16608) );
  NAND2_X1 U16762 ( .A1(n16752), .A2(n16598), .ZN(n16751) );
  NAND2_X1 U16763 ( .A1(n16753), .A2(n16754), .ZN(n16598) );
  INV_X1 U16764 ( .A(n16755), .ZN(n16754) );
  NOR3_X1 U16765 ( .A1(n8551), .A2(n16756), .A3(n8590), .ZN(n16755) );
  NOR2_X1 U16766 ( .A1(n16596), .A2(n16597), .ZN(n16756) );
  NAND2_X1 U16767 ( .A1(n16597), .A2(n16596), .ZN(n16753) );
  NAND2_X1 U16768 ( .A1(n16757), .A2(n16758), .ZN(n16596) );
  NAND2_X1 U16769 ( .A1(n16759), .A2(n16587), .ZN(n16758) );
  NAND2_X1 U16770 ( .A1(n16760), .A2(n16761), .ZN(n16587) );
  NAND3_X1 U16771 ( .A1(n9107), .A2(n16762), .A3(n16285), .ZN(n16761) );
  INV_X1 U16772 ( .A(n16763), .ZN(n16762) );
  NOR2_X1 U16773 ( .A1(n16586), .A2(n16585), .ZN(n16763) );
  NAND2_X1 U16774 ( .A1(n16585), .A2(n16586), .ZN(n16760) );
  NAND2_X1 U16775 ( .A1(n16764), .A2(n16765), .ZN(n16586) );
  NAND2_X1 U16776 ( .A1(n16766), .A2(n16576), .ZN(n16765) );
  NAND2_X1 U16777 ( .A1(n16767), .A2(n16768), .ZN(n16576) );
  INV_X1 U16778 ( .A(n16769), .ZN(n16768) );
  NOR3_X1 U16779 ( .A1(n8535), .A2(n16770), .A3(n8590), .ZN(n16769) );
  NOR2_X1 U16780 ( .A1(n16574), .A2(n16575), .ZN(n16770) );
  NAND2_X1 U16781 ( .A1(n16575), .A2(n16574), .ZN(n16767) );
  NAND2_X1 U16782 ( .A1(n16771), .A2(n16772), .ZN(n16574) );
  NAND3_X1 U16783 ( .A1(n9373), .A2(n16773), .A3(n16285), .ZN(n16772) );
  INV_X1 U16784 ( .A(n16774), .ZN(n16773) );
  NOR2_X1 U16785 ( .A1(n16571), .A2(n16570), .ZN(n16774) );
  INV_X1 U16786 ( .A(n9126), .ZN(n9373) );
  NAND2_X1 U16787 ( .A1(n16570), .A2(n16571), .ZN(n16771) );
  NAND2_X1 U16788 ( .A1(n16564), .A2(n16775), .ZN(n16571) );
  NAND2_X1 U16789 ( .A1(n16776), .A2(n16563), .ZN(n16775) );
  NAND2_X1 U16790 ( .A1(n16777), .A2(n16778), .ZN(n16563) );
  NAND3_X1 U16791 ( .A1(n9138), .A2(n16779), .A3(n16285), .ZN(n16778) );
  INV_X1 U16792 ( .A(n16780), .ZN(n16779) );
  NOR2_X1 U16793 ( .A1(n16560), .A2(n16561), .ZN(n16780) );
  NAND2_X1 U16794 ( .A1(n16561), .A2(n16560), .ZN(n16777) );
  NAND2_X1 U16795 ( .A1(n16556), .A2(n16781), .ZN(n16560) );
  NAND3_X1 U16796 ( .A1(n8874), .A2(n8585), .A3(n16557), .ZN(n16781) );
  NOR2_X1 U16797 ( .A1(n8590), .A2(n9146), .ZN(n16557) );
  NAND3_X1 U16798 ( .A1(n8537), .A2(n8874), .A3(n16285), .ZN(n16556) );
  NOR2_X1 U16799 ( .A1(n8538), .A2(n16551), .ZN(n9149) );
  INV_X1 U16800 ( .A(n8627), .ZN(n16551) );
  XOR2_X1 U16801 ( .A(n16782), .B(n16783), .Z(n8627) );
  NOR2_X1 U16802 ( .A1(n16785), .A2(n16782), .ZN(n8632) );
  NOR2_X1 U16803 ( .A1(b_31_), .A2(a_31_), .ZN(n16785) );
  NOR2_X1 U16804 ( .A1(n9146), .A2(n16404), .ZN(n16561) );
  XNOR2_X1 U16805 ( .A(n16786), .B(n16787), .ZN(n9146) );
  XOR2_X1 U16806 ( .A(b_29_), .B(a_29_), .Z(n16787) );
  NAND2_X1 U16807 ( .A1(n8574), .A2(n16567), .ZN(n16776) );
  INV_X1 U16808 ( .A(n16788), .ZN(n16564) );
  NOR3_X1 U16809 ( .A1(n16284), .A2(n9378), .A3(n16567), .ZN(n16788) );
  NAND2_X1 U16810 ( .A1(n9138), .A2(n8874), .ZN(n16567) );
  INV_X1 U16811 ( .A(n9383), .ZN(n9138) );
  XOR2_X1 U16812 ( .A(n16789), .B(n16790), .Z(n9383) );
  XNOR2_X1 U16813 ( .A(a_28_), .B(b_28_), .ZN(n16789) );
  NOR2_X1 U16814 ( .A1(n9378), .A2(n16404), .ZN(n16570) );
  XNOR2_X1 U16815 ( .A(n16791), .B(n16792), .ZN(n9378) );
  XOR2_X1 U16816 ( .A(b_27_), .B(a_27_), .Z(n16792) );
  NOR2_X1 U16817 ( .A1(n9126), .A2(n16404), .ZN(n16575) );
  XNOR2_X1 U16818 ( .A(n16793), .B(n16794), .ZN(n9126) );
  XOR2_X1 U16819 ( .A(b_26_), .B(a_26_), .Z(n16794) );
  NAND2_X1 U16820 ( .A1(n8584), .A2(n16582), .ZN(n16766) );
  INV_X1 U16821 ( .A(n16579), .ZN(n16764) );
  NOR3_X1 U16822 ( .A1(n16284), .A2(n8584), .A3(n16582), .ZN(n16579) );
  NAND2_X1 U16823 ( .A1(n9121), .A2(n8874), .ZN(n16582) );
  INV_X1 U16824 ( .A(n8535), .ZN(n9121) );
  XOR2_X1 U16825 ( .A(b_25_), .B(a_25_), .Z(n16796) );
  NOR2_X1 U16826 ( .A1(n9176), .A2(n16404), .ZN(n16585) );
  XNOR2_X1 U16827 ( .A(n16797), .B(n16798), .ZN(n9176) );
  XOR2_X1 U16828 ( .A(b_24_), .B(a_24_), .Z(n16798) );
  NAND2_X1 U16829 ( .A1(n8563), .A2(n16593), .ZN(n16759) );
  INV_X1 U16830 ( .A(n16590), .ZN(n16757) );
  NOR3_X1 U16831 ( .A1(n16284), .A2(n8563), .A3(n16593), .ZN(n16590) );
  NAND2_X1 U16832 ( .A1(n9107), .A2(n8874), .ZN(n16593) );
  INV_X1 U16833 ( .A(n8548), .ZN(n9107) );
  XOR2_X1 U16834 ( .A(b_23_), .B(a_23_), .Z(n16800) );
  NOR2_X1 U16835 ( .A1(n9094), .A2(n16404), .ZN(n16597) );
  XNOR2_X1 U16836 ( .A(n16801), .B(n16802), .ZN(n9094) );
  XOR2_X1 U16837 ( .A(b_22_), .B(a_22_), .Z(n16802) );
  NAND2_X1 U16838 ( .A1(n8588), .A2(n16604), .ZN(n16752) );
  INV_X1 U16839 ( .A(n16601), .ZN(n16750) );
  NOR3_X1 U16840 ( .A1(n16284), .A2(n8588), .A3(n16604), .ZN(n16601) );
  NAND2_X1 U16841 ( .A1(n8515), .A2(n8874), .ZN(n16604) );
  XOR2_X1 U16842 ( .A(b_21_), .B(a_21_), .Z(n16804) );
  NOR2_X1 U16843 ( .A1(n9076), .A2(n16404), .ZN(n16607) );
  XNOR2_X1 U16844 ( .A(n16805), .B(n16806), .ZN(n9076) );
  XOR2_X1 U16845 ( .A(b_20_), .B(a_20_), .Z(n16806) );
  NAND2_X1 U16846 ( .A1(n8583), .A2(n16614), .ZN(n16745) );
  INV_X1 U16847 ( .A(n16807), .ZN(n16611) );
  NOR3_X1 U16848 ( .A1(n16284), .A2(n8583), .A3(n16614), .ZN(n16807) );
  NAND2_X1 U16849 ( .A1(n9070), .A2(n8874), .ZN(n16614) );
  INV_X1 U16850 ( .A(n9066), .ZN(n9070) );
  XNOR2_X1 U16851 ( .A(n16808), .B(n16809), .ZN(n9066) );
  XOR2_X1 U16852 ( .A(b_19_), .B(a_19_), .Z(n16809) );
  NOR2_X1 U16853 ( .A1(n9061), .A2(n16404), .ZN(n16617) );
  XNOR2_X1 U16854 ( .A(n16810), .B(n16811), .ZN(n9061) );
  XOR2_X1 U16855 ( .A(b_18_), .B(a_18_), .Z(n16811) );
  NAND2_X1 U16856 ( .A1(n8569), .A2(n16625), .ZN(n16739) );
  INV_X1 U16857 ( .A(n16622), .ZN(n16737) );
  NOR3_X1 U16858 ( .A1(n16284), .A2(n8569), .A3(n16625), .ZN(n16622) );
  NAND2_X1 U16859 ( .A1(n10722), .A2(n8874), .ZN(n16625) );
  INV_X1 U16860 ( .A(n9056), .ZN(n10722) );
  XNOR2_X1 U16861 ( .A(n16812), .B(n16813), .ZN(n9056) );
  XOR2_X1 U16862 ( .A(b_17_), .B(a_17_), .Z(n16813) );
  NOR2_X1 U16863 ( .A1(n9050), .A2(n16404), .ZN(n16628) );
  XNOR2_X1 U16864 ( .A(n16814), .B(n16815), .ZN(n9050) );
  XOR2_X1 U16865 ( .A(b_16_), .B(a_16_), .Z(n16815) );
  NAND2_X1 U16866 ( .A1(n8562), .A2(n16635), .ZN(n16732) );
  INV_X1 U16867 ( .A(n16816), .ZN(n16632) );
  NOR3_X1 U16868 ( .A1(n16284), .A2(n8562), .A3(n16635), .ZN(n16816) );
  NAND2_X1 U16869 ( .A1(n10222), .A2(n8874), .ZN(n16635) );
  INV_X1 U16870 ( .A(n8545), .ZN(n10222) );
  XOR2_X1 U16871 ( .A(b_15_), .B(a_15_), .Z(n16818) );
  NOR2_X1 U16872 ( .A1(n9041), .A2(n16404), .ZN(n16638) );
  XNOR2_X1 U16873 ( .A(n16819), .B(n16820), .ZN(n9041) );
  XOR2_X1 U16874 ( .A(b_14_), .B(a_14_), .Z(n16820) );
  NAND2_X1 U16875 ( .A1(n8582), .A2(n16646), .ZN(n16726) );
  INV_X1 U16876 ( .A(n16643), .ZN(n16724) );
  NOR3_X1 U16877 ( .A1(n16284), .A2(n8582), .A3(n16646), .ZN(n16643) );
  NAND2_X1 U16878 ( .A1(n9721), .A2(n8874), .ZN(n16646) );
  INV_X1 U16879 ( .A(n9036), .ZN(n9721) );
  XNOR2_X1 U16880 ( .A(n16821), .B(n16822), .ZN(n9036) );
  XOR2_X1 U16881 ( .A(b_13_), .B(a_13_), .Z(n16822) );
  NOR2_X1 U16882 ( .A1(n9031), .A2(n16404), .ZN(n16649) );
  XNOR2_X1 U16883 ( .A(n16823), .B(n16824), .ZN(n9031) );
  XOR2_X1 U16884 ( .A(b_12_), .B(a_12_), .Z(n16824) );
  NAND2_X1 U16885 ( .A1(n8556), .A2(n16656), .ZN(n16719) );
  INV_X1 U16886 ( .A(n16825), .ZN(n16653) );
  NOR3_X1 U16887 ( .A1(n9020), .A2(n8590), .A3(n16656), .ZN(n16825) );
  NAND2_X1 U16888 ( .A1(n9209), .A2(n8874), .ZN(n16656) );
  INV_X1 U16889 ( .A(n9025), .ZN(n9209) );
  XNOR2_X1 U16890 ( .A(n16826), .B(n16827), .ZN(n9025) );
  XOR2_X1 U16891 ( .A(b_11_), .B(a_11_), .Z(n16827) );
  NOR2_X1 U16892 ( .A1(n9020), .A2(n16404), .ZN(n16716) );
  XNOR2_X1 U16893 ( .A(n16828), .B(n16829), .ZN(n9020) );
  XOR2_X1 U16894 ( .A(b_10_), .B(a_10_), .Z(n16829) );
  NAND2_X1 U16895 ( .A1(n8560), .A2(n16830), .ZN(n16712) );
  NOR3_X1 U16896 ( .A1(n9010), .A2(n8590), .A3(n16830), .ZN(n16664) );
  INV_X1 U16897 ( .A(n16665), .ZN(n16830) );
  NOR2_X1 U16898 ( .A1(n9014), .A2(n16404), .ZN(n16665) );
  XNOR2_X1 U16899 ( .A(n16831), .B(n16832), .ZN(n9014) );
  XOR2_X1 U16900 ( .A(b_9_), .B(a_9_), .Z(n16832) );
  NAND2_X1 U16901 ( .A1(n9295), .A2(n8874), .ZN(n16670) );
  INV_X1 U16902 ( .A(n9010), .ZN(n9295) );
  XNOR2_X1 U16903 ( .A(n16833), .B(n16834), .ZN(n9010) );
  XOR2_X1 U16904 ( .A(b_8_), .B(a_8_), .Z(n16834) );
  NAND2_X1 U16905 ( .A1(n8555), .A2(n16676), .ZN(n16705) );
  INV_X1 U16906 ( .A(n16835), .ZN(n16673) );
  NOR3_X1 U16907 ( .A1(n9000), .A2(n8590), .A3(n16676), .ZN(n16835) );
  NAND2_X1 U16908 ( .A1(n8543), .A2(n8874), .ZN(n16676) );
  XNOR2_X1 U16909 ( .A(n16836), .B(n16837), .ZN(n9005) );
  XOR2_X1 U16910 ( .A(b_7_), .B(a_7_), .Z(n16837) );
  NOR2_X1 U16911 ( .A1(n9000), .A2(n16404), .ZN(n16702) );
  XNOR2_X1 U16912 ( .A(n16838), .B(n16839), .ZN(n9000) );
  XOR2_X1 U16913 ( .A(b_6_), .B(a_6_), .Z(n16839) );
  NAND2_X1 U16914 ( .A1(n8528), .A2(n16840), .ZN(n16698) );
  NOR3_X1 U16915 ( .A1(n8528), .A2(n8590), .A3(n16840), .ZN(n16684) );
  INV_X1 U16916 ( .A(n16685), .ZN(n16840) );
  NOR2_X1 U16917 ( .A1(n8995), .A2(n16404), .ZN(n16685) );
  INV_X1 U16918 ( .A(n8874), .ZN(n16404) );
  XNOR2_X1 U16919 ( .A(n16841), .B(n16842), .ZN(n8995) );
  XOR2_X1 U16920 ( .A(b_5_), .B(a_5_), .Z(n16842) );
  NAND2_X1 U16921 ( .A1(n9277), .A2(n8874), .ZN(n16690) );
  INV_X1 U16922 ( .A(n8528), .ZN(n9277) );
  XOR2_X1 U16923 ( .A(b_4_), .B(a_4_), .Z(n16844) );
  NAND2_X1 U16924 ( .A1(n16419), .A2(n16845), .ZN(n16691) );
  NAND2_X1 U16925 ( .A1(n16846), .A2(n16423), .ZN(n16845) );
  NAND2_X1 U16926 ( .A1(n9268), .A2(n16285), .ZN(n16846) );
  INV_X1 U16927 ( .A(n16847), .ZN(n16419) );
  NOR3_X1 U16928 ( .A1(n8982), .A2(n8590), .A3(n16423), .ZN(n16847) );
  NAND2_X1 U16929 ( .A1(n9792), .A2(n8874), .ZN(n16423) );
  XOR2_X1 U16930 ( .A(d_0_), .B(c_0_), .Z(n16849) );
  NAND2_X1 U16931 ( .A1(n16850), .A2(n16851), .ZN(n16848) );
  NAND2_X1 U16932 ( .A1(n16852), .A2(n16853), .ZN(n16851) );
  NAND2_X1 U16933 ( .A1(c_1_), .A2(n16854), .ZN(n16852) );
  INV_X1 U16934 ( .A(n16855), .ZN(n16850) );
  NOR2_X1 U16935 ( .A1(n16854), .A2(c_1_), .ZN(n16855) );
  INV_X1 U16936 ( .A(n8527), .ZN(n9792) );
  XOR2_X1 U16937 ( .A(b_3_), .B(a_3_), .Z(n16857) );
  XNOR2_X1 U16938 ( .A(n16854), .B(n16858), .ZN(n16284) );
  XNOR2_X1 U16939 ( .A(n16853), .B(c_1_), .ZN(n16858) );
  INV_X1 U16940 ( .A(d_1_), .ZN(n16853) );
  NAND2_X1 U16941 ( .A1(n16859), .A2(n16860), .ZN(n16854) );
  NAND2_X1 U16942 ( .A1(d_2_), .A2(n16861), .ZN(n16860) );
  INV_X1 U16943 ( .A(n16862), .ZN(n16861) );
  NOR2_X1 U16944 ( .A1(n16552), .A2(c_2_), .ZN(n16862) );
  NAND2_X1 U16945 ( .A1(c_2_), .A2(n16552), .ZN(n16859) );
  NAND2_X1 U16946 ( .A1(d_3_), .A2(n16865), .ZN(n16864) );
  INV_X1 U16947 ( .A(n16866), .ZN(n16865) );
  NOR2_X1 U16948 ( .A1(n16288), .A2(c_3_), .ZN(n16866) );
  NAND2_X1 U16949 ( .A1(c_3_), .A2(n16288), .ZN(n16863) );
  NAND2_X1 U16950 ( .A1(n16867), .A2(n16868), .ZN(n16288) );
  NAND2_X1 U16951 ( .A1(d_4_), .A2(n16869), .ZN(n16868) );
  INV_X1 U16952 ( .A(n16870), .ZN(n16869) );
  NOR2_X1 U16953 ( .A1(n16043), .A2(c_4_), .ZN(n16870) );
  NAND2_X1 U16954 ( .A1(c_4_), .A2(n16043), .ZN(n16867) );
  NAND2_X1 U16955 ( .A1(n16871), .A2(n16872), .ZN(n16043) );
  NAND2_X1 U16956 ( .A1(d_5_), .A2(n16873), .ZN(n16872) );
  INV_X1 U16957 ( .A(n16874), .ZN(n16873) );
  NOR2_X1 U16958 ( .A1(n15777), .A2(c_5_), .ZN(n16874) );
  NAND2_X1 U16959 ( .A1(c_5_), .A2(n15777), .ZN(n16871) );
  NAND2_X1 U16960 ( .A1(n16875), .A2(n16876), .ZN(n15777) );
  NAND2_X1 U16961 ( .A1(d_6_), .A2(n16877), .ZN(n16876) );
  INV_X1 U16962 ( .A(n16878), .ZN(n16877) );
  NOR2_X1 U16963 ( .A1(n15560), .A2(c_6_), .ZN(n16878) );
  NAND2_X1 U16964 ( .A1(c_6_), .A2(n15560), .ZN(n16875) );
  NAND2_X1 U16965 ( .A1(n16879), .A2(n16880), .ZN(n15560) );
  NAND2_X1 U16966 ( .A1(d_7_), .A2(n16881), .ZN(n16880) );
  INV_X1 U16967 ( .A(n16882), .ZN(n16881) );
  NOR2_X1 U16968 ( .A1(n15271), .A2(c_7_), .ZN(n16882) );
  NAND2_X1 U16969 ( .A1(c_7_), .A2(n15271), .ZN(n16879) );
  NAND2_X1 U16970 ( .A1(n16883), .A2(n16884), .ZN(n15271) );
  NAND2_X1 U16971 ( .A1(d_8_), .A2(n16885), .ZN(n16884) );
  INV_X1 U16972 ( .A(n16886), .ZN(n16885) );
  NOR2_X1 U16973 ( .A1(n15050), .A2(c_8_), .ZN(n16886) );
  NAND2_X1 U16974 ( .A1(c_8_), .A2(n15050), .ZN(n16883) );
  NAND2_X1 U16975 ( .A1(n16887), .A2(n16888), .ZN(n15050) );
  NAND2_X1 U16976 ( .A1(d_9_), .A2(n16889), .ZN(n16888) );
  INV_X1 U16977 ( .A(n16890), .ZN(n16889) );
  NOR2_X1 U16978 ( .A1(n14764), .A2(c_9_), .ZN(n16890) );
  NAND2_X1 U16979 ( .A1(c_9_), .A2(n14764), .ZN(n16887) );
  NAND2_X1 U16980 ( .A1(n16891), .A2(n16892), .ZN(n14764) );
  NAND2_X1 U16981 ( .A1(d_10_), .A2(n16893), .ZN(n16892) );
  INV_X1 U16982 ( .A(n16894), .ZN(n16893) );
  NOR2_X1 U16983 ( .A1(n14546), .A2(c_10_), .ZN(n16894) );
  NAND2_X1 U16984 ( .A1(c_10_), .A2(n14546), .ZN(n16891) );
  NAND2_X1 U16985 ( .A1(n16895), .A2(n16896), .ZN(n14546) );
  NAND2_X1 U16986 ( .A1(d_11_), .A2(n16897), .ZN(n16896) );
  INV_X1 U16987 ( .A(n16898), .ZN(n16897) );
  NOR2_X1 U16988 ( .A1(n14251), .A2(c_11_), .ZN(n16898) );
  NAND2_X1 U16989 ( .A1(c_11_), .A2(n14251), .ZN(n16895) );
  NAND2_X1 U16990 ( .A1(n16899), .A2(n16900), .ZN(n14251) );
  NAND2_X1 U16991 ( .A1(d_12_), .A2(n16901), .ZN(n16900) );
  INV_X1 U16992 ( .A(n16902), .ZN(n16901) );
  NOR2_X1 U16993 ( .A1(n14034), .A2(c_12_), .ZN(n16902) );
  NAND2_X1 U16994 ( .A1(c_12_), .A2(n14034), .ZN(n16899) );
  NAND2_X1 U16995 ( .A1(n16903), .A2(n16904), .ZN(n14034) );
  NAND2_X1 U16996 ( .A1(d_13_), .A2(n16905), .ZN(n16904) );
  INV_X1 U16997 ( .A(n16906), .ZN(n16905) );
  NOR2_X1 U16998 ( .A1(n13742), .A2(c_13_), .ZN(n16906) );
  NAND2_X1 U16999 ( .A1(c_13_), .A2(n13742), .ZN(n16903) );
  NAND2_X1 U17000 ( .A1(n16907), .A2(n16908), .ZN(n13742) );
  NAND2_X1 U17001 ( .A1(d_14_), .A2(n16909), .ZN(n16908) );
  INV_X1 U17002 ( .A(n16910), .ZN(n16909) );
  NOR2_X1 U17003 ( .A1(n13507), .A2(c_14_), .ZN(n16910) );
  NAND2_X1 U17004 ( .A1(c_14_), .A2(n13507), .ZN(n16907) );
  NAND2_X1 U17005 ( .A1(n16911), .A2(n16912), .ZN(n13507) );
  NAND2_X1 U17006 ( .A1(d_15_), .A2(n16913), .ZN(n16912) );
  INV_X1 U17007 ( .A(n16914), .ZN(n16913) );
  NOR2_X1 U17008 ( .A1(n13223), .A2(c_15_), .ZN(n16914) );
  NAND2_X1 U17009 ( .A1(c_15_), .A2(n13223), .ZN(n16911) );
  NAND2_X1 U17010 ( .A1(n16915), .A2(n16916), .ZN(n13223) );
  NAND2_X1 U17011 ( .A1(d_16_), .A2(n16917), .ZN(n16916) );
  INV_X1 U17012 ( .A(n16918), .ZN(n16917) );
  NOR2_X1 U17013 ( .A1(n12984), .A2(c_16_), .ZN(n16918) );
  NAND2_X1 U17014 ( .A1(c_16_), .A2(n12984), .ZN(n16915) );
  NAND2_X1 U17015 ( .A1(d_17_), .A2(n16921), .ZN(n16920) );
  INV_X1 U17016 ( .A(n16922), .ZN(n16921) );
  NOR2_X1 U17017 ( .A1(n12731), .A2(c_17_), .ZN(n16922) );
  NAND2_X1 U17018 ( .A1(c_17_), .A2(n12731), .ZN(n16919) );
  NAND2_X1 U17019 ( .A1(d_18_), .A2(n16925), .ZN(n16924) );
  INV_X1 U17020 ( .A(n16926), .ZN(n16925) );
  NOR2_X1 U17021 ( .A1(n12460), .A2(c_18_), .ZN(n16926) );
  NAND2_X1 U17022 ( .A1(c_18_), .A2(n12460), .ZN(n16923) );
  NAND2_X1 U17023 ( .A1(d_19_), .A2(n16929), .ZN(n16928) );
  INV_X1 U17024 ( .A(n16930), .ZN(n16929) );
  NOR2_X1 U17025 ( .A1(n12199), .A2(c_19_), .ZN(n16930) );
  NAND2_X1 U17026 ( .A1(c_19_), .A2(n12199), .ZN(n16927) );
  NAND2_X1 U17027 ( .A1(n16931), .A2(n16932), .ZN(n12199) );
  NAND2_X1 U17028 ( .A1(d_20_), .A2(n16933), .ZN(n16932) );
  INV_X1 U17029 ( .A(n16934), .ZN(n16933) );
  NOR2_X1 U17030 ( .A1(n11939), .A2(c_20_), .ZN(n16934) );
  NAND2_X1 U17031 ( .A1(c_20_), .A2(n11939), .ZN(n16931) );
  NAND2_X1 U17032 ( .A1(d_21_), .A2(n16937), .ZN(n16936) );
  INV_X1 U17033 ( .A(n16938), .ZN(n16937) );
  NOR2_X1 U17034 ( .A1(n11689), .A2(c_21_), .ZN(n16938) );
  NAND2_X1 U17035 ( .A1(c_21_), .A2(n11689), .ZN(n16935) );
  NAND2_X1 U17036 ( .A1(n16939), .A2(n16940), .ZN(n11689) );
  NAND2_X1 U17037 ( .A1(d_22_), .A2(n16941), .ZN(n16940) );
  INV_X1 U17038 ( .A(n16942), .ZN(n16941) );
  NOR2_X1 U17039 ( .A1(n11435), .A2(c_22_), .ZN(n16942) );
  NAND2_X1 U17040 ( .A1(c_22_), .A2(n11435), .ZN(n16939) );
  NAND2_X1 U17041 ( .A1(n16943), .A2(n16944), .ZN(n11435) );
  NAND2_X1 U17042 ( .A1(d_23_), .A2(n16945), .ZN(n16944) );
  INV_X1 U17043 ( .A(n16946), .ZN(n16945) );
  NOR2_X1 U17044 ( .A1(n11185), .A2(c_23_), .ZN(n16946) );
  NAND2_X1 U17045 ( .A1(c_23_), .A2(n11185), .ZN(n16943) );
  NAND2_X1 U17046 ( .A1(d_24_), .A2(n16949), .ZN(n16948) );
  INV_X1 U17047 ( .A(n16950), .ZN(n16949) );
  NOR2_X1 U17048 ( .A1(n11048), .A2(c_24_), .ZN(n16950) );
  NAND2_X1 U17049 ( .A1(c_24_), .A2(n11048), .ZN(n16947) );
  NAND2_X1 U17050 ( .A1(n16951), .A2(n16952), .ZN(n11048) );
  NAND2_X1 U17051 ( .A1(d_25_), .A2(n16953), .ZN(n16952) );
  INV_X1 U17052 ( .A(n16954), .ZN(n16953) );
  NOR2_X1 U17053 ( .A1(n10764), .A2(c_25_), .ZN(n16954) );
  NAND2_X1 U17054 ( .A1(c_25_), .A2(n10764), .ZN(n16951) );
  NAND2_X1 U17055 ( .A1(n16955), .A2(n16956), .ZN(n10764) );
  NAND2_X1 U17056 ( .A1(d_26_), .A2(n16957), .ZN(n16956) );
  INV_X1 U17057 ( .A(n16958), .ZN(n16957) );
  NOR2_X1 U17058 ( .A1(n10505), .A2(c_26_), .ZN(n16958) );
  NAND2_X1 U17059 ( .A1(c_26_), .A2(n10505), .ZN(n16955) );
  NAND2_X1 U17060 ( .A1(n16959), .A2(n16960), .ZN(n10505) );
  NAND2_X1 U17061 ( .A1(d_27_), .A2(n16961), .ZN(n16960) );
  INV_X1 U17062 ( .A(n16962), .ZN(n16961) );
  NOR2_X1 U17063 ( .A1(n10256), .A2(c_27_), .ZN(n16962) );
  NAND2_X1 U17064 ( .A1(c_27_), .A2(n10256), .ZN(n16959) );
  NAND2_X1 U17065 ( .A1(d_28_), .A2(n16965), .ZN(n16964) );
  INV_X1 U17066 ( .A(n16966), .ZN(n16965) );
  NOR2_X1 U17067 ( .A1(n9907), .A2(c_28_), .ZN(n16966) );
  NAND2_X1 U17068 ( .A1(c_28_), .A2(n9907), .ZN(n16963) );
  NAND2_X1 U17069 ( .A1(n16967), .A2(n16968), .ZN(n9907) );
  NAND2_X1 U17070 ( .A1(d_29_), .A2(n16969), .ZN(n16968) );
  INV_X1 U17071 ( .A(n16970), .ZN(n16969) );
  NOR2_X1 U17072 ( .A1(n9762), .A2(c_29_), .ZN(n16970) );
  NAND2_X1 U17073 ( .A1(c_29_), .A2(n9762), .ZN(n16967) );
  NAND2_X1 U17074 ( .A1(n16971), .A2(n16972), .ZN(n9762) );
  NAND2_X1 U17075 ( .A1(d_30_), .A2(n16973), .ZN(n16972) );
  INV_X1 U17076 ( .A(n16974), .ZN(n16973) );
  NOR2_X1 U17077 ( .A1(c_30_), .A2(n9151), .ZN(n16974) );
  NAND2_X1 U17078 ( .A1(c_30_), .A2(n9151), .ZN(n16971) );
  INV_X1 U17079 ( .A(n9396), .ZN(n9151) );
  NAND2_X1 U17080 ( .A1(d_31_), .A2(c_31_), .ZN(n9396) );
  XOR2_X1 U17081 ( .A(b_2_), .B(a_2_), .Z(n16976) );
  XNOR2_X1 U17082 ( .A(n16977), .B(n16978), .ZN(n8872) );
  XOR2_X1 U17083 ( .A(b_0_), .B(a_0_), .Z(n16978) );
  NAND2_X1 U17084 ( .A1(n16979), .A2(n16980), .ZN(n16977) );
  NAND2_X1 U17085 ( .A1(n16981), .A2(n16430), .ZN(n16980) );
  INV_X1 U17086 ( .A(b_1_), .ZN(n16430) );
  NAND2_X1 U17087 ( .A1(a_1_), .A2(n16428), .ZN(n16981) );
  INV_X1 U17088 ( .A(n16982), .ZN(n16979) );
  NOR2_X1 U17089 ( .A1(n16428), .A2(a_1_), .ZN(n16982) );
  NAND2_X1 U17090 ( .A1(b_2_), .A2(n16985), .ZN(n16984) );
  INV_X1 U17091 ( .A(n16986), .ZN(n16985) );
  NOR2_X1 U17092 ( .A1(n16975), .A2(a_2_), .ZN(n16986) );
  NAND2_X1 U17093 ( .A1(a_2_), .A2(n16975), .ZN(n16983) );
  NAND2_X1 U17094 ( .A1(n16987), .A2(n16988), .ZN(n16975) );
  NAND2_X1 U17095 ( .A1(b_3_), .A2(n16989), .ZN(n16988) );
  INV_X1 U17096 ( .A(n16990), .ZN(n16989) );
  NOR2_X1 U17097 ( .A1(n16856), .A2(a_3_), .ZN(n16990) );
  NAND2_X1 U17098 ( .A1(a_3_), .A2(n16856), .ZN(n16987) );
  NAND2_X1 U17099 ( .A1(n16991), .A2(n16992), .ZN(n16856) );
  NAND2_X1 U17100 ( .A1(b_4_), .A2(n16993), .ZN(n16992) );
  INV_X1 U17101 ( .A(n16994), .ZN(n16993) );
  NOR2_X1 U17102 ( .A1(n16843), .A2(a_4_), .ZN(n16994) );
  NAND2_X1 U17103 ( .A1(a_4_), .A2(n16843), .ZN(n16991) );
  NAND2_X1 U17104 ( .A1(n16995), .A2(n16996), .ZN(n16843) );
  NAND2_X1 U17105 ( .A1(b_5_), .A2(n16997), .ZN(n16996) );
  INV_X1 U17106 ( .A(n16998), .ZN(n16997) );
  NOR2_X1 U17107 ( .A1(n16841), .A2(a_5_), .ZN(n16998) );
  NAND2_X1 U17108 ( .A1(a_5_), .A2(n16841), .ZN(n16995) );
  NAND2_X1 U17109 ( .A1(n16999), .A2(n17000), .ZN(n16841) );
  NAND2_X1 U17110 ( .A1(b_6_), .A2(n17001), .ZN(n17000) );
  INV_X1 U17111 ( .A(n17002), .ZN(n17001) );
  NOR2_X1 U17112 ( .A1(n16838), .A2(a_6_), .ZN(n17002) );
  NAND2_X1 U17113 ( .A1(a_6_), .A2(n16838), .ZN(n16999) );
  NAND2_X1 U17114 ( .A1(n17003), .A2(n17004), .ZN(n16838) );
  NAND2_X1 U17115 ( .A1(b_7_), .A2(n17005), .ZN(n17004) );
  INV_X1 U17116 ( .A(n17006), .ZN(n17005) );
  NOR2_X1 U17117 ( .A1(n16836), .A2(a_7_), .ZN(n17006) );
  NAND2_X1 U17118 ( .A1(a_7_), .A2(n16836), .ZN(n17003) );
  NAND2_X1 U17119 ( .A1(n17007), .A2(n17008), .ZN(n16836) );
  NAND2_X1 U17120 ( .A1(b_8_), .A2(n17009), .ZN(n17008) );
  INV_X1 U17121 ( .A(n17010), .ZN(n17009) );
  NOR2_X1 U17122 ( .A1(n16833), .A2(a_8_), .ZN(n17010) );
  NAND2_X1 U17123 ( .A1(a_8_), .A2(n16833), .ZN(n17007) );
  NAND2_X1 U17124 ( .A1(n17011), .A2(n17012), .ZN(n16833) );
  NAND2_X1 U17125 ( .A1(b_9_), .A2(n17013), .ZN(n17012) );
  INV_X1 U17126 ( .A(n17014), .ZN(n17013) );
  NOR2_X1 U17127 ( .A1(n16831), .A2(a_9_), .ZN(n17014) );
  NAND2_X1 U17128 ( .A1(a_9_), .A2(n16831), .ZN(n17011) );
  NAND2_X1 U17129 ( .A1(b_10_), .A2(n17017), .ZN(n17016) );
  INV_X1 U17130 ( .A(n17018), .ZN(n17017) );
  NOR2_X1 U17131 ( .A1(n16828), .A2(a_10_), .ZN(n17018) );
  NAND2_X1 U17132 ( .A1(a_10_), .A2(n16828), .ZN(n17015) );
  NAND2_X1 U17133 ( .A1(n17019), .A2(n17020), .ZN(n16828) );
  NAND2_X1 U17134 ( .A1(b_11_), .A2(n17021), .ZN(n17020) );
  INV_X1 U17135 ( .A(n17022), .ZN(n17021) );
  NOR2_X1 U17136 ( .A1(n16826), .A2(a_11_), .ZN(n17022) );
  NAND2_X1 U17137 ( .A1(a_11_), .A2(n16826), .ZN(n17019) );
  NAND2_X1 U17138 ( .A1(n17023), .A2(n17024), .ZN(n16826) );
  NAND2_X1 U17139 ( .A1(b_12_), .A2(n17025), .ZN(n17024) );
  INV_X1 U17140 ( .A(n17026), .ZN(n17025) );
  NOR2_X1 U17141 ( .A1(n16823), .A2(a_12_), .ZN(n17026) );
  NAND2_X1 U17142 ( .A1(a_12_), .A2(n16823), .ZN(n17023) );
  NAND2_X1 U17143 ( .A1(b_13_), .A2(n17029), .ZN(n17028) );
  INV_X1 U17144 ( .A(n17030), .ZN(n17029) );
  NOR2_X1 U17145 ( .A1(n16821), .A2(a_13_), .ZN(n17030) );
  NAND2_X1 U17146 ( .A1(a_13_), .A2(n16821), .ZN(n17027) );
  NAND2_X1 U17147 ( .A1(b_14_), .A2(n17033), .ZN(n17032) );
  INV_X1 U17148 ( .A(n17034), .ZN(n17033) );
  NOR2_X1 U17149 ( .A1(n16819), .A2(a_14_), .ZN(n17034) );
  NAND2_X1 U17150 ( .A1(a_14_), .A2(n16819), .ZN(n17031) );
  NAND2_X1 U17151 ( .A1(n17035), .A2(n17036), .ZN(n16819) );
  NAND2_X1 U17152 ( .A1(b_15_), .A2(n17037), .ZN(n17036) );
  INV_X1 U17153 ( .A(n17038), .ZN(n17037) );
  NOR2_X1 U17154 ( .A1(n16817), .A2(a_15_), .ZN(n17038) );
  NAND2_X1 U17155 ( .A1(a_15_), .A2(n16817), .ZN(n17035) );
  NAND2_X1 U17156 ( .A1(n17039), .A2(n17040), .ZN(n16817) );
  NAND2_X1 U17157 ( .A1(b_16_), .A2(n17041), .ZN(n17040) );
  INV_X1 U17158 ( .A(n17042), .ZN(n17041) );
  NOR2_X1 U17159 ( .A1(n16814), .A2(a_16_), .ZN(n17042) );
  NAND2_X1 U17160 ( .A1(a_16_), .A2(n16814), .ZN(n17039) );
  NAND2_X1 U17161 ( .A1(n17043), .A2(n17044), .ZN(n16814) );
  NAND2_X1 U17162 ( .A1(b_17_), .A2(n17045), .ZN(n17044) );
  INV_X1 U17163 ( .A(n17046), .ZN(n17045) );
  NOR2_X1 U17164 ( .A1(n16812), .A2(a_17_), .ZN(n17046) );
  NAND2_X1 U17165 ( .A1(a_17_), .A2(n16812), .ZN(n17043) );
  NAND2_X1 U17166 ( .A1(b_18_), .A2(n17049), .ZN(n17048) );
  INV_X1 U17167 ( .A(n17050), .ZN(n17049) );
  NOR2_X1 U17168 ( .A1(n16810), .A2(a_18_), .ZN(n17050) );
  NAND2_X1 U17169 ( .A1(a_18_), .A2(n16810), .ZN(n17047) );
  NAND2_X1 U17170 ( .A1(b_19_), .A2(n17053), .ZN(n17052) );
  INV_X1 U17171 ( .A(n17054), .ZN(n17053) );
  NOR2_X1 U17172 ( .A1(n16808), .A2(a_19_), .ZN(n17054) );
  NAND2_X1 U17173 ( .A1(a_19_), .A2(n16808), .ZN(n17051) );
  NAND2_X1 U17174 ( .A1(b_20_), .A2(n17057), .ZN(n17056) );
  INV_X1 U17175 ( .A(n17058), .ZN(n17057) );
  NOR2_X1 U17176 ( .A1(n16805), .A2(a_20_), .ZN(n17058) );
  NAND2_X1 U17177 ( .A1(a_20_), .A2(n16805), .ZN(n17055) );
  NAND2_X1 U17178 ( .A1(b_21_), .A2(n17061), .ZN(n17060) );
  INV_X1 U17179 ( .A(n17062), .ZN(n17061) );
  NOR2_X1 U17180 ( .A1(n16803), .A2(a_21_), .ZN(n17062) );
  NAND2_X1 U17181 ( .A1(a_21_), .A2(n16803), .ZN(n17059) );
  NAND2_X1 U17182 ( .A1(n17063), .A2(n17064), .ZN(n16803) );
  NAND2_X1 U17183 ( .A1(b_22_), .A2(n17065), .ZN(n17064) );
  INV_X1 U17184 ( .A(n17066), .ZN(n17065) );
  NOR2_X1 U17185 ( .A1(n16801), .A2(a_22_), .ZN(n17066) );
  NAND2_X1 U17186 ( .A1(a_22_), .A2(n16801), .ZN(n17063) );
  NAND2_X1 U17187 ( .A1(n17067), .A2(n17068), .ZN(n16801) );
  NAND2_X1 U17188 ( .A1(b_23_), .A2(n17069), .ZN(n17068) );
  INV_X1 U17189 ( .A(n17070), .ZN(n17069) );
  NOR2_X1 U17190 ( .A1(n16799), .A2(a_23_), .ZN(n17070) );
  NAND2_X1 U17191 ( .A1(a_23_), .A2(n16799), .ZN(n17067) );
  NAND2_X1 U17192 ( .A1(n17071), .A2(n17072), .ZN(n16799) );
  NAND2_X1 U17193 ( .A1(b_24_), .A2(n17073), .ZN(n17072) );
  INV_X1 U17194 ( .A(n17074), .ZN(n17073) );
  NOR2_X1 U17195 ( .A1(n16797), .A2(a_24_), .ZN(n17074) );
  NAND2_X1 U17196 ( .A1(a_24_), .A2(n16797), .ZN(n17071) );
  NAND2_X1 U17197 ( .A1(b_25_), .A2(n17077), .ZN(n17076) );
  INV_X1 U17198 ( .A(n17078), .ZN(n17077) );
  NOR2_X1 U17199 ( .A1(n16795), .A2(a_25_), .ZN(n17078) );
  NAND2_X1 U17200 ( .A1(a_25_), .A2(n16795), .ZN(n17075) );
  NAND2_X1 U17201 ( .A1(n17079), .A2(n17080), .ZN(n16795) );
  NAND2_X1 U17202 ( .A1(b_26_), .A2(n17081), .ZN(n17080) );
  INV_X1 U17203 ( .A(n17082), .ZN(n17081) );
  NOR2_X1 U17204 ( .A1(n16793), .A2(a_26_), .ZN(n17082) );
  NAND2_X1 U17205 ( .A1(a_26_), .A2(n16793), .ZN(n17079) );
  NAND2_X1 U17206 ( .A1(n17083), .A2(n17084), .ZN(n16793) );
  NAND2_X1 U17207 ( .A1(b_27_), .A2(n17085), .ZN(n17084) );
  INV_X1 U17208 ( .A(n17086), .ZN(n17085) );
  NOR2_X1 U17209 ( .A1(n16791), .A2(a_27_), .ZN(n17086) );
  NAND2_X1 U17210 ( .A1(a_27_), .A2(n16791), .ZN(n17083) );
  NAND2_X1 U17211 ( .A1(b_28_), .A2(n17089), .ZN(n17088) );
  INV_X1 U17212 ( .A(n17090), .ZN(n17089) );
  NOR2_X1 U17213 ( .A1(n16790), .A2(a_28_), .ZN(n17090) );
  NAND2_X1 U17214 ( .A1(a_28_), .A2(n16790), .ZN(n17087) );
  NAND2_X1 U17215 ( .A1(n17091), .A2(n17092), .ZN(n16790) );
  NAND2_X1 U17216 ( .A1(b_29_), .A2(n17093), .ZN(n17092) );
  INV_X1 U17217 ( .A(n17094), .ZN(n17093) );
  NOR2_X1 U17218 ( .A1(n16786), .A2(a_29_), .ZN(n17094) );
  NAND2_X1 U17219 ( .A1(a_29_), .A2(n16786), .ZN(n17091) );
  NAND2_X1 U17220 ( .A1(n17095), .A2(n17096), .ZN(n16786) );
  NAND2_X1 U17221 ( .A1(b_30_), .A2(n17097), .ZN(n17096) );
  NAND2_X1 U17222 ( .A1(n16784), .A2(n17098), .ZN(n17097) );
  INV_X1 U17223 ( .A(a_30_), .ZN(n16784) );
  NAND2_X1 U17224 ( .A1(a_30_), .A2(n16782), .ZN(n17095) );
  INV_X1 U17225 ( .A(n17098), .ZN(n16782) );
  NAND2_X1 U17226 ( .A1(b_31_), .A2(a_31_), .ZN(n17098) );
endmodule

