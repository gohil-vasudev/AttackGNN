module locked_c1355 (  G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,  G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT  );
  input  G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n311_, new_n313_, new_n314_, new_n316_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n328_, new_n330_, new_n331_, new_n333_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n342_, new_n344_, new_n346_, new_n347_, new_n349_, new_n350_, new_n352_, new_n354_, new_n356_, new_n357_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n392_, new_n393_, new_n395_, new_n396_, new_n398_, new_n399_, new_n401_, new_n402_, new_n404_, new_n405_, new_n406_, new_n408_, new_n410_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n437_, new_n438_, new_n439_, new_n440_, new_n442_, new_n444_, new_n445_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n453_, new_n454_, new_n456_, new_n458_, new_n459_;
  INV_X1 g000 ( .A(G1GAT), .ZN(new_n138_) );
  XNOR2_X1 g001 ( .A(G120GAT), .B(G127GAT), .ZN(new_n139_) );
  XNOR2_X1 g002 ( .A(G113GAT), .B(KEYINPUT0), .ZN(new_n140_) );
  XNOR2_X1 g003 ( .A(new_n139_), .B(new_n140_), .ZN(new_n141_) );
  XNOR2_X1 g004 ( .A(new_n141_), .B(new_n138_), .ZN(new_n142_) );
  XNOR2_X1 g005 ( .A(G155GAT), .B(KEYINPUT3), .ZN(new_n143_) );
  XNOR2_X1 g006 ( .A(G141GAT), .B(KEYINPUT2), .ZN(new_n144_) );
  XNOR2_X1 g007 ( .A(new_n143_), .B(new_n144_), .ZN(new_n145_) );
  XNOR2_X1 g008 ( .A(G57GAT), .B(KEYINPUT1), .ZN(new_n146_) );
  AND2_X1 g009 ( .A1(G225GAT), .A2(G233GAT), .ZN(new_n147_) );
  XNOR2_X1 g010 ( .A(new_n146_), .B(new_n147_), .ZN(new_n148_) );
  XOR2_X1 g011 ( .A(new_n145_), .B(new_n148_), .Z(new_n149_) );
  XNOR2_X1 g012 ( .A(new_n149_), .B(new_n142_), .ZN(new_n150_) );
  XOR2_X1 g013 ( .A(G29GAT), .B(G134GAT), .Z(new_n151_) );
  XOR2_X1 g014 ( .A(new_n150_), .B(new_n151_), .Z(new_n152_) );
  XNOR2_X1 g015 ( .A(G85GAT), .B(G162GAT), .ZN(new_n153_) );
  XNOR2_X1 g016 ( .A(new_n152_), .B(new_n153_), .ZN(new_n154_) );
  XOR2_X1 g017 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(new_n155_) );
  XNOR2_X1 g018 ( .A(G148GAT), .B(KEYINPUT6), .ZN(new_n156_) );
  XNOR2_X1 g019 ( .A(new_n155_), .B(new_n156_), .ZN(new_n157_) );
  XOR2_X1 g020 ( .A(new_n154_), .B(new_n157_), .Z(new_n158_) );
  INV_X1 g021 ( .A(new_n158_), .ZN(new_n159_) );
  XNOR2_X1 g022 ( .A(G211GAT), .B(G218GAT), .ZN(new_n160_) );
  XNOR2_X1 g023 ( .A(G204GAT), .B(KEYINPUT21), .ZN(new_n161_) );
  XOR2_X1 g024 ( .A(new_n160_), .B(new_n161_), .Z(new_n162_) );
  XNOR2_X1 g025 ( .A(new_n162_), .B(G197GAT), .ZN(new_n163_) );
  XOR2_X1 g026 ( .A(new_n163_), .B(new_n145_), .Z(new_n164_) );
  XNOR2_X1 g027 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(new_n165_) );
  XNOR2_X1 g028 ( .A(G22GAT), .B(KEYINPUT22), .ZN(new_n166_) );
  XNOR2_X1 g029 ( .A(new_n165_), .B(new_n166_), .ZN(new_n167_) );
  INV_X1 g030 ( .A(G148GAT), .ZN(new_n168_) );
  XOR2_X1 g031 ( .A(G78GAT), .B(G106GAT), .Z(new_n169_) );
  OR2_X1 g032 ( .A1(new_n169_), .A2(new_n168_), .ZN(new_n170_) );
  INV_X1 g033 ( .A(G78GAT), .ZN(new_n171_) );
  INV_X1 g034 ( .A(G106GAT), .ZN(new_n172_) );
  AND2_X1 g035 ( .A1(new_n171_), .A2(new_n172_), .ZN(new_n173_) );
  AND2_X1 g036 ( .A1(G78GAT), .A2(G106GAT), .ZN(new_n174_) );
  OR2_X1 g037 ( .A1(new_n174_), .A2(G148GAT), .ZN(new_n175_) );
  OR2_X1 g038 ( .A1(new_n175_), .A2(new_n173_), .ZN(new_n176_) );
  AND2_X1 g039 ( .A1(new_n176_), .A2(new_n170_), .ZN(new_n177_) );
  XOR2_X1 g040 ( .A(new_n177_), .B(new_n167_), .Z(new_n178_) );
  XNOR2_X1 g041 ( .A(new_n164_), .B(new_n178_), .ZN(new_n179_) );
  XOR2_X1 g042 ( .A(G50GAT), .B(G162GAT), .Z(new_n180_) );
  INV_X1 g043 ( .A(new_n180_), .ZN(new_n181_) );
  XNOR2_X1 g044 ( .A(new_n179_), .B(new_n181_), .ZN(new_n182_) );
  AND2_X1 g045 ( .A1(G228GAT), .A2(G233GAT), .ZN(new_n183_) );
  XNOR2_X1 g046 ( .A(new_n182_), .B(new_n183_), .ZN(new_n184_) );
  XNOR2_X1 g047 ( .A(new_n141_), .B(G15GAT), .ZN(new_n185_) );
  AND2_X1 g048 ( .A1(G227GAT), .A2(G233GAT), .ZN(new_n186_) );
  XOR2_X1 g049 ( .A(new_n185_), .B(new_n186_), .Z(new_n187_) );
  XNOR2_X1 g050 ( .A(G176GAT), .B(G183GAT), .ZN(new_n188_) );
  XNOR2_X1 g051 ( .A(G71GAT), .B(KEYINPUT20), .ZN(new_n189_) );
  XOR2_X1 g052 ( .A(new_n188_), .B(new_n189_), .Z(new_n190_) );
  XNOR2_X1 g053 ( .A(new_n187_), .B(new_n190_), .ZN(new_n191_) );
  XNOR2_X1 g054 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(new_n192_) );
  XNOR2_X1 g055 ( .A(G169GAT), .B(KEYINPUT19), .ZN(new_n193_) );
  XNOR2_X1 g056 ( .A(new_n192_), .B(new_n193_), .ZN(new_n194_) );
  XOR2_X1 g057 ( .A(G134GAT), .B(G190GAT), .Z(new_n195_) );
  XNOR2_X1 g058 ( .A(G43GAT), .B(G99GAT), .ZN(new_n196_) );
  XNOR2_X1 g059 ( .A(new_n195_), .B(new_n196_), .ZN(new_n197_) );
  XNOR2_X1 g060 ( .A(new_n197_), .B(new_n194_), .ZN(new_n198_) );
  XOR2_X1 g061 ( .A(new_n191_), .B(new_n198_), .Z(new_n199_) );
  OR2_X1 g062 ( .A1(new_n184_), .A2(new_n199_), .ZN(new_n200_) );
  XOR2_X1 g063 ( .A(new_n200_), .B(KEYINPUT26), .Z(new_n201_) );
  XNOR2_X1 g064 ( .A(G36GAT), .B(G190GAT), .ZN(new_n202_) );
  INV_X1 g065 ( .A(new_n202_), .ZN(new_n203_) );
  XNOR2_X1 g066 ( .A(new_n163_), .B(new_n203_), .ZN(new_n204_) );
  INV_X1 g067 ( .A(G92GAT), .ZN(new_n205_) );
  XNOR2_X1 g068 ( .A(G64GAT), .B(G176GAT), .ZN(new_n206_) );
  XNOR2_X1 g069 ( .A(new_n206_), .B(new_n205_), .ZN(new_n207_) );
  AND2_X1 g070 ( .A1(G226GAT), .A2(G233GAT), .ZN(new_n208_) );
  XNOR2_X1 g071 ( .A(new_n207_), .B(new_n208_), .ZN(new_n209_) );
  XNOR2_X1 g072 ( .A(G8GAT), .B(G183GAT), .ZN(new_n210_) );
  XNOR2_X1 g073 ( .A(new_n209_), .B(new_n210_), .ZN(new_n211_) );
  XNOR2_X1 g074 ( .A(new_n204_), .B(new_n211_), .ZN(new_n212_) );
  XNOR2_X1 g075 ( .A(new_n212_), .B(new_n194_), .ZN(new_n213_) );
  XNOR2_X1 g076 ( .A(new_n213_), .B(KEYINPUT27), .ZN(new_n214_) );
  AND2_X1 g077 ( .A1(new_n201_), .A2(new_n214_), .ZN(new_n215_) );
  INV_X1 g078 ( .A(new_n199_), .ZN(new_n216_) );
  INV_X1 g079 ( .A(new_n213_), .ZN(new_n217_) );
  OR2_X1 g080 ( .A1(new_n216_), .A2(new_n217_), .ZN(new_n218_) );
  AND2_X1 g081 ( .A1(new_n184_), .A2(new_n218_), .ZN(new_n219_) );
  XOR2_X1 g082 ( .A(new_n219_), .B(KEYINPUT25), .Z(new_n220_) );
  OR2_X1 g083 ( .A1(new_n215_), .A2(new_n220_), .ZN(new_n221_) );
  AND2_X1 g084 ( .A1(new_n221_), .A2(new_n158_), .ZN(new_n222_) );
  XOR2_X1 g085 ( .A(new_n184_), .B(KEYINPUT28), .Z(new_n223_) );
  INV_X1 g086 ( .A(new_n223_), .ZN(new_n224_) );
  AND2_X1 g087 ( .A1(new_n159_), .A2(new_n214_), .ZN(new_n225_) );
  AND2_X1 g088 ( .A1(new_n225_), .A2(new_n216_), .ZN(new_n226_) );
  AND2_X1 g089 ( .A1(new_n226_), .A2(new_n224_), .ZN(new_n227_) );
  OR2_X1 g090 ( .A1(new_n222_), .A2(new_n227_), .ZN(new_n228_) );
  XNOR2_X1 g091 ( .A(G106GAT), .B(G218GAT), .ZN(new_n229_) );
  XNOR2_X1 g092 ( .A(new_n151_), .B(new_n229_), .ZN(new_n230_) );
  XOR2_X1 g093 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(new_n231_) );
  AND2_X1 g094 ( .A1(G232GAT), .A2(G233GAT), .ZN(new_n232_) );
  XNOR2_X1 g095 ( .A(new_n231_), .B(new_n232_), .ZN(new_n233_) );
  XNOR2_X1 g096 ( .A(new_n233_), .B(KEYINPUT9), .ZN(new_n234_) );
  INV_X1 g097 ( .A(KEYINPUT7), .ZN(new_n235_) );
  XOR2_X1 g098 ( .A(G43GAT), .B(KEYINPUT8), .Z(new_n236_) );
  OR2_X1 g099 ( .A1(new_n236_), .A2(new_n235_), .ZN(new_n237_) );
  INV_X1 g100 ( .A(G43GAT), .ZN(new_n238_) );
  INV_X1 g101 ( .A(KEYINPUT8), .ZN(new_n239_) );
  AND2_X1 g102 ( .A1(new_n238_), .A2(new_n239_), .ZN(new_n240_) );
  AND2_X1 g103 ( .A1(G43GAT), .A2(KEYINPUT8), .ZN(new_n241_) );
  OR2_X1 g104 ( .A1(new_n241_), .A2(KEYINPUT7), .ZN(new_n242_) );
  OR2_X1 g105 ( .A1(new_n242_), .A2(new_n240_), .ZN(new_n243_) );
  AND2_X1 g106 ( .A1(new_n243_), .A2(new_n237_), .ZN(new_n244_) );
  XOR2_X1 g107 ( .A(G85GAT), .B(G99GAT), .Z(new_n245_) );
  OR2_X1 g108 ( .A1(new_n245_), .A2(new_n205_), .ZN(new_n246_) );
  INV_X1 g109 ( .A(G85GAT), .ZN(new_n247_) );
  INV_X1 g110 ( .A(G99GAT), .ZN(new_n248_) );
  AND2_X1 g111 ( .A1(new_n247_), .A2(new_n248_), .ZN(new_n249_) );
  AND2_X1 g112 ( .A1(G85GAT), .A2(G99GAT), .ZN(new_n250_) );
  OR2_X1 g113 ( .A1(new_n250_), .A2(G92GAT), .ZN(new_n251_) );
  OR2_X1 g114 ( .A1(new_n251_), .A2(new_n249_), .ZN(new_n252_) );
  AND2_X1 g115 ( .A1(new_n252_), .A2(new_n246_), .ZN(new_n253_) );
  XNOR2_X1 g116 ( .A(new_n244_), .B(new_n253_), .ZN(new_n254_) );
  XNOR2_X1 g117 ( .A(new_n254_), .B(new_n234_), .ZN(new_n255_) );
  XNOR2_X1 g118 ( .A(new_n255_), .B(new_n230_), .ZN(new_n256_) );
  XNOR2_X1 g119 ( .A(new_n256_), .B(new_n181_), .ZN(new_n257_) );
  XNOR2_X1 g120 ( .A(new_n257_), .B(new_n203_), .ZN(new_n258_) );
  INV_X1 g121 ( .A(new_n258_), .ZN(new_n259_) );
  XNOR2_X1 g122 ( .A(G78GAT), .B(G155GAT), .ZN(new_n260_) );
  XNOR2_X1 g123 ( .A(G127GAT), .B(G211GAT), .ZN(new_n261_) );
  XOR2_X1 g124 ( .A(new_n260_), .B(new_n261_), .Z(new_n262_) );
  XNOR2_X1 g125 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(new_n263_) );
  XNOR2_X1 g126 ( .A(G64GAT), .B(KEYINPUT15), .ZN(new_n264_) );
  XNOR2_X1 g127 ( .A(new_n263_), .B(new_n264_), .ZN(new_n265_) );
  XNOR2_X1 g128 ( .A(new_n262_), .B(new_n265_), .ZN(new_n266_) );
  XNOR2_X1 g129 ( .A(G15GAT), .B(G22GAT), .ZN(new_n267_) );
  XNOR2_X1 g130 ( .A(new_n267_), .B(new_n138_), .ZN(new_n268_) );
  XNOR2_X1 g131 ( .A(G57GAT), .B(G71GAT), .ZN(new_n269_) );
  XOR2_X1 g132 ( .A(new_n269_), .B(KEYINPUT13), .Z(new_n270_) );
  XNOR2_X1 g133 ( .A(new_n270_), .B(new_n268_), .ZN(new_n271_) );
  XOR2_X1 g134 ( .A(new_n266_), .B(new_n271_), .Z(new_n272_) );
  XNOR2_X1 g135 ( .A(new_n272_), .B(new_n210_), .ZN(new_n273_) );
  AND2_X1 g136 ( .A1(G231GAT), .A2(G233GAT), .ZN(new_n274_) );
  XOR2_X1 g137 ( .A(new_n273_), .B(new_n274_), .Z(new_n275_) );
  INV_X1 g138 ( .A(new_n275_), .ZN(new_n276_) );
  AND2_X1 g139 ( .A1(new_n259_), .A2(new_n276_), .ZN(new_n277_) );
  XNOR2_X1 g140 ( .A(new_n277_), .B(KEYINPUT16), .ZN(new_n278_) );
  AND2_X1 g141 ( .A1(new_n228_), .A2(new_n278_), .ZN(new_n279_) );
  XNOR2_X1 g142 ( .A(G8GAT), .B(G169GAT), .ZN(new_n280_) );
  XNOR2_X1 g143 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(new_n281_) );
  XNOR2_X1 g144 ( .A(new_n280_), .B(new_n281_), .ZN(new_n282_) );
  XNOR2_X1 g145 ( .A(G113GAT), .B(G197GAT), .ZN(new_n283_) );
  XNOR2_X1 g146 ( .A(G29GAT), .B(G141GAT), .ZN(new_n284_) );
  XOR2_X1 g147 ( .A(new_n283_), .B(new_n284_), .Z(new_n285_) );
  XNOR2_X1 g148 ( .A(new_n285_), .B(new_n282_), .ZN(new_n286_) );
  XNOR2_X1 g149 ( .A(new_n244_), .B(new_n268_), .ZN(new_n287_) );
  XOR2_X1 g150 ( .A(new_n287_), .B(new_n286_), .Z(new_n288_) );
  XNOR2_X1 g151 ( .A(G36GAT), .B(G50GAT), .ZN(new_n289_) );
  AND2_X1 g152 ( .A1(G229GAT), .A2(G233GAT), .ZN(new_n290_) );
  XNOR2_X1 g153 ( .A(new_n289_), .B(new_n290_), .ZN(new_n291_) );
  XOR2_X1 g154 ( .A(new_n288_), .B(new_n291_), .Z(new_n292_) );
  INV_X1 g155 ( .A(new_n292_), .ZN(new_n293_) );
  INV_X1 g156 ( .A(new_n270_), .ZN(new_n294_) );
  XOR2_X1 g157 ( .A(G120GAT), .B(G204GAT), .Z(new_n295_) );
  XNOR2_X1 g158 ( .A(new_n177_), .B(new_n253_), .ZN(new_n296_) );
  XNOR2_X1 g159 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(new_n297_) );
  AND2_X1 g160 ( .A1(G230GAT), .A2(G233GAT), .ZN(new_n298_) );
  XNOR2_X1 g161 ( .A(new_n297_), .B(new_n298_), .ZN(new_n299_) );
  XNOR2_X1 g162 ( .A(new_n299_), .B(KEYINPUT32), .ZN(new_n300_) );
  XNOR2_X1 g163 ( .A(new_n296_), .B(new_n300_), .ZN(new_n301_) );
  XNOR2_X1 g164 ( .A(new_n301_), .B(new_n206_), .ZN(new_n302_) );
  XNOR2_X1 g165 ( .A(new_n302_), .B(new_n295_), .ZN(new_n303_) );
  XNOR2_X1 g166 ( .A(new_n303_), .B(new_n294_), .ZN(new_n304_) );
  INV_X1 g167 ( .A(new_n304_), .ZN(new_n305_) );
  AND2_X1 g168 ( .A1(new_n305_), .A2(new_n293_), .ZN(new_n306_) );
  AND2_X1 g169 ( .A1(new_n279_), .A2(new_n306_), .ZN(new_n307_) );
  AND2_X1 g170 ( .A1(new_n307_), .A2(new_n159_), .ZN(new_n308_) );
  XNOR2_X1 g171 ( .A(new_n308_), .B(KEYINPUT34), .ZN(new_n309_) );
  XNOR2_X1 g172 ( .A(new_n309_), .B(new_n138_), .ZN(G1324GAT) );
  AND2_X1 g173 ( .A1(new_n307_), .A2(new_n213_), .ZN(new_n311_) );
  XOR2_X1 g174 ( .A(new_n311_), .B(G8GAT), .Z(G1325GAT) );
  AND2_X1 g175 ( .A1(new_n307_), .A2(new_n199_), .ZN(new_n313_) );
  XNOR2_X1 g176 ( .A(G15GAT), .B(KEYINPUT35), .ZN(new_n314_) );
  XNOR2_X1 g177 ( .A(new_n313_), .B(new_n314_), .ZN(G1326GAT) );
  AND2_X1 g178 ( .A1(new_n307_), .A2(new_n223_), .ZN(new_n316_) );
  XOR2_X1 g179 ( .A(new_n316_), .B(G22GAT), .Z(G1327GAT) );
  XOR2_X1 g180 ( .A(new_n258_), .B(KEYINPUT36), .Z(new_n318_) );
  INV_X1 g181 ( .A(new_n318_), .ZN(new_n319_) );
  AND2_X1 g182 ( .A1(new_n319_), .A2(new_n275_), .ZN(new_n320_) );
  AND2_X1 g183 ( .A1(new_n228_), .A2(new_n320_), .ZN(new_n321_) );
  XOR2_X1 g184 ( .A(new_n321_), .B(KEYINPUT37), .Z(new_n322_) );
  AND2_X1 g185 ( .A1(new_n322_), .A2(new_n306_), .ZN(new_n323_) );
  XNOR2_X1 g186 ( .A(new_n323_), .B(KEYINPUT38), .ZN(new_n324_) );
  AND2_X1 g187 ( .A1(new_n324_), .A2(new_n159_), .ZN(new_n325_) );
  XNOR2_X1 g188 ( .A(G29GAT), .B(KEYINPUT39), .ZN(new_n326_) );
  XNOR2_X1 g189 ( .A(new_n325_), .B(new_n326_), .ZN(G1328GAT) );
  AND2_X1 g190 ( .A1(new_n324_), .A2(new_n213_), .ZN(new_n328_) );
  XOR2_X1 g191 ( .A(new_n328_), .B(G36GAT), .Z(G1329GAT) );
  AND2_X1 g192 ( .A1(new_n324_), .A2(new_n199_), .ZN(new_n330_) );
  XNOR2_X1 g193 ( .A(new_n330_), .B(KEYINPUT40), .ZN(new_n331_) );
  XNOR2_X1 g194 ( .A(new_n331_), .B(new_n238_), .ZN(G1330GAT) );
  AND2_X1 g195 ( .A1(new_n324_), .A2(new_n223_), .ZN(new_n333_) );
  XOR2_X1 g196 ( .A(new_n333_), .B(G50GAT), .Z(G1331GAT) );
  INV_X1 g197 ( .A(KEYINPUT41), .ZN(new_n335_) );
  XNOR2_X1 g198 ( .A(new_n304_), .B(new_n335_), .ZN(new_n336_) );
  AND2_X1 g199 ( .A1(new_n336_), .A2(new_n292_), .ZN(new_n337_) );
  AND2_X1 g200 ( .A1(new_n279_), .A2(new_n337_), .ZN(new_n338_) );
  AND2_X1 g201 ( .A1(new_n338_), .A2(new_n159_), .ZN(new_n339_) );
  XOR2_X1 g202 ( .A(G57GAT), .B(KEYINPUT42), .Z(new_n340_) );
  XNOR2_X1 g203 ( .A(new_n339_), .B(new_n340_), .ZN(G1332GAT) );
  AND2_X1 g204 ( .A1(new_n338_), .A2(new_n213_), .ZN(new_n342_) );
  XOR2_X1 g205 ( .A(new_n342_), .B(G64GAT), .Z(G1333GAT) );
  AND2_X1 g206 ( .A1(new_n338_), .A2(new_n199_), .ZN(new_n344_) );
  XOR2_X1 g207 ( .A(new_n344_), .B(G71GAT), .Z(G1334GAT) );
  AND2_X1 g208 ( .A1(new_n338_), .A2(new_n223_), .ZN(new_n346_) );
  XNOR2_X1 g209 ( .A(G78GAT), .B(KEYINPUT43), .ZN(new_n347_) );
  XNOR2_X1 g210 ( .A(new_n346_), .B(new_n347_), .ZN(G1335GAT) );
  AND2_X1 g211 ( .A1(new_n322_), .A2(new_n337_), .ZN(new_n349_) );
  AND2_X1 g212 ( .A1(new_n349_), .A2(new_n159_), .ZN(new_n350_) );
  XNOR2_X1 g213 ( .A(new_n350_), .B(new_n247_), .ZN(G1336GAT) );
  AND2_X1 g214 ( .A1(new_n349_), .A2(new_n213_), .ZN(new_n352_) );
  XNOR2_X1 g215 ( .A(new_n352_), .B(new_n205_), .ZN(G1337GAT) );
  AND2_X1 g216 ( .A1(new_n349_), .A2(new_n199_), .ZN(new_n354_) );
  XNOR2_X1 g217 ( .A(new_n354_), .B(new_n248_), .ZN(G1338GAT) );
  AND2_X1 g218 ( .A1(new_n349_), .A2(new_n223_), .ZN(new_n356_) );
  XNOR2_X1 g219 ( .A(new_n356_), .B(KEYINPUT44), .ZN(new_n357_) );
  XNOR2_X1 g220 ( .A(new_n357_), .B(new_n172_), .ZN(G1339GAT) );
  AND2_X1 g221 ( .A1(new_n336_), .A2(new_n293_), .ZN(new_n359_) );
  AND2_X1 g222 ( .A1(new_n359_), .A2(KEYINPUT46), .ZN(new_n360_) );
  INV_X1 g223 ( .A(KEYINPUT46), .ZN(new_n361_) );
  XNOR2_X1 g224 ( .A(new_n304_), .B(KEYINPUT41), .ZN(new_n362_) );
  OR2_X1 g225 ( .A1(new_n362_), .A2(new_n292_), .ZN(new_n363_) );
  AND2_X1 g226 ( .A1(new_n363_), .A2(new_n361_), .ZN(new_n364_) );
  AND2_X1 g227 ( .A1(new_n259_), .A2(new_n275_), .ZN(new_n365_) );
  INV_X1 g228 ( .A(new_n365_), .ZN(new_n366_) );
  OR2_X1 g229 ( .A1(new_n364_), .A2(new_n366_), .ZN(new_n367_) );
  OR2_X1 g230 ( .A1(new_n367_), .A2(new_n360_), .ZN(new_n368_) );
  AND2_X1 g231 ( .A1(new_n368_), .A2(KEYINPUT47), .ZN(new_n369_) );
  INV_X1 g232 ( .A(new_n369_), .ZN(new_n370_) );
  OR2_X1 g233 ( .A1(new_n368_), .A2(KEYINPUT47), .ZN(new_n371_) );
  INV_X1 g234 ( .A(KEYINPUT45), .ZN(new_n372_) );
  OR2_X1 g235 ( .A1(new_n318_), .A2(new_n275_), .ZN(new_n373_) );
  INV_X1 g236 ( .A(new_n373_), .ZN(new_n374_) );
  OR2_X1 g237 ( .A1(new_n374_), .A2(new_n372_), .ZN(new_n375_) );
  OR2_X1 g238 ( .A1(new_n373_), .A2(KEYINPUT45), .ZN(new_n376_) );
  AND2_X1 g239 ( .A1(new_n305_), .A2(new_n292_), .ZN(new_n377_) );
  AND2_X1 g240 ( .A1(new_n376_), .A2(new_n377_), .ZN(new_n378_) );
  AND2_X1 g241 ( .A1(new_n378_), .A2(new_n375_), .ZN(new_n379_) );
  INV_X1 g242 ( .A(new_n379_), .ZN(new_n380_) );
  AND2_X1 g243 ( .A1(new_n371_), .A2(new_n380_), .ZN(new_n381_) );
  AND2_X1 g244 ( .A1(new_n381_), .A2(new_n370_), .ZN(new_n382_) );
  AND2_X1 g245 ( .A1(new_n382_), .A2(KEYINPUT48), .ZN(new_n383_) );
  INV_X1 g246 ( .A(new_n383_), .ZN(new_n384_) );
  OR2_X1 g247 ( .A1(new_n382_), .A2(KEYINPUT48), .ZN(new_n385_) );
  AND2_X1 g248 ( .A1(new_n385_), .A2(new_n225_), .ZN(new_n386_) );
  AND2_X1 g249 ( .A1(new_n386_), .A2(new_n384_), .ZN(new_n387_) );
  AND2_X1 g250 ( .A1(new_n224_), .A2(new_n199_), .ZN(new_n388_) );
  AND2_X1 g251 ( .A1(new_n387_), .A2(new_n388_), .ZN(new_n389_) );
  AND2_X1 g252 ( .A1(new_n389_), .A2(new_n293_), .ZN(new_n390_) );
  XOR2_X1 g253 ( .A(new_n390_), .B(G113GAT), .Z(G1340GAT) );
  AND2_X1 g254 ( .A1(new_n389_), .A2(new_n336_), .ZN(new_n392_) );
  XNOR2_X1 g255 ( .A(G120GAT), .B(KEYINPUT49), .ZN(new_n393_) );
  XNOR2_X1 g256 ( .A(new_n392_), .B(new_n393_), .ZN(G1341GAT) );
  AND2_X1 g257 ( .A1(new_n389_), .A2(new_n276_), .ZN(new_n395_) );
  XOR2_X1 g258 ( .A(new_n395_), .B(KEYINPUT50), .Z(new_n396_) );
  XNOR2_X1 g259 ( .A(new_n396_), .B(G127GAT), .ZN(G1342GAT) );
  AND2_X1 g260 ( .A1(new_n389_), .A2(new_n258_), .ZN(new_n398_) );
  XNOR2_X1 g261 ( .A(G134GAT), .B(KEYINPUT51), .ZN(new_n399_) );
  XNOR2_X1 g262 ( .A(new_n398_), .B(new_n399_), .ZN(G1343GAT) );
  AND2_X1 g263 ( .A1(new_n387_), .A2(new_n201_), .ZN(new_n401_) );
  AND2_X1 g264 ( .A1(new_n401_), .A2(new_n293_), .ZN(new_n402_) );
  XOR2_X1 g265 ( .A(new_n402_), .B(G141GAT), .Z(G1344GAT) );
  AND2_X1 g266 ( .A1(new_n401_), .A2(new_n336_), .ZN(new_n404_) );
  XNOR2_X1 g267 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(new_n405_) );
  XNOR2_X1 g268 ( .A(new_n404_), .B(new_n405_), .ZN(new_n406_) );
  XNOR2_X1 g269 ( .A(new_n406_), .B(G148GAT), .ZN(G1345GAT) );
  AND2_X1 g270 ( .A1(new_n401_), .A2(new_n276_), .ZN(new_n408_) );
  XOR2_X1 g271 ( .A(new_n408_), .B(G155GAT), .Z(G1346GAT) );
  AND2_X1 g272 ( .A1(new_n401_), .A2(new_n258_), .ZN(new_n410_) );
  XOR2_X1 g273 ( .A(new_n410_), .B(G162GAT), .Z(G1347GAT) );
  INV_X1 g274 ( .A(KEYINPUT55), .ZN(new_n412_) );
  INV_X1 g275 ( .A(KEYINPUT54), .ZN(new_n413_) );
  AND2_X1 g276 ( .A1(new_n385_), .A2(new_n213_), .ZN(new_n414_) );
  AND2_X1 g277 ( .A1(new_n414_), .A2(new_n384_), .ZN(new_n415_) );
  OR2_X1 g278 ( .A1(new_n415_), .A2(new_n413_), .ZN(new_n416_) );
  AND2_X1 g279 ( .A1(new_n416_), .A2(new_n158_), .ZN(new_n417_) );
  INV_X1 g280 ( .A(KEYINPUT48), .ZN(new_n418_) );
  INV_X1 g281 ( .A(KEYINPUT47), .ZN(new_n419_) );
  INV_X1 g282 ( .A(new_n360_), .ZN(new_n420_) );
  OR2_X1 g283 ( .A1(new_n359_), .A2(KEYINPUT46), .ZN(new_n421_) );
  AND2_X1 g284 ( .A1(new_n421_), .A2(new_n365_), .ZN(new_n422_) );
  AND2_X1 g285 ( .A1(new_n422_), .A2(new_n420_), .ZN(new_n423_) );
  AND2_X1 g286 ( .A1(new_n423_), .A2(new_n419_), .ZN(new_n424_) );
  OR2_X1 g287 ( .A1(new_n424_), .A2(new_n379_), .ZN(new_n425_) );
  OR2_X1 g288 ( .A1(new_n425_), .A2(new_n369_), .ZN(new_n426_) );
  AND2_X1 g289 ( .A1(new_n426_), .A2(new_n418_), .ZN(new_n427_) );
  OR2_X1 g290 ( .A1(new_n427_), .A2(new_n217_), .ZN(new_n428_) );
  OR2_X1 g291 ( .A1(new_n428_), .A2(new_n383_), .ZN(new_n429_) );
  OR2_X1 g292 ( .A1(new_n429_), .A2(KEYINPUT54), .ZN(new_n430_) );
  AND2_X1 g293 ( .A1(new_n430_), .A2(new_n184_), .ZN(new_n431_) );
  AND2_X1 g294 ( .A1(new_n417_), .A2(new_n431_), .ZN(new_n432_) );
  XNOR2_X1 g295 ( .A(new_n432_), .B(new_n412_), .ZN(new_n433_) );
  AND2_X1 g296 ( .A1(new_n433_), .A2(new_n199_), .ZN(new_n434_) );
  AND2_X1 g297 ( .A1(new_n434_), .A2(new_n293_), .ZN(new_n435_) );
  XOR2_X1 g298 ( .A(new_n435_), .B(G169GAT), .Z(G1348GAT) );
  INV_X1 g299 ( .A(G176GAT), .ZN(new_n437_) );
  AND2_X1 g300 ( .A1(new_n434_), .A2(new_n336_), .ZN(new_n438_) );
  XOR2_X1 g301 ( .A(KEYINPUT57), .B(KEYINPUT56), .Z(new_n439_) );
  XNOR2_X1 g302 ( .A(new_n438_), .B(new_n439_), .ZN(new_n440_) );
  XNOR2_X1 g303 ( .A(new_n440_), .B(new_n437_), .ZN(G1349GAT) );
  AND2_X1 g304 ( .A1(new_n434_), .A2(new_n276_), .ZN(new_n442_) );
  XOR2_X1 g305 ( .A(new_n442_), .B(G183GAT), .Z(G1350GAT) );
  AND2_X1 g306 ( .A1(new_n434_), .A2(new_n258_), .ZN(new_n444_) );
  XOR2_X1 g307 ( .A(G190GAT), .B(KEYINPUT58), .Z(new_n445_) );
  XNOR2_X1 g308 ( .A(new_n444_), .B(new_n445_), .ZN(G1351GAT) );
  AND2_X1 g309 ( .A1(new_n430_), .A2(new_n201_), .ZN(new_n447_) );
  AND2_X1 g310 ( .A1(new_n417_), .A2(new_n447_), .ZN(new_n448_) );
  AND2_X1 g311 ( .A1(new_n448_), .A2(new_n293_), .ZN(new_n449_) );
  XNOR2_X1 g312 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(new_n450_) );
  XNOR2_X1 g313 ( .A(new_n449_), .B(new_n450_), .ZN(new_n451_) );
  XNOR2_X1 g314 ( .A(new_n451_), .B(G197GAT), .ZN(G1352GAT) );
  AND2_X1 g315 ( .A1(new_n448_), .A2(new_n304_), .ZN(new_n453_) );
  XNOR2_X1 g316 ( .A(G204GAT), .B(KEYINPUT61), .ZN(new_n454_) );
  XNOR2_X1 g317 ( .A(new_n453_), .B(new_n454_), .ZN(G1353GAT) );
  AND2_X1 g318 ( .A1(new_n448_), .A2(new_n276_), .ZN(new_n456_) );
  XOR2_X1 g319 ( .A(new_n456_), .B(G211GAT), .Z(G1354GAT) );
  AND2_X1 g320 ( .A1(new_n448_), .A2(new_n319_), .ZN(new_n458_) );
  XNOR2_X1 g321 ( .A(new_n458_), .B(KEYINPUT62), .ZN(new_n459_) );
  XOR2_X1 g322 ( .A(new_n459_), .B(G218GAT), .Z(G1355GAT) );
endmodule


