module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n595_, new_n1233_, new_n445_, new_n1009_, new_n238_, new_n479_, new_n1105_, new_n1215_, new_n608_, new_n501_, new_n1157_, new_n421_, new_n777_, new_n1048_, new_n885_, new_n439_, new_n283_, new_n223_, new_n390_, new_n743_, new_n241_, new_n566_, new_n186_, new_n339_, new_n641_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n1024_, new_n1125_, new_n246_, new_n911_, new_n679_, new_n937_, new_n667_, new_n367_, new_n1237_, new_n173_, new_n728_, new_n1071_, new_n214_, new_n894_, new_n853_, new_n695_, new_n660_, new_n526_, new_n908_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n1119_, new_n752_, new_n1045_, new_n500_, new_n1163_, new_n786_, new_n317_, new_n1188_, new_n721_, new_n504_, new_n742_, new_n892_, new_n234_, new_n472_, new_n873_, new_n1167_, new_n774_, new_n792_, new_n953_, new_n257_, new_n481_, new_n1073_, new_n1110_, new_n449_, new_n580_, new_n639_, new_n484_, new_n766_, new_n272_, new_n282_, new_n1212_, new_n1059_, new_n634_, new_n192_, new_n635_, new_n685_, new_n326_, new_n648_, new_n903_, new_n983_, new_n822_, new_n1082_, new_n1018_, new_n606_, new_n796_, new_n655_, new_n1054_, new_n630_, new_n385_, new_n1049_, new_n694_, new_n461_, new_n297_, new_n565_, new_n1196_, new_n183_, new_n511_, new_n303_, new_n325_, new_n1031_, new_n1216_, new_n629_, new_n1214_, new_n883_, new_n1005_, new_n999_, new_n321_, new_n324_, new_n960_, new_n491_, new_n549_, new_n676_, new_n995_, new_n1035_, new_n271_, new_n674_, new_n274_, new_n991_, new_n1044_, new_n497_, new_n816_, new_n568_, new_n420_, new_n876_, new_n423_, new_n498_, new_n496_, new_n1217_, new_n1046_, new_n1182_, new_n708_, new_n206_, new_n429_, new_n1222_, new_n353_, new_n734_, new_n912_, new_n1062_, new_n506_, new_n680_, new_n872_, new_n981_, new_n1198_, new_n656_, new_n1127_, new_n388_, new_n1028_, new_n1168_, new_n194_, new_n483_, new_n1004_, new_n1152_, new_n394_, new_n299_, new_n935_, new_n657_, new_n1150_, new_n652_, new_n582_, new_n1020_, new_n363_, new_n1113_, new_n441_, new_n785_, new_n477_, new_n664_, new_n600_, new_n280_, new_n1041_, new_n426_, new_n1036_, new_n235_, new_n398_, new_n301_, new_n1132_, new_n395_, new_n383_, new_n343_, new_n854_, new_n458_, new_n1106_, new_n207_, new_n267_, new_n473_, new_n1147_, new_n1229_, new_n187_, new_n969_, new_n334_, new_n331_, new_n835_, new_n1234_, new_n378_, new_n621_, new_n244_, new_n172_, new_n705_, new_n943_, new_n874_, new_n402_, new_n1209_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n1003_, new_n696_, new_n208_, new_n1039_, new_n1239_, new_n528_, new_n952_, new_n179_, new_n729_, new_n1111_, new_n1218_, new_n559_, new_n1201_, new_n762_, new_n1193_, new_n1187_, new_n1205_, new_n1154_, new_n295_, new_n628_, new_n409_, new_n1090_, new_n745_, new_n553_, new_n1114_, new_n1084_, new_n1061_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n1032_, new_n867_, new_n954_, new_n901_, new_n1171_, new_n276_, new_n688_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n886_, new_n371_, new_n509_, new_n202_, new_n296_, new_n661_, new_n797_, new_n232_, new_n724_, new_n1070_, new_n1109_, new_n261_, new_n672_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n938_, new_n362_, new_n809_, new_n1142_, new_n1104_, new_n571_, new_n758_, new_n328_, new_n460_, new_n268_, new_n380_, new_n1079_, new_n861_, new_n352_, new_n931_, new_n575_, new_n562_, new_n944_, new_n1064_, new_n1065_, new_n177_, new_n1118_, new_n493_, new_n547_, new_n264_, new_n379_, new_n273_, new_n224_, new_n586_, new_n963_, new_n993_, new_n1191_, new_n824_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n858_, new_n936_, new_n189_, new_n411_, new_n1016_, new_n673_, new_n1144_, new_n182_, new_n407_, new_n666_, new_n736_, new_n879_, new_n513_, new_n558_, new_n219_, new_n313_, new_n382_, new_n239_, new_n718_, new_n1126_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n302_, new_n755_, new_n1040_, new_n544_, new_n615_, new_n722_, new_n856_, new_n415_, new_n537_, new_n345_, new_n499_, new_n255_, new_n533_, new_n1130_, new_n795_, new_n459_, new_n1122_, new_n1185_, new_n1240_, new_n354_, new_n1174_, new_n968_, new_n613_, new_n337_, new_n1195_, new_n417_, new_n658_, new_n591_, new_n837_, new_n801_, new_n631_, new_n453_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n531_, new_n593_, new_n974_, new_n252_, new_n751_, new_n1038_, new_n372_, new_n852_, new_n978_, new_n408_, new_n470_, new_n213_, new_n769_, new_n433_, new_n871_, new_n992_, new_n1098_, new_n265_, new_n732_, new_n689_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n1052_, new_n857_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n269_, new_n512_, new_n1220_, new_n989_, new_n1117_, new_n644_, new_n836_, new_n1116_, new_n904_, new_n913_, new_n327_, new_n681_, new_n594_, new_n561_, new_n495_, new_n927_, new_n431_, new_n1206_, new_n196_, new_n818_, new_n881_, new_n640_, new_n684_, new_n754_, new_n653_, new_n377_, new_n905_, new_n375_, new_n962_, new_n760_, new_n627_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n1153_, new_n357_, new_n320_, new_n780_, new_n984_, new_n1183_, new_n245_, new_n643_, new_n1194_, new_n1230_, new_n1027_, new_n348_, new_n610_, new_n843_, new_n322_, new_n703_, new_n698_, new_n1165_, new_n175_, new_n226_, new_n1208_, new_n697_, new_n1099_, new_n185_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n1235_, new_n540_, new_n1149_, new_n1066_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n770_, new_n757_, new_n1225_, new_n521_, new_n793_, new_n406_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n1089_, new_n1192_, new_n405_, new_n942_, new_n614_, new_n895_, new_n958_, new_n976_, new_n699_, new_n236_, new_n955_, new_n847_, new_n250_, new_n288_, new_n798_, new_n1180_, new_n817_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n941_, new_n827_, new_n366_, new_n779_, new_n1232_, new_n1025_, new_n365_, new_n859_, new_n197_, new_n1211_, new_n1207_, new_n1176_, new_n601_, new_n842_, new_n1057_, new_n682_, new_n1075_, new_n812_, new_n266_, new_n821_, new_n542_, new_n548_, new_n669_, new_n220_, new_n1172_, new_n419_, new_n624_, new_n534_, new_n1131_, new_n1120_, new_n819_, new_n637_, new_n451_, new_n489_, new_n424_, new_n804_, new_n602_, new_n1210_, new_n188_, new_n1060_, new_n240_, new_n413_, new_n442_, new_n677_, new_n642_, new_n211_, new_n462_, new_n603_, new_n564_, new_n761_, new_n840_, new_n735_, new_n898_, new_n799_, new_n946_, new_n344_, new_n287_, new_n1108_, new_n862_, new_n427_, new_n532_, new_n393_, new_n418_, new_n746_, new_n1221_, new_n292_, new_n215_, new_n626_, new_n959_, new_n990_, new_n716_, new_n701_, new_n1238_, new_n1058_, new_n1162_, new_n212_, new_n902_, new_n364_, new_n832_, new_n201_, new_n414_, new_n1101_, new_n315_, new_n1050_, new_n554_, new_n230_, new_n1151_, new_n281_, new_n430_, new_n844_, new_n482_, new_n849_, new_n1203_, new_n855_, new_n1037_, new_n589_, new_n248_, new_n350_, new_n759_, new_n1083_, new_n829_, new_n988_, new_n478_, new_n1228_, new_n710_, new_n971_, new_n906_, new_n361_, new_n764_, new_n683_, new_n463_, new_n510_, new_n966_, new_n351_, new_n1184_, new_n517_, new_n609_, new_n180_, new_n961_, new_n530_, new_n890_, new_n318_, new_n1006_, new_n622_, new_n702_, new_n833_, new_n715_, new_n811_, new_n443_, new_n1086_, new_n956_, new_n763_, new_n1138_, new_n486_, new_n970_, new_n466_, new_n262_, new_n218_, new_n1170_, new_n845_, new_n768_, new_n773_, new_n1051_, new_n899_, new_n1053_, new_n205_, new_n492_, new_n1200_, new_n650_, new_n750_, new_n887_, new_n254_, new_n355_, new_n926_, new_n432_, new_n925_, new_n875_, new_n256_, new_n1226_, new_n778_, new_n452_, new_n381_, new_n1219_, new_n920_, new_n1121_, new_n820_, new_n771_, new_n979_, new_n508_, new_n714_, new_n1007_, new_n882_, new_n1145_, new_n929_, new_n986_, new_n314_, new_n1159_, new_n216_, new_n917_, new_n1133_, new_n1177_, new_n646_, new_n538_, new_n1026_, new_n210_, new_n541_, new_n447_, new_n790_, new_n1081_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n263_, new_n341_, new_n996_, new_n846_, new_n915_, new_n349_, new_n488_, new_n524_, new_n848_, new_n277_, new_n663_, new_n579_, new_n286_, new_n198_, new_n438_, new_n939_, new_n632_, new_n671_, new_n965_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n1202_, new_n397_, new_n975_, new_n1199_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n1115_, new_n948_, new_n1231_, new_n1055_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n1085_, new_n359_, new_n794_, new_n457_, new_n1128_, new_n1002_, new_n1169_, new_n448_, new_n384_, new_n900_, new_n1161_, new_n924_, new_n775_, new_n454_, new_n1034_, new_n1124_, new_n308_, new_n1000_, new_n633_, new_n784_, new_n258_, new_n176_, new_n860_, new_n306_, new_n494_, new_n291_, new_n309_, new_n1160_, new_n1166_, new_n259_, new_n654_, new_n713_, new_n880_, new_n1102_, new_n227_, new_n690_, new_n416_, new_n222_, new_n1043_, new_n744_, new_n400_, new_n1175_, new_n693_, new_n505_, new_n619_, new_n471_, new_n967_, new_n577_, new_n374_, new_n1135_, new_n376_, new_n747_, new_n749_, new_n1091_, new_n310_, new_n1095_, new_n275_, new_n998_, new_n1056_, new_n1094_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n578_, new_n918_, new_n940_, new_n810_, new_n808_, new_n907_, new_n665_, new_n800_, new_n897_, new_n1012_, new_n719_, new_n869_, new_n1178_, new_n270_, new_n570_, new_n598_, new_n893_, new_n1063_, new_n520_, new_n1001_, new_n253_, new_n825_, new_n557_, new_n260_, new_n251_, new_n300_, new_n507_, new_n741_, new_n806_, new_n605_, new_n1224_, new_n1074_, new_n748_, new_n1137_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n1141_, new_n807_, new_n592_, new_n726_, new_n1123_, new_n231_, new_n583_, new_n617_, new_n1080_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n199_, new_n487_, new_n360_, new_n675_, new_n1155_, new_n1186_, new_n191_, new_n225_, new_n922_, new_n387_, new_n476_, new_n987_, new_n949_, new_n221_, new_n243_, new_n450_, new_n1179_, new_n298_, new_n184_, new_n1088_, new_n1148_, new_n1146_, new_n569_, new_n555_, new_n174_, new_n468_, new_n977_, new_n1139_, new_n782_, new_n444_, new_n392_, new_n518_, new_n950_, new_n737_, new_n1022_, new_n340_, new_n285_, new_n692_, new_n502_, new_n209_, new_n623_, new_n446_, new_n203_, new_n316_, new_n590_, new_n826_, new_n789_, new_n515_, new_n332_, new_n972_, new_n1067_, new_n891_, new_n516_, new_n1227_, new_n733_, new_n1021_, new_n1076_, new_n585_, new_n312_, new_n535_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n307_, new_n190_, new_n1181_, new_n597_, new_n1093_, new_n1092_, new_n1143_, new_n1072_, new_n1190_, new_n1097_, new_n1069_, new_n651_, new_n1164_, new_n435_, new_n1010_, new_n776_, new_n687_, new_n370_, new_n1029_, new_n638_, new_n523_, new_n909_, new_n217_, new_n788_, new_n841_, new_n1204_, new_n1112_, new_n711_, new_n1156_, new_n731_, new_n599_, new_n930_, new_n973_, new_n412_, new_n607_, new_n645_, new_n1096_, new_n1087_, new_n723_, new_n756_, new_n823_, new_n574_, new_n928_, new_n319_, new_n1008_, new_n338_, new_n707_, new_n740_, new_n957_, new_n1047_, new_n787_, new_n1134_, new_n336_, new_n247_, new_n539_, new_n803_, new_n330_, new_n727_, new_n294_, new_n1173_, new_n704_, new_n1189_, new_n1197_, new_n474_, new_n1223_, new_n1129_, new_n467_, new_n1013_, new_n404_, new_n1077_, new_n193_, new_n490_, new_n560_, new_n1100_, new_n865_, new_n358_, new_n877_, new_n545_, new_n228_, new_n611_, new_n289_, new_n1011_, new_n425_, new_n896_, new_n802_, new_n1236_, new_n866_, new_n947_, new_n994_, new_n982_, new_n964_, new_n1078_, new_n551_, new_n279_, new_n455_, new_n618_, new_n1140_, new_n1042_, new_n863_, new_n828_, new_n980_, new_n464_, new_n204_, new_n181_, new_n573_, new_n765_, new_n1103_;

not g0000 ( new_n172_, keyIn_0_14 );
and g0001 ( new_n173_, keyIn_0_0, N1 );
not g0002 ( new_n174_, new_n173_ );
or g0003 ( new_n175_, keyIn_0_0, N1 );
and g0004 ( new_n176_, new_n174_, new_n175_ );
not g0005 ( new_n177_, new_n176_ );
and g0006 ( new_n178_, new_n177_, N4 );
or g0007 ( new_n179_, new_n178_, new_n172_ );
not g0008 ( new_n180_, new_n179_ );
and g0009 ( new_n181_, new_n178_, new_n172_ );
or g0010 ( new_n182_, new_n180_, new_n181_ );
not g0011 ( new_n183_, N95 );
not g0012 ( new_n184_, keyIn_0_11 );
or g0013 ( new_n185_, new_n184_, N89 );
not g0014 ( new_n186_, N89 );
or g0015 ( new_n187_, new_n186_, keyIn_0_11 );
and g0016 ( new_n188_, new_n185_, new_n187_ );
or g0017 ( new_n189_, new_n188_, new_n183_ );
and g0018 ( new_n190_, new_n189_, keyIn_0_20 );
not g0019 ( new_n191_, keyIn_0_20 );
and g0020 ( new_n192_, new_n186_, keyIn_0_11 );
and g0021 ( new_n193_, new_n184_, N89 );
or g0022 ( new_n194_, new_n192_, new_n193_ );
and g0023 ( new_n195_, new_n194_, N95 );
and g0024 ( new_n196_, new_n195_, new_n191_ );
or g0025 ( new_n197_, new_n190_, new_n196_ );
not g0026 ( new_n198_, keyIn_0_19 );
or g0027 ( new_n199_, keyIn_0_7, N50 );
not g0028 ( new_n200_, new_n199_ );
not g0029 ( new_n201_, N56 );
and g0030 ( new_n202_, keyIn_0_7, N50 );
or g0031 ( new_n203_, new_n202_, new_n201_ );
or g0032 ( new_n204_, new_n203_, new_n200_ );
and g0033 ( new_n205_, new_n204_, new_n198_ );
not g0034 ( new_n206_, new_n205_ );
or g0035 ( new_n207_, new_n204_, new_n198_ );
and g0036 ( new_n208_, new_n206_, new_n207_ );
or g0037 ( new_n209_, new_n197_, new_n208_ );
or g0038 ( new_n210_, new_n209_, new_n182_ );
not g0039 ( new_n211_, keyIn_0_18 );
not g0040 ( new_n212_, N43 );
not g0041 ( new_n213_, keyIn_0_6 );
or g0042 ( new_n214_, new_n213_, N37 );
not g0043 ( new_n215_, N37 );
or g0044 ( new_n216_, new_n215_, keyIn_0_6 );
and g0045 ( new_n217_, new_n214_, new_n216_ );
or g0046 ( new_n218_, new_n217_, new_n212_ );
or g0047 ( new_n219_, new_n218_, new_n211_ );
and g0048 ( new_n220_, new_n215_, keyIn_0_6 );
and g0049 ( new_n221_, new_n213_, N37 );
or g0050 ( new_n222_, new_n220_, new_n221_ );
and g0051 ( new_n223_, new_n222_, N43 );
or g0052 ( new_n224_, new_n223_, keyIn_0_18 );
and g0053 ( new_n225_, new_n219_, new_n224_ );
not g0054 ( new_n226_, keyIn_0_9 );
and g0055 ( new_n227_, new_n226_, N76 );
not g0056 ( new_n228_, new_n227_ );
or g0057 ( new_n229_, new_n226_, N76 );
and g0058 ( new_n230_, new_n229_, N82 );
and g0059 ( new_n231_, new_n230_, new_n228_ );
not g0060 ( new_n232_, keyIn_0_2 );
not g0061 ( new_n233_, N11 );
and g0062 ( new_n234_, new_n232_, new_n233_ );
and g0063 ( new_n235_, keyIn_0_2, N11 );
or g0064 ( new_n236_, new_n234_, new_n235_ );
and g0065 ( new_n237_, new_n236_, N17 );
not g0066 ( new_n238_, N63 );
and g0067 ( new_n239_, new_n238_, N69 );
or g0068 ( new_n240_, new_n237_, new_n239_ );
or g0069 ( new_n241_, new_n240_, new_n231_ );
or g0070 ( new_n242_, new_n225_, new_n241_ );
not g0071 ( new_n243_, keyIn_0_21 );
or g0072 ( new_n244_, keyIn_0_12, N102 );
not g0073 ( new_n245_, new_n244_ );
not g0074 ( new_n246_, N108 );
and g0075 ( new_n247_, keyIn_0_12, N102 );
or g0076 ( new_n248_, new_n247_, new_n246_ );
or g0077 ( new_n249_, new_n248_, new_n245_ );
not g0078 ( new_n250_, new_n249_ );
and g0079 ( new_n251_, new_n250_, new_n243_ );
and g0080 ( new_n252_, new_n249_, keyIn_0_21 );
or g0081 ( new_n253_, new_n251_, new_n252_ );
not g0082 ( new_n254_, keyIn_0_17 );
or g0083 ( new_n255_, keyIn_0_4, N24 );
not g0084 ( new_n256_, new_n255_ );
not g0085 ( new_n257_, N30 );
and g0086 ( new_n258_, keyIn_0_4, N24 );
or g0087 ( new_n259_, new_n258_, new_n257_ );
or g0088 ( new_n260_, new_n259_, new_n256_ );
and g0089 ( new_n261_, new_n260_, new_n254_ );
not g0090 ( new_n262_, new_n261_ );
or g0091 ( new_n263_, new_n260_, new_n254_ );
and g0092 ( new_n264_, new_n262_, new_n263_ );
or g0093 ( new_n265_, new_n253_, new_n264_ );
or g0094 ( new_n266_, new_n242_, new_n265_ );
or g0095 ( new_n267_, new_n266_, new_n210_ );
and g0096 ( new_n268_, new_n267_, keyIn_0_38 );
not g0097 ( new_n269_, keyIn_0_38 );
not g0098 ( new_n270_, new_n181_ );
and g0099 ( new_n271_, new_n270_, new_n179_ );
or g0100 ( new_n272_, new_n195_, new_n191_ );
or g0101 ( new_n273_, new_n189_, keyIn_0_20 );
and g0102 ( new_n274_, new_n273_, new_n272_ );
not g0103 ( new_n275_, new_n203_ );
and g0104 ( new_n276_, new_n275_, new_n199_ );
and g0105 ( new_n277_, new_n276_, keyIn_0_19 );
or g0106 ( new_n278_, new_n277_, new_n205_ );
and g0107 ( new_n279_, new_n274_, new_n278_ );
and g0108 ( new_n280_, new_n279_, new_n271_ );
and g0109 ( new_n281_, new_n223_, keyIn_0_18 );
and g0110 ( new_n282_, new_n218_, new_n211_ );
or g0111 ( new_n283_, new_n282_, new_n281_ );
not g0112 ( new_n284_, new_n231_ );
not g0113 ( new_n285_, N17 );
or g0114 ( new_n286_, keyIn_0_2, N11 );
not g0115 ( new_n287_, new_n235_ );
and g0116 ( new_n288_, new_n287_, new_n286_ );
or g0117 ( new_n289_, new_n288_, new_n285_ );
not g0118 ( new_n290_, new_n239_ );
and g0119 ( new_n291_, new_n289_, new_n290_ );
and g0120 ( new_n292_, new_n291_, new_n284_ );
and g0121 ( new_n293_, new_n283_, new_n292_ );
or g0122 ( new_n294_, new_n249_, keyIn_0_21 );
not g0123 ( new_n295_, new_n252_ );
and g0124 ( new_n296_, new_n295_, new_n294_ );
not g0125 ( new_n297_, new_n259_ );
and g0126 ( new_n298_, new_n297_, new_n255_ );
and g0127 ( new_n299_, new_n298_, keyIn_0_17 );
or g0128 ( new_n300_, new_n299_, new_n261_ );
and g0129 ( new_n301_, new_n296_, new_n300_ );
and g0130 ( new_n302_, new_n293_, new_n301_ );
and g0131 ( new_n303_, new_n302_, new_n280_ );
and g0132 ( new_n304_, new_n303_, new_n269_ );
or g0133 ( N223, new_n268_, new_n304_ );
not g0134 ( new_n306_, keyIn_0_80 );
not g0135 ( new_n307_, keyIn_0_71 );
not g0136 ( new_n308_, keyIn_0_43 );
not g0137 ( new_n309_, keyIn_0_37 );
and g0138 ( new_n310_, new_n303_, new_n309_ );
and g0139 ( new_n311_, new_n267_, keyIn_0_37 );
or g0140 ( new_n312_, new_n311_, new_n310_ );
and g0141 ( new_n313_, new_n312_, new_n290_ );
not g0142 ( new_n314_, new_n310_ );
or g0143 ( new_n315_, new_n303_, new_n309_ );
and g0144 ( new_n316_, new_n314_, new_n315_ );
and g0145 ( new_n317_, new_n316_, new_n239_ );
or g0146 ( new_n318_, new_n313_, new_n317_ );
not g0147 ( new_n319_, new_n318_ );
and g0148 ( new_n320_, new_n319_, new_n308_ );
and g0149 ( new_n321_, new_n318_, keyIn_0_43 );
or g0150 ( new_n322_, new_n320_, new_n321_ );
not g0151 ( new_n323_, N73 );
and g0152 ( new_n324_, new_n323_, N69 );
not g0153 ( new_n325_, new_n324_ );
and g0154 ( new_n326_, new_n325_, keyIn_0_29 );
not g0155 ( new_n327_, new_n326_ );
or g0156 ( new_n328_, new_n325_, keyIn_0_29 );
and g0157 ( new_n329_, new_n327_, new_n328_ );
and g0158 ( new_n330_, new_n322_, new_n329_ );
and g0159 ( new_n331_, new_n330_, keyIn_0_59 );
not g0160 ( new_n332_, new_n331_ );
or g0161 ( new_n333_, new_n330_, keyIn_0_59 );
and g0162 ( new_n334_, new_n332_, new_n333_ );
and g0163 ( new_n335_, new_n312_, new_n283_ );
and g0164 ( new_n336_, new_n316_, new_n225_ );
or g0165 ( new_n337_, new_n335_, new_n336_ );
and g0166 ( new_n338_, new_n337_, keyIn_0_41 );
not g0167 ( new_n339_, keyIn_0_41 );
or g0168 ( new_n340_, new_n316_, new_n225_ );
or g0169 ( new_n341_, new_n312_, new_n283_ );
and g0170 ( new_n342_, new_n341_, new_n340_ );
and g0171 ( new_n343_, new_n342_, new_n339_ );
or g0172 ( new_n344_, new_n338_, new_n343_ );
not g0173 ( new_n345_, N47 );
and g0174 ( new_n346_, new_n345_, N43 );
and g0175 ( new_n347_, new_n346_, keyIn_0_25 );
not g0176 ( new_n348_, new_n347_ );
or g0177 ( new_n349_, new_n346_, keyIn_0_25 );
and g0178 ( new_n350_, new_n348_, new_n349_ );
or g0179 ( new_n351_, new_n344_, new_n350_ );
or g0180 ( new_n352_, new_n351_, keyIn_0_58 );
not g0181 ( new_n353_, keyIn_0_58 );
or g0182 ( new_n354_, new_n342_, new_n339_ );
or g0183 ( new_n355_, new_n337_, keyIn_0_41 );
and g0184 ( new_n356_, new_n355_, new_n354_ );
not g0185 ( new_n357_, new_n350_ );
and g0186 ( new_n358_, new_n356_, new_n357_ );
or g0187 ( new_n359_, new_n358_, new_n353_ );
and g0188 ( new_n360_, new_n352_, new_n359_ );
not g0189 ( new_n361_, keyIn_0_47 );
and g0190 ( new_n362_, new_n312_, new_n296_ );
and g0191 ( new_n363_, new_n316_, new_n253_ );
or g0192 ( new_n364_, new_n362_, new_n363_ );
or g0193 ( new_n365_, new_n364_, new_n361_ );
or g0194 ( new_n366_, new_n316_, new_n253_ );
or g0195 ( new_n367_, new_n312_, new_n296_ );
and g0196 ( new_n368_, new_n367_, new_n366_ );
or g0197 ( new_n369_, new_n368_, keyIn_0_47 );
and g0198 ( new_n370_, new_n365_, new_n369_ );
not g0199 ( new_n371_, N112 );
and g0200 ( new_n372_, keyIn_0_13, N108 );
not g0201 ( new_n373_, new_n372_ );
or g0202 ( new_n374_, keyIn_0_13, N108 );
and g0203 ( new_n375_, new_n373_, new_n374_ );
not g0204 ( new_n376_, new_n375_ );
and g0205 ( new_n377_, new_n376_, new_n371_ );
and g0206 ( new_n378_, new_n377_, keyIn_0_35 );
not g0207 ( new_n379_, new_n378_ );
or g0208 ( new_n380_, new_n377_, keyIn_0_35 );
and g0209 ( new_n381_, new_n379_, new_n380_ );
or g0210 ( new_n382_, new_n370_, new_n381_ );
or g0211 ( new_n383_, new_n382_, keyIn_0_62 );
not g0212 ( new_n384_, keyIn_0_62 );
and g0213 ( new_n385_, new_n368_, keyIn_0_47 );
and g0214 ( new_n386_, new_n364_, new_n361_ );
or g0215 ( new_n387_, new_n386_, new_n385_ );
not g0216 ( new_n388_, new_n381_ );
and g0217 ( new_n389_, new_n387_, new_n388_ );
or g0218 ( new_n390_, new_n389_, new_n384_ );
and g0219 ( new_n391_, new_n383_, new_n390_ );
or g0220 ( new_n392_, new_n360_, new_n391_ );
or g0221 ( new_n393_, new_n392_, new_n334_ );
not g0222 ( new_n394_, keyIn_0_61 );
and g0223 ( new_n395_, new_n312_, new_n274_ );
and g0224 ( new_n396_, new_n316_, new_n197_ );
or g0225 ( new_n397_, new_n395_, new_n396_ );
or g0226 ( new_n398_, new_n397_, keyIn_0_45 );
not g0227 ( new_n399_, keyIn_0_45 );
or g0228 ( new_n400_, new_n316_, new_n197_ );
or g0229 ( new_n401_, new_n312_, new_n274_ );
and g0230 ( new_n402_, new_n401_, new_n400_ );
or g0231 ( new_n403_, new_n402_, new_n399_ );
and g0232 ( new_n404_, new_n398_, new_n403_ );
not g0233 ( new_n405_, keyIn_0_33 );
not g0234 ( new_n406_, N99 );
and g0235 ( new_n407_, new_n406_, N95 );
not g0236 ( new_n408_, new_n407_ );
and g0237 ( new_n409_, new_n408_, new_n405_ );
and g0238 ( new_n410_, new_n407_, keyIn_0_33 );
or g0239 ( new_n411_, new_n409_, new_n410_ );
or g0240 ( new_n412_, new_n404_, new_n411_ );
or g0241 ( new_n413_, new_n412_, new_n394_ );
and g0242 ( new_n414_, new_n402_, new_n399_ );
and g0243 ( new_n415_, new_n397_, keyIn_0_45 );
or g0244 ( new_n416_, new_n415_, new_n414_ );
not g0245 ( new_n417_, new_n411_ );
and g0246 ( new_n418_, new_n416_, new_n417_ );
or g0247 ( new_n419_, new_n418_, keyIn_0_61 );
and g0248 ( new_n420_, new_n413_, new_n419_ );
and g0249 ( new_n421_, new_n312_, new_n284_ );
and g0250 ( new_n422_, new_n316_, new_n231_ );
or g0251 ( new_n423_, new_n421_, new_n422_ );
not g0252 ( new_n424_, new_n423_ );
not g0253 ( new_n425_, N86 );
and g0254 ( new_n426_, keyIn_0_10, N82 );
not g0255 ( new_n427_, new_n426_ );
or g0256 ( new_n428_, keyIn_0_10, N82 );
and g0257 ( new_n429_, new_n427_, new_n428_ );
not g0258 ( new_n430_, new_n429_ );
and g0259 ( new_n431_, new_n430_, new_n425_ );
and g0260 ( new_n432_, new_n431_, keyIn_0_31 );
not g0261 ( new_n433_, new_n432_ );
or g0262 ( new_n434_, new_n431_, keyIn_0_31 );
and g0263 ( new_n435_, new_n433_, new_n434_ );
or g0264 ( new_n436_, new_n424_, new_n435_ );
not g0265 ( new_n437_, new_n436_ );
and g0266 ( new_n438_, new_n437_, keyIn_0_60 );
not g0267 ( new_n439_, keyIn_0_60 );
and g0268 ( new_n440_, new_n436_, new_n439_ );
or g0269 ( new_n441_, new_n438_, new_n440_ );
or g0270 ( new_n442_, new_n316_, new_n182_ );
and g0271 ( new_n443_, new_n182_, new_n309_ );
not g0272 ( new_n444_, new_n443_ );
and g0273 ( new_n445_, new_n442_, new_n444_ );
not g0274 ( new_n446_, keyIn_0_15 );
not g0275 ( new_n447_, N8 );
and g0276 ( new_n448_, keyIn_0_1, N4 );
not g0277 ( new_n449_, new_n448_ );
or g0278 ( new_n450_, keyIn_0_1, N4 );
and g0279 ( new_n451_, new_n449_, new_n450_ );
not g0280 ( new_n452_, new_n451_ );
and g0281 ( new_n453_, new_n452_, new_n447_ );
and g0282 ( new_n454_, new_n453_, new_n446_ );
not g0283 ( new_n455_, new_n454_ );
or g0284 ( new_n456_, new_n453_, new_n446_ );
and g0285 ( new_n457_, new_n455_, new_n456_ );
or g0286 ( new_n458_, new_n445_, new_n457_ );
and g0287 ( new_n459_, new_n458_, keyIn_0_54 );
not g0288 ( new_n460_, keyIn_0_54 );
and g0289 ( new_n461_, new_n312_, new_n271_ );
or g0290 ( new_n462_, new_n461_, new_n443_ );
not g0291 ( new_n463_, new_n457_ );
and g0292 ( new_n464_, new_n462_, new_n463_ );
and g0293 ( new_n465_, new_n464_, new_n460_ );
or g0294 ( new_n466_, new_n459_, new_n465_ );
not g0295 ( new_n467_, keyIn_0_42 );
and g0296 ( new_n468_, new_n312_, new_n278_ );
and g0297 ( new_n469_, new_n316_, new_n208_ );
or g0298 ( new_n470_, new_n468_, new_n469_ );
or g0299 ( new_n471_, new_n470_, new_n467_ );
or g0300 ( new_n472_, new_n316_, new_n208_ );
or g0301 ( new_n473_, new_n312_, new_n278_ );
and g0302 ( new_n474_, new_n473_, new_n472_ );
or g0303 ( new_n475_, new_n474_, keyIn_0_42 );
and g0304 ( new_n476_, new_n471_, new_n475_ );
not g0305 ( new_n477_, keyIn_0_27 );
not g0306 ( new_n478_, N60 );
and g0307 ( new_n479_, keyIn_0_8, N56 );
not g0308 ( new_n480_, new_n479_ );
or g0309 ( new_n481_, keyIn_0_8, N56 );
and g0310 ( new_n482_, new_n480_, new_n481_ );
not g0311 ( new_n483_, new_n482_ );
and g0312 ( new_n484_, new_n483_, new_n478_ );
and g0313 ( new_n485_, new_n484_, new_n477_ );
not g0314 ( new_n486_, new_n485_ );
or g0315 ( new_n487_, new_n484_, new_n477_ );
and g0316 ( new_n488_, new_n486_, new_n487_ );
not g0317 ( new_n489_, new_n488_ );
and g0318 ( new_n490_, new_n476_, new_n489_ );
or g0319 ( new_n491_, new_n466_, new_n490_ );
or g0320 ( new_n492_, new_n491_, new_n441_ );
or g0321 ( new_n493_, new_n492_, new_n420_ );
not g0322 ( new_n494_, keyIn_0_39 );
and g0323 ( new_n495_, new_n312_, new_n289_ );
and g0324 ( new_n496_, new_n316_, new_n237_ );
or g0325 ( new_n497_, new_n495_, new_n496_ );
or g0326 ( new_n498_, new_n497_, new_n494_ );
or g0327 ( new_n499_, new_n316_, new_n237_ );
or g0328 ( new_n500_, new_n312_, new_n289_ );
and g0329 ( new_n501_, new_n500_, new_n499_ );
or g0330 ( new_n502_, new_n501_, keyIn_0_39 );
and g0331 ( new_n503_, new_n498_, new_n502_ );
not g0332 ( new_n504_, keyIn_0_22 );
not g0333 ( new_n505_, N21 );
and g0334 ( new_n506_, new_n285_, keyIn_0_3 );
not g0335 ( new_n507_, new_n506_ );
or g0336 ( new_n508_, new_n285_, keyIn_0_3 );
and g0337 ( new_n509_, new_n507_, new_n508_ );
not g0338 ( new_n510_, new_n509_ );
and g0339 ( new_n511_, new_n510_, new_n505_ );
not g0340 ( new_n512_, new_n511_ );
and g0341 ( new_n513_, new_n512_, new_n504_ );
and g0342 ( new_n514_, new_n511_, keyIn_0_22 );
or g0343 ( new_n515_, new_n513_, new_n514_ );
or g0344 ( new_n516_, new_n503_, new_n515_ );
or g0345 ( new_n517_, new_n516_, keyIn_0_56 );
not g0346 ( new_n518_, keyIn_0_56 );
and g0347 ( new_n519_, new_n501_, keyIn_0_39 );
and g0348 ( new_n520_, new_n497_, new_n494_ );
or g0349 ( new_n521_, new_n520_, new_n519_ );
not g0350 ( new_n522_, new_n515_ );
and g0351 ( new_n523_, new_n521_, new_n522_ );
or g0352 ( new_n524_, new_n523_, new_n518_ );
and g0353 ( new_n525_, new_n517_, new_n524_ );
not g0354 ( new_n526_, keyIn_0_57 );
and g0355 ( new_n527_, new_n312_, new_n300_ );
and g0356 ( new_n528_, new_n264_, new_n309_ );
or g0357 ( new_n529_, new_n527_, new_n528_ );
and g0358 ( new_n530_, new_n529_, keyIn_0_40 );
not g0359 ( new_n531_, keyIn_0_40 );
or g0360 ( new_n532_, new_n316_, new_n264_ );
not g0361 ( new_n533_, new_n528_ );
and g0362 ( new_n534_, new_n532_, new_n533_ );
and g0363 ( new_n535_, new_n534_, new_n531_ );
or g0364 ( new_n536_, new_n530_, new_n535_ );
not g0365 ( new_n537_, N34 );
and g0366 ( new_n538_, new_n257_, keyIn_0_5 );
not g0367 ( new_n539_, new_n538_ );
or g0368 ( new_n540_, new_n257_, keyIn_0_5 );
and g0369 ( new_n541_, new_n539_, new_n540_ );
not g0370 ( new_n542_, new_n541_ );
and g0371 ( new_n543_, new_n542_, new_n537_ );
not g0372 ( new_n544_, new_n543_ );
and g0373 ( new_n545_, new_n544_, keyIn_0_23 );
not g0374 ( new_n546_, new_n545_ );
or g0375 ( new_n547_, new_n544_, keyIn_0_23 );
and g0376 ( new_n548_, new_n546_, new_n547_ );
or g0377 ( new_n549_, new_n536_, new_n548_ );
or g0378 ( new_n550_, new_n549_, new_n526_ );
or g0379 ( new_n551_, new_n534_, new_n531_ );
or g0380 ( new_n552_, new_n529_, keyIn_0_40 );
and g0381 ( new_n553_, new_n552_, new_n551_ );
not g0382 ( new_n554_, new_n548_ );
and g0383 ( new_n555_, new_n553_, new_n554_ );
or g0384 ( new_n556_, new_n555_, keyIn_0_57 );
and g0385 ( new_n557_, new_n550_, new_n556_ );
or g0386 ( new_n558_, new_n525_, new_n557_ );
or g0387 ( new_n559_, new_n493_, new_n558_ );
or g0388 ( new_n560_, new_n559_, new_n393_ );
and g0389 ( new_n561_, new_n560_, new_n307_ );
not g0390 ( new_n562_, new_n333_ );
or g0391 ( new_n563_, new_n562_, new_n331_ );
and g0392 ( new_n564_, new_n358_, new_n353_ );
and g0393 ( new_n565_, new_n351_, keyIn_0_58 );
or g0394 ( new_n566_, new_n565_, new_n564_ );
and g0395 ( new_n567_, new_n389_, new_n384_ );
and g0396 ( new_n568_, new_n382_, keyIn_0_62 );
or g0397 ( new_n569_, new_n568_, new_n567_ );
and g0398 ( new_n570_, new_n569_, new_n566_ );
and g0399 ( new_n571_, new_n570_, new_n563_ );
and g0400 ( new_n572_, new_n418_, keyIn_0_61 );
and g0401 ( new_n573_, new_n412_, new_n394_ );
or g0402 ( new_n574_, new_n573_, new_n572_ );
or g0403 ( new_n575_, new_n436_, new_n439_ );
not g0404 ( new_n576_, new_n440_ );
and g0405 ( new_n577_, new_n576_, new_n575_ );
or g0406 ( new_n578_, new_n464_, new_n460_ );
or g0407 ( new_n579_, new_n458_, keyIn_0_54 );
and g0408 ( new_n580_, new_n579_, new_n578_ );
and g0409 ( new_n581_, new_n474_, keyIn_0_42 );
and g0410 ( new_n582_, new_n470_, new_n467_ );
or g0411 ( new_n583_, new_n582_, new_n581_ );
or g0412 ( new_n584_, new_n583_, new_n488_ );
and g0413 ( new_n585_, new_n584_, new_n580_ );
and g0414 ( new_n586_, new_n585_, new_n577_ );
and g0415 ( new_n587_, new_n574_, new_n586_ );
and g0416 ( new_n588_, new_n523_, new_n518_ );
and g0417 ( new_n589_, new_n516_, keyIn_0_56 );
or g0418 ( new_n590_, new_n589_, new_n588_ );
and g0419 ( new_n591_, new_n555_, keyIn_0_57 );
and g0420 ( new_n592_, new_n549_, new_n526_ );
or g0421 ( new_n593_, new_n592_, new_n591_ );
and g0422 ( new_n594_, new_n590_, new_n593_ );
and g0423 ( new_n595_, new_n587_, new_n594_ );
and g0424 ( new_n596_, new_n595_, new_n571_ );
and g0425 ( new_n597_, new_n596_, keyIn_0_71 );
or g0426 ( new_n598_, new_n561_, new_n597_ );
and g0427 ( new_n599_, new_n598_, new_n306_ );
or g0428 ( new_n600_, new_n596_, keyIn_0_71 );
not g0429 ( new_n601_, new_n597_ );
and g0430 ( new_n602_, new_n601_, new_n600_ );
and g0431 ( new_n603_, new_n602_, keyIn_0_80 );
or g0432 ( N329, new_n599_, new_n603_ );
not g0433 ( new_n605_, keyIn_0_83 );
and g0434 ( new_n606_, new_n598_, keyIn_0_78 );
not g0435 ( new_n607_, keyIn_0_78 );
and g0436 ( new_n608_, new_n602_, new_n607_ );
or g0437 ( new_n609_, new_n606_, new_n608_ );
and g0438 ( new_n610_, new_n609_, new_n584_ );
or g0439 ( new_n611_, new_n602_, new_n607_ );
or g0440 ( new_n612_, new_n598_, keyIn_0_78 );
and g0441 ( new_n613_, new_n612_, new_n611_ );
and g0442 ( new_n614_, new_n613_, new_n490_ );
or g0443 ( new_n615_, new_n610_, new_n614_ );
and g0444 ( new_n616_, new_n615_, new_n605_ );
not g0445 ( new_n617_, new_n616_ );
or g0446 ( new_n618_, new_n615_, new_n605_ );
and g0447 ( new_n619_, new_n617_, new_n618_ );
not g0448 ( new_n620_, keyIn_0_66 );
not g0449 ( new_n621_, N66 );
and g0450 ( new_n622_, new_n483_, new_n621_ );
and g0451 ( new_n623_, new_n622_, keyIn_0_28 );
not g0452 ( new_n624_, new_n623_ );
or g0453 ( new_n625_, new_n622_, keyIn_0_28 );
and g0454 ( new_n626_, new_n624_, new_n625_ );
or g0455 ( new_n627_, new_n583_, new_n626_ );
and g0456 ( new_n628_, new_n627_, new_n620_ );
not g0457 ( new_n629_, new_n628_ );
or g0458 ( new_n630_, new_n627_, new_n620_ );
and g0459 ( new_n631_, new_n629_, new_n630_ );
or g0460 ( new_n632_, new_n619_, new_n631_ );
not g0461 ( new_n633_, keyIn_0_86 );
and g0462 ( new_n634_, new_n609_, new_n577_ );
and g0463 ( new_n635_, new_n613_, new_n441_ );
or g0464 ( new_n636_, new_n634_, new_n635_ );
not g0465 ( new_n637_, new_n636_ );
and g0466 ( new_n638_, new_n637_, new_n633_ );
and g0467 ( new_n639_, new_n636_, keyIn_0_86 );
or g0468 ( new_n640_, new_n638_, new_n639_ );
not g0469 ( new_n641_, N92 );
and g0470 ( new_n642_, new_n430_, new_n641_ );
and g0471 ( new_n643_, new_n642_, keyIn_0_32 );
not g0472 ( new_n644_, new_n643_ );
or g0473 ( new_n645_, new_n642_, keyIn_0_32 );
and g0474 ( new_n646_, new_n644_, new_n645_ );
or g0475 ( new_n647_, new_n424_, new_n646_ );
and g0476 ( new_n648_, new_n647_, keyIn_0_68 );
not g0477 ( new_n649_, new_n648_ );
or g0478 ( new_n650_, new_n647_, keyIn_0_68 );
and g0479 ( new_n651_, new_n649_, new_n650_ );
not g0480 ( new_n652_, new_n651_ );
and g0481 ( new_n653_, new_n652_, keyIn_0_75 );
not g0482 ( new_n654_, new_n653_ );
or g0483 ( new_n655_, new_n652_, keyIn_0_75 );
and g0484 ( new_n656_, new_n654_, new_n655_ );
not g0485 ( new_n657_, new_n656_ );
and g0486 ( new_n658_, new_n640_, new_n657_ );
not g0487 ( new_n659_, new_n658_ );
and g0488 ( new_n660_, new_n659_, new_n632_ );
not g0489 ( new_n661_, keyIn_0_95 );
and g0490 ( new_n662_, new_n609_, new_n593_ );
and g0491 ( new_n663_, new_n613_, new_n557_ );
or g0492 ( new_n664_, new_n662_, new_n663_ );
not g0493 ( new_n665_, keyIn_0_64 );
not g0494 ( new_n666_, N40 );
and g0495 ( new_n667_, new_n542_, new_n666_ );
not g0496 ( new_n668_, new_n667_ );
and g0497 ( new_n669_, new_n668_, keyIn_0_24 );
not g0498 ( new_n670_, new_n669_ );
or g0499 ( new_n671_, new_n668_, keyIn_0_24 );
and g0500 ( new_n672_, new_n670_, new_n671_ );
or g0501 ( new_n673_, new_n536_, new_n672_ );
not g0502 ( new_n674_, new_n673_ );
and g0503 ( new_n675_, new_n674_, new_n665_ );
and g0504 ( new_n676_, new_n673_, keyIn_0_64 );
or g0505 ( new_n677_, new_n675_, new_n676_ );
and g0506 ( new_n678_, new_n677_, keyIn_0_73 );
not g0507 ( new_n679_, new_n678_ );
or g0508 ( new_n680_, new_n677_, keyIn_0_73 );
and g0509 ( new_n681_, new_n679_, new_n680_ );
not g0510 ( new_n682_, new_n681_ );
and g0511 ( new_n683_, new_n664_, new_n682_ );
not g0512 ( new_n684_, new_n683_ );
and g0513 ( new_n685_, new_n684_, new_n661_ );
and g0514 ( new_n686_, new_n683_, keyIn_0_95 );
or g0515 ( new_n687_, new_n685_, new_n686_ );
and g0516 ( new_n688_, new_n609_, new_n566_ );
and g0517 ( new_n689_, new_n613_, new_n360_ );
or g0518 ( new_n690_, new_n688_, new_n689_ );
not g0519 ( new_n691_, keyIn_0_65 );
not g0520 ( new_n692_, keyIn_0_26 );
not g0521 ( new_n693_, N53 );
and g0522 ( new_n694_, new_n693_, N43 );
and g0523 ( new_n695_, new_n694_, new_n692_ );
not g0524 ( new_n696_, new_n695_ );
or g0525 ( new_n697_, new_n694_, new_n692_ );
and g0526 ( new_n698_, new_n696_, new_n697_ );
or g0527 ( new_n699_, new_n344_, new_n698_ );
not g0528 ( new_n700_, new_n699_ );
and g0529 ( new_n701_, new_n700_, new_n691_ );
and g0530 ( new_n702_, new_n699_, keyIn_0_65 );
or g0531 ( new_n703_, new_n701_, new_n702_ );
and g0532 ( new_n704_, new_n690_, new_n703_ );
not g0533 ( new_n705_, new_n704_ );
and g0534 ( new_n706_, new_n705_, keyIn_0_96 );
or g0535 ( new_n707_, new_n705_, keyIn_0_96 );
not g0536 ( new_n708_, new_n707_ );
or g0537 ( new_n709_, new_n708_, new_n706_ );
and g0538 ( new_n710_, new_n709_, new_n687_ );
and g0539 ( new_n711_, new_n710_, new_n660_ );
and g0540 ( new_n712_, new_n609_, new_n590_ );
and g0541 ( new_n713_, new_n613_, new_n525_ );
or g0542 ( new_n714_, new_n712_, new_n713_ );
not g0543 ( new_n715_, new_n714_ );
and g0544 ( new_n716_, new_n715_, keyIn_0_82 );
not g0545 ( new_n717_, new_n716_ );
or g0546 ( new_n718_, new_n715_, keyIn_0_82 );
not g0547 ( new_n719_, keyIn_0_63 );
not g0548 ( new_n720_, N27 );
and g0549 ( new_n721_, new_n510_, new_n720_ );
and g0550 ( new_n722_, new_n521_, new_n721_ );
not g0551 ( new_n723_, new_n722_ );
and g0552 ( new_n724_, new_n723_, new_n719_ );
and g0553 ( new_n725_, new_n722_, keyIn_0_63 );
or g0554 ( new_n726_, new_n724_, new_n725_ );
and g0555 ( new_n727_, new_n718_, new_n726_ );
and g0556 ( new_n728_, new_n727_, new_n717_ );
or g0557 ( new_n729_, new_n728_, keyIn_0_94 );
and g0558 ( new_n730_, new_n728_, keyIn_0_94 );
not g0559 ( new_n731_, new_n730_ );
and g0560 ( new_n732_, new_n731_, new_n729_ );
and g0561 ( new_n733_, new_n711_, new_n732_ );
not g0562 ( new_n734_, new_n733_ );
not g0563 ( new_n735_, keyIn_0_98 );
and g0564 ( new_n736_, new_n609_, new_n574_ );
and g0565 ( new_n737_, new_n613_, new_n420_ );
or g0566 ( new_n738_, new_n736_, new_n737_ );
or g0567 ( new_n739_, new_n738_, keyIn_0_88 );
not g0568 ( new_n740_, keyIn_0_88 );
or g0569 ( new_n741_, new_n613_, new_n420_ );
or g0570 ( new_n742_, new_n609_, new_n574_ );
and g0571 ( new_n743_, new_n742_, new_n741_ );
or g0572 ( new_n744_, new_n743_, new_n740_ );
and g0573 ( new_n745_, new_n739_, new_n744_ );
not g0574 ( new_n746_, keyIn_0_76 );
not g0575 ( new_n747_, keyIn_0_34 );
not g0576 ( new_n748_, N105 );
and g0577 ( new_n749_, new_n748_, N95 );
and g0578 ( new_n750_, new_n749_, new_n747_ );
not g0579 ( new_n751_, new_n750_ );
or g0580 ( new_n752_, new_n749_, new_n747_ );
and g0581 ( new_n753_, new_n751_, new_n752_ );
and g0582 ( new_n754_, new_n416_, new_n753_ );
not g0583 ( new_n755_, new_n754_ );
and g0584 ( new_n756_, new_n755_, keyIn_0_69 );
not g0585 ( new_n757_, new_n756_ );
or g0586 ( new_n758_, new_n755_, keyIn_0_69 );
and g0587 ( new_n759_, new_n757_, new_n758_ );
and g0588 ( new_n760_, new_n759_, new_n746_ );
not g0589 ( new_n761_, new_n760_ );
or g0590 ( new_n762_, new_n759_, new_n746_ );
and g0591 ( new_n763_, new_n761_, new_n762_ );
or g0592 ( new_n764_, new_n745_, new_n763_ );
or g0593 ( new_n765_, new_n764_, new_n735_ );
and g0594 ( new_n766_, new_n743_, new_n740_ );
and g0595 ( new_n767_, new_n738_, keyIn_0_88 );
or g0596 ( new_n768_, new_n767_, new_n766_ );
not g0597 ( new_n769_, new_n763_ );
and g0598 ( new_n770_, new_n768_, new_n769_ );
or g0599 ( new_n771_, new_n770_, keyIn_0_98 );
and g0600 ( new_n772_, new_n765_, new_n771_ );
not g0601 ( new_n773_, keyIn_0_90 );
and g0602 ( new_n774_, new_n609_, new_n569_ );
and g0603 ( new_n775_, new_n613_, new_n391_ );
or g0604 ( new_n776_, new_n774_, new_n775_ );
or g0605 ( new_n777_, new_n776_, new_n773_ );
or g0606 ( new_n778_, new_n613_, new_n391_ );
or g0607 ( new_n779_, new_n609_, new_n569_ );
and g0608 ( new_n780_, new_n779_, new_n778_ );
or g0609 ( new_n781_, new_n780_, keyIn_0_90 );
and g0610 ( new_n782_, new_n777_, new_n781_ );
not g0611 ( new_n783_, keyIn_0_77 );
not g0612 ( new_n784_, keyIn_0_70 );
not g0613 ( new_n785_, keyIn_0_36 );
not g0614 ( new_n786_, N115 );
and g0615 ( new_n787_, new_n376_, new_n786_ );
and g0616 ( new_n788_, new_n787_, new_n785_ );
not g0617 ( new_n789_, new_n788_ );
or g0618 ( new_n790_, new_n787_, new_n785_ );
and g0619 ( new_n791_, new_n789_, new_n790_ );
or g0620 ( new_n792_, new_n370_, new_n791_ );
and g0621 ( new_n793_, new_n792_, new_n784_ );
not g0622 ( new_n794_, new_n793_ );
or g0623 ( new_n795_, new_n792_, new_n784_ );
and g0624 ( new_n796_, new_n794_, new_n795_ );
and g0625 ( new_n797_, new_n796_, new_n783_ );
not g0626 ( new_n798_, new_n797_ );
or g0627 ( new_n799_, new_n796_, new_n783_ );
and g0628 ( new_n800_, new_n798_, new_n799_ );
or g0629 ( new_n801_, new_n782_, new_n800_ );
or g0630 ( new_n802_, new_n801_, keyIn_0_99 );
not g0631 ( new_n803_, keyIn_0_99 );
and g0632 ( new_n804_, new_n780_, keyIn_0_90 );
and g0633 ( new_n805_, new_n776_, new_n773_ );
or g0634 ( new_n806_, new_n805_, new_n804_ );
not g0635 ( new_n807_, new_n800_ );
and g0636 ( new_n808_, new_n806_, new_n807_ );
or g0637 ( new_n809_, new_n808_, new_n803_ );
and g0638 ( new_n810_, new_n802_, new_n809_ );
or g0639 ( new_n811_, new_n772_, new_n810_ );
not g0640 ( new_n812_, keyIn_0_93 );
or g0641 ( new_n813_, new_n613_, new_n466_ );
or g0642 ( new_n814_, new_n609_, new_n580_ );
and g0643 ( new_n815_, new_n814_, new_n813_ );
and g0644 ( new_n816_, new_n815_, keyIn_0_81 );
not g0645 ( new_n817_, keyIn_0_81 );
and g0646 ( new_n818_, new_n609_, new_n580_ );
and g0647 ( new_n819_, new_n613_, new_n466_ );
or g0648 ( new_n820_, new_n818_, new_n819_ );
and g0649 ( new_n821_, new_n820_, new_n817_ );
not g0650 ( new_n822_, keyIn_0_16 );
not g0651 ( new_n823_, N14 );
and g0652 ( new_n824_, new_n452_, new_n823_ );
and g0653 ( new_n825_, new_n824_, new_n822_ );
not g0654 ( new_n826_, new_n825_ );
or g0655 ( new_n827_, new_n824_, new_n822_ );
and g0656 ( new_n828_, new_n826_, new_n827_ );
or g0657 ( new_n829_, new_n445_, new_n828_ );
and g0658 ( new_n830_, new_n829_, keyIn_0_55 );
not g0659 ( new_n831_, new_n830_ );
or g0660 ( new_n832_, new_n829_, keyIn_0_55 );
and g0661 ( new_n833_, new_n831_, new_n832_ );
not g0662 ( new_n834_, new_n833_ );
and g0663 ( new_n835_, new_n834_, keyIn_0_72 );
not g0664 ( new_n836_, new_n835_ );
or g0665 ( new_n837_, new_n834_, keyIn_0_72 );
and g0666 ( new_n838_, new_n836_, new_n837_ );
or g0667 ( new_n839_, new_n821_, new_n838_ );
or g0668 ( new_n840_, new_n839_, new_n816_ );
or g0669 ( new_n841_, new_n840_, new_n812_ );
not g0670 ( new_n842_, new_n816_ );
or g0671 ( new_n843_, new_n815_, keyIn_0_81 );
not g0672 ( new_n844_, new_n838_ );
and g0673 ( new_n845_, new_n843_, new_n844_ );
and g0674 ( new_n846_, new_n845_, new_n842_ );
or g0675 ( new_n847_, new_n846_, keyIn_0_93 );
and g0676 ( new_n848_, new_n841_, new_n847_ );
or g0677 ( new_n849_, new_n613_, new_n334_ );
or g0678 ( new_n850_, new_n609_, new_n563_ );
and g0679 ( new_n851_, new_n850_, new_n849_ );
and g0680 ( new_n852_, new_n851_, keyIn_0_85 );
not g0681 ( new_n853_, keyIn_0_85 );
and g0682 ( new_n854_, new_n609_, new_n563_ );
and g0683 ( new_n855_, new_n613_, new_n334_ );
or g0684 ( new_n856_, new_n854_, new_n855_ );
and g0685 ( new_n857_, new_n856_, new_n853_ );
not g0686 ( new_n858_, keyIn_0_67 );
not g0687 ( new_n859_, keyIn_0_30 );
not g0688 ( new_n860_, N79 );
and g0689 ( new_n861_, new_n860_, N69 );
and g0690 ( new_n862_, new_n861_, new_n859_ );
not g0691 ( new_n863_, new_n862_ );
or g0692 ( new_n864_, new_n861_, new_n859_ );
and g0693 ( new_n865_, new_n863_, new_n864_ );
and g0694 ( new_n866_, new_n322_, new_n865_ );
not g0695 ( new_n867_, new_n866_ );
and g0696 ( new_n868_, new_n867_, new_n858_ );
and g0697 ( new_n869_, new_n866_, keyIn_0_67 );
or g0698 ( new_n870_, new_n868_, new_n869_ );
and g0699 ( new_n871_, new_n870_, keyIn_0_74 );
not g0700 ( new_n872_, new_n871_ );
or g0701 ( new_n873_, new_n870_, keyIn_0_74 );
and g0702 ( new_n874_, new_n872_, new_n873_ );
or g0703 ( new_n875_, new_n857_, new_n874_ );
or g0704 ( new_n876_, new_n875_, new_n852_ );
or g0705 ( new_n877_, new_n876_, keyIn_0_97 );
not g0706 ( new_n878_, keyIn_0_97 );
not g0707 ( new_n879_, new_n852_ );
or g0708 ( new_n880_, new_n851_, keyIn_0_85 );
not g0709 ( new_n881_, new_n874_ );
and g0710 ( new_n882_, new_n880_, new_n881_ );
and g0711 ( new_n883_, new_n882_, new_n879_ );
or g0712 ( new_n884_, new_n883_, new_n878_ );
and g0713 ( new_n885_, new_n877_, new_n884_ );
or g0714 ( new_n886_, new_n848_, new_n885_ );
or g0715 ( new_n887_, new_n811_, new_n886_ );
or g0716 ( N370, new_n887_, new_n734_ );
not g0717 ( new_n889_, keyIn_0_120 );
not g0718 ( new_n890_, keyIn_0_115 );
not g0719 ( new_n891_, keyIn_0_106 );
not g0720 ( new_n892_, keyIn_0_100 );
and g0721 ( new_n893_, new_n770_, keyIn_0_98 );
and g0722 ( new_n894_, new_n764_, new_n735_ );
or g0723 ( new_n895_, new_n894_, new_n893_ );
and g0724 ( new_n896_, new_n808_, new_n803_ );
and g0725 ( new_n897_, new_n801_, keyIn_0_99 );
or g0726 ( new_n898_, new_n897_, new_n896_ );
and g0727 ( new_n899_, new_n895_, new_n898_ );
and g0728 ( new_n900_, new_n846_, keyIn_0_93 );
and g0729 ( new_n901_, new_n840_, new_n812_ );
or g0730 ( new_n902_, new_n901_, new_n900_ );
and g0731 ( new_n903_, new_n883_, new_n878_ );
and g0732 ( new_n904_, new_n876_, keyIn_0_97 );
or g0733 ( new_n905_, new_n904_, new_n903_ );
and g0734 ( new_n906_, new_n902_, new_n905_ );
and g0735 ( new_n907_, new_n899_, new_n906_ );
and g0736 ( new_n908_, new_n907_, new_n733_ );
and g0737 ( new_n909_, new_n908_, new_n892_ );
and g0738 ( new_n910_, N370, keyIn_0_100 );
or g0739 ( new_n911_, new_n910_, new_n909_ );
or g0740 ( new_n912_, new_n911_, new_n860_ );
or g0741 ( new_n913_, new_n912_, new_n891_ );
not g0742 ( new_n914_, new_n909_ );
or g0743 ( new_n915_, new_n908_, new_n892_ );
and g0744 ( new_n916_, new_n914_, new_n915_ );
and g0745 ( new_n917_, new_n916_, N79 );
or g0746 ( new_n918_, new_n917_, keyIn_0_106 );
and g0747 ( new_n919_, new_n913_, new_n918_ );
and g0748 ( new_n920_, new_n598_, keyIn_0_79 );
not g0749 ( new_n921_, new_n920_ );
or g0750 ( new_n922_, new_n598_, keyIn_0_79 );
and g0751 ( new_n923_, new_n921_, new_n922_ );
not g0752 ( new_n924_, new_n923_ );
and g0753 ( new_n925_, new_n924_, N73 );
and g0754 ( new_n926_, new_n925_, keyIn_0_91 );
not g0755 ( new_n927_, new_n926_ );
or g0756 ( new_n928_, new_n925_, keyIn_0_91 );
and g0757 ( new_n929_, new_n267_, N63 );
and g0758 ( new_n930_, new_n929_, keyIn_0_50 );
not g0759 ( new_n931_, new_n930_ );
or g0760 ( new_n932_, new_n929_, keyIn_0_50 );
and g0761 ( new_n933_, new_n932_, N69 );
and g0762 ( new_n934_, new_n933_, new_n931_ );
and g0763 ( new_n935_, new_n928_, new_n934_ );
and g0764 ( new_n936_, new_n935_, new_n927_ );
not g0765 ( new_n937_, new_n936_ );
or g0766 ( new_n938_, new_n919_, new_n937_ );
or g0767 ( new_n939_, new_n938_, keyIn_0_113 );
not g0768 ( new_n940_, keyIn_0_113 );
and g0769 ( new_n941_, new_n917_, keyIn_0_106 );
and g0770 ( new_n942_, new_n912_, new_n891_ );
or g0771 ( new_n943_, new_n942_, new_n941_ );
and g0772 ( new_n944_, new_n943_, new_n936_ );
or g0773 ( new_n945_, new_n944_, new_n940_ );
and g0774 ( new_n946_, new_n939_, new_n945_ );
not g0775 ( new_n947_, keyIn_0_107 );
and g0776 ( new_n948_, new_n916_, N92 );
and g0777 ( new_n949_, new_n948_, new_n947_ );
not g0778 ( new_n950_, new_n949_ );
or g0779 ( new_n951_, new_n948_, new_n947_ );
and g0780 ( new_n952_, new_n950_, new_n951_ );
and g0781 ( new_n953_, new_n924_, N86 );
not g0782 ( new_n954_, N82 );
not g0783 ( new_n955_, keyIn_0_51 );
and g0784 ( new_n956_, new_n267_, N76 );
and g0785 ( new_n957_, new_n956_, new_n955_ );
not g0786 ( new_n958_, new_n957_ );
or g0787 ( new_n959_, new_n956_, new_n955_ );
and g0788 ( new_n960_, new_n958_, new_n959_ );
or g0789 ( new_n961_, new_n960_, new_n954_ );
or g0790 ( new_n962_, new_n953_, new_n961_ );
or g0791 ( new_n963_, new_n952_, new_n962_ );
not g0792 ( new_n964_, new_n963_ );
and g0793 ( new_n965_, new_n964_, keyIn_0_114 );
not g0794 ( new_n966_, keyIn_0_114 );
and g0795 ( new_n967_, new_n963_, new_n966_ );
or g0796 ( new_n968_, new_n965_, new_n967_ );
and g0797 ( new_n969_, new_n916_, N105 );
and g0798 ( new_n970_, new_n969_, keyIn_0_108 );
not g0799 ( new_n971_, new_n970_ );
or g0800 ( new_n972_, new_n969_, keyIn_0_108 );
and g0801 ( new_n973_, new_n971_, new_n972_ );
not g0802 ( new_n974_, new_n973_ );
and g0803 ( new_n975_, new_n924_, N99 );
and g0804 ( new_n976_, new_n975_, keyIn_0_92 );
not g0805 ( new_n977_, new_n976_ );
or g0806 ( new_n978_, new_n975_, keyIn_0_92 );
not g0807 ( new_n979_, keyIn_0_52 );
and g0808 ( new_n980_, new_n267_, N89 );
and g0809 ( new_n981_, new_n980_, new_n979_ );
not g0810 ( new_n982_, new_n981_ );
or g0811 ( new_n983_, new_n980_, new_n979_ );
and g0812 ( new_n984_, new_n983_, N95 );
and g0813 ( new_n985_, new_n984_, new_n982_ );
and g0814 ( new_n986_, new_n978_, new_n985_ );
and g0815 ( new_n987_, new_n986_, new_n977_ );
and g0816 ( new_n988_, new_n974_, new_n987_ );
not g0817 ( new_n989_, new_n988_ );
and g0818 ( new_n990_, new_n916_, N115 );
and g0819 ( new_n991_, new_n924_, N112 );
and g0820 ( new_n992_, new_n267_, N102 );
and g0821 ( new_n993_, new_n992_, keyIn_0_53 );
not g0822 ( new_n994_, new_n993_ );
or g0823 ( new_n995_, new_n992_, keyIn_0_53 );
and g0824 ( new_n996_, new_n994_, new_n995_ );
or g0825 ( new_n997_, new_n996_, new_n246_ );
or g0826 ( new_n998_, new_n991_, new_n997_ );
or g0827 ( new_n999_, new_n990_, new_n998_ );
and g0828 ( new_n1000_, new_n989_, new_n999_ );
and g0829 ( new_n1001_, new_n968_, new_n1000_ );
and g0830 ( new_n1002_, new_n1001_, new_n946_ );
not g0831 ( new_n1003_, keyIn_0_102 );
and g0832 ( new_n1004_, new_n916_, N27 );
and g0833 ( new_n1005_, new_n1004_, new_n1003_ );
not g0834 ( new_n1006_, new_n1005_ );
or g0835 ( new_n1007_, new_n1004_, new_n1003_ );
and g0836 ( new_n1008_, new_n1006_, new_n1007_ );
not g0837 ( new_n1009_, new_n1008_ );
not g0838 ( new_n1010_, keyIn_0_84 );
and g0839 ( new_n1011_, new_n924_, N21 );
and g0840 ( new_n1012_, new_n1011_, new_n1010_ );
not g0841 ( new_n1013_, new_n1012_ );
or g0842 ( new_n1014_, new_n1011_, new_n1010_ );
and g0843 ( new_n1015_, new_n267_, N11 );
or g0844 ( new_n1016_, new_n1015_, new_n285_ );
not g0845 ( new_n1017_, new_n1016_ );
and g0846 ( new_n1018_, new_n1014_, new_n1017_ );
and g0847 ( new_n1019_, new_n1018_, new_n1013_ );
and g0848 ( new_n1020_, new_n1009_, new_n1019_ );
not g0849 ( new_n1021_, new_n1020_ );
and g0850 ( new_n1022_, new_n1021_, keyIn_0_110 );
not g0851 ( new_n1023_, keyIn_0_110 );
and g0852 ( new_n1024_, new_n1020_, new_n1023_ );
or g0853 ( new_n1025_, new_n1022_, new_n1024_ );
or g0854 ( new_n1026_, new_n911_, new_n666_ );
or g0855 ( new_n1027_, new_n1026_, keyIn_0_103 );
not g0856 ( new_n1028_, keyIn_0_103 );
and g0857 ( new_n1029_, new_n916_, N40 );
or g0858 ( new_n1030_, new_n1029_, new_n1028_ );
and g0859 ( new_n1031_, new_n1027_, new_n1030_ );
and g0860 ( new_n1032_, new_n924_, N34 );
not g0861 ( new_n1033_, new_n1032_ );
not g0862 ( new_n1034_, keyIn_0_46 );
and g0863 ( new_n1035_, new_n267_, N24 );
and g0864 ( new_n1036_, new_n1035_, new_n1034_ );
not g0865 ( new_n1037_, new_n1036_ );
or g0866 ( new_n1038_, new_n1035_, new_n1034_ );
and g0867 ( new_n1039_, new_n1038_, N30 );
and g0868 ( new_n1040_, new_n1039_, new_n1037_ );
and g0869 ( new_n1041_, new_n1033_, new_n1040_ );
not g0870 ( new_n1042_, new_n1041_ );
or g0871 ( new_n1043_, new_n1031_, new_n1042_ );
or g0872 ( new_n1044_, new_n1043_, keyIn_0_111 );
not g0873 ( new_n1045_, keyIn_0_111 );
and g0874 ( new_n1046_, new_n1029_, new_n1028_ );
and g0875 ( new_n1047_, new_n1026_, keyIn_0_103 );
or g0876 ( new_n1048_, new_n1047_, new_n1046_ );
and g0877 ( new_n1049_, new_n1048_, new_n1041_ );
or g0878 ( new_n1050_, new_n1049_, new_n1045_ );
and g0879 ( new_n1051_, new_n1044_, new_n1050_ );
and g0880 ( new_n1052_, new_n1025_, new_n1051_ );
not g0881 ( new_n1053_, keyIn_0_112 );
not g0882 ( new_n1054_, keyIn_0_105 );
and g0883 ( new_n1055_, new_n916_, N66 );
and g0884 ( new_n1056_, new_n1055_, new_n1054_ );
not g0885 ( new_n1057_, new_n1056_ );
or g0886 ( new_n1058_, new_n1055_, new_n1054_ );
and g0887 ( new_n1059_, new_n924_, N60 );
and g0888 ( new_n1060_, new_n1059_, keyIn_0_89 );
not g0889 ( new_n1061_, new_n1060_ );
or g0890 ( new_n1062_, new_n1059_, keyIn_0_89 );
not g0891 ( new_n1063_, keyIn_0_49 );
and g0892 ( new_n1064_, new_n267_, N50 );
not g0893 ( new_n1065_, new_n1064_ );
and g0894 ( new_n1066_, new_n1065_, new_n1063_ );
and g0895 ( new_n1067_, new_n1064_, keyIn_0_49 );
or g0896 ( new_n1068_, new_n1067_, new_n201_ );
or g0897 ( new_n1069_, new_n1068_, new_n1066_ );
not g0898 ( new_n1070_, new_n1069_ );
and g0899 ( new_n1071_, new_n1062_, new_n1070_ );
and g0900 ( new_n1072_, new_n1071_, new_n1061_ );
and g0901 ( new_n1073_, new_n1058_, new_n1072_ );
and g0902 ( new_n1074_, new_n1073_, new_n1057_ );
and g0903 ( new_n1075_, new_n1074_, new_n1053_ );
not g0904 ( new_n1076_, new_n1075_ );
or g0905 ( new_n1077_, new_n1074_, new_n1053_ );
and g0906 ( new_n1078_, new_n1076_, new_n1077_ );
not g0907 ( new_n1079_, new_n1078_ );
not g0908 ( new_n1080_, keyIn_0_104 );
and g0909 ( new_n1081_, new_n916_, N53 );
not g0910 ( new_n1082_, new_n1081_ );
and g0911 ( new_n1083_, new_n1082_, new_n1080_ );
and g0912 ( new_n1084_, new_n1081_, keyIn_0_104 );
or g0913 ( new_n1085_, new_n1083_, new_n1084_ );
and g0914 ( new_n1086_, new_n924_, N47 );
and g0915 ( new_n1087_, new_n1086_, keyIn_0_87 );
not g0916 ( new_n1088_, new_n1087_ );
or g0917 ( new_n1089_, new_n1086_, keyIn_0_87 );
not g0918 ( new_n1090_, keyIn_0_48 );
and g0919 ( new_n1091_, new_n267_, N37 );
and g0920 ( new_n1092_, new_n1091_, new_n1090_ );
not g0921 ( new_n1093_, new_n1092_ );
or g0922 ( new_n1094_, new_n1091_, new_n1090_ );
and g0923 ( new_n1095_, new_n1094_, N43 );
and g0924 ( new_n1096_, new_n1095_, new_n1093_ );
and g0925 ( new_n1097_, new_n1089_, new_n1096_ );
and g0926 ( new_n1098_, new_n1097_, new_n1088_ );
and g0927 ( new_n1099_, new_n1085_, new_n1098_ );
not g0928 ( new_n1100_, new_n1099_ );
and g0929 ( new_n1101_, new_n1079_, new_n1100_ );
and g0930 ( new_n1102_, new_n1052_, new_n1101_ );
and g0931 ( new_n1103_, new_n1102_, new_n1002_ );
and g0932 ( new_n1104_, new_n1103_, new_n890_ );
not g0933 ( new_n1105_, new_n1104_ );
or g0934 ( new_n1106_, new_n1103_, new_n890_ );
and g0935 ( new_n1107_, new_n1105_, new_n1106_ );
and g0936 ( new_n1108_, new_n916_, N14 );
and g0937 ( new_n1109_, new_n1108_, keyIn_0_101 );
not g0938 ( new_n1110_, new_n1109_ );
or g0939 ( new_n1111_, new_n1108_, keyIn_0_101 );
and g0940 ( new_n1112_, new_n924_, N8 );
not g0941 ( new_n1113_, new_n1112_ );
and g0942 ( new_n1114_, new_n267_, N1 );
and g0943 ( new_n1115_, new_n1114_, keyIn_0_44 );
not g0944 ( new_n1116_, new_n1115_ );
or g0945 ( new_n1117_, new_n1114_, keyIn_0_44 );
and g0946 ( new_n1118_, new_n1117_, N4 );
and g0947 ( new_n1119_, new_n1118_, new_n1116_ );
and g0948 ( new_n1120_, new_n1113_, new_n1119_ );
and g0949 ( new_n1121_, new_n1111_, new_n1120_ );
and g0950 ( new_n1122_, new_n1121_, new_n1110_ );
not g0951 ( new_n1123_, new_n1122_ );
and g0952 ( new_n1124_, new_n1123_, keyIn_0_109 );
not g0953 ( new_n1125_, new_n1124_ );
or g0954 ( new_n1126_, new_n1123_, keyIn_0_109 );
and g0955 ( new_n1127_, new_n1125_, new_n1126_ );
or g0956 ( new_n1128_, new_n1107_, new_n1127_ );
or g0957 ( new_n1129_, new_n1128_, new_n889_ );
not g0958 ( new_n1130_, new_n1103_ );
and g0959 ( new_n1131_, new_n1130_, keyIn_0_115 );
or g0960 ( new_n1132_, new_n1131_, new_n1104_ );
not g0961 ( new_n1133_, new_n1127_ );
and g0962 ( new_n1134_, new_n1132_, new_n1133_ );
or g0963 ( new_n1135_, new_n1134_, keyIn_0_120 );
and g0964 ( N421, new_n1129_, new_n1135_ );
not g0965 ( new_n1137_, keyIn_0_125 );
and g0966 ( new_n1138_, new_n1049_, new_n1045_ );
and g0967 ( new_n1139_, new_n1043_, keyIn_0_111 );
or g0968 ( new_n1140_, new_n1139_, new_n1138_ );
and g0969 ( new_n1141_, new_n1099_, keyIn_0_116 );
not g0970 ( new_n1142_, new_n1141_ );
or g0971 ( new_n1143_, new_n1099_, keyIn_0_116 );
and g0972 ( new_n1144_, new_n1142_, new_n1143_ );
or g0973 ( new_n1145_, new_n1144_, new_n1140_ );
not g0974 ( new_n1146_, new_n1145_ );
and g0975 ( new_n1147_, new_n1146_, keyIn_0_121 );
not g0976 ( new_n1148_, new_n1147_ );
not g0977 ( new_n1149_, keyIn_0_121 );
and g0978 ( new_n1150_, new_n1145_, new_n1149_ );
not g0979 ( new_n1151_, new_n1150_ );
and g0980 ( new_n1152_, new_n1052_, new_n1079_ );
and g0981 ( new_n1153_, new_n1151_, new_n1152_ );
and g0982 ( new_n1154_, new_n1153_, new_n1148_ );
not g0983 ( new_n1155_, new_n1154_ );
and g0984 ( new_n1156_, new_n1155_, new_n1137_ );
and g0985 ( new_n1157_, new_n1154_, keyIn_0_125 );
or g0986 ( N430, new_n1156_, new_n1157_ );
not g0987 ( new_n1159_, new_n965_ );
not g0988 ( new_n1160_, new_n967_ );
and g0989 ( new_n1161_, new_n1159_, new_n1160_ );
and g0990 ( new_n1162_, new_n1161_, keyIn_0_118 );
not g0991 ( new_n1163_, new_n1162_ );
not g0992 ( new_n1164_, keyIn_0_118 );
and g0993 ( new_n1165_, new_n968_, new_n1164_ );
not g0994 ( new_n1166_, new_n1165_ );
and g0995 ( new_n1167_, new_n1166_, new_n1101_ );
and g0996 ( new_n1168_, new_n1167_, new_n1163_ );
or g0997 ( new_n1169_, new_n1168_, keyIn_0_123 );
not g0998 ( new_n1170_, keyIn_0_123 );
not g0999 ( new_n1171_, new_n1101_ );
or g1000 ( new_n1172_, new_n1171_, new_n1165_ );
or g1001 ( new_n1173_, new_n1172_, new_n1162_ );
or g1002 ( new_n1174_, new_n1173_, new_n1170_ );
and g1003 ( new_n1175_, new_n1174_, new_n1169_ );
or g1004 ( new_n1176_, new_n1020_, new_n1023_ );
not g1005 ( new_n1177_, new_n1024_ );
and g1006 ( new_n1178_, new_n1177_, new_n1176_ );
or g1007 ( new_n1179_, new_n1178_, new_n1140_ );
not g1008 ( new_n1180_, keyIn_0_117 );
and g1009 ( new_n1181_, new_n944_, new_n940_ );
and g1010 ( new_n1182_, new_n938_, keyIn_0_113 );
or g1011 ( new_n1183_, new_n1182_, new_n1181_ );
or g1012 ( new_n1184_, new_n1183_, new_n1180_ );
or g1013 ( new_n1185_, new_n946_, keyIn_0_117 );
and g1014 ( new_n1186_, new_n1184_, new_n1185_ );
or g1015 ( new_n1187_, new_n1140_, new_n1099_ );
or g1016 ( new_n1188_, new_n1187_, new_n1078_ );
or g1017 ( new_n1189_, new_n1188_, new_n1186_ );
and g1018 ( new_n1190_, new_n1189_, keyIn_0_122 );
not g1019 ( new_n1191_, keyIn_0_122 );
and g1020 ( new_n1192_, new_n946_, keyIn_0_117 );
and g1021 ( new_n1193_, new_n1183_, new_n1180_ );
or g1022 ( new_n1194_, new_n1193_, new_n1192_ );
and g1023 ( new_n1195_, new_n1051_, new_n1100_ );
and g1024 ( new_n1196_, new_n1195_, new_n1079_ );
and g1025 ( new_n1197_, new_n1194_, new_n1196_ );
and g1026 ( new_n1198_, new_n1197_, new_n1191_ );
or g1027 ( new_n1199_, new_n1190_, new_n1198_ );
or g1028 ( new_n1200_, new_n1199_, new_n1179_ );
or g1029 ( new_n1201_, new_n1200_, new_n1175_ );
and g1030 ( new_n1202_, new_n1201_, keyIn_0_126 );
not g1031 ( new_n1203_, keyIn_0_126 );
and g1032 ( new_n1204_, new_n1173_, new_n1170_ );
and g1033 ( new_n1205_, new_n1168_, keyIn_0_123 );
or g1034 ( new_n1206_, new_n1204_, new_n1205_ );
or g1035 ( new_n1207_, new_n1197_, new_n1191_ );
or g1036 ( new_n1208_, new_n1189_, keyIn_0_122 );
and g1037 ( new_n1209_, new_n1208_, new_n1207_ );
and g1038 ( new_n1210_, new_n1209_, new_n1052_ );
and g1039 ( new_n1211_, new_n1210_, new_n1206_ );
and g1040 ( new_n1212_, new_n1211_, new_n1203_ );
or g1041 ( N431, new_n1202_, new_n1212_ );
not g1042 ( new_n1214_, keyIn_0_124 );
or g1043 ( new_n1215_, new_n988_, keyIn_0_119 );
and g1044 ( new_n1216_, new_n988_, keyIn_0_119 );
not g1045 ( new_n1217_, new_n1216_ );
and g1046 ( new_n1218_, new_n1217_, new_n1215_ );
or g1047 ( new_n1219_, new_n1161_, new_n1218_ );
or g1048 ( new_n1220_, new_n1219_, new_n1187_ );
or g1049 ( new_n1221_, new_n1220_, new_n1214_ );
not g1050 ( new_n1222_, new_n1215_ );
or g1051 ( new_n1223_, new_n1222_, new_n1216_ );
and g1052 ( new_n1224_, new_n1223_, new_n968_ );
and g1053 ( new_n1225_, new_n1224_, new_n1195_ );
or g1054 ( new_n1226_, new_n1225_, keyIn_0_124 );
and g1055 ( new_n1227_, new_n1221_, new_n1226_ );
or g1056 ( new_n1228_, new_n1150_, new_n1178_ );
or g1057 ( new_n1229_, new_n1228_, new_n1147_ );
or g1058 ( new_n1230_, new_n1227_, new_n1229_ );
or g1059 ( new_n1231_, new_n1230_, new_n1199_ );
and g1060 ( new_n1232_, new_n1231_, keyIn_0_127 );
not g1061 ( new_n1233_, keyIn_0_127 );
and g1062 ( new_n1234_, new_n1225_, keyIn_0_124 );
and g1063 ( new_n1235_, new_n1220_, new_n1214_ );
or g1064 ( new_n1236_, new_n1235_, new_n1234_ );
not g1065 ( new_n1237_, new_n1229_ );
and g1066 ( new_n1238_, new_n1236_, new_n1237_ );
and g1067 ( new_n1239_, new_n1238_, new_n1209_ );
and g1068 ( new_n1240_, new_n1239_, new_n1233_ );
or g1069 ( N432, new_n1232_, new_n1240_ );
endmodule