module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129, keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134, keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139, keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144, keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149, keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154, keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159, keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164, keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169, keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174, keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179, keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184, keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189, keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194, keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199, keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204, keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209, keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214, keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219, keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224, keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229, keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234, keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239, keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244, keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249, keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254, keyIn_0_255, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129, keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134, keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139, keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144, keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149, keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154, keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159, keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164, keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169, keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174, keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179, keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184, keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189, keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194, keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199, keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204, keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209, keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214, keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219, keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224, keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229, keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234, keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239, keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244, keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249, keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254, keyIn_0_255, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n976_, new_n1009_, new_n479_, new_n1105_, new_n955_, new_n608_, new_n888_, new_n847_, new_n1157_, new_n501_, new_n798_, new_n1180_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1048_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n390_, new_n743_, new_n779_, new_n1025_, new_n566_, new_n641_, new_n365_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n1176_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n1057_, new_n670_, new_n1024_, new_n456_, new_n691_, new_n1125_, new_n682_, new_n1075_, new_n812_, new_n911_, new_n679_, new_n937_, new_n667_, new_n821_, new_n542_, new_n548_, new_n669_, new_n1172_, new_n419_, new_n728_, new_n624_, new_n534_, new_n1071_, new_n1120_, new_n819_, new_n637_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n695_, new_n660_, new_n1060_, new_n413_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n552_, new_n678_, new_n649_, new_n706_, new_n1119_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n1045_, new_n500_, new_n898_, new_n1163_, new_n786_, new_n799_, new_n946_, new_n1188_, new_n721_, new_n504_, new_n1108_, new_n862_, new_n742_, new_n892_, new_n427_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n1167_, new_n626_, new_n959_, new_n990_, new_n774_, new_n716_, new_n701_, new_n792_, new_n1058_, new_n953_, new_n1162_, new_n481_, new_n1073_, new_n1110_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n1059_, new_n634_, new_n414_, new_n1101_, new_n635_, new_n685_, new_n1050_, new_n554_, new_n648_, new_n903_, new_n983_, new_n1151_, new_n844_, new_n430_, new_n822_, new_n482_, new_n1082_, new_n849_, new_n1018_, new_n855_, new_n606_, new_n1037_, new_n589_, new_n796_, new_n1083_, new_n655_, new_n759_, new_n1054_, new_n630_, new_n385_, new_n1049_, new_n988_, new_n478_, new_n694_, new_n461_, new_n710_, new_n971_, new_n565_, new_n764_, new_n906_, new_n683_, new_n511_, new_n463_, new_n510_, new_n966_, new_n351_, new_n1184_, new_n517_, new_n609_, new_n1031_, new_n961_, new_n890_, new_n530_, new_n1006_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n1005_, new_n999_, new_n715_, new_n811_, new_n443_, new_n1086_, new_n956_, new_n763_, new_n960_, new_n1138_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n970_, new_n995_, new_n1035_, new_n674_, new_n991_, new_n1044_, new_n497_, new_n1170_, new_n816_, new_n845_, new_n768_, new_n773_, new_n568_, new_n420_, new_n1051_, new_n876_, new_n899_, new_n1053_, new_n423_, new_n498_, new_n492_, new_n496_, new_n1046_, new_n1182_, new_n650_, new_n708_, new_n750_, new_n887_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n734_, new_n912_, new_n1062_, new_n925_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n452_, new_n920_, new_n656_, new_n1121_, new_n820_, new_n1127_, new_n771_, new_n388_, new_n979_, new_n1028_, new_n1168_, new_n508_, new_n714_, new_n483_, new_n1004_, new_n1152_, new_n394_, new_n1007_, new_n935_, new_n882_, new_n1145_, new_n657_, new_n1150_, new_n929_, new_n652_, new_n582_, new_n986_, new_n1159_, new_n1020_, new_n363_, new_n1113_, new_n441_, new_n785_, new_n477_, new_n664_, new_n600_, new_n1041_, new_n917_, new_n426_, new_n1036_, new_n1133_, new_n398_, new_n1177_, new_n646_, new_n1132_, new_n538_, new_n383_, new_n343_, new_n541_, new_n458_, new_n854_, new_n447_, new_n1026_, new_n1106_, new_n473_, new_n1147_, new_n790_, new_n1081_, new_n587_, new_n465_, new_n739_, new_n783_, new_n969_, new_n835_, new_n996_, new_n378_, new_n621_, new_n846_, new_n915_, new_n349_, new_n488_, new_n524_, new_n705_, new_n848_, new_n943_, new_n874_, new_n402_, new_n663_, new_n347_, new_n659_, new_n700_, new_n921_, new_n396_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n632_, new_n1039_, new_n671_, new_n965_, new_n528_, new_n952_, new_n1158_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n397_, new_n729_, new_n1111_, new_n975_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n1115_, new_n559_, new_n948_, new_n762_, new_n1055_, new_n838_, new_n923_, new_n1187_, new_n469_, new_n391_, new_n1154_, new_n437_, new_n1085_, new_n794_, new_n628_, new_n409_, new_n1090_, new_n745_, new_n457_, new_n553_, new_n1114_, new_n1084_, new_n1061_, new_n668_, new_n1128_, new_n1002_, new_n834_, new_n1169_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n1032_, new_n1171_, new_n688_, new_n384_, new_n900_, new_n1161_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n1034_, new_n661_, new_n1124_, new_n1000_, new_n633_, new_n797_, new_n784_, new_n724_, new_n1070_, new_n1109_, new_n860_, new_n494_, new_n672_, new_n616_, new_n529_, new_n884_, new_n914_, new_n938_, new_n1160_, new_n1166_, new_n809_, new_n1142_, new_n654_, new_n713_, new_n880_, new_n1102_, new_n604_, new_n1104_, new_n690_, new_n416_, new_n1043_, new_n744_, new_n571_, new_n400_, new_n758_, new_n460_, new_n1175_, new_n1136_, new_n693_, new_n505_, new_n619_, new_n471_, new_n967_, new_n577_, new_n374_, new_n1135_, new_n376_, new_n380_, new_n1079_, new_n747_, new_n749_, new_n861_, new_n1091_, new_n1095_, new_n998_, new_n352_, new_n1094_, new_n931_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n1064_, new_n1065_, new_n1118_, new_n493_, new_n547_, new_n907_, new_n665_, new_n800_, new_n897_, new_n1012_, new_n719_, new_n869_, new_n1178_, new_n586_, new_n570_, new_n598_, new_n893_, new_n993_, new_n1063_, new_n824_, new_n520_, new_n717_, new_n403_, new_n475_, new_n868_, new_n825_, new_n858_, new_n557_, new_n936_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1016_, new_n1074_, new_n748_, new_n1144_, new_n1137_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n1141_, new_n807_, new_n736_, new_n879_, new_n513_, new_n592_, new_n726_, new_n1123_, new_n558_, new_n382_, new_n583_, new_n617_, new_n1080_, new_n718_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n487_, new_n675_, new_n1126_, new_n1155_, new_n546_, new_n1186_, new_n612_, new_n919_, new_n1015_, new_n755_, new_n1040_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n450_, new_n345_, new_n1179_, new_n499_, new_n533_, new_n1088_, new_n1130_, new_n1148_, new_n795_, new_n1146_, new_n459_, new_n569_, new_n555_, new_n468_, new_n1122_, new_n977_, new_n1139_, new_n782_, new_n1185_, new_n444_, new_n392_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n1174_, new_n692_, new_n502_, new_n613_, new_n623_, new_n446_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n972_, new_n1067_, new_n891_, new_n631_, new_n453_, new_n516_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n1076_, new_n585_, new_n751_, new_n535_, new_n1038_, new_n372_, new_n725_, new_n814_, new_n503_, new_n527_, new_n772_, new_n852_, new_n1181_, new_n597_, new_n978_, new_n1093_, new_n1092_, new_n408_, new_n1143_, new_n470_, new_n1072_, new_n769_, new_n1190_, new_n1097_, new_n1069_, new_n651_, new_n433_, new_n1164_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n992_, new_n1098_, new_n732_, new_n687_, new_n370_, new_n1029_, new_n689_, new_n584_, new_n815_, new_n933_, new_n1052_, new_n638_, new_n523_, new_n909_, new_n857_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n512_, new_n788_, new_n841_, new_n989_, new_n1117_, new_n1112_, new_n711_, new_n1156_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n1116_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n1096_, new_n681_, new_n1087_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n1008_, new_n640_, new_n684_, new_n707_, new_n740_, new_n957_, new_n754_, new_n1047_, new_n787_, new_n653_, new_n1134_, new_n905_, new_n539_, new_n803_, new_n727_, new_n375_, new_n962_, new_n760_, new_n627_, new_n1173_, new_n704_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n1189_, new_n1153_, new_n357_, new_n780_, new_n984_, new_n1183_, new_n643_, new_n474_, new_n1129_, new_n467_, new_n1013_, new_n1077_, new_n490_, new_n560_, new_n1100_, new_n865_, new_n1027_, new_n358_, new_n877_, new_n610_, new_n843_, new_n545_, new_n611_, new_n703_, new_n698_, new_n1011_, new_n1165_, new_n425_, new_n896_, new_n802_, new_n697_, new_n1099_, new_n1023_, new_n951_, new_n709_, new_n866_, new_n540_, new_n1149_, new_n1066_, new_n434_, new_n947_, new_n994_, new_n982_, new_n422_, new_n964_, new_n1078_, new_n581_, new_n686_, new_n934_, new_n551_, new_n455_, new_n770_, new_n757_, new_n618_, new_n1140_, new_n521_, new_n1042_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n356_, new_n647_, new_n889_, new_n536_, new_n464_, new_n1089_, new_n573_, new_n765_, new_n405_, new_n1103_;

nand g000 ( new_n343_, N29, N42, N75 );
not g001 ( N388, new_n343_ );
nand g002 ( new_n345_, N29, N36, N80 );
not g003 ( N389, new_n345_ );
nand g004 ( new_n347_, N29, N36, N42 );
not g005 ( N390, new_n347_ );
nand g006 ( new_n349_, N85, N86 );
not g007 ( N391, new_n349_ );
nand g008 ( new_n351_, N1, N8 );
not g009 ( new_n352_, new_n351_ );
nand g010 ( new_n353_, new_n352_, N13, N17 );
not g011 ( N418, new_n353_ );
not g012 ( new_n355_, N13 );
not g013 ( new_n356_, N17 );
nand g014 ( new_n357_, N1, N26 );
nor g015 ( new_n358_, new_n357_, new_n355_, new_n356_ );
nand g016 ( N419, new_n358_, new_n347_ );
nand g017 ( N420, N59, N75, N80 );
nand g018 ( N421, N36, N59, N80 );
nand g019 ( N422, N36, N42, N59 );
not g020 ( new_n363_, N90 );
nor g021 ( new_n364_, N87, N88 );
nor g022 ( new_n365_, new_n364_, new_n363_ );
xnor g023 ( N423, new_n365_, keyIn_0_22 );
nand g024 ( N446, new_n358_, N390 );
nand g025 ( new_n368_, N1, N26, N51 );
nand g026 ( new_n369_, new_n368_, keyIn_0_0 );
not g027 ( new_n370_, keyIn_0_0 );
nand g028 ( new_n371_, new_n370_, N1, N26, N51 );
nand g029 ( new_n372_, new_n369_, new_n371_ );
xnor g030 ( N447, new_n372_, keyIn_0_26 );
nand g031 ( new_n374_, new_n352_, N13, N55 );
xor g032 ( new_n375_, new_n374_, keyIn_0_2 );
nand g033 ( new_n376_, N29, N68 );
nor g034 ( N448, new_n375_, new_n376_ );
nand g035 ( new_n378_, N59, N68, N74 );
nor g036 ( N449, new_n375_, new_n378_ );
not g037 ( new_n380_, N89 );
nor g038 ( N450, new_n364_, new_n380_ );
nand g039 ( new_n382_, N111, N116 );
nand g040 ( new_n383_, new_n382_, keyIn_0_6 );
nor g041 ( new_n384_, N111, N116 );
nor g042 ( new_n385_, new_n382_, keyIn_0_6 );
nor g043 ( new_n386_, new_n385_, new_n384_ );
nand g044 ( new_n387_, new_n386_, new_n383_ );
xor g045 ( new_n388_, N121, N126 );
xnor g046 ( new_n389_, new_n387_, new_n388_ );
xnor g047 ( new_n390_, new_n389_, N135 );
xnor g048 ( new_n391_, N91, N96 );
xnor g049 ( new_n392_, N101, N106 );
xnor g050 ( new_n393_, new_n391_, new_n392_ );
xnor g051 ( new_n394_, new_n393_, N130 );
xnor g052 ( N767, new_n390_, new_n394_ );
xor g053 ( new_n396_, N159, N165 );
xnor g054 ( new_n397_, N171, N177 );
xnor g055 ( new_n398_, new_n396_, new_n397_ );
xnor g056 ( new_n399_, new_n398_, N130 );
xnor g057 ( new_n400_, N183, N189 );
xnor g058 ( new_n401_, N195, N201 );
xnor g059 ( new_n402_, new_n400_, new_n401_ );
xnor g060 ( new_n403_, new_n402_, N207 );
xnor g061 ( N768, new_n399_, new_n403_ );
not g062 ( new_n405_, N261 );
not g063 ( new_n406_, keyIn_0_110 );
not g064 ( new_n407_, keyIn_0_65 );
not g065 ( new_n408_, keyIn_0_25 );
nand g066 ( new_n409_, new_n372_, keyIn_0_18 );
not g067 ( new_n410_, keyIn_0_18 );
nand g068 ( new_n411_, new_n369_, new_n410_, new_n371_ );
nand g069 ( new_n412_, new_n409_, new_n411_ );
nand g070 ( new_n413_, new_n412_, new_n408_ );
nand g071 ( new_n414_, new_n409_, keyIn_0_25, new_n411_ );
nand g072 ( new_n415_, new_n413_, new_n414_ );
nand g073 ( new_n416_, N59, N156 );
xor g074 ( new_n417_, new_n416_, keyIn_0_12 );
nand g075 ( new_n418_, new_n415_, keyIn_0_35, N17, new_n417_ );
not g076 ( new_n419_, keyIn_0_35 );
nand g077 ( new_n420_, new_n415_, N17, new_n417_ );
nand g078 ( new_n421_, new_n420_, new_n419_ );
nand g079 ( new_n422_, new_n421_, keyIn_0_46, N1, new_n418_ );
not g080 ( new_n423_, keyIn_0_46 );
nand g081 ( new_n424_, new_n421_, N1, new_n418_ );
nand g082 ( new_n425_, new_n424_, new_n423_ );
nand g083 ( new_n426_, new_n425_, N153, new_n422_ );
nand g084 ( new_n427_, new_n426_, new_n407_ );
nand g085 ( new_n428_, new_n425_, keyIn_0_65, N153, new_n422_ );
nand g086 ( new_n429_, new_n427_, new_n428_ );
not g087 ( new_n430_, keyIn_0_66 );
nor g088 ( new_n431_, N17, N42 );
nor g089 ( new_n432_, new_n431_, keyIn_0_13 );
not g090 ( new_n433_, keyIn_0_13 );
nor g091 ( new_n434_, new_n433_, N17, N42 );
nor g092 ( new_n435_, new_n432_, new_n434_ );
nand g093 ( new_n436_, N17, N42 );
xnor g094 ( new_n437_, new_n436_, keyIn_0_14 );
nor g095 ( new_n438_, new_n435_, new_n437_ );
nor g096 ( new_n439_, new_n438_, keyIn_0_24 );
not g097 ( new_n440_, new_n416_ );
not g098 ( new_n441_, N42 );
nand g099 ( new_n442_, new_n356_, new_n441_ );
nand g100 ( new_n443_, new_n442_, new_n433_ );
nand g101 ( new_n444_, new_n431_, keyIn_0_13 );
nand g102 ( new_n445_, new_n443_, new_n444_ );
nand g103 ( new_n446_, keyIn_0_14, N17, N42 );
not g104 ( new_n447_, keyIn_0_14 );
nand g105 ( new_n448_, new_n436_, new_n447_ );
nand g106 ( new_n449_, new_n448_, new_n446_ );
nand g107 ( new_n450_, new_n445_, keyIn_0_24, new_n449_ );
nand g108 ( new_n451_, new_n450_, new_n440_ );
nor g109 ( new_n452_, new_n439_, new_n451_ );
nand g110 ( new_n453_, new_n452_, new_n415_, keyIn_0_34 );
not g111 ( new_n454_, keyIn_0_34 );
nand g112 ( new_n455_, new_n452_, new_n415_ );
nand g113 ( new_n456_, new_n455_, new_n454_ );
not g114 ( new_n457_, keyIn_0_1 );
nand g115 ( new_n458_, N1, N8, N17, N51 );
nand g116 ( new_n459_, new_n458_, new_n457_ );
nand g117 ( new_n460_, new_n352_, keyIn_0_1, N17, N51 );
nand g118 ( new_n461_, new_n460_, new_n459_ );
nand g119 ( new_n462_, new_n461_, keyIn_0_19 );
not g120 ( new_n463_, keyIn_0_19 );
nand g121 ( new_n464_, new_n460_, new_n463_, new_n459_ );
nand g122 ( new_n465_, new_n462_, new_n464_ );
nand g123 ( new_n466_, N42, N59, N75 );
xnor g124 ( new_n467_, new_n466_, keyIn_0_5 );
nand g125 ( new_n468_, new_n467_, keyIn_0_21 );
not g126 ( new_n469_, keyIn_0_21 );
not g127 ( new_n470_, keyIn_0_5 );
xnor g128 ( new_n471_, new_n466_, new_n470_ );
nand g129 ( new_n472_, new_n471_, new_n469_ );
nand g130 ( new_n473_, new_n468_, new_n472_ );
nand g131 ( new_n474_, new_n465_, new_n473_ );
nand g132 ( new_n475_, new_n474_, keyIn_0_28 );
not g133 ( new_n476_, keyIn_0_28 );
nand g134 ( new_n477_, new_n465_, new_n473_, new_n476_ );
nand g135 ( new_n478_, new_n475_, new_n477_ );
nand g136 ( new_n479_, new_n456_, new_n453_, new_n478_ );
nand g137 ( new_n480_, new_n479_, keyIn_0_37 );
not g138 ( new_n481_, keyIn_0_37 );
nand g139 ( new_n482_, new_n456_, new_n478_, new_n481_, new_n453_ );
nand g140 ( new_n483_, new_n480_, new_n482_ );
nand g141 ( new_n484_, new_n483_, N126 );
nand g142 ( new_n485_, new_n484_, new_n430_ );
nand g143 ( new_n486_, new_n483_, keyIn_0_66, N126 );
nand g144 ( new_n487_, new_n485_, new_n486_ );
nand g145 ( new_n488_, new_n487_, new_n429_ );
nand g146 ( new_n489_, new_n488_, keyIn_0_80 );
nand g147 ( new_n490_, N29, N75, N80 );
xor g148 ( new_n491_, new_n490_, keyIn_0_4 );
nand g149 ( new_n492_, new_n415_, new_n491_ );
not g150 ( new_n493_, new_n492_ );
nand g151 ( new_n494_, new_n493_, N55 );
nand g152 ( new_n495_, new_n494_, keyIn_0_33 );
xnor g153 ( new_n496_, keyIn_0_8, N268 );
xnor g154 ( new_n497_, new_n496_, keyIn_0_23 );
not g155 ( new_n498_, new_n497_ );
not g156 ( new_n499_, keyIn_0_33 );
nand g157 ( new_n500_, new_n493_, new_n499_, N55 );
nand g158 ( new_n501_, new_n495_, new_n498_, new_n500_ );
xor g159 ( new_n502_, new_n501_, keyIn_0_50 );
not g160 ( new_n503_, keyIn_0_80 );
nand g161 ( new_n504_, new_n487_, new_n503_, new_n429_ );
nand g162 ( new_n505_, new_n489_, new_n502_, new_n504_ );
nand g163 ( new_n506_, new_n505_, keyIn_0_88 );
not g164 ( new_n507_, keyIn_0_88 );
nand g165 ( new_n508_, new_n489_, new_n507_, new_n502_, new_n504_ );
nand g166 ( new_n509_, new_n506_, new_n508_ );
nand g167 ( new_n510_, new_n509_, N201 );
nand g168 ( new_n511_, new_n510_, new_n406_ );
nand g169 ( new_n512_, new_n509_, keyIn_0_110, N201 );
not g170 ( new_n513_, N201 );
nand g171 ( new_n514_, new_n506_, new_n513_, new_n508_ );
xnor g172 ( new_n515_, new_n514_, keyIn_0_111 );
nand g173 ( new_n516_, new_n515_, new_n511_, new_n512_ );
xnor g174 ( new_n517_, new_n516_, keyIn_0_135 );
nand g175 ( new_n518_, new_n517_, keyIn_0_162, new_n405_ );
not g176 ( new_n519_, new_n517_ );
nand g177 ( new_n520_, new_n519_, keyIn_0_163, N261 );
not g178 ( new_n521_, keyIn_0_163 );
nand g179 ( new_n522_, new_n519_, N261 );
nand g180 ( new_n523_, new_n522_, new_n521_ );
not g181 ( new_n524_, keyIn_0_162 );
nand g182 ( new_n525_, new_n517_, new_n405_ );
nand g183 ( new_n526_, new_n525_, new_n524_ );
nand g184 ( new_n527_, new_n523_, new_n518_, new_n520_, new_n526_ );
nand g185 ( new_n528_, new_n527_, keyIn_0_182 );
not g186 ( new_n529_, keyIn_0_182 );
not g187 ( new_n530_, new_n527_ );
nand g188 ( new_n531_, new_n530_, new_n529_ );
nand g189 ( new_n532_, new_n531_, keyIn_0_190, N219, new_n528_ );
nand g190 ( new_n533_, N121, N210 );
xor g191 ( new_n534_, new_n533_, keyIn_0_17 );
not g192 ( new_n535_, keyIn_0_190 );
nand g193 ( new_n536_, new_n531_, N219, new_n528_ );
nand g194 ( new_n537_, new_n536_, new_n535_ );
nand g195 ( new_n538_, new_n537_, new_n532_, new_n534_ );
nand g196 ( new_n539_, new_n538_, keyIn_0_196 );
not g197 ( new_n540_, keyIn_0_196 );
nand g198 ( new_n541_, new_n537_, new_n540_, new_n532_, new_n534_ );
nand g199 ( new_n542_, new_n519_, keyIn_0_164, N228 );
not g200 ( new_n543_, keyIn_0_164 );
nand g201 ( new_n544_, new_n519_, N228 );
nand g202 ( new_n545_, new_n544_, new_n543_ );
nand g203 ( new_n546_, new_n511_, new_n512_ );
nand g204 ( new_n547_, new_n546_, keyIn_0_134 );
not g205 ( new_n548_, keyIn_0_134 );
nand g206 ( new_n549_, new_n511_, new_n548_, new_n512_ );
nand g207 ( new_n550_, new_n547_, new_n549_ );
nand g208 ( new_n551_, new_n550_, N237 );
xnor g209 ( new_n552_, new_n551_, keyIn_0_165 );
nand g210 ( new_n553_, new_n545_, new_n542_, new_n552_ );
nand g211 ( new_n554_, new_n553_, keyIn_0_183 );
nor g212 ( new_n555_, new_n553_, keyIn_0_183 );
nand g213 ( new_n556_, new_n509_, keyIn_0_112, N246 );
nand g214 ( new_n557_, N255, N267 );
not g215 ( new_n558_, keyIn_0_112 );
nand g216 ( new_n559_, new_n509_, N246 );
nand g217 ( new_n560_, new_n559_, new_n558_ );
nand g218 ( new_n561_, new_n560_, new_n556_, new_n557_ );
nand g219 ( new_n562_, new_n561_, keyIn_0_136 );
nand g220 ( new_n563_, N42, N59, N68, N72 );
xor g221 ( new_n564_, new_n563_, keyIn_0_3 );
nor g222 ( new_n565_, new_n375_, new_n564_ );
xor g223 ( new_n566_, new_n565_, keyIn_0_20 );
nand g224 ( new_n567_, new_n566_, N73 );
xnor g225 ( new_n568_, new_n567_, keyIn_0_27 );
xnor g226 ( new_n569_, new_n568_, keyIn_0_30 );
xor g227 ( new_n570_, new_n569_, keyIn_0_36 );
nand g228 ( new_n571_, new_n570_, N201 );
not g229 ( new_n572_, keyIn_0_136 );
nand g230 ( new_n573_, new_n560_, new_n572_, new_n556_, new_n557_ );
nand g231 ( new_n574_, new_n562_, new_n571_, new_n573_ );
nor g232 ( new_n575_, new_n555_, new_n574_ );
nand g233 ( new_n576_, new_n539_, new_n541_, new_n554_, new_n575_ );
xnor g234 ( new_n577_, new_n576_, keyIn_0_202 );
xor g235 ( new_n578_, new_n577_, keyIn_0_213 );
xnor g236 ( N850, new_n578_, keyIn_0_224 );
nand g237 ( new_n580_, new_n483_, N111 );
xnor g238 ( new_n581_, new_n580_, keyIn_0_60 );
xnor g239 ( new_n582_, new_n424_, keyIn_0_46 );
nand g240 ( new_n583_, new_n582_, N143 );
xor g241 ( new_n584_, new_n583_, keyIn_0_59 );
nand g242 ( new_n585_, new_n584_, new_n581_ );
nand g243 ( new_n586_, new_n585_, keyIn_0_77 );
xnor g244 ( new_n587_, new_n501_, keyIn_0_47 );
not g245 ( new_n588_, keyIn_0_77 );
nand g246 ( new_n589_, new_n584_, new_n588_, new_n581_ );
nand g247 ( new_n590_, new_n586_, new_n587_, new_n589_ );
xnor g248 ( new_n591_, new_n590_, keyIn_0_85 );
nand g249 ( new_n592_, new_n591_, N183 );
xnor g250 ( new_n593_, new_n592_, keyIn_0_101 );
not g251 ( new_n594_, N183 );
not g252 ( new_n595_, new_n591_ );
nand g253 ( new_n596_, new_n595_, new_n594_ );
xor g254 ( new_n597_, new_n596_, keyIn_0_102 );
nand g255 ( new_n598_, new_n597_, new_n593_ );
xnor g256 ( new_n599_, new_n598_, keyIn_0_126 );
not g257 ( new_n600_, keyIn_0_176 );
not g258 ( new_n601_, keyIn_0_155 );
not g259 ( new_n602_, keyIn_0_61 );
nand g260 ( new_n603_, new_n425_, N146, new_n422_ );
xnor g261 ( new_n604_, new_n603_, new_n602_ );
not g262 ( new_n605_, keyIn_0_62 );
nand g263 ( new_n606_, new_n483_, N116 );
nand g264 ( new_n607_, new_n606_, new_n605_ );
nand g265 ( new_n608_, new_n483_, keyIn_0_62, N116 );
nand g266 ( new_n609_, new_n604_, keyIn_0_78, new_n607_, new_n608_ );
xor g267 ( new_n610_, new_n501_, keyIn_0_48 );
not g268 ( new_n611_, keyIn_0_78 );
nand g269 ( new_n612_, new_n582_, new_n602_, N146 );
nand g270 ( new_n613_, new_n603_, keyIn_0_61 );
nand g271 ( new_n614_, new_n607_, new_n612_, new_n613_, new_n608_ );
nand g272 ( new_n615_, new_n614_, new_n611_ );
nand g273 ( new_n616_, new_n615_, new_n609_, keyIn_0_86, new_n610_ );
not g274 ( new_n617_, keyIn_0_86 );
nand g275 ( new_n618_, new_n615_, new_n609_, new_n610_ );
nand g276 ( new_n619_, new_n618_, new_n617_ );
nand g277 ( new_n620_, new_n619_, new_n616_ );
nand g278 ( new_n621_, new_n620_, keyIn_0_104, N189 );
not g279 ( new_n622_, keyIn_0_104 );
nand g280 ( new_n623_, new_n620_, N189 );
nand g281 ( new_n624_, new_n623_, new_n622_ );
nand g282 ( new_n625_, new_n624_, new_n621_ );
nand g283 ( new_n626_, new_n625_, keyIn_0_128 );
not g284 ( new_n627_, keyIn_0_128 );
nand g285 ( new_n628_, new_n624_, new_n627_, new_n621_ );
nand g286 ( new_n629_, new_n626_, new_n628_ );
nand g287 ( new_n630_, new_n629_, new_n601_ );
nand g288 ( new_n631_, new_n626_, keyIn_0_155, new_n628_ );
nand g289 ( new_n632_, new_n630_, new_n631_ );
not g290 ( new_n633_, N189 );
nand g291 ( new_n634_, new_n619_, new_n633_, new_n616_ );
xnor g292 ( new_n635_, new_n634_, keyIn_0_105 );
not g293 ( new_n636_, N195 );
not g294 ( new_n637_, keyIn_0_64 );
nand g295 ( new_n638_, new_n483_, new_n637_, N121 );
nand g296 ( new_n639_, new_n483_, N121 );
nand g297 ( new_n640_, new_n639_, keyIn_0_64 );
nand g298 ( new_n641_, new_n640_, new_n638_ );
nand g299 ( new_n642_, new_n425_, N149, new_n422_ );
xnor g300 ( new_n643_, new_n642_, keyIn_0_63 );
nand g301 ( new_n644_, new_n641_, new_n643_ );
nand g302 ( new_n645_, new_n644_, keyIn_0_79 );
xnor g303 ( new_n646_, new_n501_, keyIn_0_49 );
not g304 ( new_n647_, keyIn_0_79 );
nand g305 ( new_n648_, new_n641_, new_n643_, new_n647_ );
nand g306 ( new_n649_, new_n645_, keyIn_0_87, new_n646_, new_n648_ );
not g307 ( new_n650_, keyIn_0_87 );
nand g308 ( new_n651_, new_n645_, new_n646_, new_n648_ );
nand g309 ( new_n652_, new_n651_, new_n650_ );
nand g310 ( new_n653_, new_n652_, new_n649_ );
nand g311 ( new_n654_, new_n653_, new_n636_ );
nand g312 ( new_n655_, new_n654_, keyIn_0_108 );
not g313 ( new_n656_, keyIn_0_108 );
nand g314 ( new_n657_, new_n653_, new_n656_, new_n636_ );
nand g315 ( new_n658_, new_n655_, new_n657_ );
nand g316 ( new_n659_, new_n658_, new_n515_, N261, new_n635_ );
nand g317 ( new_n660_, new_n659_, keyIn_0_139 );
not g318 ( new_n661_, keyIn_0_139 );
nand g319 ( new_n662_, new_n515_, N261 );
not g320 ( new_n663_, new_n662_ );
nand g321 ( new_n664_, new_n663_, new_n661_, new_n635_, new_n658_ );
nand g322 ( new_n665_, new_n664_, new_n660_ );
nand g323 ( new_n666_, new_n665_, new_n632_ );
not g324 ( new_n667_, new_n666_ );
nand g325 ( new_n668_, new_n658_, new_n635_ );
not g326 ( new_n669_, new_n668_ );
nand g327 ( new_n670_, new_n550_, new_n669_ );
nand g328 ( new_n671_, new_n670_, keyIn_0_168 );
not g329 ( new_n672_, keyIn_0_168 );
nand g330 ( new_n673_, new_n550_, new_n669_, new_n672_ );
nand g331 ( new_n674_, new_n671_, new_n673_ );
not g332 ( new_n675_, keyIn_0_167 );
not g333 ( new_n676_, keyIn_0_131 );
nand g334 ( new_n677_, new_n652_, N195, new_n649_ );
nand g335 ( new_n678_, new_n677_, keyIn_0_107 );
not g336 ( new_n679_, keyIn_0_107 );
nand g337 ( new_n680_, new_n652_, new_n679_, N195, new_n649_ );
nand g338 ( new_n681_, new_n678_, new_n676_, new_n680_ );
nand g339 ( new_n682_, new_n678_, new_n680_ );
nand g340 ( new_n683_, new_n682_, keyIn_0_131 );
nand g341 ( new_n684_, new_n683_, new_n681_ );
nand g342 ( new_n685_, new_n684_, new_n635_ );
nand g343 ( new_n686_, new_n685_, new_n675_ );
nand g344 ( new_n687_, new_n684_, keyIn_0_167, new_n635_ );
nand g345 ( new_n688_, new_n686_, new_n687_ );
nand g346 ( new_n689_, new_n667_, new_n600_, new_n674_, new_n688_ );
nand g347 ( new_n690_, new_n674_, new_n632_, new_n665_, new_n688_ );
nand g348 ( new_n691_, new_n690_, keyIn_0_176 );
nand g349 ( new_n692_, new_n691_, new_n689_ );
nand g350 ( new_n693_, new_n692_, new_n599_ );
xnor g351 ( new_n694_, new_n693_, keyIn_0_185 );
not g352 ( new_n695_, new_n599_ );
nand g353 ( new_n696_, new_n695_, new_n689_, new_n691_ );
xor g354 ( new_n697_, new_n696_, keyIn_0_184 );
nand g355 ( new_n698_, new_n697_, new_n694_ );
xor g356 ( new_n699_, new_n698_, keyIn_0_193 );
nand g357 ( new_n700_, new_n699_, N219 );
nand g358 ( new_n701_, new_n700_, keyIn_0_199 );
nand g359 ( new_n702_, N106, N210 );
not g360 ( new_n703_, keyIn_0_199 );
nand g361 ( new_n704_, new_n699_, new_n703_, N219 );
nand g362 ( new_n705_, new_n701_, new_n702_, new_n704_ );
xnor g363 ( new_n706_, new_n705_, keyIn_0_210 );
not g364 ( new_n707_, keyIn_0_177 );
not g365 ( new_n708_, keyIn_0_153 );
nand g366 ( new_n709_, new_n599_, new_n708_, N228 );
nand g367 ( new_n710_, new_n599_, N228 );
nand g368 ( new_n711_, new_n710_, keyIn_0_153 );
xnor g369 ( new_n712_, new_n593_, keyIn_0_125 );
nand g370 ( new_n713_, new_n712_, N237 );
xnor g371 ( new_n714_, new_n713_, keyIn_0_154 );
nand g372 ( new_n715_, new_n711_, new_n709_, new_n714_ );
nand g373 ( new_n716_, new_n715_, new_n707_ );
not g374 ( new_n717_, keyIn_0_103 );
nand g375 ( new_n718_, new_n591_, new_n717_, N246 );
nand g376 ( new_n719_, new_n570_, N183 );
xor g377 ( new_n720_, new_n719_, keyIn_0_71 );
nand g378 ( new_n721_, new_n591_, N246 );
nand g379 ( new_n722_, new_n721_, keyIn_0_103 );
nand g380 ( new_n723_, new_n722_, new_n720_, new_n718_ );
xor g381 ( new_n724_, new_n723_, keyIn_0_127 );
nor g382 ( new_n725_, new_n715_, new_n707_ );
nor g383 ( new_n726_, new_n725_, new_n724_ );
nand g384 ( new_n727_, new_n706_, new_n716_, new_n726_ );
xnor g385 ( new_n728_, new_n727_, keyIn_0_221 );
xnor g386 ( new_n729_, new_n728_, keyIn_0_230 );
xnor g387 ( N863, new_n729_, keyIn_0_238 );
nand g388 ( new_n731_, new_n550_, new_n658_ );
xor g389 ( new_n732_, new_n731_, keyIn_0_166 );
nand g390 ( new_n733_, new_n663_, new_n658_ );
xnor g391 ( new_n734_, new_n733_, keyIn_0_138 );
xnor g392 ( new_n735_, new_n684_, keyIn_0_158 );
nand g393 ( new_n736_, new_n732_, new_n734_, new_n735_ );
xnor g394 ( new_n737_, new_n736_, keyIn_0_178 );
not g395 ( new_n738_, new_n737_ );
nand g396 ( new_n739_, new_n635_, new_n621_, new_n624_ );
xor g397 ( new_n740_, new_n739_, keyIn_0_129 );
not g398 ( new_n741_, new_n740_ );
nand g399 ( new_n742_, new_n738_, new_n741_ );
xor g400 ( new_n743_, new_n742_, keyIn_0_187 );
nand g401 ( new_n744_, new_n737_, new_n740_ );
xor g402 ( new_n745_, new_n744_, keyIn_0_186 );
nand g403 ( new_n746_, new_n743_, new_n745_ );
xor g404 ( new_n747_, new_n746_, keyIn_0_194 );
nand g405 ( new_n748_, new_n747_, keyIn_0_200, N219 );
not g406 ( new_n749_, keyIn_0_200 );
nand g407 ( new_n750_, new_n747_, N219 );
nand g408 ( new_n751_, new_n750_, new_n749_ );
nand g409 ( new_n752_, N111, N210 );
xnor g410 ( new_n753_, new_n752_, keyIn_0_16 );
nand g411 ( new_n754_, new_n751_, new_n748_, new_n753_ );
xnor g412 ( new_n755_, new_n754_, keyIn_0_211 );
nand g413 ( new_n756_, new_n741_, N228 );
xor g414 ( new_n757_, new_n756_, keyIn_0_156 );
nand g415 ( new_n758_, new_n626_, N237, new_n628_ );
xor g416 ( new_n759_, new_n758_, keyIn_0_157 );
nand g417 ( new_n760_, new_n757_, new_n759_ );
xor g418 ( new_n761_, new_n760_, keyIn_0_179 );
not g419 ( new_n762_, keyIn_0_130 );
nand g420 ( new_n763_, new_n620_, keyIn_0_106, N246 );
nand g421 ( new_n764_, N255, N259 );
not g422 ( new_n765_, keyIn_0_106 );
nand g423 ( new_n766_, new_n620_, N246 );
nand g424 ( new_n767_, new_n766_, new_n765_ );
nand g425 ( new_n768_, new_n767_, new_n762_, new_n763_, new_n764_ );
nand g426 ( new_n769_, new_n570_, N189 );
xor g427 ( new_n770_, new_n769_, keyIn_0_72 );
nand g428 ( new_n771_, new_n767_, new_n763_, new_n764_ );
nand g429 ( new_n772_, new_n771_, keyIn_0_130 );
nand g430 ( new_n773_, new_n772_, new_n768_, new_n770_ );
not g431 ( new_n774_, new_n773_ );
nand g432 ( new_n775_, new_n755_, new_n761_, new_n774_ );
xor g433 ( new_n776_, new_n775_, keyIn_0_222 );
xnor g434 ( new_n777_, new_n776_, keyIn_0_231 );
xnor g435 ( N864, new_n777_, keyIn_0_239 );
not g436 ( new_n779_, keyIn_0_212 );
not g437 ( new_n780_, keyIn_0_195 );
nand g438 ( new_n781_, new_n658_, new_n682_ );
xnor g439 ( new_n782_, new_n781_, keyIn_0_132 );
not g440 ( new_n783_, new_n782_ );
nand g441 ( new_n784_, new_n550_, keyIn_0_161 );
not g442 ( new_n785_, keyIn_0_161 );
nand g443 ( new_n786_, new_n547_, new_n785_, new_n549_ );
xor g444 ( new_n787_, new_n662_, keyIn_0_137 );
nand g445 ( new_n788_, new_n787_, new_n784_, new_n786_ );
xor g446 ( new_n789_, new_n788_, keyIn_0_180 );
nand g447 ( new_n790_, new_n789_, new_n783_ );
xor g448 ( new_n791_, new_n790_, keyIn_0_188 );
not g449 ( new_n792_, new_n789_ );
nand g450 ( new_n793_, new_n792_, new_n782_ );
xor g451 ( new_n794_, new_n793_, keyIn_0_189 );
nand g452 ( new_n795_, new_n794_, new_n780_, new_n791_ );
nand g453 ( new_n796_, new_n794_, new_n791_ );
nand g454 ( new_n797_, new_n796_, keyIn_0_195 );
nand g455 ( new_n798_, new_n797_, keyIn_0_201, N219, new_n795_ );
nand g456 ( new_n799_, N116, N210 );
not g457 ( new_n800_, keyIn_0_201 );
nand g458 ( new_n801_, new_n797_, N219, new_n795_ );
nand g459 ( new_n802_, new_n801_, new_n800_ );
nand g460 ( new_n803_, new_n802_, new_n798_, new_n799_ );
nand g461 ( new_n804_, new_n803_, new_n779_ );
nand g462 ( new_n805_, new_n802_, keyIn_0_212, new_n798_, new_n799_ );
nand g463 ( new_n806_, new_n782_, N228 );
nand g464 ( new_n807_, new_n806_, keyIn_0_159 );
not g465 ( new_n808_, keyIn_0_159 );
nand g466 ( new_n809_, new_n782_, new_n808_, N228 );
nand g467 ( new_n810_, new_n684_, N237 );
xnor g468 ( new_n811_, new_n810_, keyIn_0_160 );
nand g469 ( new_n812_, new_n807_, new_n809_, new_n811_ );
nand g470 ( new_n813_, new_n812_, keyIn_0_181 );
nor g471 ( new_n814_, new_n812_, keyIn_0_181 );
nand g472 ( new_n815_, new_n570_, N195 );
not g473 ( new_n816_, new_n815_ );
not g474 ( new_n817_, keyIn_0_109 );
not g475 ( new_n818_, new_n653_ );
nand g476 ( new_n819_, new_n818_, new_n817_, N246 );
nand g477 ( new_n820_, N255, N260 );
nand g478 ( new_n821_, new_n818_, N246 );
nand g479 ( new_n822_, new_n821_, keyIn_0_109 );
nand g480 ( new_n823_, new_n822_, new_n819_, new_n820_ );
xnor g481 ( new_n824_, new_n823_, keyIn_0_133 );
nor g482 ( new_n825_, new_n814_, new_n816_, new_n824_ );
nand g483 ( new_n826_, new_n804_, new_n805_, new_n813_, new_n825_ );
xor g484 ( new_n827_, new_n826_, keyIn_0_223 );
xnor g485 ( new_n828_, new_n827_, keyIn_0_232 );
xnor g486 ( N865, new_n828_, keyIn_0_240 );
not g487 ( new_n830_, keyIn_0_206 );
not g488 ( new_n831_, N165 );
nand g489 ( new_n832_, new_n483_, keyIn_0_53, N96 );
not g490 ( new_n833_, keyIn_0_53 );
nand g491 ( new_n834_, new_n483_, N96 );
nand g492 ( new_n835_, new_n834_, new_n833_ );
nand g493 ( new_n836_, N51, N138 );
xor g494 ( new_n837_, new_n836_, keyIn_0_9 );
nand g495 ( new_n838_, new_n835_, new_n832_, new_n837_ );
nand g496 ( new_n839_, new_n838_, keyIn_0_74 );
not g497 ( new_n840_, keyIn_0_74 );
nand g498 ( new_n841_, new_n835_, new_n840_, new_n832_, new_n837_ );
nand g499 ( new_n842_, new_n493_, N17 );
xor g500 ( new_n843_, new_n842_, keyIn_0_32 );
nand g501 ( new_n844_, new_n843_, new_n496_ );
xnor g502 ( new_n845_, new_n844_, keyIn_0_41 );
nand g503 ( new_n846_, new_n415_, N55, new_n417_ );
xor g504 ( new_n847_, new_n846_, keyIn_0_31 );
nand g505 ( new_n848_, new_n847_, N146 );
xor g506 ( new_n849_, new_n848_, keyIn_0_40 );
nand g507 ( new_n850_, new_n845_, new_n849_ );
xor g508 ( new_n851_, new_n850_, keyIn_0_54 );
nand g509 ( new_n852_, new_n851_, new_n839_, new_n841_ );
xnor g510 ( new_n853_, new_n852_, keyIn_0_82 );
not g511 ( new_n854_, new_n853_ );
nand g512 ( new_n855_, new_n854_, new_n831_ );
xor g513 ( new_n856_, new_n855_, keyIn_0_93 );
not g514 ( new_n857_, N171 );
nand g515 ( new_n858_, new_n483_, keyIn_0_55, N101 );
nand g516 ( new_n859_, N17, N138 );
xnor g517 ( new_n860_, new_n859_, keyIn_0_10 );
not g518 ( new_n861_, keyIn_0_55 );
nand g519 ( new_n862_, new_n483_, N101 );
nand g520 ( new_n863_, new_n862_, new_n861_ );
nand g521 ( new_n864_, new_n863_, new_n858_, new_n860_ );
xor g522 ( new_n865_, new_n864_, keyIn_0_75 );
nand g523 ( new_n866_, new_n843_, keyIn_0_43, new_n496_ );
not g524 ( new_n867_, keyIn_0_43 );
nand g525 ( new_n868_, new_n844_, new_n867_ );
nand g526 ( new_n869_, new_n847_, N149 );
xor g527 ( new_n870_, new_n869_, keyIn_0_42 );
nand g528 ( new_n871_, new_n870_, new_n866_, new_n868_ );
xnor g529 ( new_n872_, new_n871_, keyIn_0_56 );
nand g530 ( new_n873_, new_n872_, new_n865_ );
xor g531 ( new_n874_, new_n873_, keyIn_0_83 );
nand g532 ( new_n875_, new_n874_, new_n857_ );
xnor g533 ( new_n876_, new_n875_, keyIn_0_96 );
nand g534 ( new_n877_, new_n856_, new_n876_ );
not g535 ( new_n878_, new_n877_ );
not g536 ( new_n879_, keyIn_0_192 );
nand g537 ( new_n880_, new_n692_, new_n597_ );
nand g538 ( new_n881_, new_n880_, keyIn_0_191 );
not g539 ( new_n882_, keyIn_0_191 );
nand g540 ( new_n883_, new_n692_, new_n882_, new_n597_ );
nand g541 ( new_n884_, new_n881_, new_n883_ );
xnor g542 ( new_n885_, new_n712_, keyIn_0_152 );
nand g543 ( new_n886_, new_n884_, new_n885_ );
nand g544 ( new_n887_, new_n886_, new_n879_ );
nand g545 ( new_n888_, new_n884_, keyIn_0_192, new_n885_ );
nand g546 ( new_n889_, new_n887_, new_n888_ );
not g547 ( new_n890_, N177 );
nand g548 ( new_n891_, new_n847_, N153 );
xnor g549 ( new_n892_, new_n891_, keyIn_0_44 );
xor g550 ( new_n893_, new_n844_, keyIn_0_45 );
nand g551 ( new_n894_, new_n893_, new_n892_ );
xnor g552 ( new_n895_, new_n894_, keyIn_0_58 );
nand g553 ( new_n896_, new_n483_, N106 );
xor g554 ( new_n897_, new_n896_, keyIn_0_57 );
nand g555 ( new_n898_, N138, N152 );
xnor g556 ( new_n899_, new_n898_, keyIn_0_11 );
nand g557 ( new_n900_, new_n897_, new_n899_ );
xor g558 ( new_n901_, new_n900_, keyIn_0_76 );
nand g559 ( new_n902_, new_n901_, new_n895_ );
xnor g560 ( new_n903_, new_n902_, keyIn_0_84 );
not g561 ( new_n904_, new_n903_ );
nand g562 ( new_n905_, new_n904_, new_n890_ );
xor g563 ( new_n906_, new_n905_, keyIn_0_99 );
nand g564 ( new_n907_, new_n889_, new_n878_, new_n906_ );
nand g565 ( new_n908_, new_n907_, keyIn_0_205 );
not g566 ( new_n909_, keyIn_0_205 );
nand g567 ( new_n910_, new_n889_, new_n909_, new_n878_, new_n906_ );
nand g568 ( new_n911_, new_n908_, new_n910_ );
nand g569 ( new_n912_, new_n903_, N177 );
xnor g570 ( new_n913_, new_n912_, keyIn_0_98 );
xor g571 ( new_n914_, new_n913_, keyIn_0_122 );
nand g572 ( new_n915_, new_n878_, new_n914_ );
xor g573 ( new_n916_, new_n915_, keyIn_0_171 );
nand g574 ( new_n917_, new_n853_, N165 );
xor g575 ( new_n918_, new_n917_, keyIn_0_92 );
xnor g576 ( new_n919_, new_n918_, keyIn_0_116 );
xor g577 ( new_n920_, new_n919_, keyIn_0_143 );
not g578 ( new_n921_, new_n874_ );
nand g579 ( new_n922_, new_n921_, N171 );
xor g580 ( new_n923_, new_n922_, keyIn_0_95 );
xor g581 ( new_n924_, new_n923_, keyIn_0_119 );
nand g582 ( new_n925_, new_n924_, new_n856_ );
xor g583 ( new_n926_, new_n925_, keyIn_0_170 );
nor g584 ( new_n927_, new_n926_, new_n916_, new_n920_ );
nand g585 ( new_n928_, new_n911_, new_n927_ );
nand g586 ( new_n929_, new_n928_, new_n830_ );
nand g587 ( new_n930_, new_n911_, keyIn_0_206, new_n927_ );
nand g588 ( new_n931_, new_n929_, new_n930_ );
not g589 ( new_n932_, N159 );
not g590 ( new_n933_, keyIn_0_51 );
nand g591 ( new_n934_, new_n483_, new_n933_, N91 );
nand g592 ( new_n935_, new_n483_, N91 );
nand g593 ( new_n936_, new_n935_, keyIn_0_51 );
nand g594 ( new_n937_, N8, N138 );
xnor g595 ( new_n938_, new_n937_, keyIn_0_7 );
nand g596 ( new_n939_, new_n936_, new_n934_, new_n938_ );
nand g597 ( new_n940_, new_n939_, keyIn_0_73 );
not g598 ( new_n941_, keyIn_0_73 );
nand g599 ( new_n942_, new_n936_, new_n941_, new_n934_, new_n938_ );
nand g600 ( new_n943_, new_n847_, N143 );
xnor g601 ( new_n944_, new_n943_, keyIn_0_38 );
xor g602 ( new_n945_, new_n844_, keyIn_0_39 );
nand g603 ( new_n946_, new_n945_, new_n944_ );
xnor g604 ( new_n947_, new_n946_, keyIn_0_52 );
nand g605 ( new_n948_, new_n947_, new_n940_, new_n942_ );
xnor g606 ( new_n949_, new_n948_, keyIn_0_81 );
nand g607 ( new_n950_, new_n949_, new_n932_ );
xor g608 ( new_n951_, new_n950_, keyIn_0_90 );
nand g609 ( new_n952_, new_n931_, keyIn_0_225, new_n951_ );
not g610 ( new_n953_, new_n949_ );
nand g611 ( new_n954_, new_n953_, N159 );
xor g612 ( new_n955_, new_n954_, keyIn_0_89 );
xnor g613 ( new_n956_, new_n955_, keyIn_0_113 );
xor g614 ( new_n957_, new_n956_, keyIn_0_140 );
not g615 ( new_n958_, keyIn_0_225 );
nand g616 ( new_n959_, new_n931_, new_n951_ );
nand g617 ( new_n960_, new_n959_, new_n958_ );
nand g618 ( new_n961_, new_n960_, new_n952_, new_n957_ );
xor g619 ( new_n962_, new_n961_, keyIn_0_233 );
xnor g620 ( N866, new_n962_, keyIn_0_241 );
not g621 ( new_n964_, keyIn_0_220 );
not g622 ( new_n965_, keyIn_0_209 );
nand g623 ( new_n966_, new_n906_, new_n913_ );
xor g624 ( new_n967_, new_n966_, keyIn_0_123 );
nand g625 ( new_n968_, new_n887_, new_n888_, new_n967_ );
xor g626 ( new_n969_, new_n968_, keyIn_0_197 );
not g627 ( new_n970_, new_n967_ );
nand g628 ( new_n971_, new_n889_, new_n970_ );
xor g629 ( new_n972_, new_n971_, keyIn_0_198 );
nand g630 ( new_n973_, new_n972_, new_n969_ );
nand g631 ( new_n974_, new_n973_, new_n965_ );
nand g632 ( new_n975_, new_n972_, keyIn_0_209, new_n969_ );
nand g633 ( new_n976_, new_n974_, new_n964_, N219, new_n975_ );
nand g634 ( new_n977_, N101, N210 );
nand g635 ( new_n978_, new_n974_, N219, new_n975_ );
nand g636 ( new_n979_, new_n978_, keyIn_0_220 );
nand g637 ( new_n980_, new_n979_, new_n976_, new_n977_ );
nand g638 ( new_n981_, new_n980_, keyIn_0_229 );
not g639 ( new_n982_, keyIn_0_229 );
nand g640 ( new_n983_, new_n979_, new_n982_, new_n976_, new_n977_ );
not g641 ( new_n984_, keyIn_0_100 );
nand g642 ( new_n985_, new_n903_, new_n984_, N246 );
nand g643 ( new_n986_, new_n570_, N177 );
xor g644 ( new_n987_, new_n986_, keyIn_0_70 );
nand g645 ( new_n988_, new_n903_, N246 );
nand g646 ( new_n989_, new_n988_, keyIn_0_100 );
nand g647 ( new_n990_, new_n989_, new_n985_, new_n987_ );
xor g648 ( new_n991_, new_n990_, keyIn_0_124 );
nand g649 ( new_n992_, new_n970_, N228 );
xnor g650 ( new_n993_, new_n992_, keyIn_0_150 );
nand g651 ( new_n994_, new_n914_, N237 );
xor g652 ( new_n995_, new_n994_, keyIn_0_151 );
nand g653 ( new_n996_, new_n993_, new_n995_ );
xor g654 ( new_n997_, new_n996_, keyIn_0_175 );
nand g655 ( new_n998_, new_n981_, new_n983_, new_n991_, new_n997_ );
xor g656 ( new_n999_, new_n998_, keyIn_0_237 );
xnor g657 ( new_n1000_, new_n999_, keyIn_0_245 );
xnor g658 ( N874, new_n1000_, keyIn_0_249 );
not g659 ( new_n1002_, keyIn_0_246 );
not g660 ( new_n1003_, keyIn_0_234 );
not g661 ( new_n1004_, keyIn_0_226 );
not g662 ( new_n1005_, keyIn_0_215 );
nand g663 ( new_n1006_, new_n955_, new_n951_ );
xor g664 ( new_n1007_, new_n1006_, keyIn_0_114 );
nand g665 ( new_n1008_, new_n931_, new_n1007_ );
nand g666 ( new_n1009_, new_n1008_, new_n1005_ );
nand g667 ( new_n1010_, new_n931_, keyIn_0_215, new_n1007_ );
nand g668 ( new_n1011_, new_n1009_, new_n1010_ );
not g669 ( new_n1012_, keyIn_0_214 );
not g670 ( new_n1013_, new_n1007_ );
nand g671 ( new_n1014_, new_n929_, new_n930_, new_n1013_ );
xnor g672 ( new_n1015_, new_n1014_, new_n1012_ );
nand g673 ( new_n1016_, new_n1011_, new_n1015_, new_n1004_ );
nand g674 ( new_n1017_, new_n1011_, new_n1015_ );
nand g675 ( new_n1018_, new_n1017_, keyIn_0_226 );
nand g676 ( new_n1019_, new_n1018_, new_n1003_, N219, new_n1016_ );
nand g677 ( new_n1020_, new_n497_, N210 );
xor g678 ( new_n1021_, new_n1020_, keyIn_0_29 );
nand g679 ( new_n1022_, new_n1018_, N219, new_n1016_ );
nand g680 ( new_n1023_, new_n1022_, keyIn_0_234 );
nand g681 ( new_n1024_, new_n1023_, new_n1019_, new_n1021_ );
nand g682 ( new_n1025_, new_n1024_, keyIn_0_242 );
not g683 ( new_n1026_, keyIn_0_242 );
nand g684 ( new_n1027_, new_n1023_, new_n1026_, new_n1019_, new_n1021_ );
nand g685 ( new_n1028_, new_n1025_, new_n1027_ );
nand g686 ( new_n1029_, new_n1007_, N228 );
xor g687 ( new_n1030_, new_n1029_, keyIn_0_141 );
nand g688 ( new_n1031_, new_n956_, N237 );
xor g689 ( new_n1032_, new_n1031_, keyIn_0_142 );
nand g690 ( new_n1033_, new_n1030_, new_n1032_ );
xor g691 ( new_n1034_, new_n1033_, keyIn_0_172 );
not g692 ( new_n1035_, keyIn_0_91 );
nand g693 ( new_n1036_, new_n953_, new_n1035_, N246 );
nand g694 ( new_n1037_, new_n570_, N159 );
xnor g695 ( new_n1038_, new_n1037_, keyIn_0_67 );
nand g696 ( new_n1039_, new_n953_, N246 );
nand g697 ( new_n1040_, new_n1039_, keyIn_0_91 );
nand g698 ( new_n1041_, new_n1040_, new_n1036_, new_n1038_ );
xnor g699 ( new_n1042_, new_n1041_, keyIn_0_115 );
nand g700 ( new_n1043_, new_n1034_, new_n1042_ );
not g701 ( new_n1044_, new_n1043_ );
nand g702 ( new_n1045_, new_n1028_, new_n1044_ );
nand g703 ( new_n1046_, new_n1045_, new_n1002_ );
nand g704 ( new_n1047_, new_n1028_, keyIn_0_246, new_n1044_ );
nand g705 ( new_n1048_, new_n1046_, new_n1047_ );
nand g706 ( new_n1049_, new_n1048_, keyIn_0_250 );
not g707 ( new_n1050_, keyIn_0_250 );
nand g708 ( new_n1051_, new_n1046_, new_n1050_, new_n1047_ );
nand g709 ( new_n1052_, new_n1049_, new_n1051_ );
nand g710 ( new_n1053_, new_n1052_, keyIn_0_253 );
not g711 ( new_n1054_, keyIn_0_253 );
nand g712 ( new_n1055_, new_n1049_, new_n1054_, new_n1051_ );
nand g713 ( N878, new_n1053_, new_n1055_ );
not g714 ( new_n1057_, keyIn_0_251 );
not g715 ( new_n1058_, keyIn_0_227 );
nand g716 ( new_n1059_, new_n856_, new_n918_ );
xor g717 ( new_n1060_, new_n1059_, keyIn_0_117 );
not g718 ( new_n1061_, new_n1060_ );
not g719 ( new_n1062_, keyIn_0_204 );
nand g720 ( new_n1063_, new_n889_, new_n1062_, new_n876_, new_n906_ );
nand g721 ( new_n1064_, new_n889_, new_n876_, new_n906_ );
nand g722 ( new_n1065_, new_n1064_, keyIn_0_204 );
not g723 ( new_n1066_, keyIn_0_169 );
nand g724 ( new_n1067_, new_n914_, new_n876_ );
nand g725 ( new_n1068_, new_n1067_, new_n1066_ );
nand g726 ( new_n1069_, new_n914_, keyIn_0_169, new_n876_ );
xor g727 ( new_n1070_, new_n924_, keyIn_0_146 );
nand g728 ( new_n1071_, new_n1070_, new_n1068_, new_n1069_ );
not g729 ( new_n1072_, new_n1071_ );
nand g730 ( new_n1073_, new_n1065_, new_n1063_, new_n1072_ );
xnor g731 ( new_n1074_, new_n1073_, keyIn_0_207 );
nand g732 ( new_n1075_, new_n1074_, new_n1061_ );
nand g733 ( new_n1076_, new_n1075_, keyIn_0_217 );
not g734 ( new_n1077_, keyIn_0_217 );
nand g735 ( new_n1078_, new_n1074_, new_n1077_, new_n1061_ );
nand g736 ( new_n1079_, new_n1076_, new_n1078_ );
not g737 ( new_n1080_, keyIn_0_216 );
not g738 ( new_n1081_, keyIn_0_207 );
xnor g739 ( new_n1082_, new_n1073_, new_n1081_ );
nand g740 ( new_n1083_, new_n1082_, new_n1080_, new_n1060_ );
nand g741 ( new_n1084_, new_n1082_, new_n1060_ );
nand g742 ( new_n1085_, new_n1084_, keyIn_0_216 );
nand g743 ( new_n1086_, new_n1085_, new_n1083_ );
nand g744 ( new_n1087_, new_n1079_, new_n1086_, new_n1058_ );
nand g745 ( new_n1088_, new_n1079_, new_n1086_ );
nand g746 ( new_n1089_, new_n1088_, keyIn_0_227 );
nand g747 ( new_n1090_, new_n1089_, new_n1087_ );
nand g748 ( new_n1091_, new_n1090_, keyIn_0_235, N219 );
not g749 ( new_n1092_, keyIn_0_235 );
nand g750 ( new_n1093_, new_n1090_, N219 );
nand g751 ( new_n1094_, new_n1093_, new_n1092_ );
nand g752 ( new_n1095_, N91, N210 );
xor g753 ( new_n1096_, new_n1095_, keyIn_0_15 );
nand g754 ( new_n1097_, new_n1094_, keyIn_0_243, new_n1091_, new_n1096_ );
not g755 ( new_n1098_, keyIn_0_243 );
nand g756 ( new_n1099_, new_n1094_, new_n1091_, new_n1096_ );
nand g757 ( new_n1100_, new_n1099_, new_n1098_ );
nand g758 ( new_n1101_, new_n919_, N237 );
xor g759 ( new_n1102_, new_n1101_, keyIn_0_145 );
not g760 ( new_n1103_, keyIn_0_144 );
nand g761 ( new_n1104_, new_n1061_, new_n1103_, N228 );
nand g762 ( new_n1105_, new_n1061_, N228 );
nand g763 ( new_n1106_, new_n1105_, keyIn_0_144 );
nand g764 ( new_n1107_, new_n1106_, new_n1102_, new_n1104_ );
nand g765 ( new_n1108_, new_n1107_, keyIn_0_173 );
not g766 ( new_n1109_, new_n1108_ );
nand g767 ( new_n1110_, new_n853_, N246 );
xnor g768 ( new_n1111_, new_n1110_, keyIn_0_94 );
nand g769 ( new_n1112_, new_n570_, N165 );
xnor g770 ( new_n1113_, new_n1112_, keyIn_0_68 );
nand g771 ( new_n1114_, new_n1111_, new_n1113_ );
xnor g772 ( new_n1115_, new_n1114_, keyIn_0_118 );
not g773 ( new_n1116_, keyIn_0_173 );
nand g774 ( new_n1117_, new_n1106_, new_n1116_, new_n1102_, new_n1104_ );
not g775 ( new_n1118_, new_n1117_ );
nor g776 ( new_n1119_, new_n1109_, new_n1115_, new_n1118_ );
nand g777 ( new_n1120_, new_n1100_, keyIn_0_247, new_n1097_, new_n1119_ );
not g778 ( new_n1121_, keyIn_0_247 );
nand g779 ( new_n1122_, new_n1100_, new_n1097_, new_n1119_ );
nand g780 ( new_n1123_, new_n1122_, new_n1121_ );
nand g781 ( new_n1124_, new_n1123_, new_n1120_ );
nand g782 ( new_n1125_, new_n1124_, new_n1057_ );
nand g783 ( new_n1126_, new_n1123_, keyIn_0_251, new_n1120_ );
nand g784 ( new_n1127_, new_n1125_, new_n1126_ );
nand g785 ( new_n1128_, new_n1127_, keyIn_0_254 );
not g786 ( new_n1129_, keyIn_0_254 );
nand g787 ( new_n1130_, new_n1125_, new_n1129_, new_n1126_ );
nand g788 ( N879, new_n1128_, new_n1130_ );
not g789 ( new_n1132_, keyIn_0_244 );
nand g790 ( new_n1133_, new_n923_, new_n876_ );
xor g791 ( new_n1134_, new_n1133_, keyIn_0_120 );
not g792 ( new_n1135_, keyIn_0_203 );
nand g793 ( new_n1136_, new_n889_, new_n1135_, new_n906_ );
xnor g794 ( new_n1137_, new_n914_, keyIn_0_149 );
nand g795 ( new_n1138_, new_n889_, new_n906_ );
nand g796 ( new_n1139_, new_n1138_, keyIn_0_203 );
nand g797 ( new_n1140_, new_n1139_, new_n1136_, new_n1137_ );
xnor g798 ( new_n1141_, new_n1140_, keyIn_0_208 );
nand g799 ( new_n1142_, new_n1141_, new_n1134_ );
nand g800 ( new_n1143_, new_n1142_, keyIn_0_218 );
not g801 ( new_n1144_, keyIn_0_219 );
not g802 ( new_n1145_, new_n1134_ );
not g803 ( new_n1146_, new_n1141_ );
nand g804 ( new_n1147_, new_n1146_, new_n1145_ );
nand g805 ( new_n1148_, new_n1147_, new_n1144_ );
not g806 ( new_n1149_, keyIn_0_218 );
nand g807 ( new_n1150_, new_n1141_, new_n1149_, new_n1134_ );
nand g808 ( new_n1151_, new_n1146_, keyIn_0_219, new_n1145_ );
nand g809 ( new_n1152_, new_n1151_, new_n1150_ );
not g810 ( new_n1153_, new_n1152_ );
nand g811 ( new_n1154_, new_n1153_, keyIn_0_228, new_n1143_, new_n1148_ );
not g812 ( new_n1155_, keyIn_0_228 );
nand g813 ( new_n1156_, new_n1148_, new_n1143_, new_n1150_, new_n1151_ );
nand g814 ( new_n1157_, new_n1156_, new_n1155_ );
nand g815 ( new_n1158_, new_n1154_, new_n1157_, N219 );
nand g816 ( new_n1159_, new_n1158_, keyIn_0_236 );
nand g817 ( new_n1160_, N96, N210 );
not g818 ( new_n1161_, keyIn_0_236 );
nand g819 ( new_n1162_, new_n1154_, new_n1157_, new_n1161_, N219 );
nand g820 ( new_n1163_, new_n1159_, new_n1132_, new_n1160_, new_n1162_ );
nand g821 ( new_n1164_, new_n1159_, new_n1160_, new_n1162_ );
nand g822 ( new_n1165_, new_n1164_, keyIn_0_244 );
nand g823 ( new_n1166_, new_n1145_, N228 );
xor g824 ( new_n1167_, new_n1166_, keyIn_0_147 );
nand g825 ( new_n1168_, new_n924_, N237 );
xor g826 ( new_n1169_, new_n1168_, keyIn_0_148 );
nand g827 ( new_n1170_, new_n1167_, new_n1169_ );
xor g828 ( new_n1171_, new_n1170_, keyIn_0_174 );
not g829 ( new_n1172_, keyIn_0_97 );
nand g830 ( new_n1173_, new_n921_, new_n1172_, N246 );
nand g831 ( new_n1174_, new_n570_, N171 );
xnor g832 ( new_n1175_, new_n1174_, keyIn_0_69 );
nand g833 ( new_n1176_, new_n921_, N246 );
nand g834 ( new_n1177_, new_n1176_, keyIn_0_97 );
nand g835 ( new_n1178_, new_n1177_, new_n1173_, new_n1175_ );
xnor g836 ( new_n1179_, new_n1178_, keyIn_0_121 );
nand g837 ( new_n1180_, new_n1171_, new_n1179_ );
not g838 ( new_n1181_, new_n1180_ );
nand g839 ( new_n1182_, new_n1165_, keyIn_0_248, new_n1163_, new_n1181_ );
not g840 ( new_n1183_, keyIn_0_248 );
nand g841 ( new_n1184_, new_n1165_, new_n1163_, new_n1181_ );
nand g842 ( new_n1185_, new_n1184_, new_n1183_ );
nand g843 ( new_n1186_, new_n1185_, new_n1182_ );
nand g844 ( new_n1187_, new_n1186_, keyIn_0_252 );
not g845 ( new_n1188_, keyIn_0_252 );
nand g846 ( new_n1189_, new_n1185_, new_n1188_, new_n1182_ );
nand g847 ( new_n1190_, new_n1187_, new_n1189_ );
xnor g848 ( N880, new_n1190_, keyIn_0_255 );
endmodule