module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n595_, new_n445_, new_n1009_, new_n238_, new_n479_, new_n1105_, new_n608_, new_n501_, new_n1157_, new_n421_, new_n777_, new_n1048_, new_n885_, new_n439_, new_n283_, new_n223_, new_n390_, new_n743_, new_n241_, new_n566_, new_n186_, new_n339_, new_n641_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n1024_, new_n1125_, new_n246_, new_n911_, new_n679_, new_n937_, new_n667_, new_n367_, new_n173_, new_n728_, new_n1071_, new_n214_, new_n894_, new_n853_, new_n695_, new_n660_, new_n526_, new_n908_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n752_, new_n1045_, new_n500_, new_n1163_, new_n786_, new_n317_, new_n1188_, new_n721_, new_n504_, new_n742_, new_n892_, new_n234_, new_n472_, new_n873_, new_n1167_, new_n774_, new_n792_, new_n953_, new_n257_, new_n481_, new_n1073_, new_n1110_, new_n449_, new_n580_, new_n639_, new_n484_, new_n766_, new_n272_, new_n282_, new_n1059_, new_n634_, new_n192_, new_n635_, new_n685_, new_n326_, new_n648_, new_n903_, new_n983_, new_n822_, new_n1082_, new_n1018_, new_n606_, new_n796_, new_n655_, new_n1054_, new_n630_, new_n385_, new_n1049_, new_n694_, new_n461_, new_n297_, new_n565_, new_n1196_, new_n183_, new_n511_, new_n303_, new_n325_, new_n1031_, new_n629_, new_n883_, new_n1005_, new_n999_, new_n324_, new_n960_, new_n491_, new_n549_, new_n676_, new_n995_, new_n1035_, new_n271_, new_n674_, new_n274_, new_n991_, new_n1044_, new_n497_, new_n816_, new_n568_, new_n420_, new_n876_, new_n423_, new_n498_, new_n496_, new_n1046_, new_n1182_, new_n708_, new_n206_, new_n429_, new_n353_, new_n734_, new_n912_, new_n1062_, new_n506_, new_n680_, new_n872_, new_n981_, new_n1198_, new_n656_, new_n1127_, new_n388_, new_n1028_, new_n1168_, new_n194_, new_n483_, new_n1004_, new_n1152_, new_n394_, new_n299_, new_n935_, new_n657_, new_n1150_, new_n652_, new_n582_, new_n1020_, new_n363_, new_n1113_, new_n441_, new_n785_, new_n477_, new_n664_, new_n600_, new_n280_, new_n1041_, new_n426_, new_n1036_, new_n235_, new_n398_, new_n301_, new_n1132_, new_n395_, new_n383_, new_n343_, new_n854_, new_n458_, new_n1106_, new_n207_, new_n267_, new_n473_, new_n1147_, new_n187_, new_n969_, new_n334_, new_n331_, new_n835_, new_n378_, new_n621_, new_n244_, new_n172_, new_n705_, new_n943_, new_n874_, new_n402_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n1003_, new_n696_, new_n208_, new_n1039_, new_n528_, new_n952_, new_n179_, new_n1158_, new_n729_, new_n1111_, new_n559_, new_n1201_, new_n762_, new_n1193_, new_n1187_, new_n1205_, new_n1154_, new_n295_, new_n628_, new_n409_, new_n1090_, new_n745_, new_n553_, new_n1114_, new_n1084_, new_n1061_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n1032_, new_n867_, new_n954_, new_n901_, new_n1171_, new_n276_, new_n688_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n886_, new_n371_, new_n509_, new_n202_, new_n296_, new_n661_, new_n797_, new_n232_, new_n724_, new_n1070_, new_n1109_, new_n261_, new_n672_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n938_, new_n362_, new_n809_, new_n1142_, new_n604_, new_n1104_, new_n571_, new_n758_, new_n328_, new_n460_, new_n268_, new_n380_, new_n1079_, new_n861_, new_n352_, new_n931_, new_n575_, new_n562_, new_n944_, new_n1064_, new_n1065_, new_n177_, new_n1118_, new_n493_, new_n547_, new_n264_, new_n379_, new_n273_, new_n224_, new_n586_, new_n963_, new_n993_, new_n1191_, new_n824_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n858_, new_n936_, new_n189_, new_n411_, new_n1016_, new_n673_, new_n1144_, new_n182_, new_n407_, new_n666_, new_n736_, new_n879_, new_n513_, new_n558_, new_n219_, new_n313_, new_n382_, new_n239_, new_n718_, new_n1126_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n302_, new_n755_, new_n1040_, new_n544_, new_n615_, new_n722_, new_n856_, new_n415_, new_n537_, new_n345_, new_n499_, new_n255_, new_n533_, new_n1130_, new_n795_, new_n459_, new_n1122_, new_n1185_, new_n354_, new_n1174_, new_n968_, new_n613_, new_n337_, new_n1195_, new_n417_, new_n658_, new_n591_, new_n837_, new_n801_, new_n631_, new_n453_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n531_, new_n593_, new_n974_, new_n252_, new_n751_, new_n1038_, new_n372_, new_n852_, new_n978_, new_n408_, new_n470_, new_n213_, new_n769_, new_n433_, new_n871_, new_n992_, new_n1098_, new_n265_, new_n732_, new_n689_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n1052_, new_n857_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n269_, new_n512_, new_n989_, new_n1117_, new_n644_, new_n836_, new_n1116_, new_n904_, new_n913_, new_n327_, new_n681_, new_n594_, new_n561_, new_n495_, new_n927_, new_n431_, new_n1206_, new_n196_, new_n818_, new_n881_, new_n640_, new_n684_, new_n754_, new_n653_, new_n377_, new_n905_, new_n375_, new_n962_, new_n760_, new_n627_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n1153_, new_n357_, new_n320_, new_n780_, new_n984_, new_n1183_, new_n245_, new_n643_, new_n1194_, new_n1027_, new_n348_, new_n610_, new_n843_, new_n322_, new_n703_, new_n698_, new_n1165_, new_n175_, new_n226_, new_n1208_, new_n697_, new_n1099_, new_n185_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n540_, new_n1149_, new_n1066_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n770_, new_n757_, new_n521_, new_n793_, new_n406_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n1089_, new_n1192_, new_n405_, new_n942_, new_n614_, new_n895_, new_n958_, new_n976_, new_n699_, new_n236_, new_n955_, new_n847_, new_n250_, new_n888_, new_n288_, new_n798_, new_n1180_, new_n817_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n941_, new_n827_, new_n366_, new_n779_, new_n1025_, new_n365_, new_n859_, new_n197_, new_n1207_, new_n1176_, new_n601_, new_n842_, new_n1057_, new_n682_, new_n1075_, new_n812_, new_n266_, new_n821_, new_n542_, new_n548_, new_n669_, new_n220_, new_n419_, new_n624_, new_n534_, new_n1131_, new_n1120_, new_n819_, new_n637_, new_n451_, new_n489_, new_n424_, new_n804_, new_n602_, new_n188_, new_n1060_, new_n240_, new_n413_, new_n442_, new_n677_, new_n642_, new_n211_, new_n462_, new_n603_, new_n564_, new_n761_, new_n840_, new_n735_, new_n898_, new_n799_, new_n946_, new_n344_, new_n287_, new_n1108_, new_n862_, new_n427_, new_n532_, new_n393_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n959_, new_n990_, new_n716_, new_n701_, new_n1058_, new_n1162_, new_n212_, new_n902_, new_n364_, new_n832_, new_n201_, new_n414_, new_n1101_, new_n315_, new_n1050_, new_n554_, new_n230_, new_n1151_, new_n281_, new_n430_, new_n844_, new_n482_, new_n849_, new_n1203_, new_n855_, new_n1037_, new_n589_, new_n248_, new_n350_, new_n759_, new_n1083_, new_n829_, new_n988_, new_n478_, new_n710_, new_n971_, new_n906_, new_n361_, new_n764_, new_n683_, new_n463_, new_n510_, new_n966_, new_n351_, new_n1184_, new_n517_, new_n609_, new_n180_, new_n961_, new_n530_, new_n890_, new_n318_, new_n1006_, new_n622_, new_n702_, new_n833_, new_n715_, new_n811_, new_n443_, new_n1086_, new_n956_, new_n763_, new_n1138_, new_n486_, new_n970_, new_n466_, new_n262_, new_n218_, new_n1170_, new_n845_, new_n768_, new_n773_, new_n305_, new_n1051_, new_n899_, new_n1053_, new_n205_, new_n492_, new_n1200_, new_n650_, new_n750_, new_n887_, new_n254_, new_n355_, new_n926_, new_n432_, new_n925_, new_n875_, new_n256_, new_n778_, new_n452_, new_n381_, new_n920_, new_n1121_, new_n820_, new_n771_, new_n979_, new_n508_, new_n714_, new_n1007_, new_n882_, new_n1145_, new_n929_, new_n986_, new_n314_, new_n1159_, new_n216_, new_n917_, new_n1133_, new_n1177_, new_n646_, new_n538_, new_n1026_, new_n210_, new_n541_, new_n447_, new_n790_, new_n1081_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n263_, new_n341_, new_n996_, new_n846_, new_n915_, new_n349_, new_n488_, new_n524_, new_n848_, new_n277_, new_n663_, new_n579_, new_n286_, new_n198_, new_n438_, new_n939_, new_n632_, new_n671_, new_n965_, new_n572_, new_n1019_, new_n1202_, new_n436_, new_n397_, new_n975_, new_n1199_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n1115_, new_n948_, new_n1055_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n1085_, new_n359_, new_n794_, new_n457_, new_n1128_, new_n1002_, new_n1169_, new_n448_, new_n384_, new_n900_, new_n1161_, new_n924_, new_n775_, new_n454_, new_n1034_, new_n1124_, new_n308_, new_n1000_, new_n633_, new_n784_, new_n258_, new_n176_, new_n860_, new_n306_, new_n494_, new_n291_, new_n309_, new_n1160_, new_n1166_, new_n259_, new_n654_, new_n713_, new_n880_, new_n1102_, new_n227_, new_n690_, new_n416_, new_n222_, new_n1043_, new_n744_, new_n400_, new_n1175_, new_n1136_, new_n693_, new_n505_, new_n619_, new_n471_, new_n967_, new_n577_, new_n374_, new_n1135_, new_n376_, new_n747_, new_n749_, new_n1091_, new_n310_, new_n1095_, new_n275_, new_n998_, new_n1056_, new_n1094_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n578_, new_n918_, new_n940_, new_n810_, new_n808_, new_n907_, new_n665_, new_n800_, new_n897_, new_n1012_, new_n719_, new_n869_, new_n1178_, new_n270_, new_n570_, new_n598_, new_n893_, new_n1063_, new_n520_, new_n1001_, new_n253_, new_n825_, new_n557_, new_n260_, new_n251_, new_n300_, new_n507_, new_n741_, new_n806_, new_n605_, new_n1074_, new_n748_, new_n1137_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n1141_, new_n807_, new_n592_, new_n726_, new_n1123_, new_n231_, new_n583_, new_n617_, new_n1080_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n199_, new_n487_, new_n360_, new_n675_, new_n1155_, new_n1186_, new_n191_, new_n225_, new_n922_, new_n387_, new_n476_, new_n987_, new_n949_, new_n221_, new_n243_, new_n450_, new_n1179_, new_n298_, new_n184_, new_n1088_, new_n1148_, new_n1146_, new_n569_, new_n555_, new_n174_, new_n468_, new_n977_, new_n1139_, new_n782_, new_n444_, new_n392_, new_n518_, new_n950_, new_n737_, new_n1022_, new_n340_, new_n285_, new_n692_, new_n502_, new_n209_, new_n623_, new_n446_, new_n203_, new_n316_, new_n590_, new_n826_, new_n789_, new_n515_, new_n332_, new_n972_, new_n1067_, new_n891_, new_n516_, new_n733_, new_n1021_, new_n1076_, new_n585_, new_n312_, new_n535_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n307_, new_n190_, new_n1181_, new_n597_, new_n1093_, new_n1092_, new_n1143_, new_n1072_, new_n1190_, new_n1097_, new_n1069_, new_n651_, new_n1164_, new_n435_, new_n1010_, new_n776_, new_n687_, new_n370_, new_n1029_, new_n638_, new_n523_, new_n909_, new_n217_, new_n788_, new_n841_, new_n1204_, new_n1112_, new_n711_, new_n1156_, new_n731_, new_n930_, new_n973_, new_n412_, new_n607_, new_n645_, new_n1087_, new_n723_, new_n756_, new_n823_, new_n574_, new_n928_, new_n319_, new_n1008_, new_n338_, new_n707_, new_n740_, new_n957_, new_n1047_, new_n787_, new_n1134_, new_n336_, new_n247_, new_n539_, new_n803_, new_n330_, new_n727_, new_n294_, new_n1173_, new_n704_, new_n1189_, new_n1197_, new_n474_, new_n1129_, new_n467_, new_n1013_, new_n404_, new_n1077_, new_n193_, new_n490_, new_n560_, new_n1100_, new_n865_, new_n358_, new_n877_, new_n545_, new_n228_, new_n611_, new_n289_, new_n1011_, new_n425_, new_n896_, new_n802_, new_n866_, new_n947_, new_n994_, new_n982_, new_n964_, new_n1078_, new_n551_, new_n279_, new_n455_, new_n618_, new_n1140_, new_n1042_, new_n863_, new_n828_, new_n980_, new_n464_, new_n204_, new_n181_, new_n573_, new_n765_, new_n1103_;

not g0000 ( new_n172_, keyIn_0_36 );
not g0001 ( new_n173_, keyIn_0_27 );
not g0002 ( new_n174_, N108 );
and g0003 ( new_n175_, keyIn_0_16, N102 );
not g0004 ( new_n176_, new_n175_ );
or g0005 ( new_n177_, keyIn_0_16, N102 );
and g0006 ( new_n178_, new_n176_, new_n177_ );
or g0007 ( new_n179_, new_n178_, new_n174_ );
or g0008 ( new_n180_, new_n179_, new_n173_ );
and g0009 ( new_n181_, new_n179_, new_n173_ );
not g0010 ( new_n182_, new_n181_ );
and g0011 ( new_n183_, new_n182_, new_n180_ );
not g0012 ( new_n184_, keyIn_0_25 );
not g0013 ( new_n185_, N82 );
not g0014 ( new_n186_, N76 );
and g0015 ( new_n187_, new_n186_, keyIn_0_12 );
not g0016 ( new_n188_, new_n187_ );
or g0017 ( new_n189_, new_n186_, keyIn_0_12 );
and g0018 ( new_n190_, new_n188_, new_n189_ );
or g0019 ( new_n191_, new_n190_, new_n185_ );
or g0020 ( new_n192_, new_n191_, new_n184_ );
and g0021 ( new_n193_, new_n191_, new_n184_ );
not g0022 ( new_n194_, new_n193_ );
and g0023 ( new_n195_, new_n194_, new_n192_ );
not g0024 ( new_n196_, N89 );
and g0025 ( new_n197_, new_n196_, keyIn_0_14 );
not g0026 ( new_n198_, new_n197_ );
or g0027 ( new_n199_, new_n196_, keyIn_0_14 );
and g0028 ( new_n200_, new_n199_, N95 );
and g0029 ( new_n201_, new_n200_, new_n198_ );
not g0030 ( new_n202_, new_n201_ );
and g0031 ( new_n203_, new_n202_, keyIn_0_26 );
not g0032 ( new_n204_, keyIn_0_26 );
and g0033 ( new_n205_, new_n201_, new_n204_ );
or g0034 ( new_n206_, new_n203_, new_n205_ );
not g0035 ( new_n207_, new_n206_ );
or g0036 ( new_n208_, new_n207_, new_n195_ );
or g0037 ( new_n209_, new_n208_, new_n183_ );
not g0038 ( new_n210_, keyIn_0_21 );
not g0039 ( new_n211_, N30 );
or g0040 ( new_n212_, keyIn_0_4, N24 );
and g0041 ( new_n213_, keyIn_0_4, N24 );
not g0042 ( new_n214_, new_n213_ );
and g0043 ( new_n215_, new_n214_, new_n212_ );
or g0044 ( new_n216_, new_n215_, new_n211_ );
and g0045 ( new_n217_, new_n216_, new_n210_ );
not g0046 ( new_n218_, new_n217_ );
or g0047 ( new_n219_, new_n216_, new_n210_ );
and g0048 ( new_n220_, new_n218_, new_n219_ );
not g0049 ( new_n221_, keyIn_0_23 );
not g0050 ( new_n222_, N56 );
or g0051 ( new_n223_, keyIn_0_8, N50 );
and g0052 ( new_n224_, keyIn_0_8, N50 );
not g0053 ( new_n225_, new_n224_ );
and g0054 ( new_n226_, new_n225_, new_n223_ );
or g0055 ( new_n227_, new_n226_, new_n222_ );
and g0056 ( new_n228_, new_n227_, new_n221_ );
not g0057 ( new_n229_, new_n228_ );
or g0058 ( new_n230_, new_n227_, new_n221_ );
and g0059 ( new_n231_, new_n229_, new_n230_ );
and g0060 ( new_n232_, new_n220_, new_n231_ );
not g0061 ( new_n233_, new_n232_ );
not g0062 ( new_n234_, N37 );
and g0063 ( new_n235_, new_n234_, keyIn_0_6 );
not g0064 ( new_n236_, new_n235_ );
or g0065 ( new_n237_, new_n234_, keyIn_0_6 );
and g0066 ( new_n238_, new_n237_, N43 );
and g0067 ( new_n239_, new_n238_, new_n236_ );
or g0068 ( new_n240_, new_n239_, keyIn_0_22 );
not g0069 ( new_n241_, keyIn_0_22 );
not g0070 ( new_n242_, N43 );
not g0071 ( new_n243_, keyIn_0_6 );
and g0072 ( new_n244_, new_n243_, N37 );
or g0073 ( new_n245_, new_n244_, new_n242_ );
or g0074 ( new_n246_, new_n245_, new_n235_ );
or g0075 ( new_n247_, new_n246_, new_n241_ );
and g0076 ( new_n248_, new_n247_, new_n240_ );
or g0077 ( new_n249_, keyIn_0_10, N63 );
not g0078 ( new_n250_, new_n249_ );
not g0079 ( new_n251_, N69 );
and g0080 ( new_n252_, keyIn_0_10, N63 );
or g0081 ( new_n253_, new_n252_, new_n251_ );
or g0082 ( new_n254_, new_n253_, new_n250_ );
or g0083 ( new_n255_, new_n254_, keyIn_0_24 );
not g0084 ( new_n256_, keyIn_0_24 );
not g0085 ( new_n257_, new_n252_ );
and g0086 ( new_n258_, new_n257_, N69 );
and g0087 ( new_n259_, new_n258_, new_n249_ );
or g0088 ( new_n260_, new_n259_, new_n256_ );
and g0089 ( new_n261_, new_n260_, new_n255_ );
or g0090 ( new_n262_, new_n248_, new_n261_ );
not g0091 ( new_n263_, N4 );
not g0092 ( new_n264_, keyIn_0_0 );
or g0093 ( new_n265_, new_n264_, N1 );
not g0094 ( new_n266_, N1 );
or g0095 ( new_n267_, new_n266_, keyIn_0_0 );
and g0096 ( new_n268_, new_n265_, new_n267_ );
or g0097 ( new_n269_, new_n268_, new_n263_ );
and g0098 ( new_n270_, new_n269_, keyIn_0_18 );
not g0099 ( new_n271_, keyIn_0_18 );
and g0100 ( new_n272_, new_n266_, keyIn_0_0 );
and g0101 ( new_n273_, new_n264_, N1 );
or g0102 ( new_n274_, new_n272_, new_n273_ );
and g0103 ( new_n275_, new_n274_, N4 );
and g0104 ( new_n276_, new_n275_, new_n271_ );
or g0105 ( new_n277_, new_n270_, new_n276_ );
and g0106 ( new_n278_, keyIn_0_2, N11 );
not g0107 ( new_n279_, keyIn_0_2 );
not g0108 ( new_n280_, N11 );
and g0109 ( new_n281_, new_n279_, new_n280_ );
or g0110 ( new_n282_, new_n281_, new_n278_ );
and g0111 ( new_n283_, new_n282_, N17 );
or g0112 ( new_n284_, new_n283_, keyIn_0_20 );
not g0113 ( new_n285_, keyIn_0_20 );
not g0114 ( new_n286_, N17 );
not g0115 ( new_n287_, new_n278_ );
or g0116 ( new_n288_, keyIn_0_2, N11 );
and g0117 ( new_n289_, new_n287_, new_n288_ );
or g0118 ( new_n290_, new_n289_, new_n286_ );
or g0119 ( new_n291_, new_n290_, new_n285_ );
and g0120 ( new_n292_, new_n284_, new_n291_ );
or g0121 ( new_n293_, new_n277_, new_n292_ );
or g0122 ( new_n294_, new_n293_, new_n262_ );
or g0123 ( new_n295_, new_n294_, new_n233_ );
or g0124 ( new_n296_, new_n295_, new_n209_ );
and g0125 ( new_n297_, new_n296_, new_n172_ );
not g0126 ( new_n298_, new_n183_ );
not g0127 ( new_n299_, new_n192_ );
or g0128 ( new_n300_, new_n299_, new_n193_ );
and g0129 ( new_n301_, new_n300_, new_n206_ );
and g0130 ( new_n302_, new_n301_, new_n298_ );
and g0131 ( new_n303_, new_n246_, new_n241_ );
and g0132 ( new_n304_, new_n239_, keyIn_0_22 );
or g0133 ( new_n305_, new_n303_, new_n304_ );
and g0134 ( new_n306_, new_n259_, new_n256_ );
and g0135 ( new_n307_, new_n254_, keyIn_0_24 );
or g0136 ( new_n308_, new_n306_, new_n307_ );
and g0137 ( new_n309_, new_n305_, new_n308_ );
or g0138 ( new_n310_, new_n275_, new_n271_ );
or g0139 ( new_n311_, new_n269_, keyIn_0_18 );
and g0140 ( new_n312_, new_n311_, new_n310_ );
and g0141 ( new_n313_, new_n290_, new_n285_ );
and g0142 ( new_n314_, new_n283_, keyIn_0_20 );
or g0143 ( new_n315_, new_n313_, new_n314_ );
and g0144 ( new_n316_, new_n312_, new_n315_ );
and g0145 ( new_n317_, new_n316_, new_n309_ );
and g0146 ( new_n318_, new_n317_, new_n232_ );
and g0147 ( new_n319_, new_n318_, new_n302_ );
and g0148 ( new_n320_, new_n319_, keyIn_0_36 );
or g0149 ( N223, new_n297_, new_n320_ );
not g0150 ( new_n322_, keyIn_0_60 );
not g0151 ( new_n323_, keyIn_0_42 );
and g0152 ( new_n324_, N223, keyIn_0_37 );
not g0153 ( new_n325_, keyIn_0_37 );
or g0154 ( new_n326_, new_n319_, keyIn_0_36 );
not g0155 ( new_n327_, new_n320_ );
and g0156 ( new_n328_, new_n327_, new_n326_ );
and g0157 ( new_n329_, new_n328_, new_n325_ );
or g0158 ( new_n330_, new_n324_, new_n329_ );
and g0159 ( new_n331_, new_n330_, new_n231_ );
not g0160 ( new_n332_, new_n231_ );
or g0161 ( new_n333_, new_n328_, new_n325_ );
or g0162 ( new_n334_, N223, keyIn_0_37 );
and g0163 ( new_n335_, new_n334_, new_n333_ );
and g0164 ( new_n336_, new_n335_, new_n332_ );
or g0165 ( new_n337_, new_n331_, new_n336_ );
and g0166 ( new_n338_, new_n337_, new_n323_ );
not g0167 ( new_n339_, new_n338_ );
or g0168 ( new_n340_, new_n337_, new_n323_ );
and g0169 ( new_n341_, new_n339_, new_n340_ );
or g0170 ( new_n342_, keyIn_0_9, N56 );
not g0171 ( new_n343_, N60 );
and g0172 ( new_n344_, keyIn_0_9, N56 );
not g0173 ( new_n345_, new_n344_ );
and g0174 ( new_n346_, new_n345_, new_n343_ );
and g0175 ( new_n347_, new_n346_, new_n342_ );
and g0176 ( new_n348_, new_n347_, keyIn_0_31 );
not g0177 ( new_n349_, new_n348_ );
or g0178 ( new_n350_, new_n347_, keyIn_0_31 );
and g0179 ( new_n351_, new_n349_, new_n350_ );
or g0180 ( new_n352_, new_n341_, new_n351_ );
not g0181 ( new_n353_, new_n352_ );
or g0182 ( new_n354_, new_n353_, keyIn_0_52 );
not g0183 ( new_n355_, keyIn_0_52 );
or g0184 ( new_n356_, new_n352_, new_n355_ );
and g0185 ( new_n357_, new_n354_, new_n356_ );
and g0186 ( new_n358_, new_n330_, new_n308_ );
and g0187 ( new_n359_, new_n335_, new_n261_ );
or g0188 ( new_n360_, new_n358_, new_n359_ );
and g0189 ( new_n361_, new_n360_, keyIn_0_43 );
not g0190 ( new_n362_, new_n361_ );
or g0191 ( new_n363_, new_n360_, keyIn_0_43 );
and g0192 ( new_n364_, new_n362_, new_n363_ );
not g0193 ( new_n365_, N73 );
and g0194 ( new_n366_, new_n251_, keyIn_0_11 );
not g0195 ( new_n367_, new_n366_ );
or g0196 ( new_n368_, new_n251_, keyIn_0_11 );
and g0197 ( new_n369_, new_n367_, new_n368_ );
not g0198 ( new_n370_, new_n369_ );
and g0199 ( new_n371_, new_n370_, new_n365_ );
not g0200 ( new_n372_, new_n371_ );
and g0201 ( new_n373_, new_n372_, keyIn_0_32 );
not g0202 ( new_n374_, new_n373_ );
or g0203 ( new_n375_, new_n372_, keyIn_0_32 );
and g0204 ( new_n376_, new_n374_, new_n375_ );
or g0205 ( new_n377_, new_n364_, new_n376_ );
not g0206 ( new_n378_, new_n377_ );
and g0207 ( new_n379_, new_n378_, keyIn_0_53 );
not g0208 ( new_n380_, keyIn_0_53 );
and g0209 ( new_n381_, new_n377_, new_n380_ );
or g0210 ( new_n382_, new_n379_, new_n381_ );
not g0211 ( new_n383_, keyIn_0_51 );
not g0212 ( new_n384_, keyIn_0_41 );
and g0213 ( new_n385_, new_n330_, new_n305_ );
and g0214 ( new_n386_, new_n335_, new_n248_ );
or g0215 ( new_n387_, new_n385_, new_n386_ );
and g0216 ( new_n388_, new_n387_, new_n384_ );
not g0217 ( new_n389_, new_n388_ );
or g0218 ( new_n390_, new_n387_, new_n384_ );
and g0219 ( new_n391_, new_n389_, new_n390_ );
not g0220 ( new_n392_, keyIn_0_30 );
not g0221 ( new_n393_, N47 );
and g0222 ( new_n394_, new_n242_, keyIn_0_7 );
not g0223 ( new_n395_, new_n394_ );
or g0224 ( new_n396_, new_n242_, keyIn_0_7 );
and g0225 ( new_n397_, new_n395_, new_n396_ );
not g0226 ( new_n398_, new_n397_ );
and g0227 ( new_n399_, new_n398_, new_n393_ );
and g0228 ( new_n400_, new_n399_, new_n392_ );
not g0229 ( new_n401_, new_n400_ );
or g0230 ( new_n402_, new_n399_, new_n392_ );
and g0231 ( new_n403_, new_n401_, new_n402_ );
not g0232 ( new_n404_, new_n403_ );
or g0233 ( new_n405_, new_n391_, new_n404_ );
not g0234 ( new_n406_, new_n405_ );
or g0235 ( new_n407_, new_n406_, new_n383_ );
or g0236 ( new_n408_, new_n405_, keyIn_0_51 );
and g0237 ( new_n409_, new_n407_, new_n408_ );
and g0238 ( new_n410_, new_n382_, new_n409_ );
and g0239 ( new_n411_, new_n410_, new_n357_ );
and g0240 ( new_n412_, new_n330_, new_n300_ );
and g0241 ( new_n413_, new_n335_, new_n195_ );
or g0242 ( new_n414_, new_n412_, new_n413_ );
not g0243 ( new_n415_, new_n414_ );
and g0244 ( new_n416_, new_n415_, keyIn_0_44 );
not g0245 ( new_n417_, keyIn_0_44 );
and g0246 ( new_n418_, new_n414_, new_n417_ );
or g0247 ( new_n419_, new_n416_, new_n418_ );
not g0248 ( new_n420_, keyIn_0_33 );
not g0249 ( new_n421_, N86 );
and g0250 ( new_n422_, new_n185_, keyIn_0_13 );
not g0251 ( new_n423_, new_n422_ );
or g0252 ( new_n424_, new_n185_, keyIn_0_13 );
and g0253 ( new_n425_, new_n423_, new_n424_ );
and g0254 ( new_n426_, new_n425_, new_n421_ );
not g0255 ( new_n427_, new_n426_ );
and g0256 ( new_n428_, new_n427_, new_n420_ );
and g0257 ( new_n429_, new_n426_, keyIn_0_33 );
or g0258 ( new_n430_, new_n428_, new_n429_ );
not g0259 ( new_n431_, new_n430_ );
and g0260 ( new_n432_, new_n419_, new_n431_ );
not g0261 ( new_n433_, new_n432_ );
and g0262 ( new_n434_, new_n433_, keyIn_0_54 );
not g0263 ( new_n435_, keyIn_0_54 );
and g0264 ( new_n436_, new_n432_, new_n435_ );
or g0265 ( new_n437_, new_n434_, new_n436_ );
and g0266 ( new_n438_, new_n330_, new_n298_ );
and g0267 ( new_n439_, new_n335_, new_n183_ );
or g0268 ( new_n440_, new_n438_, new_n439_ );
and g0269 ( new_n441_, new_n440_, keyIn_0_47 );
not g0270 ( new_n442_, new_n441_ );
or g0271 ( new_n443_, new_n440_, keyIn_0_47 );
and g0272 ( new_n444_, new_n442_, new_n443_ );
not g0273 ( new_n445_, keyIn_0_35 );
not g0274 ( new_n446_, N112 );
and g0275 ( new_n447_, new_n174_, keyIn_0_17 );
not g0276 ( new_n448_, new_n447_ );
or g0277 ( new_n449_, new_n174_, keyIn_0_17 );
and g0278 ( new_n450_, new_n448_, new_n449_ );
and g0279 ( new_n451_, new_n450_, new_n446_ );
and g0280 ( new_n452_, new_n451_, new_n445_ );
not g0281 ( new_n453_, new_n452_ );
or g0282 ( new_n454_, new_n451_, new_n445_ );
and g0283 ( new_n455_, new_n453_, new_n454_ );
and g0284 ( new_n456_, new_n444_, new_n455_ );
not g0285 ( new_n457_, new_n456_ );
and g0286 ( new_n458_, new_n457_, keyIn_0_56 );
not g0287 ( new_n459_, keyIn_0_56 );
and g0288 ( new_n460_, new_n456_, new_n459_ );
or g0289 ( new_n461_, new_n458_, new_n460_ );
and g0290 ( new_n462_, new_n437_, new_n461_ );
and g0291 ( new_n463_, new_n330_, new_n220_ );
not g0292 ( new_n464_, new_n220_ );
and g0293 ( new_n465_, new_n335_, new_n464_ );
or g0294 ( new_n466_, new_n463_, new_n465_ );
or g0295 ( new_n467_, new_n466_, keyIn_0_40 );
not g0296 ( new_n468_, keyIn_0_40 );
or g0297 ( new_n469_, new_n335_, new_n464_ );
or g0298 ( new_n470_, new_n330_, new_n220_ );
and g0299 ( new_n471_, new_n470_, new_n469_ );
or g0300 ( new_n472_, new_n471_, new_n468_ );
and g0301 ( new_n473_, new_n467_, new_n472_ );
not g0302 ( new_n474_, N34 );
and g0303 ( new_n475_, keyIn_0_5, N30 );
not g0304 ( new_n476_, new_n475_ );
or g0305 ( new_n477_, keyIn_0_5, N30 );
and g0306 ( new_n478_, new_n476_, new_n477_ );
not g0307 ( new_n479_, new_n478_ );
and g0308 ( new_n480_, new_n479_, new_n474_ );
not g0309 ( new_n481_, new_n480_ );
and g0310 ( new_n482_, new_n481_, keyIn_0_29 );
not g0311 ( new_n483_, new_n482_ );
or g0312 ( new_n484_, new_n481_, keyIn_0_29 );
and g0313 ( new_n485_, new_n483_, new_n484_ );
not g0314 ( new_n486_, new_n485_ );
or g0315 ( new_n487_, new_n473_, new_n486_ );
and g0316 ( new_n488_, new_n487_, keyIn_0_50 );
not g0317 ( new_n489_, keyIn_0_50 );
and g0318 ( new_n490_, new_n471_, new_n468_ );
and g0319 ( new_n491_, new_n466_, keyIn_0_40 );
or g0320 ( new_n492_, new_n491_, new_n490_ );
and g0321 ( new_n493_, new_n492_, new_n485_ );
and g0322 ( new_n494_, new_n493_, new_n489_ );
or g0323 ( new_n495_, new_n488_, new_n494_ );
not g0324 ( new_n496_, keyIn_0_55 );
not g0325 ( new_n497_, keyIn_0_46 );
and g0326 ( new_n498_, new_n330_, new_n206_ );
and g0327 ( new_n499_, new_n335_, new_n207_ );
or g0328 ( new_n500_, new_n498_, new_n499_ );
or g0329 ( new_n501_, new_n500_, new_n497_ );
or g0330 ( new_n502_, new_n335_, new_n207_ );
or g0331 ( new_n503_, new_n330_, new_n206_ );
and g0332 ( new_n504_, new_n503_, new_n502_ );
or g0333 ( new_n505_, new_n504_, keyIn_0_46 );
and g0334 ( new_n506_, new_n501_, new_n505_ );
not g0335 ( new_n507_, N99 );
not g0336 ( new_n508_, N95 );
and g0337 ( new_n509_, new_n508_, keyIn_0_15 );
not g0338 ( new_n510_, new_n509_ );
or g0339 ( new_n511_, new_n508_, keyIn_0_15 );
and g0340 ( new_n512_, new_n510_, new_n511_ );
not g0341 ( new_n513_, new_n512_ );
and g0342 ( new_n514_, new_n513_, new_n507_ );
not g0343 ( new_n515_, new_n514_ );
and g0344 ( new_n516_, new_n515_, keyIn_0_34 );
not g0345 ( new_n517_, new_n516_ );
or g0346 ( new_n518_, new_n515_, keyIn_0_34 );
and g0347 ( new_n519_, new_n517_, new_n518_ );
or g0348 ( new_n520_, new_n506_, new_n519_ );
or g0349 ( new_n521_, new_n520_, new_n496_ );
and g0350 ( new_n522_, new_n504_, keyIn_0_46 );
and g0351 ( new_n523_, new_n500_, new_n497_ );
or g0352 ( new_n524_, new_n523_, new_n522_ );
not g0353 ( new_n525_, new_n519_ );
and g0354 ( new_n526_, new_n524_, new_n525_ );
or g0355 ( new_n527_, new_n526_, keyIn_0_55 );
and g0356 ( new_n528_, new_n521_, new_n527_ );
and g0357 ( new_n529_, new_n495_, new_n528_ );
not g0358 ( new_n530_, keyIn_0_48 );
not g0359 ( new_n531_, keyIn_0_38 );
and g0360 ( new_n532_, new_n330_, new_n312_ );
and g0361 ( new_n533_, new_n335_, new_n277_ );
or g0362 ( new_n534_, new_n532_, new_n533_ );
or g0363 ( new_n535_, new_n534_, new_n531_ );
or g0364 ( new_n536_, new_n335_, new_n277_ );
or g0365 ( new_n537_, new_n330_, new_n312_ );
and g0366 ( new_n538_, new_n537_, new_n536_ );
or g0367 ( new_n539_, new_n538_, keyIn_0_38 );
and g0368 ( new_n540_, new_n535_, new_n539_ );
not g0369 ( new_n541_, N8 );
and g0370 ( new_n542_, new_n263_, keyIn_0_1 );
not g0371 ( new_n543_, new_n542_ );
or g0372 ( new_n544_, new_n263_, keyIn_0_1 );
and g0373 ( new_n545_, new_n543_, new_n544_ );
and g0374 ( new_n546_, new_n545_, new_n541_ );
and g0375 ( new_n547_, new_n546_, keyIn_0_19 );
not g0376 ( new_n548_, new_n547_ );
or g0377 ( new_n549_, new_n546_, keyIn_0_19 );
and g0378 ( new_n550_, new_n548_, new_n549_ );
and g0379 ( new_n551_, new_n540_, new_n550_ );
and g0380 ( new_n552_, new_n551_, new_n530_ );
and g0381 ( new_n553_, new_n538_, keyIn_0_38 );
and g0382 ( new_n554_, new_n534_, new_n531_ );
or g0383 ( new_n555_, new_n554_, new_n553_ );
not g0384 ( new_n556_, new_n550_ );
or g0385 ( new_n557_, new_n555_, new_n556_ );
and g0386 ( new_n558_, new_n557_, keyIn_0_48 );
or g0387 ( new_n559_, new_n558_, new_n552_ );
not g0388 ( new_n560_, keyIn_0_39 );
and g0389 ( new_n561_, new_n330_, new_n315_ );
and g0390 ( new_n562_, new_n335_, new_n292_ );
or g0391 ( new_n563_, new_n561_, new_n562_ );
or g0392 ( new_n564_, new_n563_, new_n560_ );
or g0393 ( new_n565_, new_n335_, new_n292_ );
or g0394 ( new_n566_, new_n330_, new_n315_ );
and g0395 ( new_n567_, new_n566_, new_n565_ );
or g0396 ( new_n568_, new_n567_, keyIn_0_39 );
and g0397 ( new_n569_, new_n564_, new_n568_ );
not g0398 ( new_n570_, N21 );
and g0399 ( new_n571_, keyIn_0_3, N17 );
not g0400 ( new_n572_, new_n571_ );
or g0401 ( new_n573_, keyIn_0_3, N17 );
and g0402 ( new_n574_, new_n572_, new_n573_ );
not g0403 ( new_n575_, new_n574_ );
and g0404 ( new_n576_, new_n575_, new_n570_ );
not g0405 ( new_n577_, new_n576_ );
and g0406 ( new_n578_, new_n577_, keyIn_0_28 );
not g0407 ( new_n579_, new_n578_ );
or g0408 ( new_n580_, new_n577_, keyIn_0_28 );
and g0409 ( new_n581_, new_n579_, new_n580_ );
and g0410 ( new_n582_, new_n569_, new_n581_ );
and g0411 ( new_n583_, new_n582_, keyIn_0_49 );
not g0412 ( new_n584_, keyIn_0_49 );
and g0413 ( new_n585_, new_n567_, keyIn_0_39 );
and g0414 ( new_n586_, new_n563_, new_n560_ );
or g0415 ( new_n587_, new_n586_, new_n585_ );
not g0416 ( new_n588_, new_n581_ );
or g0417 ( new_n589_, new_n587_, new_n588_ );
and g0418 ( new_n590_, new_n589_, new_n584_ );
or g0419 ( new_n591_, new_n590_, new_n583_ );
and g0420 ( new_n592_, new_n559_, new_n591_ );
and g0421 ( new_n593_, new_n592_, new_n529_ );
and g0422 ( new_n594_, new_n593_, new_n462_ );
and g0423 ( new_n595_, new_n594_, new_n411_ );
not g0424 ( new_n596_, new_n595_ );
and g0425 ( new_n597_, new_n596_, new_n322_ );
and g0426 ( new_n598_, new_n595_, keyIn_0_60 );
or g0427 ( N329, new_n597_, new_n598_ );
not g0428 ( new_n600_, keyIn_0_95 );
not g0429 ( new_n601_, keyIn_0_66 );
not g0430 ( new_n602_, new_n559_ );
not g0431 ( new_n603_, keyIn_0_64 );
and g0432 ( new_n604_, N329, new_n603_ );
or g0433 ( new_n605_, new_n595_, keyIn_0_60 );
not g0434 ( new_n606_, new_n598_ );
and g0435 ( new_n607_, new_n606_, new_n605_ );
and g0436 ( new_n608_, new_n607_, keyIn_0_64 );
or g0437 ( new_n609_, new_n604_, new_n608_ );
and g0438 ( new_n610_, new_n609_, new_n602_ );
or g0439 ( new_n611_, new_n607_, keyIn_0_64 );
or g0440 ( new_n612_, N329, new_n603_ );
and g0441 ( new_n613_, new_n612_, new_n611_ );
and g0442 ( new_n614_, new_n613_, new_n559_ );
or g0443 ( new_n615_, new_n610_, new_n614_ );
and g0444 ( new_n616_, new_n615_, new_n601_ );
not g0445 ( new_n617_, new_n616_ );
or g0446 ( new_n618_, new_n615_, new_n601_ );
and g0447 ( new_n619_, new_n617_, new_n618_ );
not g0448 ( new_n620_, new_n619_ );
not g0449 ( new_n621_, N14 );
and g0450 ( new_n622_, new_n545_, new_n621_ );
and g0451 ( new_n623_, new_n540_, new_n622_ );
and g0452 ( new_n624_, new_n620_, new_n623_ );
not g0453 ( new_n625_, new_n624_ );
and g0454 ( new_n626_, new_n625_, keyIn_0_84 );
not g0455 ( new_n627_, keyIn_0_84 );
and g0456 ( new_n628_, new_n624_, new_n627_ );
or g0457 ( new_n629_, new_n626_, new_n628_ );
not g0458 ( new_n630_, keyIn_0_77 );
not g0459 ( new_n631_, new_n528_ );
and g0460 ( new_n632_, new_n609_, new_n631_ );
and g0461 ( new_n633_, new_n613_, new_n528_ );
or g0462 ( new_n634_, new_n632_, new_n633_ );
and g0463 ( new_n635_, new_n634_, new_n630_ );
not g0464 ( new_n636_, new_n635_ );
or g0465 ( new_n637_, new_n634_, new_n630_ );
and g0466 ( new_n638_, new_n636_, new_n637_ );
not g0467 ( new_n639_, N105 );
and g0468 ( new_n640_, new_n513_, new_n639_ );
and g0469 ( new_n641_, new_n524_, new_n640_ );
and g0470 ( new_n642_, new_n641_, keyIn_0_59 );
not g0471 ( new_n643_, new_n642_ );
or g0472 ( new_n644_, new_n641_, keyIn_0_59 );
and g0473 ( new_n645_, new_n643_, new_n644_ );
not g0474 ( new_n646_, new_n645_ );
and g0475 ( new_n647_, new_n646_, keyIn_0_63 );
not g0476 ( new_n648_, new_n647_ );
or g0477 ( new_n649_, new_n646_, keyIn_0_63 );
and g0478 ( new_n650_, new_n648_, new_n649_ );
or g0479 ( new_n651_, new_n638_, new_n650_ );
not g0480 ( new_n652_, new_n651_ );
and g0481 ( new_n653_, new_n652_, keyIn_0_91 );
not g0482 ( new_n654_, keyIn_0_91 );
and g0483 ( new_n655_, new_n651_, new_n654_ );
or g0484 ( new_n656_, new_n653_, new_n655_ );
not g0485 ( new_n657_, keyIn_0_85 );
not g0486 ( new_n658_, keyIn_0_67 );
and g0487 ( new_n659_, new_n613_, new_n591_ );
not g0488 ( new_n660_, new_n659_ );
or g0489 ( new_n661_, new_n613_, new_n591_ );
and g0490 ( new_n662_, new_n660_, new_n661_ );
and g0491 ( new_n663_, new_n662_, new_n658_ );
not g0492 ( new_n664_, new_n663_ );
or g0493 ( new_n665_, new_n662_, new_n658_ );
not g0494 ( new_n666_, N27 );
and g0495 ( new_n667_, new_n575_, new_n666_ );
and g0496 ( new_n668_, new_n569_, new_n667_ );
and g0497 ( new_n669_, new_n665_, new_n668_ );
and g0498 ( new_n670_, new_n669_, new_n664_ );
not g0499 ( new_n671_, new_n670_ );
and g0500 ( new_n672_, new_n671_, new_n657_ );
and g0501 ( new_n673_, new_n670_, keyIn_0_85 );
or g0502 ( new_n674_, new_n672_, new_n673_ );
and g0503 ( new_n675_, new_n656_, new_n674_ );
and g0504 ( new_n676_, new_n675_, new_n629_ );
not g0505 ( new_n677_, keyIn_0_86 );
not g0506 ( new_n678_, new_n495_ );
and g0507 ( new_n679_, new_n609_, new_n678_ );
and g0508 ( new_n680_, new_n613_, new_n495_ );
or g0509 ( new_n681_, new_n679_, new_n680_ );
and g0510 ( new_n682_, new_n681_, keyIn_0_68 );
not g0511 ( new_n683_, new_n682_ );
or g0512 ( new_n684_, new_n681_, keyIn_0_68 );
and g0513 ( new_n685_, new_n683_, new_n684_ );
not g0514 ( new_n686_, N40 );
and g0515 ( new_n687_, new_n479_, new_n686_ );
and g0516 ( new_n688_, new_n492_, new_n687_ );
not g0517 ( new_n689_, new_n688_ );
or g0518 ( new_n690_, new_n685_, new_n689_ );
not g0519 ( new_n691_, new_n690_ );
or g0520 ( new_n692_, new_n691_, new_n677_ );
and g0521 ( new_n693_, new_n613_, new_n409_ );
not g0522 ( new_n694_, new_n693_ );
or g0523 ( new_n695_, new_n613_, new_n409_ );
and g0524 ( new_n696_, new_n694_, new_n695_ );
not g0525 ( new_n697_, new_n696_ );
and g0526 ( new_n698_, new_n697_, keyIn_0_69 );
not g0527 ( new_n699_, keyIn_0_69 );
and g0528 ( new_n700_, new_n696_, new_n699_ );
not g0529 ( new_n701_, new_n391_ );
not g0530 ( new_n702_, N53 );
and g0531 ( new_n703_, new_n398_, new_n702_ );
and g0532 ( new_n704_, new_n701_, new_n703_ );
not g0533 ( new_n705_, new_n704_ );
or g0534 ( new_n706_, new_n700_, new_n705_ );
or g0535 ( new_n707_, new_n706_, new_n698_ );
not g0536 ( new_n708_, new_n707_ );
or g0537 ( new_n709_, new_n708_, keyIn_0_87 );
and g0538 ( new_n710_, new_n692_, new_n709_ );
or g0539 ( new_n711_, new_n690_, keyIn_0_86 );
not g0540 ( new_n712_, keyIn_0_87 );
or g0541 ( new_n713_, new_n707_, new_n712_ );
and g0542 ( new_n714_, new_n711_, new_n713_ );
and g0543 ( new_n715_, new_n710_, new_n714_ );
not g0544 ( new_n716_, keyIn_0_90 );
or g0545 ( new_n717_, new_n613_, new_n437_ );
not g0546 ( new_n718_, new_n437_ );
or g0547 ( new_n719_, new_n609_, new_n718_ );
and g0548 ( new_n720_, new_n719_, new_n717_ );
and g0549 ( new_n721_, new_n720_, keyIn_0_75 );
not g0550 ( new_n722_, keyIn_0_75 );
and g0551 ( new_n723_, new_n609_, new_n718_ );
and g0552 ( new_n724_, new_n613_, new_n437_ );
or g0553 ( new_n725_, new_n723_, new_n724_ );
and g0554 ( new_n726_, new_n725_, new_n722_ );
not g0555 ( new_n727_, N92 );
and g0556 ( new_n728_, new_n425_, new_n727_ );
and g0557 ( new_n729_, new_n419_, new_n728_ );
not g0558 ( new_n730_, new_n729_ );
or g0559 ( new_n731_, new_n726_, new_n730_ );
or g0560 ( new_n732_, new_n731_, new_n721_ );
or g0561 ( new_n733_, new_n732_, new_n716_ );
not g0562 ( new_n734_, keyIn_0_92 );
not g0563 ( new_n735_, new_n461_ );
and g0564 ( new_n736_, new_n609_, new_n735_ );
and g0565 ( new_n737_, new_n613_, new_n461_ );
or g0566 ( new_n738_, new_n736_, new_n737_ );
or g0567 ( new_n739_, new_n738_, keyIn_0_79 );
not g0568 ( new_n740_, keyIn_0_79 );
or g0569 ( new_n741_, new_n613_, new_n461_ );
or g0570 ( new_n742_, new_n609_, new_n735_ );
and g0571 ( new_n743_, new_n742_, new_n741_ );
or g0572 ( new_n744_, new_n743_, new_n740_ );
and g0573 ( new_n745_, new_n739_, new_n744_ );
not g0574 ( new_n746_, N115 );
and g0575 ( new_n747_, new_n450_, new_n746_ );
and g0576 ( new_n748_, new_n444_, new_n747_ );
not g0577 ( new_n749_, new_n748_ );
or g0578 ( new_n750_, new_n745_, new_n749_ );
or g0579 ( new_n751_, new_n750_, new_n734_ );
and g0580 ( new_n752_, new_n733_, new_n751_ );
and g0581 ( new_n753_, new_n743_, new_n740_ );
and g0582 ( new_n754_, new_n738_, keyIn_0_79 );
or g0583 ( new_n755_, new_n754_, new_n753_ );
and g0584 ( new_n756_, new_n755_, new_n748_ );
or g0585 ( new_n757_, new_n756_, keyIn_0_92 );
not g0586 ( new_n758_, new_n721_ );
or g0587 ( new_n759_, new_n720_, keyIn_0_75 );
and g0588 ( new_n760_, new_n759_, new_n729_ );
and g0589 ( new_n761_, new_n760_, new_n758_ );
or g0590 ( new_n762_, new_n761_, keyIn_0_90 );
and g0591 ( new_n763_, new_n757_, new_n762_ );
and g0592 ( new_n764_, new_n752_, new_n763_ );
not g0593 ( new_n765_, keyIn_0_71 );
or g0594 ( new_n766_, new_n613_, new_n357_ );
not g0595 ( new_n767_, new_n357_ );
or g0596 ( new_n768_, new_n609_, new_n767_ );
and g0597 ( new_n769_, new_n768_, new_n766_ );
and g0598 ( new_n770_, new_n769_, new_n765_ );
and g0599 ( new_n771_, new_n609_, new_n767_ );
and g0600 ( new_n772_, new_n613_, new_n357_ );
or g0601 ( new_n773_, new_n771_, new_n772_ );
and g0602 ( new_n774_, new_n773_, keyIn_0_71 );
not g0603 ( new_n775_, keyIn_0_61 );
not g0604 ( new_n776_, new_n341_ );
not g0605 ( new_n777_, N66 );
and g0606 ( new_n778_, new_n345_, new_n777_ );
and g0607 ( new_n779_, new_n778_, new_n342_ );
and g0608 ( new_n780_, new_n776_, new_n779_ );
not g0609 ( new_n781_, new_n780_ );
and g0610 ( new_n782_, new_n781_, keyIn_0_57 );
not g0611 ( new_n783_, new_n782_ );
or g0612 ( new_n784_, new_n781_, keyIn_0_57 );
and g0613 ( new_n785_, new_n783_, new_n784_ );
not g0614 ( new_n786_, new_n785_ );
and g0615 ( new_n787_, new_n786_, new_n775_ );
and g0616 ( new_n788_, new_n785_, keyIn_0_61 );
or g0617 ( new_n789_, new_n787_, new_n788_ );
not g0618 ( new_n790_, new_n789_ );
or g0619 ( new_n791_, new_n774_, new_n790_ );
or g0620 ( new_n792_, new_n791_, new_n770_ );
or g0621 ( new_n793_, new_n792_, keyIn_0_88 );
not g0622 ( new_n794_, keyIn_0_73 );
not g0623 ( new_n795_, new_n382_ );
and g0624 ( new_n796_, new_n609_, new_n795_ );
and g0625 ( new_n797_, new_n613_, new_n382_ );
or g0626 ( new_n798_, new_n796_, new_n797_ );
and g0627 ( new_n799_, new_n798_, new_n794_ );
or g0628 ( new_n800_, new_n613_, new_n382_ );
or g0629 ( new_n801_, new_n609_, new_n795_ );
and g0630 ( new_n802_, new_n801_, new_n800_ );
and g0631 ( new_n803_, new_n802_, keyIn_0_73 );
or g0632 ( new_n804_, new_n799_, new_n803_ );
not g0633 ( new_n805_, new_n364_ );
not g0634 ( new_n806_, N79 );
and g0635 ( new_n807_, new_n370_, new_n806_ );
and g0636 ( new_n808_, new_n805_, new_n807_ );
not g0637 ( new_n809_, new_n808_ );
and g0638 ( new_n810_, new_n809_, keyIn_0_58 );
not g0639 ( new_n811_, new_n810_ );
or g0640 ( new_n812_, new_n809_, keyIn_0_58 );
and g0641 ( new_n813_, new_n811_, new_n812_ );
not g0642 ( new_n814_, new_n813_ );
and g0643 ( new_n815_, new_n814_, keyIn_0_62 );
not g0644 ( new_n816_, new_n815_ );
or g0645 ( new_n817_, new_n814_, keyIn_0_62 );
and g0646 ( new_n818_, new_n816_, new_n817_ );
not g0647 ( new_n819_, new_n818_ );
and g0648 ( new_n820_, new_n804_, new_n819_ );
or g0649 ( new_n821_, new_n820_, keyIn_0_89 );
and g0650 ( new_n822_, new_n793_, new_n821_ );
not g0651 ( new_n823_, keyIn_0_89 );
or g0652 ( new_n824_, new_n802_, keyIn_0_73 );
or g0653 ( new_n825_, new_n798_, new_n794_ );
and g0654 ( new_n826_, new_n825_, new_n824_ );
or g0655 ( new_n827_, new_n826_, new_n818_ );
or g0656 ( new_n828_, new_n827_, new_n823_ );
not g0657 ( new_n829_, keyIn_0_88 );
not g0658 ( new_n830_, new_n770_ );
or g0659 ( new_n831_, new_n769_, new_n765_ );
and g0660 ( new_n832_, new_n831_, new_n789_ );
and g0661 ( new_n833_, new_n832_, new_n830_ );
or g0662 ( new_n834_, new_n833_, new_n829_ );
and g0663 ( new_n835_, new_n828_, new_n834_ );
and g0664 ( new_n836_, new_n822_, new_n835_ );
and g0665 ( new_n837_, new_n764_, new_n836_ );
and g0666 ( new_n838_, new_n837_, new_n715_ );
and g0667 ( new_n839_, new_n838_, new_n676_ );
not g0668 ( new_n840_, new_n839_ );
and g0669 ( new_n841_, new_n840_, keyIn_0_93 );
not g0670 ( new_n842_, keyIn_0_93 );
and g0671 ( new_n843_, new_n839_, new_n842_ );
or g0672 ( new_n844_, new_n841_, new_n843_ );
or g0673 ( new_n845_, new_n844_, new_n600_ );
or g0674 ( new_n846_, new_n839_, new_n842_ );
not g0675 ( new_n847_, new_n843_ );
and g0676 ( new_n848_, new_n847_, new_n846_ );
or g0677 ( new_n849_, new_n848_, keyIn_0_95 );
and g0678 ( N370, new_n845_, new_n849_ );
not g0679 ( new_n851_, keyIn_0_115 );
not g0680 ( new_n852_, keyIn_0_102 );
and g0681 ( new_n853_, new_n848_, keyIn_0_94 );
not g0682 ( new_n854_, keyIn_0_94 );
and g0683 ( new_n855_, new_n844_, new_n854_ );
or g0684 ( new_n856_, new_n855_, new_n853_ );
or g0685 ( new_n857_, new_n856_, new_n727_ );
and g0686 ( new_n858_, new_n857_, new_n852_ );
or g0687 ( new_n859_, new_n844_, new_n854_ );
or g0688 ( new_n860_, new_n848_, keyIn_0_94 );
and g0689 ( new_n861_, new_n859_, new_n860_ );
and g0690 ( new_n862_, new_n861_, N92 );
and g0691 ( new_n863_, new_n862_, keyIn_0_102 );
or g0692 ( new_n864_, new_n858_, new_n863_ );
and g0693 ( new_n865_, new_n607_, keyIn_0_65 );
not g0694 ( new_n866_, new_n865_ );
or g0695 ( new_n867_, new_n607_, keyIn_0_65 );
and g0696 ( new_n868_, new_n866_, new_n867_ );
and g0697 ( new_n869_, new_n868_, N86 );
and g0698 ( new_n870_, new_n869_, keyIn_0_81 );
not g0699 ( new_n871_, new_n870_ );
or g0700 ( new_n872_, new_n869_, keyIn_0_81 );
and g0701 ( new_n873_, new_n871_, new_n872_ );
and g0702 ( new_n874_, N223, N76 );
or g0703 ( new_n875_, new_n874_, new_n185_ );
or g0704 ( new_n876_, new_n873_, new_n875_ );
not g0705 ( new_n877_, new_n876_ );
and g0706 ( new_n878_, new_n864_, new_n877_ );
and g0707 ( new_n879_, new_n878_, keyIn_0_111 );
not g0708 ( new_n880_, keyIn_0_111 );
or g0709 ( new_n881_, new_n862_, keyIn_0_102 );
or g0710 ( new_n882_, new_n857_, new_n852_ );
and g0711 ( new_n883_, new_n882_, new_n881_ );
or g0712 ( new_n884_, new_n883_, new_n876_ );
and g0713 ( new_n885_, new_n884_, new_n880_ );
or g0714 ( new_n886_, new_n885_, new_n879_ );
not g0715 ( new_n887_, keyIn_0_113 );
not g0716 ( new_n888_, keyIn_0_104 );
and g0717 ( new_n889_, new_n861_, N115 );
and g0718 ( new_n890_, new_n889_, new_n888_ );
not g0719 ( new_n891_, new_n890_ );
or g0720 ( new_n892_, new_n889_, new_n888_ );
and g0721 ( new_n893_, new_n891_, new_n892_ );
and g0722 ( new_n894_, new_n868_, N112 );
and g0723 ( new_n895_, new_n894_, keyIn_0_83 );
not g0724 ( new_n896_, new_n895_ );
or g0725 ( new_n897_, new_n894_, keyIn_0_83 );
and g0726 ( new_n898_, new_n896_, new_n897_ );
and g0727 ( new_n899_, N223, N102 );
or g0728 ( new_n900_, new_n899_, new_n174_ );
or g0729 ( new_n901_, new_n898_, new_n900_ );
or g0730 ( new_n902_, new_n893_, new_n901_ );
not g0731 ( new_n903_, new_n902_ );
or g0732 ( new_n904_, new_n903_, new_n887_ );
or g0733 ( new_n905_, new_n902_, keyIn_0_113 );
and g0734 ( new_n906_, new_n904_, new_n905_ );
and g0735 ( new_n907_, new_n906_, new_n886_ );
not g0736 ( new_n908_, keyIn_0_110 );
and g0737 ( new_n909_, new_n861_, N79 );
and g0738 ( new_n910_, new_n909_, keyIn_0_101 );
not g0739 ( new_n911_, keyIn_0_101 );
or g0740 ( new_n912_, new_n856_, new_n806_ );
and g0741 ( new_n913_, new_n912_, new_n911_ );
not g0742 ( new_n914_, keyIn_0_80 );
and g0743 ( new_n915_, new_n868_, N73 );
and g0744 ( new_n916_, new_n915_, new_n914_ );
not g0745 ( new_n917_, new_n916_ );
or g0746 ( new_n918_, new_n915_, new_n914_ );
and g0747 ( new_n919_, N223, N63 );
or g0748 ( new_n920_, new_n919_, new_n251_ );
not g0749 ( new_n921_, new_n920_ );
and g0750 ( new_n922_, new_n918_, new_n921_ );
and g0751 ( new_n923_, new_n922_, new_n917_ );
not g0752 ( new_n924_, new_n923_ );
or g0753 ( new_n925_, new_n913_, new_n924_ );
or g0754 ( new_n926_, new_n925_, new_n910_ );
or g0755 ( new_n927_, new_n926_, new_n908_ );
not g0756 ( new_n928_, new_n910_ );
or g0757 ( new_n929_, new_n909_, keyIn_0_101 );
and g0758 ( new_n930_, new_n929_, new_n923_ );
and g0759 ( new_n931_, new_n930_, new_n928_ );
or g0760 ( new_n932_, new_n931_, keyIn_0_110 );
and g0761 ( new_n933_, new_n927_, new_n932_ );
and g0762 ( new_n934_, new_n861_, N105 );
and g0763 ( new_n935_, new_n934_, keyIn_0_103 );
not g0764 ( new_n936_, keyIn_0_103 );
or g0765 ( new_n937_, new_n856_, new_n639_ );
and g0766 ( new_n938_, new_n937_, new_n936_ );
and g0767 ( new_n939_, new_n868_, N99 );
not g0768 ( new_n940_, new_n939_ );
and g0769 ( new_n941_, new_n940_, keyIn_0_82 );
not g0770 ( new_n942_, new_n941_ );
or g0771 ( new_n943_, new_n940_, keyIn_0_82 );
and g0772 ( new_n944_, new_n942_, new_n943_ );
and g0773 ( new_n945_, N223, N89 );
or g0774 ( new_n946_, new_n945_, new_n508_ );
or g0775 ( new_n947_, new_n944_, new_n946_ );
or g0776 ( new_n948_, new_n938_, new_n947_ );
or g0777 ( new_n949_, new_n948_, new_n935_ );
or g0778 ( new_n950_, new_n949_, keyIn_0_112 );
not g0779 ( new_n951_, keyIn_0_112 );
not g0780 ( new_n952_, new_n935_ );
or g0781 ( new_n953_, new_n934_, keyIn_0_103 );
not g0782 ( new_n954_, new_n947_ );
and g0783 ( new_n955_, new_n953_, new_n954_ );
and g0784 ( new_n956_, new_n955_, new_n952_ );
or g0785 ( new_n957_, new_n956_, new_n951_ );
and g0786 ( new_n958_, new_n950_, new_n957_ );
and g0787 ( new_n959_, new_n933_, new_n958_ );
and g0788 ( new_n960_, new_n907_, new_n959_ );
not g0789 ( new_n961_, keyIn_0_107 );
or g0790 ( new_n962_, new_n856_, new_n686_ );
or g0791 ( new_n963_, new_n962_, keyIn_0_98 );
not g0792 ( new_n964_, keyIn_0_98 );
and g0793 ( new_n965_, new_n861_, N40 );
or g0794 ( new_n966_, new_n965_, new_n964_ );
and g0795 ( new_n967_, new_n963_, new_n966_ );
and g0796 ( new_n968_, new_n868_, N34 );
and g0797 ( new_n969_, new_n968_, keyIn_0_74 );
not g0798 ( new_n970_, new_n969_ );
or g0799 ( new_n971_, new_n968_, keyIn_0_74 );
and g0800 ( new_n972_, new_n970_, new_n971_ );
and g0801 ( new_n973_, N223, N24 );
or g0802 ( new_n974_, new_n973_, new_n211_ );
or g0803 ( new_n975_, new_n972_, new_n974_ );
or g0804 ( new_n976_, new_n967_, new_n975_ );
and g0805 ( new_n977_, new_n976_, new_n961_ );
and g0806 ( new_n978_, new_n965_, new_n964_ );
and g0807 ( new_n979_, new_n962_, keyIn_0_98 );
or g0808 ( new_n980_, new_n979_, new_n978_ );
not g0809 ( new_n981_, new_n975_ );
and g0810 ( new_n982_, new_n980_, new_n981_ );
and g0811 ( new_n983_, new_n982_, keyIn_0_107 );
or g0812 ( new_n984_, new_n977_, new_n983_ );
not g0813 ( new_n985_, new_n984_ );
and g0814 ( new_n986_, new_n861_, N27 );
and g0815 ( new_n987_, new_n986_, keyIn_0_97 );
not g0816 ( new_n988_, new_n987_ );
or g0817 ( new_n989_, new_n986_, keyIn_0_97 );
not g0818 ( new_n990_, keyIn_0_72 );
and g0819 ( new_n991_, new_n868_, N21 );
and g0820 ( new_n992_, new_n991_, new_n990_ );
not g0821 ( new_n993_, new_n992_ );
or g0822 ( new_n994_, new_n991_, new_n990_ );
and g0823 ( new_n995_, N223, N11 );
and g0824 ( new_n996_, new_n995_, keyIn_0_45 );
not g0825 ( new_n997_, new_n996_ );
or g0826 ( new_n998_, new_n995_, keyIn_0_45 );
and g0827 ( new_n999_, new_n998_, N17 );
and g0828 ( new_n1000_, new_n999_, new_n997_ );
and g0829 ( new_n1001_, new_n994_, new_n1000_ );
and g0830 ( new_n1002_, new_n1001_, new_n993_ );
and g0831 ( new_n1003_, new_n989_, new_n1002_ );
and g0832 ( new_n1004_, new_n1003_, new_n988_ );
not g0833 ( new_n1005_, new_n1004_ );
and g0834 ( new_n1006_, new_n1005_, keyIn_0_106 );
not g0835 ( new_n1007_, keyIn_0_106 );
and g0836 ( new_n1008_, new_n1004_, new_n1007_ );
or g0837 ( new_n1009_, new_n1006_, new_n1008_ );
and g0838 ( new_n1010_, new_n985_, new_n1009_ );
not g0839 ( new_n1011_, keyIn_0_100 );
or g0840 ( new_n1012_, new_n856_, new_n777_ );
or g0841 ( new_n1013_, new_n1012_, new_n1011_ );
and g0842 ( new_n1014_, new_n861_, N66 );
or g0843 ( new_n1015_, new_n1014_, keyIn_0_100 );
and g0844 ( new_n1016_, new_n1013_, new_n1015_ );
not g0845 ( new_n1017_, keyIn_0_78 );
and g0846 ( new_n1018_, new_n868_, N60 );
and g0847 ( new_n1019_, new_n1018_, new_n1017_ );
not g0848 ( new_n1020_, new_n1019_ );
or g0849 ( new_n1021_, new_n1018_, new_n1017_ );
and g0850 ( new_n1022_, new_n1020_, new_n1021_ );
and g0851 ( new_n1023_, N223, N50 );
or g0852 ( new_n1024_, new_n1023_, new_n222_ );
or g0853 ( new_n1025_, new_n1022_, new_n1024_ );
or g0854 ( new_n1026_, new_n1016_, new_n1025_ );
and g0855 ( new_n1027_, new_n1026_, keyIn_0_109 );
not g0856 ( new_n1028_, keyIn_0_109 );
and g0857 ( new_n1029_, new_n1014_, keyIn_0_100 );
and g0858 ( new_n1030_, new_n1012_, new_n1011_ );
or g0859 ( new_n1031_, new_n1030_, new_n1029_ );
not g0860 ( new_n1032_, new_n1025_ );
and g0861 ( new_n1033_, new_n1031_, new_n1032_ );
and g0862 ( new_n1034_, new_n1033_, new_n1028_ );
or g0863 ( new_n1035_, new_n1027_, new_n1034_ );
not g0864 ( new_n1036_, keyIn_0_108 );
or g0865 ( new_n1037_, new_n856_, new_n702_ );
or g0866 ( new_n1038_, new_n1037_, keyIn_0_99 );
not g0867 ( new_n1039_, keyIn_0_99 );
and g0868 ( new_n1040_, new_n861_, N53 );
or g0869 ( new_n1041_, new_n1040_, new_n1039_ );
and g0870 ( new_n1042_, new_n1038_, new_n1041_ );
and g0871 ( new_n1043_, new_n868_, N47 );
and g0872 ( new_n1044_, new_n1043_, keyIn_0_76 );
not g0873 ( new_n1045_, new_n1044_ );
or g0874 ( new_n1046_, new_n1043_, keyIn_0_76 );
and g0875 ( new_n1047_, new_n1045_, new_n1046_ );
and g0876 ( new_n1048_, N223, N37 );
or g0877 ( new_n1049_, new_n1048_, new_n242_ );
or g0878 ( new_n1050_, new_n1047_, new_n1049_ );
or g0879 ( new_n1051_, new_n1042_, new_n1050_ );
and g0880 ( new_n1052_, new_n1051_, new_n1036_ );
and g0881 ( new_n1053_, new_n1040_, new_n1039_ );
and g0882 ( new_n1054_, new_n1037_, keyIn_0_99 );
or g0883 ( new_n1055_, new_n1054_, new_n1053_ );
not g0884 ( new_n1056_, new_n1050_ );
and g0885 ( new_n1057_, new_n1055_, new_n1056_ );
and g0886 ( new_n1058_, new_n1057_, keyIn_0_108 );
or g0887 ( new_n1059_, new_n1052_, new_n1058_ );
and g0888 ( new_n1060_, new_n1035_, new_n1059_ );
and g0889 ( new_n1061_, new_n1010_, new_n1060_ );
and g0890 ( new_n1062_, new_n960_, new_n1061_ );
or g0891 ( new_n1063_, new_n1062_, new_n851_ );
and g0892 ( new_n1064_, new_n1062_, new_n851_ );
not g0893 ( new_n1065_, new_n1064_ );
not g0894 ( new_n1066_, keyIn_0_114 );
not g0895 ( new_n1067_, keyIn_0_96 );
and g0896 ( new_n1068_, new_n861_, N14 );
and g0897 ( new_n1069_, new_n1068_, new_n1067_ );
not g0898 ( new_n1070_, new_n1069_ );
or g0899 ( new_n1071_, new_n1068_, new_n1067_ );
and g0900 ( new_n1072_, new_n1070_, new_n1071_ );
and g0901 ( new_n1073_, new_n868_, N8 );
and g0902 ( new_n1074_, new_n1073_, keyIn_0_70 );
not g0903 ( new_n1075_, new_n1074_ );
or g0904 ( new_n1076_, new_n1073_, keyIn_0_70 );
and g0905 ( new_n1077_, new_n1075_, new_n1076_ );
and g0906 ( new_n1078_, N223, N1 );
or g0907 ( new_n1079_, new_n1078_, new_n263_ );
or g0908 ( new_n1080_, new_n1077_, new_n1079_ );
or g0909 ( new_n1081_, new_n1072_, new_n1080_ );
and g0910 ( new_n1082_, new_n1081_, keyIn_0_105 );
not g0911 ( new_n1083_, new_n1082_ );
or g0912 ( new_n1084_, new_n1081_, keyIn_0_105 );
and g0913 ( new_n1085_, new_n1083_, new_n1084_ );
not g0914 ( new_n1086_, new_n1085_ );
and g0915 ( new_n1087_, new_n1086_, new_n1066_ );
and g0916 ( new_n1088_, new_n1085_, keyIn_0_114 );
or g0917 ( new_n1089_, new_n1087_, new_n1088_ );
and g0918 ( new_n1090_, new_n1065_, new_n1089_ );
and g0919 ( new_n1091_, new_n1090_, new_n1063_ );
or g0920 ( new_n1092_, new_n1091_, keyIn_0_120 );
not g0921 ( new_n1093_, keyIn_0_120 );
not g0922 ( new_n1094_, new_n1091_ );
or g0923 ( new_n1095_, new_n1094_, new_n1093_ );
and g0924 ( N421, new_n1095_, new_n1092_ );
or g0925 ( new_n1097_, new_n1059_, keyIn_0_116 );
not g0926 ( new_n1098_, keyIn_0_116 );
or g0927 ( new_n1099_, new_n1057_, keyIn_0_108 );
or g0928 ( new_n1100_, new_n1051_, new_n1036_ );
and g0929 ( new_n1101_, new_n1100_, new_n1099_ );
or g0930 ( new_n1102_, new_n1101_, new_n1098_ );
and g0931 ( new_n1103_, new_n1097_, new_n1102_ );
or g0932 ( new_n1104_, new_n1103_, new_n984_ );
and g0933 ( new_n1105_, new_n1104_, keyIn_0_121 );
not g0934 ( new_n1106_, keyIn_0_121 );
and g0935 ( new_n1107_, new_n1101_, new_n1098_ );
and g0936 ( new_n1108_, new_n1059_, keyIn_0_116 );
or g0937 ( new_n1109_, new_n1108_, new_n1107_ );
and g0938 ( new_n1110_, new_n1109_, new_n985_ );
and g0939 ( new_n1111_, new_n1110_, new_n1106_ );
or g0940 ( new_n1112_, new_n1105_, new_n1111_ );
and g0941 ( new_n1113_, new_n1010_, new_n1035_ );
and g0942 ( new_n1114_, new_n1112_, new_n1113_ );
not g0943 ( new_n1115_, new_n1114_ );
or g0944 ( new_n1116_, new_n1115_, keyIn_0_125 );
not g0945 ( new_n1117_, keyIn_0_125 );
or g0946 ( new_n1118_, new_n1114_, new_n1117_ );
and g0947 ( N430, new_n1116_, new_n1118_ );
not g0948 ( new_n1120_, keyIn_0_126 );
not g0949 ( new_n1121_, keyIn_0_122 );
or g0950 ( new_n1122_, new_n933_, keyIn_0_117 );
not g0951 ( new_n1123_, keyIn_0_117 );
and g0952 ( new_n1124_, new_n931_, keyIn_0_110 );
and g0953 ( new_n1125_, new_n926_, new_n908_ );
or g0954 ( new_n1126_, new_n1125_, new_n1124_ );
or g0955 ( new_n1127_, new_n1126_, new_n1123_ );
and g0956 ( new_n1128_, new_n1122_, new_n1127_ );
or g0957 ( new_n1129_, new_n1033_, new_n1028_ );
or g0958 ( new_n1130_, new_n1026_, keyIn_0_109 );
and g0959 ( new_n1131_, new_n1130_, new_n1129_ );
or g0960 ( new_n1132_, new_n1131_, new_n1101_ );
or g0961 ( new_n1133_, new_n1132_, new_n984_ );
or g0962 ( new_n1134_, new_n1133_, new_n1128_ );
and g0963 ( new_n1135_, new_n1134_, new_n1121_ );
and g0964 ( new_n1136_, new_n1126_, new_n1123_ );
and g0965 ( new_n1137_, new_n933_, keyIn_0_117 );
or g0966 ( new_n1138_, new_n1136_, new_n1137_ );
and g0967 ( new_n1139_, new_n1060_, new_n985_ );
and g0968 ( new_n1140_, new_n1138_, new_n1139_ );
and g0969 ( new_n1141_, new_n1140_, keyIn_0_122 );
or g0970 ( new_n1142_, new_n1135_, new_n1141_ );
not g0971 ( new_n1143_, new_n1010_ );
or g0972 ( new_n1144_, new_n884_, new_n880_ );
or g0973 ( new_n1145_, new_n878_, keyIn_0_111 );
and g0974 ( new_n1146_, new_n1144_, new_n1145_ );
and g0975 ( new_n1147_, new_n1146_, keyIn_0_118 );
not g0976 ( new_n1148_, keyIn_0_118 );
and g0977 ( new_n1149_, new_n886_, new_n1148_ );
or g0978 ( new_n1150_, new_n1149_, new_n1147_ );
and g0979 ( new_n1151_, new_n1150_, new_n1060_ );
or g0980 ( new_n1152_, new_n1151_, keyIn_0_123 );
not g0981 ( new_n1153_, keyIn_0_123 );
or g0982 ( new_n1154_, new_n886_, new_n1148_ );
or g0983 ( new_n1155_, new_n1146_, keyIn_0_118 );
and g0984 ( new_n1156_, new_n1154_, new_n1155_ );
or g0985 ( new_n1157_, new_n1156_, new_n1132_ );
or g0986 ( new_n1158_, new_n1157_, new_n1153_ );
and g0987 ( new_n1159_, new_n1158_, new_n1152_ );
or g0988 ( new_n1160_, new_n1159_, new_n1143_ );
or g0989 ( new_n1161_, new_n1160_, new_n1142_ );
or g0990 ( new_n1162_, new_n1161_, new_n1120_ );
or g0991 ( new_n1163_, new_n1140_, keyIn_0_122 );
not g0992 ( new_n1164_, new_n1141_ );
and g0993 ( new_n1165_, new_n1164_, new_n1163_ );
and g0994 ( new_n1166_, new_n1157_, new_n1153_ );
and g0995 ( new_n1167_, new_n1151_, keyIn_0_123 );
or g0996 ( new_n1168_, new_n1166_, new_n1167_ );
and g0997 ( new_n1169_, new_n1168_, new_n1010_ );
and g0998 ( new_n1170_, new_n1169_, new_n1165_ );
or g0999 ( new_n1171_, new_n1170_, keyIn_0_126 );
and g1000 ( N431, new_n1162_, new_n1171_ );
not g1001 ( new_n1173_, keyIn_0_124 );
and g1002 ( new_n1174_, new_n985_, new_n886_ );
and g1003 ( new_n1175_, new_n1174_, new_n1059_ );
and g1004 ( new_n1176_, new_n956_, new_n951_ );
and g1005 ( new_n1177_, new_n949_, keyIn_0_112 );
or g1006 ( new_n1178_, new_n1177_, new_n1176_ );
and g1007 ( new_n1179_, new_n1178_, keyIn_0_119 );
not g1008 ( new_n1180_, new_n1179_ );
not g1009 ( new_n1181_, keyIn_0_119 );
and g1010 ( new_n1182_, new_n958_, new_n1181_ );
not g1011 ( new_n1183_, new_n1182_ );
and g1012 ( new_n1184_, new_n1180_, new_n1183_ );
and g1013 ( new_n1185_, new_n1184_, new_n1175_ );
and g1014 ( new_n1186_, new_n1185_, new_n1173_ );
not g1015 ( new_n1187_, new_n1009_ );
or g1016 ( new_n1188_, new_n984_, new_n1146_ );
or g1017 ( new_n1189_, new_n1188_, new_n1101_ );
or g1018 ( new_n1190_, new_n1179_, new_n1182_ );
or g1019 ( new_n1191_, new_n1189_, new_n1190_ );
and g1020 ( new_n1192_, new_n1191_, keyIn_0_124 );
or g1021 ( new_n1193_, new_n1192_, new_n1187_ );
or g1022 ( new_n1194_, new_n1193_, new_n1186_ );
or g1023 ( new_n1195_, new_n1110_, new_n1106_ );
or g1024 ( new_n1196_, new_n1104_, keyIn_0_121 );
and g1025 ( new_n1197_, new_n1196_, new_n1195_ );
or g1026 ( new_n1198_, new_n1142_, new_n1197_ );
or g1027 ( new_n1199_, new_n1194_, new_n1198_ );
and g1028 ( new_n1200_, new_n1199_, keyIn_0_127 );
not g1029 ( new_n1201_, keyIn_0_127 );
not g1030 ( new_n1202_, new_n1186_ );
or g1031 ( new_n1203_, new_n1185_, new_n1173_ );
and g1032 ( new_n1204_, new_n1203_, new_n1009_ );
and g1033 ( new_n1205_, new_n1204_, new_n1202_ );
and g1034 ( new_n1206_, new_n1165_, new_n1112_ );
and g1035 ( new_n1207_, new_n1206_, new_n1205_ );
and g1036 ( new_n1208_, new_n1207_, new_n1201_ );
or g1037 ( N432, new_n1200_, new_n1208_ );
endmodule