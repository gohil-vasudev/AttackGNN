module add_mul_combine_16_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, 
        b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, 
        b_14_, b_15_, Result_mul_0_, Result_mul_1_, Result_mul_2_, 
        Result_mul_3_, Result_mul_4_, Result_mul_5_, Result_mul_6_, 
        Result_mul_7_, Result_mul_8_, Result_mul_9_, Result_mul_10_, 
        Result_mul_11_, Result_mul_12_, Result_mul_13_, Result_mul_14_, 
        Result_mul_15_, Result_mul_16_, Result_mul_17_, Result_mul_18_, 
        Result_mul_19_, Result_mul_20_, Result_mul_21_, Result_mul_22_, 
        Result_mul_23_, Result_mul_24_, Result_mul_25_, Result_mul_26_, 
        Result_mul_27_, Result_mul_28_, Result_mul_29_, Result_mul_30_, 
        Result_mul_31_, Result_add_0_, Result_add_1_, Result_add_2_, 
        Result_add_3_, Result_add_4_, Result_add_5_, Result_add_6_, 
        Result_add_7_, Result_add_8_, Result_add_9_, Result_add_10_, 
        Result_add_11_, Result_add_12_, Result_add_13_, Result_add_14_, 
        Result_add_15_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_,
         b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_;
  output Result_mul_0_, Result_mul_1_, Result_mul_2_, Result_mul_3_,
         Result_mul_4_, Result_mul_5_, Result_mul_6_, Result_mul_7_,
         Result_mul_8_, Result_mul_9_, Result_mul_10_, Result_mul_11_,
         Result_mul_12_, Result_mul_13_, Result_mul_14_, Result_mul_15_,
         Result_mul_16_, Result_mul_17_, Result_mul_18_, Result_mul_19_,
         Result_mul_20_, Result_mul_21_, Result_mul_22_, Result_mul_23_,
         Result_mul_24_, Result_mul_25_, Result_mul_26_, Result_mul_27_,
         Result_mul_28_, Result_mul_29_, Result_mul_30_, Result_mul_31_,
         Result_add_0_, Result_add_1_, Result_add_2_, Result_add_3_,
         Result_add_4_, Result_add_5_, Result_add_6_, Result_add_7_,
         Result_add_8_, Result_add_9_, Result_add_10_, Result_add_11_,
         Result_add_12_, Result_add_13_, Result_add_14_, Result_add_15_;
  wire   n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844;

  XOR2_X1 U1873 ( .A(n1826), .B(n1827), .Z(Result_mul_9_) );
  AND2_X1 U1874 ( .A1(n1828), .A2(n1829), .ZN(n1827) );
  XOR2_X1 U1875 ( .A(n1830), .B(n1831), .Z(Result_mul_8_) );
  AND2_X1 U1876 ( .A1(n1832), .A2(n1833), .ZN(n1831) );
  XOR2_X1 U1877 ( .A(n1834), .B(n1835), .Z(Result_mul_7_) );
  AND2_X1 U1878 ( .A1(n1836), .A2(n1837), .ZN(n1835) );
  XOR2_X1 U1879 ( .A(n1838), .B(n1839), .Z(Result_mul_6_) );
  AND2_X1 U1880 ( .A1(n1840), .A2(n1841), .ZN(n1839) );
  XOR2_X1 U1881 ( .A(n1842), .B(n1843), .Z(Result_mul_5_) );
  AND2_X1 U1882 ( .A1(n1844), .A2(n1845), .ZN(n1843) );
  XOR2_X1 U1883 ( .A(n1846), .B(n1847), .Z(Result_mul_4_) );
  AND2_X1 U1884 ( .A1(n1848), .A2(n1849), .ZN(n1847) );
  XOR2_X1 U1885 ( .A(n1850), .B(n1851), .Z(Result_mul_3_) );
  AND2_X1 U1886 ( .A1(n1852), .A2(n1853), .ZN(n1851) );
  NAND2_X1 U1887 ( .A1(n1854), .A2(n1855), .ZN(Result_mul_30_) );
  NAND2_X1 U1888 ( .A1(b_14_), .A2(n1856), .ZN(n1855) );
  NAND2_X1 U1889 ( .A1(n1857), .A2(n1858), .ZN(n1856) );
  NAND2_X1 U1890 ( .A1(a_15_), .A2(n1859), .ZN(n1858) );
  NAND2_X1 U1891 ( .A1(b_15_), .A2(n1860), .ZN(n1854) );
  NAND2_X1 U1892 ( .A1(n1861), .A2(n1862), .ZN(n1860) );
  NAND2_X1 U1893 ( .A1(a_14_), .A2(n1863), .ZN(n1862) );
  XOR2_X1 U1894 ( .A(n1864), .B(n1865), .Z(Result_mul_2_) );
  AND2_X1 U1895 ( .A1(n1866), .A2(n1867), .ZN(n1865) );
  XOR2_X1 U1896 ( .A(n1868), .B(n1869), .Z(Result_mul_29_) );
  NOR2_X1 U1897 ( .A1(n1870), .A2(n1859), .ZN(n1869) );
  XOR2_X1 U1898 ( .A(n1871), .B(n1872), .Z(n1868) );
  XOR2_X1 U1899 ( .A(n1873), .B(n1874), .Z(Result_mul_28_) );
  XNOR2_X1 U1900 ( .A(n1875), .B(n1876), .ZN(n1874) );
  NAND2_X1 U1901 ( .A1(b_15_), .A2(a_12_), .ZN(n1875) );
  XNOR2_X1 U1902 ( .A(n1877), .B(n1878), .ZN(Result_mul_27_) );
  NAND2_X1 U1903 ( .A1(n1879), .A2(n1880), .ZN(n1877) );
  XOR2_X1 U1904 ( .A(n1881), .B(n1882), .Z(Result_mul_26_) );
  XOR2_X1 U1905 ( .A(n1883), .B(n1884), .Z(n1881) );
  NOR2_X1 U1906 ( .A1(n1885), .A2(n1859), .ZN(n1884) );
  XNOR2_X1 U1907 ( .A(n1886), .B(n1887), .ZN(Result_mul_25_) );
  NAND2_X1 U1908 ( .A1(n1888), .A2(n1889), .ZN(n1886) );
  XNOR2_X1 U1909 ( .A(n1890), .B(n1891), .ZN(Result_mul_24_) );
  XOR2_X1 U1910 ( .A(n1892), .B(n1893), .Z(n1891) );
  NAND2_X1 U1911 ( .A1(b_15_), .A2(a_8_), .ZN(n1893) );
  XNOR2_X1 U1912 ( .A(n1894), .B(n1895), .ZN(Result_mul_23_) );
  NAND2_X1 U1913 ( .A1(n1896), .A2(n1897), .ZN(n1894) );
  XNOR2_X1 U1914 ( .A(n1898), .B(n1899), .ZN(Result_mul_22_) );
  XOR2_X1 U1915 ( .A(n1900), .B(n1901), .Z(n1899) );
  NAND2_X1 U1916 ( .A1(b_15_), .A2(a_6_), .ZN(n1901) );
  XNOR2_X1 U1917 ( .A(n1902), .B(n1903), .ZN(Result_mul_21_) );
  XOR2_X1 U1918 ( .A(n1904), .B(n1905), .Z(n1903) );
  NAND2_X1 U1919 ( .A1(b_15_), .A2(a_5_), .ZN(n1905) );
  XNOR2_X1 U1920 ( .A(n1906), .B(n1907), .ZN(Result_mul_20_) );
  XOR2_X1 U1921 ( .A(n1908), .B(n1909), .Z(n1907) );
  NAND2_X1 U1922 ( .A1(b_15_), .A2(a_4_), .ZN(n1909) );
  XOR2_X1 U1923 ( .A(n1910), .B(n1911), .Z(Result_mul_1_) );
  NOR2_X1 U1924 ( .A1(n1912), .A2(n1913), .ZN(n1911) );
  INV_X1 U1925 ( .A(n1914), .ZN(n1912) );
  XOR2_X1 U1926 ( .A(n1915), .B(n1916), .Z(Result_mul_19_) );
  XOR2_X1 U1927 ( .A(n1917), .B(n1918), .Z(n1915) );
  NOR2_X1 U1928 ( .A1(n1919), .A2(n1859), .ZN(n1918) );
  INV_X1 U1929 ( .A(b_15_), .ZN(n1859) );
  XNOR2_X1 U1930 ( .A(n1920), .B(n1921), .ZN(Result_mul_18_) );
  XOR2_X1 U1931 ( .A(n1922), .B(n1923), .Z(n1921) );
  NAND2_X1 U1932 ( .A1(b_15_), .A2(a_2_), .ZN(n1923) );
  XNOR2_X1 U1933 ( .A(n1924), .B(n1925), .ZN(Result_mul_17_) );
  XOR2_X1 U1934 ( .A(n1926), .B(n1927), .Z(n1925) );
  NAND2_X1 U1935 ( .A1(b_15_), .A2(a_1_), .ZN(n1927) );
  XNOR2_X1 U1936 ( .A(n1928), .B(n1929), .ZN(Result_mul_16_) );
  XOR2_X1 U1937 ( .A(n1930), .B(n1931), .Z(n1929) );
  NAND2_X1 U1938 ( .A1(b_15_), .A2(a_0_), .ZN(n1931) );
  XOR2_X1 U1939 ( .A(n1932), .B(n1933), .Z(Result_mul_15_) );
  NOR2_X1 U1940 ( .A1(n1934), .A2(n1935), .ZN(Result_mul_14_) );
  NOR2_X1 U1941 ( .A1(n1936), .A2(n1937), .ZN(n1935) );
  AND2_X1 U1942 ( .A1(n1932), .A2(n1933), .ZN(n1936) );
  XNOR2_X1 U1943 ( .A(n1934), .B(n1938), .ZN(Result_mul_13_) );
  NAND2_X1 U1944 ( .A1(n1939), .A2(n1940), .ZN(n1938) );
  NAND2_X1 U1945 ( .A1(n1941), .A2(n1942), .ZN(n1940) );
  INV_X1 U1946 ( .A(n1943), .ZN(n1942) );
  NAND2_X1 U1947 ( .A1(n1944), .A2(n1945), .ZN(n1941) );
  XOR2_X1 U1948 ( .A(n1946), .B(n1947), .Z(Result_mul_12_) );
  XNOR2_X1 U1949 ( .A(n1948), .B(n1949), .ZN(Result_mul_11_) );
  NAND2_X1 U1950 ( .A1(n1950), .A2(n1951), .ZN(n1949) );
  XNOR2_X1 U1951 ( .A(n1952), .B(n1953), .ZN(Result_mul_10_) );
  NAND2_X1 U1952 ( .A1(n1954), .A2(n1955), .ZN(n1952) );
  NAND2_X1 U1953 ( .A1(n1956), .A2(n1957), .ZN(Result_mul_0_) );
  NAND2_X1 U1954 ( .A1(n1914), .A2(n1910), .ZN(n1957) );
  NAND2_X1 U1955 ( .A1(n1867), .A2(n1958), .ZN(n1910) );
  NAND2_X1 U1956 ( .A1(n1866), .A2(n1864), .ZN(n1958) );
  NAND2_X1 U1957 ( .A1(n1853), .A2(n1959), .ZN(n1864) );
  NAND2_X1 U1958 ( .A1(n1852), .A2(n1850), .ZN(n1959) );
  NAND2_X1 U1959 ( .A1(n1849), .A2(n1960), .ZN(n1850) );
  NAND2_X1 U1960 ( .A1(n1848), .A2(n1846), .ZN(n1960) );
  NAND2_X1 U1961 ( .A1(n1845), .A2(n1961), .ZN(n1846) );
  NAND2_X1 U1962 ( .A1(n1844), .A2(n1842), .ZN(n1961) );
  NAND2_X1 U1963 ( .A1(n1841), .A2(n1962), .ZN(n1842) );
  NAND2_X1 U1964 ( .A1(n1840), .A2(n1838), .ZN(n1962) );
  NAND2_X1 U1965 ( .A1(n1837), .A2(n1963), .ZN(n1838) );
  NAND2_X1 U1966 ( .A1(n1836), .A2(n1834), .ZN(n1963) );
  NAND2_X1 U1967 ( .A1(n1833), .A2(n1964), .ZN(n1834) );
  NAND2_X1 U1968 ( .A1(n1832), .A2(n1830), .ZN(n1964) );
  NAND2_X1 U1969 ( .A1(n1829), .A2(n1965), .ZN(n1830) );
  NAND2_X1 U1970 ( .A1(n1828), .A2(n1826), .ZN(n1965) );
  NAND2_X1 U1971 ( .A1(n1954), .A2(n1966), .ZN(n1826) );
  NAND2_X1 U1972 ( .A1(n1953), .A2(n1955), .ZN(n1966) );
  NAND2_X1 U1973 ( .A1(n1967), .A2(n1968), .ZN(n1955) );
  XNOR2_X1 U1974 ( .A(n1969), .B(n1970), .ZN(n1967) );
  NAND2_X1 U1975 ( .A1(n1950), .A2(n1971), .ZN(n1953) );
  NAND2_X1 U1976 ( .A1(n1948), .A2(n1951), .ZN(n1971) );
  NAND2_X1 U1977 ( .A1(n1972), .A2(n1973), .ZN(n1951) );
  NAND2_X1 U1978 ( .A1(n1974), .A2(n1968), .ZN(n1973) );
  NAND2_X1 U1979 ( .A1(n1975), .A2(n1976), .ZN(n1974) );
  NAND2_X1 U1980 ( .A1(n1977), .A2(n1978), .ZN(n1972) );
  AND2_X1 U1981 ( .A1(n1947), .A2(n1946), .ZN(n1948) );
  NAND2_X1 U1982 ( .A1(n1979), .A2(n1980), .ZN(n1946) );
  NAND2_X1 U1983 ( .A1(n1934), .A2(n1943), .ZN(n1980) );
  AND2_X1 U1984 ( .A1(n1981), .A2(n1933), .ZN(n1934) );
  XOR2_X1 U1985 ( .A(n1982), .B(n1983), .Z(n1933) );
  XOR2_X1 U1986 ( .A(n1984), .B(n1985), .Z(n1982) );
  NOR2_X1 U1987 ( .A1(n1986), .A2(n1863), .ZN(n1985) );
  AND2_X1 U1988 ( .A1(n1932), .A2(n1937), .ZN(n1981) );
  XOR2_X1 U1989 ( .A(n1945), .B(n1944), .Z(n1937) );
  NAND2_X1 U1990 ( .A1(n1987), .A2(n1988), .ZN(n1932) );
  NAND2_X1 U1991 ( .A1(n1989), .A2(b_15_), .ZN(n1988) );
  NOR2_X1 U1992 ( .A1(n1990), .A2(n1986), .ZN(n1989) );
  NOR2_X1 U1993 ( .A1(n1928), .A2(n1930), .ZN(n1990) );
  NAND2_X1 U1994 ( .A1(n1928), .A2(n1930), .ZN(n1987) );
  NAND2_X1 U1995 ( .A1(n1991), .A2(n1992), .ZN(n1930) );
  NAND2_X1 U1996 ( .A1(n1993), .A2(b_15_), .ZN(n1992) );
  NOR2_X1 U1997 ( .A1(n1994), .A2(n1995), .ZN(n1993) );
  NOR2_X1 U1998 ( .A1(n1924), .A2(n1926), .ZN(n1994) );
  NAND2_X1 U1999 ( .A1(n1924), .A2(n1926), .ZN(n1991) );
  NAND2_X1 U2000 ( .A1(n1996), .A2(n1997), .ZN(n1926) );
  NAND2_X1 U2001 ( .A1(n1998), .A2(b_15_), .ZN(n1997) );
  NOR2_X1 U2002 ( .A1(n1999), .A2(n2000), .ZN(n1998) );
  NOR2_X1 U2003 ( .A1(n1920), .A2(n1922), .ZN(n1999) );
  NAND2_X1 U2004 ( .A1(n1920), .A2(n1922), .ZN(n1996) );
  NAND2_X1 U2005 ( .A1(n2001), .A2(n2002), .ZN(n1922) );
  NAND2_X1 U2006 ( .A1(n2003), .A2(b_15_), .ZN(n2002) );
  NOR2_X1 U2007 ( .A1(n2004), .A2(n1919), .ZN(n2003) );
  NOR2_X1 U2008 ( .A1(n1916), .A2(n1917), .ZN(n2004) );
  NAND2_X1 U2009 ( .A1(n1916), .A2(n1917), .ZN(n2001) );
  NAND2_X1 U2010 ( .A1(n2005), .A2(n2006), .ZN(n1917) );
  NAND2_X1 U2011 ( .A1(n2007), .A2(b_15_), .ZN(n2006) );
  NOR2_X1 U2012 ( .A1(n2008), .A2(n2009), .ZN(n2007) );
  NOR2_X1 U2013 ( .A1(n1906), .A2(n1908), .ZN(n2008) );
  NAND2_X1 U2014 ( .A1(n1906), .A2(n1908), .ZN(n2005) );
  NAND2_X1 U2015 ( .A1(n2010), .A2(n2011), .ZN(n1908) );
  NAND2_X1 U2016 ( .A1(n2012), .A2(b_15_), .ZN(n2011) );
  NOR2_X1 U2017 ( .A1(n2013), .A2(n2014), .ZN(n2012) );
  NOR2_X1 U2018 ( .A1(n1902), .A2(n1904), .ZN(n2013) );
  NAND2_X1 U2019 ( .A1(n1902), .A2(n1904), .ZN(n2010) );
  NAND2_X1 U2020 ( .A1(n2015), .A2(n2016), .ZN(n1904) );
  NAND2_X1 U2021 ( .A1(n2017), .A2(b_15_), .ZN(n2016) );
  NOR2_X1 U2022 ( .A1(n2018), .A2(n2019), .ZN(n2017) );
  NOR2_X1 U2023 ( .A1(n1898), .A2(n1900), .ZN(n2018) );
  NAND2_X1 U2024 ( .A1(n1898), .A2(n1900), .ZN(n2015) );
  NAND2_X1 U2025 ( .A1(n1896), .A2(n2020), .ZN(n1900) );
  NAND2_X1 U2026 ( .A1(n1895), .A2(n1897), .ZN(n2020) );
  NAND2_X1 U2027 ( .A1(n2021), .A2(n2022), .ZN(n1897) );
  NAND2_X1 U2028 ( .A1(b_15_), .A2(a_7_), .ZN(n2022) );
  INV_X1 U2029 ( .A(n2023), .ZN(n2021) );
  XOR2_X1 U2030 ( .A(n2024), .B(n2025), .Z(n1895) );
  XOR2_X1 U2031 ( .A(n2026), .B(n2027), .Z(n2024) );
  NOR2_X1 U2032 ( .A1(n2028), .A2(n1863), .ZN(n2027) );
  NAND2_X1 U2033 ( .A1(a_7_), .A2(n2023), .ZN(n1896) );
  NAND2_X1 U2034 ( .A1(n2029), .A2(n2030), .ZN(n2023) );
  NAND2_X1 U2035 ( .A1(n2031), .A2(b_15_), .ZN(n2030) );
  NOR2_X1 U2036 ( .A1(n2032), .A2(n2028), .ZN(n2031) );
  NOR2_X1 U2037 ( .A1(n1890), .A2(n1892), .ZN(n2032) );
  NAND2_X1 U2038 ( .A1(n1890), .A2(n1892), .ZN(n2029) );
  NAND2_X1 U2039 ( .A1(n1888), .A2(n2033), .ZN(n1892) );
  NAND2_X1 U2040 ( .A1(n1887), .A2(n1889), .ZN(n2033) );
  NAND2_X1 U2041 ( .A1(n2034), .A2(n2035), .ZN(n1889) );
  NAND2_X1 U2042 ( .A1(b_15_), .A2(a_9_), .ZN(n2035) );
  INV_X1 U2043 ( .A(n2036), .ZN(n2034) );
  XNOR2_X1 U2044 ( .A(n2037), .B(n2038), .ZN(n1887) );
  NAND2_X1 U2045 ( .A1(n2039), .A2(n2040), .ZN(n2037) );
  NAND2_X1 U2046 ( .A1(a_9_), .A2(n2036), .ZN(n1888) );
  NAND2_X1 U2047 ( .A1(n2041), .A2(n2042), .ZN(n2036) );
  NAND2_X1 U2048 ( .A1(n2043), .A2(b_15_), .ZN(n2042) );
  NOR2_X1 U2049 ( .A1(n2044), .A2(n1885), .ZN(n2043) );
  NOR2_X1 U2050 ( .A1(n1882), .A2(n1883), .ZN(n2044) );
  NAND2_X1 U2051 ( .A1(n1882), .A2(n1883), .ZN(n2041) );
  NAND2_X1 U2052 ( .A1(n1879), .A2(n2045), .ZN(n1883) );
  NAND2_X1 U2053 ( .A1(n1878), .A2(n1880), .ZN(n2045) );
  NAND2_X1 U2054 ( .A1(n2046), .A2(n2047), .ZN(n1880) );
  NAND2_X1 U2055 ( .A1(b_15_), .A2(a_11_), .ZN(n2047) );
  INV_X1 U2056 ( .A(n2048), .ZN(n2046) );
  XNOR2_X1 U2057 ( .A(n2049), .B(n2050), .ZN(n1878) );
  XOR2_X1 U2058 ( .A(n2051), .B(n2052), .Z(n2050) );
  NAND2_X1 U2059 ( .A1(b_14_), .A2(a_12_), .ZN(n2052) );
  NAND2_X1 U2060 ( .A1(a_11_), .A2(n2048), .ZN(n1879) );
  NAND2_X1 U2061 ( .A1(n2053), .A2(n2054), .ZN(n2048) );
  NAND2_X1 U2062 ( .A1(n2055), .A2(b_15_), .ZN(n2054) );
  NOR2_X1 U2063 ( .A1(n2056), .A2(n2057), .ZN(n2055) );
  NOR2_X1 U2064 ( .A1(n1873), .A2(n1876), .ZN(n2056) );
  NAND2_X1 U2065 ( .A1(n1873), .A2(n1876), .ZN(n2053) );
  NAND2_X1 U2066 ( .A1(n2058), .A2(n2059), .ZN(n1876) );
  NAND2_X1 U2067 ( .A1(n2060), .A2(b_15_), .ZN(n2059) );
  NOR2_X1 U2068 ( .A1(n2061), .A2(n1870), .ZN(n2060) );
  NOR2_X1 U2069 ( .A1(n1871), .A2(n1872), .ZN(n2061) );
  NAND2_X1 U2070 ( .A1(n1871), .A2(n1872), .ZN(n2058) );
  NAND2_X1 U2071 ( .A1(n2062), .A2(n2063), .ZN(n1872) );
  NAND2_X1 U2072 ( .A1(n2064), .A2(b_14_), .ZN(n2063) );
  NOR2_X1 U2073 ( .A1(n2065), .A2(n2066), .ZN(n2062) );
  NOR2_X1 U2074 ( .A1(n2067), .A2(n2068), .ZN(n2066) );
  NOR2_X1 U2075 ( .A1(n2069), .A2(n2070), .ZN(n2067) );
  NOR2_X1 U2076 ( .A1(b_14_), .A2(n2071), .ZN(n2069) );
  NOR2_X1 U2077 ( .A1(b_13_), .A2(n2072), .ZN(n2065) );
  XOR2_X1 U2078 ( .A(n2073), .B(n2074), .Z(n1873) );
  XOR2_X1 U2079 ( .A(n2075), .B(n2076), .Z(n2073) );
  XNOR2_X1 U2080 ( .A(n2077), .B(n2078), .ZN(n1882) );
  NAND2_X1 U2081 ( .A1(n2079), .A2(n2080), .ZN(n2077) );
  XNOR2_X1 U2082 ( .A(n2081), .B(n2082), .ZN(n1890) );
  XNOR2_X1 U2083 ( .A(n2083), .B(n2084), .ZN(n2082) );
  XOR2_X1 U2084 ( .A(n2085), .B(n2086), .Z(n1898) );
  XOR2_X1 U2085 ( .A(n2087), .B(n2088), .Z(n2085) );
  XOR2_X1 U2086 ( .A(n2089), .B(n2090), .Z(n1902) );
  XOR2_X1 U2087 ( .A(n2091), .B(n2092), .Z(n2089) );
  NOR2_X1 U2088 ( .A1(n2019), .A2(n1863), .ZN(n2092) );
  XOR2_X1 U2089 ( .A(n2093), .B(n2094), .Z(n1906) );
  XOR2_X1 U2090 ( .A(n2095), .B(n2096), .Z(n2093) );
  XOR2_X1 U2091 ( .A(n2097), .B(n2098), .Z(n1916) );
  XOR2_X1 U2092 ( .A(n2099), .B(n2100), .Z(n2097) );
  NOR2_X1 U2093 ( .A1(n2009), .A2(n1863), .ZN(n2100) );
  XNOR2_X1 U2094 ( .A(n2101), .B(n2102), .ZN(n1920) );
  XNOR2_X1 U2095 ( .A(n2103), .B(n2104), .ZN(n2102) );
  XOR2_X1 U2096 ( .A(n2105), .B(n2106), .Z(n1924) );
  XOR2_X1 U2097 ( .A(n2107), .B(n2108), .Z(n2105) );
  NOR2_X1 U2098 ( .A1(n2000), .A2(n1863), .ZN(n2108) );
  XOR2_X1 U2099 ( .A(n2109), .B(n2110), .Z(n1928) );
  XOR2_X1 U2100 ( .A(n2111), .B(n2112), .Z(n2109) );
  NOR2_X1 U2101 ( .A1(n1995), .A2(n1863), .ZN(n2112) );
  NOR2_X1 U2102 ( .A1(n2113), .A2(n2114), .ZN(n1979) );
  INV_X1 U2103 ( .A(n1939), .ZN(n2113) );
  NAND2_X1 U2104 ( .A1(n2115), .A2(n1943), .ZN(n1939) );
  NOR2_X1 U2105 ( .A1(n2114), .A2(n2116), .ZN(n1943) );
  AND2_X1 U2106 ( .A1(n2117), .A2(n2118), .ZN(n2116) );
  NOR2_X1 U2107 ( .A1(n2118), .A2(n2117), .ZN(n2114) );
  XNOR2_X1 U2108 ( .A(n2119), .B(n2120), .ZN(n2117) );
  XOR2_X1 U2109 ( .A(n2121), .B(n2122), .Z(n2119) );
  NOR2_X1 U2110 ( .A1(n1986), .A2(n2123), .ZN(n2122) );
  NAND2_X1 U2111 ( .A1(n2124), .A2(n2125), .ZN(n2118) );
  NAND2_X1 U2112 ( .A1(n2126), .A2(n2127), .ZN(n2125) );
  NAND2_X1 U2113 ( .A1(n2128), .A2(n2129), .ZN(n2127) );
  OR2_X1 U2114 ( .A1(n2129), .A2(n2128), .ZN(n2124) );
  AND2_X1 U2115 ( .A1(n1945), .A2(n1944), .ZN(n2115) );
  XNOR2_X1 U2116 ( .A(n2130), .B(n2126), .ZN(n1944) );
  XOR2_X1 U2117 ( .A(n2131), .B(n2132), .Z(n2126) );
  XNOR2_X1 U2118 ( .A(n2133), .B(n2134), .ZN(n2131) );
  XOR2_X1 U2119 ( .A(n2129), .B(n2128), .Z(n2130) );
  NOR2_X1 U2120 ( .A1(n2068), .A2(n1986), .ZN(n2128) );
  NAND2_X1 U2121 ( .A1(n2135), .A2(n2136), .ZN(n2129) );
  NAND2_X1 U2122 ( .A1(n2137), .A2(b_13_), .ZN(n2136) );
  NOR2_X1 U2123 ( .A1(n2138), .A2(n1995), .ZN(n2137) );
  NOR2_X1 U2124 ( .A1(n2139), .A2(n2140), .ZN(n2138) );
  NAND2_X1 U2125 ( .A1(n2139), .A2(n2140), .ZN(n2135) );
  NAND2_X1 U2126 ( .A1(n2141), .A2(n2142), .ZN(n1945) );
  NAND2_X1 U2127 ( .A1(n2143), .A2(b_14_), .ZN(n2142) );
  NOR2_X1 U2128 ( .A1(n2144), .A2(n1986), .ZN(n2143) );
  NOR2_X1 U2129 ( .A1(n1983), .A2(n1984), .ZN(n2144) );
  NAND2_X1 U2130 ( .A1(n1983), .A2(n1984), .ZN(n2141) );
  NAND2_X1 U2131 ( .A1(n2145), .A2(n2146), .ZN(n1984) );
  NAND2_X1 U2132 ( .A1(n2147), .A2(b_14_), .ZN(n2146) );
  NOR2_X1 U2133 ( .A1(n2148), .A2(n1995), .ZN(n2147) );
  NOR2_X1 U2134 ( .A1(n2110), .A2(n2111), .ZN(n2148) );
  NAND2_X1 U2135 ( .A1(n2110), .A2(n2111), .ZN(n2145) );
  NAND2_X1 U2136 ( .A1(n2149), .A2(n2150), .ZN(n2111) );
  NAND2_X1 U2137 ( .A1(n2151), .A2(b_14_), .ZN(n2150) );
  NOR2_X1 U2138 ( .A1(n2152), .A2(n2000), .ZN(n2151) );
  NOR2_X1 U2139 ( .A1(n2106), .A2(n2107), .ZN(n2152) );
  NAND2_X1 U2140 ( .A1(n2106), .A2(n2107), .ZN(n2149) );
  NAND2_X1 U2141 ( .A1(n2153), .A2(n2154), .ZN(n2107) );
  NAND2_X1 U2142 ( .A1(n2104), .A2(n2155), .ZN(n2154) );
  OR2_X1 U2143 ( .A1(n2103), .A2(n2101), .ZN(n2155) );
  NOR2_X1 U2144 ( .A1(n1863), .A2(n1919), .ZN(n2104) );
  NAND2_X1 U2145 ( .A1(n2101), .A2(n2103), .ZN(n2153) );
  NAND2_X1 U2146 ( .A1(n2156), .A2(n2157), .ZN(n2103) );
  NAND2_X1 U2147 ( .A1(n2158), .A2(b_14_), .ZN(n2157) );
  NOR2_X1 U2148 ( .A1(n2159), .A2(n2009), .ZN(n2158) );
  NOR2_X1 U2149 ( .A1(n2098), .A2(n2099), .ZN(n2159) );
  NAND2_X1 U2150 ( .A1(n2098), .A2(n2099), .ZN(n2156) );
  NAND2_X1 U2151 ( .A1(n2160), .A2(n2161), .ZN(n2099) );
  NAND2_X1 U2152 ( .A1(n2096), .A2(n2162), .ZN(n2161) );
  OR2_X1 U2153 ( .A1(n2095), .A2(n2094), .ZN(n2162) );
  NOR2_X1 U2154 ( .A1(n1863), .A2(n2014), .ZN(n2096) );
  NAND2_X1 U2155 ( .A1(n2094), .A2(n2095), .ZN(n2160) );
  NAND2_X1 U2156 ( .A1(n2163), .A2(n2164), .ZN(n2095) );
  NAND2_X1 U2157 ( .A1(n2165), .A2(b_14_), .ZN(n2164) );
  NOR2_X1 U2158 ( .A1(n2166), .A2(n2019), .ZN(n2165) );
  NOR2_X1 U2159 ( .A1(n2090), .A2(n2091), .ZN(n2166) );
  NAND2_X1 U2160 ( .A1(n2090), .A2(n2091), .ZN(n2163) );
  NAND2_X1 U2161 ( .A1(n2167), .A2(n2168), .ZN(n2091) );
  NAND2_X1 U2162 ( .A1(n2088), .A2(n2169), .ZN(n2168) );
  OR2_X1 U2163 ( .A1(n2087), .A2(n2086), .ZN(n2169) );
  NOR2_X1 U2164 ( .A1(n1863), .A2(n2170), .ZN(n2088) );
  NAND2_X1 U2165 ( .A1(n2086), .A2(n2087), .ZN(n2167) );
  NAND2_X1 U2166 ( .A1(n2171), .A2(n2172), .ZN(n2087) );
  NAND2_X1 U2167 ( .A1(n2173), .A2(b_14_), .ZN(n2172) );
  NOR2_X1 U2168 ( .A1(n2174), .A2(n2028), .ZN(n2173) );
  NOR2_X1 U2169 ( .A1(n2025), .A2(n2026), .ZN(n2174) );
  NAND2_X1 U2170 ( .A1(n2025), .A2(n2026), .ZN(n2171) );
  NAND2_X1 U2171 ( .A1(n2175), .A2(n2176), .ZN(n2026) );
  NAND2_X1 U2172 ( .A1(n2084), .A2(n2177), .ZN(n2176) );
  OR2_X1 U2173 ( .A1(n2083), .A2(n2081), .ZN(n2177) );
  NOR2_X1 U2174 ( .A1(n1863), .A2(n2178), .ZN(n2084) );
  NAND2_X1 U2175 ( .A1(n2081), .A2(n2083), .ZN(n2175) );
  NAND2_X1 U2176 ( .A1(n2039), .A2(n2179), .ZN(n2083) );
  NAND2_X1 U2177 ( .A1(n2038), .A2(n2040), .ZN(n2179) );
  NAND2_X1 U2178 ( .A1(n2180), .A2(n2181), .ZN(n2040) );
  NAND2_X1 U2179 ( .A1(b_14_), .A2(a_10_), .ZN(n2181) );
  INV_X1 U2180 ( .A(n2182), .ZN(n2180) );
  XNOR2_X1 U2181 ( .A(n2183), .B(n2184), .ZN(n2038) );
  NAND2_X1 U2182 ( .A1(n2185), .A2(n2186), .ZN(n2183) );
  NAND2_X1 U2183 ( .A1(a_10_), .A2(n2182), .ZN(n2039) );
  NAND2_X1 U2184 ( .A1(n2079), .A2(n2187), .ZN(n2182) );
  NAND2_X1 U2185 ( .A1(n2078), .A2(n2080), .ZN(n2187) );
  NAND2_X1 U2186 ( .A1(n2188), .A2(n2189), .ZN(n2080) );
  NAND2_X1 U2187 ( .A1(b_14_), .A2(a_11_), .ZN(n2189) );
  INV_X1 U2188 ( .A(n2190), .ZN(n2188) );
  XNOR2_X1 U2189 ( .A(n2191), .B(n2192), .ZN(n2078) );
  XOR2_X1 U2190 ( .A(n2193), .B(n2194), .Z(n2192) );
  NAND2_X1 U2191 ( .A1(b_13_), .A2(a_12_), .ZN(n2194) );
  NAND2_X1 U2192 ( .A1(a_11_), .A2(n2190), .ZN(n2079) );
  NAND2_X1 U2193 ( .A1(n2195), .A2(n2196), .ZN(n2190) );
  NAND2_X1 U2194 ( .A1(n2197), .A2(b_14_), .ZN(n2196) );
  NOR2_X1 U2195 ( .A1(n2198), .A2(n2057), .ZN(n2197) );
  NOR2_X1 U2196 ( .A1(n2049), .A2(n2051), .ZN(n2198) );
  NAND2_X1 U2197 ( .A1(n2049), .A2(n2051), .ZN(n2195) );
  NAND2_X1 U2198 ( .A1(n2199), .A2(n2200), .ZN(n2051) );
  NAND2_X1 U2199 ( .A1(n2074), .A2(n2201), .ZN(n2200) );
  NAND2_X1 U2200 ( .A1(n2076), .A2(n2075), .ZN(n2201) );
  NOR2_X1 U2201 ( .A1(n1863), .A2(n1870), .ZN(n2074) );
  OR2_X1 U2202 ( .A1(n2075), .A2(n2076), .ZN(n2199) );
  AND2_X1 U2203 ( .A1(n2202), .A2(n2203), .ZN(n2076) );
  NAND2_X1 U2204 ( .A1(n2204), .A2(b_12_), .ZN(n2203) );
  NOR2_X1 U2205 ( .A1(n2205), .A2(n2071), .ZN(n2204) );
  NOR2_X1 U2206 ( .A1(n2070), .A2(n2068), .ZN(n2205) );
  NAND2_X1 U2207 ( .A1(n2206), .A2(b_13_), .ZN(n2202) );
  NOR2_X1 U2208 ( .A1(n2207), .A2(n2208), .ZN(n2206) );
  NOR2_X1 U2209 ( .A1(n2064), .A2(n2123), .ZN(n2207) );
  NAND2_X1 U2210 ( .A1(n2209), .A2(b_14_), .ZN(n2075) );
  NOR2_X1 U2211 ( .A1(n2210), .A2(n2068), .ZN(n2209) );
  XOR2_X1 U2212 ( .A(n2211), .B(n2212), .Z(n2049) );
  XOR2_X1 U2213 ( .A(n2213), .B(n2214), .Z(n2211) );
  XNOR2_X1 U2214 ( .A(n2215), .B(n2216), .ZN(n2081) );
  NAND2_X1 U2215 ( .A1(n2217), .A2(n2218), .ZN(n2215) );
  XNOR2_X1 U2216 ( .A(n2219), .B(n2220), .ZN(n2025) );
  XNOR2_X1 U2217 ( .A(n2221), .B(n2222), .ZN(n2219) );
  XNOR2_X1 U2218 ( .A(n2223), .B(n2224), .ZN(n2086) );
  XOR2_X1 U2219 ( .A(n2225), .B(n2226), .Z(n2224) );
  NAND2_X1 U2220 ( .A1(b_13_), .A2(a_8_), .ZN(n2226) );
  XNOR2_X1 U2221 ( .A(n2227), .B(n2228), .ZN(n2090) );
  XNOR2_X1 U2222 ( .A(n2229), .B(n2230), .ZN(n2227) );
  XNOR2_X1 U2223 ( .A(n2231), .B(n2232), .ZN(n2094) );
  XOR2_X1 U2224 ( .A(n2233), .B(n2234), .Z(n2232) );
  NAND2_X1 U2225 ( .A1(b_13_), .A2(a_6_), .ZN(n2234) );
  XNOR2_X1 U2226 ( .A(n2235), .B(n2236), .ZN(n2098) );
  XNOR2_X1 U2227 ( .A(n2237), .B(n2238), .ZN(n2236) );
  XNOR2_X1 U2228 ( .A(n2239), .B(n2240), .ZN(n2101) );
  XOR2_X1 U2229 ( .A(n2241), .B(n2242), .Z(n2240) );
  NAND2_X1 U2230 ( .A1(b_13_), .A2(a_4_), .ZN(n2242) );
  XNOR2_X1 U2231 ( .A(n2243), .B(n2244), .ZN(n2106) );
  XNOR2_X1 U2232 ( .A(n2245), .B(n2246), .ZN(n2244) );
  XOR2_X1 U2233 ( .A(n2247), .B(n2248), .Z(n2110) );
  XOR2_X1 U2234 ( .A(n2249), .B(n2250), .Z(n2247) );
  NOR2_X1 U2235 ( .A1(n2000), .A2(n2068), .ZN(n2250) );
  XNOR2_X1 U2236 ( .A(n2139), .B(n2251), .ZN(n1983) );
  XOR2_X1 U2237 ( .A(n2140), .B(n2252), .Z(n2251) );
  NAND2_X1 U2238 ( .A1(b_13_), .A2(a_1_), .ZN(n2252) );
  NAND2_X1 U2239 ( .A1(n2253), .A2(n2254), .ZN(n2140) );
  NAND2_X1 U2240 ( .A1(n2255), .A2(b_13_), .ZN(n2254) );
  NOR2_X1 U2241 ( .A1(n2256), .A2(n2000), .ZN(n2255) );
  NOR2_X1 U2242 ( .A1(n2248), .A2(n2249), .ZN(n2256) );
  NAND2_X1 U2243 ( .A1(n2248), .A2(n2249), .ZN(n2253) );
  NAND2_X1 U2244 ( .A1(n2257), .A2(n2258), .ZN(n2249) );
  NAND2_X1 U2245 ( .A1(n2246), .A2(n2259), .ZN(n2258) );
  OR2_X1 U2246 ( .A1(n2245), .A2(n2243), .ZN(n2259) );
  NOR2_X1 U2247 ( .A1(n2068), .A2(n1919), .ZN(n2246) );
  NAND2_X1 U2248 ( .A1(n2243), .A2(n2245), .ZN(n2257) );
  NAND2_X1 U2249 ( .A1(n2260), .A2(n2261), .ZN(n2245) );
  NAND2_X1 U2250 ( .A1(n2262), .A2(b_13_), .ZN(n2261) );
  NOR2_X1 U2251 ( .A1(n2263), .A2(n2009), .ZN(n2262) );
  NOR2_X1 U2252 ( .A1(n2239), .A2(n2241), .ZN(n2263) );
  NAND2_X1 U2253 ( .A1(n2239), .A2(n2241), .ZN(n2260) );
  NAND2_X1 U2254 ( .A1(n2264), .A2(n2265), .ZN(n2241) );
  NAND2_X1 U2255 ( .A1(n2238), .A2(n2266), .ZN(n2265) );
  OR2_X1 U2256 ( .A1(n2237), .A2(n2235), .ZN(n2266) );
  NOR2_X1 U2257 ( .A1(n2068), .A2(n2014), .ZN(n2238) );
  NAND2_X1 U2258 ( .A1(n2235), .A2(n2237), .ZN(n2264) );
  NAND2_X1 U2259 ( .A1(n2267), .A2(n2268), .ZN(n2237) );
  NAND2_X1 U2260 ( .A1(n2269), .A2(b_13_), .ZN(n2268) );
  NOR2_X1 U2261 ( .A1(n2270), .A2(n2019), .ZN(n2269) );
  NOR2_X1 U2262 ( .A1(n2231), .A2(n2233), .ZN(n2270) );
  NAND2_X1 U2263 ( .A1(n2231), .A2(n2233), .ZN(n2267) );
  NAND2_X1 U2264 ( .A1(n2271), .A2(n2272), .ZN(n2233) );
  NAND2_X1 U2265 ( .A1(n2230), .A2(n2273), .ZN(n2272) );
  NAND2_X1 U2266 ( .A1(n2229), .A2(n2228), .ZN(n2273) );
  NOR2_X1 U2267 ( .A1(n2068), .A2(n2170), .ZN(n2230) );
  OR2_X1 U2268 ( .A1(n2228), .A2(n2229), .ZN(n2271) );
  AND2_X1 U2269 ( .A1(n2274), .A2(n2275), .ZN(n2229) );
  NAND2_X1 U2270 ( .A1(n2276), .A2(b_13_), .ZN(n2275) );
  NOR2_X1 U2271 ( .A1(n2277), .A2(n2028), .ZN(n2276) );
  NOR2_X1 U2272 ( .A1(n2223), .A2(n2225), .ZN(n2277) );
  NAND2_X1 U2273 ( .A1(n2223), .A2(n2225), .ZN(n2274) );
  NAND2_X1 U2274 ( .A1(n2278), .A2(n2279), .ZN(n2225) );
  NAND2_X1 U2275 ( .A1(n2222), .A2(n2280), .ZN(n2279) );
  NAND2_X1 U2276 ( .A1(n2221), .A2(n2220), .ZN(n2280) );
  NOR2_X1 U2277 ( .A1(n2068), .A2(n2178), .ZN(n2222) );
  OR2_X1 U2278 ( .A1(n2220), .A2(n2221), .ZN(n2278) );
  AND2_X1 U2279 ( .A1(n2217), .A2(n2281), .ZN(n2221) );
  NAND2_X1 U2280 ( .A1(n2216), .A2(n2218), .ZN(n2281) );
  NAND2_X1 U2281 ( .A1(n2282), .A2(n2283), .ZN(n2218) );
  NAND2_X1 U2282 ( .A1(b_13_), .A2(a_10_), .ZN(n2283) );
  INV_X1 U2283 ( .A(n2284), .ZN(n2282) );
  XNOR2_X1 U2284 ( .A(n2285), .B(n2286), .ZN(n2216) );
  NAND2_X1 U2285 ( .A1(n2287), .A2(n2288), .ZN(n2285) );
  NAND2_X1 U2286 ( .A1(a_10_), .A2(n2284), .ZN(n2217) );
  NAND2_X1 U2287 ( .A1(n2185), .A2(n2289), .ZN(n2284) );
  NAND2_X1 U2288 ( .A1(n2184), .A2(n2186), .ZN(n2289) );
  NAND2_X1 U2289 ( .A1(n2290), .A2(n2291), .ZN(n2186) );
  NAND2_X1 U2290 ( .A1(b_13_), .A2(a_11_), .ZN(n2291) );
  INV_X1 U2291 ( .A(n2292), .ZN(n2290) );
  XNOR2_X1 U2292 ( .A(n2293), .B(n2294), .ZN(n2184) );
  XNOR2_X1 U2293 ( .A(n2295), .B(n2296), .ZN(n2294) );
  NAND2_X1 U2294 ( .A1(a_11_), .A2(n2292), .ZN(n2185) );
  NAND2_X1 U2295 ( .A1(n2297), .A2(n2298), .ZN(n2292) );
  NAND2_X1 U2296 ( .A1(n2299), .A2(b_13_), .ZN(n2298) );
  NOR2_X1 U2297 ( .A1(n2300), .A2(n2057), .ZN(n2299) );
  NOR2_X1 U2298 ( .A1(n2191), .A2(n2193), .ZN(n2300) );
  NAND2_X1 U2299 ( .A1(n2191), .A2(n2193), .ZN(n2297) );
  NAND2_X1 U2300 ( .A1(n2301), .A2(n2302), .ZN(n2193) );
  NAND2_X1 U2301 ( .A1(n2212), .A2(n2303), .ZN(n2302) );
  NAND2_X1 U2302 ( .A1(n2214), .A2(n2213), .ZN(n2303) );
  OR2_X1 U2303 ( .A1(n2213), .A2(n2214), .ZN(n2301) );
  AND2_X1 U2304 ( .A1(n2304), .A2(n2305), .ZN(n2214) );
  NAND2_X1 U2305 ( .A1(n2306), .A2(a_15_), .ZN(n2305) );
  NOR2_X1 U2306 ( .A1(n2307), .A2(n2308), .ZN(n2306) );
  NOR2_X1 U2307 ( .A1(n2070), .A2(n2123), .ZN(n2307) );
  NAND2_X1 U2308 ( .A1(n2309), .A2(b_12_), .ZN(n2304) );
  NOR2_X1 U2309 ( .A1(n2310), .A2(n2208), .ZN(n2309) );
  NOR2_X1 U2310 ( .A1(n2064), .A2(n2308), .ZN(n2310) );
  NAND2_X1 U2311 ( .A1(n2311), .A2(b_13_), .ZN(n2213) );
  NOR2_X1 U2312 ( .A1(n2210), .A2(n2123), .ZN(n2311) );
  XOR2_X1 U2313 ( .A(n2312), .B(n2313), .Z(n2191) );
  XOR2_X1 U2314 ( .A(n2314), .B(n2315), .Z(n2312) );
  XNOR2_X1 U2315 ( .A(n2316), .B(n2317), .ZN(n2220) );
  NOR2_X1 U2316 ( .A1(n2318), .A2(n2319), .ZN(n2317) );
  NOR2_X1 U2317 ( .A1(n2320), .A2(n2321), .ZN(n2318) );
  NOR2_X1 U2318 ( .A1(n1885), .A2(n2123), .ZN(n2320) );
  XOR2_X1 U2319 ( .A(n2322), .B(n2323), .Z(n2223) );
  XOR2_X1 U2320 ( .A(n2324), .B(n2325), .Z(n2322) );
  XNOR2_X1 U2321 ( .A(n2326), .B(n2327), .ZN(n2228) );
  XNOR2_X1 U2322 ( .A(n2328), .B(n2329), .ZN(n2326) );
  NAND2_X1 U2323 ( .A1(b_12_), .A2(a_8_), .ZN(n2328) );
  XNOR2_X1 U2324 ( .A(n2330), .B(n2331), .ZN(n2231) );
  XNOR2_X1 U2325 ( .A(n2332), .B(n2333), .ZN(n2331) );
  XNOR2_X1 U2326 ( .A(n2334), .B(n2335), .ZN(n2235) );
  XOR2_X1 U2327 ( .A(n2336), .B(n2337), .Z(n2335) );
  NAND2_X1 U2328 ( .A1(b_12_), .A2(a_6_), .ZN(n2337) );
  XOR2_X1 U2329 ( .A(n2338), .B(n2339), .Z(n2239) );
  XOR2_X1 U2330 ( .A(n2340), .B(n2341), .Z(n2338) );
  XNOR2_X1 U2331 ( .A(n2342), .B(n2343), .ZN(n2243) );
  XOR2_X1 U2332 ( .A(n2344), .B(n2345), .Z(n2343) );
  NAND2_X1 U2333 ( .A1(b_12_), .A2(a_4_), .ZN(n2345) );
  XNOR2_X1 U2334 ( .A(n2346), .B(n2347), .ZN(n2248) );
  XOR2_X1 U2335 ( .A(n2348), .B(n2349), .Z(n2347) );
  NAND2_X1 U2336 ( .A1(b_12_), .A2(a_3_), .ZN(n2349) );
  XNOR2_X1 U2337 ( .A(n2350), .B(n2351), .ZN(n2139) );
  XNOR2_X1 U2338 ( .A(n2352), .B(n2353), .ZN(n2351) );
  XOR2_X1 U2339 ( .A(n1978), .B(n1977), .Z(n1947) );
  INV_X1 U2340 ( .A(n2354), .ZN(n1977) );
  NAND2_X1 U2341 ( .A1(n2355), .A2(n2356), .ZN(n1950) );
  AND2_X1 U2342 ( .A1(n1968), .A2(n1978), .ZN(n2356) );
  NAND2_X1 U2343 ( .A1(n2357), .A2(n2358), .ZN(n1978) );
  NAND2_X1 U2344 ( .A1(n2359), .A2(b_12_), .ZN(n2358) );
  NOR2_X1 U2345 ( .A1(n2360), .A2(n1986), .ZN(n2359) );
  NOR2_X1 U2346 ( .A1(n2120), .A2(n2121), .ZN(n2360) );
  NAND2_X1 U2347 ( .A1(n2120), .A2(n2121), .ZN(n2357) );
  NAND2_X1 U2348 ( .A1(n2361), .A2(n2362), .ZN(n2121) );
  NAND2_X1 U2349 ( .A1(n2134), .A2(n2363), .ZN(n2362) );
  NAND2_X1 U2350 ( .A1(n2133), .A2(n2132), .ZN(n2363) );
  NOR2_X1 U2351 ( .A1(n2123), .A2(n1995), .ZN(n2134) );
  OR2_X1 U2352 ( .A1(n2132), .A2(n2133), .ZN(n2361) );
  AND2_X1 U2353 ( .A1(n2364), .A2(n2365), .ZN(n2133) );
  NAND2_X1 U2354 ( .A1(n2353), .A2(n2366), .ZN(n2365) );
  OR2_X1 U2355 ( .A1(n2352), .A2(n2350), .ZN(n2366) );
  NOR2_X1 U2356 ( .A1(n2123), .A2(n2000), .ZN(n2353) );
  NAND2_X1 U2357 ( .A1(n2350), .A2(n2352), .ZN(n2364) );
  NAND2_X1 U2358 ( .A1(n2367), .A2(n2368), .ZN(n2352) );
  NAND2_X1 U2359 ( .A1(n2369), .A2(b_12_), .ZN(n2368) );
  NOR2_X1 U2360 ( .A1(n2370), .A2(n1919), .ZN(n2369) );
  NOR2_X1 U2361 ( .A1(n2346), .A2(n2348), .ZN(n2370) );
  NAND2_X1 U2362 ( .A1(n2346), .A2(n2348), .ZN(n2367) );
  NAND2_X1 U2363 ( .A1(n2371), .A2(n2372), .ZN(n2348) );
  NAND2_X1 U2364 ( .A1(n2373), .A2(b_12_), .ZN(n2372) );
  NOR2_X1 U2365 ( .A1(n2374), .A2(n2009), .ZN(n2373) );
  NOR2_X1 U2366 ( .A1(n2342), .A2(n2344), .ZN(n2374) );
  NAND2_X1 U2367 ( .A1(n2342), .A2(n2344), .ZN(n2371) );
  NAND2_X1 U2368 ( .A1(n2375), .A2(n2376), .ZN(n2344) );
  NAND2_X1 U2369 ( .A1(n2341), .A2(n2377), .ZN(n2376) );
  OR2_X1 U2370 ( .A1(n2340), .A2(n2339), .ZN(n2377) );
  NOR2_X1 U2371 ( .A1(n2123), .A2(n2014), .ZN(n2341) );
  NAND2_X1 U2372 ( .A1(n2339), .A2(n2340), .ZN(n2375) );
  NAND2_X1 U2373 ( .A1(n2378), .A2(n2379), .ZN(n2340) );
  NAND2_X1 U2374 ( .A1(n2380), .A2(b_12_), .ZN(n2379) );
  NOR2_X1 U2375 ( .A1(n2381), .A2(n2019), .ZN(n2380) );
  NOR2_X1 U2376 ( .A1(n2334), .A2(n2336), .ZN(n2381) );
  NAND2_X1 U2377 ( .A1(n2334), .A2(n2336), .ZN(n2378) );
  NAND2_X1 U2378 ( .A1(n2382), .A2(n2383), .ZN(n2336) );
  NAND2_X1 U2379 ( .A1(n2333), .A2(n2384), .ZN(n2383) );
  OR2_X1 U2380 ( .A1(n2332), .A2(n2330), .ZN(n2384) );
  NOR2_X1 U2381 ( .A1(n2123), .A2(n2170), .ZN(n2333) );
  NAND2_X1 U2382 ( .A1(n2330), .A2(n2332), .ZN(n2382) );
  NAND2_X1 U2383 ( .A1(n2385), .A2(n2386), .ZN(n2332) );
  NAND2_X1 U2384 ( .A1(n2387), .A2(b_12_), .ZN(n2386) );
  NOR2_X1 U2385 ( .A1(n2388), .A2(n2028), .ZN(n2387) );
  NOR2_X1 U2386 ( .A1(n2327), .A2(n2329), .ZN(n2388) );
  NAND2_X1 U2387 ( .A1(n2327), .A2(n2329), .ZN(n2385) );
  NAND2_X1 U2388 ( .A1(n2389), .A2(n2390), .ZN(n2329) );
  NAND2_X1 U2389 ( .A1(n2325), .A2(n2391), .ZN(n2390) );
  OR2_X1 U2390 ( .A1(n2324), .A2(n2323), .ZN(n2391) );
  NOR2_X1 U2391 ( .A1(n2123), .A2(n2178), .ZN(n2325) );
  NAND2_X1 U2392 ( .A1(n2323), .A2(n2324), .ZN(n2389) );
  OR2_X1 U2393 ( .A1(n2319), .A2(n2392), .ZN(n2324) );
  AND2_X1 U2394 ( .A1(n2316), .A2(n2393), .ZN(n2392) );
  NAND2_X1 U2395 ( .A1(n2394), .A2(n2395), .ZN(n2393) );
  NAND2_X1 U2396 ( .A1(b_12_), .A2(a_10_), .ZN(n2395) );
  XOR2_X1 U2397 ( .A(n2396), .B(n2397), .Z(n2316) );
  XOR2_X1 U2398 ( .A(n2398), .B(n2399), .Z(n2396) );
  NOR2_X1 U2399 ( .A1(n1885), .A2(n2394), .ZN(n2319) );
  INV_X1 U2400 ( .A(n2321), .ZN(n2394) );
  NAND2_X1 U2401 ( .A1(n2287), .A2(n2400), .ZN(n2321) );
  NAND2_X1 U2402 ( .A1(n2286), .A2(n2288), .ZN(n2400) );
  NAND2_X1 U2403 ( .A1(n2401), .A2(n2402), .ZN(n2288) );
  NAND2_X1 U2404 ( .A1(b_12_), .A2(a_11_), .ZN(n2402) );
  INV_X1 U2405 ( .A(n2403), .ZN(n2401) );
  XNOR2_X1 U2406 ( .A(n2404), .B(n2405), .ZN(n2286) );
  XOR2_X1 U2407 ( .A(n2406), .B(n2407), .Z(n2405) );
  NAND2_X1 U2408 ( .A1(a_12_), .A2(b_11_), .ZN(n2407) );
  NAND2_X1 U2409 ( .A1(a_11_), .A2(n2403), .ZN(n2287) );
  NAND2_X1 U2410 ( .A1(n2408), .A2(n2409), .ZN(n2403) );
  NAND2_X1 U2411 ( .A1(n2296), .A2(n2410), .ZN(n2409) );
  OR2_X1 U2412 ( .A1(n2295), .A2(n2293), .ZN(n2410) );
  NAND2_X1 U2413 ( .A1(n2293), .A2(n2295), .ZN(n2408) );
  NAND2_X1 U2414 ( .A1(n2411), .A2(n2412), .ZN(n2295) );
  NAND2_X1 U2415 ( .A1(n2313), .A2(n2413), .ZN(n2412) );
  NAND2_X1 U2416 ( .A1(n2315), .A2(n2314), .ZN(n2413) );
  NOR2_X1 U2417 ( .A1(n2123), .A2(n1870), .ZN(n2313) );
  OR2_X1 U2418 ( .A1(n2314), .A2(n2315), .ZN(n2411) );
  AND2_X1 U2419 ( .A1(n2414), .A2(n2415), .ZN(n2315) );
  NAND2_X1 U2420 ( .A1(n2416), .A2(a_15_), .ZN(n2415) );
  NOR2_X1 U2421 ( .A1(n2417), .A2(n2418), .ZN(n2416) );
  NOR2_X1 U2422 ( .A1(n2070), .A2(n2308), .ZN(n2417) );
  NAND2_X1 U2423 ( .A1(n2419), .A2(a_14_), .ZN(n2414) );
  NOR2_X1 U2424 ( .A1(n2420), .A2(n2308), .ZN(n2419) );
  NOR2_X1 U2425 ( .A1(n2064), .A2(n2418), .ZN(n2420) );
  NAND2_X1 U2426 ( .A1(n2421), .A2(b_12_), .ZN(n2314) );
  NOR2_X1 U2427 ( .A1(n2308), .A2(n2210), .ZN(n2421) );
  XOR2_X1 U2428 ( .A(n2422), .B(n2423), .Z(n2293) );
  XOR2_X1 U2429 ( .A(n2424), .B(n2425), .Z(n2422) );
  XNOR2_X1 U2430 ( .A(n2426), .B(n2427), .ZN(n2323) );
  NAND2_X1 U2431 ( .A1(n2428), .A2(n2429), .ZN(n2426) );
  XNOR2_X1 U2432 ( .A(n2430), .B(n2431), .ZN(n2327) );
  XNOR2_X1 U2433 ( .A(n2432), .B(n2433), .ZN(n2431) );
  XNOR2_X1 U2434 ( .A(n2434), .B(n2435), .ZN(n2330) );
  XOR2_X1 U2435 ( .A(n2436), .B(n2437), .Z(n2435) );
  NAND2_X1 U2436 ( .A1(a_8_), .A2(b_11_), .ZN(n2437) );
  XOR2_X1 U2437 ( .A(n2438), .B(n2439), .Z(n2334) );
  XOR2_X1 U2438 ( .A(n2440), .B(n2441), .Z(n2438) );
  XNOR2_X1 U2439 ( .A(n2442), .B(n2443), .ZN(n2339) );
  XOR2_X1 U2440 ( .A(n2444), .B(n2445), .Z(n2443) );
  NAND2_X1 U2441 ( .A1(a_6_), .A2(b_11_), .ZN(n2445) );
  XNOR2_X1 U2442 ( .A(n2446), .B(n2447), .ZN(n2342) );
  XNOR2_X1 U2443 ( .A(n2448), .B(n2449), .ZN(n2447) );
  XNOR2_X1 U2444 ( .A(n2450), .B(n2451), .ZN(n2346) );
  XNOR2_X1 U2445 ( .A(n2452), .B(n2453), .ZN(n2450) );
  XOR2_X1 U2446 ( .A(n2454), .B(n2455), .Z(n2350) );
  XOR2_X1 U2447 ( .A(n2456), .B(n2457), .Z(n2454) );
  NOR2_X1 U2448 ( .A1(n2308), .A2(n1919), .ZN(n2457) );
  XOR2_X1 U2449 ( .A(n2458), .B(n2459), .Z(n2132) );
  XOR2_X1 U2450 ( .A(n2460), .B(n2461), .Z(n2459) );
  NAND2_X1 U2451 ( .A1(a_2_), .A2(b_11_), .ZN(n2461) );
  XNOR2_X1 U2452 ( .A(n2462), .B(n2463), .ZN(n2120) );
  XOR2_X1 U2453 ( .A(n2464), .B(n2465), .Z(n2463) );
  NAND2_X1 U2454 ( .A1(a_1_), .A2(b_11_), .ZN(n2465) );
  INV_X1 U2455 ( .A(n2466), .ZN(n1968) );
  NOR2_X1 U2456 ( .A1(n2467), .A2(n2354), .ZN(n2355) );
  XOR2_X1 U2457 ( .A(n2468), .B(n2469), .Z(n2354) );
  XOR2_X1 U2458 ( .A(n2470), .B(n2471), .Z(n2468) );
  AND2_X1 U2459 ( .A1(n1976), .A2(n1975), .ZN(n2467) );
  NAND2_X1 U2460 ( .A1(n2472), .A2(n2466), .ZN(n1954) );
  NOR2_X1 U2461 ( .A1(n1976), .A2(n1975), .ZN(n2466) );
  XOR2_X1 U2462 ( .A(n2473), .B(n2474), .Z(n1975) );
  NAND2_X1 U2463 ( .A1(n2475), .A2(n2476), .ZN(n2473) );
  NAND2_X1 U2464 ( .A1(n2477), .A2(n2478), .ZN(n1976) );
  NAND2_X1 U2465 ( .A1(n2469), .A2(n2479), .ZN(n2478) );
  NAND2_X1 U2466 ( .A1(n2471), .A2(n2470), .ZN(n2479) );
  XNOR2_X1 U2467 ( .A(n2480), .B(n2481), .ZN(n2469) );
  XOR2_X1 U2468 ( .A(n2482), .B(n2483), .Z(n2480) );
  OR2_X1 U2469 ( .A1(n2470), .A2(n2471), .ZN(n2477) );
  NOR2_X1 U2470 ( .A1(n1986), .A2(n2308), .ZN(n2471) );
  NAND2_X1 U2471 ( .A1(n2484), .A2(n2485), .ZN(n2470) );
  NAND2_X1 U2472 ( .A1(n2486), .A2(a_1_), .ZN(n2485) );
  NOR2_X1 U2473 ( .A1(n2487), .A2(n2308), .ZN(n2486) );
  NOR2_X1 U2474 ( .A1(n2462), .A2(n2464), .ZN(n2487) );
  NAND2_X1 U2475 ( .A1(n2462), .A2(n2464), .ZN(n2484) );
  NAND2_X1 U2476 ( .A1(n2488), .A2(n2489), .ZN(n2464) );
  NAND2_X1 U2477 ( .A1(n2490), .A2(a_2_), .ZN(n2489) );
  NOR2_X1 U2478 ( .A1(n2491), .A2(n2308), .ZN(n2490) );
  NOR2_X1 U2479 ( .A1(n2458), .A2(n2460), .ZN(n2491) );
  NAND2_X1 U2480 ( .A1(n2458), .A2(n2460), .ZN(n2488) );
  NAND2_X1 U2481 ( .A1(n2492), .A2(n2493), .ZN(n2460) );
  NAND2_X1 U2482 ( .A1(n2494), .A2(a_3_), .ZN(n2493) );
  NOR2_X1 U2483 ( .A1(n2495), .A2(n2308), .ZN(n2494) );
  NOR2_X1 U2484 ( .A1(n2455), .A2(n2456), .ZN(n2495) );
  NAND2_X1 U2485 ( .A1(n2455), .A2(n2456), .ZN(n2492) );
  NAND2_X1 U2486 ( .A1(n2496), .A2(n2497), .ZN(n2456) );
  NAND2_X1 U2487 ( .A1(n2453), .A2(n2498), .ZN(n2497) );
  NAND2_X1 U2488 ( .A1(n2452), .A2(n2451), .ZN(n2498) );
  NOR2_X1 U2489 ( .A1(n2308), .A2(n2009), .ZN(n2453) );
  OR2_X1 U2490 ( .A1(n2451), .A2(n2452), .ZN(n2496) );
  AND2_X1 U2491 ( .A1(n2499), .A2(n2500), .ZN(n2452) );
  NAND2_X1 U2492 ( .A1(n2449), .A2(n2501), .ZN(n2500) );
  OR2_X1 U2493 ( .A1(n2448), .A2(n2446), .ZN(n2501) );
  NOR2_X1 U2494 ( .A1(n2014), .A2(n2308), .ZN(n2449) );
  NAND2_X1 U2495 ( .A1(n2446), .A2(n2448), .ZN(n2499) );
  NAND2_X1 U2496 ( .A1(n2502), .A2(n2503), .ZN(n2448) );
  NAND2_X1 U2497 ( .A1(n2504), .A2(a_6_), .ZN(n2503) );
  NOR2_X1 U2498 ( .A1(n2505), .A2(n2308), .ZN(n2504) );
  NOR2_X1 U2499 ( .A1(n2442), .A2(n2444), .ZN(n2505) );
  NAND2_X1 U2500 ( .A1(n2442), .A2(n2444), .ZN(n2502) );
  NAND2_X1 U2501 ( .A1(n2506), .A2(n2507), .ZN(n2444) );
  NAND2_X1 U2502 ( .A1(n2441), .A2(n2508), .ZN(n2507) );
  OR2_X1 U2503 ( .A1(n2440), .A2(n2439), .ZN(n2508) );
  NOR2_X1 U2504 ( .A1(n2170), .A2(n2308), .ZN(n2441) );
  NAND2_X1 U2505 ( .A1(n2439), .A2(n2440), .ZN(n2506) );
  NAND2_X1 U2506 ( .A1(n2509), .A2(n2510), .ZN(n2440) );
  NAND2_X1 U2507 ( .A1(n2511), .A2(a_8_), .ZN(n2510) );
  NOR2_X1 U2508 ( .A1(n2512), .A2(n2308), .ZN(n2511) );
  NOR2_X1 U2509 ( .A1(n2434), .A2(n2436), .ZN(n2512) );
  NAND2_X1 U2510 ( .A1(n2434), .A2(n2436), .ZN(n2509) );
  NAND2_X1 U2511 ( .A1(n2513), .A2(n2514), .ZN(n2436) );
  NAND2_X1 U2512 ( .A1(n2433), .A2(n2515), .ZN(n2514) );
  OR2_X1 U2513 ( .A1(n2432), .A2(n2430), .ZN(n2515) );
  NOR2_X1 U2514 ( .A1(n2178), .A2(n2308), .ZN(n2433) );
  NAND2_X1 U2515 ( .A1(n2430), .A2(n2432), .ZN(n2513) );
  NAND2_X1 U2516 ( .A1(n2428), .A2(n2516), .ZN(n2432) );
  NAND2_X1 U2517 ( .A1(n2427), .A2(n2429), .ZN(n2516) );
  NAND2_X1 U2518 ( .A1(n2517), .A2(n2518), .ZN(n2429) );
  NAND2_X1 U2519 ( .A1(a_10_), .A2(b_11_), .ZN(n2518) );
  INV_X1 U2520 ( .A(n2519), .ZN(n2517) );
  XNOR2_X1 U2521 ( .A(n2520), .B(n2521), .ZN(n2427) );
  NAND2_X1 U2522 ( .A1(n2522), .A2(n2523), .ZN(n2520) );
  NAND2_X1 U2523 ( .A1(a_10_), .A2(n2519), .ZN(n2428) );
  NAND2_X1 U2524 ( .A1(n2524), .A2(n2525), .ZN(n2519) );
  NAND2_X1 U2525 ( .A1(n2397), .A2(n2526), .ZN(n2525) );
  OR2_X1 U2526 ( .A1(n2398), .A2(n2399), .ZN(n2526) );
  XNOR2_X1 U2527 ( .A(n2527), .B(n2528), .ZN(n2397) );
  XOR2_X1 U2528 ( .A(n2529), .B(n2530), .Z(n2528) );
  NAND2_X1 U2529 ( .A1(a_12_), .A2(b_10_), .ZN(n2530) );
  NAND2_X1 U2530 ( .A1(n2399), .A2(n2398), .ZN(n2524) );
  NAND2_X1 U2531 ( .A1(n2531), .A2(n2532), .ZN(n2398) );
  NAND2_X1 U2532 ( .A1(n2533), .A2(a_12_), .ZN(n2532) );
  NOR2_X1 U2533 ( .A1(n2534), .A2(n2308), .ZN(n2533) );
  NOR2_X1 U2534 ( .A1(n2404), .A2(n2406), .ZN(n2534) );
  NAND2_X1 U2535 ( .A1(n2404), .A2(n2406), .ZN(n2531) );
  NAND2_X1 U2536 ( .A1(n2535), .A2(n2536), .ZN(n2406) );
  NAND2_X1 U2537 ( .A1(n2423), .A2(n2537), .ZN(n2536) );
  NAND2_X1 U2538 ( .A1(n2425), .A2(n2424), .ZN(n2537) );
  NOR2_X1 U2539 ( .A1(n1870), .A2(n2308), .ZN(n2423) );
  OR2_X1 U2540 ( .A1(n2424), .A2(n2425), .ZN(n2535) );
  AND2_X1 U2541 ( .A1(n2538), .A2(n2539), .ZN(n2425) );
  NAND2_X1 U2542 ( .A1(n2540), .A2(b_10_), .ZN(n2539) );
  NOR2_X1 U2543 ( .A1(n2541), .A2(n2208), .ZN(n2540) );
  NOR2_X1 U2544 ( .A1(n2064), .A2(n2542), .ZN(n2541) );
  NAND2_X1 U2545 ( .A1(n2543), .A2(a_15_), .ZN(n2538) );
  NOR2_X1 U2546 ( .A1(n2544), .A2(n2542), .ZN(n2543) );
  NOR2_X1 U2547 ( .A1(n2070), .A2(n2418), .ZN(n2544) );
  NAND2_X1 U2548 ( .A1(n2545), .A2(n2546), .ZN(n2424) );
  NOR2_X1 U2549 ( .A1(n2308), .A2(n2418), .ZN(n2545) );
  XOR2_X1 U2550 ( .A(n2547), .B(n2548), .Z(n2404) );
  XOR2_X1 U2551 ( .A(n2549), .B(n2550), .Z(n2547) );
  XOR2_X1 U2552 ( .A(n2551), .B(n2552), .Z(n2430) );
  XOR2_X1 U2553 ( .A(n2553), .B(n2554), .Z(n2551) );
  XOR2_X1 U2554 ( .A(n2555), .B(n2556), .Z(n2434) );
  XOR2_X1 U2555 ( .A(n2557), .B(n2558), .Z(n2555) );
  XOR2_X1 U2556 ( .A(n2559), .B(n2560), .Z(n2439) );
  XOR2_X1 U2557 ( .A(n2561), .B(n2562), .Z(n2559) );
  NOR2_X1 U2558 ( .A1(n2418), .A2(n2028), .ZN(n2562) );
  XNOR2_X1 U2559 ( .A(n2563), .B(n2564), .ZN(n2442) );
  XNOR2_X1 U2560 ( .A(n2565), .B(n2566), .ZN(n2564) );
  XOR2_X1 U2561 ( .A(n2567), .B(n2568), .Z(n2446) );
  XOR2_X1 U2562 ( .A(n2569), .B(n2570), .Z(n2567) );
  NOR2_X1 U2563 ( .A1(n2418), .A2(n2019), .ZN(n2570) );
  XOR2_X1 U2564 ( .A(n2571), .B(n2572), .Z(n2451) );
  XOR2_X1 U2565 ( .A(n2573), .B(n2574), .Z(n2572) );
  NAND2_X1 U2566 ( .A1(b_10_), .A2(a_5_), .ZN(n2574) );
  XNOR2_X1 U2567 ( .A(n2575), .B(n2576), .ZN(n2455) );
  XNOR2_X1 U2568 ( .A(n2577), .B(n2578), .ZN(n2576) );
  XNOR2_X1 U2569 ( .A(n2579), .B(n2580), .ZN(n2458) );
  XNOR2_X1 U2570 ( .A(n2581), .B(n2582), .ZN(n2579) );
  XOR2_X1 U2571 ( .A(n2583), .B(n2584), .Z(n2462) );
  XOR2_X1 U2572 ( .A(n2585), .B(n2586), .Z(n2583) );
  NOR2_X1 U2573 ( .A1(n2418), .A2(n2000), .ZN(n2586) );
  XOR2_X1 U2574 ( .A(n1969), .B(n1970), .Z(n2472) );
  NAND2_X1 U2575 ( .A1(n2587), .A2(n2588), .ZN(n1828) );
  NAND2_X1 U2576 ( .A1(n1970), .A2(n1969), .ZN(n2588) );
  XOR2_X1 U2577 ( .A(n2589), .B(n2590), .Z(n2587) );
  NAND2_X1 U2578 ( .A1(n2591), .A2(n2592), .ZN(n1829) );
  XOR2_X1 U2579 ( .A(n2593), .B(n2590), .Z(n2592) );
  AND2_X1 U2580 ( .A1(n1969), .A2(n1970), .ZN(n2591) );
  XNOR2_X1 U2581 ( .A(n2594), .B(n2595), .ZN(n1970) );
  XOR2_X1 U2582 ( .A(n2596), .B(n2597), .Z(n2595) );
  NAND2_X1 U2583 ( .A1(a_0_), .A2(b_9_), .ZN(n2597) );
  NAND2_X1 U2584 ( .A1(n2475), .A2(n2598), .ZN(n1969) );
  NAND2_X1 U2585 ( .A1(n2474), .A2(n2476), .ZN(n2598) );
  NAND2_X1 U2586 ( .A1(n2599), .A2(n2600), .ZN(n2476) );
  NAND2_X1 U2587 ( .A1(a_0_), .A2(b_10_), .ZN(n2600) );
  INV_X1 U2588 ( .A(n2601), .ZN(n2599) );
  XNOR2_X1 U2589 ( .A(n2602), .B(n2603), .ZN(n2474) );
  XOR2_X1 U2590 ( .A(n2604), .B(n2605), .Z(n2603) );
  NAND2_X1 U2591 ( .A1(a_1_), .A2(b_9_), .ZN(n2605) );
  NAND2_X1 U2592 ( .A1(a_0_), .A2(n2601), .ZN(n2475) );
  NAND2_X1 U2593 ( .A1(n2606), .A2(n2607), .ZN(n2601) );
  NAND2_X1 U2594 ( .A1(n2483), .A2(n2608), .ZN(n2607) );
  OR2_X1 U2595 ( .A1(n2481), .A2(n2482), .ZN(n2608) );
  NOR2_X1 U2596 ( .A1(n1995), .A2(n2418), .ZN(n2483) );
  NAND2_X1 U2597 ( .A1(n2481), .A2(n2482), .ZN(n2606) );
  NAND2_X1 U2598 ( .A1(n2609), .A2(n2610), .ZN(n2482) );
  NAND2_X1 U2599 ( .A1(n2611), .A2(a_2_), .ZN(n2610) );
  NOR2_X1 U2600 ( .A1(n2612), .A2(n2418), .ZN(n2611) );
  NOR2_X1 U2601 ( .A1(n2584), .A2(n2585), .ZN(n2612) );
  NAND2_X1 U2602 ( .A1(n2584), .A2(n2585), .ZN(n2609) );
  NAND2_X1 U2603 ( .A1(n2613), .A2(n2614), .ZN(n2585) );
  NAND2_X1 U2604 ( .A1(n2581), .A2(n2615), .ZN(n2614) );
  NAND2_X1 U2605 ( .A1(n2582), .A2(n2580), .ZN(n2615) );
  NOR2_X1 U2606 ( .A1(n1919), .A2(n2418), .ZN(n2581) );
  OR2_X1 U2607 ( .A1(n2580), .A2(n2582), .ZN(n2613) );
  AND2_X1 U2608 ( .A1(n2616), .A2(n2617), .ZN(n2582) );
  NAND2_X1 U2609 ( .A1(n2578), .A2(n2618), .ZN(n2617) );
  OR2_X1 U2610 ( .A1(n2575), .A2(n2577), .ZN(n2618) );
  NOR2_X1 U2611 ( .A1(n2418), .A2(n2009), .ZN(n2578) );
  NAND2_X1 U2612 ( .A1(n2575), .A2(n2577), .ZN(n2616) );
  NAND2_X1 U2613 ( .A1(n2619), .A2(n2620), .ZN(n2577) );
  NAND2_X1 U2614 ( .A1(n2621), .A2(b_10_), .ZN(n2620) );
  NOR2_X1 U2615 ( .A1(n2622), .A2(n2014), .ZN(n2621) );
  NOR2_X1 U2616 ( .A1(n2573), .A2(n2571), .ZN(n2622) );
  NAND2_X1 U2617 ( .A1(n2571), .A2(n2573), .ZN(n2619) );
  NAND2_X1 U2618 ( .A1(n2623), .A2(n2624), .ZN(n2573) );
  NAND2_X1 U2619 ( .A1(n2625), .A2(a_6_), .ZN(n2624) );
  NOR2_X1 U2620 ( .A1(n2626), .A2(n2418), .ZN(n2625) );
  NOR2_X1 U2621 ( .A1(n2569), .A2(n2568), .ZN(n2626) );
  NAND2_X1 U2622 ( .A1(n2568), .A2(n2569), .ZN(n2623) );
  NAND2_X1 U2623 ( .A1(n2627), .A2(n2628), .ZN(n2569) );
  NAND2_X1 U2624 ( .A1(n2566), .A2(n2629), .ZN(n2628) );
  OR2_X1 U2625 ( .A1(n2563), .A2(n2565), .ZN(n2629) );
  NOR2_X1 U2626 ( .A1(n2418), .A2(n2170), .ZN(n2566) );
  NAND2_X1 U2627 ( .A1(n2563), .A2(n2565), .ZN(n2627) );
  NAND2_X1 U2628 ( .A1(n2630), .A2(n2631), .ZN(n2565) );
  NAND2_X1 U2629 ( .A1(n2632), .A2(a_8_), .ZN(n2631) );
  NOR2_X1 U2630 ( .A1(n2633), .A2(n2418), .ZN(n2632) );
  NOR2_X1 U2631 ( .A1(n2560), .A2(n2561), .ZN(n2633) );
  NAND2_X1 U2632 ( .A1(n2560), .A2(n2561), .ZN(n2630) );
  NAND2_X1 U2633 ( .A1(n2634), .A2(n2635), .ZN(n2561) );
  NAND2_X1 U2634 ( .A1(n2558), .A2(n2636), .ZN(n2635) );
  OR2_X1 U2635 ( .A1(n2556), .A2(n2557), .ZN(n2636) );
  NOR2_X1 U2636 ( .A1(n2418), .A2(n2178), .ZN(n2558) );
  NAND2_X1 U2637 ( .A1(n2556), .A2(n2557), .ZN(n2634) );
  NAND2_X1 U2638 ( .A1(n2637), .A2(n2638), .ZN(n2557) );
  NAND2_X1 U2639 ( .A1(n2554), .A2(n2639), .ZN(n2638) );
  OR2_X1 U2640 ( .A1(n2552), .A2(n2553), .ZN(n2639) );
  INV_X1 U2641 ( .A(n2640), .ZN(n2554) );
  NAND2_X1 U2642 ( .A1(n2552), .A2(n2553), .ZN(n2637) );
  NAND2_X1 U2643 ( .A1(n2522), .A2(n2641), .ZN(n2553) );
  NAND2_X1 U2644 ( .A1(n2521), .A2(n2523), .ZN(n2641) );
  NAND2_X1 U2645 ( .A1(n2642), .A2(n2643), .ZN(n2523) );
  NAND2_X1 U2646 ( .A1(b_10_), .A2(a_11_), .ZN(n2643) );
  INV_X1 U2647 ( .A(n2644), .ZN(n2642) );
  XNOR2_X1 U2648 ( .A(n2645), .B(n2646), .ZN(n2521) );
  XOR2_X1 U2649 ( .A(n2647), .B(n2648), .Z(n2646) );
  NAND2_X1 U2650 ( .A1(a_12_), .A2(b_9_), .ZN(n2648) );
  NAND2_X1 U2651 ( .A1(a_11_), .A2(n2644), .ZN(n2522) );
  NAND2_X1 U2652 ( .A1(n2649), .A2(n2650), .ZN(n2644) );
  NAND2_X1 U2653 ( .A1(n2651), .A2(a_12_), .ZN(n2650) );
  NOR2_X1 U2654 ( .A1(n2652), .A2(n2418), .ZN(n2651) );
  NOR2_X1 U2655 ( .A1(n2527), .A2(n2529), .ZN(n2652) );
  NAND2_X1 U2656 ( .A1(n2527), .A2(n2529), .ZN(n2649) );
  NAND2_X1 U2657 ( .A1(n2653), .A2(n2654), .ZN(n2529) );
  NAND2_X1 U2658 ( .A1(n2548), .A2(n2655), .ZN(n2654) );
  NAND2_X1 U2659 ( .A1(n2550), .A2(n2549), .ZN(n2655) );
  NOR2_X1 U2660 ( .A1(n2418), .A2(n1870), .ZN(n2548) );
  OR2_X1 U2661 ( .A1(n2549), .A2(n2550), .ZN(n2653) );
  AND2_X1 U2662 ( .A1(n2656), .A2(n2657), .ZN(n2550) );
  NAND2_X1 U2663 ( .A1(n2658), .A2(b_8_), .ZN(n2657) );
  NOR2_X1 U2664 ( .A1(n2659), .A2(n2071), .ZN(n2658) );
  NOR2_X1 U2665 ( .A1(n2070), .A2(n2542), .ZN(n2659) );
  NAND2_X1 U2666 ( .A1(n2660), .A2(b_9_), .ZN(n2656) );
  NOR2_X1 U2667 ( .A1(n2661), .A2(n2208), .ZN(n2660) );
  NOR2_X1 U2668 ( .A1(n2064), .A2(n2662), .ZN(n2661) );
  NAND2_X1 U2669 ( .A1(n2663), .A2(n2546), .ZN(n2549) );
  INV_X1 U2670 ( .A(n2210), .ZN(n2546) );
  NOR2_X1 U2671 ( .A1(n2542), .A2(n2418), .ZN(n2663) );
  XOR2_X1 U2672 ( .A(n2664), .B(n2665), .Z(n2527) );
  XOR2_X1 U2673 ( .A(n2666), .B(n2667), .Z(n2664) );
  XNOR2_X1 U2674 ( .A(n2668), .B(n2669), .ZN(n2552) );
  NAND2_X1 U2675 ( .A1(n2670), .A2(n2671), .ZN(n2668) );
  XNOR2_X1 U2676 ( .A(n2672), .B(n2673), .ZN(n2556) );
  NAND2_X1 U2677 ( .A1(n2674), .A2(n2675), .ZN(n2672) );
  XNOR2_X1 U2678 ( .A(n2676), .B(n2677), .ZN(n2560) );
  XOR2_X1 U2679 ( .A(n2678), .B(n2679), .Z(n2677) );
  XOR2_X1 U2680 ( .A(n2680), .B(n2681), .Z(n2563) );
  XOR2_X1 U2681 ( .A(n2682), .B(n2683), .Z(n2680) );
  NOR2_X1 U2682 ( .A1(n2542), .A2(n2028), .ZN(n2683) );
  XNOR2_X1 U2683 ( .A(n2684), .B(n2685), .ZN(n2568) );
  XNOR2_X1 U2684 ( .A(n2686), .B(n2687), .ZN(n2685) );
  XNOR2_X1 U2685 ( .A(n2688), .B(n2689), .ZN(n2571) );
  XNOR2_X1 U2686 ( .A(n2690), .B(n2691), .ZN(n2689) );
  XNOR2_X1 U2687 ( .A(n2692), .B(n2693), .ZN(n2575) );
  XOR2_X1 U2688 ( .A(n2694), .B(n2695), .Z(n2693) );
  NAND2_X1 U2689 ( .A1(b_9_), .A2(a_5_), .ZN(n2695) );
  XOR2_X1 U2690 ( .A(n2696), .B(n2697), .Z(n2580) );
  NAND2_X1 U2691 ( .A1(n2698), .A2(n2699), .ZN(n2696) );
  XOR2_X1 U2692 ( .A(n2700), .B(n2701), .Z(n2584) );
  XOR2_X1 U2693 ( .A(n2702), .B(n2703), .Z(n2700) );
  NOR2_X1 U2694 ( .A1(n2542), .A2(n1919), .ZN(n2703) );
  XNOR2_X1 U2695 ( .A(n2704), .B(n2705), .ZN(n2481) );
  XOR2_X1 U2696 ( .A(n2706), .B(n2707), .Z(n2705) );
  NAND2_X1 U2697 ( .A1(a_2_), .A2(b_9_), .ZN(n2707) );
  NAND2_X1 U2698 ( .A1(n2708), .A2(n2709), .ZN(n1832) );
  NAND2_X1 U2699 ( .A1(n2590), .A2(n2593), .ZN(n2709) );
  NAND2_X1 U2700 ( .A1(n2710), .A2(n2590), .ZN(n1833) );
  XOR2_X1 U2701 ( .A(n2711), .B(n2712), .Z(n2590) );
  XOR2_X1 U2702 ( .A(n2713), .B(n2714), .Z(n2711) );
  NOR2_X1 U2703 ( .A1(n2589), .A2(n2708), .ZN(n2710) );
  XOR2_X1 U2704 ( .A(n2715), .B(n2716), .Z(n2708) );
  INV_X1 U2705 ( .A(n2717), .ZN(n2716) );
  INV_X1 U2706 ( .A(n2593), .ZN(n2589) );
  NAND2_X1 U2707 ( .A1(n2718), .A2(n2719), .ZN(n2593) );
  NAND2_X1 U2708 ( .A1(n2720), .A2(a_0_), .ZN(n2719) );
  NOR2_X1 U2709 ( .A1(n2721), .A2(n2542), .ZN(n2720) );
  NOR2_X1 U2710 ( .A1(n2594), .A2(n2596), .ZN(n2721) );
  NAND2_X1 U2711 ( .A1(n2594), .A2(n2596), .ZN(n2718) );
  NAND2_X1 U2712 ( .A1(n2722), .A2(n2723), .ZN(n2596) );
  NAND2_X1 U2713 ( .A1(n2724), .A2(a_1_), .ZN(n2723) );
  NOR2_X1 U2714 ( .A1(n2725), .A2(n2542), .ZN(n2724) );
  NOR2_X1 U2715 ( .A1(n2604), .A2(n2602), .ZN(n2725) );
  NAND2_X1 U2716 ( .A1(n2602), .A2(n2604), .ZN(n2722) );
  NAND2_X1 U2717 ( .A1(n2726), .A2(n2727), .ZN(n2604) );
  NAND2_X1 U2718 ( .A1(n2728), .A2(a_2_), .ZN(n2727) );
  NOR2_X1 U2719 ( .A1(n2729), .A2(n2542), .ZN(n2728) );
  NOR2_X1 U2720 ( .A1(n2704), .A2(n2706), .ZN(n2729) );
  NAND2_X1 U2721 ( .A1(n2704), .A2(n2706), .ZN(n2726) );
  NAND2_X1 U2722 ( .A1(n2730), .A2(n2731), .ZN(n2706) );
  NAND2_X1 U2723 ( .A1(n2732), .A2(a_3_), .ZN(n2731) );
  NOR2_X1 U2724 ( .A1(n2733), .A2(n2542), .ZN(n2732) );
  NOR2_X1 U2725 ( .A1(n2702), .A2(n2701), .ZN(n2733) );
  NAND2_X1 U2726 ( .A1(n2701), .A2(n2702), .ZN(n2730) );
  NAND2_X1 U2727 ( .A1(n2698), .A2(n2734), .ZN(n2702) );
  NAND2_X1 U2728 ( .A1(n2697), .A2(n2699), .ZN(n2734) );
  NAND2_X1 U2729 ( .A1(n2735), .A2(n2736), .ZN(n2699) );
  NAND2_X1 U2730 ( .A1(b_9_), .A2(a_4_), .ZN(n2736) );
  INV_X1 U2731 ( .A(n2737), .ZN(n2735) );
  XNOR2_X1 U2732 ( .A(n2738), .B(n2739), .ZN(n2697) );
  XOR2_X1 U2733 ( .A(n2740), .B(n2741), .Z(n2739) );
  NAND2_X1 U2734 ( .A1(b_8_), .A2(a_5_), .ZN(n2741) );
  NAND2_X1 U2735 ( .A1(a_4_), .A2(n2737), .ZN(n2698) );
  NAND2_X1 U2736 ( .A1(n2742), .A2(n2743), .ZN(n2737) );
  NAND2_X1 U2737 ( .A1(n2744), .A2(b_9_), .ZN(n2743) );
  NOR2_X1 U2738 ( .A1(n2745), .A2(n2014), .ZN(n2744) );
  NOR2_X1 U2739 ( .A1(n2692), .A2(n2694), .ZN(n2745) );
  NAND2_X1 U2740 ( .A1(n2692), .A2(n2694), .ZN(n2742) );
  NAND2_X1 U2741 ( .A1(n2746), .A2(n2747), .ZN(n2694) );
  NAND2_X1 U2742 ( .A1(n2691), .A2(n2748), .ZN(n2747) );
  OR2_X1 U2743 ( .A1(n2690), .A2(n2688), .ZN(n2748) );
  NOR2_X1 U2744 ( .A1(n2019), .A2(n2542), .ZN(n2691) );
  NAND2_X1 U2745 ( .A1(n2688), .A2(n2690), .ZN(n2746) );
  NAND2_X1 U2746 ( .A1(n2749), .A2(n2750), .ZN(n2690) );
  NAND2_X1 U2747 ( .A1(n2687), .A2(n2751), .ZN(n2750) );
  OR2_X1 U2748 ( .A1(n2686), .A2(n2684), .ZN(n2751) );
  NOR2_X1 U2749 ( .A1(n2542), .A2(n2170), .ZN(n2687) );
  NAND2_X1 U2750 ( .A1(n2684), .A2(n2686), .ZN(n2749) );
  NAND2_X1 U2751 ( .A1(n2752), .A2(n2753), .ZN(n2686) );
  NAND2_X1 U2752 ( .A1(n2754), .A2(a_8_), .ZN(n2753) );
  NOR2_X1 U2753 ( .A1(n2755), .A2(n2542), .ZN(n2754) );
  NOR2_X1 U2754 ( .A1(n2681), .A2(n2682), .ZN(n2755) );
  NAND2_X1 U2755 ( .A1(n2681), .A2(n2682), .ZN(n2752) );
  NAND2_X1 U2756 ( .A1(n2756), .A2(n2757), .ZN(n2682) );
  NAND2_X1 U2757 ( .A1(n2758), .A2(n2759), .ZN(n2757) );
  OR2_X1 U2758 ( .A1(n2676), .A2(n2678), .ZN(n2759) );
  NAND2_X1 U2759 ( .A1(n2676), .A2(n2678), .ZN(n2756) );
  NAND2_X1 U2760 ( .A1(n2674), .A2(n2760), .ZN(n2678) );
  NAND2_X1 U2761 ( .A1(n2673), .A2(n2675), .ZN(n2760) );
  NAND2_X1 U2762 ( .A1(n2761), .A2(n2762), .ZN(n2675) );
  NAND2_X1 U2763 ( .A1(a_10_), .A2(b_9_), .ZN(n2762) );
  INV_X1 U2764 ( .A(n2763), .ZN(n2761) );
  XNOR2_X1 U2765 ( .A(n2764), .B(n2765), .ZN(n2673) );
  NAND2_X1 U2766 ( .A1(n2766), .A2(n2767), .ZN(n2764) );
  NAND2_X1 U2767 ( .A1(a_10_), .A2(n2763), .ZN(n2674) );
  NAND2_X1 U2768 ( .A1(n2670), .A2(n2768), .ZN(n2763) );
  NAND2_X1 U2769 ( .A1(n2669), .A2(n2671), .ZN(n2768) );
  NAND2_X1 U2770 ( .A1(n2769), .A2(n2770), .ZN(n2671) );
  NAND2_X1 U2771 ( .A1(b_9_), .A2(a_11_), .ZN(n2770) );
  INV_X1 U2772 ( .A(n2771), .ZN(n2769) );
  XNOR2_X1 U2773 ( .A(n2772), .B(n2773), .ZN(n2669) );
  XOR2_X1 U2774 ( .A(n2774), .B(n2775), .Z(n2773) );
  NAND2_X1 U2775 ( .A1(a_12_), .A2(b_8_), .ZN(n2775) );
  NAND2_X1 U2776 ( .A1(a_11_), .A2(n2771), .ZN(n2670) );
  NAND2_X1 U2777 ( .A1(n2776), .A2(n2777), .ZN(n2771) );
  NAND2_X1 U2778 ( .A1(n2778), .A2(a_12_), .ZN(n2777) );
  NOR2_X1 U2779 ( .A1(n2779), .A2(n2542), .ZN(n2778) );
  NOR2_X1 U2780 ( .A1(n2645), .A2(n2647), .ZN(n2779) );
  NAND2_X1 U2781 ( .A1(n2645), .A2(n2647), .ZN(n2776) );
  NAND2_X1 U2782 ( .A1(n2780), .A2(n2781), .ZN(n2647) );
  NAND2_X1 U2783 ( .A1(n2665), .A2(n2782), .ZN(n2781) );
  NAND2_X1 U2784 ( .A1(n2667), .A2(n2666), .ZN(n2782) );
  NOR2_X1 U2785 ( .A1(n2542), .A2(n1870), .ZN(n2665) );
  OR2_X1 U2786 ( .A1(n2666), .A2(n2667), .ZN(n2780) );
  AND2_X1 U2787 ( .A1(n2783), .A2(n2784), .ZN(n2667) );
  NAND2_X1 U2788 ( .A1(n2785), .A2(b_7_), .ZN(n2784) );
  NOR2_X1 U2789 ( .A1(n2786), .A2(n2071), .ZN(n2785) );
  NOR2_X1 U2790 ( .A1(n2070), .A2(n2662), .ZN(n2786) );
  NAND2_X1 U2791 ( .A1(n2787), .A2(b_8_), .ZN(n2783) );
  NOR2_X1 U2792 ( .A1(n2788), .A2(n2208), .ZN(n2787) );
  NOR2_X1 U2793 ( .A1(n2064), .A2(n2789), .ZN(n2788) );
  NAND2_X1 U2794 ( .A1(n2790), .A2(b_8_), .ZN(n2666) );
  NOR2_X1 U2795 ( .A1(n2542), .A2(n2210), .ZN(n2790) );
  XOR2_X1 U2796 ( .A(n2791), .B(n2792), .Z(n2645) );
  XOR2_X1 U2797 ( .A(n2793), .B(n2794), .Z(n2791) );
  XNOR2_X1 U2798 ( .A(n2795), .B(n2796), .ZN(n2676) );
  NAND2_X1 U2799 ( .A1(n2797), .A2(n2798), .ZN(n2795) );
  XNOR2_X1 U2800 ( .A(n2799), .B(n2800), .ZN(n2681) );
  XNOR2_X1 U2801 ( .A(n2801), .B(n2802), .ZN(n2800) );
  XOR2_X1 U2802 ( .A(n2803), .B(n2804), .Z(n2684) );
  XOR2_X1 U2803 ( .A(n2805), .B(n2806), .Z(n2803) );
  XOR2_X1 U2804 ( .A(n2807), .B(n2808), .Z(n2688) );
  XOR2_X1 U2805 ( .A(n2809), .B(n2810), .Z(n2807) );
  NOR2_X1 U2806 ( .A1(n2170), .A2(n2662), .ZN(n2810) );
  XOR2_X1 U2807 ( .A(n2811), .B(n2812), .Z(n2692) );
  XNOR2_X1 U2808 ( .A(n2813), .B(n2814), .ZN(n2811) );
  NAND2_X1 U2809 ( .A1(a_6_), .A2(b_8_), .ZN(n2813) );
  XNOR2_X1 U2810 ( .A(n2815), .B(n2816), .ZN(n2701) );
  XOR2_X1 U2811 ( .A(n2817), .B(n2818), .Z(n2816) );
  NAND2_X1 U2812 ( .A1(b_8_), .A2(a_4_), .ZN(n2818) );
  XNOR2_X1 U2813 ( .A(n2819), .B(n2820), .ZN(n2704) );
  XNOR2_X1 U2814 ( .A(n2821), .B(n2822), .ZN(n2820) );
  XOR2_X1 U2815 ( .A(n2823), .B(n2824), .Z(n2602) );
  XOR2_X1 U2816 ( .A(n2825), .B(n2826), .Z(n2823) );
  XOR2_X1 U2817 ( .A(n2827), .B(n2828), .Z(n2594) );
  XOR2_X1 U2818 ( .A(n2829), .B(n2830), .Z(n2827) );
  NAND2_X1 U2819 ( .A1(n2831), .A2(n2832), .ZN(n1836) );
  NAND2_X1 U2820 ( .A1(n2717), .A2(n2715), .ZN(n2832) );
  NAND2_X1 U2821 ( .A1(n2833), .A2(n2717), .ZN(n1837) );
  XNOR2_X1 U2822 ( .A(n2834), .B(n2835), .ZN(n2717) );
  XOR2_X1 U2823 ( .A(n2836), .B(n2837), .Z(n2835) );
  NAND2_X1 U2824 ( .A1(a_0_), .A2(b_7_), .ZN(n2837) );
  NOR2_X1 U2825 ( .A1(n2838), .A2(n2831), .ZN(n2833) );
  XOR2_X1 U2826 ( .A(n2839), .B(n2840), .Z(n2831) );
  INV_X1 U2827 ( .A(n2841), .ZN(n2840) );
  INV_X1 U2828 ( .A(n2715), .ZN(n2838) );
  NAND2_X1 U2829 ( .A1(n2842), .A2(n2843), .ZN(n2715) );
  NAND2_X1 U2830 ( .A1(n2714), .A2(n2844), .ZN(n2843) );
  OR2_X1 U2831 ( .A1(n2712), .A2(n2713), .ZN(n2844) );
  NOR2_X1 U2832 ( .A1(n1986), .A2(n2662), .ZN(n2714) );
  NAND2_X1 U2833 ( .A1(n2712), .A2(n2713), .ZN(n2842) );
  NAND2_X1 U2834 ( .A1(n2845), .A2(n2846), .ZN(n2713) );
  NAND2_X1 U2835 ( .A1(n2829), .A2(n2847), .ZN(n2846) );
  OR2_X1 U2836 ( .A1(n2828), .A2(n2830), .ZN(n2847) );
  NOR2_X1 U2837 ( .A1(n1995), .A2(n2662), .ZN(n2829) );
  NAND2_X1 U2838 ( .A1(n2828), .A2(n2830), .ZN(n2845) );
  NAND2_X1 U2839 ( .A1(n2848), .A2(n2849), .ZN(n2830) );
  NAND2_X1 U2840 ( .A1(n2826), .A2(n2850), .ZN(n2849) );
  OR2_X1 U2841 ( .A1(n2825), .A2(n2824), .ZN(n2850) );
  NOR2_X1 U2842 ( .A1(n2000), .A2(n2662), .ZN(n2826) );
  NAND2_X1 U2843 ( .A1(n2824), .A2(n2825), .ZN(n2848) );
  NAND2_X1 U2844 ( .A1(n2851), .A2(n2852), .ZN(n2825) );
  NAND2_X1 U2845 ( .A1(n2822), .A2(n2853), .ZN(n2852) );
  OR2_X1 U2846 ( .A1(n2819), .A2(n2821), .ZN(n2853) );
  NOR2_X1 U2847 ( .A1(n1919), .A2(n2662), .ZN(n2822) );
  NAND2_X1 U2848 ( .A1(n2819), .A2(n2821), .ZN(n2851) );
  NAND2_X1 U2849 ( .A1(n2854), .A2(n2855), .ZN(n2821) );
  NAND2_X1 U2850 ( .A1(n2856), .A2(b_8_), .ZN(n2855) );
  NOR2_X1 U2851 ( .A1(n2857), .A2(n2009), .ZN(n2856) );
  NOR2_X1 U2852 ( .A1(n2815), .A2(n2817), .ZN(n2857) );
  NAND2_X1 U2853 ( .A1(n2815), .A2(n2817), .ZN(n2854) );
  NAND2_X1 U2854 ( .A1(n2858), .A2(n2859), .ZN(n2817) );
  NAND2_X1 U2855 ( .A1(n2860), .A2(b_8_), .ZN(n2859) );
  NOR2_X1 U2856 ( .A1(n2861), .A2(n2014), .ZN(n2860) );
  NOR2_X1 U2857 ( .A1(n2740), .A2(n2738), .ZN(n2861) );
  NAND2_X1 U2858 ( .A1(n2738), .A2(n2740), .ZN(n2858) );
  NAND2_X1 U2859 ( .A1(n2862), .A2(n2863), .ZN(n2740) );
  NAND2_X1 U2860 ( .A1(n2864), .A2(a_6_), .ZN(n2863) );
  NOR2_X1 U2861 ( .A1(n2865), .A2(n2662), .ZN(n2864) );
  NOR2_X1 U2862 ( .A1(n2814), .A2(n2812), .ZN(n2865) );
  NAND2_X1 U2863 ( .A1(n2812), .A2(n2814), .ZN(n2862) );
  NAND2_X1 U2864 ( .A1(n2866), .A2(n2867), .ZN(n2814) );
  NAND2_X1 U2865 ( .A1(n2868), .A2(b_8_), .ZN(n2867) );
  NOR2_X1 U2866 ( .A1(n2869), .A2(n2170), .ZN(n2868) );
  NOR2_X1 U2867 ( .A1(n2809), .A2(n2808), .ZN(n2869) );
  NAND2_X1 U2868 ( .A1(n2808), .A2(n2809), .ZN(n2866) );
  NAND2_X1 U2869 ( .A1(n2870), .A2(n2871), .ZN(n2809) );
  NAND2_X1 U2870 ( .A1(n2806), .A2(n2872), .ZN(n2871) );
  OR2_X1 U2871 ( .A1(n2804), .A2(n2805), .ZN(n2872) );
  INV_X1 U2872 ( .A(n2873), .ZN(n2806) );
  NAND2_X1 U2873 ( .A1(n2804), .A2(n2805), .ZN(n2870) );
  NAND2_X1 U2874 ( .A1(n2874), .A2(n2875), .ZN(n2805) );
  NAND2_X1 U2875 ( .A1(n2802), .A2(n2876), .ZN(n2875) );
  OR2_X1 U2876 ( .A1(n2799), .A2(n2801), .ZN(n2876) );
  NOR2_X1 U2877 ( .A1(n2662), .A2(n2178), .ZN(n2802) );
  NAND2_X1 U2878 ( .A1(n2799), .A2(n2801), .ZN(n2874) );
  NAND2_X1 U2879 ( .A1(n2797), .A2(n2877), .ZN(n2801) );
  NAND2_X1 U2880 ( .A1(n2796), .A2(n2798), .ZN(n2877) );
  NAND2_X1 U2881 ( .A1(n2878), .A2(n2879), .ZN(n2798) );
  NAND2_X1 U2882 ( .A1(a_10_), .A2(b_8_), .ZN(n2879) );
  INV_X1 U2883 ( .A(n2880), .ZN(n2878) );
  XNOR2_X1 U2884 ( .A(n2881), .B(n2882), .ZN(n2796) );
  NAND2_X1 U2885 ( .A1(n2883), .A2(n2884), .ZN(n2881) );
  NAND2_X1 U2886 ( .A1(a_10_), .A2(n2880), .ZN(n2797) );
  NAND2_X1 U2887 ( .A1(n2766), .A2(n2885), .ZN(n2880) );
  NAND2_X1 U2888 ( .A1(n2765), .A2(n2767), .ZN(n2885) );
  NAND2_X1 U2889 ( .A1(n2886), .A2(n2887), .ZN(n2767) );
  NAND2_X1 U2890 ( .A1(b_8_), .A2(a_11_), .ZN(n2887) );
  INV_X1 U2891 ( .A(n2888), .ZN(n2886) );
  XNOR2_X1 U2892 ( .A(n2889), .B(n2890), .ZN(n2765) );
  XOR2_X1 U2893 ( .A(n2891), .B(n2892), .Z(n2890) );
  NAND2_X1 U2894 ( .A1(b_7_), .A2(a_12_), .ZN(n2892) );
  NAND2_X1 U2895 ( .A1(a_11_), .A2(n2888), .ZN(n2766) );
  NAND2_X1 U2896 ( .A1(n2893), .A2(n2894), .ZN(n2888) );
  NAND2_X1 U2897 ( .A1(n2895), .A2(a_12_), .ZN(n2894) );
  NOR2_X1 U2898 ( .A1(n2896), .A2(n2662), .ZN(n2895) );
  NOR2_X1 U2899 ( .A1(n2772), .A2(n2774), .ZN(n2896) );
  NAND2_X1 U2900 ( .A1(n2772), .A2(n2774), .ZN(n2893) );
  NAND2_X1 U2901 ( .A1(n2897), .A2(n2898), .ZN(n2774) );
  NAND2_X1 U2902 ( .A1(n2792), .A2(n2899), .ZN(n2898) );
  NAND2_X1 U2903 ( .A1(n2794), .A2(n2793), .ZN(n2899) );
  NOR2_X1 U2904 ( .A1(n2662), .A2(n1870), .ZN(n2792) );
  OR2_X1 U2905 ( .A1(n2793), .A2(n2794), .ZN(n2897) );
  AND2_X1 U2906 ( .A1(n2900), .A2(n2901), .ZN(n2794) );
  NAND2_X1 U2907 ( .A1(n2902), .A2(b_6_), .ZN(n2901) );
  NOR2_X1 U2908 ( .A1(n2903), .A2(n2071), .ZN(n2902) );
  NOR2_X1 U2909 ( .A1(n2070), .A2(n2789), .ZN(n2903) );
  NAND2_X1 U2910 ( .A1(n2904), .A2(b_7_), .ZN(n2900) );
  NOR2_X1 U2911 ( .A1(n2905), .A2(n2208), .ZN(n2904) );
  NOR2_X1 U2912 ( .A1(n2064), .A2(n2906), .ZN(n2905) );
  NAND2_X1 U2913 ( .A1(n2907), .A2(b_7_), .ZN(n2793) );
  NOR2_X1 U2914 ( .A1(n2210), .A2(n2662), .ZN(n2907) );
  XOR2_X1 U2915 ( .A(n2908), .B(n2909), .Z(n2772) );
  XOR2_X1 U2916 ( .A(n2910), .B(n2911), .Z(n2908) );
  XNOR2_X1 U2917 ( .A(n2912), .B(n2913), .ZN(n2799) );
  NAND2_X1 U2918 ( .A1(n2914), .A2(n2915), .ZN(n2912) );
  XNOR2_X1 U2919 ( .A(n2916), .B(n2917), .ZN(n2804) );
  XNOR2_X1 U2920 ( .A(n2918), .B(n2919), .ZN(n2917) );
  XOR2_X1 U2921 ( .A(n2920), .B(n2921), .Z(n2808) );
  XOR2_X1 U2922 ( .A(n2922), .B(n2923), .Z(n2920) );
  NOR2_X1 U2923 ( .A1(n2789), .A2(n2028), .ZN(n2923) );
  XOR2_X1 U2924 ( .A(n2924), .B(n2925), .Z(n2812) );
  XOR2_X1 U2925 ( .A(n2926), .B(n2927), .Z(n2924) );
  XOR2_X1 U2926 ( .A(n2928), .B(n2929), .Z(n2738) );
  XOR2_X1 U2927 ( .A(n2930), .B(n2931), .Z(n2928) );
  NOR2_X1 U2928 ( .A1(n2789), .A2(n2019), .ZN(n2931) );
  XNOR2_X1 U2929 ( .A(n2932), .B(n2933), .ZN(n2815) );
  XOR2_X1 U2930 ( .A(n2934), .B(n2935), .Z(n2933) );
  NAND2_X1 U2931 ( .A1(b_7_), .A2(a_5_), .ZN(n2935) );
  XNOR2_X1 U2932 ( .A(n2936), .B(n2937), .ZN(n2819) );
  XOR2_X1 U2933 ( .A(n2938), .B(n2939), .Z(n2937) );
  NAND2_X1 U2934 ( .A1(b_7_), .A2(a_4_), .ZN(n2939) );
  XNOR2_X1 U2935 ( .A(n2940), .B(n2941), .ZN(n2824) );
  XOR2_X1 U2936 ( .A(n2942), .B(n2943), .Z(n2941) );
  NAND2_X1 U2937 ( .A1(a_3_), .A2(b_7_), .ZN(n2943) );
  XNOR2_X1 U2938 ( .A(n2944), .B(n2945), .ZN(n2828) );
  XOR2_X1 U2939 ( .A(n2946), .B(n2947), .Z(n2945) );
  NAND2_X1 U2940 ( .A1(a_2_), .A2(b_7_), .ZN(n2947) );
  XNOR2_X1 U2941 ( .A(n2948), .B(n2949), .ZN(n2712) );
  XOR2_X1 U2942 ( .A(n2950), .B(n2951), .Z(n2949) );
  NAND2_X1 U2943 ( .A1(a_1_), .A2(b_7_), .ZN(n2951) );
  NAND2_X1 U2944 ( .A1(n2952), .A2(n2953), .ZN(n1840) );
  NAND2_X1 U2945 ( .A1(n2841), .A2(n2839), .ZN(n2953) );
  NAND2_X1 U2946 ( .A1(n2954), .A2(n2841), .ZN(n1841) );
  XNOR2_X1 U2947 ( .A(n2955), .B(n2956), .ZN(n2841) );
  XOR2_X1 U2948 ( .A(n2957), .B(n2958), .Z(n2956) );
  NAND2_X1 U2949 ( .A1(a_0_), .A2(b_6_), .ZN(n2958) );
  NOR2_X1 U2950 ( .A1(n2959), .A2(n2952), .ZN(n2954) );
  XNOR2_X1 U2951 ( .A(n2960), .B(n2961), .ZN(n2952) );
  INV_X1 U2952 ( .A(n2839), .ZN(n2959) );
  NAND2_X1 U2953 ( .A1(n2962), .A2(n2963), .ZN(n2839) );
  NAND2_X1 U2954 ( .A1(n2964), .A2(a_0_), .ZN(n2963) );
  NOR2_X1 U2955 ( .A1(n2965), .A2(n2789), .ZN(n2964) );
  NOR2_X1 U2956 ( .A1(n2836), .A2(n2834), .ZN(n2965) );
  NAND2_X1 U2957 ( .A1(n2834), .A2(n2836), .ZN(n2962) );
  NAND2_X1 U2958 ( .A1(n2966), .A2(n2967), .ZN(n2836) );
  NAND2_X1 U2959 ( .A1(n2968), .A2(a_1_), .ZN(n2967) );
  NOR2_X1 U2960 ( .A1(n2969), .A2(n2789), .ZN(n2968) );
  NOR2_X1 U2961 ( .A1(n2948), .A2(n2950), .ZN(n2969) );
  NAND2_X1 U2962 ( .A1(n2948), .A2(n2950), .ZN(n2966) );
  NAND2_X1 U2963 ( .A1(n2970), .A2(n2971), .ZN(n2950) );
  NAND2_X1 U2964 ( .A1(n2972), .A2(a_2_), .ZN(n2971) );
  NOR2_X1 U2965 ( .A1(n2973), .A2(n2789), .ZN(n2972) );
  NOR2_X1 U2966 ( .A1(n2944), .A2(n2946), .ZN(n2973) );
  NAND2_X1 U2967 ( .A1(n2944), .A2(n2946), .ZN(n2970) );
  NAND2_X1 U2968 ( .A1(n2974), .A2(n2975), .ZN(n2946) );
  NAND2_X1 U2969 ( .A1(n2976), .A2(a_3_), .ZN(n2975) );
  NOR2_X1 U2970 ( .A1(n2977), .A2(n2789), .ZN(n2976) );
  NOR2_X1 U2971 ( .A1(n2942), .A2(n2940), .ZN(n2977) );
  NAND2_X1 U2972 ( .A1(n2940), .A2(n2942), .ZN(n2974) );
  NAND2_X1 U2973 ( .A1(n2978), .A2(n2979), .ZN(n2942) );
  NAND2_X1 U2974 ( .A1(n2980), .A2(b_7_), .ZN(n2979) );
  NOR2_X1 U2975 ( .A1(n2981), .A2(n2009), .ZN(n2980) );
  NOR2_X1 U2976 ( .A1(n2936), .A2(n2938), .ZN(n2981) );
  NAND2_X1 U2977 ( .A1(n2936), .A2(n2938), .ZN(n2978) );
  NAND2_X1 U2978 ( .A1(n2982), .A2(n2983), .ZN(n2938) );
  NAND2_X1 U2979 ( .A1(n2984), .A2(b_7_), .ZN(n2983) );
  NOR2_X1 U2980 ( .A1(n2985), .A2(n2014), .ZN(n2984) );
  NOR2_X1 U2981 ( .A1(n2934), .A2(n2932), .ZN(n2985) );
  NAND2_X1 U2982 ( .A1(n2932), .A2(n2934), .ZN(n2982) );
  NAND2_X1 U2983 ( .A1(n2986), .A2(n2987), .ZN(n2934) );
  NAND2_X1 U2984 ( .A1(n2988), .A2(a_6_), .ZN(n2987) );
  NOR2_X1 U2985 ( .A1(n2989), .A2(n2789), .ZN(n2988) );
  NOR2_X1 U2986 ( .A1(n2929), .A2(n2930), .ZN(n2989) );
  NAND2_X1 U2987 ( .A1(n2929), .A2(n2930), .ZN(n2986) );
  NAND2_X1 U2988 ( .A1(n2990), .A2(n2991), .ZN(n2930) );
  NAND2_X1 U2989 ( .A1(n2925), .A2(n2992), .ZN(n2991) );
  OR2_X1 U2990 ( .A1(n2926), .A2(n2927), .ZN(n2992) );
  XOR2_X1 U2991 ( .A(n2993), .B(n2994), .Z(n2925) );
  XOR2_X1 U2992 ( .A(n2995), .B(n2996), .Z(n2993) );
  NAND2_X1 U2993 ( .A1(n2927), .A2(n2926), .ZN(n2990) );
  NAND2_X1 U2994 ( .A1(n2997), .A2(n2998), .ZN(n2926) );
  NAND2_X1 U2995 ( .A1(n2999), .A2(a_8_), .ZN(n2998) );
  NOR2_X1 U2996 ( .A1(n3000), .A2(n2789), .ZN(n2999) );
  NOR2_X1 U2997 ( .A1(n2921), .A2(n2922), .ZN(n3000) );
  NAND2_X1 U2998 ( .A1(n2921), .A2(n2922), .ZN(n2997) );
  NAND2_X1 U2999 ( .A1(n3001), .A2(n3002), .ZN(n2922) );
  NAND2_X1 U3000 ( .A1(n2919), .A2(n3003), .ZN(n3002) );
  OR2_X1 U3001 ( .A1(n2918), .A2(n2916), .ZN(n3003) );
  NOR2_X1 U3002 ( .A1(n2789), .A2(n2178), .ZN(n2919) );
  NAND2_X1 U3003 ( .A1(n2916), .A2(n2918), .ZN(n3001) );
  NAND2_X1 U3004 ( .A1(n2914), .A2(n3004), .ZN(n2918) );
  NAND2_X1 U3005 ( .A1(n2913), .A2(n2915), .ZN(n3004) );
  NAND2_X1 U3006 ( .A1(n3005), .A2(n3006), .ZN(n2915) );
  NAND2_X1 U3007 ( .A1(a_10_), .A2(b_7_), .ZN(n3006) );
  INV_X1 U3008 ( .A(n3007), .ZN(n3005) );
  XNOR2_X1 U3009 ( .A(n3008), .B(n3009), .ZN(n2913) );
  NAND2_X1 U3010 ( .A1(n3010), .A2(n3011), .ZN(n3008) );
  NAND2_X1 U3011 ( .A1(a_10_), .A2(n3007), .ZN(n2914) );
  NAND2_X1 U3012 ( .A1(n2883), .A2(n3012), .ZN(n3007) );
  NAND2_X1 U3013 ( .A1(n2882), .A2(n2884), .ZN(n3012) );
  NAND2_X1 U3014 ( .A1(n3013), .A2(n3014), .ZN(n2884) );
  NAND2_X1 U3015 ( .A1(b_7_), .A2(a_11_), .ZN(n3014) );
  INV_X1 U3016 ( .A(n3015), .ZN(n3013) );
  XNOR2_X1 U3017 ( .A(n3016), .B(n3017), .ZN(n2882) );
  XOR2_X1 U3018 ( .A(n3018), .B(n3019), .Z(n3017) );
  NAND2_X1 U3019 ( .A1(b_6_), .A2(a_12_), .ZN(n3019) );
  NAND2_X1 U3020 ( .A1(a_11_), .A2(n3015), .ZN(n2883) );
  NAND2_X1 U3021 ( .A1(n3020), .A2(n3021), .ZN(n3015) );
  NAND2_X1 U3022 ( .A1(n3022), .A2(b_7_), .ZN(n3021) );
  NOR2_X1 U3023 ( .A1(n3023), .A2(n2057), .ZN(n3022) );
  NOR2_X1 U3024 ( .A1(n2889), .A2(n2891), .ZN(n3023) );
  NAND2_X1 U3025 ( .A1(n2889), .A2(n2891), .ZN(n3020) );
  NAND2_X1 U3026 ( .A1(n3024), .A2(n3025), .ZN(n2891) );
  NAND2_X1 U3027 ( .A1(n2909), .A2(n3026), .ZN(n3025) );
  NAND2_X1 U3028 ( .A1(n2911), .A2(n2910), .ZN(n3026) );
  NOR2_X1 U3029 ( .A1(n2789), .A2(n1870), .ZN(n2909) );
  OR2_X1 U3030 ( .A1(n2910), .A2(n2911), .ZN(n3024) );
  AND2_X1 U3031 ( .A1(n3027), .A2(n3028), .ZN(n2911) );
  NAND2_X1 U3032 ( .A1(n3029), .A2(b_5_), .ZN(n3028) );
  NOR2_X1 U3033 ( .A1(n3030), .A2(n2071), .ZN(n3029) );
  NOR2_X1 U3034 ( .A1(n2070), .A2(n2906), .ZN(n3030) );
  NAND2_X1 U3035 ( .A1(n3031), .A2(b_6_), .ZN(n3027) );
  NOR2_X1 U3036 ( .A1(n3032), .A2(n2208), .ZN(n3031) );
  NOR2_X1 U3037 ( .A1(n2064), .A2(n3033), .ZN(n3032) );
  NAND2_X1 U3038 ( .A1(n3034), .A2(b_6_), .ZN(n2910) );
  NOR2_X1 U3039 ( .A1(n2210), .A2(n2789), .ZN(n3034) );
  XOR2_X1 U3040 ( .A(n3035), .B(n3036), .Z(n2889) );
  XOR2_X1 U3041 ( .A(n3037), .B(n3038), .Z(n3035) );
  XNOR2_X1 U3042 ( .A(n3039), .B(n3040), .ZN(n2916) );
  NAND2_X1 U3043 ( .A1(n3041), .A2(n3042), .ZN(n3039) );
  XNOR2_X1 U3044 ( .A(n3043), .B(n3044), .ZN(n2921) );
  NAND2_X1 U3045 ( .A1(n3045), .A2(n3046), .ZN(n3043) );
  XNOR2_X1 U3046 ( .A(n3047), .B(n3048), .ZN(n2929) );
  NAND2_X1 U3047 ( .A1(n3049), .A2(n3050), .ZN(n3047) );
  XOR2_X1 U3048 ( .A(n3051), .B(n3052), .Z(n2932) );
  XNOR2_X1 U3049 ( .A(n3053), .B(n3054), .ZN(n3051) );
  XNOR2_X1 U3050 ( .A(n3055), .B(n3056), .ZN(n2936) );
  NAND2_X1 U3051 ( .A1(n3057), .A2(n3058), .ZN(n3055) );
  XOR2_X1 U3052 ( .A(n3059), .B(n3060), .Z(n2940) );
  XOR2_X1 U3053 ( .A(n3061), .B(n3062), .Z(n3060) );
  XNOR2_X1 U3054 ( .A(n3063), .B(n3064), .ZN(n2944) );
  NAND2_X1 U3055 ( .A1(n3065), .A2(n3066), .ZN(n3063) );
  XOR2_X1 U3056 ( .A(n3067), .B(n3068), .Z(n2948) );
  XOR2_X1 U3057 ( .A(n3069), .B(n3070), .Z(n3067) );
  NOR2_X1 U3058 ( .A1(n2906), .A2(n2000), .ZN(n3070) );
  XNOR2_X1 U3059 ( .A(n3071), .B(n3072), .ZN(n2834) );
  XOR2_X1 U3060 ( .A(n3073), .B(n3074), .Z(n3072) );
  NAND2_X1 U3061 ( .A1(a_1_), .A2(b_6_), .ZN(n3074) );
  NAND2_X1 U3062 ( .A1(n3075), .A2(n3076), .ZN(n1844) );
  OR2_X1 U3063 ( .A1(n2961), .A2(n2960), .ZN(n3076) );
  XNOR2_X1 U3064 ( .A(n3077), .B(n3078), .ZN(n3075) );
  NAND2_X1 U3065 ( .A1(n3079), .A2(n3080), .ZN(n1845) );
  XOR2_X1 U3066 ( .A(n3077), .B(n3078), .Z(n3080) );
  NOR2_X1 U3067 ( .A1(n2960), .A2(n2961), .ZN(n3079) );
  XOR2_X1 U3068 ( .A(n3081), .B(n3082), .Z(n2961) );
  XOR2_X1 U3069 ( .A(n3083), .B(n3084), .Z(n3082) );
  NAND2_X1 U3070 ( .A1(a_0_), .A2(b_5_), .ZN(n3084) );
  AND2_X1 U3071 ( .A1(n3085), .A2(n3086), .ZN(n2960) );
  NAND2_X1 U3072 ( .A1(n3087), .A2(a_0_), .ZN(n3086) );
  NOR2_X1 U3073 ( .A1(n3088), .A2(n2906), .ZN(n3087) );
  NOR2_X1 U3074 ( .A1(n2957), .A2(n2955), .ZN(n3088) );
  NAND2_X1 U3075 ( .A1(n2955), .A2(n2957), .ZN(n3085) );
  NAND2_X1 U3076 ( .A1(n3089), .A2(n3090), .ZN(n2957) );
  NAND2_X1 U3077 ( .A1(n3091), .A2(a_1_), .ZN(n3090) );
  NOR2_X1 U3078 ( .A1(n3092), .A2(n2906), .ZN(n3091) );
  NOR2_X1 U3079 ( .A1(n3071), .A2(n3073), .ZN(n3092) );
  NAND2_X1 U3080 ( .A1(n3071), .A2(n3073), .ZN(n3089) );
  NAND2_X1 U3081 ( .A1(n3093), .A2(n3094), .ZN(n3073) );
  NAND2_X1 U3082 ( .A1(n3095), .A2(a_2_), .ZN(n3094) );
  NOR2_X1 U3083 ( .A1(n3096), .A2(n2906), .ZN(n3095) );
  NOR2_X1 U3084 ( .A1(n3069), .A2(n3068), .ZN(n3096) );
  NAND2_X1 U3085 ( .A1(n3068), .A2(n3069), .ZN(n3093) );
  NAND2_X1 U3086 ( .A1(n3065), .A2(n3097), .ZN(n3069) );
  NAND2_X1 U3087 ( .A1(n3064), .A2(n3066), .ZN(n3097) );
  NAND2_X1 U3088 ( .A1(n3098), .A2(n3099), .ZN(n3066) );
  NAND2_X1 U3089 ( .A1(a_3_), .A2(b_6_), .ZN(n3099) );
  INV_X1 U3090 ( .A(n3100), .ZN(n3098) );
  XOR2_X1 U3091 ( .A(n3101), .B(n3102), .Z(n3064) );
  XNOR2_X1 U3092 ( .A(n3103), .B(n3104), .ZN(n3101) );
  NAND2_X1 U3093 ( .A1(b_5_), .A2(a_4_), .ZN(n3103) );
  NAND2_X1 U3094 ( .A1(a_3_), .A2(n3100), .ZN(n3065) );
  NAND2_X1 U3095 ( .A1(n3105), .A2(n3106), .ZN(n3100) );
  NAND2_X1 U3096 ( .A1(n3062), .A2(n3107), .ZN(n3106) );
  NAND2_X1 U3097 ( .A1(n3061), .A2(n3059), .ZN(n3107) );
  NOR2_X1 U3098 ( .A1(n2906), .A2(n2009), .ZN(n3062) );
  OR2_X1 U3099 ( .A1(n3059), .A2(n3061), .ZN(n3105) );
  AND2_X1 U3100 ( .A1(n3057), .A2(n3108), .ZN(n3061) );
  NAND2_X1 U3101 ( .A1(n3056), .A2(n3058), .ZN(n3108) );
  NAND2_X1 U3102 ( .A1(n3109), .A2(n3110), .ZN(n3058) );
  NAND2_X1 U3103 ( .A1(b_6_), .A2(a_5_), .ZN(n3110) );
  XNOR2_X1 U3104 ( .A(n3111), .B(n3112), .ZN(n3056) );
  XOR2_X1 U3105 ( .A(n3113), .B(n3114), .Z(n3112) );
  NAND2_X1 U3106 ( .A1(a_6_), .A2(b_5_), .ZN(n3114) );
  OR2_X1 U3107 ( .A1(n3109), .A2(n2014), .ZN(n3057) );
  NAND2_X1 U3108 ( .A1(n3115), .A2(n3116), .ZN(n3109) );
  NAND2_X1 U3109 ( .A1(n3117), .A2(n3054), .ZN(n3116) );
  NAND2_X1 U3110 ( .A1(n3052), .A2(n3053), .ZN(n3117) );
  OR2_X1 U3111 ( .A1(n3053), .A2(n3052), .ZN(n3115) );
  XOR2_X1 U3112 ( .A(n3118), .B(n3119), .Z(n3052) );
  XOR2_X1 U3113 ( .A(n3120), .B(n3121), .Z(n3118) );
  NOR2_X1 U3114 ( .A1(n2170), .A2(n3033), .ZN(n3121) );
  NAND2_X1 U3115 ( .A1(n3049), .A2(n3122), .ZN(n3053) );
  NAND2_X1 U3116 ( .A1(n3048), .A2(n3050), .ZN(n3122) );
  NAND2_X1 U3117 ( .A1(n3123), .A2(n3124), .ZN(n3050) );
  NAND2_X1 U3118 ( .A1(b_6_), .A2(a_7_), .ZN(n3124) );
  INV_X1 U3119 ( .A(n3125), .ZN(n3123) );
  XOR2_X1 U3120 ( .A(n3126), .B(n3127), .Z(n3048) );
  XOR2_X1 U3121 ( .A(n3128), .B(n3129), .Z(n3126) );
  NOR2_X1 U3122 ( .A1(n3033), .A2(n2028), .ZN(n3129) );
  NAND2_X1 U3123 ( .A1(a_7_), .A2(n3125), .ZN(n3049) );
  NAND2_X1 U3124 ( .A1(n3130), .A2(n3131), .ZN(n3125) );
  NAND2_X1 U3125 ( .A1(n2996), .A2(n3132), .ZN(n3131) );
  OR2_X1 U3126 ( .A1(n2994), .A2(n2995), .ZN(n3132) );
  NOR2_X1 U3127 ( .A1(n2028), .A2(n2906), .ZN(n2996) );
  NAND2_X1 U3128 ( .A1(n2994), .A2(n2995), .ZN(n3130) );
  NAND2_X1 U3129 ( .A1(n3045), .A2(n3133), .ZN(n2995) );
  NAND2_X1 U3130 ( .A1(n3044), .A2(n3046), .ZN(n3133) );
  NAND2_X1 U3131 ( .A1(n3134), .A2(n3135), .ZN(n3046) );
  NAND2_X1 U3132 ( .A1(b_6_), .A2(a_9_), .ZN(n3135) );
  INV_X1 U3133 ( .A(n3136), .ZN(n3134) );
  XOR2_X1 U3134 ( .A(n3137), .B(n3138), .Z(n3044) );
  XOR2_X1 U3135 ( .A(n3139), .B(n3140), .Z(n3137) );
  NAND2_X1 U3136 ( .A1(a_9_), .A2(n3136), .ZN(n3045) );
  NAND2_X1 U3137 ( .A1(n3041), .A2(n3141), .ZN(n3136) );
  NAND2_X1 U3138 ( .A1(n3040), .A2(n3042), .ZN(n3141) );
  NAND2_X1 U3139 ( .A1(n3142), .A2(n3143), .ZN(n3042) );
  NAND2_X1 U3140 ( .A1(b_6_), .A2(a_10_), .ZN(n3143) );
  INV_X1 U3141 ( .A(n3144), .ZN(n3142) );
  XOR2_X1 U3142 ( .A(n3145), .B(n3146), .Z(n3040) );
  XOR2_X1 U3143 ( .A(n3147), .B(n3148), .Z(n3145) );
  NAND2_X1 U3144 ( .A1(a_10_), .A2(n3144), .ZN(n3041) );
  NAND2_X1 U3145 ( .A1(n3010), .A2(n3149), .ZN(n3144) );
  NAND2_X1 U3146 ( .A1(n3009), .A2(n3011), .ZN(n3149) );
  NAND2_X1 U3147 ( .A1(n3150), .A2(n3151), .ZN(n3011) );
  NAND2_X1 U3148 ( .A1(b_6_), .A2(a_11_), .ZN(n3151) );
  INV_X1 U3149 ( .A(n3152), .ZN(n3150) );
  XNOR2_X1 U3150 ( .A(n3153), .B(n3154), .ZN(n3009) );
  XOR2_X1 U3151 ( .A(n3155), .B(n3156), .Z(n3154) );
  NAND2_X1 U3152 ( .A1(b_5_), .A2(a_12_), .ZN(n3156) );
  NAND2_X1 U3153 ( .A1(a_11_), .A2(n3152), .ZN(n3010) );
  NAND2_X1 U3154 ( .A1(n3157), .A2(n3158), .ZN(n3152) );
  NAND2_X1 U3155 ( .A1(n3159), .A2(b_6_), .ZN(n3158) );
  NOR2_X1 U3156 ( .A1(n3160), .A2(n2057), .ZN(n3159) );
  NOR2_X1 U3157 ( .A1(n3016), .A2(n3018), .ZN(n3160) );
  NAND2_X1 U3158 ( .A1(n3016), .A2(n3018), .ZN(n3157) );
  NAND2_X1 U3159 ( .A1(n3161), .A2(n3162), .ZN(n3018) );
  NAND2_X1 U3160 ( .A1(n3036), .A2(n3163), .ZN(n3162) );
  NAND2_X1 U3161 ( .A1(n3038), .A2(n3037), .ZN(n3163) );
  NOR2_X1 U3162 ( .A1(n2906), .A2(n1870), .ZN(n3036) );
  OR2_X1 U3163 ( .A1(n3037), .A2(n3038), .ZN(n3161) );
  AND2_X1 U3164 ( .A1(n3164), .A2(n3165), .ZN(n3038) );
  NAND2_X1 U3165 ( .A1(n3166), .A2(b_4_), .ZN(n3165) );
  NOR2_X1 U3166 ( .A1(n3167), .A2(n2071), .ZN(n3166) );
  NOR2_X1 U3167 ( .A1(n2070), .A2(n3033), .ZN(n3167) );
  NAND2_X1 U3168 ( .A1(n3168), .A2(b_5_), .ZN(n3164) );
  NOR2_X1 U3169 ( .A1(n3169), .A2(n2208), .ZN(n3168) );
  NOR2_X1 U3170 ( .A1(n2064), .A2(n3170), .ZN(n3169) );
  NAND2_X1 U3171 ( .A1(n3171), .A2(b_5_), .ZN(n3037) );
  NOR2_X1 U3172 ( .A1(n2210), .A2(n2906), .ZN(n3171) );
  XOR2_X1 U3173 ( .A(n3172), .B(n3173), .Z(n3016) );
  XOR2_X1 U3174 ( .A(n3174), .B(n3175), .Z(n3172) );
  XNOR2_X1 U3175 ( .A(n3176), .B(n3177), .ZN(n2994) );
  NAND2_X1 U3176 ( .A1(n3178), .A2(n3179), .ZN(n3176) );
  XOR2_X1 U3177 ( .A(n3180), .B(n3181), .Z(n3059) );
  XNOR2_X1 U3178 ( .A(n3182), .B(n3183), .ZN(n3181) );
  XNOR2_X1 U3179 ( .A(n3184), .B(n3185), .ZN(n3068) );
  XOR2_X1 U3180 ( .A(n3186), .B(n3187), .Z(n3185) );
  NAND2_X1 U3181 ( .A1(a_3_), .A2(b_5_), .ZN(n3187) );
  XNOR2_X1 U3182 ( .A(n3188), .B(n3189), .ZN(n3071) );
  XOR2_X1 U3183 ( .A(n3190), .B(n3191), .Z(n3189) );
  NAND2_X1 U3184 ( .A1(a_2_), .A2(b_5_), .ZN(n3191) );
  XNOR2_X1 U3185 ( .A(n3192), .B(n3193), .ZN(n2955) );
  XOR2_X1 U3186 ( .A(n3194), .B(n3195), .Z(n3193) );
  NAND2_X1 U3187 ( .A1(a_1_), .A2(b_5_), .ZN(n3195) );
  NAND2_X1 U3188 ( .A1(n3196), .A2(n3197), .ZN(n1848) );
  NAND2_X1 U3189 ( .A1(n3078), .A2(n3077), .ZN(n3197) );
  XOR2_X1 U3190 ( .A(n3198), .B(n3199), .Z(n3196) );
  NAND2_X1 U3191 ( .A1(n3200), .A2(n3201), .ZN(n1849) );
  XOR2_X1 U3192 ( .A(n3202), .B(n3199), .Z(n3201) );
  AND2_X1 U3193 ( .A1(n3077), .A2(n3078), .ZN(n3200) );
  XOR2_X1 U3194 ( .A(n3203), .B(n3204), .Z(n3078) );
  XOR2_X1 U3195 ( .A(n3205), .B(n3206), .Z(n3203) );
  NOR2_X1 U3196 ( .A1(n3170), .A2(n1986), .ZN(n3206) );
  NAND2_X1 U3197 ( .A1(n3207), .A2(n3208), .ZN(n3077) );
  NAND2_X1 U3198 ( .A1(n3209), .A2(a_0_), .ZN(n3208) );
  NOR2_X1 U3199 ( .A1(n3210), .A2(n3033), .ZN(n3209) );
  NOR2_X1 U3200 ( .A1(n3083), .A2(n3081), .ZN(n3210) );
  NAND2_X1 U3201 ( .A1(n3081), .A2(n3083), .ZN(n3207) );
  NAND2_X1 U3202 ( .A1(n3211), .A2(n3212), .ZN(n3083) );
  NAND2_X1 U3203 ( .A1(n3213), .A2(a_1_), .ZN(n3212) );
  NOR2_X1 U3204 ( .A1(n3214), .A2(n3033), .ZN(n3213) );
  NOR2_X1 U3205 ( .A1(n3192), .A2(n3194), .ZN(n3214) );
  NAND2_X1 U3206 ( .A1(n3192), .A2(n3194), .ZN(n3211) );
  NAND2_X1 U3207 ( .A1(n3215), .A2(n3216), .ZN(n3194) );
  NAND2_X1 U3208 ( .A1(n3217), .A2(a_2_), .ZN(n3216) );
  NOR2_X1 U3209 ( .A1(n3218), .A2(n3033), .ZN(n3217) );
  NOR2_X1 U3210 ( .A1(n3190), .A2(n3188), .ZN(n3218) );
  NAND2_X1 U3211 ( .A1(n3188), .A2(n3190), .ZN(n3215) );
  NAND2_X1 U3212 ( .A1(n3219), .A2(n3220), .ZN(n3190) );
  NAND2_X1 U3213 ( .A1(n3221), .A2(a_3_), .ZN(n3220) );
  NOR2_X1 U3214 ( .A1(n3222), .A2(n3033), .ZN(n3221) );
  NOR2_X1 U3215 ( .A1(n3184), .A2(n3186), .ZN(n3222) );
  NAND2_X1 U3216 ( .A1(n3184), .A2(n3186), .ZN(n3219) );
  NAND2_X1 U3217 ( .A1(n3223), .A2(n3224), .ZN(n3186) );
  NAND2_X1 U3218 ( .A1(n3225), .A2(b_5_), .ZN(n3224) );
  NOR2_X1 U3219 ( .A1(n3226), .A2(n2009), .ZN(n3225) );
  NOR2_X1 U3220 ( .A1(n3104), .A2(n3102), .ZN(n3226) );
  NAND2_X1 U3221 ( .A1(n3102), .A2(n3104), .ZN(n3223) );
  NAND2_X1 U3222 ( .A1(n3227), .A2(n3228), .ZN(n3104) );
  NAND2_X1 U3223 ( .A1(n3180), .A2(n3229), .ZN(n3228) );
  OR2_X1 U3224 ( .A1(n3183), .A2(n3182), .ZN(n3229) );
  XNOR2_X1 U3225 ( .A(n3230), .B(n3231), .ZN(n3180) );
  XOR2_X1 U3226 ( .A(n3232), .B(n3233), .Z(n3231) );
  NAND2_X1 U3227 ( .A1(a_6_), .A2(b_4_), .ZN(n3233) );
  NAND2_X1 U3228 ( .A1(n3182), .A2(n3183), .ZN(n3227) );
  NAND2_X1 U3229 ( .A1(n3234), .A2(n3235), .ZN(n3183) );
  NAND2_X1 U3230 ( .A1(n3236), .A2(a_6_), .ZN(n3235) );
  NOR2_X1 U3231 ( .A1(n3237), .A2(n3033), .ZN(n3236) );
  NOR2_X1 U3232 ( .A1(n3113), .A2(n3111), .ZN(n3237) );
  NAND2_X1 U3233 ( .A1(n3111), .A2(n3113), .ZN(n3234) );
  NAND2_X1 U3234 ( .A1(n3238), .A2(n3239), .ZN(n3113) );
  NAND2_X1 U3235 ( .A1(n3240), .A2(b_5_), .ZN(n3239) );
  NOR2_X1 U3236 ( .A1(n3241), .A2(n2170), .ZN(n3240) );
  NOR2_X1 U3237 ( .A1(n3120), .A2(n3119), .ZN(n3241) );
  NAND2_X1 U3238 ( .A1(n3119), .A2(n3120), .ZN(n3238) );
  NAND2_X1 U3239 ( .A1(n3242), .A2(n3243), .ZN(n3120) );
  NAND2_X1 U3240 ( .A1(n3244), .A2(a_8_), .ZN(n3243) );
  NOR2_X1 U3241 ( .A1(n3245), .A2(n3033), .ZN(n3244) );
  NOR2_X1 U3242 ( .A1(n3128), .A2(n3127), .ZN(n3245) );
  NAND2_X1 U3243 ( .A1(n3127), .A2(n3128), .ZN(n3242) );
  NAND2_X1 U3244 ( .A1(n3178), .A2(n3246), .ZN(n3128) );
  NAND2_X1 U3245 ( .A1(n3177), .A2(n3179), .ZN(n3246) );
  NAND2_X1 U3246 ( .A1(n3247), .A2(n3248), .ZN(n3179) );
  NAND2_X1 U3247 ( .A1(b_5_), .A2(a_9_), .ZN(n3248) );
  INV_X1 U3248 ( .A(n3249), .ZN(n3247) );
  XNOR2_X1 U3249 ( .A(n3250), .B(n3251), .ZN(n3177) );
  XNOR2_X1 U3250 ( .A(n3252), .B(n3253), .ZN(n3250) );
  NAND2_X1 U3251 ( .A1(a_9_), .A2(n3249), .ZN(n3178) );
  NAND2_X1 U3252 ( .A1(n3254), .A2(n3255), .ZN(n3249) );
  NAND2_X1 U3253 ( .A1(n3140), .A2(n3256), .ZN(n3255) );
  OR2_X1 U3254 ( .A1(n3138), .A2(n3139), .ZN(n3256) );
  NOR2_X1 U3255 ( .A1(n3033), .A2(n1885), .ZN(n3140) );
  NAND2_X1 U3256 ( .A1(n3138), .A2(n3139), .ZN(n3254) );
  NAND2_X1 U3257 ( .A1(n3257), .A2(n3258), .ZN(n3139) );
  NAND2_X1 U3258 ( .A1(n3148), .A2(n3259), .ZN(n3258) );
  OR2_X1 U3259 ( .A1(n3146), .A2(n3147), .ZN(n3259) );
  NOR2_X1 U3260 ( .A1(n3033), .A2(n3260), .ZN(n3148) );
  NAND2_X1 U3261 ( .A1(n3146), .A2(n3147), .ZN(n3257) );
  NAND2_X1 U3262 ( .A1(n3261), .A2(n3262), .ZN(n3147) );
  NAND2_X1 U3263 ( .A1(n3263), .A2(b_5_), .ZN(n3262) );
  NOR2_X1 U3264 ( .A1(n3264), .A2(n2057), .ZN(n3263) );
  NOR2_X1 U3265 ( .A1(n3153), .A2(n3155), .ZN(n3264) );
  NAND2_X1 U3266 ( .A1(n3153), .A2(n3155), .ZN(n3261) );
  NAND2_X1 U3267 ( .A1(n3265), .A2(n3266), .ZN(n3155) );
  NAND2_X1 U3268 ( .A1(n3173), .A2(n3267), .ZN(n3266) );
  NAND2_X1 U3269 ( .A1(n3175), .A2(n3174), .ZN(n3267) );
  NOR2_X1 U3270 ( .A1(n3033), .A2(n1870), .ZN(n3173) );
  OR2_X1 U3271 ( .A1(n3174), .A2(n3175), .ZN(n3265) );
  AND2_X1 U3272 ( .A1(n3268), .A2(n3269), .ZN(n3175) );
  NAND2_X1 U3273 ( .A1(n3270), .A2(b_3_), .ZN(n3269) );
  NOR2_X1 U3274 ( .A1(n3271), .A2(n2071), .ZN(n3270) );
  NOR2_X1 U3275 ( .A1(n2070), .A2(n3170), .ZN(n3271) );
  NAND2_X1 U3276 ( .A1(n3272), .A2(b_4_), .ZN(n3268) );
  NOR2_X1 U3277 ( .A1(n3273), .A2(n2208), .ZN(n3272) );
  NOR2_X1 U3278 ( .A1(n2064), .A2(n3274), .ZN(n3273) );
  NAND2_X1 U3279 ( .A1(n3275), .A2(b_4_), .ZN(n3174) );
  NOR2_X1 U3280 ( .A1(n2210), .A2(n3033), .ZN(n3275) );
  XOR2_X1 U3281 ( .A(n3276), .B(n3277), .Z(n3153) );
  XOR2_X1 U3282 ( .A(n3278), .B(n3279), .Z(n3276) );
  XNOR2_X1 U3283 ( .A(n3280), .B(n3281), .ZN(n3146) );
  XOR2_X1 U3284 ( .A(n3282), .B(n3283), .Z(n3281) );
  NAND2_X1 U3285 ( .A1(b_4_), .A2(a_12_), .ZN(n3283) );
  XNOR2_X1 U3286 ( .A(n3284), .B(n3285), .ZN(n3138) );
  NAND2_X1 U3287 ( .A1(n3286), .A2(n3287), .ZN(n3284) );
  XNOR2_X1 U3288 ( .A(n3288), .B(n3289), .ZN(n3127) );
  NAND2_X1 U3289 ( .A1(n3290), .A2(n3291), .ZN(n3288) );
  XOR2_X1 U3290 ( .A(n3292), .B(n3293), .Z(n3119) );
  XOR2_X1 U3291 ( .A(n3294), .B(n3295), .Z(n3292) );
  NOR2_X1 U3292 ( .A1(n3170), .A2(n2028), .ZN(n3295) );
  XNOR2_X1 U3293 ( .A(n3296), .B(n3297), .ZN(n3111) );
  XOR2_X1 U3294 ( .A(n3298), .B(n3299), .Z(n3297) );
  NAND2_X1 U3295 ( .A1(b_4_), .A2(a_7_), .ZN(n3299) );
  XNOR2_X1 U3296 ( .A(n3300), .B(n3301), .ZN(n3102) );
  XOR2_X1 U3297 ( .A(n3302), .B(n3303), .Z(n3301) );
  NAND2_X1 U3298 ( .A1(b_4_), .A2(a_5_), .ZN(n3303) );
  XNOR2_X1 U3299 ( .A(n3304), .B(n3305), .ZN(n3184) );
  XNOR2_X1 U3300 ( .A(n3306), .B(n3307), .ZN(n3305) );
  XOR2_X1 U3301 ( .A(n3308), .B(n3309), .Z(n3188) );
  XNOR2_X1 U3302 ( .A(n3310), .B(n3311), .ZN(n3308) );
  NAND2_X1 U3303 ( .A1(a_3_), .A2(b_4_), .ZN(n3310) );
  XOR2_X1 U3304 ( .A(n3312), .B(n3313), .Z(n3192) );
  XNOR2_X1 U3305 ( .A(n3314), .B(n3315), .ZN(n3312) );
  NAND2_X1 U3306 ( .A1(a_2_), .A2(b_4_), .ZN(n3314) );
  XOR2_X1 U3307 ( .A(n3316), .B(n3317), .Z(n3081) );
  XOR2_X1 U3308 ( .A(n3318), .B(n3319), .Z(n3316) );
  NOR2_X1 U3309 ( .A1(n3170), .A2(n1995), .ZN(n3319) );
  NAND2_X1 U3310 ( .A1(n3320), .A2(n3321), .ZN(n1852) );
  NAND2_X1 U3311 ( .A1(n3199), .A2(n3202), .ZN(n3321) );
  NAND2_X1 U3312 ( .A1(n3322), .A2(n3199), .ZN(n1853) );
  XOR2_X1 U3313 ( .A(n3323), .B(n3324), .Z(n3199) );
  XOR2_X1 U3314 ( .A(n3325), .B(n3326), .Z(n3323) );
  NOR2_X1 U3315 ( .A1(n3274), .A2(n1986), .ZN(n3326) );
  NOR2_X1 U3316 ( .A1(n3198), .A2(n3320), .ZN(n3322) );
  XNOR2_X1 U3317 ( .A(n3327), .B(n3328), .ZN(n3320) );
  INV_X1 U3318 ( .A(n3202), .ZN(n3198) );
  NAND2_X1 U3319 ( .A1(n3329), .A2(n3330), .ZN(n3202) );
  NAND2_X1 U3320 ( .A1(n3331), .A2(a_0_), .ZN(n3330) );
  NOR2_X1 U3321 ( .A1(n3332), .A2(n3170), .ZN(n3331) );
  NOR2_X1 U3322 ( .A1(n3204), .A2(n3205), .ZN(n3332) );
  NAND2_X1 U3323 ( .A1(n3204), .A2(n3205), .ZN(n3329) );
  NAND2_X1 U3324 ( .A1(n3333), .A2(n3334), .ZN(n3205) );
  NAND2_X1 U3325 ( .A1(n3335), .A2(a_1_), .ZN(n3334) );
  NOR2_X1 U3326 ( .A1(n3336), .A2(n3170), .ZN(n3335) );
  NOR2_X1 U3327 ( .A1(n3317), .A2(n3318), .ZN(n3336) );
  NAND2_X1 U3328 ( .A1(n3317), .A2(n3318), .ZN(n3333) );
  NAND2_X1 U3329 ( .A1(n3337), .A2(n3338), .ZN(n3318) );
  NAND2_X1 U3330 ( .A1(n3339), .A2(a_2_), .ZN(n3338) );
  NOR2_X1 U3331 ( .A1(n3340), .A2(n3170), .ZN(n3339) );
  NOR2_X1 U3332 ( .A1(n3315), .A2(n3313), .ZN(n3340) );
  NAND2_X1 U3333 ( .A1(n3313), .A2(n3315), .ZN(n3337) );
  NAND2_X1 U3334 ( .A1(n3341), .A2(n3342), .ZN(n3315) );
  NAND2_X1 U3335 ( .A1(n3343), .A2(a_3_), .ZN(n3342) );
  NOR2_X1 U3336 ( .A1(n3344), .A2(n3170), .ZN(n3343) );
  NOR2_X1 U3337 ( .A1(n3309), .A2(n3311), .ZN(n3344) );
  NAND2_X1 U3338 ( .A1(n3309), .A2(n3311), .ZN(n3341) );
  NAND2_X1 U3339 ( .A1(n3345), .A2(n3346), .ZN(n3311) );
  NAND2_X1 U3340 ( .A1(n3306), .A2(n3347), .ZN(n3346) );
  OR2_X1 U3341 ( .A1(n3304), .A2(n3307), .ZN(n3347) );
  NAND2_X1 U3342 ( .A1(n3304), .A2(n3307), .ZN(n3345) );
  NAND2_X1 U3343 ( .A1(n3348), .A2(n3349), .ZN(n3307) );
  NAND2_X1 U3344 ( .A1(n3350), .A2(b_4_), .ZN(n3349) );
  NOR2_X1 U3345 ( .A1(n3351), .A2(n2014), .ZN(n3350) );
  NOR2_X1 U3346 ( .A1(n3300), .A2(n3302), .ZN(n3351) );
  NAND2_X1 U3347 ( .A1(n3300), .A2(n3302), .ZN(n3348) );
  NAND2_X1 U3348 ( .A1(n3352), .A2(n3353), .ZN(n3302) );
  NAND2_X1 U3349 ( .A1(n3354), .A2(a_6_), .ZN(n3353) );
  NOR2_X1 U3350 ( .A1(n3355), .A2(n3170), .ZN(n3354) );
  NOR2_X1 U3351 ( .A1(n3230), .A2(n3232), .ZN(n3355) );
  NAND2_X1 U3352 ( .A1(n3230), .A2(n3232), .ZN(n3352) );
  NAND2_X1 U3353 ( .A1(n3356), .A2(n3357), .ZN(n3232) );
  NAND2_X1 U3354 ( .A1(n3358), .A2(b_4_), .ZN(n3357) );
  NOR2_X1 U3355 ( .A1(n3359), .A2(n2170), .ZN(n3358) );
  NOR2_X1 U3356 ( .A1(n3296), .A2(n3298), .ZN(n3359) );
  NAND2_X1 U3357 ( .A1(n3296), .A2(n3298), .ZN(n3356) );
  NAND2_X1 U3358 ( .A1(n3360), .A2(n3361), .ZN(n3298) );
  NAND2_X1 U3359 ( .A1(n3362), .A2(a_8_), .ZN(n3361) );
  NOR2_X1 U3360 ( .A1(n3363), .A2(n3170), .ZN(n3362) );
  NOR2_X1 U3361 ( .A1(n3293), .A2(n3294), .ZN(n3363) );
  NAND2_X1 U3362 ( .A1(n3293), .A2(n3294), .ZN(n3360) );
  NAND2_X1 U3363 ( .A1(n3290), .A2(n3364), .ZN(n3294) );
  NAND2_X1 U3364 ( .A1(n3289), .A2(n3291), .ZN(n3364) );
  NAND2_X1 U3365 ( .A1(n3365), .A2(n3366), .ZN(n3291) );
  NAND2_X1 U3366 ( .A1(b_4_), .A2(a_9_), .ZN(n3366) );
  INV_X1 U3367 ( .A(n3367), .ZN(n3365) );
  XNOR2_X1 U3368 ( .A(n3368), .B(n3369), .ZN(n3289) );
  NAND2_X1 U3369 ( .A1(n3370), .A2(n3371), .ZN(n3368) );
  NAND2_X1 U3370 ( .A1(a_9_), .A2(n3367), .ZN(n3290) );
  NAND2_X1 U3371 ( .A1(n3372), .A2(n3373), .ZN(n3367) );
  NAND2_X1 U3372 ( .A1(n3253), .A2(n3374), .ZN(n3373) );
  NAND2_X1 U3373 ( .A1(n3252), .A2(n3251), .ZN(n3374) );
  NOR2_X1 U3374 ( .A1(n3170), .A2(n1885), .ZN(n3253) );
  OR2_X1 U3375 ( .A1(n3251), .A2(n3252), .ZN(n3372) );
  AND2_X1 U3376 ( .A1(n3286), .A2(n3375), .ZN(n3252) );
  NAND2_X1 U3377 ( .A1(n3285), .A2(n3287), .ZN(n3375) );
  NAND2_X1 U3378 ( .A1(n3376), .A2(n3377), .ZN(n3287) );
  NAND2_X1 U3379 ( .A1(b_4_), .A2(a_11_), .ZN(n3377) );
  INV_X1 U3380 ( .A(n3378), .ZN(n3376) );
  XNOR2_X1 U3381 ( .A(n3379), .B(n3380), .ZN(n3285) );
  XNOR2_X1 U3382 ( .A(n3381), .B(n3382), .ZN(n3379) );
  NAND2_X1 U3383 ( .A1(a_11_), .A2(n3378), .ZN(n3286) );
  NAND2_X1 U3384 ( .A1(n3383), .A2(n3384), .ZN(n3378) );
  NAND2_X1 U3385 ( .A1(n3385), .A2(b_4_), .ZN(n3384) );
  NOR2_X1 U3386 ( .A1(n3386), .A2(n2057), .ZN(n3385) );
  NOR2_X1 U3387 ( .A1(n3280), .A2(n3282), .ZN(n3386) );
  NAND2_X1 U3388 ( .A1(n3280), .A2(n3282), .ZN(n3383) );
  NAND2_X1 U3389 ( .A1(n3387), .A2(n3388), .ZN(n3282) );
  NAND2_X1 U3390 ( .A1(n3277), .A2(n3389), .ZN(n3388) );
  NAND2_X1 U3391 ( .A1(n3279), .A2(n3278), .ZN(n3389) );
  NOR2_X1 U3392 ( .A1(n3170), .A2(n1870), .ZN(n3277) );
  OR2_X1 U3393 ( .A1(n3278), .A2(n3279), .ZN(n3387) );
  AND2_X1 U3394 ( .A1(n3390), .A2(n3391), .ZN(n3279) );
  NAND2_X1 U3395 ( .A1(n3392), .A2(b_2_), .ZN(n3391) );
  NOR2_X1 U3396 ( .A1(n3393), .A2(n2071), .ZN(n3392) );
  NOR2_X1 U3397 ( .A1(n2070), .A2(n3274), .ZN(n3393) );
  NAND2_X1 U3398 ( .A1(n3394), .A2(b_3_), .ZN(n3390) );
  NOR2_X1 U3399 ( .A1(n3395), .A2(n2208), .ZN(n3394) );
  NOR2_X1 U3400 ( .A1(n2064), .A2(n3396), .ZN(n3395) );
  NAND2_X1 U3401 ( .A1(n3397), .A2(b_3_), .ZN(n3278) );
  NOR2_X1 U3402 ( .A1(n2210), .A2(n3170), .ZN(n3397) );
  XOR2_X1 U3403 ( .A(n3398), .B(n3399), .Z(n3280) );
  NOR2_X1 U3404 ( .A1(n1870), .A2(n3274), .ZN(n3399) );
  XOR2_X1 U3405 ( .A(n3400), .B(n3401), .Z(n3398) );
  XOR2_X1 U3406 ( .A(n3402), .B(n3403), .Z(n3251) );
  NAND2_X1 U3407 ( .A1(n3404), .A2(n3405), .ZN(n3402) );
  XNOR2_X1 U3408 ( .A(n3406), .B(n3407), .ZN(n3293) );
  NAND2_X1 U3409 ( .A1(n3408), .A2(n3409), .ZN(n3406) );
  XOR2_X1 U3410 ( .A(n3410), .B(n3411), .Z(n3296) );
  XOR2_X1 U3411 ( .A(n3412), .B(n3413), .Z(n3410) );
  NOR2_X1 U3412 ( .A1(n2028), .A2(n3274), .ZN(n3413) );
  XNOR2_X1 U3413 ( .A(n3414), .B(n3415), .ZN(n3230) );
  NAND2_X1 U3414 ( .A1(n3416), .A2(n3417), .ZN(n3414) );
  XOR2_X1 U3415 ( .A(n3418), .B(n3419), .Z(n3300) );
  XOR2_X1 U3416 ( .A(n3420), .B(n3421), .Z(n3418) );
  NOR2_X1 U3417 ( .A1(n3274), .A2(n2019), .ZN(n3421) );
  XOR2_X1 U3418 ( .A(n3422), .B(n3423), .Z(n3304) );
  XOR2_X1 U3419 ( .A(n3424), .B(n3425), .Z(n3422) );
  NOR2_X1 U3420 ( .A1(n2014), .A2(n3274), .ZN(n3425) );
  XOR2_X1 U3421 ( .A(n3426), .B(n3427), .Z(n3309) );
  XOR2_X1 U3422 ( .A(n3428), .B(n3429), .Z(n3426) );
  NOR2_X1 U3423 ( .A1(n2009), .A2(n3274), .ZN(n3429) );
  XOR2_X1 U3424 ( .A(n3430), .B(n3431), .Z(n3313) );
  XOR2_X1 U3425 ( .A(n3432), .B(n3433), .Z(n3430) );
  XOR2_X1 U3426 ( .A(n3434), .B(n3435), .Z(n3317) );
  XNOR2_X1 U3427 ( .A(n3436), .B(n3437), .ZN(n3434) );
  NAND2_X1 U3428 ( .A1(a_2_), .A2(b_3_), .ZN(n3436) );
  XOR2_X1 U3429 ( .A(n3438), .B(n3439), .Z(n3204) );
  XOR2_X1 U3430 ( .A(n3440), .B(n3441), .Z(n3438) );
  NOR2_X1 U3431 ( .A1(n3274), .A2(n1995), .ZN(n3441) );
  NAND2_X1 U3432 ( .A1(n3442), .A2(n3443), .ZN(n1866) );
  OR2_X1 U3433 ( .A1(n3328), .A2(n3327), .ZN(n3443) );
  XNOR2_X1 U3434 ( .A(n3444), .B(n3445), .ZN(n3442) );
  NAND2_X1 U3435 ( .A1(n3446), .A2(n3447), .ZN(n1867) );
  NOR2_X1 U3436 ( .A1(n3448), .A2(n3327), .ZN(n3447) );
  AND2_X1 U3437 ( .A1(n3449), .A2(n3450), .ZN(n3327) );
  NAND2_X1 U3438 ( .A1(n3451), .A2(a_0_), .ZN(n3450) );
  NOR2_X1 U3439 ( .A1(n3452), .A2(n3274), .ZN(n3451) );
  NOR2_X1 U3440 ( .A1(n3325), .A2(n3324), .ZN(n3452) );
  NAND2_X1 U3441 ( .A1(n3324), .A2(n3325), .ZN(n3449) );
  NAND2_X1 U3442 ( .A1(n3453), .A2(n3454), .ZN(n3325) );
  NAND2_X1 U3443 ( .A1(n3455), .A2(a_1_), .ZN(n3454) );
  NOR2_X1 U3444 ( .A1(n3456), .A2(n3274), .ZN(n3455) );
  NOR2_X1 U3445 ( .A1(n3440), .A2(n3439), .ZN(n3456) );
  NAND2_X1 U3446 ( .A1(n3439), .A2(n3440), .ZN(n3453) );
  NAND2_X1 U3447 ( .A1(n3457), .A2(n3458), .ZN(n3440) );
  NAND2_X1 U3448 ( .A1(n3459), .A2(a_2_), .ZN(n3458) );
  NOR2_X1 U3449 ( .A1(n3460), .A2(n3274), .ZN(n3459) );
  NOR2_X1 U3450 ( .A1(n3437), .A2(n3435), .ZN(n3460) );
  NAND2_X1 U3451 ( .A1(n3435), .A2(n3437), .ZN(n3457) );
  NAND2_X1 U3452 ( .A1(n3461), .A2(n3462), .ZN(n3437) );
  NAND2_X1 U3453 ( .A1(n3431), .A2(n3463), .ZN(n3462) );
  OR2_X1 U3454 ( .A1(n3432), .A2(n3433), .ZN(n3463) );
  XNOR2_X1 U3455 ( .A(n3464), .B(n3465), .ZN(n3431) );
  NAND2_X1 U3456 ( .A1(n3466), .A2(n3467), .ZN(n3464) );
  NAND2_X1 U3457 ( .A1(n3433), .A2(n3432), .ZN(n3461) );
  NAND2_X1 U3458 ( .A1(n3468), .A2(n3469), .ZN(n3432) );
  NAND2_X1 U3459 ( .A1(n3470), .A2(b_3_), .ZN(n3469) );
  NOR2_X1 U3460 ( .A1(n3471), .A2(n2009), .ZN(n3470) );
  NOR2_X1 U3461 ( .A1(n3428), .A2(n3427), .ZN(n3471) );
  NAND2_X1 U3462 ( .A1(n3427), .A2(n3428), .ZN(n3468) );
  NAND2_X1 U3463 ( .A1(n3472), .A2(n3473), .ZN(n3428) );
  NAND2_X1 U3464 ( .A1(n3474), .A2(b_3_), .ZN(n3473) );
  NOR2_X1 U3465 ( .A1(n3475), .A2(n2014), .ZN(n3474) );
  NOR2_X1 U3466 ( .A1(n3423), .A2(n3424), .ZN(n3475) );
  NAND2_X1 U3467 ( .A1(n3423), .A2(n3424), .ZN(n3472) );
  NAND2_X1 U3468 ( .A1(n3476), .A2(n3477), .ZN(n3424) );
  NAND2_X1 U3469 ( .A1(n3478), .A2(a_6_), .ZN(n3477) );
  NOR2_X1 U3470 ( .A1(n3479), .A2(n3274), .ZN(n3478) );
  NOR2_X1 U3471 ( .A1(n3420), .A2(n3419), .ZN(n3479) );
  NAND2_X1 U3472 ( .A1(n3419), .A2(n3420), .ZN(n3476) );
  NAND2_X1 U3473 ( .A1(n3416), .A2(n3480), .ZN(n3420) );
  NAND2_X1 U3474 ( .A1(n3415), .A2(n3417), .ZN(n3480) );
  NAND2_X1 U3475 ( .A1(n3481), .A2(n3482), .ZN(n3417) );
  NAND2_X1 U3476 ( .A1(b_3_), .A2(a_7_), .ZN(n3482) );
  INV_X1 U3477 ( .A(n3483), .ZN(n3481) );
  XNOR2_X1 U3478 ( .A(n3484), .B(n3485), .ZN(n3415) );
  NAND2_X1 U3479 ( .A1(n3486), .A2(n3487), .ZN(n3484) );
  NAND2_X1 U3480 ( .A1(a_7_), .A2(n3483), .ZN(n3416) );
  NAND2_X1 U3481 ( .A1(n3488), .A2(n3489), .ZN(n3483) );
  NAND2_X1 U3482 ( .A1(n3490), .A2(b_3_), .ZN(n3489) );
  NOR2_X1 U3483 ( .A1(n3491), .A2(n2028), .ZN(n3490) );
  NOR2_X1 U3484 ( .A1(n3412), .A2(n3411), .ZN(n3491) );
  NAND2_X1 U3485 ( .A1(n3411), .A2(n3412), .ZN(n3488) );
  NAND2_X1 U3486 ( .A1(n3408), .A2(n3492), .ZN(n3412) );
  NAND2_X1 U3487 ( .A1(n3407), .A2(n3409), .ZN(n3492) );
  NAND2_X1 U3488 ( .A1(n3493), .A2(n3494), .ZN(n3409) );
  NAND2_X1 U3489 ( .A1(b_3_), .A2(a_9_), .ZN(n3494) );
  INV_X1 U3490 ( .A(n3495), .ZN(n3493) );
  XNOR2_X1 U3491 ( .A(n3496), .B(n3497), .ZN(n3407) );
  NAND2_X1 U3492 ( .A1(n3498), .A2(n3499), .ZN(n3496) );
  NAND2_X1 U3493 ( .A1(a_9_), .A2(n3495), .ZN(n3408) );
  NAND2_X1 U3494 ( .A1(n3370), .A2(n3500), .ZN(n3495) );
  NAND2_X1 U3495 ( .A1(n3369), .A2(n3371), .ZN(n3500) );
  NAND2_X1 U3496 ( .A1(n3501), .A2(n3502), .ZN(n3371) );
  NAND2_X1 U3497 ( .A1(b_3_), .A2(a_10_), .ZN(n3502) );
  INV_X1 U3498 ( .A(n3503), .ZN(n3501) );
  XNOR2_X1 U3499 ( .A(n3504), .B(n3505), .ZN(n3369) );
  XNOR2_X1 U3500 ( .A(n3506), .B(n3507), .ZN(n3505) );
  NAND2_X1 U3501 ( .A1(a_10_), .A2(n3503), .ZN(n3370) );
  NAND2_X1 U3502 ( .A1(n3404), .A2(n3508), .ZN(n3503) );
  NAND2_X1 U3503 ( .A1(n3403), .A2(n3405), .ZN(n3508) );
  NAND2_X1 U3504 ( .A1(n3509), .A2(n3510), .ZN(n3405) );
  NAND2_X1 U3505 ( .A1(b_3_), .A2(a_11_), .ZN(n3510) );
  INV_X1 U3506 ( .A(n3511), .ZN(n3509) );
  XNOR2_X1 U3507 ( .A(n3512), .B(n3513), .ZN(n3403) );
  XNOR2_X1 U3508 ( .A(n3514), .B(n3515), .ZN(n3512) );
  NAND2_X1 U3509 ( .A1(a_11_), .A2(n3511), .ZN(n3404) );
  NAND2_X1 U3510 ( .A1(n3516), .A2(n3517), .ZN(n3511) );
  NAND2_X1 U3511 ( .A1(n3381), .A2(n3518), .ZN(n3517) );
  NAND2_X1 U3512 ( .A1(n3382), .A2(n3380), .ZN(n3518) );
  NOR2_X1 U3513 ( .A1(n3274), .A2(n2057), .ZN(n3381) );
  OR2_X1 U3514 ( .A1(n3380), .A2(n3382), .ZN(n3516) );
  AND2_X1 U3515 ( .A1(n3519), .A2(n3520), .ZN(n3382) );
  NAND2_X1 U3516 ( .A1(n3521), .A2(b_3_), .ZN(n3520) );
  NOR2_X1 U3517 ( .A1(n3522), .A2(n1870), .ZN(n3521) );
  NOR2_X1 U3518 ( .A1(n3400), .A2(n3401), .ZN(n3522) );
  NAND2_X1 U3519 ( .A1(n3400), .A2(n3401), .ZN(n3519) );
  NAND2_X1 U3520 ( .A1(n3523), .A2(n3524), .ZN(n3401) );
  NAND2_X1 U3521 ( .A1(n3525), .A2(b_1_), .ZN(n3524) );
  NOR2_X1 U3522 ( .A1(n3526), .A2(n2071), .ZN(n3525) );
  NOR2_X1 U3523 ( .A1(n2070), .A2(n3396), .ZN(n3526) );
  NAND2_X1 U3524 ( .A1(n3527), .A2(b_2_), .ZN(n3523) );
  NOR2_X1 U3525 ( .A1(n3528), .A2(n2208), .ZN(n3527) );
  NOR2_X1 U3526 ( .A1(n2064), .A2(n3529), .ZN(n3528) );
  AND2_X1 U3527 ( .A1(n3530), .A2(b_2_), .ZN(n3400) );
  NOR2_X1 U3528 ( .A1(n2210), .A2(n3274), .ZN(n3530) );
  XNOR2_X1 U3529 ( .A(n3531), .B(n3532), .ZN(n3380) );
  NOR2_X1 U3530 ( .A1(n1870), .A2(n3396), .ZN(n3532) );
  XOR2_X1 U3531 ( .A(n3533), .B(n3534), .Z(n3531) );
  XNOR2_X1 U3532 ( .A(n3535), .B(n3536), .ZN(n3411) );
  XNOR2_X1 U3533 ( .A(n3537), .B(n3538), .ZN(n3535) );
  XNOR2_X1 U3534 ( .A(n3539), .B(n3540), .ZN(n3419) );
  XNOR2_X1 U3535 ( .A(n3541), .B(n3542), .ZN(n3539) );
  XNOR2_X1 U3536 ( .A(n3543), .B(n3544), .ZN(n3423) );
  NAND2_X1 U3537 ( .A1(n3545), .A2(n3546), .ZN(n3543) );
  XNOR2_X1 U3538 ( .A(n3547), .B(n3548), .ZN(n3427) );
  XNOR2_X1 U3539 ( .A(n3549), .B(n3550), .ZN(n3547) );
  XNOR2_X1 U3540 ( .A(n3551), .B(n3552), .ZN(n3435) );
  XNOR2_X1 U3541 ( .A(n3553), .B(n3554), .ZN(n3551) );
  XNOR2_X1 U3542 ( .A(n3555), .B(n3556), .ZN(n3439) );
  XNOR2_X1 U3543 ( .A(n3557), .B(n3558), .ZN(n3555) );
  XNOR2_X1 U3544 ( .A(n3559), .B(n3560), .ZN(n3324) );
  XNOR2_X1 U3545 ( .A(n3561), .B(n3562), .ZN(n3559) );
  NOR2_X1 U3546 ( .A1(n3563), .A2(n3328), .ZN(n3446) );
  XOR2_X1 U3547 ( .A(n3564), .B(n3565), .Z(n3328) );
  NAND2_X1 U3548 ( .A1(n3566), .A2(n3567), .ZN(n3564) );
  NOR2_X1 U3549 ( .A1(n3445), .A2(n3444), .ZN(n3563) );
  NAND2_X1 U3550 ( .A1(n3568), .A2(n3569), .ZN(n1914) );
  XOR2_X1 U3551 ( .A(n3570), .B(n3571), .Z(n3568) );
  NOR2_X1 U3552 ( .A1(n1913), .A2(n3572), .ZN(n1956) );
  AND2_X1 U3553 ( .A1(n3573), .A2(n3448), .ZN(n1913) );
  INV_X1 U3554 ( .A(n3569), .ZN(n3448) );
  NAND2_X1 U3555 ( .A1(n3445), .A2(n3444), .ZN(n3569) );
  NAND2_X1 U3556 ( .A1(n3566), .A2(n3574), .ZN(n3444) );
  NAND2_X1 U3557 ( .A1(n3565), .A2(n3567), .ZN(n3574) );
  NAND2_X1 U3558 ( .A1(n3575), .A2(n3576), .ZN(n3567) );
  NAND2_X1 U3559 ( .A1(a_0_), .A2(b_2_), .ZN(n3576) );
  INV_X1 U3560 ( .A(n3577), .ZN(n3575) );
  XOR2_X1 U3561 ( .A(n3578), .B(n3579), .Z(n3565) );
  NOR2_X1 U3562 ( .A1(n3580), .A2(n2000), .ZN(n3579) );
  XOR2_X1 U3563 ( .A(n3581), .B(n3582), .Z(n3578) );
  NAND2_X1 U3564 ( .A1(a_0_), .A2(n3577), .ZN(n3566) );
  NAND2_X1 U3565 ( .A1(n3583), .A2(n3584), .ZN(n3577) );
  NAND2_X1 U3566 ( .A1(n3562), .A2(n3585), .ZN(n3584) );
  NAND2_X1 U3567 ( .A1(n3561), .A2(n3560), .ZN(n3585) );
  NOR2_X1 U3568 ( .A1(n1995), .A2(n3396), .ZN(n3562) );
  OR2_X1 U3569 ( .A1(n3560), .A2(n3561), .ZN(n3583) );
  AND2_X1 U3570 ( .A1(n3586), .A2(n3587), .ZN(n3561) );
  NAND2_X1 U3571 ( .A1(n3558), .A2(n3588), .ZN(n3587) );
  NAND2_X1 U3572 ( .A1(n3557), .A2(n3556), .ZN(n3588) );
  OR2_X1 U3573 ( .A1(n3556), .A2(n3557), .ZN(n3586) );
  AND2_X1 U3574 ( .A1(n3589), .A2(n3590), .ZN(n3557) );
  NAND2_X1 U3575 ( .A1(n3554), .A2(n3591), .ZN(n3590) );
  NAND2_X1 U3576 ( .A1(n3553), .A2(n3552), .ZN(n3591) );
  NOR2_X1 U3577 ( .A1(n1919), .A2(n3396), .ZN(n3554) );
  OR2_X1 U3578 ( .A1(n3552), .A2(n3553), .ZN(n3589) );
  AND2_X1 U3579 ( .A1(n3466), .A2(n3592), .ZN(n3553) );
  NAND2_X1 U3580 ( .A1(n3465), .A2(n3467), .ZN(n3592) );
  NAND2_X1 U3581 ( .A1(n3593), .A2(n3594), .ZN(n3467) );
  NAND2_X1 U3582 ( .A1(b_2_), .A2(a_4_), .ZN(n3594) );
  INV_X1 U3583 ( .A(n3595), .ZN(n3593) );
  XOR2_X1 U3584 ( .A(n3596), .B(n3597), .Z(n3465) );
  NOR2_X1 U3585 ( .A1(n2014), .A2(n3529), .ZN(n3597) );
  XOR2_X1 U3586 ( .A(n3598), .B(n3599), .Z(n3596) );
  NAND2_X1 U3587 ( .A1(a_4_), .A2(n3595), .ZN(n3466) );
  NAND2_X1 U3588 ( .A1(n3600), .A2(n3601), .ZN(n3595) );
  NAND2_X1 U3589 ( .A1(n3550), .A2(n3602), .ZN(n3601) );
  NAND2_X1 U3590 ( .A1(n3549), .A2(n3548), .ZN(n3602) );
  NOR2_X1 U3591 ( .A1(n3396), .A2(n2014), .ZN(n3550) );
  OR2_X1 U3592 ( .A1(n3548), .A2(n3549), .ZN(n3600) );
  AND2_X1 U3593 ( .A1(n3545), .A2(n3603), .ZN(n3549) );
  NAND2_X1 U3594 ( .A1(n3544), .A2(n3546), .ZN(n3603) );
  NAND2_X1 U3595 ( .A1(n3604), .A2(n3605), .ZN(n3546) );
  NAND2_X1 U3596 ( .A1(a_6_), .A2(b_2_), .ZN(n3605) );
  INV_X1 U3597 ( .A(n3606), .ZN(n3604) );
  XOR2_X1 U3598 ( .A(n3607), .B(n3608), .Z(n3544) );
  NOR2_X1 U3599 ( .A1(n2170), .A2(n3529), .ZN(n3608) );
  XOR2_X1 U3600 ( .A(n3609), .B(n3610), .Z(n3607) );
  NAND2_X1 U3601 ( .A1(a_6_), .A2(n3606), .ZN(n3545) );
  NAND2_X1 U3602 ( .A1(n3611), .A2(n3612), .ZN(n3606) );
  NAND2_X1 U3603 ( .A1(n3542), .A2(n3613), .ZN(n3612) );
  NAND2_X1 U3604 ( .A1(n3541), .A2(n3540), .ZN(n3613) );
  NOR2_X1 U3605 ( .A1(n3396), .A2(n2170), .ZN(n3542) );
  OR2_X1 U3606 ( .A1(n3540), .A2(n3541), .ZN(n3611) );
  AND2_X1 U3607 ( .A1(n3486), .A2(n3614), .ZN(n3541) );
  NAND2_X1 U3608 ( .A1(n3485), .A2(n3487), .ZN(n3614) );
  NAND2_X1 U3609 ( .A1(n3615), .A2(n3616), .ZN(n3487) );
  NAND2_X1 U3610 ( .A1(b_2_), .A2(a_8_), .ZN(n3616) );
  INV_X1 U3611 ( .A(n3617), .ZN(n3615) );
  XOR2_X1 U3612 ( .A(n3618), .B(n3619), .Z(n3485) );
  XNOR2_X1 U3613 ( .A(n3620), .B(n3621), .ZN(n3619) );
  NAND2_X1 U3614 ( .A1(b_1_), .A2(a_9_), .ZN(n3618) );
  NAND2_X1 U3615 ( .A1(a_8_), .A2(n3617), .ZN(n3486) );
  NAND2_X1 U3616 ( .A1(n3622), .A2(n3623), .ZN(n3617) );
  NAND2_X1 U3617 ( .A1(n3538), .A2(n3624), .ZN(n3623) );
  NAND2_X1 U3618 ( .A1(n3537), .A2(n3536), .ZN(n3624) );
  NOR2_X1 U3619 ( .A1(n3396), .A2(n2178), .ZN(n3538) );
  OR2_X1 U3620 ( .A1(n3536), .A2(n3537), .ZN(n3622) );
  AND2_X1 U3621 ( .A1(n3498), .A2(n3625), .ZN(n3537) );
  NAND2_X1 U3622 ( .A1(n3497), .A2(n3499), .ZN(n3625) );
  NAND2_X1 U3623 ( .A1(n3626), .A2(n3627), .ZN(n3499) );
  NAND2_X1 U3624 ( .A1(b_2_), .A2(a_10_), .ZN(n3627) );
  INV_X1 U3625 ( .A(n3628), .ZN(n3626) );
  XOR2_X1 U3626 ( .A(n3629), .B(n3630), .Z(n3497) );
  NOR2_X1 U3627 ( .A1(n3260), .A2(n3529), .ZN(n3630) );
  XOR2_X1 U3628 ( .A(n3631), .B(n3632), .Z(n3629) );
  NAND2_X1 U3629 ( .A1(a_10_), .A2(n3628), .ZN(n3498) );
  NAND2_X1 U3630 ( .A1(n3633), .A2(n3634), .ZN(n3628) );
  NAND2_X1 U3631 ( .A1(n3507), .A2(n3635), .ZN(n3634) );
  OR2_X1 U3632 ( .A1(n3506), .A2(n3504), .ZN(n3635) );
  NOR2_X1 U3633 ( .A1(n3396), .A2(n3260), .ZN(n3507) );
  NAND2_X1 U3634 ( .A1(n3504), .A2(n3506), .ZN(n3633) );
  NAND2_X1 U3635 ( .A1(n3636), .A2(n3637), .ZN(n3506) );
  NAND2_X1 U3636 ( .A1(n3514), .A2(n3638), .ZN(n3637) );
  NAND2_X1 U3637 ( .A1(n3513), .A2(n3515), .ZN(n3638) );
  NOR2_X1 U3638 ( .A1(n3396), .A2(n2057), .ZN(n3514) );
  OR2_X1 U3639 ( .A1(n3513), .A2(n3515), .ZN(n3636) );
  AND2_X1 U3640 ( .A1(n3639), .A2(n3640), .ZN(n3515) );
  NAND2_X1 U3641 ( .A1(n3641), .A2(b_2_), .ZN(n3640) );
  NOR2_X1 U3642 ( .A1(n3642), .A2(n1870), .ZN(n3641) );
  NOR2_X1 U3643 ( .A1(n3533), .A2(n3534), .ZN(n3642) );
  NAND2_X1 U3644 ( .A1(n3533), .A2(n3534), .ZN(n3639) );
  NAND2_X1 U3645 ( .A1(n3643), .A2(n3644), .ZN(n3534) );
  NAND2_X1 U3646 ( .A1(n3645), .A2(b_0_), .ZN(n3644) );
  NOR2_X1 U3647 ( .A1(n3646), .A2(n2071), .ZN(n3645) );
  NOR2_X1 U3648 ( .A1(n2070), .A2(n3529), .ZN(n3646) );
  INV_X1 U3649 ( .A(n1857), .ZN(n2070) );
  NAND2_X1 U3650 ( .A1(a_15_), .A2(n2208), .ZN(n1857) );
  NAND2_X1 U3651 ( .A1(n3647), .A2(b_1_), .ZN(n3643) );
  NOR2_X1 U3652 ( .A1(n3648), .A2(n2208), .ZN(n3647) );
  NOR2_X1 U3653 ( .A1(n2064), .A2(n3580), .ZN(n3648) );
  INV_X1 U3654 ( .A(n1861), .ZN(n2064) );
  NAND2_X1 U3655 ( .A1(a_14_), .A2(n2071), .ZN(n1861) );
  INV_X1 U3656 ( .A(a_15_), .ZN(n2071) );
  AND2_X1 U3657 ( .A1(n3649), .A2(b_1_), .ZN(n3533) );
  NOR2_X1 U3658 ( .A1(n2210), .A2(n3396), .ZN(n3649) );
  XNOR2_X1 U3659 ( .A(n3650), .B(n3651), .ZN(n3513) );
  XNOR2_X1 U3660 ( .A(n3652), .B(n3653), .ZN(n3651) );
  XOR2_X1 U3661 ( .A(n3654), .B(n3655), .Z(n3504) );
  XOR2_X1 U3662 ( .A(n3656), .B(n3657), .Z(n3654) );
  XNOR2_X1 U3663 ( .A(n3658), .B(n3659), .ZN(n3536) );
  XOR2_X1 U3664 ( .A(n3660), .B(n3661), .Z(n3658) );
  XOR2_X1 U3665 ( .A(n3662), .B(n3663), .Z(n3540) );
  XNOR2_X1 U3666 ( .A(n3664), .B(n3665), .ZN(n3663) );
  XOR2_X1 U3667 ( .A(n3666), .B(n3667), .Z(n3548) );
  XOR2_X1 U3668 ( .A(n3668), .B(n3669), .Z(n3667) );
  XNOR2_X1 U3669 ( .A(n3670), .B(n3671), .ZN(n3552) );
  XOR2_X1 U3670 ( .A(n3672), .B(n3673), .Z(n3670) );
  XNOR2_X1 U3671 ( .A(n3674), .B(n3675), .ZN(n3556) );
  NOR2_X1 U3672 ( .A1(n3529), .A2(n1919), .ZN(n3675) );
  XOR2_X1 U3673 ( .A(n3676), .B(n3677), .Z(n3674) );
  XNOR2_X1 U3674 ( .A(n3678), .B(n3679), .ZN(n3560) );
  NOR2_X1 U3675 ( .A1(n3680), .A2(n3681), .ZN(n3679) );
  INV_X1 U3676 ( .A(n3682), .ZN(n3681) );
  NOR2_X1 U3677 ( .A1(n3683), .A2(n3684), .ZN(n3680) );
  XOR2_X1 U3678 ( .A(n3685), .B(n3686), .Z(n3445) );
  NOR2_X1 U3679 ( .A1(n3687), .A2(n3688), .ZN(n3686) );
  INV_X1 U3680 ( .A(n3689), .ZN(n3688) );
  NOR2_X1 U3681 ( .A1(n3690), .A2(n3691), .ZN(n3687) );
  NOR2_X1 U3682 ( .A1(n3572), .A2(n3570), .ZN(n3573) );
  AND2_X1 U3683 ( .A1(a_0_), .A2(n3571), .ZN(n3572) );
  NAND2_X1 U3684 ( .A1(n3689), .A2(n3692), .ZN(n3571) );
  NAND2_X1 U3685 ( .A1(n3693), .A2(n3685), .ZN(n3692) );
  NAND2_X1 U3686 ( .A1(n3694), .A2(n3695), .ZN(n3685) );
  NAND2_X1 U3687 ( .A1(n3696), .A2(a_2_), .ZN(n3695) );
  NOR2_X1 U3688 ( .A1(n3697), .A2(n3580), .ZN(n3696) );
  NOR2_X1 U3689 ( .A1(n3582), .A2(n3581), .ZN(n3697) );
  NAND2_X1 U3690 ( .A1(n3582), .A2(n3581), .ZN(n3694) );
  NAND2_X1 U3691 ( .A1(n3682), .A2(n3698), .ZN(n3581) );
  NAND2_X1 U3692 ( .A1(n3699), .A2(n3678), .ZN(n3698) );
  NAND2_X1 U3693 ( .A1(n3700), .A2(n3701), .ZN(n3678) );
  NAND2_X1 U3694 ( .A1(n3702), .A2(a_3_), .ZN(n3701) );
  NOR2_X1 U3695 ( .A1(n3703), .A2(n3529), .ZN(n3702) );
  NOR2_X1 U3696 ( .A1(n3676), .A2(n3677), .ZN(n3703) );
  NAND2_X1 U3697 ( .A1(n3676), .A2(n3677), .ZN(n3700) );
  NAND2_X1 U3698 ( .A1(n3704), .A2(n3705), .ZN(n3677) );
  NAND2_X1 U3699 ( .A1(n3671), .A2(n3706), .ZN(n3705) );
  OR2_X1 U3700 ( .A1(n3672), .A2(n3673), .ZN(n3706) );
  NOR2_X1 U3701 ( .A1(n3529), .A2(n2009), .ZN(n3671) );
  NAND2_X1 U3702 ( .A1(n3673), .A2(n3672), .ZN(n3704) );
  NAND2_X1 U3703 ( .A1(n3707), .A2(n3708), .ZN(n3672) );
  NAND2_X1 U3704 ( .A1(n3709), .A2(b_1_), .ZN(n3708) );
  NOR2_X1 U3705 ( .A1(n3710), .A2(n2014), .ZN(n3709) );
  NOR2_X1 U3706 ( .A1(n3599), .A2(n3598), .ZN(n3710) );
  NAND2_X1 U3707 ( .A1(n3599), .A2(n3598), .ZN(n3707) );
  NAND2_X1 U3708 ( .A1(n3711), .A2(n3712), .ZN(n3598) );
  NAND2_X1 U3709 ( .A1(n3666), .A2(n3713), .ZN(n3712) );
  NAND2_X1 U3710 ( .A1(n3669), .A2(n3714), .ZN(n3713) );
  INV_X1 U3711 ( .A(n3715), .ZN(n3669) );
  NOR2_X1 U3712 ( .A1(n3529), .A2(n2019), .ZN(n3666) );
  NAND2_X1 U3713 ( .A1(n3668), .A2(n3715), .ZN(n3711) );
  NAND2_X1 U3714 ( .A1(n3716), .A2(n3717), .ZN(n3715) );
  NAND2_X1 U3715 ( .A1(n3718), .A2(b_1_), .ZN(n3717) );
  NOR2_X1 U3716 ( .A1(n3719), .A2(n2170), .ZN(n3718) );
  NOR2_X1 U3717 ( .A1(n3609), .A2(n3610), .ZN(n3719) );
  NAND2_X1 U3718 ( .A1(n3609), .A2(n3610), .ZN(n3716) );
  NAND2_X1 U3719 ( .A1(n3720), .A2(n3721), .ZN(n3610) );
  NAND2_X1 U3720 ( .A1(n3662), .A2(n3722), .ZN(n3721) );
  OR2_X1 U3721 ( .A1(n3665), .A2(n3664), .ZN(n3722) );
  NOR2_X1 U3722 ( .A1(n3529), .A2(n2028), .ZN(n3662) );
  NAND2_X1 U3723 ( .A1(n3664), .A2(n3665), .ZN(n3720) );
  NAND2_X1 U3724 ( .A1(n3723), .A2(n3724), .ZN(n3665) );
  NAND2_X1 U3725 ( .A1(n3725), .A2(b_1_), .ZN(n3724) );
  NOR2_X1 U3726 ( .A1(n3726), .A2(n2178), .ZN(n3725) );
  NOR2_X1 U3727 ( .A1(n3621), .A2(n3620), .ZN(n3726) );
  NAND2_X1 U3728 ( .A1(n3621), .A2(n3620), .ZN(n3723) );
  NAND2_X1 U3729 ( .A1(n3727), .A2(n3728), .ZN(n3620) );
  NAND2_X1 U3730 ( .A1(n3659), .A2(n3729), .ZN(n3728) );
  OR2_X1 U3731 ( .A1(n3661), .A2(n3660), .ZN(n3729) );
  NOR2_X1 U3732 ( .A1(n3529), .A2(n1885), .ZN(n3659) );
  NAND2_X1 U3733 ( .A1(n3660), .A2(n3661), .ZN(n3727) );
  NAND2_X1 U3734 ( .A1(n3730), .A2(n3731), .ZN(n3661) );
  NAND2_X1 U3735 ( .A1(n3732), .A2(b_1_), .ZN(n3731) );
  NOR2_X1 U3736 ( .A1(n3733), .A2(n3260), .ZN(n3732) );
  NOR2_X1 U3737 ( .A1(n3631), .A2(n3632), .ZN(n3733) );
  NAND2_X1 U3738 ( .A1(n3631), .A2(n3632), .ZN(n3730) );
  NAND2_X1 U3739 ( .A1(n3734), .A2(n3735), .ZN(n3632) );
  NAND2_X1 U3740 ( .A1(n3655), .A2(n3736), .ZN(n3735) );
  OR2_X1 U3741 ( .A1(n3656), .A2(n3657), .ZN(n3736) );
  NOR2_X1 U3742 ( .A1(n3529), .A2(n2057), .ZN(n3655) );
  NAND2_X1 U3743 ( .A1(n3657), .A2(n3656), .ZN(n3734) );
  NAND2_X1 U3744 ( .A1(n3737), .A2(n3653), .ZN(n3656) );
  NAND2_X1 U3745 ( .A1(n3738), .A2(b_0_), .ZN(n3653) );
  NOR2_X1 U3746 ( .A1(n2210), .A2(n3529), .ZN(n3738) );
  NAND2_X1 U3747 ( .A1(a_15_), .A2(a_14_), .ZN(n2210) );
  NAND2_X1 U3748 ( .A1(n3650), .A2(n3652), .ZN(n3737) );
  NOR2_X1 U3749 ( .A1(n3529), .A2(n1870), .ZN(n3652) );
  NOR2_X1 U3750 ( .A1(n3580), .A2(n2208), .ZN(n3650) );
  NOR2_X1 U3751 ( .A1(n3580), .A2(n1870), .ZN(n3657) );
  NOR2_X1 U3752 ( .A1(n3580), .A2(n2057), .ZN(n3631) );
  NOR2_X1 U3753 ( .A1(n3580), .A2(n3260), .ZN(n3660) );
  NOR2_X1 U3754 ( .A1(n3580), .A2(n1885), .ZN(n3621) );
  NOR2_X1 U3755 ( .A1(n3580), .A2(n2178), .ZN(n3664) );
  NOR2_X1 U3756 ( .A1(n3580), .A2(n2028), .ZN(n3609) );
  INV_X1 U3757 ( .A(n3714), .ZN(n3668) );
  NAND2_X1 U3758 ( .A1(b_0_), .A2(a_7_), .ZN(n3714) );
  NOR2_X1 U3759 ( .A1(n3580), .A2(n2019), .ZN(n3599) );
  NOR2_X1 U3760 ( .A1(n3580), .A2(n2014), .ZN(n3673) );
  NOR2_X1 U3761 ( .A1(n3580), .A2(n2009), .ZN(n3676) );
  OR2_X1 U3762 ( .A1(n3683), .A2(a_2_), .ZN(n3699) );
  NAND2_X1 U3763 ( .A1(n3684), .A2(n3683), .ZN(n3682) );
  NOR2_X1 U3764 ( .A1(n1919), .A2(n3580), .ZN(n3683) );
  NOR2_X1 U3765 ( .A1(n3529), .A2(n2000), .ZN(n3684) );
  OR2_X1 U3766 ( .A1(n3690), .A2(a_0_), .ZN(n3693) );
  NAND2_X1 U3767 ( .A1(n3691), .A2(n3690), .ZN(n3689) );
  NOR2_X1 U3768 ( .A1(n1995), .A2(n3580), .ZN(n3690) );
  INV_X1 U3769 ( .A(b_0_), .ZN(n3580) );
  NOR2_X1 U3770 ( .A1(n3529), .A2(n1986), .ZN(n3691) );
  INV_X1 U3771 ( .A(a_0_), .ZN(n1986) );
  NAND2_X1 U3772 ( .A1(n3739), .A2(n3740), .ZN(Result_add_9_) );
  NAND2_X1 U3773 ( .A1(n2758), .A2(n3741), .ZN(n3740) );
  INV_X1 U3774 ( .A(n2679), .ZN(n2758) );
  NOR2_X1 U3775 ( .A1(n3742), .A2(n3743), .ZN(n3739) );
  NOR2_X1 U3776 ( .A1(b_9_), .A2(n3744), .ZN(n3743) );
  XOR2_X1 U3777 ( .A(n2178), .B(n3741), .Z(n3744) );
  NOR2_X1 U3778 ( .A1(n2542), .A2(n3745), .ZN(n3742) );
  OR2_X1 U3779 ( .A1(n3741), .A2(a_9_), .ZN(n3745) );
  XOR2_X1 U3780 ( .A(n3746), .B(n3747), .Z(Result_add_8_) );
  AND2_X1 U3781 ( .A1(n3748), .A2(n2873), .ZN(n3747) );
  NAND2_X1 U3782 ( .A1(n3749), .A2(n3750), .ZN(Result_add_7_) );
  NAND2_X1 U3783 ( .A1(n2927), .A2(n3751), .ZN(n3750) );
  INV_X1 U3784 ( .A(n3752), .ZN(n2927) );
  NOR2_X1 U3785 ( .A1(n3753), .A2(n3754), .ZN(n3749) );
  NOR2_X1 U3786 ( .A1(b_7_), .A2(n3755), .ZN(n3754) );
  XOR2_X1 U3787 ( .A(n2170), .B(n3751), .Z(n3755) );
  NOR2_X1 U3788 ( .A1(n2789), .A2(n3756), .ZN(n3753) );
  OR2_X1 U3789 ( .A1(n3751), .A2(a_7_), .ZN(n3756) );
  XOR2_X1 U3790 ( .A(n3757), .B(n3758), .Z(Result_add_6_) );
  AND2_X1 U3791 ( .A1(n3759), .A2(n3054), .ZN(n3758) );
  NAND2_X1 U3792 ( .A1(n3760), .A2(n3761), .ZN(Result_add_5_) );
  NAND2_X1 U3793 ( .A1(n3182), .A2(n3762), .ZN(n3761) );
  NOR2_X1 U3794 ( .A1(n3763), .A2(n3764), .ZN(n3760) );
  NOR2_X1 U3795 ( .A1(b_5_), .A2(n3765), .ZN(n3764) );
  XOR2_X1 U3796 ( .A(n2014), .B(n3762), .Z(n3765) );
  NOR2_X1 U3797 ( .A1(n3033), .A2(n3766), .ZN(n3763) );
  OR2_X1 U3798 ( .A1(n3762), .A2(a_5_), .ZN(n3766) );
  XNOR2_X1 U3799 ( .A(n3767), .B(n3768), .ZN(Result_add_4_) );
  NOR2_X1 U3800 ( .A1(n3769), .A2(n3306), .ZN(n3768) );
  NAND2_X1 U3801 ( .A1(n3770), .A2(n3771), .ZN(Result_add_3_) );
  NAND2_X1 U3802 ( .A1(n3433), .A2(n3772), .ZN(n3771) );
  INV_X1 U3803 ( .A(n3773), .ZN(n3433) );
  NOR2_X1 U3804 ( .A1(n3774), .A2(n3775), .ZN(n3770) );
  NOR2_X1 U3805 ( .A1(b_3_), .A2(n3776), .ZN(n3775) );
  XOR2_X1 U3806 ( .A(n1919), .B(n3772), .Z(n3776) );
  NOR2_X1 U3807 ( .A1(n3274), .A2(n3777), .ZN(n3774) );
  NAND2_X1 U3808 ( .A1(n3778), .A2(n1919), .ZN(n3777) );
  XNOR2_X1 U3809 ( .A(n3779), .B(n3780), .ZN(Result_add_2_) );
  NOR2_X1 U3810 ( .A1(n3781), .A2(n3558), .ZN(n3780) );
  NAND2_X1 U3811 ( .A1(n3782), .A2(n3783), .ZN(Result_add_1_) );
  NAND2_X1 U3812 ( .A1(n3784), .A2(n3785), .ZN(n3783) );
  OR2_X1 U3813 ( .A1(n3582), .A2(n3786), .ZN(n3784) );
  NAND2_X1 U3814 ( .A1(n3787), .A2(n3788), .ZN(n3782) );
  XOR2_X1 U3815 ( .A(b_1_), .B(a_1_), .Z(n3787) );
  XOR2_X1 U3816 ( .A(b_15_), .B(a_15_), .Z(Result_add_15_) );
  NAND2_X1 U3817 ( .A1(n3789), .A2(n3790), .ZN(Result_add_14_) );
  INV_X1 U3818 ( .A(n1871), .ZN(n3790) );
  NOR2_X1 U3819 ( .A1(n2072), .A2(n3791), .ZN(n1871) );
  NOR2_X1 U3820 ( .A1(n3792), .A2(n3793), .ZN(n3789) );
  NOR2_X1 U3821 ( .A1(n1863), .A2(n3794), .ZN(n3793) );
  NAND2_X1 U3822 ( .A1(n3791), .A2(n2208), .ZN(n3794) );
  NOR2_X1 U3823 ( .A1(b_14_), .A2(n3795), .ZN(n3792) );
  XOR2_X1 U3824 ( .A(n3791), .B(a_14_), .Z(n3795) );
  NAND2_X1 U3825 ( .A1(n3796), .A2(n3797), .ZN(Result_add_13_) );
  NAND2_X1 U3826 ( .A1(n2212), .A2(n3798), .ZN(n3797) );
  INV_X1 U3827 ( .A(n3799), .ZN(n2212) );
  NOR2_X1 U3828 ( .A1(n3800), .A2(n3801), .ZN(n3796) );
  NOR2_X1 U3829 ( .A1(b_13_), .A2(n3802), .ZN(n3801) );
  XOR2_X1 U3830 ( .A(a_13_), .B(n3803), .Z(n3802) );
  NOR2_X1 U3831 ( .A1(n2068), .A2(n3804), .ZN(n3800) );
  NAND2_X1 U3832 ( .A1(n3803), .A2(n1870), .ZN(n3804) );
  INV_X1 U3833 ( .A(n3798), .ZN(n3803) );
  XNOR2_X1 U3834 ( .A(n3805), .B(n3806), .ZN(Result_add_12_) );
  NOR2_X1 U3835 ( .A1(n3807), .A2(n2296), .ZN(n3806) );
  NAND2_X1 U3836 ( .A1(n3808), .A2(n3809), .ZN(Result_add_11_) );
  NAND2_X1 U3837 ( .A1(n2399), .A2(n3810), .ZN(n3809) );
  INV_X1 U3838 ( .A(n3811), .ZN(n2399) );
  NOR2_X1 U3839 ( .A1(n3812), .A2(n3813), .ZN(n3808) );
  NOR2_X1 U3840 ( .A1(b_11_), .A2(n3814), .ZN(n3813) );
  XOR2_X1 U3841 ( .A(n3260), .B(n3810), .Z(n3814) );
  NOR2_X1 U3842 ( .A1(n2308), .A2(n3815), .ZN(n3812) );
  NAND2_X1 U3843 ( .A1(n3816), .A2(n3260), .ZN(n3815) );
  XOR2_X1 U3844 ( .A(n3817), .B(n3818), .Z(Result_add_10_) );
  AND2_X1 U3845 ( .A1(n3819), .A2(n2640), .ZN(n3818) );
  XOR2_X1 U3846 ( .A(n3820), .B(n3821), .Z(Result_add_0_) );
  NOR2_X1 U3847 ( .A1(n3822), .A2(n3823), .ZN(n3821) );
  INV_X1 U3848 ( .A(n3570), .ZN(n3823) );
  NAND2_X1 U3849 ( .A1(a_0_), .A2(b_0_), .ZN(n3570) );
  NOR2_X1 U3850 ( .A1(b_0_), .A2(a_0_), .ZN(n3822) );
  NOR2_X1 U3851 ( .A1(n3786), .A2(n3824), .ZN(n3820) );
  NOR2_X1 U3852 ( .A1(n3582), .A2(n3785), .ZN(n3824) );
  INV_X1 U3853 ( .A(n3788), .ZN(n3785) );
  NOR2_X1 U3854 ( .A1(n3558), .A2(n3825), .ZN(n3788) );
  NOR2_X1 U3855 ( .A1(n3781), .A2(n3779), .ZN(n3825) );
  AND2_X1 U3856 ( .A1(n3773), .A2(n3826), .ZN(n3779) );
  NAND2_X1 U3857 ( .A1(n3827), .A2(n3772), .ZN(n3826) );
  INV_X1 U3858 ( .A(n3778), .ZN(n3772) );
  NOR2_X1 U3859 ( .A1(n3306), .A2(n3828), .ZN(n3778) );
  NOR2_X1 U3860 ( .A1(n3769), .A2(n3767), .ZN(n3828) );
  NOR2_X1 U3861 ( .A1(n3182), .A2(n3829), .ZN(n3767) );
  AND2_X1 U3862 ( .A1(n3830), .A2(n3762), .ZN(n3829) );
  NAND2_X1 U3863 ( .A1(n3054), .A2(n3831), .ZN(n3762) );
  NAND2_X1 U3864 ( .A1(n3759), .A2(n3757), .ZN(n3831) );
  NAND2_X1 U3865 ( .A1(n3752), .A2(n3832), .ZN(n3757) );
  NAND2_X1 U3866 ( .A1(n3833), .A2(n3751), .ZN(n3832) );
  NAND2_X1 U3867 ( .A1(n2873), .A2(n3834), .ZN(n3751) );
  NAND2_X1 U3868 ( .A1(n3748), .A2(n3746), .ZN(n3834) );
  NAND2_X1 U3869 ( .A1(n2679), .A2(n3835), .ZN(n3746) );
  NAND2_X1 U3870 ( .A1(n3836), .A2(n3741), .ZN(n3835) );
  NAND2_X1 U3871 ( .A1(n2640), .A2(n3837), .ZN(n3741) );
  NAND2_X1 U3872 ( .A1(n3819), .A2(n3817), .ZN(n3837) );
  NAND2_X1 U3873 ( .A1(n3811), .A2(n3838), .ZN(n3817) );
  NAND2_X1 U3874 ( .A1(n3839), .A2(n3810), .ZN(n3838) );
  INV_X1 U3875 ( .A(n3816), .ZN(n3810) );
  NOR2_X1 U3876 ( .A1(n2296), .A2(n3840), .ZN(n3816) );
  NOR2_X1 U3877 ( .A1(n3807), .A2(n3805), .ZN(n3840) );
  AND2_X1 U3878 ( .A1(n3799), .A2(n3841), .ZN(n3805) );
  NAND2_X1 U3879 ( .A1(n3842), .A2(n3798), .ZN(n3841) );
  NAND2_X1 U3880 ( .A1(n2072), .A2(n3843), .ZN(n3798) );
  NAND2_X1 U3881 ( .A1(Result_mul_31_), .A2(n3844), .ZN(n3843) );
  NAND2_X1 U3882 ( .A1(n1863), .A2(n2208), .ZN(n3844) );
  INV_X1 U3883 ( .A(a_14_), .ZN(n2208) );
  INV_X1 U3884 ( .A(b_14_), .ZN(n1863) );
  INV_X1 U3885 ( .A(n3791), .ZN(Result_mul_31_) );
  NAND2_X1 U3886 ( .A1(b_15_), .A2(a_15_), .ZN(n3791) );
  NAND2_X1 U3887 ( .A1(b_14_), .A2(a_14_), .ZN(n2072) );
  NAND2_X1 U3888 ( .A1(n2068), .A2(n1870), .ZN(n3842) );
  INV_X1 U3889 ( .A(a_13_), .ZN(n1870) );
  INV_X1 U3890 ( .A(b_13_), .ZN(n2068) );
  NAND2_X1 U3891 ( .A1(b_13_), .A2(a_13_), .ZN(n3799) );
  NOR2_X1 U3892 ( .A1(b_12_), .A2(a_12_), .ZN(n3807) );
  NOR2_X1 U3893 ( .A1(n2123), .A2(n2057), .ZN(n2296) );
  INV_X1 U3894 ( .A(a_12_), .ZN(n2057) );
  INV_X1 U3895 ( .A(b_12_), .ZN(n2123) );
  NAND2_X1 U3896 ( .A1(n2308), .A2(n3260), .ZN(n3839) );
  INV_X1 U3897 ( .A(a_11_), .ZN(n3260) );
  INV_X1 U3898 ( .A(b_11_), .ZN(n2308) );
  NAND2_X1 U3899 ( .A1(a_11_), .A2(b_11_), .ZN(n3811) );
  NAND2_X1 U3900 ( .A1(n2418), .A2(n1885), .ZN(n3819) );
  INV_X1 U3901 ( .A(a_10_), .ZN(n1885) );
  INV_X1 U3902 ( .A(b_10_), .ZN(n2418) );
  NAND2_X1 U3903 ( .A1(a_10_), .A2(b_10_), .ZN(n2640) );
  NAND2_X1 U3904 ( .A1(n2542), .A2(n2178), .ZN(n3836) );
  INV_X1 U3905 ( .A(a_9_), .ZN(n2178) );
  INV_X1 U3906 ( .A(b_9_), .ZN(n2542) );
  NAND2_X1 U3907 ( .A1(b_9_), .A2(a_9_), .ZN(n2679) );
  NAND2_X1 U3908 ( .A1(n2662), .A2(n2028), .ZN(n3748) );
  INV_X1 U3909 ( .A(a_8_), .ZN(n2028) );
  INV_X1 U3910 ( .A(b_8_), .ZN(n2662) );
  NAND2_X1 U3911 ( .A1(a_8_), .A2(b_8_), .ZN(n2873) );
  NAND2_X1 U3912 ( .A1(n2789), .A2(n2170), .ZN(n3833) );
  INV_X1 U3913 ( .A(a_7_), .ZN(n2170) );
  INV_X1 U3914 ( .A(b_7_), .ZN(n2789) );
  NAND2_X1 U3915 ( .A1(b_7_), .A2(a_7_), .ZN(n3752) );
  NAND2_X1 U3916 ( .A1(n2906), .A2(n2019), .ZN(n3759) );
  INV_X1 U3917 ( .A(a_6_), .ZN(n2019) );
  INV_X1 U3918 ( .A(b_6_), .ZN(n2906) );
  NAND2_X1 U3919 ( .A1(a_6_), .A2(b_6_), .ZN(n3054) );
  NAND2_X1 U3920 ( .A1(n3033), .A2(n2014), .ZN(n3830) );
  NOR2_X1 U3921 ( .A1(n3033), .A2(n2014), .ZN(n3182) );
  INV_X1 U3922 ( .A(a_5_), .ZN(n2014) );
  INV_X1 U3923 ( .A(b_5_), .ZN(n3033) );
  NOR2_X1 U3924 ( .A1(b_4_), .A2(a_4_), .ZN(n3769) );
  NOR2_X1 U3925 ( .A1(n3170), .A2(n2009), .ZN(n3306) );
  INV_X1 U3926 ( .A(a_4_), .ZN(n2009) );
  INV_X1 U3927 ( .A(b_4_), .ZN(n3170) );
  NAND2_X1 U3928 ( .A1(n3274), .A2(n1919), .ZN(n3827) );
  INV_X1 U3929 ( .A(a_3_), .ZN(n1919) );
  INV_X1 U3930 ( .A(b_3_), .ZN(n3274) );
  NAND2_X1 U3931 ( .A1(a_3_), .A2(b_3_), .ZN(n3773) );
  NOR2_X1 U3932 ( .A1(b_2_), .A2(a_2_), .ZN(n3781) );
  NOR2_X1 U3933 ( .A1(n2000), .A2(n3396), .ZN(n3558) );
  INV_X1 U3934 ( .A(b_2_), .ZN(n3396) );
  INV_X1 U3935 ( .A(a_2_), .ZN(n2000) );
  NOR2_X1 U3936 ( .A1(n1995), .A2(n3529), .ZN(n3582) );
  INV_X1 U3937 ( .A(b_1_), .ZN(n3529) );
  INV_X1 U3938 ( .A(a_1_), .ZN(n1995) );
  NOR2_X1 U3939 ( .A1(b_1_), .A2(a_1_), .ZN(n3786) );
endmodule

