module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n614_, new_n445_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n421_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n456_, new_n246_, new_n170_, new_n266_, new_n367_, new_n542_, new_n548_, new_n173_, new_n220_, new_n419_, new_n534_, new_n214_, new_n451_, new_n489_, new_n602_, new_n188_, new_n240_, new_n413_, new_n442_, new_n211_, new_n552_, new_n342_, new_n462_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n234_, new_n532_, new_n393_, new_n292_, new_n215_, new_n152_, new_n157_, new_n153_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n484_, new_n272_, new_n282_, new_n201_, new_n192_, new_n315_, new_n326_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n167_, new_n385_, new_n478_, new_n297_, new_n361_, new_n565_, new_n150_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n321_, new_n324_, new_n158_, new_n486_, new_n491_, new_n549_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n506_, new_n256_, new_n452_, new_n381_, new_n388_, new_n508_, new_n194_, new_n483_, new_n394_, new_n299_, new_n142_, new_n139_, new_n314_, new_n363_, new_n165_, new_n441_, new_n477_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n187_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n579_, new_n286_, new_n335_, new_n347_, new_n346_, new_n396_, new_n198_, new_n438_, new_n208_, new_n179_, new_n572_, new_n436_, new_n397_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n166_, new_n162_, new_n457_, new_n161_, new_n553_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n155_, new_n384_, new_n410_, new_n543_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n308_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n309_, new_n529_, new_n323_, new_n259_, new_n362_, new_n604_, new_n227_, new_n416_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n505_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n138_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n177_, new_n493_, new_n547_, new_n264_, new_n379_, new_n273_, new_n224_, new_n270_, new_n598_, new_n143_, new_n520_, new_n145_, new_n253_, new_n403_, new_n475_, new_n237_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n605_, new_n182_, new_n407_, new_n480_, new_n151_, new_n513_, new_n592_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n522_, new_n588_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n612_, new_n302_, new_n191_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n415_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n340_, new_n147_, new_n285_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n203_, new_n316_, new_n417_, new_n591_, new_n515_, new_n332_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n440_, new_n531_, new_n593_, new_n252_, new_n585_, new_n160_, new_n312_, new_n535_, new_n372_, new_n242_, new_n503_, new_n527_, new_n307_, new_n190_, new_n597_, new_n408_, new_n213_, new_n433_, new_n435_, new_n265_, new_n370_, new_n584_, new_n278_, new_n304_, new_n523_, new_n550_, new_n217_, new_n269_, new_n512_, new_n599_, new_n607_, new_n327_, new_n594_, new_n561_, new_n495_, new_n196_, new_n574_, new_n319_, new_n338_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n195_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n358_, new_n348_, new_n610_, new_n159_, new_n322_, new_n228_, new_n545_, new_n611_, new_n289_, new_n425_, new_n175_, new_n226_, new_n185_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n551_, new_n168_, new_n279_, new_n455_, new_n521_, new_n406_, new_n356_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n573_;

not g000 ( new_n138_, keyIn_0_41 );
not g001 ( new_n139_, keyIn_0_21 );
not g002 ( new_n140_, N37 );
xnor g003 ( new_n141_, keyIn_0_2, N33 );
xnor g004 ( new_n142_, new_n141_, new_n140_ );
xnor g005 ( new_n143_, N41, N45 );
xnor g006 ( new_n144_, new_n143_, keyIn_0_3 );
nand g007 ( new_n145_, new_n142_, new_n144_ );
xnor g008 ( new_n146_, new_n141_, N37 );
not g009 ( new_n147_, keyIn_0_3 );
xnor g010 ( new_n148_, new_n143_, new_n147_ );
nand g011 ( new_n149_, new_n146_, new_n148_ );
nand g012 ( new_n150_, new_n145_, new_n149_ );
nand g013 ( new_n151_, new_n150_, keyIn_0_17 );
not g014 ( new_n152_, keyIn_0_17 );
nand g015 ( new_n153_, new_n145_, new_n149_, new_n152_ );
nand g016 ( new_n154_, new_n151_, new_n153_ );
xnor g017 ( new_n155_, N1, N5 );
xnor g018 ( new_n156_, N9, N13 );
xnor g019 ( new_n157_, new_n155_, new_n156_ );
xnor g020 ( new_n158_, new_n157_, keyIn_0_16 );
nand g021 ( new_n159_, new_n154_, new_n158_ );
not g022 ( new_n160_, keyIn_0_16 );
xnor g023 ( new_n161_, new_n157_, new_n160_ );
nand g024 ( new_n162_, new_n151_, new_n153_, new_n161_ );
nand g025 ( new_n163_, new_n159_, new_n162_ );
nand g026 ( new_n164_, new_n163_, new_n139_ );
nand g027 ( new_n165_, new_n159_, keyIn_0_21, new_n162_ );
nand g028 ( new_n166_, new_n164_, new_n165_ );
nand g029 ( new_n167_, N135, N137 );
xnor g030 ( new_n168_, new_n167_, keyIn_0_10 );
nand g031 ( new_n169_, new_n166_, new_n168_ );
not g032 ( new_n170_, new_n168_ );
nand g033 ( new_n171_, new_n164_, new_n165_, new_n170_ );
nand g034 ( new_n172_, new_n169_, new_n171_ );
xor g035 ( new_n173_, N73, N89 );
xnor g036 ( new_n174_, N105, N121 );
xnor g037 ( new_n175_, new_n173_, new_n174_ );
xor g038 ( new_n176_, new_n175_, keyIn_0_20 );
nand g039 ( new_n177_, new_n172_, new_n176_ );
not g040 ( new_n178_, new_n176_ );
nand g041 ( new_n179_, new_n169_, new_n171_, new_n178_ );
nand g042 ( new_n180_, new_n177_, new_n179_ );
not g043 ( new_n181_, new_n180_ );
not g044 ( new_n182_, keyIn_0_4 );
xnor g045 ( new_n183_, N57, N61 );
xnor g046 ( new_n184_, new_n183_, new_n182_ );
xor g047 ( new_n185_, N49, N53 );
not g048 ( new_n186_, new_n185_ );
xnor g049 ( new_n187_, new_n184_, new_n186_ );
nand g050 ( new_n188_, new_n154_, new_n187_ );
xnor g051 ( new_n189_, new_n184_, new_n185_ );
nand g052 ( new_n190_, new_n151_, new_n153_, new_n189_ );
nand g053 ( new_n191_, N134, N137 );
nand g054 ( new_n192_, new_n188_, new_n190_, new_n191_ );
nand g055 ( new_n193_, new_n188_, new_n190_ );
not g056 ( new_n194_, new_n191_ );
nand g057 ( new_n195_, new_n193_, new_n194_ );
nand g058 ( new_n196_, new_n195_, new_n192_ );
xor g059 ( new_n197_, N69, N85 );
xnor g060 ( new_n198_, N101, N117 );
xor g061 ( new_n199_, new_n197_, new_n198_ );
nand g062 ( new_n200_, new_n196_, new_n199_ );
not g063 ( new_n201_, new_n199_ );
nand g064 ( new_n202_, new_n195_, new_n192_, new_n201_ );
nand g065 ( new_n203_, new_n200_, new_n202_ );
xnor g066 ( new_n204_, N25, N29 );
xnor g067 ( new_n205_, new_n204_, keyIn_0_1 );
xnor g068 ( new_n206_, N17, N21 );
xnor g069 ( new_n207_, new_n206_, keyIn_0_0 );
or g070 ( new_n208_, new_n205_, new_n207_ );
nand g071 ( new_n209_, new_n205_, new_n207_ );
nand g072 ( new_n210_, new_n208_, new_n209_ );
nand g073 ( new_n211_, new_n210_, new_n158_ );
nand g074 ( new_n212_, new_n161_, new_n208_, new_n209_ );
nand g075 ( new_n213_, N133, N137 );
nand g076 ( new_n214_, new_n212_, new_n211_, new_n213_ );
nand g077 ( new_n215_, new_n212_, new_n211_ );
nand g078 ( new_n216_, new_n215_, N133, N137 );
nand g079 ( new_n217_, new_n216_, new_n214_ );
xnor g080 ( new_n218_, N97, N113 );
xnor g081 ( new_n219_, new_n218_, keyIn_0_15 );
xnor g082 ( new_n220_, N65, N81 );
xnor g083 ( new_n221_, new_n219_, new_n220_ );
not g084 ( new_n222_, new_n221_ );
nand g085 ( new_n223_, new_n217_, new_n222_ );
nand g086 ( new_n224_, new_n216_, new_n214_, new_n221_ );
nand g087 ( new_n225_, new_n223_, new_n224_ );
not g088 ( new_n226_, new_n225_ );
nor g089 ( new_n227_, new_n203_, new_n226_ );
not g090 ( new_n228_, new_n227_ );
nand g091 ( new_n229_, new_n210_, new_n187_ );
nand g092 ( new_n230_, new_n189_, new_n208_, new_n209_ );
nand g093 ( new_n231_, new_n229_, new_n230_ );
nand g094 ( new_n232_, N136, N137 );
xnor g095 ( new_n233_, new_n232_, keyIn_0_11 );
not g096 ( new_n234_, new_n233_ );
nand g097 ( new_n235_, new_n231_, new_n234_ );
nand g098 ( new_n236_, new_n229_, new_n230_, new_n233_ );
xor g099 ( new_n237_, N77, N93 );
xnor g100 ( new_n238_, N109, N125 );
xor g101 ( new_n239_, new_n237_, new_n238_ );
nand g102 ( new_n240_, new_n235_, new_n236_, new_n239_ );
nand g103 ( new_n241_, new_n235_, new_n236_ );
not g104 ( new_n242_, new_n239_ );
nand g105 ( new_n243_, new_n241_, new_n242_ );
and g106 ( new_n244_, new_n243_, new_n240_ );
not g107 ( new_n245_, new_n244_ );
nor g108 ( new_n246_, new_n181_, new_n228_, new_n245_ );
nand g109 ( new_n247_, N65, N69 );
not g110 ( new_n248_, N65 );
not g111 ( new_n249_, N69 );
nand g112 ( new_n250_, new_n248_, new_n249_ );
nand g113 ( new_n251_, new_n250_, new_n247_ );
nand g114 ( new_n252_, new_n251_, keyIn_0_5 );
not g115 ( new_n253_, keyIn_0_5 );
nand g116 ( new_n254_, new_n250_, new_n253_, new_n247_ );
nand g117 ( new_n255_, new_n252_, new_n254_ );
nand g118 ( new_n256_, new_n255_, keyIn_0_6 );
not g119 ( new_n257_, keyIn_0_6 );
nand g120 ( new_n258_, new_n252_, new_n257_, new_n254_ );
nand g121 ( new_n259_, new_n256_, new_n258_ );
xnor g122 ( new_n260_, N73, N77 );
nand g123 ( new_n261_, new_n259_, new_n260_ );
not g124 ( new_n262_, new_n260_ );
nand g125 ( new_n263_, new_n256_, new_n258_, new_n262_ );
nand g126 ( new_n264_, new_n261_, new_n263_ );
xor g127 ( new_n265_, N81, N85 );
xnor g128 ( new_n266_, N89, N93 );
xnor g129 ( new_n267_, new_n265_, new_n266_ );
xnor g130 ( new_n268_, new_n264_, new_n267_ );
nand g131 ( new_n269_, N129, N137 );
or g132 ( new_n270_, new_n268_, new_n269_ );
nand g133 ( new_n271_, new_n268_, new_n269_ );
nand g134 ( new_n272_, new_n270_, new_n271_ );
xnor g135 ( new_n273_, N1, N17 );
xnor g136 ( new_n274_, N33, N49 );
xor g137 ( new_n275_, new_n273_, new_n274_ );
not g138 ( new_n276_, new_n275_ );
nand g139 ( new_n277_, new_n272_, new_n276_ );
nand g140 ( new_n278_, new_n270_, new_n271_, new_n275_ );
nand g141 ( new_n279_, new_n277_, new_n278_ );
not g142 ( new_n280_, keyIn_0_36 );
xnor g143 ( new_n281_, N121, N125 );
nand g144 ( new_n282_, new_n281_, keyIn_0_7 );
not g145 ( new_n283_, keyIn_0_7 );
nand g146 ( new_n284_, N121, N125 );
not g147 ( new_n285_, N121 );
not g148 ( new_n286_, N125 );
nand g149 ( new_n287_, new_n285_, new_n286_ );
nand g150 ( new_n288_, new_n287_, new_n283_, new_n284_ );
nand g151 ( new_n289_, new_n282_, new_n288_ );
xor g152 ( new_n290_, N113, N117 );
nand g153 ( new_n291_, new_n289_, new_n290_ );
not g154 ( new_n292_, new_n290_ );
nand g155 ( new_n293_, new_n292_, new_n282_, new_n288_ );
nand g156 ( new_n294_, new_n291_, new_n293_ );
nand g157 ( new_n295_, new_n294_, keyIn_0_19 );
not g158 ( new_n296_, keyIn_0_19 );
nand g159 ( new_n297_, new_n291_, new_n296_, new_n293_ );
nand g160 ( new_n298_, new_n295_, new_n297_ );
not g161 ( new_n299_, keyIn_0_18 );
xnor g162 ( new_n300_, N97, N101 );
xnor g163 ( new_n301_, N105, N109 );
xnor g164 ( new_n302_, new_n300_, new_n301_ );
xnor g165 ( new_n303_, new_n302_, new_n299_ );
nand g166 ( new_n304_, new_n298_, new_n303_ );
xnor g167 ( new_n305_, new_n302_, keyIn_0_18 );
nand g168 ( new_n306_, new_n305_, new_n295_, new_n297_ );
nand g169 ( new_n307_, new_n304_, new_n306_ );
nand g170 ( new_n308_, new_n307_, keyIn_0_22 );
not g171 ( new_n309_, keyIn_0_22 );
nand g172 ( new_n310_, new_n304_, new_n309_, new_n306_ );
nand g173 ( new_n311_, new_n308_, new_n310_ );
nand g174 ( new_n312_, new_n311_, keyIn_0_8 );
not g175 ( new_n313_, keyIn_0_8 );
nand g176 ( new_n314_, new_n308_, new_n313_, new_n310_ );
nand g177 ( new_n315_, new_n312_, new_n314_ );
nand g178 ( new_n316_, N130, N137 );
nand g179 ( new_n317_, new_n315_, new_n316_ );
nand g180 ( new_n318_, new_n312_, N130, N137, new_n314_ );
nand g181 ( new_n319_, new_n317_, new_n318_ );
xor g182 ( new_n320_, N37, N53 );
xnor g183 ( new_n321_, new_n320_, keyIn_0_13 );
xor g184 ( new_n322_, N5, N21 );
xnor g185 ( new_n323_, new_n322_, keyIn_0_12 );
xnor g186 ( new_n324_, new_n321_, new_n323_ );
nand g187 ( new_n325_, new_n319_, new_n324_ );
not g188 ( new_n326_, new_n324_ );
nand g189 ( new_n327_, new_n317_, new_n318_, new_n326_ );
and g190 ( new_n328_, new_n325_, new_n327_ );
not g191 ( new_n329_, new_n267_ );
nand g192 ( new_n330_, new_n298_, new_n329_ );
nand g193 ( new_n331_, new_n295_, new_n267_, new_n297_ );
nand g194 ( new_n332_, new_n330_, new_n331_ );
nand g195 ( new_n333_, new_n332_, keyIn_0_9 );
not g196 ( new_n334_, keyIn_0_9 );
nand g197 ( new_n335_, new_n330_, new_n334_, new_n331_ );
nand g198 ( new_n336_, new_n333_, new_n335_ );
nand g199 ( new_n337_, N132, N137 );
nand g200 ( new_n338_, new_n336_, new_n337_ );
nand g201 ( new_n339_, new_n333_, N132, N137, new_n335_ );
nand g202 ( new_n340_, new_n338_, new_n339_ );
nand g203 ( new_n341_, new_n340_, keyIn_0_23 );
not g204 ( new_n342_, keyIn_0_23 );
nand g205 ( new_n343_, new_n338_, new_n342_, new_n339_ );
nand g206 ( new_n344_, new_n341_, new_n343_ );
xor g207 ( new_n345_, N13, N29 );
xnor g208 ( new_n346_, new_n345_, keyIn_0_14 );
xor g209 ( new_n347_, N45, N61 );
xnor g210 ( new_n348_, new_n346_, new_n347_ );
not g211 ( new_n349_, new_n348_ );
nand g212 ( new_n350_, new_n344_, new_n349_ );
nand g213 ( new_n351_, new_n341_, new_n343_, new_n348_ );
nand g214 ( new_n352_, new_n350_, new_n351_ );
not g215 ( new_n353_, keyIn_0_26 );
nand g216 ( new_n354_, new_n264_, new_n305_ );
nand g217 ( new_n355_, new_n303_, new_n261_, new_n263_ );
nand g218 ( new_n356_, new_n354_, new_n355_ );
nand g219 ( new_n357_, N131, N137 );
nand g220 ( new_n358_, new_n356_, new_n357_ );
nand g221 ( new_n359_, new_n354_, N131, new_n355_, N137 );
nand g222 ( new_n360_, new_n358_, new_n359_ );
xor g223 ( new_n361_, N9, N25 );
xnor g224 ( new_n362_, N41, N57 );
xor g225 ( new_n363_, new_n361_, new_n362_ );
nand g226 ( new_n364_, new_n360_, new_n363_ );
not g227 ( new_n365_, new_n363_ );
nand g228 ( new_n366_, new_n358_, new_n359_, new_n365_ );
nand g229 ( new_n367_, new_n364_, new_n366_ );
nand g230 ( new_n368_, new_n367_, keyIn_0_24 );
not g231 ( new_n369_, keyIn_0_24 );
nand g232 ( new_n370_, new_n364_, new_n369_, new_n366_ );
nand g233 ( new_n371_, new_n368_, new_n370_ );
nand g234 ( new_n372_, new_n371_, new_n353_ );
nand g235 ( new_n373_, new_n368_, keyIn_0_26, new_n370_ );
nand g236 ( new_n374_, new_n372_, new_n373_ );
nand g237 ( new_n375_, new_n328_, new_n279_, new_n352_, new_n374_ );
nand g238 ( new_n376_, new_n375_, new_n280_ );
not g239 ( new_n377_, new_n279_ );
nand g240 ( new_n378_, new_n325_, new_n327_ );
nor g241 ( new_n379_, new_n378_, new_n377_ );
nand g242 ( new_n380_, new_n379_, keyIn_0_36, new_n352_, new_n374_ );
nand g243 ( new_n381_, new_n376_, new_n380_ );
not g244 ( new_n382_, new_n371_ );
xnor g245 ( new_n383_, new_n279_, keyIn_0_25 );
nand g246 ( new_n384_, new_n328_, new_n382_, new_n383_ );
nor g247 ( new_n385_, new_n382_, new_n279_ );
nand g248 ( new_n386_, new_n385_, new_n378_ );
nand g249 ( new_n387_, new_n384_, new_n386_ );
nand g250 ( new_n388_, new_n387_, new_n352_ );
not g251 ( new_n389_, new_n352_ );
nand g252 ( new_n390_, new_n389_, new_n328_, new_n385_ );
nand g253 ( new_n391_, new_n381_, new_n388_, new_n390_ );
and g254 ( new_n392_, new_n391_, new_n279_ );
nand g255 ( new_n393_, new_n392_, new_n246_ );
xnor g256 ( new_n394_, new_n393_, new_n138_ );
xnor g257 ( N724, new_n394_, N1 );
and g258 ( new_n396_, new_n391_, new_n378_ );
nand g259 ( new_n397_, new_n396_, new_n246_ );
xnor g260 ( new_n398_, new_n397_, keyIn_0_42 );
xnor g261 ( N725, new_n398_, N5 );
and g262 ( new_n400_, new_n391_, new_n382_ );
nand g263 ( new_n401_, new_n400_, new_n246_ );
xnor g264 ( N726, new_n401_, N9 );
and g265 ( new_n403_, new_n391_, new_n389_ );
nand g266 ( new_n404_, new_n403_, new_n246_ );
xnor g267 ( N727, new_n404_, N13 );
nor g268 ( new_n406_, new_n228_, new_n180_, new_n244_ );
nand g269 ( new_n407_, new_n392_, new_n406_ );
xnor g270 ( new_n408_, new_n407_, N17 );
xnor g271 ( N728, new_n408_, keyIn_0_54 );
nand g272 ( new_n410_, new_n396_, new_n406_ );
xnor g273 ( new_n411_, new_n410_, N21 );
xnor g274 ( N729, new_n411_, keyIn_0_55 );
nand g275 ( new_n413_, new_n400_, new_n406_ );
xnor g276 ( N730, new_n413_, N25 );
not g277 ( new_n415_, keyIn_0_43 );
nand g278 ( new_n416_, new_n403_, new_n406_ );
xnor g279 ( new_n417_, new_n416_, new_n415_ );
xnor g280 ( N731, new_n417_, N29 );
not g281 ( new_n419_, new_n203_ );
nor g282 ( new_n420_, new_n419_, new_n225_, new_n245_ );
and g283 ( new_n421_, new_n420_, new_n180_ );
nand g284 ( new_n422_, new_n392_, new_n421_ );
xnor g285 ( new_n423_, new_n422_, N33 );
xnor g286 ( N732, new_n423_, keyIn_0_56 );
nand g287 ( new_n425_, new_n396_, new_n421_ );
xnor g288 ( new_n426_, new_n425_, new_n140_ );
xnor g289 ( N733, new_n426_, keyIn_0_57 );
not g290 ( new_n428_, keyIn_0_44 );
nand g291 ( new_n429_, new_n400_, new_n421_ );
xnor g292 ( new_n430_, new_n429_, new_n428_ );
xnor g293 ( N734, new_n430_, N41 );
not g294 ( new_n432_, keyIn_0_58 );
nand g295 ( new_n433_, new_n391_, new_n389_, new_n421_ );
xnor g296 ( new_n434_, new_n433_, keyIn_0_45 );
nand g297 ( new_n435_, new_n434_, N45 );
not g298 ( new_n436_, N45 );
nand g299 ( new_n437_, new_n433_, keyIn_0_45 );
or g300 ( new_n438_, new_n433_, keyIn_0_45 );
nand g301 ( new_n439_, new_n438_, new_n436_, new_n437_ );
nand g302 ( new_n440_, new_n435_, new_n439_ );
nand g303 ( new_n441_, new_n440_, new_n432_ );
nand g304 ( new_n442_, new_n435_, keyIn_0_58, new_n439_ );
nand g305 ( N735, new_n441_, new_n442_ );
not g306 ( new_n444_, keyIn_0_59 );
not g307 ( new_n445_, N49 );
not g308 ( new_n446_, keyIn_0_39 );
nand g309 ( new_n447_, new_n181_, keyIn_0_27 );
or g310 ( new_n448_, new_n181_, keyIn_0_27 );
nor g311 ( new_n449_, new_n244_, new_n225_ );
and g312 ( new_n450_, new_n203_, new_n448_, new_n447_, new_n449_ );
nand g313 ( new_n451_, new_n391_, new_n450_ );
nand g314 ( new_n452_, new_n451_, new_n446_ );
nand g315 ( new_n453_, new_n391_, keyIn_0_39, new_n450_ );
nand g316 ( new_n454_, new_n452_, new_n453_ );
nand g317 ( new_n455_, new_n454_, new_n279_ );
nand g318 ( new_n456_, new_n455_, new_n445_ );
nand g319 ( new_n457_, new_n454_, N49, new_n279_ );
nand g320 ( new_n458_, new_n456_, new_n457_ );
nand g321 ( new_n459_, new_n458_, new_n444_ );
nand g322 ( new_n460_, new_n456_, keyIn_0_59, new_n457_ );
nand g323 ( N736, new_n459_, new_n460_ );
not g324 ( new_n462_, N53 );
not g325 ( new_n463_, keyIn_0_46 );
nand g326 ( new_n464_, new_n454_, new_n378_ );
nand g327 ( new_n465_, new_n464_, new_n463_ );
nand g328 ( new_n466_, new_n454_, keyIn_0_46, new_n378_ );
nand g329 ( new_n467_, new_n465_, new_n466_ );
nand g330 ( new_n468_, new_n467_, new_n462_ );
nand g331 ( new_n469_, new_n465_, N53, new_n466_ );
nand g332 ( N737, new_n468_, new_n469_ );
nand g333 ( new_n471_, new_n454_, new_n382_ );
xnor g334 ( N738, new_n471_, N57 );
nand g335 ( new_n473_, new_n454_, new_n389_ );
xnor g336 ( N739, new_n473_, N61 );
not g337 ( new_n475_, keyIn_0_37 );
not g338 ( new_n476_, keyIn_0_31 );
nand g339 ( new_n477_, new_n177_, new_n476_, new_n179_ );
nand g340 ( new_n478_, new_n180_, keyIn_0_31 );
nand g341 ( new_n479_, new_n478_, new_n475_, new_n420_, new_n477_ );
not g342 ( new_n480_, keyIn_0_32 );
nand g343 ( new_n481_, new_n180_, new_n480_ );
nand g344 ( new_n482_, new_n177_, keyIn_0_32, new_n179_ );
nand g345 ( new_n483_, new_n481_, new_n482_ );
xor g346 ( new_n484_, new_n244_, keyIn_0_33 );
nand g347 ( new_n485_, new_n483_, new_n227_, new_n484_ );
xnor g348 ( new_n486_, new_n244_, keyIn_0_30 );
not g349 ( new_n487_, keyIn_0_29 );
xnor g350 ( new_n488_, new_n225_, new_n487_ );
nand g351 ( new_n489_, new_n180_, new_n486_, new_n419_, new_n488_ );
nand g352 ( new_n490_, new_n203_, keyIn_0_28 );
not g353 ( new_n491_, keyIn_0_28 );
nand g354 ( new_n492_, new_n200_, new_n491_, new_n202_ );
nand g355 ( new_n493_, new_n490_, new_n492_ );
nand g356 ( new_n494_, new_n493_, new_n177_, new_n179_, new_n449_ );
and g357 ( new_n495_, new_n489_, new_n494_ );
and g358 ( new_n496_, new_n485_, new_n495_, new_n479_ );
not g359 ( new_n497_, keyIn_0_38 );
nand g360 ( new_n498_, new_n478_, new_n420_, new_n477_ );
nand g361 ( new_n499_, new_n498_, keyIn_0_37 );
and g362 ( new_n500_, new_n499_, new_n497_ );
nand g363 ( new_n501_, new_n496_, new_n500_ );
nand g364 ( new_n502_, new_n485_, new_n499_, new_n495_, new_n479_ );
nand g365 ( new_n503_, new_n502_, keyIn_0_38 );
nand g366 ( new_n504_, new_n352_, new_n382_ );
nor g367 ( new_n505_, new_n504_, new_n377_, new_n378_ );
nand g368 ( new_n506_, new_n501_, new_n503_, new_n505_ );
nand g369 ( new_n507_, new_n506_, keyIn_0_40 );
not g370 ( new_n508_, keyIn_0_40 );
nand g371 ( new_n509_, new_n501_, new_n503_, new_n508_, new_n505_ );
nand g372 ( new_n510_, new_n507_, new_n509_ );
nand g373 ( new_n511_, new_n510_, new_n225_ );
nand g374 ( new_n512_, new_n511_, keyIn_0_47 );
not g375 ( new_n513_, keyIn_0_47 );
nand g376 ( new_n514_, new_n510_, new_n513_, new_n225_ );
nand g377 ( new_n515_, new_n512_, new_n514_ );
nand g378 ( new_n516_, new_n515_, new_n248_ );
nand g379 ( new_n517_, new_n512_, N65, new_n514_ );
nand g380 ( N740, new_n516_, new_n517_ );
not g381 ( new_n519_, keyIn_0_48 );
nand g382 ( new_n520_, new_n510_, new_n203_ );
nand g383 ( new_n521_, new_n520_, new_n519_ );
nand g384 ( new_n522_, new_n510_, keyIn_0_48, new_n203_ );
nand g385 ( new_n523_, new_n521_, new_n522_ );
nand g386 ( new_n524_, new_n523_, N69 );
nand g387 ( new_n525_, new_n521_, new_n249_, new_n522_ );
nand g388 ( N741, new_n524_, new_n525_ );
nand g389 ( new_n527_, new_n510_, new_n180_ );
xnor g390 ( N742, new_n527_, N73 );
nand g391 ( new_n529_, new_n510_, new_n245_ );
nand g392 ( new_n530_, new_n529_, N77 );
not g393 ( new_n531_, N77 );
nand g394 ( new_n532_, new_n510_, new_n531_, new_n245_ );
nand g395 ( new_n533_, new_n530_, new_n532_ );
nand g396 ( new_n534_, new_n533_, keyIn_0_60 );
not g397 ( new_n535_, keyIn_0_60 );
nand g398 ( new_n536_, new_n530_, new_n535_, new_n532_ );
nand g399 ( N743, new_n534_, new_n536_ );
and g400 ( new_n538_, new_n501_, new_n503_ );
nor g401 ( new_n539_, new_n378_, keyIn_0_34 );
and g402 ( new_n540_, new_n378_, keyIn_0_34 );
nand g403 ( new_n541_, new_n371_, new_n279_ );
nor g404 ( new_n542_, new_n540_, new_n539_, new_n352_, new_n541_ );
nand g405 ( new_n543_, new_n538_, new_n542_ );
not g406 ( new_n544_, new_n543_ );
nand g407 ( new_n545_, new_n544_, new_n225_ );
xnor g408 ( N744, new_n545_, N81 );
nand g409 ( new_n547_, new_n544_, new_n203_ );
nand g410 ( new_n548_, new_n547_, keyIn_0_49 );
or g411 ( new_n549_, new_n543_, keyIn_0_49, new_n419_ );
nand g412 ( new_n550_, new_n548_, new_n549_ );
nand g413 ( new_n551_, new_n550_, N85 );
not g414 ( new_n552_, N85 );
nand g415 ( new_n553_, new_n548_, new_n552_, new_n549_ );
nand g416 ( N745, new_n551_, new_n553_ );
nand g417 ( new_n555_, new_n544_, new_n180_ );
nand g418 ( new_n556_, new_n555_, N89 );
or g419 ( new_n557_, new_n543_, N89, new_n181_ );
nand g420 ( new_n558_, new_n556_, new_n557_ );
nand g421 ( new_n559_, new_n558_, keyIn_0_61 );
not g422 ( new_n560_, keyIn_0_61 );
nand g423 ( new_n561_, new_n556_, new_n560_, new_n557_ );
nand g424 ( N746, new_n559_, new_n561_ );
nand g425 ( new_n563_, new_n544_, new_n245_ );
xnor g426 ( N747, new_n563_, N93 );
xor g427 ( new_n565_, new_n279_, keyIn_0_35 );
nor g428 ( new_n566_, new_n504_, new_n565_, new_n328_ );
nand g429 ( new_n567_, new_n538_, new_n566_ );
not g430 ( new_n568_, new_n567_ );
nand g431 ( new_n569_, new_n568_, new_n225_ );
xnor g432 ( N748, new_n569_, N97 );
nand g433 ( new_n571_, new_n568_, new_n203_ );
nand g434 ( new_n572_, new_n571_, keyIn_0_50 );
or g435 ( new_n573_, new_n567_, keyIn_0_50, new_n419_ );
nand g436 ( new_n574_, new_n572_, new_n573_ );
nand g437 ( new_n575_, new_n574_, N101 );
not g438 ( new_n576_, N101 );
nand g439 ( new_n577_, new_n572_, new_n576_, new_n573_ );
nand g440 ( N749, new_n575_, new_n577_ );
nand g441 ( new_n579_, new_n568_, new_n180_ );
xnor g442 ( N750, new_n579_, N105 );
nand g443 ( new_n581_, new_n568_, new_n245_ );
xnor g444 ( N751, new_n581_, N109 );
nand g445 ( new_n583_, new_n389_, new_n378_, new_n385_ );
nor g446 ( new_n584_, new_n583_, new_n226_ );
nand g447 ( new_n585_, new_n538_, new_n584_ );
xnor g448 ( N752, new_n585_, N113 );
nor g449 ( new_n587_, new_n583_, new_n419_ );
nand g450 ( new_n588_, new_n538_, new_n587_ );
xnor g451 ( new_n589_, new_n588_, keyIn_0_51 );
xor g452 ( N753, new_n589_, N117 );
nor g453 ( new_n591_, new_n583_, new_n181_ );
nand g454 ( new_n592_, new_n538_, keyIn_0_52, new_n591_ );
not g455 ( new_n593_, keyIn_0_52 );
nand g456 ( new_n594_, new_n501_, new_n503_, new_n591_ );
nand g457 ( new_n595_, new_n594_, new_n593_ );
nand g458 ( new_n596_, new_n592_, new_n595_ );
nand g459 ( new_n597_, new_n596_, new_n285_ );
nand g460 ( new_n598_, new_n592_, N121, new_n595_ );
nand g461 ( new_n599_, new_n597_, new_n598_ );
nand g462 ( new_n600_, new_n599_, keyIn_0_62 );
not g463 ( new_n601_, keyIn_0_62 );
nand g464 ( new_n602_, new_n597_, new_n601_, new_n598_ );
nand g465 ( N754, new_n600_, new_n602_ );
not g466 ( new_n604_, keyIn_0_63 );
nor g467 ( new_n605_, new_n583_, new_n244_ );
nand g468 ( new_n606_, new_n538_, keyIn_0_53, new_n605_ );
not g469 ( new_n607_, keyIn_0_53 );
nand g470 ( new_n608_, new_n501_, new_n503_, new_n605_ );
nand g471 ( new_n609_, new_n608_, new_n607_ );
nand g472 ( new_n610_, new_n606_, new_n609_ );
nand g473 ( new_n611_, new_n610_, new_n286_ );
nand g474 ( new_n612_, new_n606_, N125, new_n609_ );
nand g475 ( new_n613_, new_n611_, new_n612_ );
nand g476 ( new_n614_, new_n613_, new_n604_ );
nand g477 ( new_n615_, new_n611_, keyIn_0_63, new_n612_ );
nand g478 ( N755, new_n614_, new_n615_ );
endmodule