module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n595_, new_n614_, new_n445_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n421_, new_n620_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n170_, new_n246_, new_n682_, new_n679_, new_n266_, new_n667_, new_n367_, new_n542_, new_n548_, new_n669_, new_n220_, new_n419_, new_n624_, new_n534_, new_n637_, new_n214_, new_n489_, new_n424_, new_n602_, new_n188_, new_n695_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n649_, new_n678_, new_n462_, new_n603_, new_n564_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n626_, new_n152_, new_n157_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n272_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n655_, new_n167_, new_n385_, new_n478_, new_n694_, new_n461_, new_n297_, new_n361_, new_n565_, new_n683_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n622_, new_n629_, new_n321_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n650_, new_n206_, new_n254_, new_n429_, new_n353_, new_n432_, new_n506_, new_n680_, new_n256_, new_n452_, new_n381_, new_n656_, new_n388_, new_n508_, new_n194_, new_n483_, new_n394_, new_n299_, new_n142_, new_n139_, new_n657_, new_n652_, new_n314_, new_n582_, new_n363_, new_n165_, new_n441_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n187_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n399_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n628_, new_n162_, new_n409_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n688_, new_n155_, new_n384_, new_n410_, new_n543_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n232_, new_n258_, new_n176_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n654_, new_n227_, new_n690_, new_n416_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n693_, new_n130_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n138_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n562_, new_n578_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n379_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n520_, new_n125_, new_n145_, new_n253_, new_n403_, new_n475_, new_n237_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n605_, new_n182_, new_n407_, new_n666_, new_n625_, new_n151_, new_n513_, new_n592_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n522_, new_n588_, new_n428_, new_n199_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n191_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n131_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n662_, new_n440_, new_n122_, new_n531_, new_n593_, new_n252_, new_n585_, new_n160_, new_n312_, new_n535_, new_n372_, new_n242_, new_n503_, new_n527_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n134_, new_n651_, new_n433_, new_n435_, new_n265_, new_n687_, new_n370_, new_n689_, new_n278_, new_n304_, new_n523_, new_n638_, new_n550_, new_n217_, new_n269_, new_n512_, new_n129_, new_n644_, new_n599_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n594_, new_n561_, new_n495_, new_n431_, new_n196_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n627_, new_n195_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n358_, new_n348_, new_n610_, new_n159_, new_n322_, new_n228_, new_n545_, new_n611_, new_n289_, new_n425_, new_n175_, new_n226_, new_n185_, new_n373_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n618_, new_n120_, new_n521_, new_n406_, new_n356_, new_n647_, new_n536_, new_n464_, new_n204_, new_n181_, new_n135_, new_n573_, new_n405_;

not g000 ( new_n119_, N75 );
nand g001 ( new_n120_, N29, N42 );
nor g002 ( N388, new_n120_, new_n119_ );
not g003 ( new_n122_, N80 );
nand g004 ( new_n123_, N29, N36 );
nor g005 ( N389, new_n123_, new_n122_ );
not g006 ( new_n125_, N42 );
nor g007 ( N390, new_n123_, new_n125_ );
nand g008 ( new_n127_, N85, N86 );
not g009 ( N391, new_n127_ );
not g010 ( new_n129_, N17 );
nand g011 ( new_n130_, N1, N8 );
not g012 ( new_n131_, new_n130_ );
nand g013 ( new_n132_, new_n131_, N13 );
nor g014 ( N418, new_n132_, new_n129_ );
not g015 ( new_n134_, N390 );
nor g016 ( new_n135_, new_n134_, keyIn_0_0 );
nand g017 ( new_n136_, new_n134_, keyIn_0_0 );
not g018 ( new_n137_, new_n136_ );
nor g019 ( new_n138_, new_n137_, new_n135_ );
not g020 ( new_n139_, new_n138_ );
nand g021 ( new_n140_, N1, N26 );
nand g022 ( new_n141_, N13, N17 );
nor g023 ( new_n142_, new_n140_, new_n141_ );
nand g024 ( N419, new_n139_, new_n142_ );
nand g025 ( new_n144_, N59, N75 );
not g026 ( new_n145_, new_n144_ );
nand g027 ( N420, new_n145_, N80 );
nand g028 ( new_n147_, N36, N59 );
not g029 ( new_n148_, new_n147_ );
nand g030 ( N421, new_n148_, N80 );
nand g031 ( N422, new_n148_, N42 );
not g032 ( new_n151_, N90 );
nor g033 ( new_n152_, N87, N88 );
nor g034 ( N423, new_n152_, new_n151_ );
nand g035 ( N446, new_n138_, new_n142_ );
not g036 ( new_n155_, N51 );
nor g037 ( N447, new_n140_, new_n155_ );
not g038 ( new_n157_, N55 );
nor g039 ( new_n158_, new_n132_, new_n157_ );
not g040 ( new_n159_, new_n158_ );
nand g041 ( new_n160_, N29, N68 );
nand g042 ( new_n161_, new_n160_, keyIn_0_1 );
not g043 ( new_n162_, keyIn_0_1 );
not g044 ( new_n163_, new_n160_ );
nand g045 ( new_n164_, new_n163_, new_n162_ );
nand g046 ( new_n165_, new_n164_, new_n161_ );
nor g047 ( N448, new_n159_, new_n165_ );
not g048 ( new_n167_, N74 );
nand g049 ( new_n168_, N59, N68 );
nor g050 ( new_n169_, new_n159_, new_n168_ );
not g051 ( new_n170_, new_n169_ );
nor g052 ( N449, new_n170_, new_n167_ );
not g053 ( new_n172_, N89 );
nor g054 ( N450, new_n152_, new_n172_ );
not g055 ( new_n174_, keyIn_0_7 );
nand g056 ( new_n175_, N101, N106 );
nor g057 ( new_n176_, new_n175_, keyIn_0_2 );
nand g058 ( new_n177_, new_n175_, keyIn_0_2 );
not g059 ( new_n178_, N101 );
not g060 ( new_n179_, N106 );
nand g061 ( new_n180_, new_n178_, new_n179_ );
nand g062 ( new_n181_, new_n177_, new_n180_ );
nor g063 ( new_n182_, new_n181_, new_n176_ );
not g064 ( new_n183_, new_n182_ );
not g065 ( new_n184_, N91 );
nor g066 ( new_n185_, new_n184_, N96 );
not g067 ( new_n186_, N96 );
nor g068 ( new_n187_, new_n186_, N91 );
nor g069 ( new_n188_, new_n185_, new_n187_ );
nor g070 ( new_n189_, new_n183_, new_n188_ );
not g071 ( new_n190_, new_n189_ );
nor g072 ( new_n191_, new_n190_, new_n174_ );
nand g073 ( new_n192_, new_n190_, new_n174_ );
nand g074 ( new_n193_, new_n183_, new_n188_ );
nand g075 ( new_n194_, new_n192_, new_n193_ );
nor g076 ( new_n195_, new_n194_, new_n191_ );
nor g077 ( new_n196_, new_n195_, N130 );
not g078 ( new_n197_, new_n196_ );
nor g079 ( new_n198_, new_n197_, keyIn_0_10 );
nand g080 ( new_n199_, new_n197_, keyIn_0_10 );
not g081 ( new_n200_, new_n199_ );
nor g082 ( new_n201_, new_n200_, new_n198_ );
nand g083 ( new_n202_, new_n195_, N130 );
nand g084 ( new_n203_, new_n202_, keyIn_0_9 );
not g085 ( new_n204_, new_n203_ );
nor g086 ( new_n205_, new_n202_, keyIn_0_9 );
nor g087 ( new_n206_, new_n204_, new_n205_ );
nor g088 ( new_n207_, new_n201_, new_n206_ );
not g089 ( new_n208_, new_n207_ );
nand g090 ( new_n209_, N111, N116 );
not g091 ( new_n210_, new_n209_ );
nor g092 ( new_n211_, N111, N116 );
nor g093 ( new_n212_, new_n210_, new_n211_ );
nand g094 ( new_n213_, N121, N126 );
not g095 ( new_n214_, new_n213_ );
nor g096 ( new_n215_, N121, N126 );
nor g097 ( new_n216_, new_n214_, new_n215_ );
nor g098 ( new_n217_, new_n212_, new_n216_ );
nand g099 ( new_n218_, new_n212_, new_n216_ );
not g100 ( new_n219_, new_n218_ );
nor g101 ( new_n220_, new_n219_, new_n217_ );
not g102 ( new_n221_, new_n220_ );
nand g103 ( new_n222_, new_n221_, N135 );
not g104 ( new_n223_, new_n222_ );
nor g105 ( new_n224_, new_n221_, N135 );
nor g106 ( new_n225_, new_n223_, new_n224_ );
not g107 ( new_n226_, new_n225_ );
nand g108 ( new_n227_, new_n208_, new_n226_ );
nand g109 ( new_n228_, new_n207_, new_n225_ );
nand g110 ( N767, new_n227_, new_n228_ );
not g111 ( new_n230_, keyIn_0_12 );
not g112 ( new_n231_, N159 );
nor g113 ( new_n232_, new_n231_, N165 );
not g114 ( new_n233_, N165 );
nor g115 ( new_n234_, new_n233_, N159 );
nor g116 ( new_n235_, new_n232_, new_n234_ );
nand g117 ( new_n236_, N171, N177 );
not g118 ( new_n237_, new_n236_ );
nor g119 ( new_n238_, N171, N177 );
nor g120 ( new_n239_, new_n237_, new_n238_ );
nor g121 ( new_n240_, new_n235_, new_n239_ );
nand g122 ( new_n241_, new_n235_, new_n239_ );
not g123 ( new_n242_, new_n241_ );
nor g124 ( new_n243_, new_n242_, new_n240_ );
not g125 ( new_n244_, new_n243_ );
nor g126 ( new_n245_, new_n244_, N130 );
not g127 ( new_n246_, new_n245_ );
nor g128 ( new_n247_, new_n246_, new_n230_ );
nor g129 ( new_n248_, new_n245_, keyIn_0_12 );
not g130 ( new_n249_, keyIn_0_15 );
nand g131 ( new_n250_, new_n244_, N130 );
nand g132 ( new_n251_, new_n250_, new_n249_ );
nor g133 ( new_n252_, new_n248_, new_n251_ );
not g134 ( new_n253_, new_n252_ );
nor g135 ( new_n254_, new_n253_, new_n247_ );
not g136 ( new_n255_, new_n254_ );
not g137 ( new_n256_, N207 );
not g138 ( new_n257_, keyIn_0_5 );
nand g139 ( new_n258_, N195, N201 );
not g140 ( new_n259_, new_n258_ );
nor g141 ( new_n260_, N195, N201 );
nor g142 ( new_n261_, new_n259_, new_n260_ );
not g143 ( new_n262_, new_n261_ );
nand g144 ( new_n263_, new_n262_, keyIn_0_6 );
nand g145 ( new_n264_, new_n263_, new_n257_ );
nand g146 ( new_n265_, N183, N189 );
not g147 ( new_n266_, new_n265_ );
nor g148 ( new_n267_, N183, N189 );
nor g149 ( new_n268_, new_n266_, new_n267_ );
nand g150 ( new_n269_, new_n264_, new_n268_ );
not g151 ( new_n270_, new_n268_ );
nand g152 ( new_n271_, new_n270_, new_n257_ );
nand g153 ( new_n272_, new_n271_, keyIn_0_6 );
nand g154 ( new_n273_, new_n272_, new_n261_ );
nand g155 ( new_n274_, new_n269_, new_n273_ );
nor g156 ( new_n275_, new_n274_, new_n256_ );
nand g157 ( new_n276_, new_n274_, new_n256_ );
not g158 ( new_n277_, new_n276_ );
nor g159 ( new_n278_, new_n277_, new_n275_ );
not g160 ( new_n279_, new_n278_ );
nand g161 ( new_n280_, new_n255_, new_n279_ );
nand g162 ( new_n281_, new_n254_, new_n278_ );
nand g163 ( N768, new_n280_, new_n281_ );
not g164 ( new_n283_, N126 );
nand g165 ( new_n284_, N17, N51 );
nor g166 ( new_n285_, new_n130_, new_n284_ );
nor g167 ( new_n286_, new_n285_, keyIn_0_4 );
nand g168 ( new_n287_, new_n285_, keyIn_0_4 );
nand g169 ( new_n288_, new_n145_, N42 );
nand g170 ( new_n289_, new_n287_, new_n288_ );
nor g171 ( new_n290_, new_n289_, new_n286_ );
not g172 ( new_n291_, N447 );
nand g173 ( new_n292_, N17, N42 );
nor g174 ( new_n293_, N17, N42 );
nand g175 ( new_n294_, N59, N156 );
nor g176 ( new_n295_, new_n293_, new_n294_ );
nand g177 ( new_n296_, new_n295_, new_n292_ );
nor g178 ( new_n297_, new_n296_, new_n291_ );
nor g179 ( new_n298_, new_n290_, new_n297_ );
nor g180 ( new_n299_, new_n298_, new_n283_ );
nand g181 ( new_n300_, new_n299_, keyIn_0_11 );
not g182 ( new_n301_, keyIn_0_11 );
not g183 ( new_n302_, new_n286_ );
not g184 ( new_n303_, new_n289_ );
nand g185 ( new_n304_, new_n303_, new_n302_ );
not g186 ( new_n305_, new_n297_ );
nand g187 ( new_n306_, new_n304_, new_n305_ );
nand g188 ( new_n307_, new_n306_, N126 );
nand g189 ( new_n308_, new_n307_, new_n301_ );
nand g190 ( new_n309_, new_n308_, new_n300_ );
nand g191 ( new_n310_, new_n294_, N17 );
not g192 ( new_n311_, new_n310_ );
nand g193 ( new_n312_, new_n311_, N447 );
nand g194 ( new_n313_, new_n312_, N1 );
nand g195 ( new_n314_, new_n313_, N153 );
nand g196 ( new_n315_, N29, N75 );
nor g197 ( new_n316_, new_n315_, new_n122_ );
nand g198 ( new_n317_, N447, new_n316_ );
not g199 ( new_n318_, new_n317_ );
nor g200 ( new_n319_, new_n157_, N268 );
nand g201 ( new_n320_, new_n318_, new_n319_ );
nand g202 ( new_n321_, new_n314_, new_n320_ );
not g203 ( new_n322_, new_n321_ );
nand g204 ( new_n323_, new_n309_, new_n322_ );
nand g205 ( new_n324_, new_n323_, N201 );
not g206 ( new_n325_, new_n324_ );
nor g207 ( new_n326_, new_n323_, N201 );
nor g208 ( new_n327_, new_n325_, new_n326_ );
nand g209 ( new_n328_, new_n327_, N261 );
not g210 ( new_n329_, N219 );
nor g211 ( new_n330_, new_n327_, N261 );
nor g212 ( new_n331_, new_n330_, new_n329_ );
nand g213 ( new_n332_, new_n331_, new_n328_ );
nand g214 ( new_n333_, new_n327_, N228 );
not g215 ( new_n334_, N237 );
nor g216 ( new_n335_, new_n324_, new_n334_ );
not g217 ( new_n336_, N73 );
nand g218 ( new_n337_, N42, N72 );
nor g219 ( new_n338_, new_n337_, new_n336_ );
nand g220 ( new_n339_, new_n169_, new_n338_ );
not g221 ( new_n340_, new_n339_ );
nand g222 ( new_n341_, new_n340_, N201 );
nand g223 ( new_n342_, N121, N210 );
nand g224 ( new_n343_, new_n341_, new_n342_ );
nor g225 ( new_n344_, new_n335_, new_n343_ );
nand g226 ( new_n345_, new_n333_, new_n344_ );
nand g227 ( new_n346_, new_n323_, N246 );
nand g228 ( new_n347_, N255, N267 );
nand g229 ( new_n348_, new_n346_, new_n347_ );
nand g230 ( new_n349_, new_n348_, keyIn_0_19 );
not g231 ( new_n350_, keyIn_0_19 );
not g232 ( new_n351_, new_n348_ );
nand g233 ( new_n352_, new_n351_, new_n350_ );
nand g234 ( new_n353_, new_n352_, new_n349_ );
nor g235 ( new_n354_, new_n345_, new_n353_ );
nand g236 ( N850, new_n332_, new_n354_ );
not g237 ( new_n356_, N183 );
nand g238 ( new_n357_, new_n306_, N111 );
not g239 ( new_n358_, new_n357_ );
nand g240 ( new_n359_, new_n313_, N143 );
nand g241 ( new_n360_, new_n359_, new_n320_ );
nor g242 ( new_n361_, new_n358_, new_n360_ );
nor g243 ( new_n362_, new_n361_, new_n356_ );
not g244 ( new_n363_, new_n362_ );
not g245 ( new_n364_, N261 );
nor g246 ( new_n365_, new_n326_, new_n364_ );
nor g247 ( new_n366_, new_n365_, new_n325_ );
not g248 ( new_n367_, keyIn_0_14 );
nand g249 ( new_n368_, new_n306_, N121 );
nand g250 ( new_n369_, new_n313_, N149 );
nand g251 ( new_n370_, new_n369_, new_n320_ );
not g252 ( new_n371_, new_n370_ );
nand g253 ( new_n372_, new_n368_, new_n371_ );
not g254 ( new_n373_, new_n372_ );
nor g255 ( new_n374_, new_n373_, new_n367_ );
nor g256 ( new_n375_, new_n372_, keyIn_0_14 );
nor g257 ( new_n376_, new_n374_, new_n375_ );
not g258 ( new_n377_, new_n376_ );
nor g259 ( new_n378_, new_n377_, N195 );
nor g260 ( new_n379_, new_n366_, new_n378_ );
not g261 ( new_n380_, N189 );
nand g262 ( new_n381_, new_n306_, N116 );
nand g263 ( new_n382_, new_n313_, N146 );
nand g264 ( new_n383_, new_n382_, new_n320_ );
not g265 ( new_n384_, new_n383_ );
nand g266 ( new_n385_, new_n381_, new_n384_ );
nand g267 ( new_n386_, new_n385_, keyIn_0_13 );
not g268 ( new_n387_, keyIn_0_13 );
not g269 ( new_n388_, N116 );
nor g270 ( new_n389_, new_n298_, new_n388_ );
nor g271 ( new_n390_, new_n389_, new_n383_ );
nand g272 ( new_n391_, new_n390_, new_n387_ );
nand g273 ( new_n392_, new_n391_, new_n386_ );
nor g274 ( new_n393_, new_n382_, new_n387_ );
nor g275 ( new_n394_, new_n392_, new_n393_ );
not g276 ( new_n395_, new_n394_ );
nand g277 ( new_n396_, new_n395_, new_n380_ );
nand g278 ( new_n397_, new_n379_, new_n396_ );
not g279 ( new_n398_, keyIn_0_24 );
nand g280 ( new_n399_, new_n394_, N189 );
nand g281 ( new_n400_, new_n399_, keyIn_0_22 );
nand g282 ( new_n401_, new_n400_, new_n398_ );
not g283 ( new_n402_, N195 );
nor g284 ( new_n403_, new_n376_, new_n402_ );
nand g285 ( new_n404_, new_n396_, new_n403_ );
nor g286 ( new_n405_, new_n399_, keyIn_0_22 );
not g287 ( new_n406_, new_n405_ );
nand g288 ( new_n407_, new_n406_, new_n404_ );
nor g289 ( new_n408_, new_n407_, new_n401_ );
nand g290 ( new_n409_, new_n408_, new_n397_ );
nand g291 ( new_n410_, new_n392_, new_n380_ );
nand g292 ( new_n411_, new_n379_, new_n410_ );
nand g293 ( new_n412_, new_n403_, new_n410_ );
nand g294 ( new_n413_, new_n412_, new_n400_ );
nor g295 ( new_n414_, new_n413_, new_n405_ );
nand g296 ( new_n415_, new_n411_, new_n414_ );
nand g297 ( new_n416_, new_n415_, keyIn_0_24 );
nand g298 ( new_n417_, new_n416_, new_n409_ );
not g299 ( new_n418_, keyIn_0_17 );
nand g300 ( new_n419_, new_n361_, new_n356_ );
nor g301 ( new_n420_, new_n419_, new_n418_ );
nand g302 ( new_n421_, new_n419_, new_n418_ );
not g303 ( new_n422_, new_n421_ );
nor g304 ( new_n423_, new_n422_, new_n420_ );
nand g305 ( new_n424_, new_n417_, new_n423_ );
not g306 ( new_n425_, new_n424_ );
nand g307 ( new_n426_, new_n425_, new_n363_ );
nand g308 ( new_n427_, new_n423_, new_n363_ );
not g309 ( new_n428_, new_n427_ );
nor g310 ( new_n429_, new_n417_, new_n428_ );
nor g311 ( new_n430_, new_n429_, new_n329_ );
nand g312 ( new_n431_, new_n426_, new_n430_ );
not g313 ( new_n432_, N228 );
nor g314 ( new_n433_, new_n427_, new_n432_ );
nor g315 ( new_n434_, new_n362_, keyIn_0_18 );
nand g316 ( new_n435_, new_n362_, keyIn_0_18 );
not g317 ( new_n436_, new_n435_ );
nor g318 ( new_n437_, new_n436_, new_n434_ );
nand g319 ( new_n438_, new_n437_, N237 );
not g320 ( new_n439_, N246 );
nor g321 ( new_n440_, new_n361_, new_n439_ );
nand g322 ( new_n441_, new_n340_, N183 );
nand g323 ( new_n442_, N106, N210 );
nand g324 ( new_n443_, new_n442_, keyIn_0_3 );
not g325 ( new_n444_, new_n443_ );
nor g326 ( new_n445_, new_n442_, keyIn_0_3 );
nor g327 ( new_n446_, new_n444_, new_n445_ );
nand g328 ( new_n447_, new_n441_, new_n446_ );
nor g329 ( new_n448_, new_n440_, new_n447_ );
nand g330 ( new_n449_, new_n438_, new_n448_ );
nor g331 ( new_n450_, new_n433_, new_n449_ );
nand g332 ( N863, new_n431_, new_n450_ );
nor g333 ( new_n452_, new_n379_, new_n403_ );
nor g334 ( new_n453_, new_n392_, new_n380_ );
not g335 ( new_n454_, new_n453_ );
nand g336 ( new_n455_, new_n396_, new_n454_ );
nor g337 ( new_n456_, new_n452_, new_n455_ );
nand g338 ( new_n457_, new_n452_, new_n455_ );
nand g339 ( new_n458_, new_n457_, N219 );
nor g340 ( new_n459_, new_n458_, new_n456_ );
nor g341 ( new_n460_, new_n455_, new_n432_ );
nor g342 ( new_n461_, new_n454_, new_n334_ );
nor g343 ( new_n462_, new_n395_, new_n439_ );
nor g344 ( new_n463_, new_n339_, new_n380_ );
nand g345 ( new_n464_, N111, N210 );
nand g346 ( new_n465_, N255, N259 );
nand g347 ( new_n466_, new_n464_, new_n465_ );
nor g348 ( new_n467_, new_n463_, new_n466_ );
not g349 ( new_n468_, new_n467_ );
nor g350 ( new_n469_, new_n462_, new_n468_ );
not g351 ( new_n470_, new_n469_ );
nor g352 ( new_n471_, new_n470_, new_n461_ );
not g353 ( new_n472_, new_n471_ );
nor g354 ( new_n473_, new_n472_, new_n460_ );
not g355 ( new_n474_, new_n473_ );
nor g356 ( new_n475_, new_n459_, new_n474_ );
not g357 ( new_n476_, new_n475_ );
nand g358 ( new_n477_, new_n476_, keyIn_0_27 );
not g359 ( new_n478_, keyIn_0_27 );
nand g360 ( new_n479_, new_n475_, new_n478_ );
nand g361 ( N864, new_n477_, new_n479_ );
nor g362 ( new_n481_, new_n378_, new_n403_ );
not g363 ( new_n482_, new_n481_ );
nor g364 ( new_n483_, new_n482_, new_n366_ );
not g365 ( new_n484_, new_n483_ );
nand g366 ( new_n485_, new_n484_, keyIn_0_25 );
not g367 ( new_n486_, keyIn_0_25 );
nand g368 ( new_n487_, new_n483_, new_n486_ );
nand g369 ( new_n488_, new_n485_, new_n487_ );
not g370 ( new_n489_, new_n366_ );
nor g371 ( new_n490_, new_n489_, new_n481_ );
nor g372 ( new_n491_, new_n490_, new_n329_ );
nand g373 ( new_n492_, new_n488_, new_n491_ );
nor g374 ( new_n493_, new_n482_, new_n432_ );
nand g375 ( new_n494_, new_n403_, N237 );
nand g376 ( new_n495_, new_n377_, N246 );
nor g377 ( new_n496_, new_n339_, new_n402_ );
nand g378 ( new_n497_, N116, N210 );
nand g379 ( new_n498_, N255, N260 );
nand g380 ( new_n499_, new_n497_, new_n498_ );
nor g381 ( new_n500_, new_n496_, new_n499_ );
nand g382 ( new_n501_, new_n495_, new_n500_ );
not g383 ( new_n502_, new_n501_ );
nand g384 ( new_n503_, new_n502_, new_n494_ );
nor g385 ( new_n504_, new_n493_, new_n503_ );
nand g386 ( new_n505_, new_n492_, new_n504_ );
nand g387 ( new_n506_, new_n505_, keyIn_0_28 );
not g388 ( new_n507_, keyIn_0_28 );
not g389 ( new_n508_, new_n505_ );
nand g390 ( new_n509_, new_n508_, new_n507_ );
nand g391 ( N865, new_n509_, new_n506_ );
not g392 ( new_n511_, new_n437_ );
nand g393 ( new_n512_, new_n424_, new_n511_ );
nor g394 ( new_n513_, new_n298_, new_n179_ );
nor g395 ( new_n514_, new_n129_, N268 );
nand g396 ( new_n515_, new_n318_, new_n514_ );
not g397 ( new_n516_, new_n515_ );
nand g398 ( new_n517_, new_n294_, N55 );
nor g399 ( new_n518_, new_n291_, new_n517_ );
nand g400 ( new_n519_, new_n518_, N153 );
nand g401 ( new_n520_, N138, N152 );
nand g402 ( new_n521_, new_n519_, new_n520_ );
nor g403 ( new_n522_, new_n521_, new_n516_ );
not g404 ( new_n523_, new_n522_ );
nor g405 ( new_n524_, new_n523_, new_n513_ );
not g406 ( new_n525_, new_n524_ );
nor g407 ( new_n526_, new_n525_, N177 );
not g408 ( new_n527_, new_n526_ );
nand g409 ( new_n528_, new_n512_, new_n527_ );
nand g410 ( new_n529_, new_n525_, N177 );
nand g411 ( new_n530_, new_n528_, new_n529_ );
nor g412 ( new_n531_, new_n298_, new_n178_ );
nand g413 ( new_n532_, new_n518_, N149 );
not g414 ( new_n533_, new_n532_ );
nand g415 ( new_n534_, N17, N138 );
nand g416 ( new_n535_, new_n515_, new_n534_ );
nor g417 ( new_n536_, new_n535_, new_n533_ );
not g418 ( new_n537_, new_n536_ );
nor g419 ( new_n538_, new_n537_, new_n531_ );
not g420 ( new_n539_, new_n538_ );
nor g421 ( new_n540_, new_n539_, N171 );
nor g422 ( new_n541_, new_n298_, new_n186_ );
nand g423 ( new_n542_, new_n518_, N146 );
not g424 ( new_n543_, new_n542_ );
nand g425 ( new_n544_, N51, N138 );
nand g426 ( new_n545_, new_n515_, new_n544_ );
nor g427 ( new_n546_, new_n545_, new_n543_ );
not g428 ( new_n547_, new_n546_ );
nor g429 ( new_n548_, new_n547_, new_n541_ );
not g430 ( new_n549_, new_n548_ );
nor g431 ( new_n550_, new_n549_, N165 );
nor g432 ( new_n551_, new_n540_, new_n550_ );
nand g433 ( new_n552_, new_n530_, new_n551_ );
not g434 ( new_n553_, keyIn_0_16 );
nor g435 ( new_n554_, new_n548_, new_n233_ );
nor g436 ( new_n555_, new_n554_, new_n553_ );
nand g437 ( new_n556_, new_n554_, new_n553_ );
not g438 ( new_n557_, new_n556_ );
nor g439 ( new_n558_, new_n557_, new_n555_ );
not g440 ( new_n559_, new_n558_ );
not g441 ( new_n560_, N171 );
nor g442 ( new_n561_, new_n538_, new_n560_ );
not g443 ( new_n562_, new_n561_ );
nor g444 ( new_n563_, new_n550_, new_n562_ );
nor g445 ( new_n564_, new_n559_, new_n563_ );
nand g446 ( new_n565_, new_n552_, new_n564_ );
nor g447 ( new_n566_, new_n298_, new_n184_ );
nor g448 ( new_n567_, new_n516_, keyIn_0_8 );
nand g449 ( new_n568_, new_n516_, keyIn_0_8 );
not g450 ( new_n569_, new_n568_ );
nand g451 ( new_n570_, new_n518_, N143 );
nand g452 ( new_n571_, N8, N138 );
nand g453 ( new_n572_, new_n570_, new_n571_ );
nor g454 ( new_n573_, new_n569_, new_n572_ );
not g455 ( new_n574_, new_n573_ );
nor g456 ( new_n575_, new_n574_, new_n567_ );
not g457 ( new_n576_, new_n575_ );
nor g458 ( new_n577_, new_n576_, new_n566_ );
not g459 ( new_n578_, new_n577_ );
nor g460 ( new_n579_, new_n578_, N159 );
not g461 ( new_n580_, new_n579_ );
nand g462 ( new_n581_, new_n565_, new_n580_ );
nor g463 ( new_n582_, new_n577_, new_n231_ );
not g464 ( new_n583_, new_n582_ );
nand g465 ( N866, new_n581_, new_n583_ );
not g466 ( new_n585_, new_n528_ );
nand g467 ( new_n586_, new_n585_, new_n529_ );
not g468 ( new_n587_, new_n529_ );
nor g469 ( new_n588_, new_n587_, new_n526_ );
nor g470 ( new_n589_, new_n512_, new_n588_ );
nor g471 ( new_n590_, new_n589_, new_n329_ );
nand g472 ( new_n591_, new_n586_, new_n590_ );
nand g473 ( new_n592_, new_n588_, N228 );
nand g474 ( new_n593_, new_n587_, N237 );
nand g475 ( new_n594_, new_n592_, new_n593_ );
nor g476 ( new_n595_, new_n594_, keyIn_0_23 );
nand g477 ( new_n596_, new_n594_, keyIn_0_23 );
nor g478 ( new_n597_, new_n524_, new_n439_ );
nand g479 ( new_n598_, new_n340_, N177 );
nand g480 ( new_n599_, N101, N210 );
nand g481 ( new_n600_, new_n598_, new_n599_ );
nor g482 ( new_n601_, new_n597_, new_n600_ );
nand g483 ( new_n602_, new_n596_, new_n601_ );
nor g484 ( new_n603_, new_n602_, new_n595_ );
nand g485 ( N874, new_n591_, new_n603_ );
nor g486 ( new_n605_, new_n579_, new_n582_ );
nand g487 ( new_n606_, new_n565_, new_n605_ );
nor g488 ( new_n607_, new_n565_, new_n605_ );
nor g489 ( new_n608_, new_n607_, new_n329_ );
nand g490 ( new_n609_, new_n608_, new_n606_ );
not g491 ( new_n610_, new_n605_ );
nor g492 ( new_n611_, new_n610_, new_n432_ );
not g493 ( new_n612_, new_n611_ );
nor g494 ( new_n613_, new_n612_, keyIn_0_20 );
nand g495 ( new_n614_, new_n612_, keyIn_0_20 );
nor g496 ( new_n615_, new_n583_, new_n334_ );
nand g497 ( new_n616_, new_n578_, N246 );
nor g498 ( new_n617_, new_n339_, new_n231_ );
nand g499 ( new_n618_, N210, N268 );
not g500 ( new_n619_, new_n618_ );
nor g501 ( new_n620_, new_n617_, new_n619_ );
nand g502 ( new_n621_, new_n616_, new_n620_ );
nor g503 ( new_n622_, new_n615_, new_n621_ );
nand g504 ( new_n623_, new_n614_, new_n622_ );
nor g505 ( new_n624_, new_n623_, new_n613_ );
nand g506 ( new_n625_, new_n609_, new_n624_ );
nand g507 ( new_n626_, new_n625_, keyIn_0_31 );
not g508 ( new_n627_, keyIn_0_31 );
not g509 ( new_n628_, new_n625_ );
nand g510 ( new_n629_, new_n628_, new_n627_ );
nand g511 ( N878, new_n629_, new_n626_ );
not g512 ( new_n631_, keyIn_0_29 );
not g513 ( new_n632_, new_n540_ );
nand g514 ( new_n633_, new_n530_, new_n632_ );
nand g515 ( new_n634_, new_n633_, new_n562_ );
nor g516 ( new_n635_, new_n559_, new_n550_ );
nand g517 ( new_n636_, new_n634_, new_n635_ );
nor g518 ( new_n637_, new_n634_, new_n635_ );
nor g519 ( new_n638_, new_n637_, new_n329_ );
nand g520 ( new_n639_, new_n638_, new_n636_ );
not g521 ( new_n640_, new_n639_ );
nand g522 ( new_n641_, new_n640_, new_n631_ );
nand g523 ( new_n642_, new_n639_, keyIn_0_29 );
not g524 ( new_n643_, keyIn_0_21 );
nand g525 ( new_n644_, new_n635_, N228 );
nor g526 ( new_n645_, new_n644_, new_n643_ );
nand g527 ( new_n646_, new_n644_, new_n643_ );
nand g528 ( new_n647_, new_n559_, N237 );
nor g529 ( new_n648_, new_n548_, new_n439_ );
nand g530 ( new_n649_, new_n340_, N165 );
nand g531 ( new_n650_, N91, N210 );
nand g532 ( new_n651_, new_n649_, new_n650_ );
nor g533 ( new_n652_, new_n648_, new_n651_ );
nand g534 ( new_n653_, new_n647_, new_n652_ );
not g535 ( new_n654_, new_n653_ );
nand g536 ( new_n655_, new_n646_, new_n654_ );
nor g537 ( new_n656_, new_n655_, new_n645_ );
nand g538 ( new_n657_, new_n642_, new_n656_ );
not g539 ( new_n658_, new_n657_ );
nand g540 ( N879, new_n658_, new_n641_ );
not g541 ( new_n660_, keyIn_0_26 );
not g542 ( new_n661_, new_n530_ );
nor g543 ( new_n662_, new_n540_, new_n561_ );
not g544 ( new_n663_, new_n662_ );
nand g545 ( new_n664_, new_n661_, new_n663_ );
nand g546 ( new_n665_, new_n530_, new_n662_ );
nand g547 ( new_n666_, new_n664_, new_n665_ );
nor g548 ( new_n667_, new_n666_, new_n660_ );
not g549 ( new_n668_, new_n667_ );
nor g550 ( new_n669_, new_n530_, new_n662_ );
not g551 ( new_n670_, new_n665_ );
nor g552 ( new_n671_, new_n670_, new_n669_ );
nor g553 ( new_n672_, new_n671_, keyIn_0_26 );
nor g554 ( new_n673_, new_n672_, new_n329_ );
nand g555 ( new_n674_, new_n673_, new_n668_ );
nor g556 ( new_n675_, new_n663_, new_n432_ );
nor g557 ( new_n676_, new_n562_, new_n334_ );
nor g558 ( new_n677_, new_n538_, new_n439_ );
nor g559 ( new_n678_, new_n339_, new_n560_ );
nand g560 ( new_n679_, N96, N210 );
not g561 ( new_n680_, new_n679_ );
nor g562 ( new_n681_, new_n678_, new_n680_ );
not g563 ( new_n682_, new_n681_ );
nor g564 ( new_n683_, new_n677_, new_n682_ );
not g565 ( new_n684_, new_n683_ );
nor g566 ( new_n685_, new_n676_, new_n684_ );
not g567 ( new_n686_, new_n685_ );
nor g568 ( new_n687_, new_n686_, new_n675_ );
nand g569 ( new_n688_, new_n674_, new_n687_ );
nand g570 ( new_n689_, new_n688_, keyIn_0_30 );
not g571 ( new_n690_, keyIn_0_30 );
nand g572 ( new_n691_, new_n666_, new_n660_ );
nand g573 ( new_n692_, new_n691_, N219 );
nor g574 ( new_n693_, new_n692_, new_n667_ );
not g575 ( new_n694_, new_n687_ );
nor g576 ( new_n695_, new_n693_, new_n694_ );
nand g577 ( new_n696_, new_n695_, new_n690_ );
nand g578 ( N880, new_n689_, new_n696_ );
endmodule