module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n595_, new_n614_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n421_, new_n720_, new_n620_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n241_, new_n566_, new_n641_, new_n339_, new_n365_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n246_, new_n170_, new_n682_, new_n679_, new_n266_, new_n667_, new_n367_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n534_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n602_, new_n188_, new_n695_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n735_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n742_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n157_, new_n716_, new_n153_, new_n701_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n655_, new_n630_, new_n385_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n683_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n622_, new_n629_, new_n702_, new_n321_, new_n715_, new_n443_, new_n324_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n650_, new_n708_, new_n750_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n506_, new_n680_, new_n256_, new_n452_, new_n381_, new_n656_, new_n388_, new_n508_, new_n714_, new_n194_, new_n483_, new_n394_, new_n299_, new_n657_, new_n652_, new_n314_, new_n582_, new_n363_, new_n441_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n488_, new_n524_, new_n705_, new_n277_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n437_, new_n295_, new_n359_, new_n628_, new_n162_, new_n409_, new_n745_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n688_, new_n155_, new_n384_, new_n410_, new_n543_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n232_, new_n258_, new_n724_, new_n176_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n654_, new_n713_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n749_, new_n310_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n562_, new_n578_, new_n177_, new_n493_, new_n264_, new_n665_, new_n379_, new_n719_, new_n273_, new_n224_, new_n586_, new_n570_, new_n598_, new_n520_, new_n253_, new_n717_, new_n403_, new_n475_, new_n237_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n605_, new_n748_, new_n182_, new_n407_, new_n666_, new_n480_, new_n625_, new_n730_, new_n736_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n231_, new_n219_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n428_, new_n199_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n191_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n499_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n737_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n662_, new_n440_, new_n733_, new_n531_, new_n593_, new_n252_, new_n585_, new_n312_, new_n535_, new_n372_, new_n725_, new_n242_, new_n503_, new_n527_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n651_, new_n433_, new_n435_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n278_, new_n304_, new_n638_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n711_, new_n644_, new_n731_, new_n599_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n723_, new_n594_, new_n495_, new_n431_, new_n196_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n727_, new_n375_, new_n294_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n358_, new_n348_, new_n610_, new_n159_, new_n322_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n697_, new_n185_, new_n709_, new_n373_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n551_, new_n279_, new_n455_, new_n618_, new_n521_, new_n406_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n573_, new_n405_;

nand g000 ( new_n151_, N29, N42, N75 );
not g001 ( N388, new_n151_ );
nand g002 ( new_n153_, N29, N36, N80 );
not g003 ( N389, new_n153_ );
nand g004 ( new_n155_, N29, N36, N42 );
not g005 ( N390, new_n155_ );
nand g006 ( new_n157_, N85, N86 );
not g007 ( N391, new_n157_ );
nand g008 ( new_n159_, N1, N8, N13, N17 );
not g009 ( N418, new_n159_ );
not g010 ( new_n161_, N13 );
not g011 ( new_n162_, N17 );
nand g012 ( new_n163_, N1, N26 );
nor g013 ( new_n164_, new_n163_, new_n161_, new_n162_ );
nand g014 ( N419, new_n164_, new_n155_ );
nand g015 ( N420, N59, N75, N80 );
nand g016 ( N421, N36, N59, N80 );
nand g017 ( N422, N36, N42, N59 );
not g018 ( new_n169_, N90 );
nor g019 ( new_n170_, N87, N88 );
nor g020 ( N423, new_n170_, new_n169_ );
nand g021 ( N446, new_n164_, N390 );
not g022 ( new_n173_, keyIn_0_0 );
nand g023 ( new_n174_, N1, N26, N51 );
nand g024 ( new_n175_, new_n174_, new_n173_ );
nand g025 ( new_n176_, keyIn_0_0, N1, N26, N51 );
nand g026 ( new_n177_, new_n175_, new_n176_ );
not g027 ( N447, new_n177_ );
nand g028 ( new_n179_, N1, N8, N13, N55 );
nand g029 ( new_n180_, N29, N68 );
nor g030 ( N448, new_n179_, new_n180_ );
not g031 ( new_n182_, N74 );
nand g032 ( new_n183_, N59, N68 );
nor g033 ( N449, new_n179_, new_n182_, new_n183_ );
not g034 ( new_n185_, N89 );
nor g035 ( N450, new_n170_, new_n185_ );
not g036 ( new_n187_, N135 );
not g037 ( new_n188_, N111 );
not g038 ( new_n189_, N116 );
nand g039 ( new_n190_, new_n188_, new_n189_ );
nand g040 ( new_n191_, N111, N116 );
nand g041 ( new_n192_, new_n190_, new_n191_ );
not g042 ( new_n193_, N121 );
not g043 ( new_n194_, N126 );
nand g044 ( new_n195_, new_n193_, new_n194_ );
nand g045 ( new_n196_, N121, N126 );
nand g046 ( new_n197_, new_n195_, new_n196_ );
nand g047 ( new_n198_, new_n192_, new_n197_ );
nand g048 ( new_n199_, new_n190_, new_n195_, new_n191_, new_n196_ );
nand g049 ( new_n200_, new_n198_, new_n199_ );
nand g050 ( new_n201_, new_n200_, new_n187_ );
nand g051 ( new_n202_, new_n201_, keyIn_0_21 );
not g052 ( new_n203_, keyIn_0_21 );
nand g053 ( new_n204_, new_n200_, new_n203_, new_n187_ );
nand g054 ( new_n205_, new_n202_, new_n204_ );
nand g055 ( new_n206_, new_n198_, N135, new_n199_ );
nand g056 ( new_n207_, new_n205_, new_n206_ );
not g057 ( new_n208_, N130 );
not g058 ( new_n209_, N91 );
not g059 ( new_n210_, N96 );
nand g060 ( new_n211_, new_n209_, new_n210_ );
nand g061 ( new_n212_, N91, N96 );
nand g062 ( new_n213_, new_n211_, new_n212_ );
not g063 ( new_n214_, N101 );
not g064 ( new_n215_, N106 );
nand g065 ( new_n216_, new_n214_, new_n215_ );
nand g066 ( new_n217_, N101, N106 );
nand g067 ( new_n218_, new_n216_, new_n217_ );
nand g068 ( new_n219_, new_n213_, new_n218_ );
nand g069 ( new_n220_, new_n211_, new_n216_, new_n212_, new_n217_ );
nand g070 ( new_n221_, new_n219_, new_n220_ );
nand g071 ( new_n222_, new_n221_, new_n208_ );
nand g072 ( new_n223_, new_n219_, N130, new_n220_ );
nand g073 ( new_n224_, new_n222_, new_n223_ );
nand g074 ( new_n225_, new_n207_, new_n224_ );
nand g075 ( new_n226_, new_n205_, new_n206_, new_n222_, new_n223_ );
nand g076 ( new_n227_, new_n225_, new_n226_ );
not g077 ( N767, new_n227_ );
not g078 ( new_n229_, N207 );
nor g079 ( new_n230_, N195, N201 );
not g080 ( new_n231_, new_n230_ );
nand g081 ( new_n232_, N195, N201 );
nand g082 ( new_n233_, new_n231_, new_n232_ );
not g083 ( new_n234_, new_n233_ );
nand g084 ( new_n235_, keyIn_0_6, N183 );
nand g085 ( new_n236_, new_n234_, new_n235_ );
not g086 ( new_n237_, new_n236_ );
nor g087 ( new_n238_, new_n234_, new_n235_ );
nor g088 ( new_n239_, new_n237_, new_n238_ );
not g089 ( new_n240_, new_n239_ );
not g090 ( new_n241_, N189 );
nor g091 ( new_n242_, keyIn_0_6, N183 );
nor g092 ( new_n243_, new_n242_, new_n241_ );
nand g093 ( new_n244_, new_n240_, new_n243_ );
not g094 ( new_n245_, new_n243_ );
nand g095 ( new_n246_, new_n239_, new_n245_ );
nand g096 ( new_n247_, new_n244_, new_n246_ );
nand g097 ( new_n248_, new_n247_, new_n229_ );
nand g098 ( new_n249_, new_n244_, N207, new_n246_ );
nand g099 ( new_n250_, new_n248_, new_n249_ );
not g100 ( new_n251_, N159 );
not g101 ( new_n252_, N165 );
nand g102 ( new_n253_, new_n251_, new_n252_ );
nand g103 ( new_n254_, N159, N165 );
nand g104 ( new_n255_, new_n253_, new_n254_ );
not g105 ( new_n256_, N171 );
not g106 ( new_n257_, N177 );
nand g107 ( new_n258_, new_n256_, new_n257_ );
nand g108 ( new_n259_, N171, N177 );
nand g109 ( new_n260_, new_n258_, new_n259_ );
nand g110 ( new_n261_, new_n255_, new_n260_ );
nand g111 ( new_n262_, new_n253_, new_n258_, new_n254_, new_n259_ );
nand g112 ( new_n263_, new_n261_, new_n262_ );
nand g113 ( new_n264_, new_n263_, new_n208_ );
nand g114 ( new_n265_, new_n261_, N130, new_n262_ );
nand g115 ( new_n266_, new_n264_, new_n265_ );
nand g116 ( new_n267_, new_n250_, new_n266_ );
nand g117 ( new_n268_, new_n248_, new_n249_, new_n264_, new_n265_ );
nand g118 ( new_n269_, new_n267_, new_n268_ );
not g119 ( N768, new_n269_ );
not g120 ( new_n271_, keyIn_0_30 );
not g121 ( new_n272_, keyIn_0_18 );
not g122 ( new_n273_, keyIn_0_12 );
nand g123 ( new_n274_, new_n177_, keyIn_0_8 );
not g124 ( new_n275_, keyIn_0_8 );
nand g125 ( new_n276_, new_n175_, new_n275_, new_n176_ );
nand g126 ( new_n277_, new_n274_, new_n276_ );
nand g127 ( new_n278_, new_n277_, new_n273_ );
nand g128 ( new_n279_, new_n274_, keyIn_0_12, new_n276_ );
nand g129 ( new_n280_, new_n278_, new_n279_ );
nand g130 ( new_n281_, N59, N156 );
not g131 ( new_n282_, new_n281_ );
nand g132 ( new_n283_, new_n282_, keyIn_0_3 );
not g133 ( new_n284_, keyIn_0_3 );
nand g134 ( new_n285_, new_n281_, new_n284_ );
nand g135 ( new_n286_, new_n283_, new_n285_ );
nand g136 ( new_n287_, new_n280_, keyIn_0_16, N17, new_n286_ );
not g137 ( new_n288_, keyIn_0_16 );
nand g138 ( new_n289_, new_n280_, N17, new_n286_ );
nand g139 ( new_n290_, new_n289_, new_n288_ );
nand g140 ( new_n291_, new_n290_, N1, new_n287_ );
nand g141 ( new_n292_, new_n291_, new_n272_ );
nand g142 ( new_n293_, new_n290_, keyIn_0_18, N1, new_n287_ );
nand g143 ( new_n294_, new_n292_, new_n293_ );
not g144 ( new_n295_, new_n294_ );
nand g145 ( new_n296_, new_n295_, N153 );
not g146 ( new_n297_, keyIn_0_11 );
nor g147 ( new_n298_, N17, N42 );
nor g148 ( new_n299_, new_n298_, keyIn_0_4 );
not g149 ( new_n300_, keyIn_0_4 );
nor g150 ( new_n301_, new_n300_, N17, N42 );
nor g151 ( new_n302_, new_n299_, new_n301_ );
not g152 ( new_n303_, keyIn_0_5 );
nand g153 ( new_n304_, N17, N42 );
nand g154 ( new_n305_, new_n304_, new_n303_ );
nand g155 ( new_n306_, keyIn_0_5, N17, N42 );
nand g156 ( new_n307_, new_n305_, new_n306_ );
not g157 ( new_n308_, new_n307_ );
nand g158 ( new_n309_, new_n302_, new_n308_, new_n297_ );
not g159 ( new_n310_, N42 );
nand g160 ( new_n311_, new_n162_, new_n310_ );
nand g161 ( new_n312_, new_n311_, new_n300_ );
nand g162 ( new_n313_, new_n298_, keyIn_0_4 );
nand g163 ( new_n314_, new_n312_, new_n313_, new_n305_, new_n306_ );
nand g164 ( new_n315_, new_n314_, keyIn_0_11 );
nand g165 ( new_n316_, new_n315_, new_n309_, new_n282_ );
not g166 ( new_n317_, new_n316_ );
nand g167 ( new_n318_, new_n280_, new_n317_ );
nand g168 ( new_n319_, new_n318_, keyIn_0_15 );
not g169 ( new_n320_, keyIn_0_15 );
nand g170 ( new_n321_, new_n280_, new_n317_, new_n320_ );
nand g171 ( new_n322_, new_n319_, new_n321_ );
not g172 ( new_n323_, keyIn_0_13 );
not g173 ( new_n324_, keyIn_0_2 );
nand g174 ( new_n325_, N42, N59, N75 );
nand g175 ( new_n326_, new_n325_, new_n324_ );
nand g176 ( new_n327_, keyIn_0_2, N42, N59, N75 );
nand g177 ( new_n328_, new_n326_, new_n327_ );
nand g178 ( new_n329_, new_n328_, keyIn_0_10 );
not g179 ( new_n330_, keyIn_0_10 );
nand g180 ( new_n331_, new_n326_, new_n330_, new_n327_ );
nand g181 ( new_n332_, new_n329_, new_n331_ );
not g182 ( new_n333_, new_n332_ );
not g183 ( new_n334_, keyIn_0_1 );
nand g184 ( new_n335_, N17, N51 );
not g185 ( new_n336_, new_n335_ );
nand g186 ( new_n337_, new_n336_, N1, N8 );
nand g187 ( new_n338_, new_n337_, new_n334_ );
nand g188 ( new_n339_, new_n336_, keyIn_0_1, N1, N8 );
nand g189 ( new_n340_, new_n338_, new_n339_ );
nand g190 ( new_n341_, new_n340_, keyIn_0_9 );
not g191 ( new_n342_, keyIn_0_9 );
nand g192 ( new_n343_, new_n338_, new_n342_, new_n339_ );
nand g193 ( new_n344_, new_n333_, new_n341_, new_n343_ );
nand g194 ( new_n345_, new_n344_, new_n323_ );
nand g195 ( new_n346_, new_n333_, new_n341_, keyIn_0_13, new_n343_ );
nand g196 ( new_n347_, new_n345_, new_n346_ );
nand g197 ( new_n348_, new_n322_, new_n347_ );
nand g198 ( new_n349_, new_n348_, keyIn_0_17 );
not g199 ( new_n350_, keyIn_0_17 );
nand g200 ( new_n351_, new_n322_, new_n350_, new_n347_ );
nand g201 ( new_n352_, new_n349_, new_n351_ );
nand g202 ( new_n353_, new_n352_, N126 );
nand g203 ( new_n354_, new_n296_, new_n353_ );
nand g204 ( new_n355_, new_n354_, keyIn_0_27 );
not g205 ( new_n356_, keyIn_0_27 );
nand g206 ( new_n357_, new_n296_, new_n353_, new_n356_ );
nand g207 ( new_n358_, new_n355_, new_n357_ );
not g208 ( new_n359_, N268 );
not g209 ( new_n360_, keyIn_0_14 );
nand g210 ( new_n361_, new_n280_, N29, N75, N80 );
not g211 ( new_n362_, new_n361_ );
nand g212 ( new_n363_, new_n362_, N55 );
nand g213 ( new_n364_, new_n363_, new_n360_ );
nand g214 ( new_n365_, new_n362_, keyIn_0_14, N55 );
nand g215 ( new_n366_, new_n364_, new_n365_ );
nand g216 ( new_n367_, new_n366_, new_n359_ );
nand g217 ( new_n368_, new_n358_, new_n367_ );
nand g218 ( new_n369_, new_n368_, new_n271_ );
nand g219 ( new_n370_, new_n358_, keyIn_0_30, new_n367_ );
nand g220 ( new_n371_, new_n369_, new_n370_ );
not g221 ( new_n372_, new_n371_ );
nand g222 ( new_n373_, new_n372_, N201 );
not g223 ( new_n374_, N201 );
nand g224 ( new_n375_, new_n371_, new_n374_ );
nand g225 ( new_n376_, new_n375_, keyIn_0_35 );
not g226 ( new_n377_, keyIn_0_35 );
nand g227 ( new_n378_, new_n371_, new_n377_, new_n374_ );
nand g228 ( new_n379_, new_n376_, new_n378_ );
nand g229 ( new_n380_, new_n379_, new_n373_ );
not g230 ( new_n381_, new_n380_ );
nand g231 ( new_n382_, new_n381_, N261 );
not g232 ( new_n383_, N261 );
nand g233 ( new_n384_, new_n380_, new_n383_ );
nand g234 ( new_n385_, new_n382_, N219, new_n384_ );
nand g235 ( new_n386_, new_n381_, N228 );
not g236 ( new_n387_, new_n373_ );
nand g237 ( new_n388_, new_n387_, N237 );
nand g238 ( new_n389_, new_n372_, N246 );
nand g239 ( new_n390_, N42, N72, N73 );
nor g240 ( new_n391_, new_n179_, new_n390_, new_n183_ );
nand g241 ( new_n392_, new_n391_, N201 );
nand g242 ( new_n393_, keyIn_0_7, N121, N210 );
nand g243 ( new_n394_, N255, N267 );
not g244 ( new_n395_, keyIn_0_7 );
nand g245 ( new_n396_, N121, N210 );
nand g246 ( new_n397_, new_n396_, new_n395_ );
nand g247 ( new_n398_, new_n397_, new_n393_, new_n394_ );
not g248 ( new_n399_, new_n398_ );
nand g249 ( new_n400_, new_n388_, new_n389_, new_n392_, new_n399_ );
not g250 ( new_n401_, new_n400_ );
nand g251 ( N850, new_n385_, new_n386_, new_n401_ );
not g252 ( new_n403_, keyIn_0_32 );
not g253 ( new_n404_, keyIn_0_25 );
nand g254 ( new_n405_, new_n292_, N146, new_n293_ );
nand g255 ( new_n406_, new_n405_, keyIn_0_22 );
not g256 ( new_n407_, keyIn_0_22 );
nand g257 ( new_n408_, new_n292_, new_n407_, N146, new_n293_ );
nand g258 ( new_n409_, new_n406_, new_n408_ );
not g259 ( new_n410_, keyIn_0_23 );
nand g260 ( new_n411_, new_n352_, N116 );
nand g261 ( new_n412_, new_n411_, new_n410_ );
nand g262 ( new_n413_, new_n352_, keyIn_0_23, N116 );
nand g263 ( new_n414_, new_n412_, new_n409_, new_n413_ );
nand g264 ( new_n415_, new_n414_, new_n404_ );
nand g265 ( new_n416_, new_n412_, keyIn_0_25, new_n409_, new_n413_ );
nand g266 ( new_n417_, new_n415_, new_n416_ );
not g267 ( new_n418_, new_n367_ );
nand g268 ( new_n419_, new_n418_, keyIn_0_20 );
not g269 ( new_n420_, keyIn_0_20 );
nand g270 ( new_n421_, new_n367_, new_n420_ );
nand g271 ( new_n422_, new_n419_, new_n421_ );
nand g272 ( new_n423_, new_n417_, new_n422_ );
nand g273 ( new_n424_, new_n423_, keyIn_0_28 );
not g274 ( new_n425_, keyIn_0_28 );
nand g275 ( new_n426_, new_n417_, new_n425_, new_n422_ );
nand g276 ( new_n427_, new_n424_, new_n426_ );
nand g277 ( new_n428_, new_n427_, new_n241_ );
nand g278 ( new_n429_, new_n428_, new_n403_ );
nand g279 ( new_n430_, new_n427_, keyIn_0_32, new_n241_ );
nand g280 ( new_n431_, new_n429_, new_n430_ );
not g281 ( new_n432_, keyIn_0_34 );
not g282 ( new_n433_, N195 );
not g283 ( new_n434_, keyIn_0_29 );
not g284 ( new_n435_, keyIn_0_26 );
nand g285 ( new_n436_, new_n352_, keyIn_0_24, N121 );
nand g286 ( new_n437_, new_n295_, N149 );
not g287 ( new_n438_, keyIn_0_24 );
nand g288 ( new_n439_, new_n352_, N121 );
nand g289 ( new_n440_, new_n439_, new_n438_ );
nand g290 ( new_n441_, new_n440_, new_n435_, new_n436_, new_n437_ );
nand g291 ( new_n442_, new_n440_, new_n436_, new_n437_ );
nand g292 ( new_n443_, new_n442_, keyIn_0_26 );
nand g293 ( new_n444_, new_n443_, new_n367_, new_n441_ );
nand g294 ( new_n445_, new_n444_, new_n434_ );
nand g295 ( new_n446_, new_n443_, keyIn_0_29, new_n367_, new_n441_ );
nand g296 ( new_n447_, new_n445_, new_n446_ );
nand g297 ( new_n448_, new_n447_, new_n433_ );
nand g298 ( new_n449_, new_n448_, new_n432_ );
nand g299 ( new_n450_, new_n447_, keyIn_0_34, new_n433_ );
nand g300 ( new_n451_, new_n449_, new_n450_ );
nand g301 ( new_n452_, new_n431_, new_n387_, new_n451_ );
nand g302 ( new_n453_, new_n452_, keyIn_0_41 );
not g303 ( new_n454_, keyIn_0_41 );
nand g304 ( new_n455_, new_n431_, new_n454_, new_n387_, new_n451_ );
nand g305 ( new_n456_, new_n453_, new_n455_ );
nand g306 ( new_n457_, new_n431_, N261, new_n379_, new_n451_ );
nand g307 ( new_n458_, new_n457_, keyIn_0_38 );
not g308 ( new_n459_, keyIn_0_38 );
nand g309 ( new_n460_, new_n379_, N261 );
not g310 ( new_n461_, new_n460_ );
nand g311 ( new_n462_, new_n461_, new_n459_, new_n431_, new_n451_ );
nand g312 ( new_n463_, new_n458_, new_n462_ );
not g313 ( new_n464_, new_n463_ );
not g314 ( new_n465_, keyIn_0_36 );
nand g315 ( new_n466_, new_n424_, N189, new_n426_ );
nand g316 ( new_n467_, new_n466_, keyIn_0_31 );
not g317 ( new_n468_, keyIn_0_31 );
nand g318 ( new_n469_, new_n424_, new_n468_, N189, new_n426_ );
nand g319 ( new_n470_, new_n467_, new_n469_ );
nand g320 ( new_n471_, new_n470_, new_n465_ );
nand g321 ( new_n472_, new_n467_, keyIn_0_36, new_n469_ );
nand g322 ( new_n473_, new_n471_, new_n472_ );
nand g323 ( new_n474_, new_n473_, keyIn_0_39 );
not g324 ( new_n475_, keyIn_0_39 );
nand g325 ( new_n476_, new_n471_, new_n475_, new_n472_ );
nand g326 ( new_n477_, new_n474_, new_n476_ );
not g327 ( new_n478_, keyIn_0_40 );
not g328 ( new_n479_, keyIn_0_33 );
nand g329 ( new_n480_, new_n445_, N195, new_n446_ );
nand g330 ( new_n481_, new_n480_, new_n479_ );
nand g331 ( new_n482_, new_n445_, keyIn_0_33, N195, new_n446_ );
nand g332 ( new_n483_, new_n481_, new_n482_ );
nand g333 ( new_n484_, new_n483_, keyIn_0_37 );
not g334 ( new_n485_, keyIn_0_37 );
nand g335 ( new_n486_, new_n481_, new_n485_, new_n482_ );
nand g336 ( new_n487_, new_n431_, new_n484_, new_n486_ );
nand g337 ( new_n488_, new_n487_, new_n478_ );
nand g338 ( new_n489_, new_n431_, keyIn_0_40, new_n484_, new_n486_ );
nand g339 ( new_n490_, new_n488_, new_n489_ );
not g340 ( new_n491_, new_n490_ );
nand g341 ( new_n492_, new_n464_, new_n491_, new_n456_, new_n477_ );
nand g342 ( new_n493_, new_n492_, keyIn_0_42 );
not g343 ( new_n494_, keyIn_0_42 );
not g344 ( new_n495_, new_n456_ );
nor g345 ( new_n496_, new_n495_, new_n463_ );
not g346 ( new_n497_, new_n477_ );
nor g347 ( new_n498_, new_n497_, new_n490_ );
nand g348 ( new_n499_, new_n496_, new_n498_, new_n494_ );
nand g349 ( new_n500_, new_n493_, new_n499_ );
nand g350 ( new_n501_, new_n295_, N143 );
nand g351 ( new_n502_, new_n352_, N111 );
nand g352 ( new_n503_, new_n418_, keyIn_0_19 );
not g353 ( new_n504_, keyIn_0_19 );
nand g354 ( new_n505_, new_n367_, new_n504_ );
nand g355 ( new_n506_, new_n503_, new_n505_ );
nand g356 ( new_n507_, new_n506_, new_n501_, new_n502_ );
nand g357 ( new_n508_, new_n507_, N183 );
not g358 ( new_n509_, N183 );
nand g359 ( new_n510_, new_n506_, new_n509_, new_n501_, new_n502_ );
nand g360 ( new_n511_, new_n508_, new_n510_ );
not g361 ( new_n512_, new_n511_ );
nand g362 ( new_n513_, new_n500_, new_n512_ );
nand g363 ( new_n514_, new_n493_, new_n499_, new_n511_ );
nand g364 ( new_n515_, new_n513_, N219, new_n514_ );
nand g365 ( new_n516_, new_n512_, N228 );
nand g366 ( new_n517_, new_n507_, N183, N237 );
nand g367 ( new_n518_, new_n507_, N246 );
nand g368 ( new_n519_, new_n391_, N183 );
nand g369 ( new_n520_, N106, N210 );
nand g370 ( new_n521_, new_n517_, new_n518_, new_n519_, new_n520_ );
not g371 ( new_n522_, new_n521_ );
nand g372 ( N863, new_n515_, new_n516_, new_n522_ );
not g373 ( new_n524_, keyIn_0_50 );
not g374 ( new_n525_, new_n470_ );
nand g375 ( new_n526_, new_n525_, new_n431_ );
not g376 ( new_n527_, new_n526_ );
nand g377 ( new_n528_, new_n484_, new_n486_ );
nand g378 ( new_n529_, new_n460_, new_n373_ );
nand g379 ( new_n530_, new_n529_, new_n451_ );
nand g380 ( new_n531_, new_n530_, new_n528_ );
nand g381 ( new_n532_, new_n531_, new_n527_ );
nand g382 ( new_n533_, new_n530_, new_n528_, new_n526_ );
nand g383 ( new_n534_, new_n532_, N219, new_n533_ );
nand g384 ( new_n535_, N111, N210 );
nand g385 ( new_n536_, new_n534_, new_n535_ );
nand g386 ( new_n537_, new_n536_, new_n524_ );
nand g387 ( new_n538_, new_n534_, keyIn_0_50, new_n535_ );
nand g388 ( new_n539_, new_n537_, new_n538_ );
nand g389 ( new_n540_, new_n471_, N237, new_n472_ );
nand g390 ( new_n541_, new_n527_, N228 );
nand g391 ( new_n542_, new_n424_, N246, new_n426_ );
nand g392 ( new_n543_, new_n391_, N189 );
nand g393 ( new_n544_, N255, N259 );
nand g394 ( new_n545_, new_n542_, new_n543_, new_n544_ );
not g395 ( new_n546_, new_n545_ );
nand g396 ( N864, new_n539_, new_n540_, new_n541_, new_n546_ );
nand g397 ( new_n548_, new_n451_, new_n483_ );
nand g398 ( new_n549_, new_n548_, new_n373_, new_n460_ );
not g399 ( new_n550_, new_n548_ );
nand g400 ( new_n551_, new_n550_, new_n529_ );
nand g401 ( new_n552_, new_n551_, N219, new_n549_ );
nand g402 ( new_n553_, new_n484_, N237, new_n486_ );
nand g403 ( new_n554_, new_n550_, N228 );
nand g404 ( new_n555_, new_n445_, N246, new_n446_ );
nand g405 ( new_n556_, new_n391_, N195 );
nand g406 ( new_n557_, N116, N210 );
nand g407 ( new_n558_, N255, N260 );
nand g408 ( new_n559_, new_n555_, new_n556_, new_n557_, new_n558_ );
not g409 ( new_n560_, new_n559_ );
nand g410 ( N865, new_n552_, new_n553_, new_n554_, new_n560_ );
not g411 ( new_n562_, keyIn_0_48 );
not g412 ( new_n563_, keyIn_0_47 );
not g413 ( new_n564_, keyIn_0_44 );
nand g414 ( new_n565_, new_n500_, new_n510_ );
nand g415 ( new_n566_, new_n565_, keyIn_0_43 );
not g416 ( new_n567_, keyIn_0_43 );
nand g417 ( new_n568_, new_n500_, new_n567_, new_n510_ );
nand g418 ( new_n569_, new_n566_, new_n568_ );
nand g419 ( new_n570_, new_n569_, new_n508_ );
nand g420 ( new_n571_, new_n570_, new_n564_ );
nand g421 ( new_n572_, new_n569_, keyIn_0_44, new_n508_ );
nand g422 ( new_n573_, new_n352_, N96 );
nand g423 ( new_n574_, new_n280_, N55, new_n286_ );
not g424 ( new_n575_, new_n574_ );
nand g425 ( new_n576_, new_n575_, N146 );
nand g426 ( new_n577_, N51, N138 );
nand g427 ( new_n578_, new_n362_, N17, new_n359_ );
nand g428 ( new_n579_, new_n578_, new_n576_, new_n577_ );
not g429 ( new_n580_, new_n579_ );
nand g430 ( new_n581_, new_n573_, new_n252_, new_n580_ );
nand g431 ( new_n582_, new_n352_, N101 );
nand g432 ( new_n583_, new_n575_, N149 );
nand g433 ( new_n584_, N17, N138 );
nand g434 ( new_n585_, new_n578_, new_n583_, new_n584_ );
not g435 ( new_n586_, new_n585_ );
nand g436 ( new_n587_, new_n582_, new_n256_, new_n586_ );
nand g437 ( new_n588_, new_n581_, new_n587_ );
not g438 ( new_n589_, new_n588_ );
nand g439 ( new_n590_, new_n352_, N106 );
nand g440 ( new_n591_, new_n575_, N153 );
nand g441 ( new_n592_, N138, N152 );
nand g442 ( new_n593_, new_n578_, new_n591_, new_n592_ );
not g443 ( new_n594_, new_n593_ );
nand g444 ( new_n595_, new_n590_, new_n257_, new_n594_ );
nand g445 ( new_n596_, new_n589_, new_n595_ );
not g446 ( new_n597_, new_n596_ );
nand g447 ( new_n598_, new_n571_, new_n563_, new_n572_, new_n597_ );
nand g448 ( new_n599_, new_n571_, new_n572_, new_n597_ );
nand g449 ( new_n600_, new_n599_, keyIn_0_47 );
nand g450 ( new_n601_, new_n590_, new_n594_ );
nand g451 ( new_n602_, new_n601_, N177 );
nand g452 ( new_n603_, new_n582_, new_n586_ );
nand g453 ( new_n604_, new_n603_, N171 );
nand g454 ( new_n605_, new_n602_, new_n604_ );
nand g455 ( new_n606_, new_n589_, new_n605_ );
nand g456 ( new_n607_, new_n573_, new_n580_ );
nand g457 ( new_n608_, new_n607_, N165 );
nand g458 ( new_n609_, new_n606_, new_n608_ );
not g459 ( new_n610_, new_n609_ );
nand g460 ( new_n611_, new_n600_, new_n598_, new_n610_ );
nand g461 ( new_n612_, new_n611_, new_n562_ );
nand g462 ( new_n613_, new_n600_, keyIn_0_48, new_n598_, new_n610_ );
nand g463 ( new_n614_, new_n612_, new_n613_ );
nand g464 ( new_n615_, new_n352_, N91 );
nand g465 ( new_n616_, new_n575_, N143 );
nand g466 ( new_n617_, N8, N138 );
nand g467 ( new_n618_, new_n578_, new_n616_, new_n617_ );
not g468 ( new_n619_, new_n618_ );
nand g469 ( new_n620_, new_n615_, new_n251_, new_n619_ );
nand g470 ( new_n621_, new_n614_, new_n620_ );
nand g471 ( new_n622_, new_n615_, new_n619_ );
nand g472 ( new_n623_, new_n622_, N159 );
nand g473 ( N866, new_n621_, new_n623_ );
not g474 ( new_n625_, keyIn_0_61 );
nand g475 ( new_n626_, new_n571_, new_n572_ );
not g476 ( new_n627_, new_n626_ );
nand g477 ( new_n628_, new_n602_, new_n595_ );
not g478 ( new_n629_, new_n628_ );
nand g479 ( new_n630_, new_n627_, new_n629_ );
nand g480 ( new_n631_, new_n630_, keyIn_0_46 );
nand g481 ( new_n632_, new_n626_, new_n628_ );
nand g482 ( new_n633_, new_n632_, keyIn_0_45 );
nand g483 ( new_n634_, new_n631_, new_n633_ );
not g484 ( new_n635_, new_n634_ );
not g485 ( new_n636_, keyIn_0_45 );
nand g486 ( new_n637_, new_n626_, new_n636_, new_n628_ );
not g487 ( new_n638_, keyIn_0_46 );
nand g488 ( new_n639_, new_n627_, new_n638_, new_n629_ );
nand g489 ( new_n640_, new_n635_, keyIn_0_49, new_n637_, new_n639_ );
not g490 ( new_n641_, keyIn_0_49 );
nand g491 ( new_n642_, new_n635_, new_n637_, new_n639_ );
nand g492 ( new_n643_, new_n642_, new_n641_ );
nand g493 ( new_n644_, new_n643_, N219, new_n640_ );
nand g494 ( new_n645_, new_n644_, keyIn_0_53 );
not g495 ( new_n646_, keyIn_0_53 );
nand g496 ( new_n647_, new_n643_, new_n646_, N219, new_n640_ );
nand g497 ( new_n648_, new_n645_, new_n647_ );
nand g498 ( new_n649_, N101, N210 );
nand g499 ( new_n650_, new_n648_, new_n649_ );
nand g500 ( new_n651_, new_n650_, keyIn_0_55 );
not g501 ( new_n652_, keyIn_0_55 );
nand g502 ( new_n653_, new_n648_, new_n652_, new_n649_ );
nand g503 ( new_n654_, new_n651_, new_n653_ );
nand g504 ( new_n655_, new_n629_, N228 );
not g505 ( new_n656_, new_n655_ );
nand g506 ( new_n657_, new_n601_, N177, N237 );
nand g507 ( new_n658_, new_n601_, N246 );
nand g508 ( new_n659_, new_n391_, N177 );
nand g509 ( new_n660_, new_n657_, new_n658_, new_n659_ );
nor g510 ( new_n661_, new_n656_, new_n660_ );
nand g511 ( new_n662_, new_n654_, new_n661_ );
nand g512 ( new_n663_, new_n662_, keyIn_0_57 );
not g513 ( new_n664_, keyIn_0_57 );
nand g514 ( new_n665_, new_n654_, new_n664_, new_n661_ );
nand g515 ( new_n666_, new_n663_, new_n665_ );
nand g516 ( new_n667_, new_n666_, keyIn_0_59 );
not g517 ( new_n668_, keyIn_0_59 );
nand g518 ( new_n669_, new_n663_, new_n668_, new_n665_ );
nand g519 ( new_n670_, new_n667_, new_n669_ );
nand g520 ( new_n671_, new_n670_, new_n625_ );
nand g521 ( new_n672_, new_n667_, keyIn_0_61, new_n669_ );
nand g522 ( new_n673_, new_n671_, new_n672_ );
not g523 ( N874, new_n673_ );
not g524 ( new_n675_, keyIn_0_62 );
not g525 ( new_n676_, keyIn_0_58 );
not g526 ( new_n677_, keyIn_0_54 );
not g527 ( new_n678_, keyIn_0_52 );
nand g528 ( new_n679_, new_n623_, new_n620_ );
not g529 ( new_n680_, new_n679_ );
nand g530 ( new_n681_, new_n614_, new_n678_, new_n680_ );
not g531 ( new_n682_, keyIn_0_51 );
nand g532 ( new_n683_, new_n612_, new_n682_, new_n613_, new_n679_ );
nand g533 ( new_n684_, new_n612_, new_n613_, new_n679_ );
nand g534 ( new_n685_, new_n684_, keyIn_0_51 );
nand g535 ( new_n686_, new_n614_, new_n680_ );
nand g536 ( new_n687_, new_n686_, keyIn_0_52 );
nand g537 ( new_n688_, new_n687_, new_n681_, new_n683_, new_n685_ );
nand g538 ( new_n689_, new_n688_, new_n677_ );
nand g539 ( new_n690_, new_n681_, new_n683_ );
not g540 ( new_n691_, new_n690_ );
nand g541 ( new_n692_, new_n691_, keyIn_0_54, new_n685_, new_n687_ );
nand g542 ( new_n693_, new_n692_, new_n689_ );
nand g543 ( new_n694_, new_n693_, N219 );
nand g544 ( new_n695_, new_n694_, keyIn_0_56 );
not g545 ( new_n696_, keyIn_0_56 );
nand g546 ( new_n697_, new_n693_, new_n696_, N219 );
nand g547 ( new_n698_, new_n695_, new_n697_ );
nand g548 ( new_n699_, N210, N268 );
nand g549 ( new_n700_, new_n698_, new_n676_, new_n699_ );
nand g550 ( new_n701_, new_n698_, new_n699_ );
nand g551 ( new_n702_, new_n701_, keyIn_0_58 );
nand g552 ( new_n703_, new_n680_, N228 );
not g553 ( new_n704_, new_n703_ );
nand g554 ( new_n705_, new_n622_, N159, N237 );
nand g555 ( new_n706_, new_n622_, N246 );
nand g556 ( new_n707_, new_n391_, N159 );
nand g557 ( new_n708_, new_n705_, new_n706_, new_n707_ );
nor g558 ( new_n709_, new_n704_, new_n708_ );
nand g559 ( new_n710_, new_n702_, new_n700_, new_n709_ );
nand g560 ( new_n711_, new_n710_, keyIn_0_60 );
not g561 ( new_n712_, keyIn_0_60 );
nand g562 ( new_n713_, new_n702_, new_n712_, new_n700_, new_n709_ );
nand g563 ( new_n714_, new_n711_, new_n713_ );
nand g564 ( new_n715_, new_n714_, new_n675_ );
nand g565 ( new_n716_, new_n711_, keyIn_0_62, new_n713_ );
nand g566 ( new_n717_, new_n715_, new_n716_ );
nand g567 ( new_n718_, new_n717_, keyIn_0_63 );
not g568 ( new_n719_, keyIn_0_63 );
nand g569 ( new_n720_, new_n715_, new_n719_, new_n716_ );
nand g570 ( N878, new_n718_, new_n720_ );
nand g571 ( new_n722_, new_n627_, new_n595_ );
nand g572 ( new_n723_, new_n722_, new_n602_ );
nand g573 ( new_n724_, new_n723_, new_n587_ );
nand g574 ( new_n725_, new_n724_, new_n604_ );
nand g575 ( new_n726_, new_n608_, new_n581_ );
not g576 ( new_n727_, new_n726_ );
nand g577 ( new_n728_, new_n725_, new_n727_ );
nand g578 ( new_n729_, new_n724_, new_n604_, new_n726_ );
nand g579 ( new_n730_, new_n728_, N219, new_n729_ );
nand g580 ( new_n731_, new_n727_, N228 );
nand g581 ( new_n732_, new_n607_, N165, N237 );
nand g582 ( new_n733_, new_n607_, N246 );
nand g583 ( new_n734_, new_n391_, N165 );
nand g584 ( new_n735_, N91, N210 );
nand g585 ( new_n736_, new_n732_, new_n733_, new_n734_, new_n735_ );
not g586 ( new_n737_, new_n736_ );
nand g587 ( N879, new_n730_, new_n731_, new_n737_ );
nand g588 ( new_n739_, new_n604_, new_n587_ );
not g589 ( new_n740_, new_n739_ );
nand g590 ( new_n741_, new_n723_, new_n740_ );
nand g591 ( new_n742_, new_n722_, new_n602_, new_n739_ );
nand g592 ( new_n743_, new_n741_, N219, new_n742_ );
nand g593 ( new_n744_, new_n740_, N228 );
nand g594 ( new_n745_, new_n603_, N171, N237 );
nand g595 ( new_n746_, new_n603_, N246 );
nand g596 ( new_n747_, new_n391_, N171 );
nand g597 ( new_n748_, N96, N210 );
nand g598 ( new_n749_, new_n745_, new_n746_, new_n747_, new_n748_ );
not g599 ( new_n750_, new_n749_ );
nand g600 ( N880, new_n743_, new_n744_, new_n750_ );
endmodule