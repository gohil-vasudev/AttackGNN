module locked_c1908 (  G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,  G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n123_, new_n124_, new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_, new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_, new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n377_, new_n378_, new_n379_, new_n380_, new_n382_, new_n383_, new_n384_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n425_, new_n426_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n438_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n484_, new_n485_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_;
  INV_X1 g000 ( .A(G101), .ZN(new_n123_) );
  INV_X1 g001 ( .A(KEYINPUT22), .ZN(new_n124_) );
  INV_X1 g002 ( .A(KEYINPUT19), .ZN(new_n125_) );
  INV_X1 g003 ( .A(G116), .ZN(new_n126_) );
  NAND2_X1 g004 ( .A1(new_n126_), .A2(G113), .ZN(new_n127_) );
  INV_X1 g005 ( .A(G113), .ZN(new_n128_) );
  NAND2_X1 g006 ( .A1(new_n128_), .A2(G116), .ZN(new_n129_) );
  NAND2_X1 g007 ( .A1(new_n127_), .A2(new_n129_), .ZN(new_n130_) );
  XNOR2_X1 g008 ( .A(G119), .B(KEYINPUT3), .ZN(new_n131_) );
  NAND2_X1 g009 ( .A1(new_n130_), .A2(new_n131_), .ZN(new_n132_) );
  XNOR2_X1 g010 ( .A(G113), .B(G116), .ZN(new_n133_) );
  XOR2_X1 g011 ( .A(G119), .B(KEYINPUT3), .Z(new_n134_) );
  NAND2_X1 g012 ( .A1(new_n134_), .A2(new_n133_), .ZN(new_n135_) );
  NAND2_X1 g013 ( .A1(new_n135_), .A2(new_n132_), .ZN(new_n136_) );
  XNOR2_X1 g014 ( .A(G122), .B(KEYINPUT16), .ZN(new_n137_) );
  NAND2_X1 g015 ( .A1(new_n136_), .A2(new_n137_), .ZN(new_n138_) );
  XNOR2_X1 g016 ( .A(new_n133_), .B(new_n131_), .ZN(new_n139_) );
  INV_X1 g017 ( .A(new_n137_), .ZN(new_n140_) );
  NAND2_X1 g018 ( .A1(new_n139_), .A2(new_n140_), .ZN(new_n141_) );
  NAND2_X1 g019 ( .A1(new_n141_), .A2(new_n138_), .ZN(new_n142_) );
  INV_X1 g020 ( .A(KEYINPUT18), .ZN(new_n143_) );
  NAND2_X1 g021 ( .A1(new_n143_), .A2(KEYINPUT17), .ZN(new_n144_) );
  INV_X1 g022 ( .A(KEYINPUT17), .ZN(new_n145_) );
  NAND2_X1 g023 ( .A1(new_n145_), .A2(KEYINPUT18), .ZN(new_n146_) );
  NAND2_X1 g024 ( .A1(new_n144_), .A2(new_n146_), .ZN(new_n147_) );
  INV_X1 g025 ( .A(G953), .ZN(new_n148_) );
  NAND2_X1 g026 ( .A1(new_n148_), .A2(G224), .ZN(new_n149_) );
  NAND2_X1 g027 ( .A1(new_n147_), .A2(new_n149_), .ZN(new_n150_) );
  XNOR2_X1 g028 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(new_n151_) );
  INV_X1 g029 ( .A(new_n149_), .ZN(new_n152_) );
  NAND2_X1 g030 ( .A1(new_n151_), .A2(new_n152_), .ZN(new_n153_) );
  NAND2_X1 g031 ( .A1(new_n150_), .A2(new_n153_), .ZN(new_n154_) );
  XOR2_X1 g032 ( .A(G125), .B(G146), .Z(new_n155_) );
  INV_X1 g033 ( .A(new_n155_), .ZN(new_n156_) );
  XNOR2_X1 g034 ( .A(new_n154_), .B(new_n156_), .ZN(new_n157_) );
  XNOR2_X1 g035 ( .A(new_n142_), .B(new_n157_), .ZN(new_n158_) );
  INV_X1 g036 ( .A(KEYINPUT4), .ZN(new_n159_) );
  INV_X1 g037 ( .A(G128), .ZN(new_n160_) );
  NAND2_X1 g038 ( .A1(new_n160_), .A2(G143), .ZN(new_n161_) );
  INV_X1 g039 ( .A(G143), .ZN(new_n162_) );
  NAND2_X1 g040 ( .A1(new_n162_), .A2(G128), .ZN(new_n163_) );
  NAND2_X1 g041 ( .A1(new_n161_), .A2(new_n163_), .ZN(new_n164_) );
  NAND2_X1 g042 ( .A1(new_n164_), .A2(new_n159_), .ZN(new_n165_) );
  XNOR2_X1 g043 ( .A(G128), .B(G143), .ZN(new_n166_) );
  NAND2_X1 g044 ( .A1(new_n166_), .A2(KEYINPUT4), .ZN(new_n167_) );
  NAND2_X1 g045 ( .A1(new_n165_), .A2(new_n167_), .ZN(new_n168_) );
  XNOR2_X1 g046 ( .A(new_n168_), .B(new_n123_), .ZN(new_n169_) );
  INV_X1 g047 ( .A(G107), .ZN(new_n170_) );
  XNOR2_X1 g048 ( .A(G104), .B(G110), .ZN(new_n171_) );
  XNOR2_X1 g049 ( .A(new_n171_), .B(new_n170_), .ZN(new_n172_) );
  INV_X1 g050 ( .A(new_n172_), .ZN(new_n173_) );
  XNOR2_X1 g051 ( .A(new_n169_), .B(new_n173_), .ZN(new_n174_) );
  NAND2_X1 g052 ( .A1(new_n158_), .A2(new_n174_), .ZN(new_n175_) );
  XNOR2_X1 g053 ( .A(new_n154_), .B(new_n155_), .ZN(new_n176_) );
  NAND2_X1 g054 ( .A1(new_n142_), .A2(new_n176_), .ZN(new_n177_) );
  XNOR2_X1 g055 ( .A(new_n136_), .B(new_n140_), .ZN(new_n178_) );
  NAND2_X1 g056 ( .A1(new_n178_), .A2(new_n157_), .ZN(new_n179_) );
  NAND2_X1 g057 ( .A1(new_n179_), .A2(new_n177_), .ZN(new_n180_) );
  NAND2_X1 g058 ( .A1(new_n169_), .A2(new_n172_), .ZN(new_n181_) );
  XNOR2_X1 g059 ( .A(new_n168_), .B(G101), .ZN(new_n182_) );
  NAND2_X1 g060 ( .A1(new_n182_), .A2(new_n173_), .ZN(new_n183_) );
  NAND2_X1 g061 ( .A1(new_n181_), .A2(new_n183_), .ZN(new_n184_) );
  NAND2_X1 g062 ( .A1(new_n180_), .A2(new_n184_), .ZN(new_n185_) );
  NAND2_X1 g063 ( .A1(new_n175_), .A2(new_n185_), .ZN(new_n186_) );
  XOR2_X1 g064 ( .A(G902), .B(KEYINPUT15), .Z(new_n187_) );
  INV_X1 g065 ( .A(new_n187_), .ZN(new_n188_) );
  NAND2_X1 g066 ( .A1(new_n186_), .A2(new_n188_), .ZN(new_n189_) );
  INV_X1 g067 ( .A(G210), .ZN(new_n190_) );
  NOR2_X1 g068 ( .A1(G237), .A2(G902), .ZN(new_n191_) );
  NOR2_X1 g069 ( .A1(new_n191_), .A2(new_n190_), .ZN(new_n192_) );
  XNOR2_X1 g070 ( .A(new_n189_), .B(new_n192_), .ZN(new_n193_) );
  INV_X1 g071 ( .A(G214), .ZN(new_n194_) );
  NOR2_X1 g072 ( .A1(new_n191_), .A2(new_n194_), .ZN(new_n195_) );
  INV_X1 g073 ( .A(new_n195_), .ZN(new_n196_) );
  NAND2_X1 g074 ( .A1(new_n193_), .A2(new_n196_), .ZN(new_n197_) );
  NAND2_X1 g075 ( .A1(new_n197_), .A2(new_n125_), .ZN(new_n198_) );
  INV_X1 g076 ( .A(new_n192_), .ZN(new_n199_) );
  XNOR2_X1 g077 ( .A(new_n189_), .B(new_n199_), .ZN(new_n200_) );
  NOR2_X1 g078 ( .A1(new_n200_), .A2(new_n195_), .ZN(new_n201_) );
  NAND2_X1 g079 ( .A1(new_n201_), .A2(KEYINPUT19), .ZN(new_n202_) );
  NAND2_X1 g080 ( .A1(new_n202_), .A2(new_n198_), .ZN(new_n203_) );
  INV_X1 g081 ( .A(G952), .ZN(new_n204_) );
  NAND2_X1 g082 ( .A1(G234), .A2(G237), .ZN(new_n205_) );
  XOR2_X1 g083 ( .A(new_n205_), .B(KEYINPUT14), .Z(new_n206_) );
  NOR2_X1 g084 ( .A1(new_n206_), .A2(new_n204_), .ZN(new_n207_) );
  INV_X1 g085 ( .A(new_n207_), .ZN(new_n208_) );
  NOR2_X1 g086 ( .A1(new_n208_), .A2(G953), .ZN(new_n209_) );
  INV_X1 g087 ( .A(G902), .ZN(new_n210_) );
  NOR2_X1 g088 ( .A1(new_n206_), .A2(new_n210_), .ZN(new_n211_) );
  INV_X1 g089 ( .A(new_n211_), .ZN(new_n212_) );
  NOR2_X1 g090 ( .A1(new_n148_), .A2(G898), .ZN(new_n213_) );
  INV_X1 g091 ( .A(new_n213_), .ZN(new_n214_) );
  NOR2_X1 g092 ( .A1(new_n212_), .A2(new_n214_), .ZN(new_n215_) );
  NOR2_X1 g093 ( .A1(new_n209_), .A2(new_n215_), .ZN(new_n216_) );
  NOR2_X1 g094 ( .A1(new_n203_), .A2(new_n216_), .ZN(new_n217_) );
  NAND2_X1 g095 ( .A1(new_n217_), .A2(KEYINPUT0), .ZN(new_n218_) );
  INV_X1 g096 ( .A(KEYINPUT0), .ZN(new_n219_) );
  XNOR2_X1 g097 ( .A(new_n197_), .B(KEYINPUT19), .ZN(new_n220_) );
  INV_X1 g098 ( .A(new_n216_), .ZN(new_n221_) );
  NAND2_X1 g099 ( .A1(new_n220_), .A2(new_n221_), .ZN(new_n222_) );
  NAND2_X1 g100 ( .A1(new_n222_), .A2(new_n219_), .ZN(new_n223_) );
  NAND2_X1 g101 ( .A1(new_n223_), .A2(new_n218_), .ZN(new_n224_) );
  INV_X1 g102 ( .A(G234), .ZN(new_n225_) );
  NOR2_X1 g103 ( .A1(new_n225_), .A2(G953), .ZN(new_n226_) );
  NAND2_X1 g104 ( .A1(new_n226_), .A2(KEYINPUT8), .ZN(new_n227_) );
  INV_X1 g105 ( .A(KEYINPUT8), .ZN(new_n228_) );
  NAND2_X1 g106 ( .A1(new_n148_), .A2(G234), .ZN(new_n229_) );
  NAND2_X1 g107 ( .A1(new_n229_), .A2(new_n228_), .ZN(new_n230_) );
  NAND2_X1 g108 ( .A1(new_n227_), .A2(new_n230_), .ZN(new_n231_) );
  NAND2_X1 g109 ( .A1(new_n231_), .A2(G217), .ZN(new_n232_) );
  XOR2_X1 g110 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(new_n233_) );
  XNOR2_X1 g111 ( .A(new_n232_), .B(new_n233_), .ZN(new_n234_) );
  NAND2_X1 g112 ( .A1(new_n234_), .A2(new_n126_), .ZN(new_n235_) );
  INV_X1 g113 ( .A(new_n233_), .ZN(new_n236_) );
  XNOR2_X1 g114 ( .A(new_n232_), .B(new_n236_), .ZN(new_n237_) );
  NAND2_X1 g115 ( .A1(new_n237_), .A2(G116), .ZN(new_n238_) );
  NAND2_X1 g116 ( .A1(new_n235_), .A2(new_n238_), .ZN(new_n239_) );
  XNOR2_X1 g117 ( .A(new_n166_), .B(new_n170_), .ZN(new_n240_) );
  INV_X1 g118 ( .A(new_n240_), .ZN(new_n241_) );
  XNOR2_X1 g119 ( .A(new_n239_), .B(new_n241_), .ZN(new_n242_) );
  XOR2_X1 g120 ( .A(G122), .B(G134), .Z(new_n243_) );
  INV_X1 g121 ( .A(new_n243_), .ZN(new_n244_) );
  NAND2_X1 g122 ( .A1(new_n242_), .A2(new_n244_), .ZN(new_n245_) );
  XNOR2_X1 g123 ( .A(new_n239_), .B(new_n240_), .ZN(new_n246_) );
  NAND2_X1 g124 ( .A1(new_n246_), .A2(new_n243_), .ZN(new_n247_) );
  NAND2_X1 g125 ( .A1(new_n245_), .A2(new_n247_), .ZN(new_n248_) );
  NOR2_X1 g126 ( .A1(new_n248_), .A2(G902), .ZN(new_n249_) );
  XNOR2_X1 g127 ( .A(new_n249_), .B(G478), .ZN(new_n250_) );
  XOR2_X1 g128 ( .A(G140), .B(KEYINPUT11), .Z(new_n251_) );
  XNOR2_X1 g129 ( .A(G113), .B(G122), .ZN(new_n252_) );
  XNOR2_X1 g130 ( .A(new_n251_), .B(new_n252_), .ZN(new_n253_) );
  XNOR2_X1 g131 ( .A(G125), .B(KEYINPUT10), .ZN(new_n254_) );
  XNOR2_X1 g132 ( .A(new_n253_), .B(new_n254_), .ZN(new_n255_) );
  XNOR2_X1 g133 ( .A(G104), .B(G143), .ZN(new_n256_) );
  XNOR2_X1 g134 ( .A(new_n255_), .B(new_n256_), .ZN(new_n257_) );
  XNOR2_X1 g135 ( .A(G131), .B(G146), .ZN(new_n258_) );
  XNOR2_X1 g136 ( .A(new_n258_), .B(KEYINPUT12), .ZN(new_n259_) );
  INV_X1 g137 ( .A(G237), .ZN(new_n260_) );
  NAND2_X1 g138 ( .A1(new_n260_), .A2(G214), .ZN(new_n261_) );
  NOR2_X1 g139 ( .A1(new_n261_), .A2(G953), .ZN(new_n262_) );
  XNOR2_X1 g140 ( .A(new_n259_), .B(new_n262_), .ZN(new_n263_) );
  XNOR2_X1 g141 ( .A(new_n257_), .B(new_n263_), .ZN(new_n264_) );
  NAND2_X1 g142 ( .A1(new_n264_), .A2(new_n210_), .ZN(new_n265_) );
  XOR2_X1 g143 ( .A(G475), .B(KEYINPUT13), .Z(new_n266_) );
  XNOR2_X1 g144 ( .A(new_n265_), .B(new_n266_), .ZN(new_n267_) );
  INV_X1 g145 ( .A(new_n267_), .ZN(new_n268_) );
  NAND2_X1 g146 ( .A1(new_n250_), .A2(new_n268_), .ZN(new_n269_) );
  NAND2_X1 g147 ( .A1(new_n188_), .A2(G234), .ZN(new_n270_) );
  XNOR2_X1 g148 ( .A(new_n270_), .B(KEYINPUT20), .ZN(new_n271_) );
  NAND2_X1 g149 ( .A1(new_n271_), .A2(G221), .ZN(new_n272_) );
  XOR2_X1 g150 ( .A(new_n272_), .B(KEYINPUT21), .Z(new_n273_) );
  INV_X1 g151 ( .A(new_n273_), .ZN(new_n274_) );
  NOR2_X1 g152 ( .A1(new_n269_), .A2(new_n274_), .ZN(new_n275_) );
  NAND2_X1 g153 ( .A1(new_n224_), .A2(new_n275_), .ZN(new_n276_) );
  XNOR2_X1 g154 ( .A(new_n276_), .B(new_n124_), .ZN(new_n277_) );
  INV_X1 g155 ( .A(KEYINPUT1), .ZN(new_n278_) );
  INV_X1 g156 ( .A(G469), .ZN(new_n279_) );
  INV_X1 g157 ( .A(G134), .ZN(new_n280_) );
  NAND2_X1 g158 ( .A1(new_n258_), .A2(new_n280_), .ZN(new_n281_) );
  NOR2_X1 g159 ( .A1(G131), .A2(G146), .ZN(new_n282_) );
  NAND2_X1 g160 ( .A1(G131), .A2(G146), .ZN(new_n283_) );
  INV_X1 g161 ( .A(new_n283_), .ZN(new_n284_) );
  NOR2_X1 g162 ( .A1(new_n284_), .A2(new_n282_), .ZN(new_n285_) );
  NAND2_X1 g163 ( .A1(new_n285_), .A2(G134), .ZN(new_n286_) );
  NAND2_X1 g164 ( .A1(new_n286_), .A2(new_n281_), .ZN(new_n287_) );
  XOR2_X1 g165 ( .A(G137), .B(G140), .Z(new_n288_) );
  NAND2_X1 g166 ( .A1(new_n287_), .A2(new_n288_), .ZN(new_n289_) );
  XNOR2_X1 g167 ( .A(new_n258_), .B(G134), .ZN(new_n290_) );
  XNOR2_X1 g168 ( .A(G137), .B(G140), .ZN(new_n291_) );
  NAND2_X1 g169 ( .A1(new_n290_), .A2(new_n291_), .ZN(new_n292_) );
  NAND2_X1 g170 ( .A1(new_n292_), .A2(new_n289_), .ZN(new_n293_) );
  NAND2_X1 g171 ( .A1(new_n148_), .A2(G227), .ZN(new_n294_) );
  INV_X1 g172 ( .A(new_n294_), .ZN(new_n295_) );
  XNOR2_X1 g173 ( .A(new_n293_), .B(new_n295_), .ZN(new_n296_) );
  NAND2_X1 g174 ( .A1(new_n296_), .A2(new_n184_), .ZN(new_n297_) );
  XNOR2_X1 g175 ( .A(new_n293_), .B(new_n294_), .ZN(new_n298_) );
  NAND2_X1 g176 ( .A1(new_n174_), .A2(new_n298_), .ZN(new_n299_) );
  NAND2_X1 g177 ( .A1(new_n299_), .A2(new_n297_), .ZN(new_n300_) );
  NOR2_X1 g178 ( .A1(new_n300_), .A2(G902), .ZN(new_n301_) );
  NAND2_X1 g179 ( .A1(new_n301_), .A2(new_n279_), .ZN(new_n302_) );
  XNOR2_X1 g180 ( .A(new_n298_), .B(new_n184_), .ZN(new_n303_) );
  NAND2_X1 g181 ( .A1(new_n303_), .A2(new_n210_), .ZN(new_n304_) );
  NAND2_X1 g182 ( .A1(new_n304_), .A2(G469), .ZN(new_n305_) );
  NAND2_X1 g183 ( .A1(new_n305_), .A2(new_n302_), .ZN(new_n306_) );
  XNOR2_X1 g184 ( .A(new_n306_), .B(new_n278_), .ZN(new_n307_) );
  NAND2_X1 g185 ( .A1(new_n277_), .A2(new_n307_), .ZN(new_n308_) );
  INV_X1 g186 ( .A(G472), .ZN(new_n309_) );
  XNOR2_X1 g187 ( .A(G137), .B(KEYINPUT5), .ZN(new_n310_) );
  NOR2_X1 g188 ( .A1(new_n190_), .A2(G237), .ZN(new_n311_) );
  NAND2_X1 g189 ( .A1(new_n311_), .A2(new_n148_), .ZN(new_n312_) );
  XNOR2_X1 g190 ( .A(new_n312_), .B(new_n310_), .ZN(new_n313_) );
  NAND2_X1 g191 ( .A1(new_n139_), .A2(new_n313_), .ZN(new_n314_) );
  NAND2_X1 g192 ( .A1(new_n260_), .A2(G210), .ZN(new_n315_) );
  NOR2_X1 g193 ( .A1(new_n315_), .A2(G953), .ZN(new_n316_) );
  NAND2_X1 g194 ( .A1(new_n316_), .A2(new_n310_), .ZN(new_n317_) );
  XOR2_X1 g195 ( .A(G137), .B(KEYINPUT5), .Z(new_n318_) );
  NAND2_X1 g196 ( .A1(new_n318_), .A2(new_n312_), .ZN(new_n319_) );
  NAND2_X1 g197 ( .A1(new_n319_), .A2(new_n317_), .ZN(new_n320_) );
  NAND2_X1 g198 ( .A1(new_n136_), .A2(new_n320_), .ZN(new_n321_) );
  NAND2_X1 g199 ( .A1(new_n314_), .A2(new_n321_), .ZN(new_n322_) );
  NAND2_X1 g200 ( .A1(new_n322_), .A2(new_n287_), .ZN(new_n323_) );
  XNOR2_X1 g201 ( .A(new_n313_), .B(new_n136_), .ZN(new_n324_) );
  NAND2_X1 g202 ( .A1(new_n324_), .A2(new_n290_), .ZN(new_n325_) );
  NAND2_X1 g203 ( .A1(new_n325_), .A2(new_n323_), .ZN(new_n326_) );
  NAND2_X1 g204 ( .A1(new_n326_), .A2(new_n169_), .ZN(new_n327_) );
  XNOR2_X1 g205 ( .A(new_n322_), .B(new_n290_), .ZN(new_n328_) );
  NAND2_X1 g206 ( .A1(new_n328_), .A2(new_n182_), .ZN(new_n329_) );
  NAND2_X1 g207 ( .A1(new_n329_), .A2(new_n327_), .ZN(new_n330_) );
  NOR2_X1 g208 ( .A1(new_n330_), .A2(G902), .ZN(new_n331_) );
  XNOR2_X1 g209 ( .A(new_n331_), .B(new_n309_), .ZN(new_n332_) );
  XNOR2_X1 g210 ( .A(new_n332_), .B(KEYINPUT6), .ZN(new_n333_) );
  NAND2_X1 g211 ( .A1(new_n271_), .A2(G217), .ZN(new_n334_) );
  INV_X1 g212 ( .A(new_n334_), .ZN(new_n335_) );
  XNOR2_X1 g213 ( .A(G110), .B(G128), .ZN(new_n336_) );
  XNOR2_X1 g214 ( .A(G119), .B(G146), .ZN(new_n337_) );
  XNOR2_X1 g215 ( .A(new_n336_), .B(new_n337_), .ZN(new_n338_) );
  XNOR2_X1 g216 ( .A(new_n288_), .B(new_n254_), .ZN(new_n339_) );
  NAND2_X1 g217 ( .A1(new_n339_), .A2(new_n338_), .ZN(new_n340_) );
  XOR2_X1 g218 ( .A(new_n336_), .B(new_n337_), .Z(new_n341_) );
  XNOR2_X1 g219 ( .A(new_n254_), .B(new_n291_), .ZN(new_n342_) );
  NAND2_X1 g220 ( .A1(new_n341_), .A2(new_n342_), .ZN(new_n343_) );
  NAND2_X1 g221 ( .A1(new_n343_), .A2(new_n340_), .ZN(new_n344_) );
  NAND2_X1 g222 ( .A1(new_n231_), .A2(G221), .ZN(new_n345_) );
  XOR2_X1 g223 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(new_n346_) );
  XNOR2_X1 g224 ( .A(new_n345_), .B(new_n346_), .ZN(new_n347_) );
  INV_X1 g225 ( .A(new_n347_), .ZN(new_n348_) );
  XNOR2_X1 g226 ( .A(new_n348_), .B(new_n344_), .ZN(new_n349_) );
  NAND2_X1 g227 ( .A1(new_n349_), .A2(new_n210_), .ZN(new_n350_) );
  NAND2_X1 g228 ( .A1(new_n350_), .A2(new_n335_), .ZN(new_n351_) );
  XNOR2_X1 g229 ( .A(new_n344_), .B(new_n347_), .ZN(new_n352_) );
  NOR2_X1 g230 ( .A1(new_n352_), .A2(G902), .ZN(new_n353_) );
  NAND2_X1 g231 ( .A1(new_n353_), .A2(new_n334_), .ZN(new_n354_) );
  NAND2_X1 g232 ( .A1(new_n354_), .A2(new_n351_), .ZN(new_n355_) );
  XNOR2_X1 g233 ( .A(new_n355_), .B(KEYINPUT25), .ZN(new_n356_) );
  NAND2_X1 g234 ( .A1(new_n333_), .A2(new_n356_), .ZN(new_n357_) );
  NOR2_X1 g235 ( .A1(new_n308_), .A2(new_n357_), .ZN(new_n358_) );
  XNOR2_X1 g236 ( .A(new_n358_), .B(new_n123_), .ZN(G3) );
  INV_X1 g237 ( .A(new_n224_), .ZN(new_n360_) );
  XNOR2_X1 g238 ( .A(new_n301_), .B(G469), .ZN(new_n361_) );
  NAND2_X1 g239 ( .A1(new_n356_), .A2(new_n273_), .ZN(new_n362_) );
  NOR2_X1 g240 ( .A1(new_n362_), .A2(new_n361_), .ZN(new_n363_) );
  INV_X1 g241 ( .A(new_n363_), .ZN(new_n364_) );
  NOR2_X1 g242 ( .A1(new_n364_), .A2(new_n332_), .ZN(new_n365_) );
  INV_X1 g243 ( .A(new_n365_), .ZN(new_n366_) );
  NOR2_X1 g244 ( .A1(new_n360_), .A2(new_n366_), .ZN(new_n367_) );
  INV_X1 g245 ( .A(G478), .ZN(new_n368_) );
  NAND2_X1 g246 ( .A1(new_n249_), .A2(new_n368_), .ZN(new_n369_) );
  XNOR2_X1 g247 ( .A(new_n246_), .B(new_n244_), .ZN(new_n370_) );
  NAND2_X1 g248 ( .A1(new_n370_), .A2(new_n210_), .ZN(new_n371_) );
  NAND2_X1 g249 ( .A1(new_n371_), .A2(G478), .ZN(new_n372_) );
  NAND2_X1 g250 ( .A1(new_n372_), .A2(new_n369_), .ZN(new_n373_) );
  NOR2_X1 g251 ( .A1(new_n268_), .A2(new_n373_), .ZN(new_n374_) );
  NAND2_X1 g252 ( .A1(new_n367_), .A2(new_n374_), .ZN(new_n375_) );
  XNOR2_X1 g253 ( .A(new_n375_), .B(G104), .ZN(G6) );
  NOR2_X1 g254 ( .A1(new_n250_), .A2(new_n267_), .ZN(new_n377_) );
  NAND2_X1 g255 ( .A1(new_n367_), .A2(new_n377_), .ZN(new_n378_) );
  XOR2_X1 g256 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(new_n379_) );
  XNOR2_X1 g257 ( .A(new_n378_), .B(new_n379_), .ZN(new_n380_) );
  XNOR2_X1 g258 ( .A(new_n380_), .B(G107), .ZN(G9) );
  NOR2_X1 g259 ( .A1(new_n356_), .A2(new_n332_), .ZN(new_n382_) );
  INV_X1 g260 ( .A(new_n382_), .ZN(new_n383_) );
  NOR2_X1 g261 ( .A1(new_n308_), .A2(new_n383_), .ZN(new_n384_) );
  XOR2_X1 g262 ( .A(new_n384_), .B(G110), .Z(G12) );
  INV_X1 g263 ( .A(new_n377_), .ZN(new_n386_) );
  NAND2_X1 g264 ( .A1(new_n331_), .A2(G472), .ZN(new_n387_) );
  XNOR2_X1 g265 ( .A(new_n326_), .B(new_n182_), .ZN(new_n388_) );
  NAND2_X1 g266 ( .A1(new_n388_), .A2(new_n210_), .ZN(new_n389_) );
  NAND2_X1 g267 ( .A1(new_n389_), .A2(new_n309_), .ZN(new_n390_) );
  NAND2_X1 g268 ( .A1(new_n390_), .A2(new_n387_), .ZN(new_n391_) );
  INV_X1 g269 ( .A(KEYINPUT25), .ZN(new_n392_) );
  XNOR2_X1 g270 ( .A(new_n355_), .B(new_n392_), .ZN(new_n393_) );
  NOR2_X1 g271 ( .A1(new_n148_), .A2(G900), .ZN(new_n394_) );
  NAND2_X1 g272 ( .A1(new_n211_), .A2(new_n394_), .ZN(new_n395_) );
  INV_X1 g273 ( .A(new_n395_), .ZN(new_n396_) );
  NOR2_X1 g274 ( .A1(new_n209_), .A2(new_n396_), .ZN(new_n397_) );
  NOR2_X1 g275 ( .A1(new_n274_), .A2(new_n397_), .ZN(new_n398_) );
  NAND2_X1 g276 ( .A1(new_n393_), .A2(new_n398_), .ZN(new_n399_) );
  NOR2_X1 g277 ( .A1(new_n399_), .A2(new_n391_), .ZN(new_n400_) );
  INV_X1 g278 ( .A(new_n400_), .ZN(new_n401_) );
  NOR2_X1 g279 ( .A1(new_n401_), .A2(KEYINPUT28), .ZN(new_n402_) );
  NAND2_X1 g280 ( .A1(new_n401_), .A2(KEYINPUT28), .ZN(new_n403_) );
  NAND2_X1 g281 ( .A1(new_n403_), .A2(new_n306_), .ZN(new_n404_) );
  NOR2_X1 g282 ( .A1(new_n404_), .A2(new_n402_), .ZN(new_n405_) );
  NAND2_X1 g283 ( .A1(new_n405_), .A2(new_n220_), .ZN(new_n406_) );
  NOR2_X1 g284 ( .A1(new_n406_), .A2(new_n386_), .ZN(new_n407_) );
  XNOR2_X1 g285 ( .A(G128), .B(KEYINPUT29), .ZN(new_n408_) );
  XNOR2_X1 g286 ( .A(new_n407_), .B(new_n408_), .ZN(G30) );
  INV_X1 g287 ( .A(KEYINPUT30), .ZN(new_n410_) );
  NAND2_X1 g288 ( .A1(new_n332_), .A2(new_n196_), .ZN(new_n411_) );
  NAND2_X1 g289 ( .A1(new_n411_), .A2(new_n410_), .ZN(new_n412_) );
  NOR2_X1 g290 ( .A1(new_n391_), .A2(new_n195_), .ZN(new_n413_) );
  NAND2_X1 g291 ( .A1(new_n413_), .A2(KEYINPUT30), .ZN(new_n414_) );
  NAND2_X1 g292 ( .A1(new_n412_), .A2(new_n414_), .ZN(new_n415_) );
  NAND2_X1 g293 ( .A1(new_n415_), .A2(new_n193_), .ZN(new_n416_) );
  NOR2_X1 g294 ( .A1(new_n250_), .A2(new_n268_), .ZN(new_n417_) );
  INV_X1 g295 ( .A(new_n417_), .ZN(new_n418_) );
  INV_X1 g296 ( .A(new_n397_), .ZN(new_n419_) );
  NAND2_X1 g297 ( .A1(new_n363_), .A2(new_n419_), .ZN(new_n420_) );
  NOR2_X1 g298 ( .A1(new_n418_), .A2(new_n420_), .ZN(new_n421_) );
  INV_X1 g299 ( .A(new_n421_), .ZN(new_n422_) );
  NOR2_X1 g300 ( .A1(new_n422_), .A2(new_n416_), .ZN(new_n423_) );
  XNOR2_X1 g301 ( .A(new_n423_), .B(new_n162_), .ZN(G45) );
  INV_X1 g302 ( .A(new_n374_), .ZN(new_n425_) );
  NOR2_X1 g303 ( .A1(new_n406_), .A2(new_n425_), .ZN(new_n426_) );
  XOR2_X1 g304 ( .A(new_n426_), .B(G146), .Z(G48) );
  NAND2_X1 g305 ( .A1(new_n306_), .A2(KEYINPUT1), .ZN(new_n428_) );
  NAND2_X1 g306 ( .A1(new_n361_), .A2(new_n278_), .ZN(new_n429_) );
  NAND2_X1 g307 ( .A1(new_n429_), .A2(new_n428_), .ZN(new_n430_) );
  NOR2_X1 g308 ( .A1(new_n393_), .A2(new_n274_), .ZN(new_n431_) );
  NAND2_X1 g309 ( .A1(new_n430_), .A2(new_n431_), .ZN(new_n432_) );
  NOR2_X1 g310 ( .A1(new_n432_), .A2(new_n391_), .ZN(new_n433_) );
  NAND2_X1 g311 ( .A1(new_n224_), .A2(new_n433_), .ZN(new_n434_) );
  XNOR2_X1 g312 ( .A(new_n434_), .B(KEYINPUT31), .ZN(new_n435_) );
  NAND2_X1 g313 ( .A1(new_n435_), .A2(new_n374_), .ZN(new_n436_) );
  XNOR2_X1 g314 ( .A(new_n436_), .B(G113), .ZN(G15) );
  NAND2_X1 g315 ( .A1(new_n435_), .A2(new_n377_), .ZN(new_n438_) );
  XNOR2_X1 g316 ( .A(new_n438_), .B(G116), .ZN(G18) );
  NOR2_X1 g317 ( .A1(new_n307_), .A2(new_n356_), .ZN(new_n440_) );
  NAND2_X1 g318 ( .A1(new_n440_), .A2(new_n333_), .ZN(new_n441_) );
  INV_X1 g319 ( .A(new_n441_), .ZN(new_n442_) );
  NAND2_X1 g320 ( .A1(new_n277_), .A2(new_n442_), .ZN(new_n443_) );
  NAND2_X1 g321 ( .A1(new_n443_), .A2(KEYINPUT32), .ZN(new_n444_) );
  INV_X1 g322 ( .A(KEYINPUT32), .ZN(new_n445_) );
  XNOR2_X1 g323 ( .A(new_n276_), .B(KEYINPUT22), .ZN(new_n446_) );
  NOR2_X1 g324 ( .A1(new_n446_), .A2(new_n441_), .ZN(new_n447_) );
  NAND2_X1 g325 ( .A1(new_n447_), .A2(new_n445_), .ZN(new_n448_) );
  NAND2_X1 g326 ( .A1(new_n448_), .A2(new_n444_), .ZN(new_n449_) );
  XNOR2_X1 g327 ( .A(new_n449_), .B(G119), .ZN(G21) );
  INV_X1 g328 ( .A(KEYINPUT35), .ZN(new_n451_) );
  INV_X1 g329 ( .A(KEYINPUT34), .ZN(new_n452_) );
  INV_X1 g330 ( .A(KEYINPUT33), .ZN(new_n453_) );
  NOR2_X1 g331 ( .A1(new_n432_), .A2(new_n333_), .ZN(new_n454_) );
  NAND2_X1 g332 ( .A1(new_n454_), .A2(new_n453_), .ZN(new_n455_) );
  XNOR2_X1 g333 ( .A(new_n391_), .B(KEYINPUT6), .ZN(new_n456_) );
  NOR2_X1 g334 ( .A1(new_n307_), .A2(new_n362_), .ZN(new_n457_) );
  NAND2_X1 g335 ( .A1(new_n457_), .A2(new_n456_), .ZN(new_n458_) );
  NAND2_X1 g336 ( .A1(new_n458_), .A2(KEYINPUT33), .ZN(new_n459_) );
  NAND2_X1 g337 ( .A1(new_n459_), .A2(new_n455_), .ZN(new_n460_) );
  NAND2_X1 g338 ( .A1(new_n224_), .A2(new_n460_), .ZN(new_n461_) );
  XNOR2_X1 g339 ( .A(new_n461_), .B(new_n452_), .ZN(new_n462_) );
  NAND2_X1 g340 ( .A1(new_n462_), .A2(new_n417_), .ZN(new_n463_) );
  XNOR2_X1 g341 ( .A(new_n463_), .B(new_n451_), .ZN(new_n464_) );
  XNOR2_X1 g342 ( .A(new_n464_), .B(G122), .ZN(G24) );
  NOR2_X1 g343 ( .A1(new_n333_), .A2(new_n399_), .ZN(new_n466_) );
  NAND2_X1 g344 ( .A1(new_n466_), .A2(new_n374_), .ZN(new_n467_) );
  NOR2_X1 g345 ( .A1(new_n467_), .A2(new_n197_), .ZN(new_n468_) );
  INV_X1 g346 ( .A(new_n468_), .ZN(new_n469_) );
  NOR2_X1 g347 ( .A1(new_n469_), .A2(KEYINPUT36), .ZN(new_n470_) );
  NAND2_X1 g348 ( .A1(new_n469_), .A2(KEYINPUT36), .ZN(new_n471_) );
  NAND2_X1 g349 ( .A1(new_n471_), .A2(new_n430_), .ZN(new_n472_) );
  NOR2_X1 g350 ( .A1(new_n472_), .A2(new_n470_), .ZN(new_n473_) );
  XNOR2_X1 g351 ( .A(new_n473_), .B(G125), .ZN(new_n474_) );
  XNOR2_X1 g352 ( .A(new_n474_), .B(KEYINPUT37), .ZN(G27) );
  INV_X1 g353 ( .A(KEYINPUT39), .ZN(new_n476_) );
  XNOR2_X1 g354 ( .A(new_n200_), .B(KEYINPUT38), .ZN(new_n477_) );
  NAND2_X1 g355 ( .A1(new_n415_), .A2(new_n477_), .ZN(new_n478_) );
  NOR2_X1 g356 ( .A1(new_n478_), .A2(new_n420_), .ZN(new_n479_) );
  XNOR2_X1 g357 ( .A(new_n479_), .B(new_n476_), .ZN(new_n480_) );
  NAND2_X1 g358 ( .A1(new_n480_), .A2(new_n374_), .ZN(new_n481_) );
  XNOR2_X1 g359 ( .A(new_n481_), .B(KEYINPUT40), .ZN(new_n482_) );
  XNOR2_X1 g360 ( .A(new_n482_), .B(G131), .ZN(G33) );
  XNOR2_X1 g361 ( .A(new_n479_), .B(KEYINPUT39), .ZN(new_n484_) );
  NOR2_X1 g362 ( .A1(new_n484_), .A2(new_n386_), .ZN(new_n485_) );
  XNOR2_X1 g363 ( .A(new_n485_), .B(new_n280_), .ZN(G36) );
  INV_X1 g364 ( .A(KEYINPUT42), .ZN(new_n487_) );
  INV_X1 g365 ( .A(new_n402_), .ZN(new_n488_) );
  INV_X1 g366 ( .A(new_n404_), .ZN(new_n489_) );
  NAND2_X1 g367 ( .A1(new_n489_), .A2(new_n488_), .ZN(new_n490_) );
  INV_X1 g368 ( .A(KEYINPUT41), .ZN(new_n491_) );
  NOR2_X1 g369 ( .A1(new_n269_), .A2(new_n195_), .ZN(new_n492_) );
  NAND2_X1 g370 ( .A1(new_n492_), .A2(new_n477_), .ZN(new_n493_) );
  NAND2_X1 g371 ( .A1(new_n493_), .A2(new_n491_), .ZN(new_n494_) );
  INV_X1 g372 ( .A(new_n477_), .ZN(new_n495_) );
  NOR2_X1 g373 ( .A1(new_n373_), .A2(new_n267_), .ZN(new_n496_) );
  NAND2_X1 g374 ( .A1(new_n496_), .A2(new_n196_), .ZN(new_n497_) );
  NOR2_X1 g375 ( .A1(new_n497_), .A2(new_n495_), .ZN(new_n498_) );
  NAND2_X1 g376 ( .A1(new_n498_), .A2(KEYINPUT41), .ZN(new_n499_) );
  NAND2_X1 g377 ( .A1(new_n494_), .A2(new_n499_), .ZN(new_n500_) );
  NOR2_X1 g378 ( .A1(new_n500_), .A2(new_n490_), .ZN(new_n501_) );
  XNOR2_X1 g379 ( .A(new_n501_), .B(new_n487_), .ZN(new_n502_) );
  XNOR2_X1 g380 ( .A(new_n502_), .B(G137), .ZN(G39) );
  INV_X1 g381 ( .A(KEYINPUT43), .ZN(new_n504_) );
  INV_X1 g382 ( .A(new_n467_), .ZN(new_n505_) );
  NOR2_X1 g383 ( .A1(new_n430_), .A2(new_n195_), .ZN(new_n506_) );
  NAND2_X1 g384 ( .A1(new_n505_), .A2(new_n506_), .ZN(new_n507_) );
  NOR2_X1 g385 ( .A1(new_n507_), .A2(new_n504_), .ZN(new_n508_) );
  NAND2_X1 g386 ( .A1(new_n507_), .A2(new_n504_), .ZN(new_n509_) );
  NAND2_X1 g387 ( .A1(new_n509_), .A2(new_n200_), .ZN(new_n510_) );
  NOR2_X1 g388 ( .A1(new_n510_), .A2(new_n508_), .ZN(new_n511_) );
  XOR2_X1 g389 ( .A(new_n511_), .B(G140), .Z(G42) );
  INV_X1 g390 ( .A(KEYINPUT45), .ZN(new_n513_) );
  INV_X1 g391 ( .A(new_n384_), .ZN(new_n514_) );
  NAND2_X1 g392 ( .A1(new_n449_), .A2(new_n514_), .ZN(new_n515_) );
  NAND2_X1 g393 ( .A1(new_n515_), .A2(KEYINPUT44), .ZN(new_n516_) );
  INV_X1 g394 ( .A(KEYINPUT44), .ZN(new_n517_) );
  NAND2_X1 g395 ( .A1(new_n464_), .A2(new_n517_), .ZN(new_n518_) );
  NOR2_X1 g396 ( .A1(new_n518_), .A2(new_n515_), .ZN(new_n519_) );
  NAND2_X1 g397 ( .A1(new_n463_), .A2(KEYINPUT35), .ZN(new_n520_) );
  XNOR2_X1 g398 ( .A(new_n461_), .B(KEYINPUT34), .ZN(new_n521_) );
  NOR2_X1 g399 ( .A1(new_n521_), .A2(new_n418_), .ZN(new_n522_) );
  NAND2_X1 g400 ( .A1(new_n522_), .A2(new_n451_), .ZN(new_n523_) );
  NAND2_X1 g401 ( .A1(new_n523_), .A2(new_n520_), .ZN(new_n524_) );
  NAND2_X1 g402 ( .A1(new_n524_), .A2(KEYINPUT44), .ZN(new_n525_) );
  NOR2_X1 g403 ( .A1(new_n377_), .A2(new_n374_), .ZN(new_n526_) );
  NOR2_X1 g404 ( .A1(new_n435_), .A2(new_n367_), .ZN(new_n527_) );
  NOR2_X1 g405 ( .A1(new_n527_), .A2(new_n526_), .ZN(new_n528_) );
  NOR2_X1 g406 ( .A1(new_n528_), .A2(new_n358_), .ZN(new_n529_) );
  NAND2_X1 g407 ( .A1(new_n525_), .A2(new_n529_), .ZN(new_n530_) );
  NOR2_X1 g408 ( .A1(new_n519_), .A2(new_n530_), .ZN(new_n531_) );
  NAND2_X1 g409 ( .A1(new_n531_), .A2(new_n516_), .ZN(new_n532_) );
  NOR2_X1 g410 ( .A1(new_n532_), .A2(new_n513_), .ZN(new_n533_) );
  NAND2_X1 g411 ( .A1(new_n482_), .A2(new_n502_), .ZN(new_n534_) );
  NOR2_X1 g412 ( .A1(new_n534_), .A2(KEYINPUT46), .ZN(new_n535_) );
  INV_X1 g413 ( .A(new_n535_), .ZN(new_n536_) );
  INV_X1 g414 ( .A(KEYINPUT46), .ZN(new_n537_) );
  INV_X1 g415 ( .A(KEYINPUT40), .ZN(new_n538_) );
  NAND2_X1 g416 ( .A1(new_n481_), .A2(new_n538_), .ZN(new_n539_) );
  NOR2_X1 g417 ( .A1(new_n484_), .A2(new_n425_), .ZN(new_n540_) );
  NAND2_X1 g418 ( .A1(new_n540_), .A2(KEYINPUT40), .ZN(new_n541_) );
  NAND2_X1 g419 ( .A1(new_n541_), .A2(new_n539_), .ZN(new_n542_) );
  XNOR2_X1 g420 ( .A(new_n498_), .B(new_n491_), .ZN(new_n543_) );
  NAND2_X1 g421 ( .A1(new_n543_), .A2(new_n405_), .ZN(new_n544_) );
  NAND2_X1 g422 ( .A1(new_n544_), .A2(new_n487_), .ZN(new_n545_) );
  NAND2_X1 g423 ( .A1(new_n501_), .A2(KEYINPUT42), .ZN(new_n546_) );
  NAND2_X1 g424 ( .A1(new_n545_), .A2(new_n546_), .ZN(new_n547_) );
  NOR2_X1 g425 ( .A1(new_n542_), .A2(new_n547_), .ZN(new_n548_) );
  NOR2_X1 g426 ( .A1(new_n548_), .A2(new_n537_), .ZN(new_n549_) );
  NOR2_X1 g427 ( .A1(new_n473_), .A2(new_n423_), .ZN(new_n550_) );
  NOR2_X1 g428 ( .A1(new_n406_), .A2(new_n526_), .ZN(new_n551_) );
  XNOR2_X1 g429 ( .A(new_n551_), .B(KEYINPUT47), .ZN(new_n552_) );
  NAND2_X1 g430 ( .A1(new_n552_), .A2(new_n550_), .ZN(new_n553_) );
  NOR2_X1 g431 ( .A1(new_n549_), .A2(new_n553_), .ZN(new_n554_) );
  NAND2_X1 g432 ( .A1(new_n554_), .A2(new_n536_), .ZN(new_n555_) );
  NOR2_X1 g433 ( .A1(new_n555_), .A2(KEYINPUT48), .ZN(new_n556_) );
  NAND2_X1 g434 ( .A1(new_n555_), .A2(KEYINPUT48), .ZN(new_n557_) );
  NOR2_X1 g435 ( .A1(new_n511_), .A2(new_n485_), .ZN(new_n558_) );
  NAND2_X1 g436 ( .A1(new_n557_), .A2(new_n558_), .ZN(new_n559_) );
  NOR2_X1 g437 ( .A1(new_n559_), .A2(new_n556_), .ZN(new_n560_) );
  NAND2_X1 g438 ( .A1(new_n532_), .A2(new_n513_), .ZN(new_n561_) );
  NAND2_X1 g439 ( .A1(new_n561_), .A2(new_n560_), .ZN(new_n562_) );
  NOR2_X1 g440 ( .A1(new_n562_), .A2(new_n533_), .ZN(new_n563_) );
  NAND2_X1 g441 ( .A1(new_n563_), .A2(KEYINPUT2), .ZN(new_n564_) );
  INV_X1 g442 ( .A(KEYINPUT2), .ZN(new_n565_) );
  INV_X1 g443 ( .A(new_n533_), .ZN(new_n566_) );
  INV_X1 g444 ( .A(new_n556_), .ZN(new_n567_) );
  INV_X1 g445 ( .A(KEYINPUT48), .ZN(new_n568_) );
  NAND2_X1 g446 ( .A1(new_n534_), .A2(KEYINPUT46), .ZN(new_n569_) );
  INV_X1 g447 ( .A(new_n553_), .ZN(new_n570_) );
  NAND2_X1 g448 ( .A1(new_n569_), .A2(new_n570_), .ZN(new_n571_) );
  NOR2_X1 g449 ( .A1(new_n571_), .A2(new_n535_), .ZN(new_n572_) );
  NOR2_X1 g450 ( .A1(new_n572_), .A2(new_n568_), .ZN(new_n573_) );
  INV_X1 g451 ( .A(new_n558_), .ZN(new_n574_) );
  NOR2_X1 g452 ( .A1(new_n573_), .A2(new_n574_), .ZN(new_n575_) );
  NAND2_X1 g453 ( .A1(new_n575_), .A2(new_n567_), .ZN(new_n576_) );
  INV_X1 g454 ( .A(new_n516_), .ZN(new_n577_) );
  XNOR2_X1 g455 ( .A(new_n443_), .B(new_n445_), .ZN(new_n578_) );
  NOR2_X1 g456 ( .A1(new_n578_), .A2(new_n384_), .ZN(new_n579_) );
  NOR2_X1 g457 ( .A1(new_n524_), .A2(KEYINPUT44), .ZN(new_n580_) );
  NAND2_X1 g458 ( .A1(new_n579_), .A2(new_n580_), .ZN(new_n581_) );
  INV_X1 g459 ( .A(new_n530_), .ZN(new_n582_) );
  NAND2_X1 g460 ( .A1(new_n582_), .A2(new_n581_), .ZN(new_n583_) );
  NOR2_X1 g461 ( .A1(new_n583_), .A2(new_n577_), .ZN(new_n584_) );
  NOR2_X1 g462 ( .A1(new_n584_), .A2(KEYINPUT45), .ZN(new_n585_) );
  NOR2_X1 g463 ( .A1(new_n585_), .A2(new_n576_), .ZN(new_n586_) );
  NAND2_X1 g464 ( .A1(new_n586_), .A2(new_n566_), .ZN(new_n587_) );
  NAND2_X1 g465 ( .A1(new_n587_), .A2(new_n565_), .ZN(new_n588_) );
  NAND2_X1 g466 ( .A1(new_n588_), .A2(new_n564_), .ZN(new_n589_) );
  NOR2_X1 g467 ( .A1(new_n430_), .A2(new_n431_), .ZN(new_n590_) );
  NOR2_X1 g468 ( .A1(new_n590_), .A2(KEYINPUT50), .ZN(new_n591_) );
  NAND2_X1 g469 ( .A1(new_n590_), .A2(KEYINPUT50), .ZN(new_n592_) );
  NAND2_X1 g470 ( .A1(new_n393_), .A2(new_n274_), .ZN(new_n593_) );
  XNOR2_X1 g471 ( .A(new_n593_), .B(KEYINPUT49), .ZN(new_n594_) );
  NOR2_X1 g472 ( .A1(new_n594_), .A2(new_n332_), .ZN(new_n595_) );
  NAND2_X1 g473 ( .A1(new_n595_), .A2(new_n592_), .ZN(new_n596_) );
  NOR2_X1 g474 ( .A1(new_n596_), .A2(new_n591_), .ZN(new_n597_) );
  NOR2_X1 g475 ( .A1(new_n597_), .A2(new_n433_), .ZN(new_n598_) );
  INV_X1 g476 ( .A(new_n598_), .ZN(new_n599_) );
  NOR2_X1 g477 ( .A1(new_n599_), .A2(KEYINPUT51), .ZN(new_n600_) );
  NAND2_X1 g478 ( .A1(new_n599_), .A2(KEYINPUT51), .ZN(new_n601_) );
  NAND2_X1 g479 ( .A1(new_n601_), .A2(new_n543_), .ZN(new_n602_) );
  NOR2_X1 g480 ( .A1(new_n602_), .A2(new_n600_), .ZN(new_n603_) );
  NOR2_X1 g481 ( .A1(new_n526_), .A2(new_n195_), .ZN(new_n604_) );
  NOR2_X1 g482 ( .A1(new_n604_), .A2(new_n496_), .ZN(new_n605_) );
  NAND2_X1 g483 ( .A1(new_n497_), .A2(new_n495_), .ZN(new_n606_) );
  NAND2_X1 g484 ( .A1(new_n460_), .A2(new_n606_), .ZN(new_n607_) );
  NOR2_X1 g485 ( .A1(new_n607_), .A2(new_n605_), .ZN(new_n608_) );
  NOR2_X1 g486 ( .A1(new_n603_), .A2(new_n608_), .ZN(new_n609_) );
  NOR2_X1 g487 ( .A1(new_n609_), .A2(KEYINPUT52), .ZN(new_n610_) );
  NAND2_X1 g488 ( .A1(new_n609_), .A2(KEYINPUT52), .ZN(new_n611_) );
  NAND2_X1 g489 ( .A1(new_n611_), .A2(new_n207_), .ZN(new_n612_) );
  NOR2_X1 g490 ( .A1(new_n612_), .A2(new_n610_), .ZN(new_n613_) );
  NAND2_X1 g491 ( .A1(new_n543_), .A2(new_n460_), .ZN(new_n614_) );
  NAND2_X1 g492 ( .A1(new_n614_), .A2(new_n148_), .ZN(new_n615_) );
  NOR2_X1 g493 ( .A1(new_n613_), .A2(new_n615_), .ZN(new_n616_) );
  NAND2_X1 g494 ( .A1(new_n589_), .A2(new_n616_), .ZN(new_n617_) );
  XOR2_X1 g495 ( .A(new_n617_), .B(KEYINPUT53), .Z(G75) );
  INV_X1 g496 ( .A(KEYINPUT56), .ZN(new_n619_) );
  XNOR2_X1 g497 ( .A(new_n563_), .B(new_n565_), .ZN(new_n620_) );
  NOR2_X1 g498 ( .A1(new_n188_), .A2(new_n190_), .ZN(new_n621_) );
  NAND2_X1 g499 ( .A1(new_n620_), .A2(new_n621_), .ZN(new_n622_) );
  XNOR2_X1 g500 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(new_n623_) );
  XNOR2_X1 g501 ( .A(new_n186_), .B(new_n623_), .ZN(new_n624_) );
  NOR2_X1 g502 ( .A1(new_n622_), .A2(new_n624_), .ZN(new_n625_) );
  INV_X1 g503 ( .A(new_n625_), .ZN(new_n626_) );
  INV_X1 g504 ( .A(new_n621_), .ZN(new_n627_) );
  NOR2_X1 g505 ( .A1(new_n589_), .A2(new_n627_), .ZN(new_n628_) );
  INV_X1 g506 ( .A(new_n624_), .ZN(new_n629_) );
  NOR2_X1 g507 ( .A1(new_n628_), .A2(new_n629_), .ZN(new_n630_) );
  NOR2_X1 g508 ( .A1(new_n148_), .A2(G952), .ZN(new_n631_) );
  NOR2_X1 g509 ( .A1(new_n630_), .A2(new_n631_), .ZN(new_n632_) );
  NAND2_X1 g510 ( .A1(new_n632_), .A2(new_n626_), .ZN(new_n633_) );
  NAND2_X1 g511 ( .A1(new_n633_), .A2(new_n619_), .ZN(new_n634_) );
  NAND2_X1 g512 ( .A1(new_n622_), .A2(new_n624_), .ZN(new_n635_) );
  INV_X1 g513 ( .A(new_n631_), .ZN(new_n636_) );
  NAND2_X1 g514 ( .A1(new_n635_), .A2(new_n636_), .ZN(new_n637_) );
  NOR2_X1 g515 ( .A1(new_n637_), .A2(new_n625_), .ZN(new_n638_) );
  NAND2_X1 g516 ( .A1(new_n638_), .A2(KEYINPUT56), .ZN(new_n639_) );
  NAND2_X1 g517 ( .A1(new_n634_), .A2(new_n639_), .ZN(G51) );
  NOR2_X1 g518 ( .A1(new_n188_), .A2(new_n279_), .ZN(new_n641_) );
  INV_X1 g519 ( .A(new_n641_), .ZN(new_n642_) );
  NOR2_X1 g520 ( .A1(new_n589_), .A2(new_n642_), .ZN(new_n643_) );
  XOR2_X1 g521 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(new_n644_) );
  INV_X1 g522 ( .A(new_n644_), .ZN(new_n645_) );
  NAND2_X1 g523 ( .A1(new_n643_), .A2(new_n645_), .ZN(new_n646_) );
  NAND2_X1 g524 ( .A1(new_n620_), .A2(new_n641_), .ZN(new_n647_) );
  NAND2_X1 g525 ( .A1(new_n647_), .A2(new_n644_), .ZN(new_n648_) );
  NAND2_X1 g526 ( .A1(new_n648_), .A2(new_n646_), .ZN(new_n649_) );
  NOR2_X1 g527 ( .A1(new_n649_), .A2(new_n300_), .ZN(new_n650_) );
  NAND2_X1 g528 ( .A1(new_n649_), .A2(new_n300_), .ZN(new_n651_) );
  NAND2_X1 g529 ( .A1(new_n651_), .A2(new_n636_), .ZN(new_n652_) );
  NOR2_X1 g530 ( .A1(new_n652_), .A2(new_n650_), .ZN(G54) );
  INV_X1 g531 ( .A(KEYINPUT60), .ZN(new_n654_) );
  NAND2_X1 g532 ( .A1(new_n187_), .A2(G475), .ZN(new_n655_) );
  INV_X1 g533 ( .A(new_n655_), .ZN(new_n656_) );
  NAND2_X1 g534 ( .A1(new_n620_), .A2(new_n656_), .ZN(new_n657_) );
  XNOR2_X1 g535 ( .A(new_n264_), .B(KEYINPUT59), .ZN(new_n658_) );
  NOR2_X1 g536 ( .A1(new_n657_), .A2(new_n658_), .ZN(new_n659_) );
  INV_X1 g537 ( .A(new_n659_), .ZN(new_n660_) );
  NOR2_X1 g538 ( .A1(new_n589_), .A2(new_n655_), .ZN(new_n661_) );
  INV_X1 g539 ( .A(new_n658_), .ZN(new_n662_) );
  NOR2_X1 g540 ( .A1(new_n661_), .A2(new_n662_), .ZN(new_n663_) );
  NOR2_X1 g541 ( .A1(new_n663_), .A2(new_n631_), .ZN(new_n664_) );
  NAND2_X1 g542 ( .A1(new_n664_), .A2(new_n660_), .ZN(new_n665_) );
  NAND2_X1 g543 ( .A1(new_n665_), .A2(new_n654_), .ZN(new_n666_) );
  NAND2_X1 g544 ( .A1(new_n657_), .A2(new_n658_), .ZN(new_n667_) );
  NAND2_X1 g545 ( .A1(new_n667_), .A2(new_n636_), .ZN(new_n668_) );
  NOR2_X1 g546 ( .A1(new_n668_), .A2(new_n659_), .ZN(new_n669_) );
  NAND2_X1 g547 ( .A1(new_n669_), .A2(KEYINPUT60), .ZN(new_n670_) );
  NAND2_X1 g548 ( .A1(new_n666_), .A2(new_n670_), .ZN(G60) );
  NOR2_X1 g549 ( .A1(new_n188_), .A2(new_n368_), .ZN(new_n672_) );
  NAND2_X1 g550 ( .A1(new_n620_), .A2(new_n672_), .ZN(new_n673_) );
  NOR2_X1 g551 ( .A1(new_n673_), .A2(new_n248_), .ZN(new_n674_) );
  NAND2_X1 g552 ( .A1(new_n673_), .A2(new_n248_), .ZN(new_n675_) );
  NAND2_X1 g553 ( .A1(new_n675_), .A2(new_n636_), .ZN(new_n676_) );
  NOR2_X1 g554 ( .A1(new_n676_), .A2(new_n674_), .ZN(G63) );
  INV_X1 g555 ( .A(G217), .ZN(new_n678_) );
  NOR2_X1 g556 ( .A1(new_n188_), .A2(new_n678_), .ZN(new_n679_) );
  NAND2_X1 g557 ( .A1(new_n620_), .A2(new_n679_), .ZN(new_n680_) );
  NOR2_X1 g558 ( .A1(new_n680_), .A2(new_n352_), .ZN(new_n681_) );
  NAND2_X1 g559 ( .A1(new_n680_), .A2(new_n352_), .ZN(new_n682_) );
  NAND2_X1 g560 ( .A1(new_n682_), .A2(new_n636_), .ZN(new_n683_) );
  NOR2_X1 g561 ( .A1(new_n683_), .A2(new_n681_), .ZN(G66) );
  NOR2_X1 g562 ( .A1(new_n585_), .A2(G953), .ZN(new_n685_) );
  NAND2_X1 g563 ( .A1(new_n685_), .A2(new_n566_), .ZN(new_n686_) );
  INV_X1 g564 ( .A(KEYINPUT61), .ZN(new_n687_) );
  NAND2_X1 g565 ( .A1(G224), .A2(G953), .ZN(new_n688_) );
  NAND2_X1 g566 ( .A1(new_n688_), .A2(new_n687_), .ZN(new_n689_) );
  INV_X1 g567 ( .A(G898), .ZN(new_n690_) );
  NOR2_X1 g568 ( .A1(new_n688_), .A2(new_n687_), .ZN(new_n691_) );
  NOR2_X1 g569 ( .A1(new_n691_), .A2(new_n690_), .ZN(new_n692_) );
  NAND2_X1 g570 ( .A1(new_n692_), .A2(new_n689_), .ZN(new_n693_) );
  NAND2_X1 g571 ( .A1(new_n686_), .A2(new_n693_), .ZN(new_n694_) );
  XNOR2_X1 g572 ( .A(new_n172_), .B(G101), .ZN(new_n695_) );
  XNOR2_X1 g573 ( .A(new_n695_), .B(new_n142_), .ZN(new_n696_) );
  NOR2_X1 g574 ( .A1(new_n696_), .A2(new_n213_), .ZN(new_n697_) );
  XNOR2_X1 g575 ( .A(new_n694_), .B(new_n697_), .ZN(G69) );
  XOR2_X1 g576 ( .A(new_n168_), .B(new_n254_), .Z(new_n699_) );
  XNOR2_X1 g577 ( .A(new_n699_), .B(new_n293_), .ZN(new_n700_) );
  XNOR2_X1 g578 ( .A(new_n576_), .B(new_n700_), .ZN(new_n701_) );
  NAND2_X1 g579 ( .A1(new_n701_), .A2(new_n148_), .ZN(new_n702_) );
  XNOR2_X1 g580 ( .A(new_n700_), .B(G227), .ZN(new_n703_) );
  NAND2_X1 g581 ( .A1(new_n703_), .A2(G900), .ZN(new_n704_) );
  NAND2_X1 g582 ( .A1(new_n704_), .A2(G953), .ZN(new_n705_) );
  NAND2_X1 g583 ( .A1(new_n702_), .A2(new_n705_), .ZN(G72) );
  NOR2_X1 g584 ( .A1(new_n188_), .A2(new_n309_), .ZN(new_n707_) );
  NAND2_X1 g585 ( .A1(new_n620_), .A2(new_n707_), .ZN(new_n708_) );
  XNOR2_X1 g586 ( .A(new_n330_), .B(KEYINPUT62), .ZN(new_n709_) );
  NOR2_X1 g587 ( .A1(new_n708_), .A2(new_n709_), .ZN(new_n710_) );
  INV_X1 g588 ( .A(new_n710_), .ZN(new_n711_) );
  INV_X1 g589 ( .A(new_n707_), .ZN(new_n712_) );
  NOR2_X1 g590 ( .A1(new_n589_), .A2(new_n712_), .ZN(new_n713_) );
  INV_X1 g591 ( .A(new_n709_), .ZN(new_n714_) );
  NOR2_X1 g592 ( .A1(new_n713_), .A2(new_n714_), .ZN(new_n715_) );
  NOR2_X1 g593 ( .A1(new_n715_), .A2(new_n631_), .ZN(new_n716_) );
  NAND2_X1 g594 ( .A1(new_n716_), .A2(new_n711_), .ZN(new_n717_) );
  NAND2_X1 g595 ( .A1(new_n717_), .A2(KEYINPUT63), .ZN(new_n718_) );
  INV_X1 g596 ( .A(KEYINPUT63), .ZN(new_n719_) );
  NAND2_X1 g597 ( .A1(new_n708_), .A2(new_n709_), .ZN(new_n720_) );
  NAND2_X1 g598 ( .A1(new_n720_), .A2(new_n636_), .ZN(new_n721_) );
  NOR2_X1 g599 ( .A1(new_n721_), .A2(new_n710_), .ZN(new_n722_) );
  NAND2_X1 g600 ( .A1(new_n722_), .A2(new_n719_), .ZN(new_n723_) );
  NAND2_X1 g601 ( .A1(new_n718_), .A2(new_n723_), .ZN(G57) );
endmodule


