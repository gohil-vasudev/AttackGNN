module locked_c1908 (  G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,  G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n123_, new_n124_, new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_, new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_, new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n631_, new_n632_, new_n633_, new_n634_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n653_, new_n654_, new_n655_, new_n656_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_;
  INV_X1 g000 ( .A(G101), .ZN(new_n123_) );
  INV_X1 g001 ( .A(KEYINPUT22), .ZN(new_n124_) );
  INV_X1 g002 ( .A(KEYINPUT21), .ZN(new_n125_) );
  INV_X1 g003 ( .A(KEYINPUT20), .ZN(new_n126_) );
  OR2_X1 g004 ( .A1(G902), .A2(KEYINPUT15), .ZN(new_n127_) );
  AND2_X1 g005 ( .A1(G902), .A2(KEYINPUT15), .ZN(new_n128_) );
  INV_X1 g006 ( .A(new_n128_), .ZN(new_n129_) );
  AND2_X1 g007 ( .A1(new_n129_), .A2(new_n127_), .ZN(new_n130_) );
  INV_X1 g008 ( .A(new_n130_), .ZN(new_n131_) );
  AND2_X1 g009 ( .A1(new_n131_), .A2(G234), .ZN(new_n132_) );
  INV_X1 g010 ( .A(new_n132_), .ZN(new_n133_) );
  AND2_X1 g011 ( .A1(new_n133_), .A2(new_n126_), .ZN(new_n134_) );
  AND2_X1 g012 ( .A1(new_n132_), .A2(KEYINPUT20), .ZN(new_n135_) );
  OR2_X1 g013 ( .A1(new_n134_), .A2(new_n135_), .ZN(new_n136_) );
  INV_X1 g014 ( .A(new_n136_), .ZN(new_n137_) );
  AND2_X1 g015 ( .A1(new_n137_), .A2(G221), .ZN(new_n138_) );
  INV_X1 g016 ( .A(new_n138_), .ZN(new_n139_) );
  AND2_X1 g017 ( .A1(new_n139_), .A2(new_n125_), .ZN(new_n140_) );
  AND2_X1 g018 ( .A1(new_n138_), .A2(KEYINPUT21), .ZN(new_n141_) );
  OR2_X1 g019 ( .A1(new_n140_), .A2(new_n141_), .ZN(new_n142_) );
  INV_X1 g020 ( .A(G478), .ZN(new_n143_) );
  INV_X1 g021 ( .A(G116), .ZN(new_n144_) );
  INV_X1 g022 ( .A(G953), .ZN(new_n145_) );
  AND2_X1 g023 ( .A1(new_n145_), .A2(G234), .ZN(new_n146_) );
  OR2_X1 g024 ( .A1(new_n146_), .A2(KEYINPUT8), .ZN(new_n147_) );
  AND2_X1 g025 ( .A1(new_n146_), .A2(KEYINPUT8), .ZN(new_n148_) );
  INV_X1 g026 ( .A(new_n148_), .ZN(new_n149_) );
  AND2_X1 g027 ( .A1(new_n149_), .A2(new_n147_), .ZN(new_n150_) );
  INV_X1 g028 ( .A(new_n150_), .ZN(new_n151_) );
  AND2_X1 g029 ( .A1(new_n151_), .A2(G217), .ZN(new_n152_) );
  INV_X1 g030 ( .A(new_n152_), .ZN(new_n153_) );
  OR2_X1 g031 ( .A1(KEYINPUT9), .A2(KEYINPUT7), .ZN(new_n154_) );
  AND2_X1 g032 ( .A1(KEYINPUT9), .A2(KEYINPUT7), .ZN(new_n155_) );
  INV_X1 g033 ( .A(new_n155_), .ZN(new_n156_) );
  AND2_X1 g034 ( .A1(new_n156_), .A2(new_n154_), .ZN(new_n157_) );
  INV_X1 g035 ( .A(new_n157_), .ZN(new_n158_) );
  AND2_X1 g036 ( .A1(new_n153_), .A2(new_n158_), .ZN(new_n159_) );
  AND2_X1 g037 ( .A1(new_n152_), .A2(new_n157_), .ZN(new_n160_) );
  OR2_X1 g038 ( .A1(new_n159_), .A2(new_n160_), .ZN(new_n161_) );
  AND2_X1 g039 ( .A1(new_n161_), .A2(new_n144_), .ZN(new_n162_) );
  INV_X1 g040 ( .A(new_n162_), .ZN(new_n163_) );
  OR2_X1 g041 ( .A1(new_n161_), .A2(new_n144_), .ZN(new_n164_) );
  AND2_X1 g042 ( .A1(new_n163_), .A2(new_n164_), .ZN(new_n165_) );
  INV_X1 g043 ( .A(G107), .ZN(new_n166_) );
  INV_X1 g044 ( .A(G128), .ZN(new_n167_) );
  INV_X1 g045 ( .A(G143), .ZN(new_n168_) );
  AND2_X1 g046 ( .A1(new_n167_), .A2(new_n168_), .ZN(new_n169_) );
  AND2_X1 g047 ( .A1(G128), .A2(G143), .ZN(new_n170_) );
  OR2_X1 g048 ( .A1(new_n169_), .A2(new_n170_), .ZN(new_n171_) );
  AND2_X1 g049 ( .A1(new_n171_), .A2(new_n166_), .ZN(new_n172_) );
  OR2_X1 g050 ( .A1(G128), .A2(G143), .ZN(new_n173_) );
  INV_X1 g051 ( .A(new_n170_), .ZN(new_n174_) );
  AND2_X1 g052 ( .A1(new_n174_), .A2(new_n173_), .ZN(new_n175_) );
  AND2_X1 g053 ( .A1(new_n175_), .A2(G107), .ZN(new_n176_) );
  OR2_X1 g054 ( .A1(new_n172_), .A2(new_n176_), .ZN(new_n177_) );
  INV_X1 g055 ( .A(new_n177_), .ZN(new_n178_) );
  OR2_X1 g056 ( .A1(new_n165_), .A2(new_n178_), .ZN(new_n179_) );
  AND2_X1 g057 ( .A1(new_n165_), .A2(new_n178_), .ZN(new_n180_) );
  INV_X1 g058 ( .A(new_n180_), .ZN(new_n181_) );
  AND2_X1 g059 ( .A1(new_n181_), .A2(new_n179_), .ZN(new_n182_) );
  INV_X1 g060 ( .A(G134), .ZN(new_n183_) );
  AND2_X1 g061 ( .A1(new_n183_), .A2(G122), .ZN(new_n184_) );
  INV_X1 g062 ( .A(G122), .ZN(new_n185_) );
  AND2_X1 g063 ( .A1(new_n185_), .A2(G134), .ZN(new_n186_) );
  OR2_X1 g064 ( .A1(new_n184_), .A2(new_n186_), .ZN(new_n187_) );
  INV_X1 g065 ( .A(new_n187_), .ZN(new_n188_) );
  OR2_X1 g066 ( .A1(new_n182_), .A2(new_n188_), .ZN(new_n189_) );
  AND2_X1 g067 ( .A1(new_n182_), .A2(new_n188_), .ZN(new_n190_) );
  INV_X1 g068 ( .A(new_n190_), .ZN(new_n191_) );
  AND2_X1 g069 ( .A1(new_n191_), .A2(new_n189_), .ZN(new_n192_) );
  OR2_X1 g070 ( .A1(new_n192_), .A2(G902), .ZN(new_n193_) );
  AND2_X1 g071 ( .A1(new_n193_), .A2(new_n143_), .ZN(new_n194_) );
  INV_X1 g072 ( .A(G902), .ZN(new_n195_) );
  INV_X1 g073 ( .A(new_n179_), .ZN(new_n196_) );
  OR2_X1 g074 ( .A1(new_n196_), .A2(new_n180_), .ZN(new_n197_) );
  AND2_X1 g075 ( .A1(new_n197_), .A2(new_n187_), .ZN(new_n198_) );
  OR2_X1 g076 ( .A1(new_n198_), .A2(new_n190_), .ZN(new_n199_) );
  AND2_X1 g077 ( .A1(new_n199_), .A2(new_n195_), .ZN(new_n200_) );
  AND2_X1 g078 ( .A1(new_n200_), .A2(G478), .ZN(new_n201_) );
  OR2_X1 g079 ( .A1(new_n194_), .A2(new_n201_), .ZN(new_n202_) );
  INV_X1 g080 ( .A(G125), .ZN(new_n203_) );
  AND2_X1 g081 ( .A1(new_n203_), .A2(KEYINPUT10), .ZN(new_n204_) );
  INV_X1 g082 ( .A(KEYINPUT10), .ZN(new_n205_) );
  AND2_X1 g083 ( .A1(new_n205_), .A2(G125), .ZN(new_n206_) );
  OR2_X1 g084 ( .A1(new_n204_), .A2(new_n206_), .ZN(new_n207_) );
  INV_X1 g085 ( .A(G140), .ZN(new_n208_) );
  AND2_X1 g086 ( .A1(new_n208_), .A2(KEYINPUT11), .ZN(new_n209_) );
  INV_X1 g087 ( .A(new_n209_), .ZN(new_n210_) );
  OR2_X1 g088 ( .A1(new_n208_), .A2(KEYINPUT11), .ZN(new_n211_) );
  AND2_X1 g089 ( .A1(new_n210_), .A2(new_n211_), .ZN(new_n212_) );
  INV_X1 g090 ( .A(new_n212_), .ZN(new_n213_) );
  INV_X1 g091 ( .A(G113), .ZN(new_n214_) );
  AND2_X1 g092 ( .A1(new_n214_), .A2(new_n185_), .ZN(new_n215_) );
  AND2_X1 g093 ( .A1(G113), .A2(G122), .ZN(new_n216_) );
  OR2_X1 g094 ( .A1(new_n215_), .A2(new_n216_), .ZN(new_n217_) );
  AND2_X1 g095 ( .A1(new_n213_), .A2(new_n217_), .ZN(new_n218_) );
  INV_X1 g096 ( .A(new_n218_), .ZN(new_n219_) );
  OR2_X1 g097 ( .A1(new_n213_), .A2(new_n217_), .ZN(new_n220_) );
  AND2_X1 g098 ( .A1(new_n219_), .A2(new_n220_), .ZN(new_n221_) );
  INV_X1 g099 ( .A(new_n221_), .ZN(new_n222_) );
  AND2_X1 g100 ( .A1(new_n222_), .A2(new_n207_), .ZN(new_n223_) );
  INV_X1 g101 ( .A(new_n207_), .ZN(new_n224_) );
  AND2_X1 g102 ( .A1(new_n221_), .A2(new_n224_), .ZN(new_n225_) );
  OR2_X1 g103 ( .A1(new_n223_), .A2(new_n225_), .ZN(new_n226_) );
  AND2_X1 g104 ( .A1(new_n168_), .A2(G104), .ZN(new_n227_) );
  INV_X1 g105 ( .A(G104), .ZN(new_n228_) );
  AND2_X1 g106 ( .A1(new_n228_), .A2(G143), .ZN(new_n229_) );
  OR2_X1 g107 ( .A1(new_n227_), .A2(new_n229_), .ZN(new_n230_) );
  AND2_X1 g108 ( .A1(new_n226_), .A2(new_n230_), .ZN(new_n231_) );
  INV_X1 g109 ( .A(new_n231_), .ZN(new_n232_) );
  OR2_X1 g110 ( .A1(new_n226_), .A2(new_n230_), .ZN(new_n233_) );
  AND2_X1 g111 ( .A1(new_n232_), .A2(new_n233_), .ZN(new_n234_) );
  INV_X1 g112 ( .A(G131), .ZN(new_n235_) );
  INV_X1 g113 ( .A(G146), .ZN(new_n236_) );
  AND2_X1 g114 ( .A1(new_n235_), .A2(new_n236_), .ZN(new_n237_) );
  AND2_X1 g115 ( .A1(G131), .A2(G146), .ZN(new_n238_) );
  OR2_X1 g116 ( .A1(new_n237_), .A2(new_n238_), .ZN(new_n239_) );
  AND2_X1 g117 ( .A1(new_n239_), .A2(KEYINPUT12), .ZN(new_n240_) );
  INV_X1 g118 ( .A(new_n238_), .ZN(new_n241_) );
  INV_X1 g119 ( .A(KEYINPUT12), .ZN(new_n242_) );
  INV_X1 g120 ( .A(new_n237_), .ZN(new_n243_) );
  AND2_X1 g121 ( .A1(new_n243_), .A2(new_n242_), .ZN(new_n244_) );
  AND2_X1 g122 ( .A1(new_n244_), .A2(new_n241_), .ZN(new_n245_) );
  OR2_X1 g123 ( .A1(new_n245_), .A2(new_n240_), .ZN(new_n246_) );
  INV_X1 g124 ( .A(new_n246_), .ZN(new_n247_) );
  INV_X1 g125 ( .A(G237), .ZN(new_n248_) );
  AND2_X1 g126 ( .A1(new_n248_), .A2(G214), .ZN(new_n249_) );
  AND2_X1 g127 ( .A1(new_n249_), .A2(new_n145_), .ZN(new_n250_) );
  INV_X1 g128 ( .A(new_n250_), .ZN(new_n251_) );
  AND2_X1 g129 ( .A1(new_n247_), .A2(new_n251_), .ZN(new_n252_) );
  AND2_X1 g130 ( .A1(new_n246_), .A2(new_n250_), .ZN(new_n253_) );
  OR2_X1 g131 ( .A1(new_n252_), .A2(new_n253_), .ZN(new_n254_) );
  INV_X1 g132 ( .A(new_n254_), .ZN(new_n255_) );
  OR2_X1 g133 ( .A1(new_n234_), .A2(new_n255_), .ZN(new_n256_) );
  AND2_X1 g134 ( .A1(new_n234_), .A2(new_n255_), .ZN(new_n257_) );
  INV_X1 g135 ( .A(new_n257_), .ZN(new_n258_) );
  AND2_X1 g136 ( .A1(new_n258_), .A2(new_n256_), .ZN(new_n259_) );
  OR2_X1 g137 ( .A1(new_n259_), .A2(G902), .ZN(new_n260_) );
  INV_X1 g138 ( .A(G475), .ZN(new_n261_) );
  AND2_X1 g139 ( .A1(new_n261_), .A2(KEYINPUT13), .ZN(new_n262_) );
  INV_X1 g140 ( .A(new_n262_), .ZN(new_n263_) );
  OR2_X1 g141 ( .A1(new_n261_), .A2(KEYINPUT13), .ZN(new_n264_) );
  AND2_X1 g142 ( .A1(new_n263_), .A2(new_n264_), .ZN(new_n265_) );
  AND2_X1 g143 ( .A1(new_n260_), .A2(new_n265_), .ZN(new_n266_) );
  INV_X1 g144 ( .A(new_n266_), .ZN(new_n267_) );
  OR2_X1 g145 ( .A1(new_n260_), .A2(new_n265_), .ZN(new_n268_) );
  AND2_X1 g146 ( .A1(new_n267_), .A2(new_n268_), .ZN(new_n269_) );
  INV_X1 g147 ( .A(new_n269_), .ZN(new_n270_) );
  AND2_X1 g148 ( .A1(new_n202_), .A2(new_n270_), .ZN(new_n271_) );
  AND2_X1 g149 ( .A1(new_n271_), .A2(new_n142_), .ZN(new_n272_) );
  INV_X1 g150 ( .A(G119), .ZN(new_n273_) );
  INV_X1 g151 ( .A(KEYINPUT3), .ZN(new_n274_) );
  AND2_X1 g152 ( .A1(new_n273_), .A2(new_n274_), .ZN(new_n275_) );
  AND2_X1 g153 ( .A1(G119), .A2(KEYINPUT3), .ZN(new_n276_) );
  OR2_X1 g154 ( .A1(new_n275_), .A2(new_n276_), .ZN(new_n277_) );
  AND2_X1 g155 ( .A1(new_n214_), .A2(new_n144_), .ZN(new_n278_) );
  AND2_X1 g156 ( .A1(G113), .A2(G116), .ZN(new_n279_) );
  OR2_X1 g157 ( .A1(new_n278_), .A2(new_n279_), .ZN(new_n280_) );
  AND2_X1 g158 ( .A1(new_n277_), .A2(new_n280_), .ZN(new_n281_) );
  OR2_X1 g159 ( .A1(G119), .A2(KEYINPUT3), .ZN(new_n282_) );
  INV_X1 g160 ( .A(new_n276_), .ZN(new_n283_) );
  AND2_X1 g161 ( .A1(new_n283_), .A2(new_n282_), .ZN(new_n284_) );
  OR2_X1 g162 ( .A1(G113), .A2(G116), .ZN(new_n285_) );
  INV_X1 g163 ( .A(new_n279_), .ZN(new_n286_) );
  AND2_X1 g164 ( .A1(new_n286_), .A2(new_n285_), .ZN(new_n287_) );
  AND2_X1 g165 ( .A1(new_n284_), .A2(new_n287_), .ZN(new_n288_) );
  OR2_X1 g166 ( .A1(new_n281_), .A2(new_n288_), .ZN(new_n289_) );
  AND2_X1 g167 ( .A1(G122), .A2(KEYINPUT16), .ZN(new_n290_) );
  INV_X1 g168 ( .A(new_n290_), .ZN(new_n291_) );
  OR2_X1 g169 ( .A1(G122), .A2(KEYINPUT16), .ZN(new_n292_) );
  AND2_X1 g170 ( .A1(new_n291_), .A2(new_n292_), .ZN(new_n293_) );
  AND2_X1 g171 ( .A1(new_n289_), .A2(new_n293_), .ZN(new_n294_) );
  OR2_X1 g172 ( .A1(new_n284_), .A2(new_n287_), .ZN(new_n295_) );
  OR2_X1 g173 ( .A1(new_n277_), .A2(new_n280_), .ZN(new_n296_) );
  AND2_X1 g174 ( .A1(new_n296_), .A2(new_n295_), .ZN(new_n297_) );
  INV_X1 g175 ( .A(new_n293_), .ZN(new_n298_) );
  AND2_X1 g176 ( .A1(new_n297_), .A2(new_n298_), .ZN(new_n299_) );
  OR2_X1 g177 ( .A1(new_n299_), .A2(new_n294_), .ZN(new_n300_) );
  INV_X1 g178 ( .A(KEYINPUT18), .ZN(new_n301_) );
  INV_X1 g179 ( .A(KEYINPUT17), .ZN(new_n302_) );
  AND2_X1 g180 ( .A1(new_n301_), .A2(new_n302_), .ZN(new_n303_) );
  AND2_X1 g181 ( .A1(KEYINPUT18), .A2(KEYINPUT17), .ZN(new_n304_) );
  OR2_X1 g182 ( .A1(new_n303_), .A2(new_n304_), .ZN(new_n305_) );
  AND2_X1 g183 ( .A1(new_n145_), .A2(G224), .ZN(new_n306_) );
  AND2_X1 g184 ( .A1(new_n305_), .A2(new_n306_), .ZN(new_n307_) );
  OR2_X1 g185 ( .A1(KEYINPUT18), .A2(KEYINPUT17), .ZN(new_n308_) );
  INV_X1 g186 ( .A(new_n304_), .ZN(new_n309_) );
  AND2_X1 g187 ( .A1(new_n309_), .A2(new_n308_), .ZN(new_n310_) );
  INV_X1 g188 ( .A(new_n306_), .ZN(new_n311_) );
  AND2_X1 g189 ( .A1(new_n310_), .A2(new_n311_), .ZN(new_n312_) );
  OR2_X1 g190 ( .A1(new_n307_), .A2(new_n312_), .ZN(new_n313_) );
  AND2_X1 g191 ( .A1(new_n236_), .A2(G125), .ZN(new_n314_) );
  AND2_X1 g192 ( .A1(new_n203_), .A2(G146), .ZN(new_n315_) );
  OR2_X1 g193 ( .A1(new_n314_), .A2(new_n315_), .ZN(new_n316_) );
  INV_X1 g194 ( .A(new_n316_), .ZN(new_n317_) );
  AND2_X1 g195 ( .A1(new_n313_), .A2(new_n317_), .ZN(new_n318_) );
  OR2_X1 g196 ( .A1(new_n310_), .A2(new_n311_), .ZN(new_n319_) );
  OR2_X1 g197 ( .A1(new_n305_), .A2(new_n306_), .ZN(new_n320_) );
  AND2_X1 g198 ( .A1(new_n320_), .A2(new_n319_), .ZN(new_n321_) );
  AND2_X1 g199 ( .A1(new_n321_), .A2(new_n316_), .ZN(new_n322_) );
  OR2_X1 g200 ( .A1(new_n318_), .A2(new_n322_), .ZN(new_n323_) );
  AND2_X1 g201 ( .A1(new_n300_), .A2(new_n323_), .ZN(new_n324_) );
  OR2_X1 g202 ( .A1(new_n297_), .A2(new_n298_), .ZN(new_n325_) );
  OR2_X1 g203 ( .A1(new_n289_), .A2(new_n293_), .ZN(new_n326_) );
  AND2_X1 g204 ( .A1(new_n325_), .A2(new_n326_), .ZN(new_n327_) );
  OR2_X1 g205 ( .A1(new_n321_), .A2(new_n316_), .ZN(new_n328_) );
  OR2_X1 g206 ( .A1(new_n313_), .A2(new_n317_), .ZN(new_n329_) );
  AND2_X1 g207 ( .A1(new_n329_), .A2(new_n328_), .ZN(new_n330_) );
  AND2_X1 g208 ( .A1(new_n327_), .A2(new_n330_), .ZN(new_n331_) );
  OR2_X1 g209 ( .A1(new_n324_), .A2(new_n331_), .ZN(new_n332_) );
  AND2_X1 g210 ( .A1(new_n171_), .A2(KEYINPUT4), .ZN(new_n333_) );
  INV_X1 g211 ( .A(KEYINPUT4), .ZN(new_n334_) );
  AND2_X1 g212 ( .A1(new_n173_), .A2(new_n334_), .ZN(new_n335_) );
  AND2_X1 g213 ( .A1(new_n335_), .A2(new_n174_), .ZN(new_n336_) );
  OR2_X1 g214 ( .A1(new_n333_), .A2(new_n336_), .ZN(new_n337_) );
  AND2_X1 g215 ( .A1(new_n337_), .A2(new_n123_), .ZN(new_n338_) );
  OR2_X1 g216 ( .A1(new_n175_), .A2(new_n334_), .ZN(new_n339_) );
  INV_X1 g217 ( .A(new_n336_), .ZN(new_n340_) );
  AND2_X1 g218 ( .A1(new_n340_), .A2(new_n339_), .ZN(new_n341_) );
  AND2_X1 g219 ( .A1(new_n341_), .A2(G101), .ZN(new_n342_) );
  OR2_X1 g220 ( .A1(new_n338_), .A2(new_n342_), .ZN(new_n343_) );
  AND2_X1 g221 ( .A1(G104), .A2(G110), .ZN(new_n344_) );
  INV_X1 g222 ( .A(G110), .ZN(new_n345_) );
  AND2_X1 g223 ( .A1(new_n228_), .A2(new_n345_), .ZN(new_n346_) );
  OR2_X1 g224 ( .A1(new_n346_), .A2(new_n344_), .ZN(new_n347_) );
  OR2_X1 g225 ( .A1(new_n347_), .A2(G107), .ZN(new_n348_) );
  AND2_X1 g226 ( .A1(new_n347_), .A2(G107), .ZN(new_n349_) );
  INV_X1 g227 ( .A(new_n349_), .ZN(new_n350_) );
  AND2_X1 g228 ( .A1(new_n350_), .A2(new_n348_), .ZN(new_n351_) );
  AND2_X1 g229 ( .A1(new_n343_), .A2(new_n351_), .ZN(new_n352_) );
  OR2_X1 g230 ( .A1(new_n341_), .A2(G101), .ZN(new_n353_) );
  OR2_X1 g231 ( .A1(new_n337_), .A2(new_n123_), .ZN(new_n354_) );
  AND2_X1 g232 ( .A1(new_n354_), .A2(new_n353_), .ZN(new_n355_) );
  INV_X1 g233 ( .A(new_n351_), .ZN(new_n356_) );
  AND2_X1 g234 ( .A1(new_n355_), .A2(new_n356_), .ZN(new_n357_) );
  OR2_X1 g235 ( .A1(new_n352_), .A2(new_n357_), .ZN(new_n358_) );
  AND2_X1 g236 ( .A1(new_n332_), .A2(new_n358_), .ZN(new_n359_) );
  OR2_X1 g237 ( .A1(new_n327_), .A2(new_n330_), .ZN(new_n360_) );
  OR2_X1 g238 ( .A1(new_n300_), .A2(new_n323_), .ZN(new_n361_) );
  AND2_X1 g239 ( .A1(new_n361_), .A2(new_n360_), .ZN(new_n362_) );
  OR2_X1 g240 ( .A1(new_n355_), .A2(new_n356_), .ZN(new_n363_) );
  OR2_X1 g241 ( .A1(new_n343_), .A2(new_n351_), .ZN(new_n364_) );
  AND2_X1 g242 ( .A1(new_n364_), .A2(new_n363_), .ZN(new_n365_) );
  AND2_X1 g243 ( .A1(new_n362_), .A2(new_n365_), .ZN(new_n366_) );
  OR2_X1 g244 ( .A1(new_n359_), .A2(new_n366_), .ZN(new_n367_) );
  OR2_X1 g245 ( .A1(new_n367_), .A2(new_n130_), .ZN(new_n368_) );
  AND2_X1 g246 ( .A1(new_n248_), .A2(new_n195_), .ZN(new_n369_) );
  INV_X1 g247 ( .A(new_n369_), .ZN(new_n370_) );
  AND2_X1 g248 ( .A1(new_n370_), .A2(G210), .ZN(new_n371_) );
  AND2_X1 g249 ( .A1(new_n368_), .A2(new_n371_), .ZN(new_n372_) );
  OR2_X1 g250 ( .A1(new_n362_), .A2(new_n365_), .ZN(new_n373_) );
  OR2_X1 g251 ( .A1(new_n332_), .A2(new_n358_), .ZN(new_n374_) );
  AND2_X1 g252 ( .A1(new_n374_), .A2(new_n373_), .ZN(new_n375_) );
  AND2_X1 g253 ( .A1(new_n375_), .A2(new_n131_), .ZN(new_n376_) );
  INV_X1 g254 ( .A(new_n371_), .ZN(new_n377_) );
  AND2_X1 g255 ( .A1(new_n376_), .A2(new_n377_), .ZN(new_n378_) );
  OR2_X1 g256 ( .A1(new_n372_), .A2(new_n378_), .ZN(new_n379_) );
  AND2_X1 g257 ( .A1(new_n370_), .A2(G214), .ZN(new_n380_) );
  INV_X1 g258 ( .A(new_n380_), .ZN(new_n381_) );
  AND2_X1 g259 ( .A1(new_n379_), .A2(new_n381_), .ZN(new_n382_) );
  AND2_X1 g260 ( .A1(new_n382_), .A2(KEYINPUT19), .ZN(new_n383_) );
  AND2_X1 g261 ( .A1(new_n383_), .A2(KEYINPUT0), .ZN(new_n384_) );
  INV_X1 g262 ( .A(new_n384_), .ZN(new_n385_) );
  INV_X1 g263 ( .A(KEYINPUT0), .ZN(new_n386_) );
  INV_X1 g264 ( .A(KEYINPUT14), .ZN(new_n387_) );
  AND2_X1 g265 ( .A1(G234), .A2(G237), .ZN(new_n388_) );
  OR2_X1 g266 ( .A1(new_n388_), .A2(new_n387_), .ZN(new_n389_) );
  AND2_X1 g267 ( .A1(new_n388_), .A2(new_n387_), .ZN(new_n390_) );
  INV_X1 g268 ( .A(new_n390_), .ZN(new_n391_) );
  AND2_X1 g269 ( .A1(new_n391_), .A2(new_n389_), .ZN(new_n392_) );
  INV_X1 g270 ( .A(new_n392_), .ZN(new_n393_) );
  AND2_X1 g271 ( .A1(new_n393_), .A2(G952), .ZN(new_n394_) );
  AND2_X1 g272 ( .A1(new_n394_), .A2(new_n145_), .ZN(new_n395_) );
  AND2_X1 g273 ( .A1(new_n393_), .A2(G902), .ZN(new_n396_) );
  INV_X1 g274 ( .A(G898), .ZN(new_n397_) );
  AND2_X1 g275 ( .A1(new_n397_), .A2(G953), .ZN(new_n398_) );
  AND2_X1 g276 ( .A1(new_n396_), .A2(new_n398_), .ZN(new_n399_) );
  OR2_X1 g277 ( .A1(new_n395_), .A2(new_n399_), .ZN(new_n400_) );
  INV_X1 g278 ( .A(KEYINPUT19), .ZN(new_n401_) );
  OR2_X1 g279 ( .A1(new_n376_), .A2(new_n377_), .ZN(new_n402_) );
  OR2_X1 g280 ( .A1(new_n368_), .A2(new_n371_), .ZN(new_n403_) );
  AND2_X1 g281 ( .A1(new_n403_), .A2(new_n402_), .ZN(new_n404_) );
  OR2_X1 g282 ( .A1(new_n404_), .A2(new_n380_), .ZN(new_n405_) );
  OR2_X1 g283 ( .A1(new_n405_), .A2(new_n401_), .ZN(new_n406_) );
  OR2_X1 g284 ( .A1(new_n382_), .A2(KEYINPUT19), .ZN(new_n407_) );
  AND2_X1 g285 ( .A1(new_n406_), .A2(new_n407_), .ZN(new_n408_) );
  AND2_X1 g286 ( .A1(new_n408_), .A2(new_n400_), .ZN(new_n409_) );
  OR2_X1 g287 ( .A1(new_n409_), .A2(new_n386_), .ZN(new_n410_) );
  INV_X1 g288 ( .A(new_n400_), .ZN(new_n411_) );
  AND2_X1 g289 ( .A1(new_n405_), .A2(new_n401_), .ZN(new_n412_) );
  OR2_X1 g290 ( .A1(new_n412_), .A2(new_n383_), .ZN(new_n413_) );
  OR2_X1 g291 ( .A1(new_n413_), .A2(new_n411_), .ZN(new_n414_) );
  OR2_X1 g292 ( .A1(new_n414_), .A2(KEYINPUT0), .ZN(new_n415_) );
  AND2_X1 g293 ( .A1(new_n415_), .A2(new_n410_), .ZN(new_n416_) );
  AND2_X1 g294 ( .A1(new_n416_), .A2(new_n385_), .ZN(new_n417_) );
  AND2_X1 g295 ( .A1(new_n417_), .A2(new_n272_), .ZN(new_n418_) );
  AND2_X1 g296 ( .A1(new_n418_), .A2(new_n124_), .ZN(new_n419_) );
  INV_X1 g297 ( .A(new_n419_), .ZN(new_n420_) );
  OR2_X1 g298 ( .A1(new_n418_), .A2(new_n124_), .ZN(new_n421_) );
  INV_X1 g299 ( .A(G469), .ZN(new_n422_) );
  AND2_X1 g300 ( .A1(new_n145_), .A2(G227), .ZN(new_n423_) );
  INV_X1 g301 ( .A(new_n423_), .ZN(new_n424_) );
  INV_X1 g302 ( .A(G137), .ZN(new_n425_) );
  AND2_X1 g303 ( .A1(new_n425_), .A2(new_n208_), .ZN(new_n426_) );
  AND2_X1 g304 ( .A1(G137), .A2(G140), .ZN(new_n427_) );
  OR2_X1 g305 ( .A1(new_n426_), .A2(new_n427_), .ZN(new_n428_) );
  AND2_X1 g306 ( .A1(new_n239_), .A2(G134), .ZN(new_n429_) );
  INV_X1 g307 ( .A(new_n429_), .ZN(new_n430_) );
  OR2_X1 g308 ( .A1(new_n239_), .A2(G134), .ZN(new_n431_) );
  AND2_X1 g309 ( .A1(new_n430_), .A2(new_n431_), .ZN(new_n432_) );
  AND2_X1 g310 ( .A1(new_n432_), .A2(new_n428_), .ZN(new_n433_) );
  INV_X1 g311 ( .A(new_n428_), .ZN(new_n434_) );
  INV_X1 g312 ( .A(new_n432_), .ZN(new_n435_) );
  AND2_X1 g313 ( .A1(new_n435_), .A2(new_n434_), .ZN(new_n436_) );
  OR2_X1 g314 ( .A1(new_n436_), .A2(new_n433_), .ZN(new_n437_) );
  INV_X1 g315 ( .A(new_n437_), .ZN(new_n438_) );
  AND2_X1 g316 ( .A1(new_n438_), .A2(new_n424_), .ZN(new_n439_) );
  AND2_X1 g317 ( .A1(new_n437_), .A2(new_n423_), .ZN(new_n440_) );
  OR2_X1 g318 ( .A1(new_n439_), .A2(new_n440_), .ZN(new_n441_) );
  INV_X1 g319 ( .A(new_n441_), .ZN(new_n442_) );
  AND2_X1 g320 ( .A1(new_n442_), .A2(new_n358_), .ZN(new_n443_) );
  AND2_X1 g321 ( .A1(new_n441_), .A2(new_n365_), .ZN(new_n444_) );
  OR2_X1 g322 ( .A1(new_n443_), .A2(new_n444_), .ZN(new_n445_) );
  OR2_X1 g323 ( .A1(new_n445_), .A2(G902), .ZN(new_n446_) );
  AND2_X1 g324 ( .A1(new_n446_), .A2(new_n422_), .ZN(new_n447_) );
  OR2_X1 g325 ( .A1(new_n446_), .A2(new_n422_), .ZN(new_n448_) );
  INV_X1 g326 ( .A(new_n448_), .ZN(new_n449_) );
  OR2_X1 g327 ( .A1(new_n449_), .A2(new_n447_), .ZN(new_n450_) );
  AND2_X1 g328 ( .A1(new_n450_), .A2(KEYINPUT1), .ZN(new_n451_) );
  INV_X1 g329 ( .A(KEYINPUT1), .ZN(new_n452_) );
  INV_X1 g330 ( .A(new_n447_), .ZN(new_n453_) );
  AND2_X1 g331 ( .A1(new_n453_), .A2(new_n448_), .ZN(new_n454_) );
  AND2_X1 g332 ( .A1(new_n454_), .A2(new_n452_), .ZN(new_n455_) );
  OR2_X1 g333 ( .A1(new_n451_), .A2(new_n455_), .ZN(new_n456_) );
  AND2_X1 g334 ( .A1(new_n421_), .A2(new_n456_), .ZN(new_n457_) );
  AND2_X1 g335 ( .A1(new_n457_), .A2(new_n420_), .ZN(new_n458_) );
  INV_X1 g336 ( .A(KEYINPUT25), .ZN(new_n459_) );
  AND2_X1 g337 ( .A1(new_n207_), .A2(new_n428_), .ZN(new_n460_) );
  AND2_X1 g338 ( .A1(new_n224_), .A2(new_n434_), .ZN(new_n461_) );
  OR2_X1 g339 ( .A1(new_n461_), .A2(new_n460_), .ZN(new_n462_) );
  AND2_X1 g340 ( .A1(new_n273_), .A2(new_n236_), .ZN(new_n463_) );
  AND2_X1 g341 ( .A1(G119), .A2(G146), .ZN(new_n464_) );
  OR2_X1 g342 ( .A1(new_n463_), .A2(new_n464_), .ZN(new_n465_) );
  AND2_X1 g343 ( .A1(new_n345_), .A2(new_n167_), .ZN(new_n466_) );
  AND2_X1 g344 ( .A1(G110), .A2(G128), .ZN(new_n467_) );
  OR2_X1 g345 ( .A1(new_n466_), .A2(new_n467_), .ZN(new_n468_) );
  AND2_X1 g346 ( .A1(new_n465_), .A2(new_n468_), .ZN(new_n469_) );
  INV_X1 g347 ( .A(new_n469_), .ZN(new_n470_) );
  OR2_X1 g348 ( .A1(new_n465_), .A2(new_n468_), .ZN(new_n471_) );
  AND2_X1 g349 ( .A1(new_n470_), .A2(new_n471_), .ZN(new_n472_) );
  INV_X1 g350 ( .A(new_n472_), .ZN(new_n473_) );
  AND2_X1 g351 ( .A1(new_n473_), .A2(new_n462_), .ZN(new_n474_) );
  INV_X1 g352 ( .A(new_n474_), .ZN(new_n475_) );
  OR2_X1 g353 ( .A1(new_n473_), .A2(new_n462_), .ZN(new_n476_) );
  AND2_X1 g354 ( .A1(new_n475_), .A2(new_n476_), .ZN(new_n477_) );
  AND2_X1 g355 ( .A1(new_n151_), .A2(G221), .ZN(new_n478_) );
  INV_X1 g356 ( .A(new_n478_), .ZN(new_n479_) );
  INV_X1 g357 ( .A(KEYINPUT24), .ZN(new_n480_) );
  AND2_X1 g358 ( .A1(new_n480_), .A2(KEYINPUT23), .ZN(new_n481_) );
  INV_X1 g359 ( .A(new_n481_), .ZN(new_n482_) );
  OR2_X1 g360 ( .A1(new_n480_), .A2(KEYINPUT23), .ZN(new_n483_) );
  AND2_X1 g361 ( .A1(new_n482_), .A2(new_n483_), .ZN(new_n484_) );
  INV_X1 g362 ( .A(new_n484_), .ZN(new_n485_) );
  AND2_X1 g363 ( .A1(new_n479_), .A2(new_n485_), .ZN(new_n486_) );
  AND2_X1 g364 ( .A1(new_n478_), .A2(new_n484_), .ZN(new_n487_) );
  OR2_X1 g365 ( .A1(new_n486_), .A2(new_n487_), .ZN(new_n488_) );
  OR2_X1 g366 ( .A1(new_n477_), .A2(new_n488_), .ZN(new_n489_) );
  AND2_X1 g367 ( .A1(new_n477_), .A2(new_n488_), .ZN(new_n490_) );
  INV_X1 g368 ( .A(new_n490_), .ZN(new_n491_) );
  AND2_X1 g369 ( .A1(new_n491_), .A2(new_n489_), .ZN(new_n492_) );
  OR2_X1 g370 ( .A1(new_n492_), .A2(G902), .ZN(new_n493_) );
  AND2_X1 g371 ( .A1(new_n137_), .A2(G217), .ZN(new_n494_) );
  AND2_X1 g372 ( .A1(new_n493_), .A2(new_n494_), .ZN(new_n495_) );
  INV_X1 g373 ( .A(new_n492_), .ZN(new_n496_) );
  AND2_X1 g374 ( .A1(new_n496_), .A2(new_n195_), .ZN(new_n497_) );
  INV_X1 g375 ( .A(new_n494_), .ZN(new_n498_) );
  AND2_X1 g376 ( .A1(new_n497_), .A2(new_n498_), .ZN(new_n499_) );
  OR2_X1 g377 ( .A1(new_n499_), .A2(new_n495_), .ZN(new_n500_) );
  AND2_X1 g378 ( .A1(new_n500_), .A2(new_n459_), .ZN(new_n501_) );
  INV_X1 g379 ( .A(new_n495_), .ZN(new_n502_) );
  OR2_X1 g380 ( .A1(new_n493_), .A2(new_n494_), .ZN(new_n503_) );
  AND2_X1 g381 ( .A1(new_n502_), .A2(new_n503_), .ZN(new_n504_) );
  AND2_X1 g382 ( .A1(new_n504_), .A2(KEYINPUT25), .ZN(new_n505_) );
  OR2_X1 g383 ( .A1(new_n501_), .A2(new_n505_), .ZN(new_n506_) );
  INV_X1 g384 ( .A(new_n506_), .ZN(new_n507_) );
  INV_X1 g385 ( .A(KEYINPUT6), .ZN(new_n508_) );
  OR2_X1 g386 ( .A1(G137), .A2(KEYINPUT5), .ZN(new_n509_) );
  AND2_X1 g387 ( .A1(G137), .A2(KEYINPUT5), .ZN(new_n510_) );
  INV_X1 g388 ( .A(new_n510_), .ZN(new_n511_) );
  AND2_X1 g389 ( .A1(new_n511_), .A2(new_n509_), .ZN(new_n512_) );
  INV_X1 g390 ( .A(new_n512_), .ZN(new_n513_) );
  AND2_X1 g391 ( .A1(new_n248_), .A2(G210), .ZN(new_n514_) );
  AND2_X1 g392 ( .A1(new_n514_), .A2(new_n145_), .ZN(new_n515_) );
  INV_X1 g393 ( .A(new_n515_), .ZN(new_n516_) );
  AND2_X1 g394 ( .A1(new_n513_), .A2(new_n516_), .ZN(new_n517_) );
  AND2_X1 g395 ( .A1(new_n512_), .A2(new_n515_), .ZN(new_n518_) );
  OR2_X1 g396 ( .A1(new_n517_), .A2(new_n518_), .ZN(new_n519_) );
  AND2_X1 g397 ( .A1(new_n519_), .A2(new_n289_), .ZN(new_n520_) );
  INV_X1 g398 ( .A(new_n520_), .ZN(new_n521_) );
  OR2_X1 g399 ( .A1(new_n519_), .A2(new_n289_), .ZN(new_n522_) );
  AND2_X1 g400 ( .A1(new_n521_), .A2(new_n522_), .ZN(new_n523_) );
  OR2_X1 g401 ( .A1(new_n523_), .A2(new_n435_), .ZN(new_n524_) );
  AND2_X1 g402 ( .A1(new_n523_), .A2(new_n435_), .ZN(new_n525_) );
  INV_X1 g403 ( .A(new_n525_), .ZN(new_n526_) );
  AND2_X1 g404 ( .A1(new_n526_), .A2(new_n524_), .ZN(new_n527_) );
  OR2_X1 g405 ( .A1(new_n527_), .A2(new_n355_), .ZN(new_n528_) );
  INV_X1 g406 ( .A(new_n523_), .ZN(new_n529_) );
  AND2_X1 g407 ( .A1(new_n529_), .A2(new_n432_), .ZN(new_n530_) );
  OR2_X1 g408 ( .A1(new_n530_), .A2(new_n525_), .ZN(new_n531_) );
  OR2_X1 g409 ( .A1(new_n531_), .A2(new_n343_), .ZN(new_n532_) );
  AND2_X1 g410 ( .A1(new_n532_), .A2(new_n528_), .ZN(new_n533_) );
  AND2_X1 g411 ( .A1(new_n533_), .A2(new_n195_), .ZN(new_n534_) );
  OR2_X1 g412 ( .A1(new_n534_), .A2(G472), .ZN(new_n535_) );
  INV_X1 g413 ( .A(G472), .ZN(new_n536_) );
  AND2_X1 g414 ( .A1(new_n531_), .A2(new_n343_), .ZN(new_n537_) );
  AND2_X1 g415 ( .A1(new_n527_), .A2(new_n355_), .ZN(new_n538_) );
  OR2_X1 g416 ( .A1(new_n537_), .A2(new_n538_), .ZN(new_n539_) );
  OR2_X1 g417 ( .A1(new_n539_), .A2(G902), .ZN(new_n540_) );
  OR2_X1 g418 ( .A1(new_n540_), .A2(new_n536_), .ZN(new_n541_) );
  AND2_X1 g419 ( .A1(new_n541_), .A2(new_n535_), .ZN(new_n542_) );
  OR2_X1 g420 ( .A1(new_n542_), .A2(new_n508_), .ZN(new_n543_) );
  AND2_X1 g421 ( .A1(new_n540_), .A2(new_n536_), .ZN(new_n544_) );
  AND2_X1 g422 ( .A1(new_n534_), .A2(G472), .ZN(new_n545_) );
  OR2_X1 g423 ( .A1(new_n544_), .A2(new_n545_), .ZN(new_n546_) );
  OR2_X1 g424 ( .A1(new_n546_), .A2(KEYINPUT6), .ZN(new_n547_) );
  AND2_X1 g425 ( .A1(new_n543_), .A2(new_n547_), .ZN(new_n548_) );
  AND2_X1 g426 ( .A1(new_n548_), .A2(new_n507_), .ZN(new_n549_) );
  AND2_X1 g427 ( .A1(new_n458_), .A2(new_n549_), .ZN(new_n550_) );
  AND2_X1 g428 ( .A1(new_n550_), .A2(new_n123_), .ZN(new_n551_) );
  INV_X1 g429 ( .A(new_n550_), .ZN(new_n552_) );
  AND2_X1 g430 ( .A1(new_n552_), .A2(G101), .ZN(new_n553_) );
  OR2_X1 g431 ( .A1(new_n553_), .A2(new_n551_), .ZN(G3) );
  INV_X1 g432 ( .A(new_n142_), .ZN(new_n555_) );
  OR2_X1 g433 ( .A1(new_n506_), .A2(new_n555_), .ZN(new_n556_) );
  OR2_X1 g434 ( .A1(new_n556_), .A2(new_n450_), .ZN(new_n557_) );
  INV_X1 g435 ( .A(new_n557_), .ZN(new_n558_) );
  AND2_X1 g436 ( .A1(new_n558_), .A2(new_n546_), .ZN(new_n559_) );
  AND2_X1 g437 ( .A1(new_n417_), .A2(new_n559_), .ZN(new_n560_) );
  AND2_X1 g438 ( .A1(new_n202_), .A2(new_n269_), .ZN(new_n561_) );
  AND2_X1 g439 ( .A1(new_n560_), .A2(new_n561_), .ZN(new_n562_) );
  INV_X1 g440 ( .A(new_n562_), .ZN(new_n563_) );
  AND2_X1 g441 ( .A1(new_n563_), .A2(G104), .ZN(new_n564_) );
  AND2_X1 g442 ( .A1(new_n562_), .A2(new_n228_), .ZN(new_n565_) );
  OR2_X1 g443 ( .A1(new_n564_), .A2(new_n565_), .ZN(G6) );
  OR2_X1 g444 ( .A1(new_n200_), .A2(G478), .ZN(new_n567_) );
  OR2_X1 g445 ( .A1(new_n193_), .A2(new_n143_), .ZN(new_n568_) );
  AND2_X1 g446 ( .A1(new_n568_), .A2(new_n567_), .ZN(new_n569_) );
  AND2_X1 g447 ( .A1(new_n569_), .A2(new_n270_), .ZN(new_n570_) );
  AND2_X1 g448 ( .A1(new_n560_), .A2(new_n570_), .ZN(new_n571_) );
  INV_X1 g449 ( .A(new_n571_), .ZN(new_n572_) );
  INV_X1 g450 ( .A(KEYINPUT26), .ZN(new_n573_) );
  AND2_X1 g451 ( .A1(new_n573_), .A2(KEYINPUT27), .ZN(new_n574_) );
  INV_X1 g452 ( .A(new_n574_), .ZN(new_n575_) );
  OR2_X1 g453 ( .A1(new_n573_), .A2(KEYINPUT27), .ZN(new_n576_) );
  AND2_X1 g454 ( .A1(new_n575_), .A2(new_n576_), .ZN(new_n577_) );
  INV_X1 g455 ( .A(new_n577_), .ZN(new_n578_) );
  AND2_X1 g456 ( .A1(new_n572_), .A2(new_n578_), .ZN(new_n579_) );
  AND2_X1 g457 ( .A1(new_n571_), .A2(new_n577_), .ZN(new_n580_) );
  OR2_X1 g458 ( .A1(new_n579_), .A2(new_n580_), .ZN(new_n581_) );
  AND2_X1 g459 ( .A1(new_n581_), .A2(G107), .ZN(new_n582_) );
  INV_X1 g460 ( .A(new_n581_), .ZN(new_n583_) );
  AND2_X1 g461 ( .A1(new_n583_), .A2(new_n166_), .ZN(new_n584_) );
  OR2_X1 g462 ( .A1(new_n584_), .A2(new_n582_), .ZN(G9) );
  AND2_X1 g463 ( .A1(new_n506_), .A2(new_n546_), .ZN(new_n586_) );
  AND2_X1 g464 ( .A1(new_n458_), .A2(new_n586_), .ZN(new_n587_) );
  INV_X1 g465 ( .A(new_n587_), .ZN(new_n588_) );
  AND2_X1 g466 ( .A1(new_n588_), .A2(G110), .ZN(new_n589_) );
  AND2_X1 g467 ( .A1(new_n587_), .A2(new_n345_), .ZN(new_n590_) );
  OR2_X1 g468 ( .A1(new_n589_), .A2(new_n590_), .ZN(G12) );
  INV_X1 g469 ( .A(KEYINPUT28), .ZN(new_n592_) );
  INV_X1 g470 ( .A(G900), .ZN(new_n593_) );
  AND2_X1 g471 ( .A1(new_n593_), .A2(G953), .ZN(new_n594_) );
  AND2_X1 g472 ( .A1(new_n396_), .A2(new_n594_), .ZN(new_n595_) );
  OR2_X1 g473 ( .A1(new_n395_), .A2(new_n595_), .ZN(new_n596_) );
  AND2_X1 g474 ( .A1(new_n142_), .A2(new_n596_), .ZN(new_n597_) );
  AND2_X1 g475 ( .A1(new_n506_), .A2(new_n597_), .ZN(new_n598_) );
  AND2_X1 g476 ( .A1(new_n598_), .A2(new_n542_), .ZN(new_n599_) );
  AND2_X1 g477 ( .A1(new_n599_), .A2(new_n592_), .ZN(new_n600_) );
  INV_X1 g478 ( .A(new_n600_), .ZN(new_n601_) );
  OR2_X1 g479 ( .A1(new_n599_), .A2(new_n592_), .ZN(new_n602_) );
  AND2_X1 g480 ( .A1(new_n602_), .A2(new_n454_), .ZN(new_n603_) );
  AND2_X1 g481 ( .A1(new_n603_), .A2(new_n601_), .ZN(new_n604_) );
  AND2_X1 g482 ( .A1(new_n604_), .A2(new_n408_), .ZN(new_n605_) );
  AND2_X1 g483 ( .A1(new_n605_), .A2(new_n570_), .ZN(new_n606_) );
  INV_X1 g484 ( .A(new_n606_), .ZN(new_n607_) );
  AND2_X1 g485 ( .A1(new_n167_), .A2(KEYINPUT29), .ZN(new_n608_) );
  INV_X1 g486 ( .A(new_n608_), .ZN(new_n609_) );
  OR2_X1 g487 ( .A1(new_n167_), .A2(KEYINPUT29), .ZN(new_n610_) );
  AND2_X1 g488 ( .A1(new_n609_), .A2(new_n610_), .ZN(new_n611_) );
  INV_X1 g489 ( .A(new_n611_), .ZN(new_n612_) );
  AND2_X1 g490 ( .A1(new_n607_), .A2(new_n612_), .ZN(new_n613_) );
  AND2_X1 g491 ( .A1(new_n606_), .A2(new_n611_), .ZN(new_n614_) );
  OR2_X1 g492 ( .A1(new_n613_), .A2(new_n614_), .ZN(G30) );
  AND2_X1 g493 ( .A1(new_n542_), .A2(new_n381_), .ZN(new_n616_) );
  OR2_X1 g494 ( .A1(new_n616_), .A2(KEYINPUT30), .ZN(new_n617_) );
  AND2_X1 g495 ( .A1(new_n616_), .A2(KEYINPUT30), .ZN(new_n618_) );
  INV_X1 g496 ( .A(new_n618_), .ZN(new_n619_) );
  AND2_X1 g497 ( .A1(new_n619_), .A2(new_n617_), .ZN(new_n620_) );
  INV_X1 g498 ( .A(new_n620_), .ZN(new_n621_) );
  AND2_X1 g499 ( .A1(new_n558_), .A2(new_n596_), .ZN(new_n622_) );
  AND2_X1 g500 ( .A1(new_n622_), .A2(new_n621_), .ZN(new_n623_) );
  AND2_X1 g501 ( .A1(new_n569_), .A2(new_n269_), .ZN(new_n624_) );
  AND2_X1 g502 ( .A1(new_n624_), .A2(new_n379_), .ZN(new_n625_) );
  AND2_X1 g503 ( .A1(new_n623_), .A2(new_n625_), .ZN(new_n626_) );
  AND2_X1 g504 ( .A1(new_n626_), .A2(new_n168_), .ZN(new_n627_) );
  INV_X1 g505 ( .A(new_n626_), .ZN(new_n628_) );
  AND2_X1 g506 ( .A1(new_n628_), .A2(G143), .ZN(new_n629_) );
  OR2_X1 g507 ( .A1(new_n629_), .A2(new_n627_), .ZN(G45) );
  AND2_X1 g508 ( .A1(new_n605_), .A2(new_n561_), .ZN(new_n631_) );
  INV_X1 g509 ( .A(new_n631_), .ZN(new_n632_) );
  AND2_X1 g510 ( .A1(new_n632_), .A2(G146), .ZN(new_n633_) );
  AND2_X1 g511 ( .A1(new_n631_), .A2(new_n236_), .ZN(new_n634_) );
  OR2_X1 g512 ( .A1(new_n633_), .A2(new_n634_), .ZN(G48) );
  OR2_X1 g513 ( .A1(new_n454_), .A2(new_n452_), .ZN(new_n636_) );
  OR2_X1 g514 ( .A1(new_n450_), .A2(KEYINPUT1), .ZN(new_n637_) );
  AND2_X1 g515 ( .A1(new_n637_), .A2(new_n636_), .ZN(new_n638_) );
  AND2_X1 g516 ( .A1(new_n507_), .A2(new_n142_), .ZN(new_n639_) );
  AND2_X1 g517 ( .A1(new_n639_), .A2(new_n542_), .ZN(new_n640_) );
  AND2_X1 g518 ( .A1(new_n640_), .A2(new_n638_), .ZN(new_n641_) );
  AND2_X1 g519 ( .A1(new_n417_), .A2(new_n641_), .ZN(new_n642_) );
  INV_X1 g520 ( .A(new_n642_), .ZN(new_n643_) );
  AND2_X1 g521 ( .A1(new_n643_), .A2(KEYINPUT31), .ZN(new_n644_) );
  INV_X1 g522 ( .A(KEYINPUT31), .ZN(new_n645_) );
  AND2_X1 g523 ( .A1(new_n642_), .A2(new_n645_), .ZN(new_n646_) );
  OR2_X1 g524 ( .A1(new_n644_), .A2(new_n646_), .ZN(new_n647_) );
  AND2_X1 g525 ( .A1(new_n647_), .A2(new_n561_), .ZN(new_n648_) );
  INV_X1 g526 ( .A(new_n648_), .ZN(new_n649_) );
  AND2_X1 g527 ( .A1(new_n649_), .A2(G113), .ZN(new_n650_) );
  AND2_X1 g528 ( .A1(new_n648_), .A2(new_n214_), .ZN(new_n651_) );
  OR2_X1 g529 ( .A1(new_n650_), .A2(new_n651_), .ZN(G15) );
  AND2_X1 g530 ( .A1(new_n647_), .A2(new_n570_), .ZN(new_n653_) );
  INV_X1 g531 ( .A(new_n653_), .ZN(new_n654_) );
  AND2_X1 g532 ( .A1(new_n654_), .A2(G116), .ZN(new_n655_) );
  AND2_X1 g533 ( .A1(new_n653_), .A2(new_n144_), .ZN(new_n656_) );
  OR2_X1 g534 ( .A1(new_n655_), .A2(new_n656_), .ZN(G18) );
  OR2_X1 g535 ( .A1(new_n569_), .A2(new_n269_), .ZN(new_n658_) );
  OR2_X1 g536 ( .A1(new_n658_), .A2(new_n555_), .ZN(new_n659_) );
  AND2_X1 g537 ( .A1(new_n414_), .A2(KEYINPUT0), .ZN(new_n660_) );
  AND2_X1 g538 ( .A1(new_n409_), .A2(new_n386_), .ZN(new_n661_) );
  OR2_X1 g539 ( .A1(new_n660_), .A2(new_n661_), .ZN(new_n662_) );
  OR2_X1 g540 ( .A1(new_n662_), .A2(new_n384_), .ZN(new_n663_) );
  OR2_X1 g541 ( .A1(new_n663_), .A2(new_n659_), .ZN(new_n664_) );
  AND2_X1 g542 ( .A1(new_n664_), .A2(KEYINPUT22), .ZN(new_n665_) );
  AND2_X1 g543 ( .A1(new_n272_), .A2(new_n124_), .ZN(new_n666_) );
  AND2_X1 g544 ( .A1(new_n666_), .A2(new_n416_), .ZN(new_n667_) );
  AND2_X1 g545 ( .A1(new_n548_), .A2(new_n506_), .ZN(new_n668_) );
  AND2_X1 g546 ( .A1(new_n638_), .A2(new_n668_), .ZN(new_n669_) );
  INV_X1 g547 ( .A(new_n669_), .ZN(new_n670_) );
  OR2_X1 g548 ( .A1(new_n667_), .A2(new_n670_), .ZN(new_n671_) );
  OR2_X1 g549 ( .A1(new_n665_), .A2(new_n671_), .ZN(new_n672_) );
  AND2_X1 g550 ( .A1(new_n672_), .A2(KEYINPUT32), .ZN(new_n673_) );
  INV_X1 g551 ( .A(KEYINPUT32), .ZN(new_n674_) );
  INV_X1 g552 ( .A(new_n671_), .ZN(new_n675_) );
  AND2_X1 g553 ( .A1(new_n675_), .A2(new_n421_), .ZN(new_n676_) );
  AND2_X1 g554 ( .A1(new_n676_), .A2(new_n674_), .ZN(new_n677_) );
  OR2_X1 g555 ( .A1(new_n673_), .A2(new_n677_), .ZN(new_n678_) );
  AND2_X1 g556 ( .A1(new_n678_), .A2(G119), .ZN(new_n679_) );
  OR2_X1 g557 ( .A1(new_n676_), .A2(new_n674_), .ZN(new_n680_) );
  OR2_X1 g558 ( .A1(new_n672_), .A2(KEYINPUT32), .ZN(new_n681_) );
  AND2_X1 g559 ( .A1(new_n681_), .A2(new_n680_), .ZN(new_n682_) );
  AND2_X1 g560 ( .A1(new_n682_), .A2(new_n273_), .ZN(new_n683_) );
  OR2_X1 g561 ( .A1(new_n679_), .A2(new_n683_), .ZN(G21) );
  INV_X1 g562 ( .A(KEYINPUT35), .ZN(new_n685_) );
  INV_X1 g563 ( .A(new_n624_), .ZN(new_n686_) );
  OR2_X1 g564 ( .A1(new_n548_), .A2(new_n556_), .ZN(new_n687_) );
  OR2_X1 g565 ( .A1(new_n456_), .A2(new_n687_), .ZN(new_n688_) );
  AND2_X1 g566 ( .A1(new_n688_), .A2(KEYINPUT33), .ZN(new_n689_) );
  INV_X1 g567 ( .A(KEYINPUT33), .ZN(new_n690_) );
  AND2_X1 g568 ( .A1(new_n546_), .A2(KEYINPUT6), .ZN(new_n691_) );
  AND2_X1 g569 ( .A1(new_n542_), .A2(new_n508_), .ZN(new_n692_) );
  OR2_X1 g570 ( .A1(new_n691_), .A2(new_n692_), .ZN(new_n693_) );
  AND2_X1 g571 ( .A1(new_n639_), .A2(new_n693_), .ZN(new_n694_) );
  AND2_X1 g572 ( .A1(new_n694_), .A2(new_n638_), .ZN(new_n695_) );
  AND2_X1 g573 ( .A1(new_n695_), .A2(new_n690_), .ZN(new_n696_) );
  OR2_X1 g574 ( .A1(new_n689_), .A2(new_n696_), .ZN(new_n697_) );
  AND2_X1 g575 ( .A1(new_n697_), .A2(new_n417_), .ZN(new_n698_) );
  OR2_X1 g576 ( .A1(new_n698_), .A2(KEYINPUT34), .ZN(new_n699_) );
  INV_X1 g577 ( .A(KEYINPUT34), .ZN(new_n700_) );
  OR2_X1 g578 ( .A1(new_n695_), .A2(new_n690_), .ZN(new_n701_) );
  OR2_X1 g579 ( .A1(new_n688_), .A2(KEYINPUT33), .ZN(new_n702_) );
  AND2_X1 g580 ( .A1(new_n702_), .A2(new_n701_), .ZN(new_n703_) );
  OR2_X1 g581 ( .A1(new_n663_), .A2(new_n703_), .ZN(new_n704_) );
  OR2_X1 g582 ( .A1(new_n704_), .A2(new_n700_), .ZN(new_n705_) );
  AND2_X1 g583 ( .A1(new_n705_), .A2(new_n699_), .ZN(new_n706_) );
  OR2_X1 g584 ( .A1(new_n706_), .A2(new_n686_), .ZN(new_n707_) );
  AND2_X1 g585 ( .A1(new_n707_), .A2(new_n685_), .ZN(new_n708_) );
  AND2_X1 g586 ( .A1(new_n704_), .A2(new_n700_), .ZN(new_n709_) );
  AND2_X1 g587 ( .A1(new_n698_), .A2(KEYINPUT34), .ZN(new_n710_) );
  OR2_X1 g588 ( .A1(new_n709_), .A2(new_n710_), .ZN(new_n711_) );
  AND2_X1 g589 ( .A1(new_n711_), .A2(new_n624_), .ZN(new_n712_) );
  AND2_X1 g590 ( .A1(new_n712_), .A2(KEYINPUT35), .ZN(new_n713_) );
  OR2_X1 g591 ( .A1(new_n708_), .A2(new_n713_), .ZN(new_n714_) );
  AND2_X1 g592 ( .A1(new_n714_), .A2(G122), .ZN(new_n715_) );
  OR2_X1 g593 ( .A1(new_n712_), .A2(KEYINPUT35), .ZN(new_n716_) );
  OR2_X1 g594 ( .A1(new_n707_), .A2(new_n685_), .ZN(new_n717_) );
  AND2_X1 g595 ( .A1(new_n717_), .A2(new_n716_), .ZN(new_n718_) );
  AND2_X1 g596 ( .A1(new_n718_), .A2(new_n185_), .ZN(new_n719_) );
  OR2_X1 g597 ( .A1(new_n715_), .A2(new_n719_), .ZN(G24) );
  INV_X1 g598 ( .A(KEYINPUT37), .ZN(new_n721_) );
  AND2_X1 g599 ( .A1(new_n693_), .A2(new_n598_), .ZN(new_n722_) );
  AND2_X1 g600 ( .A1(new_n561_), .A2(new_n722_), .ZN(new_n723_) );
  AND2_X1 g601 ( .A1(new_n723_), .A2(new_n382_), .ZN(new_n724_) );
  INV_X1 g602 ( .A(new_n724_), .ZN(new_n725_) );
  AND2_X1 g603 ( .A1(new_n725_), .A2(KEYINPUT36), .ZN(new_n726_) );
  INV_X1 g604 ( .A(new_n726_), .ZN(new_n727_) );
  OR2_X1 g605 ( .A1(new_n725_), .A2(KEYINPUT36), .ZN(new_n728_) );
  AND2_X1 g606 ( .A1(new_n728_), .A2(new_n638_), .ZN(new_n729_) );
  AND2_X1 g607 ( .A1(new_n729_), .A2(new_n727_), .ZN(new_n730_) );
  INV_X1 g608 ( .A(new_n730_), .ZN(new_n731_) );
  AND2_X1 g609 ( .A1(new_n731_), .A2(G125), .ZN(new_n732_) );
  AND2_X1 g610 ( .A1(new_n730_), .A2(new_n203_), .ZN(new_n733_) );
  OR2_X1 g611 ( .A1(new_n732_), .A2(new_n733_), .ZN(new_n734_) );
  AND2_X1 g612 ( .A1(new_n734_), .A2(new_n721_), .ZN(new_n735_) );
  INV_X1 g613 ( .A(new_n734_), .ZN(new_n736_) );
  AND2_X1 g614 ( .A1(new_n736_), .A2(KEYINPUT37), .ZN(new_n737_) );
  OR2_X1 g615 ( .A1(new_n737_), .A2(new_n735_), .ZN(G27) );
  INV_X1 g616 ( .A(new_n561_), .ZN(new_n739_) );
  INV_X1 g617 ( .A(KEYINPUT39), .ZN(new_n740_) );
  AND2_X1 g618 ( .A1(new_n404_), .A2(KEYINPUT38), .ZN(new_n741_) );
  INV_X1 g619 ( .A(new_n741_), .ZN(new_n742_) );
  OR2_X1 g620 ( .A1(new_n404_), .A2(KEYINPUT38), .ZN(new_n743_) );
  AND2_X1 g621 ( .A1(new_n742_), .A2(new_n743_), .ZN(new_n744_) );
  INV_X1 g622 ( .A(new_n744_), .ZN(new_n745_) );
  AND2_X1 g623 ( .A1(new_n623_), .A2(new_n745_), .ZN(new_n746_) );
  OR2_X1 g624 ( .A1(new_n746_), .A2(new_n740_), .ZN(new_n747_) );
  INV_X1 g625 ( .A(new_n596_), .ZN(new_n748_) );
  OR2_X1 g626 ( .A1(new_n557_), .A2(new_n748_), .ZN(new_n749_) );
  OR2_X1 g627 ( .A1(new_n749_), .A2(new_n620_), .ZN(new_n750_) );
  OR2_X1 g628 ( .A1(new_n750_), .A2(new_n744_), .ZN(new_n751_) );
  OR2_X1 g629 ( .A1(new_n751_), .A2(KEYINPUT39), .ZN(new_n752_) );
  AND2_X1 g630 ( .A1(new_n747_), .A2(new_n752_), .ZN(new_n753_) );
  OR2_X1 g631 ( .A1(new_n753_), .A2(new_n739_), .ZN(new_n754_) );
  AND2_X1 g632 ( .A1(new_n754_), .A2(KEYINPUT40), .ZN(new_n755_) );
  INV_X1 g633 ( .A(KEYINPUT40), .ZN(new_n756_) );
  AND2_X1 g634 ( .A1(new_n751_), .A2(KEYINPUT39), .ZN(new_n757_) );
  AND2_X1 g635 ( .A1(new_n746_), .A2(new_n740_), .ZN(new_n758_) );
  OR2_X1 g636 ( .A1(new_n758_), .A2(new_n757_), .ZN(new_n759_) );
  AND2_X1 g637 ( .A1(new_n759_), .A2(new_n561_), .ZN(new_n760_) );
  AND2_X1 g638 ( .A1(new_n760_), .A2(new_n756_), .ZN(new_n761_) );
  OR2_X1 g639 ( .A1(new_n755_), .A2(new_n761_), .ZN(new_n762_) );
  AND2_X1 g640 ( .A1(new_n762_), .A2(G131), .ZN(new_n763_) );
  OR2_X1 g641 ( .A1(new_n760_), .A2(new_n756_), .ZN(new_n764_) );
  OR2_X1 g642 ( .A1(new_n754_), .A2(KEYINPUT40), .ZN(new_n765_) );
  AND2_X1 g643 ( .A1(new_n765_), .A2(new_n764_), .ZN(new_n766_) );
  AND2_X1 g644 ( .A1(new_n766_), .A2(new_n235_), .ZN(new_n767_) );
  OR2_X1 g645 ( .A1(new_n763_), .A2(new_n767_), .ZN(G33) );
  AND2_X1 g646 ( .A1(new_n759_), .A2(new_n570_), .ZN(new_n769_) );
  INV_X1 g647 ( .A(new_n769_), .ZN(new_n770_) );
  AND2_X1 g648 ( .A1(new_n770_), .A2(G134), .ZN(new_n771_) );
  AND2_X1 g649 ( .A1(new_n769_), .A2(new_n183_), .ZN(new_n772_) );
  OR2_X1 g650 ( .A1(new_n771_), .A2(new_n772_), .ZN(G36) );
  INV_X1 g651 ( .A(KEYINPUT42), .ZN(new_n774_) );
  INV_X1 g652 ( .A(new_n604_), .ZN(new_n775_) );
  INV_X1 g653 ( .A(KEYINPUT41), .ZN(new_n776_) );
  AND2_X1 g654 ( .A1(new_n745_), .A2(new_n381_), .ZN(new_n777_) );
  AND2_X1 g655 ( .A1(new_n271_), .A2(new_n777_), .ZN(new_n778_) );
  INV_X1 g656 ( .A(new_n778_), .ZN(new_n779_) );
  AND2_X1 g657 ( .A1(new_n779_), .A2(new_n776_), .ZN(new_n780_) );
  AND2_X1 g658 ( .A1(new_n778_), .A2(KEYINPUT41), .ZN(new_n781_) );
  OR2_X1 g659 ( .A1(new_n780_), .A2(new_n781_), .ZN(new_n782_) );
  OR2_X1 g660 ( .A1(new_n782_), .A2(new_n775_), .ZN(new_n783_) );
  AND2_X1 g661 ( .A1(new_n783_), .A2(new_n774_), .ZN(new_n784_) );
  INV_X1 g662 ( .A(new_n784_), .ZN(new_n785_) );
  OR2_X1 g663 ( .A1(new_n783_), .A2(new_n774_), .ZN(new_n786_) );
  AND2_X1 g664 ( .A1(new_n785_), .A2(new_n786_), .ZN(new_n787_) );
  INV_X1 g665 ( .A(new_n787_), .ZN(new_n788_) );
  AND2_X1 g666 ( .A1(new_n788_), .A2(new_n425_), .ZN(new_n789_) );
  AND2_X1 g667 ( .A1(new_n787_), .A2(G137), .ZN(new_n790_) );
  OR2_X1 g668 ( .A1(new_n789_), .A2(new_n790_), .ZN(G39) );
  AND2_X1 g669 ( .A1(new_n456_), .A2(new_n381_), .ZN(new_n792_) );
  AND2_X1 g670 ( .A1(new_n723_), .A2(new_n792_), .ZN(new_n793_) );
  AND2_X1 g671 ( .A1(new_n793_), .A2(KEYINPUT43), .ZN(new_n794_) );
  INV_X1 g672 ( .A(new_n794_), .ZN(new_n795_) );
  OR2_X1 g673 ( .A1(new_n793_), .A2(KEYINPUT43), .ZN(new_n796_) );
  AND2_X1 g674 ( .A1(new_n796_), .A2(new_n404_), .ZN(new_n797_) );
  AND2_X1 g675 ( .A1(new_n797_), .A2(new_n795_), .ZN(new_n798_) );
  INV_X1 g676 ( .A(new_n798_), .ZN(new_n799_) );
  AND2_X1 g677 ( .A1(new_n799_), .A2(G140), .ZN(new_n800_) );
  AND2_X1 g678 ( .A1(new_n798_), .A2(new_n208_), .ZN(new_n801_) );
  OR2_X1 g679 ( .A1(new_n800_), .A2(new_n801_), .ZN(G42) );
  INV_X1 g680 ( .A(KEYINPUT53), .ZN(new_n803_) );
  INV_X1 g681 ( .A(KEYINPUT44), .ZN(new_n804_) );
  AND2_X1 g682 ( .A1(new_n588_), .A2(new_n678_), .ZN(new_n805_) );
  AND2_X1 g683 ( .A1(new_n714_), .A2(new_n805_), .ZN(new_n806_) );
  AND2_X1 g684 ( .A1(new_n806_), .A2(new_n804_), .ZN(new_n807_) );
  OR2_X1 g685 ( .A1(new_n682_), .A2(new_n587_), .ZN(new_n808_) );
  OR2_X1 g686 ( .A1(new_n718_), .A2(new_n808_), .ZN(new_n809_) );
  AND2_X1 g687 ( .A1(new_n809_), .A2(KEYINPUT44), .ZN(new_n810_) );
  OR2_X1 g688 ( .A1(new_n570_), .A2(new_n561_), .ZN(new_n811_) );
  OR2_X1 g689 ( .A1(new_n647_), .A2(new_n560_), .ZN(new_n812_) );
  AND2_X1 g690 ( .A1(new_n812_), .A2(new_n811_), .ZN(new_n813_) );
  OR2_X1 g691 ( .A1(new_n813_), .A2(new_n550_), .ZN(new_n814_) );
  OR2_X1 g692 ( .A1(new_n810_), .A2(new_n814_), .ZN(new_n815_) );
  OR2_X1 g693 ( .A1(new_n815_), .A2(new_n807_), .ZN(new_n816_) );
  AND2_X1 g694 ( .A1(new_n816_), .A2(KEYINPUT45), .ZN(new_n817_) );
  INV_X1 g695 ( .A(KEYINPUT45), .ZN(new_n818_) );
  INV_X1 g696 ( .A(new_n807_), .ZN(new_n819_) );
  OR2_X1 g697 ( .A1(new_n806_), .A2(new_n804_), .ZN(new_n820_) );
  INV_X1 g698 ( .A(new_n814_), .ZN(new_n821_) );
  AND2_X1 g699 ( .A1(new_n820_), .A2(new_n821_), .ZN(new_n822_) );
  AND2_X1 g700 ( .A1(new_n822_), .A2(new_n819_), .ZN(new_n823_) );
  AND2_X1 g701 ( .A1(new_n823_), .A2(new_n818_), .ZN(new_n824_) );
  OR2_X1 g702 ( .A1(new_n817_), .A2(new_n824_), .ZN(new_n825_) );
  INV_X1 g703 ( .A(KEYINPUT48), .ZN(new_n826_) );
  INV_X1 g704 ( .A(KEYINPUT46), .ZN(new_n827_) );
  OR2_X1 g705 ( .A1(new_n766_), .A2(new_n788_), .ZN(new_n828_) );
  AND2_X1 g706 ( .A1(new_n828_), .A2(new_n827_), .ZN(new_n829_) );
  AND2_X1 g707 ( .A1(new_n762_), .A2(new_n787_), .ZN(new_n830_) );
  AND2_X1 g708 ( .A1(new_n830_), .A2(KEYINPUT46), .ZN(new_n831_) );
  OR2_X1 g709 ( .A1(new_n829_), .A2(new_n831_), .ZN(new_n832_) );
  AND2_X1 g710 ( .A1(new_n731_), .A2(new_n628_), .ZN(new_n833_) );
  INV_X1 g711 ( .A(KEYINPUT47), .ZN(new_n834_) );
  AND2_X1 g712 ( .A1(new_n605_), .A2(new_n811_), .ZN(new_n835_) );
  OR2_X1 g713 ( .A1(new_n835_), .A2(new_n834_), .ZN(new_n836_) );
  AND2_X1 g714 ( .A1(new_n835_), .A2(new_n834_), .ZN(new_n837_) );
  INV_X1 g715 ( .A(new_n837_), .ZN(new_n838_) );
  AND2_X1 g716 ( .A1(new_n838_), .A2(new_n836_), .ZN(new_n839_) );
  AND2_X1 g717 ( .A1(new_n833_), .A2(new_n839_), .ZN(new_n840_) );
  AND2_X1 g718 ( .A1(new_n832_), .A2(new_n840_), .ZN(new_n841_) );
  AND2_X1 g719 ( .A1(new_n841_), .A2(new_n826_), .ZN(new_n842_) );
  INV_X1 g720 ( .A(new_n842_), .ZN(new_n843_) );
  OR2_X1 g721 ( .A1(new_n841_), .A2(new_n826_), .ZN(new_n844_) );
  AND2_X1 g722 ( .A1(new_n770_), .A2(new_n799_), .ZN(new_n845_) );
  AND2_X1 g723 ( .A1(new_n844_), .A2(new_n845_), .ZN(new_n846_) );
  AND2_X1 g724 ( .A1(new_n846_), .A2(new_n843_), .ZN(new_n847_) );
  AND2_X1 g725 ( .A1(new_n825_), .A2(new_n847_), .ZN(new_n848_) );
  OR2_X1 g726 ( .A1(new_n848_), .A2(KEYINPUT2), .ZN(new_n849_) );
  INV_X1 g727 ( .A(KEYINPUT2), .ZN(new_n850_) );
  OR2_X1 g728 ( .A1(new_n823_), .A2(new_n818_), .ZN(new_n851_) );
  OR2_X1 g729 ( .A1(new_n816_), .A2(KEYINPUT45), .ZN(new_n852_) );
  AND2_X1 g730 ( .A1(new_n852_), .A2(new_n851_), .ZN(new_n853_) );
  OR2_X1 g731 ( .A1(new_n830_), .A2(KEYINPUT46), .ZN(new_n854_) );
  OR2_X1 g732 ( .A1(new_n828_), .A2(new_n827_), .ZN(new_n855_) );
  AND2_X1 g733 ( .A1(new_n855_), .A2(new_n854_), .ZN(new_n856_) );
  INV_X1 g734 ( .A(new_n840_), .ZN(new_n857_) );
  OR2_X1 g735 ( .A1(new_n856_), .A2(new_n857_), .ZN(new_n858_) );
  AND2_X1 g736 ( .A1(new_n858_), .A2(KEYINPUT48), .ZN(new_n859_) );
  INV_X1 g737 ( .A(new_n845_), .ZN(new_n860_) );
  OR2_X1 g738 ( .A1(new_n859_), .A2(new_n860_), .ZN(new_n861_) );
  OR2_X1 g739 ( .A1(new_n861_), .A2(new_n842_), .ZN(new_n862_) );
  OR2_X1 g740 ( .A1(new_n853_), .A2(new_n862_), .ZN(new_n863_) );
  OR2_X1 g741 ( .A1(new_n863_), .A2(new_n850_), .ZN(new_n864_) );
  AND2_X1 g742 ( .A1(new_n864_), .A2(new_n849_), .ZN(new_n865_) );
  INV_X1 g743 ( .A(KEYINPUT51), .ZN(new_n866_) );
  AND2_X1 g744 ( .A1(new_n456_), .A2(new_n556_), .ZN(new_n867_) );
  AND2_X1 g745 ( .A1(new_n867_), .A2(KEYINPUT50), .ZN(new_n868_) );
  INV_X1 g746 ( .A(new_n868_), .ZN(new_n869_) );
  OR2_X1 g747 ( .A1(new_n867_), .A2(KEYINPUT50), .ZN(new_n870_) );
  INV_X1 g748 ( .A(KEYINPUT49), .ZN(new_n871_) );
  AND2_X1 g749 ( .A1(new_n506_), .A2(new_n555_), .ZN(new_n872_) );
  AND2_X1 g750 ( .A1(new_n872_), .A2(new_n871_), .ZN(new_n873_) );
  INV_X1 g751 ( .A(new_n873_), .ZN(new_n874_) );
  OR2_X1 g752 ( .A1(new_n872_), .A2(new_n871_), .ZN(new_n875_) );
  AND2_X1 g753 ( .A1(new_n875_), .A2(new_n546_), .ZN(new_n876_) );
  AND2_X1 g754 ( .A1(new_n876_), .A2(new_n874_), .ZN(new_n877_) );
  AND2_X1 g755 ( .A1(new_n870_), .A2(new_n877_), .ZN(new_n878_) );
  AND2_X1 g756 ( .A1(new_n878_), .A2(new_n869_), .ZN(new_n879_) );
  OR2_X1 g757 ( .A1(new_n879_), .A2(new_n641_), .ZN(new_n880_) );
  INV_X1 g758 ( .A(new_n880_), .ZN(new_n881_) );
  AND2_X1 g759 ( .A1(new_n881_), .A2(new_n866_), .ZN(new_n882_) );
  AND2_X1 g760 ( .A1(new_n880_), .A2(KEYINPUT51), .ZN(new_n883_) );
  OR2_X1 g761 ( .A1(new_n883_), .A2(new_n782_), .ZN(new_n884_) );
  OR2_X1 g762 ( .A1(new_n884_), .A2(new_n882_), .ZN(new_n885_) );
  AND2_X1 g763 ( .A1(new_n811_), .A2(new_n777_), .ZN(new_n886_) );
  INV_X1 g764 ( .A(new_n886_), .ZN(new_n887_) );
  AND2_X1 g765 ( .A1(new_n744_), .A2(new_n380_), .ZN(new_n888_) );
  OR2_X1 g766 ( .A1(new_n658_), .A2(new_n888_), .ZN(new_n889_) );
  AND2_X1 g767 ( .A1(new_n887_), .A2(new_n889_), .ZN(new_n890_) );
  OR2_X1 g768 ( .A1(new_n890_), .A2(new_n703_), .ZN(new_n891_) );
  AND2_X1 g769 ( .A1(new_n885_), .A2(new_n891_), .ZN(new_n892_) );
  AND2_X1 g770 ( .A1(new_n892_), .A2(KEYINPUT52), .ZN(new_n893_) );
  INV_X1 g771 ( .A(new_n893_), .ZN(new_n894_) );
  OR2_X1 g772 ( .A1(new_n892_), .A2(KEYINPUT52), .ZN(new_n895_) );
  AND2_X1 g773 ( .A1(new_n895_), .A2(new_n394_), .ZN(new_n896_) );
  AND2_X1 g774 ( .A1(new_n896_), .A2(new_n894_), .ZN(new_n897_) );
  INV_X1 g775 ( .A(new_n782_), .ZN(new_n898_) );
  AND2_X1 g776 ( .A1(new_n898_), .A2(new_n697_), .ZN(new_n899_) );
  OR2_X1 g777 ( .A1(new_n899_), .A2(G953), .ZN(new_n900_) );
  OR2_X1 g778 ( .A1(new_n897_), .A2(new_n900_), .ZN(new_n901_) );
  OR2_X1 g779 ( .A1(new_n865_), .A2(new_n901_), .ZN(new_n902_) );
  AND2_X1 g780 ( .A1(new_n902_), .A2(new_n803_), .ZN(new_n903_) );
  INV_X1 g781 ( .A(new_n902_), .ZN(new_n904_) );
  AND2_X1 g782 ( .A1(new_n904_), .A2(KEYINPUT53), .ZN(new_n905_) );
  OR2_X1 g783 ( .A1(new_n905_), .A2(new_n903_), .ZN(G75) );
  INV_X1 g784 ( .A(KEYINPUT56), .ZN(new_n907_) );
  AND2_X1 g785 ( .A1(new_n130_), .A2(G210), .ZN(new_n908_) );
  AND2_X1 g786 ( .A1(new_n865_), .A2(new_n908_), .ZN(new_n909_) );
  AND2_X1 g787 ( .A1(KEYINPUT55), .A2(KEYINPUT54), .ZN(new_n910_) );
  INV_X1 g788 ( .A(new_n910_), .ZN(new_n911_) );
  OR2_X1 g789 ( .A1(KEYINPUT55), .A2(KEYINPUT54), .ZN(new_n912_) );
  AND2_X1 g790 ( .A1(new_n911_), .A2(new_n912_), .ZN(new_n913_) );
  AND2_X1 g791 ( .A1(new_n367_), .A2(new_n913_), .ZN(new_n914_) );
  INV_X1 g792 ( .A(new_n914_), .ZN(new_n915_) );
  OR2_X1 g793 ( .A1(new_n367_), .A2(new_n913_), .ZN(new_n916_) );
  AND2_X1 g794 ( .A1(new_n915_), .A2(new_n916_), .ZN(new_n917_) );
  AND2_X1 g795 ( .A1(new_n909_), .A2(new_n917_), .ZN(new_n918_) );
  OR2_X1 g796 ( .A1(new_n145_), .A2(G952), .ZN(new_n919_) );
  INV_X1 g797 ( .A(new_n919_), .ZN(new_n920_) );
  AND2_X1 g798 ( .A1(new_n863_), .A2(new_n850_), .ZN(new_n921_) );
  AND2_X1 g799 ( .A1(new_n848_), .A2(KEYINPUT2), .ZN(new_n922_) );
  OR2_X1 g800 ( .A1(new_n921_), .A2(new_n922_), .ZN(new_n923_) );
  INV_X1 g801 ( .A(new_n908_), .ZN(new_n924_) );
  OR2_X1 g802 ( .A1(new_n923_), .A2(new_n924_), .ZN(new_n925_) );
  INV_X1 g803 ( .A(new_n917_), .ZN(new_n926_) );
  AND2_X1 g804 ( .A1(new_n925_), .A2(new_n926_), .ZN(new_n927_) );
  OR2_X1 g805 ( .A1(new_n927_), .A2(new_n920_), .ZN(new_n928_) );
  OR2_X1 g806 ( .A1(new_n928_), .A2(new_n918_), .ZN(new_n929_) );
  AND2_X1 g807 ( .A1(new_n929_), .A2(new_n907_), .ZN(new_n930_) );
  INV_X1 g808 ( .A(new_n918_), .ZN(new_n931_) );
  OR2_X1 g809 ( .A1(new_n909_), .A2(new_n917_), .ZN(new_n932_) );
  AND2_X1 g810 ( .A1(new_n932_), .A2(new_n919_), .ZN(new_n933_) );
  AND2_X1 g811 ( .A1(new_n933_), .A2(new_n931_), .ZN(new_n934_) );
  AND2_X1 g812 ( .A1(new_n934_), .A2(KEYINPUT56), .ZN(new_n935_) );
  OR2_X1 g813 ( .A1(new_n930_), .A2(new_n935_), .ZN(G51) );
  AND2_X1 g814 ( .A1(new_n130_), .A2(G469), .ZN(new_n937_) );
  AND2_X1 g815 ( .A1(new_n865_), .A2(new_n937_), .ZN(new_n938_) );
  INV_X1 g816 ( .A(KEYINPUT57), .ZN(new_n939_) );
  AND2_X1 g817 ( .A1(new_n939_), .A2(KEYINPUT58), .ZN(new_n940_) );
  INV_X1 g818 ( .A(new_n940_), .ZN(new_n941_) );
  OR2_X1 g819 ( .A1(new_n939_), .A2(KEYINPUT58), .ZN(new_n942_) );
  AND2_X1 g820 ( .A1(new_n941_), .A2(new_n942_), .ZN(new_n943_) );
  OR2_X1 g821 ( .A1(new_n938_), .A2(new_n943_), .ZN(new_n944_) );
  INV_X1 g822 ( .A(new_n937_), .ZN(new_n945_) );
  OR2_X1 g823 ( .A1(new_n923_), .A2(new_n945_), .ZN(new_n946_) );
  INV_X1 g824 ( .A(new_n943_), .ZN(new_n947_) );
  OR2_X1 g825 ( .A1(new_n946_), .A2(new_n947_), .ZN(new_n948_) );
  AND2_X1 g826 ( .A1(new_n948_), .A2(new_n944_), .ZN(new_n949_) );
  INV_X1 g827 ( .A(new_n949_), .ZN(new_n950_) );
  OR2_X1 g828 ( .A1(new_n950_), .A2(new_n445_), .ZN(new_n951_) );
  INV_X1 g829 ( .A(new_n445_), .ZN(new_n952_) );
  OR2_X1 g830 ( .A1(new_n949_), .A2(new_n952_), .ZN(new_n953_) );
  AND2_X1 g831 ( .A1(new_n953_), .A2(new_n919_), .ZN(new_n954_) );
  AND2_X1 g832 ( .A1(new_n954_), .A2(new_n951_), .ZN(G54) );
  INV_X1 g833 ( .A(KEYINPUT60), .ZN(new_n956_) );
  AND2_X1 g834 ( .A1(new_n130_), .A2(G475), .ZN(new_n957_) );
  INV_X1 g835 ( .A(new_n957_), .ZN(new_n958_) );
  OR2_X1 g836 ( .A1(new_n923_), .A2(new_n958_), .ZN(new_n959_) );
  INV_X1 g837 ( .A(new_n259_), .ZN(new_n960_) );
  AND2_X1 g838 ( .A1(new_n960_), .A2(KEYINPUT59), .ZN(new_n961_) );
  INV_X1 g839 ( .A(new_n961_), .ZN(new_n962_) );
  OR2_X1 g840 ( .A1(new_n960_), .A2(KEYINPUT59), .ZN(new_n963_) );
  AND2_X1 g841 ( .A1(new_n962_), .A2(new_n963_), .ZN(new_n964_) );
  INV_X1 g842 ( .A(new_n964_), .ZN(new_n965_) );
  AND2_X1 g843 ( .A1(new_n959_), .A2(new_n965_), .ZN(new_n966_) );
  AND2_X1 g844 ( .A1(new_n865_), .A2(new_n957_), .ZN(new_n967_) );
  AND2_X1 g845 ( .A1(new_n967_), .A2(new_n964_), .ZN(new_n968_) );
  OR2_X1 g846 ( .A1(new_n968_), .A2(new_n920_), .ZN(new_n969_) );
  OR2_X1 g847 ( .A1(new_n969_), .A2(new_n966_), .ZN(new_n970_) );
  AND2_X1 g848 ( .A1(new_n970_), .A2(new_n956_), .ZN(new_n971_) );
  INV_X1 g849 ( .A(new_n966_), .ZN(new_n972_) );
  OR2_X1 g850 ( .A1(new_n959_), .A2(new_n965_), .ZN(new_n973_) );
  AND2_X1 g851 ( .A1(new_n973_), .A2(new_n919_), .ZN(new_n974_) );
  AND2_X1 g852 ( .A1(new_n974_), .A2(new_n972_), .ZN(new_n975_) );
  AND2_X1 g853 ( .A1(new_n975_), .A2(KEYINPUT60), .ZN(new_n976_) );
  OR2_X1 g854 ( .A1(new_n976_), .A2(new_n971_), .ZN(G60) );
  AND2_X1 g855 ( .A1(new_n130_), .A2(G478), .ZN(new_n978_) );
  AND2_X1 g856 ( .A1(new_n865_), .A2(new_n978_), .ZN(new_n979_) );
  OR2_X1 g857 ( .A1(new_n979_), .A2(new_n199_), .ZN(new_n980_) );
  INV_X1 g858 ( .A(new_n979_), .ZN(new_n981_) );
  OR2_X1 g859 ( .A1(new_n981_), .A2(new_n192_), .ZN(new_n982_) );
  AND2_X1 g860 ( .A1(new_n982_), .A2(new_n919_), .ZN(new_n983_) );
  AND2_X1 g861 ( .A1(new_n983_), .A2(new_n980_), .ZN(G63) );
  AND2_X1 g862 ( .A1(new_n130_), .A2(G217), .ZN(new_n985_) );
  AND2_X1 g863 ( .A1(new_n865_), .A2(new_n985_), .ZN(new_n986_) );
  OR2_X1 g864 ( .A1(new_n986_), .A2(new_n496_), .ZN(new_n987_) );
  INV_X1 g865 ( .A(new_n986_), .ZN(new_n988_) );
  OR2_X1 g866 ( .A1(new_n988_), .A2(new_n492_), .ZN(new_n989_) );
  AND2_X1 g867 ( .A1(new_n989_), .A2(new_n919_), .ZN(new_n990_) );
  AND2_X1 g868 ( .A1(new_n990_), .A2(new_n987_), .ZN(G66) );
  AND2_X1 g869 ( .A1(new_n825_), .A2(new_n145_), .ZN(new_n992_) );
  AND2_X1 g870 ( .A1(G224), .A2(G953), .ZN(new_n993_) );
  OR2_X1 g871 ( .A1(new_n993_), .A2(KEYINPUT61), .ZN(new_n994_) );
  AND2_X1 g872 ( .A1(new_n993_), .A2(KEYINPUT61), .ZN(new_n995_) );
  OR2_X1 g873 ( .A1(new_n995_), .A2(new_n397_), .ZN(new_n996_) );
  INV_X1 g874 ( .A(new_n996_), .ZN(new_n997_) );
  AND2_X1 g875 ( .A1(new_n997_), .A2(new_n994_), .ZN(new_n998_) );
  OR2_X1 g876 ( .A1(new_n992_), .A2(new_n998_), .ZN(new_n999_) );
  AND2_X1 g877 ( .A1(new_n351_), .A2(G101), .ZN(new_n1000_) );
  AND2_X1 g878 ( .A1(new_n356_), .A2(new_n123_), .ZN(new_n1001_) );
  OR2_X1 g879 ( .A1(new_n1001_), .A2(new_n1000_), .ZN(new_n1002_) );
  INV_X1 g880 ( .A(new_n1002_), .ZN(new_n1003_) );
  AND2_X1 g881 ( .A1(new_n1003_), .A2(new_n327_), .ZN(new_n1004_) );
  AND2_X1 g882 ( .A1(new_n1002_), .A2(new_n300_), .ZN(new_n1005_) );
  OR2_X1 g883 ( .A1(new_n1005_), .A2(new_n398_), .ZN(new_n1006_) );
  OR2_X1 g884 ( .A1(new_n1006_), .A2(new_n1004_), .ZN(new_n1007_) );
  INV_X1 g885 ( .A(new_n1007_), .ZN(new_n1008_) );
  AND2_X1 g886 ( .A1(new_n999_), .A2(new_n1008_), .ZN(new_n1009_) );
  INV_X1 g887 ( .A(new_n999_), .ZN(new_n1010_) );
  AND2_X1 g888 ( .A1(new_n1010_), .A2(new_n1007_), .ZN(new_n1011_) );
  OR2_X1 g889 ( .A1(new_n1011_), .A2(new_n1009_), .ZN(G69) );
  AND2_X1 g890 ( .A1(new_n337_), .A2(new_n207_), .ZN(new_n1013_) );
  AND2_X1 g891 ( .A1(new_n341_), .A2(new_n224_), .ZN(new_n1014_) );
  OR2_X1 g892 ( .A1(new_n1013_), .A2(new_n1014_), .ZN(new_n1015_) );
  INV_X1 g893 ( .A(new_n1015_), .ZN(new_n1016_) );
  AND2_X1 g894 ( .A1(new_n437_), .A2(new_n1016_), .ZN(new_n1017_) );
  AND2_X1 g895 ( .A1(new_n438_), .A2(new_n1015_), .ZN(new_n1018_) );
  OR2_X1 g896 ( .A1(new_n1018_), .A2(new_n1017_), .ZN(new_n1019_) );
  INV_X1 g897 ( .A(new_n1019_), .ZN(new_n1020_) );
  AND2_X1 g898 ( .A1(new_n847_), .A2(new_n1020_), .ZN(new_n1021_) );
  AND2_X1 g899 ( .A1(new_n862_), .A2(new_n1019_), .ZN(new_n1022_) );
  OR2_X1 g900 ( .A1(new_n1022_), .A2(new_n1021_), .ZN(new_n1023_) );
  AND2_X1 g901 ( .A1(new_n1023_), .A2(new_n145_), .ZN(new_n1024_) );
  AND2_X1 g902 ( .A1(new_n1020_), .A2(G227), .ZN(new_n1025_) );
  INV_X1 g903 ( .A(G227), .ZN(new_n1026_) );
  AND2_X1 g904 ( .A1(new_n1019_), .A2(new_n1026_), .ZN(new_n1027_) );
  OR2_X1 g905 ( .A1(new_n1027_), .A2(new_n593_), .ZN(new_n1028_) );
  OR2_X1 g906 ( .A1(new_n1028_), .A2(new_n1025_), .ZN(new_n1029_) );
  AND2_X1 g907 ( .A1(new_n1029_), .A2(G953), .ZN(new_n1030_) );
  OR2_X1 g908 ( .A1(new_n1024_), .A2(new_n1030_), .ZN(G72) );
  AND2_X1 g909 ( .A1(new_n130_), .A2(G472), .ZN(new_n1032_) );
  INV_X1 g910 ( .A(new_n1032_), .ZN(new_n1033_) );
  OR2_X1 g911 ( .A1(new_n923_), .A2(new_n1033_), .ZN(new_n1034_) );
  AND2_X1 g912 ( .A1(new_n539_), .A2(KEYINPUT62), .ZN(new_n1035_) );
  INV_X1 g913 ( .A(new_n1035_), .ZN(new_n1036_) );
  OR2_X1 g914 ( .A1(new_n539_), .A2(KEYINPUT62), .ZN(new_n1037_) );
  AND2_X1 g915 ( .A1(new_n1036_), .A2(new_n1037_), .ZN(new_n1038_) );
  INV_X1 g916 ( .A(new_n1038_), .ZN(new_n1039_) );
  AND2_X1 g917 ( .A1(new_n1034_), .A2(new_n1039_), .ZN(new_n1040_) );
  AND2_X1 g918 ( .A1(new_n865_), .A2(new_n1032_), .ZN(new_n1041_) );
  AND2_X1 g919 ( .A1(new_n1041_), .A2(new_n1038_), .ZN(new_n1042_) );
  OR2_X1 g920 ( .A1(new_n1042_), .A2(new_n920_), .ZN(new_n1043_) );
  OR2_X1 g921 ( .A1(new_n1043_), .A2(new_n1040_), .ZN(new_n1044_) );
  AND2_X1 g922 ( .A1(new_n1044_), .A2(KEYINPUT63), .ZN(new_n1045_) );
  INV_X1 g923 ( .A(KEYINPUT63), .ZN(new_n1046_) );
  INV_X1 g924 ( .A(new_n1040_), .ZN(new_n1047_) );
  OR2_X1 g925 ( .A1(new_n1034_), .A2(new_n1039_), .ZN(new_n1048_) );
  AND2_X1 g926 ( .A1(new_n1048_), .A2(new_n919_), .ZN(new_n1049_) );
  AND2_X1 g927 ( .A1(new_n1049_), .A2(new_n1047_), .ZN(new_n1050_) );
  AND2_X1 g928 ( .A1(new_n1050_), .A2(new_n1046_), .ZN(new_n1051_) );
  OR2_X1 g929 ( .A1(new_n1051_), .A2(new_n1045_), .ZN(G57) );
endmodule


