module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129, keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134, keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139, keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144, keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149, keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154, keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159, keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164, keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169, keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174, keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179, keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184, keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189, keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194, keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199, keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204, keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209, keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214, keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219, keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224, keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229, keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234, keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239, keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244, keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249, keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254, keyIn_0_255, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129, keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134, keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139, keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144, keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149, keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154, keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159, keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164, keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169, keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174, keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179, keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184, keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189, keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194, keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199, keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204, keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209, keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214, keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219, keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224, keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229, keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234, keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239, keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244, keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249, keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254, keyIn_0_255, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n1668_, new_n1359_, new_n595_, new_n1233_, new_n2051_, new_n1839_, new_n445_, new_n1009_, new_n479_, new_n1105_, new_n1215_, new_n1448_, new_n608_, new_n1743_, new_n501_, new_n1157_, new_n1442_, new_n1345_, new_n421_, new_n777_, new_n1988_, new_n1433_, new_n1517_, new_n1575_, new_n1472_, new_n1048_, new_n1785_, new_n885_, new_n439_, new_n1532_, new_n1808_, new_n390_, new_n1910_, new_n743_, new_n1962_, new_n1327_, new_n1535_, new_n2041_, new_n1922_, new_n566_, new_n641_, new_n1849_, new_n386_, new_n767_, new_n389_, new_n514_, new_n1865_, new_n1351_, new_n556_, new_n636_, new_n1899_, new_n691_, new_n1024_, new_n670_, new_n456_, new_n1125_, new_n1590_, new_n1881_, new_n911_, new_n679_, new_n937_, new_n667_, new_n1879_, new_n1237_, new_n2054_, new_n2026_, new_n1837_, new_n1568_, new_n728_, new_n1479_, new_n1071_, new_n1294_, new_n894_, new_n853_, new_n695_, new_n660_, new_n2038_, new_n1311_, new_n526_, new_n908_, new_n1886_, new_n2023_, new_n552_, new_n678_, new_n1662_, new_n706_, new_n649_, new_n1119_, new_n1213_, new_n752_, new_n2063_, new_n1524_, new_n1045_, new_n1305_, new_n500_, new_n2033_, new_n1163_, new_n786_, new_n2045_, new_n1769_, new_n1103_, new_n1188_, new_n1415_, new_n1390_, new_n721_, new_n504_, new_n1414_, new_n742_, new_n892_, new_n1368_, new_n472_, new_n873_, new_n1919_, new_n1985_, new_n1768_, new_n1167_, new_n1530_, new_n1300_, new_n2070_, new_n1898_, new_n1490_, new_n774_, new_n1777_, new_n792_, new_n1620_, new_n953_, new_n1786_, new_n1946_, new_n481_, new_n1265_, new_n1073_, new_n1110_, new_n1580_, new_n449_, new_n580_, new_n639_, new_n484_, new_n766_, new_n1973_, new_n1212_, new_n1059_, new_n634_, new_n1332_, new_n1851_, new_n1447_, new_n635_, new_n1774_, new_n685_, new_n648_, new_n903_, new_n1595_, new_n1803_, new_n983_, new_n822_, new_n1406_, new_n1990_, new_n1082_, new_n1760_, new_n1018_, new_n1884_, new_n1864_, new_n606_, new_n796_, new_n1054_, new_n655_, new_n1288_, new_n630_, new_n1717_, new_n385_, new_n1670_, new_n1049_, new_n1330_, new_n694_, new_n461_, new_n1323_, new_n565_, new_n1979_, new_n1196_, new_n1366_, new_n1984_, new_n511_, new_n1714_, new_n2034_, new_n1640_, new_n1285_, new_n1031_, new_n1733_, new_n1842_, new_n1216_, new_n1632_, new_n1889_, new_n1987_, new_n1281_, new_n629_, new_n1214_, new_n883_, new_n1911_, new_n1005_, new_n999_, new_n1647_, new_n1816_, new_n1713_, new_n960_, new_n1377_, new_n1522_, new_n549_, new_n491_, new_n676_, new_n995_, new_n1035_, new_n674_, new_n991_, new_n1044_, new_n1362_, new_n1404_, new_n1443_, new_n1484_, new_n2072_, new_n1512_, new_n497_, new_n816_, new_n1355_, new_n1678_, new_n568_, new_n420_, new_n876_, new_n1894_, new_n1900_, new_n1950_, new_n1936_, new_n423_, new_n498_, new_n496_, new_n1217_, new_n1046_, new_n1182_, new_n708_, new_n2032_, new_n1463_, new_n429_, new_n1222_, new_n353_, new_n734_, new_n912_, new_n1424_, new_n1062_, new_n680_, new_n981_, new_n506_, new_n872_, new_n1527_, new_n1275_, new_n1277_, new_n1800_, new_n1198_, new_n1428_, new_n1440_, new_n656_, new_n1127_, new_n388_, new_n1028_, new_n1168_, new_n2012_, new_n483_, new_n1004_, new_n1152_, new_n1558_, new_n394_, new_n935_, new_n1972_, new_n657_, new_n1150_, new_n652_, new_n582_, new_n1020_, new_n363_, new_n1266_, new_n1735_, new_n1113_, new_n785_, new_n1501_, new_n441_, new_n477_, new_n664_, new_n1752_, new_n600_, new_n1737_, new_n1930_, new_n1041_, new_n1657_, new_n1989_, new_n1797_, new_n426_, new_n1036_, new_n1562_, new_n1939_, new_n1953_, new_n398_, new_n1576_, new_n1718_, new_n1333_, new_n395_, new_n1132_, new_n343_, new_n854_, new_n458_, new_n1106_, new_n1740_, new_n1395_, new_n473_, new_n1624_, new_n1147_, new_n1682_, new_n1795_, new_n1373_, new_n1229_, new_n1827_, new_n1422_, new_n1523_, new_n1698_, new_n1468_, new_n1679_, new_n969_, new_n835_, new_n1234_, new_n1360_, new_n378_, new_n1574_, new_n1614_, new_n621_, new_n1423_, new_n1637_, new_n1732_, new_n705_, new_n943_, new_n874_, new_n402_, new_n1798_, new_n1321_, new_n1690_, new_n1209_, new_n1709_, new_n347_, new_n2084_, new_n659_, new_n700_, new_n1419_, new_n921_, new_n346_, new_n396_, new_n1954_, new_n1315_, new_n1003_, new_n696_, new_n1868_, new_n1039_, new_n1507_, new_n1439_, new_n1658_, new_n1952_, new_n1671_, new_n1239_, new_n528_, new_n952_, new_n1870_, new_n1158_, new_n1667_, new_n729_, new_n1111_, new_n1413_, new_n1218_, new_n1385_, new_n1346_, new_n1201_, new_n559_, new_n1282_, new_n1630_, new_n762_, new_n1349_, new_n1193_, new_n1547_, new_n1780_, new_n1994_, new_n1437_, new_n1598_, new_n1187_, new_n1205_, new_n1966_, new_n1154_, new_n1253_, new_n1546_, new_n1453_, new_n1256_, new_n1850_, new_n628_, new_n1513_, new_n409_, new_n1090_, new_n1669_, new_n1489_, new_n553_, new_n745_, new_n1114_, new_n1084_, new_n1061_, new_n668_, new_n834_, new_n1991_, new_n1573_, new_n1781_, new_n1738_, new_n369_, new_n1693_, new_n1171_, new_n867_, new_n954_, new_n1591_, new_n1626_, new_n1032_, new_n1545_, new_n901_, new_n1757_, new_n688_, new_n1255_, new_n1704_, new_n985_, new_n2074_, new_n1995_, new_n851_, new_n1518_, new_n932_, new_n878_, new_n1981_, new_n543_, new_n1943_, new_n1975_, new_n886_, new_n371_, new_n1712_, new_n509_, new_n1761_, new_n2058_, new_n2075_, new_n661_, new_n797_, new_n1358_, new_n724_, new_n1070_, new_n1686_, new_n1416_, new_n1109_, new_n1496_, new_n672_, new_n1269_, new_n616_, new_n1653_, new_n529_, new_n884_, new_n914_, new_n1875_, new_n938_, new_n362_, new_n1600_, new_n1592_, new_n809_, new_n1631_, new_n1142_, new_n1623_, new_n604_, new_n1461_, new_n1104_, new_n1703_, new_n1771_, new_n1511_, new_n571_, new_n1859_, new_n1504_, new_n758_, new_n1802_, new_n460_, new_n1267_, new_n2015_, new_n1794_, new_n1705_, new_n1466_, new_n1707_, new_n1716_, new_n1516_, new_n1299_, new_n380_, new_n1477_, new_n1079_, new_n861_, new_n1564_, new_n1656_, new_n1252_, new_n1993_, new_n1804_, new_n1553_, new_n931_, new_n575_, new_n1493_, new_n1593_, new_n944_, new_n1929_, new_n1638_, new_n1542_, new_n1064_, new_n1949_, new_n1065_, new_n1118_, new_n1645_, new_n493_, new_n547_, new_n1480_, new_n1934_, new_n1745_, new_n1860_, new_n379_, new_n1825_, new_n963_, new_n586_, new_n1481_, new_n1325_, new_n993_, new_n1625_, new_n1357_, new_n1191_, new_n1931_, new_n824_, new_n1628_, new_n717_, new_n1455_, new_n403_, new_n868_, new_n1242_, new_n475_, new_n858_, new_n1612_, new_n1384_, new_n1343_, new_n936_, new_n1459_, new_n1434_, new_n1438_, new_n1016_, new_n411_, new_n673_, new_n1766_, new_n1904_, new_n1144_, new_n2025_, new_n1465_, new_n2082_, new_n666_, new_n1290_, new_n2065_, new_n407_, new_n1897_, new_n1833_, new_n1519_, new_n1407_, new_n1692_, new_n1726_, new_n879_, new_n1417_, new_n1700_, new_n736_, new_n513_, new_n1903_, new_n558_, new_n382_, new_n1370_, new_n718_, new_n1310_, new_n2042_, new_n1710_, new_n1398_, new_n1126_, new_n2047_, new_n546_, new_n612_, new_n1015_, new_n919_, new_n755_, new_n2017_, new_n1040_, new_n1635_, new_n1509_, new_n1559_, new_n1789_, new_n544_, new_n615_, new_n722_, new_n1941_, new_n856_, new_n415_, new_n1324_, new_n1293_, new_n537_, new_n1336_, new_n2068_, new_n2066_, new_n499_, new_n533_, new_n1130_, new_n2064_, new_n795_, new_n459_, new_n1441_, new_n1122_, new_n1728_, new_n1185_, new_n1240_, new_n2031_, new_n1510_, new_n354_, new_n1174_, new_n968_, new_n2001_, new_n2055_, new_n1655_, new_n1464_, new_n613_, new_n1508_, new_n1195_, new_n417_, new_n658_, new_n837_, new_n591_, new_n801_, new_n2039_, new_n1458_, new_n631_, new_n453_, new_n1723_, new_n1818_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n1521_, new_n1334_, new_n2044_, new_n531_, new_n1826_, new_n1675_, new_n593_, new_n1543_, new_n1765_, new_n1907_, new_n1565_, new_n1248_, new_n1812_, new_n751_, new_n1978_, new_n1038_, new_n372_, new_n1758_, new_n852_, new_n1454_, new_n1474_, new_n1328_, new_n978_, new_n1308_, new_n408_, new_n1430_, new_n470_, new_n769_, new_n1660_, new_n433_, new_n871_, new_n1956_, new_n1450_, new_n992_, new_n1098_, new_n1729_, new_n2069_, new_n732_, new_n1832_, new_n689_, new_n933_, new_n584_, new_n815_, new_n1608_, new_n1492_, new_n1367_, new_n1619_, new_n1052_, new_n1425_, new_n1980_, new_n857_, new_n1379_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n1853_, new_n512_, new_n1471_, new_n1673_, new_n1220_, new_n989_, new_n1741_, new_n1117_, new_n1421_, new_n644_, new_n1594_, new_n836_, new_n1856_, new_n1116_, new_n1684_, new_n904_, new_n1392_, new_n1276_, new_n1444_, new_n913_, new_n681_, new_n594_, new_n561_, new_n495_, new_n927_, new_n431_, new_n1206_, new_n1427_, new_n818_, new_n881_, new_n1815_, new_n1268_, new_n2052_, new_n1376_, new_n1381_, new_n1876_, new_n1566_, new_n1534_, new_n684_, new_n640_, new_n1274_, new_n1893_, new_n1665_, new_n754_, new_n1787_, new_n653_, new_n1659_, new_n905_, new_n1258_, new_n1539_, new_n1643_, new_n375_, new_n1958_, new_n962_, new_n1841_, new_n760_, new_n627_, new_n1391_, new_n1724_, new_n1436_, new_n1986_, new_n567_, new_n1353_, new_n1033_, new_n576_, new_n831_, new_n791_, new_n2050_, new_n1153_, new_n1339_, new_n1784_, new_n1970_, new_n984_, new_n780_, new_n1183_, new_n643_, new_n1316_, new_n1194_, new_n1338_, new_n1460_, new_n1878_, new_n1230_, new_n1602_, new_n1027_, new_n610_, new_n1369_, new_n1694_, new_n843_, new_n703_, new_n698_, new_n1639_, new_n1165_, new_n1401_, new_n1259_, new_n1208_, new_n697_, new_n1099_, new_n1023_, new_n951_, new_n1942_, new_n709_, new_n1235_, new_n1320_, new_n540_, new_n1149_, new_n1928_, new_n1066_, new_n1861_, new_n434_, new_n2021_, new_n422_, new_n1944_, new_n581_, new_n1664_, new_n686_, new_n934_, new_n1567_, new_n1651_, new_n770_, new_n1389_, new_n1400_, new_n757_, new_n1225_, new_n521_, new_n793_, new_n406_, new_n1597_, new_n356_, new_n647_, new_n889_, new_n536_, new_n2083_, new_n1616_, new_n1089_, new_n1192_, new_n405_, new_n942_, new_n1806_, new_n614_, new_n895_, new_n958_, new_n976_, new_n699_, new_n1405_, new_n1249_, new_n1354_, new_n955_, new_n1895_, new_n847_, new_n888_, new_n1505_, new_n1340_, new_n798_, new_n1180_, new_n1926_, new_n1969_, new_n1948_, new_n817_, new_n720_, new_n1801_, new_n753_, new_n620_, new_n368_, new_n1361_, new_n941_, new_n1410_, new_n738_, new_n2073_, new_n827_, new_n1356_, new_n1363_, new_n1747_, new_n1317_, new_n366_, new_n779_, new_n1232_, new_n1025_, new_n365_, new_n859_, new_n1211_, new_n1412_, new_n1207_, new_n1176_, new_n1374_, new_n1799_, new_n601_, new_n842_, new_n1552_, new_n1057_, new_n1644_, new_n1677_, new_n682_, new_n1075_, new_n1790_, new_n812_, new_n2030_, new_n1563_, new_n821_, new_n1937_, new_n542_, new_n548_, new_n669_, new_n1397_, new_n1402_, new_n1313_, new_n1172_, new_n419_, new_n624_, new_n534_, new_n1131_, new_n1120_, new_n819_, new_n637_, new_n1603_, new_n1971_, new_n451_, new_n489_, new_n804_, new_n1342_, new_n424_, new_n602_, new_n1210_, new_n1060_, new_n1303_, new_n413_, new_n1906_, new_n1544_, new_n1382_, new_n1896_, new_n442_, new_n677_, new_n1843_, new_n1487_, new_n1646_, new_n642_, new_n1418_, new_n462_, new_n603_, new_n564_, new_n1528_, new_n1814_, new_n1871_, new_n761_, new_n2027_, new_n735_, new_n840_, new_n1283_, new_n1913_, new_n1873_, new_n898_, new_n1734_, new_n799_, new_n1304_, new_n1537_, new_n946_, new_n1764_, new_n1834_, new_n344_, new_n1977_, new_n1108_, new_n1469_, new_n862_, new_n1749_, new_n1606_, new_n1838_, new_n427_, new_n532_, new_n1739_, new_n393_, new_n1617_, new_n418_, new_n746_, new_n1221_, new_n1585_, new_n1587_, new_n1264_, new_n1319_, new_n626_, new_n1680_, new_n1473_, new_n959_, new_n990_, new_n1629_, new_n2005_, new_n716_, new_n701_, new_n1238_, new_n2062_, new_n1676_, new_n1058_, new_n2037_, new_n1880_, new_n1162_, new_n1730_, new_n2018_, new_n2003_, new_n1278_, new_n902_, new_n364_, new_n832_, new_n1996_, new_n1696_, new_n414_, new_n2028_, new_n1968_, new_n1101_, new_n1250_, new_n2011_, new_n1681_, new_n1482_, new_n1050_, new_n554_, new_n1151_, new_n844_, new_n1302_, new_n430_, new_n482_, new_n849_, new_n1203_, new_n855_, new_n1037_, new_n589_, new_n1083_, new_n759_, new_n1297_, new_n1959_, new_n829_, new_n1257_, new_n1306_, new_n1720_, new_n988_, new_n1858_, new_n478_, new_n1307_, new_n1228_, new_n710_, new_n971_, new_n1486_, new_n361_, new_n764_, new_n906_, new_n683_, new_n2081_, new_n1409_, new_n2007_, new_n1429_, new_n1955_, new_n463_, new_n1683_, new_n1372_, new_n510_, new_n966_, new_n1685_, new_n1721_, new_n351_, new_n1877_, new_n1184_, new_n1960_, new_n1292_, new_n1426_, new_n2036_, new_n609_, new_n517_, new_n2077_, new_n1759_, new_n961_, new_n530_, new_n890_, new_n1992_, new_n1006_, new_n1836_, new_n622_, new_n1706_, new_n2006_, new_n702_, new_n2014_, new_n833_, new_n1560_, new_n1701_, new_n1905_, new_n715_, new_n811_, new_n1445_, new_n1371_, new_n443_, new_n1086_, new_n1902_, new_n956_, new_n763_, new_n1622_, new_n1138_, new_n486_, new_n970_, new_n466_, new_n1618_, new_n1652_, new_n1847_, new_n2057_, new_n1170_, new_n845_, new_n768_, new_n1691_, new_n773_, new_n1051_, new_n899_, new_n1053_, new_n1540_, new_n1611_, new_n1823_, new_n1708_, new_n492_, new_n1200_, new_n1533_, new_n650_, new_n750_, new_n1754_, new_n1750_, new_n1767_, new_n887_, new_n355_, new_n926_, new_n432_, new_n925_, new_n2060_, new_n875_, new_n2040_, new_n1226_, new_n1940_, new_n778_, new_n452_, new_n1727_, new_n381_, new_n1483_, new_n1219_, new_n920_, new_n1121_, new_n1495_, new_n1341_, new_n820_, new_n1386_, new_n771_, new_n979_, new_n1819_, new_n508_, new_n1435_, new_n1844_, new_n1748_, new_n1280_, new_n1007_, new_n1613_, new_n1241_, new_n882_, new_n1145_, new_n1557_, new_n929_, new_n986_, new_n1159_, new_n1584_, new_n1337_, new_n1782_, new_n1348_, new_n917_, new_n2071_, new_n1555_, new_n1636_, new_n1322_, new_n1751_, new_n1133_, new_n1822_, new_n1887_, new_n1177_, new_n646_, new_n538_, new_n1026_, new_n2019_, new_n541_, new_n447_, new_n1967_, new_n1388_, new_n1550_, new_n790_, new_n1081_, new_n587_, new_n2010_, new_n1247_, new_n1411_, new_n465_, new_n783_, new_n1380_, new_n2016_, new_n2000_, new_n739_, new_n996_, new_n2080_, new_n1601_, new_n1318_, new_n846_, new_n915_, new_n488_, new_n524_, new_n349_, new_n848_, new_n1921_, new_n1725_, new_n1245_, new_n1772_, new_n663_, new_n1499_, new_n1497_, new_n579_, new_n1791_, new_n2035_, new_n1375_, new_n1908_, new_n1711_, new_n1254_, new_n1689_, new_n438_, new_n1344_, new_n1857_, new_n939_, new_n1393_, new_n632_, new_n1335_, new_n1364_, new_n671_, new_n965_, new_n1514_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n1202_, new_n1526_, new_n397_, new_n1446_, new_n975_, new_n1199_, new_n399_, new_n1581_, new_n596_, new_n945_, new_n870_, new_n805_, new_n1420_, new_n1882_, new_n1115_, new_n1846_, new_n1403_, new_n1866_, new_n1383_, new_n1231_, new_n948_, new_n1520_, new_n1055_, new_n2043_, new_n1431_, new_n838_, new_n1609_, new_n923_, new_n1755_, new_n1674_, new_n469_, new_n437_, new_n1085_, new_n1633_, new_n1607_, new_n359_, new_n794_, new_n1924_, new_n457_, new_n1852_, new_n1301_, new_n1128_, new_n1582_, new_n2056_, new_n1002_, new_n2009_, new_n1169_, new_n1702_, new_n1909_, new_n1810_, new_n448_, new_n1932_, new_n384_, new_n900_, new_n1722_, new_n1824_, new_n1329_, new_n1161_, new_n1788_, new_n1648_, new_n1914_, new_n924_, new_n775_, new_n1867_, new_n454_, new_n1034_, new_n1872_, new_n1124_, new_n1957_, new_n1663_, new_n1000_, new_n1947_, new_n633_, new_n784_, new_n1273_, new_n1396_, new_n1491_, new_n1554_, new_n1923_, new_n2013_, new_n860_, new_n494_, new_n1160_, new_n1166_, new_n1536_, new_n654_, new_n1456_, new_n713_, new_n880_, new_n1102_, new_n1920_, new_n690_, new_n416_, new_n1043_, new_n744_, new_n400_, new_n1175_, new_n1136_, new_n1272_, new_n693_, new_n1287_, new_n1485_, new_n505_, new_n1462_, new_n619_, new_n1890_, new_n471_, new_n967_, new_n577_, new_n1135_, new_n376_, new_n1538_, new_n1579_, new_n1289_, new_n1561_, new_n1271_, new_n1251_, new_n747_, new_n749_, new_n1091_, new_n1095_, new_n998_, new_n1056_, new_n1331_, new_n1094_, new_n1776_, new_n1621_, new_n839_, new_n1030_, new_n2078_, new_n485_, new_n578_, new_n525_, new_n1695_, new_n918_, new_n1586_, new_n1805_, new_n940_, new_n810_, new_n808_, new_n1284_, new_n1572_, new_n907_, new_n665_, new_n800_, new_n897_, new_n1012_, new_n1387_, new_n719_, new_n869_, new_n1178_, new_n1775_, new_n1525_, new_n570_, new_n598_, new_n893_, new_n1935_, new_n1063_, new_n520_, new_n1347_, new_n1001_, new_n1917_, new_n825_, new_n1627_, new_n557_, new_n1642_, new_n1807_, new_n1503_, new_n1742_, new_n507_, new_n741_, new_n806_, new_n1699_, new_n605_, new_n1224_, new_n2008_, new_n748_, new_n1074_, new_n1137_, new_n1286_, new_n1551_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n1141_, new_n1650_, new_n807_, new_n1326_, new_n592_, new_n1820_, new_n726_, new_n1763_, new_n1263_, new_n1123_, new_n2020_, new_n1080_, new_n583_, new_n617_, new_n1279_, new_n1467_, new_n522_, new_n588_, new_n1762_, new_n1997_, new_n916_, new_n781_, new_n1014_, new_n428_, new_n1855_, new_n487_, new_n675_, new_n1155_, new_n360_, new_n1186_, new_n1915_, new_n1596_, new_n1848_, new_n1261_, new_n2022_, new_n2002_, new_n1863_, new_n1246_, new_n1488_, new_n2024_, new_n922_, new_n2029_, new_n387_, new_n476_, new_n987_, new_n1641_, new_n1951_, new_n949_, new_n2048_, new_n450_, new_n1394_, new_n1179_, new_n1088_, new_n1148_, new_n1146_, new_n1756_, new_n569_, new_n555_, new_n468_, new_n977_, new_n2049_, new_n1139_, new_n782_, new_n1793_, new_n444_, new_n392_, new_n518_, new_n950_, new_n1845_, new_n737_, new_n1022_, new_n692_, new_n502_, new_n1821_, new_n1888_, new_n623_, new_n446_, new_n590_, new_n826_, new_n2079_, new_n789_, new_n1476_, new_n515_, new_n1854_, new_n972_, new_n1634_, new_n1067_, new_n891_, new_n516_, new_n1227_, new_n1352_, new_n1835_, new_n1916_, new_n2046_, new_n733_, new_n1983_, new_n1021_, new_n1076_, new_n585_, new_n2076_, new_n1350_, new_n535_, new_n1976_, new_n725_, new_n814_, new_n503_, new_n527_, new_n772_, new_n1244_, new_n1736_, new_n1945_, new_n1378_, new_n1478_, new_n1181_, new_n1093_, new_n597_, new_n1451_, new_n1092_, new_n1783_, new_n1143_, new_n1072_, new_n1190_, new_n1097_, new_n1069_, new_n651_, new_n1164_, new_n1779_, new_n1869_, new_n1296_, new_n435_, new_n1891_, new_n1719_, new_n1883_, new_n1309_, new_n1796_, new_n1010_, new_n776_, new_n1830_, new_n2053_, new_n1885_, new_n687_, new_n1029_, new_n1649_, new_n1862_, new_n1654_, new_n1515_, new_n1746_, new_n638_, new_n523_, new_n909_, new_n1840_, new_n1688_, new_n1963_, new_n1571_, new_n1773_, new_n788_, new_n841_, new_n1457_, new_n1204_, new_n1610_, new_n1470_, new_n1112_, new_n1715_, new_n1156_, new_n711_, new_n1938_, new_n1298_, new_n731_, new_n599_, new_n930_, new_n1475_, new_n1604_, new_n1260_, new_n973_, new_n1529_, new_n607_, new_n1731_, new_n1541_, new_n645_, new_n1087_, new_n1096_, new_n723_, new_n1599_, new_n756_, new_n823_, new_n1549_, new_n1933_, new_n1577_, new_n574_, new_n1500_, new_n928_, new_n1548_, new_n1578_, new_n1008_, new_n2059_, new_n1687_, new_n1661_, new_n1615_, new_n707_, new_n740_, new_n957_, new_n1047_, new_n787_, new_n1134_, new_n1291_, new_n539_, new_n1399_, new_n803_, new_n1270_, new_n1817_, new_n727_, new_n1531_, new_n1672_, new_n1927_, new_n1589_, new_n2061_, new_n1792_, new_n1965_, new_n1295_, new_n1173_, new_n704_, new_n1809_, new_n1432_, new_n1570_, new_n1811_, new_n2004_, new_n1189_, new_n1197_, new_n1912_, new_n1312_, new_n1502_, new_n1778_, new_n1874_, new_n474_, new_n1223_, new_n1129_, new_n1013_, new_n467_, new_n404_, new_n1243_, new_n1077_, new_n2067_, new_n490_, new_n560_, new_n1100_, new_n1666_, new_n865_, new_n1744_, new_n358_, new_n877_, new_n1506_, new_n1583_, new_n2085_, new_n1697_, new_n545_, new_n611_, new_n1998_, new_n1011_, new_n425_, new_n896_, new_n1831_, new_n802_, new_n1925_, new_n1236_, new_n1829_, new_n1770_, new_n866_, new_n1556_, new_n947_, new_n994_, new_n1813_, new_n982_, new_n1494_, new_n1449_, new_n964_, new_n1078_, new_n1961_, new_n551_, new_n1408_, new_n455_, new_n1982_, new_n1569_, new_n618_, new_n1140_, new_n1042_, new_n863_, new_n828_, new_n980_, new_n1918_, new_n1605_, new_n464_, new_n1498_, new_n1588_, new_n1974_, new_n573_, new_n765_, new_n1964_, new_n1314_, new_n1892_;

not g0000 ( new_n343_, N75 );
nand g0001 ( new_n344_, N29, N42 );
nor g0002 ( N388, new_n344_, new_n343_ );
not g0003 ( new_n346_, N80 );
nand g0004 ( new_n347_, N29, N36 );
nor g0005 ( N389, new_n347_, new_n346_ );
not g0006 ( new_n349_, N42 );
nor g0007 ( N390, new_n347_, new_n349_ );
nand g0008 ( new_n351_, N85, N86 );
not g0009 ( N391, new_n351_ );
not g0010 ( new_n353_, N17 );
nand g0011 ( new_n354_, N1, N8 );
not g0012 ( new_n355_, new_n354_ );
nand g0013 ( new_n356_, new_n355_, N13 );
nor g0014 ( N418, new_n356_, new_n353_ );
nand g0015 ( new_n358_, N1, N26 );
nand g0016 ( new_n359_, N13, N17 );
nor g0017 ( new_n360_, new_n358_, new_n359_ );
not g0018 ( new_n361_, new_n360_ );
nor g0019 ( new_n362_, new_n361_, N390 );
not g0020 ( new_n363_, new_n362_ );
nand g0021 ( new_n364_, new_n363_, keyIn_0_8 );
not g0022 ( new_n365_, keyIn_0_8 );
nand g0023 ( new_n366_, new_n362_, new_n365_ );
nand g0024 ( N419, new_n364_, new_n366_ );
nand g0025 ( new_n368_, N59, N75 );
not g0026 ( new_n369_, new_n368_ );
nand g0027 ( N420, new_n369_, N80 );
nand g0028 ( new_n371_, N36, N59 );
not g0029 ( new_n372_, new_n371_ );
nand g0030 ( N421, new_n372_, N80 );
nand g0031 ( N422, new_n372_, N42 );
not g0032 ( new_n375_, N90 );
nor g0033 ( new_n376_, N87, N88 );
nor g0034 ( N423, new_n376_, new_n375_ );
nand g0035 ( new_n378_, new_n360_, N390 );
nand g0036 ( new_n379_, new_n378_, keyIn_0_25 );
not g0037 ( new_n380_, keyIn_0_25 );
not g0038 ( new_n381_, new_n378_ );
nand g0039 ( new_n382_, new_n381_, new_n380_ );
nand g0040 ( N446, new_n382_, new_n379_ );
not g0041 ( new_n384_, keyIn_0_0 );
not g0042 ( new_n385_, N51 );
nor g0043 ( new_n386_, new_n358_, new_n385_ );
nor g0044 ( new_n387_, new_n386_, new_n384_ );
not g0045 ( new_n388_, new_n358_ );
nand g0046 ( new_n389_, new_n388_, N51 );
nor g0047 ( new_n390_, new_n389_, keyIn_0_0 );
nor g0048 ( N447, new_n390_, new_n387_ );
not g0049 ( new_n392_, N55 );
nor g0050 ( new_n393_, new_n356_, new_n392_ );
not g0051 ( new_n394_, new_n393_ );
nand g0052 ( new_n395_, N29, N68 );
nor g0053 ( new_n396_, new_n394_, new_n395_ );
not g0054 ( new_n397_, new_n396_ );
nand g0055 ( new_n398_, new_n397_, keyIn_0_12 );
not g0056 ( new_n399_, keyIn_0_12 );
nand g0057 ( new_n400_, new_n396_, new_n399_ );
nand g0058 ( N448, new_n398_, new_n400_ );
nand g0059 ( new_n402_, N59, N68 );
not g0060 ( new_n403_, new_n402_ );
nand g0061 ( new_n404_, new_n403_, N74 );
nor g0062 ( new_n405_, new_n394_, new_n404_ );
not g0063 ( new_n406_, new_n405_ );
nand g0064 ( new_n407_, new_n406_, keyIn_0_13 );
not g0065 ( new_n408_, keyIn_0_13 );
nand g0066 ( new_n409_, new_n405_, new_n408_ );
nand g0067 ( N449, new_n407_, new_n409_ );
not g0068 ( new_n411_, N89 );
nor g0069 ( N450, new_n376_, new_n411_ );
not g0070 ( new_n413_, keyIn_0_139 );
not g0071 ( new_n414_, keyIn_0_95 );
not g0072 ( new_n415_, keyIn_0_73 );
not g0073 ( new_n416_, keyIn_0_43 );
not g0074 ( new_n417_, keyIn_0_18 );
nor g0075 ( new_n418_, N121, N126 );
nand g0076 ( new_n419_, N121, N126 );
not g0077 ( new_n420_, new_n419_ );
nor g0078 ( new_n421_, new_n420_, new_n418_ );
nor g0079 ( new_n422_, new_n421_, new_n417_ );
nand g0080 ( new_n423_, new_n421_, new_n417_ );
not g0081 ( new_n424_, new_n423_ );
nor g0082 ( new_n425_, new_n424_, new_n422_ );
nor g0083 ( new_n426_, new_n425_, keyIn_0_32 );
nand g0084 ( new_n427_, new_n425_, keyIn_0_32 );
not g0085 ( new_n428_, new_n427_ );
nor g0086 ( new_n429_, new_n428_, new_n426_ );
not g0087 ( new_n430_, N111 );
nor g0088 ( new_n431_, new_n430_, N116 );
not g0089 ( new_n432_, N116 );
nor g0090 ( new_n433_, new_n432_, N111 );
nor g0091 ( new_n434_, new_n431_, new_n433_ );
not g0092 ( new_n435_, new_n434_ );
nand g0093 ( new_n436_, new_n435_, keyIn_0_17 );
not g0094 ( new_n437_, new_n436_ );
nor g0095 ( new_n438_, new_n435_, keyIn_0_17 );
nor g0096 ( new_n439_, new_n437_, new_n438_ );
nor g0097 ( new_n440_, new_n439_, keyIn_0_31 );
nand g0098 ( new_n441_, new_n439_, keyIn_0_31 );
not g0099 ( new_n442_, new_n441_ );
nor g0100 ( new_n443_, new_n442_, new_n440_ );
nor g0101 ( new_n444_, new_n443_, new_n429_ );
not g0102 ( new_n445_, new_n444_ );
nand g0103 ( new_n446_, new_n445_, new_n416_ );
not g0104 ( new_n447_, new_n446_ );
nor g0105 ( new_n448_, new_n445_, new_n416_ );
nor g0106 ( new_n449_, new_n447_, new_n448_ );
not g0107 ( new_n450_, keyIn_0_33 );
nor g0108 ( new_n451_, new_n439_, new_n425_ );
not g0109 ( new_n452_, new_n451_ );
nand g0110 ( new_n453_, new_n452_, new_n450_ );
not g0111 ( new_n454_, new_n453_ );
nor g0112 ( new_n455_, new_n452_, new_n450_ );
nor g0113 ( new_n456_, new_n454_, new_n455_ );
nor g0114 ( new_n457_, new_n449_, new_n456_ );
nor g0115 ( new_n458_, new_n457_, keyIn_0_53 );
nand g0116 ( new_n459_, new_n457_, keyIn_0_53 );
not g0117 ( new_n460_, new_n459_ );
nor g0118 ( new_n461_, new_n460_, new_n458_ );
not g0119 ( new_n462_, new_n461_ );
nor g0120 ( new_n463_, new_n462_, N135 );
nor g0121 ( new_n464_, new_n463_, new_n415_ );
nand g0122 ( new_n465_, new_n463_, new_n415_ );
not g0123 ( new_n466_, new_n465_ );
nor g0124 ( new_n467_, new_n466_, new_n464_ );
nand g0125 ( new_n468_, new_n462_, N135 );
nand g0126 ( new_n469_, new_n468_, keyIn_0_72 );
not g0127 ( new_n470_, new_n469_ );
nor g0128 ( new_n471_, new_n468_, keyIn_0_72 );
nor g0129 ( new_n472_, new_n470_, new_n471_ );
nor g0130 ( new_n473_, new_n467_, new_n472_ );
not g0131 ( new_n474_, new_n473_ );
nand g0132 ( new_n475_, new_n474_, new_n414_ );
not g0133 ( new_n476_, new_n475_ );
nor g0134 ( new_n477_, new_n474_, new_n414_ );
nor g0135 ( new_n478_, new_n476_, new_n477_ );
not g0136 ( new_n479_, keyIn_0_94 );
not g0137 ( new_n480_, keyIn_0_71 );
not g0138 ( new_n481_, keyIn_0_52 );
not g0139 ( new_n482_, keyIn_0_15 );
nor g0140 ( new_n483_, N91, N96 );
nand g0141 ( new_n484_, N91, N96 );
not g0142 ( new_n485_, new_n484_ );
nor g0143 ( new_n486_, new_n485_, new_n483_ );
nor g0144 ( new_n487_, new_n486_, new_n482_ );
nand g0145 ( new_n488_, new_n486_, new_n482_ );
not g0146 ( new_n489_, new_n488_ );
nor g0147 ( new_n490_, new_n489_, new_n487_ );
nor g0148 ( new_n491_, new_n490_, keyIn_0_28 );
nand g0149 ( new_n492_, new_n490_, keyIn_0_28 );
not g0150 ( new_n493_, new_n492_ );
nor g0151 ( new_n494_, new_n493_, new_n491_ );
not g0152 ( new_n495_, N101 );
nor g0153 ( new_n496_, new_n495_, N106 );
not g0154 ( new_n497_, N106 );
nor g0155 ( new_n498_, new_n497_, N101 );
nor g0156 ( new_n499_, new_n496_, new_n498_ );
not g0157 ( new_n500_, new_n499_ );
nand g0158 ( new_n501_, new_n500_, keyIn_0_16 );
not g0159 ( new_n502_, new_n501_ );
nor g0160 ( new_n503_, new_n500_, keyIn_0_16 );
nor g0161 ( new_n504_, new_n502_, new_n503_ );
nor g0162 ( new_n505_, new_n504_, keyIn_0_29 );
nand g0163 ( new_n506_, new_n504_, keyIn_0_29 );
not g0164 ( new_n507_, new_n506_ );
nor g0165 ( new_n508_, new_n507_, new_n505_ );
nor g0166 ( new_n509_, new_n508_, new_n494_ );
not g0167 ( new_n510_, new_n509_ );
nor g0168 ( new_n511_, new_n510_, keyIn_0_42 );
nor g0169 ( new_n512_, new_n504_, new_n490_ );
not g0170 ( new_n513_, new_n512_ );
nand g0171 ( new_n514_, new_n513_, keyIn_0_30 );
not g0172 ( new_n515_, keyIn_0_30 );
nand g0173 ( new_n516_, new_n512_, new_n515_ );
nand g0174 ( new_n517_, new_n514_, new_n516_ );
nand g0175 ( new_n518_, new_n510_, keyIn_0_42 );
nand g0176 ( new_n519_, new_n518_, new_n517_ );
nor g0177 ( new_n520_, new_n519_, new_n511_ );
nor g0178 ( new_n521_, new_n520_, new_n481_ );
nand g0179 ( new_n522_, new_n520_, new_n481_ );
not g0180 ( new_n523_, new_n522_ );
nor g0181 ( new_n524_, new_n523_, new_n521_ );
not g0182 ( new_n525_, new_n524_ );
nor g0183 ( new_n526_, new_n525_, N130 );
nor g0184 ( new_n527_, new_n526_, new_n480_ );
nand g0185 ( new_n528_, new_n526_, new_n480_ );
not g0186 ( new_n529_, new_n528_ );
nor g0187 ( new_n530_, new_n529_, new_n527_ );
not g0188 ( new_n531_, keyIn_0_70 );
not g0189 ( new_n532_, N130 );
nor g0190 ( new_n533_, new_n524_, new_n532_ );
not g0191 ( new_n534_, new_n533_ );
nand g0192 ( new_n535_, new_n534_, new_n531_ );
not g0193 ( new_n536_, new_n535_ );
nor g0194 ( new_n537_, new_n534_, new_n531_ );
nor g0195 ( new_n538_, new_n536_, new_n537_ );
nor g0196 ( new_n539_, new_n538_, new_n530_ );
not g0197 ( new_n540_, new_n539_ );
nand g0198 ( new_n541_, new_n540_, new_n479_ );
not g0199 ( new_n542_, new_n541_ );
nor g0200 ( new_n543_, new_n540_, new_n479_ );
nor g0201 ( new_n544_, new_n542_, new_n543_ );
not g0202 ( new_n545_, new_n544_ );
nor g0203 ( new_n546_, new_n478_, new_n545_ );
not g0204 ( new_n547_, new_n546_ );
nand g0205 ( new_n548_, new_n547_, keyIn_0_106 );
not g0206 ( new_n549_, new_n548_ );
nand g0207 ( new_n550_, new_n478_, new_n545_ );
not g0208 ( new_n551_, new_n550_ );
nor g0209 ( new_n552_, new_n551_, keyIn_0_116 );
nor g0210 ( new_n553_, new_n549_, new_n552_ );
nor g0211 ( new_n554_, new_n547_, keyIn_0_106 );
nand g0212 ( new_n555_, new_n551_, keyIn_0_116 );
not g0213 ( new_n556_, new_n555_ );
nor g0214 ( new_n557_, new_n556_, new_n554_ );
nand g0215 ( new_n558_, new_n553_, new_n557_ );
not g0216 ( new_n559_, new_n558_ );
nand g0217 ( new_n560_, new_n559_, new_n413_ );
nand g0218 ( new_n561_, new_n558_, keyIn_0_139 );
nand g0219 ( N767, new_n560_, new_n561_ );
not g0220 ( new_n563_, keyIn_0_104 );
not g0221 ( new_n564_, keyIn_0_91 );
not g0222 ( new_n565_, keyIn_0_68 );
not g0223 ( new_n566_, keyIn_0_35 );
nand g0224 ( new_n567_, N159, N165 );
not g0225 ( new_n568_, new_n567_ );
nor g0226 ( new_n569_, N159, N165 );
nor g0227 ( new_n570_, new_n568_, new_n569_ );
not g0228 ( new_n571_, new_n570_ );
nor g0229 ( new_n572_, new_n571_, keyIn_0_21 );
nand g0230 ( new_n573_, new_n571_, keyIn_0_21 );
not g0231 ( new_n574_, new_n573_ );
nor g0232 ( new_n575_, new_n574_, new_n572_ );
nor g0233 ( new_n576_, new_n575_, new_n566_ );
not g0234 ( new_n577_, new_n575_ );
nor g0235 ( new_n578_, new_n577_, keyIn_0_35 );
nor g0236 ( new_n579_, new_n578_, new_n576_ );
not g0237 ( new_n580_, N171 );
nor g0238 ( new_n581_, new_n580_, N177 );
not g0239 ( new_n582_, N177 );
nor g0240 ( new_n583_, new_n582_, N171 );
nor g0241 ( new_n584_, new_n581_, new_n583_ );
not g0242 ( new_n585_, new_n584_ );
nand g0243 ( new_n586_, new_n585_, keyIn_0_22 );
not g0244 ( new_n587_, new_n586_ );
nor g0245 ( new_n588_, new_n585_, keyIn_0_22 );
nor g0246 ( new_n589_, new_n587_, new_n588_ );
not g0247 ( new_n590_, new_n589_ );
nor g0248 ( new_n591_, new_n590_, keyIn_0_36 );
nand g0249 ( new_n592_, new_n590_, keyIn_0_36 );
not g0250 ( new_n593_, new_n592_ );
nor g0251 ( new_n594_, new_n593_, new_n591_ );
nor g0252 ( new_n595_, new_n594_, new_n579_ );
not g0253 ( new_n596_, new_n595_ );
nand g0254 ( new_n597_, new_n596_, keyIn_0_49 );
not g0255 ( new_n598_, new_n597_ );
nor g0256 ( new_n599_, new_n596_, keyIn_0_49 );
nor g0257 ( new_n600_, new_n598_, new_n599_ );
nor g0258 ( new_n601_, new_n590_, new_n577_ );
nor g0259 ( new_n602_, new_n601_, keyIn_0_37 );
nand g0260 ( new_n603_, new_n601_, keyIn_0_37 );
not g0261 ( new_n604_, new_n603_ );
nor g0262 ( new_n605_, new_n604_, new_n602_ );
nor g0263 ( new_n606_, new_n600_, new_n605_ );
nor g0264 ( new_n607_, new_n606_, new_n565_ );
nand g0265 ( new_n608_, new_n606_, new_n565_ );
not g0266 ( new_n609_, new_n608_ );
nor g0267 ( new_n610_, new_n609_, new_n607_ );
not g0268 ( new_n611_, new_n610_ );
nor g0269 ( new_n612_, new_n611_, N130 );
nor g0270 ( new_n613_, new_n612_, new_n564_ );
nand g0271 ( new_n614_, new_n612_, new_n564_ );
not g0272 ( new_n615_, new_n614_ );
nor g0273 ( new_n616_, new_n615_, new_n613_ );
nor g0274 ( new_n617_, new_n610_, new_n532_ );
not g0275 ( new_n618_, new_n617_ );
nand g0276 ( new_n619_, new_n618_, keyIn_0_90 );
not g0277 ( new_n620_, new_n619_ );
nor g0278 ( new_n621_, new_n618_, keyIn_0_90 );
nor g0279 ( new_n622_, new_n620_, new_n621_ );
nor g0280 ( new_n623_, new_n622_, new_n616_ );
not g0281 ( new_n624_, new_n623_ );
nand g0282 ( new_n625_, new_n624_, new_n563_ );
not g0283 ( new_n626_, new_n625_ );
nor g0284 ( new_n627_, new_n624_, new_n563_ );
nor g0285 ( new_n628_, new_n626_, new_n627_ );
not g0286 ( new_n629_, new_n628_ );
not g0287 ( new_n630_, keyIn_0_92 );
not g0288 ( new_n631_, N207 );
not g0289 ( new_n632_, N195 );
nor g0290 ( new_n633_, new_n632_, N201 );
not g0291 ( new_n634_, N201 );
nor g0292 ( new_n635_, new_n634_, N195 );
nor g0293 ( new_n636_, new_n633_, new_n635_ );
not g0294 ( new_n637_, new_n636_ );
nand g0295 ( new_n638_, new_n637_, keyIn_0_24 );
not g0296 ( new_n639_, new_n638_ );
nor g0297 ( new_n640_, new_n637_, keyIn_0_24 );
nor g0298 ( new_n641_, new_n639_, new_n640_ );
not g0299 ( new_n642_, new_n641_ );
nand g0300 ( new_n643_, new_n642_, keyIn_0_39 );
not g0301 ( new_n644_, keyIn_0_39 );
nand g0302 ( new_n645_, new_n641_, new_n644_ );
nand g0303 ( new_n646_, new_n643_, new_n645_ );
not g0304 ( new_n647_, N183 );
nor g0305 ( new_n648_, new_n647_, N189 );
not g0306 ( new_n649_, N189 );
nor g0307 ( new_n650_, new_n649_, N183 );
nor g0308 ( new_n651_, new_n648_, new_n650_ );
not g0309 ( new_n652_, new_n651_ );
nand g0310 ( new_n653_, new_n652_, keyIn_0_23 );
not g0311 ( new_n654_, new_n653_ );
nor g0312 ( new_n655_, new_n652_, keyIn_0_23 );
nor g0313 ( new_n656_, new_n654_, new_n655_ );
not g0314 ( new_n657_, new_n656_ );
nand g0315 ( new_n658_, new_n657_, keyIn_0_38 );
not g0316 ( new_n659_, keyIn_0_38 );
nand g0317 ( new_n660_, new_n656_, new_n659_ );
nand g0318 ( new_n661_, new_n658_, new_n660_ );
nand g0319 ( new_n662_, new_n646_, new_n661_ );
nor g0320 ( new_n663_, new_n662_, keyIn_0_50 );
nor g0321 ( new_n664_, new_n641_, new_n656_ );
not g0322 ( new_n665_, new_n664_ );
nand g0323 ( new_n666_, new_n665_, keyIn_0_40 );
not g0324 ( new_n667_, keyIn_0_40 );
nand g0325 ( new_n668_, new_n664_, new_n667_ );
nand g0326 ( new_n669_, new_n666_, new_n668_ );
nand g0327 ( new_n670_, new_n662_, keyIn_0_50 );
nand g0328 ( new_n671_, new_n670_, new_n669_ );
nor g0329 ( new_n672_, new_n671_, new_n663_ );
nor g0330 ( new_n673_, new_n672_, keyIn_0_69 );
nand g0331 ( new_n674_, new_n672_, keyIn_0_69 );
not g0332 ( new_n675_, new_n674_ );
nor g0333 ( new_n676_, new_n675_, new_n673_ );
not g0334 ( new_n677_, new_n676_ );
nor g0335 ( new_n678_, new_n677_, new_n631_ );
nor g0336 ( new_n679_, new_n678_, new_n630_ );
nand g0337 ( new_n680_, new_n678_, new_n630_ );
not g0338 ( new_n681_, new_n680_ );
nor g0339 ( new_n682_, new_n681_, new_n679_ );
not g0340 ( new_n683_, keyIn_0_93 );
nor g0341 ( new_n684_, new_n676_, N207 );
not g0342 ( new_n685_, new_n684_ );
nand g0343 ( new_n686_, new_n685_, new_n683_ );
not g0344 ( new_n687_, new_n686_ );
nor g0345 ( new_n688_, new_n685_, new_n683_ );
nor g0346 ( new_n689_, new_n687_, new_n688_ );
nor g0347 ( new_n690_, new_n689_, new_n682_ );
not g0348 ( new_n691_, new_n690_ );
nand g0349 ( new_n692_, new_n691_, keyIn_0_105 );
not g0350 ( new_n693_, new_n692_ );
nor g0351 ( new_n694_, new_n691_, keyIn_0_105 );
nor g0352 ( new_n695_, new_n693_, new_n694_ );
not g0353 ( new_n696_, new_n695_ );
nor g0354 ( new_n697_, new_n629_, new_n696_ );
not g0355 ( new_n698_, new_n697_ );
nand g0356 ( new_n699_, new_n698_, keyIn_0_115 );
not g0357 ( new_n700_, keyIn_0_115 );
nand g0358 ( new_n701_, new_n697_, new_n700_ );
nand g0359 ( new_n702_, new_n699_, new_n701_ );
nor g0360 ( new_n703_, new_n628_, new_n695_ );
not g0361 ( new_n704_, new_n703_ );
nand g0362 ( new_n705_, new_n704_, keyIn_0_117 );
not g0363 ( new_n706_, keyIn_0_117 );
nand g0364 ( new_n707_, new_n703_, new_n706_ );
nand g0365 ( new_n708_, new_n705_, new_n707_ );
nand g0366 ( new_n709_, new_n702_, new_n708_ );
nand g0367 ( new_n710_, new_n709_, keyIn_0_140 );
not g0368 ( new_n711_, keyIn_0_140 );
not g0369 ( new_n712_, new_n709_ );
nand g0370 ( new_n713_, new_n712_, new_n711_ );
nand g0371 ( N768, new_n713_, new_n710_ );
not g0372 ( new_n715_, keyIn_0_210 );
not g0373 ( new_n716_, keyIn_0_202 );
not g0374 ( new_n717_, keyIn_0_184 );
not g0375 ( new_n718_, keyIn_0_103 );
not g0376 ( new_n719_, keyIn_0_63 );
not g0377 ( new_n720_, keyIn_0_9 );
nor g0378 ( new_n721_, N447, new_n720_ );
nand g0379 ( new_n722_, new_n389_, keyIn_0_0 );
nand g0380 ( new_n723_, new_n386_, new_n384_ );
nand g0381 ( new_n724_, new_n722_, new_n723_ );
nor g0382 ( new_n725_, new_n724_, keyIn_0_9 );
nor g0383 ( new_n726_, new_n721_, new_n725_ );
nor g0384 ( new_n727_, new_n726_, keyIn_0_26 );
not g0385 ( new_n728_, keyIn_0_26 );
nand g0386 ( new_n729_, new_n724_, keyIn_0_9 );
nand g0387 ( new_n730_, N447, new_n720_ );
nand g0388 ( new_n731_, new_n730_, new_n729_ );
nor g0389 ( new_n732_, new_n731_, new_n728_ );
nor g0390 ( new_n733_, new_n727_, new_n732_ );
not g0391 ( new_n734_, keyIn_0_5 );
nand g0392 ( new_n735_, N59, N156 );
nand g0393 ( new_n736_, new_n735_, new_n734_ );
not g0394 ( new_n737_, new_n736_ );
nor g0395 ( new_n738_, new_n735_, new_n734_ );
nor g0396 ( new_n739_, new_n737_, new_n738_ );
not g0397 ( new_n740_, new_n739_ );
nor g0398 ( new_n741_, new_n733_, new_n740_ );
nand g0399 ( new_n742_, new_n741_, N17 );
nand g0400 ( new_n743_, new_n742_, keyIn_0_48 );
not g0401 ( new_n744_, keyIn_0_48 );
nand g0402 ( new_n745_, new_n731_, new_n728_ );
nand g0403 ( new_n746_, new_n726_, keyIn_0_26 );
nand g0404 ( new_n747_, new_n746_, new_n745_ );
nand g0405 ( new_n748_, new_n747_, new_n739_ );
nor g0406 ( new_n749_, new_n748_, new_n353_ );
nand g0407 ( new_n750_, new_n749_, new_n744_ );
nand g0408 ( new_n751_, new_n743_, new_n750_ );
nand g0409 ( new_n752_, new_n751_, N1 );
nand g0410 ( new_n753_, new_n752_, new_n719_ );
nor g0411 ( new_n754_, new_n752_, new_n719_ );
not g0412 ( new_n755_, new_n754_ );
nand g0413 ( new_n756_, new_n755_, new_n753_ );
nand g0414 ( new_n757_, new_n756_, N153 );
nand g0415 ( new_n758_, new_n757_, keyIn_0_88 );
not g0416 ( new_n759_, keyIn_0_88 );
not g0417 ( new_n760_, N153 );
not g0418 ( new_n761_, new_n753_ );
nor g0419 ( new_n762_, new_n761_, new_n754_ );
nor g0420 ( new_n763_, new_n762_, new_n760_ );
nand g0421 ( new_n764_, new_n763_, new_n759_ );
nand g0422 ( new_n765_, new_n764_, new_n758_ );
not g0423 ( new_n766_, keyIn_0_89 );
not g0424 ( new_n767_, keyIn_0_54 );
nand g0425 ( new_n768_, N17, N42 );
nand g0426 ( new_n769_, new_n768_, keyIn_0_7 );
nor g0427 ( new_n770_, N17, N42 );
nor g0428 ( new_n771_, new_n770_, keyIn_0_6 );
not g0429 ( new_n772_, new_n771_ );
nand g0430 ( new_n773_, new_n772_, new_n769_ );
nor g0431 ( new_n774_, new_n768_, keyIn_0_7 );
not g0432 ( new_n775_, new_n774_ );
nand g0433 ( new_n776_, new_n770_, keyIn_0_6 );
nand g0434 ( new_n777_, new_n775_, new_n776_ );
nor g0435 ( new_n778_, new_n773_, new_n777_ );
nor g0436 ( new_n779_, new_n778_, keyIn_0_20 );
not g0437 ( new_n780_, new_n735_ );
nand g0438 ( new_n781_, new_n778_, keyIn_0_20 );
nand g0439 ( new_n782_, new_n781_, new_n780_ );
nor g0440 ( new_n783_, new_n782_, new_n779_ );
nand g0441 ( new_n784_, new_n747_, new_n783_ );
nor g0442 ( new_n785_, new_n784_, keyIn_0_47 );
nand g0443 ( new_n786_, new_n784_, keyIn_0_47 );
nand g0444 ( new_n787_, N17, N51 );
nor g0445 ( new_n788_, new_n354_, new_n787_ );
nor g0446 ( new_n789_, new_n788_, keyIn_0_1 );
nand g0447 ( new_n790_, new_n788_, keyIn_0_1 );
not g0448 ( new_n791_, new_n790_ );
nor g0449 ( new_n792_, new_n791_, new_n789_ );
not g0450 ( new_n793_, new_n792_ );
nand g0451 ( new_n794_, new_n793_, keyIn_0_10 );
not g0452 ( new_n795_, keyIn_0_10 );
nand g0453 ( new_n796_, new_n792_, new_n795_ );
nand g0454 ( new_n797_, new_n794_, new_n796_ );
nor g0455 ( new_n798_, new_n368_, new_n349_ );
nor g0456 ( new_n799_, new_n798_, keyIn_0_3 );
nand g0457 ( new_n800_, new_n798_, keyIn_0_3 );
not g0458 ( new_n801_, new_n800_ );
nor g0459 ( new_n802_, new_n801_, new_n799_ );
not g0460 ( new_n803_, new_n802_ );
nand g0461 ( new_n804_, new_n803_, keyIn_0_14 );
not g0462 ( new_n805_, keyIn_0_14 );
nand g0463 ( new_n806_, new_n802_, new_n805_ );
nand g0464 ( new_n807_, new_n804_, new_n806_ );
nand g0465 ( new_n808_, new_n797_, new_n807_ );
nand g0466 ( new_n809_, new_n808_, keyIn_0_34 );
not g0467 ( new_n810_, keyIn_0_34 );
not g0468 ( new_n811_, new_n808_ );
nand g0469 ( new_n812_, new_n811_, new_n810_ );
nand g0470 ( new_n813_, new_n812_, new_n809_ );
nand g0471 ( new_n814_, new_n813_, new_n786_ );
nor g0472 ( new_n815_, new_n814_, new_n785_ );
nor g0473 ( new_n816_, new_n815_, new_n767_ );
nand g0474 ( new_n817_, new_n815_, new_n767_ );
not g0475 ( new_n818_, new_n817_ );
nor g0476 ( new_n819_, new_n818_, new_n816_ );
nand g0477 ( new_n820_, new_n819_, N126 );
nand g0478 ( new_n821_, new_n820_, new_n766_ );
nor g0479 ( new_n822_, new_n820_, new_n766_ );
not g0480 ( new_n823_, new_n822_ );
nand g0481 ( new_n824_, new_n823_, new_n821_ );
nand g0482 ( new_n825_, new_n765_, new_n824_ );
nor g0483 ( new_n826_, new_n825_, new_n718_ );
not g0484 ( new_n827_, new_n826_ );
not g0485 ( new_n828_, keyIn_0_67 );
nand g0486 ( new_n829_, N29, N75 );
nor g0487 ( new_n830_, new_n829_, new_n346_ );
nor g0488 ( new_n831_, new_n830_, keyIn_0_2 );
nand g0489 ( new_n832_, new_n830_, keyIn_0_2 );
not g0490 ( new_n833_, new_n832_ );
nor g0491 ( new_n834_, new_n833_, new_n831_ );
nor g0492 ( new_n835_, new_n733_, new_n834_ );
not g0493 ( new_n836_, new_n835_ );
nor g0494 ( new_n837_, new_n836_, new_n392_ );
not g0495 ( new_n838_, new_n837_ );
nor g0496 ( new_n839_, new_n838_, keyIn_0_46 );
not g0497 ( new_n840_, keyIn_0_19 );
nand g0498 ( new_n841_, keyIn_0_4, N268 );
not g0499 ( new_n842_, new_n841_ );
nor g0500 ( new_n843_, keyIn_0_4, N268 );
nor g0501 ( new_n844_, new_n842_, new_n843_ );
not g0502 ( new_n845_, new_n844_ );
nor g0503 ( new_n846_, new_n845_, new_n840_ );
nor g0504 ( new_n847_, new_n844_, keyIn_0_19 );
nor g0505 ( new_n848_, new_n846_, new_n847_ );
nand g0506 ( new_n849_, new_n838_, keyIn_0_46 );
nand g0507 ( new_n850_, new_n849_, new_n848_ );
nor g0508 ( new_n851_, new_n850_, new_n839_ );
nand g0509 ( new_n852_, new_n851_, new_n828_ );
not g0510 ( new_n853_, new_n851_ );
nand g0511 ( new_n854_, new_n853_, keyIn_0_67 );
nand g0512 ( new_n855_, new_n854_, new_n852_ );
nand g0513 ( new_n856_, new_n825_, new_n718_ );
nand g0514 ( new_n857_, new_n856_, new_n855_ );
not g0515 ( new_n858_, new_n857_ );
nand g0516 ( new_n859_, new_n858_, new_n827_ );
nand g0517 ( new_n860_, new_n859_, keyIn_0_114 );
not g0518 ( new_n861_, keyIn_0_114 );
nor g0519 ( new_n862_, new_n857_, new_n826_ );
nand g0520 ( new_n863_, new_n862_, new_n861_ );
nand g0521 ( new_n864_, new_n860_, new_n863_ );
nand g0522 ( new_n865_, new_n864_, new_n634_ );
nand g0523 ( new_n866_, new_n865_, keyIn_0_138 );
nor g0524 ( new_n867_, new_n865_, keyIn_0_138 );
not g0525 ( new_n868_, new_n867_ );
nand g0526 ( new_n869_, new_n868_, new_n866_ );
not g0527 ( new_n870_, keyIn_0_137 );
nor g0528 ( new_n871_, new_n864_, new_n634_ );
nor g0529 ( new_n872_, new_n871_, new_n870_ );
nor g0530 ( new_n873_, new_n862_, new_n861_ );
not g0531 ( new_n874_, new_n863_ );
nor g0532 ( new_n875_, new_n874_, new_n873_ );
nand g0533 ( new_n876_, new_n875_, N201 );
nor g0534 ( new_n877_, new_n876_, keyIn_0_137 );
nor g0535 ( new_n878_, new_n877_, new_n872_ );
nor g0536 ( new_n879_, new_n869_, new_n878_ );
nor g0537 ( new_n880_, new_n879_, keyIn_0_163 );
nand g0538 ( new_n881_, new_n879_, keyIn_0_163 );
not g0539 ( new_n882_, new_n881_ );
nor g0540 ( new_n883_, new_n882_, new_n880_ );
not g0541 ( new_n884_, new_n883_ );
nor g0542 ( new_n885_, new_n884_, N261 );
nor g0543 ( new_n886_, new_n885_, new_n717_ );
nand g0544 ( new_n887_, new_n885_, new_n717_ );
not g0545 ( new_n888_, new_n887_ );
nor g0546 ( new_n889_, new_n888_, new_n886_ );
not g0547 ( new_n890_, keyIn_0_185 );
not g0548 ( new_n891_, N261 );
nor g0549 ( new_n892_, new_n883_, new_n891_ );
not g0550 ( new_n893_, new_n892_ );
nand g0551 ( new_n894_, new_n893_, new_n890_ );
not g0552 ( new_n895_, new_n894_ );
nor g0553 ( new_n896_, new_n893_, new_n890_ );
nor g0554 ( new_n897_, new_n895_, new_n896_ );
nor g0555 ( new_n898_, new_n897_, new_n889_ );
not g0556 ( new_n899_, new_n898_ );
nor g0557 ( new_n900_, new_n899_, new_n716_ );
nand g0558 ( new_n901_, new_n899_, new_n716_ );
nand g0559 ( new_n902_, new_n901_, N219 );
nor g0560 ( new_n903_, new_n902_, new_n900_ );
nor g0561 ( new_n904_, new_n903_, new_n715_ );
nand g0562 ( new_n905_, new_n903_, new_n715_ );
not g0563 ( new_n906_, new_n905_ );
nor g0564 ( new_n907_, new_n906_, new_n904_ );
nand g0565 ( new_n908_, N121, N210 );
not g0566 ( new_n909_, new_n908_ );
nor g0567 ( new_n910_, new_n907_, new_n909_ );
not g0568 ( new_n911_, new_n910_ );
nor g0569 ( new_n912_, new_n911_, keyIn_0_216 );
nand g0570 ( new_n913_, new_n911_, keyIn_0_216 );
not g0571 ( new_n914_, keyIn_0_203 );
nand g0572 ( new_n915_, new_n884_, N228 );
not g0573 ( new_n916_, keyIn_0_162 );
nand g0574 ( new_n917_, new_n876_, keyIn_0_137 );
nand g0575 ( new_n918_, new_n871_, new_n870_ );
nand g0576 ( new_n919_, new_n917_, new_n918_ );
nand g0577 ( new_n920_, new_n919_, new_n916_ );
nand g0578 ( new_n921_, new_n878_, keyIn_0_162 );
nand g0579 ( new_n922_, new_n921_, new_n920_ );
nand g0580 ( new_n923_, new_n922_, N237 );
nand g0581 ( new_n924_, new_n915_, new_n923_ );
nor g0582 ( new_n925_, new_n924_, new_n914_ );
nand g0583 ( new_n926_, new_n924_, new_n914_ );
not g0584 ( new_n927_, keyIn_0_51 );
not g0585 ( new_n928_, keyIn_0_41 );
not g0586 ( new_n929_, N73 );
nand g0587 ( new_n930_, N42, N72 );
nor g0588 ( new_n931_, new_n402_, new_n930_ );
nand g0589 ( new_n932_, new_n393_, new_n931_ );
not g0590 ( new_n933_, new_n932_ );
nor g0591 ( new_n934_, new_n933_, keyIn_0_11 );
nand g0592 ( new_n935_, new_n933_, keyIn_0_11 );
not g0593 ( new_n936_, new_n935_ );
nor g0594 ( new_n937_, new_n936_, new_n934_ );
nor g0595 ( new_n938_, new_n937_, new_n929_ );
not g0596 ( new_n939_, new_n938_ );
nand g0597 ( new_n940_, new_n939_, keyIn_0_27 );
not g0598 ( new_n941_, new_n940_ );
nor g0599 ( new_n942_, new_n939_, keyIn_0_27 );
nor g0600 ( new_n943_, new_n941_, new_n942_ );
nor g0601 ( new_n944_, new_n943_, new_n928_ );
nand g0602 ( new_n945_, new_n943_, new_n928_ );
not g0603 ( new_n946_, new_n945_ );
nor g0604 ( new_n947_, new_n946_, new_n944_ );
nor g0605 ( new_n948_, new_n947_, new_n927_ );
nand g0606 ( new_n949_, new_n947_, new_n927_ );
not g0607 ( new_n950_, new_n949_ );
nor g0608 ( new_n951_, new_n950_, new_n948_ );
not g0609 ( new_n952_, new_n951_ );
nand g0610 ( new_n953_, new_n952_, N201 );
nand g0611 ( new_n954_, N255, N267 );
not g0612 ( new_n955_, new_n954_ );
not g0613 ( new_n956_, N246 );
nor g0614 ( new_n957_, new_n864_, new_n956_ );
nor g0615 ( new_n958_, new_n957_, new_n955_ );
not g0616 ( new_n959_, new_n958_ );
nand g0617 ( new_n960_, new_n959_, keyIn_0_164 );
not g0618 ( new_n961_, keyIn_0_164 );
nand g0619 ( new_n962_, new_n958_, new_n961_ );
nand g0620 ( new_n963_, new_n960_, new_n962_ );
nand g0621 ( new_n964_, new_n963_, new_n953_ );
not g0622 ( new_n965_, new_n964_ );
nand g0623 ( new_n966_, new_n926_, new_n965_ );
nor g0624 ( new_n967_, new_n966_, new_n925_ );
nand g0625 ( new_n968_, new_n913_, new_n967_ );
nor g0626 ( new_n969_, new_n968_, new_n912_ );
not g0627 ( new_n970_, new_n969_ );
nand g0628 ( new_n971_, new_n970_, keyIn_0_222 );
not g0629 ( new_n972_, keyIn_0_222 );
nand g0630 ( new_n973_, new_n969_, new_n972_ );
nand g0631 ( N850, new_n971_, new_n973_ );
not g0632 ( new_n975_, keyIn_0_240 );
not g0633 ( new_n976_, keyIn_0_219 );
not g0634 ( new_n977_, N219 );
not g0635 ( new_n978_, keyIn_0_131 );
not g0636 ( new_n979_, keyIn_0_111 );
not g0637 ( new_n980_, keyIn_0_100 );
not g0638 ( new_n981_, new_n819_ );
nor g0639 ( new_n982_, new_n981_, new_n430_ );
nor g0640 ( new_n983_, new_n982_, keyIn_0_83 );
nand g0641 ( new_n984_, new_n982_, keyIn_0_83 );
not g0642 ( new_n985_, new_n984_ );
nor g0643 ( new_n986_, new_n985_, new_n983_ );
not g0644 ( new_n987_, N143 );
nor g0645 ( new_n988_, new_n762_, new_n987_ );
nor g0646 ( new_n989_, new_n988_, keyIn_0_82 );
nand g0647 ( new_n990_, new_n988_, keyIn_0_82 );
not g0648 ( new_n991_, new_n990_ );
nor g0649 ( new_n992_, new_n991_, new_n989_ );
nor g0650 ( new_n993_, new_n992_, new_n986_ );
not g0651 ( new_n994_, new_n993_ );
nand g0652 ( new_n995_, new_n994_, new_n980_ );
not g0653 ( new_n996_, new_n995_ );
nor g0654 ( new_n997_, new_n994_, new_n980_ );
nor g0655 ( new_n998_, new_n996_, new_n997_ );
nor g0656 ( new_n999_, new_n853_, keyIn_0_64 );
nand g0657 ( new_n1000_, new_n853_, keyIn_0_64 );
not g0658 ( new_n1001_, new_n1000_ );
nor g0659 ( new_n1002_, new_n1001_, new_n999_ );
nor g0660 ( new_n1003_, new_n998_, new_n1002_ );
nor g0661 ( new_n1004_, new_n1003_, new_n979_ );
nand g0662 ( new_n1005_, new_n1003_, new_n979_ );
not g0663 ( new_n1006_, new_n1005_ );
nor g0664 ( new_n1007_, new_n1006_, new_n1004_ );
not g0665 ( new_n1008_, new_n1007_ );
nor g0666 ( new_n1009_, new_n1008_, N183 );
nor g0667 ( new_n1010_, new_n1009_, new_n978_ );
nand g0668 ( new_n1011_, new_n1009_, new_n978_ );
not g0669 ( new_n1012_, new_n1011_ );
nor g0670 ( new_n1013_, new_n1012_, new_n1010_ );
not g0671 ( new_n1014_, new_n1013_ );
nor g0672 ( new_n1015_, new_n1007_, new_n647_ );
not g0673 ( new_n1016_, new_n1015_ );
nand g0674 ( new_n1017_, new_n1016_, keyIn_0_130 );
not g0675 ( new_n1018_, new_n1017_ );
nor g0676 ( new_n1019_, new_n1016_, keyIn_0_130 );
nor g0677 ( new_n1020_, new_n1018_, new_n1019_ );
nor g0678 ( new_n1021_, new_n1014_, new_n1020_ );
nor g0679 ( new_n1022_, new_n1021_, keyIn_0_154 );
nand g0680 ( new_n1023_, new_n1021_, keyIn_0_154 );
not g0681 ( new_n1024_, new_n1023_ );
nor g0682 ( new_n1025_, new_n1024_, new_n1022_ );
not g0683 ( new_n1026_, keyIn_0_196 );
not g0684 ( new_n1027_, keyIn_0_187 );
not g0685 ( new_n1028_, keyIn_0_112 );
nand g0686 ( new_n1029_, new_n756_, N146 );
nand g0687 ( new_n1030_, new_n1029_, keyIn_0_84 );
not g0688 ( new_n1031_, keyIn_0_84 );
not g0689 ( new_n1032_, N146 );
nor g0690 ( new_n1033_, new_n762_, new_n1032_ );
nand g0691 ( new_n1034_, new_n1033_, new_n1031_ );
nand g0692 ( new_n1035_, new_n1034_, new_n1030_ );
not g0693 ( new_n1036_, keyIn_0_85 );
nand g0694 ( new_n1037_, new_n819_, N116 );
nand g0695 ( new_n1038_, new_n1037_, new_n1036_ );
nor g0696 ( new_n1039_, new_n1037_, new_n1036_ );
not g0697 ( new_n1040_, new_n1039_ );
nand g0698 ( new_n1041_, new_n1040_, new_n1038_ );
nand g0699 ( new_n1042_, new_n1035_, new_n1041_ );
nor g0700 ( new_n1043_, new_n1042_, keyIn_0_101 );
not g0701 ( new_n1044_, new_n1043_ );
not g0702 ( new_n1045_, keyIn_0_65 );
nand g0703 ( new_n1046_, new_n851_, new_n1045_ );
nand g0704 ( new_n1047_, new_n853_, keyIn_0_65 );
nand g0705 ( new_n1048_, new_n1047_, new_n1046_ );
nand g0706 ( new_n1049_, new_n1042_, keyIn_0_101 );
nand g0707 ( new_n1050_, new_n1049_, new_n1048_ );
not g0708 ( new_n1051_, new_n1050_ );
nand g0709 ( new_n1052_, new_n1051_, new_n1044_ );
nand g0710 ( new_n1053_, new_n1052_, new_n1028_ );
nor g0711 ( new_n1054_, new_n1050_, new_n1043_ );
nand g0712 ( new_n1055_, new_n1054_, keyIn_0_112 );
nand g0713 ( new_n1056_, new_n1053_, new_n1055_ );
nor g0714 ( new_n1057_, new_n1056_, N189 );
nor g0715 ( new_n1058_, new_n1057_, keyIn_0_134 );
not g0716 ( new_n1059_, keyIn_0_134 );
nor g0717 ( new_n1060_, new_n1054_, keyIn_0_112 );
not g0718 ( new_n1061_, new_n1055_ );
nor g0719 ( new_n1062_, new_n1061_, new_n1060_ );
nand g0720 ( new_n1063_, new_n1062_, new_n649_ );
nor g0721 ( new_n1064_, new_n1063_, new_n1059_ );
nor g0722 ( new_n1065_, new_n1064_, new_n1058_ );
not g0723 ( new_n1066_, keyIn_0_159 );
not g0724 ( new_n1067_, keyIn_0_113 );
not g0725 ( new_n1068_, keyIn_0_102 );
not g0726 ( new_n1069_, keyIn_0_86 );
nand g0727 ( new_n1070_, new_n756_, N149 );
nand g0728 ( new_n1071_, new_n1070_, new_n1069_ );
not g0729 ( new_n1072_, N149 );
nor g0730 ( new_n1073_, new_n762_, new_n1072_ );
nand g0731 ( new_n1074_, new_n1073_, keyIn_0_86 );
nand g0732 ( new_n1075_, new_n1074_, new_n1071_ );
not g0733 ( new_n1076_, keyIn_0_87 );
nand g0734 ( new_n1077_, new_n819_, N121 );
nand g0735 ( new_n1078_, new_n1077_, new_n1076_ );
nor g0736 ( new_n1079_, new_n1077_, new_n1076_ );
not g0737 ( new_n1080_, new_n1079_ );
nand g0738 ( new_n1081_, new_n1080_, new_n1078_ );
nand g0739 ( new_n1082_, new_n1075_, new_n1081_ );
nor g0740 ( new_n1083_, new_n1082_, new_n1068_ );
not g0741 ( new_n1084_, new_n1083_ );
nand g0742 ( new_n1085_, new_n1082_, new_n1068_ );
not g0743 ( new_n1086_, keyIn_0_66 );
nor g0744 ( new_n1087_, new_n853_, new_n1086_ );
nor g0745 ( new_n1088_, new_n851_, keyIn_0_66 );
nor g0746 ( new_n1089_, new_n1087_, new_n1088_ );
nand g0747 ( new_n1090_, new_n1085_, new_n1089_ );
not g0748 ( new_n1091_, new_n1090_ );
nand g0749 ( new_n1092_, new_n1091_, new_n1084_ );
nand g0750 ( new_n1093_, new_n1092_, new_n1067_ );
nor g0751 ( new_n1094_, new_n1090_, new_n1083_ );
nand g0752 ( new_n1095_, new_n1094_, keyIn_0_113 );
nand g0753 ( new_n1096_, new_n1093_, new_n1095_ );
nand g0754 ( new_n1097_, new_n1096_, N195 );
nand g0755 ( new_n1098_, new_n1097_, keyIn_0_135 );
not g0756 ( new_n1099_, new_n1098_ );
nor g0757 ( new_n1100_, new_n1097_, keyIn_0_135 );
nor g0758 ( new_n1101_, new_n1099_, new_n1100_ );
not g0759 ( new_n1102_, new_n1101_ );
nand g0760 ( new_n1103_, new_n1102_, new_n1066_ );
nand g0761 ( new_n1104_, new_n1101_, keyIn_0_159 );
nand g0762 ( new_n1105_, new_n1103_, new_n1104_ );
nand g0763 ( new_n1106_, new_n1105_, new_n1065_ );
nand g0764 ( new_n1107_, new_n1106_, new_n1027_ );
not g0765 ( new_n1108_, new_n1106_ );
nand g0766 ( new_n1109_, new_n1108_, keyIn_0_187 );
nand g0767 ( new_n1110_, new_n1109_, new_n1107_ );
nand g0768 ( new_n1111_, new_n1063_, new_n1059_ );
nand g0769 ( new_n1112_, new_n1057_, keyIn_0_134 );
nand g0770 ( new_n1113_, new_n1111_, new_n1112_ );
not g0771 ( new_n1114_, keyIn_0_136 );
nor g0772 ( new_n1115_, new_n1094_, keyIn_0_113 );
not g0773 ( new_n1116_, new_n1095_ );
nor g0774 ( new_n1117_, new_n1116_, new_n1115_ );
nand g0775 ( new_n1118_, new_n1117_, new_n632_ );
nand g0776 ( new_n1119_, new_n1118_, new_n1114_ );
nor g0777 ( new_n1120_, new_n1096_, N195 );
nand g0778 ( new_n1121_, new_n1120_, keyIn_0_136 );
nand g0779 ( new_n1122_, new_n1119_, new_n1121_ );
nor g0780 ( new_n1123_, new_n1113_, new_n1122_ );
nand g0781 ( new_n1124_, new_n922_, new_n1123_ );
nand g0782 ( new_n1125_, new_n1124_, keyIn_0_188 );
not g0783 ( new_n1126_, keyIn_0_167 );
nor g0784 ( new_n1127_, new_n869_, new_n891_ );
nand g0785 ( new_n1128_, new_n1127_, new_n1123_ );
nand g0786 ( new_n1129_, new_n1128_, new_n1126_ );
nor g0787 ( new_n1130_, new_n1120_, keyIn_0_136 );
nor g0788 ( new_n1131_, new_n1118_, new_n1114_ );
nor g0789 ( new_n1132_, new_n1131_, new_n1130_ );
nand g0790 ( new_n1133_, new_n1065_, new_n1132_ );
not g0791 ( new_n1134_, new_n866_ );
nor g0792 ( new_n1135_, new_n1134_, new_n867_ );
nand g0793 ( new_n1136_, new_n1135_, N261 );
nor g0794 ( new_n1137_, new_n1133_, new_n1136_ );
nand g0795 ( new_n1138_, new_n1137_, keyIn_0_167 );
nand g0796 ( new_n1139_, new_n1138_, new_n1129_ );
nand g0797 ( new_n1140_, new_n1139_, new_n1125_ );
not g0798 ( new_n1141_, keyIn_0_156 );
not g0799 ( new_n1142_, keyIn_0_133 );
nand g0800 ( new_n1143_, new_n1056_, N189 );
nand g0801 ( new_n1144_, new_n1143_, new_n1142_ );
not g0802 ( new_n1145_, new_n1143_ );
nand g0803 ( new_n1146_, new_n1145_, keyIn_0_133 );
nand g0804 ( new_n1147_, new_n1146_, new_n1144_ );
nand g0805 ( new_n1148_, new_n1147_, new_n1141_ );
not g0806 ( new_n1149_, new_n1144_ );
nor g0807 ( new_n1150_, new_n1143_, new_n1142_ );
nor g0808 ( new_n1151_, new_n1149_, new_n1150_ );
nand g0809 ( new_n1152_, new_n1151_, keyIn_0_156 );
nand g0810 ( new_n1153_, new_n1152_, new_n1148_ );
nand g0811 ( new_n1154_, new_n1153_, keyIn_0_177 );
not g0812 ( new_n1155_, keyIn_0_177 );
nor g0813 ( new_n1156_, new_n1151_, keyIn_0_156 );
nor g0814 ( new_n1157_, new_n1147_, new_n1141_ );
nor g0815 ( new_n1158_, new_n1156_, new_n1157_ );
nand g0816 ( new_n1159_, new_n1158_, new_n1155_ );
nand g0817 ( new_n1160_, new_n1159_, new_n1154_ );
not g0818 ( new_n1161_, keyIn_0_188 );
nor g0819 ( new_n1162_, new_n878_, keyIn_0_162 );
nor g0820 ( new_n1163_, new_n919_, new_n916_ );
nor g0821 ( new_n1164_, new_n1162_, new_n1163_ );
nor g0822 ( new_n1165_, new_n1164_, new_n1133_ );
nand g0823 ( new_n1166_, new_n1165_, new_n1161_ );
nand g0824 ( new_n1167_, new_n1166_, new_n1160_ );
nor g0825 ( new_n1168_, new_n1167_, new_n1140_ );
nand g0826 ( new_n1169_, new_n1168_, new_n1110_ );
nand g0827 ( new_n1170_, new_n1169_, new_n1026_ );
not g0828 ( new_n1171_, new_n1107_ );
nor g0829 ( new_n1172_, new_n1106_, new_n1027_ );
nor g0830 ( new_n1173_, new_n1171_, new_n1172_ );
not g0831 ( new_n1174_, new_n1125_ );
nor g0832 ( new_n1175_, new_n1137_, keyIn_0_167 );
nor g0833 ( new_n1176_, new_n1128_, new_n1126_ );
nor g0834 ( new_n1177_, new_n1175_, new_n1176_ );
nor g0835 ( new_n1178_, new_n1177_, new_n1174_ );
not g0836 ( new_n1179_, new_n1154_ );
nor g0837 ( new_n1180_, new_n1153_, keyIn_0_177 );
nor g0838 ( new_n1181_, new_n1179_, new_n1180_ );
nor g0839 ( new_n1182_, new_n1124_, keyIn_0_188 );
nor g0840 ( new_n1183_, new_n1181_, new_n1182_ );
nand g0841 ( new_n1184_, new_n1183_, new_n1178_ );
nor g0842 ( new_n1185_, new_n1184_, new_n1173_ );
nand g0843 ( new_n1186_, new_n1185_, keyIn_0_196 );
nand g0844 ( new_n1187_, new_n1186_, new_n1170_ );
nor g0845 ( new_n1188_, new_n1187_, new_n1025_ );
nor g0846 ( new_n1189_, new_n1188_, keyIn_0_205 );
nand g0847 ( new_n1190_, new_n1188_, keyIn_0_205 );
not g0848 ( new_n1191_, new_n1190_ );
nor g0849 ( new_n1192_, new_n1191_, new_n1189_ );
not g0850 ( new_n1193_, new_n1025_ );
not g0851 ( new_n1194_, new_n1170_ );
nor g0852 ( new_n1195_, new_n1169_, new_n1026_ );
nor g0853 ( new_n1196_, new_n1194_, new_n1195_ );
nor g0854 ( new_n1197_, new_n1196_, new_n1193_ );
not g0855 ( new_n1198_, new_n1197_ );
nand g0856 ( new_n1199_, new_n1198_, keyIn_0_204 );
not g0857 ( new_n1200_, new_n1199_ );
nor g0858 ( new_n1201_, new_n1198_, keyIn_0_204 );
nor g0859 ( new_n1202_, new_n1200_, new_n1201_ );
nor g0860 ( new_n1203_, new_n1202_, new_n1192_ );
not g0861 ( new_n1204_, new_n1203_ );
nand g0862 ( new_n1205_, new_n1204_, keyIn_0_213 );
not g0863 ( new_n1206_, new_n1205_ );
nor g0864 ( new_n1207_, new_n1204_, keyIn_0_213 );
nor g0865 ( new_n1208_, new_n1206_, new_n1207_ );
nor g0866 ( new_n1209_, new_n1208_, new_n977_ );
nor g0867 ( new_n1210_, new_n1209_, new_n976_ );
nand g0868 ( new_n1211_, new_n1209_, new_n976_ );
not g0869 ( new_n1212_, new_n1211_ );
nor g0870 ( new_n1213_, new_n1212_, new_n1210_ );
nand g0871 ( new_n1214_, N106, N210 );
not g0872 ( new_n1215_, new_n1214_ );
nor g0873 ( new_n1216_, new_n1213_, new_n1215_ );
not g0874 ( new_n1217_, new_n1216_ );
nor g0875 ( new_n1218_, new_n1217_, keyIn_0_230 );
nand g0876 ( new_n1219_, new_n1217_, keyIn_0_230 );
not g0877 ( new_n1220_, keyIn_0_197 );
not g0878 ( new_n1221_, N228 );
nor g0879 ( new_n1222_, new_n1025_, new_n1221_ );
not g0880 ( new_n1223_, new_n1222_ );
nand g0881 ( new_n1224_, new_n1223_, keyIn_0_175 );
not g0882 ( new_n1225_, keyIn_0_175 );
nand g0883 ( new_n1226_, new_n1222_, new_n1225_ );
nand g0884 ( new_n1227_, new_n1224_, new_n1226_ );
not g0885 ( new_n1228_, N237 );
nor g0886 ( new_n1229_, new_n1020_, keyIn_0_153 );
nand g0887 ( new_n1230_, new_n1020_, keyIn_0_153 );
not g0888 ( new_n1231_, new_n1230_ );
nor g0889 ( new_n1232_, new_n1231_, new_n1229_ );
nor g0890 ( new_n1233_, new_n1232_, new_n1228_ );
not g0891 ( new_n1234_, new_n1233_ );
nand g0892 ( new_n1235_, new_n1234_, keyIn_0_176 );
not g0893 ( new_n1236_, keyIn_0_176 );
nand g0894 ( new_n1237_, new_n1233_, new_n1236_ );
nand g0895 ( new_n1238_, new_n1235_, new_n1237_ );
nand g0896 ( new_n1239_, new_n1227_, new_n1238_ );
nor g0897 ( new_n1240_, new_n1239_, new_n1220_ );
nand g0898 ( new_n1241_, new_n1239_, new_n1220_ );
not g0899 ( new_n1242_, keyIn_0_155 );
not g0900 ( new_n1243_, keyIn_0_132 );
nor g0901 ( new_n1244_, new_n1007_, new_n956_ );
not g0902 ( new_n1245_, new_n1244_ );
nor g0903 ( new_n1246_, new_n1245_, new_n1243_ );
nand g0904 ( new_n1247_, new_n952_, N183 );
nand g0905 ( new_n1248_, new_n1245_, new_n1243_ );
nand g0906 ( new_n1249_, new_n1248_, new_n1247_ );
nor g0907 ( new_n1250_, new_n1249_, new_n1246_ );
nor g0908 ( new_n1251_, new_n1250_, new_n1242_ );
not g0909 ( new_n1252_, new_n1250_ );
nor g0910 ( new_n1253_, new_n1252_, keyIn_0_155 );
nor g0911 ( new_n1254_, new_n1253_, new_n1251_ );
nand g0912 ( new_n1255_, new_n1241_, new_n1254_ );
nor g0913 ( new_n1256_, new_n1255_, new_n1240_ );
nand g0914 ( new_n1257_, new_n1219_, new_n1256_ );
nor g0915 ( new_n1258_, new_n1257_, new_n1218_ );
not g0916 ( new_n1259_, new_n1258_ );
nand g0917 ( new_n1260_, new_n1259_, new_n975_ );
nand g0918 ( new_n1261_, new_n1258_, keyIn_0_240 );
nand g0919 ( N863, new_n1260_, new_n1261_ );
not g0920 ( new_n1263_, keyIn_0_241 );
not g0921 ( new_n1264_, keyIn_0_220 );
not g0922 ( new_n1265_, keyIn_0_214 );
not g0923 ( new_n1266_, keyIn_0_157 );
nor g0924 ( new_n1267_, new_n1151_, new_n1113_ );
nor g0925 ( new_n1268_, new_n1267_, new_n1266_ );
nand g0926 ( new_n1269_, new_n1267_, new_n1266_ );
not g0927 ( new_n1270_, new_n1269_ );
nor g0928 ( new_n1271_, new_n1270_, new_n1268_ );
not g0929 ( new_n1272_, new_n1271_ );
not g0930 ( new_n1273_, keyIn_0_198 );
not g0931 ( new_n1274_, keyIn_0_186 );
nor g0932 ( new_n1275_, new_n1164_, new_n1122_ );
not g0933 ( new_n1276_, new_n1275_ );
nand g0934 ( new_n1277_, new_n1276_, new_n1274_ );
not g0935 ( new_n1278_, new_n1277_ );
nor g0936 ( new_n1279_, new_n1276_, new_n1274_ );
nor g0937 ( new_n1280_, new_n1278_, new_n1279_ );
not g0938 ( new_n1281_, keyIn_0_180 );
nor g0939 ( new_n1282_, new_n1101_, keyIn_0_159 );
not g0940 ( new_n1283_, new_n1104_ );
nor g0941 ( new_n1284_, new_n1283_, new_n1282_ );
nor g0942 ( new_n1285_, new_n1284_, new_n1281_ );
nor g0943 ( new_n1286_, new_n1105_, keyIn_0_180 );
nor g0944 ( new_n1287_, new_n1285_, new_n1286_ );
not g0945 ( new_n1288_, keyIn_0_166 );
nor g0946 ( new_n1289_, new_n1136_, new_n1122_ );
nor g0947 ( new_n1290_, new_n1289_, new_n1288_ );
nand g0948 ( new_n1291_, new_n1289_, new_n1288_ );
not g0949 ( new_n1292_, new_n1291_ );
nor g0950 ( new_n1293_, new_n1292_, new_n1290_ );
nand g0951 ( new_n1294_, new_n1287_, new_n1293_ );
nor g0952 ( new_n1295_, new_n1280_, new_n1294_ );
not g0953 ( new_n1296_, new_n1295_ );
nand g0954 ( new_n1297_, new_n1296_, new_n1273_ );
not g0955 ( new_n1298_, new_n1297_ );
nor g0956 ( new_n1299_, new_n1296_, new_n1273_ );
nor g0957 ( new_n1300_, new_n1298_, new_n1299_ );
not g0958 ( new_n1301_, new_n1300_ );
nor g0959 ( new_n1302_, new_n1301_, new_n1272_ );
nor g0960 ( new_n1303_, new_n1302_, keyIn_0_206 );
nand g0961 ( new_n1304_, new_n1302_, keyIn_0_206 );
not g0962 ( new_n1305_, new_n1304_ );
nor g0963 ( new_n1306_, new_n1305_, new_n1303_ );
nor g0964 ( new_n1307_, new_n1300_, new_n1271_ );
not g0965 ( new_n1308_, new_n1307_ );
nand g0966 ( new_n1309_, new_n1308_, keyIn_0_207 );
not g0967 ( new_n1310_, new_n1309_ );
nor g0968 ( new_n1311_, new_n1308_, keyIn_0_207 );
nor g0969 ( new_n1312_, new_n1310_, new_n1311_ );
nor g0970 ( new_n1313_, new_n1312_, new_n1306_ );
not g0971 ( new_n1314_, new_n1313_ );
nand g0972 ( new_n1315_, new_n1314_, new_n1265_ );
not g0973 ( new_n1316_, new_n1315_ );
nor g0974 ( new_n1317_, new_n1314_, new_n1265_ );
nor g0975 ( new_n1318_, new_n1316_, new_n1317_ );
nor g0976 ( new_n1319_, new_n1318_, new_n977_ );
nor g0977 ( new_n1320_, new_n1319_, new_n1264_ );
nand g0978 ( new_n1321_, new_n1319_, new_n1264_ );
not g0979 ( new_n1322_, new_n1321_ );
nor g0980 ( new_n1323_, new_n1322_, new_n1320_ );
nand g0981 ( new_n1324_, N111, N210 );
not g0982 ( new_n1325_, new_n1324_ );
nor g0983 ( new_n1326_, new_n1323_, new_n1325_ );
not g0984 ( new_n1327_, new_n1326_ );
nor g0985 ( new_n1328_, new_n1327_, keyIn_0_231 );
nand g0986 ( new_n1329_, new_n1327_, keyIn_0_231 );
not g0987 ( new_n1330_, keyIn_0_199 );
not g0988 ( new_n1331_, keyIn_0_178 );
nor g0989 ( new_n1332_, new_n1271_, new_n1221_ );
not g0990 ( new_n1333_, new_n1332_ );
nand g0991 ( new_n1334_, new_n1333_, new_n1331_ );
not g0992 ( new_n1335_, new_n1334_ );
nor g0993 ( new_n1336_, new_n1333_, new_n1331_ );
nor g0994 ( new_n1337_, new_n1335_, new_n1336_ );
nor g0995 ( new_n1338_, new_n1153_, new_n1228_ );
nor g0996 ( new_n1339_, new_n1338_, keyIn_0_179 );
nand g0997 ( new_n1340_, new_n1338_, keyIn_0_179 );
not g0998 ( new_n1341_, new_n1340_ );
nor g0999 ( new_n1342_, new_n1341_, new_n1339_ );
nor g1000 ( new_n1343_, new_n1337_, new_n1342_ );
nor g1001 ( new_n1344_, new_n1343_, new_n1330_ );
not g1002 ( new_n1345_, new_n1343_ );
nor g1003 ( new_n1346_, new_n1345_, keyIn_0_199 );
nor g1004 ( new_n1347_, new_n1346_, new_n1344_ );
not g1005 ( new_n1348_, keyIn_0_158 );
nand g1006 ( new_n1349_, new_n1056_, N246 );
nand g1007 ( new_n1350_, N255, N259 );
nand g1008 ( new_n1351_, new_n1349_, new_n1350_ );
not g1009 ( new_n1352_, new_n1351_ );
nand g1010 ( new_n1353_, new_n1352_, new_n1348_ );
nand g1011 ( new_n1354_, new_n952_, N189 );
nand g1012 ( new_n1355_, new_n1351_, keyIn_0_158 );
nand g1013 ( new_n1356_, new_n1355_, new_n1354_ );
not g1014 ( new_n1357_, new_n1356_ );
nand g1015 ( new_n1358_, new_n1357_, new_n1353_ );
nor g1016 ( new_n1359_, new_n1347_, new_n1358_ );
nand g1017 ( new_n1360_, new_n1329_, new_n1359_ );
nor g1018 ( new_n1361_, new_n1360_, new_n1328_ );
not g1019 ( new_n1362_, new_n1361_ );
nand g1020 ( new_n1363_, new_n1362_, new_n1263_ );
nand g1021 ( new_n1364_, new_n1361_, keyIn_0_241 );
nand g1022 ( N864, new_n1363_, new_n1364_ );
not g1023 ( new_n1366_, keyIn_0_242 );
not g1024 ( new_n1367_, keyIn_0_215 );
not g1025 ( new_n1368_, keyIn_0_209 );
not g1026 ( new_n1369_, keyIn_0_183 );
nor g1027 ( new_n1370_, new_n1164_, new_n1369_ );
nor g1028 ( new_n1371_, new_n922_, keyIn_0_183 );
nor g1029 ( new_n1372_, new_n1370_, new_n1371_ );
not g1030 ( new_n1373_, keyIn_0_165 );
nor g1031 ( new_n1374_, new_n1127_, new_n1373_ );
nor g1032 ( new_n1375_, new_n1136_, keyIn_0_165 );
nor g1033 ( new_n1376_, new_n1374_, new_n1375_ );
nor g1034 ( new_n1377_, new_n1372_, new_n1376_ );
not g1035 ( new_n1378_, new_n1377_ );
nand g1036 ( new_n1379_, new_n1378_, keyIn_0_200 );
not g1037 ( new_n1380_, new_n1379_ );
nor g1038 ( new_n1381_, new_n1378_, keyIn_0_200 );
nor g1039 ( new_n1382_, new_n1380_, new_n1381_ );
not g1040 ( new_n1383_, new_n1382_ );
not g1041 ( new_n1384_, keyIn_0_160 );
nor g1042 ( new_n1385_, new_n1101_, new_n1122_ );
nor g1043 ( new_n1386_, new_n1385_, new_n1384_ );
nand g1044 ( new_n1387_, new_n1385_, new_n1384_ );
not g1045 ( new_n1388_, new_n1387_ );
nor g1046 ( new_n1389_, new_n1388_, new_n1386_ );
not g1047 ( new_n1390_, new_n1389_ );
nor g1048 ( new_n1391_, new_n1383_, new_n1390_ );
not g1049 ( new_n1392_, new_n1391_ );
nand g1050 ( new_n1393_, new_n1392_, new_n1368_ );
nand g1051 ( new_n1394_, new_n1391_, keyIn_0_209 );
nand g1052 ( new_n1395_, new_n1393_, new_n1394_ );
not g1053 ( new_n1396_, keyIn_0_208 );
nor g1054 ( new_n1397_, new_n1382_, new_n1389_ );
not g1055 ( new_n1398_, new_n1397_ );
nand g1056 ( new_n1399_, new_n1398_, new_n1396_ );
nand g1057 ( new_n1400_, new_n1397_, keyIn_0_208 );
nand g1058 ( new_n1401_, new_n1399_, new_n1400_ );
nand g1059 ( new_n1402_, new_n1395_, new_n1401_ );
nor g1060 ( new_n1403_, new_n1402_, new_n1367_ );
nand g1061 ( new_n1404_, new_n1402_, new_n1367_ );
nand g1062 ( new_n1405_, new_n1404_, N219 );
nor g1063 ( new_n1406_, new_n1405_, new_n1403_ );
nor g1064 ( new_n1407_, new_n1406_, keyIn_0_221 );
nand g1065 ( new_n1408_, new_n1406_, keyIn_0_221 );
not g1066 ( new_n1409_, new_n1408_ );
nor g1067 ( new_n1410_, new_n1409_, new_n1407_ );
nand g1068 ( new_n1411_, N116, N210 );
not g1069 ( new_n1412_, new_n1411_ );
nor g1070 ( new_n1413_, new_n1410_, new_n1412_ );
not g1071 ( new_n1414_, new_n1413_ );
nand g1072 ( new_n1415_, new_n1414_, keyIn_0_232 );
not g1073 ( new_n1416_, new_n1415_ );
nor g1074 ( new_n1417_, new_n1414_, keyIn_0_232 );
nor g1075 ( new_n1418_, new_n1416_, new_n1417_ );
nor g1076 ( new_n1419_, new_n1390_, new_n1221_ );
nor g1077 ( new_n1420_, new_n1419_, keyIn_0_181 );
nand g1078 ( new_n1421_, new_n1419_, keyIn_0_181 );
not g1079 ( new_n1422_, new_n1421_ );
nor g1080 ( new_n1423_, new_n1422_, new_n1420_ );
not g1081 ( new_n1424_, keyIn_0_182 );
nor g1082 ( new_n1425_, new_n1284_, new_n1228_ );
not g1083 ( new_n1426_, new_n1425_ );
nand g1084 ( new_n1427_, new_n1426_, new_n1424_ );
not g1085 ( new_n1428_, new_n1427_ );
nor g1086 ( new_n1429_, new_n1426_, new_n1424_ );
nor g1087 ( new_n1430_, new_n1428_, new_n1429_ );
nor g1088 ( new_n1431_, new_n1423_, new_n1430_ );
not g1089 ( new_n1432_, new_n1431_ );
nand g1090 ( new_n1433_, new_n1432_, keyIn_0_201 );
not g1091 ( new_n1434_, new_n1433_ );
nor g1092 ( new_n1435_, new_n1432_, keyIn_0_201 );
nor g1093 ( new_n1436_, new_n1434_, new_n1435_ );
nand g1094 ( new_n1437_, new_n1096_, N246 );
nand g1095 ( new_n1438_, N255, N260 );
nand g1096 ( new_n1439_, new_n1437_, new_n1438_ );
nor g1097 ( new_n1440_, new_n1439_, keyIn_0_161 );
nand g1098 ( new_n1441_, new_n952_, N195 );
nand g1099 ( new_n1442_, new_n1439_, keyIn_0_161 );
nand g1100 ( new_n1443_, new_n1442_, new_n1441_ );
nor g1101 ( new_n1444_, new_n1443_, new_n1440_ );
not g1102 ( new_n1445_, new_n1444_ );
nor g1103 ( new_n1446_, new_n1436_, new_n1445_ );
not g1104 ( new_n1447_, new_n1446_ );
nor g1105 ( new_n1448_, new_n1418_, new_n1447_ );
not g1106 ( new_n1449_, new_n1448_ );
nand g1107 ( new_n1450_, new_n1449_, new_n1366_ );
nand g1108 ( new_n1451_, new_n1448_, keyIn_0_242 );
nand g1109 ( N865, new_n1450_, new_n1451_ );
not g1110 ( new_n1453_, keyIn_0_248 );
not g1111 ( new_n1454_, keyIn_0_212 );
nand g1112 ( new_n1455_, new_n1196_, new_n1013_ );
nand g1113 ( new_n1456_, new_n1455_, keyIn_0_211 );
not g1114 ( new_n1457_, keyIn_0_211 );
nor g1115 ( new_n1458_, new_n1187_, new_n1014_ );
nand g1116 ( new_n1459_, new_n1458_, new_n1457_ );
nand g1117 ( new_n1460_, new_n1456_, new_n1459_ );
not g1118 ( new_n1461_, keyIn_0_174 );
not g1119 ( new_n1462_, new_n1232_ );
nand g1120 ( new_n1463_, new_n1462_, new_n1461_ );
nand g1121 ( new_n1464_, new_n1232_, keyIn_0_174 );
nand g1122 ( new_n1465_, new_n1463_, new_n1464_ );
nand g1123 ( new_n1466_, new_n1460_, new_n1465_ );
nand g1124 ( new_n1467_, new_n1466_, new_n1454_ );
not g1125 ( new_n1468_, new_n1467_ );
nor g1126 ( new_n1469_, new_n1466_, new_n1454_ );
nor g1127 ( new_n1470_, new_n1468_, new_n1469_ );
not g1128 ( new_n1471_, keyIn_0_108 );
not g1129 ( new_n1472_, keyIn_0_97 );
nand g1130 ( new_n1473_, new_n819_, N96 );
not g1131 ( new_n1474_, new_n1473_ );
nor g1132 ( new_n1475_, new_n1474_, keyIn_0_76 );
nand g1133 ( new_n1476_, new_n1474_, keyIn_0_76 );
not g1134 ( new_n1477_, new_n1476_ );
nor g1135 ( new_n1478_, new_n1477_, new_n1475_ );
nand g1136 ( new_n1479_, N51, N138 );
not g1137 ( new_n1480_, new_n1479_ );
nor g1138 ( new_n1481_, new_n1478_, new_n1480_ );
not g1139 ( new_n1482_, new_n1481_ );
nand g1140 ( new_n1483_, new_n1482_, new_n1472_ );
not g1141 ( new_n1484_, new_n1483_ );
nor g1142 ( new_n1485_, new_n1482_, new_n1472_ );
nor g1143 ( new_n1486_, new_n1484_, new_n1485_ );
not g1144 ( new_n1487_, keyIn_0_58 );
nor g1145 ( new_n1488_, new_n836_, new_n353_ );
not g1146 ( new_n1489_, new_n1488_ );
nor g1147 ( new_n1490_, new_n1489_, keyIn_0_45 );
nand g1148 ( new_n1491_, new_n1489_, keyIn_0_45 );
nand g1149 ( new_n1492_, new_n1491_, new_n844_ );
nor g1150 ( new_n1493_, new_n1492_, new_n1490_ );
not g1151 ( new_n1494_, new_n1493_ );
nor g1152 ( new_n1495_, new_n1494_, new_n1487_ );
nor g1153 ( new_n1496_, new_n1493_, keyIn_0_58 );
nor g1154 ( new_n1497_, new_n1495_, new_n1496_ );
not g1155 ( new_n1498_, keyIn_0_57 );
nor g1156 ( new_n1499_, new_n748_, new_n392_ );
nor g1157 ( new_n1500_, new_n1499_, keyIn_0_44 );
nand g1158 ( new_n1501_, new_n1499_, keyIn_0_44 );
not g1159 ( new_n1502_, new_n1501_ );
nor g1160 ( new_n1503_, new_n1502_, new_n1500_ );
nor g1161 ( new_n1504_, new_n1503_, new_n1032_ );
not g1162 ( new_n1505_, new_n1504_ );
nand g1163 ( new_n1506_, new_n1505_, new_n1498_ );
not g1164 ( new_n1507_, new_n1506_ );
nor g1165 ( new_n1508_, new_n1505_, new_n1498_ );
nor g1166 ( new_n1509_, new_n1507_, new_n1508_ );
nor g1167 ( new_n1510_, new_n1497_, new_n1509_ );
nor g1168 ( new_n1511_, new_n1510_, keyIn_0_77 );
nand g1169 ( new_n1512_, new_n1510_, keyIn_0_77 );
not g1170 ( new_n1513_, new_n1512_ );
nor g1171 ( new_n1514_, new_n1513_, new_n1511_ );
nor g1172 ( new_n1515_, new_n1486_, new_n1514_ );
nor g1173 ( new_n1516_, new_n1515_, new_n1471_ );
nand g1174 ( new_n1517_, new_n1515_, new_n1471_ );
not g1175 ( new_n1518_, new_n1517_ );
nor g1176 ( new_n1519_, new_n1518_, new_n1516_ );
not g1177 ( new_n1520_, new_n1519_ );
nor g1178 ( new_n1521_, new_n1520_, N165 );
nor g1179 ( new_n1522_, new_n1521_, keyIn_0_122 );
nand g1180 ( new_n1523_, new_n1521_, keyIn_0_122 );
not g1181 ( new_n1524_, new_n1523_ );
nor g1182 ( new_n1525_, new_n1524_, new_n1522_ );
not g1183 ( new_n1526_, new_n1525_ );
not g1184 ( new_n1527_, keyIn_0_125 );
not g1185 ( new_n1528_, keyIn_0_109 );
nor g1186 ( new_n1529_, new_n981_, new_n495_ );
nor g1187 ( new_n1530_, new_n1529_, keyIn_0_78 );
nand g1188 ( new_n1531_, new_n1529_, keyIn_0_78 );
not g1189 ( new_n1532_, new_n1531_ );
nor g1190 ( new_n1533_, new_n1532_, new_n1530_ );
nand g1191 ( new_n1534_, N17, N138 );
not g1192 ( new_n1535_, new_n1534_ );
nor g1193 ( new_n1536_, new_n1533_, new_n1535_ );
not g1194 ( new_n1537_, new_n1536_ );
nand g1195 ( new_n1538_, new_n1537_, keyIn_0_98 );
not g1196 ( new_n1539_, new_n1538_ );
nor g1197 ( new_n1540_, new_n1537_, keyIn_0_98 );
nor g1198 ( new_n1541_, new_n1539_, new_n1540_ );
not g1199 ( new_n1542_, keyIn_0_60 );
nor g1200 ( new_n1543_, new_n1494_, new_n1542_ );
nor g1201 ( new_n1544_, new_n1493_, keyIn_0_60 );
nor g1202 ( new_n1545_, new_n1543_, new_n1544_ );
nor g1203 ( new_n1546_, new_n1503_, new_n1072_ );
not g1204 ( new_n1547_, new_n1546_ );
nand g1205 ( new_n1548_, new_n1547_, keyIn_0_59 );
not g1206 ( new_n1549_, new_n1548_ );
nor g1207 ( new_n1550_, new_n1547_, keyIn_0_59 );
nor g1208 ( new_n1551_, new_n1549_, new_n1550_ );
nor g1209 ( new_n1552_, new_n1545_, new_n1551_ );
nor g1210 ( new_n1553_, new_n1552_, keyIn_0_79 );
nand g1211 ( new_n1554_, new_n1552_, keyIn_0_79 );
not g1212 ( new_n1555_, new_n1554_ );
nor g1213 ( new_n1556_, new_n1555_, new_n1553_ );
nor g1214 ( new_n1557_, new_n1541_, new_n1556_ );
nor g1215 ( new_n1558_, new_n1557_, new_n1528_ );
nand g1216 ( new_n1559_, new_n1557_, new_n1528_ );
not g1217 ( new_n1560_, new_n1559_ );
nor g1218 ( new_n1561_, new_n1560_, new_n1558_ );
nor g1219 ( new_n1562_, new_n1561_, N171 );
not g1220 ( new_n1563_, new_n1562_ );
nand g1221 ( new_n1564_, new_n1563_, new_n1527_ );
not g1222 ( new_n1565_, new_n1564_ );
nor g1223 ( new_n1566_, new_n1563_, new_n1527_ );
nor g1224 ( new_n1567_, new_n1565_, new_n1566_ );
nor g1225 ( new_n1568_, new_n1526_, new_n1567_ );
not g1226 ( new_n1569_, new_n1568_ );
not g1227 ( new_n1570_, keyIn_0_128 );
not g1228 ( new_n1571_, keyIn_0_110 );
not g1229 ( new_n1572_, keyIn_0_99 );
nor g1230 ( new_n1573_, new_n981_, new_n497_ );
not g1231 ( new_n1574_, new_n1573_ );
nor g1232 ( new_n1575_, new_n1574_, keyIn_0_80 );
nand g1233 ( new_n1576_, N138, N152 );
nand g1234 ( new_n1577_, new_n1574_, keyIn_0_80 );
nand g1235 ( new_n1578_, new_n1577_, new_n1576_ );
nor g1236 ( new_n1579_, new_n1578_, new_n1575_ );
not g1237 ( new_n1580_, new_n1579_ );
nor g1238 ( new_n1581_, new_n1580_, new_n1572_ );
not g1239 ( new_n1582_, keyIn_0_81 );
not g1240 ( new_n1583_, keyIn_0_62 );
nor g1241 ( new_n1584_, new_n1494_, new_n1583_ );
nor g1242 ( new_n1585_, new_n1493_, keyIn_0_62 );
nor g1243 ( new_n1586_, new_n1584_, new_n1585_ );
nor g1244 ( new_n1587_, new_n1503_, new_n760_ );
not g1245 ( new_n1588_, new_n1587_ );
nand g1246 ( new_n1589_, new_n1588_, keyIn_0_61 );
not g1247 ( new_n1590_, new_n1589_ );
nor g1248 ( new_n1591_, new_n1588_, keyIn_0_61 );
nor g1249 ( new_n1592_, new_n1590_, new_n1591_ );
nor g1250 ( new_n1593_, new_n1586_, new_n1592_ );
nor g1251 ( new_n1594_, new_n1593_, new_n1582_ );
nand g1252 ( new_n1595_, new_n1593_, new_n1582_ );
not g1253 ( new_n1596_, new_n1595_ );
nor g1254 ( new_n1597_, new_n1596_, new_n1594_ );
nor g1255 ( new_n1598_, new_n1579_, keyIn_0_99 );
nor g1256 ( new_n1599_, new_n1597_, new_n1598_ );
not g1257 ( new_n1600_, new_n1599_ );
nor g1258 ( new_n1601_, new_n1600_, new_n1581_ );
nor g1259 ( new_n1602_, new_n1601_, new_n1571_ );
nand g1260 ( new_n1603_, new_n1601_, new_n1571_ );
not g1261 ( new_n1604_, new_n1603_ );
nor g1262 ( new_n1605_, new_n1604_, new_n1602_ );
not g1263 ( new_n1606_, new_n1605_ );
nor g1264 ( new_n1607_, new_n1606_, N177 );
nor g1265 ( new_n1608_, new_n1607_, new_n1570_ );
nand g1266 ( new_n1609_, new_n1607_, new_n1570_ );
not g1267 ( new_n1610_, new_n1609_ );
nor g1268 ( new_n1611_, new_n1610_, new_n1608_ );
not g1269 ( new_n1612_, new_n1611_ );
nor g1270 ( new_n1613_, new_n1569_, new_n1612_ );
nand g1271 ( new_n1614_, new_n1470_, new_n1613_ );
nor g1272 ( new_n1615_, new_n1614_, keyIn_0_225 );
nand g1273 ( new_n1616_, new_n1614_, keyIn_0_225 );
not g1274 ( new_n1617_, keyIn_0_127 );
nor g1275 ( new_n1618_, new_n1605_, new_n582_ );
not g1276 ( new_n1619_, new_n1618_ );
nand g1277 ( new_n1620_, new_n1619_, new_n1617_ );
not g1278 ( new_n1621_, new_n1620_ );
nor g1279 ( new_n1622_, new_n1619_, new_n1617_ );
nor g1280 ( new_n1623_, new_n1621_, new_n1622_ );
nor g1281 ( new_n1624_, new_n1623_, keyIn_0_150 );
nand g1282 ( new_n1625_, new_n1623_, keyIn_0_150 );
not g1283 ( new_n1626_, new_n1625_ );
nor g1284 ( new_n1627_, new_n1626_, new_n1624_ );
nor g1285 ( new_n1628_, new_n1627_, new_n1569_ );
not g1286 ( new_n1629_, new_n1628_ );
nand g1287 ( new_n1630_, new_n1629_, keyIn_0_191 );
not g1288 ( new_n1631_, new_n1630_ );
nor g1289 ( new_n1632_, new_n1629_, keyIn_0_191 );
nor g1290 ( new_n1633_, new_n1631_, new_n1632_ );
not g1291 ( new_n1634_, keyIn_0_190 );
not g1292 ( new_n1635_, keyIn_0_147 );
not g1293 ( new_n1636_, new_n1561_ );
nor g1294 ( new_n1637_, new_n1636_, new_n580_ );
nor g1295 ( new_n1638_, new_n1637_, keyIn_0_124 );
nand g1296 ( new_n1639_, new_n1637_, keyIn_0_124 );
not g1297 ( new_n1640_, new_n1639_ );
nor g1298 ( new_n1641_, new_n1640_, new_n1638_ );
nor g1299 ( new_n1642_, new_n1641_, new_n1635_ );
not g1300 ( new_n1643_, new_n1641_ );
nor g1301 ( new_n1644_, new_n1643_, keyIn_0_147 );
nor g1302 ( new_n1645_, new_n1644_, new_n1642_ );
nor g1303 ( new_n1646_, new_n1645_, new_n1526_ );
not g1304 ( new_n1647_, new_n1646_ );
nor g1305 ( new_n1648_, new_n1647_, new_n1634_ );
nand g1306 ( new_n1649_, new_n1647_, new_n1634_ );
not g1307 ( new_n1650_, new_n1649_ );
not g1308 ( new_n1651_, keyIn_0_144 );
not g1309 ( new_n1652_, keyIn_0_121 );
not g1310 ( new_n1653_, N165 );
nor g1311 ( new_n1654_, new_n1519_, new_n1653_ );
not g1312 ( new_n1655_, new_n1654_ );
nand g1313 ( new_n1656_, new_n1655_, new_n1652_ );
not g1314 ( new_n1657_, new_n1656_ );
nor g1315 ( new_n1658_, new_n1655_, new_n1652_ );
nor g1316 ( new_n1659_, new_n1657_, new_n1658_ );
nor g1317 ( new_n1660_, new_n1659_, new_n1651_ );
not g1318 ( new_n1661_, new_n1659_ );
nor g1319 ( new_n1662_, new_n1661_, keyIn_0_144 );
nor g1320 ( new_n1663_, new_n1662_, new_n1660_ );
nor g1321 ( new_n1664_, new_n1663_, keyIn_0_168 );
nand g1322 ( new_n1665_, new_n1663_, keyIn_0_168 );
not g1323 ( new_n1666_, new_n1665_ );
nor g1324 ( new_n1667_, new_n1666_, new_n1664_ );
nor g1325 ( new_n1668_, new_n1650_, new_n1667_ );
not g1326 ( new_n1669_, new_n1668_ );
nor g1327 ( new_n1670_, new_n1669_, new_n1648_ );
not g1328 ( new_n1671_, new_n1670_ );
nor g1329 ( new_n1672_, new_n1671_, new_n1633_ );
nand g1330 ( new_n1673_, new_n1616_, new_n1672_ );
nor g1331 ( new_n1674_, new_n1673_, new_n1615_ );
nor g1332 ( new_n1675_, new_n1674_, keyIn_0_226 );
not g1333 ( new_n1676_, keyIn_0_226 );
not g1334 ( new_n1677_, new_n1615_ );
not g1335 ( new_n1678_, keyIn_0_225 );
not g1336 ( new_n1679_, new_n1466_ );
nand g1337 ( new_n1680_, new_n1679_, keyIn_0_212 );
nand g1338 ( new_n1681_, new_n1680_, new_n1467_ );
not g1339 ( new_n1682_, new_n1613_ );
nor g1340 ( new_n1683_, new_n1681_, new_n1682_ );
nor g1341 ( new_n1684_, new_n1683_, new_n1678_ );
not g1342 ( new_n1685_, new_n1672_ );
nor g1343 ( new_n1686_, new_n1684_, new_n1685_ );
nand g1344 ( new_n1687_, new_n1686_, new_n1677_ );
nor g1345 ( new_n1688_, new_n1687_, new_n1676_ );
nor g1346 ( new_n1689_, new_n1688_, new_n1675_ );
not g1347 ( new_n1690_, keyIn_0_107 );
nand g1348 ( new_n1691_, new_n819_, N91 );
not g1349 ( new_n1692_, new_n1691_ );
nor g1350 ( new_n1693_, new_n1692_, keyIn_0_74 );
nand g1351 ( new_n1694_, new_n1692_, keyIn_0_74 );
not g1352 ( new_n1695_, new_n1694_ );
nor g1353 ( new_n1696_, new_n1695_, new_n1693_ );
nand g1354 ( new_n1697_, N8, N138 );
not g1355 ( new_n1698_, new_n1697_ );
nor g1356 ( new_n1699_, new_n1696_, new_n1698_ );
not g1357 ( new_n1700_, new_n1699_ );
nor g1358 ( new_n1701_, new_n1700_, keyIn_0_96 );
not g1359 ( new_n1702_, keyIn_0_75 );
not g1360 ( new_n1703_, keyIn_0_56 );
nor g1361 ( new_n1704_, new_n1494_, new_n1703_ );
nor g1362 ( new_n1705_, new_n1493_, keyIn_0_56 );
nor g1363 ( new_n1706_, new_n1704_, new_n1705_ );
not g1364 ( new_n1707_, keyIn_0_55 );
nor g1365 ( new_n1708_, new_n1503_, new_n987_ );
not g1366 ( new_n1709_, new_n1708_ );
nand g1367 ( new_n1710_, new_n1709_, new_n1707_ );
not g1368 ( new_n1711_, new_n1710_ );
nor g1369 ( new_n1712_, new_n1709_, new_n1707_ );
nor g1370 ( new_n1713_, new_n1711_, new_n1712_ );
nor g1371 ( new_n1714_, new_n1706_, new_n1713_ );
not g1372 ( new_n1715_, new_n1714_ );
nand g1373 ( new_n1716_, new_n1715_, new_n1702_ );
nand g1374 ( new_n1717_, new_n1714_, keyIn_0_75 );
nand g1375 ( new_n1718_, new_n1716_, new_n1717_ );
nand g1376 ( new_n1719_, new_n1700_, keyIn_0_96 );
nand g1377 ( new_n1720_, new_n1719_, new_n1718_ );
nor g1378 ( new_n1721_, new_n1720_, new_n1701_ );
nor g1379 ( new_n1722_, new_n1721_, new_n1690_ );
nand g1380 ( new_n1723_, new_n1721_, new_n1690_ );
not g1381 ( new_n1724_, new_n1723_ );
nor g1382 ( new_n1725_, new_n1724_, new_n1722_ );
not g1383 ( new_n1726_, new_n1725_ );
nor g1384 ( new_n1727_, new_n1726_, N159 );
nor g1385 ( new_n1728_, new_n1727_, keyIn_0_119 );
nand g1386 ( new_n1729_, new_n1727_, keyIn_0_119 );
not g1387 ( new_n1730_, new_n1729_ );
nor g1388 ( new_n1731_, new_n1730_, new_n1728_ );
nor g1389 ( new_n1732_, new_n1689_, new_n1731_ );
not g1390 ( new_n1733_, new_n1732_ );
nor g1391 ( new_n1734_, new_n1733_, keyIn_0_243 );
not g1392 ( new_n1735_, keyIn_0_141 );
not g1393 ( new_n1736_, N159 );
nor g1394 ( new_n1737_, new_n1725_, new_n1736_ );
not g1395 ( new_n1738_, new_n1737_ );
nand g1396 ( new_n1739_, new_n1738_, keyIn_0_118 );
not g1397 ( new_n1740_, new_n1739_ );
nor g1398 ( new_n1741_, new_n1738_, keyIn_0_118 );
nor g1399 ( new_n1742_, new_n1740_, new_n1741_ );
nor g1400 ( new_n1743_, new_n1742_, new_n1735_ );
not g1401 ( new_n1744_, new_n1742_ );
nor g1402 ( new_n1745_, new_n1744_, keyIn_0_141 );
nor g1403 ( new_n1746_, new_n1745_, new_n1743_ );
nand g1404 ( new_n1747_, new_n1733_, keyIn_0_243 );
nand g1405 ( new_n1748_, new_n1747_, new_n1746_ );
nor g1406 ( new_n1749_, new_n1748_, new_n1734_ );
not g1407 ( new_n1750_, new_n1749_ );
nand g1408 ( new_n1751_, new_n1750_, new_n1453_ );
nand g1409 ( new_n1752_, new_n1749_, keyIn_0_248 );
nand g1410 ( N866, new_n1751_, new_n1752_ );
not g1411 ( new_n1754_, keyIn_0_247 );
not g1412 ( new_n1755_, keyIn_0_239 );
nor g1413 ( new_n1756_, new_n1612_, new_n1623_ );
nor g1414 ( new_n1757_, new_n1756_, keyIn_0_151 );
nand g1415 ( new_n1758_, new_n1756_, keyIn_0_151 );
not g1416 ( new_n1759_, new_n1758_ );
nor g1417 ( new_n1760_, new_n1759_, new_n1757_ );
not g1418 ( new_n1761_, new_n1760_ );
nor g1419 ( new_n1762_, new_n1681_, new_n1761_ );
not g1420 ( new_n1763_, new_n1762_ );
nand g1421 ( new_n1764_, new_n1763_, keyIn_0_218 );
not g1422 ( new_n1765_, keyIn_0_218 );
nand g1423 ( new_n1766_, new_n1762_, new_n1765_ );
nand g1424 ( new_n1767_, new_n1764_, new_n1766_ );
nor g1425 ( new_n1768_, new_n1470_, new_n1760_ );
not g1426 ( new_n1769_, new_n1768_ );
nand g1427 ( new_n1770_, new_n1769_, keyIn_0_217 );
not g1428 ( new_n1771_, keyIn_0_217 );
nand g1429 ( new_n1772_, new_n1768_, new_n1771_ );
nand g1430 ( new_n1773_, new_n1770_, new_n1772_ );
nand g1431 ( new_n1774_, new_n1773_, new_n1767_ );
nor g1432 ( new_n1775_, new_n1774_, keyIn_0_229 );
nand g1433 ( new_n1776_, new_n1774_, keyIn_0_229 );
nand g1434 ( new_n1777_, new_n1776_, N219 );
nor g1435 ( new_n1778_, new_n1777_, new_n1775_ );
nor g1436 ( new_n1779_, new_n1778_, new_n1755_ );
nand g1437 ( new_n1780_, new_n1778_, new_n1755_ );
not g1438 ( new_n1781_, new_n1780_ );
nor g1439 ( new_n1782_, new_n1781_, new_n1779_ );
nand g1440 ( new_n1783_, N101, N210 );
not g1441 ( new_n1784_, new_n1783_ );
nor g1442 ( new_n1785_, new_n1782_, new_n1784_ );
not g1443 ( new_n1786_, new_n1785_ );
nand g1444 ( new_n1787_, new_n1786_, new_n1754_ );
not g1445 ( new_n1788_, new_n1787_ );
nor g1446 ( new_n1789_, new_n1786_, new_n1754_ );
nor g1447 ( new_n1790_, new_n1788_, new_n1789_ );
not g1448 ( new_n1791_, keyIn_0_172 );
nor g1449 ( new_n1792_, new_n1761_, new_n1221_ );
nor g1450 ( new_n1793_, new_n1792_, new_n1791_ );
nand g1451 ( new_n1794_, new_n1792_, new_n1791_ );
not g1452 ( new_n1795_, new_n1794_ );
nor g1453 ( new_n1796_, new_n1795_, new_n1793_ );
not g1454 ( new_n1797_, keyIn_0_173 );
nor g1455 ( new_n1798_, new_n1627_, new_n1228_ );
not g1456 ( new_n1799_, new_n1798_ );
nand g1457 ( new_n1800_, new_n1799_, new_n1797_ );
not g1458 ( new_n1801_, new_n1800_ );
nor g1459 ( new_n1802_, new_n1799_, new_n1797_ );
nor g1460 ( new_n1803_, new_n1801_, new_n1802_ );
nor g1461 ( new_n1804_, new_n1796_, new_n1803_ );
not g1462 ( new_n1805_, new_n1804_ );
nor g1463 ( new_n1806_, new_n1805_, keyIn_0_195 );
nand g1464 ( new_n1807_, new_n1805_, keyIn_0_195 );
nor g1465 ( new_n1808_, new_n1605_, new_n956_ );
not g1466 ( new_n1809_, new_n1808_ );
nor g1467 ( new_n1810_, new_n1809_, keyIn_0_129 );
nand g1468 ( new_n1811_, new_n952_, N177 );
nand g1469 ( new_n1812_, new_n1809_, keyIn_0_129 );
nand g1470 ( new_n1813_, new_n1812_, new_n1811_ );
nor g1471 ( new_n1814_, new_n1813_, new_n1810_ );
nor g1472 ( new_n1815_, new_n1814_, keyIn_0_152 );
not g1473 ( new_n1816_, keyIn_0_152 );
not g1474 ( new_n1817_, new_n1814_ );
nor g1475 ( new_n1818_, new_n1817_, new_n1816_ );
nor g1476 ( new_n1819_, new_n1818_, new_n1815_ );
nand g1477 ( new_n1820_, new_n1807_, new_n1819_ );
nor g1478 ( new_n1821_, new_n1820_, new_n1806_ );
not g1479 ( new_n1822_, new_n1821_ );
nor g1480 ( new_n1823_, new_n1790_, new_n1822_ );
not g1481 ( new_n1824_, new_n1823_ );
nand g1482 ( new_n1825_, new_n1824_, keyIn_0_249 );
not g1483 ( new_n1826_, keyIn_0_249 );
nand g1484 ( new_n1827_, new_n1823_, new_n1826_ );
nand g1485 ( N874, new_n1825_, new_n1827_ );
not g1486 ( new_n1829_, keyIn_0_250 );
not g1487 ( new_n1830_, keyIn_0_244 );
nand g1488 ( new_n1831_, new_n1687_, new_n1676_ );
nand g1489 ( new_n1832_, new_n1674_, keyIn_0_226 );
nand g1490 ( new_n1833_, new_n1831_, new_n1832_ );
nor g1491 ( new_n1834_, new_n1742_, new_n1731_ );
not g1492 ( new_n1835_, new_n1834_ );
nand g1493 ( new_n1836_, new_n1835_, keyIn_0_142 );
not g1494 ( new_n1837_, new_n1836_ );
nor g1495 ( new_n1838_, new_n1835_, keyIn_0_142 );
nor g1496 ( new_n1839_, new_n1837_, new_n1838_ );
nand g1497 ( new_n1840_, new_n1833_, new_n1839_ );
nand g1498 ( new_n1841_, new_n1840_, keyIn_0_234 );
not g1499 ( new_n1842_, keyIn_0_234 );
not g1500 ( new_n1843_, new_n1840_ );
nand g1501 ( new_n1844_, new_n1843_, new_n1842_ );
nand g1502 ( new_n1845_, new_n1844_, new_n1841_ );
not g1503 ( new_n1846_, new_n1839_ );
nand g1504 ( new_n1847_, new_n1689_, new_n1846_ );
nand g1505 ( new_n1848_, new_n1847_, keyIn_0_233 );
not g1506 ( new_n1849_, keyIn_0_233 );
nor g1507 ( new_n1850_, new_n1833_, new_n1839_ );
nand g1508 ( new_n1851_, new_n1850_, new_n1849_ );
nand g1509 ( new_n1852_, new_n1848_, new_n1851_ );
nand g1510 ( new_n1853_, new_n1845_, new_n1852_ );
nor g1511 ( new_n1854_, new_n1853_, new_n1830_ );
nand g1512 ( new_n1855_, new_n1853_, new_n1830_ );
nand g1513 ( new_n1856_, new_n1855_, N219 );
nor g1514 ( new_n1857_, new_n1856_, new_n1854_ );
not g1515 ( new_n1858_, N210 );
nor g1516 ( new_n1859_, new_n848_, new_n1858_ );
nor g1517 ( new_n1860_, new_n1857_, new_n1859_ );
nor g1518 ( new_n1861_, new_n1860_, new_n1829_ );
not g1519 ( new_n1862_, new_n1861_ );
nand g1520 ( new_n1863_, new_n1860_, new_n1829_ );
nand g1521 ( new_n1864_, new_n1862_, new_n1863_ );
nor g1522 ( new_n1865_, new_n1846_, new_n1221_ );
nor g1523 ( new_n1866_, new_n1746_, new_n1228_ );
nor g1524 ( new_n1867_, new_n1865_, new_n1866_ );
not g1525 ( new_n1868_, new_n1867_ );
nor g1526 ( new_n1869_, new_n1868_, keyIn_0_192 );
not g1527 ( new_n1870_, keyIn_0_120 );
nor g1528 ( new_n1871_, new_n1725_, new_n956_ );
not g1529 ( new_n1872_, new_n1871_ );
nand g1530 ( new_n1873_, new_n1872_, new_n1870_ );
not g1531 ( new_n1874_, new_n1873_ );
nor g1532 ( new_n1875_, new_n1872_, new_n1870_ );
nor g1533 ( new_n1876_, new_n1874_, new_n1875_ );
nor g1534 ( new_n1877_, new_n951_, new_n1736_ );
nor g1535 ( new_n1878_, new_n1876_, new_n1877_ );
nor g1536 ( new_n1879_, new_n1878_, keyIn_0_143 );
nand g1537 ( new_n1880_, new_n1878_, keyIn_0_143 );
not g1538 ( new_n1881_, new_n1880_ );
nor g1539 ( new_n1882_, new_n1881_, new_n1879_ );
nand g1540 ( new_n1883_, new_n1868_, keyIn_0_192 );
not g1541 ( new_n1884_, new_n1883_ );
nor g1542 ( new_n1885_, new_n1884_, new_n1882_ );
not g1543 ( new_n1886_, new_n1885_ );
nor g1544 ( new_n1887_, new_n1886_, new_n1869_ );
nand g1545 ( new_n1888_, new_n1864_, new_n1887_ );
nand g1546 ( new_n1889_, new_n1888_, keyIn_0_253 );
not g1547 ( new_n1890_, keyIn_0_253 );
not g1548 ( new_n1891_, new_n1854_ );
not g1549 ( new_n1892_, new_n1856_ );
nand g1550 ( new_n1893_, new_n1892_, new_n1891_ );
not g1551 ( new_n1894_, new_n1859_ );
nand g1552 ( new_n1895_, new_n1893_, new_n1894_ );
nor g1553 ( new_n1896_, new_n1895_, keyIn_0_250 );
nor g1554 ( new_n1897_, new_n1896_, new_n1861_ );
not g1555 ( new_n1898_, new_n1887_ );
nor g1556 ( new_n1899_, new_n1897_, new_n1898_ );
nand g1557 ( new_n1900_, new_n1899_, new_n1890_ );
nand g1558 ( N878, new_n1900_, new_n1889_ );
not g1559 ( new_n1902_, keyIn_0_254 );
not g1560 ( new_n1903_, keyIn_0_251 );
not g1561 ( new_n1904_, keyIn_0_236 );
not g1562 ( new_n1905_, keyIn_0_224 );
nor g1563 ( new_n1906_, new_n1612_, new_n1567_ );
nand g1564 ( new_n1907_, new_n1470_, new_n1906_ );
nand g1565 ( new_n1908_, new_n1907_, new_n1905_ );
not g1566 ( new_n1909_, new_n1906_ );
nor g1567 ( new_n1910_, new_n1681_, new_n1909_ );
nand g1568 ( new_n1911_, new_n1910_, keyIn_0_224 );
nand g1569 ( new_n1912_, new_n1908_, new_n1911_ );
not g1570 ( new_n1913_, keyIn_0_189 );
not g1571 ( new_n1914_, new_n1567_ );
not g1572 ( new_n1915_, new_n1627_ );
nand g1573 ( new_n1916_, new_n1915_, new_n1914_ );
nor g1574 ( new_n1917_, new_n1916_, new_n1913_ );
nand g1575 ( new_n1918_, new_n1916_, new_n1913_ );
nor g1576 ( new_n1919_, new_n1645_, keyIn_0_169 );
not g1577 ( new_n1920_, keyIn_0_169 );
not g1578 ( new_n1921_, new_n1645_ );
nor g1579 ( new_n1922_, new_n1921_, new_n1920_ );
nor g1580 ( new_n1923_, new_n1922_, new_n1919_ );
nand g1581 ( new_n1924_, new_n1923_, new_n1918_ );
nor g1582 ( new_n1925_, new_n1924_, new_n1917_ );
nand g1583 ( new_n1926_, new_n1912_, new_n1925_ );
nand g1584 ( new_n1927_, new_n1926_, keyIn_0_227 );
not g1585 ( new_n1928_, keyIn_0_227 );
not g1586 ( new_n1929_, new_n1926_ );
nand g1587 ( new_n1930_, new_n1929_, new_n1928_ );
nand g1588 ( new_n1931_, new_n1930_, new_n1927_ );
not g1589 ( new_n1932_, keyIn_0_145 );
nor g1590 ( new_n1933_, new_n1661_, new_n1526_ );
nor g1591 ( new_n1934_, new_n1933_, new_n1932_ );
nand g1592 ( new_n1935_, new_n1933_, new_n1932_ );
not g1593 ( new_n1936_, new_n1935_ );
nor g1594 ( new_n1937_, new_n1936_, new_n1934_ );
nand g1595 ( new_n1938_, new_n1931_, new_n1937_ );
nand g1596 ( new_n1939_, new_n1938_, new_n1904_ );
not g1597 ( new_n1940_, new_n1927_ );
nor g1598 ( new_n1941_, new_n1926_, keyIn_0_227 );
nor g1599 ( new_n1942_, new_n1940_, new_n1941_ );
not g1600 ( new_n1943_, new_n1937_ );
nor g1601 ( new_n1944_, new_n1942_, new_n1943_ );
nand g1602 ( new_n1945_, new_n1944_, keyIn_0_236 );
nand g1603 ( new_n1946_, new_n1945_, new_n1939_ );
nand g1604 ( new_n1947_, new_n1942_, new_n1943_ );
nand g1605 ( new_n1948_, new_n1947_, keyIn_0_235 );
not g1606 ( new_n1949_, keyIn_0_235 );
nor g1607 ( new_n1950_, new_n1931_, new_n1937_ );
nand g1608 ( new_n1951_, new_n1950_, new_n1949_ );
nand g1609 ( new_n1952_, new_n1948_, new_n1951_ );
nand g1610 ( new_n1953_, new_n1946_, new_n1952_ );
nor g1611 ( new_n1954_, new_n1953_, keyIn_0_245 );
not g1612 ( new_n1955_, new_n1954_ );
nand g1613 ( new_n1956_, new_n1953_, keyIn_0_245 );
nand g1614 ( new_n1957_, new_n1956_, N219 );
not g1615 ( new_n1958_, new_n1957_ );
nand g1616 ( new_n1959_, new_n1958_, new_n1955_ );
nand g1617 ( new_n1960_, N91, N210 );
nand g1618 ( new_n1961_, new_n1959_, new_n1960_ );
nand g1619 ( new_n1962_, new_n1961_, new_n1903_ );
nor g1620 ( new_n1963_, new_n1957_, new_n1954_ );
not g1621 ( new_n1964_, new_n1960_ );
nor g1622 ( new_n1965_, new_n1963_, new_n1964_ );
nand g1623 ( new_n1966_, new_n1965_, keyIn_0_251 );
nand g1624 ( new_n1967_, new_n1962_, new_n1966_ );
nor g1625 ( new_n1968_, new_n1943_, new_n1221_ );
nor g1626 ( new_n1969_, new_n1663_, new_n1228_ );
nor g1627 ( new_n1970_, new_n1968_, new_n1969_ );
not g1628 ( new_n1971_, new_n1970_ );
nor g1629 ( new_n1972_, new_n1971_, keyIn_0_193 );
not g1630 ( new_n1973_, keyIn_0_146 );
nor g1631 ( new_n1974_, new_n1519_, new_n956_ );
not g1632 ( new_n1975_, new_n1974_ );
nand g1633 ( new_n1976_, new_n1975_, keyIn_0_123 );
not g1634 ( new_n1977_, new_n1976_ );
nor g1635 ( new_n1978_, new_n1975_, keyIn_0_123 );
nor g1636 ( new_n1979_, new_n1977_, new_n1978_ );
nor g1637 ( new_n1980_, new_n951_, new_n1653_ );
nor g1638 ( new_n1981_, new_n1979_, new_n1980_ );
nor g1639 ( new_n1982_, new_n1981_, new_n1973_ );
nand g1640 ( new_n1983_, new_n1981_, new_n1973_ );
not g1641 ( new_n1984_, new_n1983_ );
nor g1642 ( new_n1985_, new_n1984_, new_n1982_ );
nand g1643 ( new_n1986_, new_n1971_, keyIn_0_193 );
not g1644 ( new_n1987_, new_n1986_ );
nor g1645 ( new_n1988_, new_n1987_, new_n1985_ );
not g1646 ( new_n1989_, new_n1988_ );
nor g1647 ( new_n1990_, new_n1989_, new_n1972_ );
nand g1648 ( new_n1991_, new_n1967_, new_n1990_ );
nand g1649 ( new_n1992_, new_n1991_, new_n1902_ );
nor g1650 ( new_n1993_, new_n1965_, keyIn_0_251 );
nor g1651 ( new_n1994_, new_n1961_, new_n1903_ );
nor g1652 ( new_n1995_, new_n1994_, new_n1993_ );
not g1653 ( new_n1996_, new_n1990_ );
nor g1654 ( new_n1997_, new_n1995_, new_n1996_ );
nand g1655 ( new_n1998_, new_n1997_, keyIn_0_254 );
nand g1656 ( N879, new_n1998_, new_n1992_ );
not g1657 ( new_n2000_, keyIn_0_252 );
not g1658 ( new_n2001_, keyIn_0_148 );
nor g1659 ( new_n2002_, new_n1567_, new_n1641_ );
not g1660 ( new_n2003_, new_n2002_ );
nand g1661 ( new_n2004_, new_n2003_, new_n2001_ );
not g1662 ( new_n2005_, new_n2004_ );
nor g1663 ( new_n2006_, new_n2003_, new_n2001_ );
nor g1664 ( new_n2007_, new_n2005_, new_n2006_ );
not g1665 ( new_n2008_, new_n2007_ );
nand g1666 ( new_n2009_, new_n1470_, new_n1611_ );
nor g1667 ( new_n2010_, new_n2009_, keyIn_0_223 );
not g1668 ( new_n2011_, keyIn_0_171 );
nor g1669 ( new_n2012_, new_n1915_, new_n2011_ );
nor g1670 ( new_n2013_, new_n1627_, keyIn_0_171 );
nor g1671 ( new_n2014_, new_n2012_, new_n2013_ );
not g1672 ( new_n2015_, new_n2014_ );
nand g1673 ( new_n2016_, new_n2009_, keyIn_0_223 );
nand g1674 ( new_n2017_, new_n2016_, new_n2015_ );
nor g1675 ( new_n2018_, new_n2017_, new_n2010_ );
nor g1676 ( new_n2019_, new_n2018_, keyIn_0_228 );
not g1677 ( new_n2020_, new_n2019_ );
nand g1678 ( new_n2021_, new_n2018_, keyIn_0_228 );
nand g1679 ( new_n2022_, new_n2020_, new_n2021_ );
nand g1680 ( new_n2023_, new_n2022_, new_n2008_ );
nand g1681 ( new_n2024_, new_n2023_, keyIn_0_237 );
not g1682 ( new_n2025_, keyIn_0_237 );
not g1683 ( new_n2026_, new_n2021_ );
nor g1684 ( new_n2027_, new_n2026_, new_n2019_ );
nor g1685 ( new_n2028_, new_n2027_, new_n2007_ );
nand g1686 ( new_n2029_, new_n2028_, new_n2025_ );
nand g1687 ( new_n2030_, new_n2029_, new_n2024_ );
not g1688 ( new_n2031_, keyIn_0_238 );
nand g1689 ( new_n2032_, new_n2027_, new_n2007_ );
nand g1690 ( new_n2033_, new_n2032_, new_n2031_ );
nor g1691 ( new_n2034_, new_n2022_, new_n2008_ );
nand g1692 ( new_n2035_, new_n2034_, keyIn_0_238 );
nand g1693 ( new_n2036_, new_n2035_, new_n2033_ );
nand g1694 ( new_n2037_, new_n2030_, new_n2036_ );
nor g1695 ( new_n2038_, new_n2037_, keyIn_0_246 );
nand g1696 ( new_n2039_, new_n2037_, keyIn_0_246 );
nand g1697 ( new_n2040_, new_n2039_, N219 );
nor g1698 ( new_n2041_, new_n2040_, new_n2038_ );
not g1699 ( new_n2042_, new_n2041_ );
nand g1700 ( new_n2043_, N96, N210 );
nand g1701 ( new_n2044_, new_n2042_, new_n2043_ );
nor g1702 ( new_n2045_, new_n2044_, new_n2000_ );
not g1703 ( new_n2046_, new_n2045_ );
not g1704 ( new_n2047_, new_n2043_ );
nor g1705 ( new_n2048_, new_n2041_, new_n2047_ );
nor g1706 ( new_n2049_, new_n2048_, keyIn_0_252 );
nor g1707 ( new_n2050_, new_n1645_, new_n1228_ );
not g1708 ( new_n2051_, new_n2050_ );
nand g1709 ( new_n2052_, new_n2051_, keyIn_0_170 );
not g1710 ( new_n2053_, new_n2052_ );
nor g1711 ( new_n2054_, new_n2051_, keyIn_0_170 );
nor g1712 ( new_n2055_, new_n2053_, new_n2054_ );
nor g1713 ( new_n2056_, new_n2008_, new_n1221_ );
nor g1714 ( new_n2057_, new_n2055_, new_n2056_ );
not g1715 ( new_n2058_, new_n2057_ );
nor g1716 ( new_n2059_, new_n2058_, keyIn_0_194 );
not g1717 ( new_n2060_, keyIn_0_149 );
not g1718 ( new_n2061_, keyIn_0_126 );
nor g1719 ( new_n2062_, new_n1636_, new_n956_ );
not g1720 ( new_n2063_, new_n2062_ );
nor g1721 ( new_n2064_, new_n2063_, new_n2061_ );
nor g1722 ( new_n2065_, new_n951_, new_n580_ );
nor g1723 ( new_n2066_, new_n2062_, keyIn_0_126 );
nor g1724 ( new_n2067_, new_n2066_, new_n2065_ );
not g1725 ( new_n2068_, new_n2067_ );
nor g1726 ( new_n2069_, new_n2068_, new_n2064_ );
not g1727 ( new_n2070_, new_n2069_ );
nand g1728 ( new_n2071_, new_n2070_, new_n2060_ );
nand g1729 ( new_n2072_, new_n2069_, keyIn_0_149 );
nand g1730 ( new_n2073_, new_n2071_, new_n2072_ );
nand g1731 ( new_n2074_, new_n2058_, keyIn_0_194 );
nand g1732 ( new_n2075_, new_n2074_, new_n2073_ );
nor g1733 ( new_n2076_, new_n2075_, new_n2059_ );
not g1734 ( new_n2077_, new_n2076_ );
nor g1735 ( new_n2078_, new_n2049_, new_n2077_ );
nand g1736 ( new_n2079_, new_n2046_, new_n2078_ );
nand g1737 ( new_n2080_, new_n2079_, keyIn_0_255 );
not g1738 ( new_n2081_, keyIn_0_255 );
nand g1739 ( new_n2082_, new_n2044_, new_n2000_ );
nand g1740 ( new_n2083_, new_n2082_, new_n2076_ );
nor g1741 ( new_n2084_, new_n2083_, new_n2045_ );
nand g1742 ( new_n2085_, new_n2084_, new_n2081_ );
nand g1743 ( N880, new_n2085_, new_n2080_ );
endmodule