module add_mul_combine_32_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, 
        a_18_, a_19_, a_20_, a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, 
        a_28_, a_29_, a_30_, a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, 
        b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, 
        b_17_, b_18_, b_19_, b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, 
        b_27_, b_28_, b_29_, b_30_, b_31_, Result_mul_0_, Result_mul_1_, 
        Result_mul_2_, Result_mul_3_, Result_mul_4_, Result_mul_5_, 
        Result_mul_6_, Result_mul_7_, Result_mul_8_, Result_mul_9_, 
        Result_mul_10_, Result_mul_11_, Result_mul_12_, Result_mul_13_, 
        Result_mul_14_, Result_mul_15_, Result_mul_16_, Result_mul_17_, 
        Result_mul_18_, Result_mul_19_, Result_mul_20_, Result_mul_21_, 
        Result_mul_22_, Result_mul_23_, Result_mul_24_, Result_mul_25_, 
        Result_mul_26_, Result_mul_27_, Result_mul_28_, Result_mul_29_, 
        Result_mul_30_, Result_mul_31_, Result_mul_32_, Result_mul_33_, 
        Result_mul_34_, Result_mul_35_, Result_mul_36_, Result_mul_37_, 
        Result_mul_38_, Result_mul_39_, Result_mul_40_, Result_mul_41_, 
        Result_mul_42_, Result_mul_43_, Result_mul_44_, Result_mul_45_, 
        Result_mul_46_, Result_mul_47_, Result_mul_48_, Result_mul_49_, 
        Result_mul_50_, Result_mul_51_, Result_mul_52_, Result_mul_53_, 
        Result_mul_54_, Result_mul_55_, Result_mul_56_, Result_mul_57_, 
        Result_mul_58_, Result_mul_59_, Result_mul_60_, Result_mul_61_, 
        Result_mul_62_, Result_mul_63_, Result_add_0_, Result_add_1_, 
        Result_add_2_, Result_add_3_, Result_add_4_, Result_add_5_, 
        Result_add_6_, Result_add_7_, Result_add_8_, Result_add_9_, 
        Result_add_10_, Result_add_11_, Result_add_12_, Result_add_13_, 
        Result_add_14_, Result_add_15_, Result_add_16_, Result_add_17_, 
        Result_add_18_, Result_add_19_, Result_add_20_, Result_add_21_, 
        Result_add_22_, Result_add_23_, Result_add_24_, Result_add_25_, 
        Result_add_26_, Result_add_27_, Result_add_28_, Result_add_29_, 
        Result_add_30_, Result_add_31_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, a_19_, a_20_,
         a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, a_29_, a_30_,
         a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_,
         b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, b_18_, b_19_,
         b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, b_28_, b_29_,
         b_30_, b_31_;
  output Result_mul_0_, Result_mul_1_, Result_mul_2_, Result_mul_3_,
         Result_mul_4_, Result_mul_5_, Result_mul_6_, Result_mul_7_,
         Result_mul_8_, Result_mul_9_, Result_mul_10_, Result_mul_11_,
         Result_mul_12_, Result_mul_13_, Result_mul_14_, Result_mul_15_,
         Result_mul_16_, Result_mul_17_, Result_mul_18_, Result_mul_19_,
         Result_mul_20_, Result_mul_21_, Result_mul_22_, Result_mul_23_,
         Result_mul_24_, Result_mul_25_, Result_mul_26_, Result_mul_27_,
         Result_mul_28_, Result_mul_29_, Result_mul_30_, Result_mul_31_,
         Result_mul_32_, Result_mul_33_, Result_mul_34_, Result_mul_35_,
         Result_mul_36_, Result_mul_37_, Result_mul_38_, Result_mul_39_,
         Result_mul_40_, Result_mul_41_, Result_mul_42_, Result_mul_43_,
         Result_mul_44_, Result_mul_45_, Result_mul_46_, Result_mul_47_,
         Result_mul_48_, Result_mul_49_, Result_mul_50_, Result_mul_51_,
         Result_mul_52_, Result_mul_53_, Result_mul_54_, Result_mul_55_,
         Result_mul_56_, Result_mul_57_, Result_mul_58_, Result_mul_59_,
         Result_mul_60_, Result_mul_61_, Result_mul_62_, Result_mul_63_,
         Result_add_0_, Result_add_1_, Result_add_2_, Result_add_3_,
         Result_add_4_, Result_add_5_, Result_add_6_, Result_add_7_,
         Result_add_8_, Result_add_9_, Result_add_10_, Result_add_11_,
         Result_add_12_, Result_add_13_, Result_add_14_, Result_add_15_,
         Result_add_16_, Result_add_17_, Result_add_18_, Result_add_19_,
         Result_add_20_, Result_add_21_, Result_add_22_, Result_add_23_,
         Result_add_24_, Result_add_25_, Result_add_26_, Result_add_27_,
         Result_add_28_, Result_add_29_, Result_add_30_, Result_add_31_;
  wire   n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301;

  NAND2_X2 U7404 ( .A1(a_31_), .A2(a_30_), .ZN(n8055) );
  INV_X2 U7405 ( .A(b_19_), .ZN(n10207) );
  INV_X2 U7406 ( .A(b_21_), .ZN(n9734) );
  INV_X2 U7407 ( .A(b_27_), .ZN(n8292) );
  INV_X2 U7408 ( .A(b_10_), .ZN(n12422) );
  INV_X2 U7409 ( .A(a_31_), .ZN(n7817) );
  INV_X2 U7410 ( .A(b_17_), .ZN(n10693) );
  INV_X2 U7411 ( .A(b_3_), .ZN(n14110) );
  INV_X2 U7412 ( .A(a_2_), .ZN(n7469) );
  INV_X2 U7413 ( .A(a_25_), .ZN(n8022) );
  INV_X2 U7414 ( .A(a_28_), .ZN(n7803) );
  INV_X2 U7415 ( .A(a_3_), .ZN(n7464) );
  INV_X2 U7416 ( .A(n7332), .ZN(n7810) );
  INV_X2 U7417 ( .A(n7328), .ZN(n7816) );
  INV_X2 U7418 ( .A(a_6_), .ZN(n7450) );
  INV_X2 U7419 ( .A(a_4_), .ZN(n7682) );
  INV_X2 U7420 ( .A(a_9_), .ZN(n7704) );
  INV_X2 U7421 ( .A(a_19_), .ZN(n7750) );
  INV_X2 U7422 ( .A(a_30_), .ZN(n8052) );
  INV_X2 U7423 ( .A(b_0_), .ZN(n14859) );
  INV_X2 U7424 ( .A(b_6_), .ZN(n13377) );
  INV_X2 U7425 ( .A(a_17_), .ZN(n7397) );
  INV_X2 U7426 ( .A(a_7_), .ZN(n7445) );
  INV_X2 U7427 ( .A(a_22_), .ZN(n7765) );
  INV_X2 U7428 ( .A(a_1_), .ZN(n7669) );
  INV_X2 U7429 ( .A(a_13_), .ZN(n7415) );
  INV_X2 U7430 ( .A(a_15_), .ZN(n7406) );
  INV_X2 U7431 ( .A(b_8_), .ZN(n12909) );
  INV_X2 U7432 ( .A(a_29_), .ZN(n7337) );
  INV_X2 U7433 ( .A(a_12_), .ZN(n7718) );
  INV_X2 U7434 ( .A(a_14_), .ZN(n7727) );
  INV_X2 U7435 ( .A(a_5_), .ZN(n7455) );
  INV_X2 U7436 ( .A(a_10_), .ZN(n7709) );
  INV_X2 U7437 ( .A(b_4_), .ZN(n13861) );
  INV_X2 U7438 ( .A(a_23_), .ZN(n8014) );
  INV_X2 U7439 ( .A(a_24_), .ZN(n7774) );
  INV_X2 U7440 ( .A(a_8_), .ZN(n7699) );
  INV_X2 U7441 ( .A(a_21_), .ZN(n7760) );
  INV_X2 U7442 ( .A(a_11_), .ZN(n7424) );
  INV_X2 U7443 ( .A(a_16_), .ZN(n7736) );
  INV_X2 U7444 ( .A(b_1_), .ZN(n14645) );
  INV_X2 U7445 ( .A(b_7_), .ZN(n13127) );
  INV_X2 U7446 ( .A(a_0_), .ZN(n7478) );
  INV_X2 U7447 ( .A(a_18_), .ZN(n7745) );
  INV_X2 U7448 ( .A(b_11_), .ZN(n12145) );
  INV_X2 U7449 ( .A(b_9_), .ZN(n12638) );
  INV_X2 U7450 ( .A(b_5_), .ZN(n13620) );
  INV_X2 U7451 ( .A(a_20_), .ZN(n7755) );
  XOR2_X1 U7452 ( .A(n7309), .B(n7310), .Z(Result_mul_9_) );
  AND2_X1 U7453 ( .A1(n7311), .A2(n7312), .ZN(n7310) );
  XOR2_X1 U7454 ( .A(n7313), .B(n7314), .Z(Result_mul_8_) );
  AND2_X1 U7455 ( .A1(n7315), .A2(n7316), .ZN(n7314) );
  XOR2_X1 U7456 ( .A(n7317), .B(n7318), .Z(Result_mul_7_) );
  AND2_X1 U7457 ( .A1(n7319), .A2(n7320), .ZN(n7318) );
  XOR2_X1 U7458 ( .A(n7321), .B(n7322), .Z(Result_mul_6_) );
  AND2_X1 U7459 ( .A1(n7323), .A2(n7324), .ZN(n7322) );
  NAND2_X1 U7460 ( .A1(n7325), .A2(n7326), .ZN(Result_mul_62_) );
  NAND2_X1 U7461 ( .A1(b_30_), .A2(n7327), .ZN(n7326) );
  NAND2_X1 U7462 ( .A1(n7328), .A2(n7329), .ZN(n7327) );
  NAND2_X1 U7463 ( .A1(a_31_), .A2(n7330), .ZN(n7329) );
  NAND2_X1 U7464 ( .A1(b_31_), .A2(n7331), .ZN(n7325) );
  NAND2_X1 U7465 ( .A1(n7332), .A2(n7333), .ZN(n7331) );
  NAND2_X1 U7466 ( .A1(a_30_), .A2(n7334), .ZN(n7333) );
  XOR2_X1 U7467 ( .A(n7335), .B(n7336), .Z(Result_mul_61_) );
  NOR2_X1 U7468 ( .A1(n7337), .A2(n7330), .ZN(n7336) );
  XOR2_X1 U7469 ( .A(n7338), .B(n7339), .Z(n7335) );
  XOR2_X1 U7470 ( .A(n7340), .B(n7341), .Z(Result_mul_60_) );
  XNOR2_X1 U7471 ( .A(n7342), .B(n7343), .ZN(n7341) );
  NAND2_X1 U7472 ( .A1(b_31_), .A2(a_28_), .ZN(n7342) );
  XOR2_X1 U7473 ( .A(n7344), .B(n7345), .Z(Result_mul_5_) );
  AND2_X1 U7474 ( .A1(n7346), .A2(n7347), .ZN(n7345) );
  XNOR2_X1 U7475 ( .A(n7348), .B(n7349), .ZN(Result_mul_59_) );
  NAND2_X1 U7476 ( .A1(n7350), .A2(n7351), .ZN(n7348) );
  XOR2_X1 U7477 ( .A(n7352), .B(n7353), .Z(Result_mul_58_) );
  XOR2_X1 U7478 ( .A(n7354), .B(n7355), .Z(n7352) );
  NOR2_X1 U7479 ( .A1(n7356), .A2(n7330), .ZN(n7355) );
  XNOR2_X1 U7480 ( .A(n7357), .B(n7358), .ZN(Result_mul_57_) );
  NAND2_X1 U7481 ( .A1(n7359), .A2(n7360), .ZN(n7357) );
  XNOR2_X1 U7482 ( .A(n7361), .B(n7362), .ZN(Result_mul_56_) );
  XOR2_X1 U7483 ( .A(n7363), .B(n7364), .Z(n7362) );
  NAND2_X1 U7484 ( .A1(b_31_), .A2(a_24_), .ZN(n7364) );
  XNOR2_X1 U7485 ( .A(n7365), .B(n7366), .ZN(Result_mul_55_) );
  NAND2_X1 U7486 ( .A1(n7367), .A2(n7368), .ZN(n7365) );
  XNOR2_X1 U7487 ( .A(n7369), .B(n7370), .ZN(Result_mul_54_) );
  XOR2_X1 U7488 ( .A(n7371), .B(n7372), .Z(n7370) );
  NAND2_X1 U7489 ( .A1(b_31_), .A2(a_22_), .ZN(n7372) );
  XNOR2_X1 U7490 ( .A(n7373), .B(n7374), .ZN(Result_mul_53_) );
  XOR2_X1 U7491 ( .A(n7375), .B(n7376), .Z(n7374) );
  NAND2_X1 U7492 ( .A1(b_31_), .A2(a_21_), .ZN(n7376) );
  XNOR2_X1 U7493 ( .A(n7377), .B(n7378), .ZN(Result_mul_52_) );
  XOR2_X1 U7494 ( .A(n7379), .B(n7380), .Z(n7378) );
  NAND2_X1 U7495 ( .A1(b_31_), .A2(a_20_), .ZN(n7380) );
  XNOR2_X1 U7496 ( .A(n7381), .B(n7382), .ZN(Result_mul_51_) );
  XOR2_X1 U7497 ( .A(n7383), .B(n7384), .Z(n7382) );
  NAND2_X1 U7498 ( .A1(b_31_), .A2(a_19_), .ZN(n7384) );
  XNOR2_X1 U7499 ( .A(n7385), .B(n7386), .ZN(Result_mul_50_) );
  XOR2_X1 U7500 ( .A(n7387), .B(n7388), .Z(n7386) );
  NAND2_X1 U7501 ( .A1(b_31_), .A2(a_18_), .ZN(n7388) );
  XOR2_X1 U7502 ( .A(n7389), .B(n7390), .Z(Result_mul_4_) );
  AND2_X1 U7503 ( .A1(n7391), .A2(n7392), .ZN(n7390) );
  XOR2_X1 U7504 ( .A(n7393), .B(n7394), .Z(Result_mul_49_) );
  XOR2_X1 U7505 ( .A(n7395), .B(n7396), .Z(n7393) );
  NOR2_X1 U7506 ( .A1(n7397), .A2(n7330), .ZN(n7396) );
  XNOR2_X1 U7507 ( .A(n7398), .B(n7399), .ZN(Result_mul_48_) );
  XOR2_X1 U7508 ( .A(n7400), .B(n7401), .Z(n7399) );
  NAND2_X1 U7509 ( .A1(b_31_), .A2(a_16_), .ZN(n7401) );
  XOR2_X1 U7510 ( .A(n7402), .B(n7403), .Z(Result_mul_47_) );
  XOR2_X1 U7511 ( .A(n7404), .B(n7405), .Z(n7402) );
  NOR2_X1 U7512 ( .A1(n7406), .A2(n7330), .ZN(n7405) );
  XNOR2_X1 U7513 ( .A(n7407), .B(n7408), .ZN(Result_mul_46_) );
  XOR2_X1 U7514 ( .A(n7409), .B(n7410), .Z(n7408) );
  NAND2_X1 U7515 ( .A1(b_31_), .A2(a_14_), .ZN(n7410) );
  XOR2_X1 U7516 ( .A(n7411), .B(n7412), .Z(Result_mul_45_) );
  XOR2_X1 U7517 ( .A(n7413), .B(n7414), .Z(n7411) );
  NOR2_X1 U7518 ( .A1(n7415), .A2(n7330), .ZN(n7414) );
  XNOR2_X1 U7519 ( .A(n7416), .B(n7417), .ZN(Result_mul_44_) );
  XOR2_X1 U7520 ( .A(n7418), .B(n7419), .Z(n7417) );
  NAND2_X1 U7521 ( .A1(b_31_), .A2(a_12_), .ZN(n7419) );
  XOR2_X1 U7522 ( .A(n7420), .B(n7421), .Z(Result_mul_43_) );
  XOR2_X1 U7523 ( .A(n7422), .B(n7423), .Z(n7420) );
  NOR2_X1 U7524 ( .A1(n7424), .A2(n7330), .ZN(n7423) );
  XNOR2_X1 U7525 ( .A(n7425), .B(n7426), .ZN(Result_mul_42_) );
  XOR2_X1 U7526 ( .A(n7427), .B(n7428), .Z(n7426) );
  NAND2_X1 U7527 ( .A1(b_31_), .A2(a_10_), .ZN(n7428) );
  XNOR2_X1 U7528 ( .A(n7429), .B(n7430), .ZN(Result_mul_41_) );
  XOR2_X1 U7529 ( .A(n7431), .B(n7432), .Z(n7430) );
  NAND2_X1 U7530 ( .A1(b_31_), .A2(a_9_), .ZN(n7432) );
  XNOR2_X1 U7531 ( .A(n7433), .B(n7434), .ZN(Result_mul_40_) );
  XOR2_X1 U7532 ( .A(n7435), .B(n7436), .Z(n7434) );
  NAND2_X1 U7533 ( .A1(b_31_), .A2(a_8_), .ZN(n7436) );
  XOR2_X1 U7534 ( .A(n7437), .B(n7438), .Z(Result_mul_3_) );
  AND2_X1 U7535 ( .A1(n7439), .A2(n7440), .ZN(n7438) );
  XOR2_X1 U7536 ( .A(n7441), .B(n7442), .Z(Result_mul_39_) );
  XOR2_X1 U7537 ( .A(n7443), .B(n7444), .Z(n7441) );
  NOR2_X1 U7538 ( .A1(n7445), .A2(n7330), .ZN(n7444) );
  XOR2_X1 U7539 ( .A(n7446), .B(n7447), .Z(Result_mul_38_) );
  XOR2_X1 U7540 ( .A(n7448), .B(n7449), .Z(n7446) );
  NOR2_X1 U7541 ( .A1(n7450), .A2(n7330), .ZN(n7449) );
  XOR2_X1 U7542 ( .A(n7451), .B(n7452), .Z(Result_mul_37_) );
  XOR2_X1 U7543 ( .A(n7453), .B(n7454), .Z(n7451) );
  NOR2_X1 U7544 ( .A1(n7455), .A2(n7330), .ZN(n7454) );
  XNOR2_X1 U7545 ( .A(n7456), .B(n7457), .ZN(Result_mul_36_) );
  XOR2_X1 U7546 ( .A(n7458), .B(n7459), .Z(n7457) );
  NAND2_X1 U7547 ( .A1(b_31_), .A2(a_4_), .ZN(n7459) );
  XOR2_X1 U7548 ( .A(n7460), .B(n7461), .Z(Result_mul_35_) );
  XOR2_X1 U7549 ( .A(n7462), .B(n7463), .Z(n7460) );
  NOR2_X1 U7550 ( .A1(n7464), .A2(n7330), .ZN(n7463) );
  XOR2_X1 U7551 ( .A(n7465), .B(n7466), .Z(Result_mul_34_) );
  XOR2_X1 U7552 ( .A(n7467), .B(n7468), .Z(n7465) );
  NOR2_X1 U7553 ( .A1(n7469), .A2(n7330), .ZN(n7468) );
  XNOR2_X1 U7554 ( .A(n7470), .B(n7471), .ZN(Result_mul_33_) );
  XOR2_X1 U7555 ( .A(n7472), .B(n7473), .Z(n7471) );
  NAND2_X1 U7556 ( .A1(b_31_), .A2(a_1_), .ZN(n7473) );
  XOR2_X1 U7557 ( .A(n7474), .B(n7475), .Z(Result_mul_32_) );
  XOR2_X1 U7558 ( .A(n7476), .B(n7477), .Z(n7474) );
  NOR2_X1 U7559 ( .A1(n7478), .A2(n7330), .ZN(n7477) );
  INV_X1 U7560 ( .A(b_31_), .ZN(n7330) );
  XOR2_X1 U7561 ( .A(n7479), .B(n7480), .Z(Result_mul_31_) );
  NOR2_X1 U7562 ( .A1(n7481), .A2(n7482), .ZN(Result_mul_30_) );
  NOR2_X1 U7563 ( .A1(n7483), .A2(n7484), .ZN(n7482) );
  XOR2_X1 U7564 ( .A(n7485), .B(n7486), .Z(Result_mul_2_) );
  AND2_X1 U7565 ( .A1(n7487), .A2(n7488), .ZN(n7486) );
  XNOR2_X1 U7566 ( .A(n7481), .B(n7489), .ZN(Result_mul_29_) );
  NAND2_X1 U7567 ( .A1(n7490), .A2(n7491), .ZN(n7489) );
  XNOR2_X1 U7568 ( .A(n7492), .B(n7493), .ZN(Result_mul_28_) );
  NAND2_X1 U7569 ( .A1(n7494), .A2(n7495), .ZN(n7492) );
  XOR2_X1 U7570 ( .A(n7496), .B(n7497), .Z(Result_mul_27_) );
  AND2_X1 U7571 ( .A1(n7498), .A2(n7499), .ZN(n7497) );
  XOR2_X1 U7572 ( .A(n7500), .B(n7501), .Z(Result_mul_26_) );
  AND2_X1 U7573 ( .A1(n7502), .A2(n7503), .ZN(n7501) );
  XOR2_X1 U7574 ( .A(n7504), .B(n7505), .Z(Result_mul_25_) );
  AND2_X1 U7575 ( .A1(n7506), .A2(n7507), .ZN(n7505) );
  XOR2_X1 U7576 ( .A(n7508), .B(n7509), .Z(Result_mul_24_) );
  AND2_X1 U7577 ( .A1(n7510), .A2(n7511), .ZN(n7509) );
  XOR2_X1 U7578 ( .A(n7512), .B(n7513), .Z(Result_mul_23_) );
  AND2_X1 U7579 ( .A1(n7514), .A2(n7515), .ZN(n7513) );
  XOR2_X1 U7580 ( .A(n7516), .B(n7517), .Z(Result_mul_22_) );
  AND2_X1 U7581 ( .A1(n7518), .A2(n7519), .ZN(n7517) );
  XOR2_X1 U7582 ( .A(n7520), .B(n7521), .Z(Result_mul_21_) );
  AND2_X1 U7583 ( .A1(n7522), .A2(n7523), .ZN(n7521) );
  XOR2_X1 U7584 ( .A(n7524), .B(n7525), .Z(Result_mul_20_) );
  AND2_X1 U7585 ( .A1(n7526), .A2(n7527), .ZN(n7525) );
  XOR2_X1 U7586 ( .A(n7528), .B(n7529), .Z(Result_mul_1_) );
  NOR2_X1 U7587 ( .A1(n7530), .A2(n7531), .ZN(n7529) );
  INV_X1 U7588 ( .A(n7532), .ZN(n7530) );
  XOR2_X1 U7589 ( .A(n7533), .B(n7534), .Z(Result_mul_19_) );
  AND2_X1 U7590 ( .A1(n7535), .A2(n7536), .ZN(n7534) );
  XOR2_X1 U7591 ( .A(n7537), .B(n7538), .Z(Result_mul_18_) );
  AND2_X1 U7592 ( .A1(n7539), .A2(n7540), .ZN(n7538) );
  XOR2_X1 U7593 ( .A(n7541), .B(n7542), .Z(Result_mul_17_) );
  AND2_X1 U7594 ( .A1(n7543), .A2(n7544), .ZN(n7542) );
  XOR2_X1 U7595 ( .A(n7545), .B(n7546), .Z(Result_mul_16_) );
  AND2_X1 U7596 ( .A1(n7547), .A2(n7548), .ZN(n7546) );
  XOR2_X1 U7597 ( .A(n7549), .B(n7550), .Z(Result_mul_15_) );
  AND2_X1 U7598 ( .A1(n7551), .A2(n7552), .ZN(n7550) );
  XOR2_X1 U7599 ( .A(n7553), .B(n7554), .Z(Result_mul_14_) );
  AND2_X1 U7600 ( .A1(n7555), .A2(n7556), .ZN(n7554) );
  XOR2_X1 U7601 ( .A(n7557), .B(n7558), .Z(Result_mul_13_) );
  AND2_X1 U7602 ( .A1(n7559), .A2(n7560), .ZN(n7558) );
  XOR2_X1 U7603 ( .A(n7561), .B(n7562), .Z(Result_mul_12_) );
  AND2_X1 U7604 ( .A1(n7563), .A2(n7564), .ZN(n7562) );
  XOR2_X1 U7605 ( .A(n7565), .B(n7566), .Z(Result_mul_11_) );
  AND2_X1 U7606 ( .A1(n7567), .A2(n7568), .ZN(n7566) );
  XOR2_X1 U7607 ( .A(n7569), .B(n7570), .Z(Result_mul_10_) );
  AND2_X1 U7608 ( .A1(n7571), .A2(n7572), .ZN(n7570) );
  NAND2_X1 U7609 ( .A1(n7573), .A2(n7574), .ZN(Result_mul_0_) );
  NAND2_X1 U7610 ( .A1(n7532), .A2(n7528), .ZN(n7574) );
  NAND2_X1 U7611 ( .A1(n7488), .A2(n7575), .ZN(n7528) );
  NAND2_X1 U7612 ( .A1(n7487), .A2(n7485), .ZN(n7575) );
  NAND2_X1 U7613 ( .A1(n7439), .A2(n7576), .ZN(n7485) );
  NAND2_X1 U7614 ( .A1(n7440), .A2(n7437), .ZN(n7576) );
  NAND2_X1 U7615 ( .A1(n7392), .A2(n7577), .ZN(n7437) );
  NAND2_X1 U7616 ( .A1(n7391), .A2(n7389), .ZN(n7577) );
  NAND2_X1 U7617 ( .A1(n7346), .A2(n7578), .ZN(n7389) );
  NAND2_X1 U7618 ( .A1(n7347), .A2(n7344), .ZN(n7578) );
  NAND2_X1 U7619 ( .A1(n7324), .A2(n7579), .ZN(n7344) );
  NAND2_X1 U7620 ( .A1(n7323), .A2(n7321), .ZN(n7579) );
  NAND2_X1 U7621 ( .A1(n7319), .A2(n7580), .ZN(n7321) );
  NAND2_X1 U7622 ( .A1(n7320), .A2(n7317), .ZN(n7580) );
  NAND2_X1 U7623 ( .A1(n7316), .A2(n7581), .ZN(n7317) );
  NAND2_X1 U7624 ( .A1(n7315), .A2(n7313), .ZN(n7581) );
  NAND2_X1 U7625 ( .A1(n7311), .A2(n7582), .ZN(n7313) );
  NAND2_X1 U7626 ( .A1(n7312), .A2(n7309), .ZN(n7582) );
  NAND2_X1 U7627 ( .A1(n7572), .A2(n7583), .ZN(n7309) );
  NAND2_X1 U7628 ( .A1(n7569), .A2(n7571), .ZN(n7583) );
  NAND2_X1 U7629 ( .A1(n7584), .A2(n7585), .ZN(n7571) );
  NAND2_X1 U7630 ( .A1(n7567), .A2(n7586), .ZN(n7569) );
  NAND2_X1 U7631 ( .A1(n7565), .A2(n7568), .ZN(n7586) );
  NAND2_X1 U7632 ( .A1(n7587), .A2(n7588), .ZN(n7568) );
  NAND2_X1 U7633 ( .A1(n7564), .A2(n7589), .ZN(n7565) );
  NAND2_X1 U7634 ( .A1(n7561), .A2(n7563), .ZN(n7589) );
  NAND2_X1 U7635 ( .A1(n7590), .A2(n7591), .ZN(n7563) );
  XNOR2_X1 U7636 ( .A(n7592), .B(n7593), .ZN(n7590) );
  NAND2_X1 U7637 ( .A1(n7559), .A2(n7594), .ZN(n7561) );
  NAND2_X1 U7638 ( .A1(n7557), .A2(n7560), .ZN(n7594) );
  NAND2_X1 U7639 ( .A1(n7595), .A2(n7596), .ZN(n7560) );
  NAND2_X1 U7640 ( .A1(n7556), .A2(n7597), .ZN(n7557) );
  NAND2_X1 U7641 ( .A1(n7555), .A2(n7553), .ZN(n7597) );
  NAND2_X1 U7642 ( .A1(n7552), .A2(n7598), .ZN(n7553) );
  NAND2_X1 U7643 ( .A1(n7551), .A2(n7549), .ZN(n7598) );
  NAND2_X1 U7644 ( .A1(n7548), .A2(n7599), .ZN(n7549) );
  NAND2_X1 U7645 ( .A1(n7545), .A2(n7547), .ZN(n7599) );
  NAND2_X1 U7646 ( .A1(n7600), .A2(n7601), .ZN(n7547) );
  NAND2_X1 U7647 ( .A1(n7602), .A2(n7603), .ZN(n7601) );
  XOR2_X1 U7648 ( .A(n7604), .B(n7605), .Z(n7600) );
  NAND2_X1 U7649 ( .A1(n7544), .A2(n7606), .ZN(n7545) );
  NAND2_X1 U7650 ( .A1(n7543), .A2(n7541), .ZN(n7606) );
  NAND2_X1 U7651 ( .A1(n7539), .A2(n7607), .ZN(n7541) );
  NAND2_X1 U7652 ( .A1(n7537), .A2(n7540), .ZN(n7607) );
  NAND2_X1 U7653 ( .A1(n7608), .A2(n7609), .ZN(n7540) );
  NAND2_X1 U7654 ( .A1(n7610), .A2(n7611), .ZN(n7609) );
  XOR2_X1 U7655 ( .A(n7612), .B(n7613), .Z(n7608) );
  NAND2_X1 U7656 ( .A1(n7536), .A2(n7614), .ZN(n7537) );
  NAND2_X1 U7657 ( .A1(n7533), .A2(n7535), .ZN(n7614) );
  NAND2_X1 U7658 ( .A1(n7615), .A2(n7616), .ZN(n7535) );
  NAND2_X1 U7659 ( .A1(n7617), .A2(n7618), .ZN(n7616) );
  XNOR2_X1 U7660 ( .A(n7611), .B(n7610), .ZN(n7615) );
  NAND2_X1 U7661 ( .A1(n7527), .A2(n7619), .ZN(n7533) );
  NAND2_X1 U7662 ( .A1(n7524), .A2(n7526), .ZN(n7619) );
  NAND2_X1 U7663 ( .A1(n7620), .A2(n7621), .ZN(n7526) );
  NAND2_X1 U7664 ( .A1(n7522), .A2(n7622), .ZN(n7524) );
  NAND2_X1 U7665 ( .A1(n7523), .A2(n7520), .ZN(n7622) );
  NAND2_X1 U7666 ( .A1(n7518), .A2(n7623), .ZN(n7520) );
  NAND2_X1 U7667 ( .A1(n7516), .A2(n7519), .ZN(n7623) );
  NAND2_X1 U7668 ( .A1(n7624), .A2(n7625), .ZN(n7519) );
  NAND2_X1 U7669 ( .A1(n7626), .A2(n7627), .ZN(n7625) );
  XNOR2_X1 U7670 ( .A(n7628), .B(n7629), .ZN(n7624) );
  NAND2_X1 U7671 ( .A1(n7515), .A2(n7630), .ZN(n7516) );
  NAND2_X1 U7672 ( .A1(n7512), .A2(n7514), .ZN(n7630) );
  NAND2_X1 U7673 ( .A1(n7631), .A2(n7632), .ZN(n7514) );
  NAND2_X1 U7674 ( .A1(n7633), .A2(n7634), .ZN(n7632) );
  XOR2_X1 U7675 ( .A(n7627), .B(n7635), .Z(n7631) );
  NAND2_X1 U7676 ( .A1(n7511), .A2(n7636), .ZN(n7512) );
  NAND2_X1 U7677 ( .A1(n7508), .A2(n7510), .ZN(n7636) );
  NAND2_X1 U7678 ( .A1(n7637), .A2(n7638), .ZN(n7510) );
  NAND2_X1 U7679 ( .A1(n7506), .A2(n7639), .ZN(n7508) );
  NAND2_X1 U7680 ( .A1(n7507), .A2(n7504), .ZN(n7639) );
  NAND2_X1 U7681 ( .A1(n7640), .A2(n7502), .ZN(n7504) );
  NAND2_X1 U7682 ( .A1(n7641), .A2(n7642), .ZN(n7502) );
  XOR2_X1 U7683 ( .A(n7643), .B(n7644), .Z(n7641) );
  NAND2_X1 U7684 ( .A1(n7503), .A2(n7500), .ZN(n7640) );
  NAND2_X1 U7685 ( .A1(n7499), .A2(n7645), .ZN(n7500) );
  NAND2_X1 U7686 ( .A1(n7498), .A2(n7496), .ZN(n7645) );
  NAND2_X1 U7687 ( .A1(n7494), .A2(n7646), .ZN(n7496) );
  NAND2_X1 U7688 ( .A1(n7493), .A2(n7495), .ZN(n7646) );
  NAND2_X1 U7689 ( .A1(n7647), .A2(n7648), .ZN(n7495) );
  NAND2_X1 U7690 ( .A1(n7649), .A2(n7650), .ZN(n7648) );
  NAND2_X1 U7691 ( .A1(n7491), .A2(n7651), .ZN(n7493) );
  NAND2_X1 U7692 ( .A1(n7481), .A2(n7490), .ZN(n7651) );
  NAND2_X1 U7693 ( .A1(n7652), .A2(n7653), .ZN(n7490) );
  NAND2_X1 U7694 ( .A1(n7654), .A2(n7655), .ZN(n7653) );
  XOR2_X1 U7695 ( .A(n7656), .B(n7649), .Z(n7652) );
  AND2_X1 U7696 ( .A1(n7483), .A2(n7484), .ZN(n7481) );
  XOR2_X1 U7697 ( .A(n7655), .B(n7654), .Z(n7484) );
  NOR2_X1 U7698 ( .A1(n7479), .A2(n7480), .ZN(n7483) );
  XNOR2_X1 U7699 ( .A(n7657), .B(n7658), .ZN(n7480) );
  XOR2_X1 U7700 ( .A(n7659), .B(n7660), .Z(n7657) );
  NOR2_X1 U7701 ( .A1(n7478), .A2(n7334), .ZN(n7660) );
  AND2_X1 U7702 ( .A1(n7661), .A2(n7662), .ZN(n7479) );
  NAND2_X1 U7703 ( .A1(n7663), .A2(b_31_), .ZN(n7662) );
  NOR2_X1 U7704 ( .A1(n7664), .A2(n7478), .ZN(n7663) );
  NOR2_X1 U7705 ( .A1(n7475), .A2(n7476), .ZN(n7664) );
  NAND2_X1 U7706 ( .A1(n7475), .A2(n7476), .ZN(n7661) );
  NAND2_X1 U7707 ( .A1(n7665), .A2(n7666), .ZN(n7476) );
  NAND2_X1 U7708 ( .A1(n7667), .A2(b_31_), .ZN(n7666) );
  NOR2_X1 U7709 ( .A1(n7668), .A2(n7669), .ZN(n7667) );
  NOR2_X1 U7710 ( .A1(n7470), .A2(n7472), .ZN(n7668) );
  NAND2_X1 U7711 ( .A1(n7470), .A2(n7472), .ZN(n7665) );
  NAND2_X1 U7712 ( .A1(n7670), .A2(n7671), .ZN(n7472) );
  NAND2_X1 U7713 ( .A1(n7672), .A2(b_31_), .ZN(n7671) );
  NOR2_X1 U7714 ( .A1(n7673), .A2(n7469), .ZN(n7672) );
  NOR2_X1 U7715 ( .A1(n7466), .A2(n7467), .ZN(n7673) );
  NAND2_X1 U7716 ( .A1(n7466), .A2(n7467), .ZN(n7670) );
  NAND2_X1 U7717 ( .A1(n7674), .A2(n7675), .ZN(n7467) );
  NAND2_X1 U7718 ( .A1(n7676), .A2(b_31_), .ZN(n7675) );
  NOR2_X1 U7719 ( .A1(n7677), .A2(n7464), .ZN(n7676) );
  NOR2_X1 U7720 ( .A1(n7461), .A2(n7462), .ZN(n7677) );
  NAND2_X1 U7721 ( .A1(n7461), .A2(n7462), .ZN(n7674) );
  NAND2_X1 U7722 ( .A1(n7678), .A2(n7679), .ZN(n7462) );
  NAND2_X1 U7723 ( .A1(n7680), .A2(b_31_), .ZN(n7679) );
  NOR2_X1 U7724 ( .A1(n7681), .A2(n7682), .ZN(n7680) );
  NOR2_X1 U7725 ( .A1(n7456), .A2(n7458), .ZN(n7681) );
  NAND2_X1 U7726 ( .A1(n7456), .A2(n7458), .ZN(n7678) );
  NAND2_X1 U7727 ( .A1(n7683), .A2(n7684), .ZN(n7458) );
  NAND2_X1 U7728 ( .A1(n7685), .A2(b_31_), .ZN(n7684) );
  NOR2_X1 U7729 ( .A1(n7686), .A2(n7455), .ZN(n7685) );
  NOR2_X1 U7730 ( .A1(n7452), .A2(n7453), .ZN(n7686) );
  NAND2_X1 U7731 ( .A1(n7452), .A2(n7453), .ZN(n7683) );
  NAND2_X1 U7732 ( .A1(n7687), .A2(n7688), .ZN(n7453) );
  NAND2_X1 U7733 ( .A1(n7689), .A2(b_31_), .ZN(n7688) );
  NOR2_X1 U7734 ( .A1(n7690), .A2(n7450), .ZN(n7689) );
  NOR2_X1 U7735 ( .A1(n7447), .A2(n7448), .ZN(n7690) );
  NAND2_X1 U7736 ( .A1(n7447), .A2(n7448), .ZN(n7687) );
  NAND2_X1 U7737 ( .A1(n7691), .A2(n7692), .ZN(n7448) );
  NAND2_X1 U7738 ( .A1(n7693), .A2(b_31_), .ZN(n7692) );
  NOR2_X1 U7739 ( .A1(n7694), .A2(n7445), .ZN(n7693) );
  NOR2_X1 U7740 ( .A1(n7442), .A2(n7443), .ZN(n7694) );
  NAND2_X1 U7741 ( .A1(n7442), .A2(n7443), .ZN(n7691) );
  NAND2_X1 U7742 ( .A1(n7695), .A2(n7696), .ZN(n7443) );
  NAND2_X1 U7743 ( .A1(n7697), .A2(b_31_), .ZN(n7696) );
  NOR2_X1 U7744 ( .A1(n7698), .A2(n7699), .ZN(n7697) );
  NOR2_X1 U7745 ( .A1(n7433), .A2(n7435), .ZN(n7698) );
  NAND2_X1 U7746 ( .A1(n7433), .A2(n7435), .ZN(n7695) );
  NAND2_X1 U7747 ( .A1(n7700), .A2(n7701), .ZN(n7435) );
  NAND2_X1 U7748 ( .A1(n7702), .A2(b_31_), .ZN(n7701) );
  NOR2_X1 U7749 ( .A1(n7703), .A2(n7704), .ZN(n7702) );
  NOR2_X1 U7750 ( .A1(n7429), .A2(n7431), .ZN(n7703) );
  NAND2_X1 U7751 ( .A1(n7429), .A2(n7431), .ZN(n7700) );
  NAND2_X1 U7752 ( .A1(n7705), .A2(n7706), .ZN(n7431) );
  NAND2_X1 U7753 ( .A1(n7707), .A2(b_31_), .ZN(n7706) );
  NOR2_X1 U7754 ( .A1(n7708), .A2(n7709), .ZN(n7707) );
  NOR2_X1 U7755 ( .A1(n7425), .A2(n7427), .ZN(n7708) );
  NAND2_X1 U7756 ( .A1(n7425), .A2(n7427), .ZN(n7705) );
  NAND2_X1 U7757 ( .A1(n7710), .A2(n7711), .ZN(n7427) );
  NAND2_X1 U7758 ( .A1(n7712), .A2(b_31_), .ZN(n7711) );
  NOR2_X1 U7759 ( .A1(n7713), .A2(n7424), .ZN(n7712) );
  NOR2_X1 U7760 ( .A1(n7421), .A2(n7422), .ZN(n7713) );
  NAND2_X1 U7761 ( .A1(n7421), .A2(n7422), .ZN(n7710) );
  NAND2_X1 U7762 ( .A1(n7714), .A2(n7715), .ZN(n7422) );
  NAND2_X1 U7763 ( .A1(n7716), .A2(b_31_), .ZN(n7715) );
  NOR2_X1 U7764 ( .A1(n7717), .A2(n7718), .ZN(n7716) );
  NOR2_X1 U7765 ( .A1(n7416), .A2(n7418), .ZN(n7717) );
  NAND2_X1 U7766 ( .A1(n7416), .A2(n7418), .ZN(n7714) );
  NAND2_X1 U7767 ( .A1(n7719), .A2(n7720), .ZN(n7418) );
  NAND2_X1 U7768 ( .A1(n7721), .A2(b_31_), .ZN(n7720) );
  NOR2_X1 U7769 ( .A1(n7722), .A2(n7415), .ZN(n7721) );
  NOR2_X1 U7770 ( .A1(n7412), .A2(n7413), .ZN(n7722) );
  NAND2_X1 U7771 ( .A1(n7412), .A2(n7413), .ZN(n7719) );
  NAND2_X1 U7772 ( .A1(n7723), .A2(n7724), .ZN(n7413) );
  NAND2_X1 U7773 ( .A1(n7725), .A2(b_31_), .ZN(n7724) );
  NOR2_X1 U7774 ( .A1(n7726), .A2(n7727), .ZN(n7725) );
  NOR2_X1 U7775 ( .A1(n7407), .A2(n7409), .ZN(n7726) );
  NAND2_X1 U7776 ( .A1(n7407), .A2(n7409), .ZN(n7723) );
  NAND2_X1 U7777 ( .A1(n7728), .A2(n7729), .ZN(n7409) );
  NAND2_X1 U7778 ( .A1(n7730), .A2(b_31_), .ZN(n7729) );
  NOR2_X1 U7779 ( .A1(n7731), .A2(n7406), .ZN(n7730) );
  NOR2_X1 U7780 ( .A1(n7403), .A2(n7404), .ZN(n7731) );
  NAND2_X1 U7781 ( .A1(n7403), .A2(n7404), .ZN(n7728) );
  NAND2_X1 U7782 ( .A1(n7732), .A2(n7733), .ZN(n7404) );
  NAND2_X1 U7783 ( .A1(n7734), .A2(b_31_), .ZN(n7733) );
  NOR2_X1 U7784 ( .A1(n7735), .A2(n7736), .ZN(n7734) );
  NOR2_X1 U7785 ( .A1(n7398), .A2(n7400), .ZN(n7735) );
  NAND2_X1 U7786 ( .A1(n7398), .A2(n7400), .ZN(n7732) );
  NAND2_X1 U7787 ( .A1(n7737), .A2(n7738), .ZN(n7400) );
  NAND2_X1 U7788 ( .A1(n7739), .A2(b_31_), .ZN(n7738) );
  NOR2_X1 U7789 ( .A1(n7740), .A2(n7397), .ZN(n7739) );
  NOR2_X1 U7790 ( .A1(n7394), .A2(n7395), .ZN(n7740) );
  NAND2_X1 U7791 ( .A1(n7394), .A2(n7395), .ZN(n7737) );
  NAND2_X1 U7792 ( .A1(n7741), .A2(n7742), .ZN(n7395) );
  NAND2_X1 U7793 ( .A1(n7743), .A2(b_31_), .ZN(n7742) );
  NOR2_X1 U7794 ( .A1(n7744), .A2(n7745), .ZN(n7743) );
  NOR2_X1 U7795 ( .A1(n7385), .A2(n7387), .ZN(n7744) );
  NAND2_X1 U7796 ( .A1(n7385), .A2(n7387), .ZN(n7741) );
  NAND2_X1 U7797 ( .A1(n7746), .A2(n7747), .ZN(n7387) );
  NAND2_X1 U7798 ( .A1(n7748), .A2(b_31_), .ZN(n7747) );
  NOR2_X1 U7799 ( .A1(n7749), .A2(n7750), .ZN(n7748) );
  NOR2_X1 U7800 ( .A1(n7381), .A2(n7383), .ZN(n7749) );
  NAND2_X1 U7801 ( .A1(n7381), .A2(n7383), .ZN(n7746) );
  NAND2_X1 U7802 ( .A1(n7751), .A2(n7752), .ZN(n7383) );
  NAND2_X1 U7803 ( .A1(n7753), .A2(b_31_), .ZN(n7752) );
  NOR2_X1 U7804 ( .A1(n7754), .A2(n7755), .ZN(n7753) );
  NOR2_X1 U7805 ( .A1(n7377), .A2(n7379), .ZN(n7754) );
  NAND2_X1 U7806 ( .A1(n7377), .A2(n7379), .ZN(n7751) );
  NAND2_X1 U7807 ( .A1(n7756), .A2(n7757), .ZN(n7379) );
  NAND2_X1 U7808 ( .A1(n7758), .A2(b_31_), .ZN(n7757) );
  NOR2_X1 U7809 ( .A1(n7759), .A2(n7760), .ZN(n7758) );
  NOR2_X1 U7810 ( .A1(n7373), .A2(n7375), .ZN(n7759) );
  NAND2_X1 U7811 ( .A1(n7373), .A2(n7375), .ZN(n7756) );
  NAND2_X1 U7812 ( .A1(n7761), .A2(n7762), .ZN(n7375) );
  NAND2_X1 U7813 ( .A1(n7763), .A2(b_31_), .ZN(n7762) );
  NOR2_X1 U7814 ( .A1(n7764), .A2(n7765), .ZN(n7763) );
  NOR2_X1 U7815 ( .A1(n7369), .A2(n7371), .ZN(n7764) );
  NAND2_X1 U7816 ( .A1(n7369), .A2(n7371), .ZN(n7761) );
  NAND2_X1 U7817 ( .A1(n7367), .A2(n7766), .ZN(n7371) );
  NAND2_X1 U7818 ( .A1(n7366), .A2(n7368), .ZN(n7766) );
  NAND2_X1 U7819 ( .A1(n7767), .A2(n7768), .ZN(n7368) );
  NAND2_X1 U7820 ( .A1(b_31_), .A2(a_23_), .ZN(n7768) );
  INV_X1 U7821 ( .A(n7769), .ZN(n7767) );
  XOR2_X1 U7822 ( .A(n7770), .B(n7771), .Z(n7366) );
  XOR2_X1 U7823 ( .A(n7772), .B(n7773), .Z(n7770) );
  NOR2_X1 U7824 ( .A1(n7774), .A2(n7334), .ZN(n7773) );
  NAND2_X1 U7825 ( .A1(a_23_), .A2(n7769), .ZN(n7367) );
  NAND2_X1 U7826 ( .A1(n7775), .A2(n7776), .ZN(n7769) );
  NAND2_X1 U7827 ( .A1(n7777), .A2(b_31_), .ZN(n7776) );
  NOR2_X1 U7828 ( .A1(n7778), .A2(n7774), .ZN(n7777) );
  NOR2_X1 U7829 ( .A1(n7361), .A2(n7363), .ZN(n7778) );
  NAND2_X1 U7830 ( .A1(n7361), .A2(n7363), .ZN(n7775) );
  NAND2_X1 U7831 ( .A1(n7359), .A2(n7779), .ZN(n7363) );
  NAND2_X1 U7832 ( .A1(n7358), .A2(n7360), .ZN(n7779) );
  NAND2_X1 U7833 ( .A1(n7780), .A2(n7781), .ZN(n7360) );
  NAND2_X1 U7834 ( .A1(b_31_), .A2(a_25_), .ZN(n7781) );
  INV_X1 U7835 ( .A(n7782), .ZN(n7780) );
  XNOR2_X1 U7836 ( .A(n7783), .B(n7784), .ZN(n7358) );
  NAND2_X1 U7837 ( .A1(n7785), .A2(n7786), .ZN(n7783) );
  NAND2_X1 U7838 ( .A1(a_25_), .A2(n7782), .ZN(n7359) );
  NAND2_X1 U7839 ( .A1(n7787), .A2(n7788), .ZN(n7782) );
  NAND2_X1 U7840 ( .A1(n7789), .A2(b_31_), .ZN(n7788) );
  NOR2_X1 U7841 ( .A1(n7790), .A2(n7356), .ZN(n7789) );
  NOR2_X1 U7842 ( .A1(n7353), .A2(n7354), .ZN(n7790) );
  NAND2_X1 U7843 ( .A1(n7353), .A2(n7354), .ZN(n7787) );
  NAND2_X1 U7844 ( .A1(n7350), .A2(n7791), .ZN(n7354) );
  NAND2_X1 U7845 ( .A1(n7349), .A2(n7351), .ZN(n7791) );
  NAND2_X1 U7846 ( .A1(n7792), .A2(n7793), .ZN(n7351) );
  NAND2_X1 U7847 ( .A1(b_31_), .A2(a_27_), .ZN(n7793) );
  INV_X1 U7848 ( .A(n7794), .ZN(n7792) );
  XNOR2_X1 U7849 ( .A(n7795), .B(n7796), .ZN(n7349) );
  XOR2_X1 U7850 ( .A(n7797), .B(n7798), .Z(n7796) );
  NAND2_X1 U7851 ( .A1(b_30_), .A2(a_28_), .ZN(n7798) );
  NAND2_X1 U7852 ( .A1(a_27_), .A2(n7794), .ZN(n7350) );
  NAND2_X1 U7853 ( .A1(n7799), .A2(n7800), .ZN(n7794) );
  NAND2_X1 U7854 ( .A1(n7801), .A2(b_31_), .ZN(n7800) );
  NOR2_X1 U7855 ( .A1(n7802), .A2(n7803), .ZN(n7801) );
  NOR2_X1 U7856 ( .A1(n7340), .A2(n7343), .ZN(n7802) );
  NAND2_X1 U7857 ( .A1(n7340), .A2(n7343), .ZN(n7799) );
  NAND2_X1 U7858 ( .A1(n7804), .A2(n7805), .ZN(n7343) );
  NAND2_X1 U7859 ( .A1(n7806), .A2(b_31_), .ZN(n7805) );
  NOR2_X1 U7860 ( .A1(n7807), .A2(n7337), .ZN(n7806) );
  NOR2_X1 U7861 ( .A1(n7338), .A2(n7339), .ZN(n7807) );
  NAND2_X1 U7862 ( .A1(n7338), .A2(n7339), .ZN(n7804) );
  NAND2_X1 U7863 ( .A1(n7808), .A2(n7809), .ZN(n7339) );
  NAND2_X1 U7864 ( .A1(n7810), .A2(b_30_), .ZN(n7809) );
  NOR2_X1 U7865 ( .A1(n7811), .A2(n7812), .ZN(n7808) );
  NOR2_X1 U7866 ( .A1(n7813), .A2(n7814), .ZN(n7812) );
  NOR2_X1 U7867 ( .A1(n7815), .A2(n7816), .ZN(n7813) );
  NOR2_X1 U7868 ( .A1(b_30_), .A2(n7817), .ZN(n7815) );
  NOR2_X1 U7869 ( .A1(b_29_), .A2(n7818), .ZN(n7811) );
  XOR2_X1 U7870 ( .A(n7819), .B(n7820), .Z(n7340) );
  XOR2_X1 U7871 ( .A(n7821), .B(n7822), .Z(n7819) );
  XNOR2_X1 U7872 ( .A(n7823), .B(n7824), .ZN(n7353) );
  NAND2_X1 U7873 ( .A1(n7825), .A2(n7826), .ZN(n7823) );
  XOR2_X1 U7874 ( .A(n7827), .B(n7828), .Z(n7361) );
  XOR2_X1 U7875 ( .A(n7829), .B(n7830), .Z(n7827) );
  XOR2_X1 U7876 ( .A(n7831), .B(n7832), .Z(n7369) );
  XOR2_X1 U7877 ( .A(n7833), .B(n7834), .Z(n7831) );
  XOR2_X1 U7878 ( .A(n7835), .B(n7836), .Z(n7373) );
  XOR2_X1 U7879 ( .A(n7837), .B(n7838), .Z(n7835) );
  NOR2_X1 U7880 ( .A1(n7765), .A2(n7334), .ZN(n7838) );
  XOR2_X1 U7881 ( .A(n7839), .B(n7840), .Z(n7377) );
  XOR2_X1 U7882 ( .A(n7841), .B(n7842), .Z(n7839) );
  XOR2_X1 U7883 ( .A(n7843), .B(n7844), .Z(n7381) );
  XOR2_X1 U7884 ( .A(n7845), .B(n7846), .Z(n7843) );
  NOR2_X1 U7885 ( .A1(n7755), .A2(n7334), .ZN(n7846) );
  XOR2_X1 U7886 ( .A(n7847), .B(n7848), .Z(n7385) );
  XOR2_X1 U7887 ( .A(n7849), .B(n7850), .Z(n7847) );
  XNOR2_X1 U7888 ( .A(n7851), .B(n7852), .ZN(n7394) );
  XOR2_X1 U7889 ( .A(n7853), .B(n7854), .Z(n7852) );
  NAND2_X1 U7890 ( .A1(b_30_), .A2(a_18_), .ZN(n7854) );
  XOR2_X1 U7891 ( .A(n7855), .B(n7856), .Z(n7398) );
  XOR2_X1 U7892 ( .A(n7857), .B(n7858), .Z(n7855) );
  XOR2_X1 U7893 ( .A(n7859), .B(n7860), .Z(n7403) );
  XOR2_X1 U7894 ( .A(n7861), .B(n7862), .Z(n7859) );
  NOR2_X1 U7895 ( .A1(n7736), .A2(n7334), .ZN(n7862) );
  XOR2_X1 U7896 ( .A(n7863), .B(n7864), .Z(n7407) );
  XOR2_X1 U7897 ( .A(n7865), .B(n7866), .Z(n7863) );
  XOR2_X1 U7898 ( .A(n7867), .B(n7868), .Z(n7412) );
  XOR2_X1 U7899 ( .A(n7869), .B(n7870), .Z(n7867) );
  NOR2_X1 U7900 ( .A1(n7727), .A2(n7334), .ZN(n7870) );
  XOR2_X1 U7901 ( .A(n7871), .B(n7872), .Z(n7416) );
  XOR2_X1 U7902 ( .A(n7873), .B(n7874), .Z(n7871) );
  XOR2_X1 U7903 ( .A(n7875), .B(n7876), .Z(n7421) );
  XOR2_X1 U7904 ( .A(n7877), .B(n7878), .Z(n7875) );
  NOR2_X1 U7905 ( .A1(n7718), .A2(n7334), .ZN(n7878) );
  XOR2_X1 U7906 ( .A(n7879), .B(n7880), .Z(n7425) );
  XOR2_X1 U7907 ( .A(n7881), .B(n7882), .Z(n7879) );
  XNOR2_X1 U7908 ( .A(n7883), .B(n7884), .ZN(n7429) );
  XOR2_X1 U7909 ( .A(n7885), .B(n7886), .Z(n7884) );
  NAND2_X1 U7910 ( .A1(b_30_), .A2(a_10_), .ZN(n7886) );
  XOR2_X1 U7911 ( .A(n7887), .B(n7888), .Z(n7433) );
  XOR2_X1 U7912 ( .A(n7889), .B(n7890), .Z(n7887) );
  XOR2_X1 U7913 ( .A(n7891), .B(n7892), .Z(n7442) );
  XOR2_X1 U7914 ( .A(n7893), .B(n7894), .Z(n7891) );
  NOR2_X1 U7915 ( .A1(n7699), .A2(n7334), .ZN(n7894) );
  XNOR2_X1 U7916 ( .A(n7895), .B(n7896), .ZN(n7447) );
  XNOR2_X1 U7917 ( .A(n7897), .B(n7898), .ZN(n7895) );
  XOR2_X1 U7918 ( .A(n7899), .B(n7900), .Z(n7452) );
  XOR2_X1 U7919 ( .A(n7901), .B(n7902), .Z(n7899) );
  NOR2_X1 U7920 ( .A1(n7450), .A2(n7334), .ZN(n7902) );
  XOR2_X1 U7921 ( .A(n7903), .B(n7904), .Z(n7456) );
  XOR2_X1 U7922 ( .A(n7905), .B(n7906), .Z(n7903) );
  XNOR2_X1 U7923 ( .A(n7907), .B(n7908), .ZN(n7461) );
  XOR2_X1 U7924 ( .A(n7909), .B(n7910), .Z(n7908) );
  NAND2_X1 U7925 ( .A1(b_30_), .A2(a_4_), .ZN(n7910) );
  XNOR2_X1 U7926 ( .A(n7911), .B(n7912), .ZN(n7466) );
  XNOR2_X1 U7927 ( .A(n7913), .B(n7914), .ZN(n7911) );
  XNOR2_X1 U7928 ( .A(n7915), .B(n7916), .ZN(n7470) );
  XOR2_X1 U7929 ( .A(n7917), .B(n7918), .Z(n7916) );
  NAND2_X1 U7930 ( .A1(b_30_), .A2(a_2_), .ZN(n7918) );
  XOR2_X1 U7931 ( .A(n7919), .B(n7920), .Z(n7475) );
  XNOR2_X1 U7932 ( .A(n7921), .B(n7922), .ZN(n7919) );
  NAND2_X1 U7933 ( .A1(b_30_), .A2(a_1_), .ZN(n7921) );
  NAND2_X1 U7934 ( .A1(n7923), .A2(n7924), .ZN(n7491) );
  XOR2_X1 U7935 ( .A(n7650), .B(n7649), .Z(n7924) );
  AND2_X1 U7936 ( .A1(n7655), .A2(n7654), .ZN(n7923) );
  XOR2_X1 U7937 ( .A(n7925), .B(n7926), .Z(n7654) );
  XOR2_X1 U7938 ( .A(n7927), .B(n7928), .Z(n7925) );
  NOR2_X1 U7939 ( .A1(n7478), .A2(n7814), .ZN(n7928) );
  NAND2_X1 U7940 ( .A1(n7929), .A2(n7930), .ZN(n7655) );
  NAND2_X1 U7941 ( .A1(n7931), .A2(b_30_), .ZN(n7930) );
  NOR2_X1 U7942 ( .A1(n7932), .A2(n7478), .ZN(n7931) );
  NOR2_X1 U7943 ( .A1(n7658), .A2(n7659), .ZN(n7932) );
  NAND2_X1 U7944 ( .A1(n7658), .A2(n7659), .ZN(n7929) );
  NAND2_X1 U7945 ( .A1(n7933), .A2(n7934), .ZN(n7659) );
  NAND2_X1 U7946 ( .A1(n7935), .A2(b_30_), .ZN(n7934) );
  NOR2_X1 U7947 ( .A1(n7936), .A2(n7669), .ZN(n7935) );
  NOR2_X1 U7948 ( .A1(n7920), .A2(n7922), .ZN(n7936) );
  NAND2_X1 U7949 ( .A1(n7920), .A2(n7922), .ZN(n7933) );
  NAND2_X1 U7950 ( .A1(n7937), .A2(n7938), .ZN(n7922) );
  NAND2_X1 U7951 ( .A1(n7939), .A2(b_30_), .ZN(n7938) );
  NOR2_X1 U7952 ( .A1(n7940), .A2(n7469), .ZN(n7939) );
  NOR2_X1 U7953 ( .A1(n7917), .A2(n7915), .ZN(n7940) );
  NAND2_X1 U7954 ( .A1(n7915), .A2(n7917), .ZN(n7937) );
  NAND2_X1 U7955 ( .A1(n7941), .A2(n7942), .ZN(n7917) );
  NAND2_X1 U7956 ( .A1(n7914), .A2(n7943), .ZN(n7942) );
  NAND2_X1 U7957 ( .A1(n7913), .A2(n7912), .ZN(n7943) );
  NOR2_X1 U7958 ( .A1(n7334), .A2(n7464), .ZN(n7914) );
  OR2_X1 U7959 ( .A1(n7912), .A2(n7913), .ZN(n7941) );
  AND2_X1 U7960 ( .A1(n7944), .A2(n7945), .ZN(n7913) );
  NAND2_X1 U7961 ( .A1(n7946), .A2(b_30_), .ZN(n7945) );
  NOR2_X1 U7962 ( .A1(n7947), .A2(n7682), .ZN(n7946) );
  NOR2_X1 U7963 ( .A1(n7907), .A2(n7909), .ZN(n7947) );
  NAND2_X1 U7964 ( .A1(n7907), .A2(n7909), .ZN(n7944) );
  NAND2_X1 U7965 ( .A1(n7948), .A2(n7949), .ZN(n7909) );
  NAND2_X1 U7966 ( .A1(n7906), .A2(n7950), .ZN(n7949) );
  OR2_X1 U7967 ( .A1(n7904), .A2(n7905), .ZN(n7950) );
  NOR2_X1 U7968 ( .A1(n7334), .A2(n7455), .ZN(n7906) );
  NAND2_X1 U7969 ( .A1(n7904), .A2(n7905), .ZN(n7948) );
  NAND2_X1 U7970 ( .A1(n7951), .A2(n7952), .ZN(n7905) );
  NAND2_X1 U7971 ( .A1(n7953), .A2(b_30_), .ZN(n7952) );
  NOR2_X1 U7972 ( .A1(n7954), .A2(n7450), .ZN(n7953) );
  NOR2_X1 U7973 ( .A1(n7900), .A2(n7901), .ZN(n7954) );
  NAND2_X1 U7974 ( .A1(n7900), .A2(n7901), .ZN(n7951) );
  NAND2_X1 U7975 ( .A1(n7955), .A2(n7956), .ZN(n7901) );
  NAND2_X1 U7976 ( .A1(n7898), .A2(n7957), .ZN(n7956) );
  NAND2_X1 U7977 ( .A1(n7897), .A2(n7896), .ZN(n7957) );
  NOR2_X1 U7978 ( .A1(n7334), .A2(n7445), .ZN(n7898) );
  OR2_X1 U7979 ( .A1(n7896), .A2(n7897), .ZN(n7955) );
  AND2_X1 U7980 ( .A1(n7958), .A2(n7959), .ZN(n7897) );
  NAND2_X1 U7981 ( .A1(n7960), .A2(b_30_), .ZN(n7959) );
  NOR2_X1 U7982 ( .A1(n7961), .A2(n7699), .ZN(n7960) );
  NOR2_X1 U7983 ( .A1(n7892), .A2(n7893), .ZN(n7961) );
  NAND2_X1 U7984 ( .A1(n7892), .A2(n7893), .ZN(n7958) );
  NAND2_X1 U7985 ( .A1(n7962), .A2(n7963), .ZN(n7893) );
  NAND2_X1 U7986 ( .A1(n7890), .A2(n7964), .ZN(n7963) );
  OR2_X1 U7987 ( .A1(n7888), .A2(n7889), .ZN(n7964) );
  NOR2_X1 U7988 ( .A1(n7334), .A2(n7704), .ZN(n7890) );
  NAND2_X1 U7989 ( .A1(n7888), .A2(n7889), .ZN(n7962) );
  NAND2_X1 U7990 ( .A1(n7965), .A2(n7966), .ZN(n7889) );
  NAND2_X1 U7991 ( .A1(n7967), .A2(b_30_), .ZN(n7966) );
  NOR2_X1 U7992 ( .A1(n7968), .A2(n7709), .ZN(n7967) );
  NOR2_X1 U7993 ( .A1(n7885), .A2(n7883), .ZN(n7968) );
  NAND2_X1 U7994 ( .A1(n7883), .A2(n7885), .ZN(n7965) );
  NAND2_X1 U7995 ( .A1(n7969), .A2(n7970), .ZN(n7885) );
  NAND2_X1 U7996 ( .A1(n7882), .A2(n7971), .ZN(n7970) );
  OR2_X1 U7997 ( .A1(n7880), .A2(n7881), .ZN(n7971) );
  NOR2_X1 U7998 ( .A1(n7334), .A2(n7424), .ZN(n7882) );
  NAND2_X1 U7999 ( .A1(n7880), .A2(n7881), .ZN(n7969) );
  NAND2_X1 U8000 ( .A1(n7972), .A2(n7973), .ZN(n7881) );
  NAND2_X1 U8001 ( .A1(n7974), .A2(b_30_), .ZN(n7973) );
  NOR2_X1 U8002 ( .A1(n7975), .A2(n7718), .ZN(n7974) );
  NOR2_X1 U8003 ( .A1(n7876), .A2(n7877), .ZN(n7975) );
  NAND2_X1 U8004 ( .A1(n7876), .A2(n7877), .ZN(n7972) );
  NAND2_X1 U8005 ( .A1(n7976), .A2(n7977), .ZN(n7877) );
  NAND2_X1 U8006 ( .A1(n7874), .A2(n7978), .ZN(n7977) );
  OR2_X1 U8007 ( .A1(n7872), .A2(n7873), .ZN(n7978) );
  NOR2_X1 U8008 ( .A1(n7334), .A2(n7415), .ZN(n7874) );
  NAND2_X1 U8009 ( .A1(n7872), .A2(n7873), .ZN(n7976) );
  NAND2_X1 U8010 ( .A1(n7979), .A2(n7980), .ZN(n7873) );
  NAND2_X1 U8011 ( .A1(n7981), .A2(b_30_), .ZN(n7980) );
  NOR2_X1 U8012 ( .A1(n7982), .A2(n7727), .ZN(n7981) );
  NOR2_X1 U8013 ( .A1(n7868), .A2(n7869), .ZN(n7982) );
  NAND2_X1 U8014 ( .A1(n7868), .A2(n7869), .ZN(n7979) );
  NAND2_X1 U8015 ( .A1(n7983), .A2(n7984), .ZN(n7869) );
  NAND2_X1 U8016 ( .A1(n7866), .A2(n7985), .ZN(n7984) );
  OR2_X1 U8017 ( .A1(n7864), .A2(n7865), .ZN(n7985) );
  NOR2_X1 U8018 ( .A1(n7334), .A2(n7406), .ZN(n7866) );
  NAND2_X1 U8019 ( .A1(n7864), .A2(n7865), .ZN(n7983) );
  NAND2_X1 U8020 ( .A1(n7986), .A2(n7987), .ZN(n7865) );
  NAND2_X1 U8021 ( .A1(n7988), .A2(b_30_), .ZN(n7987) );
  NOR2_X1 U8022 ( .A1(n7989), .A2(n7736), .ZN(n7988) );
  NOR2_X1 U8023 ( .A1(n7860), .A2(n7861), .ZN(n7989) );
  NAND2_X1 U8024 ( .A1(n7860), .A2(n7861), .ZN(n7986) );
  NAND2_X1 U8025 ( .A1(n7990), .A2(n7991), .ZN(n7861) );
  NAND2_X1 U8026 ( .A1(n7858), .A2(n7992), .ZN(n7991) );
  OR2_X1 U8027 ( .A1(n7856), .A2(n7857), .ZN(n7992) );
  NOR2_X1 U8028 ( .A1(n7334), .A2(n7397), .ZN(n7858) );
  NAND2_X1 U8029 ( .A1(n7856), .A2(n7857), .ZN(n7990) );
  NAND2_X1 U8030 ( .A1(n7993), .A2(n7994), .ZN(n7857) );
  NAND2_X1 U8031 ( .A1(n7995), .A2(b_30_), .ZN(n7994) );
  NOR2_X1 U8032 ( .A1(n7996), .A2(n7745), .ZN(n7995) );
  NOR2_X1 U8033 ( .A1(n7851), .A2(n7853), .ZN(n7996) );
  NAND2_X1 U8034 ( .A1(n7851), .A2(n7853), .ZN(n7993) );
  NAND2_X1 U8035 ( .A1(n7997), .A2(n7998), .ZN(n7853) );
  NAND2_X1 U8036 ( .A1(n7850), .A2(n7999), .ZN(n7998) );
  OR2_X1 U8037 ( .A1(n7848), .A2(n7849), .ZN(n7999) );
  NOR2_X1 U8038 ( .A1(n7334), .A2(n7750), .ZN(n7850) );
  NAND2_X1 U8039 ( .A1(n7848), .A2(n7849), .ZN(n7997) );
  NAND2_X1 U8040 ( .A1(n8000), .A2(n8001), .ZN(n7849) );
  NAND2_X1 U8041 ( .A1(n8002), .A2(b_30_), .ZN(n8001) );
  NOR2_X1 U8042 ( .A1(n8003), .A2(n7755), .ZN(n8002) );
  NOR2_X1 U8043 ( .A1(n7844), .A2(n7845), .ZN(n8003) );
  NAND2_X1 U8044 ( .A1(n7844), .A2(n7845), .ZN(n8000) );
  NAND2_X1 U8045 ( .A1(n8004), .A2(n8005), .ZN(n7845) );
  NAND2_X1 U8046 ( .A1(n7841), .A2(n8006), .ZN(n8005) );
  OR2_X1 U8047 ( .A1(n7840), .A2(n7842), .ZN(n8006) );
  NOR2_X1 U8048 ( .A1(n7334), .A2(n7760), .ZN(n7841) );
  NAND2_X1 U8049 ( .A1(n7840), .A2(n7842), .ZN(n8004) );
  NAND2_X1 U8050 ( .A1(n8007), .A2(n8008), .ZN(n7842) );
  NAND2_X1 U8051 ( .A1(n8009), .A2(b_30_), .ZN(n8008) );
  NOR2_X1 U8052 ( .A1(n8010), .A2(n7765), .ZN(n8009) );
  NOR2_X1 U8053 ( .A1(n7837), .A2(n7836), .ZN(n8010) );
  NAND2_X1 U8054 ( .A1(n7836), .A2(n7837), .ZN(n8007) );
  NAND2_X1 U8055 ( .A1(n8011), .A2(n8012), .ZN(n7837) );
  NAND2_X1 U8056 ( .A1(n7833), .A2(n8013), .ZN(n8012) );
  OR2_X1 U8057 ( .A1(n7832), .A2(n7834), .ZN(n8013) );
  NOR2_X1 U8058 ( .A1(n7334), .A2(n8014), .ZN(n7833) );
  NAND2_X1 U8059 ( .A1(n7832), .A2(n7834), .ZN(n8011) );
  NAND2_X1 U8060 ( .A1(n8015), .A2(n8016), .ZN(n7834) );
  NAND2_X1 U8061 ( .A1(n8017), .A2(b_30_), .ZN(n8016) );
  NOR2_X1 U8062 ( .A1(n8018), .A2(n7774), .ZN(n8017) );
  NOR2_X1 U8063 ( .A1(n7772), .A2(n7771), .ZN(n8018) );
  NAND2_X1 U8064 ( .A1(n7771), .A2(n7772), .ZN(n8015) );
  NAND2_X1 U8065 ( .A1(n8019), .A2(n8020), .ZN(n7772) );
  NAND2_X1 U8066 ( .A1(n7830), .A2(n8021), .ZN(n8020) );
  OR2_X1 U8067 ( .A1(n7828), .A2(n7829), .ZN(n8021) );
  NOR2_X1 U8068 ( .A1(n7334), .A2(n8022), .ZN(n7830) );
  NAND2_X1 U8069 ( .A1(n7828), .A2(n7829), .ZN(n8019) );
  NAND2_X1 U8070 ( .A1(n7785), .A2(n8023), .ZN(n7829) );
  NAND2_X1 U8071 ( .A1(n7784), .A2(n7786), .ZN(n8023) );
  NAND2_X1 U8072 ( .A1(n8024), .A2(n8025), .ZN(n7786) );
  NAND2_X1 U8073 ( .A1(b_30_), .A2(a_26_), .ZN(n8025) );
  INV_X1 U8074 ( .A(n8026), .ZN(n8024) );
  XNOR2_X1 U8075 ( .A(n8027), .B(n8028), .ZN(n7784) );
  NAND2_X1 U8076 ( .A1(n8029), .A2(n8030), .ZN(n8027) );
  NAND2_X1 U8077 ( .A1(a_26_), .A2(n8026), .ZN(n7785) );
  NAND2_X1 U8078 ( .A1(n7825), .A2(n8031), .ZN(n8026) );
  NAND2_X1 U8079 ( .A1(n7824), .A2(n7826), .ZN(n8031) );
  NAND2_X1 U8080 ( .A1(n8032), .A2(n8033), .ZN(n7826) );
  NAND2_X1 U8081 ( .A1(b_30_), .A2(a_27_), .ZN(n8033) );
  INV_X1 U8082 ( .A(n8034), .ZN(n8032) );
  XNOR2_X1 U8083 ( .A(n8035), .B(n8036), .ZN(n7824) );
  XOR2_X1 U8084 ( .A(n8037), .B(n8038), .Z(n8036) );
  NAND2_X1 U8085 ( .A1(b_29_), .A2(a_28_), .ZN(n8038) );
  NAND2_X1 U8086 ( .A1(a_27_), .A2(n8034), .ZN(n7825) );
  NAND2_X1 U8087 ( .A1(n8039), .A2(n8040), .ZN(n8034) );
  NAND2_X1 U8088 ( .A1(n8041), .A2(b_30_), .ZN(n8040) );
  NOR2_X1 U8089 ( .A1(n8042), .A2(n7803), .ZN(n8041) );
  NOR2_X1 U8090 ( .A1(n7795), .A2(n7797), .ZN(n8042) );
  NAND2_X1 U8091 ( .A1(n7795), .A2(n7797), .ZN(n8039) );
  NAND2_X1 U8092 ( .A1(n8043), .A2(n8044), .ZN(n7797) );
  NAND2_X1 U8093 ( .A1(n7820), .A2(n8045), .ZN(n8044) );
  NAND2_X1 U8094 ( .A1(n7822), .A2(n7821), .ZN(n8045) );
  NOR2_X1 U8095 ( .A1(n7334), .A2(n7337), .ZN(n7820) );
  OR2_X1 U8096 ( .A1(n7821), .A2(n7822), .ZN(n8043) );
  AND2_X1 U8097 ( .A1(n8046), .A2(n8047), .ZN(n7822) );
  NAND2_X1 U8098 ( .A1(n8048), .A2(b_28_), .ZN(n8047) );
  NOR2_X1 U8099 ( .A1(n8049), .A2(n7817), .ZN(n8048) );
  NOR2_X1 U8100 ( .A1(n7816), .A2(n7814), .ZN(n8049) );
  NAND2_X1 U8101 ( .A1(n8050), .A2(b_29_), .ZN(n8046) );
  NOR2_X1 U8102 ( .A1(n8051), .A2(n8052), .ZN(n8050) );
  NOR2_X1 U8103 ( .A1(n7810), .A2(n8053), .ZN(n8051) );
  NAND2_X1 U8104 ( .A1(n8054), .A2(b_30_), .ZN(n7821) );
  NOR2_X1 U8105 ( .A1(n8055), .A2(n7814), .ZN(n8054) );
  XOR2_X1 U8106 ( .A(n8056), .B(n8057), .Z(n7795) );
  XOR2_X1 U8107 ( .A(n8058), .B(n8059), .Z(n8056) );
  XNOR2_X1 U8108 ( .A(n8060), .B(n8061), .ZN(n7828) );
  NAND2_X1 U8109 ( .A1(n8062), .A2(n8063), .ZN(n8060) );
  XNOR2_X1 U8110 ( .A(n8064), .B(n8065), .ZN(n7771) );
  XNOR2_X1 U8111 ( .A(n8066), .B(n8067), .ZN(n8064) );
  XNOR2_X1 U8112 ( .A(n8068), .B(n8069), .ZN(n7832) );
  XOR2_X1 U8113 ( .A(n8070), .B(n8071), .Z(n8069) );
  NAND2_X1 U8114 ( .A1(b_29_), .A2(a_24_), .ZN(n8071) );
  XNOR2_X1 U8115 ( .A(n8072), .B(n8073), .ZN(n7836) );
  XNOR2_X1 U8116 ( .A(n8074), .B(n8075), .ZN(n8072) );
  XNOR2_X1 U8117 ( .A(n8076), .B(n8077), .ZN(n7840) );
  XOR2_X1 U8118 ( .A(n8078), .B(n8079), .Z(n8077) );
  NAND2_X1 U8119 ( .A1(b_29_), .A2(a_22_), .ZN(n8079) );
  XOR2_X1 U8120 ( .A(n8080), .B(n8081), .Z(n7844) );
  XOR2_X1 U8121 ( .A(n8082), .B(n8083), .Z(n8080) );
  XNOR2_X1 U8122 ( .A(n8084), .B(n8085), .ZN(n7848) );
  XOR2_X1 U8123 ( .A(n8086), .B(n8087), .Z(n8085) );
  NAND2_X1 U8124 ( .A1(b_29_), .A2(a_20_), .ZN(n8087) );
  XOR2_X1 U8125 ( .A(n8088), .B(n8089), .Z(n7851) );
  XOR2_X1 U8126 ( .A(n8090), .B(n8091), .Z(n8088) );
  XOR2_X1 U8127 ( .A(n8092), .B(n8093), .Z(n7856) );
  XOR2_X1 U8128 ( .A(n8094), .B(n8095), .Z(n8092) );
  NOR2_X1 U8129 ( .A1(n7745), .A2(n7814), .ZN(n8095) );
  XNOR2_X1 U8130 ( .A(n8096), .B(n8097), .ZN(n7860) );
  XNOR2_X1 U8131 ( .A(n8098), .B(n8099), .ZN(n8097) );
  XOR2_X1 U8132 ( .A(n8100), .B(n8101), .Z(n7864) );
  XOR2_X1 U8133 ( .A(n8102), .B(n8103), .Z(n8100) );
  NOR2_X1 U8134 ( .A1(n7736), .A2(n7814), .ZN(n8103) );
  XOR2_X1 U8135 ( .A(n8104), .B(n8105), .Z(n7868) );
  XOR2_X1 U8136 ( .A(n8106), .B(n8107), .Z(n8104) );
  XOR2_X1 U8137 ( .A(n8108), .B(n8109), .Z(n7872) );
  XOR2_X1 U8138 ( .A(n8110), .B(n8111), .Z(n8108) );
  NOR2_X1 U8139 ( .A1(n7727), .A2(n7814), .ZN(n8111) );
  XOR2_X1 U8140 ( .A(n8112), .B(n8113), .Z(n7876) );
  XOR2_X1 U8141 ( .A(n8114), .B(n8115), .Z(n8112) );
  XNOR2_X1 U8142 ( .A(n8116), .B(n8117), .ZN(n7880) );
  XOR2_X1 U8143 ( .A(n8118), .B(n8119), .Z(n8117) );
  NAND2_X1 U8144 ( .A1(b_29_), .A2(a_12_), .ZN(n8119) );
  XNOR2_X1 U8145 ( .A(n8120), .B(n8121), .ZN(n7883) );
  XNOR2_X1 U8146 ( .A(n8122), .B(n8123), .ZN(n8120) );
  XOR2_X1 U8147 ( .A(n8124), .B(n8125), .Z(n7888) );
  XOR2_X1 U8148 ( .A(n8126), .B(n8127), .Z(n8124) );
  NOR2_X1 U8149 ( .A1(n7709), .A2(n7814), .ZN(n8127) );
  XOR2_X1 U8150 ( .A(n8128), .B(n8129), .Z(n7892) );
  XOR2_X1 U8151 ( .A(n8130), .B(n8131), .Z(n8128) );
  XNOR2_X1 U8152 ( .A(n8132), .B(n8133), .ZN(n7896) );
  XOR2_X1 U8153 ( .A(n8134), .B(n8135), .Z(n8132) );
  NOR2_X1 U8154 ( .A1(n7699), .A2(n7814), .ZN(n8135) );
  XOR2_X1 U8155 ( .A(n8136), .B(n8137), .Z(n7900) );
  XOR2_X1 U8156 ( .A(n8138), .B(n8139), .Z(n8136) );
  XNOR2_X1 U8157 ( .A(n8140), .B(n8141), .ZN(n7904) );
  XOR2_X1 U8158 ( .A(n8142), .B(n8143), .Z(n8141) );
  NAND2_X1 U8159 ( .A1(b_29_), .A2(a_6_), .ZN(n8143) );
  XOR2_X1 U8160 ( .A(n8144), .B(n8145), .Z(n7907) );
  XOR2_X1 U8161 ( .A(n8146), .B(n8147), .Z(n8144) );
  XNOR2_X1 U8162 ( .A(n8148), .B(n8149), .ZN(n7912) );
  XOR2_X1 U8163 ( .A(n8150), .B(n8151), .Z(n8148) );
  NOR2_X1 U8164 ( .A1(n7682), .A2(n7814), .ZN(n8151) );
  XNOR2_X1 U8165 ( .A(n8152), .B(n8153), .ZN(n7915) );
  XOR2_X1 U8166 ( .A(n8154), .B(n8155), .Z(n8153) );
  NAND2_X1 U8167 ( .A1(b_29_), .A2(a_3_), .ZN(n8155) );
  XOR2_X1 U8168 ( .A(n8156), .B(n8157), .Z(n7920) );
  XOR2_X1 U8169 ( .A(n8158), .B(n8159), .Z(n8156) );
  XOR2_X1 U8170 ( .A(n8160), .B(n8161), .Z(n7658) );
  XOR2_X1 U8171 ( .A(n8162), .B(n8163), .Z(n8160) );
  NOR2_X1 U8172 ( .A1(n7669), .A2(n7814), .ZN(n8163) );
  NAND2_X1 U8173 ( .A1(n8164), .A2(n7649), .ZN(n7494) );
  XOR2_X1 U8174 ( .A(n8165), .B(n8166), .Z(n7649) );
  XOR2_X1 U8175 ( .A(n8167), .B(n8168), .Z(n8165) );
  NOR2_X1 U8176 ( .A1(n7656), .A2(n7647), .ZN(n8164) );
  XNOR2_X1 U8177 ( .A(n8169), .B(n8170), .ZN(n7647) );
  INV_X1 U8178 ( .A(n7650), .ZN(n7656) );
  NAND2_X1 U8179 ( .A1(n8171), .A2(n8172), .ZN(n7650) );
  NAND2_X1 U8180 ( .A1(n8173), .A2(b_29_), .ZN(n8172) );
  NOR2_X1 U8181 ( .A1(n8174), .A2(n7478), .ZN(n8173) );
  NOR2_X1 U8182 ( .A1(n7926), .A2(n7927), .ZN(n8174) );
  NAND2_X1 U8183 ( .A1(n7926), .A2(n7927), .ZN(n8171) );
  NAND2_X1 U8184 ( .A1(n8175), .A2(n8176), .ZN(n7927) );
  NAND2_X1 U8185 ( .A1(n8177), .A2(b_29_), .ZN(n8176) );
  NOR2_X1 U8186 ( .A1(n8178), .A2(n7669), .ZN(n8177) );
  NOR2_X1 U8187 ( .A1(n8161), .A2(n8162), .ZN(n8178) );
  NAND2_X1 U8188 ( .A1(n8161), .A2(n8162), .ZN(n8175) );
  NAND2_X1 U8189 ( .A1(n8179), .A2(n8180), .ZN(n8162) );
  NAND2_X1 U8190 ( .A1(n8158), .A2(n8181), .ZN(n8180) );
  OR2_X1 U8191 ( .A1(n8157), .A2(n8159), .ZN(n8181) );
  NAND2_X1 U8192 ( .A1(n8182), .A2(n8183), .ZN(n8158) );
  NAND2_X1 U8193 ( .A1(n8184), .A2(b_29_), .ZN(n8183) );
  NOR2_X1 U8194 ( .A1(n8185), .A2(n7464), .ZN(n8184) );
  NOR2_X1 U8195 ( .A1(n8152), .A2(n8154), .ZN(n8185) );
  NAND2_X1 U8196 ( .A1(n8152), .A2(n8154), .ZN(n8182) );
  NAND2_X1 U8197 ( .A1(n8186), .A2(n8187), .ZN(n8154) );
  NAND2_X1 U8198 ( .A1(n8188), .A2(b_29_), .ZN(n8187) );
  NOR2_X1 U8199 ( .A1(n8189), .A2(n7682), .ZN(n8188) );
  NOR2_X1 U8200 ( .A1(n8149), .A2(n8150), .ZN(n8189) );
  NAND2_X1 U8201 ( .A1(n8149), .A2(n8150), .ZN(n8186) );
  NAND2_X1 U8202 ( .A1(n8190), .A2(n8191), .ZN(n8150) );
  NAND2_X1 U8203 ( .A1(n8147), .A2(n8192), .ZN(n8191) );
  OR2_X1 U8204 ( .A1(n8146), .A2(n8145), .ZN(n8192) );
  NOR2_X1 U8205 ( .A1(n7814), .A2(n7455), .ZN(n8147) );
  NAND2_X1 U8206 ( .A1(n8145), .A2(n8146), .ZN(n8190) );
  NAND2_X1 U8207 ( .A1(n8193), .A2(n8194), .ZN(n8146) );
  NAND2_X1 U8208 ( .A1(n8195), .A2(b_29_), .ZN(n8194) );
  NOR2_X1 U8209 ( .A1(n8196), .A2(n7450), .ZN(n8195) );
  NOR2_X1 U8210 ( .A1(n8140), .A2(n8142), .ZN(n8196) );
  NAND2_X1 U8211 ( .A1(n8140), .A2(n8142), .ZN(n8193) );
  NAND2_X1 U8212 ( .A1(n8197), .A2(n8198), .ZN(n8142) );
  NAND2_X1 U8213 ( .A1(n8138), .A2(n8199), .ZN(n8198) );
  OR2_X1 U8214 ( .A1(n8139), .A2(n8137), .ZN(n8199) );
  NOR2_X1 U8215 ( .A1(n7814), .A2(n7445), .ZN(n8138) );
  NAND2_X1 U8216 ( .A1(n8137), .A2(n8139), .ZN(n8197) );
  NAND2_X1 U8217 ( .A1(n8200), .A2(n8201), .ZN(n8139) );
  NAND2_X1 U8218 ( .A1(n8202), .A2(b_29_), .ZN(n8201) );
  NOR2_X1 U8219 ( .A1(n8203), .A2(n7699), .ZN(n8202) );
  NOR2_X1 U8220 ( .A1(n8133), .A2(n8134), .ZN(n8203) );
  NAND2_X1 U8221 ( .A1(n8133), .A2(n8134), .ZN(n8200) );
  NAND2_X1 U8222 ( .A1(n8204), .A2(n8205), .ZN(n8134) );
  NAND2_X1 U8223 ( .A1(n8131), .A2(n8206), .ZN(n8205) );
  OR2_X1 U8224 ( .A1(n8130), .A2(n8129), .ZN(n8206) );
  NOR2_X1 U8225 ( .A1(n7814), .A2(n7704), .ZN(n8131) );
  NAND2_X1 U8226 ( .A1(n8129), .A2(n8130), .ZN(n8204) );
  NAND2_X1 U8227 ( .A1(n8207), .A2(n8208), .ZN(n8130) );
  NAND2_X1 U8228 ( .A1(n8209), .A2(b_29_), .ZN(n8208) );
  NOR2_X1 U8229 ( .A1(n8210), .A2(n7709), .ZN(n8209) );
  NOR2_X1 U8230 ( .A1(n8125), .A2(n8126), .ZN(n8210) );
  NAND2_X1 U8231 ( .A1(n8125), .A2(n8126), .ZN(n8207) );
  NAND2_X1 U8232 ( .A1(n8211), .A2(n8212), .ZN(n8126) );
  NAND2_X1 U8233 ( .A1(n8123), .A2(n8213), .ZN(n8212) );
  NAND2_X1 U8234 ( .A1(n8122), .A2(n8121), .ZN(n8213) );
  NOR2_X1 U8235 ( .A1(n7814), .A2(n7424), .ZN(n8123) );
  OR2_X1 U8236 ( .A1(n8121), .A2(n8122), .ZN(n8211) );
  AND2_X1 U8237 ( .A1(n8214), .A2(n8215), .ZN(n8122) );
  NAND2_X1 U8238 ( .A1(n8216), .A2(b_29_), .ZN(n8215) );
  NOR2_X1 U8239 ( .A1(n8217), .A2(n7718), .ZN(n8216) );
  NOR2_X1 U8240 ( .A1(n8116), .A2(n8118), .ZN(n8217) );
  NAND2_X1 U8241 ( .A1(n8116), .A2(n8118), .ZN(n8214) );
  NAND2_X1 U8242 ( .A1(n8218), .A2(n8219), .ZN(n8118) );
  NAND2_X1 U8243 ( .A1(n8115), .A2(n8220), .ZN(n8219) );
  OR2_X1 U8244 ( .A1(n8114), .A2(n8113), .ZN(n8220) );
  NOR2_X1 U8245 ( .A1(n7814), .A2(n7415), .ZN(n8115) );
  NAND2_X1 U8246 ( .A1(n8113), .A2(n8114), .ZN(n8218) );
  NAND2_X1 U8247 ( .A1(n8221), .A2(n8222), .ZN(n8114) );
  NAND2_X1 U8248 ( .A1(n8223), .A2(b_29_), .ZN(n8222) );
  NOR2_X1 U8249 ( .A1(n8224), .A2(n7727), .ZN(n8223) );
  NOR2_X1 U8250 ( .A1(n8109), .A2(n8110), .ZN(n8224) );
  NAND2_X1 U8251 ( .A1(n8109), .A2(n8110), .ZN(n8221) );
  NAND2_X1 U8252 ( .A1(n8225), .A2(n8226), .ZN(n8110) );
  NAND2_X1 U8253 ( .A1(n8107), .A2(n8227), .ZN(n8226) );
  OR2_X1 U8254 ( .A1(n8106), .A2(n8105), .ZN(n8227) );
  NOR2_X1 U8255 ( .A1(n7814), .A2(n7406), .ZN(n8107) );
  NAND2_X1 U8256 ( .A1(n8105), .A2(n8106), .ZN(n8225) );
  NAND2_X1 U8257 ( .A1(n8228), .A2(n8229), .ZN(n8106) );
  NAND2_X1 U8258 ( .A1(n8230), .A2(b_29_), .ZN(n8229) );
  NOR2_X1 U8259 ( .A1(n8231), .A2(n7736), .ZN(n8230) );
  NOR2_X1 U8260 ( .A1(n8101), .A2(n8102), .ZN(n8231) );
  NAND2_X1 U8261 ( .A1(n8101), .A2(n8102), .ZN(n8228) );
  NAND2_X1 U8262 ( .A1(n8232), .A2(n8233), .ZN(n8102) );
  NAND2_X1 U8263 ( .A1(n8099), .A2(n8234), .ZN(n8233) );
  OR2_X1 U8264 ( .A1(n8098), .A2(n8096), .ZN(n8234) );
  NOR2_X1 U8265 ( .A1(n7814), .A2(n7397), .ZN(n8099) );
  NAND2_X1 U8266 ( .A1(n8096), .A2(n8098), .ZN(n8232) );
  NAND2_X1 U8267 ( .A1(n8235), .A2(n8236), .ZN(n8098) );
  NAND2_X1 U8268 ( .A1(n8237), .A2(b_29_), .ZN(n8236) );
  NOR2_X1 U8269 ( .A1(n8238), .A2(n7745), .ZN(n8237) );
  NOR2_X1 U8270 ( .A1(n8093), .A2(n8094), .ZN(n8238) );
  NAND2_X1 U8271 ( .A1(n8093), .A2(n8094), .ZN(n8235) );
  NAND2_X1 U8272 ( .A1(n8239), .A2(n8240), .ZN(n8094) );
  NAND2_X1 U8273 ( .A1(n8091), .A2(n8241), .ZN(n8240) );
  OR2_X1 U8274 ( .A1(n8090), .A2(n8089), .ZN(n8241) );
  NOR2_X1 U8275 ( .A1(n7814), .A2(n7750), .ZN(n8091) );
  NAND2_X1 U8276 ( .A1(n8089), .A2(n8090), .ZN(n8239) );
  NAND2_X1 U8277 ( .A1(n8242), .A2(n8243), .ZN(n8090) );
  NAND2_X1 U8278 ( .A1(n8244), .A2(b_29_), .ZN(n8243) );
  NOR2_X1 U8279 ( .A1(n8245), .A2(n7755), .ZN(n8244) );
  NOR2_X1 U8280 ( .A1(n8084), .A2(n8086), .ZN(n8245) );
  NAND2_X1 U8281 ( .A1(n8084), .A2(n8086), .ZN(n8242) );
  NAND2_X1 U8282 ( .A1(n8246), .A2(n8247), .ZN(n8086) );
  NAND2_X1 U8283 ( .A1(n8083), .A2(n8248), .ZN(n8247) );
  OR2_X1 U8284 ( .A1(n8082), .A2(n8081), .ZN(n8248) );
  NOR2_X1 U8285 ( .A1(n7814), .A2(n7760), .ZN(n8083) );
  NAND2_X1 U8286 ( .A1(n8081), .A2(n8082), .ZN(n8246) );
  NAND2_X1 U8287 ( .A1(n8249), .A2(n8250), .ZN(n8082) );
  NAND2_X1 U8288 ( .A1(n8251), .A2(b_29_), .ZN(n8250) );
  NOR2_X1 U8289 ( .A1(n8252), .A2(n7765), .ZN(n8251) );
  NOR2_X1 U8290 ( .A1(n8076), .A2(n8078), .ZN(n8252) );
  NAND2_X1 U8291 ( .A1(n8076), .A2(n8078), .ZN(n8249) );
  NAND2_X1 U8292 ( .A1(n8253), .A2(n8254), .ZN(n8078) );
  NAND2_X1 U8293 ( .A1(n8075), .A2(n8255), .ZN(n8254) );
  NAND2_X1 U8294 ( .A1(n8074), .A2(n8073), .ZN(n8255) );
  NOR2_X1 U8295 ( .A1(n7814), .A2(n8014), .ZN(n8075) );
  OR2_X1 U8296 ( .A1(n8073), .A2(n8074), .ZN(n8253) );
  AND2_X1 U8297 ( .A1(n8256), .A2(n8257), .ZN(n8074) );
  NAND2_X1 U8298 ( .A1(n8258), .A2(b_29_), .ZN(n8257) );
  NOR2_X1 U8299 ( .A1(n8259), .A2(n7774), .ZN(n8258) );
  NOR2_X1 U8300 ( .A1(n8068), .A2(n8070), .ZN(n8259) );
  NAND2_X1 U8301 ( .A1(n8068), .A2(n8070), .ZN(n8256) );
  NAND2_X1 U8302 ( .A1(n8260), .A2(n8261), .ZN(n8070) );
  NAND2_X1 U8303 ( .A1(n8067), .A2(n8262), .ZN(n8261) );
  NAND2_X1 U8304 ( .A1(n8066), .A2(n8065), .ZN(n8262) );
  NOR2_X1 U8305 ( .A1(n7814), .A2(n8022), .ZN(n8067) );
  OR2_X1 U8306 ( .A1(n8065), .A2(n8066), .ZN(n8260) );
  AND2_X1 U8307 ( .A1(n8062), .A2(n8263), .ZN(n8066) );
  NAND2_X1 U8308 ( .A1(n8061), .A2(n8063), .ZN(n8263) );
  NAND2_X1 U8309 ( .A1(n8264), .A2(n8265), .ZN(n8063) );
  NAND2_X1 U8310 ( .A1(b_29_), .A2(a_26_), .ZN(n8265) );
  INV_X1 U8311 ( .A(n8266), .ZN(n8264) );
  XNOR2_X1 U8312 ( .A(n8267), .B(n8268), .ZN(n8061) );
  NAND2_X1 U8313 ( .A1(n8269), .A2(n8270), .ZN(n8267) );
  NAND2_X1 U8314 ( .A1(a_26_), .A2(n8266), .ZN(n8062) );
  NAND2_X1 U8315 ( .A1(n8029), .A2(n8271), .ZN(n8266) );
  NAND2_X1 U8316 ( .A1(n8028), .A2(n8030), .ZN(n8271) );
  NAND2_X1 U8317 ( .A1(n8272), .A2(n8273), .ZN(n8030) );
  NAND2_X1 U8318 ( .A1(b_29_), .A2(a_27_), .ZN(n8273) );
  INV_X1 U8319 ( .A(n8274), .ZN(n8272) );
  XNOR2_X1 U8320 ( .A(n8275), .B(n8276), .ZN(n8028) );
  XOR2_X1 U8321 ( .A(n8277), .B(n8278), .Z(n8276) );
  NAND2_X1 U8322 ( .A1(a_27_), .A2(n8274), .ZN(n8029) );
  NAND2_X1 U8323 ( .A1(n8279), .A2(n8280), .ZN(n8274) );
  NAND2_X1 U8324 ( .A1(n8281), .A2(b_29_), .ZN(n8280) );
  NOR2_X1 U8325 ( .A1(n8282), .A2(n7803), .ZN(n8281) );
  NOR2_X1 U8326 ( .A1(n8035), .A2(n8037), .ZN(n8282) );
  NAND2_X1 U8327 ( .A1(n8035), .A2(n8037), .ZN(n8279) );
  NAND2_X1 U8328 ( .A1(n8283), .A2(n8284), .ZN(n8037) );
  NAND2_X1 U8329 ( .A1(n8057), .A2(n8285), .ZN(n8284) );
  NAND2_X1 U8330 ( .A1(n8059), .A2(n8058), .ZN(n8285) );
  OR2_X1 U8331 ( .A1(n8058), .A2(n8059), .ZN(n8283) );
  AND2_X1 U8332 ( .A1(n8286), .A2(n8287), .ZN(n8059) );
  NAND2_X1 U8333 ( .A1(n8288), .A2(b_27_), .ZN(n8287) );
  NOR2_X1 U8334 ( .A1(n8289), .A2(n7817), .ZN(n8288) );
  NOR2_X1 U8335 ( .A1(n7816), .A2(n8053), .ZN(n8289) );
  NAND2_X1 U8336 ( .A1(n8290), .A2(b_28_), .ZN(n8286) );
  NOR2_X1 U8337 ( .A1(n8291), .A2(n8052), .ZN(n8290) );
  NOR2_X1 U8338 ( .A1(n7810), .A2(n8292), .ZN(n8291) );
  NAND2_X1 U8339 ( .A1(n8293), .A2(b_29_), .ZN(n8058) );
  NOR2_X1 U8340 ( .A1(n8055), .A2(n8053), .ZN(n8293) );
  XOR2_X1 U8341 ( .A(n8294), .B(n8295), .Z(n8035) );
  XOR2_X1 U8342 ( .A(n8296), .B(n8297), .Z(n8294) );
  XOR2_X1 U8343 ( .A(n8298), .B(n8299), .Z(n8065) );
  NAND2_X1 U8344 ( .A1(n8300), .A2(n8301), .ZN(n8298) );
  XOR2_X1 U8345 ( .A(n8302), .B(n8303), .Z(n8068) );
  XOR2_X1 U8346 ( .A(n8304), .B(n8305), .Z(n8302) );
  XNOR2_X1 U8347 ( .A(n8306), .B(n8307), .ZN(n8073) );
  XNOR2_X1 U8348 ( .A(n8308), .B(n8309), .ZN(n8306) );
  NAND2_X1 U8349 ( .A1(b_28_), .A2(a_24_), .ZN(n8308) );
  XOR2_X1 U8350 ( .A(n8310), .B(n8311), .Z(n8076) );
  XOR2_X1 U8351 ( .A(n8312), .B(n8313), .Z(n8310) );
  XNOR2_X1 U8352 ( .A(n8314), .B(n8315), .ZN(n8081) );
  XOR2_X1 U8353 ( .A(n8316), .B(n8317), .Z(n8315) );
  NAND2_X1 U8354 ( .A1(b_28_), .A2(a_22_), .ZN(n8317) );
  XOR2_X1 U8355 ( .A(n8318), .B(n8319), .Z(n8084) );
  XOR2_X1 U8356 ( .A(n8320), .B(n8321), .Z(n8318) );
  XOR2_X1 U8357 ( .A(n8322), .B(n8323), .Z(n8089) );
  XOR2_X1 U8358 ( .A(n8324), .B(n8325), .Z(n8322) );
  NOR2_X1 U8359 ( .A1(n7755), .A2(n8053), .ZN(n8325) );
  XOR2_X1 U8360 ( .A(n8326), .B(n8327), .Z(n8093) );
  XOR2_X1 U8361 ( .A(n8328), .B(n8329), .Z(n8326) );
  XOR2_X1 U8362 ( .A(n8330), .B(n8331), .Z(n8096) );
  XOR2_X1 U8363 ( .A(n8332), .B(n8333), .Z(n8330) );
  NOR2_X1 U8364 ( .A1(n7745), .A2(n8053), .ZN(n8333) );
  XOR2_X1 U8365 ( .A(n8334), .B(n8335), .Z(n8101) );
  XOR2_X1 U8366 ( .A(n8336), .B(n8337), .Z(n8334) );
  XOR2_X1 U8367 ( .A(n8338), .B(n8339), .Z(n8105) );
  XOR2_X1 U8368 ( .A(n8340), .B(n8341), .Z(n8338) );
  NOR2_X1 U8369 ( .A1(n7736), .A2(n8053), .ZN(n8341) );
  XOR2_X1 U8370 ( .A(n8342), .B(n8343), .Z(n8109) );
  XOR2_X1 U8371 ( .A(n8344), .B(n8345), .Z(n8342) );
  XNOR2_X1 U8372 ( .A(n8346), .B(n8347), .ZN(n8113) );
  XOR2_X1 U8373 ( .A(n8348), .B(n8349), .Z(n8347) );
  NAND2_X1 U8374 ( .A1(b_28_), .A2(a_14_), .ZN(n8349) );
  XOR2_X1 U8375 ( .A(n8350), .B(n8351), .Z(n8116) );
  XOR2_X1 U8376 ( .A(n8352), .B(n8353), .Z(n8350) );
  XNOR2_X1 U8377 ( .A(n8354), .B(n8355), .ZN(n8121) );
  XOR2_X1 U8378 ( .A(n8356), .B(n8357), .Z(n8354) );
  NOR2_X1 U8379 ( .A1(n7718), .A2(n8053), .ZN(n8357) );
  XOR2_X1 U8380 ( .A(n8358), .B(n8359), .Z(n8125) );
  XOR2_X1 U8381 ( .A(n8360), .B(n8361), .Z(n8358) );
  XOR2_X1 U8382 ( .A(n8362), .B(n8363), .Z(n8129) );
  XOR2_X1 U8383 ( .A(n8364), .B(n8365), .Z(n8362) );
  NOR2_X1 U8384 ( .A1(n7709), .A2(n8053), .ZN(n8365) );
  XNOR2_X1 U8385 ( .A(n8366), .B(n8367), .ZN(n8133) );
  XNOR2_X1 U8386 ( .A(n8368), .B(n8369), .ZN(n8366) );
  XNOR2_X1 U8387 ( .A(n8370), .B(n8371), .ZN(n8137) );
  XOR2_X1 U8388 ( .A(n8372), .B(n8373), .Z(n8371) );
  NAND2_X1 U8389 ( .A1(b_28_), .A2(a_8_), .ZN(n8373) );
  XOR2_X1 U8390 ( .A(n8374), .B(n8375), .Z(n8140) );
  XOR2_X1 U8391 ( .A(n8376), .B(n8377), .Z(n8374) );
  XNOR2_X1 U8392 ( .A(n8378), .B(n8379), .ZN(n8145) );
  XOR2_X1 U8393 ( .A(n8380), .B(n8381), .Z(n8379) );
  NAND2_X1 U8394 ( .A1(b_28_), .A2(a_6_), .ZN(n8381) );
  XNOR2_X1 U8395 ( .A(n8382), .B(n8383), .ZN(n8149) );
  XNOR2_X1 U8396 ( .A(n8384), .B(n8385), .ZN(n8382) );
  XNOR2_X1 U8397 ( .A(n8386), .B(n8387), .ZN(n8152) );
  XOR2_X1 U8398 ( .A(n8388), .B(n8389), .Z(n8387) );
  NAND2_X1 U8399 ( .A1(b_28_), .A2(a_4_), .ZN(n8389) );
  NAND2_X1 U8400 ( .A1(n8159), .A2(n8157), .ZN(n8179) );
  XNOR2_X1 U8401 ( .A(n8390), .B(n8391), .ZN(n8157) );
  NAND2_X1 U8402 ( .A1(n8392), .A2(n8393), .ZN(n8390) );
  NOR2_X1 U8403 ( .A1(n7814), .A2(n7469), .ZN(n8159) );
  XOR2_X1 U8404 ( .A(n8394), .B(n8395), .Z(n8161) );
  XOR2_X1 U8405 ( .A(n8396), .B(n8397), .Z(n8394) );
  XOR2_X1 U8406 ( .A(n8398), .B(n8399), .Z(n7926) );
  XOR2_X1 U8407 ( .A(n8400), .B(n8401), .Z(n8398) );
  NAND2_X1 U8408 ( .A1(n8402), .A2(n8403), .ZN(n7498) );
  OR2_X1 U8409 ( .A1(n8403), .A2(n8402), .ZN(n7499) );
  NAND2_X1 U8410 ( .A1(n8404), .A2(n8405), .ZN(n8402) );
  NAND2_X1 U8411 ( .A1(n8406), .A2(n8407), .ZN(n8405) );
  OR2_X1 U8412 ( .A1(n8169), .A2(n8170), .ZN(n8403) );
  XNOR2_X1 U8413 ( .A(n8408), .B(n8409), .ZN(n8170) );
  XNOR2_X1 U8414 ( .A(n8410), .B(n8411), .ZN(n8409) );
  AND2_X1 U8415 ( .A1(n8412), .A2(n8413), .ZN(n8169) );
  NAND2_X1 U8416 ( .A1(n8168), .A2(n8414), .ZN(n8413) );
  OR2_X1 U8417 ( .A1(n8167), .A2(n8166), .ZN(n8414) );
  NOR2_X1 U8418 ( .A1(n8053), .A2(n7478), .ZN(n8168) );
  NAND2_X1 U8419 ( .A1(n8166), .A2(n8167), .ZN(n8412) );
  NAND2_X1 U8420 ( .A1(n8415), .A2(n8416), .ZN(n8167) );
  NAND2_X1 U8421 ( .A1(n8401), .A2(n8417), .ZN(n8416) );
  OR2_X1 U8422 ( .A1(n8400), .A2(n8399), .ZN(n8417) );
  NOR2_X1 U8423 ( .A1(n8053), .A2(n7669), .ZN(n8401) );
  NAND2_X1 U8424 ( .A1(n8399), .A2(n8400), .ZN(n8415) );
  NAND2_X1 U8425 ( .A1(n8418), .A2(n8419), .ZN(n8400) );
  NAND2_X1 U8426 ( .A1(n8396), .A2(n8420), .ZN(n8419) );
  OR2_X1 U8427 ( .A1(n8395), .A2(n8397), .ZN(n8420) );
  NAND2_X1 U8428 ( .A1(n8392), .A2(n8421), .ZN(n8396) );
  NAND2_X1 U8429 ( .A1(n8391), .A2(n8393), .ZN(n8421) );
  NAND2_X1 U8430 ( .A1(n8422), .A2(n8423), .ZN(n8393) );
  NAND2_X1 U8431 ( .A1(b_28_), .A2(a_3_), .ZN(n8423) );
  INV_X1 U8432 ( .A(n8424), .ZN(n8422) );
  XOR2_X1 U8433 ( .A(n8425), .B(n8426), .Z(n8391) );
  XOR2_X1 U8434 ( .A(n8427), .B(n8428), .Z(n8425) );
  NOR2_X1 U8435 ( .A1(n7682), .A2(n8292), .ZN(n8428) );
  NAND2_X1 U8436 ( .A1(a_3_), .A2(n8424), .ZN(n8392) );
  NAND2_X1 U8437 ( .A1(n8429), .A2(n8430), .ZN(n8424) );
  NAND2_X1 U8438 ( .A1(n8431), .A2(b_28_), .ZN(n8430) );
  NOR2_X1 U8439 ( .A1(n8432), .A2(n7682), .ZN(n8431) );
  NOR2_X1 U8440 ( .A1(n8386), .A2(n8388), .ZN(n8432) );
  NAND2_X1 U8441 ( .A1(n8386), .A2(n8388), .ZN(n8429) );
  NAND2_X1 U8442 ( .A1(n8433), .A2(n8434), .ZN(n8388) );
  NAND2_X1 U8443 ( .A1(n8385), .A2(n8435), .ZN(n8434) );
  NAND2_X1 U8444 ( .A1(n8384), .A2(n8383), .ZN(n8435) );
  NOR2_X1 U8445 ( .A1(n8053), .A2(n7455), .ZN(n8385) );
  OR2_X1 U8446 ( .A1(n8383), .A2(n8384), .ZN(n8433) );
  AND2_X1 U8447 ( .A1(n8436), .A2(n8437), .ZN(n8384) );
  NAND2_X1 U8448 ( .A1(n8438), .A2(b_28_), .ZN(n8437) );
  NOR2_X1 U8449 ( .A1(n8439), .A2(n7450), .ZN(n8438) );
  NOR2_X1 U8450 ( .A1(n8378), .A2(n8380), .ZN(n8439) );
  NAND2_X1 U8451 ( .A1(n8378), .A2(n8380), .ZN(n8436) );
  NAND2_X1 U8452 ( .A1(n8440), .A2(n8441), .ZN(n8380) );
  NAND2_X1 U8453 ( .A1(n8377), .A2(n8442), .ZN(n8441) );
  OR2_X1 U8454 ( .A1(n8376), .A2(n8375), .ZN(n8442) );
  NOR2_X1 U8455 ( .A1(n8053), .A2(n7445), .ZN(n8377) );
  NAND2_X1 U8456 ( .A1(n8375), .A2(n8376), .ZN(n8440) );
  NAND2_X1 U8457 ( .A1(n8443), .A2(n8444), .ZN(n8376) );
  NAND2_X1 U8458 ( .A1(n8445), .A2(b_28_), .ZN(n8444) );
  NOR2_X1 U8459 ( .A1(n8446), .A2(n7699), .ZN(n8445) );
  NOR2_X1 U8460 ( .A1(n8370), .A2(n8372), .ZN(n8446) );
  NAND2_X1 U8461 ( .A1(n8370), .A2(n8372), .ZN(n8443) );
  NAND2_X1 U8462 ( .A1(n8447), .A2(n8448), .ZN(n8372) );
  NAND2_X1 U8463 ( .A1(n8369), .A2(n8449), .ZN(n8448) );
  NAND2_X1 U8464 ( .A1(n8368), .A2(n8367), .ZN(n8449) );
  NOR2_X1 U8465 ( .A1(n8053), .A2(n7704), .ZN(n8369) );
  OR2_X1 U8466 ( .A1(n8367), .A2(n8368), .ZN(n8447) );
  AND2_X1 U8467 ( .A1(n8450), .A2(n8451), .ZN(n8368) );
  NAND2_X1 U8468 ( .A1(n8452), .A2(b_28_), .ZN(n8451) );
  NOR2_X1 U8469 ( .A1(n8453), .A2(n7709), .ZN(n8452) );
  NOR2_X1 U8470 ( .A1(n8363), .A2(n8364), .ZN(n8453) );
  NAND2_X1 U8471 ( .A1(n8363), .A2(n8364), .ZN(n8450) );
  NAND2_X1 U8472 ( .A1(n8454), .A2(n8455), .ZN(n8364) );
  NAND2_X1 U8473 ( .A1(n8361), .A2(n8456), .ZN(n8455) );
  OR2_X1 U8474 ( .A1(n8360), .A2(n8359), .ZN(n8456) );
  NOR2_X1 U8475 ( .A1(n8053), .A2(n7424), .ZN(n8361) );
  NAND2_X1 U8476 ( .A1(n8359), .A2(n8360), .ZN(n8454) );
  NAND2_X1 U8477 ( .A1(n8457), .A2(n8458), .ZN(n8360) );
  NAND2_X1 U8478 ( .A1(n8459), .A2(b_28_), .ZN(n8458) );
  NOR2_X1 U8479 ( .A1(n8460), .A2(n7718), .ZN(n8459) );
  NOR2_X1 U8480 ( .A1(n8355), .A2(n8356), .ZN(n8460) );
  NAND2_X1 U8481 ( .A1(n8355), .A2(n8356), .ZN(n8457) );
  NAND2_X1 U8482 ( .A1(n8461), .A2(n8462), .ZN(n8356) );
  NAND2_X1 U8483 ( .A1(n8353), .A2(n8463), .ZN(n8462) );
  OR2_X1 U8484 ( .A1(n8352), .A2(n8351), .ZN(n8463) );
  NOR2_X1 U8485 ( .A1(n8053), .A2(n7415), .ZN(n8353) );
  NAND2_X1 U8486 ( .A1(n8351), .A2(n8352), .ZN(n8461) );
  NAND2_X1 U8487 ( .A1(n8464), .A2(n8465), .ZN(n8352) );
  NAND2_X1 U8488 ( .A1(n8466), .A2(b_28_), .ZN(n8465) );
  NOR2_X1 U8489 ( .A1(n8467), .A2(n7727), .ZN(n8466) );
  NOR2_X1 U8490 ( .A1(n8346), .A2(n8348), .ZN(n8467) );
  NAND2_X1 U8491 ( .A1(n8346), .A2(n8348), .ZN(n8464) );
  NAND2_X1 U8492 ( .A1(n8468), .A2(n8469), .ZN(n8348) );
  NAND2_X1 U8493 ( .A1(n8345), .A2(n8470), .ZN(n8469) );
  OR2_X1 U8494 ( .A1(n8344), .A2(n8343), .ZN(n8470) );
  NOR2_X1 U8495 ( .A1(n8053), .A2(n7406), .ZN(n8345) );
  NAND2_X1 U8496 ( .A1(n8343), .A2(n8344), .ZN(n8468) );
  NAND2_X1 U8497 ( .A1(n8471), .A2(n8472), .ZN(n8344) );
  NAND2_X1 U8498 ( .A1(n8473), .A2(b_28_), .ZN(n8472) );
  NOR2_X1 U8499 ( .A1(n8474), .A2(n7736), .ZN(n8473) );
  NOR2_X1 U8500 ( .A1(n8339), .A2(n8340), .ZN(n8474) );
  NAND2_X1 U8501 ( .A1(n8339), .A2(n8340), .ZN(n8471) );
  NAND2_X1 U8502 ( .A1(n8475), .A2(n8476), .ZN(n8340) );
  NAND2_X1 U8503 ( .A1(n8337), .A2(n8477), .ZN(n8476) );
  OR2_X1 U8504 ( .A1(n8336), .A2(n8335), .ZN(n8477) );
  NOR2_X1 U8505 ( .A1(n8053), .A2(n7397), .ZN(n8337) );
  NAND2_X1 U8506 ( .A1(n8335), .A2(n8336), .ZN(n8475) );
  NAND2_X1 U8507 ( .A1(n8478), .A2(n8479), .ZN(n8336) );
  NAND2_X1 U8508 ( .A1(n8480), .A2(b_28_), .ZN(n8479) );
  NOR2_X1 U8509 ( .A1(n8481), .A2(n7745), .ZN(n8480) );
  NOR2_X1 U8510 ( .A1(n8331), .A2(n8332), .ZN(n8481) );
  NAND2_X1 U8511 ( .A1(n8331), .A2(n8332), .ZN(n8478) );
  NAND2_X1 U8512 ( .A1(n8482), .A2(n8483), .ZN(n8332) );
  NAND2_X1 U8513 ( .A1(n8329), .A2(n8484), .ZN(n8483) );
  OR2_X1 U8514 ( .A1(n8328), .A2(n8327), .ZN(n8484) );
  NOR2_X1 U8515 ( .A1(n8053), .A2(n7750), .ZN(n8329) );
  NAND2_X1 U8516 ( .A1(n8327), .A2(n8328), .ZN(n8482) );
  NAND2_X1 U8517 ( .A1(n8485), .A2(n8486), .ZN(n8328) );
  NAND2_X1 U8518 ( .A1(n8487), .A2(b_28_), .ZN(n8486) );
  NOR2_X1 U8519 ( .A1(n8488), .A2(n7755), .ZN(n8487) );
  NOR2_X1 U8520 ( .A1(n8323), .A2(n8324), .ZN(n8488) );
  NAND2_X1 U8521 ( .A1(n8323), .A2(n8324), .ZN(n8485) );
  NAND2_X1 U8522 ( .A1(n8489), .A2(n8490), .ZN(n8324) );
  NAND2_X1 U8523 ( .A1(n8321), .A2(n8491), .ZN(n8490) );
  OR2_X1 U8524 ( .A1(n8320), .A2(n8319), .ZN(n8491) );
  NOR2_X1 U8525 ( .A1(n8053), .A2(n7760), .ZN(n8321) );
  NAND2_X1 U8526 ( .A1(n8319), .A2(n8320), .ZN(n8489) );
  NAND2_X1 U8527 ( .A1(n8492), .A2(n8493), .ZN(n8320) );
  NAND2_X1 U8528 ( .A1(n8494), .A2(b_28_), .ZN(n8493) );
  NOR2_X1 U8529 ( .A1(n8495), .A2(n7765), .ZN(n8494) );
  NOR2_X1 U8530 ( .A1(n8314), .A2(n8316), .ZN(n8495) );
  NAND2_X1 U8531 ( .A1(n8314), .A2(n8316), .ZN(n8492) );
  NAND2_X1 U8532 ( .A1(n8496), .A2(n8497), .ZN(n8316) );
  NAND2_X1 U8533 ( .A1(n8313), .A2(n8498), .ZN(n8497) );
  OR2_X1 U8534 ( .A1(n8312), .A2(n8311), .ZN(n8498) );
  NOR2_X1 U8535 ( .A1(n8053), .A2(n8014), .ZN(n8313) );
  NAND2_X1 U8536 ( .A1(n8311), .A2(n8312), .ZN(n8496) );
  NAND2_X1 U8537 ( .A1(n8499), .A2(n8500), .ZN(n8312) );
  NAND2_X1 U8538 ( .A1(n8501), .A2(b_28_), .ZN(n8500) );
  NOR2_X1 U8539 ( .A1(n8502), .A2(n7774), .ZN(n8501) );
  NOR2_X1 U8540 ( .A1(n8307), .A2(n8309), .ZN(n8502) );
  NAND2_X1 U8541 ( .A1(n8307), .A2(n8309), .ZN(n8499) );
  NAND2_X1 U8542 ( .A1(n8503), .A2(n8504), .ZN(n8309) );
  NAND2_X1 U8543 ( .A1(n8305), .A2(n8505), .ZN(n8504) );
  OR2_X1 U8544 ( .A1(n8304), .A2(n8303), .ZN(n8505) );
  NOR2_X1 U8545 ( .A1(n8053), .A2(n8022), .ZN(n8305) );
  NAND2_X1 U8546 ( .A1(n8303), .A2(n8304), .ZN(n8503) );
  NAND2_X1 U8547 ( .A1(n8300), .A2(n8506), .ZN(n8304) );
  NAND2_X1 U8548 ( .A1(n8299), .A2(n8301), .ZN(n8506) );
  NAND2_X1 U8549 ( .A1(n8507), .A2(n8508), .ZN(n8301) );
  NAND2_X1 U8550 ( .A1(b_28_), .A2(a_26_), .ZN(n8508) );
  INV_X1 U8551 ( .A(n8509), .ZN(n8507) );
  XOR2_X1 U8552 ( .A(n8510), .B(n8511), .Z(n8299) );
  XOR2_X1 U8553 ( .A(n8512), .B(n8513), .Z(n8510) );
  NAND2_X1 U8554 ( .A1(a_26_), .A2(n8509), .ZN(n8300) );
  NAND2_X1 U8555 ( .A1(n8269), .A2(n8514), .ZN(n8509) );
  NAND2_X1 U8556 ( .A1(n8268), .A2(n8270), .ZN(n8514) );
  NAND2_X1 U8557 ( .A1(n8515), .A2(n8516), .ZN(n8270) );
  NAND2_X1 U8558 ( .A1(b_28_), .A2(a_27_), .ZN(n8516) );
  INV_X1 U8559 ( .A(n8517), .ZN(n8515) );
  XNOR2_X1 U8560 ( .A(n8518), .B(n8519), .ZN(n8268) );
  XOR2_X1 U8561 ( .A(n8520), .B(n8521), .Z(n8519) );
  NAND2_X1 U8562 ( .A1(b_27_), .A2(a_28_), .ZN(n8521) );
  NAND2_X1 U8563 ( .A1(a_27_), .A2(n8517), .ZN(n8269) );
  NAND2_X1 U8564 ( .A1(n8522), .A2(n8523), .ZN(n8517) );
  NAND2_X1 U8565 ( .A1(n8524), .A2(n8525), .ZN(n8523) );
  OR2_X1 U8566 ( .A1(n8277), .A2(n8275), .ZN(n8525) );
  INV_X1 U8567 ( .A(n8278), .ZN(n8524) );
  NAND2_X1 U8568 ( .A1(n8275), .A2(n8277), .ZN(n8522) );
  NAND2_X1 U8569 ( .A1(n8526), .A2(n8527), .ZN(n8277) );
  NAND2_X1 U8570 ( .A1(n8295), .A2(n8528), .ZN(n8527) );
  NAND2_X1 U8571 ( .A1(n8297), .A2(n8296), .ZN(n8528) );
  NOR2_X1 U8572 ( .A1(n8053), .A2(n7337), .ZN(n8295) );
  OR2_X1 U8573 ( .A1(n8296), .A2(n8297), .ZN(n8526) );
  AND2_X1 U8574 ( .A1(n8529), .A2(n8530), .ZN(n8297) );
  NAND2_X1 U8575 ( .A1(n8531), .A2(b_26_), .ZN(n8530) );
  NOR2_X1 U8576 ( .A1(n8532), .A2(n7817), .ZN(n8531) );
  NOR2_X1 U8577 ( .A1(n7816), .A2(n8292), .ZN(n8532) );
  NAND2_X1 U8578 ( .A1(n8533), .A2(b_27_), .ZN(n8529) );
  NOR2_X1 U8579 ( .A1(n8534), .A2(n8052), .ZN(n8533) );
  NOR2_X1 U8580 ( .A1(n7810), .A2(n8535), .ZN(n8534) );
  NAND2_X1 U8581 ( .A1(n8536), .A2(b_28_), .ZN(n8296) );
  XOR2_X1 U8582 ( .A(n8537), .B(n8538), .Z(n8275) );
  XOR2_X1 U8583 ( .A(n8539), .B(n8540), .Z(n8537) );
  XNOR2_X1 U8584 ( .A(n8541), .B(n8542), .ZN(n8303) );
  NAND2_X1 U8585 ( .A1(n8543), .A2(n8544), .ZN(n8541) );
  XNOR2_X1 U8586 ( .A(n8545), .B(n8546), .ZN(n8307) );
  XNOR2_X1 U8587 ( .A(n8547), .B(n8548), .ZN(n8545) );
  XNOR2_X1 U8588 ( .A(n8549), .B(n8550), .ZN(n8311) );
  XOR2_X1 U8589 ( .A(n8551), .B(n8552), .Z(n8550) );
  NAND2_X1 U8590 ( .A1(b_27_), .A2(a_24_), .ZN(n8552) );
  XOR2_X1 U8591 ( .A(n8553), .B(n8554), .Z(n8314) );
  XOR2_X1 U8592 ( .A(n8555), .B(n8556), .Z(n8553) );
  XOR2_X1 U8593 ( .A(n8557), .B(n8558), .Z(n8319) );
  XOR2_X1 U8594 ( .A(n8559), .B(n8560), .Z(n8557) );
  NOR2_X1 U8595 ( .A1(n7765), .A2(n8292), .ZN(n8560) );
  XOR2_X1 U8596 ( .A(n8561), .B(n8562), .Z(n8323) );
  XOR2_X1 U8597 ( .A(n8563), .B(n8564), .Z(n8561) );
  XOR2_X1 U8598 ( .A(n8565), .B(n8566), .Z(n8327) );
  XOR2_X1 U8599 ( .A(n8567), .B(n8568), .Z(n8565) );
  NOR2_X1 U8600 ( .A1(n7755), .A2(n8292), .ZN(n8568) );
  XNOR2_X1 U8601 ( .A(n8569), .B(n8570), .ZN(n8331) );
  XNOR2_X1 U8602 ( .A(n8571), .B(n8572), .ZN(n8570) );
  XOR2_X1 U8603 ( .A(n8573), .B(n8574), .Z(n8335) );
  XOR2_X1 U8604 ( .A(n8575), .B(n8576), .Z(n8573) );
  NOR2_X1 U8605 ( .A1(n7745), .A2(n8292), .ZN(n8576) );
  XOR2_X1 U8606 ( .A(n8577), .B(n8578), .Z(n8339) );
  XOR2_X1 U8607 ( .A(n8579), .B(n8580), .Z(n8577) );
  XNOR2_X1 U8608 ( .A(n8581), .B(n8582), .ZN(n8343) );
  XOR2_X1 U8609 ( .A(n8583), .B(n8584), .Z(n8582) );
  NAND2_X1 U8610 ( .A1(b_27_), .A2(a_16_), .ZN(n8584) );
  XOR2_X1 U8611 ( .A(n8585), .B(n8586), .Z(n8346) );
  XOR2_X1 U8612 ( .A(n8587), .B(n8588), .Z(n8585) );
  XOR2_X1 U8613 ( .A(n8589), .B(n8590), .Z(n8351) );
  XOR2_X1 U8614 ( .A(n8591), .B(n8592), .Z(n8589) );
  NOR2_X1 U8615 ( .A1(n7727), .A2(n8292), .ZN(n8592) );
  XNOR2_X1 U8616 ( .A(n8593), .B(n8594), .ZN(n8355) );
  XNOR2_X1 U8617 ( .A(n8595), .B(n8596), .ZN(n8593) );
  XOR2_X1 U8618 ( .A(n8597), .B(n8598), .Z(n8359) );
  XOR2_X1 U8619 ( .A(n8599), .B(n8600), .Z(n8597) );
  NOR2_X1 U8620 ( .A1(n7718), .A2(n8292), .ZN(n8600) );
  XOR2_X1 U8621 ( .A(n8601), .B(n8602), .Z(n8363) );
  XOR2_X1 U8622 ( .A(n8603), .B(n8604), .Z(n8601) );
  XOR2_X1 U8623 ( .A(n8605), .B(n8606), .Z(n8367) );
  XOR2_X1 U8624 ( .A(n8607), .B(n8608), .Z(n8606) );
  NAND2_X1 U8625 ( .A1(b_27_), .A2(a_10_), .ZN(n8608) );
  XOR2_X1 U8626 ( .A(n8609), .B(n8610), .Z(n8370) );
  XOR2_X1 U8627 ( .A(n8611), .B(n8612), .Z(n8609) );
  XOR2_X1 U8628 ( .A(n8613), .B(n8614), .Z(n8375) );
  XOR2_X1 U8629 ( .A(n8615), .B(n8616), .Z(n8613) );
  NOR2_X1 U8630 ( .A1(n7699), .A2(n8292), .ZN(n8616) );
  XOR2_X1 U8631 ( .A(n8617), .B(n8618), .Z(n8378) );
  XOR2_X1 U8632 ( .A(n8619), .B(n8620), .Z(n8617) );
  NOR2_X1 U8633 ( .A1(n7445), .A2(n8292), .ZN(n8620) );
  XNOR2_X1 U8634 ( .A(n8621), .B(n8622), .ZN(n8383) );
  XOR2_X1 U8635 ( .A(n8623), .B(n8624), .Z(n8621) );
  NOR2_X1 U8636 ( .A1(n7450), .A2(n8292), .ZN(n8624) );
  XNOR2_X1 U8637 ( .A(n8625), .B(n8626), .ZN(n8386) );
  XNOR2_X1 U8638 ( .A(n8627), .B(n8628), .ZN(n8625) );
  NAND2_X1 U8639 ( .A1(n8397), .A2(n8395), .ZN(n8418) );
  XNOR2_X1 U8640 ( .A(n8629), .B(n8630), .ZN(n8395) );
  NAND2_X1 U8641 ( .A1(n8631), .A2(n8632), .ZN(n8629) );
  NOR2_X1 U8642 ( .A1(n8053), .A2(n7469), .ZN(n8397) );
  XNOR2_X1 U8643 ( .A(n8633), .B(n8634), .ZN(n8399) );
  NAND2_X1 U8644 ( .A1(n8635), .A2(n8636), .ZN(n8633) );
  XOR2_X1 U8645 ( .A(n8637), .B(n8638), .Z(n8166) );
  XOR2_X1 U8646 ( .A(n8639), .B(n8640), .Z(n8637) );
  NOR2_X1 U8647 ( .A1(n7669), .A2(n8292), .ZN(n8640) );
  NAND2_X1 U8648 ( .A1(n8641), .A2(n8404), .ZN(n7503) );
  INV_X1 U8649 ( .A(n7642), .ZN(n8404) );
  NOR2_X1 U8650 ( .A1(n8407), .A2(n8406), .ZN(n7642) );
  XOR2_X1 U8651 ( .A(n8642), .B(n8643), .Z(n8406) );
  XNOR2_X1 U8652 ( .A(n8644), .B(n8645), .ZN(n8643) );
  NAND2_X1 U8653 ( .A1(n8646), .A2(n8647), .ZN(n8407) );
  NAND2_X1 U8654 ( .A1(n8410), .A2(n8648), .ZN(n8647) );
  OR2_X1 U8655 ( .A1(n8411), .A2(n8408), .ZN(n8648) );
  AND2_X1 U8656 ( .A1(n8649), .A2(n8650), .ZN(n8410) );
  NAND2_X1 U8657 ( .A1(n8651), .A2(b_27_), .ZN(n8650) );
  NOR2_X1 U8658 ( .A1(n8652), .A2(n7669), .ZN(n8651) );
  NOR2_X1 U8659 ( .A1(n8638), .A2(n8639), .ZN(n8652) );
  NAND2_X1 U8660 ( .A1(n8638), .A2(n8639), .ZN(n8649) );
  NAND2_X1 U8661 ( .A1(n8635), .A2(n8653), .ZN(n8639) );
  NAND2_X1 U8662 ( .A1(n8634), .A2(n8636), .ZN(n8653) );
  NAND2_X1 U8663 ( .A1(n8654), .A2(n8655), .ZN(n8636) );
  NAND2_X1 U8664 ( .A1(b_27_), .A2(a_2_), .ZN(n8655) );
  INV_X1 U8665 ( .A(n8656), .ZN(n8654) );
  XNOR2_X1 U8666 ( .A(n8657), .B(n8658), .ZN(n8634) );
  XNOR2_X1 U8667 ( .A(n8659), .B(n8660), .ZN(n8658) );
  NAND2_X1 U8668 ( .A1(a_2_), .A2(n8656), .ZN(n8635) );
  NAND2_X1 U8669 ( .A1(n8631), .A2(n8661), .ZN(n8656) );
  NAND2_X1 U8670 ( .A1(n8630), .A2(n8632), .ZN(n8661) );
  NAND2_X1 U8671 ( .A1(n8662), .A2(n8663), .ZN(n8632) );
  NAND2_X1 U8672 ( .A1(b_27_), .A2(a_3_), .ZN(n8663) );
  INV_X1 U8673 ( .A(n8664), .ZN(n8662) );
  XNOR2_X1 U8674 ( .A(n8665), .B(n8666), .ZN(n8630) );
  XNOR2_X1 U8675 ( .A(n8667), .B(n8668), .ZN(n8666) );
  NAND2_X1 U8676 ( .A1(a_3_), .A2(n8664), .ZN(n8631) );
  NAND2_X1 U8677 ( .A1(n8669), .A2(n8670), .ZN(n8664) );
  NAND2_X1 U8678 ( .A1(n8671), .A2(b_27_), .ZN(n8670) );
  NOR2_X1 U8679 ( .A1(n8672), .A2(n7682), .ZN(n8671) );
  NOR2_X1 U8680 ( .A1(n8426), .A2(n8427), .ZN(n8672) );
  NAND2_X1 U8681 ( .A1(n8426), .A2(n8427), .ZN(n8669) );
  NAND2_X1 U8682 ( .A1(n8673), .A2(n8674), .ZN(n8427) );
  NAND2_X1 U8683 ( .A1(n8628), .A2(n8675), .ZN(n8674) );
  NAND2_X1 U8684 ( .A1(n8627), .A2(n8626), .ZN(n8675) );
  NOR2_X1 U8685 ( .A1(n8292), .A2(n7455), .ZN(n8628) );
  OR2_X1 U8686 ( .A1(n8626), .A2(n8627), .ZN(n8673) );
  AND2_X1 U8687 ( .A1(n8676), .A2(n8677), .ZN(n8627) );
  NAND2_X1 U8688 ( .A1(n8678), .A2(b_27_), .ZN(n8677) );
  NOR2_X1 U8689 ( .A1(n8679), .A2(n7450), .ZN(n8678) );
  NOR2_X1 U8690 ( .A1(n8622), .A2(n8623), .ZN(n8679) );
  NAND2_X1 U8691 ( .A1(n8622), .A2(n8623), .ZN(n8676) );
  NAND2_X1 U8692 ( .A1(n8680), .A2(n8681), .ZN(n8623) );
  NAND2_X1 U8693 ( .A1(n8682), .A2(b_27_), .ZN(n8681) );
  NOR2_X1 U8694 ( .A1(n8683), .A2(n7445), .ZN(n8682) );
  NOR2_X1 U8695 ( .A1(n8618), .A2(n8619), .ZN(n8683) );
  NAND2_X1 U8696 ( .A1(n8618), .A2(n8619), .ZN(n8680) );
  NAND2_X1 U8697 ( .A1(n8684), .A2(n8685), .ZN(n8619) );
  NAND2_X1 U8698 ( .A1(n8686), .A2(b_27_), .ZN(n8685) );
  NOR2_X1 U8699 ( .A1(n8687), .A2(n7699), .ZN(n8686) );
  NOR2_X1 U8700 ( .A1(n8614), .A2(n8615), .ZN(n8687) );
  NAND2_X1 U8701 ( .A1(n8614), .A2(n8615), .ZN(n8684) );
  NAND2_X1 U8702 ( .A1(n8688), .A2(n8689), .ZN(n8615) );
  NAND2_X1 U8703 ( .A1(n8612), .A2(n8690), .ZN(n8689) );
  OR2_X1 U8704 ( .A1(n8611), .A2(n8610), .ZN(n8690) );
  NOR2_X1 U8705 ( .A1(n8292), .A2(n7704), .ZN(n8612) );
  NAND2_X1 U8706 ( .A1(n8610), .A2(n8611), .ZN(n8688) );
  NAND2_X1 U8707 ( .A1(n8691), .A2(n8692), .ZN(n8611) );
  NAND2_X1 U8708 ( .A1(n8693), .A2(b_27_), .ZN(n8692) );
  NOR2_X1 U8709 ( .A1(n8694), .A2(n7709), .ZN(n8693) );
  NOR2_X1 U8710 ( .A1(n8605), .A2(n8607), .ZN(n8694) );
  NAND2_X1 U8711 ( .A1(n8605), .A2(n8607), .ZN(n8691) );
  NAND2_X1 U8712 ( .A1(n8695), .A2(n8696), .ZN(n8607) );
  NAND2_X1 U8713 ( .A1(n8604), .A2(n8697), .ZN(n8696) );
  OR2_X1 U8714 ( .A1(n8603), .A2(n8602), .ZN(n8697) );
  NOR2_X1 U8715 ( .A1(n8292), .A2(n7424), .ZN(n8604) );
  NAND2_X1 U8716 ( .A1(n8602), .A2(n8603), .ZN(n8695) );
  NAND2_X1 U8717 ( .A1(n8698), .A2(n8699), .ZN(n8603) );
  NAND2_X1 U8718 ( .A1(n8700), .A2(b_27_), .ZN(n8699) );
  NOR2_X1 U8719 ( .A1(n8701), .A2(n7718), .ZN(n8700) );
  NOR2_X1 U8720 ( .A1(n8598), .A2(n8599), .ZN(n8701) );
  NAND2_X1 U8721 ( .A1(n8598), .A2(n8599), .ZN(n8698) );
  NAND2_X1 U8722 ( .A1(n8702), .A2(n8703), .ZN(n8599) );
  NAND2_X1 U8723 ( .A1(n8596), .A2(n8704), .ZN(n8703) );
  NAND2_X1 U8724 ( .A1(n8595), .A2(n8594), .ZN(n8704) );
  NOR2_X1 U8725 ( .A1(n8292), .A2(n7415), .ZN(n8596) );
  OR2_X1 U8726 ( .A1(n8594), .A2(n8595), .ZN(n8702) );
  AND2_X1 U8727 ( .A1(n8705), .A2(n8706), .ZN(n8595) );
  NAND2_X1 U8728 ( .A1(n8707), .A2(b_27_), .ZN(n8706) );
  NOR2_X1 U8729 ( .A1(n8708), .A2(n7727), .ZN(n8707) );
  NOR2_X1 U8730 ( .A1(n8590), .A2(n8591), .ZN(n8708) );
  NAND2_X1 U8731 ( .A1(n8590), .A2(n8591), .ZN(n8705) );
  NAND2_X1 U8732 ( .A1(n8709), .A2(n8710), .ZN(n8591) );
  NAND2_X1 U8733 ( .A1(n8588), .A2(n8711), .ZN(n8710) );
  OR2_X1 U8734 ( .A1(n8587), .A2(n8586), .ZN(n8711) );
  NOR2_X1 U8735 ( .A1(n8292), .A2(n7406), .ZN(n8588) );
  NAND2_X1 U8736 ( .A1(n8586), .A2(n8587), .ZN(n8709) );
  NAND2_X1 U8737 ( .A1(n8712), .A2(n8713), .ZN(n8587) );
  NAND2_X1 U8738 ( .A1(n8714), .A2(b_27_), .ZN(n8713) );
  NOR2_X1 U8739 ( .A1(n8715), .A2(n7736), .ZN(n8714) );
  NOR2_X1 U8740 ( .A1(n8581), .A2(n8583), .ZN(n8715) );
  NAND2_X1 U8741 ( .A1(n8581), .A2(n8583), .ZN(n8712) );
  NAND2_X1 U8742 ( .A1(n8716), .A2(n8717), .ZN(n8583) );
  NAND2_X1 U8743 ( .A1(n8580), .A2(n8718), .ZN(n8717) );
  OR2_X1 U8744 ( .A1(n8579), .A2(n8578), .ZN(n8718) );
  NOR2_X1 U8745 ( .A1(n8292), .A2(n7397), .ZN(n8580) );
  NAND2_X1 U8746 ( .A1(n8578), .A2(n8579), .ZN(n8716) );
  NAND2_X1 U8747 ( .A1(n8719), .A2(n8720), .ZN(n8579) );
  NAND2_X1 U8748 ( .A1(n8721), .A2(b_27_), .ZN(n8720) );
  NOR2_X1 U8749 ( .A1(n8722), .A2(n7745), .ZN(n8721) );
  NOR2_X1 U8750 ( .A1(n8574), .A2(n8575), .ZN(n8722) );
  NAND2_X1 U8751 ( .A1(n8574), .A2(n8575), .ZN(n8719) );
  NAND2_X1 U8752 ( .A1(n8723), .A2(n8724), .ZN(n8575) );
  NAND2_X1 U8753 ( .A1(n8572), .A2(n8725), .ZN(n8724) );
  OR2_X1 U8754 ( .A1(n8571), .A2(n8569), .ZN(n8725) );
  NOR2_X1 U8755 ( .A1(n8292), .A2(n7750), .ZN(n8572) );
  NAND2_X1 U8756 ( .A1(n8569), .A2(n8571), .ZN(n8723) );
  NAND2_X1 U8757 ( .A1(n8726), .A2(n8727), .ZN(n8571) );
  NAND2_X1 U8758 ( .A1(n8728), .A2(b_27_), .ZN(n8727) );
  NOR2_X1 U8759 ( .A1(n8729), .A2(n7755), .ZN(n8728) );
  NOR2_X1 U8760 ( .A1(n8566), .A2(n8567), .ZN(n8729) );
  NAND2_X1 U8761 ( .A1(n8566), .A2(n8567), .ZN(n8726) );
  NAND2_X1 U8762 ( .A1(n8730), .A2(n8731), .ZN(n8567) );
  NAND2_X1 U8763 ( .A1(n8564), .A2(n8732), .ZN(n8731) );
  OR2_X1 U8764 ( .A1(n8563), .A2(n8562), .ZN(n8732) );
  NOR2_X1 U8765 ( .A1(n8292), .A2(n7760), .ZN(n8564) );
  NAND2_X1 U8766 ( .A1(n8562), .A2(n8563), .ZN(n8730) );
  NAND2_X1 U8767 ( .A1(n8733), .A2(n8734), .ZN(n8563) );
  NAND2_X1 U8768 ( .A1(n8735), .A2(b_27_), .ZN(n8734) );
  NOR2_X1 U8769 ( .A1(n8736), .A2(n7765), .ZN(n8735) );
  NOR2_X1 U8770 ( .A1(n8558), .A2(n8559), .ZN(n8736) );
  NAND2_X1 U8771 ( .A1(n8558), .A2(n8559), .ZN(n8733) );
  NAND2_X1 U8772 ( .A1(n8737), .A2(n8738), .ZN(n8559) );
  NAND2_X1 U8773 ( .A1(n8556), .A2(n8739), .ZN(n8738) );
  OR2_X1 U8774 ( .A1(n8555), .A2(n8554), .ZN(n8739) );
  NOR2_X1 U8775 ( .A1(n8292), .A2(n8014), .ZN(n8556) );
  NAND2_X1 U8776 ( .A1(n8554), .A2(n8555), .ZN(n8737) );
  NAND2_X1 U8777 ( .A1(n8740), .A2(n8741), .ZN(n8555) );
  NAND2_X1 U8778 ( .A1(n8742), .A2(b_27_), .ZN(n8741) );
  NOR2_X1 U8779 ( .A1(n8743), .A2(n7774), .ZN(n8742) );
  NOR2_X1 U8780 ( .A1(n8549), .A2(n8551), .ZN(n8743) );
  NAND2_X1 U8781 ( .A1(n8549), .A2(n8551), .ZN(n8740) );
  NAND2_X1 U8782 ( .A1(n8744), .A2(n8745), .ZN(n8551) );
  NAND2_X1 U8783 ( .A1(n8548), .A2(n8746), .ZN(n8745) );
  NAND2_X1 U8784 ( .A1(n8547), .A2(n8546), .ZN(n8746) );
  NOR2_X1 U8785 ( .A1(n8292), .A2(n8022), .ZN(n8548) );
  OR2_X1 U8786 ( .A1(n8546), .A2(n8547), .ZN(n8744) );
  AND2_X1 U8787 ( .A1(n8543), .A2(n8747), .ZN(n8547) );
  NAND2_X1 U8788 ( .A1(n8542), .A2(n8544), .ZN(n8747) );
  NAND2_X1 U8789 ( .A1(n8748), .A2(n8749), .ZN(n8544) );
  NAND2_X1 U8790 ( .A1(b_27_), .A2(a_26_), .ZN(n8749) );
  INV_X1 U8791 ( .A(n8750), .ZN(n8748) );
  XNOR2_X1 U8792 ( .A(n8751), .B(n8752), .ZN(n8542) );
  NAND2_X1 U8793 ( .A1(n8753), .A2(n8754), .ZN(n8751) );
  NAND2_X1 U8794 ( .A1(a_26_), .A2(n8750), .ZN(n8543) );
  NAND2_X1 U8795 ( .A1(n8755), .A2(n8756), .ZN(n8750) );
  NAND2_X1 U8796 ( .A1(n8511), .A2(n8757), .ZN(n8756) );
  OR2_X1 U8797 ( .A1(n8512), .A2(n8513), .ZN(n8757) );
  XNOR2_X1 U8798 ( .A(n8758), .B(n8759), .ZN(n8511) );
  XOR2_X1 U8799 ( .A(n8760), .B(n8761), .Z(n8759) );
  NAND2_X1 U8800 ( .A1(b_26_), .A2(a_28_), .ZN(n8761) );
  NAND2_X1 U8801 ( .A1(n8513), .A2(n8512), .ZN(n8755) );
  NAND2_X1 U8802 ( .A1(n8762), .A2(n8763), .ZN(n8512) );
  NAND2_X1 U8803 ( .A1(n8764), .A2(b_27_), .ZN(n8763) );
  NOR2_X1 U8804 ( .A1(n8765), .A2(n7803), .ZN(n8764) );
  NOR2_X1 U8805 ( .A1(n8518), .A2(n8520), .ZN(n8765) );
  NAND2_X1 U8806 ( .A1(n8518), .A2(n8520), .ZN(n8762) );
  NAND2_X1 U8807 ( .A1(n8766), .A2(n8767), .ZN(n8520) );
  NAND2_X1 U8808 ( .A1(n8538), .A2(n8768), .ZN(n8767) );
  NAND2_X1 U8809 ( .A1(n8540), .A2(n8539), .ZN(n8768) );
  NOR2_X1 U8810 ( .A1(n8292), .A2(n7337), .ZN(n8538) );
  OR2_X1 U8811 ( .A1(n8539), .A2(n8540), .ZN(n8766) );
  AND2_X1 U8812 ( .A1(n8769), .A2(n8770), .ZN(n8540) );
  NAND2_X1 U8813 ( .A1(n8771), .A2(b_25_), .ZN(n8770) );
  NOR2_X1 U8814 ( .A1(n8772), .A2(n7817), .ZN(n8771) );
  NOR2_X1 U8815 ( .A1(n7816), .A2(n8535), .ZN(n8772) );
  NAND2_X1 U8816 ( .A1(n8773), .A2(b_26_), .ZN(n8769) );
  NOR2_X1 U8817 ( .A1(n8774), .A2(n8052), .ZN(n8773) );
  NOR2_X1 U8818 ( .A1(n7810), .A2(n8775), .ZN(n8774) );
  NAND2_X1 U8819 ( .A1(n8536), .A2(b_26_), .ZN(n8539) );
  NOR2_X1 U8820 ( .A1(n8055), .A2(n8292), .ZN(n8536) );
  XOR2_X1 U8821 ( .A(n8776), .B(n8777), .Z(n8518) );
  XOR2_X1 U8822 ( .A(n8778), .B(n8779), .Z(n8776) );
  XNOR2_X1 U8823 ( .A(n8780), .B(n8781), .ZN(n8546) );
  XOR2_X1 U8824 ( .A(n8782), .B(n8783), .Z(n8780) );
  XOR2_X1 U8825 ( .A(n8784), .B(n8785), .Z(n8549) );
  XOR2_X1 U8826 ( .A(n8786), .B(n8787), .Z(n8784) );
  XOR2_X1 U8827 ( .A(n8788), .B(n8789), .Z(n8554) );
  XOR2_X1 U8828 ( .A(n8790), .B(n8791), .Z(n8788) );
  NOR2_X1 U8829 ( .A1(n7774), .A2(n8535), .ZN(n8791) );
  XOR2_X1 U8830 ( .A(n8792), .B(n8793), .Z(n8558) );
  XOR2_X1 U8831 ( .A(n8794), .B(n8795), .Z(n8792) );
  XOR2_X1 U8832 ( .A(n8796), .B(n8797), .Z(n8562) );
  XOR2_X1 U8833 ( .A(n8798), .B(n8799), .Z(n8796) );
  NOR2_X1 U8834 ( .A1(n7765), .A2(n8535), .ZN(n8799) );
  XOR2_X1 U8835 ( .A(n8800), .B(n8801), .Z(n8566) );
  XOR2_X1 U8836 ( .A(n8802), .B(n8803), .Z(n8800) );
  XOR2_X1 U8837 ( .A(n8804), .B(n8805), .Z(n8569) );
  XOR2_X1 U8838 ( .A(n8806), .B(n8807), .Z(n8804) );
  NOR2_X1 U8839 ( .A1(n7755), .A2(n8535), .ZN(n8807) );
  XOR2_X1 U8840 ( .A(n8808), .B(n8809), .Z(n8574) );
  XOR2_X1 U8841 ( .A(n8810), .B(n8811), .Z(n8808) );
  XNOR2_X1 U8842 ( .A(n8812), .B(n8813), .ZN(n8578) );
  XOR2_X1 U8843 ( .A(n8814), .B(n8815), .Z(n8813) );
  NAND2_X1 U8844 ( .A1(b_26_), .A2(a_18_), .ZN(n8815) );
  XOR2_X1 U8845 ( .A(n8816), .B(n8817), .Z(n8581) );
  XOR2_X1 U8846 ( .A(n8818), .B(n8819), .Z(n8816) );
  XOR2_X1 U8847 ( .A(n8820), .B(n8821), .Z(n8586) );
  XOR2_X1 U8848 ( .A(n8822), .B(n8823), .Z(n8820) );
  NOR2_X1 U8849 ( .A1(n7736), .A2(n8535), .ZN(n8823) );
  XOR2_X1 U8850 ( .A(n8824), .B(n8825), .Z(n8590) );
  XOR2_X1 U8851 ( .A(n8826), .B(n8827), .Z(n8824) );
  XNOR2_X1 U8852 ( .A(n8828), .B(n8829), .ZN(n8594) );
  XOR2_X1 U8853 ( .A(n8830), .B(n8831), .Z(n8828) );
  NOR2_X1 U8854 ( .A1(n7727), .A2(n8535), .ZN(n8831) );
  XNOR2_X1 U8855 ( .A(n8832), .B(n8833), .ZN(n8598) );
  XNOR2_X1 U8856 ( .A(n8834), .B(n8835), .ZN(n8833) );
  XNOR2_X1 U8857 ( .A(n8836), .B(n8837), .ZN(n8602) );
  XOR2_X1 U8858 ( .A(n8838), .B(n8839), .Z(n8837) );
  NAND2_X1 U8859 ( .A1(b_26_), .A2(a_12_), .ZN(n8839) );
  XNOR2_X1 U8860 ( .A(n8840), .B(n8841), .ZN(n8605) );
  XNOR2_X1 U8861 ( .A(n8842), .B(n8843), .ZN(n8840) );
  XNOR2_X1 U8862 ( .A(n8844), .B(n8845), .ZN(n8610) );
  XOR2_X1 U8863 ( .A(n8846), .B(n8847), .Z(n8845) );
  NAND2_X1 U8864 ( .A1(b_26_), .A2(a_10_), .ZN(n8847) );
  XOR2_X1 U8865 ( .A(n8848), .B(n8849), .Z(n8614) );
  XOR2_X1 U8866 ( .A(n8850), .B(n8851), .Z(n8848) );
  XOR2_X1 U8867 ( .A(n8852), .B(n8853), .Z(n8618) );
  XOR2_X1 U8868 ( .A(n8854), .B(n8855), .Z(n8852) );
  NOR2_X1 U8869 ( .A1(n7699), .A2(n8535), .ZN(n8855) );
  XNOR2_X1 U8870 ( .A(n8856), .B(n8857), .ZN(n8622) );
  NAND2_X1 U8871 ( .A1(n8858), .A2(n8859), .ZN(n8856) );
  XNOR2_X1 U8872 ( .A(n8860), .B(n8861), .ZN(n8626) );
  XOR2_X1 U8873 ( .A(n8862), .B(n8863), .Z(n8860) );
  NOR2_X1 U8874 ( .A1(n7450), .A2(n8535), .ZN(n8863) );
  XNOR2_X1 U8875 ( .A(n8864), .B(n8865), .ZN(n8426) );
  XOR2_X1 U8876 ( .A(n8866), .B(n8867), .Z(n8865) );
  NAND2_X1 U8877 ( .A1(b_26_), .A2(a_5_), .ZN(n8867) );
  XNOR2_X1 U8878 ( .A(n8868), .B(n8869), .ZN(n8638) );
  NAND2_X1 U8879 ( .A1(n8870), .A2(n8871), .ZN(n8868) );
  NAND2_X1 U8880 ( .A1(n8408), .A2(n8411), .ZN(n8646) );
  NAND2_X1 U8881 ( .A1(b_27_), .A2(a_0_), .ZN(n8411) );
  XNOR2_X1 U8882 ( .A(n8872), .B(n8873), .ZN(n8408) );
  XOR2_X1 U8883 ( .A(n8874), .B(n8875), .Z(n8872) );
  NOR2_X1 U8884 ( .A1(n7669), .A2(n8535), .ZN(n8875) );
  NAND2_X1 U8885 ( .A1(n8876), .A2(n8877), .ZN(n8641) );
  NAND2_X1 U8886 ( .A1(n7644), .A2(n7643), .ZN(n8877) );
  NAND2_X1 U8887 ( .A1(n8876), .A2(n8878), .ZN(n7507) );
  NAND2_X1 U8888 ( .A1(n8879), .A2(n7638), .ZN(n8878) );
  INV_X1 U8889 ( .A(n8880), .ZN(n8876) );
  NAND2_X1 U8890 ( .A1(n8881), .A2(n8880), .ZN(n7506) );
  NOR2_X1 U8891 ( .A1(n7643), .A2(n7644), .ZN(n8880) );
  AND2_X1 U8892 ( .A1(n8882), .A2(n8883), .ZN(n7644) );
  NAND2_X1 U8893 ( .A1(n8645), .A2(n8884), .ZN(n8883) );
  OR2_X1 U8894 ( .A1(n8644), .A2(n8642), .ZN(n8884) );
  NOR2_X1 U8895 ( .A1(n8535), .A2(n7478), .ZN(n8645) );
  NAND2_X1 U8896 ( .A1(n8642), .A2(n8644), .ZN(n8882) );
  NAND2_X1 U8897 ( .A1(n8885), .A2(n8886), .ZN(n8644) );
  NAND2_X1 U8898 ( .A1(n8887), .A2(b_26_), .ZN(n8886) );
  NOR2_X1 U8899 ( .A1(n8888), .A2(n7669), .ZN(n8887) );
  NOR2_X1 U8900 ( .A1(n8873), .A2(n8874), .ZN(n8888) );
  NAND2_X1 U8901 ( .A1(n8873), .A2(n8874), .ZN(n8885) );
  NAND2_X1 U8902 ( .A1(n8870), .A2(n8889), .ZN(n8874) );
  NAND2_X1 U8903 ( .A1(n8869), .A2(n8871), .ZN(n8889) );
  NAND2_X1 U8904 ( .A1(n8890), .A2(n8891), .ZN(n8871) );
  NAND2_X1 U8905 ( .A1(b_26_), .A2(a_2_), .ZN(n8891) );
  INV_X1 U8906 ( .A(n8892), .ZN(n8890) );
  XOR2_X1 U8907 ( .A(n8893), .B(n8894), .Z(n8869) );
  XOR2_X1 U8908 ( .A(n8895), .B(n8896), .Z(n8893) );
  NOR2_X1 U8909 ( .A1(n7464), .A2(n8775), .ZN(n8896) );
  NAND2_X1 U8910 ( .A1(a_2_), .A2(n8892), .ZN(n8870) );
  NAND2_X1 U8911 ( .A1(n8897), .A2(n8898), .ZN(n8892) );
  NAND2_X1 U8912 ( .A1(n8660), .A2(n8899), .ZN(n8898) );
  OR2_X1 U8913 ( .A1(n8659), .A2(n8657), .ZN(n8899) );
  NOR2_X1 U8914 ( .A1(n8535), .A2(n7464), .ZN(n8660) );
  NAND2_X1 U8915 ( .A1(n8657), .A2(n8659), .ZN(n8897) );
  NAND2_X1 U8916 ( .A1(n8900), .A2(n8901), .ZN(n8659) );
  NAND2_X1 U8917 ( .A1(n8668), .A2(n8902), .ZN(n8901) );
  OR2_X1 U8918 ( .A1(n8667), .A2(n8665), .ZN(n8902) );
  NOR2_X1 U8919 ( .A1(n8535), .A2(n7682), .ZN(n8668) );
  NAND2_X1 U8920 ( .A1(n8665), .A2(n8667), .ZN(n8900) );
  NAND2_X1 U8921 ( .A1(n8903), .A2(n8904), .ZN(n8667) );
  NAND2_X1 U8922 ( .A1(n8905), .A2(b_26_), .ZN(n8904) );
  NOR2_X1 U8923 ( .A1(n8906), .A2(n7455), .ZN(n8905) );
  NOR2_X1 U8924 ( .A1(n8866), .A2(n8864), .ZN(n8906) );
  NAND2_X1 U8925 ( .A1(n8864), .A2(n8866), .ZN(n8903) );
  NAND2_X1 U8926 ( .A1(n8907), .A2(n8908), .ZN(n8866) );
  NAND2_X1 U8927 ( .A1(n8909), .A2(b_26_), .ZN(n8908) );
  NOR2_X1 U8928 ( .A1(n8910), .A2(n7450), .ZN(n8909) );
  NOR2_X1 U8929 ( .A1(n8862), .A2(n8861), .ZN(n8910) );
  NAND2_X1 U8930 ( .A1(n8861), .A2(n8862), .ZN(n8907) );
  NAND2_X1 U8931 ( .A1(n8858), .A2(n8911), .ZN(n8862) );
  NAND2_X1 U8932 ( .A1(n8857), .A2(n8859), .ZN(n8911) );
  NAND2_X1 U8933 ( .A1(n8912), .A2(n8913), .ZN(n8859) );
  NAND2_X1 U8934 ( .A1(b_26_), .A2(a_7_), .ZN(n8913) );
  INV_X1 U8935 ( .A(n8914), .ZN(n8912) );
  XOR2_X1 U8936 ( .A(n8915), .B(n8916), .Z(n8857) );
  XOR2_X1 U8937 ( .A(n8917), .B(n8918), .Z(n8915) );
  NOR2_X1 U8938 ( .A1(n7699), .A2(n8775), .ZN(n8918) );
  NAND2_X1 U8939 ( .A1(a_7_), .A2(n8914), .ZN(n8858) );
  NAND2_X1 U8940 ( .A1(n8919), .A2(n8920), .ZN(n8914) );
  NAND2_X1 U8941 ( .A1(n8921), .A2(b_26_), .ZN(n8920) );
  NOR2_X1 U8942 ( .A1(n8922), .A2(n7699), .ZN(n8921) );
  NOR2_X1 U8943 ( .A1(n8853), .A2(n8854), .ZN(n8922) );
  NAND2_X1 U8944 ( .A1(n8853), .A2(n8854), .ZN(n8919) );
  NAND2_X1 U8945 ( .A1(n8923), .A2(n8924), .ZN(n8854) );
  NAND2_X1 U8946 ( .A1(n8851), .A2(n8925), .ZN(n8924) );
  OR2_X1 U8947 ( .A1(n8849), .A2(n8850), .ZN(n8925) );
  NOR2_X1 U8948 ( .A1(n8535), .A2(n7704), .ZN(n8851) );
  NAND2_X1 U8949 ( .A1(n8849), .A2(n8850), .ZN(n8923) );
  NAND2_X1 U8950 ( .A1(n8926), .A2(n8927), .ZN(n8850) );
  NAND2_X1 U8951 ( .A1(n8928), .A2(b_26_), .ZN(n8927) );
  NOR2_X1 U8952 ( .A1(n8929), .A2(n7709), .ZN(n8928) );
  NOR2_X1 U8953 ( .A1(n8844), .A2(n8846), .ZN(n8929) );
  NAND2_X1 U8954 ( .A1(n8844), .A2(n8846), .ZN(n8926) );
  NAND2_X1 U8955 ( .A1(n8930), .A2(n8931), .ZN(n8846) );
  NAND2_X1 U8956 ( .A1(n8843), .A2(n8932), .ZN(n8931) );
  NAND2_X1 U8957 ( .A1(n8842), .A2(n8841), .ZN(n8932) );
  NOR2_X1 U8958 ( .A1(n8535), .A2(n7424), .ZN(n8843) );
  OR2_X1 U8959 ( .A1(n8841), .A2(n8842), .ZN(n8930) );
  AND2_X1 U8960 ( .A1(n8933), .A2(n8934), .ZN(n8842) );
  NAND2_X1 U8961 ( .A1(n8935), .A2(b_26_), .ZN(n8934) );
  NOR2_X1 U8962 ( .A1(n8936), .A2(n7718), .ZN(n8935) );
  NOR2_X1 U8963 ( .A1(n8836), .A2(n8838), .ZN(n8936) );
  NAND2_X1 U8964 ( .A1(n8836), .A2(n8838), .ZN(n8933) );
  NAND2_X1 U8965 ( .A1(n8937), .A2(n8938), .ZN(n8838) );
  NAND2_X1 U8966 ( .A1(n8835), .A2(n8939), .ZN(n8938) );
  OR2_X1 U8967 ( .A1(n8832), .A2(n8834), .ZN(n8939) );
  NOR2_X1 U8968 ( .A1(n8535), .A2(n7415), .ZN(n8835) );
  NAND2_X1 U8969 ( .A1(n8832), .A2(n8834), .ZN(n8937) );
  NAND2_X1 U8970 ( .A1(n8940), .A2(n8941), .ZN(n8834) );
  NAND2_X1 U8971 ( .A1(n8942), .A2(b_26_), .ZN(n8941) );
  NOR2_X1 U8972 ( .A1(n8943), .A2(n7727), .ZN(n8942) );
  NOR2_X1 U8973 ( .A1(n8830), .A2(n8829), .ZN(n8943) );
  NAND2_X1 U8974 ( .A1(n8829), .A2(n8830), .ZN(n8940) );
  NAND2_X1 U8975 ( .A1(n8944), .A2(n8945), .ZN(n8830) );
  NAND2_X1 U8976 ( .A1(n8827), .A2(n8946), .ZN(n8945) );
  OR2_X1 U8977 ( .A1(n8825), .A2(n8826), .ZN(n8946) );
  NOR2_X1 U8978 ( .A1(n8535), .A2(n7406), .ZN(n8827) );
  NAND2_X1 U8979 ( .A1(n8825), .A2(n8826), .ZN(n8944) );
  NAND2_X1 U8980 ( .A1(n8947), .A2(n8948), .ZN(n8826) );
  NAND2_X1 U8981 ( .A1(n8949), .A2(b_26_), .ZN(n8948) );
  NOR2_X1 U8982 ( .A1(n8950), .A2(n7736), .ZN(n8949) );
  NOR2_X1 U8983 ( .A1(n8821), .A2(n8822), .ZN(n8950) );
  NAND2_X1 U8984 ( .A1(n8821), .A2(n8822), .ZN(n8947) );
  NAND2_X1 U8985 ( .A1(n8951), .A2(n8952), .ZN(n8822) );
  NAND2_X1 U8986 ( .A1(n8819), .A2(n8953), .ZN(n8952) );
  OR2_X1 U8987 ( .A1(n8817), .A2(n8818), .ZN(n8953) );
  NOR2_X1 U8988 ( .A1(n8535), .A2(n7397), .ZN(n8819) );
  NAND2_X1 U8989 ( .A1(n8817), .A2(n8818), .ZN(n8951) );
  NAND2_X1 U8990 ( .A1(n8954), .A2(n8955), .ZN(n8818) );
  NAND2_X1 U8991 ( .A1(n8956), .A2(b_26_), .ZN(n8955) );
  NOR2_X1 U8992 ( .A1(n8957), .A2(n7745), .ZN(n8956) );
  NOR2_X1 U8993 ( .A1(n8812), .A2(n8814), .ZN(n8957) );
  NAND2_X1 U8994 ( .A1(n8812), .A2(n8814), .ZN(n8954) );
  NAND2_X1 U8995 ( .A1(n8958), .A2(n8959), .ZN(n8814) );
  NAND2_X1 U8996 ( .A1(n8811), .A2(n8960), .ZN(n8959) );
  OR2_X1 U8997 ( .A1(n8809), .A2(n8810), .ZN(n8960) );
  NOR2_X1 U8998 ( .A1(n8535), .A2(n7750), .ZN(n8811) );
  NAND2_X1 U8999 ( .A1(n8809), .A2(n8810), .ZN(n8958) );
  NAND2_X1 U9000 ( .A1(n8961), .A2(n8962), .ZN(n8810) );
  NAND2_X1 U9001 ( .A1(n8963), .A2(b_26_), .ZN(n8962) );
  NOR2_X1 U9002 ( .A1(n8964), .A2(n7755), .ZN(n8963) );
  NOR2_X1 U9003 ( .A1(n8805), .A2(n8806), .ZN(n8964) );
  NAND2_X1 U9004 ( .A1(n8805), .A2(n8806), .ZN(n8961) );
  NAND2_X1 U9005 ( .A1(n8965), .A2(n8966), .ZN(n8806) );
  NAND2_X1 U9006 ( .A1(n8803), .A2(n8967), .ZN(n8966) );
  OR2_X1 U9007 ( .A1(n8801), .A2(n8802), .ZN(n8967) );
  NOR2_X1 U9008 ( .A1(n8535), .A2(n7760), .ZN(n8803) );
  NAND2_X1 U9009 ( .A1(n8801), .A2(n8802), .ZN(n8965) );
  NAND2_X1 U9010 ( .A1(n8968), .A2(n8969), .ZN(n8802) );
  NAND2_X1 U9011 ( .A1(n8970), .A2(b_26_), .ZN(n8969) );
  NOR2_X1 U9012 ( .A1(n8971), .A2(n7765), .ZN(n8970) );
  NOR2_X1 U9013 ( .A1(n8797), .A2(n8798), .ZN(n8971) );
  NAND2_X1 U9014 ( .A1(n8797), .A2(n8798), .ZN(n8968) );
  NAND2_X1 U9015 ( .A1(n8972), .A2(n8973), .ZN(n8798) );
  NAND2_X1 U9016 ( .A1(n8795), .A2(n8974), .ZN(n8973) );
  OR2_X1 U9017 ( .A1(n8793), .A2(n8794), .ZN(n8974) );
  NOR2_X1 U9018 ( .A1(n8535), .A2(n8014), .ZN(n8795) );
  NAND2_X1 U9019 ( .A1(n8793), .A2(n8794), .ZN(n8972) );
  NAND2_X1 U9020 ( .A1(n8975), .A2(n8976), .ZN(n8794) );
  NAND2_X1 U9021 ( .A1(n8977), .A2(b_26_), .ZN(n8976) );
  NOR2_X1 U9022 ( .A1(n8978), .A2(n7774), .ZN(n8977) );
  NOR2_X1 U9023 ( .A1(n8789), .A2(n8790), .ZN(n8978) );
  NAND2_X1 U9024 ( .A1(n8789), .A2(n8790), .ZN(n8975) );
  NAND2_X1 U9025 ( .A1(n8979), .A2(n8980), .ZN(n8790) );
  NAND2_X1 U9026 ( .A1(n8787), .A2(n8981), .ZN(n8980) );
  OR2_X1 U9027 ( .A1(n8785), .A2(n8786), .ZN(n8981) );
  NOR2_X1 U9028 ( .A1(n8535), .A2(n8022), .ZN(n8787) );
  NAND2_X1 U9029 ( .A1(n8785), .A2(n8786), .ZN(n8979) );
  NAND2_X1 U9030 ( .A1(n8982), .A2(n8983), .ZN(n8786) );
  NAND2_X1 U9031 ( .A1(n8783), .A2(n8984), .ZN(n8983) );
  OR2_X1 U9032 ( .A1(n8781), .A2(n8782), .ZN(n8984) );
  INV_X1 U9033 ( .A(n8985), .ZN(n8783) );
  NAND2_X1 U9034 ( .A1(n8781), .A2(n8782), .ZN(n8982) );
  NAND2_X1 U9035 ( .A1(n8753), .A2(n8986), .ZN(n8782) );
  NAND2_X1 U9036 ( .A1(n8752), .A2(n8754), .ZN(n8986) );
  NAND2_X1 U9037 ( .A1(n8987), .A2(n8988), .ZN(n8754) );
  NAND2_X1 U9038 ( .A1(b_26_), .A2(a_27_), .ZN(n8988) );
  INV_X1 U9039 ( .A(n8989), .ZN(n8987) );
  XNOR2_X1 U9040 ( .A(n8990), .B(n8991), .ZN(n8752) );
  XOR2_X1 U9041 ( .A(n8992), .B(n8993), .Z(n8991) );
  NAND2_X1 U9042 ( .A1(b_25_), .A2(a_28_), .ZN(n8993) );
  NAND2_X1 U9043 ( .A1(a_27_), .A2(n8989), .ZN(n8753) );
  NAND2_X1 U9044 ( .A1(n8994), .A2(n8995), .ZN(n8989) );
  NAND2_X1 U9045 ( .A1(n8996), .A2(b_26_), .ZN(n8995) );
  NOR2_X1 U9046 ( .A1(n8997), .A2(n7803), .ZN(n8996) );
  NOR2_X1 U9047 ( .A1(n8758), .A2(n8760), .ZN(n8997) );
  NAND2_X1 U9048 ( .A1(n8758), .A2(n8760), .ZN(n8994) );
  NAND2_X1 U9049 ( .A1(n8998), .A2(n8999), .ZN(n8760) );
  NAND2_X1 U9050 ( .A1(n8777), .A2(n9000), .ZN(n8999) );
  NAND2_X1 U9051 ( .A1(n8779), .A2(n8778), .ZN(n9000) );
  NOR2_X1 U9052 ( .A1(n8535), .A2(n7337), .ZN(n8777) );
  OR2_X1 U9053 ( .A1(n8778), .A2(n8779), .ZN(n8998) );
  AND2_X1 U9054 ( .A1(n9001), .A2(n9002), .ZN(n8779) );
  NAND2_X1 U9055 ( .A1(n9003), .A2(b_24_), .ZN(n9002) );
  NOR2_X1 U9056 ( .A1(n9004), .A2(n7817), .ZN(n9003) );
  NOR2_X1 U9057 ( .A1(n7816), .A2(n8775), .ZN(n9004) );
  NAND2_X1 U9058 ( .A1(n9005), .A2(b_25_), .ZN(n9001) );
  NOR2_X1 U9059 ( .A1(n9006), .A2(n8052), .ZN(n9005) );
  NOR2_X1 U9060 ( .A1(n7810), .A2(n9007), .ZN(n9006) );
  NAND2_X1 U9061 ( .A1(n9008), .A2(b_26_), .ZN(n8778) );
  NOR2_X1 U9062 ( .A1(n8055), .A2(n8775), .ZN(n9008) );
  XOR2_X1 U9063 ( .A(n9009), .B(n9010), .Z(n8758) );
  XOR2_X1 U9064 ( .A(n9011), .B(n9012), .Z(n9009) );
  XNOR2_X1 U9065 ( .A(n9013), .B(n9014), .ZN(n8781) );
  NAND2_X1 U9066 ( .A1(n9015), .A2(n9016), .ZN(n9013) );
  XNOR2_X1 U9067 ( .A(n9017), .B(n9018), .ZN(n8785) );
  NAND2_X1 U9068 ( .A1(n9019), .A2(n9020), .ZN(n9017) );
  XOR2_X1 U9069 ( .A(n9021), .B(n9022), .Z(n8789) );
  XOR2_X1 U9070 ( .A(n9023), .B(n9024), .Z(n9021) );
  XOR2_X1 U9071 ( .A(n9025), .B(n9026), .Z(n8793) );
  XNOR2_X1 U9072 ( .A(n9027), .B(n9028), .ZN(n9025) );
  NAND2_X1 U9073 ( .A1(b_25_), .A2(a_24_), .ZN(n9027) );
  XOR2_X1 U9074 ( .A(n9029), .B(n9030), .Z(n8797) );
  XOR2_X1 U9075 ( .A(n9031), .B(n9032), .Z(n9029) );
  XNOR2_X1 U9076 ( .A(n9033), .B(n9034), .ZN(n8801) );
  XOR2_X1 U9077 ( .A(n9035), .B(n9036), .Z(n9034) );
  NAND2_X1 U9078 ( .A1(b_25_), .A2(a_22_), .ZN(n9036) );
  XNOR2_X1 U9079 ( .A(n9037), .B(n9038), .ZN(n8805) );
  XNOR2_X1 U9080 ( .A(n9039), .B(n9040), .ZN(n9038) );
  XNOR2_X1 U9081 ( .A(n9041), .B(n9042), .ZN(n8809) );
  XOR2_X1 U9082 ( .A(n9043), .B(n9044), .Z(n9042) );
  NAND2_X1 U9083 ( .A1(b_25_), .A2(a_20_), .ZN(n9044) );
  XNOR2_X1 U9084 ( .A(n9045), .B(n9046), .ZN(n8812) );
  XNOR2_X1 U9085 ( .A(n9047), .B(n9048), .ZN(n9046) );
  XOR2_X1 U9086 ( .A(n9049), .B(n9050), .Z(n8817) );
  XOR2_X1 U9087 ( .A(n9051), .B(n9052), .Z(n9049) );
  NOR2_X1 U9088 ( .A1(n7745), .A2(n8775), .ZN(n9052) );
  XNOR2_X1 U9089 ( .A(n9053), .B(n9054), .ZN(n8821) );
  XNOR2_X1 U9090 ( .A(n9055), .B(n9056), .ZN(n9054) );
  XOR2_X1 U9091 ( .A(n9057), .B(n9058), .Z(n8825) );
  XOR2_X1 U9092 ( .A(n9059), .B(n9060), .Z(n9057) );
  NOR2_X1 U9093 ( .A1(n7736), .A2(n8775), .ZN(n9060) );
  XNOR2_X1 U9094 ( .A(n9061), .B(n9062), .ZN(n8829) );
  XNOR2_X1 U9095 ( .A(n9063), .B(n9064), .ZN(n9061) );
  XNOR2_X1 U9096 ( .A(n9065), .B(n9066), .ZN(n8832) );
  XOR2_X1 U9097 ( .A(n9067), .B(n9068), .Z(n9066) );
  NAND2_X1 U9098 ( .A1(b_25_), .A2(a_14_), .ZN(n9068) );
  XOR2_X1 U9099 ( .A(n9069), .B(n9070), .Z(n8836) );
  XOR2_X1 U9100 ( .A(n9071), .B(n9072), .Z(n9069) );
  XNOR2_X1 U9101 ( .A(n9073), .B(n9074), .ZN(n8841) );
  XOR2_X1 U9102 ( .A(n9075), .B(n9076), .Z(n9073) );
  NOR2_X1 U9103 ( .A1(n7718), .A2(n8775), .ZN(n9076) );
  XOR2_X1 U9104 ( .A(n9077), .B(n9078), .Z(n8844) );
  XOR2_X1 U9105 ( .A(n9079), .B(n9080), .Z(n9077) );
  NOR2_X1 U9106 ( .A1(n7424), .A2(n8775), .ZN(n9080) );
  XOR2_X1 U9107 ( .A(n9081), .B(n9082), .Z(n8849) );
  XOR2_X1 U9108 ( .A(n9083), .B(n9084), .Z(n9081) );
  NOR2_X1 U9109 ( .A1(n7709), .A2(n8775), .ZN(n9084) );
  XOR2_X1 U9110 ( .A(n9085), .B(n9086), .Z(n8853) );
  XOR2_X1 U9111 ( .A(n9087), .B(n9088), .Z(n9085) );
  XNOR2_X1 U9112 ( .A(n9089), .B(n9090), .ZN(n8861) );
  NAND2_X1 U9113 ( .A1(n9091), .A2(n9092), .ZN(n9089) );
  XNOR2_X1 U9114 ( .A(n9093), .B(n9094), .ZN(n8864) );
  XNOR2_X1 U9115 ( .A(n9095), .B(n9096), .ZN(n9093) );
  XOR2_X1 U9116 ( .A(n9097), .B(n9098), .Z(n8665) );
  XOR2_X1 U9117 ( .A(n9099), .B(n9100), .Z(n9097) );
  NOR2_X1 U9118 ( .A1(n7455), .A2(n8775), .ZN(n9100) );
  XOR2_X1 U9119 ( .A(n9101), .B(n9102), .Z(n8657) );
  XOR2_X1 U9120 ( .A(n9103), .B(n9104), .Z(n9101) );
  NOR2_X1 U9121 ( .A1(n7682), .A2(n8775), .ZN(n9104) );
  XNOR2_X1 U9122 ( .A(n9105), .B(n9106), .ZN(n8873) );
  NAND2_X1 U9123 ( .A1(n9107), .A2(n9108), .ZN(n9105) );
  XOR2_X1 U9124 ( .A(n9109), .B(n9110), .Z(n8642) );
  XOR2_X1 U9125 ( .A(n9111), .B(n9112), .Z(n9109) );
  NOR2_X1 U9126 ( .A1(n7669), .A2(n8775), .ZN(n9112) );
  XOR2_X1 U9127 ( .A(n9113), .B(n9114), .Z(n7643) );
  XNOR2_X1 U9128 ( .A(n9115), .B(n9116), .ZN(n9113) );
  AND2_X1 U9129 ( .A1(n7638), .A2(n8879), .ZN(n8881) );
  NAND2_X1 U9130 ( .A1(n9117), .A2(n9118), .ZN(n8879) );
  XOR2_X1 U9131 ( .A(n9119), .B(n9120), .Z(n9118) );
  NOR2_X1 U9132 ( .A1(n9121), .A2(n9122), .ZN(n9117) );
  NOR2_X1 U9133 ( .A1(n9115), .A2(n9114), .ZN(n9122) );
  INV_X1 U9134 ( .A(n9123), .ZN(n9121) );
  OR2_X1 U9135 ( .A1(n7638), .A2(n7637), .ZN(n7511) );
  XNOR2_X1 U9136 ( .A(n7634), .B(n7633), .ZN(n7637) );
  NAND2_X1 U9137 ( .A1(n9124), .A2(n9125), .ZN(n7638) );
  NAND2_X1 U9138 ( .A1(n9126), .A2(n9123), .ZN(n9125) );
  NAND2_X1 U9139 ( .A1(n9116), .A2(n9127), .ZN(n9123) );
  NAND2_X1 U9140 ( .A1(n9115), .A2(n9114), .ZN(n9127) );
  NOR2_X1 U9141 ( .A1(n8775), .A2(n7478), .ZN(n9116) );
  OR2_X1 U9142 ( .A1(n9114), .A2(n9115), .ZN(n9126) );
  AND2_X1 U9143 ( .A1(n9128), .A2(n9129), .ZN(n9115) );
  NAND2_X1 U9144 ( .A1(n9130), .A2(b_25_), .ZN(n9129) );
  NOR2_X1 U9145 ( .A1(n9131), .A2(n7669), .ZN(n9130) );
  NOR2_X1 U9146 ( .A1(n9110), .A2(n9111), .ZN(n9131) );
  NAND2_X1 U9147 ( .A1(n9110), .A2(n9111), .ZN(n9128) );
  NAND2_X1 U9148 ( .A1(n9107), .A2(n9132), .ZN(n9111) );
  NAND2_X1 U9149 ( .A1(n9106), .A2(n9108), .ZN(n9132) );
  NAND2_X1 U9150 ( .A1(n9133), .A2(n9134), .ZN(n9108) );
  NAND2_X1 U9151 ( .A1(b_25_), .A2(a_2_), .ZN(n9134) );
  INV_X1 U9152 ( .A(n9135), .ZN(n9133) );
  XNOR2_X1 U9153 ( .A(n9136), .B(n9137), .ZN(n9106) );
  NAND2_X1 U9154 ( .A1(n9138), .A2(n9139), .ZN(n9136) );
  NAND2_X1 U9155 ( .A1(a_2_), .A2(n9135), .ZN(n9107) );
  NAND2_X1 U9156 ( .A1(n9140), .A2(n9141), .ZN(n9135) );
  NAND2_X1 U9157 ( .A1(n9142), .A2(b_25_), .ZN(n9141) );
  NOR2_X1 U9158 ( .A1(n9143), .A2(n7464), .ZN(n9142) );
  NOR2_X1 U9159 ( .A1(n8894), .A2(n8895), .ZN(n9143) );
  NAND2_X1 U9160 ( .A1(n8894), .A2(n8895), .ZN(n9140) );
  NAND2_X1 U9161 ( .A1(n9144), .A2(n9145), .ZN(n8895) );
  NAND2_X1 U9162 ( .A1(n9146), .A2(b_25_), .ZN(n9145) );
  NOR2_X1 U9163 ( .A1(n9147), .A2(n7682), .ZN(n9146) );
  NOR2_X1 U9164 ( .A1(n9102), .A2(n9103), .ZN(n9147) );
  NAND2_X1 U9165 ( .A1(n9102), .A2(n9103), .ZN(n9144) );
  NAND2_X1 U9166 ( .A1(n9148), .A2(n9149), .ZN(n9103) );
  NAND2_X1 U9167 ( .A1(n9150), .A2(b_25_), .ZN(n9149) );
  NOR2_X1 U9168 ( .A1(n9151), .A2(n7455), .ZN(n9150) );
  NOR2_X1 U9169 ( .A1(n9098), .A2(n9099), .ZN(n9151) );
  NAND2_X1 U9170 ( .A1(n9098), .A2(n9099), .ZN(n9148) );
  NAND2_X1 U9171 ( .A1(n9152), .A2(n9153), .ZN(n9099) );
  NAND2_X1 U9172 ( .A1(n9095), .A2(n9154), .ZN(n9153) );
  NAND2_X1 U9173 ( .A1(n9094), .A2(n9096), .ZN(n9154) );
  NAND2_X1 U9174 ( .A1(n9091), .A2(n9155), .ZN(n9095) );
  NAND2_X1 U9175 ( .A1(n9090), .A2(n9092), .ZN(n9155) );
  NAND2_X1 U9176 ( .A1(n9156), .A2(n9157), .ZN(n9092) );
  NAND2_X1 U9177 ( .A1(b_25_), .A2(a_7_), .ZN(n9157) );
  INV_X1 U9178 ( .A(n9158), .ZN(n9156) );
  XNOR2_X1 U9179 ( .A(n9159), .B(n9160), .ZN(n9090) );
  XOR2_X1 U9180 ( .A(n9161), .B(n9162), .Z(n9160) );
  NAND2_X1 U9181 ( .A1(b_24_), .A2(a_8_), .ZN(n9162) );
  NAND2_X1 U9182 ( .A1(a_7_), .A2(n9158), .ZN(n9091) );
  NAND2_X1 U9183 ( .A1(n9163), .A2(n9164), .ZN(n9158) );
  NAND2_X1 U9184 ( .A1(n9165), .A2(b_25_), .ZN(n9164) );
  NOR2_X1 U9185 ( .A1(n9166), .A2(n7699), .ZN(n9165) );
  NOR2_X1 U9186 ( .A1(n8916), .A2(n8917), .ZN(n9166) );
  NAND2_X1 U9187 ( .A1(n8916), .A2(n8917), .ZN(n9163) );
  NAND2_X1 U9188 ( .A1(n9167), .A2(n9168), .ZN(n8917) );
  NAND2_X1 U9189 ( .A1(n9088), .A2(n9169), .ZN(n9168) );
  OR2_X1 U9190 ( .A1(n9087), .A2(n9086), .ZN(n9169) );
  NOR2_X1 U9191 ( .A1(n8775), .A2(n7704), .ZN(n9088) );
  NAND2_X1 U9192 ( .A1(n9086), .A2(n9087), .ZN(n9167) );
  NAND2_X1 U9193 ( .A1(n9170), .A2(n9171), .ZN(n9087) );
  NAND2_X1 U9194 ( .A1(n9172), .A2(b_25_), .ZN(n9171) );
  NOR2_X1 U9195 ( .A1(n9173), .A2(n7709), .ZN(n9172) );
  NOR2_X1 U9196 ( .A1(n9082), .A2(n9083), .ZN(n9173) );
  NAND2_X1 U9197 ( .A1(n9082), .A2(n9083), .ZN(n9170) );
  NAND2_X1 U9198 ( .A1(n9174), .A2(n9175), .ZN(n9083) );
  NAND2_X1 U9199 ( .A1(n9176), .A2(b_25_), .ZN(n9175) );
  NOR2_X1 U9200 ( .A1(n9177), .A2(n7424), .ZN(n9176) );
  NOR2_X1 U9201 ( .A1(n9078), .A2(n9079), .ZN(n9177) );
  NAND2_X1 U9202 ( .A1(n9078), .A2(n9079), .ZN(n9174) );
  NAND2_X1 U9203 ( .A1(n9178), .A2(n9179), .ZN(n9079) );
  NAND2_X1 U9204 ( .A1(n9180), .A2(b_25_), .ZN(n9179) );
  NOR2_X1 U9205 ( .A1(n9181), .A2(n7718), .ZN(n9180) );
  NOR2_X1 U9206 ( .A1(n9074), .A2(n9075), .ZN(n9181) );
  NAND2_X1 U9207 ( .A1(n9074), .A2(n9075), .ZN(n9178) );
  NAND2_X1 U9208 ( .A1(n9182), .A2(n9183), .ZN(n9075) );
  NAND2_X1 U9209 ( .A1(n9072), .A2(n9184), .ZN(n9183) );
  OR2_X1 U9210 ( .A1(n9071), .A2(n9070), .ZN(n9184) );
  NOR2_X1 U9211 ( .A1(n8775), .A2(n7415), .ZN(n9072) );
  NAND2_X1 U9212 ( .A1(n9070), .A2(n9071), .ZN(n9182) );
  NAND2_X1 U9213 ( .A1(n9185), .A2(n9186), .ZN(n9071) );
  NAND2_X1 U9214 ( .A1(n9187), .A2(b_25_), .ZN(n9186) );
  NOR2_X1 U9215 ( .A1(n9188), .A2(n7727), .ZN(n9187) );
  NOR2_X1 U9216 ( .A1(n9065), .A2(n9067), .ZN(n9188) );
  NAND2_X1 U9217 ( .A1(n9065), .A2(n9067), .ZN(n9185) );
  NAND2_X1 U9218 ( .A1(n9189), .A2(n9190), .ZN(n9067) );
  NAND2_X1 U9219 ( .A1(n9064), .A2(n9191), .ZN(n9190) );
  NAND2_X1 U9220 ( .A1(n9063), .A2(n9062), .ZN(n9191) );
  NOR2_X1 U9221 ( .A1(n8775), .A2(n7406), .ZN(n9064) );
  OR2_X1 U9222 ( .A1(n9062), .A2(n9063), .ZN(n9189) );
  AND2_X1 U9223 ( .A1(n9192), .A2(n9193), .ZN(n9063) );
  NAND2_X1 U9224 ( .A1(n9194), .A2(b_25_), .ZN(n9193) );
  NOR2_X1 U9225 ( .A1(n9195), .A2(n7736), .ZN(n9194) );
  NOR2_X1 U9226 ( .A1(n9058), .A2(n9059), .ZN(n9195) );
  NAND2_X1 U9227 ( .A1(n9058), .A2(n9059), .ZN(n9192) );
  NAND2_X1 U9228 ( .A1(n9196), .A2(n9197), .ZN(n9059) );
  NAND2_X1 U9229 ( .A1(n9056), .A2(n9198), .ZN(n9197) );
  OR2_X1 U9230 ( .A1(n9055), .A2(n9053), .ZN(n9198) );
  NOR2_X1 U9231 ( .A1(n8775), .A2(n7397), .ZN(n9056) );
  NAND2_X1 U9232 ( .A1(n9053), .A2(n9055), .ZN(n9196) );
  NAND2_X1 U9233 ( .A1(n9199), .A2(n9200), .ZN(n9055) );
  NAND2_X1 U9234 ( .A1(n9201), .A2(b_25_), .ZN(n9200) );
  NOR2_X1 U9235 ( .A1(n9202), .A2(n7745), .ZN(n9201) );
  NOR2_X1 U9236 ( .A1(n9050), .A2(n9051), .ZN(n9202) );
  NAND2_X1 U9237 ( .A1(n9050), .A2(n9051), .ZN(n9199) );
  NAND2_X1 U9238 ( .A1(n9203), .A2(n9204), .ZN(n9051) );
  NAND2_X1 U9239 ( .A1(n9048), .A2(n9205), .ZN(n9204) );
  OR2_X1 U9240 ( .A1(n9047), .A2(n9045), .ZN(n9205) );
  NOR2_X1 U9241 ( .A1(n8775), .A2(n7750), .ZN(n9048) );
  NAND2_X1 U9242 ( .A1(n9045), .A2(n9047), .ZN(n9203) );
  NAND2_X1 U9243 ( .A1(n9206), .A2(n9207), .ZN(n9047) );
  NAND2_X1 U9244 ( .A1(n9208), .A2(b_25_), .ZN(n9207) );
  NOR2_X1 U9245 ( .A1(n9209), .A2(n7755), .ZN(n9208) );
  NOR2_X1 U9246 ( .A1(n9041), .A2(n9043), .ZN(n9209) );
  NAND2_X1 U9247 ( .A1(n9041), .A2(n9043), .ZN(n9206) );
  NAND2_X1 U9248 ( .A1(n9210), .A2(n9211), .ZN(n9043) );
  NAND2_X1 U9249 ( .A1(n9040), .A2(n9212), .ZN(n9211) );
  OR2_X1 U9250 ( .A1(n9039), .A2(n9037), .ZN(n9212) );
  NOR2_X1 U9251 ( .A1(n8775), .A2(n7760), .ZN(n9040) );
  NAND2_X1 U9252 ( .A1(n9037), .A2(n9039), .ZN(n9210) );
  NAND2_X1 U9253 ( .A1(n9213), .A2(n9214), .ZN(n9039) );
  NAND2_X1 U9254 ( .A1(n9215), .A2(b_25_), .ZN(n9214) );
  NOR2_X1 U9255 ( .A1(n9216), .A2(n7765), .ZN(n9215) );
  NOR2_X1 U9256 ( .A1(n9033), .A2(n9035), .ZN(n9216) );
  NAND2_X1 U9257 ( .A1(n9033), .A2(n9035), .ZN(n9213) );
  NAND2_X1 U9258 ( .A1(n9217), .A2(n9218), .ZN(n9035) );
  NAND2_X1 U9259 ( .A1(n9032), .A2(n9219), .ZN(n9218) );
  OR2_X1 U9260 ( .A1(n9031), .A2(n9030), .ZN(n9219) );
  NOR2_X1 U9261 ( .A1(n8775), .A2(n8014), .ZN(n9032) );
  NAND2_X1 U9262 ( .A1(n9030), .A2(n9031), .ZN(n9217) );
  NAND2_X1 U9263 ( .A1(n9220), .A2(n9221), .ZN(n9031) );
  NAND2_X1 U9264 ( .A1(n9222), .A2(b_25_), .ZN(n9221) );
  NOR2_X1 U9265 ( .A1(n9223), .A2(n7774), .ZN(n9222) );
  NOR2_X1 U9266 ( .A1(n9026), .A2(n9028), .ZN(n9223) );
  NAND2_X1 U9267 ( .A1(n9026), .A2(n9028), .ZN(n9220) );
  NAND2_X1 U9268 ( .A1(n9224), .A2(n9225), .ZN(n9028) );
  NAND2_X1 U9269 ( .A1(n9024), .A2(n9226), .ZN(n9225) );
  OR2_X1 U9270 ( .A1(n9023), .A2(n9022), .ZN(n9226) );
  NAND2_X1 U9271 ( .A1(n9022), .A2(n9023), .ZN(n9224) );
  NAND2_X1 U9272 ( .A1(n9019), .A2(n9227), .ZN(n9023) );
  NAND2_X1 U9273 ( .A1(n9018), .A2(n9020), .ZN(n9227) );
  NAND2_X1 U9274 ( .A1(n9228), .A2(n9229), .ZN(n9020) );
  NAND2_X1 U9275 ( .A1(b_25_), .A2(a_26_), .ZN(n9229) );
  INV_X1 U9276 ( .A(n9230), .ZN(n9228) );
  XNOR2_X1 U9277 ( .A(n9231), .B(n9232), .ZN(n9018) );
  NAND2_X1 U9278 ( .A1(n9233), .A2(n9234), .ZN(n9231) );
  NAND2_X1 U9279 ( .A1(a_26_), .A2(n9230), .ZN(n9019) );
  NAND2_X1 U9280 ( .A1(n9015), .A2(n9235), .ZN(n9230) );
  NAND2_X1 U9281 ( .A1(n9014), .A2(n9016), .ZN(n9235) );
  NAND2_X1 U9282 ( .A1(n9236), .A2(n9237), .ZN(n9016) );
  NAND2_X1 U9283 ( .A1(b_25_), .A2(a_27_), .ZN(n9237) );
  INV_X1 U9284 ( .A(n9238), .ZN(n9236) );
  XNOR2_X1 U9285 ( .A(n9239), .B(n9240), .ZN(n9014) );
  XOR2_X1 U9286 ( .A(n9241), .B(n9242), .Z(n9240) );
  NAND2_X1 U9287 ( .A1(b_24_), .A2(a_28_), .ZN(n9242) );
  NAND2_X1 U9288 ( .A1(a_27_), .A2(n9238), .ZN(n9015) );
  NAND2_X1 U9289 ( .A1(n9243), .A2(n9244), .ZN(n9238) );
  NAND2_X1 U9290 ( .A1(n9245), .A2(b_25_), .ZN(n9244) );
  NOR2_X1 U9291 ( .A1(n9246), .A2(n7803), .ZN(n9245) );
  NOR2_X1 U9292 ( .A1(n8990), .A2(n8992), .ZN(n9246) );
  NAND2_X1 U9293 ( .A1(n8990), .A2(n8992), .ZN(n9243) );
  NAND2_X1 U9294 ( .A1(n9247), .A2(n9248), .ZN(n8992) );
  NAND2_X1 U9295 ( .A1(n9010), .A2(n9249), .ZN(n9248) );
  NAND2_X1 U9296 ( .A1(n9012), .A2(n9011), .ZN(n9249) );
  NOR2_X1 U9297 ( .A1(n8775), .A2(n7337), .ZN(n9010) );
  OR2_X1 U9298 ( .A1(n9011), .A2(n9012), .ZN(n9247) );
  AND2_X1 U9299 ( .A1(n9250), .A2(n9251), .ZN(n9012) );
  NAND2_X1 U9300 ( .A1(n9252), .A2(b_23_), .ZN(n9251) );
  NOR2_X1 U9301 ( .A1(n9253), .A2(n7817), .ZN(n9252) );
  NOR2_X1 U9302 ( .A1(n7816), .A2(n9007), .ZN(n9253) );
  NAND2_X1 U9303 ( .A1(n9254), .A2(b_24_), .ZN(n9250) );
  NOR2_X1 U9304 ( .A1(n9255), .A2(n8052), .ZN(n9254) );
  NOR2_X1 U9305 ( .A1(n7810), .A2(n9256), .ZN(n9255) );
  NAND2_X1 U9306 ( .A1(n9257), .A2(b_25_), .ZN(n9011) );
  NOR2_X1 U9307 ( .A1(n8055), .A2(n9007), .ZN(n9257) );
  XOR2_X1 U9308 ( .A(n9258), .B(n9259), .Z(n8990) );
  XOR2_X1 U9309 ( .A(n9260), .B(n9261), .Z(n9258) );
  XNOR2_X1 U9310 ( .A(n9262), .B(n9263), .ZN(n9022) );
  NAND2_X1 U9311 ( .A1(n9264), .A2(n9265), .ZN(n9262) );
  XOR2_X1 U9312 ( .A(n9266), .B(n9267), .Z(n9026) );
  XOR2_X1 U9313 ( .A(n9268), .B(n9269), .Z(n9266) );
  XNOR2_X1 U9314 ( .A(n9270), .B(n9271), .ZN(n9030) );
  XNOR2_X1 U9315 ( .A(n9272), .B(n9273), .ZN(n9270) );
  XNOR2_X1 U9316 ( .A(n9274), .B(n9275), .ZN(n9033) );
  XNOR2_X1 U9317 ( .A(n9276), .B(n9277), .ZN(n9275) );
  XNOR2_X1 U9318 ( .A(n9278), .B(n9279), .ZN(n9037) );
  XOR2_X1 U9319 ( .A(n9280), .B(n9281), .Z(n9279) );
  NAND2_X1 U9320 ( .A1(b_24_), .A2(a_22_), .ZN(n9281) );
  XOR2_X1 U9321 ( .A(n9282), .B(n9283), .Z(n9041) );
  XOR2_X1 U9322 ( .A(n9284), .B(n9285), .Z(n9282) );
  XOR2_X1 U9323 ( .A(n9286), .B(n9287), .Z(n9045) );
  XOR2_X1 U9324 ( .A(n9288), .B(n9289), .Z(n9286) );
  NOR2_X1 U9325 ( .A1(n7755), .A2(n9007), .ZN(n9289) );
  XOR2_X1 U9326 ( .A(n9290), .B(n9291), .Z(n9050) );
  XOR2_X1 U9327 ( .A(n9292), .B(n9293), .Z(n9290) );
  XOR2_X1 U9328 ( .A(n9294), .B(n9295), .Z(n9053) );
  XOR2_X1 U9329 ( .A(n9296), .B(n9297), .Z(n9294) );
  NOR2_X1 U9330 ( .A1(n7745), .A2(n9007), .ZN(n9297) );
  XOR2_X1 U9331 ( .A(n9298), .B(n9299), .Z(n9058) );
  XOR2_X1 U9332 ( .A(n9300), .B(n9301), .Z(n9298) );
  XOR2_X1 U9333 ( .A(n9302), .B(n9303), .Z(n9062) );
  XOR2_X1 U9334 ( .A(n9304), .B(n9305), .Z(n9303) );
  NAND2_X1 U9335 ( .A1(b_24_), .A2(a_16_), .ZN(n9305) );
  XOR2_X1 U9336 ( .A(n9306), .B(n9307), .Z(n9065) );
  XOR2_X1 U9337 ( .A(n9308), .B(n9309), .Z(n9306) );
  XOR2_X1 U9338 ( .A(n9310), .B(n9311), .Z(n9070) );
  XOR2_X1 U9339 ( .A(n9312), .B(n9313), .Z(n9310) );
  NOR2_X1 U9340 ( .A1(n7727), .A2(n9007), .ZN(n9313) );
  XNOR2_X1 U9341 ( .A(n9314), .B(n9315), .ZN(n9074) );
  XNOR2_X1 U9342 ( .A(n9316), .B(n9317), .ZN(n9314) );
  XOR2_X1 U9343 ( .A(n9318), .B(n9319), .Z(n9078) );
  XOR2_X1 U9344 ( .A(n9320), .B(n9321), .Z(n9318) );
  NOR2_X1 U9345 ( .A1(n7718), .A2(n9007), .ZN(n9321) );
  XOR2_X1 U9346 ( .A(n9322), .B(n9323), .Z(n9082) );
  XOR2_X1 U9347 ( .A(n9324), .B(n9325), .Z(n9322) );
  NOR2_X1 U9348 ( .A1(n7424), .A2(n9007), .ZN(n9325) );
  XOR2_X1 U9349 ( .A(n9326), .B(n9327), .Z(n9086) );
  XOR2_X1 U9350 ( .A(n9328), .B(n9329), .Z(n9326) );
  NOR2_X1 U9351 ( .A1(n7709), .A2(n9007), .ZN(n9329) );
  XOR2_X1 U9352 ( .A(n9330), .B(n9331), .Z(n8916) );
  XOR2_X1 U9353 ( .A(n9332), .B(n9333), .Z(n9330) );
  OR2_X1 U9354 ( .A1(n9096), .A2(n9094), .ZN(n9152) );
  XOR2_X1 U9355 ( .A(n9334), .B(n9335), .Z(n9094) );
  NAND2_X1 U9356 ( .A1(n9336), .A2(n9337), .ZN(n9334) );
  NAND2_X1 U9357 ( .A1(b_25_), .A2(a_6_), .ZN(n9096) );
  XNOR2_X1 U9358 ( .A(n9338), .B(n9339), .ZN(n9098) );
  XNOR2_X1 U9359 ( .A(n9340), .B(n9341), .ZN(n9338) );
  XNOR2_X1 U9360 ( .A(n9342), .B(n9343), .ZN(n9102) );
  XNOR2_X1 U9361 ( .A(n9344), .B(n9345), .ZN(n9343) );
  XOR2_X1 U9362 ( .A(n9346), .B(n9347), .Z(n8894) );
  XOR2_X1 U9363 ( .A(n9348), .B(n9349), .Z(n9346) );
  NOR2_X1 U9364 ( .A1(n7682), .A2(n9007), .ZN(n9349) );
  XNOR2_X1 U9365 ( .A(n9350), .B(n9351), .ZN(n9110) );
  NAND2_X1 U9366 ( .A1(n9352), .A2(n9353), .ZN(n9350) );
  XNOR2_X1 U9367 ( .A(n9354), .B(n9355), .ZN(n9114) );
  XOR2_X1 U9368 ( .A(n9356), .B(n9357), .Z(n9354) );
  XOR2_X1 U9369 ( .A(n9358), .B(n9119), .Z(n9124) );
  XNOR2_X1 U9370 ( .A(n9359), .B(n9360), .ZN(n9119) );
  NOR2_X1 U9371 ( .A1(n7478), .A2(n9007), .ZN(n9360) );
  INV_X1 U9372 ( .A(n9120), .ZN(n9358) );
  NAND2_X1 U9373 ( .A1(n9361), .A2(n9362), .ZN(n7515) );
  XOR2_X1 U9374 ( .A(n7627), .B(n7626), .Z(n9362) );
  INV_X1 U9375 ( .A(n7635), .ZN(n7626) );
  AND2_X1 U9376 ( .A1(n7634), .A2(n7633), .ZN(n9361) );
  XOR2_X1 U9377 ( .A(n9363), .B(n9364), .Z(n7633) );
  XOR2_X1 U9378 ( .A(n9365), .B(n9366), .Z(n9363) );
  NOR2_X1 U9379 ( .A1(n7478), .A2(n9256), .ZN(n9366) );
  NAND2_X1 U9380 ( .A1(n9367), .A2(n9368), .ZN(n7634) );
  NAND2_X1 U9381 ( .A1(n9369), .A2(b_24_), .ZN(n9368) );
  NOR2_X1 U9382 ( .A1(n9370), .A2(n7478), .ZN(n9369) );
  NOR2_X1 U9383 ( .A1(n9120), .A2(n9359), .ZN(n9370) );
  NAND2_X1 U9384 ( .A1(n9120), .A2(n9359), .ZN(n9367) );
  NAND2_X1 U9385 ( .A1(n9371), .A2(n9372), .ZN(n9359) );
  NAND2_X1 U9386 ( .A1(n9356), .A2(n9373), .ZN(n9372) );
  OR2_X1 U9387 ( .A1(n9355), .A2(n9357), .ZN(n9373) );
  NAND2_X1 U9388 ( .A1(n9352), .A2(n9374), .ZN(n9356) );
  NAND2_X1 U9389 ( .A1(n9351), .A2(n9353), .ZN(n9374) );
  NAND2_X1 U9390 ( .A1(n9375), .A2(n9376), .ZN(n9353) );
  NAND2_X1 U9391 ( .A1(b_24_), .A2(a_2_), .ZN(n9376) );
  INV_X1 U9392 ( .A(n9377), .ZN(n9375) );
  XNOR2_X1 U9393 ( .A(n9378), .B(n9379), .ZN(n9351) );
  XOR2_X1 U9394 ( .A(n9380), .B(n9381), .Z(n9379) );
  NAND2_X1 U9395 ( .A1(b_23_), .A2(a_3_), .ZN(n9381) );
  NAND2_X1 U9396 ( .A1(a_2_), .A2(n9377), .ZN(n9352) );
  NAND2_X1 U9397 ( .A1(n9138), .A2(n9382), .ZN(n9377) );
  NAND2_X1 U9398 ( .A1(n9137), .A2(n9139), .ZN(n9382) );
  NAND2_X1 U9399 ( .A1(n9383), .A2(n9384), .ZN(n9139) );
  NAND2_X1 U9400 ( .A1(b_24_), .A2(a_3_), .ZN(n9384) );
  INV_X1 U9401 ( .A(n9385), .ZN(n9383) );
  XNOR2_X1 U9402 ( .A(n9386), .B(n9387), .ZN(n9137) );
  XOR2_X1 U9403 ( .A(n9388), .B(n9389), .Z(n9387) );
  NAND2_X1 U9404 ( .A1(b_23_), .A2(a_4_), .ZN(n9389) );
  NAND2_X1 U9405 ( .A1(a_3_), .A2(n9385), .ZN(n9138) );
  NAND2_X1 U9406 ( .A1(n9390), .A2(n9391), .ZN(n9385) );
  NAND2_X1 U9407 ( .A1(n9392), .A2(b_24_), .ZN(n9391) );
  NOR2_X1 U9408 ( .A1(n9393), .A2(n7682), .ZN(n9392) );
  NOR2_X1 U9409 ( .A1(n9347), .A2(n9348), .ZN(n9393) );
  NAND2_X1 U9410 ( .A1(n9347), .A2(n9348), .ZN(n9390) );
  NAND2_X1 U9411 ( .A1(n9394), .A2(n9395), .ZN(n9348) );
  NAND2_X1 U9412 ( .A1(n9345), .A2(n9396), .ZN(n9395) );
  OR2_X1 U9413 ( .A1(n9344), .A2(n9342), .ZN(n9396) );
  NOR2_X1 U9414 ( .A1(n9007), .A2(n7455), .ZN(n9345) );
  NAND2_X1 U9415 ( .A1(n9342), .A2(n9344), .ZN(n9394) );
  NAND2_X1 U9416 ( .A1(n9397), .A2(n9398), .ZN(n9344) );
  NAND2_X1 U9417 ( .A1(n9340), .A2(n9399), .ZN(n9398) );
  NAND2_X1 U9418 ( .A1(n9339), .A2(n9341), .ZN(n9399) );
  NAND2_X1 U9419 ( .A1(n9336), .A2(n9400), .ZN(n9340) );
  NAND2_X1 U9420 ( .A1(n9335), .A2(n9337), .ZN(n9400) );
  NAND2_X1 U9421 ( .A1(n9401), .A2(n9402), .ZN(n9337) );
  NAND2_X1 U9422 ( .A1(b_24_), .A2(a_7_), .ZN(n9402) );
  INV_X1 U9423 ( .A(n9403), .ZN(n9401) );
  XOR2_X1 U9424 ( .A(n9404), .B(n9405), .Z(n9335) );
  XOR2_X1 U9425 ( .A(n9406), .B(n9407), .Z(n9404) );
  NAND2_X1 U9426 ( .A1(a_7_), .A2(n9403), .ZN(n9336) );
  NAND2_X1 U9427 ( .A1(n9408), .A2(n9409), .ZN(n9403) );
  NAND2_X1 U9428 ( .A1(n9410), .A2(b_24_), .ZN(n9409) );
  NOR2_X1 U9429 ( .A1(n9411), .A2(n7699), .ZN(n9410) );
  NOR2_X1 U9430 ( .A1(n9159), .A2(n9161), .ZN(n9411) );
  NAND2_X1 U9431 ( .A1(n9159), .A2(n9161), .ZN(n9408) );
  NAND2_X1 U9432 ( .A1(n9412), .A2(n9413), .ZN(n9161) );
  NAND2_X1 U9433 ( .A1(n9333), .A2(n9414), .ZN(n9413) );
  OR2_X1 U9434 ( .A1(n9332), .A2(n9331), .ZN(n9414) );
  NOR2_X1 U9435 ( .A1(n9007), .A2(n7704), .ZN(n9333) );
  NAND2_X1 U9436 ( .A1(n9331), .A2(n9332), .ZN(n9412) );
  NAND2_X1 U9437 ( .A1(n9415), .A2(n9416), .ZN(n9332) );
  NAND2_X1 U9438 ( .A1(n9417), .A2(b_24_), .ZN(n9416) );
  NOR2_X1 U9439 ( .A1(n9418), .A2(n7709), .ZN(n9417) );
  NOR2_X1 U9440 ( .A1(n9327), .A2(n9328), .ZN(n9418) );
  NAND2_X1 U9441 ( .A1(n9327), .A2(n9328), .ZN(n9415) );
  NAND2_X1 U9442 ( .A1(n9419), .A2(n9420), .ZN(n9328) );
  NAND2_X1 U9443 ( .A1(n9421), .A2(b_24_), .ZN(n9420) );
  NOR2_X1 U9444 ( .A1(n9422), .A2(n7424), .ZN(n9421) );
  NOR2_X1 U9445 ( .A1(n9323), .A2(n9324), .ZN(n9422) );
  NAND2_X1 U9446 ( .A1(n9323), .A2(n9324), .ZN(n9419) );
  NAND2_X1 U9447 ( .A1(n9423), .A2(n9424), .ZN(n9324) );
  NAND2_X1 U9448 ( .A1(n9425), .A2(b_24_), .ZN(n9424) );
  NOR2_X1 U9449 ( .A1(n9426), .A2(n7718), .ZN(n9425) );
  NOR2_X1 U9450 ( .A1(n9319), .A2(n9320), .ZN(n9426) );
  NAND2_X1 U9451 ( .A1(n9319), .A2(n9320), .ZN(n9423) );
  NAND2_X1 U9452 ( .A1(n9427), .A2(n9428), .ZN(n9320) );
  NAND2_X1 U9453 ( .A1(n9317), .A2(n9429), .ZN(n9428) );
  NAND2_X1 U9454 ( .A1(n9316), .A2(n9315), .ZN(n9429) );
  NOR2_X1 U9455 ( .A1(n9007), .A2(n7415), .ZN(n9317) );
  OR2_X1 U9456 ( .A1(n9315), .A2(n9316), .ZN(n9427) );
  AND2_X1 U9457 ( .A1(n9430), .A2(n9431), .ZN(n9316) );
  NAND2_X1 U9458 ( .A1(n9432), .A2(b_24_), .ZN(n9431) );
  NOR2_X1 U9459 ( .A1(n9433), .A2(n7727), .ZN(n9432) );
  NOR2_X1 U9460 ( .A1(n9311), .A2(n9312), .ZN(n9433) );
  NAND2_X1 U9461 ( .A1(n9311), .A2(n9312), .ZN(n9430) );
  NAND2_X1 U9462 ( .A1(n9434), .A2(n9435), .ZN(n9312) );
  NAND2_X1 U9463 ( .A1(n9309), .A2(n9436), .ZN(n9435) );
  OR2_X1 U9464 ( .A1(n9308), .A2(n9307), .ZN(n9436) );
  NOR2_X1 U9465 ( .A1(n9007), .A2(n7406), .ZN(n9309) );
  NAND2_X1 U9466 ( .A1(n9307), .A2(n9308), .ZN(n9434) );
  NAND2_X1 U9467 ( .A1(n9437), .A2(n9438), .ZN(n9308) );
  NAND2_X1 U9468 ( .A1(n9439), .A2(b_24_), .ZN(n9438) );
  NOR2_X1 U9469 ( .A1(n9440), .A2(n7736), .ZN(n9439) );
  NOR2_X1 U9470 ( .A1(n9302), .A2(n9304), .ZN(n9440) );
  NAND2_X1 U9471 ( .A1(n9302), .A2(n9304), .ZN(n9437) );
  NAND2_X1 U9472 ( .A1(n9441), .A2(n9442), .ZN(n9304) );
  NAND2_X1 U9473 ( .A1(n9301), .A2(n9443), .ZN(n9442) );
  OR2_X1 U9474 ( .A1(n9300), .A2(n9299), .ZN(n9443) );
  NOR2_X1 U9475 ( .A1(n9007), .A2(n7397), .ZN(n9301) );
  NAND2_X1 U9476 ( .A1(n9299), .A2(n9300), .ZN(n9441) );
  NAND2_X1 U9477 ( .A1(n9444), .A2(n9445), .ZN(n9300) );
  NAND2_X1 U9478 ( .A1(n9446), .A2(b_24_), .ZN(n9445) );
  NOR2_X1 U9479 ( .A1(n9447), .A2(n7745), .ZN(n9446) );
  NOR2_X1 U9480 ( .A1(n9295), .A2(n9296), .ZN(n9447) );
  NAND2_X1 U9481 ( .A1(n9295), .A2(n9296), .ZN(n9444) );
  NAND2_X1 U9482 ( .A1(n9448), .A2(n9449), .ZN(n9296) );
  NAND2_X1 U9483 ( .A1(n9293), .A2(n9450), .ZN(n9449) );
  OR2_X1 U9484 ( .A1(n9292), .A2(n9291), .ZN(n9450) );
  NOR2_X1 U9485 ( .A1(n9007), .A2(n7750), .ZN(n9293) );
  NAND2_X1 U9486 ( .A1(n9291), .A2(n9292), .ZN(n9448) );
  NAND2_X1 U9487 ( .A1(n9451), .A2(n9452), .ZN(n9292) );
  NAND2_X1 U9488 ( .A1(n9453), .A2(b_24_), .ZN(n9452) );
  NOR2_X1 U9489 ( .A1(n9454), .A2(n7755), .ZN(n9453) );
  NOR2_X1 U9490 ( .A1(n9287), .A2(n9288), .ZN(n9454) );
  NAND2_X1 U9491 ( .A1(n9287), .A2(n9288), .ZN(n9451) );
  NAND2_X1 U9492 ( .A1(n9455), .A2(n9456), .ZN(n9288) );
  NAND2_X1 U9493 ( .A1(n9285), .A2(n9457), .ZN(n9456) );
  OR2_X1 U9494 ( .A1(n9284), .A2(n9283), .ZN(n9457) );
  NOR2_X1 U9495 ( .A1(n9007), .A2(n7760), .ZN(n9285) );
  NAND2_X1 U9496 ( .A1(n9283), .A2(n9284), .ZN(n9455) );
  NAND2_X1 U9497 ( .A1(n9458), .A2(n9459), .ZN(n9284) );
  NAND2_X1 U9498 ( .A1(n9460), .A2(b_24_), .ZN(n9459) );
  NOR2_X1 U9499 ( .A1(n9461), .A2(n7765), .ZN(n9460) );
  NOR2_X1 U9500 ( .A1(n9278), .A2(n9280), .ZN(n9461) );
  NAND2_X1 U9501 ( .A1(n9278), .A2(n9280), .ZN(n9458) );
  NAND2_X1 U9502 ( .A1(n9462), .A2(n9463), .ZN(n9280) );
  NAND2_X1 U9503 ( .A1(n9277), .A2(n9464), .ZN(n9463) );
  OR2_X1 U9504 ( .A1(n9276), .A2(n9274), .ZN(n9464) );
  NOR2_X1 U9505 ( .A1(n9007), .A2(n8014), .ZN(n9277) );
  NAND2_X1 U9506 ( .A1(n9274), .A2(n9276), .ZN(n9462) );
  NAND2_X1 U9507 ( .A1(n9465), .A2(n9466), .ZN(n9276) );
  NAND2_X1 U9508 ( .A1(n9272), .A2(n9467), .ZN(n9466) );
  NAND2_X1 U9509 ( .A1(n9273), .A2(n9271), .ZN(n9467) );
  OR2_X1 U9510 ( .A1(n9271), .A2(n9273), .ZN(n9465) );
  AND2_X1 U9511 ( .A1(n9468), .A2(n9469), .ZN(n9273) );
  NAND2_X1 U9512 ( .A1(n9269), .A2(n9470), .ZN(n9469) );
  OR2_X1 U9513 ( .A1(n9268), .A2(n9267), .ZN(n9470) );
  NOR2_X1 U9514 ( .A1(n9007), .A2(n8022), .ZN(n9269) );
  NAND2_X1 U9515 ( .A1(n9267), .A2(n9268), .ZN(n9468) );
  NAND2_X1 U9516 ( .A1(n9264), .A2(n9471), .ZN(n9268) );
  NAND2_X1 U9517 ( .A1(n9263), .A2(n9265), .ZN(n9471) );
  NAND2_X1 U9518 ( .A1(n9472), .A2(n9473), .ZN(n9265) );
  NAND2_X1 U9519 ( .A1(b_24_), .A2(a_26_), .ZN(n9473) );
  INV_X1 U9520 ( .A(n9474), .ZN(n9472) );
  XNOR2_X1 U9521 ( .A(n9475), .B(n9476), .ZN(n9263) );
  NAND2_X1 U9522 ( .A1(n9477), .A2(n9478), .ZN(n9475) );
  NAND2_X1 U9523 ( .A1(a_26_), .A2(n9474), .ZN(n9264) );
  NAND2_X1 U9524 ( .A1(n9233), .A2(n9479), .ZN(n9474) );
  NAND2_X1 U9525 ( .A1(n9232), .A2(n9234), .ZN(n9479) );
  NAND2_X1 U9526 ( .A1(n9480), .A2(n9481), .ZN(n9234) );
  NAND2_X1 U9527 ( .A1(b_24_), .A2(a_27_), .ZN(n9481) );
  INV_X1 U9528 ( .A(n9482), .ZN(n9480) );
  XNOR2_X1 U9529 ( .A(n9483), .B(n9484), .ZN(n9232) );
  XOR2_X1 U9530 ( .A(n9485), .B(n9486), .Z(n9484) );
  NAND2_X1 U9531 ( .A1(b_23_), .A2(a_28_), .ZN(n9486) );
  NAND2_X1 U9532 ( .A1(a_27_), .A2(n9482), .ZN(n9233) );
  NAND2_X1 U9533 ( .A1(n9487), .A2(n9488), .ZN(n9482) );
  NAND2_X1 U9534 ( .A1(n9489), .A2(b_24_), .ZN(n9488) );
  NOR2_X1 U9535 ( .A1(n9490), .A2(n7803), .ZN(n9489) );
  NOR2_X1 U9536 ( .A1(n9239), .A2(n9241), .ZN(n9490) );
  NAND2_X1 U9537 ( .A1(n9239), .A2(n9241), .ZN(n9487) );
  NAND2_X1 U9538 ( .A1(n9491), .A2(n9492), .ZN(n9241) );
  NAND2_X1 U9539 ( .A1(n9259), .A2(n9493), .ZN(n9492) );
  NAND2_X1 U9540 ( .A1(n9261), .A2(n9260), .ZN(n9493) );
  NOR2_X1 U9541 ( .A1(n9007), .A2(n7337), .ZN(n9259) );
  OR2_X1 U9542 ( .A1(n9260), .A2(n9261), .ZN(n9491) );
  AND2_X1 U9543 ( .A1(n9494), .A2(n9495), .ZN(n9261) );
  NAND2_X1 U9544 ( .A1(n9496), .A2(b_22_), .ZN(n9495) );
  NOR2_X1 U9545 ( .A1(n9497), .A2(n7817), .ZN(n9496) );
  NOR2_X1 U9546 ( .A1(n7816), .A2(n9256), .ZN(n9497) );
  NAND2_X1 U9547 ( .A1(n9498), .A2(b_23_), .ZN(n9494) );
  NOR2_X1 U9548 ( .A1(n9499), .A2(n8052), .ZN(n9498) );
  NOR2_X1 U9549 ( .A1(n7810), .A2(n9500), .ZN(n9499) );
  NAND2_X1 U9550 ( .A1(n9501), .A2(b_24_), .ZN(n9260) );
  XOR2_X1 U9551 ( .A(n9502), .B(n9503), .Z(n9239) );
  XOR2_X1 U9552 ( .A(n9504), .B(n9505), .Z(n9502) );
  XNOR2_X1 U9553 ( .A(n9506), .B(n9507), .ZN(n9267) );
  NAND2_X1 U9554 ( .A1(n9508), .A2(n9509), .ZN(n9506) );
  XNOR2_X1 U9555 ( .A(n9510), .B(n9511), .ZN(n9271) );
  XOR2_X1 U9556 ( .A(n9512), .B(n9513), .Z(n9510) );
  XOR2_X1 U9557 ( .A(n9514), .B(n9515), .Z(n9274) );
  XNOR2_X1 U9558 ( .A(n9516), .B(n9517), .ZN(n9514) );
  NAND2_X1 U9559 ( .A1(b_23_), .A2(a_24_), .ZN(n9516) );
  XOR2_X1 U9560 ( .A(n9518), .B(n9519), .Z(n9278) );
  XOR2_X1 U9561 ( .A(n9520), .B(n9521), .Z(n9518) );
  XNOR2_X1 U9562 ( .A(n9522), .B(n9523), .ZN(n9283) );
  XOR2_X1 U9563 ( .A(n9524), .B(n9525), .Z(n9523) );
  NAND2_X1 U9564 ( .A1(b_23_), .A2(a_22_), .ZN(n9525) );
  XOR2_X1 U9565 ( .A(n9526), .B(n9527), .Z(n9287) );
  XOR2_X1 U9566 ( .A(n9528), .B(n9529), .Z(n9526) );
  XOR2_X1 U9567 ( .A(n9530), .B(n9531), .Z(n9291) );
  XOR2_X1 U9568 ( .A(n9532), .B(n9533), .Z(n9530) );
  NOR2_X1 U9569 ( .A1(n7755), .A2(n9256), .ZN(n9533) );
  XNOR2_X1 U9570 ( .A(n9534), .B(n9535), .ZN(n9295) );
  XNOR2_X1 U9571 ( .A(n9536), .B(n9537), .ZN(n9535) );
  XNOR2_X1 U9572 ( .A(n9538), .B(n9539), .ZN(n9299) );
  XOR2_X1 U9573 ( .A(n9540), .B(n9541), .Z(n9539) );
  NAND2_X1 U9574 ( .A1(b_23_), .A2(a_18_), .ZN(n9541) );
  XNOR2_X1 U9575 ( .A(n9542), .B(n9543), .ZN(n9302) );
  XNOR2_X1 U9576 ( .A(n9544), .B(n9545), .ZN(n9543) );
  XOR2_X1 U9577 ( .A(n9546), .B(n9547), .Z(n9307) );
  XOR2_X1 U9578 ( .A(n9548), .B(n9549), .Z(n9546) );
  NOR2_X1 U9579 ( .A1(n7736), .A2(n9256), .ZN(n9549) );
  XOR2_X1 U9580 ( .A(n9550), .B(n9551), .Z(n9311) );
  XOR2_X1 U9581 ( .A(n9552), .B(n9553), .Z(n9550) );
  NOR2_X1 U9582 ( .A1(n7406), .A2(n9256), .ZN(n9553) );
  XOR2_X1 U9583 ( .A(n9554), .B(n9555), .Z(n9315) );
  NAND2_X1 U9584 ( .A1(n9556), .A2(n9557), .ZN(n9554) );
  XOR2_X1 U9585 ( .A(n9558), .B(n9559), .Z(n9319) );
  XOR2_X1 U9586 ( .A(n9560), .B(n9561), .Z(n9558) );
  XOR2_X1 U9587 ( .A(n9562), .B(n9563), .Z(n9323) );
  XOR2_X1 U9588 ( .A(n9564), .B(n9565), .Z(n9562) );
  NOR2_X1 U9589 ( .A1(n7718), .A2(n9256), .ZN(n9565) );
  XOR2_X1 U9590 ( .A(n9566), .B(n9567), .Z(n9327) );
  XOR2_X1 U9591 ( .A(n9568), .B(n9569), .Z(n9566) );
  NOR2_X1 U9592 ( .A1(n7424), .A2(n9256), .ZN(n9569) );
  XNOR2_X1 U9593 ( .A(n9570), .B(n9571), .ZN(n9331) );
  XOR2_X1 U9594 ( .A(n9572), .B(n9573), .Z(n9571) );
  NAND2_X1 U9595 ( .A1(b_23_), .A2(a_10_), .ZN(n9573) );
  XOR2_X1 U9596 ( .A(n9574), .B(n9575), .Z(n9159) );
  XOR2_X1 U9597 ( .A(n9576), .B(n9577), .Z(n9574) );
  OR2_X1 U9598 ( .A1(n9341), .A2(n9339), .ZN(n9397) );
  XNOR2_X1 U9599 ( .A(n9578), .B(n9579), .ZN(n9339) );
  XOR2_X1 U9600 ( .A(n9580), .B(n9581), .Z(n9578) );
  NOR2_X1 U9601 ( .A1(n7445), .A2(n9256), .ZN(n9581) );
  NAND2_X1 U9602 ( .A1(b_24_), .A2(a_6_), .ZN(n9341) );
  XNOR2_X1 U9603 ( .A(n9582), .B(n9583), .ZN(n9342) );
  NAND2_X1 U9604 ( .A1(n9584), .A2(n9585), .ZN(n9582) );
  XOR2_X1 U9605 ( .A(n9586), .B(n9587), .Z(n9347) );
  XOR2_X1 U9606 ( .A(n9588), .B(n9589), .Z(n9586) );
  NOR2_X1 U9607 ( .A1(n7455), .A2(n9256), .ZN(n9589) );
  NAND2_X1 U9608 ( .A1(n9357), .A2(n9355), .ZN(n9371) );
  XNOR2_X1 U9609 ( .A(n9590), .B(n9591), .ZN(n9355) );
  XOR2_X1 U9610 ( .A(n9592), .B(n9593), .Z(n9591) );
  NAND2_X1 U9611 ( .A1(b_23_), .A2(a_2_), .ZN(n9593) );
  NOR2_X1 U9612 ( .A1(n9007), .A2(n7669), .ZN(n9357) );
  XNOR2_X1 U9613 ( .A(n9594), .B(n9595), .ZN(n9120) );
  XOR2_X1 U9614 ( .A(n9596), .B(n9597), .Z(n9595) );
  NAND2_X1 U9615 ( .A1(b_23_), .A2(a_1_), .ZN(n9597) );
  NAND2_X1 U9616 ( .A1(n9598), .A2(n9599), .ZN(n7518) );
  AND2_X1 U9617 ( .A1(n9600), .A2(n7627), .ZN(n9599) );
  NAND2_X1 U9618 ( .A1(n9601), .A2(n9602), .ZN(n7627) );
  NAND2_X1 U9619 ( .A1(n9603), .A2(b_23_), .ZN(n9602) );
  NOR2_X1 U9620 ( .A1(n9604), .A2(n7478), .ZN(n9603) );
  NOR2_X1 U9621 ( .A1(n9364), .A2(n9365), .ZN(n9604) );
  NAND2_X1 U9622 ( .A1(n9364), .A2(n9365), .ZN(n9601) );
  NAND2_X1 U9623 ( .A1(n9605), .A2(n9606), .ZN(n9365) );
  NAND2_X1 U9624 ( .A1(n9607), .A2(b_23_), .ZN(n9606) );
  NOR2_X1 U9625 ( .A1(n9608), .A2(n7669), .ZN(n9607) );
  NOR2_X1 U9626 ( .A1(n9594), .A2(n9596), .ZN(n9608) );
  NAND2_X1 U9627 ( .A1(n9594), .A2(n9596), .ZN(n9605) );
  NAND2_X1 U9628 ( .A1(n9609), .A2(n9610), .ZN(n9596) );
  NAND2_X1 U9629 ( .A1(n9611), .A2(b_23_), .ZN(n9610) );
  NOR2_X1 U9630 ( .A1(n9612), .A2(n7469), .ZN(n9611) );
  NOR2_X1 U9631 ( .A1(n9590), .A2(n9592), .ZN(n9612) );
  NAND2_X1 U9632 ( .A1(n9590), .A2(n9592), .ZN(n9609) );
  NAND2_X1 U9633 ( .A1(n9613), .A2(n9614), .ZN(n9592) );
  NAND2_X1 U9634 ( .A1(n9615), .A2(b_23_), .ZN(n9614) );
  NOR2_X1 U9635 ( .A1(n9616), .A2(n7464), .ZN(n9615) );
  NOR2_X1 U9636 ( .A1(n9378), .A2(n9380), .ZN(n9616) );
  NAND2_X1 U9637 ( .A1(n9378), .A2(n9380), .ZN(n9613) );
  NAND2_X1 U9638 ( .A1(n9617), .A2(n9618), .ZN(n9380) );
  NAND2_X1 U9639 ( .A1(n9619), .A2(b_23_), .ZN(n9618) );
  NOR2_X1 U9640 ( .A1(n9620), .A2(n7682), .ZN(n9619) );
  NOR2_X1 U9641 ( .A1(n9386), .A2(n9388), .ZN(n9620) );
  NAND2_X1 U9642 ( .A1(n9386), .A2(n9388), .ZN(n9617) );
  NAND2_X1 U9643 ( .A1(n9621), .A2(n9622), .ZN(n9388) );
  NAND2_X1 U9644 ( .A1(n9623), .A2(b_23_), .ZN(n9622) );
  NOR2_X1 U9645 ( .A1(n9624), .A2(n7455), .ZN(n9623) );
  NOR2_X1 U9646 ( .A1(n9587), .A2(n9588), .ZN(n9624) );
  NAND2_X1 U9647 ( .A1(n9587), .A2(n9588), .ZN(n9621) );
  NAND2_X1 U9648 ( .A1(n9584), .A2(n9625), .ZN(n9588) );
  NAND2_X1 U9649 ( .A1(n9583), .A2(n9585), .ZN(n9625) );
  NAND2_X1 U9650 ( .A1(n9626), .A2(n9627), .ZN(n9585) );
  NAND2_X1 U9651 ( .A1(b_23_), .A2(a_6_), .ZN(n9627) );
  INV_X1 U9652 ( .A(n9628), .ZN(n9626) );
  XNOR2_X1 U9653 ( .A(n9629), .B(n9630), .ZN(n9583) );
  XNOR2_X1 U9654 ( .A(n9631), .B(n9632), .ZN(n9630) );
  NAND2_X1 U9655 ( .A1(a_6_), .A2(n9628), .ZN(n9584) );
  NAND2_X1 U9656 ( .A1(n9633), .A2(n9634), .ZN(n9628) );
  NAND2_X1 U9657 ( .A1(n9635), .A2(b_23_), .ZN(n9634) );
  NOR2_X1 U9658 ( .A1(n9636), .A2(n7445), .ZN(n9635) );
  NOR2_X1 U9659 ( .A1(n9579), .A2(n9580), .ZN(n9636) );
  NAND2_X1 U9660 ( .A1(n9579), .A2(n9580), .ZN(n9633) );
  NAND2_X1 U9661 ( .A1(n9637), .A2(n9638), .ZN(n9580) );
  NAND2_X1 U9662 ( .A1(n9407), .A2(n9639), .ZN(n9638) );
  OR2_X1 U9663 ( .A1(n9406), .A2(n9405), .ZN(n9639) );
  NOR2_X1 U9664 ( .A1(n9256), .A2(n7699), .ZN(n9407) );
  NAND2_X1 U9665 ( .A1(n9405), .A2(n9406), .ZN(n9637) );
  NAND2_X1 U9666 ( .A1(n9640), .A2(n9641), .ZN(n9406) );
  NAND2_X1 U9667 ( .A1(n9577), .A2(n9642), .ZN(n9641) );
  OR2_X1 U9668 ( .A1(n9576), .A2(n9575), .ZN(n9642) );
  NOR2_X1 U9669 ( .A1(n9256), .A2(n7704), .ZN(n9577) );
  NAND2_X1 U9670 ( .A1(n9575), .A2(n9576), .ZN(n9640) );
  NAND2_X1 U9671 ( .A1(n9643), .A2(n9644), .ZN(n9576) );
  NAND2_X1 U9672 ( .A1(n9645), .A2(b_23_), .ZN(n9644) );
  NOR2_X1 U9673 ( .A1(n9646), .A2(n7709), .ZN(n9645) );
  NOR2_X1 U9674 ( .A1(n9570), .A2(n9572), .ZN(n9646) );
  NAND2_X1 U9675 ( .A1(n9570), .A2(n9572), .ZN(n9643) );
  NAND2_X1 U9676 ( .A1(n9647), .A2(n9648), .ZN(n9572) );
  NAND2_X1 U9677 ( .A1(n9649), .A2(b_23_), .ZN(n9648) );
  NOR2_X1 U9678 ( .A1(n9650), .A2(n7424), .ZN(n9649) );
  NOR2_X1 U9679 ( .A1(n9567), .A2(n9568), .ZN(n9650) );
  NAND2_X1 U9680 ( .A1(n9567), .A2(n9568), .ZN(n9647) );
  NAND2_X1 U9681 ( .A1(n9651), .A2(n9652), .ZN(n9568) );
  NAND2_X1 U9682 ( .A1(n9653), .A2(b_23_), .ZN(n9652) );
  NOR2_X1 U9683 ( .A1(n9654), .A2(n7718), .ZN(n9653) );
  NOR2_X1 U9684 ( .A1(n9563), .A2(n9564), .ZN(n9654) );
  NAND2_X1 U9685 ( .A1(n9563), .A2(n9564), .ZN(n9651) );
  NAND2_X1 U9686 ( .A1(n9655), .A2(n9656), .ZN(n9564) );
  NAND2_X1 U9687 ( .A1(n9561), .A2(n9657), .ZN(n9656) );
  OR2_X1 U9688 ( .A1(n9560), .A2(n9559), .ZN(n9657) );
  NOR2_X1 U9689 ( .A1(n9256), .A2(n7415), .ZN(n9561) );
  NAND2_X1 U9690 ( .A1(n9559), .A2(n9560), .ZN(n9655) );
  NAND2_X1 U9691 ( .A1(n9556), .A2(n9658), .ZN(n9560) );
  NAND2_X1 U9692 ( .A1(n9555), .A2(n9557), .ZN(n9658) );
  NAND2_X1 U9693 ( .A1(n9659), .A2(n9660), .ZN(n9557) );
  NAND2_X1 U9694 ( .A1(b_23_), .A2(a_14_), .ZN(n9660) );
  INV_X1 U9695 ( .A(n9661), .ZN(n9659) );
  XOR2_X1 U9696 ( .A(n9662), .B(n9663), .Z(n9555) );
  XOR2_X1 U9697 ( .A(n9664), .B(n9665), .Z(n9662) );
  NAND2_X1 U9698 ( .A1(a_14_), .A2(n9661), .ZN(n9556) );
  NAND2_X1 U9699 ( .A1(n9666), .A2(n9667), .ZN(n9661) );
  NAND2_X1 U9700 ( .A1(n9668), .A2(b_23_), .ZN(n9667) );
  NOR2_X1 U9701 ( .A1(n9669), .A2(n7406), .ZN(n9668) );
  NOR2_X1 U9702 ( .A1(n9551), .A2(n9552), .ZN(n9669) );
  NAND2_X1 U9703 ( .A1(n9551), .A2(n9552), .ZN(n9666) );
  NAND2_X1 U9704 ( .A1(n9670), .A2(n9671), .ZN(n9552) );
  NAND2_X1 U9705 ( .A1(n9672), .A2(b_23_), .ZN(n9671) );
  NOR2_X1 U9706 ( .A1(n9673), .A2(n7736), .ZN(n9672) );
  NOR2_X1 U9707 ( .A1(n9547), .A2(n9548), .ZN(n9673) );
  NAND2_X1 U9708 ( .A1(n9547), .A2(n9548), .ZN(n9670) );
  NAND2_X1 U9709 ( .A1(n9674), .A2(n9675), .ZN(n9548) );
  NAND2_X1 U9710 ( .A1(n9545), .A2(n9676), .ZN(n9675) );
  OR2_X1 U9711 ( .A1(n9544), .A2(n9542), .ZN(n9676) );
  NOR2_X1 U9712 ( .A1(n9256), .A2(n7397), .ZN(n9545) );
  NAND2_X1 U9713 ( .A1(n9542), .A2(n9544), .ZN(n9674) );
  NAND2_X1 U9714 ( .A1(n9677), .A2(n9678), .ZN(n9544) );
  NAND2_X1 U9715 ( .A1(n9679), .A2(b_23_), .ZN(n9678) );
  NOR2_X1 U9716 ( .A1(n9680), .A2(n7745), .ZN(n9679) );
  NOR2_X1 U9717 ( .A1(n9538), .A2(n9540), .ZN(n9680) );
  NAND2_X1 U9718 ( .A1(n9538), .A2(n9540), .ZN(n9677) );
  NAND2_X1 U9719 ( .A1(n9681), .A2(n9682), .ZN(n9540) );
  NAND2_X1 U9720 ( .A1(n9537), .A2(n9683), .ZN(n9682) );
  OR2_X1 U9721 ( .A1(n9536), .A2(n9534), .ZN(n9683) );
  NOR2_X1 U9722 ( .A1(n9256), .A2(n7750), .ZN(n9537) );
  NAND2_X1 U9723 ( .A1(n9534), .A2(n9536), .ZN(n9681) );
  NAND2_X1 U9724 ( .A1(n9684), .A2(n9685), .ZN(n9536) );
  NAND2_X1 U9725 ( .A1(n9686), .A2(b_23_), .ZN(n9685) );
  NOR2_X1 U9726 ( .A1(n9687), .A2(n7755), .ZN(n9686) );
  NOR2_X1 U9727 ( .A1(n9531), .A2(n9532), .ZN(n9687) );
  NAND2_X1 U9728 ( .A1(n9531), .A2(n9532), .ZN(n9684) );
  NAND2_X1 U9729 ( .A1(n9688), .A2(n9689), .ZN(n9532) );
  NAND2_X1 U9730 ( .A1(n9529), .A2(n9690), .ZN(n9689) );
  OR2_X1 U9731 ( .A1(n9528), .A2(n9527), .ZN(n9690) );
  NOR2_X1 U9732 ( .A1(n9256), .A2(n7760), .ZN(n9529) );
  NAND2_X1 U9733 ( .A1(n9527), .A2(n9528), .ZN(n9688) );
  NAND2_X1 U9734 ( .A1(n9691), .A2(n9692), .ZN(n9528) );
  NAND2_X1 U9735 ( .A1(n9693), .A2(b_23_), .ZN(n9692) );
  NOR2_X1 U9736 ( .A1(n9694), .A2(n7765), .ZN(n9693) );
  NOR2_X1 U9737 ( .A1(n9522), .A2(n9524), .ZN(n9694) );
  NAND2_X1 U9738 ( .A1(n9522), .A2(n9524), .ZN(n9691) );
  NAND2_X1 U9739 ( .A1(n9695), .A2(n9696), .ZN(n9524) );
  NAND2_X1 U9740 ( .A1(n9521), .A2(n9697), .ZN(n9696) );
  OR2_X1 U9741 ( .A1(n9520), .A2(n9519), .ZN(n9697) );
  NAND2_X1 U9742 ( .A1(n9519), .A2(n9520), .ZN(n9695) );
  NAND2_X1 U9743 ( .A1(n9698), .A2(n9699), .ZN(n9520) );
  NAND2_X1 U9744 ( .A1(n9700), .A2(b_23_), .ZN(n9699) );
  NOR2_X1 U9745 ( .A1(n9701), .A2(n7774), .ZN(n9700) );
  NOR2_X1 U9746 ( .A1(n9515), .A2(n9517), .ZN(n9701) );
  NAND2_X1 U9747 ( .A1(n9515), .A2(n9517), .ZN(n9698) );
  NAND2_X1 U9748 ( .A1(n9702), .A2(n9703), .ZN(n9517) );
  NAND2_X1 U9749 ( .A1(n9513), .A2(n9704), .ZN(n9703) );
  OR2_X1 U9750 ( .A1(n9512), .A2(n9511), .ZN(n9704) );
  NOR2_X1 U9751 ( .A1(n9256), .A2(n8022), .ZN(n9513) );
  NAND2_X1 U9752 ( .A1(n9511), .A2(n9512), .ZN(n9702) );
  NAND2_X1 U9753 ( .A1(n9508), .A2(n9705), .ZN(n9512) );
  NAND2_X1 U9754 ( .A1(n9507), .A2(n9509), .ZN(n9705) );
  NAND2_X1 U9755 ( .A1(n9706), .A2(n9707), .ZN(n9509) );
  NAND2_X1 U9756 ( .A1(b_23_), .A2(a_26_), .ZN(n9707) );
  INV_X1 U9757 ( .A(n9708), .ZN(n9706) );
  XNOR2_X1 U9758 ( .A(n9709), .B(n9710), .ZN(n9507) );
  NAND2_X1 U9759 ( .A1(n9711), .A2(n9712), .ZN(n9709) );
  NAND2_X1 U9760 ( .A1(a_26_), .A2(n9708), .ZN(n9508) );
  NAND2_X1 U9761 ( .A1(n9477), .A2(n9713), .ZN(n9708) );
  NAND2_X1 U9762 ( .A1(n9476), .A2(n9478), .ZN(n9713) );
  NAND2_X1 U9763 ( .A1(n9714), .A2(n9715), .ZN(n9478) );
  NAND2_X1 U9764 ( .A1(b_23_), .A2(a_27_), .ZN(n9715) );
  INV_X1 U9765 ( .A(n9716), .ZN(n9714) );
  XNOR2_X1 U9766 ( .A(n9717), .B(n9718), .ZN(n9476) );
  XOR2_X1 U9767 ( .A(n9719), .B(n9720), .Z(n9718) );
  NAND2_X1 U9768 ( .A1(b_22_), .A2(a_28_), .ZN(n9720) );
  NAND2_X1 U9769 ( .A1(a_27_), .A2(n9716), .ZN(n9477) );
  NAND2_X1 U9770 ( .A1(n9721), .A2(n9722), .ZN(n9716) );
  NAND2_X1 U9771 ( .A1(n9723), .A2(b_23_), .ZN(n9722) );
  NOR2_X1 U9772 ( .A1(n9724), .A2(n7803), .ZN(n9723) );
  NOR2_X1 U9773 ( .A1(n9483), .A2(n9485), .ZN(n9724) );
  NAND2_X1 U9774 ( .A1(n9483), .A2(n9485), .ZN(n9721) );
  NAND2_X1 U9775 ( .A1(n9725), .A2(n9726), .ZN(n9485) );
  NAND2_X1 U9776 ( .A1(n9503), .A2(n9727), .ZN(n9726) );
  NAND2_X1 U9777 ( .A1(n9505), .A2(n9504), .ZN(n9727) );
  NOR2_X1 U9778 ( .A1(n9256), .A2(n7337), .ZN(n9503) );
  OR2_X1 U9779 ( .A1(n9504), .A2(n9505), .ZN(n9725) );
  AND2_X1 U9780 ( .A1(n9728), .A2(n9729), .ZN(n9505) );
  NAND2_X1 U9781 ( .A1(n9730), .A2(b_21_), .ZN(n9729) );
  NOR2_X1 U9782 ( .A1(n9731), .A2(n7817), .ZN(n9730) );
  NOR2_X1 U9783 ( .A1(n7816), .A2(n9500), .ZN(n9731) );
  NAND2_X1 U9784 ( .A1(n9732), .A2(b_22_), .ZN(n9728) );
  NOR2_X1 U9785 ( .A1(n9733), .A2(n8052), .ZN(n9732) );
  NOR2_X1 U9786 ( .A1(n7810), .A2(n9734), .ZN(n9733) );
  NAND2_X1 U9787 ( .A1(n9501), .A2(b_22_), .ZN(n9504) );
  NOR2_X1 U9788 ( .A1(n8055), .A2(n9256), .ZN(n9501) );
  XOR2_X1 U9789 ( .A(n9735), .B(n9736), .Z(n9483) );
  XOR2_X1 U9790 ( .A(n9737), .B(n9738), .Z(n9735) );
  XNOR2_X1 U9791 ( .A(n9739), .B(n9740), .ZN(n9511) );
  NAND2_X1 U9792 ( .A1(n9741), .A2(n9742), .ZN(n9739) );
  XOR2_X1 U9793 ( .A(n9743), .B(n9744), .Z(n9515) );
  XOR2_X1 U9794 ( .A(n9745), .B(n9746), .Z(n9743) );
  XOR2_X1 U9795 ( .A(n9747), .B(n9748), .Z(n9519) );
  XOR2_X1 U9796 ( .A(n9749), .B(n9750), .Z(n9747) );
  NOR2_X1 U9797 ( .A1(n7774), .A2(n9500), .ZN(n9750) );
  XOR2_X1 U9798 ( .A(n9751), .B(n9752), .Z(n9522) );
  XOR2_X1 U9799 ( .A(n9753), .B(n9754), .Z(n9751) );
  XNOR2_X1 U9800 ( .A(n9755), .B(n9756), .ZN(n9527) );
  XNOR2_X1 U9801 ( .A(n9757), .B(n9758), .ZN(n9755) );
  XNOR2_X1 U9802 ( .A(n9759), .B(n9760), .ZN(n9531) );
  XNOR2_X1 U9803 ( .A(n9761), .B(n9762), .ZN(n9760) );
  XNOR2_X1 U9804 ( .A(n9763), .B(n9764), .ZN(n9534) );
  XOR2_X1 U9805 ( .A(n9765), .B(n9766), .Z(n9764) );
  NAND2_X1 U9806 ( .A1(b_22_), .A2(a_20_), .ZN(n9766) );
  XOR2_X1 U9807 ( .A(n9767), .B(n9768), .Z(n9538) );
  XOR2_X1 U9808 ( .A(n9769), .B(n9770), .Z(n9767) );
  XOR2_X1 U9809 ( .A(n9771), .B(n9772), .Z(n9542) );
  XOR2_X1 U9810 ( .A(n9773), .B(n9774), .Z(n9771) );
  NOR2_X1 U9811 ( .A1(n7745), .A2(n9500), .ZN(n9774) );
  XOR2_X1 U9812 ( .A(n9775), .B(n9776), .Z(n9547) );
  XOR2_X1 U9813 ( .A(n9777), .B(n9778), .Z(n9775) );
  XOR2_X1 U9814 ( .A(n9779), .B(n9780), .Z(n9551) );
  XOR2_X1 U9815 ( .A(n9781), .B(n9782), .Z(n9779) );
  NOR2_X1 U9816 ( .A1(n7736), .A2(n9500), .ZN(n9782) );
  XOR2_X1 U9817 ( .A(n9783), .B(n9784), .Z(n9559) );
  XOR2_X1 U9818 ( .A(n9785), .B(n9786), .Z(n9783) );
  NOR2_X1 U9819 ( .A1(n7727), .A2(n9500), .ZN(n9786) );
  XOR2_X1 U9820 ( .A(n9787), .B(n9788), .Z(n9563) );
  XOR2_X1 U9821 ( .A(n9789), .B(n9790), .Z(n9787) );
  XNOR2_X1 U9822 ( .A(n9791), .B(n9792), .ZN(n9567) );
  XOR2_X1 U9823 ( .A(n9793), .B(n9794), .Z(n9792) );
  NAND2_X1 U9824 ( .A1(b_22_), .A2(a_12_), .ZN(n9794) );
  XOR2_X1 U9825 ( .A(n9795), .B(n9796), .Z(n9570) );
  XOR2_X1 U9826 ( .A(n9797), .B(n9798), .Z(n9795) );
  XOR2_X1 U9827 ( .A(n9799), .B(n9800), .Z(n9575) );
  XOR2_X1 U9828 ( .A(n9801), .B(n9802), .Z(n9799) );
  NOR2_X1 U9829 ( .A1(n7709), .A2(n9500), .ZN(n9802) );
  XOR2_X1 U9830 ( .A(n9803), .B(n9804), .Z(n9405) );
  XOR2_X1 U9831 ( .A(n9805), .B(n9806), .Z(n9803) );
  NOR2_X1 U9832 ( .A1(n7704), .A2(n9500), .ZN(n9806) );
  XNOR2_X1 U9833 ( .A(n9807), .B(n9808), .ZN(n9579) );
  XNOR2_X1 U9834 ( .A(n9809), .B(n9810), .ZN(n9807) );
  XNOR2_X1 U9835 ( .A(n9811), .B(n9812), .ZN(n9587) );
  XNOR2_X1 U9836 ( .A(n9813), .B(n9814), .ZN(n9812) );
  XNOR2_X1 U9837 ( .A(n9815), .B(n9816), .ZN(n9386) );
  XOR2_X1 U9838 ( .A(n9817), .B(n9818), .Z(n9816) );
  NAND2_X1 U9839 ( .A1(b_22_), .A2(a_5_), .ZN(n9818) );
  XNOR2_X1 U9840 ( .A(n9819), .B(n9820), .ZN(n9378) );
  NAND2_X1 U9841 ( .A1(n9821), .A2(n9822), .ZN(n9819) );
  XNOR2_X1 U9842 ( .A(n9823), .B(n9824), .ZN(n9590) );
  XNOR2_X1 U9843 ( .A(n9825), .B(n9826), .ZN(n9824) );
  XNOR2_X1 U9844 ( .A(n9827), .B(n9828), .ZN(n9594) );
  XNOR2_X1 U9845 ( .A(n9829), .B(n9830), .ZN(n9827) );
  XNOR2_X1 U9846 ( .A(n9831), .B(n9832), .ZN(n9364) );
  XOR2_X1 U9847 ( .A(n9833), .B(n9834), .Z(n9832) );
  NAND2_X1 U9848 ( .A1(b_22_), .A2(a_1_), .ZN(n9834) );
  NOR2_X1 U9849 ( .A1(n9835), .A2(n7635), .ZN(n9598) );
  XOR2_X1 U9850 ( .A(n9836), .B(n9837), .Z(n7635) );
  XNOR2_X1 U9851 ( .A(n9838), .B(n9839), .ZN(n9836) );
  NOR2_X1 U9852 ( .A1(n7628), .A2(n7629), .ZN(n9835) );
  NAND2_X1 U9853 ( .A1(n9600), .A2(n9840), .ZN(n7523) );
  NAND2_X1 U9854 ( .A1(n9841), .A2(n7621), .ZN(n9840) );
  NAND2_X1 U9855 ( .A1(n9842), .A2(n9843), .ZN(n7522) );
  INV_X1 U9856 ( .A(n9600), .ZN(n9843) );
  NAND2_X1 U9857 ( .A1(n7628), .A2(n7629), .ZN(n9600) );
  NAND2_X1 U9858 ( .A1(n9844), .A2(n9845), .ZN(n7629) );
  NAND2_X1 U9859 ( .A1(n9839), .A2(n9846), .ZN(n9845) );
  NAND2_X1 U9860 ( .A1(n9838), .A2(n9837), .ZN(n9846) );
  NOR2_X1 U9861 ( .A1(n9500), .A2(n7478), .ZN(n9839) );
  OR2_X1 U9862 ( .A1(n9837), .A2(n9838), .ZN(n9844) );
  AND2_X1 U9863 ( .A1(n9847), .A2(n9848), .ZN(n9838) );
  NAND2_X1 U9864 ( .A1(n9849), .A2(b_22_), .ZN(n9848) );
  NOR2_X1 U9865 ( .A1(n9850), .A2(n7669), .ZN(n9849) );
  NOR2_X1 U9866 ( .A1(n9831), .A2(n9833), .ZN(n9850) );
  NAND2_X1 U9867 ( .A1(n9831), .A2(n9833), .ZN(n9847) );
  NAND2_X1 U9868 ( .A1(n9851), .A2(n9852), .ZN(n9833) );
  NAND2_X1 U9869 ( .A1(n9830), .A2(n9853), .ZN(n9852) );
  NAND2_X1 U9870 ( .A1(n9829), .A2(n9828), .ZN(n9853) );
  NOR2_X1 U9871 ( .A1(n9500), .A2(n7469), .ZN(n9830) );
  OR2_X1 U9872 ( .A1(n9828), .A2(n9829), .ZN(n9851) );
  AND2_X1 U9873 ( .A1(n9854), .A2(n9855), .ZN(n9829) );
  NAND2_X1 U9874 ( .A1(n9826), .A2(n9856), .ZN(n9855) );
  OR2_X1 U9875 ( .A1(n9823), .A2(n9825), .ZN(n9856) );
  NOR2_X1 U9876 ( .A1(n9500), .A2(n7464), .ZN(n9826) );
  NAND2_X1 U9877 ( .A1(n9823), .A2(n9825), .ZN(n9854) );
  NAND2_X1 U9878 ( .A1(n9821), .A2(n9857), .ZN(n9825) );
  NAND2_X1 U9879 ( .A1(n9820), .A2(n9822), .ZN(n9857) );
  NAND2_X1 U9880 ( .A1(n9858), .A2(n9859), .ZN(n9822) );
  NAND2_X1 U9881 ( .A1(b_22_), .A2(a_4_), .ZN(n9859) );
  INV_X1 U9882 ( .A(n9860), .ZN(n9858) );
  XOR2_X1 U9883 ( .A(n9861), .B(n9862), .Z(n9820) );
  XOR2_X1 U9884 ( .A(n9863), .B(n9864), .Z(n9861) );
  NOR2_X1 U9885 ( .A1(n7455), .A2(n9734), .ZN(n9864) );
  NAND2_X1 U9886 ( .A1(a_4_), .A2(n9860), .ZN(n9821) );
  NAND2_X1 U9887 ( .A1(n9865), .A2(n9866), .ZN(n9860) );
  NAND2_X1 U9888 ( .A1(n9867), .A2(b_22_), .ZN(n9866) );
  NOR2_X1 U9889 ( .A1(n9868), .A2(n7455), .ZN(n9867) );
  NOR2_X1 U9890 ( .A1(n9815), .A2(n9817), .ZN(n9868) );
  NAND2_X1 U9891 ( .A1(n9815), .A2(n9817), .ZN(n9865) );
  NAND2_X1 U9892 ( .A1(n9869), .A2(n9870), .ZN(n9817) );
  NAND2_X1 U9893 ( .A1(n9814), .A2(n9871), .ZN(n9870) );
  OR2_X1 U9894 ( .A1(n9813), .A2(n9811), .ZN(n9871) );
  NOR2_X1 U9895 ( .A1(n9500), .A2(n7450), .ZN(n9814) );
  NAND2_X1 U9896 ( .A1(n9811), .A2(n9813), .ZN(n9869) );
  NAND2_X1 U9897 ( .A1(n9872), .A2(n9873), .ZN(n9813) );
  NAND2_X1 U9898 ( .A1(n9632), .A2(n9874), .ZN(n9873) );
  OR2_X1 U9899 ( .A1(n9629), .A2(n9631), .ZN(n9874) );
  NOR2_X1 U9900 ( .A1(n9500), .A2(n7445), .ZN(n9632) );
  NAND2_X1 U9901 ( .A1(n9629), .A2(n9631), .ZN(n9872) );
  NAND2_X1 U9902 ( .A1(n9875), .A2(n9876), .ZN(n9631) );
  NAND2_X1 U9903 ( .A1(n9810), .A2(n9877), .ZN(n9876) );
  NAND2_X1 U9904 ( .A1(n9809), .A2(n9808), .ZN(n9877) );
  NOR2_X1 U9905 ( .A1(n9500), .A2(n7699), .ZN(n9810) );
  OR2_X1 U9906 ( .A1(n9808), .A2(n9809), .ZN(n9875) );
  AND2_X1 U9907 ( .A1(n9878), .A2(n9879), .ZN(n9809) );
  NAND2_X1 U9908 ( .A1(n9880), .A2(b_22_), .ZN(n9879) );
  NOR2_X1 U9909 ( .A1(n9881), .A2(n7704), .ZN(n9880) );
  NOR2_X1 U9910 ( .A1(n9804), .A2(n9805), .ZN(n9881) );
  NAND2_X1 U9911 ( .A1(n9804), .A2(n9805), .ZN(n9878) );
  NAND2_X1 U9912 ( .A1(n9882), .A2(n9883), .ZN(n9805) );
  NAND2_X1 U9913 ( .A1(n9884), .A2(b_22_), .ZN(n9883) );
  NOR2_X1 U9914 ( .A1(n9885), .A2(n7709), .ZN(n9884) );
  NOR2_X1 U9915 ( .A1(n9800), .A2(n9801), .ZN(n9885) );
  NAND2_X1 U9916 ( .A1(n9800), .A2(n9801), .ZN(n9882) );
  NAND2_X1 U9917 ( .A1(n9886), .A2(n9887), .ZN(n9801) );
  NAND2_X1 U9918 ( .A1(n9798), .A2(n9888), .ZN(n9887) );
  OR2_X1 U9919 ( .A1(n9796), .A2(n9797), .ZN(n9888) );
  NOR2_X1 U9920 ( .A1(n9500), .A2(n7424), .ZN(n9798) );
  NAND2_X1 U9921 ( .A1(n9796), .A2(n9797), .ZN(n9886) );
  NAND2_X1 U9922 ( .A1(n9889), .A2(n9890), .ZN(n9797) );
  NAND2_X1 U9923 ( .A1(n9891), .A2(b_22_), .ZN(n9890) );
  NOR2_X1 U9924 ( .A1(n9892), .A2(n7718), .ZN(n9891) );
  NOR2_X1 U9925 ( .A1(n9791), .A2(n9793), .ZN(n9892) );
  NAND2_X1 U9926 ( .A1(n9791), .A2(n9793), .ZN(n9889) );
  NAND2_X1 U9927 ( .A1(n9893), .A2(n9894), .ZN(n9793) );
  NAND2_X1 U9928 ( .A1(n9790), .A2(n9895), .ZN(n9894) );
  OR2_X1 U9929 ( .A1(n9788), .A2(n9789), .ZN(n9895) );
  NOR2_X1 U9930 ( .A1(n9500), .A2(n7415), .ZN(n9790) );
  NAND2_X1 U9931 ( .A1(n9788), .A2(n9789), .ZN(n9893) );
  NAND2_X1 U9932 ( .A1(n9896), .A2(n9897), .ZN(n9789) );
  NAND2_X1 U9933 ( .A1(n9898), .A2(b_22_), .ZN(n9897) );
  NOR2_X1 U9934 ( .A1(n9899), .A2(n7727), .ZN(n9898) );
  NOR2_X1 U9935 ( .A1(n9784), .A2(n9785), .ZN(n9899) );
  NAND2_X1 U9936 ( .A1(n9784), .A2(n9785), .ZN(n9896) );
  NAND2_X1 U9937 ( .A1(n9900), .A2(n9901), .ZN(n9785) );
  NAND2_X1 U9938 ( .A1(n9665), .A2(n9902), .ZN(n9901) );
  OR2_X1 U9939 ( .A1(n9663), .A2(n9664), .ZN(n9902) );
  NOR2_X1 U9940 ( .A1(n9500), .A2(n7406), .ZN(n9665) );
  NAND2_X1 U9941 ( .A1(n9663), .A2(n9664), .ZN(n9900) );
  NAND2_X1 U9942 ( .A1(n9903), .A2(n9904), .ZN(n9664) );
  NAND2_X1 U9943 ( .A1(n9905), .A2(b_22_), .ZN(n9904) );
  NOR2_X1 U9944 ( .A1(n9906), .A2(n7736), .ZN(n9905) );
  NOR2_X1 U9945 ( .A1(n9780), .A2(n9781), .ZN(n9906) );
  NAND2_X1 U9946 ( .A1(n9780), .A2(n9781), .ZN(n9903) );
  NAND2_X1 U9947 ( .A1(n9907), .A2(n9908), .ZN(n9781) );
  NAND2_X1 U9948 ( .A1(n9778), .A2(n9909), .ZN(n9908) );
  OR2_X1 U9949 ( .A1(n9776), .A2(n9777), .ZN(n9909) );
  NOR2_X1 U9950 ( .A1(n9500), .A2(n7397), .ZN(n9778) );
  NAND2_X1 U9951 ( .A1(n9776), .A2(n9777), .ZN(n9907) );
  NAND2_X1 U9952 ( .A1(n9910), .A2(n9911), .ZN(n9777) );
  NAND2_X1 U9953 ( .A1(n9912), .A2(b_22_), .ZN(n9911) );
  NOR2_X1 U9954 ( .A1(n9913), .A2(n7745), .ZN(n9912) );
  NOR2_X1 U9955 ( .A1(n9773), .A2(n9772), .ZN(n9913) );
  NAND2_X1 U9956 ( .A1(n9772), .A2(n9773), .ZN(n9910) );
  NAND2_X1 U9957 ( .A1(n9914), .A2(n9915), .ZN(n9773) );
  NAND2_X1 U9958 ( .A1(n9770), .A2(n9916), .ZN(n9915) );
  OR2_X1 U9959 ( .A1(n9768), .A2(n9769), .ZN(n9916) );
  NOR2_X1 U9960 ( .A1(n9500), .A2(n7750), .ZN(n9770) );
  NAND2_X1 U9961 ( .A1(n9768), .A2(n9769), .ZN(n9914) );
  NAND2_X1 U9962 ( .A1(n9917), .A2(n9918), .ZN(n9769) );
  NAND2_X1 U9963 ( .A1(n9919), .A2(b_22_), .ZN(n9918) );
  NOR2_X1 U9964 ( .A1(n9920), .A2(n7755), .ZN(n9919) );
  NOR2_X1 U9965 ( .A1(n9763), .A2(n9765), .ZN(n9920) );
  NAND2_X1 U9966 ( .A1(n9763), .A2(n9765), .ZN(n9917) );
  NAND2_X1 U9967 ( .A1(n9921), .A2(n9922), .ZN(n9765) );
  NAND2_X1 U9968 ( .A1(n9762), .A2(n9923), .ZN(n9922) );
  OR2_X1 U9969 ( .A1(n9759), .A2(n9761), .ZN(n9923) );
  NOR2_X1 U9970 ( .A1(n9500), .A2(n7760), .ZN(n9762) );
  NAND2_X1 U9971 ( .A1(n9759), .A2(n9761), .ZN(n9921) );
  NAND2_X1 U9972 ( .A1(n9924), .A2(n9925), .ZN(n9761) );
  NAND2_X1 U9973 ( .A1(n9758), .A2(n9926), .ZN(n9925) );
  NAND2_X1 U9974 ( .A1(n9757), .A2(n9756), .ZN(n9926) );
  OR2_X1 U9975 ( .A1(n9756), .A2(n9757), .ZN(n9924) );
  AND2_X1 U9976 ( .A1(n9927), .A2(n9928), .ZN(n9757) );
  NAND2_X1 U9977 ( .A1(n9754), .A2(n9929), .ZN(n9928) );
  OR2_X1 U9978 ( .A1(n9752), .A2(n9753), .ZN(n9929) );
  NOR2_X1 U9979 ( .A1(n9500), .A2(n8014), .ZN(n9754) );
  NAND2_X1 U9980 ( .A1(n9752), .A2(n9753), .ZN(n9927) );
  NAND2_X1 U9981 ( .A1(n9930), .A2(n9931), .ZN(n9753) );
  NAND2_X1 U9982 ( .A1(n9932), .A2(b_22_), .ZN(n9931) );
  NOR2_X1 U9983 ( .A1(n9933), .A2(n7774), .ZN(n9932) );
  NOR2_X1 U9984 ( .A1(n9748), .A2(n9749), .ZN(n9933) );
  NAND2_X1 U9985 ( .A1(n9748), .A2(n9749), .ZN(n9930) );
  NAND2_X1 U9986 ( .A1(n9934), .A2(n9935), .ZN(n9749) );
  NAND2_X1 U9987 ( .A1(n9746), .A2(n9936), .ZN(n9935) );
  OR2_X1 U9988 ( .A1(n9744), .A2(n9745), .ZN(n9936) );
  NOR2_X1 U9989 ( .A1(n9500), .A2(n8022), .ZN(n9746) );
  NAND2_X1 U9990 ( .A1(n9744), .A2(n9745), .ZN(n9934) );
  NAND2_X1 U9991 ( .A1(n9741), .A2(n9937), .ZN(n9745) );
  NAND2_X1 U9992 ( .A1(n9740), .A2(n9742), .ZN(n9937) );
  NAND2_X1 U9993 ( .A1(n9938), .A2(n9939), .ZN(n9742) );
  NAND2_X1 U9994 ( .A1(b_22_), .A2(a_26_), .ZN(n9939) );
  INV_X1 U9995 ( .A(n9940), .ZN(n9938) );
  XNOR2_X1 U9996 ( .A(n9941), .B(n9942), .ZN(n9740) );
  NAND2_X1 U9997 ( .A1(n9943), .A2(n9944), .ZN(n9941) );
  NAND2_X1 U9998 ( .A1(a_26_), .A2(n9940), .ZN(n9741) );
  NAND2_X1 U9999 ( .A1(n9711), .A2(n9945), .ZN(n9940) );
  NAND2_X1 U10000 ( .A1(n9710), .A2(n9712), .ZN(n9945) );
  NAND2_X1 U10001 ( .A1(n9946), .A2(n9947), .ZN(n9712) );
  NAND2_X1 U10002 ( .A1(b_22_), .A2(a_27_), .ZN(n9947) );
  INV_X1 U10003 ( .A(n9948), .ZN(n9946) );
  XNOR2_X1 U10004 ( .A(n9949), .B(n9950), .ZN(n9710) );
  XOR2_X1 U10005 ( .A(n9951), .B(n9952), .Z(n9950) );
  NAND2_X1 U10006 ( .A1(b_21_), .A2(a_28_), .ZN(n9952) );
  NAND2_X1 U10007 ( .A1(a_27_), .A2(n9948), .ZN(n9711) );
  NAND2_X1 U10008 ( .A1(n9953), .A2(n9954), .ZN(n9948) );
  NAND2_X1 U10009 ( .A1(n9955), .A2(b_22_), .ZN(n9954) );
  NOR2_X1 U10010 ( .A1(n9956), .A2(n7803), .ZN(n9955) );
  NOR2_X1 U10011 ( .A1(n9717), .A2(n9719), .ZN(n9956) );
  NAND2_X1 U10012 ( .A1(n9717), .A2(n9719), .ZN(n9953) );
  NAND2_X1 U10013 ( .A1(n9957), .A2(n9958), .ZN(n9719) );
  NAND2_X1 U10014 ( .A1(n9736), .A2(n9959), .ZN(n9958) );
  NAND2_X1 U10015 ( .A1(n9738), .A2(n9737), .ZN(n9959) );
  NOR2_X1 U10016 ( .A1(n9500), .A2(n7337), .ZN(n9736) );
  OR2_X1 U10017 ( .A1(n9737), .A2(n9738), .ZN(n9957) );
  AND2_X1 U10018 ( .A1(n9960), .A2(n9961), .ZN(n9738) );
  NAND2_X1 U10019 ( .A1(n9962), .A2(b_20_), .ZN(n9961) );
  NOR2_X1 U10020 ( .A1(n9963), .A2(n7817), .ZN(n9962) );
  NOR2_X1 U10021 ( .A1(n7816), .A2(n9734), .ZN(n9963) );
  NAND2_X1 U10022 ( .A1(n9964), .A2(b_21_), .ZN(n9960) );
  NOR2_X1 U10023 ( .A1(n9965), .A2(n8052), .ZN(n9964) );
  NOR2_X1 U10024 ( .A1(n7810), .A2(n9966), .ZN(n9965) );
  NAND2_X1 U10025 ( .A1(n9967), .A2(b_22_), .ZN(n9737) );
  NOR2_X1 U10026 ( .A1(n8055), .A2(n9734), .ZN(n9967) );
  XOR2_X1 U10027 ( .A(n9968), .B(n9969), .Z(n9717) );
  XOR2_X1 U10028 ( .A(n9970), .B(n9971), .Z(n9968) );
  XNOR2_X1 U10029 ( .A(n9972), .B(n9973), .ZN(n9744) );
  NAND2_X1 U10030 ( .A1(n9974), .A2(n9975), .ZN(n9972) );
  XOR2_X1 U10031 ( .A(n9976), .B(n9977), .Z(n9748) );
  XOR2_X1 U10032 ( .A(n9978), .B(n9979), .Z(n9976) );
  XOR2_X1 U10033 ( .A(n9980), .B(n9981), .Z(n9752) );
  XNOR2_X1 U10034 ( .A(n9982), .B(n9983), .ZN(n9980) );
  NAND2_X1 U10035 ( .A1(b_21_), .A2(a_24_), .ZN(n9982) );
  XNOR2_X1 U10036 ( .A(n9984), .B(n9985), .ZN(n9756) );
  XOR2_X1 U10037 ( .A(n9986), .B(n9987), .Z(n9984) );
  XNOR2_X1 U10038 ( .A(n9988), .B(n9989), .ZN(n9759) );
  XOR2_X1 U10039 ( .A(n9990), .B(n9991), .Z(n9989) );
  NAND2_X1 U10040 ( .A1(b_21_), .A2(a_22_), .ZN(n9991) );
  XOR2_X1 U10041 ( .A(n9992), .B(n9993), .Z(n9763) );
  XOR2_X1 U10042 ( .A(n9994), .B(n9995), .Z(n9992) );
  XOR2_X1 U10043 ( .A(n9996), .B(n9997), .Z(n9768) );
  XOR2_X1 U10044 ( .A(n9998), .B(n9999), .Z(n9996) );
  NOR2_X1 U10045 ( .A1(n7755), .A2(n9734), .ZN(n9999) );
  XNOR2_X1 U10046 ( .A(n10000), .B(n10001), .ZN(n9772) );
  XNOR2_X1 U10047 ( .A(n10002), .B(n10003), .ZN(n10001) );
  XOR2_X1 U10048 ( .A(n10004), .B(n10005), .Z(n9776) );
  XOR2_X1 U10049 ( .A(n10006), .B(n10007), .Z(n10004) );
  NOR2_X1 U10050 ( .A1(n7745), .A2(n9734), .ZN(n10007) );
  XNOR2_X1 U10051 ( .A(n10008), .B(n10009), .ZN(n9780) );
  XNOR2_X1 U10052 ( .A(n10010), .B(n10011), .ZN(n10009) );
  XOR2_X1 U10053 ( .A(n10012), .B(n10013), .Z(n9663) );
  XOR2_X1 U10054 ( .A(n10014), .B(n10015), .Z(n10012) );
  NOR2_X1 U10055 ( .A1(n7736), .A2(n9734), .ZN(n10015) );
  XOR2_X1 U10056 ( .A(n10016), .B(n10017), .Z(n9784) );
  XOR2_X1 U10057 ( .A(n10018), .B(n10019), .Z(n10016) );
  XNOR2_X1 U10058 ( .A(n10020), .B(n10021), .ZN(n9788) );
  XOR2_X1 U10059 ( .A(n10022), .B(n10023), .Z(n10021) );
  NAND2_X1 U10060 ( .A1(b_21_), .A2(a_14_), .ZN(n10023) );
  XOR2_X1 U10061 ( .A(n10024), .B(n10025), .Z(n9791) );
  XOR2_X1 U10062 ( .A(n10026), .B(n10027), .Z(n10024) );
  XOR2_X1 U10063 ( .A(n10028), .B(n10029), .Z(n9796) );
  XOR2_X1 U10064 ( .A(n10030), .B(n10031), .Z(n10028) );
  NOR2_X1 U10065 ( .A1(n7718), .A2(n9734), .ZN(n10031) );
  XOR2_X1 U10066 ( .A(n10032), .B(n10033), .Z(n9800) );
  XOR2_X1 U10067 ( .A(n10034), .B(n10035), .Z(n10032) );
  XNOR2_X1 U10068 ( .A(n10036), .B(n10037), .ZN(n9804) );
  XNOR2_X1 U10069 ( .A(n10038), .B(n10039), .ZN(n10037) );
  XOR2_X1 U10070 ( .A(n10040), .B(n10041), .Z(n9808) );
  XOR2_X1 U10071 ( .A(n10042), .B(n10043), .Z(n10041) );
  NAND2_X1 U10072 ( .A1(b_21_), .A2(a_9_), .ZN(n10043) );
  XOR2_X1 U10073 ( .A(n10044), .B(n10045), .Z(n9629) );
  XOR2_X1 U10074 ( .A(n10046), .B(n10047), .Z(n10044) );
  NOR2_X1 U10075 ( .A1(n7699), .A2(n9734), .ZN(n10047) );
  XOR2_X1 U10076 ( .A(n10048), .B(n10049), .Z(n9811) );
  XOR2_X1 U10077 ( .A(n10050), .B(n10051), .Z(n10048) );
  NOR2_X1 U10078 ( .A1(n7445), .A2(n9734), .ZN(n10051) );
  XOR2_X1 U10079 ( .A(n10052), .B(n10053), .Z(n9815) );
  XOR2_X1 U10080 ( .A(n10054), .B(n10055), .Z(n10052) );
  NOR2_X1 U10081 ( .A1(n7450), .A2(n9734), .ZN(n10055) );
  XNOR2_X1 U10082 ( .A(n10056), .B(n10057), .ZN(n9823) );
  XOR2_X1 U10083 ( .A(n10058), .B(n10059), .Z(n10057) );
  NAND2_X1 U10084 ( .A1(b_21_), .A2(a_4_), .ZN(n10059) );
  XNOR2_X1 U10085 ( .A(n10060), .B(n10061), .ZN(n9828) );
  XOR2_X1 U10086 ( .A(n10062), .B(n10063), .Z(n10060) );
  NOR2_X1 U10087 ( .A1(n7464), .A2(n9734), .ZN(n10063) );
  XOR2_X1 U10088 ( .A(n10064), .B(n10065), .Z(n9831) );
  XOR2_X1 U10089 ( .A(n10066), .B(n10067), .Z(n10064) );
  NOR2_X1 U10090 ( .A1(n7469), .A2(n9734), .ZN(n10067) );
  XNOR2_X1 U10091 ( .A(n10068), .B(n10069), .ZN(n9837) );
  XOR2_X1 U10092 ( .A(n10070), .B(n10071), .Z(n10068) );
  NOR2_X1 U10093 ( .A1(n7669), .A2(n9734), .ZN(n10071) );
  XNOR2_X1 U10094 ( .A(n10072), .B(n10073), .ZN(n7628) );
  XNOR2_X1 U10095 ( .A(n10074), .B(n10075), .ZN(n10072) );
  AND2_X1 U10096 ( .A1(n7621), .A2(n9841), .ZN(n9842) );
  NAND2_X1 U10097 ( .A1(n10076), .A2(n10077), .ZN(n9841) );
  XOR2_X1 U10098 ( .A(n10078), .B(n10079), .Z(n10077) );
  NOR2_X1 U10099 ( .A1(n10080), .A2(n10081), .ZN(n10076) );
  NOR2_X1 U10100 ( .A1(n10074), .A2(n10073), .ZN(n10081) );
  INV_X1 U10101 ( .A(n10082), .ZN(n10080) );
  OR2_X1 U10102 ( .A1(n7621), .A2(n7620), .ZN(n7527) );
  XNOR2_X1 U10103 ( .A(n7618), .B(n7617), .ZN(n7620) );
  NAND2_X1 U10104 ( .A1(n10083), .A2(n10084), .ZN(n7621) );
  NAND2_X1 U10105 ( .A1(n10085), .A2(n10082), .ZN(n10084) );
  NAND2_X1 U10106 ( .A1(n10075), .A2(n10086), .ZN(n10082) );
  NAND2_X1 U10107 ( .A1(n10074), .A2(n10073), .ZN(n10086) );
  NOR2_X1 U10108 ( .A1(n9734), .A2(n7478), .ZN(n10075) );
  OR2_X1 U10109 ( .A1(n10073), .A2(n10074), .ZN(n10085) );
  AND2_X1 U10110 ( .A1(n10087), .A2(n10088), .ZN(n10074) );
  NAND2_X1 U10111 ( .A1(n10089), .A2(b_21_), .ZN(n10088) );
  NOR2_X1 U10112 ( .A1(n10090), .A2(n7669), .ZN(n10089) );
  NOR2_X1 U10113 ( .A1(n10069), .A2(n10070), .ZN(n10090) );
  NAND2_X1 U10114 ( .A1(n10069), .A2(n10070), .ZN(n10087) );
  NAND2_X1 U10115 ( .A1(n10091), .A2(n10092), .ZN(n10070) );
  NAND2_X1 U10116 ( .A1(n10093), .A2(b_21_), .ZN(n10092) );
  NOR2_X1 U10117 ( .A1(n10094), .A2(n7469), .ZN(n10093) );
  NOR2_X1 U10118 ( .A1(n10065), .A2(n10066), .ZN(n10094) );
  NAND2_X1 U10119 ( .A1(n10065), .A2(n10066), .ZN(n10091) );
  NAND2_X1 U10120 ( .A1(n10095), .A2(n10096), .ZN(n10066) );
  NAND2_X1 U10121 ( .A1(n10097), .A2(b_21_), .ZN(n10096) );
  NOR2_X1 U10122 ( .A1(n10098), .A2(n7464), .ZN(n10097) );
  NOR2_X1 U10123 ( .A1(n10061), .A2(n10062), .ZN(n10098) );
  NAND2_X1 U10124 ( .A1(n10061), .A2(n10062), .ZN(n10095) );
  NAND2_X1 U10125 ( .A1(n10099), .A2(n10100), .ZN(n10062) );
  NAND2_X1 U10126 ( .A1(n10101), .A2(b_21_), .ZN(n10100) );
  NOR2_X1 U10127 ( .A1(n10102), .A2(n7682), .ZN(n10101) );
  NOR2_X1 U10128 ( .A1(n10056), .A2(n10058), .ZN(n10102) );
  NAND2_X1 U10129 ( .A1(n10056), .A2(n10058), .ZN(n10099) );
  NAND2_X1 U10130 ( .A1(n10103), .A2(n10104), .ZN(n10058) );
  NAND2_X1 U10131 ( .A1(n10105), .A2(b_21_), .ZN(n10104) );
  NOR2_X1 U10132 ( .A1(n10106), .A2(n7455), .ZN(n10105) );
  NOR2_X1 U10133 ( .A1(n9862), .A2(n9863), .ZN(n10106) );
  NAND2_X1 U10134 ( .A1(n9862), .A2(n9863), .ZN(n10103) );
  NAND2_X1 U10135 ( .A1(n10107), .A2(n10108), .ZN(n9863) );
  NAND2_X1 U10136 ( .A1(n10109), .A2(b_21_), .ZN(n10108) );
  NOR2_X1 U10137 ( .A1(n10110), .A2(n7450), .ZN(n10109) );
  NOR2_X1 U10138 ( .A1(n10053), .A2(n10054), .ZN(n10110) );
  NAND2_X1 U10139 ( .A1(n10053), .A2(n10054), .ZN(n10107) );
  NAND2_X1 U10140 ( .A1(n10111), .A2(n10112), .ZN(n10054) );
  NAND2_X1 U10141 ( .A1(n10113), .A2(b_21_), .ZN(n10112) );
  NOR2_X1 U10142 ( .A1(n10114), .A2(n7445), .ZN(n10113) );
  NOR2_X1 U10143 ( .A1(n10049), .A2(n10050), .ZN(n10114) );
  NAND2_X1 U10144 ( .A1(n10049), .A2(n10050), .ZN(n10111) );
  NAND2_X1 U10145 ( .A1(n10115), .A2(n10116), .ZN(n10050) );
  NAND2_X1 U10146 ( .A1(n10117), .A2(b_21_), .ZN(n10116) );
  NOR2_X1 U10147 ( .A1(n10118), .A2(n7699), .ZN(n10117) );
  NOR2_X1 U10148 ( .A1(n10045), .A2(n10046), .ZN(n10118) );
  NAND2_X1 U10149 ( .A1(n10045), .A2(n10046), .ZN(n10115) );
  NAND2_X1 U10150 ( .A1(n10119), .A2(n10120), .ZN(n10046) );
  NAND2_X1 U10151 ( .A1(n10121), .A2(b_21_), .ZN(n10120) );
  NOR2_X1 U10152 ( .A1(n10122), .A2(n7704), .ZN(n10121) );
  NOR2_X1 U10153 ( .A1(n10040), .A2(n10042), .ZN(n10122) );
  NAND2_X1 U10154 ( .A1(n10040), .A2(n10042), .ZN(n10119) );
  NAND2_X1 U10155 ( .A1(n10123), .A2(n10124), .ZN(n10042) );
  NAND2_X1 U10156 ( .A1(n10039), .A2(n10125), .ZN(n10124) );
  OR2_X1 U10157 ( .A1(n10038), .A2(n10036), .ZN(n10125) );
  NOR2_X1 U10158 ( .A1(n9734), .A2(n7709), .ZN(n10039) );
  NAND2_X1 U10159 ( .A1(n10036), .A2(n10038), .ZN(n10123) );
  NAND2_X1 U10160 ( .A1(n10126), .A2(n10127), .ZN(n10038) );
  NAND2_X1 U10161 ( .A1(n10035), .A2(n10128), .ZN(n10127) );
  OR2_X1 U10162 ( .A1(n10034), .A2(n10033), .ZN(n10128) );
  NOR2_X1 U10163 ( .A1(n9734), .A2(n7424), .ZN(n10035) );
  NAND2_X1 U10164 ( .A1(n10033), .A2(n10034), .ZN(n10126) );
  NAND2_X1 U10165 ( .A1(n10129), .A2(n10130), .ZN(n10034) );
  NAND2_X1 U10166 ( .A1(n10131), .A2(b_21_), .ZN(n10130) );
  NOR2_X1 U10167 ( .A1(n10132), .A2(n7718), .ZN(n10131) );
  NOR2_X1 U10168 ( .A1(n10029), .A2(n10030), .ZN(n10132) );
  NAND2_X1 U10169 ( .A1(n10029), .A2(n10030), .ZN(n10129) );
  NAND2_X1 U10170 ( .A1(n10133), .A2(n10134), .ZN(n10030) );
  NAND2_X1 U10171 ( .A1(n10027), .A2(n10135), .ZN(n10134) );
  OR2_X1 U10172 ( .A1(n10026), .A2(n10025), .ZN(n10135) );
  NOR2_X1 U10173 ( .A1(n9734), .A2(n7415), .ZN(n10027) );
  NAND2_X1 U10174 ( .A1(n10025), .A2(n10026), .ZN(n10133) );
  NAND2_X1 U10175 ( .A1(n10136), .A2(n10137), .ZN(n10026) );
  NAND2_X1 U10176 ( .A1(n10138), .A2(b_21_), .ZN(n10137) );
  NOR2_X1 U10177 ( .A1(n10139), .A2(n7727), .ZN(n10138) );
  NOR2_X1 U10178 ( .A1(n10020), .A2(n10022), .ZN(n10139) );
  NAND2_X1 U10179 ( .A1(n10020), .A2(n10022), .ZN(n10136) );
  NAND2_X1 U10180 ( .A1(n10140), .A2(n10141), .ZN(n10022) );
  NAND2_X1 U10181 ( .A1(n10019), .A2(n10142), .ZN(n10141) );
  OR2_X1 U10182 ( .A1(n10018), .A2(n10017), .ZN(n10142) );
  NOR2_X1 U10183 ( .A1(n9734), .A2(n7406), .ZN(n10019) );
  NAND2_X1 U10184 ( .A1(n10017), .A2(n10018), .ZN(n10140) );
  NAND2_X1 U10185 ( .A1(n10143), .A2(n10144), .ZN(n10018) );
  NAND2_X1 U10186 ( .A1(n10145), .A2(b_21_), .ZN(n10144) );
  NOR2_X1 U10187 ( .A1(n10146), .A2(n7736), .ZN(n10145) );
  NOR2_X1 U10188 ( .A1(n10013), .A2(n10014), .ZN(n10146) );
  NAND2_X1 U10189 ( .A1(n10013), .A2(n10014), .ZN(n10143) );
  NAND2_X1 U10190 ( .A1(n10147), .A2(n10148), .ZN(n10014) );
  NAND2_X1 U10191 ( .A1(n10011), .A2(n10149), .ZN(n10148) );
  OR2_X1 U10192 ( .A1(n10010), .A2(n10008), .ZN(n10149) );
  NOR2_X1 U10193 ( .A1(n9734), .A2(n7397), .ZN(n10011) );
  NAND2_X1 U10194 ( .A1(n10008), .A2(n10010), .ZN(n10147) );
  NAND2_X1 U10195 ( .A1(n10150), .A2(n10151), .ZN(n10010) );
  NAND2_X1 U10196 ( .A1(n10152), .A2(b_21_), .ZN(n10151) );
  NOR2_X1 U10197 ( .A1(n10153), .A2(n7745), .ZN(n10152) );
  NOR2_X1 U10198 ( .A1(n10005), .A2(n10006), .ZN(n10153) );
  NAND2_X1 U10199 ( .A1(n10005), .A2(n10006), .ZN(n10150) );
  NAND2_X1 U10200 ( .A1(n10154), .A2(n10155), .ZN(n10006) );
  NAND2_X1 U10201 ( .A1(n10003), .A2(n10156), .ZN(n10155) );
  OR2_X1 U10202 ( .A1(n10002), .A2(n10000), .ZN(n10156) );
  NOR2_X1 U10203 ( .A1(n9734), .A2(n7750), .ZN(n10003) );
  NAND2_X1 U10204 ( .A1(n10000), .A2(n10002), .ZN(n10154) );
  NAND2_X1 U10205 ( .A1(n10157), .A2(n10158), .ZN(n10002) );
  NAND2_X1 U10206 ( .A1(n10159), .A2(b_21_), .ZN(n10158) );
  NOR2_X1 U10207 ( .A1(n10160), .A2(n7755), .ZN(n10159) );
  NOR2_X1 U10208 ( .A1(n9997), .A2(n9998), .ZN(n10160) );
  NAND2_X1 U10209 ( .A1(n9997), .A2(n9998), .ZN(n10157) );
  NAND2_X1 U10210 ( .A1(n10161), .A2(n10162), .ZN(n9998) );
  NAND2_X1 U10211 ( .A1(n9995), .A2(n10163), .ZN(n10162) );
  OR2_X1 U10212 ( .A1(n9994), .A2(n9993), .ZN(n10163) );
  NAND2_X1 U10213 ( .A1(n9993), .A2(n9994), .ZN(n10161) );
  NAND2_X1 U10214 ( .A1(n10164), .A2(n10165), .ZN(n9994) );
  NAND2_X1 U10215 ( .A1(n10166), .A2(b_21_), .ZN(n10165) );
  NOR2_X1 U10216 ( .A1(n10167), .A2(n7765), .ZN(n10166) );
  NOR2_X1 U10217 ( .A1(n9988), .A2(n9990), .ZN(n10167) );
  NAND2_X1 U10218 ( .A1(n9988), .A2(n9990), .ZN(n10164) );
  NAND2_X1 U10219 ( .A1(n10168), .A2(n10169), .ZN(n9990) );
  NAND2_X1 U10220 ( .A1(n9987), .A2(n10170), .ZN(n10169) );
  OR2_X1 U10221 ( .A1(n9986), .A2(n9985), .ZN(n10170) );
  NOR2_X1 U10222 ( .A1(n9734), .A2(n8014), .ZN(n9987) );
  NAND2_X1 U10223 ( .A1(n9985), .A2(n9986), .ZN(n10168) );
  NAND2_X1 U10224 ( .A1(n10171), .A2(n10172), .ZN(n9986) );
  NAND2_X1 U10225 ( .A1(n10173), .A2(b_21_), .ZN(n10172) );
  NOR2_X1 U10226 ( .A1(n10174), .A2(n7774), .ZN(n10173) );
  NOR2_X1 U10227 ( .A1(n9981), .A2(n9983), .ZN(n10174) );
  NAND2_X1 U10228 ( .A1(n9981), .A2(n9983), .ZN(n10171) );
  NAND2_X1 U10229 ( .A1(n10175), .A2(n10176), .ZN(n9983) );
  NAND2_X1 U10230 ( .A1(n9979), .A2(n10177), .ZN(n10176) );
  OR2_X1 U10231 ( .A1(n9978), .A2(n9977), .ZN(n10177) );
  NOR2_X1 U10232 ( .A1(n9734), .A2(n8022), .ZN(n9979) );
  NAND2_X1 U10233 ( .A1(n9977), .A2(n9978), .ZN(n10175) );
  NAND2_X1 U10234 ( .A1(n9974), .A2(n10178), .ZN(n9978) );
  NAND2_X1 U10235 ( .A1(n9973), .A2(n9975), .ZN(n10178) );
  NAND2_X1 U10236 ( .A1(n10179), .A2(n10180), .ZN(n9975) );
  NAND2_X1 U10237 ( .A1(b_21_), .A2(a_26_), .ZN(n10180) );
  INV_X1 U10238 ( .A(n10181), .ZN(n10179) );
  XNOR2_X1 U10239 ( .A(n10182), .B(n10183), .ZN(n9973) );
  NAND2_X1 U10240 ( .A1(n10184), .A2(n10185), .ZN(n10182) );
  NAND2_X1 U10241 ( .A1(a_26_), .A2(n10181), .ZN(n9974) );
  NAND2_X1 U10242 ( .A1(n9943), .A2(n10186), .ZN(n10181) );
  NAND2_X1 U10243 ( .A1(n9942), .A2(n9944), .ZN(n10186) );
  NAND2_X1 U10244 ( .A1(n10187), .A2(n10188), .ZN(n9944) );
  NAND2_X1 U10245 ( .A1(b_21_), .A2(a_27_), .ZN(n10188) );
  INV_X1 U10246 ( .A(n10189), .ZN(n10187) );
  XNOR2_X1 U10247 ( .A(n10190), .B(n10191), .ZN(n9942) );
  XOR2_X1 U10248 ( .A(n10192), .B(n10193), .Z(n10191) );
  NAND2_X1 U10249 ( .A1(b_20_), .A2(a_28_), .ZN(n10193) );
  NAND2_X1 U10250 ( .A1(a_27_), .A2(n10189), .ZN(n9943) );
  NAND2_X1 U10251 ( .A1(n10194), .A2(n10195), .ZN(n10189) );
  NAND2_X1 U10252 ( .A1(n10196), .A2(b_21_), .ZN(n10195) );
  NOR2_X1 U10253 ( .A1(n10197), .A2(n7803), .ZN(n10196) );
  NOR2_X1 U10254 ( .A1(n9949), .A2(n9951), .ZN(n10197) );
  NAND2_X1 U10255 ( .A1(n9949), .A2(n9951), .ZN(n10194) );
  NAND2_X1 U10256 ( .A1(n10198), .A2(n10199), .ZN(n9951) );
  NAND2_X1 U10257 ( .A1(n9969), .A2(n10200), .ZN(n10199) );
  NAND2_X1 U10258 ( .A1(n9971), .A2(n9970), .ZN(n10200) );
  NOR2_X1 U10259 ( .A1(n9734), .A2(n7337), .ZN(n9969) );
  OR2_X1 U10260 ( .A1(n9970), .A2(n9971), .ZN(n10198) );
  AND2_X1 U10261 ( .A1(n10201), .A2(n10202), .ZN(n9971) );
  NAND2_X1 U10262 ( .A1(n10203), .A2(b_19_), .ZN(n10202) );
  NOR2_X1 U10263 ( .A1(n10204), .A2(n7817), .ZN(n10203) );
  NOR2_X1 U10264 ( .A1(n7816), .A2(n9966), .ZN(n10204) );
  NAND2_X1 U10265 ( .A1(n10205), .A2(b_20_), .ZN(n10201) );
  NOR2_X1 U10266 ( .A1(n10206), .A2(n8052), .ZN(n10205) );
  NOR2_X1 U10267 ( .A1(n7810), .A2(n10207), .ZN(n10206) );
  NAND2_X1 U10268 ( .A1(n10208), .A2(b_21_), .ZN(n9970) );
  NOR2_X1 U10269 ( .A1(n8055), .A2(n9966), .ZN(n10208) );
  XOR2_X1 U10270 ( .A(n10209), .B(n10210), .Z(n9949) );
  XOR2_X1 U10271 ( .A(n10211), .B(n10212), .Z(n10209) );
  XNOR2_X1 U10272 ( .A(n10213), .B(n10214), .ZN(n9977) );
  NAND2_X1 U10273 ( .A1(n10215), .A2(n10216), .ZN(n10213) );
  XOR2_X1 U10274 ( .A(n10217), .B(n10218), .Z(n9981) );
  XOR2_X1 U10275 ( .A(n10219), .B(n10220), .Z(n10217) );
  XOR2_X1 U10276 ( .A(n10221), .B(n10222), .Z(n9985) );
  XNOR2_X1 U10277 ( .A(n10223), .B(n10224), .ZN(n10221) );
  NAND2_X1 U10278 ( .A1(b_20_), .A2(a_24_), .ZN(n10223) );
  XOR2_X1 U10279 ( .A(n10225), .B(n10226), .Z(n9988) );
  XOR2_X1 U10280 ( .A(n10227), .B(n10228), .Z(n10225) );
  XNOR2_X1 U10281 ( .A(n10229), .B(n10230), .ZN(n9993) );
  XOR2_X1 U10282 ( .A(n10231), .B(n10232), .Z(n10230) );
  NAND2_X1 U10283 ( .A1(b_20_), .A2(a_22_), .ZN(n10232) );
  XOR2_X1 U10284 ( .A(n10233), .B(n10234), .Z(n9997) );
  XOR2_X1 U10285 ( .A(n10235), .B(n10236), .Z(n10233) );
  XOR2_X1 U10286 ( .A(n10237), .B(n10238), .Z(n10000) );
  XOR2_X1 U10287 ( .A(n10239), .B(n10240), .Z(n10237) );
  XOR2_X1 U10288 ( .A(n10241), .B(n10242), .Z(n10005) );
  XOR2_X1 U10289 ( .A(n10243), .B(n10244), .Z(n10241) );
  XOR2_X1 U10290 ( .A(n10245), .B(n10246), .Z(n10008) );
  XOR2_X1 U10291 ( .A(n10247), .B(n10248), .Z(n10245) );
  NOR2_X1 U10292 ( .A1(n7745), .A2(n9966), .ZN(n10248) );
  XOR2_X1 U10293 ( .A(n10249), .B(n10250), .Z(n10013) );
  XOR2_X1 U10294 ( .A(n10251), .B(n10252), .Z(n10249) );
  XNOR2_X1 U10295 ( .A(n10253), .B(n10254), .ZN(n10017) );
  XOR2_X1 U10296 ( .A(n10255), .B(n10256), .Z(n10254) );
  NAND2_X1 U10297 ( .A1(b_20_), .A2(a_16_), .ZN(n10256) );
  XOR2_X1 U10298 ( .A(n10257), .B(n10258), .Z(n10020) );
  XOR2_X1 U10299 ( .A(n10259), .B(n10260), .Z(n10257) );
  XOR2_X1 U10300 ( .A(n10261), .B(n10262), .Z(n10025) );
  XOR2_X1 U10301 ( .A(n10263), .B(n10264), .Z(n10261) );
  NOR2_X1 U10302 ( .A1(n7727), .A2(n9966), .ZN(n10264) );
  XOR2_X1 U10303 ( .A(n10265), .B(n10266), .Z(n10029) );
  XOR2_X1 U10304 ( .A(n10267), .B(n10268), .Z(n10265) );
  XNOR2_X1 U10305 ( .A(n10269), .B(n10270), .ZN(n10033) );
  XOR2_X1 U10306 ( .A(n10271), .B(n10272), .Z(n10270) );
  NAND2_X1 U10307 ( .A1(b_20_), .A2(a_12_), .ZN(n10272) );
  XOR2_X1 U10308 ( .A(n10273), .B(n10274), .Z(n10036) );
  XOR2_X1 U10309 ( .A(n10275), .B(n10276), .Z(n10273) );
  NOR2_X1 U10310 ( .A1(n7424), .A2(n9966), .ZN(n10276) );
  XNOR2_X1 U10311 ( .A(n10277), .B(n10278), .ZN(n10040) );
  XNOR2_X1 U10312 ( .A(n10279), .B(n10280), .ZN(n10277) );
  XOR2_X1 U10313 ( .A(n10281), .B(n10282), .Z(n10045) );
  XOR2_X1 U10314 ( .A(n10283), .B(n10284), .Z(n10281) );
  XNOR2_X1 U10315 ( .A(n10285), .B(n10286), .ZN(n10049) );
  XNOR2_X1 U10316 ( .A(n10287), .B(n10288), .ZN(n10286) );
  XNOR2_X1 U10317 ( .A(n10289), .B(n10290), .ZN(n10053) );
  XOR2_X1 U10318 ( .A(n10291), .B(n10292), .Z(n10290) );
  NAND2_X1 U10319 ( .A1(b_20_), .A2(a_7_), .ZN(n10292) );
  XNOR2_X1 U10320 ( .A(n10293), .B(n10294), .ZN(n9862) );
  NAND2_X1 U10321 ( .A1(n10295), .A2(n10296), .ZN(n10293) );
  XNOR2_X1 U10322 ( .A(n10297), .B(n10298), .ZN(n10056) );
  NAND2_X1 U10323 ( .A1(n10299), .A2(n10300), .ZN(n10297) );
  XNOR2_X1 U10324 ( .A(n10301), .B(n10302), .ZN(n10061) );
  XNOR2_X1 U10325 ( .A(n10303), .B(n10304), .ZN(n10301) );
  XNOR2_X1 U10326 ( .A(n10305), .B(n10306), .ZN(n10065) );
  XOR2_X1 U10327 ( .A(n10307), .B(n10308), .Z(n10306) );
  NAND2_X1 U10328 ( .A1(b_20_), .A2(a_3_), .ZN(n10308) );
  XNOR2_X1 U10329 ( .A(n10309), .B(n10310), .ZN(n10069) );
  NAND2_X1 U10330 ( .A1(n10311), .A2(n10312), .ZN(n10309) );
  XOR2_X1 U10331 ( .A(n10313), .B(n10314), .Z(n10073) );
  XNOR2_X1 U10332 ( .A(n10315), .B(n10316), .ZN(n10313) );
  XOR2_X1 U10333 ( .A(n10317), .B(n10078), .Z(n10083) );
  XNOR2_X1 U10334 ( .A(n10318), .B(n10319), .ZN(n10078) );
  NOR2_X1 U10335 ( .A1(n7478), .A2(n9966), .ZN(n10319) );
  INV_X1 U10336 ( .A(n10079), .ZN(n10317) );
  NAND2_X1 U10337 ( .A1(n10320), .A2(n10321), .ZN(n7536) );
  XOR2_X1 U10338 ( .A(n7611), .B(n7610), .Z(n10321) );
  AND2_X1 U10339 ( .A1(n7618), .A2(n7617), .ZN(n10320) );
  XOR2_X1 U10340 ( .A(n10322), .B(n10323), .Z(n7617) );
  XOR2_X1 U10341 ( .A(n10324), .B(n10325), .Z(n10322) );
  NOR2_X1 U10342 ( .A1(n7478), .A2(n10207), .ZN(n10325) );
  NAND2_X1 U10343 ( .A1(n10326), .A2(n10327), .ZN(n7618) );
  NAND2_X1 U10344 ( .A1(n10328), .A2(b_20_), .ZN(n10327) );
  NOR2_X1 U10345 ( .A1(n10329), .A2(n7478), .ZN(n10328) );
  NOR2_X1 U10346 ( .A1(n10079), .A2(n10318), .ZN(n10329) );
  NAND2_X1 U10347 ( .A1(n10079), .A2(n10318), .ZN(n10326) );
  NAND2_X1 U10348 ( .A1(n10330), .A2(n10331), .ZN(n10318) );
  NAND2_X1 U10349 ( .A1(n10316), .A2(n10332), .ZN(n10331) );
  NAND2_X1 U10350 ( .A1(n10315), .A2(n10314), .ZN(n10332) );
  NOR2_X1 U10351 ( .A1(n9966), .A2(n7669), .ZN(n10316) );
  OR2_X1 U10352 ( .A1(n10314), .A2(n10315), .ZN(n10330) );
  AND2_X1 U10353 ( .A1(n10311), .A2(n10333), .ZN(n10315) );
  NAND2_X1 U10354 ( .A1(n10310), .A2(n10312), .ZN(n10333) );
  NAND2_X1 U10355 ( .A1(n10334), .A2(n10335), .ZN(n10312) );
  NAND2_X1 U10356 ( .A1(b_20_), .A2(a_2_), .ZN(n10335) );
  INV_X1 U10357 ( .A(n10336), .ZN(n10334) );
  XOR2_X1 U10358 ( .A(n10337), .B(n10338), .Z(n10310) );
  XOR2_X1 U10359 ( .A(n10339), .B(n10340), .Z(n10337) );
  NOR2_X1 U10360 ( .A1(n7464), .A2(n10207), .ZN(n10340) );
  NAND2_X1 U10361 ( .A1(a_2_), .A2(n10336), .ZN(n10311) );
  NAND2_X1 U10362 ( .A1(n10341), .A2(n10342), .ZN(n10336) );
  NAND2_X1 U10363 ( .A1(n10343), .A2(b_20_), .ZN(n10342) );
  NOR2_X1 U10364 ( .A1(n10344), .A2(n7464), .ZN(n10343) );
  NOR2_X1 U10365 ( .A1(n10305), .A2(n10307), .ZN(n10344) );
  NAND2_X1 U10366 ( .A1(n10305), .A2(n10307), .ZN(n10341) );
  NAND2_X1 U10367 ( .A1(n10345), .A2(n10346), .ZN(n10307) );
  NAND2_X1 U10368 ( .A1(n10304), .A2(n10347), .ZN(n10346) );
  NAND2_X1 U10369 ( .A1(n10303), .A2(n10302), .ZN(n10347) );
  NOR2_X1 U10370 ( .A1(n9966), .A2(n7682), .ZN(n10304) );
  OR2_X1 U10371 ( .A1(n10302), .A2(n10303), .ZN(n10345) );
  AND2_X1 U10372 ( .A1(n10299), .A2(n10348), .ZN(n10303) );
  NAND2_X1 U10373 ( .A1(n10298), .A2(n10300), .ZN(n10348) );
  NAND2_X1 U10374 ( .A1(n10349), .A2(n10350), .ZN(n10300) );
  NAND2_X1 U10375 ( .A1(b_20_), .A2(a_5_), .ZN(n10350) );
  INV_X1 U10376 ( .A(n10351), .ZN(n10349) );
  XOR2_X1 U10377 ( .A(n10352), .B(n10353), .Z(n10298) );
  XOR2_X1 U10378 ( .A(n10354), .B(n10355), .Z(n10352) );
  NOR2_X1 U10379 ( .A1(n7450), .A2(n10207), .ZN(n10355) );
  NAND2_X1 U10380 ( .A1(a_5_), .A2(n10351), .ZN(n10299) );
  NAND2_X1 U10381 ( .A1(n10295), .A2(n10356), .ZN(n10351) );
  NAND2_X1 U10382 ( .A1(n10294), .A2(n10296), .ZN(n10356) );
  NAND2_X1 U10383 ( .A1(n10357), .A2(n10358), .ZN(n10296) );
  NAND2_X1 U10384 ( .A1(b_20_), .A2(a_6_), .ZN(n10358) );
  INV_X1 U10385 ( .A(n10359), .ZN(n10357) );
  XOR2_X1 U10386 ( .A(n10360), .B(n10361), .Z(n10294) );
  XOR2_X1 U10387 ( .A(n10362), .B(n10363), .Z(n10360) );
  NOR2_X1 U10388 ( .A1(n7445), .A2(n10207), .ZN(n10363) );
  NAND2_X1 U10389 ( .A1(a_6_), .A2(n10359), .ZN(n10295) );
  NAND2_X1 U10390 ( .A1(n10364), .A2(n10365), .ZN(n10359) );
  NAND2_X1 U10391 ( .A1(n10366), .A2(b_20_), .ZN(n10365) );
  NOR2_X1 U10392 ( .A1(n10367), .A2(n7445), .ZN(n10366) );
  NOR2_X1 U10393 ( .A1(n10289), .A2(n10291), .ZN(n10367) );
  NAND2_X1 U10394 ( .A1(n10289), .A2(n10291), .ZN(n10364) );
  NAND2_X1 U10395 ( .A1(n10368), .A2(n10369), .ZN(n10291) );
  NAND2_X1 U10396 ( .A1(n10288), .A2(n10370), .ZN(n10369) );
  OR2_X1 U10397 ( .A1(n10287), .A2(n10285), .ZN(n10370) );
  NOR2_X1 U10398 ( .A1(n9966), .A2(n7699), .ZN(n10288) );
  NAND2_X1 U10399 ( .A1(n10285), .A2(n10287), .ZN(n10368) );
  NAND2_X1 U10400 ( .A1(n10371), .A2(n10372), .ZN(n10287) );
  NAND2_X1 U10401 ( .A1(n10284), .A2(n10373), .ZN(n10372) );
  OR2_X1 U10402 ( .A1(n10283), .A2(n10282), .ZN(n10373) );
  NOR2_X1 U10403 ( .A1(n9966), .A2(n7704), .ZN(n10284) );
  NAND2_X1 U10404 ( .A1(n10282), .A2(n10283), .ZN(n10371) );
  NAND2_X1 U10405 ( .A1(n10374), .A2(n10375), .ZN(n10283) );
  NAND2_X1 U10406 ( .A1(n10280), .A2(n10376), .ZN(n10375) );
  NAND2_X1 U10407 ( .A1(n10279), .A2(n10278), .ZN(n10376) );
  NOR2_X1 U10408 ( .A1(n9966), .A2(n7709), .ZN(n10280) );
  OR2_X1 U10409 ( .A1(n10278), .A2(n10279), .ZN(n10374) );
  AND2_X1 U10410 ( .A1(n10377), .A2(n10378), .ZN(n10279) );
  NAND2_X1 U10411 ( .A1(n10379), .A2(b_20_), .ZN(n10378) );
  NOR2_X1 U10412 ( .A1(n10380), .A2(n7424), .ZN(n10379) );
  NOR2_X1 U10413 ( .A1(n10274), .A2(n10275), .ZN(n10380) );
  NAND2_X1 U10414 ( .A1(n10274), .A2(n10275), .ZN(n10377) );
  NAND2_X1 U10415 ( .A1(n10381), .A2(n10382), .ZN(n10275) );
  NAND2_X1 U10416 ( .A1(n10383), .A2(b_20_), .ZN(n10382) );
  NOR2_X1 U10417 ( .A1(n10384), .A2(n7718), .ZN(n10383) );
  NOR2_X1 U10418 ( .A1(n10269), .A2(n10271), .ZN(n10384) );
  NAND2_X1 U10419 ( .A1(n10269), .A2(n10271), .ZN(n10381) );
  NAND2_X1 U10420 ( .A1(n10385), .A2(n10386), .ZN(n10271) );
  NAND2_X1 U10421 ( .A1(n10268), .A2(n10387), .ZN(n10386) );
  OR2_X1 U10422 ( .A1(n10267), .A2(n10266), .ZN(n10387) );
  NOR2_X1 U10423 ( .A1(n9966), .A2(n7415), .ZN(n10268) );
  NAND2_X1 U10424 ( .A1(n10266), .A2(n10267), .ZN(n10385) );
  NAND2_X1 U10425 ( .A1(n10388), .A2(n10389), .ZN(n10267) );
  NAND2_X1 U10426 ( .A1(n10390), .A2(b_20_), .ZN(n10389) );
  NOR2_X1 U10427 ( .A1(n10391), .A2(n7727), .ZN(n10390) );
  NOR2_X1 U10428 ( .A1(n10262), .A2(n10263), .ZN(n10391) );
  NAND2_X1 U10429 ( .A1(n10262), .A2(n10263), .ZN(n10388) );
  NAND2_X1 U10430 ( .A1(n10392), .A2(n10393), .ZN(n10263) );
  NAND2_X1 U10431 ( .A1(n10260), .A2(n10394), .ZN(n10393) );
  OR2_X1 U10432 ( .A1(n10259), .A2(n10258), .ZN(n10394) );
  NOR2_X1 U10433 ( .A1(n9966), .A2(n7406), .ZN(n10260) );
  NAND2_X1 U10434 ( .A1(n10258), .A2(n10259), .ZN(n10392) );
  NAND2_X1 U10435 ( .A1(n10395), .A2(n10396), .ZN(n10259) );
  NAND2_X1 U10436 ( .A1(n10397), .A2(b_20_), .ZN(n10396) );
  NOR2_X1 U10437 ( .A1(n10398), .A2(n7736), .ZN(n10397) );
  NOR2_X1 U10438 ( .A1(n10253), .A2(n10255), .ZN(n10398) );
  NAND2_X1 U10439 ( .A1(n10253), .A2(n10255), .ZN(n10395) );
  NAND2_X1 U10440 ( .A1(n10399), .A2(n10400), .ZN(n10255) );
  NAND2_X1 U10441 ( .A1(n10252), .A2(n10401), .ZN(n10400) );
  OR2_X1 U10442 ( .A1(n10251), .A2(n10250), .ZN(n10401) );
  NOR2_X1 U10443 ( .A1(n9966), .A2(n7397), .ZN(n10252) );
  NAND2_X1 U10444 ( .A1(n10250), .A2(n10251), .ZN(n10399) );
  NAND2_X1 U10445 ( .A1(n10402), .A2(n10403), .ZN(n10251) );
  NAND2_X1 U10446 ( .A1(n10404), .A2(b_20_), .ZN(n10403) );
  NOR2_X1 U10447 ( .A1(n10405), .A2(n7745), .ZN(n10404) );
  NOR2_X1 U10448 ( .A1(n10246), .A2(n10247), .ZN(n10405) );
  NAND2_X1 U10449 ( .A1(n10246), .A2(n10247), .ZN(n10402) );
  NAND2_X1 U10450 ( .A1(n10406), .A2(n10407), .ZN(n10247) );
  NAND2_X1 U10451 ( .A1(n10244), .A2(n10408), .ZN(n10407) );
  OR2_X1 U10452 ( .A1(n10243), .A2(n10242), .ZN(n10408) );
  NOR2_X1 U10453 ( .A1(n9966), .A2(n7750), .ZN(n10244) );
  NAND2_X1 U10454 ( .A1(n10242), .A2(n10243), .ZN(n10406) );
  NAND2_X1 U10455 ( .A1(n10409), .A2(n10410), .ZN(n10243) );
  NAND2_X1 U10456 ( .A1(n10240), .A2(n10411), .ZN(n10410) );
  OR2_X1 U10457 ( .A1(n10239), .A2(n10238), .ZN(n10411) );
  INV_X1 U10458 ( .A(n10412), .ZN(n10240) );
  NAND2_X1 U10459 ( .A1(n10238), .A2(n10239), .ZN(n10409) );
  NAND2_X1 U10460 ( .A1(n10413), .A2(n10414), .ZN(n10239) );
  NAND2_X1 U10461 ( .A1(n10236), .A2(n10415), .ZN(n10414) );
  OR2_X1 U10462 ( .A1(n10235), .A2(n10234), .ZN(n10415) );
  NOR2_X1 U10463 ( .A1(n9966), .A2(n7760), .ZN(n10236) );
  NAND2_X1 U10464 ( .A1(n10234), .A2(n10235), .ZN(n10413) );
  NAND2_X1 U10465 ( .A1(n10416), .A2(n10417), .ZN(n10235) );
  NAND2_X1 U10466 ( .A1(n10418), .A2(b_20_), .ZN(n10417) );
  NOR2_X1 U10467 ( .A1(n10419), .A2(n7765), .ZN(n10418) );
  NOR2_X1 U10468 ( .A1(n10229), .A2(n10231), .ZN(n10419) );
  NAND2_X1 U10469 ( .A1(n10229), .A2(n10231), .ZN(n10416) );
  NAND2_X1 U10470 ( .A1(n10420), .A2(n10421), .ZN(n10231) );
  NAND2_X1 U10471 ( .A1(n10228), .A2(n10422), .ZN(n10421) );
  OR2_X1 U10472 ( .A1(n10227), .A2(n10226), .ZN(n10422) );
  NOR2_X1 U10473 ( .A1(n9966), .A2(n8014), .ZN(n10228) );
  NAND2_X1 U10474 ( .A1(n10226), .A2(n10227), .ZN(n10420) );
  NAND2_X1 U10475 ( .A1(n10423), .A2(n10424), .ZN(n10227) );
  NAND2_X1 U10476 ( .A1(n10425), .A2(b_20_), .ZN(n10424) );
  NOR2_X1 U10477 ( .A1(n10426), .A2(n7774), .ZN(n10425) );
  NOR2_X1 U10478 ( .A1(n10222), .A2(n10224), .ZN(n10426) );
  NAND2_X1 U10479 ( .A1(n10222), .A2(n10224), .ZN(n10423) );
  NAND2_X1 U10480 ( .A1(n10427), .A2(n10428), .ZN(n10224) );
  NAND2_X1 U10481 ( .A1(n10220), .A2(n10429), .ZN(n10428) );
  OR2_X1 U10482 ( .A1(n10219), .A2(n10218), .ZN(n10429) );
  NOR2_X1 U10483 ( .A1(n9966), .A2(n8022), .ZN(n10220) );
  NAND2_X1 U10484 ( .A1(n10218), .A2(n10219), .ZN(n10427) );
  NAND2_X1 U10485 ( .A1(n10215), .A2(n10430), .ZN(n10219) );
  NAND2_X1 U10486 ( .A1(n10214), .A2(n10216), .ZN(n10430) );
  NAND2_X1 U10487 ( .A1(n10431), .A2(n10432), .ZN(n10216) );
  NAND2_X1 U10488 ( .A1(b_20_), .A2(a_26_), .ZN(n10432) );
  INV_X1 U10489 ( .A(n10433), .ZN(n10431) );
  XNOR2_X1 U10490 ( .A(n10434), .B(n10435), .ZN(n10214) );
  NAND2_X1 U10491 ( .A1(n10436), .A2(n10437), .ZN(n10434) );
  NAND2_X1 U10492 ( .A1(a_26_), .A2(n10433), .ZN(n10215) );
  NAND2_X1 U10493 ( .A1(n10184), .A2(n10438), .ZN(n10433) );
  NAND2_X1 U10494 ( .A1(n10183), .A2(n10185), .ZN(n10438) );
  NAND2_X1 U10495 ( .A1(n10439), .A2(n10440), .ZN(n10185) );
  NAND2_X1 U10496 ( .A1(b_20_), .A2(a_27_), .ZN(n10440) );
  INV_X1 U10497 ( .A(n10441), .ZN(n10439) );
  XNOR2_X1 U10498 ( .A(n10442), .B(n10443), .ZN(n10183) );
  XOR2_X1 U10499 ( .A(n10444), .B(n10445), .Z(n10443) );
  NAND2_X1 U10500 ( .A1(b_19_), .A2(a_28_), .ZN(n10445) );
  NAND2_X1 U10501 ( .A1(a_27_), .A2(n10441), .ZN(n10184) );
  NAND2_X1 U10502 ( .A1(n10446), .A2(n10447), .ZN(n10441) );
  NAND2_X1 U10503 ( .A1(n10448), .A2(b_20_), .ZN(n10447) );
  NOR2_X1 U10504 ( .A1(n10449), .A2(n7803), .ZN(n10448) );
  NOR2_X1 U10505 ( .A1(n10190), .A2(n10192), .ZN(n10449) );
  NAND2_X1 U10506 ( .A1(n10190), .A2(n10192), .ZN(n10446) );
  NAND2_X1 U10507 ( .A1(n10450), .A2(n10451), .ZN(n10192) );
  NAND2_X1 U10508 ( .A1(n10210), .A2(n10452), .ZN(n10451) );
  NAND2_X1 U10509 ( .A1(n10212), .A2(n10211), .ZN(n10452) );
  NOR2_X1 U10510 ( .A1(n9966), .A2(n7337), .ZN(n10210) );
  OR2_X1 U10511 ( .A1(n10211), .A2(n10212), .ZN(n10450) );
  AND2_X1 U10512 ( .A1(n10453), .A2(n10454), .ZN(n10212) );
  NAND2_X1 U10513 ( .A1(n10455), .A2(b_18_), .ZN(n10454) );
  NOR2_X1 U10514 ( .A1(n10456), .A2(n7817), .ZN(n10455) );
  NOR2_X1 U10515 ( .A1(n7816), .A2(n10207), .ZN(n10456) );
  NAND2_X1 U10516 ( .A1(n10457), .A2(b_19_), .ZN(n10453) );
  NOR2_X1 U10517 ( .A1(n10458), .A2(n8052), .ZN(n10457) );
  NOR2_X1 U10518 ( .A1(n7810), .A2(n10459), .ZN(n10458) );
  NAND2_X1 U10519 ( .A1(n10460), .A2(b_20_), .ZN(n10211) );
  XOR2_X1 U10520 ( .A(n10461), .B(n10462), .Z(n10190) );
  XOR2_X1 U10521 ( .A(n10463), .B(n10464), .Z(n10461) );
  XNOR2_X1 U10522 ( .A(n10465), .B(n10466), .ZN(n10218) );
  NAND2_X1 U10523 ( .A1(n10467), .A2(n10468), .ZN(n10465) );
  XOR2_X1 U10524 ( .A(n10469), .B(n10470), .Z(n10222) );
  XOR2_X1 U10525 ( .A(n10471), .B(n10472), .Z(n10469) );
  XOR2_X1 U10526 ( .A(n10473), .B(n10474), .Z(n10226) );
  XNOR2_X1 U10527 ( .A(n10475), .B(n10476), .ZN(n10473) );
  NAND2_X1 U10528 ( .A1(b_19_), .A2(a_24_), .ZN(n10475) );
  XOR2_X1 U10529 ( .A(n10477), .B(n10478), .Z(n10229) );
  XOR2_X1 U10530 ( .A(n10479), .B(n10480), .Z(n10477) );
  XNOR2_X1 U10531 ( .A(n10481), .B(n10482), .ZN(n10234) );
  XOR2_X1 U10532 ( .A(n10483), .B(n10484), .Z(n10482) );
  NAND2_X1 U10533 ( .A1(b_19_), .A2(a_22_), .ZN(n10484) );
  XNOR2_X1 U10534 ( .A(n10485), .B(n10486), .ZN(n10238) );
  XNOR2_X1 U10535 ( .A(n10487), .B(n10488), .ZN(n10485) );
  XOR2_X1 U10536 ( .A(n10489), .B(n10490), .Z(n10242) );
  XOR2_X1 U10537 ( .A(n10491), .B(n10492), .Z(n10489) );
  NOR2_X1 U10538 ( .A1(n7755), .A2(n10207), .ZN(n10492) );
  XOR2_X1 U10539 ( .A(n10493), .B(n10494), .Z(n10246) );
  XOR2_X1 U10540 ( .A(n10495), .B(n10496), .Z(n10493) );
  XNOR2_X1 U10541 ( .A(n10497), .B(n10498), .ZN(n10250) );
  XOR2_X1 U10542 ( .A(n10499), .B(n10500), .Z(n10498) );
  NAND2_X1 U10543 ( .A1(b_19_), .A2(a_18_), .ZN(n10500) );
  XNOR2_X1 U10544 ( .A(n10501), .B(n10502), .ZN(n10253) );
  XNOR2_X1 U10545 ( .A(n10503), .B(n10504), .ZN(n10502) );
  XOR2_X1 U10546 ( .A(n10505), .B(n10506), .Z(n10258) );
  XOR2_X1 U10547 ( .A(n10507), .B(n10508), .Z(n10505) );
  NOR2_X1 U10548 ( .A1(n7736), .A2(n10207), .ZN(n10508) );
  XOR2_X1 U10549 ( .A(n10509), .B(n10510), .Z(n10262) );
  XOR2_X1 U10550 ( .A(n10511), .B(n10512), .Z(n10509) );
  XNOR2_X1 U10551 ( .A(n10513), .B(n10514), .ZN(n10266) );
  XOR2_X1 U10552 ( .A(n10515), .B(n10516), .Z(n10514) );
  NAND2_X1 U10553 ( .A1(b_19_), .A2(a_14_), .ZN(n10516) );
  XOR2_X1 U10554 ( .A(n10517), .B(n10518), .Z(n10269) );
  XOR2_X1 U10555 ( .A(n10519), .B(n10520), .Z(n10517) );
  XOR2_X1 U10556 ( .A(n10521), .B(n10522), .Z(n10274) );
  XOR2_X1 U10557 ( .A(n10523), .B(n10524), .Z(n10521) );
  XNOR2_X1 U10558 ( .A(n10525), .B(n10526), .ZN(n10278) );
  XOR2_X1 U10559 ( .A(n10527), .B(n10528), .Z(n10525) );
  NOR2_X1 U10560 ( .A1(n7424), .A2(n10207), .ZN(n10528) );
  XOR2_X1 U10561 ( .A(n10529), .B(n10530), .Z(n10282) );
  XOR2_X1 U10562 ( .A(n10531), .B(n10532), .Z(n10529) );
  NOR2_X1 U10563 ( .A1(n7709), .A2(n10207), .ZN(n10532) );
  XOR2_X1 U10564 ( .A(n10533), .B(n10534), .Z(n10285) );
  XOR2_X1 U10565 ( .A(n10535), .B(n10536), .Z(n10533) );
  NOR2_X1 U10566 ( .A1(n7704), .A2(n10207), .ZN(n10536) );
  XOR2_X1 U10567 ( .A(n10537), .B(n10538), .Z(n10289) );
  XOR2_X1 U10568 ( .A(n10539), .B(n10540), .Z(n10537) );
  NOR2_X1 U10569 ( .A1(n7699), .A2(n10207), .ZN(n10540) );
  XNOR2_X1 U10570 ( .A(n10541), .B(n10542), .ZN(n10302) );
  XOR2_X1 U10571 ( .A(n10543), .B(n10544), .Z(n10541) );
  NOR2_X1 U10572 ( .A1(n7455), .A2(n10207), .ZN(n10544) );
  XOR2_X1 U10573 ( .A(n10545), .B(n10546), .Z(n10305) );
  XOR2_X1 U10574 ( .A(n10547), .B(n10548), .Z(n10545) );
  NOR2_X1 U10575 ( .A1(n7682), .A2(n10207), .ZN(n10548) );
  XOR2_X1 U10576 ( .A(n10549), .B(n10550), .Z(n10314) );
  NAND2_X1 U10577 ( .A1(n10551), .A2(n10552), .ZN(n10549) );
  XOR2_X1 U10578 ( .A(n10553), .B(n10554), .Z(n10079) );
  XOR2_X1 U10579 ( .A(n10555), .B(n10556), .Z(n10553) );
  NOR2_X1 U10580 ( .A1(n7669), .A2(n10207), .ZN(n10556) );
  NAND2_X1 U10581 ( .A1(n10557), .A2(n10558), .ZN(n7539) );
  XOR2_X1 U10582 ( .A(n7613), .B(n10559), .Z(n10558) );
  AND2_X1 U10583 ( .A1(n7611), .A2(n7610), .ZN(n10557) );
  XNOR2_X1 U10584 ( .A(n10560), .B(n10561), .ZN(n7610) );
  NAND2_X1 U10585 ( .A1(n10562), .A2(n10563), .ZN(n10560) );
  NAND2_X1 U10586 ( .A1(n10564), .A2(n10565), .ZN(n7611) );
  NAND2_X1 U10587 ( .A1(n10566), .A2(b_19_), .ZN(n10565) );
  NOR2_X1 U10588 ( .A1(n10567), .A2(n7478), .ZN(n10566) );
  NOR2_X1 U10589 ( .A1(n10323), .A2(n10324), .ZN(n10567) );
  NAND2_X1 U10590 ( .A1(n10323), .A2(n10324), .ZN(n10564) );
  NAND2_X1 U10591 ( .A1(n10568), .A2(n10569), .ZN(n10324) );
  NAND2_X1 U10592 ( .A1(n10570), .A2(b_19_), .ZN(n10569) );
  NOR2_X1 U10593 ( .A1(n10571), .A2(n7669), .ZN(n10570) );
  NOR2_X1 U10594 ( .A1(n10554), .A2(n10555), .ZN(n10571) );
  NAND2_X1 U10595 ( .A1(n10554), .A2(n10555), .ZN(n10568) );
  NAND2_X1 U10596 ( .A1(n10551), .A2(n10572), .ZN(n10555) );
  NAND2_X1 U10597 ( .A1(n10550), .A2(n10552), .ZN(n10572) );
  NAND2_X1 U10598 ( .A1(n10573), .A2(n10574), .ZN(n10552) );
  NAND2_X1 U10599 ( .A1(b_19_), .A2(a_2_), .ZN(n10574) );
  INV_X1 U10600 ( .A(n10575), .ZN(n10573) );
  XNOR2_X1 U10601 ( .A(n10576), .B(n10577), .ZN(n10550) );
  NAND2_X1 U10602 ( .A1(n10578), .A2(n10579), .ZN(n10576) );
  NAND2_X1 U10603 ( .A1(a_2_), .A2(n10575), .ZN(n10551) );
  NAND2_X1 U10604 ( .A1(n10580), .A2(n10581), .ZN(n10575) );
  NAND2_X1 U10605 ( .A1(n10582), .A2(b_19_), .ZN(n10581) );
  NOR2_X1 U10606 ( .A1(n10583), .A2(n7464), .ZN(n10582) );
  NOR2_X1 U10607 ( .A1(n10338), .A2(n10339), .ZN(n10583) );
  NAND2_X1 U10608 ( .A1(n10338), .A2(n10339), .ZN(n10580) );
  NAND2_X1 U10609 ( .A1(n10584), .A2(n10585), .ZN(n10339) );
  NAND2_X1 U10610 ( .A1(n10586), .A2(b_19_), .ZN(n10585) );
  NOR2_X1 U10611 ( .A1(n10587), .A2(n7682), .ZN(n10586) );
  NOR2_X1 U10612 ( .A1(n10546), .A2(n10547), .ZN(n10587) );
  NAND2_X1 U10613 ( .A1(n10546), .A2(n10547), .ZN(n10584) );
  NAND2_X1 U10614 ( .A1(n10588), .A2(n10589), .ZN(n10547) );
  NAND2_X1 U10615 ( .A1(n10590), .A2(b_19_), .ZN(n10589) );
  NOR2_X1 U10616 ( .A1(n10591), .A2(n7455), .ZN(n10590) );
  NOR2_X1 U10617 ( .A1(n10542), .A2(n10543), .ZN(n10591) );
  NAND2_X1 U10618 ( .A1(n10542), .A2(n10543), .ZN(n10588) );
  NAND2_X1 U10619 ( .A1(n10592), .A2(n10593), .ZN(n10543) );
  NAND2_X1 U10620 ( .A1(n10594), .A2(b_19_), .ZN(n10593) );
  NOR2_X1 U10621 ( .A1(n10595), .A2(n7450), .ZN(n10594) );
  NOR2_X1 U10622 ( .A1(n10353), .A2(n10354), .ZN(n10595) );
  NAND2_X1 U10623 ( .A1(n10353), .A2(n10354), .ZN(n10592) );
  NAND2_X1 U10624 ( .A1(n10596), .A2(n10597), .ZN(n10354) );
  NAND2_X1 U10625 ( .A1(n10598), .A2(b_19_), .ZN(n10597) );
  NOR2_X1 U10626 ( .A1(n10599), .A2(n7445), .ZN(n10598) );
  NOR2_X1 U10627 ( .A1(n10361), .A2(n10362), .ZN(n10599) );
  NAND2_X1 U10628 ( .A1(n10361), .A2(n10362), .ZN(n10596) );
  NAND2_X1 U10629 ( .A1(n10600), .A2(n10601), .ZN(n10362) );
  NAND2_X1 U10630 ( .A1(n10602), .A2(b_19_), .ZN(n10601) );
  NOR2_X1 U10631 ( .A1(n10603), .A2(n7699), .ZN(n10602) );
  NOR2_X1 U10632 ( .A1(n10538), .A2(n10539), .ZN(n10603) );
  NAND2_X1 U10633 ( .A1(n10538), .A2(n10539), .ZN(n10600) );
  NAND2_X1 U10634 ( .A1(n10604), .A2(n10605), .ZN(n10539) );
  NAND2_X1 U10635 ( .A1(n10606), .A2(b_19_), .ZN(n10605) );
  NOR2_X1 U10636 ( .A1(n10607), .A2(n7704), .ZN(n10606) );
  NOR2_X1 U10637 ( .A1(n10534), .A2(n10535), .ZN(n10607) );
  NAND2_X1 U10638 ( .A1(n10534), .A2(n10535), .ZN(n10604) );
  NAND2_X1 U10639 ( .A1(n10608), .A2(n10609), .ZN(n10535) );
  NAND2_X1 U10640 ( .A1(n10610), .A2(b_19_), .ZN(n10609) );
  NOR2_X1 U10641 ( .A1(n10611), .A2(n7709), .ZN(n10610) );
  NOR2_X1 U10642 ( .A1(n10530), .A2(n10531), .ZN(n10611) );
  NAND2_X1 U10643 ( .A1(n10530), .A2(n10531), .ZN(n10608) );
  NAND2_X1 U10644 ( .A1(n10612), .A2(n10613), .ZN(n10531) );
  NAND2_X1 U10645 ( .A1(n10614), .A2(b_19_), .ZN(n10613) );
  NOR2_X1 U10646 ( .A1(n10615), .A2(n7424), .ZN(n10614) );
  NOR2_X1 U10647 ( .A1(n10526), .A2(n10527), .ZN(n10615) );
  NAND2_X1 U10648 ( .A1(n10526), .A2(n10527), .ZN(n10612) );
  NAND2_X1 U10649 ( .A1(n10616), .A2(n10617), .ZN(n10527) );
  NAND2_X1 U10650 ( .A1(n10524), .A2(n10618), .ZN(n10617) );
  OR2_X1 U10651 ( .A1(n10523), .A2(n10522), .ZN(n10618) );
  NOR2_X1 U10652 ( .A1(n10207), .A2(n7718), .ZN(n10524) );
  NAND2_X1 U10653 ( .A1(n10522), .A2(n10523), .ZN(n10616) );
  NAND2_X1 U10654 ( .A1(n10619), .A2(n10620), .ZN(n10523) );
  NAND2_X1 U10655 ( .A1(n10520), .A2(n10621), .ZN(n10620) );
  OR2_X1 U10656 ( .A1(n10519), .A2(n10518), .ZN(n10621) );
  NOR2_X1 U10657 ( .A1(n10207), .A2(n7415), .ZN(n10520) );
  NAND2_X1 U10658 ( .A1(n10518), .A2(n10519), .ZN(n10619) );
  NAND2_X1 U10659 ( .A1(n10622), .A2(n10623), .ZN(n10519) );
  NAND2_X1 U10660 ( .A1(n10624), .A2(b_19_), .ZN(n10623) );
  NOR2_X1 U10661 ( .A1(n10625), .A2(n7727), .ZN(n10624) );
  NOR2_X1 U10662 ( .A1(n10513), .A2(n10515), .ZN(n10625) );
  NAND2_X1 U10663 ( .A1(n10513), .A2(n10515), .ZN(n10622) );
  NAND2_X1 U10664 ( .A1(n10626), .A2(n10627), .ZN(n10515) );
  NAND2_X1 U10665 ( .A1(n10512), .A2(n10628), .ZN(n10627) );
  OR2_X1 U10666 ( .A1(n10511), .A2(n10510), .ZN(n10628) );
  NOR2_X1 U10667 ( .A1(n10207), .A2(n7406), .ZN(n10512) );
  NAND2_X1 U10668 ( .A1(n10510), .A2(n10511), .ZN(n10626) );
  NAND2_X1 U10669 ( .A1(n10629), .A2(n10630), .ZN(n10511) );
  NAND2_X1 U10670 ( .A1(n10631), .A2(b_19_), .ZN(n10630) );
  NOR2_X1 U10671 ( .A1(n10632), .A2(n7736), .ZN(n10631) );
  NOR2_X1 U10672 ( .A1(n10506), .A2(n10507), .ZN(n10632) );
  NAND2_X1 U10673 ( .A1(n10506), .A2(n10507), .ZN(n10629) );
  NAND2_X1 U10674 ( .A1(n10633), .A2(n10634), .ZN(n10507) );
  NAND2_X1 U10675 ( .A1(n10504), .A2(n10635), .ZN(n10634) );
  OR2_X1 U10676 ( .A1(n10503), .A2(n10501), .ZN(n10635) );
  NOR2_X1 U10677 ( .A1(n10207), .A2(n7397), .ZN(n10504) );
  NAND2_X1 U10678 ( .A1(n10501), .A2(n10503), .ZN(n10633) );
  NAND2_X1 U10679 ( .A1(n10636), .A2(n10637), .ZN(n10503) );
  NAND2_X1 U10680 ( .A1(n10638), .A2(b_19_), .ZN(n10637) );
  NOR2_X1 U10681 ( .A1(n10639), .A2(n7745), .ZN(n10638) );
  NOR2_X1 U10682 ( .A1(n10497), .A2(n10499), .ZN(n10639) );
  NAND2_X1 U10683 ( .A1(n10497), .A2(n10499), .ZN(n10636) );
  NAND2_X1 U10684 ( .A1(n10640), .A2(n10641), .ZN(n10499) );
  NAND2_X1 U10685 ( .A1(n10496), .A2(n10642), .ZN(n10641) );
  OR2_X1 U10686 ( .A1(n10495), .A2(n10494), .ZN(n10642) );
  NAND2_X1 U10687 ( .A1(n10494), .A2(n10495), .ZN(n10640) );
  NAND2_X1 U10688 ( .A1(n10643), .A2(n10644), .ZN(n10495) );
  NAND2_X1 U10689 ( .A1(n10645), .A2(b_19_), .ZN(n10644) );
  NOR2_X1 U10690 ( .A1(n10646), .A2(n7755), .ZN(n10645) );
  NOR2_X1 U10691 ( .A1(n10490), .A2(n10491), .ZN(n10646) );
  NAND2_X1 U10692 ( .A1(n10490), .A2(n10491), .ZN(n10643) );
  NAND2_X1 U10693 ( .A1(n10647), .A2(n10648), .ZN(n10491) );
  NAND2_X1 U10694 ( .A1(n10488), .A2(n10649), .ZN(n10648) );
  NAND2_X1 U10695 ( .A1(n10487), .A2(n10486), .ZN(n10649) );
  NOR2_X1 U10696 ( .A1(n10207), .A2(n7760), .ZN(n10488) );
  OR2_X1 U10697 ( .A1(n10486), .A2(n10487), .ZN(n10647) );
  AND2_X1 U10698 ( .A1(n10650), .A2(n10651), .ZN(n10487) );
  NAND2_X1 U10699 ( .A1(n10652), .A2(b_19_), .ZN(n10651) );
  NOR2_X1 U10700 ( .A1(n10653), .A2(n7765), .ZN(n10652) );
  NOR2_X1 U10701 ( .A1(n10481), .A2(n10483), .ZN(n10653) );
  NAND2_X1 U10702 ( .A1(n10481), .A2(n10483), .ZN(n10650) );
  NAND2_X1 U10703 ( .A1(n10654), .A2(n10655), .ZN(n10483) );
  NAND2_X1 U10704 ( .A1(n10480), .A2(n10656), .ZN(n10655) );
  OR2_X1 U10705 ( .A1(n10479), .A2(n10478), .ZN(n10656) );
  NOR2_X1 U10706 ( .A1(n10207), .A2(n8014), .ZN(n10480) );
  NAND2_X1 U10707 ( .A1(n10478), .A2(n10479), .ZN(n10654) );
  NAND2_X1 U10708 ( .A1(n10657), .A2(n10658), .ZN(n10479) );
  NAND2_X1 U10709 ( .A1(n10659), .A2(b_19_), .ZN(n10658) );
  NOR2_X1 U10710 ( .A1(n10660), .A2(n7774), .ZN(n10659) );
  NOR2_X1 U10711 ( .A1(n10474), .A2(n10476), .ZN(n10660) );
  NAND2_X1 U10712 ( .A1(n10474), .A2(n10476), .ZN(n10657) );
  NAND2_X1 U10713 ( .A1(n10661), .A2(n10662), .ZN(n10476) );
  NAND2_X1 U10714 ( .A1(n10472), .A2(n10663), .ZN(n10662) );
  OR2_X1 U10715 ( .A1(n10471), .A2(n10470), .ZN(n10663) );
  NOR2_X1 U10716 ( .A1(n10207), .A2(n8022), .ZN(n10472) );
  NAND2_X1 U10717 ( .A1(n10470), .A2(n10471), .ZN(n10661) );
  NAND2_X1 U10718 ( .A1(n10467), .A2(n10664), .ZN(n10471) );
  NAND2_X1 U10719 ( .A1(n10466), .A2(n10468), .ZN(n10664) );
  NAND2_X1 U10720 ( .A1(n10665), .A2(n10666), .ZN(n10468) );
  NAND2_X1 U10721 ( .A1(b_19_), .A2(a_26_), .ZN(n10666) );
  INV_X1 U10722 ( .A(n10667), .ZN(n10665) );
  XNOR2_X1 U10723 ( .A(n10668), .B(n10669), .ZN(n10466) );
  NAND2_X1 U10724 ( .A1(n10670), .A2(n10671), .ZN(n10668) );
  NAND2_X1 U10725 ( .A1(a_26_), .A2(n10667), .ZN(n10467) );
  NAND2_X1 U10726 ( .A1(n10436), .A2(n10672), .ZN(n10667) );
  NAND2_X1 U10727 ( .A1(n10435), .A2(n10437), .ZN(n10672) );
  NAND2_X1 U10728 ( .A1(n10673), .A2(n10674), .ZN(n10437) );
  NAND2_X1 U10729 ( .A1(b_19_), .A2(a_27_), .ZN(n10674) );
  INV_X1 U10730 ( .A(n10675), .ZN(n10673) );
  XNOR2_X1 U10731 ( .A(n10676), .B(n10677), .ZN(n10435) );
  XOR2_X1 U10732 ( .A(n10678), .B(n10679), .Z(n10677) );
  NAND2_X1 U10733 ( .A1(b_18_), .A2(a_28_), .ZN(n10679) );
  NAND2_X1 U10734 ( .A1(a_27_), .A2(n10675), .ZN(n10436) );
  NAND2_X1 U10735 ( .A1(n10680), .A2(n10681), .ZN(n10675) );
  NAND2_X1 U10736 ( .A1(n10682), .A2(b_19_), .ZN(n10681) );
  NOR2_X1 U10737 ( .A1(n10683), .A2(n7803), .ZN(n10682) );
  NOR2_X1 U10738 ( .A1(n10442), .A2(n10444), .ZN(n10683) );
  NAND2_X1 U10739 ( .A1(n10442), .A2(n10444), .ZN(n10680) );
  NAND2_X1 U10740 ( .A1(n10684), .A2(n10685), .ZN(n10444) );
  NAND2_X1 U10741 ( .A1(n10462), .A2(n10686), .ZN(n10685) );
  NAND2_X1 U10742 ( .A1(n10464), .A2(n10463), .ZN(n10686) );
  NOR2_X1 U10743 ( .A1(n10207), .A2(n7337), .ZN(n10462) );
  OR2_X1 U10744 ( .A1(n10463), .A2(n10464), .ZN(n10684) );
  AND2_X1 U10745 ( .A1(n10687), .A2(n10688), .ZN(n10464) );
  NAND2_X1 U10746 ( .A1(n10689), .A2(b_17_), .ZN(n10688) );
  NOR2_X1 U10747 ( .A1(n10690), .A2(n7817), .ZN(n10689) );
  NOR2_X1 U10748 ( .A1(n7816), .A2(n10459), .ZN(n10690) );
  NAND2_X1 U10749 ( .A1(n10691), .A2(b_18_), .ZN(n10687) );
  NOR2_X1 U10750 ( .A1(n10692), .A2(n8052), .ZN(n10691) );
  NOR2_X1 U10751 ( .A1(n7810), .A2(n10693), .ZN(n10692) );
  NAND2_X1 U10752 ( .A1(n10460), .A2(b_18_), .ZN(n10463) );
  NOR2_X1 U10753 ( .A1(n8055), .A2(n10207), .ZN(n10460) );
  XOR2_X1 U10754 ( .A(n10694), .B(n10695), .Z(n10442) );
  XOR2_X1 U10755 ( .A(n10696), .B(n10697), .Z(n10694) );
  XNOR2_X1 U10756 ( .A(n10698), .B(n10699), .ZN(n10470) );
  NAND2_X1 U10757 ( .A1(n10700), .A2(n10701), .ZN(n10698) );
  XOR2_X1 U10758 ( .A(n10702), .B(n10703), .Z(n10474) );
  XOR2_X1 U10759 ( .A(n10704), .B(n10705), .Z(n10702) );
  XOR2_X1 U10760 ( .A(n10706), .B(n10707), .Z(n10478) );
  XOR2_X1 U10761 ( .A(n10708), .B(n10709), .Z(n10706) );
  NOR2_X1 U10762 ( .A1(n7774), .A2(n10459), .ZN(n10709) );
  XOR2_X1 U10763 ( .A(n10710), .B(n10711), .Z(n10481) );
  XOR2_X1 U10764 ( .A(n10712), .B(n10713), .Z(n10710) );
  NOR2_X1 U10765 ( .A1(n8014), .A2(n10459), .ZN(n10713) );
  XOR2_X1 U10766 ( .A(n10714), .B(n10715), .Z(n10486) );
  NAND2_X1 U10767 ( .A1(n10716), .A2(n10717), .ZN(n10714) );
  XOR2_X1 U10768 ( .A(n10718), .B(n10719), .Z(n10490) );
  XOR2_X1 U10769 ( .A(n10720), .B(n10721), .Z(n10718) );
  XNOR2_X1 U10770 ( .A(n10722), .B(n10723), .ZN(n10494) );
  XOR2_X1 U10771 ( .A(n10724), .B(n10725), .Z(n10723) );
  NAND2_X1 U10772 ( .A1(b_18_), .A2(a_20_), .ZN(n10725) );
  XOR2_X1 U10773 ( .A(n10726), .B(n10727), .Z(n10497) );
  XOR2_X1 U10774 ( .A(n10728), .B(n10729), .Z(n10726) );
  XNOR2_X1 U10775 ( .A(n10730), .B(n10731), .ZN(n10501) );
  XNOR2_X1 U10776 ( .A(n10732), .B(n10733), .ZN(n10730) );
  XNOR2_X1 U10777 ( .A(n10734), .B(n10735), .ZN(n10506) );
  XNOR2_X1 U10778 ( .A(n10736), .B(n10737), .ZN(n10735) );
  XNOR2_X1 U10779 ( .A(n10738), .B(n10739), .ZN(n10510) );
  XOR2_X1 U10780 ( .A(n10740), .B(n10741), .Z(n10739) );
  NAND2_X1 U10781 ( .A1(b_18_), .A2(a_16_), .ZN(n10741) );
  XOR2_X1 U10782 ( .A(n10742), .B(n10743), .Z(n10513) );
  XOR2_X1 U10783 ( .A(n10744), .B(n10745), .Z(n10742) );
  XOR2_X1 U10784 ( .A(n10746), .B(n10747), .Z(n10518) );
  XOR2_X1 U10785 ( .A(n10748), .B(n10749), .Z(n10746) );
  NOR2_X1 U10786 ( .A1(n7727), .A2(n10459), .ZN(n10749) );
  XOR2_X1 U10787 ( .A(n10750), .B(n10751), .Z(n10522) );
  XOR2_X1 U10788 ( .A(n10752), .B(n10753), .Z(n10750) );
  NOR2_X1 U10789 ( .A1(n7415), .A2(n10459), .ZN(n10753) );
  XNOR2_X1 U10790 ( .A(n10754), .B(n10755), .ZN(n10526) );
  XNOR2_X1 U10791 ( .A(n10756), .B(n10757), .ZN(n10754) );
  XOR2_X1 U10792 ( .A(n10758), .B(n10759), .Z(n10530) );
  XOR2_X1 U10793 ( .A(n10760), .B(n10761), .Z(n10758) );
  XNOR2_X1 U10794 ( .A(n10762), .B(n10763), .ZN(n10534) );
  XNOR2_X1 U10795 ( .A(n10764), .B(n10765), .ZN(n10763) );
  XNOR2_X1 U10796 ( .A(n10766), .B(n10767), .ZN(n10538) );
  XOR2_X1 U10797 ( .A(n10768), .B(n10769), .Z(n10767) );
  NAND2_X1 U10798 ( .A1(b_18_), .A2(a_9_), .ZN(n10769) );
  XNOR2_X1 U10799 ( .A(n10770), .B(n10771), .ZN(n10361) );
  NAND2_X1 U10800 ( .A1(n10772), .A2(n10773), .ZN(n10770) );
  XNOR2_X1 U10801 ( .A(n10774), .B(n10775), .ZN(n10353) );
  NAND2_X1 U10802 ( .A1(n10776), .A2(n10777), .ZN(n10774) );
  XNOR2_X1 U10803 ( .A(n10778), .B(n10779), .ZN(n10542) );
  XNOR2_X1 U10804 ( .A(n10780), .B(n10781), .ZN(n10778) );
  XOR2_X1 U10805 ( .A(n10782), .B(n10783), .Z(n10546) );
  XOR2_X1 U10806 ( .A(n10784), .B(n10785), .Z(n10782) );
  NOR2_X1 U10807 ( .A1(n7455), .A2(n10459), .ZN(n10785) );
  XNOR2_X1 U10808 ( .A(n10786), .B(n10787), .ZN(n10338) );
  NAND2_X1 U10809 ( .A1(n10788), .A2(n10789), .ZN(n10786) );
  XNOR2_X1 U10810 ( .A(n10790), .B(n10791), .ZN(n10554) );
  NAND2_X1 U10811 ( .A1(n10792), .A2(n10793), .ZN(n10790) );
  XOR2_X1 U10812 ( .A(n10794), .B(n10795), .Z(n10323) );
  NOR2_X1 U10813 ( .A1(n10796), .A2(n10797), .ZN(n10795) );
  NOR2_X1 U10814 ( .A1(n10798), .A2(n10799), .ZN(n10796) );
  NOR2_X1 U10815 ( .A1(n7669), .A2(n10459), .ZN(n10798) );
  NAND2_X1 U10816 ( .A1(n10800), .A2(n10801), .ZN(n7543) );
  NAND2_X1 U10817 ( .A1(n10802), .A2(n7612), .ZN(n10801) );
  INV_X1 U10818 ( .A(n7613), .ZN(n10802) );
  XOR2_X1 U10819 ( .A(n7603), .B(n10803), .Z(n10800) );
  NAND2_X1 U10820 ( .A1(n10804), .A2(n10805), .ZN(n7544) );
  XOR2_X1 U10821 ( .A(n7603), .B(n7602), .Z(n10805) );
  NOR2_X1 U10822 ( .A1(n10559), .A2(n7613), .ZN(n10804) );
  XNOR2_X1 U10823 ( .A(n10806), .B(n10807), .ZN(n7613) );
  XOR2_X1 U10824 ( .A(n10808), .B(n10809), .Z(n10806) );
  NOR2_X1 U10825 ( .A1(n7478), .A2(n10693), .ZN(n10809) );
  INV_X1 U10826 ( .A(n7612), .ZN(n10559) );
  NAND2_X1 U10827 ( .A1(n10562), .A2(n10810), .ZN(n7612) );
  NAND2_X1 U10828 ( .A1(n10561), .A2(n10563), .ZN(n10810) );
  NAND2_X1 U10829 ( .A1(n10811), .A2(n10812), .ZN(n10563) );
  NAND2_X1 U10830 ( .A1(b_18_), .A2(a_0_), .ZN(n10812) );
  XOR2_X1 U10831 ( .A(n10813), .B(n10814), .Z(n10561) );
  XOR2_X1 U10832 ( .A(n10815), .B(n10816), .Z(n10813) );
  NOR2_X1 U10833 ( .A1(n7669), .A2(n10693), .ZN(n10816) );
  OR2_X1 U10834 ( .A1(n7478), .A2(n10811), .ZN(n10562) );
  NOR2_X1 U10835 ( .A1(n10797), .A2(n10817), .ZN(n10811) );
  AND2_X1 U10836 ( .A1(n10794), .A2(n10818), .ZN(n10817) );
  NAND2_X1 U10837 ( .A1(n10819), .A2(n10820), .ZN(n10818) );
  NAND2_X1 U10838 ( .A1(b_18_), .A2(a_1_), .ZN(n10820) );
  XOR2_X1 U10839 ( .A(n10821), .B(n10822), .Z(n10794) );
  XOR2_X1 U10840 ( .A(n10823), .B(n10824), .Z(n10821) );
  NOR2_X1 U10841 ( .A1(n7469), .A2(n10693), .ZN(n10824) );
  NOR2_X1 U10842 ( .A1(n7669), .A2(n10819), .ZN(n10797) );
  INV_X1 U10843 ( .A(n10799), .ZN(n10819) );
  NAND2_X1 U10844 ( .A1(n10792), .A2(n10825), .ZN(n10799) );
  NAND2_X1 U10845 ( .A1(n10791), .A2(n10793), .ZN(n10825) );
  NAND2_X1 U10846 ( .A1(n10826), .A2(n10827), .ZN(n10793) );
  NAND2_X1 U10847 ( .A1(b_18_), .A2(a_2_), .ZN(n10827) );
  INV_X1 U10848 ( .A(n10828), .ZN(n10826) );
  XOR2_X1 U10849 ( .A(n10829), .B(n10830), .Z(n10791) );
  XOR2_X1 U10850 ( .A(n10831), .B(n10832), .Z(n10829) );
  NOR2_X1 U10851 ( .A1(n7464), .A2(n10693), .ZN(n10832) );
  NAND2_X1 U10852 ( .A1(a_2_), .A2(n10828), .ZN(n10792) );
  NAND2_X1 U10853 ( .A1(n10578), .A2(n10833), .ZN(n10828) );
  NAND2_X1 U10854 ( .A1(n10577), .A2(n10579), .ZN(n10833) );
  NAND2_X1 U10855 ( .A1(n10834), .A2(n10835), .ZN(n10579) );
  NAND2_X1 U10856 ( .A1(b_18_), .A2(a_3_), .ZN(n10835) );
  INV_X1 U10857 ( .A(n10836), .ZN(n10834) );
  XOR2_X1 U10858 ( .A(n10837), .B(n10838), .Z(n10577) );
  XOR2_X1 U10859 ( .A(n10839), .B(n10840), .Z(n10837) );
  NOR2_X1 U10860 ( .A1(n7682), .A2(n10693), .ZN(n10840) );
  NAND2_X1 U10861 ( .A1(a_3_), .A2(n10836), .ZN(n10578) );
  NAND2_X1 U10862 ( .A1(n10788), .A2(n10841), .ZN(n10836) );
  NAND2_X1 U10863 ( .A1(n10787), .A2(n10789), .ZN(n10841) );
  NAND2_X1 U10864 ( .A1(n10842), .A2(n10843), .ZN(n10789) );
  NAND2_X1 U10865 ( .A1(b_18_), .A2(a_4_), .ZN(n10843) );
  INV_X1 U10866 ( .A(n10844), .ZN(n10842) );
  XOR2_X1 U10867 ( .A(n10845), .B(n10846), .Z(n10787) );
  XOR2_X1 U10868 ( .A(n10847), .B(n10848), .Z(n10845) );
  NOR2_X1 U10869 ( .A1(n7455), .A2(n10693), .ZN(n10848) );
  NAND2_X1 U10870 ( .A1(a_4_), .A2(n10844), .ZN(n10788) );
  NAND2_X1 U10871 ( .A1(n10849), .A2(n10850), .ZN(n10844) );
  NAND2_X1 U10872 ( .A1(n10851), .A2(b_18_), .ZN(n10850) );
  NOR2_X1 U10873 ( .A1(n10852), .A2(n7455), .ZN(n10851) );
  NOR2_X1 U10874 ( .A1(n10783), .A2(n10784), .ZN(n10852) );
  NAND2_X1 U10875 ( .A1(n10783), .A2(n10784), .ZN(n10849) );
  NAND2_X1 U10876 ( .A1(n10853), .A2(n10854), .ZN(n10784) );
  NAND2_X1 U10877 ( .A1(n10781), .A2(n10855), .ZN(n10854) );
  NAND2_X1 U10878 ( .A1(n10780), .A2(n10779), .ZN(n10855) );
  NOR2_X1 U10879 ( .A1(n10459), .A2(n7450), .ZN(n10781) );
  OR2_X1 U10880 ( .A1(n10779), .A2(n10780), .ZN(n10853) );
  AND2_X1 U10881 ( .A1(n10776), .A2(n10856), .ZN(n10780) );
  NAND2_X1 U10882 ( .A1(n10775), .A2(n10777), .ZN(n10856) );
  NAND2_X1 U10883 ( .A1(n10857), .A2(n10858), .ZN(n10777) );
  NAND2_X1 U10884 ( .A1(b_18_), .A2(a_7_), .ZN(n10858) );
  INV_X1 U10885 ( .A(n10859), .ZN(n10857) );
  XOR2_X1 U10886 ( .A(n10860), .B(n10861), .Z(n10775) );
  XOR2_X1 U10887 ( .A(n10862), .B(n10863), .Z(n10860) );
  NOR2_X1 U10888 ( .A1(n7699), .A2(n10693), .ZN(n10863) );
  NAND2_X1 U10889 ( .A1(a_7_), .A2(n10859), .ZN(n10776) );
  NAND2_X1 U10890 ( .A1(n10772), .A2(n10864), .ZN(n10859) );
  NAND2_X1 U10891 ( .A1(n10771), .A2(n10773), .ZN(n10864) );
  NAND2_X1 U10892 ( .A1(n10865), .A2(n10866), .ZN(n10773) );
  NAND2_X1 U10893 ( .A1(b_18_), .A2(a_8_), .ZN(n10866) );
  INV_X1 U10894 ( .A(n10867), .ZN(n10865) );
  XOR2_X1 U10895 ( .A(n10868), .B(n10869), .Z(n10771) );
  XOR2_X1 U10896 ( .A(n10870), .B(n10871), .Z(n10868) );
  NOR2_X1 U10897 ( .A1(n7704), .A2(n10693), .ZN(n10871) );
  NAND2_X1 U10898 ( .A1(a_8_), .A2(n10867), .ZN(n10772) );
  NAND2_X1 U10899 ( .A1(n10872), .A2(n10873), .ZN(n10867) );
  NAND2_X1 U10900 ( .A1(n10874), .A2(b_18_), .ZN(n10873) );
  NOR2_X1 U10901 ( .A1(n10875), .A2(n7704), .ZN(n10874) );
  NOR2_X1 U10902 ( .A1(n10766), .A2(n10768), .ZN(n10875) );
  NAND2_X1 U10903 ( .A1(n10766), .A2(n10768), .ZN(n10872) );
  NAND2_X1 U10904 ( .A1(n10876), .A2(n10877), .ZN(n10768) );
  NAND2_X1 U10905 ( .A1(n10765), .A2(n10878), .ZN(n10877) );
  OR2_X1 U10906 ( .A1(n10764), .A2(n10762), .ZN(n10878) );
  NOR2_X1 U10907 ( .A1(n10459), .A2(n7709), .ZN(n10765) );
  NAND2_X1 U10908 ( .A1(n10762), .A2(n10764), .ZN(n10876) );
  NAND2_X1 U10909 ( .A1(n10879), .A2(n10880), .ZN(n10764) );
  NAND2_X1 U10910 ( .A1(n10761), .A2(n10881), .ZN(n10880) );
  OR2_X1 U10911 ( .A1(n10759), .A2(n10760), .ZN(n10881) );
  NOR2_X1 U10912 ( .A1(n10459), .A2(n7424), .ZN(n10761) );
  NAND2_X1 U10913 ( .A1(n10759), .A2(n10760), .ZN(n10879) );
  NAND2_X1 U10914 ( .A1(n10882), .A2(n10883), .ZN(n10760) );
  NAND2_X1 U10915 ( .A1(n10757), .A2(n10884), .ZN(n10883) );
  NAND2_X1 U10916 ( .A1(n10756), .A2(n10755), .ZN(n10884) );
  NOR2_X1 U10917 ( .A1(n10459), .A2(n7718), .ZN(n10757) );
  OR2_X1 U10918 ( .A1(n10755), .A2(n10756), .ZN(n10882) );
  AND2_X1 U10919 ( .A1(n10885), .A2(n10886), .ZN(n10756) );
  NAND2_X1 U10920 ( .A1(n10887), .A2(b_18_), .ZN(n10886) );
  NOR2_X1 U10921 ( .A1(n10888), .A2(n7415), .ZN(n10887) );
  NOR2_X1 U10922 ( .A1(n10751), .A2(n10752), .ZN(n10888) );
  NAND2_X1 U10923 ( .A1(n10751), .A2(n10752), .ZN(n10885) );
  NAND2_X1 U10924 ( .A1(n10889), .A2(n10890), .ZN(n10752) );
  NAND2_X1 U10925 ( .A1(n10891), .A2(b_18_), .ZN(n10890) );
  NOR2_X1 U10926 ( .A1(n10892), .A2(n7727), .ZN(n10891) );
  NOR2_X1 U10927 ( .A1(n10747), .A2(n10748), .ZN(n10892) );
  NAND2_X1 U10928 ( .A1(n10747), .A2(n10748), .ZN(n10889) );
  NAND2_X1 U10929 ( .A1(n10893), .A2(n10894), .ZN(n10748) );
  NAND2_X1 U10930 ( .A1(n10745), .A2(n10895), .ZN(n10894) );
  OR2_X1 U10931 ( .A1(n10743), .A2(n10744), .ZN(n10895) );
  NOR2_X1 U10932 ( .A1(n10459), .A2(n7406), .ZN(n10745) );
  NAND2_X1 U10933 ( .A1(n10743), .A2(n10744), .ZN(n10893) );
  NAND2_X1 U10934 ( .A1(n10896), .A2(n10897), .ZN(n10744) );
  NAND2_X1 U10935 ( .A1(n10898), .A2(b_18_), .ZN(n10897) );
  NOR2_X1 U10936 ( .A1(n10899), .A2(n7736), .ZN(n10898) );
  NOR2_X1 U10937 ( .A1(n10738), .A2(n10740), .ZN(n10899) );
  NAND2_X1 U10938 ( .A1(n10738), .A2(n10740), .ZN(n10896) );
  NAND2_X1 U10939 ( .A1(n10900), .A2(n10901), .ZN(n10740) );
  NAND2_X1 U10940 ( .A1(n10737), .A2(n10902), .ZN(n10901) );
  OR2_X1 U10941 ( .A1(n10734), .A2(n10736), .ZN(n10902) );
  NOR2_X1 U10942 ( .A1(n10459), .A2(n7397), .ZN(n10737) );
  NAND2_X1 U10943 ( .A1(n10734), .A2(n10736), .ZN(n10900) );
  NAND2_X1 U10944 ( .A1(n10903), .A2(n10904), .ZN(n10736) );
  NAND2_X1 U10945 ( .A1(n10733), .A2(n10905), .ZN(n10904) );
  NAND2_X1 U10946 ( .A1(n10732), .A2(n10731), .ZN(n10905) );
  OR2_X1 U10947 ( .A1(n10731), .A2(n10732), .ZN(n10903) );
  AND2_X1 U10948 ( .A1(n10906), .A2(n10907), .ZN(n10732) );
  NAND2_X1 U10949 ( .A1(n10729), .A2(n10908), .ZN(n10907) );
  OR2_X1 U10950 ( .A1(n10727), .A2(n10728), .ZN(n10908) );
  NOR2_X1 U10951 ( .A1(n10459), .A2(n7750), .ZN(n10729) );
  NAND2_X1 U10952 ( .A1(n10727), .A2(n10728), .ZN(n10906) );
  NAND2_X1 U10953 ( .A1(n10909), .A2(n10910), .ZN(n10728) );
  NAND2_X1 U10954 ( .A1(n10911), .A2(b_18_), .ZN(n10910) );
  NOR2_X1 U10955 ( .A1(n10912), .A2(n7755), .ZN(n10911) );
  NOR2_X1 U10956 ( .A1(n10722), .A2(n10724), .ZN(n10912) );
  NAND2_X1 U10957 ( .A1(n10722), .A2(n10724), .ZN(n10909) );
  NAND2_X1 U10958 ( .A1(n10913), .A2(n10914), .ZN(n10724) );
  NAND2_X1 U10959 ( .A1(n10721), .A2(n10915), .ZN(n10914) );
  OR2_X1 U10960 ( .A1(n10719), .A2(n10720), .ZN(n10915) );
  NOR2_X1 U10961 ( .A1(n10459), .A2(n7760), .ZN(n10721) );
  NAND2_X1 U10962 ( .A1(n10719), .A2(n10720), .ZN(n10913) );
  NAND2_X1 U10963 ( .A1(n10716), .A2(n10916), .ZN(n10720) );
  NAND2_X1 U10964 ( .A1(n10715), .A2(n10717), .ZN(n10916) );
  NAND2_X1 U10965 ( .A1(n10917), .A2(n10918), .ZN(n10717) );
  NAND2_X1 U10966 ( .A1(b_18_), .A2(a_22_), .ZN(n10918) );
  INV_X1 U10967 ( .A(n10919), .ZN(n10917) );
  XOR2_X1 U10968 ( .A(n10920), .B(n10921), .Z(n10715) );
  XOR2_X1 U10969 ( .A(n10922), .B(n10923), .Z(n10920) );
  NAND2_X1 U10970 ( .A1(a_22_), .A2(n10919), .ZN(n10716) );
  NAND2_X1 U10971 ( .A1(n10924), .A2(n10925), .ZN(n10919) );
  NAND2_X1 U10972 ( .A1(n10926), .A2(b_18_), .ZN(n10925) );
  NOR2_X1 U10973 ( .A1(n10927), .A2(n8014), .ZN(n10926) );
  NOR2_X1 U10974 ( .A1(n10712), .A2(n10711), .ZN(n10927) );
  NAND2_X1 U10975 ( .A1(n10711), .A2(n10712), .ZN(n10924) );
  NAND2_X1 U10976 ( .A1(n10928), .A2(n10929), .ZN(n10712) );
  NAND2_X1 U10977 ( .A1(n10930), .A2(b_18_), .ZN(n10929) );
  NOR2_X1 U10978 ( .A1(n10931), .A2(n7774), .ZN(n10930) );
  NOR2_X1 U10979 ( .A1(n10707), .A2(n10708), .ZN(n10931) );
  NAND2_X1 U10980 ( .A1(n10707), .A2(n10708), .ZN(n10928) );
  NAND2_X1 U10981 ( .A1(n10932), .A2(n10933), .ZN(n10708) );
  NAND2_X1 U10982 ( .A1(n10705), .A2(n10934), .ZN(n10933) );
  OR2_X1 U10983 ( .A1(n10703), .A2(n10704), .ZN(n10934) );
  NOR2_X1 U10984 ( .A1(n10459), .A2(n8022), .ZN(n10705) );
  NAND2_X1 U10985 ( .A1(n10703), .A2(n10704), .ZN(n10932) );
  NAND2_X1 U10986 ( .A1(n10700), .A2(n10935), .ZN(n10704) );
  NAND2_X1 U10987 ( .A1(n10699), .A2(n10701), .ZN(n10935) );
  NAND2_X1 U10988 ( .A1(n10936), .A2(n10937), .ZN(n10701) );
  NAND2_X1 U10989 ( .A1(b_18_), .A2(a_26_), .ZN(n10937) );
  INV_X1 U10990 ( .A(n10938), .ZN(n10936) );
  XNOR2_X1 U10991 ( .A(n10939), .B(n10940), .ZN(n10699) );
  NAND2_X1 U10992 ( .A1(n10941), .A2(n10942), .ZN(n10939) );
  NAND2_X1 U10993 ( .A1(a_26_), .A2(n10938), .ZN(n10700) );
  NAND2_X1 U10994 ( .A1(n10670), .A2(n10943), .ZN(n10938) );
  NAND2_X1 U10995 ( .A1(n10669), .A2(n10671), .ZN(n10943) );
  NAND2_X1 U10996 ( .A1(n10944), .A2(n10945), .ZN(n10671) );
  NAND2_X1 U10997 ( .A1(b_18_), .A2(a_27_), .ZN(n10945) );
  INV_X1 U10998 ( .A(n10946), .ZN(n10944) );
  XNOR2_X1 U10999 ( .A(n10947), .B(n10948), .ZN(n10669) );
  XOR2_X1 U11000 ( .A(n10949), .B(n10950), .Z(n10948) );
  NAND2_X1 U11001 ( .A1(b_17_), .A2(a_28_), .ZN(n10950) );
  NAND2_X1 U11002 ( .A1(a_27_), .A2(n10946), .ZN(n10670) );
  NAND2_X1 U11003 ( .A1(n10951), .A2(n10952), .ZN(n10946) );
  NAND2_X1 U11004 ( .A1(n10953), .A2(b_18_), .ZN(n10952) );
  NOR2_X1 U11005 ( .A1(n10954), .A2(n7803), .ZN(n10953) );
  NOR2_X1 U11006 ( .A1(n10676), .A2(n10678), .ZN(n10954) );
  NAND2_X1 U11007 ( .A1(n10676), .A2(n10678), .ZN(n10951) );
  NAND2_X1 U11008 ( .A1(n10955), .A2(n10956), .ZN(n10678) );
  NAND2_X1 U11009 ( .A1(n10695), .A2(n10957), .ZN(n10956) );
  NAND2_X1 U11010 ( .A1(n10697), .A2(n10696), .ZN(n10957) );
  NOR2_X1 U11011 ( .A1(n10459), .A2(n7337), .ZN(n10695) );
  OR2_X1 U11012 ( .A1(n10696), .A2(n10697), .ZN(n10955) );
  AND2_X1 U11013 ( .A1(n10958), .A2(n10959), .ZN(n10697) );
  NAND2_X1 U11014 ( .A1(n10960), .A2(b_16_), .ZN(n10959) );
  NOR2_X1 U11015 ( .A1(n10961), .A2(n7817), .ZN(n10960) );
  NOR2_X1 U11016 ( .A1(n7816), .A2(n10693), .ZN(n10961) );
  NAND2_X1 U11017 ( .A1(n10962), .A2(b_17_), .ZN(n10958) );
  NOR2_X1 U11018 ( .A1(n10963), .A2(n8052), .ZN(n10962) );
  NOR2_X1 U11019 ( .A1(n7810), .A2(n10964), .ZN(n10963) );
  NAND2_X1 U11020 ( .A1(n10965), .A2(b_18_), .ZN(n10696) );
  XOR2_X1 U11021 ( .A(n10966), .B(n10967), .Z(n10676) );
  XOR2_X1 U11022 ( .A(n10968), .B(n10969), .Z(n10966) );
  XNOR2_X1 U11023 ( .A(n10970), .B(n10971), .ZN(n10703) );
  NAND2_X1 U11024 ( .A1(n10972), .A2(n10973), .ZN(n10970) );
  XOR2_X1 U11025 ( .A(n10974), .B(n10975), .Z(n10707) );
  XOR2_X1 U11026 ( .A(n10976), .B(n10977), .Z(n10974) );
  XOR2_X1 U11027 ( .A(n10978), .B(n10979), .Z(n10711) );
  XNOR2_X1 U11028 ( .A(n10980), .B(n10981), .ZN(n10978) );
  NAND2_X1 U11029 ( .A1(b_17_), .A2(a_24_), .ZN(n10980) );
  XNOR2_X1 U11030 ( .A(n10982), .B(n10983), .ZN(n10719) );
  XOR2_X1 U11031 ( .A(n10984), .B(n10985), .Z(n10983) );
  NAND2_X1 U11032 ( .A1(b_17_), .A2(a_22_), .ZN(n10985) );
  XOR2_X1 U11033 ( .A(n10986), .B(n10987), .Z(n10722) );
  XOR2_X1 U11034 ( .A(n10988), .B(n10989), .Z(n10986) );
  XOR2_X1 U11035 ( .A(n10990), .B(n10991), .Z(n10727) );
  XOR2_X1 U11036 ( .A(n10992), .B(n10993), .Z(n10990) );
  NOR2_X1 U11037 ( .A1(n7755), .A2(n10693), .ZN(n10993) );
  XOR2_X1 U11038 ( .A(n10994), .B(n10995), .Z(n10731) );
  XNOR2_X1 U11039 ( .A(n10996), .B(n10997), .ZN(n10995) );
  XOR2_X1 U11040 ( .A(n10998), .B(n10999), .Z(n10734) );
  XOR2_X1 U11041 ( .A(n11000), .B(n11001), .Z(n10998) );
  NOR2_X1 U11042 ( .A1(n7745), .A2(n10693), .ZN(n11001) );
  XNOR2_X1 U11043 ( .A(n11002), .B(n11003), .ZN(n10738) );
  XNOR2_X1 U11044 ( .A(n11004), .B(n11005), .ZN(n11003) );
  XOR2_X1 U11045 ( .A(n11006), .B(n11007), .Z(n10743) );
  XOR2_X1 U11046 ( .A(n11008), .B(n11009), .Z(n11006) );
  NOR2_X1 U11047 ( .A1(n7736), .A2(n10693), .ZN(n11009) );
  XOR2_X1 U11048 ( .A(n11010), .B(n11011), .Z(n10747) );
  XOR2_X1 U11049 ( .A(n11012), .B(n11013), .Z(n11010) );
  XOR2_X1 U11050 ( .A(n11014), .B(n11015), .Z(n10751) );
  XOR2_X1 U11051 ( .A(n11016), .B(n11017), .Z(n11014) );
  XNOR2_X1 U11052 ( .A(n11018), .B(n11019), .ZN(n10755) );
  XOR2_X1 U11053 ( .A(n11020), .B(n11021), .Z(n11018) );
  NOR2_X1 U11054 ( .A1(n7415), .A2(n10693), .ZN(n11021) );
  XOR2_X1 U11055 ( .A(n11022), .B(n11023), .Z(n10759) );
  XOR2_X1 U11056 ( .A(n11024), .B(n11025), .Z(n11022) );
  NOR2_X1 U11057 ( .A1(n7718), .A2(n10693), .ZN(n11025) );
  XOR2_X1 U11058 ( .A(n11026), .B(n11027), .Z(n10762) );
  XOR2_X1 U11059 ( .A(n11028), .B(n11029), .Z(n11026) );
  NOR2_X1 U11060 ( .A1(n7424), .A2(n10693), .ZN(n11029) );
  XOR2_X1 U11061 ( .A(n11030), .B(n11031), .Z(n10766) );
  XOR2_X1 U11062 ( .A(n11032), .B(n11033), .Z(n11030) );
  NOR2_X1 U11063 ( .A1(n7709), .A2(n10693), .ZN(n11033) );
  XOR2_X1 U11064 ( .A(n11034), .B(n11035), .Z(n10779) );
  XOR2_X1 U11065 ( .A(n11036), .B(n11037), .Z(n11035) );
  NAND2_X1 U11066 ( .A1(b_17_), .A2(a_7_), .ZN(n11037) );
  XNOR2_X1 U11067 ( .A(n11038), .B(n11039), .ZN(n10783) );
  XOR2_X1 U11068 ( .A(n11040), .B(n11041), .Z(n11039) );
  NAND2_X1 U11069 ( .A1(b_17_), .A2(a_6_), .ZN(n11041) );
  NAND2_X1 U11070 ( .A1(n11042), .A2(n11043), .ZN(n7548) );
  XOR2_X1 U11071 ( .A(n7605), .B(n11044), .Z(n11043) );
  AND2_X1 U11072 ( .A1(n7603), .A2(n7602), .ZN(n11042) );
  INV_X1 U11073 ( .A(n10803), .ZN(n7602) );
  XOR2_X1 U11074 ( .A(n11045), .B(n11046), .Z(n10803) );
  NAND2_X1 U11075 ( .A1(n11047), .A2(n11048), .ZN(n11045) );
  NAND2_X1 U11076 ( .A1(n11049), .A2(n11050), .ZN(n7603) );
  NAND2_X1 U11077 ( .A1(n11051), .A2(b_17_), .ZN(n11050) );
  NOR2_X1 U11078 ( .A1(n11052), .A2(n7478), .ZN(n11051) );
  NOR2_X1 U11079 ( .A1(n10807), .A2(n10808), .ZN(n11052) );
  NAND2_X1 U11080 ( .A1(n10807), .A2(n10808), .ZN(n11049) );
  NAND2_X1 U11081 ( .A1(n11053), .A2(n11054), .ZN(n10808) );
  NAND2_X1 U11082 ( .A1(n11055), .A2(b_17_), .ZN(n11054) );
  NOR2_X1 U11083 ( .A1(n11056), .A2(n7669), .ZN(n11055) );
  NOR2_X1 U11084 ( .A1(n10814), .A2(n10815), .ZN(n11056) );
  NAND2_X1 U11085 ( .A1(n10814), .A2(n10815), .ZN(n11053) );
  NAND2_X1 U11086 ( .A1(n11057), .A2(n11058), .ZN(n10815) );
  NAND2_X1 U11087 ( .A1(n11059), .A2(b_17_), .ZN(n11058) );
  NOR2_X1 U11088 ( .A1(n11060), .A2(n7469), .ZN(n11059) );
  NOR2_X1 U11089 ( .A1(n10822), .A2(n10823), .ZN(n11060) );
  NAND2_X1 U11090 ( .A1(n10822), .A2(n10823), .ZN(n11057) );
  NAND2_X1 U11091 ( .A1(n11061), .A2(n11062), .ZN(n10823) );
  NAND2_X1 U11092 ( .A1(n11063), .A2(b_17_), .ZN(n11062) );
  NOR2_X1 U11093 ( .A1(n11064), .A2(n7464), .ZN(n11063) );
  NOR2_X1 U11094 ( .A1(n10830), .A2(n10831), .ZN(n11064) );
  NAND2_X1 U11095 ( .A1(n10830), .A2(n10831), .ZN(n11061) );
  NAND2_X1 U11096 ( .A1(n11065), .A2(n11066), .ZN(n10831) );
  NAND2_X1 U11097 ( .A1(n11067), .A2(b_17_), .ZN(n11066) );
  NOR2_X1 U11098 ( .A1(n11068), .A2(n7682), .ZN(n11067) );
  NOR2_X1 U11099 ( .A1(n10838), .A2(n10839), .ZN(n11068) );
  NAND2_X1 U11100 ( .A1(n10838), .A2(n10839), .ZN(n11065) );
  NAND2_X1 U11101 ( .A1(n11069), .A2(n11070), .ZN(n10839) );
  NAND2_X1 U11102 ( .A1(n11071), .A2(b_17_), .ZN(n11070) );
  NOR2_X1 U11103 ( .A1(n11072), .A2(n7455), .ZN(n11071) );
  NOR2_X1 U11104 ( .A1(n10846), .A2(n10847), .ZN(n11072) );
  NAND2_X1 U11105 ( .A1(n10846), .A2(n10847), .ZN(n11069) );
  NAND2_X1 U11106 ( .A1(n11073), .A2(n11074), .ZN(n10847) );
  NAND2_X1 U11107 ( .A1(n11075), .A2(b_17_), .ZN(n11074) );
  NOR2_X1 U11108 ( .A1(n11076), .A2(n7450), .ZN(n11075) );
  NOR2_X1 U11109 ( .A1(n11038), .A2(n11040), .ZN(n11076) );
  NAND2_X1 U11110 ( .A1(n11038), .A2(n11040), .ZN(n11073) );
  NAND2_X1 U11111 ( .A1(n11077), .A2(n11078), .ZN(n11040) );
  NAND2_X1 U11112 ( .A1(n11079), .A2(b_17_), .ZN(n11078) );
  NOR2_X1 U11113 ( .A1(n11080), .A2(n7445), .ZN(n11079) );
  NOR2_X1 U11114 ( .A1(n11034), .A2(n11036), .ZN(n11080) );
  NAND2_X1 U11115 ( .A1(n11034), .A2(n11036), .ZN(n11077) );
  NAND2_X1 U11116 ( .A1(n11081), .A2(n11082), .ZN(n11036) );
  NAND2_X1 U11117 ( .A1(n11083), .A2(b_17_), .ZN(n11082) );
  NOR2_X1 U11118 ( .A1(n11084), .A2(n7699), .ZN(n11083) );
  NOR2_X1 U11119 ( .A1(n10861), .A2(n10862), .ZN(n11084) );
  NAND2_X1 U11120 ( .A1(n10861), .A2(n10862), .ZN(n11081) );
  NAND2_X1 U11121 ( .A1(n11085), .A2(n11086), .ZN(n10862) );
  NAND2_X1 U11122 ( .A1(n11087), .A2(b_17_), .ZN(n11086) );
  NOR2_X1 U11123 ( .A1(n11088), .A2(n7704), .ZN(n11087) );
  NOR2_X1 U11124 ( .A1(n10869), .A2(n10870), .ZN(n11088) );
  NAND2_X1 U11125 ( .A1(n10869), .A2(n10870), .ZN(n11085) );
  NAND2_X1 U11126 ( .A1(n11089), .A2(n11090), .ZN(n10870) );
  NAND2_X1 U11127 ( .A1(n11091), .A2(b_17_), .ZN(n11090) );
  NOR2_X1 U11128 ( .A1(n11092), .A2(n7709), .ZN(n11091) );
  NOR2_X1 U11129 ( .A1(n11031), .A2(n11032), .ZN(n11092) );
  NAND2_X1 U11130 ( .A1(n11031), .A2(n11032), .ZN(n11089) );
  NAND2_X1 U11131 ( .A1(n11093), .A2(n11094), .ZN(n11032) );
  NAND2_X1 U11132 ( .A1(n11095), .A2(b_17_), .ZN(n11094) );
  NOR2_X1 U11133 ( .A1(n11096), .A2(n7424), .ZN(n11095) );
  NOR2_X1 U11134 ( .A1(n11027), .A2(n11028), .ZN(n11096) );
  NAND2_X1 U11135 ( .A1(n11027), .A2(n11028), .ZN(n11093) );
  NAND2_X1 U11136 ( .A1(n11097), .A2(n11098), .ZN(n11028) );
  NAND2_X1 U11137 ( .A1(n11099), .A2(b_17_), .ZN(n11098) );
  NOR2_X1 U11138 ( .A1(n11100), .A2(n7718), .ZN(n11099) );
  NOR2_X1 U11139 ( .A1(n11023), .A2(n11024), .ZN(n11100) );
  NAND2_X1 U11140 ( .A1(n11023), .A2(n11024), .ZN(n11097) );
  NAND2_X1 U11141 ( .A1(n11101), .A2(n11102), .ZN(n11024) );
  NAND2_X1 U11142 ( .A1(n11103), .A2(b_17_), .ZN(n11102) );
  NOR2_X1 U11143 ( .A1(n11104), .A2(n7415), .ZN(n11103) );
  NOR2_X1 U11144 ( .A1(n11019), .A2(n11020), .ZN(n11104) );
  NAND2_X1 U11145 ( .A1(n11019), .A2(n11020), .ZN(n11101) );
  NAND2_X1 U11146 ( .A1(n11105), .A2(n11106), .ZN(n11020) );
  NAND2_X1 U11147 ( .A1(n11017), .A2(n11107), .ZN(n11106) );
  OR2_X1 U11148 ( .A1(n11016), .A2(n11015), .ZN(n11107) );
  NOR2_X1 U11149 ( .A1(n10693), .A2(n7727), .ZN(n11017) );
  NAND2_X1 U11150 ( .A1(n11015), .A2(n11016), .ZN(n11105) );
  NAND2_X1 U11151 ( .A1(n11108), .A2(n11109), .ZN(n11016) );
  NAND2_X1 U11152 ( .A1(n11013), .A2(n11110), .ZN(n11109) );
  OR2_X1 U11153 ( .A1(n11012), .A2(n11011), .ZN(n11110) );
  NOR2_X1 U11154 ( .A1(n10693), .A2(n7406), .ZN(n11013) );
  NAND2_X1 U11155 ( .A1(n11011), .A2(n11012), .ZN(n11108) );
  NAND2_X1 U11156 ( .A1(n11111), .A2(n11112), .ZN(n11012) );
  NAND2_X1 U11157 ( .A1(n11113), .A2(b_17_), .ZN(n11112) );
  NOR2_X1 U11158 ( .A1(n11114), .A2(n7736), .ZN(n11113) );
  NOR2_X1 U11159 ( .A1(n11007), .A2(n11008), .ZN(n11114) );
  NAND2_X1 U11160 ( .A1(n11007), .A2(n11008), .ZN(n11111) );
  NAND2_X1 U11161 ( .A1(n11115), .A2(n11116), .ZN(n11008) );
  NAND2_X1 U11162 ( .A1(n11005), .A2(n11117), .ZN(n11116) );
  OR2_X1 U11163 ( .A1(n11004), .A2(n11002), .ZN(n11117) );
  NAND2_X1 U11164 ( .A1(n11002), .A2(n11004), .ZN(n11115) );
  NAND2_X1 U11165 ( .A1(n11118), .A2(n11119), .ZN(n11004) );
  NAND2_X1 U11166 ( .A1(n11120), .A2(b_17_), .ZN(n11119) );
  NOR2_X1 U11167 ( .A1(n11121), .A2(n7745), .ZN(n11120) );
  NOR2_X1 U11168 ( .A1(n10999), .A2(n11000), .ZN(n11121) );
  NAND2_X1 U11169 ( .A1(n10999), .A2(n11000), .ZN(n11118) );
  NAND2_X1 U11170 ( .A1(n11122), .A2(n11123), .ZN(n11000) );
  NAND2_X1 U11171 ( .A1(n10997), .A2(n11124), .ZN(n11123) );
  OR2_X1 U11172 ( .A1(n10996), .A2(n10994), .ZN(n11124) );
  NOR2_X1 U11173 ( .A1(n10693), .A2(n7750), .ZN(n10997) );
  NAND2_X1 U11174 ( .A1(n10994), .A2(n10996), .ZN(n11122) );
  NAND2_X1 U11175 ( .A1(n11125), .A2(n11126), .ZN(n10996) );
  NAND2_X1 U11176 ( .A1(n11127), .A2(b_17_), .ZN(n11126) );
  NOR2_X1 U11177 ( .A1(n11128), .A2(n7755), .ZN(n11127) );
  NOR2_X1 U11178 ( .A1(n10991), .A2(n10992), .ZN(n11128) );
  NAND2_X1 U11179 ( .A1(n10991), .A2(n10992), .ZN(n11125) );
  NAND2_X1 U11180 ( .A1(n11129), .A2(n11130), .ZN(n10992) );
  NAND2_X1 U11181 ( .A1(n10989), .A2(n11131), .ZN(n11130) );
  OR2_X1 U11182 ( .A1(n10988), .A2(n10987), .ZN(n11131) );
  NOR2_X1 U11183 ( .A1(n10693), .A2(n7760), .ZN(n10989) );
  NAND2_X1 U11184 ( .A1(n10987), .A2(n10988), .ZN(n11129) );
  NAND2_X1 U11185 ( .A1(n11132), .A2(n11133), .ZN(n10988) );
  NAND2_X1 U11186 ( .A1(n11134), .A2(b_17_), .ZN(n11133) );
  NOR2_X1 U11187 ( .A1(n11135), .A2(n7765), .ZN(n11134) );
  NOR2_X1 U11188 ( .A1(n10982), .A2(n10984), .ZN(n11135) );
  NAND2_X1 U11189 ( .A1(n10982), .A2(n10984), .ZN(n11132) );
  NAND2_X1 U11190 ( .A1(n11136), .A2(n11137), .ZN(n10984) );
  NAND2_X1 U11191 ( .A1(n10923), .A2(n11138), .ZN(n11137) );
  OR2_X1 U11192 ( .A1(n10922), .A2(n10921), .ZN(n11138) );
  NOR2_X1 U11193 ( .A1(n10693), .A2(n8014), .ZN(n10923) );
  NAND2_X1 U11194 ( .A1(n10921), .A2(n10922), .ZN(n11136) );
  NAND2_X1 U11195 ( .A1(n11139), .A2(n11140), .ZN(n10922) );
  NAND2_X1 U11196 ( .A1(n11141), .A2(b_17_), .ZN(n11140) );
  NOR2_X1 U11197 ( .A1(n11142), .A2(n7774), .ZN(n11141) );
  NOR2_X1 U11198 ( .A1(n10979), .A2(n10981), .ZN(n11142) );
  NAND2_X1 U11199 ( .A1(n10979), .A2(n10981), .ZN(n11139) );
  NAND2_X1 U11200 ( .A1(n11143), .A2(n11144), .ZN(n10981) );
  NAND2_X1 U11201 ( .A1(n10977), .A2(n11145), .ZN(n11144) );
  OR2_X1 U11202 ( .A1(n10976), .A2(n10975), .ZN(n11145) );
  NOR2_X1 U11203 ( .A1(n10693), .A2(n8022), .ZN(n10977) );
  NAND2_X1 U11204 ( .A1(n10975), .A2(n10976), .ZN(n11143) );
  NAND2_X1 U11205 ( .A1(n10972), .A2(n11146), .ZN(n10976) );
  NAND2_X1 U11206 ( .A1(n10971), .A2(n10973), .ZN(n11146) );
  NAND2_X1 U11207 ( .A1(n11147), .A2(n11148), .ZN(n10973) );
  NAND2_X1 U11208 ( .A1(b_17_), .A2(a_26_), .ZN(n11148) );
  INV_X1 U11209 ( .A(n11149), .ZN(n11147) );
  XNOR2_X1 U11210 ( .A(n11150), .B(n11151), .ZN(n10971) );
  NAND2_X1 U11211 ( .A1(n11152), .A2(n11153), .ZN(n11150) );
  NAND2_X1 U11212 ( .A1(a_26_), .A2(n11149), .ZN(n10972) );
  NAND2_X1 U11213 ( .A1(n10941), .A2(n11154), .ZN(n11149) );
  NAND2_X1 U11214 ( .A1(n10940), .A2(n10942), .ZN(n11154) );
  NAND2_X1 U11215 ( .A1(n11155), .A2(n11156), .ZN(n10942) );
  NAND2_X1 U11216 ( .A1(b_17_), .A2(a_27_), .ZN(n11156) );
  INV_X1 U11217 ( .A(n11157), .ZN(n11155) );
  XNOR2_X1 U11218 ( .A(n11158), .B(n11159), .ZN(n10940) );
  XOR2_X1 U11219 ( .A(n11160), .B(n11161), .Z(n11159) );
  NAND2_X1 U11220 ( .A1(b_16_), .A2(a_28_), .ZN(n11161) );
  NAND2_X1 U11221 ( .A1(a_27_), .A2(n11157), .ZN(n10941) );
  NAND2_X1 U11222 ( .A1(n11162), .A2(n11163), .ZN(n11157) );
  NAND2_X1 U11223 ( .A1(n11164), .A2(b_17_), .ZN(n11163) );
  NOR2_X1 U11224 ( .A1(n11165), .A2(n7803), .ZN(n11164) );
  NOR2_X1 U11225 ( .A1(n10947), .A2(n10949), .ZN(n11165) );
  NAND2_X1 U11226 ( .A1(n10947), .A2(n10949), .ZN(n11162) );
  NAND2_X1 U11227 ( .A1(n11166), .A2(n11167), .ZN(n10949) );
  NAND2_X1 U11228 ( .A1(n10967), .A2(n11168), .ZN(n11167) );
  NAND2_X1 U11229 ( .A1(n10969), .A2(n10968), .ZN(n11168) );
  NOR2_X1 U11230 ( .A1(n10693), .A2(n7337), .ZN(n10967) );
  OR2_X1 U11231 ( .A1(n10968), .A2(n10969), .ZN(n11166) );
  AND2_X1 U11232 ( .A1(n11169), .A2(n11170), .ZN(n10969) );
  NAND2_X1 U11233 ( .A1(n11171), .A2(b_15_), .ZN(n11170) );
  NOR2_X1 U11234 ( .A1(n11172), .A2(n7817), .ZN(n11171) );
  NOR2_X1 U11235 ( .A1(n7816), .A2(n10964), .ZN(n11172) );
  NAND2_X1 U11236 ( .A1(n11173), .A2(b_16_), .ZN(n11169) );
  NOR2_X1 U11237 ( .A1(n11174), .A2(n8052), .ZN(n11173) );
  NOR2_X1 U11238 ( .A1(n7810), .A2(n11175), .ZN(n11174) );
  NAND2_X1 U11239 ( .A1(n10965), .A2(b_16_), .ZN(n10968) );
  NOR2_X1 U11240 ( .A1(n8055), .A2(n10693), .ZN(n10965) );
  XOR2_X1 U11241 ( .A(n11176), .B(n11177), .Z(n10947) );
  XOR2_X1 U11242 ( .A(n11178), .B(n11179), .Z(n11176) );
  XNOR2_X1 U11243 ( .A(n11180), .B(n11181), .ZN(n10975) );
  NAND2_X1 U11244 ( .A1(n11182), .A2(n11183), .ZN(n11180) );
  XOR2_X1 U11245 ( .A(n11184), .B(n11185), .Z(n10979) );
  XOR2_X1 U11246 ( .A(n11186), .B(n11187), .Z(n11184) );
  XOR2_X1 U11247 ( .A(n11188), .B(n11189), .Z(n10921) );
  XOR2_X1 U11248 ( .A(n11190), .B(n11191), .Z(n11188) );
  NOR2_X1 U11249 ( .A1(n7774), .A2(n10964), .ZN(n11191) );
  XOR2_X1 U11250 ( .A(n11192), .B(n11193), .Z(n10982) );
  XOR2_X1 U11251 ( .A(n11194), .B(n11195), .Z(n11192) );
  XNOR2_X1 U11252 ( .A(n11196), .B(n11197), .ZN(n10987) );
  XOR2_X1 U11253 ( .A(n11198), .B(n11199), .Z(n11197) );
  NAND2_X1 U11254 ( .A1(b_16_), .A2(a_22_), .ZN(n11199) );
  XOR2_X1 U11255 ( .A(n11200), .B(n11201), .Z(n10991) );
  XOR2_X1 U11256 ( .A(n11202), .B(n11203), .Z(n11200) );
  XOR2_X1 U11257 ( .A(n11204), .B(n11205), .Z(n10994) );
  XOR2_X1 U11258 ( .A(n11206), .B(n11207), .Z(n11204) );
  NOR2_X1 U11259 ( .A1(n7755), .A2(n10964), .ZN(n11207) );
  XOR2_X1 U11260 ( .A(n11208), .B(n11209), .Z(n10999) );
  XOR2_X1 U11261 ( .A(n11210), .B(n11211), .Z(n11208) );
  XOR2_X1 U11262 ( .A(n11212), .B(n11213), .Z(n11002) );
  XOR2_X1 U11263 ( .A(n11214), .B(n11215), .Z(n11212) );
  NOR2_X1 U11264 ( .A1(n7745), .A2(n10964), .ZN(n11215) );
  XOR2_X1 U11265 ( .A(n11216), .B(n11217), .Z(n11007) );
  XOR2_X1 U11266 ( .A(n11218), .B(n11219), .Z(n11216) );
  XNOR2_X1 U11267 ( .A(n11220), .B(n11221), .ZN(n11011) );
  XNOR2_X1 U11268 ( .A(n11222), .B(n11223), .ZN(n11220) );
  XNOR2_X1 U11269 ( .A(n11224), .B(n11225), .ZN(n11015) );
  XOR2_X1 U11270 ( .A(n11226), .B(n11227), .Z(n11225) );
  NAND2_X1 U11271 ( .A1(b_16_), .A2(a_15_), .ZN(n11227) );
  XNOR2_X1 U11272 ( .A(n11228), .B(n11229), .ZN(n11019) );
  XNOR2_X1 U11273 ( .A(n11230), .B(n11231), .ZN(n11228) );
  XNOR2_X1 U11274 ( .A(n11232), .B(n11233), .ZN(n11023) );
  XNOR2_X1 U11275 ( .A(n11234), .B(n11235), .ZN(n11233) );
  XNOR2_X1 U11276 ( .A(n11236), .B(n11237), .ZN(n11027) );
  XNOR2_X1 U11277 ( .A(n11238), .B(n11239), .ZN(n11236) );
  XNOR2_X1 U11278 ( .A(n11240), .B(n11241), .ZN(n11031) );
  XNOR2_X1 U11279 ( .A(n11242), .B(n11243), .ZN(n11241) );
  XOR2_X1 U11280 ( .A(n11244), .B(n11245), .Z(n10869) );
  XOR2_X1 U11281 ( .A(n11246), .B(n11247), .Z(n11244) );
  NOR2_X1 U11282 ( .A1(n7709), .A2(n10964), .ZN(n11247) );
  XNOR2_X1 U11283 ( .A(n11248), .B(n11249), .ZN(n10861) );
  NAND2_X1 U11284 ( .A1(n11250), .A2(n11251), .ZN(n11248) );
  XNOR2_X1 U11285 ( .A(n11252), .B(n11253), .ZN(n11034) );
  XNOR2_X1 U11286 ( .A(n11254), .B(n11255), .ZN(n11252) );
  XNOR2_X1 U11287 ( .A(n11256), .B(n11257), .ZN(n11038) );
  XNOR2_X1 U11288 ( .A(n11258), .B(n11259), .ZN(n11257) );
  XNOR2_X1 U11289 ( .A(n11260), .B(n11261), .ZN(n10846) );
  XNOR2_X1 U11290 ( .A(n11262), .B(n11263), .ZN(n11261) );
  XNOR2_X1 U11291 ( .A(n11264), .B(n11265), .ZN(n10838) );
  XOR2_X1 U11292 ( .A(n11266), .B(n11267), .Z(n11265) );
  NAND2_X1 U11293 ( .A1(b_16_), .A2(a_5_), .ZN(n11267) );
  XOR2_X1 U11294 ( .A(n11268), .B(n11269), .Z(n10830) );
  XOR2_X1 U11295 ( .A(n11270), .B(n11271), .Z(n11268) );
  XNOR2_X1 U11296 ( .A(n11272), .B(n11273), .ZN(n10822) );
  XNOR2_X1 U11297 ( .A(n11274), .B(n11275), .ZN(n11272) );
  XOR2_X1 U11298 ( .A(n11276), .B(n11277), .Z(n10814) );
  XNOR2_X1 U11299 ( .A(n11278), .B(n11279), .ZN(n11276) );
  NAND2_X1 U11300 ( .A1(b_16_), .A2(a_2_), .ZN(n11278) );
  XNOR2_X1 U11301 ( .A(n11280), .B(n11281), .ZN(n10807) );
  NAND2_X1 U11302 ( .A1(n11282), .A2(n11283), .ZN(n11280) );
  NAND2_X1 U11303 ( .A1(n11284), .A2(n11285), .ZN(n7551) );
  NAND2_X1 U11304 ( .A1(n11286), .A2(n7604), .ZN(n11285) );
  INV_X1 U11305 ( .A(n7605), .ZN(n11286) );
  XOR2_X1 U11306 ( .A(n11287), .B(n11288), .Z(n11284) );
  NAND2_X1 U11307 ( .A1(n11289), .A2(n11290), .ZN(n7552) );
  XOR2_X1 U11308 ( .A(n11287), .B(n11291), .Z(n11290) );
  NOR2_X1 U11309 ( .A1(n11044), .A2(n7605), .ZN(n11289) );
  XNOR2_X1 U11310 ( .A(n11292), .B(n11293), .ZN(n7605) );
  XOR2_X1 U11311 ( .A(n11294), .B(n11295), .Z(n11292) );
  NOR2_X1 U11312 ( .A1(n7478), .A2(n11175), .ZN(n11295) );
  INV_X1 U11313 ( .A(n7604), .ZN(n11044) );
  NAND2_X1 U11314 ( .A1(n11047), .A2(n11296), .ZN(n7604) );
  NAND2_X1 U11315 ( .A1(n11046), .A2(n11048), .ZN(n11296) );
  NAND2_X1 U11316 ( .A1(n11297), .A2(n11298), .ZN(n11048) );
  NAND2_X1 U11317 ( .A1(b_16_), .A2(a_0_), .ZN(n11298) );
  INV_X1 U11318 ( .A(n11299), .ZN(n11297) );
  XNOR2_X1 U11319 ( .A(n11300), .B(n11301), .ZN(n11046) );
  NAND2_X1 U11320 ( .A1(n11302), .A2(n11303), .ZN(n11300) );
  NAND2_X1 U11321 ( .A1(a_0_), .A2(n11299), .ZN(n11047) );
  NAND2_X1 U11322 ( .A1(n11282), .A2(n11304), .ZN(n11299) );
  NAND2_X1 U11323 ( .A1(n11281), .A2(n11283), .ZN(n11304) );
  NAND2_X1 U11324 ( .A1(n11305), .A2(n11306), .ZN(n11283) );
  NAND2_X1 U11325 ( .A1(b_16_), .A2(a_1_), .ZN(n11306) );
  INV_X1 U11326 ( .A(n11307), .ZN(n11305) );
  XOR2_X1 U11327 ( .A(n11308), .B(n11309), .Z(n11281) );
  XOR2_X1 U11328 ( .A(n11310), .B(n11311), .Z(n11308) );
  NOR2_X1 U11329 ( .A1(n7469), .A2(n11175), .ZN(n11311) );
  NAND2_X1 U11330 ( .A1(a_1_), .A2(n11307), .ZN(n11282) );
  NAND2_X1 U11331 ( .A1(n11312), .A2(n11313), .ZN(n11307) );
  NAND2_X1 U11332 ( .A1(n11314), .A2(b_16_), .ZN(n11313) );
  NOR2_X1 U11333 ( .A1(n11315), .A2(n7469), .ZN(n11314) );
  NOR2_X1 U11334 ( .A1(n11277), .A2(n11279), .ZN(n11315) );
  NAND2_X1 U11335 ( .A1(n11277), .A2(n11279), .ZN(n11312) );
  NAND2_X1 U11336 ( .A1(n11316), .A2(n11317), .ZN(n11279) );
  NAND2_X1 U11337 ( .A1(n11275), .A2(n11318), .ZN(n11317) );
  NAND2_X1 U11338 ( .A1(n11274), .A2(n11273), .ZN(n11318) );
  NOR2_X1 U11339 ( .A1(n10964), .A2(n7464), .ZN(n11275) );
  OR2_X1 U11340 ( .A1(n11273), .A2(n11274), .ZN(n11316) );
  AND2_X1 U11341 ( .A1(n11319), .A2(n11320), .ZN(n11274) );
  NAND2_X1 U11342 ( .A1(n11271), .A2(n11321), .ZN(n11320) );
  OR2_X1 U11343 ( .A1(n11269), .A2(n11270), .ZN(n11321) );
  NOR2_X1 U11344 ( .A1(n10964), .A2(n7682), .ZN(n11271) );
  NAND2_X1 U11345 ( .A1(n11269), .A2(n11270), .ZN(n11319) );
  NAND2_X1 U11346 ( .A1(n11322), .A2(n11323), .ZN(n11270) );
  NAND2_X1 U11347 ( .A1(n11324), .A2(b_16_), .ZN(n11323) );
  NOR2_X1 U11348 ( .A1(n11325), .A2(n7455), .ZN(n11324) );
  NOR2_X1 U11349 ( .A1(n11264), .A2(n11266), .ZN(n11325) );
  NAND2_X1 U11350 ( .A1(n11264), .A2(n11266), .ZN(n11322) );
  NAND2_X1 U11351 ( .A1(n11326), .A2(n11327), .ZN(n11266) );
  NAND2_X1 U11352 ( .A1(n11263), .A2(n11328), .ZN(n11327) );
  OR2_X1 U11353 ( .A1(n11262), .A2(n11260), .ZN(n11328) );
  NOR2_X1 U11354 ( .A1(n10964), .A2(n7450), .ZN(n11263) );
  NAND2_X1 U11355 ( .A1(n11260), .A2(n11262), .ZN(n11326) );
  NAND2_X1 U11356 ( .A1(n11329), .A2(n11330), .ZN(n11262) );
  NAND2_X1 U11357 ( .A1(n11259), .A2(n11331), .ZN(n11330) );
  OR2_X1 U11358 ( .A1(n11258), .A2(n11256), .ZN(n11331) );
  NOR2_X1 U11359 ( .A1(n10964), .A2(n7445), .ZN(n11259) );
  NAND2_X1 U11360 ( .A1(n11256), .A2(n11258), .ZN(n11329) );
  NAND2_X1 U11361 ( .A1(n11332), .A2(n11333), .ZN(n11258) );
  NAND2_X1 U11362 ( .A1(n11255), .A2(n11334), .ZN(n11333) );
  NAND2_X1 U11363 ( .A1(n11254), .A2(n11253), .ZN(n11334) );
  NOR2_X1 U11364 ( .A1(n10964), .A2(n7699), .ZN(n11255) );
  OR2_X1 U11365 ( .A1(n11253), .A2(n11254), .ZN(n11332) );
  AND2_X1 U11366 ( .A1(n11250), .A2(n11335), .ZN(n11254) );
  NAND2_X1 U11367 ( .A1(n11249), .A2(n11251), .ZN(n11335) );
  NAND2_X1 U11368 ( .A1(n11336), .A2(n11337), .ZN(n11251) );
  NAND2_X1 U11369 ( .A1(b_16_), .A2(a_9_), .ZN(n11337) );
  INV_X1 U11370 ( .A(n11338), .ZN(n11336) );
  XOR2_X1 U11371 ( .A(n11339), .B(n11340), .Z(n11249) );
  XOR2_X1 U11372 ( .A(n11341), .B(n11342), .Z(n11339) );
  NOR2_X1 U11373 ( .A1(n7709), .A2(n11175), .ZN(n11342) );
  NAND2_X1 U11374 ( .A1(a_9_), .A2(n11338), .ZN(n11250) );
  NAND2_X1 U11375 ( .A1(n11343), .A2(n11344), .ZN(n11338) );
  NAND2_X1 U11376 ( .A1(n11345), .A2(b_16_), .ZN(n11344) );
  NOR2_X1 U11377 ( .A1(n11346), .A2(n7709), .ZN(n11345) );
  NOR2_X1 U11378 ( .A1(n11245), .A2(n11246), .ZN(n11346) );
  NAND2_X1 U11379 ( .A1(n11245), .A2(n11246), .ZN(n11343) );
  NAND2_X1 U11380 ( .A1(n11347), .A2(n11348), .ZN(n11246) );
  NAND2_X1 U11381 ( .A1(n11243), .A2(n11349), .ZN(n11348) );
  OR2_X1 U11382 ( .A1(n11242), .A2(n11240), .ZN(n11349) );
  NOR2_X1 U11383 ( .A1(n10964), .A2(n7424), .ZN(n11243) );
  NAND2_X1 U11384 ( .A1(n11240), .A2(n11242), .ZN(n11347) );
  NAND2_X1 U11385 ( .A1(n11350), .A2(n11351), .ZN(n11242) );
  NAND2_X1 U11386 ( .A1(n11239), .A2(n11352), .ZN(n11351) );
  NAND2_X1 U11387 ( .A1(n11238), .A2(n11237), .ZN(n11352) );
  NOR2_X1 U11388 ( .A1(n10964), .A2(n7718), .ZN(n11239) );
  OR2_X1 U11389 ( .A1(n11237), .A2(n11238), .ZN(n11350) );
  AND2_X1 U11390 ( .A1(n11353), .A2(n11354), .ZN(n11238) );
  NAND2_X1 U11391 ( .A1(n11235), .A2(n11355), .ZN(n11354) );
  OR2_X1 U11392 ( .A1(n11232), .A2(n11234), .ZN(n11355) );
  NOR2_X1 U11393 ( .A1(n10964), .A2(n7415), .ZN(n11235) );
  NAND2_X1 U11394 ( .A1(n11232), .A2(n11234), .ZN(n11353) );
  NAND2_X1 U11395 ( .A1(n11356), .A2(n11357), .ZN(n11234) );
  NAND2_X1 U11396 ( .A1(n11231), .A2(n11358), .ZN(n11357) );
  NAND2_X1 U11397 ( .A1(n11230), .A2(n11229), .ZN(n11358) );
  NOR2_X1 U11398 ( .A1(n10964), .A2(n7727), .ZN(n11231) );
  OR2_X1 U11399 ( .A1(n11229), .A2(n11230), .ZN(n11356) );
  AND2_X1 U11400 ( .A1(n11359), .A2(n11360), .ZN(n11230) );
  NAND2_X1 U11401 ( .A1(n11361), .A2(b_16_), .ZN(n11360) );
  NOR2_X1 U11402 ( .A1(n11362), .A2(n7406), .ZN(n11361) );
  NOR2_X1 U11403 ( .A1(n11224), .A2(n11226), .ZN(n11362) );
  NAND2_X1 U11404 ( .A1(n11224), .A2(n11226), .ZN(n11359) );
  NAND2_X1 U11405 ( .A1(n11363), .A2(n11364), .ZN(n11226) );
  NAND2_X1 U11406 ( .A1(n11223), .A2(n11365), .ZN(n11364) );
  NAND2_X1 U11407 ( .A1(n11222), .A2(n11221), .ZN(n11365) );
  OR2_X1 U11408 ( .A1(n11221), .A2(n11222), .ZN(n11363) );
  AND2_X1 U11409 ( .A1(n11366), .A2(n11367), .ZN(n11222) );
  NAND2_X1 U11410 ( .A1(n11219), .A2(n11368), .ZN(n11367) );
  OR2_X1 U11411 ( .A1(n11217), .A2(n11218), .ZN(n11368) );
  NOR2_X1 U11412 ( .A1(n10964), .A2(n7397), .ZN(n11219) );
  NAND2_X1 U11413 ( .A1(n11217), .A2(n11218), .ZN(n11366) );
  NAND2_X1 U11414 ( .A1(n11369), .A2(n11370), .ZN(n11218) );
  NAND2_X1 U11415 ( .A1(n11371), .A2(b_16_), .ZN(n11370) );
  NOR2_X1 U11416 ( .A1(n11372), .A2(n7745), .ZN(n11371) );
  NOR2_X1 U11417 ( .A1(n11213), .A2(n11214), .ZN(n11372) );
  NAND2_X1 U11418 ( .A1(n11213), .A2(n11214), .ZN(n11369) );
  NAND2_X1 U11419 ( .A1(n11373), .A2(n11374), .ZN(n11214) );
  NAND2_X1 U11420 ( .A1(n11211), .A2(n11375), .ZN(n11374) );
  OR2_X1 U11421 ( .A1(n11209), .A2(n11210), .ZN(n11375) );
  NOR2_X1 U11422 ( .A1(n10964), .A2(n7750), .ZN(n11211) );
  NAND2_X1 U11423 ( .A1(n11209), .A2(n11210), .ZN(n11373) );
  NAND2_X1 U11424 ( .A1(n11376), .A2(n11377), .ZN(n11210) );
  NAND2_X1 U11425 ( .A1(n11378), .A2(b_16_), .ZN(n11377) );
  NOR2_X1 U11426 ( .A1(n11379), .A2(n7755), .ZN(n11378) );
  NOR2_X1 U11427 ( .A1(n11205), .A2(n11206), .ZN(n11379) );
  NAND2_X1 U11428 ( .A1(n11205), .A2(n11206), .ZN(n11376) );
  NAND2_X1 U11429 ( .A1(n11380), .A2(n11381), .ZN(n11206) );
  NAND2_X1 U11430 ( .A1(n11203), .A2(n11382), .ZN(n11381) );
  OR2_X1 U11431 ( .A1(n11201), .A2(n11202), .ZN(n11382) );
  NOR2_X1 U11432 ( .A1(n10964), .A2(n7760), .ZN(n11203) );
  NAND2_X1 U11433 ( .A1(n11201), .A2(n11202), .ZN(n11380) );
  NAND2_X1 U11434 ( .A1(n11383), .A2(n11384), .ZN(n11202) );
  NAND2_X1 U11435 ( .A1(n11385), .A2(b_16_), .ZN(n11384) );
  NOR2_X1 U11436 ( .A1(n11386), .A2(n7765), .ZN(n11385) );
  NOR2_X1 U11437 ( .A1(n11196), .A2(n11198), .ZN(n11386) );
  NAND2_X1 U11438 ( .A1(n11196), .A2(n11198), .ZN(n11383) );
  NAND2_X1 U11439 ( .A1(n11387), .A2(n11388), .ZN(n11198) );
  NAND2_X1 U11440 ( .A1(n11195), .A2(n11389), .ZN(n11388) );
  OR2_X1 U11441 ( .A1(n11193), .A2(n11194), .ZN(n11389) );
  NOR2_X1 U11442 ( .A1(n10964), .A2(n8014), .ZN(n11195) );
  NAND2_X1 U11443 ( .A1(n11193), .A2(n11194), .ZN(n11387) );
  NAND2_X1 U11444 ( .A1(n11390), .A2(n11391), .ZN(n11194) );
  NAND2_X1 U11445 ( .A1(n11392), .A2(b_16_), .ZN(n11391) );
  NOR2_X1 U11446 ( .A1(n11393), .A2(n7774), .ZN(n11392) );
  NOR2_X1 U11447 ( .A1(n11189), .A2(n11190), .ZN(n11393) );
  NAND2_X1 U11448 ( .A1(n11189), .A2(n11190), .ZN(n11390) );
  NAND2_X1 U11449 ( .A1(n11394), .A2(n11395), .ZN(n11190) );
  NAND2_X1 U11450 ( .A1(n11187), .A2(n11396), .ZN(n11395) );
  OR2_X1 U11451 ( .A1(n11185), .A2(n11186), .ZN(n11396) );
  NOR2_X1 U11452 ( .A1(n10964), .A2(n8022), .ZN(n11187) );
  NAND2_X1 U11453 ( .A1(n11185), .A2(n11186), .ZN(n11394) );
  NAND2_X1 U11454 ( .A1(n11182), .A2(n11397), .ZN(n11186) );
  NAND2_X1 U11455 ( .A1(n11181), .A2(n11183), .ZN(n11397) );
  NAND2_X1 U11456 ( .A1(n11398), .A2(n11399), .ZN(n11183) );
  NAND2_X1 U11457 ( .A1(b_16_), .A2(a_26_), .ZN(n11399) );
  INV_X1 U11458 ( .A(n11400), .ZN(n11398) );
  XNOR2_X1 U11459 ( .A(n11401), .B(n11402), .ZN(n11181) );
  NAND2_X1 U11460 ( .A1(n11403), .A2(n11404), .ZN(n11401) );
  NAND2_X1 U11461 ( .A1(a_26_), .A2(n11400), .ZN(n11182) );
  NAND2_X1 U11462 ( .A1(n11152), .A2(n11405), .ZN(n11400) );
  NAND2_X1 U11463 ( .A1(n11151), .A2(n11153), .ZN(n11405) );
  NAND2_X1 U11464 ( .A1(n11406), .A2(n11407), .ZN(n11153) );
  NAND2_X1 U11465 ( .A1(b_16_), .A2(a_27_), .ZN(n11407) );
  INV_X1 U11466 ( .A(n11408), .ZN(n11406) );
  XNOR2_X1 U11467 ( .A(n11409), .B(n11410), .ZN(n11151) );
  XOR2_X1 U11468 ( .A(n11411), .B(n11412), .Z(n11410) );
  NAND2_X1 U11469 ( .A1(b_15_), .A2(a_28_), .ZN(n11412) );
  NAND2_X1 U11470 ( .A1(a_27_), .A2(n11408), .ZN(n11152) );
  NAND2_X1 U11471 ( .A1(n11413), .A2(n11414), .ZN(n11408) );
  NAND2_X1 U11472 ( .A1(n11415), .A2(b_16_), .ZN(n11414) );
  NOR2_X1 U11473 ( .A1(n11416), .A2(n7803), .ZN(n11415) );
  NOR2_X1 U11474 ( .A1(n11158), .A2(n11160), .ZN(n11416) );
  NAND2_X1 U11475 ( .A1(n11158), .A2(n11160), .ZN(n11413) );
  NAND2_X1 U11476 ( .A1(n11417), .A2(n11418), .ZN(n11160) );
  NAND2_X1 U11477 ( .A1(n11177), .A2(n11419), .ZN(n11418) );
  NAND2_X1 U11478 ( .A1(n11179), .A2(n11178), .ZN(n11419) );
  NOR2_X1 U11479 ( .A1(n10964), .A2(n7337), .ZN(n11177) );
  OR2_X1 U11480 ( .A1(n11178), .A2(n11179), .ZN(n11417) );
  AND2_X1 U11481 ( .A1(n11420), .A2(n11421), .ZN(n11179) );
  NAND2_X1 U11482 ( .A1(n11422), .A2(b_14_), .ZN(n11421) );
  NOR2_X1 U11483 ( .A1(n11423), .A2(n7817), .ZN(n11422) );
  NOR2_X1 U11484 ( .A1(n7816), .A2(n11175), .ZN(n11423) );
  NAND2_X1 U11485 ( .A1(n11424), .A2(b_15_), .ZN(n11420) );
  NOR2_X1 U11486 ( .A1(n11425), .A2(n8052), .ZN(n11424) );
  NOR2_X1 U11487 ( .A1(n7810), .A2(n11426), .ZN(n11425) );
  NAND2_X1 U11488 ( .A1(n11427), .A2(b_15_), .ZN(n11178) );
  NOR2_X1 U11489 ( .A1(n8055), .A2(n10964), .ZN(n11427) );
  XOR2_X1 U11490 ( .A(n11428), .B(n11429), .Z(n11158) );
  XOR2_X1 U11491 ( .A(n11430), .B(n11431), .Z(n11428) );
  XNOR2_X1 U11492 ( .A(n11432), .B(n11433), .ZN(n11185) );
  NAND2_X1 U11493 ( .A1(n11434), .A2(n11435), .ZN(n11432) );
  XOR2_X1 U11494 ( .A(n11436), .B(n11437), .Z(n11189) );
  XOR2_X1 U11495 ( .A(n11438), .B(n11439), .Z(n11436) );
  XOR2_X1 U11496 ( .A(n11440), .B(n11441), .Z(n11193) );
  XOR2_X1 U11497 ( .A(n11442), .B(n11443), .Z(n11440) );
  NOR2_X1 U11498 ( .A1(n7774), .A2(n11175), .ZN(n11443) );
  XOR2_X1 U11499 ( .A(n11444), .B(n11445), .Z(n11196) );
  XOR2_X1 U11500 ( .A(n11446), .B(n11447), .Z(n11444) );
  XOR2_X1 U11501 ( .A(n11448), .B(n11449), .Z(n11201) );
  XOR2_X1 U11502 ( .A(n11450), .B(n11451), .Z(n11448) );
  NOR2_X1 U11503 ( .A1(n7765), .A2(n11175), .ZN(n11451) );
  XOR2_X1 U11504 ( .A(n11452), .B(n11453), .Z(n11205) );
  XOR2_X1 U11505 ( .A(n11454), .B(n11455), .Z(n11452) );
  XOR2_X1 U11506 ( .A(n11456), .B(n11457), .Z(n11209) );
  XOR2_X1 U11507 ( .A(n11458), .B(n11459), .Z(n11456) );
  NOR2_X1 U11508 ( .A1(n7755), .A2(n11175), .ZN(n11459) );
  XOR2_X1 U11509 ( .A(n11460), .B(n11461), .Z(n11213) );
  XOR2_X1 U11510 ( .A(n11462), .B(n11463), .Z(n11460) );
  XOR2_X1 U11511 ( .A(n11464), .B(n11465), .Z(n11217) );
  XOR2_X1 U11512 ( .A(n11466), .B(n11467), .Z(n11464) );
  NOR2_X1 U11513 ( .A1(n7745), .A2(n11175), .ZN(n11467) );
  XNOR2_X1 U11514 ( .A(n11468), .B(n11469), .ZN(n11221) );
  XOR2_X1 U11515 ( .A(n11470), .B(n11471), .Z(n11468) );
  XOR2_X1 U11516 ( .A(n11472), .B(n11473), .Z(n11224) );
  XOR2_X1 U11517 ( .A(n11474), .B(n11475), .Z(n11472) );
  XNOR2_X1 U11518 ( .A(n11476), .B(n11477), .ZN(n11229) );
  XOR2_X1 U11519 ( .A(n11478), .B(n11479), .Z(n11476) );
  XOR2_X1 U11520 ( .A(n11480), .B(n11481), .Z(n11232) );
  XNOR2_X1 U11521 ( .A(n11482), .B(n11483), .ZN(n11480) );
  NAND2_X1 U11522 ( .A1(b_15_), .A2(a_14_), .ZN(n11482) );
  XNOR2_X1 U11523 ( .A(n11484), .B(n11485), .ZN(n11237) );
  XOR2_X1 U11524 ( .A(n11486), .B(n11487), .Z(n11484) );
  NOR2_X1 U11525 ( .A1(n7415), .A2(n11175), .ZN(n11487) );
  XNOR2_X1 U11526 ( .A(n11488), .B(n11489), .ZN(n11240) );
  XOR2_X1 U11527 ( .A(n11490), .B(n11491), .Z(n11489) );
  NAND2_X1 U11528 ( .A1(b_15_), .A2(a_12_), .ZN(n11491) );
  XNOR2_X1 U11529 ( .A(n11492), .B(n11493), .ZN(n11245) );
  XOR2_X1 U11530 ( .A(n11494), .B(n11495), .Z(n11493) );
  NAND2_X1 U11531 ( .A1(b_15_), .A2(a_11_), .ZN(n11495) );
  XOR2_X1 U11532 ( .A(n11496), .B(n11497), .Z(n11253) );
  XOR2_X1 U11533 ( .A(n11498), .B(n11499), .Z(n11497) );
  NAND2_X1 U11534 ( .A1(b_15_), .A2(a_9_), .ZN(n11499) );
  XOR2_X1 U11535 ( .A(n11500), .B(n11501), .Z(n11256) );
  XOR2_X1 U11536 ( .A(n11502), .B(n11503), .Z(n11500) );
  NOR2_X1 U11537 ( .A1(n7699), .A2(n11175), .ZN(n11503) );
  XOR2_X1 U11538 ( .A(n11504), .B(n11505), .Z(n11260) );
  XOR2_X1 U11539 ( .A(n11506), .B(n11507), .Z(n11504) );
  NOR2_X1 U11540 ( .A1(n7445), .A2(n11175), .ZN(n11507) );
  XOR2_X1 U11541 ( .A(n11508), .B(n11509), .Z(n11264) );
  XOR2_X1 U11542 ( .A(n11510), .B(n11511), .Z(n11508) );
  NOR2_X1 U11543 ( .A1(n7450), .A2(n11175), .ZN(n11511) );
  XNOR2_X1 U11544 ( .A(n11512), .B(n11513), .ZN(n11269) );
  XOR2_X1 U11545 ( .A(n11514), .B(n11515), .Z(n11513) );
  NAND2_X1 U11546 ( .A1(b_15_), .A2(a_5_), .ZN(n11515) );
  XOR2_X1 U11547 ( .A(n11516), .B(n11517), .Z(n11273) );
  XOR2_X1 U11548 ( .A(n11518), .B(n11519), .Z(n11517) );
  NAND2_X1 U11549 ( .A1(b_15_), .A2(a_4_), .ZN(n11519) );
  XNOR2_X1 U11550 ( .A(n11520), .B(n11521), .ZN(n11277) );
  XOR2_X1 U11551 ( .A(n11522), .B(n11523), .Z(n11521) );
  NAND2_X1 U11552 ( .A1(b_15_), .A2(a_3_), .ZN(n11523) );
  NAND2_X1 U11553 ( .A1(n11524), .A2(n11525), .ZN(n7555) );
  NAND2_X1 U11554 ( .A1(n11291), .A2(n11287), .ZN(n11525) );
  XNOR2_X1 U11555 ( .A(n11526), .B(n11527), .ZN(n11524) );
  NAND2_X1 U11556 ( .A1(n11528), .A2(n11529), .ZN(n7556) );
  AND2_X1 U11557 ( .A1(n7596), .A2(n11287), .ZN(n11529) );
  NAND2_X1 U11558 ( .A1(n11530), .A2(n11531), .ZN(n11287) );
  NAND2_X1 U11559 ( .A1(n11532), .A2(b_15_), .ZN(n11531) );
  NOR2_X1 U11560 ( .A1(n11533), .A2(n7478), .ZN(n11532) );
  NOR2_X1 U11561 ( .A1(n11293), .A2(n11294), .ZN(n11533) );
  NAND2_X1 U11562 ( .A1(n11293), .A2(n11294), .ZN(n11530) );
  NAND2_X1 U11563 ( .A1(n11302), .A2(n11534), .ZN(n11294) );
  NAND2_X1 U11564 ( .A1(n11301), .A2(n11303), .ZN(n11534) );
  NAND2_X1 U11565 ( .A1(n11535), .A2(n11536), .ZN(n11303) );
  NAND2_X1 U11566 ( .A1(b_15_), .A2(a_1_), .ZN(n11536) );
  INV_X1 U11567 ( .A(n11537), .ZN(n11535) );
  XNOR2_X1 U11568 ( .A(n11538), .B(n11539), .ZN(n11301) );
  NAND2_X1 U11569 ( .A1(n11540), .A2(n11541), .ZN(n11538) );
  NAND2_X1 U11570 ( .A1(a_1_), .A2(n11537), .ZN(n11302) );
  NAND2_X1 U11571 ( .A1(n11542), .A2(n11543), .ZN(n11537) );
  NAND2_X1 U11572 ( .A1(n11544), .A2(b_15_), .ZN(n11543) );
  NOR2_X1 U11573 ( .A1(n11545), .A2(n7469), .ZN(n11544) );
  NOR2_X1 U11574 ( .A1(n11310), .A2(n11309), .ZN(n11545) );
  NAND2_X1 U11575 ( .A1(n11309), .A2(n11310), .ZN(n11542) );
  NAND2_X1 U11576 ( .A1(n11546), .A2(n11547), .ZN(n11310) );
  NAND2_X1 U11577 ( .A1(n11548), .A2(b_15_), .ZN(n11547) );
  NOR2_X1 U11578 ( .A1(n11549), .A2(n7464), .ZN(n11548) );
  NOR2_X1 U11579 ( .A1(n11522), .A2(n11520), .ZN(n11549) );
  NAND2_X1 U11580 ( .A1(n11520), .A2(n11522), .ZN(n11546) );
  NAND2_X1 U11581 ( .A1(n11550), .A2(n11551), .ZN(n11522) );
  NAND2_X1 U11582 ( .A1(n11552), .A2(b_15_), .ZN(n11551) );
  NOR2_X1 U11583 ( .A1(n11553), .A2(n7682), .ZN(n11552) );
  NOR2_X1 U11584 ( .A1(n11518), .A2(n11516), .ZN(n11553) );
  NAND2_X1 U11585 ( .A1(n11516), .A2(n11518), .ZN(n11550) );
  NAND2_X1 U11586 ( .A1(n11554), .A2(n11555), .ZN(n11518) );
  NAND2_X1 U11587 ( .A1(n11556), .A2(b_15_), .ZN(n11555) );
  NOR2_X1 U11588 ( .A1(n11557), .A2(n7455), .ZN(n11556) );
  NOR2_X1 U11589 ( .A1(n11512), .A2(n11514), .ZN(n11557) );
  NAND2_X1 U11590 ( .A1(n11512), .A2(n11514), .ZN(n11554) );
  NAND2_X1 U11591 ( .A1(n11558), .A2(n11559), .ZN(n11514) );
  NAND2_X1 U11592 ( .A1(n11560), .A2(b_15_), .ZN(n11559) );
  NOR2_X1 U11593 ( .A1(n11561), .A2(n7450), .ZN(n11560) );
  NOR2_X1 U11594 ( .A1(n11510), .A2(n11509), .ZN(n11561) );
  NAND2_X1 U11595 ( .A1(n11509), .A2(n11510), .ZN(n11558) );
  NAND2_X1 U11596 ( .A1(n11562), .A2(n11563), .ZN(n11510) );
  NAND2_X1 U11597 ( .A1(n11564), .A2(b_15_), .ZN(n11563) );
  NOR2_X1 U11598 ( .A1(n11565), .A2(n7445), .ZN(n11564) );
  NOR2_X1 U11599 ( .A1(n11506), .A2(n11505), .ZN(n11565) );
  NAND2_X1 U11600 ( .A1(n11505), .A2(n11506), .ZN(n11562) );
  NAND2_X1 U11601 ( .A1(n11566), .A2(n11567), .ZN(n11506) );
  NAND2_X1 U11602 ( .A1(n11568), .A2(b_15_), .ZN(n11567) );
  NOR2_X1 U11603 ( .A1(n11569), .A2(n7699), .ZN(n11568) );
  NOR2_X1 U11604 ( .A1(n11502), .A2(n11501), .ZN(n11569) );
  NAND2_X1 U11605 ( .A1(n11501), .A2(n11502), .ZN(n11566) );
  NAND2_X1 U11606 ( .A1(n11570), .A2(n11571), .ZN(n11502) );
  NAND2_X1 U11607 ( .A1(n11572), .A2(b_15_), .ZN(n11571) );
  NOR2_X1 U11608 ( .A1(n11573), .A2(n7704), .ZN(n11572) );
  NOR2_X1 U11609 ( .A1(n11498), .A2(n11496), .ZN(n11573) );
  NAND2_X1 U11610 ( .A1(n11496), .A2(n11498), .ZN(n11570) );
  NAND2_X1 U11611 ( .A1(n11574), .A2(n11575), .ZN(n11498) );
  NAND2_X1 U11612 ( .A1(n11576), .A2(b_15_), .ZN(n11575) );
  NOR2_X1 U11613 ( .A1(n11577), .A2(n7709), .ZN(n11576) );
  NOR2_X1 U11614 ( .A1(n11341), .A2(n11340), .ZN(n11577) );
  NAND2_X1 U11615 ( .A1(n11340), .A2(n11341), .ZN(n11574) );
  NAND2_X1 U11616 ( .A1(n11578), .A2(n11579), .ZN(n11341) );
  NAND2_X1 U11617 ( .A1(n11580), .A2(b_15_), .ZN(n11579) );
  NOR2_X1 U11618 ( .A1(n11581), .A2(n7424), .ZN(n11580) );
  NOR2_X1 U11619 ( .A1(n11494), .A2(n11492), .ZN(n11581) );
  NAND2_X1 U11620 ( .A1(n11492), .A2(n11494), .ZN(n11578) );
  NAND2_X1 U11621 ( .A1(n11582), .A2(n11583), .ZN(n11494) );
  NAND2_X1 U11622 ( .A1(n11584), .A2(b_15_), .ZN(n11583) );
  NOR2_X1 U11623 ( .A1(n11585), .A2(n7718), .ZN(n11584) );
  NOR2_X1 U11624 ( .A1(n11490), .A2(n11488), .ZN(n11585) );
  NAND2_X1 U11625 ( .A1(n11488), .A2(n11490), .ZN(n11582) );
  NAND2_X1 U11626 ( .A1(n11586), .A2(n11587), .ZN(n11490) );
  NAND2_X1 U11627 ( .A1(n11588), .A2(b_15_), .ZN(n11587) );
  NOR2_X1 U11628 ( .A1(n11589), .A2(n7415), .ZN(n11588) );
  NOR2_X1 U11629 ( .A1(n11486), .A2(n11485), .ZN(n11589) );
  NAND2_X1 U11630 ( .A1(n11485), .A2(n11486), .ZN(n11586) );
  NAND2_X1 U11631 ( .A1(n11590), .A2(n11591), .ZN(n11486) );
  NAND2_X1 U11632 ( .A1(n11592), .A2(b_15_), .ZN(n11591) );
  NOR2_X1 U11633 ( .A1(n11593), .A2(n7727), .ZN(n11592) );
  NOR2_X1 U11634 ( .A1(n11481), .A2(n11483), .ZN(n11593) );
  NAND2_X1 U11635 ( .A1(n11481), .A2(n11483), .ZN(n11590) );
  NAND2_X1 U11636 ( .A1(n11594), .A2(n11595), .ZN(n11483) );
  NAND2_X1 U11637 ( .A1(n11477), .A2(n11596), .ZN(n11595) );
  OR2_X1 U11638 ( .A1(n11478), .A2(n11479), .ZN(n11596) );
  XNOR2_X1 U11639 ( .A(n11597), .B(n11598), .ZN(n11477) );
  XNOR2_X1 U11640 ( .A(n11599), .B(n11600), .ZN(n11597) );
  NAND2_X1 U11641 ( .A1(n11479), .A2(n11478), .ZN(n11594) );
  NAND2_X1 U11642 ( .A1(n11601), .A2(n11602), .ZN(n11478) );
  NAND2_X1 U11643 ( .A1(n11475), .A2(n11603), .ZN(n11602) );
  OR2_X1 U11644 ( .A1(n11473), .A2(n11474), .ZN(n11603) );
  NOR2_X1 U11645 ( .A1(n11175), .A2(n7736), .ZN(n11475) );
  NAND2_X1 U11646 ( .A1(n11473), .A2(n11474), .ZN(n11601) );
  NAND2_X1 U11647 ( .A1(n11604), .A2(n11605), .ZN(n11474) );
  NAND2_X1 U11648 ( .A1(n11471), .A2(n11606), .ZN(n11605) );
  OR2_X1 U11649 ( .A1(n11469), .A2(n11470), .ZN(n11606) );
  NOR2_X1 U11650 ( .A1(n11175), .A2(n7397), .ZN(n11471) );
  NAND2_X1 U11651 ( .A1(n11469), .A2(n11470), .ZN(n11604) );
  NAND2_X1 U11652 ( .A1(n11607), .A2(n11608), .ZN(n11470) );
  NAND2_X1 U11653 ( .A1(n11609), .A2(b_15_), .ZN(n11608) );
  NOR2_X1 U11654 ( .A1(n11610), .A2(n7745), .ZN(n11609) );
  NOR2_X1 U11655 ( .A1(n11465), .A2(n11466), .ZN(n11610) );
  NAND2_X1 U11656 ( .A1(n11465), .A2(n11466), .ZN(n11607) );
  NAND2_X1 U11657 ( .A1(n11611), .A2(n11612), .ZN(n11466) );
  NAND2_X1 U11658 ( .A1(n11463), .A2(n11613), .ZN(n11612) );
  OR2_X1 U11659 ( .A1(n11461), .A2(n11462), .ZN(n11613) );
  NOR2_X1 U11660 ( .A1(n11175), .A2(n7750), .ZN(n11463) );
  NAND2_X1 U11661 ( .A1(n11461), .A2(n11462), .ZN(n11611) );
  NAND2_X1 U11662 ( .A1(n11614), .A2(n11615), .ZN(n11462) );
  NAND2_X1 U11663 ( .A1(n11616), .A2(b_15_), .ZN(n11615) );
  NOR2_X1 U11664 ( .A1(n11617), .A2(n7755), .ZN(n11616) );
  NOR2_X1 U11665 ( .A1(n11457), .A2(n11458), .ZN(n11617) );
  NAND2_X1 U11666 ( .A1(n11457), .A2(n11458), .ZN(n11614) );
  NAND2_X1 U11667 ( .A1(n11618), .A2(n11619), .ZN(n11458) );
  NAND2_X1 U11668 ( .A1(n11455), .A2(n11620), .ZN(n11619) );
  OR2_X1 U11669 ( .A1(n11453), .A2(n11454), .ZN(n11620) );
  NOR2_X1 U11670 ( .A1(n11175), .A2(n7760), .ZN(n11455) );
  NAND2_X1 U11671 ( .A1(n11453), .A2(n11454), .ZN(n11618) );
  NAND2_X1 U11672 ( .A1(n11621), .A2(n11622), .ZN(n11454) );
  NAND2_X1 U11673 ( .A1(n11623), .A2(b_15_), .ZN(n11622) );
  NOR2_X1 U11674 ( .A1(n11624), .A2(n7765), .ZN(n11623) );
  NOR2_X1 U11675 ( .A1(n11449), .A2(n11450), .ZN(n11624) );
  NAND2_X1 U11676 ( .A1(n11449), .A2(n11450), .ZN(n11621) );
  NAND2_X1 U11677 ( .A1(n11625), .A2(n11626), .ZN(n11450) );
  NAND2_X1 U11678 ( .A1(n11447), .A2(n11627), .ZN(n11626) );
  OR2_X1 U11679 ( .A1(n11445), .A2(n11446), .ZN(n11627) );
  NOR2_X1 U11680 ( .A1(n11175), .A2(n8014), .ZN(n11447) );
  NAND2_X1 U11681 ( .A1(n11445), .A2(n11446), .ZN(n11625) );
  NAND2_X1 U11682 ( .A1(n11628), .A2(n11629), .ZN(n11446) );
  NAND2_X1 U11683 ( .A1(n11630), .A2(b_15_), .ZN(n11629) );
  NOR2_X1 U11684 ( .A1(n11631), .A2(n7774), .ZN(n11630) );
  NOR2_X1 U11685 ( .A1(n11441), .A2(n11442), .ZN(n11631) );
  NAND2_X1 U11686 ( .A1(n11441), .A2(n11442), .ZN(n11628) );
  NAND2_X1 U11687 ( .A1(n11632), .A2(n11633), .ZN(n11442) );
  NAND2_X1 U11688 ( .A1(n11439), .A2(n11634), .ZN(n11633) );
  OR2_X1 U11689 ( .A1(n11437), .A2(n11438), .ZN(n11634) );
  NOR2_X1 U11690 ( .A1(n11175), .A2(n8022), .ZN(n11439) );
  NAND2_X1 U11691 ( .A1(n11437), .A2(n11438), .ZN(n11632) );
  NAND2_X1 U11692 ( .A1(n11434), .A2(n11635), .ZN(n11438) );
  NAND2_X1 U11693 ( .A1(n11433), .A2(n11435), .ZN(n11635) );
  NAND2_X1 U11694 ( .A1(n11636), .A2(n11637), .ZN(n11435) );
  NAND2_X1 U11695 ( .A1(b_15_), .A2(a_26_), .ZN(n11637) );
  INV_X1 U11696 ( .A(n11638), .ZN(n11636) );
  XNOR2_X1 U11697 ( .A(n11639), .B(n11640), .ZN(n11433) );
  NAND2_X1 U11698 ( .A1(n11641), .A2(n11642), .ZN(n11639) );
  NAND2_X1 U11699 ( .A1(a_26_), .A2(n11638), .ZN(n11434) );
  NAND2_X1 U11700 ( .A1(n11403), .A2(n11643), .ZN(n11638) );
  NAND2_X1 U11701 ( .A1(n11402), .A2(n11404), .ZN(n11643) );
  NAND2_X1 U11702 ( .A1(n11644), .A2(n11645), .ZN(n11404) );
  NAND2_X1 U11703 ( .A1(b_15_), .A2(a_27_), .ZN(n11645) );
  INV_X1 U11704 ( .A(n11646), .ZN(n11644) );
  XNOR2_X1 U11705 ( .A(n11647), .B(n11648), .ZN(n11402) );
  XOR2_X1 U11706 ( .A(n11649), .B(n11650), .Z(n11648) );
  NAND2_X1 U11707 ( .A1(b_14_), .A2(a_28_), .ZN(n11650) );
  NAND2_X1 U11708 ( .A1(a_27_), .A2(n11646), .ZN(n11403) );
  NAND2_X1 U11709 ( .A1(n11651), .A2(n11652), .ZN(n11646) );
  NAND2_X1 U11710 ( .A1(n11653), .A2(b_15_), .ZN(n11652) );
  NOR2_X1 U11711 ( .A1(n11654), .A2(n7803), .ZN(n11653) );
  NOR2_X1 U11712 ( .A1(n11409), .A2(n11411), .ZN(n11654) );
  NAND2_X1 U11713 ( .A1(n11409), .A2(n11411), .ZN(n11651) );
  NAND2_X1 U11714 ( .A1(n11655), .A2(n11656), .ZN(n11411) );
  NAND2_X1 U11715 ( .A1(n11429), .A2(n11657), .ZN(n11656) );
  NAND2_X1 U11716 ( .A1(n11431), .A2(n11430), .ZN(n11657) );
  NOR2_X1 U11717 ( .A1(n11175), .A2(n7337), .ZN(n11429) );
  OR2_X1 U11718 ( .A1(n11430), .A2(n11431), .ZN(n11655) );
  AND2_X1 U11719 ( .A1(n11658), .A2(n11659), .ZN(n11431) );
  NAND2_X1 U11720 ( .A1(n11660), .A2(b_13_), .ZN(n11659) );
  NOR2_X1 U11721 ( .A1(n11661), .A2(n7817), .ZN(n11660) );
  NOR2_X1 U11722 ( .A1(n7816), .A2(n11426), .ZN(n11661) );
  NAND2_X1 U11723 ( .A1(n11662), .A2(b_14_), .ZN(n11658) );
  NOR2_X1 U11724 ( .A1(n11663), .A2(n8052), .ZN(n11662) );
  NOR2_X1 U11725 ( .A1(n7810), .A2(n11664), .ZN(n11663) );
  NAND2_X1 U11726 ( .A1(n11665), .A2(b_15_), .ZN(n11430) );
  NOR2_X1 U11727 ( .A1(n8055), .A2(n11426), .ZN(n11665) );
  XOR2_X1 U11728 ( .A(n11666), .B(n11667), .Z(n11409) );
  XOR2_X1 U11729 ( .A(n11668), .B(n11669), .Z(n11666) );
  XNOR2_X1 U11730 ( .A(n11670), .B(n11671), .ZN(n11437) );
  NAND2_X1 U11731 ( .A1(n11672), .A2(n11673), .ZN(n11670) );
  XOR2_X1 U11732 ( .A(n11674), .B(n11675), .Z(n11441) );
  XOR2_X1 U11733 ( .A(n11676), .B(n11677), .Z(n11674) );
  XOR2_X1 U11734 ( .A(n11678), .B(n11679), .Z(n11445) );
  XNOR2_X1 U11735 ( .A(n11680), .B(n11681), .ZN(n11678) );
  NAND2_X1 U11736 ( .A1(b_14_), .A2(a_24_), .ZN(n11680) );
  XOR2_X1 U11737 ( .A(n11682), .B(n11683), .Z(n11449) );
  XOR2_X1 U11738 ( .A(n11684), .B(n11685), .Z(n11682) );
  XNOR2_X1 U11739 ( .A(n11686), .B(n11687), .ZN(n11453) );
  XOR2_X1 U11740 ( .A(n11688), .B(n11689), .Z(n11687) );
  NAND2_X1 U11741 ( .A1(b_14_), .A2(a_22_), .ZN(n11689) );
  XOR2_X1 U11742 ( .A(n11690), .B(n11691), .Z(n11457) );
  XOR2_X1 U11743 ( .A(n11692), .B(n11693), .Z(n11690) );
  XOR2_X1 U11744 ( .A(n11694), .B(n11695), .Z(n11461) );
  XOR2_X1 U11745 ( .A(n11696), .B(n11697), .Z(n11694) );
  NOR2_X1 U11746 ( .A1(n7755), .A2(n11426), .ZN(n11697) );
  XNOR2_X1 U11747 ( .A(n11698), .B(n11699), .ZN(n11465) );
  XNOR2_X1 U11748 ( .A(n11700), .B(n11701), .ZN(n11699) );
  XOR2_X1 U11749 ( .A(n11702), .B(n11703), .Z(n11469) );
  XOR2_X1 U11750 ( .A(n11704), .B(n11705), .Z(n11702) );
  NOR2_X1 U11751 ( .A1(n7745), .A2(n11426), .ZN(n11705) );
  XOR2_X1 U11752 ( .A(n11706), .B(n11707), .Z(n11473) );
  XOR2_X1 U11753 ( .A(n11708), .B(n11709), .Z(n11706) );
  NOR2_X1 U11754 ( .A1(n7397), .A2(n11426), .ZN(n11709) );
  XOR2_X1 U11755 ( .A(n11710), .B(n11711), .Z(n11481) );
  XOR2_X1 U11756 ( .A(n11712), .B(n11713), .Z(n11710) );
  XNOR2_X1 U11757 ( .A(n11714), .B(n11715), .ZN(n11485) );
  XOR2_X1 U11758 ( .A(n11716), .B(n11717), .Z(n11715) );
  XOR2_X1 U11759 ( .A(n11718), .B(n11719), .Z(n11488) );
  XNOR2_X1 U11760 ( .A(n11720), .B(n11721), .ZN(n11719) );
  NAND2_X1 U11761 ( .A1(b_14_), .A2(a_13_), .ZN(n11721) );
  XNOR2_X1 U11762 ( .A(n11722), .B(n11723), .ZN(n11492) );
  NAND2_X1 U11763 ( .A1(n11724), .A2(n11725), .ZN(n11722) );
  XNOR2_X1 U11764 ( .A(n11726), .B(n11727), .ZN(n11340) );
  NAND2_X1 U11765 ( .A1(n11728), .A2(n11729), .ZN(n11726) );
  XNOR2_X1 U11766 ( .A(n11730), .B(n11731), .ZN(n11496) );
  NAND2_X1 U11767 ( .A1(n11732), .A2(n11733), .ZN(n11730) );
  XNOR2_X1 U11768 ( .A(n11734), .B(n11735), .ZN(n11501) );
  XNOR2_X1 U11769 ( .A(n11736), .B(n11737), .ZN(n11735) );
  XOR2_X1 U11770 ( .A(n11738), .B(n11739), .Z(n11505) );
  XOR2_X1 U11771 ( .A(n11740), .B(n11741), .Z(n11738) );
  NOR2_X1 U11772 ( .A1(n7699), .A2(n11426), .ZN(n11741) );
  XNOR2_X1 U11773 ( .A(n11742), .B(n11743), .ZN(n11509) );
  NAND2_X1 U11774 ( .A1(n11744), .A2(n11745), .ZN(n11742) );
  XNOR2_X1 U11775 ( .A(n11746), .B(n11747), .ZN(n11512) );
  NAND2_X1 U11776 ( .A1(n11748), .A2(n11749), .ZN(n11746) );
  XNOR2_X1 U11777 ( .A(n11750), .B(n11751), .ZN(n11516) );
  XNOR2_X1 U11778 ( .A(n11752), .B(n11753), .ZN(n11750) );
  XOR2_X1 U11779 ( .A(n11754), .B(n11755), .Z(n11520) );
  XNOR2_X1 U11780 ( .A(n11756), .B(n11757), .ZN(n11754) );
  NAND2_X1 U11781 ( .A1(b_14_), .A2(a_4_), .ZN(n11756) );
  XNOR2_X1 U11782 ( .A(n11758), .B(n11759), .ZN(n11309) );
  NAND2_X1 U11783 ( .A1(n11760), .A2(n11761), .ZN(n11758) );
  XNOR2_X1 U11784 ( .A(n11762), .B(n11763), .ZN(n11293) );
  NAND2_X1 U11785 ( .A1(n11764), .A2(n11765), .ZN(n11762) );
  NOR2_X1 U11786 ( .A1(n11766), .A2(n11288), .ZN(n11528) );
  INV_X1 U11787 ( .A(n11291), .ZN(n11288) );
  XNOR2_X1 U11788 ( .A(n11767), .B(n11768), .ZN(n11291) );
  NAND2_X1 U11789 ( .A1(n11769), .A2(n11770), .ZN(n11767) );
  NOR2_X1 U11790 ( .A1(n11526), .A2(n11527), .ZN(n11766) );
  OR2_X1 U11791 ( .A1(n7596), .A2(n7595), .ZN(n7559) );
  NAND2_X1 U11792 ( .A1(n7591), .A2(n11771), .ZN(n7595) );
  NAND2_X1 U11793 ( .A1(n11772), .A2(n11773), .ZN(n11771) );
  INV_X1 U11794 ( .A(n11774), .ZN(n11773) );
  XOR2_X1 U11795 ( .A(n11775), .B(n11776), .Z(n11772) );
  NAND2_X1 U11796 ( .A1(n11526), .A2(n11527), .ZN(n7596) );
  NAND2_X1 U11797 ( .A1(n11769), .A2(n11777), .ZN(n11527) );
  NAND2_X1 U11798 ( .A1(n11768), .A2(n11770), .ZN(n11777) );
  NAND2_X1 U11799 ( .A1(n11778), .A2(n11779), .ZN(n11770) );
  NAND2_X1 U11800 ( .A1(b_14_), .A2(a_0_), .ZN(n11779) );
  INV_X1 U11801 ( .A(n11780), .ZN(n11778) );
  XNOR2_X1 U11802 ( .A(n11781), .B(n11782), .ZN(n11768) );
  XOR2_X1 U11803 ( .A(n11783), .B(n11784), .Z(n11782) );
  NAND2_X1 U11804 ( .A1(b_13_), .A2(a_1_), .ZN(n11784) );
  NAND2_X1 U11805 ( .A1(a_0_), .A2(n11780), .ZN(n11769) );
  NAND2_X1 U11806 ( .A1(n11764), .A2(n11785), .ZN(n11780) );
  NAND2_X1 U11807 ( .A1(n11763), .A2(n11765), .ZN(n11785) );
  NAND2_X1 U11808 ( .A1(n11786), .A2(n11787), .ZN(n11765) );
  NAND2_X1 U11809 ( .A1(b_14_), .A2(a_1_), .ZN(n11787) );
  INV_X1 U11810 ( .A(n11788), .ZN(n11786) );
  XNOR2_X1 U11811 ( .A(n11789), .B(n11790), .ZN(n11763) );
  XOR2_X1 U11812 ( .A(n11791), .B(n11792), .Z(n11790) );
  NAND2_X1 U11813 ( .A1(b_13_), .A2(a_2_), .ZN(n11792) );
  NAND2_X1 U11814 ( .A1(a_1_), .A2(n11788), .ZN(n11764) );
  NAND2_X1 U11815 ( .A1(n11540), .A2(n11793), .ZN(n11788) );
  NAND2_X1 U11816 ( .A1(n11539), .A2(n11541), .ZN(n11793) );
  NAND2_X1 U11817 ( .A1(n11794), .A2(n11795), .ZN(n11541) );
  NAND2_X1 U11818 ( .A1(b_14_), .A2(a_2_), .ZN(n11795) );
  INV_X1 U11819 ( .A(n11796), .ZN(n11794) );
  XNOR2_X1 U11820 ( .A(n11797), .B(n11798), .ZN(n11539) );
  XOR2_X1 U11821 ( .A(n11799), .B(n11800), .Z(n11798) );
  NAND2_X1 U11822 ( .A1(b_13_), .A2(a_3_), .ZN(n11800) );
  NAND2_X1 U11823 ( .A1(a_2_), .A2(n11796), .ZN(n11540) );
  NAND2_X1 U11824 ( .A1(n11760), .A2(n11801), .ZN(n11796) );
  NAND2_X1 U11825 ( .A1(n11759), .A2(n11761), .ZN(n11801) );
  NAND2_X1 U11826 ( .A1(n11802), .A2(n11803), .ZN(n11761) );
  NAND2_X1 U11827 ( .A1(b_14_), .A2(a_3_), .ZN(n11803) );
  INV_X1 U11828 ( .A(n11804), .ZN(n11802) );
  XNOR2_X1 U11829 ( .A(n11805), .B(n11806), .ZN(n11759) );
  XOR2_X1 U11830 ( .A(n11807), .B(n11808), .Z(n11806) );
  NAND2_X1 U11831 ( .A1(b_13_), .A2(a_4_), .ZN(n11808) );
  NAND2_X1 U11832 ( .A1(a_3_), .A2(n11804), .ZN(n11760) );
  NAND2_X1 U11833 ( .A1(n11809), .A2(n11810), .ZN(n11804) );
  NAND2_X1 U11834 ( .A1(n11811), .A2(b_14_), .ZN(n11810) );
  NOR2_X1 U11835 ( .A1(n11812), .A2(n7682), .ZN(n11811) );
  NOR2_X1 U11836 ( .A1(n11755), .A2(n11757), .ZN(n11812) );
  NAND2_X1 U11837 ( .A1(n11755), .A2(n11757), .ZN(n11809) );
  NAND2_X1 U11838 ( .A1(n11813), .A2(n11814), .ZN(n11757) );
  NAND2_X1 U11839 ( .A1(n11753), .A2(n11815), .ZN(n11814) );
  NAND2_X1 U11840 ( .A1(n11752), .A2(n11751), .ZN(n11815) );
  NOR2_X1 U11841 ( .A1(n11426), .A2(n7455), .ZN(n11753) );
  OR2_X1 U11842 ( .A1(n11751), .A2(n11752), .ZN(n11813) );
  AND2_X1 U11843 ( .A1(n11748), .A2(n11816), .ZN(n11752) );
  NAND2_X1 U11844 ( .A1(n11747), .A2(n11749), .ZN(n11816) );
  NAND2_X1 U11845 ( .A1(n11817), .A2(n11818), .ZN(n11749) );
  NAND2_X1 U11846 ( .A1(b_14_), .A2(a_6_), .ZN(n11818) );
  INV_X1 U11847 ( .A(n11819), .ZN(n11817) );
  XNOR2_X1 U11848 ( .A(n11820), .B(n11821), .ZN(n11747) );
  XOR2_X1 U11849 ( .A(n11822), .B(n11823), .Z(n11821) );
  NAND2_X1 U11850 ( .A1(b_13_), .A2(a_7_), .ZN(n11823) );
  NAND2_X1 U11851 ( .A1(a_6_), .A2(n11819), .ZN(n11748) );
  NAND2_X1 U11852 ( .A1(n11744), .A2(n11824), .ZN(n11819) );
  NAND2_X1 U11853 ( .A1(n11743), .A2(n11745), .ZN(n11824) );
  NAND2_X1 U11854 ( .A1(n11825), .A2(n11826), .ZN(n11745) );
  NAND2_X1 U11855 ( .A1(b_14_), .A2(a_7_), .ZN(n11826) );
  INV_X1 U11856 ( .A(n11827), .ZN(n11825) );
  XNOR2_X1 U11857 ( .A(n11828), .B(n11829), .ZN(n11743) );
  XOR2_X1 U11858 ( .A(n11830), .B(n11831), .Z(n11829) );
  NAND2_X1 U11859 ( .A1(b_13_), .A2(a_8_), .ZN(n11831) );
  NAND2_X1 U11860 ( .A1(a_7_), .A2(n11827), .ZN(n11744) );
  NAND2_X1 U11861 ( .A1(n11832), .A2(n11833), .ZN(n11827) );
  NAND2_X1 U11862 ( .A1(n11834), .A2(b_14_), .ZN(n11833) );
  NOR2_X1 U11863 ( .A1(n11835), .A2(n7699), .ZN(n11834) );
  NOR2_X1 U11864 ( .A1(n11739), .A2(n11740), .ZN(n11835) );
  NAND2_X1 U11865 ( .A1(n11739), .A2(n11740), .ZN(n11832) );
  NAND2_X1 U11866 ( .A1(n11836), .A2(n11837), .ZN(n11740) );
  NAND2_X1 U11867 ( .A1(n11737), .A2(n11838), .ZN(n11837) );
  OR2_X1 U11868 ( .A1(n11736), .A2(n11734), .ZN(n11838) );
  NOR2_X1 U11869 ( .A1(n11426), .A2(n7704), .ZN(n11737) );
  NAND2_X1 U11870 ( .A1(n11734), .A2(n11736), .ZN(n11836) );
  NAND2_X1 U11871 ( .A1(n11732), .A2(n11839), .ZN(n11736) );
  NAND2_X1 U11872 ( .A1(n11731), .A2(n11733), .ZN(n11839) );
  NAND2_X1 U11873 ( .A1(n11840), .A2(n11841), .ZN(n11733) );
  NAND2_X1 U11874 ( .A1(b_14_), .A2(a_10_), .ZN(n11841) );
  INV_X1 U11875 ( .A(n11842), .ZN(n11840) );
  XNOR2_X1 U11876 ( .A(n11843), .B(n11844), .ZN(n11731) );
  XOR2_X1 U11877 ( .A(n11845), .B(n11846), .Z(n11844) );
  NAND2_X1 U11878 ( .A1(b_13_), .A2(a_11_), .ZN(n11846) );
  NAND2_X1 U11879 ( .A1(a_10_), .A2(n11842), .ZN(n11732) );
  NAND2_X1 U11880 ( .A1(n11728), .A2(n11847), .ZN(n11842) );
  NAND2_X1 U11881 ( .A1(n11727), .A2(n11729), .ZN(n11847) );
  NAND2_X1 U11882 ( .A1(n11848), .A2(n11849), .ZN(n11729) );
  NAND2_X1 U11883 ( .A1(b_14_), .A2(a_11_), .ZN(n11849) );
  INV_X1 U11884 ( .A(n11850), .ZN(n11848) );
  XOR2_X1 U11885 ( .A(n11851), .B(n11852), .Z(n11727) );
  XNOR2_X1 U11886 ( .A(n11853), .B(n11854), .ZN(n11851) );
  NAND2_X1 U11887 ( .A1(b_13_), .A2(a_12_), .ZN(n11853) );
  NAND2_X1 U11888 ( .A1(a_11_), .A2(n11850), .ZN(n11728) );
  NAND2_X1 U11889 ( .A1(n11724), .A2(n11855), .ZN(n11850) );
  NAND2_X1 U11890 ( .A1(n11723), .A2(n11725), .ZN(n11855) );
  NAND2_X1 U11891 ( .A1(n11856), .A2(n11857), .ZN(n11725) );
  NAND2_X1 U11892 ( .A1(b_14_), .A2(a_12_), .ZN(n11857) );
  INV_X1 U11893 ( .A(n11858), .ZN(n11856) );
  XOR2_X1 U11894 ( .A(n11859), .B(n11860), .Z(n11723) );
  XOR2_X1 U11895 ( .A(n11861), .B(n11862), .Z(n11859) );
  NAND2_X1 U11896 ( .A1(a_12_), .A2(n11858), .ZN(n11724) );
  NAND2_X1 U11897 ( .A1(n11863), .A2(n11864), .ZN(n11858) );
  NAND2_X1 U11898 ( .A1(n11865), .A2(b_14_), .ZN(n11864) );
  NOR2_X1 U11899 ( .A1(n11866), .A2(n7415), .ZN(n11865) );
  NOR2_X1 U11900 ( .A1(n11720), .A2(n11718), .ZN(n11866) );
  NAND2_X1 U11901 ( .A1(n11720), .A2(n11718), .ZN(n11863) );
  XOR2_X1 U11902 ( .A(n11867), .B(n11868), .Z(n11718) );
  XOR2_X1 U11903 ( .A(n11869), .B(n11870), .Z(n11867) );
  NOR2_X1 U11904 ( .A1(n7727), .A2(n11664), .ZN(n11870) );
  AND2_X1 U11905 ( .A1(n11871), .A2(n11872), .ZN(n11720) );
  NAND2_X1 U11906 ( .A1(n11873), .A2(n11717), .ZN(n11872) );
  NAND2_X1 U11907 ( .A1(n11714), .A2(n11716), .ZN(n11873) );
  OR2_X1 U11908 ( .A1(n11716), .A2(n11714), .ZN(n11871) );
  XOR2_X1 U11909 ( .A(n11874), .B(n11875), .Z(n11714) );
  XOR2_X1 U11910 ( .A(n11876), .B(n11877), .Z(n11874) );
  NOR2_X1 U11911 ( .A1(n7406), .A2(n11664), .ZN(n11877) );
  NAND2_X1 U11912 ( .A1(n11878), .A2(n11879), .ZN(n11716) );
  NAND2_X1 U11913 ( .A1(n11713), .A2(n11880), .ZN(n11879) );
  OR2_X1 U11914 ( .A1(n11712), .A2(n11711), .ZN(n11880) );
  NOR2_X1 U11915 ( .A1(n11426), .A2(n7406), .ZN(n11713) );
  NAND2_X1 U11916 ( .A1(n11711), .A2(n11712), .ZN(n11878) );
  NAND2_X1 U11917 ( .A1(n11881), .A2(n11882), .ZN(n11712) );
  NAND2_X1 U11918 ( .A1(n11600), .A2(n11883), .ZN(n11882) );
  NAND2_X1 U11919 ( .A1(n11599), .A2(n11598), .ZN(n11883) );
  NOR2_X1 U11920 ( .A1(n11426), .A2(n7736), .ZN(n11600) );
  OR2_X1 U11921 ( .A1(n11598), .A2(n11599), .ZN(n11881) );
  AND2_X1 U11922 ( .A1(n11884), .A2(n11885), .ZN(n11599) );
  NAND2_X1 U11923 ( .A1(n11886), .A2(b_14_), .ZN(n11885) );
  NOR2_X1 U11924 ( .A1(n11887), .A2(n7397), .ZN(n11886) );
  NOR2_X1 U11925 ( .A1(n11707), .A2(n11708), .ZN(n11887) );
  NAND2_X1 U11926 ( .A1(n11707), .A2(n11708), .ZN(n11884) );
  NAND2_X1 U11927 ( .A1(n11888), .A2(n11889), .ZN(n11708) );
  NAND2_X1 U11928 ( .A1(n11890), .A2(b_14_), .ZN(n11889) );
  NOR2_X1 U11929 ( .A1(n11891), .A2(n7745), .ZN(n11890) );
  NOR2_X1 U11930 ( .A1(n11703), .A2(n11704), .ZN(n11891) );
  NAND2_X1 U11931 ( .A1(n11703), .A2(n11704), .ZN(n11888) );
  NAND2_X1 U11932 ( .A1(n11892), .A2(n11893), .ZN(n11704) );
  NAND2_X1 U11933 ( .A1(n11701), .A2(n11894), .ZN(n11893) );
  OR2_X1 U11934 ( .A1(n11700), .A2(n11698), .ZN(n11894) );
  NOR2_X1 U11935 ( .A1(n11426), .A2(n7750), .ZN(n11701) );
  NAND2_X1 U11936 ( .A1(n11698), .A2(n11700), .ZN(n11892) );
  NAND2_X1 U11937 ( .A1(n11895), .A2(n11896), .ZN(n11700) );
  NAND2_X1 U11938 ( .A1(n11897), .A2(b_14_), .ZN(n11896) );
  NOR2_X1 U11939 ( .A1(n11898), .A2(n7755), .ZN(n11897) );
  NOR2_X1 U11940 ( .A1(n11695), .A2(n11696), .ZN(n11898) );
  NAND2_X1 U11941 ( .A1(n11695), .A2(n11696), .ZN(n11895) );
  NAND2_X1 U11942 ( .A1(n11899), .A2(n11900), .ZN(n11696) );
  NAND2_X1 U11943 ( .A1(n11693), .A2(n11901), .ZN(n11900) );
  OR2_X1 U11944 ( .A1(n11692), .A2(n11691), .ZN(n11901) );
  NOR2_X1 U11945 ( .A1(n11426), .A2(n7760), .ZN(n11693) );
  NAND2_X1 U11946 ( .A1(n11691), .A2(n11692), .ZN(n11899) );
  NAND2_X1 U11947 ( .A1(n11902), .A2(n11903), .ZN(n11692) );
  NAND2_X1 U11948 ( .A1(n11904), .A2(b_14_), .ZN(n11903) );
  NOR2_X1 U11949 ( .A1(n11905), .A2(n7765), .ZN(n11904) );
  NOR2_X1 U11950 ( .A1(n11686), .A2(n11688), .ZN(n11905) );
  NAND2_X1 U11951 ( .A1(n11686), .A2(n11688), .ZN(n11902) );
  NAND2_X1 U11952 ( .A1(n11906), .A2(n11907), .ZN(n11688) );
  NAND2_X1 U11953 ( .A1(n11685), .A2(n11908), .ZN(n11907) );
  OR2_X1 U11954 ( .A1(n11684), .A2(n11683), .ZN(n11908) );
  NOR2_X1 U11955 ( .A1(n11426), .A2(n8014), .ZN(n11685) );
  NAND2_X1 U11956 ( .A1(n11683), .A2(n11684), .ZN(n11906) );
  NAND2_X1 U11957 ( .A1(n11909), .A2(n11910), .ZN(n11684) );
  NAND2_X1 U11958 ( .A1(n11911), .A2(b_14_), .ZN(n11910) );
  NOR2_X1 U11959 ( .A1(n11912), .A2(n7774), .ZN(n11911) );
  NOR2_X1 U11960 ( .A1(n11679), .A2(n11681), .ZN(n11912) );
  NAND2_X1 U11961 ( .A1(n11679), .A2(n11681), .ZN(n11909) );
  NAND2_X1 U11962 ( .A1(n11913), .A2(n11914), .ZN(n11681) );
  NAND2_X1 U11963 ( .A1(n11677), .A2(n11915), .ZN(n11914) );
  OR2_X1 U11964 ( .A1(n11676), .A2(n11675), .ZN(n11915) );
  NOR2_X1 U11965 ( .A1(n11426), .A2(n8022), .ZN(n11677) );
  NAND2_X1 U11966 ( .A1(n11675), .A2(n11676), .ZN(n11913) );
  NAND2_X1 U11967 ( .A1(n11672), .A2(n11916), .ZN(n11676) );
  NAND2_X1 U11968 ( .A1(n11671), .A2(n11673), .ZN(n11916) );
  NAND2_X1 U11969 ( .A1(n11917), .A2(n11918), .ZN(n11673) );
  NAND2_X1 U11970 ( .A1(b_14_), .A2(a_26_), .ZN(n11918) );
  INV_X1 U11971 ( .A(n11919), .ZN(n11917) );
  XNOR2_X1 U11972 ( .A(n11920), .B(n11921), .ZN(n11671) );
  NAND2_X1 U11973 ( .A1(n11922), .A2(n11923), .ZN(n11920) );
  NAND2_X1 U11974 ( .A1(a_26_), .A2(n11919), .ZN(n11672) );
  NAND2_X1 U11975 ( .A1(n11641), .A2(n11924), .ZN(n11919) );
  NAND2_X1 U11976 ( .A1(n11640), .A2(n11642), .ZN(n11924) );
  NAND2_X1 U11977 ( .A1(n11925), .A2(n11926), .ZN(n11642) );
  NAND2_X1 U11978 ( .A1(b_14_), .A2(a_27_), .ZN(n11926) );
  INV_X1 U11979 ( .A(n11927), .ZN(n11925) );
  XNOR2_X1 U11980 ( .A(n11928), .B(n11929), .ZN(n11640) );
  XOR2_X1 U11981 ( .A(n11930), .B(n11931), .Z(n11929) );
  NAND2_X1 U11982 ( .A1(b_13_), .A2(a_28_), .ZN(n11931) );
  NAND2_X1 U11983 ( .A1(a_27_), .A2(n11927), .ZN(n11641) );
  NAND2_X1 U11984 ( .A1(n11932), .A2(n11933), .ZN(n11927) );
  NAND2_X1 U11985 ( .A1(n11934), .A2(b_14_), .ZN(n11933) );
  NOR2_X1 U11986 ( .A1(n11935), .A2(n7803), .ZN(n11934) );
  NOR2_X1 U11987 ( .A1(n11647), .A2(n11649), .ZN(n11935) );
  NAND2_X1 U11988 ( .A1(n11647), .A2(n11649), .ZN(n11932) );
  NAND2_X1 U11989 ( .A1(n11936), .A2(n11937), .ZN(n11649) );
  NAND2_X1 U11990 ( .A1(n11667), .A2(n11938), .ZN(n11937) );
  NAND2_X1 U11991 ( .A1(n11669), .A2(n11668), .ZN(n11938) );
  NOR2_X1 U11992 ( .A1(n11426), .A2(n7337), .ZN(n11667) );
  OR2_X1 U11993 ( .A1(n11668), .A2(n11669), .ZN(n11936) );
  AND2_X1 U11994 ( .A1(n11939), .A2(n11940), .ZN(n11669) );
  NAND2_X1 U11995 ( .A1(n11941), .A2(b_12_), .ZN(n11940) );
  NOR2_X1 U11996 ( .A1(n11942), .A2(n7817), .ZN(n11941) );
  NOR2_X1 U11997 ( .A1(n7816), .A2(n11664), .ZN(n11942) );
  NAND2_X1 U11998 ( .A1(n11943), .A2(b_13_), .ZN(n11939) );
  NOR2_X1 U11999 ( .A1(n11944), .A2(n8052), .ZN(n11943) );
  NOR2_X1 U12000 ( .A1(n7810), .A2(n11945), .ZN(n11944) );
  NAND2_X1 U12001 ( .A1(n11946), .A2(b_14_), .ZN(n11668) );
  NOR2_X1 U12002 ( .A1(n8055), .A2(n11664), .ZN(n11946) );
  XOR2_X1 U12003 ( .A(n11947), .B(n11948), .Z(n11647) );
  XOR2_X1 U12004 ( .A(n11949), .B(n11950), .Z(n11947) );
  XNOR2_X1 U12005 ( .A(n11951), .B(n11952), .ZN(n11675) );
  NAND2_X1 U12006 ( .A1(n11953), .A2(n11954), .ZN(n11951) );
  XOR2_X1 U12007 ( .A(n11955), .B(n11956), .Z(n11679) );
  XOR2_X1 U12008 ( .A(n11957), .B(n11958), .Z(n11955) );
  XOR2_X1 U12009 ( .A(n11959), .B(n11960), .Z(n11683) );
  XNOR2_X1 U12010 ( .A(n11961), .B(n11962), .ZN(n11959) );
  NAND2_X1 U12011 ( .A1(b_13_), .A2(a_24_), .ZN(n11961) );
  XOR2_X1 U12012 ( .A(n11963), .B(n11964), .Z(n11686) );
  XOR2_X1 U12013 ( .A(n11965), .B(n11966), .Z(n11963) );
  XOR2_X1 U12014 ( .A(n11967), .B(n11968), .Z(n11691) );
  XOR2_X1 U12015 ( .A(n11969), .B(n11970), .Z(n11967) );
  NOR2_X1 U12016 ( .A1(n7765), .A2(n11664), .ZN(n11970) );
  XOR2_X1 U12017 ( .A(n11971), .B(n11972), .Z(n11695) );
  XOR2_X1 U12018 ( .A(n11973), .B(n11974), .Z(n11971) );
  XOR2_X1 U12019 ( .A(n11975), .B(n11976), .Z(n11698) );
  XOR2_X1 U12020 ( .A(n11977), .B(n11978), .Z(n11975) );
  NOR2_X1 U12021 ( .A1(n7755), .A2(n11664), .ZN(n11978) );
  XOR2_X1 U12022 ( .A(n11979), .B(n11980), .Z(n11703) );
  XOR2_X1 U12023 ( .A(n11981), .B(n11982), .Z(n11979) );
  XOR2_X1 U12024 ( .A(n11983), .B(n11984), .Z(n11707) );
  XOR2_X1 U12025 ( .A(n11985), .B(n11986), .Z(n11983) );
  XOR2_X1 U12026 ( .A(n11987), .B(n11988), .Z(n11598) );
  XOR2_X1 U12027 ( .A(n11989), .B(n11990), .Z(n11988) );
  NAND2_X1 U12028 ( .A1(b_13_), .A2(a_17_), .ZN(n11990) );
  XOR2_X1 U12029 ( .A(n11991), .B(n11992), .Z(n11711) );
  XOR2_X1 U12030 ( .A(n11993), .B(n11994), .Z(n11991) );
  NOR2_X1 U12031 ( .A1(n7736), .A2(n11664), .ZN(n11994) );
  XNOR2_X1 U12032 ( .A(n11995), .B(n11996), .ZN(n11734) );
  XOR2_X1 U12033 ( .A(n11997), .B(n11998), .Z(n11996) );
  NAND2_X1 U12034 ( .A1(b_13_), .A2(a_10_), .ZN(n11998) );
  XNOR2_X1 U12035 ( .A(n11999), .B(n12000), .ZN(n11739) );
  XOR2_X1 U12036 ( .A(n12001), .B(n12002), .Z(n12000) );
  NAND2_X1 U12037 ( .A1(b_13_), .A2(a_9_), .ZN(n12002) );
  XOR2_X1 U12038 ( .A(n12003), .B(n12004), .Z(n11751) );
  XOR2_X1 U12039 ( .A(n12005), .B(n12006), .Z(n12004) );
  NAND2_X1 U12040 ( .A1(b_13_), .A2(a_6_), .ZN(n12006) );
  XNOR2_X1 U12041 ( .A(n12007), .B(n12008), .ZN(n11755) );
  XOR2_X1 U12042 ( .A(n12009), .B(n12010), .Z(n12008) );
  NAND2_X1 U12043 ( .A1(b_13_), .A2(a_5_), .ZN(n12010) );
  XNOR2_X1 U12044 ( .A(n12011), .B(n12012), .ZN(n11526) );
  XNOR2_X1 U12045 ( .A(n12013), .B(n12014), .ZN(n12012) );
  OR2_X1 U12046 ( .A1(n12015), .A2(n7591), .ZN(n7564) );
  NAND2_X1 U12047 ( .A1(n12016), .A2(n11774), .ZN(n7591) );
  NAND2_X1 U12048 ( .A1(n12017), .A2(n12018), .ZN(n11774) );
  NAND2_X1 U12049 ( .A1(n12014), .A2(n12019), .ZN(n12018) );
  OR2_X1 U12050 ( .A1(n12013), .A2(n12011), .ZN(n12019) );
  NOR2_X1 U12051 ( .A1(n11664), .A2(n7478), .ZN(n12014) );
  NAND2_X1 U12052 ( .A1(n12011), .A2(n12013), .ZN(n12017) );
  NAND2_X1 U12053 ( .A1(n12020), .A2(n12021), .ZN(n12013) );
  NAND2_X1 U12054 ( .A1(n12022), .A2(b_13_), .ZN(n12021) );
  NOR2_X1 U12055 ( .A1(n12023), .A2(n7669), .ZN(n12022) );
  NOR2_X1 U12056 ( .A1(n11781), .A2(n11783), .ZN(n12023) );
  NAND2_X1 U12057 ( .A1(n11781), .A2(n11783), .ZN(n12020) );
  NAND2_X1 U12058 ( .A1(n12024), .A2(n12025), .ZN(n11783) );
  NAND2_X1 U12059 ( .A1(n12026), .A2(b_13_), .ZN(n12025) );
  NOR2_X1 U12060 ( .A1(n12027), .A2(n7469), .ZN(n12026) );
  NOR2_X1 U12061 ( .A1(n11789), .A2(n11791), .ZN(n12027) );
  NAND2_X1 U12062 ( .A1(n11789), .A2(n11791), .ZN(n12024) );
  NAND2_X1 U12063 ( .A1(n12028), .A2(n12029), .ZN(n11791) );
  NAND2_X1 U12064 ( .A1(n12030), .A2(b_13_), .ZN(n12029) );
  NOR2_X1 U12065 ( .A1(n12031), .A2(n7464), .ZN(n12030) );
  NOR2_X1 U12066 ( .A1(n11797), .A2(n11799), .ZN(n12031) );
  NAND2_X1 U12067 ( .A1(n11797), .A2(n11799), .ZN(n12028) );
  NAND2_X1 U12068 ( .A1(n12032), .A2(n12033), .ZN(n11799) );
  NAND2_X1 U12069 ( .A1(n12034), .A2(b_13_), .ZN(n12033) );
  NOR2_X1 U12070 ( .A1(n12035), .A2(n7682), .ZN(n12034) );
  NOR2_X1 U12071 ( .A1(n11805), .A2(n11807), .ZN(n12035) );
  NAND2_X1 U12072 ( .A1(n11805), .A2(n11807), .ZN(n12032) );
  NAND2_X1 U12073 ( .A1(n12036), .A2(n12037), .ZN(n11807) );
  NAND2_X1 U12074 ( .A1(n12038), .A2(b_13_), .ZN(n12037) );
  NOR2_X1 U12075 ( .A1(n12039), .A2(n7455), .ZN(n12038) );
  NOR2_X1 U12076 ( .A1(n12007), .A2(n12009), .ZN(n12039) );
  NAND2_X1 U12077 ( .A1(n12007), .A2(n12009), .ZN(n12036) );
  NAND2_X1 U12078 ( .A1(n12040), .A2(n12041), .ZN(n12009) );
  NAND2_X1 U12079 ( .A1(n12042), .A2(b_13_), .ZN(n12041) );
  NOR2_X1 U12080 ( .A1(n12043), .A2(n7450), .ZN(n12042) );
  NOR2_X1 U12081 ( .A1(n12003), .A2(n12005), .ZN(n12043) );
  NAND2_X1 U12082 ( .A1(n12003), .A2(n12005), .ZN(n12040) );
  NAND2_X1 U12083 ( .A1(n12044), .A2(n12045), .ZN(n12005) );
  NAND2_X1 U12084 ( .A1(n12046), .A2(b_13_), .ZN(n12045) );
  NOR2_X1 U12085 ( .A1(n12047), .A2(n7445), .ZN(n12046) );
  NOR2_X1 U12086 ( .A1(n11820), .A2(n11822), .ZN(n12047) );
  NAND2_X1 U12087 ( .A1(n11820), .A2(n11822), .ZN(n12044) );
  NAND2_X1 U12088 ( .A1(n12048), .A2(n12049), .ZN(n11822) );
  NAND2_X1 U12089 ( .A1(n12050), .A2(b_13_), .ZN(n12049) );
  NOR2_X1 U12090 ( .A1(n12051), .A2(n7699), .ZN(n12050) );
  NOR2_X1 U12091 ( .A1(n11828), .A2(n11830), .ZN(n12051) );
  NAND2_X1 U12092 ( .A1(n11828), .A2(n11830), .ZN(n12048) );
  NAND2_X1 U12093 ( .A1(n12052), .A2(n12053), .ZN(n11830) );
  NAND2_X1 U12094 ( .A1(n12054), .A2(b_13_), .ZN(n12053) );
  NOR2_X1 U12095 ( .A1(n12055), .A2(n7704), .ZN(n12054) );
  NOR2_X1 U12096 ( .A1(n11999), .A2(n12001), .ZN(n12055) );
  NAND2_X1 U12097 ( .A1(n11999), .A2(n12001), .ZN(n12052) );
  NAND2_X1 U12098 ( .A1(n12056), .A2(n12057), .ZN(n12001) );
  NAND2_X1 U12099 ( .A1(n12058), .A2(b_13_), .ZN(n12057) );
  NOR2_X1 U12100 ( .A1(n12059), .A2(n7709), .ZN(n12058) );
  NOR2_X1 U12101 ( .A1(n11995), .A2(n11997), .ZN(n12059) );
  NAND2_X1 U12102 ( .A1(n11995), .A2(n11997), .ZN(n12056) );
  NAND2_X1 U12103 ( .A1(n12060), .A2(n12061), .ZN(n11997) );
  NAND2_X1 U12104 ( .A1(n12062), .A2(b_13_), .ZN(n12061) );
  NOR2_X1 U12105 ( .A1(n12063), .A2(n7424), .ZN(n12062) );
  NOR2_X1 U12106 ( .A1(n11843), .A2(n11845), .ZN(n12063) );
  NAND2_X1 U12107 ( .A1(n11843), .A2(n11845), .ZN(n12060) );
  NAND2_X1 U12108 ( .A1(n12064), .A2(n12065), .ZN(n11845) );
  NAND2_X1 U12109 ( .A1(n12066), .A2(b_13_), .ZN(n12065) );
  NOR2_X1 U12110 ( .A1(n12067), .A2(n7718), .ZN(n12066) );
  NOR2_X1 U12111 ( .A1(n11852), .A2(n11854), .ZN(n12067) );
  NAND2_X1 U12112 ( .A1(n11852), .A2(n11854), .ZN(n12064) );
  NAND2_X1 U12113 ( .A1(n12068), .A2(n12069), .ZN(n11854) );
  NAND2_X1 U12114 ( .A1(n11860), .A2(n12070), .ZN(n12069) );
  OR2_X1 U12115 ( .A1(n11861), .A2(n11862), .ZN(n12070) );
  XNOR2_X1 U12116 ( .A(n12071), .B(n12072), .ZN(n11860) );
  NAND2_X1 U12117 ( .A1(n12073), .A2(n12074), .ZN(n12071) );
  NAND2_X1 U12118 ( .A1(n11862), .A2(n11861), .ZN(n12068) );
  NAND2_X1 U12119 ( .A1(n12075), .A2(n12076), .ZN(n11861) );
  NAND2_X1 U12120 ( .A1(n12077), .A2(b_13_), .ZN(n12076) );
  NOR2_X1 U12121 ( .A1(n12078), .A2(n7727), .ZN(n12077) );
  NOR2_X1 U12122 ( .A1(n11868), .A2(n11869), .ZN(n12078) );
  NAND2_X1 U12123 ( .A1(n11868), .A2(n11869), .ZN(n12075) );
  NAND2_X1 U12124 ( .A1(n12079), .A2(n12080), .ZN(n11869) );
  NAND2_X1 U12125 ( .A1(n12081), .A2(b_13_), .ZN(n12080) );
  NOR2_X1 U12126 ( .A1(n12082), .A2(n7406), .ZN(n12081) );
  NOR2_X1 U12127 ( .A1(n11875), .A2(n11876), .ZN(n12082) );
  NAND2_X1 U12128 ( .A1(n11875), .A2(n11876), .ZN(n12079) );
  NAND2_X1 U12129 ( .A1(n12083), .A2(n12084), .ZN(n11876) );
  NAND2_X1 U12130 ( .A1(n12085), .A2(b_13_), .ZN(n12084) );
  NOR2_X1 U12131 ( .A1(n12086), .A2(n7736), .ZN(n12085) );
  NOR2_X1 U12132 ( .A1(n11992), .A2(n11993), .ZN(n12086) );
  NAND2_X1 U12133 ( .A1(n11992), .A2(n11993), .ZN(n12083) );
  NAND2_X1 U12134 ( .A1(n12087), .A2(n12088), .ZN(n11993) );
  NAND2_X1 U12135 ( .A1(n12089), .A2(b_13_), .ZN(n12088) );
  NOR2_X1 U12136 ( .A1(n12090), .A2(n7397), .ZN(n12089) );
  NOR2_X1 U12137 ( .A1(n11987), .A2(n11989), .ZN(n12090) );
  NAND2_X1 U12138 ( .A1(n11987), .A2(n11989), .ZN(n12087) );
  NAND2_X1 U12139 ( .A1(n12091), .A2(n12092), .ZN(n11989) );
  NAND2_X1 U12140 ( .A1(n11986), .A2(n12093), .ZN(n12092) );
  OR2_X1 U12141 ( .A1(n11985), .A2(n11984), .ZN(n12093) );
  NOR2_X1 U12142 ( .A1(n11664), .A2(n7745), .ZN(n11986) );
  NAND2_X1 U12143 ( .A1(n11984), .A2(n11985), .ZN(n12091) );
  NAND2_X1 U12144 ( .A1(n12094), .A2(n12095), .ZN(n11985) );
  NAND2_X1 U12145 ( .A1(n11982), .A2(n12096), .ZN(n12095) );
  OR2_X1 U12146 ( .A1(n11981), .A2(n11980), .ZN(n12096) );
  NOR2_X1 U12147 ( .A1(n11664), .A2(n7750), .ZN(n11982) );
  NAND2_X1 U12148 ( .A1(n11980), .A2(n11981), .ZN(n12094) );
  NAND2_X1 U12149 ( .A1(n12097), .A2(n12098), .ZN(n11981) );
  NAND2_X1 U12150 ( .A1(n12099), .A2(b_13_), .ZN(n12098) );
  NOR2_X1 U12151 ( .A1(n12100), .A2(n7755), .ZN(n12099) );
  NOR2_X1 U12152 ( .A1(n11976), .A2(n11977), .ZN(n12100) );
  NAND2_X1 U12153 ( .A1(n11976), .A2(n11977), .ZN(n12097) );
  NAND2_X1 U12154 ( .A1(n12101), .A2(n12102), .ZN(n11977) );
  NAND2_X1 U12155 ( .A1(n11974), .A2(n12103), .ZN(n12102) );
  OR2_X1 U12156 ( .A1(n11973), .A2(n11972), .ZN(n12103) );
  NOR2_X1 U12157 ( .A1(n11664), .A2(n7760), .ZN(n11974) );
  NAND2_X1 U12158 ( .A1(n11972), .A2(n11973), .ZN(n12101) );
  NAND2_X1 U12159 ( .A1(n12104), .A2(n12105), .ZN(n11973) );
  NAND2_X1 U12160 ( .A1(n12106), .A2(b_13_), .ZN(n12105) );
  NOR2_X1 U12161 ( .A1(n12107), .A2(n7765), .ZN(n12106) );
  NOR2_X1 U12162 ( .A1(n11968), .A2(n11969), .ZN(n12107) );
  NAND2_X1 U12163 ( .A1(n11968), .A2(n11969), .ZN(n12104) );
  NAND2_X1 U12164 ( .A1(n12108), .A2(n12109), .ZN(n11969) );
  NAND2_X1 U12165 ( .A1(n11966), .A2(n12110), .ZN(n12109) );
  OR2_X1 U12166 ( .A1(n11965), .A2(n11964), .ZN(n12110) );
  NOR2_X1 U12167 ( .A1(n11664), .A2(n8014), .ZN(n11966) );
  NAND2_X1 U12168 ( .A1(n11964), .A2(n11965), .ZN(n12108) );
  NAND2_X1 U12169 ( .A1(n12111), .A2(n12112), .ZN(n11965) );
  NAND2_X1 U12170 ( .A1(n12113), .A2(b_13_), .ZN(n12112) );
  NOR2_X1 U12171 ( .A1(n12114), .A2(n7774), .ZN(n12113) );
  NOR2_X1 U12172 ( .A1(n11960), .A2(n11962), .ZN(n12114) );
  NAND2_X1 U12173 ( .A1(n11960), .A2(n11962), .ZN(n12111) );
  NAND2_X1 U12174 ( .A1(n12115), .A2(n12116), .ZN(n11962) );
  NAND2_X1 U12175 ( .A1(n11958), .A2(n12117), .ZN(n12116) );
  OR2_X1 U12176 ( .A1(n11957), .A2(n11956), .ZN(n12117) );
  NOR2_X1 U12177 ( .A1(n11664), .A2(n8022), .ZN(n11958) );
  NAND2_X1 U12178 ( .A1(n11956), .A2(n11957), .ZN(n12115) );
  NAND2_X1 U12179 ( .A1(n11953), .A2(n12118), .ZN(n11957) );
  NAND2_X1 U12180 ( .A1(n11952), .A2(n11954), .ZN(n12118) );
  NAND2_X1 U12181 ( .A1(n12119), .A2(n12120), .ZN(n11954) );
  NAND2_X1 U12182 ( .A1(b_13_), .A2(a_26_), .ZN(n12120) );
  INV_X1 U12183 ( .A(n12121), .ZN(n12119) );
  XNOR2_X1 U12184 ( .A(n12122), .B(n12123), .ZN(n11952) );
  NAND2_X1 U12185 ( .A1(n12124), .A2(n12125), .ZN(n12122) );
  NAND2_X1 U12186 ( .A1(a_26_), .A2(n12121), .ZN(n11953) );
  NAND2_X1 U12187 ( .A1(n11922), .A2(n12126), .ZN(n12121) );
  NAND2_X1 U12188 ( .A1(n11921), .A2(n11923), .ZN(n12126) );
  NAND2_X1 U12189 ( .A1(n12127), .A2(n12128), .ZN(n11923) );
  NAND2_X1 U12190 ( .A1(b_13_), .A2(a_27_), .ZN(n12128) );
  INV_X1 U12191 ( .A(n12129), .ZN(n12127) );
  XNOR2_X1 U12192 ( .A(n12130), .B(n12131), .ZN(n11921) );
  XOR2_X1 U12193 ( .A(n12132), .B(n12133), .Z(n12131) );
  NAND2_X1 U12194 ( .A1(b_12_), .A2(a_28_), .ZN(n12133) );
  NAND2_X1 U12195 ( .A1(a_27_), .A2(n12129), .ZN(n11922) );
  NAND2_X1 U12196 ( .A1(n12134), .A2(n12135), .ZN(n12129) );
  NAND2_X1 U12197 ( .A1(n12136), .A2(b_13_), .ZN(n12135) );
  NOR2_X1 U12198 ( .A1(n12137), .A2(n7803), .ZN(n12136) );
  NOR2_X1 U12199 ( .A1(n11928), .A2(n11930), .ZN(n12137) );
  NAND2_X1 U12200 ( .A1(n11928), .A2(n11930), .ZN(n12134) );
  NAND2_X1 U12201 ( .A1(n12138), .A2(n12139), .ZN(n11930) );
  NAND2_X1 U12202 ( .A1(n11948), .A2(n12140), .ZN(n12139) );
  NAND2_X1 U12203 ( .A1(n11950), .A2(n11949), .ZN(n12140) );
  NOR2_X1 U12204 ( .A1(n11664), .A2(n7337), .ZN(n11948) );
  OR2_X1 U12205 ( .A1(n11949), .A2(n11950), .ZN(n12138) );
  AND2_X1 U12206 ( .A1(n12141), .A2(n12142), .ZN(n11950) );
  NAND2_X1 U12207 ( .A1(n12143), .A2(a_31_), .ZN(n12142) );
  NOR2_X1 U12208 ( .A1(n12144), .A2(n12145), .ZN(n12143) );
  NOR2_X1 U12209 ( .A1(n7816), .A2(n11945), .ZN(n12144) );
  NAND2_X1 U12210 ( .A1(n12146), .A2(b_12_), .ZN(n12141) );
  NOR2_X1 U12211 ( .A1(n12147), .A2(n8052), .ZN(n12146) );
  NOR2_X1 U12212 ( .A1(n7810), .A2(n12145), .ZN(n12147) );
  NAND2_X1 U12213 ( .A1(n12148), .A2(b_13_), .ZN(n11949) );
  NOR2_X1 U12214 ( .A1(n8055), .A2(n11945), .ZN(n12148) );
  XOR2_X1 U12215 ( .A(n12149), .B(n12150), .Z(n11928) );
  XOR2_X1 U12216 ( .A(n12151), .B(n12152), .Z(n12149) );
  XNOR2_X1 U12217 ( .A(n12153), .B(n12154), .ZN(n11956) );
  NAND2_X1 U12218 ( .A1(n12155), .A2(n12156), .ZN(n12153) );
  XOR2_X1 U12219 ( .A(n12157), .B(n12158), .Z(n11960) );
  XOR2_X1 U12220 ( .A(n12159), .B(n12160), .Z(n12157) );
  XOR2_X1 U12221 ( .A(n12161), .B(n12162), .Z(n11964) );
  XNOR2_X1 U12222 ( .A(n12163), .B(n12164), .ZN(n12161) );
  NAND2_X1 U12223 ( .A1(b_12_), .A2(a_24_), .ZN(n12163) );
  XOR2_X1 U12224 ( .A(n12165), .B(n12166), .Z(n11968) );
  XOR2_X1 U12225 ( .A(n12167), .B(n12168), .Z(n12165) );
  XNOR2_X1 U12226 ( .A(n12169), .B(n12170), .ZN(n11972) );
  XOR2_X1 U12227 ( .A(n12171), .B(n12172), .Z(n12170) );
  NAND2_X1 U12228 ( .A1(b_12_), .A2(a_22_), .ZN(n12172) );
  XNOR2_X1 U12229 ( .A(n12173), .B(n12174), .ZN(n11976) );
  XNOR2_X1 U12230 ( .A(n12175), .B(n12176), .ZN(n12174) );
  XOR2_X1 U12231 ( .A(n12177), .B(n12178), .Z(n11980) );
  XOR2_X1 U12232 ( .A(n12179), .B(n12180), .Z(n12177) );
  NOR2_X1 U12233 ( .A1(n7755), .A2(n11945), .ZN(n12180) );
  XOR2_X1 U12234 ( .A(n12181), .B(n12182), .Z(n11984) );
  XOR2_X1 U12235 ( .A(n12183), .B(n12184), .Z(n12181) );
  NOR2_X1 U12236 ( .A1(n7750), .A2(n11945), .ZN(n12184) );
  XNOR2_X1 U12237 ( .A(n12185), .B(n12186), .ZN(n11987) );
  XNOR2_X1 U12238 ( .A(n12187), .B(n12188), .ZN(n12185) );
  XOR2_X1 U12239 ( .A(n12189), .B(n12190), .Z(n11992) );
  XOR2_X1 U12240 ( .A(n12191), .B(n12192), .Z(n12189) );
  XNOR2_X1 U12241 ( .A(n12193), .B(n12194), .ZN(n11875) );
  XNOR2_X1 U12242 ( .A(n12195), .B(n12196), .ZN(n12193) );
  XNOR2_X1 U12243 ( .A(n12197), .B(n12198), .ZN(n11868) );
  XOR2_X1 U12244 ( .A(n12199), .B(n12200), .Z(n12198) );
  NAND2_X1 U12245 ( .A1(b_12_), .A2(a_15_), .ZN(n12200) );
  XNOR2_X1 U12246 ( .A(n12201), .B(n12202), .ZN(n11852) );
  NAND2_X1 U12247 ( .A1(n12203), .A2(n12204), .ZN(n12201) );
  XOR2_X1 U12248 ( .A(n12205), .B(n12206), .Z(n11843) );
  XOR2_X1 U12249 ( .A(n12207), .B(n12208), .Z(n12205) );
  XNOR2_X1 U12250 ( .A(n12209), .B(n12210), .ZN(n11995) );
  NAND2_X1 U12251 ( .A1(n12211), .A2(n12212), .ZN(n12209) );
  XNOR2_X1 U12252 ( .A(n12213), .B(n12214), .ZN(n11999) );
  XNOR2_X1 U12253 ( .A(n12215), .B(n12216), .ZN(n12213) );
  XNOR2_X1 U12254 ( .A(n12217), .B(n12218), .ZN(n11828) );
  XOR2_X1 U12255 ( .A(n12219), .B(n12220), .Z(n12218) );
  NAND2_X1 U12256 ( .A1(b_12_), .A2(a_9_), .ZN(n12220) );
  XNOR2_X1 U12257 ( .A(n12221), .B(n12222), .ZN(n11820) );
  NAND2_X1 U12258 ( .A1(n12223), .A2(n12224), .ZN(n12221) );
  XOR2_X1 U12259 ( .A(n12225), .B(n12226), .Z(n12003) );
  NOR2_X1 U12260 ( .A1(n12227), .A2(n12228), .ZN(n12226) );
  NOR2_X1 U12261 ( .A1(n12229), .A2(n12230), .ZN(n12227) );
  NOR2_X1 U12262 ( .A1(n7445), .A2(n11945), .ZN(n12229) );
  XNOR2_X1 U12263 ( .A(n12231), .B(n12232), .ZN(n12007) );
  NAND2_X1 U12264 ( .A1(n12233), .A2(n12234), .ZN(n12231) );
  XNOR2_X1 U12265 ( .A(n12235), .B(n12236), .ZN(n11805) );
  NAND2_X1 U12266 ( .A1(n12237), .A2(n12238), .ZN(n12235) );
  XNOR2_X1 U12267 ( .A(n12239), .B(n12240), .ZN(n11797) );
  NAND2_X1 U12268 ( .A1(n12241), .A2(n12242), .ZN(n12239) );
  XNOR2_X1 U12269 ( .A(n12243), .B(n12244), .ZN(n11789) );
  NAND2_X1 U12270 ( .A1(n12245), .A2(n12246), .ZN(n12243) );
  XNOR2_X1 U12271 ( .A(n12247), .B(n12248), .ZN(n11781) );
  XNOR2_X1 U12272 ( .A(n12249), .B(n12250), .ZN(n12248) );
  XNOR2_X1 U12273 ( .A(n12251), .B(n12252), .ZN(n12011) );
  XNOR2_X1 U12274 ( .A(n12253), .B(n12254), .ZN(n12252) );
  XOR2_X1 U12275 ( .A(n12255), .B(n11776), .Z(n12016) );
  XNOR2_X1 U12276 ( .A(n12256), .B(n12257), .ZN(n11776) );
  NOR2_X1 U12277 ( .A1(n7478), .A2(n11945), .ZN(n12257) );
  INV_X1 U12278 ( .A(n11775), .ZN(n12255) );
  NAND2_X1 U12279 ( .A1(n7588), .A2(n12258), .ZN(n12015) );
  OR2_X1 U12280 ( .A1(n7593), .A2(n7592), .ZN(n12258) );
  OR2_X1 U12281 ( .A1(n7588), .A2(n7587), .ZN(n7567) );
  NAND2_X1 U12282 ( .A1(n7585), .A2(n12259), .ZN(n7587) );
  NAND2_X1 U12283 ( .A1(n12260), .A2(n12261), .ZN(n12259) );
  INV_X1 U12284 ( .A(n12262), .ZN(n12261) );
  XOR2_X1 U12285 ( .A(n12263), .B(n12264), .Z(n12260) );
  NAND2_X1 U12286 ( .A1(n7593), .A2(n7592), .ZN(n7588) );
  NAND2_X1 U12287 ( .A1(n12265), .A2(n12266), .ZN(n7592) );
  NAND2_X1 U12288 ( .A1(n12267), .A2(b_12_), .ZN(n12266) );
  NOR2_X1 U12289 ( .A1(n12268), .A2(n7478), .ZN(n12267) );
  NOR2_X1 U12290 ( .A1(n11775), .A2(n12256), .ZN(n12268) );
  NAND2_X1 U12291 ( .A1(n11775), .A2(n12256), .ZN(n12265) );
  NAND2_X1 U12292 ( .A1(n12269), .A2(n12270), .ZN(n12256) );
  NAND2_X1 U12293 ( .A1(n12254), .A2(n12271), .ZN(n12270) );
  OR2_X1 U12294 ( .A1(n12253), .A2(n12251), .ZN(n12271) );
  NOR2_X1 U12295 ( .A1(n11945), .A2(n7669), .ZN(n12254) );
  NAND2_X1 U12296 ( .A1(n12251), .A2(n12253), .ZN(n12269) );
  NAND2_X1 U12297 ( .A1(n12272), .A2(n12273), .ZN(n12253) );
  NAND2_X1 U12298 ( .A1(n12250), .A2(n12274), .ZN(n12273) );
  OR2_X1 U12299 ( .A1(n12249), .A2(n12247), .ZN(n12274) );
  NOR2_X1 U12300 ( .A1(n11945), .A2(n7469), .ZN(n12250) );
  NAND2_X1 U12301 ( .A1(n12247), .A2(n12249), .ZN(n12272) );
  NAND2_X1 U12302 ( .A1(n12245), .A2(n12275), .ZN(n12249) );
  NAND2_X1 U12303 ( .A1(n12244), .A2(n12246), .ZN(n12275) );
  NAND2_X1 U12304 ( .A1(n12276), .A2(n12277), .ZN(n12246) );
  NAND2_X1 U12305 ( .A1(b_12_), .A2(a_3_), .ZN(n12277) );
  INV_X1 U12306 ( .A(n12278), .ZN(n12276) );
  XNOR2_X1 U12307 ( .A(n12279), .B(n12280), .ZN(n12244) );
  XOR2_X1 U12308 ( .A(n12281), .B(n12282), .Z(n12280) );
  NAND2_X1 U12309 ( .A1(a_4_), .A2(b_11_), .ZN(n12282) );
  NAND2_X1 U12310 ( .A1(a_3_), .A2(n12278), .ZN(n12245) );
  NAND2_X1 U12311 ( .A1(n12241), .A2(n12283), .ZN(n12278) );
  NAND2_X1 U12312 ( .A1(n12240), .A2(n12242), .ZN(n12283) );
  NAND2_X1 U12313 ( .A1(n12284), .A2(n12285), .ZN(n12242) );
  NAND2_X1 U12314 ( .A1(b_12_), .A2(a_4_), .ZN(n12285) );
  INV_X1 U12315 ( .A(n12286), .ZN(n12284) );
  XNOR2_X1 U12316 ( .A(n12287), .B(n12288), .ZN(n12240) );
  XOR2_X1 U12317 ( .A(n12289), .B(n12290), .Z(n12288) );
  NAND2_X1 U12318 ( .A1(a_5_), .A2(b_11_), .ZN(n12290) );
  NAND2_X1 U12319 ( .A1(a_4_), .A2(n12286), .ZN(n12241) );
  NAND2_X1 U12320 ( .A1(n12237), .A2(n12291), .ZN(n12286) );
  NAND2_X1 U12321 ( .A1(n12236), .A2(n12238), .ZN(n12291) );
  NAND2_X1 U12322 ( .A1(n12292), .A2(n12293), .ZN(n12238) );
  NAND2_X1 U12323 ( .A1(b_12_), .A2(a_5_), .ZN(n12293) );
  INV_X1 U12324 ( .A(n12294), .ZN(n12292) );
  XNOR2_X1 U12325 ( .A(n12295), .B(n12296), .ZN(n12236) );
  XOR2_X1 U12326 ( .A(n12297), .B(n12298), .Z(n12296) );
  NAND2_X1 U12327 ( .A1(a_6_), .A2(b_11_), .ZN(n12298) );
  NAND2_X1 U12328 ( .A1(a_5_), .A2(n12294), .ZN(n12237) );
  NAND2_X1 U12329 ( .A1(n12233), .A2(n12299), .ZN(n12294) );
  NAND2_X1 U12330 ( .A1(n12232), .A2(n12234), .ZN(n12299) );
  NAND2_X1 U12331 ( .A1(n12300), .A2(n12301), .ZN(n12234) );
  NAND2_X1 U12332 ( .A1(b_12_), .A2(a_6_), .ZN(n12301) );
  XNOR2_X1 U12333 ( .A(n12302), .B(n12303), .ZN(n12232) );
  XOR2_X1 U12334 ( .A(n12304), .B(n12305), .Z(n12303) );
  NAND2_X1 U12335 ( .A1(a_7_), .A2(b_11_), .ZN(n12305) );
  OR2_X1 U12336 ( .A1(n7450), .A2(n12300), .ZN(n12233) );
  NOR2_X1 U12337 ( .A1(n12228), .A2(n12306), .ZN(n12300) );
  AND2_X1 U12338 ( .A1(n12225), .A2(n12307), .ZN(n12306) );
  NAND2_X1 U12339 ( .A1(n12308), .A2(n12309), .ZN(n12307) );
  NAND2_X1 U12340 ( .A1(b_12_), .A2(a_7_), .ZN(n12309) );
  XOR2_X1 U12341 ( .A(n12310), .B(n12311), .Z(n12225) );
  XOR2_X1 U12342 ( .A(n12312), .B(n12313), .Z(n12310) );
  NOR2_X1 U12343 ( .A1(n12145), .A2(n7699), .ZN(n12313) );
  NOR2_X1 U12344 ( .A1(n7445), .A2(n12308), .ZN(n12228) );
  INV_X1 U12345 ( .A(n12230), .ZN(n12308) );
  NAND2_X1 U12346 ( .A1(n12223), .A2(n12314), .ZN(n12230) );
  NAND2_X1 U12347 ( .A1(n12222), .A2(n12224), .ZN(n12314) );
  NAND2_X1 U12348 ( .A1(n12315), .A2(n12316), .ZN(n12224) );
  NAND2_X1 U12349 ( .A1(b_12_), .A2(a_8_), .ZN(n12316) );
  INV_X1 U12350 ( .A(n12317), .ZN(n12315) );
  XOR2_X1 U12351 ( .A(n12318), .B(n12319), .Z(n12222) );
  XOR2_X1 U12352 ( .A(n12320), .B(n12321), .Z(n12318) );
  NOR2_X1 U12353 ( .A1(n12145), .A2(n7704), .ZN(n12321) );
  NAND2_X1 U12354 ( .A1(a_8_), .A2(n12317), .ZN(n12223) );
  NAND2_X1 U12355 ( .A1(n12322), .A2(n12323), .ZN(n12317) );
  NAND2_X1 U12356 ( .A1(n12324), .A2(b_12_), .ZN(n12323) );
  NOR2_X1 U12357 ( .A1(n12325), .A2(n7704), .ZN(n12324) );
  NOR2_X1 U12358 ( .A1(n12217), .A2(n12219), .ZN(n12325) );
  NAND2_X1 U12359 ( .A1(n12217), .A2(n12219), .ZN(n12322) );
  NAND2_X1 U12360 ( .A1(n12326), .A2(n12327), .ZN(n12219) );
  NAND2_X1 U12361 ( .A1(n12216), .A2(n12328), .ZN(n12327) );
  NAND2_X1 U12362 ( .A1(n12215), .A2(n12214), .ZN(n12328) );
  NOR2_X1 U12363 ( .A1(n11945), .A2(n7709), .ZN(n12216) );
  OR2_X1 U12364 ( .A1(n12214), .A2(n12215), .ZN(n12326) );
  AND2_X1 U12365 ( .A1(n12211), .A2(n12329), .ZN(n12215) );
  NAND2_X1 U12366 ( .A1(n12210), .A2(n12212), .ZN(n12329) );
  NAND2_X1 U12367 ( .A1(n12330), .A2(n12331), .ZN(n12212) );
  NAND2_X1 U12368 ( .A1(b_12_), .A2(a_11_), .ZN(n12331) );
  INV_X1 U12369 ( .A(n12332), .ZN(n12330) );
  XOR2_X1 U12370 ( .A(n12333), .B(n12334), .Z(n12210) );
  XOR2_X1 U12371 ( .A(n12335), .B(n12336), .Z(n12333) );
  NOR2_X1 U12372 ( .A1(n12145), .A2(n7718), .ZN(n12336) );
  NAND2_X1 U12373 ( .A1(a_11_), .A2(n12332), .ZN(n12211) );
  NAND2_X1 U12374 ( .A1(n12337), .A2(n12338), .ZN(n12332) );
  NAND2_X1 U12375 ( .A1(n12208), .A2(n12339), .ZN(n12338) );
  OR2_X1 U12376 ( .A1(n12207), .A2(n12206), .ZN(n12339) );
  INV_X1 U12377 ( .A(n12340), .ZN(n12208) );
  NAND2_X1 U12378 ( .A1(n12206), .A2(n12207), .ZN(n12337) );
  NAND2_X1 U12379 ( .A1(n12203), .A2(n12341), .ZN(n12207) );
  NAND2_X1 U12380 ( .A1(n12202), .A2(n12204), .ZN(n12341) );
  NAND2_X1 U12381 ( .A1(n12342), .A2(n12343), .ZN(n12204) );
  NAND2_X1 U12382 ( .A1(b_12_), .A2(a_13_), .ZN(n12343) );
  INV_X1 U12383 ( .A(n12344), .ZN(n12342) );
  XOR2_X1 U12384 ( .A(n12345), .B(n12346), .Z(n12202) );
  XOR2_X1 U12385 ( .A(n12347), .B(n12348), .Z(n12345) );
  NOR2_X1 U12386 ( .A1(n12145), .A2(n7727), .ZN(n12348) );
  NAND2_X1 U12387 ( .A1(a_13_), .A2(n12344), .ZN(n12203) );
  NAND2_X1 U12388 ( .A1(n12073), .A2(n12349), .ZN(n12344) );
  NAND2_X1 U12389 ( .A1(n12072), .A2(n12074), .ZN(n12349) );
  NAND2_X1 U12390 ( .A1(n12350), .A2(n12351), .ZN(n12074) );
  NAND2_X1 U12391 ( .A1(b_12_), .A2(a_14_), .ZN(n12351) );
  INV_X1 U12392 ( .A(n12352), .ZN(n12350) );
  XOR2_X1 U12393 ( .A(n12353), .B(n12354), .Z(n12072) );
  XOR2_X1 U12394 ( .A(n12355), .B(n12356), .Z(n12353) );
  NOR2_X1 U12395 ( .A1(n12145), .A2(n7406), .ZN(n12356) );
  NAND2_X1 U12396 ( .A1(a_14_), .A2(n12352), .ZN(n12073) );
  NAND2_X1 U12397 ( .A1(n12357), .A2(n12358), .ZN(n12352) );
  NAND2_X1 U12398 ( .A1(n12359), .A2(b_12_), .ZN(n12358) );
  NOR2_X1 U12399 ( .A1(n12360), .A2(n7406), .ZN(n12359) );
  NOR2_X1 U12400 ( .A1(n12197), .A2(n12199), .ZN(n12360) );
  NAND2_X1 U12401 ( .A1(n12197), .A2(n12199), .ZN(n12357) );
  NAND2_X1 U12402 ( .A1(n12361), .A2(n12362), .ZN(n12199) );
  NAND2_X1 U12403 ( .A1(n12196), .A2(n12363), .ZN(n12362) );
  NAND2_X1 U12404 ( .A1(n12195), .A2(n12194), .ZN(n12363) );
  NOR2_X1 U12405 ( .A1(n11945), .A2(n7736), .ZN(n12196) );
  OR2_X1 U12406 ( .A1(n12194), .A2(n12195), .ZN(n12361) );
  AND2_X1 U12407 ( .A1(n12364), .A2(n12365), .ZN(n12195) );
  NAND2_X1 U12408 ( .A1(n12192), .A2(n12366), .ZN(n12365) );
  OR2_X1 U12409 ( .A1(n12191), .A2(n12190), .ZN(n12366) );
  NOR2_X1 U12410 ( .A1(n11945), .A2(n7397), .ZN(n12192) );
  NAND2_X1 U12411 ( .A1(n12190), .A2(n12191), .ZN(n12364) );
  NAND2_X1 U12412 ( .A1(n12367), .A2(n12368), .ZN(n12191) );
  NAND2_X1 U12413 ( .A1(n12188), .A2(n12369), .ZN(n12368) );
  NAND2_X1 U12414 ( .A1(n12187), .A2(n12186), .ZN(n12369) );
  NOR2_X1 U12415 ( .A1(n11945), .A2(n7745), .ZN(n12188) );
  OR2_X1 U12416 ( .A1(n12186), .A2(n12187), .ZN(n12367) );
  AND2_X1 U12417 ( .A1(n12370), .A2(n12371), .ZN(n12187) );
  NAND2_X1 U12418 ( .A1(n12372), .A2(b_12_), .ZN(n12371) );
  NOR2_X1 U12419 ( .A1(n12373), .A2(n7750), .ZN(n12372) );
  NOR2_X1 U12420 ( .A1(n12182), .A2(n12183), .ZN(n12373) );
  NAND2_X1 U12421 ( .A1(n12182), .A2(n12183), .ZN(n12370) );
  NAND2_X1 U12422 ( .A1(n12374), .A2(n12375), .ZN(n12183) );
  NAND2_X1 U12423 ( .A1(n12376), .A2(b_12_), .ZN(n12375) );
  NOR2_X1 U12424 ( .A1(n12377), .A2(n7755), .ZN(n12376) );
  NOR2_X1 U12425 ( .A1(n12178), .A2(n12179), .ZN(n12377) );
  NAND2_X1 U12426 ( .A1(n12178), .A2(n12179), .ZN(n12374) );
  NAND2_X1 U12427 ( .A1(n12378), .A2(n12379), .ZN(n12179) );
  NAND2_X1 U12428 ( .A1(n12176), .A2(n12380), .ZN(n12379) );
  OR2_X1 U12429 ( .A1(n12175), .A2(n12173), .ZN(n12380) );
  NOR2_X1 U12430 ( .A1(n11945), .A2(n7760), .ZN(n12176) );
  NAND2_X1 U12431 ( .A1(n12173), .A2(n12175), .ZN(n12378) );
  NAND2_X1 U12432 ( .A1(n12381), .A2(n12382), .ZN(n12175) );
  NAND2_X1 U12433 ( .A1(n12383), .A2(b_12_), .ZN(n12382) );
  NOR2_X1 U12434 ( .A1(n12384), .A2(n7765), .ZN(n12383) );
  NOR2_X1 U12435 ( .A1(n12169), .A2(n12171), .ZN(n12384) );
  NAND2_X1 U12436 ( .A1(n12169), .A2(n12171), .ZN(n12381) );
  NAND2_X1 U12437 ( .A1(n12385), .A2(n12386), .ZN(n12171) );
  NAND2_X1 U12438 ( .A1(n12168), .A2(n12387), .ZN(n12386) );
  OR2_X1 U12439 ( .A1(n12167), .A2(n12166), .ZN(n12387) );
  NOR2_X1 U12440 ( .A1(n11945), .A2(n8014), .ZN(n12168) );
  NAND2_X1 U12441 ( .A1(n12166), .A2(n12167), .ZN(n12385) );
  NAND2_X1 U12442 ( .A1(n12388), .A2(n12389), .ZN(n12167) );
  NAND2_X1 U12443 ( .A1(n12390), .A2(b_12_), .ZN(n12389) );
  NOR2_X1 U12444 ( .A1(n12391), .A2(n7774), .ZN(n12390) );
  NOR2_X1 U12445 ( .A1(n12162), .A2(n12164), .ZN(n12391) );
  NAND2_X1 U12446 ( .A1(n12162), .A2(n12164), .ZN(n12388) );
  NAND2_X1 U12447 ( .A1(n12392), .A2(n12393), .ZN(n12164) );
  NAND2_X1 U12448 ( .A1(n12160), .A2(n12394), .ZN(n12393) );
  OR2_X1 U12449 ( .A1(n12159), .A2(n12158), .ZN(n12394) );
  NOR2_X1 U12450 ( .A1(n11945), .A2(n8022), .ZN(n12160) );
  NAND2_X1 U12451 ( .A1(n12158), .A2(n12159), .ZN(n12392) );
  NAND2_X1 U12452 ( .A1(n12155), .A2(n12395), .ZN(n12159) );
  NAND2_X1 U12453 ( .A1(n12154), .A2(n12156), .ZN(n12395) );
  NAND2_X1 U12454 ( .A1(n12396), .A2(n12397), .ZN(n12156) );
  NAND2_X1 U12455 ( .A1(b_12_), .A2(a_26_), .ZN(n12397) );
  INV_X1 U12456 ( .A(n12398), .ZN(n12396) );
  XNOR2_X1 U12457 ( .A(n12399), .B(n12400), .ZN(n12154) );
  NAND2_X1 U12458 ( .A1(n12401), .A2(n12402), .ZN(n12399) );
  NAND2_X1 U12459 ( .A1(a_26_), .A2(n12398), .ZN(n12155) );
  NAND2_X1 U12460 ( .A1(n12124), .A2(n12403), .ZN(n12398) );
  NAND2_X1 U12461 ( .A1(n12123), .A2(n12125), .ZN(n12403) );
  NAND2_X1 U12462 ( .A1(n12404), .A2(n12405), .ZN(n12125) );
  NAND2_X1 U12463 ( .A1(b_12_), .A2(a_27_), .ZN(n12405) );
  INV_X1 U12464 ( .A(n12406), .ZN(n12404) );
  XNOR2_X1 U12465 ( .A(n12407), .B(n12408), .ZN(n12123) );
  XOR2_X1 U12466 ( .A(n12409), .B(n12410), .Z(n12408) );
  NAND2_X1 U12467 ( .A1(a_28_), .A2(b_11_), .ZN(n12410) );
  NAND2_X1 U12468 ( .A1(a_27_), .A2(n12406), .ZN(n12124) );
  NAND2_X1 U12469 ( .A1(n12411), .A2(n12412), .ZN(n12406) );
  NAND2_X1 U12470 ( .A1(n12413), .A2(b_12_), .ZN(n12412) );
  NOR2_X1 U12471 ( .A1(n12414), .A2(n7803), .ZN(n12413) );
  NOR2_X1 U12472 ( .A1(n12130), .A2(n12132), .ZN(n12414) );
  NAND2_X1 U12473 ( .A1(n12130), .A2(n12132), .ZN(n12411) );
  NAND2_X1 U12474 ( .A1(n12415), .A2(n12416), .ZN(n12132) );
  NAND2_X1 U12475 ( .A1(n12150), .A2(n12417), .ZN(n12416) );
  NAND2_X1 U12476 ( .A1(n12152), .A2(n12151), .ZN(n12417) );
  NOR2_X1 U12477 ( .A1(n11945), .A2(n7337), .ZN(n12150) );
  OR2_X1 U12478 ( .A1(n12151), .A2(n12152), .ZN(n12415) );
  AND2_X1 U12479 ( .A1(n12418), .A2(n12419), .ZN(n12152) );
  NAND2_X1 U12480 ( .A1(n12420), .A2(a_31_), .ZN(n12419) );
  NOR2_X1 U12481 ( .A1(n12421), .A2(n12422), .ZN(n12420) );
  NOR2_X1 U12482 ( .A1(n7816), .A2(n12145), .ZN(n12421) );
  NAND2_X1 U12483 ( .A1(n12423), .A2(a_30_), .ZN(n12418) );
  NOR2_X1 U12484 ( .A1(n12424), .A2(n12145), .ZN(n12423) );
  NOR2_X1 U12485 ( .A1(n7810), .A2(n12422), .ZN(n12424) );
  NAND2_X1 U12486 ( .A1(n12425), .A2(b_12_), .ZN(n12151) );
  NOR2_X1 U12487 ( .A1(n12145), .A2(n8055), .ZN(n12425) );
  XOR2_X1 U12488 ( .A(n12426), .B(n12427), .Z(n12130) );
  XOR2_X1 U12489 ( .A(n12428), .B(n12429), .Z(n12426) );
  XNOR2_X1 U12490 ( .A(n12430), .B(n12431), .ZN(n12158) );
  NAND2_X1 U12491 ( .A1(n12432), .A2(n12433), .ZN(n12430) );
  XOR2_X1 U12492 ( .A(n12434), .B(n12435), .Z(n12162) );
  XOR2_X1 U12493 ( .A(n12436), .B(n12437), .Z(n12434) );
  XOR2_X1 U12494 ( .A(n12438), .B(n12439), .Z(n12166) );
  XNOR2_X1 U12495 ( .A(n12440), .B(n12441), .ZN(n12438) );
  NAND2_X1 U12496 ( .A1(a_24_), .A2(b_11_), .ZN(n12440) );
  XOR2_X1 U12497 ( .A(n12442), .B(n12443), .Z(n12169) );
  XOR2_X1 U12498 ( .A(n12444), .B(n12445), .Z(n12442) );
  XNOR2_X1 U12499 ( .A(n12446), .B(n12447), .ZN(n12173) );
  XOR2_X1 U12500 ( .A(n12448), .B(n12449), .Z(n12447) );
  NAND2_X1 U12501 ( .A1(a_22_), .A2(b_11_), .ZN(n12449) );
  XNOR2_X1 U12502 ( .A(n12450), .B(n12451), .ZN(n12178) );
  XNOR2_X1 U12503 ( .A(n12452), .B(n12453), .ZN(n12451) );
  XOR2_X1 U12504 ( .A(n12454), .B(n12455), .Z(n12182) );
  XOR2_X1 U12505 ( .A(n12456), .B(n12457), .Z(n12454) );
  XOR2_X1 U12506 ( .A(n12458), .B(n12459), .Z(n12186) );
  XOR2_X1 U12507 ( .A(n12460), .B(n12461), .Z(n12459) );
  NAND2_X1 U12508 ( .A1(a_19_), .A2(b_11_), .ZN(n12461) );
  XNOR2_X1 U12509 ( .A(n12462), .B(n12463), .ZN(n12190) );
  NAND2_X1 U12510 ( .A1(n12464), .A2(n12465), .ZN(n12462) );
  XNOR2_X1 U12511 ( .A(n12466), .B(n12467), .ZN(n12194) );
  XOR2_X1 U12512 ( .A(n12468), .B(n12469), .Z(n12466) );
  NOR2_X1 U12513 ( .A1(n12145), .A2(n7397), .ZN(n12469) );
  XOR2_X1 U12514 ( .A(n12470), .B(n12471), .Z(n12197) );
  XOR2_X1 U12515 ( .A(n12472), .B(n12473), .Z(n12470) );
  NOR2_X1 U12516 ( .A1(n12145), .A2(n7736), .ZN(n12473) );
  XOR2_X1 U12517 ( .A(n12474), .B(n12475), .Z(n12206) );
  XOR2_X1 U12518 ( .A(n12476), .B(n12477), .Z(n12474) );
  NOR2_X1 U12519 ( .A1(n12145), .A2(n7415), .ZN(n12477) );
  XNOR2_X1 U12520 ( .A(n12478), .B(n12479), .ZN(n12214) );
  XOR2_X1 U12521 ( .A(n12480), .B(n12481), .Z(n12478) );
  XOR2_X1 U12522 ( .A(n12482), .B(n12483), .Z(n12217) );
  XNOR2_X1 U12523 ( .A(n12484), .B(n12485), .ZN(n12482) );
  NAND2_X1 U12524 ( .A1(a_10_), .A2(b_11_), .ZN(n12484) );
  XNOR2_X1 U12525 ( .A(n12486), .B(n12487), .ZN(n12247) );
  XOR2_X1 U12526 ( .A(n12488), .B(n12489), .Z(n12487) );
  NAND2_X1 U12527 ( .A1(a_3_), .A2(b_11_), .ZN(n12489) );
  XOR2_X1 U12528 ( .A(n12490), .B(n12491), .Z(n12251) );
  XOR2_X1 U12529 ( .A(n12492), .B(n12493), .Z(n12490) );
  NOR2_X1 U12530 ( .A1(n12145), .A2(n7469), .ZN(n12493) );
  XOR2_X1 U12531 ( .A(n12494), .B(n12495), .Z(n11775) );
  XOR2_X1 U12532 ( .A(n12496), .B(n12497), .Z(n12494) );
  NOR2_X1 U12533 ( .A1(n12145), .A2(n7669), .ZN(n12497) );
  XOR2_X1 U12534 ( .A(n12498), .B(n12499), .Z(n7593) );
  XOR2_X1 U12535 ( .A(n12500), .B(n12501), .Z(n12498) );
  OR2_X1 U12536 ( .A1(n7585), .A2(n7584), .ZN(n7572) );
  XNOR2_X1 U12537 ( .A(n12502), .B(n12503), .ZN(n7584) );
  NAND2_X1 U12538 ( .A1(n12504), .A2(n12262), .ZN(n7585) );
  NAND2_X1 U12539 ( .A1(n12505), .A2(n12506), .ZN(n12262) );
  NAND2_X1 U12540 ( .A1(n12501), .A2(n12507), .ZN(n12506) );
  OR2_X1 U12541 ( .A1(n12500), .A2(n12499), .ZN(n12507) );
  NOR2_X1 U12542 ( .A1(n12145), .A2(n7478), .ZN(n12501) );
  NAND2_X1 U12543 ( .A1(n12499), .A2(n12500), .ZN(n12505) );
  NAND2_X1 U12544 ( .A1(n12508), .A2(n12509), .ZN(n12500) );
  NAND2_X1 U12545 ( .A1(n12510), .A2(a_1_), .ZN(n12509) );
  NOR2_X1 U12546 ( .A1(n12511), .A2(n12145), .ZN(n12510) );
  NOR2_X1 U12547 ( .A1(n12495), .A2(n12496), .ZN(n12511) );
  NAND2_X1 U12548 ( .A1(n12495), .A2(n12496), .ZN(n12508) );
  NAND2_X1 U12549 ( .A1(n12512), .A2(n12513), .ZN(n12496) );
  NAND2_X1 U12550 ( .A1(n12514), .A2(a_2_), .ZN(n12513) );
  NOR2_X1 U12551 ( .A1(n12515), .A2(n12145), .ZN(n12514) );
  NOR2_X1 U12552 ( .A1(n12491), .A2(n12492), .ZN(n12515) );
  NAND2_X1 U12553 ( .A1(n12491), .A2(n12492), .ZN(n12512) );
  NAND2_X1 U12554 ( .A1(n12516), .A2(n12517), .ZN(n12492) );
  NAND2_X1 U12555 ( .A1(n12518), .A2(a_3_), .ZN(n12517) );
  NOR2_X1 U12556 ( .A1(n12519), .A2(n12145), .ZN(n12518) );
  NOR2_X1 U12557 ( .A1(n12486), .A2(n12488), .ZN(n12519) );
  NAND2_X1 U12558 ( .A1(n12486), .A2(n12488), .ZN(n12516) );
  NAND2_X1 U12559 ( .A1(n12520), .A2(n12521), .ZN(n12488) );
  NAND2_X1 U12560 ( .A1(n12522), .A2(a_4_), .ZN(n12521) );
  NOR2_X1 U12561 ( .A1(n12523), .A2(n12145), .ZN(n12522) );
  NOR2_X1 U12562 ( .A1(n12279), .A2(n12281), .ZN(n12523) );
  NAND2_X1 U12563 ( .A1(n12279), .A2(n12281), .ZN(n12520) );
  NAND2_X1 U12564 ( .A1(n12524), .A2(n12525), .ZN(n12281) );
  NAND2_X1 U12565 ( .A1(n12526), .A2(a_5_), .ZN(n12525) );
  NOR2_X1 U12566 ( .A1(n12527), .A2(n12145), .ZN(n12526) );
  NOR2_X1 U12567 ( .A1(n12287), .A2(n12289), .ZN(n12527) );
  NAND2_X1 U12568 ( .A1(n12287), .A2(n12289), .ZN(n12524) );
  NAND2_X1 U12569 ( .A1(n12528), .A2(n12529), .ZN(n12289) );
  NAND2_X1 U12570 ( .A1(n12530), .A2(a_6_), .ZN(n12529) );
  NOR2_X1 U12571 ( .A1(n12531), .A2(n12145), .ZN(n12530) );
  NOR2_X1 U12572 ( .A1(n12295), .A2(n12297), .ZN(n12531) );
  NAND2_X1 U12573 ( .A1(n12295), .A2(n12297), .ZN(n12528) );
  NAND2_X1 U12574 ( .A1(n12532), .A2(n12533), .ZN(n12297) );
  NAND2_X1 U12575 ( .A1(n12534), .A2(a_7_), .ZN(n12533) );
  NOR2_X1 U12576 ( .A1(n12535), .A2(n12145), .ZN(n12534) );
  NOR2_X1 U12577 ( .A1(n12302), .A2(n12304), .ZN(n12535) );
  NAND2_X1 U12578 ( .A1(n12302), .A2(n12304), .ZN(n12532) );
  NAND2_X1 U12579 ( .A1(n12536), .A2(n12537), .ZN(n12304) );
  NAND2_X1 U12580 ( .A1(n12538), .A2(a_8_), .ZN(n12537) );
  NOR2_X1 U12581 ( .A1(n12539), .A2(n12145), .ZN(n12538) );
  NOR2_X1 U12582 ( .A1(n12311), .A2(n12312), .ZN(n12539) );
  NAND2_X1 U12583 ( .A1(n12311), .A2(n12312), .ZN(n12536) );
  NAND2_X1 U12584 ( .A1(n12540), .A2(n12541), .ZN(n12312) );
  NAND2_X1 U12585 ( .A1(n12542), .A2(a_9_), .ZN(n12541) );
  NOR2_X1 U12586 ( .A1(n12543), .A2(n12145), .ZN(n12542) );
  NOR2_X1 U12587 ( .A1(n12319), .A2(n12320), .ZN(n12543) );
  NAND2_X1 U12588 ( .A1(n12319), .A2(n12320), .ZN(n12540) );
  NAND2_X1 U12589 ( .A1(n12544), .A2(n12545), .ZN(n12320) );
  NAND2_X1 U12590 ( .A1(n12546), .A2(a_10_), .ZN(n12545) );
  NOR2_X1 U12591 ( .A1(n12547), .A2(n12145), .ZN(n12546) );
  NOR2_X1 U12592 ( .A1(n12483), .A2(n12485), .ZN(n12547) );
  NAND2_X1 U12593 ( .A1(n12483), .A2(n12485), .ZN(n12544) );
  NAND2_X1 U12594 ( .A1(n12548), .A2(n12549), .ZN(n12485) );
  NAND2_X1 U12595 ( .A1(n12479), .A2(n12550), .ZN(n12549) );
  OR2_X1 U12596 ( .A1(n12480), .A2(n12481), .ZN(n12550) );
  XNOR2_X1 U12597 ( .A(n12551), .B(n12552), .ZN(n12479) );
  NAND2_X1 U12598 ( .A1(n12553), .A2(n12554), .ZN(n12551) );
  NAND2_X1 U12599 ( .A1(n12481), .A2(n12480), .ZN(n12548) );
  NAND2_X1 U12600 ( .A1(n12555), .A2(n12556), .ZN(n12480) );
  NAND2_X1 U12601 ( .A1(n12557), .A2(a_12_), .ZN(n12556) );
  NOR2_X1 U12602 ( .A1(n12558), .A2(n12145), .ZN(n12557) );
  NOR2_X1 U12603 ( .A1(n12334), .A2(n12335), .ZN(n12558) );
  NAND2_X1 U12604 ( .A1(n12334), .A2(n12335), .ZN(n12555) );
  NAND2_X1 U12605 ( .A1(n12559), .A2(n12560), .ZN(n12335) );
  NAND2_X1 U12606 ( .A1(n12561), .A2(a_13_), .ZN(n12560) );
  NOR2_X1 U12607 ( .A1(n12562), .A2(n12145), .ZN(n12561) );
  NOR2_X1 U12608 ( .A1(n12475), .A2(n12476), .ZN(n12562) );
  NAND2_X1 U12609 ( .A1(n12475), .A2(n12476), .ZN(n12559) );
  NAND2_X1 U12610 ( .A1(n12563), .A2(n12564), .ZN(n12476) );
  NAND2_X1 U12611 ( .A1(n12565), .A2(a_14_), .ZN(n12564) );
  NOR2_X1 U12612 ( .A1(n12566), .A2(n12145), .ZN(n12565) );
  NOR2_X1 U12613 ( .A1(n12346), .A2(n12347), .ZN(n12566) );
  NAND2_X1 U12614 ( .A1(n12346), .A2(n12347), .ZN(n12563) );
  NAND2_X1 U12615 ( .A1(n12567), .A2(n12568), .ZN(n12347) );
  NAND2_X1 U12616 ( .A1(n12569), .A2(a_15_), .ZN(n12568) );
  NOR2_X1 U12617 ( .A1(n12570), .A2(n12145), .ZN(n12569) );
  NOR2_X1 U12618 ( .A1(n12354), .A2(n12355), .ZN(n12570) );
  NAND2_X1 U12619 ( .A1(n12354), .A2(n12355), .ZN(n12567) );
  NAND2_X1 U12620 ( .A1(n12571), .A2(n12572), .ZN(n12355) );
  NAND2_X1 U12621 ( .A1(n12573), .A2(a_16_), .ZN(n12572) );
  NOR2_X1 U12622 ( .A1(n12574), .A2(n12145), .ZN(n12573) );
  NOR2_X1 U12623 ( .A1(n12471), .A2(n12472), .ZN(n12574) );
  NAND2_X1 U12624 ( .A1(n12471), .A2(n12472), .ZN(n12571) );
  NAND2_X1 U12625 ( .A1(n12575), .A2(n12576), .ZN(n12472) );
  NAND2_X1 U12626 ( .A1(n12577), .A2(a_17_), .ZN(n12576) );
  NOR2_X1 U12627 ( .A1(n12578), .A2(n12145), .ZN(n12577) );
  NOR2_X1 U12628 ( .A1(n12467), .A2(n12468), .ZN(n12578) );
  NAND2_X1 U12629 ( .A1(n12467), .A2(n12468), .ZN(n12575) );
  NAND2_X1 U12630 ( .A1(n12464), .A2(n12579), .ZN(n12468) );
  NAND2_X1 U12631 ( .A1(n12463), .A2(n12465), .ZN(n12579) );
  NAND2_X1 U12632 ( .A1(n12580), .A2(n12581), .ZN(n12465) );
  NAND2_X1 U12633 ( .A1(a_18_), .A2(b_11_), .ZN(n12581) );
  INV_X1 U12634 ( .A(n12582), .ZN(n12580) );
  XNOR2_X1 U12635 ( .A(n12583), .B(n12584), .ZN(n12463) );
  XNOR2_X1 U12636 ( .A(n12585), .B(n12586), .ZN(n12583) );
  NAND2_X1 U12637 ( .A1(a_18_), .A2(n12582), .ZN(n12464) );
  NAND2_X1 U12638 ( .A1(n12587), .A2(n12588), .ZN(n12582) );
  NAND2_X1 U12639 ( .A1(n12589), .A2(a_19_), .ZN(n12588) );
  NOR2_X1 U12640 ( .A1(n12590), .A2(n12145), .ZN(n12589) );
  NOR2_X1 U12641 ( .A1(n12458), .A2(n12460), .ZN(n12590) );
  NAND2_X1 U12642 ( .A1(n12458), .A2(n12460), .ZN(n12587) );
  NAND2_X1 U12643 ( .A1(n12591), .A2(n12592), .ZN(n12460) );
  NAND2_X1 U12644 ( .A1(n12457), .A2(n12593), .ZN(n12592) );
  OR2_X1 U12645 ( .A1(n12456), .A2(n12455), .ZN(n12593) );
  NOR2_X1 U12646 ( .A1(n7755), .A2(n12145), .ZN(n12457) );
  NAND2_X1 U12647 ( .A1(n12455), .A2(n12456), .ZN(n12591) );
  NAND2_X1 U12648 ( .A1(n12594), .A2(n12595), .ZN(n12456) );
  NAND2_X1 U12649 ( .A1(n12453), .A2(n12596), .ZN(n12595) );
  OR2_X1 U12650 ( .A1(n12452), .A2(n12450), .ZN(n12596) );
  NOR2_X1 U12651 ( .A1(n7760), .A2(n12145), .ZN(n12453) );
  NAND2_X1 U12652 ( .A1(n12450), .A2(n12452), .ZN(n12594) );
  NAND2_X1 U12653 ( .A1(n12597), .A2(n12598), .ZN(n12452) );
  NAND2_X1 U12654 ( .A1(n12599), .A2(a_22_), .ZN(n12598) );
  NOR2_X1 U12655 ( .A1(n12600), .A2(n12145), .ZN(n12599) );
  NOR2_X1 U12656 ( .A1(n12446), .A2(n12448), .ZN(n12600) );
  NAND2_X1 U12657 ( .A1(n12446), .A2(n12448), .ZN(n12597) );
  NAND2_X1 U12658 ( .A1(n12601), .A2(n12602), .ZN(n12448) );
  NAND2_X1 U12659 ( .A1(n12445), .A2(n12603), .ZN(n12602) );
  OR2_X1 U12660 ( .A1(n12444), .A2(n12443), .ZN(n12603) );
  NOR2_X1 U12661 ( .A1(n8014), .A2(n12145), .ZN(n12445) );
  NAND2_X1 U12662 ( .A1(n12443), .A2(n12444), .ZN(n12601) );
  NAND2_X1 U12663 ( .A1(n12604), .A2(n12605), .ZN(n12444) );
  NAND2_X1 U12664 ( .A1(n12606), .A2(a_24_), .ZN(n12605) );
  NOR2_X1 U12665 ( .A1(n12607), .A2(n12145), .ZN(n12606) );
  NOR2_X1 U12666 ( .A1(n12439), .A2(n12441), .ZN(n12607) );
  NAND2_X1 U12667 ( .A1(n12439), .A2(n12441), .ZN(n12604) );
  NAND2_X1 U12668 ( .A1(n12608), .A2(n12609), .ZN(n12441) );
  NAND2_X1 U12669 ( .A1(n12437), .A2(n12610), .ZN(n12609) );
  OR2_X1 U12670 ( .A1(n12436), .A2(n12435), .ZN(n12610) );
  NOR2_X1 U12671 ( .A1(n8022), .A2(n12145), .ZN(n12437) );
  NAND2_X1 U12672 ( .A1(n12435), .A2(n12436), .ZN(n12608) );
  NAND2_X1 U12673 ( .A1(n12432), .A2(n12611), .ZN(n12436) );
  NAND2_X1 U12674 ( .A1(n12431), .A2(n12433), .ZN(n12611) );
  NAND2_X1 U12675 ( .A1(n12612), .A2(n12613), .ZN(n12433) );
  NAND2_X1 U12676 ( .A1(a_26_), .A2(b_11_), .ZN(n12613) );
  INV_X1 U12677 ( .A(n12614), .ZN(n12612) );
  XNOR2_X1 U12678 ( .A(n12615), .B(n12616), .ZN(n12431) );
  NAND2_X1 U12679 ( .A1(n12617), .A2(n12618), .ZN(n12615) );
  NAND2_X1 U12680 ( .A1(a_26_), .A2(n12614), .ZN(n12432) );
  NAND2_X1 U12681 ( .A1(n12401), .A2(n12619), .ZN(n12614) );
  NAND2_X1 U12682 ( .A1(n12400), .A2(n12402), .ZN(n12619) );
  NAND2_X1 U12683 ( .A1(n12620), .A2(n12621), .ZN(n12402) );
  NAND2_X1 U12684 ( .A1(a_27_), .A2(b_11_), .ZN(n12621) );
  INV_X1 U12685 ( .A(n12622), .ZN(n12620) );
  XNOR2_X1 U12686 ( .A(n12623), .B(n12624), .ZN(n12400) );
  XOR2_X1 U12687 ( .A(n12625), .B(n12626), .Z(n12624) );
  NAND2_X1 U12688 ( .A1(a_28_), .A2(b_10_), .ZN(n12626) );
  NAND2_X1 U12689 ( .A1(a_27_), .A2(n12622), .ZN(n12401) );
  NAND2_X1 U12690 ( .A1(n12627), .A2(n12628), .ZN(n12622) );
  NAND2_X1 U12691 ( .A1(n12629), .A2(a_28_), .ZN(n12628) );
  NOR2_X1 U12692 ( .A1(n12630), .A2(n12145), .ZN(n12629) );
  NOR2_X1 U12693 ( .A1(n12407), .A2(n12409), .ZN(n12630) );
  NAND2_X1 U12694 ( .A1(n12407), .A2(n12409), .ZN(n12627) );
  NAND2_X1 U12695 ( .A1(n12631), .A2(n12632), .ZN(n12409) );
  NAND2_X1 U12696 ( .A1(n12427), .A2(n12633), .ZN(n12632) );
  NAND2_X1 U12697 ( .A1(n12429), .A2(n12428), .ZN(n12633) );
  NOR2_X1 U12698 ( .A1(n7337), .A2(n12145), .ZN(n12427) );
  OR2_X1 U12699 ( .A1(n12428), .A2(n12429), .ZN(n12631) );
  AND2_X1 U12700 ( .A1(n12634), .A2(n12635), .ZN(n12429) );
  NAND2_X1 U12701 ( .A1(n12636), .A2(b_10_), .ZN(n12635) );
  NOR2_X1 U12702 ( .A1(n12637), .A2(n8052), .ZN(n12636) );
  NOR2_X1 U12703 ( .A1(n7810), .A2(n12638), .ZN(n12637) );
  NAND2_X1 U12704 ( .A1(n12639), .A2(a_31_), .ZN(n12634) );
  NOR2_X1 U12705 ( .A1(n12640), .A2(n12638), .ZN(n12639) );
  NOR2_X1 U12706 ( .A1(n7816), .A2(n12422), .ZN(n12640) );
  NAND2_X1 U12707 ( .A1(n12641), .A2(n12642), .ZN(n12428) );
  NOR2_X1 U12708 ( .A1(n12145), .A2(n12422), .ZN(n12641) );
  XOR2_X1 U12709 ( .A(n12643), .B(n12644), .Z(n12407) );
  XOR2_X1 U12710 ( .A(n12645), .B(n12646), .Z(n12643) );
  XNOR2_X1 U12711 ( .A(n12647), .B(n12648), .ZN(n12435) );
  NAND2_X1 U12712 ( .A1(n12649), .A2(n12650), .ZN(n12647) );
  XOR2_X1 U12713 ( .A(n12651), .B(n12652), .Z(n12439) );
  XOR2_X1 U12714 ( .A(n12653), .B(n12654), .Z(n12651) );
  XOR2_X1 U12715 ( .A(n12655), .B(n12656), .Z(n12443) );
  XOR2_X1 U12716 ( .A(n12657), .B(n12658), .Z(n12655) );
  NOR2_X1 U12717 ( .A1(n12422), .A2(n7774), .ZN(n12658) );
  XOR2_X1 U12718 ( .A(n12659), .B(n12660), .Z(n12446) );
  XOR2_X1 U12719 ( .A(n12661), .B(n12662), .Z(n12659) );
  XOR2_X1 U12720 ( .A(n12663), .B(n12664), .Z(n12450) );
  XOR2_X1 U12721 ( .A(n12665), .B(n12666), .Z(n12663) );
  NOR2_X1 U12722 ( .A1(n12422), .A2(n7765), .ZN(n12666) );
  XOR2_X1 U12723 ( .A(n12667), .B(n12668), .Z(n12455) );
  XOR2_X1 U12724 ( .A(n12669), .B(n12670), .Z(n12667) );
  NOR2_X1 U12725 ( .A1(n7760), .A2(n12422), .ZN(n12670) );
  XNOR2_X1 U12726 ( .A(n12671), .B(n12672), .ZN(n12458) );
  XNOR2_X1 U12727 ( .A(n12673), .B(n12674), .ZN(n12671) );
  XNOR2_X1 U12728 ( .A(n12675), .B(n12676), .ZN(n12467) );
  XNOR2_X1 U12729 ( .A(n12677), .B(n12678), .ZN(n12675) );
  XNOR2_X1 U12730 ( .A(n12679), .B(n12680), .ZN(n12471) );
  XOR2_X1 U12731 ( .A(n12681), .B(n12682), .Z(n12680) );
  NAND2_X1 U12732 ( .A1(a_17_), .A2(b_10_), .ZN(n12682) );
  XNOR2_X1 U12733 ( .A(n12683), .B(n12684), .ZN(n12354) );
  NAND2_X1 U12734 ( .A1(n12685), .A2(n12686), .ZN(n12683) );
  XNOR2_X1 U12735 ( .A(n12687), .B(n12688), .ZN(n12346) );
  NAND2_X1 U12736 ( .A1(n12689), .A2(n12690), .ZN(n12687) );
  XNOR2_X1 U12737 ( .A(n12691), .B(n12692), .ZN(n12475) );
  NAND2_X1 U12738 ( .A1(n12693), .A2(n12694), .ZN(n12691) );
  XNOR2_X1 U12739 ( .A(n12695), .B(n12696), .ZN(n12334) );
  NAND2_X1 U12740 ( .A1(n12697), .A2(n12698), .ZN(n12695) );
  XNOR2_X1 U12741 ( .A(n12699), .B(n12700), .ZN(n12483) );
  NAND2_X1 U12742 ( .A1(n12701), .A2(n12702), .ZN(n12699) );
  XOR2_X1 U12743 ( .A(n12703), .B(n12704), .Z(n12319) );
  XOR2_X1 U12744 ( .A(n12705), .B(n12706), .Z(n12703) );
  XNOR2_X1 U12745 ( .A(n12707), .B(n12708), .ZN(n12311) );
  NAND2_X1 U12746 ( .A1(n12709), .A2(n12710), .ZN(n12707) );
  XNOR2_X1 U12747 ( .A(n12711), .B(n12712), .ZN(n12302) );
  NAND2_X1 U12748 ( .A1(n12713), .A2(n12714), .ZN(n12711) );
  XNOR2_X1 U12749 ( .A(n12715), .B(n12716), .ZN(n12295) );
  XNOR2_X1 U12750 ( .A(n12717), .B(n12718), .ZN(n12715) );
  XNOR2_X1 U12751 ( .A(n12719), .B(n12720), .ZN(n12287) );
  XNOR2_X1 U12752 ( .A(n12721), .B(n12722), .ZN(n12720) );
  XNOR2_X1 U12753 ( .A(n12723), .B(n12724), .ZN(n12279) );
  XNOR2_X1 U12754 ( .A(n12725), .B(n12726), .ZN(n12724) );
  XNOR2_X1 U12755 ( .A(n12727), .B(n12728), .ZN(n12486) );
  XNOR2_X1 U12756 ( .A(n12729), .B(n12730), .ZN(n12728) );
  XNOR2_X1 U12757 ( .A(n12731), .B(n12732), .ZN(n12491) );
  XNOR2_X1 U12758 ( .A(n12733), .B(n12734), .ZN(n12732) );
  XNOR2_X1 U12759 ( .A(n12735), .B(n12736), .ZN(n12495) );
  XNOR2_X1 U12760 ( .A(n12737), .B(n12738), .ZN(n12736) );
  XOR2_X1 U12761 ( .A(n12739), .B(n12740), .Z(n12499) );
  XNOR2_X1 U12762 ( .A(n12741), .B(n12742), .ZN(n12739) );
  NAND2_X1 U12763 ( .A1(a_1_), .A2(b_10_), .ZN(n12741) );
  XOR2_X1 U12764 ( .A(n12743), .B(n12264), .Z(n12504) );
  XNOR2_X1 U12765 ( .A(n12744), .B(n12745), .ZN(n12264) );
  NOR2_X1 U12766 ( .A1(n7478), .A2(n12422), .ZN(n12745) );
  INV_X1 U12767 ( .A(n12263), .ZN(n12743) );
  NAND2_X1 U12768 ( .A1(n12746), .A2(n12747), .ZN(n7312) );
  OR2_X1 U12769 ( .A1(n12747), .A2(n12746), .ZN(n7311) );
  NAND2_X1 U12770 ( .A1(n12748), .A2(n12749), .ZN(n12746) );
  NAND2_X1 U12771 ( .A1(n12750), .A2(n12751), .ZN(n12749) );
  INV_X1 U12772 ( .A(n12752), .ZN(n12751) );
  XOR2_X1 U12773 ( .A(n12753), .B(n12754), .Z(n12750) );
  NAND2_X1 U12774 ( .A1(n12503), .A2(n12502), .ZN(n12747) );
  NAND2_X1 U12775 ( .A1(n12755), .A2(n12756), .ZN(n12502) );
  NAND2_X1 U12776 ( .A1(n12757), .A2(b_10_), .ZN(n12756) );
  NOR2_X1 U12777 ( .A1(n12758), .A2(n7478), .ZN(n12757) );
  NOR2_X1 U12778 ( .A1(n12263), .A2(n12744), .ZN(n12758) );
  NAND2_X1 U12779 ( .A1(n12263), .A2(n12744), .ZN(n12755) );
  NAND2_X1 U12780 ( .A1(n12759), .A2(n12760), .ZN(n12744) );
  NAND2_X1 U12781 ( .A1(n12761), .A2(a_1_), .ZN(n12760) );
  NOR2_X1 U12782 ( .A1(n12762), .A2(n12422), .ZN(n12761) );
  NOR2_X1 U12783 ( .A1(n12740), .A2(n12742), .ZN(n12762) );
  NAND2_X1 U12784 ( .A1(n12740), .A2(n12742), .ZN(n12759) );
  NAND2_X1 U12785 ( .A1(n12763), .A2(n12764), .ZN(n12742) );
  NAND2_X1 U12786 ( .A1(n12738), .A2(n12765), .ZN(n12764) );
  OR2_X1 U12787 ( .A1(n12737), .A2(n12735), .ZN(n12765) );
  NOR2_X1 U12788 ( .A1(n7469), .A2(n12422), .ZN(n12738) );
  NAND2_X1 U12789 ( .A1(n12735), .A2(n12737), .ZN(n12763) );
  NAND2_X1 U12790 ( .A1(n12766), .A2(n12767), .ZN(n12737) );
  NAND2_X1 U12791 ( .A1(n12734), .A2(n12768), .ZN(n12767) );
  OR2_X1 U12792 ( .A1(n12733), .A2(n12731), .ZN(n12768) );
  NOR2_X1 U12793 ( .A1(n7464), .A2(n12422), .ZN(n12734) );
  NAND2_X1 U12794 ( .A1(n12731), .A2(n12733), .ZN(n12766) );
  NAND2_X1 U12795 ( .A1(n12769), .A2(n12770), .ZN(n12733) );
  NAND2_X1 U12796 ( .A1(n12730), .A2(n12771), .ZN(n12770) );
  OR2_X1 U12797 ( .A1(n12729), .A2(n12727), .ZN(n12771) );
  NOR2_X1 U12798 ( .A1(n7682), .A2(n12422), .ZN(n12730) );
  NAND2_X1 U12799 ( .A1(n12727), .A2(n12729), .ZN(n12769) );
  NAND2_X1 U12800 ( .A1(n12772), .A2(n12773), .ZN(n12729) );
  NAND2_X1 U12801 ( .A1(n12726), .A2(n12774), .ZN(n12773) );
  OR2_X1 U12802 ( .A1(n12723), .A2(n12725), .ZN(n12774) );
  NOR2_X1 U12803 ( .A1(n7455), .A2(n12422), .ZN(n12726) );
  NAND2_X1 U12804 ( .A1(n12723), .A2(n12725), .ZN(n12772) );
  NAND2_X1 U12805 ( .A1(n12775), .A2(n12776), .ZN(n12725) );
  NAND2_X1 U12806 ( .A1(n12722), .A2(n12777), .ZN(n12776) );
  OR2_X1 U12807 ( .A1(n12721), .A2(n12719), .ZN(n12777) );
  NOR2_X1 U12808 ( .A1(n7450), .A2(n12422), .ZN(n12722) );
  NAND2_X1 U12809 ( .A1(n12719), .A2(n12721), .ZN(n12775) );
  NAND2_X1 U12810 ( .A1(n12778), .A2(n12779), .ZN(n12721) );
  NAND2_X1 U12811 ( .A1(n12718), .A2(n12780), .ZN(n12779) );
  NAND2_X1 U12812 ( .A1(n12717), .A2(n12716), .ZN(n12780) );
  NOR2_X1 U12813 ( .A1(n7445), .A2(n12422), .ZN(n12718) );
  OR2_X1 U12814 ( .A1(n12716), .A2(n12717), .ZN(n12778) );
  AND2_X1 U12815 ( .A1(n12713), .A2(n12781), .ZN(n12717) );
  NAND2_X1 U12816 ( .A1(n12712), .A2(n12714), .ZN(n12781) );
  NAND2_X1 U12817 ( .A1(n12782), .A2(n12783), .ZN(n12714) );
  NAND2_X1 U12818 ( .A1(a_8_), .A2(b_10_), .ZN(n12783) );
  INV_X1 U12819 ( .A(n12784), .ZN(n12782) );
  XOR2_X1 U12820 ( .A(n12785), .B(n12786), .Z(n12712) );
  XOR2_X1 U12821 ( .A(n12787), .B(n12788), .Z(n12785) );
  NAND2_X1 U12822 ( .A1(a_8_), .A2(n12784), .ZN(n12713) );
  NAND2_X1 U12823 ( .A1(n12709), .A2(n12789), .ZN(n12784) );
  NAND2_X1 U12824 ( .A1(n12708), .A2(n12710), .ZN(n12789) );
  NAND2_X1 U12825 ( .A1(n12790), .A2(n12791), .ZN(n12710) );
  NAND2_X1 U12826 ( .A1(a_9_), .A2(b_10_), .ZN(n12791) );
  INV_X1 U12827 ( .A(n12792), .ZN(n12790) );
  XOR2_X1 U12828 ( .A(n12793), .B(n12794), .Z(n12708) );
  XOR2_X1 U12829 ( .A(n12795), .B(n12796), .Z(n12793) );
  NOR2_X1 U12830 ( .A1(n12638), .A2(n7709), .ZN(n12796) );
  NAND2_X1 U12831 ( .A1(a_9_), .A2(n12792), .ZN(n12709) );
  NAND2_X1 U12832 ( .A1(n12797), .A2(n12798), .ZN(n12792) );
  NAND2_X1 U12833 ( .A1(n12706), .A2(n12799), .ZN(n12798) );
  OR2_X1 U12834 ( .A1(n12704), .A2(n12705), .ZN(n12799) );
  INV_X1 U12835 ( .A(n12800), .ZN(n12706) );
  NAND2_X1 U12836 ( .A1(n12704), .A2(n12705), .ZN(n12797) );
  NAND2_X1 U12837 ( .A1(n12701), .A2(n12801), .ZN(n12705) );
  NAND2_X1 U12838 ( .A1(n12700), .A2(n12702), .ZN(n12801) );
  NAND2_X1 U12839 ( .A1(n12802), .A2(n12803), .ZN(n12702) );
  NAND2_X1 U12840 ( .A1(b_10_), .A2(a_11_), .ZN(n12803) );
  INV_X1 U12841 ( .A(n12804), .ZN(n12802) );
  XNOR2_X1 U12842 ( .A(n12805), .B(n12806), .ZN(n12700) );
  XOR2_X1 U12843 ( .A(n12807), .B(n12808), .Z(n12806) );
  NAND2_X1 U12844 ( .A1(a_12_), .A2(b_9_), .ZN(n12808) );
  NAND2_X1 U12845 ( .A1(a_11_), .A2(n12804), .ZN(n12701) );
  NAND2_X1 U12846 ( .A1(n12553), .A2(n12809), .ZN(n12804) );
  NAND2_X1 U12847 ( .A1(n12552), .A2(n12554), .ZN(n12809) );
  NAND2_X1 U12848 ( .A1(n12810), .A2(n12811), .ZN(n12554) );
  NAND2_X1 U12849 ( .A1(a_12_), .A2(b_10_), .ZN(n12811) );
  INV_X1 U12850 ( .A(n12812), .ZN(n12810) );
  XOR2_X1 U12851 ( .A(n12813), .B(n12814), .Z(n12552) );
  XOR2_X1 U12852 ( .A(n12815), .B(n12816), .Z(n12813) );
  NOR2_X1 U12853 ( .A1(n12638), .A2(n7415), .ZN(n12816) );
  NAND2_X1 U12854 ( .A1(a_12_), .A2(n12812), .ZN(n12553) );
  NAND2_X1 U12855 ( .A1(n12697), .A2(n12817), .ZN(n12812) );
  NAND2_X1 U12856 ( .A1(n12696), .A2(n12698), .ZN(n12817) );
  NAND2_X1 U12857 ( .A1(n12818), .A2(n12819), .ZN(n12698) );
  NAND2_X1 U12858 ( .A1(a_13_), .A2(b_10_), .ZN(n12819) );
  INV_X1 U12859 ( .A(n12820), .ZN(n12818) );
  XOR2_X1 U12860 ( .A(n12821), .B(n12822), .Z(n12696) );
  XOR2_X1 U12861 ( .A(n12823), .B(n12824), .Z(n12821) );
  NOR2_X1 U12862 ( .A1(n12638), .A2(n7727), .ZN(n12824) );
  NAND2_X1 U12863 ( .A1(a_13_), .A2(n12820), .ZN(n12697) );
  NAND2_X1 U12864 ( .A1(n12693), .A2(n12825), .ZN(n12820) );
  NAND2_X1 U12865 ( .A1(n12692), .A2(n12694), .ZN(n12825) );
  NAND2_X1 U12866 ( .A1(n12826), .A2(n12827), .ZN(n12694) );
  NAND2_X1 U12867 ( .A1(a_14_), .A2(b_10_), .ZN(n12827) );
  INV_X1 U12868 ( .A(n12828), .ZN(n12826) );
  XNOR2_X1 U12869 ( .A(n12829), .B(n12830), .ZN(n12692) );
  XOR2_X1 U12870 ( .A(n12831), .B(n12832), .Z(n12830) );
  NAND2_X1 U12871 ( .A1(a_15_), .A2(b_9_), .ZN(n12832) );
  NAND2_X1 U12872 ( .A1(a_14_), .A2(n12828), .ZN(n12693) );
  NAND2_X1 U12873 ( .A1(n12689), .A2(n12833), .ZN(n12828) );
  NAND2_X1 U12874 ( .A1(n12688), .A2(n12690), .ZN(n12833) );
  NAND2_X1 U12875 ( .A1(n12834), .A2(n12835), .ZN(n12690) );
  NAND2_X1 U12876 ( .A1(a_15_), .A2(b_10_), .ZN(n12835) );
  INV_X1 U12877 ( .A(n12836), .ZN(n12834) );
  XOR2_X1 U12878 ( .A(n12837), .B(n12838), .Z(n12688) );
  XOR2_X1 U12879 ( .A(n12839), .B(n12840), .Z(n12837) );
  NOR2_X1 U12880 ( .A1(n12638), .A2(n7736), .ZN(n12840) );
  NAND2_X1 U12881 ( .A1(a_15_), .A2(n12836), .ZN(n12689) );
  NAND2_X1 U12882 ( .A1(n12685), .A2(n12841), .ZN(n12836) );
  NAND2_X1 U12883 ( .A1(n12684), .A2(n12686), .ZN(n12841) );
  NAND2_X1 U12884 ( .A1(n12842), .A2(n12843), .ZN(n12686) );
  NAND2_X1 U12885 ( .A1(a_16_), .A2(b_10_), .ZN(n12843) );
  INV_X1 U12886 ( .A(n12844), .ZN(n12842) );
  XOR2_X1 U12887 ( .A(n12845), .B(n12846), .Z(n12684) );
  XOR2_X1 U12888 ( .A(n12847), .B(n12848), .Z(n12845) );
  NOR2_X1 U12889 ( .A1(n12638), .A2(n7397), .ZN(n12848) );
  NAND2_X1 U12890 ( .A1(a_16_), .A2(n12844), .ZN(n12685) );
  NAND2_X1 U12891 ( .A1(n12849), .A2(n12850), .ZN(n12844) );
  NAND2_X1 U12892 ( .A1(n12851), .A2(a_17_), .ZN(n12850) );
  NOR2_X1 U12893 ( .A1(n12852), .A2(n12422), .ZN(n12851) );
  NOR2_X1 U12894 ( .A1(n12681), .A2(n12679), .ZN(n12852) );
  NAND2_X1 U12895 ( .A1(n12679), .A2(n12681), .ZN(n12849) );
  NAND2_X1 U12896 ( .A1(n12853), .A2(n12854), .ZN(n12681) );
  NAND2_X1 U12897 ( .A1(n12678), .A2(n12855), .ZN(n12854) );
  NAND2_X1 U12898 ( .A1(n12677), .A2(n12676), .ZN(n12855) );
  NOR2_X1 U12899 ( .A1(n7745), .A2(n12422), .ZN(n12678) );
  OR2_X1 U12900 ( .A1(n12676), .A2(n12677), .ZN(n12853) );
  AND2_X1 U12901 ( .A1(n12856), .A2(n12857), .ZN(n12677) );
  NAND2_X1 U12902 ( .A1(n12586), .A2(n12858), .ZN(n12857) );
  NAND2_X1 U12903 ( .A1(n12585), .A2(n12584), .ZN(n12858) );
  NOR2_X1 U12904 ( .A1(n7750), .A2(n12422), .ZN(n12586) );
  OR2_X1 U12905 ( .A1(n12584), .A2(n12585), .ZN(n12856) );
  AND2_X1 U12906 ( .A1(n12859), .A2(n12860), .ZN(n12585) );
  NAND2_X1 U12907 ( .A1(n12674), .A2(n12861), .ZN(n12860) );
  NAND2_X1 U12908 ( .A1(n12673), .A2(n12672), .ZN(n12861) );
  NOR2_X1 U12909 ( .A1(n12422), .A2(n7755), .ZN(n12674) );
  OR2_X1 U12910 ( .A1(n12672), .A2(n12673), .ZN(n12859) );
  AND2_X1 U12911 ( .A1(n12862), .A2(n12863), .ZN(n12673) );
  NAND2_X1 U12912 ( .A1(n12864), .A2(b_10_), .ZN(n12863) );
  NOR2_X1 U12913 ( .A1(n12865), .A2(n7760), .ZN(n12864) );
  NOR2_X1 U12914 ( .A1(n12668), .A2(n12669), .ZN(n12865) );
  NAND2_X1 U12915 ( .A1(n12668), .A2(n12669), .ZN(n12862) );
  NAND2_X1 U12916 ( .A1(n12866), .A2(n12867), .ZN(n12669) );
  NAND2_X1 U12917 ( .A1(n12868), .A2(a_22_), .ZN(n12867) );
  NOR2_X1 U12918 ( .A1(n12869), .A2(n12422), .ZN(n12868) );
  NOR2_X1 U12919 ( .A1(n12664), .A2(n12665), .ZN(n12869) );
  NAND2_X1 U12920 ( .A1(n12664), .A2(n12665), .ZN(n12866) );
  NAND2_X1 U12921 ( .A1(n12870), .A2(n12871), .ZN(n12665) );
  NAND2_X1 U12922 ( .A1(n12662), .A2(n12872), .ZN(n12871) );
  OR2_X1 U12923 ( .A1(n12660), .A2(n12661), .ZN(n12872) );
  NOR2_X1 U12924 ( .A1(n12422), .A2(n8014), .ZN(n12662) );
  NAND2_X1 U12925 ( .A1(n12660), .A2(n12661), .ZN(n12870) );
  NAND2_X1 U12926 ( .A1(n12873), .A2(n12874), .ZN(n12661) );
  NAND2_X1 U12927 ( .A1(n12875), .A2(a_24_), .ZN(n12874) );
  NOR2_X1 U12928 ( .A1(n12876), .A2(n12422), .ZN(n12875) );
  NOR2_X1 U12929 ( .A1(n12656), .A2(n12657), .ZN(n12876) );
  NAND2_X1 U12930 ( .A1(n12656), .A2(n12657), .ZN(n12873) );
  NAND2_X1 U12931 ( .A1(n12877), .A2(n12878), .ZN(n12657) );
  NAND2_X1 U12932 ( .A1(n12654), .A2(n12879), .ZN(n12878) );
  OR2_X1 U12933 ( .A1(n12652), .A2(n12653), .ZN(n12879) );
  NOR2_X1 U12934 ( .A1(n12422), .A2(n8022), .ZN(n12654) );
  NAND2_X1 U12935 ( .A1(n12652), .A2(n12653), .ZN(n12877) );
  NAND2_X1 U12936 ( .A1(n12649), .A2(n12880), .ZN(n12653) );
  NAND2_X1 U12937 ( .A1(n12648), .A2(n12650), .ZN(n12880) );
  NAND2_X1 U12938 ( .A1(n12881), .A2(n12882), .ZN(n12650) );
  NAND2_X1 U12939 ( .A1(a_26_), .A2(b_10_), .ZN(n12882) );
  INV_X1 U12940 ( .A(n12883), .ZN(n12881) );
  XNOR2_X1 U12941 ( .A(n12884), .B(n12885), .ZN(n12648) );
  NAND2_X1 U12942 ( .A1(n12886), .A2(n12887), .ZN(n12884) );
  NAND2_X1 U12943 ( .A1(a_26_), .A2(n12883), .ZN(n12649) );
  NAND2_X1 U12944 ( .A1(n12617), .A2(n12888), .ZN(n12883) );
  NAND2_X1 U12945 ( .A1(n12616), .A2(n12618), .ZN(n12888) );
  NAND2_X1 U12946 ( .A1(n12889), .A2(n12890), .ZN(n12618) );
  NAND2_X1 U12947 ( .A1(a_27_), .A2(b_10_), .ZN(n12890) );
  INV_X1 U12948 ( .A(n12891), .ZN(n12889) );
  XNOR2_X1 U12949 ( .A(n12892), .B(n12893), .ZN(n12616) );
  XOR2_X1 U12950 ( .A(n12894), .B(n12895), .Z(n12893) );
  NAND2_X1 U12951 ( .A1(a_28_), .A2(b_9_), .ZN(n12895) );
  NAND2_X1 U12952 ( .A1(a_27_), .A2(n12891), .ZN(n12617) );
  NAND2_X1 U12953 ( .A1(n12896), .A2(n12897), .ZN(n12891) );
  NAND2_X1 U12954 ( .A1(n12898), .A2(a_28_), .ZN(n12897) );
  NOR2_X1 U12955 ( .A1(n12899), .A2(n12422), .ZN(n12898) );
  NOR2_X1 U12956 ( .A1(n12623), .A2(n12625), .ZN(n12899) );
  NAND2_X1 U12957 ( .A1(n12623), .A2(n12625), .ZN(n12896) );
  NAND2_X1 U12958 ( .A1(n12900), .A2(n12901), .ZN(n12625) );
  NAND2_X1 U12959 ( .A1(n12644), .A2(n12902), .ZN(n12901) );
  NAND2_X1 U12960 ( .A1(n12646), .A2(n12645), .ZN(n12902) );
  NOR2_X1 U12961 ( .A1(n12422), .A2(n7337), .ZN(n12644) );
  OR2_X1 U12962 ( .A1(n12645), .A2(n12646), .ZN(n12900) );
  AND2_X1 U12963 ( .A1(n12903), .A2(n12904), .ZN(n12646) );
  NAND2_X1 U12964 ( .A1(n12905), .A2(b_8_), .ZN(n12904) );
  NOR2_X1 U12965 ( .A1(n12906), .A2(n7817), .ZN(n12905) );
  NOR2_X1 U12966 ( .A1(n7816), .A2(n12638), .ZN(n12906) );
  NAND2_X1 U12967 ( .A1(n12907), .A2(b_9_), .ZN(n12903) );
  NOR2_X1 U12968 ( .A1(n12908), .A2(n8052), .ZN(n12907) );
  NOR2_X1 U12969 ( .A1(n7810), .A2(n12909), .ZN(n12908) );
  NAND2_X1 U12970 ( .A1(n12910), .A2(n12642), .ZN(n12645) );
  INV_X1 U12971 ( .A(n8055), .ZN(n12642) );
  NOR2_X1 U12972 ( .A1(n12638), .A2(n12422), .ZN(n12910) );
  XOR2_X1 U12973 ( .A(n12911), .B(n12912), .Z(n12623) );
  XOR2_X1 U12974 ( .A(n12913), .B(n12914), .Z(n12911) );
  XNOR2_X1 U12975 ( .A(n12915), .B(n12916), .ZN(n12652) );
  NAND2_X1 U12976 ( .A1(n12917), .A2(n12918), .ZN(n12915) );
  XOR2_X1 U12977 ( .A(n12919), .B(n12920), .Z(n12656) );
  XOR2_X1 U12978 ( .A(n12921), .B(n12922), .Z(n12919) );
  XOR2_X1 U12979 ( .A(n12923), .B(n12924), .Z(n12660) );
  XOR2_X1 U12980 ( .A(n12925), .B(n12926), .Z(n12923) );
  NOR2_X1 U12981 ( .A1(n12638), .A2(n7774), .ZN(n12926) );
  XNOR2_X1 U12982 ( .A(n12927), .B(n12928), .ZN(n12664) );
  XNOR2_X1 U12983 ( .A(n12929), .B(n12930), .ZN(n12928) );
  XNOR2_X1 U12984 ( .A(n12931), .B(n12932), .ZN(n12668) );
  XNOR2_X1 U12985 ( .A(n12933), .B(n12934), .ZN(n12932) );
  XNOR2_X1 U12986 ( .A(n12935), .B(n12936), .ZN(n12672) );
  XOR2_X1 U12987 ( .A(n12937), .B(n12938), .Z(n12935) );
  NOR2_X1 U12988 ( .A1(n7760), .A2(n12638), .ZN(n12938) );
  XNOR2_X1 U12989 ( .A(n12939), .B(n12940), .ZN(n12584) );
  XNOR2_X1 U12990 ( .A(n12941), .B(n12942), .ZN(n12939) );
  NAND2_X1 U12991 ( .A1(b_9_), .A2(a_20_), .ZN(n12941) );
  XNOR2_X1 U12992 ( .A(n12943), .B(n12944), .ZN(n12676) );
  XOR2_X1 U12993 ( .A(n12945), .B(n12946), .Z(n12943) );
  NOR2_X1 U12994 ( .A1(n12638), .A2(n7750), .ZN(n12946) );
  XOR2_X1 U12995 ( .A(n12947), .B(n12948), .Z(n12679) );
  XOR2_X1 U12996 ( .A(n12949), .B(n12950), .Z(n12947) );
  NOR2_X1 U12997 ( .A1(n12638), .A2(n7745), .ZN(n12950) );
  XOR2_X1 U12998 ( .A(n12951), .B(n12952), .Z(n12704) );
  XNOR2_X1 U12999 ( .A(n12953), .B(n12954), .ZN(n12951) );
  NAND2_X1 U13000 ( .A1(b_9_), .A2(a_11_), .ZN(n12953) );
  XNOR2_X1 U13001 ( .A(n12955), .B(n12956), .ZN(n12716) );
  XOR2_X1 U13002 ( .A(n12957), .B(n12958), .Z(n12955) );
  NOR2_X1 U13003 ( .A1(n12638), .A2(n7699), .ZN(n12958) );
  XOR2_X1 U13004 ( .A(n12959), .B(n12960), .Z(n12719) );
  XOR2_X1 U13005 ( .A(n12961), .B(n12962), .Z(n12959) );
  NOR2_X1 U13006 ( .A1(n12638), .A2(n7445), .ZN(n12962) );
  XOR2_X1 U13007 ( .A(n12963), .B(n12964), .Z(n12723) );
  XOR2_X1 U13008 ( .A(n12965), .B(n12966), .Z(n12963) );
  NOR2_X1 U13009 ( .A1(n12638), .A2(n7450), .ZN(n12966) );
  XOR2_X1 U13010 ( .A(n12967), .B(n12968), .Z(n12727) );
  XOR2_X1 U13011 ( .A(n12969), .B(n12970), .Z(n12967) );
  NOR2_X1 U13012 ( .A1(n12638), .A2(n7455), .ZN(n12970) );
  XOR2_X1 U13013 ( .A(n12971), .B(n12972), .Z(n12731) );
  XOR2_X1 U13014 ( .A(n12973), .B(n12974), .Z(n12971) );
  NOR2_X1 U13015 ( .A1(n12638), .A2(n7682), .ZN(n12974) );
  XNOR2_X1 U13016 ( .A(n12975), .B(n12976), .ZN(n12735) );
  XOR2_X1 U13017 ( .A(n12977), .B(n12978), .Z(n12976) );
  NAND2_X1 U13018 ( .A1(a_3_), .A2(b_9_), .ZN(n12978) );
  XNOR2_X1 U13019 ( .A(n12979), .B(n12980), .ZN(n12740) );
  XOR2_X1 U13020 ( .A(n12981), .B(n12982), .Z(n12980) );
  NAND2_X1 U13021 ( .A1(a_2_), .A2(b_9_), .ZN(n12982) );
  XOR2_X1 U13022 ( .A(n12983), .B(n12984), .Z(n12263) );
  XOR2_X1 U13023 ( .A(n12985), .B(n12986), .Z(n12983) );
  NOR2_X1 U13024 ( .A1(n12638), .A2(n7669), .ZN(n12986) );
  XOR2_X1 U13025 ( .A(n12987), .B(n12988), .Z(n12503) );
  XOR2_X1 U13026 ( .A(n12989), .B(n12990), .Z(n12987) );
  NAND2_X1 U13027 ( .A1(n12991), .A2(n12748), .ZN(n7315) );
  OR2_X1 U13028 ( .A1(n12748), .A2(n12991), .ZN(n7316) );
  XNOR2_X1 U13029 ( .A(n12992), .B(n12993), .ZN(n12991) );
  NAND2_X1 U13030 ( .A1(n12994), .A2(n12752), .ZN(n12748) );
  NAND2_X1 U13031 ( .A1(n12995), .A2(n12996), .ZN(n12752) );
  NAND2_X1 U13032 ( .A1(n12990), .A2(n12997), .ZN(n12996) );
  OR2_X1 U13033 ( .A1(n12988), .A2(n12989), .ZN(n12997) );
  NOR2_X1 U13034 ( .A1(n12638), .A2(n7478), .ZN(n12990) );
  NAND2_X1 U13035 ( .A1(n12988), .A2(n12989), .ZN(n12995) );
  NAND2_X1 U13036 ( .A1(n12998), .A2(n12999), .ZN(n12989) );
  NAND2_X1 U13037 ( .A1(n13000), .A2(a_1_), .ZN(n12999) );
  NOR2_X1 U13038 ( .A1(n13001), .A2(n12638), .ZN(n13000) );
  NOR2_X1 U13039 ( .A1(n12985), .A2(n12984), .ZN(n13001) );
  NAND2_X1 U13040 ( .A1(n12984), .A2(n12985), .ZN(n12998) );
  NAND2_X1 U13041 ( .A1(n13002), .A2(n13003), .ZN(n12985) );
  NAND2_X1 U13042 ( .A1(n13004), .A2(a_2_), .ZN(n13003) );
  NOR2_X1 U13043 ( .A1(n13005), .A2(n12638), .ZN(n13004) );
  NOR2_X1 U13044 ( .A1(n12981), .A2(n12979), .ZN(n13005) );
  NAND2_X1 U13045 ( .A1(n12979), .A2(n12981), .ZN(n13002) );
  NAND2_X1 U13046 ( .A1(n13006), .A2(n13007), .ZN(n12981) );
  NAND2_X1 U13047 ( .A1(n13008), .A2(a_3_), .ZN(n13007) );
  NOR2_X1 U13048 ( .A1(n13009), .A2(n12638), .ZN(n13008) );
  NOR2_X1 U13049 ( .A1(n12977), .A2(n12975), .ZN(n13009) );
  NAND2_X1 U13050 ( .A1(n12975), .A2(n12977), .ZN(n13006) );
  NAND2_X1 U13051 ( .A1(n13010), .A2(n13011), .ZN(n12977) );
  NAND2_X1 U13052 ( .A1(n13012), .A2(a_4_), .ZN(n13011) );
  NOR2_X1 U13053 ( .A1(n13013), .A2(n12638), .ZN(n13012) );
  NOR2_X1 U13054 ( .A1(n12973), .A2(n12972), .ZN(n13013) );
  NAND2_X1 U13055 ( .A1(n12972), .A2(n12973), .ZN(n13010) );
  NAND2_X1 U13056 ( .A1(n13014), .A2(n13015), .ZN(n12973) );
  NAND2_X1 U13057 ( .A1(n13016), .A2(a_5_), .ZN(n13015) );
  NOR2_X1 U13058 ( .A1(n13017), .A2(n12638), .ZN(n13016) );
  NOR2_X1 U13059 ( .A1(n12969), .A2(n12968), .ZN(n13017) );
  NAND2_X1 U13060 ( .A1(n12968), .A2(n12969), .ZN(n13014) );
  NAND2_X1 U13061 ( .A1(n13018), .A2(n13019), .ZN(n12969) );
  NAND2_X1 U13062 ( .A1(n13020), .A2(a_6_), .ZN(n13019) );
  NOR2_X1 U13063 ( .A1(n13021), .A2(n12638), .ZN(n13020) );
  NOR2_X1 U13064 ( .A1(n12964), .A2(n12965), .ZN(n13021) );
  NAND2_X1 U13065 ( .A1(n12964), .A2(n12965), .ZN(n13018) );
  NAND2_X1 U13066 ( .A1(n13022), .A2(n13023), .ZN(n12965) );
  NAND2_X1 U13067 ( .A1(n13024), .A2(a_7_), .ZN(n13023) );
  NOR2_X1 U13068 ( .A1(n13025), .A2(n12638), .ZN(n13024) );
  NOR2_X1 U13069 ( .A1(n12961), .A2(n12960), .ZN(n13025) );
  NAND2_X1 U13070 ( .A1(n12960), .A2(n12961), .ZN(n13022) );
  NAND2_X1 U13071 ( .A1(n13026), .A2(n13027), .ZN(n12961) );
  NAND2_X1 U13072 ( .A1(n13028), .A2(a_8_), .ZN(n13027) );
  NOR2_X1 U13073 ( .A1(n13029), .A2(n12638), .ZN(n13028) );
  NOR2_X1 U13074 ( .A1(n12957), .A2(n12956), .ZN(n13029) );
  NAND2_X1 U13075 ( .A1(n12956), .A2(n12957), .ZN(n13026) );
  NAND2_X1 U13076 ( .A1(n13030), .A2(n13031), .ZN(n12957) );
  NAND2_X1 U13077 ( .A1(n12786), .A2(n13032), .ZN(n13031) );
  OR2_X1 U13078 ( .A1(n12787), .A2(n12788), .ZN(n13032) );
  XNOR2_X1 U13079 ( .A(n13033), .B(n13034), .ZN(n12786) );
  XNOR2_X1 U13080 ( .A(n13035), .B(n13036), .ZN(n13034) );
  NAND2_X1 U13081 ( .A1(n12788), .A2(n12787), .ZN(n13030) );
  NAND2_X1 U13082 ( .A1(n13037), .A2(n13038), .ZN(n12787) );
  NAND2_X1 U13083 ( .A1(n13039), .A2(a_10_), .ZN(n13038) );
  NOR2_X1 U13084 ( .A1(n13040), .A2(n12638), .ZN(n13039) );
  NOR2_X1 U13085 ( .A1(n12795), .A2(n12794), .ZN(n13040) );
  NAND2_X1 U13086 ( .A1(n12794), .A2(n12795), .ZN(n13037) );
  NAND2_X1 U13087 ( .A1(n13041), .A2(n13042), .ZN(n12795) );
  NAND2_X1 U13088 ( .A1(n13043), .A2(b_9_), .ZN(n13042) );
  NOR2_X1 U13089 ( .A1(n13044), .A2(n7424), .ZN(n13043) );
  NOR2_X1 U13090 ( .A1(n12952), .A2(n12954), .ZN(n13044) );
  NAND2_X1 U13091 ( .A1(n12952), .A2(n12954), .ZN(n13041) );
  NAND2_X1 U13092 ( .A1(n13045), .A2(n13046), .ZN(n12954) );
  NAND2_X1 U13093 ( .A1(n13047), .A2(a_12_), .ZN(n13046) );
  NOR2_X1 U13094 ( .A1(n13048), .A2(n12638), .ZN(n13047) );
  NOR2_X1 U13095 ( .A1(n12807), .A2(n12805), .ZN(n13048) );
  NAND2_X1 U13096 ( .A1(n12805), .A2(n12807), .ZN(n13045) );
  NAND2_X1 U13097 ( .A1(n13049), .A2(n13050), .ZN(n12807) );
  NAND2_X1 U13098 ( .A1(n13051), .A2(a_13_), .ZN(n13050) );
  NOR2_X1 U13099 ( .A1(n13052), .A2(n12638), .ZN(n13051) );
  NOR2_X1 U13100 ( .A1(n12814), .A2(n12815), .ZN(n13052) );
  NAND2_X1 U13101 ( .A1(n12814), .A2(n12815), .ZN(n13049) );
  NAND2_X1 U13102 ( .A1(n13053), .A2(n13054), .ZN(n12815) );
  NAND2_X1 U13103 ( .A1(n13055), .A2(a_14_), .ZN(n13054) );
  NOR2_X1 U13104 ( .A1(n13056), .A2(n12638), .ZN(n13055) );
  NOR2_X1 U13105 ( .A1(n12823), .A2(n12822), .ZN(n13056) );
  NAND2_X1 U13106 ( .A1(n12822), .A2(n12823), .ZN(n13053) );
  NAND2_X1 U13107 ( .A1(n13057), .A2(n13058), .ZN(n12823) );
  NAND2_X1 U13108 ( .A1(n13059), .A2(a_15_), .ZN(n13058) );
  NOR2_X1 U13109 ( .A1(n13060), .A2(n12638), .ZN(n13059) );
  NOR2_X1 U13110 ( .A1(n12831), .A2(n12829), .ZN(n13060) );
  NAND2_X1 U13111 ( .A1(n12829), .A2(n12831), .ZN(n13057) );
  NAND2_X1 U13112 ( .A1(n13061), .A2(n13062), .ZN(n12831) );
  NAND2_X1 U13113 ( .A1(n13063), .A2(a_16_), .ZN(n13062) );
  NOR2_X1 U13114 ( .A1(n13064), .A2(n12638), .ZN(n13063) );
  NOR2_X1 U13115 ( .A1(n12838), .A2(n12839), .ZN(n13064) );
  NAND2_X1 U13116 ( .A1(n12838), .A2(n12839), .ZN(n13061) );
  NAND2_X1 U13117 ( .A1(n13065), .A2(n13066), .ZN(n12839) );
  NAND2_X1 U13118 ( .A1(n13067), .A2(a_17_), .ZN(n13066) );
  NOR2_X1 U13119 ( .A1(n13068), .A2(n12638), .ZN(n13067) );
  NOR2_X1 U13120 ( .A1(n12846), .A2(n12847), .ZN(n13068) );
  NAND2_X1 U13121 ( .A1(n12846), .A2(n12847), .ZN(n13065) );
  NAND2_X1 U13122 ( .A1(n13069), .A2(n13070), .ZN(n12847) );
  NAND2_X1 U13123 ( .A1(n13071), .A2(a_18_), .ZN(n13070) );
  NOR2_X1 U13124 ( .A1(n13072), .A2(n12638), .ZN(n13071) );
  NOR2_X1 U13125 ( .A1(n12948), .A2(n12949), .ZN(n13072) );
  NAND2_X1 U13126 ( .A1(n12948), .A2(n12949), .ZN(n13069) );
  NAND2_X1 U13127 ( .A1(n13073), .A2(n13074), .ZN(n12949) );
  NAND2_X1 U13128 ( .A1(n13075), .A2(a_19_), .ZN(n13074) );
  NOR2_X1 U13129 ( .A1(n13076), .A2(n12638), .ZN(n13075) );
  NOR2_X1 U13130 ( .A1(n12945), .A2(n12944), .ZN(n13076) );
  NAND2_X1 U13131 ( .A1(n12944), .A2(n12945), .ZN(n13073) );
  NAND2_X1 U13132 ( .A1(n13077), .A2(n13078), .ZN(n12945) );
  NAND2_X1 U13133 ( .A1(n13079), .A2(b_9_), .ZN(n13078) );
  NOR2_X1 U13134 ( .A1(n13080), .A2(n7755), .ZN(n13079) );
  NOR2_X1 U13135 ( .A1(n12942), .A2(n12940), .ZN(n13080) );
  NAND2_X1 U13136 ( .A1(n12940), .A2(n12942), .ZN(n13077) );
  NAND2_X1 U13137 ( .A1(n13081), .A2(n13082), .ZN(n12942) );
  NAND2_X1 U13138 ( .A1(n13083), .A2(b_9_), .ZN(n13082) );
  NOR2_X1 U13139 ( .A1(n13084), .A2(n7760), .ZN(n13083) );
  NOR2_X1 U13140 ( .A1(n12937), .A2(n12936), .ZN(n13084) );
  NAND2_X1 U13141 ( .A1(n12936), .A2(n12937), .ZN(n13081) );
  NAND2_X1 U13142 ( .A1(n13085), .A2(n13086), .ZN(n12937) );
  NAND2_X1 U13143 ( .A1(n12934), .A2(n13087), .ZN(n13086) );
  OR2_X1 U13144 ( .A1(n12931), .A2(n12933), .ZN(n13087) );
  NOR2_X1 U13145 ( .A1(n7765), .A2(n12638), .ZN(n12934) );
  NAND2_X1 U13146 ( .A1(n12931), .A2(n12933), .ZN(n13085) );
  NAND2_X1 U13147 ( .A1(n13088), .A2(n13089), .ZN(n12933) );
  NAND2_X1 U13148 ( .A1(n12930), .A2(n13090), .ZN(n13089) );
  OR2_X1 U13149 ( .A1(n12927), .A2(n12929), .ZN(n13090) );
  NOR2_X1 U13150 ( .A1(n12638), .A2(n8014), .ZN(n12930) );
  NAND2_X1 U13151 ( .A1(n12927), .A2(n12929), .ZN(n13088) );
  NAND2_X1 U13152 ( .A1(n13091), .A2(n13092), .ZN(n12929) );
  NAND2_X1 U13153 ( .A1(n13093), .A2(a_24_), .ZN(n13092) );
  NOR2_X1 U13154 ( .A1(n13094), .A2(n12638), .ZN(n13093) );
  NOR2_X1 U13155 ( .A1(n12924), .A2(n12925), .ZN(n13094) );
  NAND2_X1 U13156 ( .A1(n12924), .A2(n12925), .ZN(n13091) );
  NAND2_X1 U13157 ( .A1(n13095), .A2(n13096), .ZN(n12925) );
  NAND2_X1 U13158 ( .A1(n12922), .A2(n13097), .ZN(n13096) );
  OR2_X1 U13159 ( .A1(n12920), .A2(n12921), .ZN(n13097) );
  NOR2_X1 U13160 ( .A1(n12638), .A2(n8022), .ZN(n12922) );
  NAND2_X1 U13161 ( .A1(n12920), .A2(n12921), .ZN(n13095) );
  NAND2_X1 U13162 ( .A1(n12917), .A2(n13098), .ZN(n12921) );
  NAND2_X1 U13163 ( .A1(n12916), .A2(n12918), .ZN(n13098) );
  NAND2_X1 U13164 ( .A1(n13099), .A2(n13100), .ZN(n12918) );
  NAND2_X1 U13165 ( .A1(a_26_), .A2(b_9_), .ZN(n13100) );
  INV_X1 U13166 ( .A(n13101), .ZN(n13099) );
  XNOR2_X1 U13167 ( .A(n13102), .B(n13103), .ZN(n12916) );
  NAND2_X1 U13168 ( .A1(n13104), .A2(n13105), .ZN(n13102) );
  NAND2_X1 U13169 ( .A1(a_26_), .A2(n13101), .ZN(n12917) );
  NAND2_X1 U13170 ( .A1(n12886), .A2(n13106), .ZN(n13101) );
  NAND2_X1 U13171 ( .A1(n12885), .A2(n12887), .ZN(n13106) );
  NAND2_X1 U13172 ( .A1(n13107), .A2(n13108), .ZN(n12887) );
  NAND2_X1 U13173 ( .A1(a_27_), .A2(b_9_), .ZN(n13108) );
  INV_X1 U13174 ( .A(n13109), .ZN(n13107) );
  XNOR2_X1 U13175 ( .A(n13110), .B(n13111), .ZN(n12885) );
  XOR2_X1 U13176 ( .A(n13112), .B(n13113), .Z(n13111) );
  NAND2_X1 U13177 ( .A1(a_28_), .A2(b_8_), .ZN(n13113) );
  NAND2_X1 U13178 ( .A1(a_27_), .A2(n13109), .ZN(n12886) );
  NAND2_X1 U13179 ( .A1(n13114), .A2(n13115), .ZN(n13109) );
  NAND2_X1 U13180 ( .A1(n13116), .A2(a_28_), .ZN(n13115) );
  NOR2_X1 U13181 ( .A1(n13117), .A2(n12638), .ZN(n13116) );
  NOR2_X1 U13182 ( .A1(n12892), .A2(n12894), .ZN(n13117) );
  NAND2_X1 U13183 ( .A1(n12892), .A2(n12894), .ZN(n13114) );
  NAND2_X1 U13184 ( .A1(n13118), .A2(n13119), .ZN(n12894) );
  NAND2_X1 U13185 ( .A1(n12912), .A2(n13120), .ZN(n13119) );
  NAND2_X1 U13186 ( .A1(n12914), .A2(n12913), .ZN(n13120) );
  NOR2_X1 U13187 ( .A1(n12638), .A2(n7337), .ZN(n12912) );
  OR2_X1 U13188 ( .A1(n12913), .A2(n12914), .ZN(n13118) );
  AND2_X1 U13189 ( .A1(n13121), .A2(n13122), .ZN(n12914) );
  NAND2_X1 U13190 ( .A1(n13123), .A2(b_7_), .ZN(n13122) );
  NOR2_X1 U13191 ( .A1(n13124), .A2(n7817), .ZN(n13123) );
  NOR2_X1 U13192 ( .A1(n7816), .A2(n12909), .ZN(n13124) );
  NAND2_X1 U13193 ( .A1(n13125), .A2(b_8_), .ZN(n13121) );
  NOR2_X1 U13194 ( .A1(n13126), .A2(n8052), .ZN(n13125) );
  NOR2_X1 U13195 ( .A1(n7810), .A2(n13127), .ZN(n13126) );
  NAND2_X1 U13196 ( .A1(n13128), .A2(b_8_), .ZN(n12913) );
  NOR2_X1 U13197 ( .A1(n12638), .A2(n8055), .ZN(n13128) );
  XOR2_X1 U13198 ( .A(n13129), .B(n13130), .Z(n12892) );
  XOR2_X1 U13199 ( .A(n13131), .B(n13132), .Z(n13129) );
  XNOR2_X1 U13200 ( .A(n13133), .B(n13134), .ZN(n12920) );
  NAND2_X1 U13201 ( .A1(n13135), .A2(n13136), .ZN(n13133) );
  XOR2_X1 U13202 ( .A(n13137), .B(n13138), .Z(n12924) );
  XOR2_X1 U13203 ( .A(n13139), .B(n13140), .Z(n13137) );
  XOR2_X1 U13204 ( .A(n13141), .B(n13142), .Z(n12927) );
  XOR2_X1 U13205 ( .A(n13143), .B(n13144), .Z(n13141) );
  NOR2_X1 U13206 ( .A1(n12909), .A2(n7774), .ZN(n13144) );
  XOR2_X1 U13207 ( .A(n13145), .B(n13146), .Z(n12931) );
  XOR2_X1 U13208 ( .A(n13147), .B(n13148), .Z(n13145) );
  NOR2_X1 U13209 ( .A1(n8014), .A2(n12909), .ZN(n13148) );
  XNOR2_X1 U13210 ( .A(n13149), .B(n13150), .ZN(n12936) );
  XNOR2_X1 U13211 ( .A(n13151), .B(n13152), .ZN(n13149) );
  XNOR2_X1 U13212 ( .A(n13153), .B(n13154), .ZN(n12940) );
  XNOR2_X1 U13213 ( .A(n13155), .B(n13156), .ZN(n13153) );
  XNOR2_X1 U13214 ( .A(n13157), .B(n13158), .ZN(n12944) );
  XNOR2_X1 U13215 ( .A(n13159), .B(n13160), .ZN(n13157) );
  XOR2_X1 U13216 ( .A(n13161), .B(n13162), .Z(n12948) );
  XOR2_X1 U13217 ( .A(n13163), .B(n13164), .Z(n13161) );
  XOR2_X1 U13218 ( .A(n13165), .B(n13166), .Z(n12846) );
  XOR2_X1 U13219 ( .A(n13167), .B(n13168), .Z(n13165) );
  NOR2_X1 U13220 ( .A1(n12909), .A2(n7745), .ZN(n13168) );
  XNOR2_X1 U13221 ( .A(n13169), .B(n13170), .ZN(n12838) );
  NAND2_X1 U13222 ( .A1(n13171), .A2(n13172), .ZN(n13169) );
  XNOR2_X1 U13223 ( .A(n13173), .B(n13174), .ZN(n12829) );
  NAND2_X1 U13224 ( .A1(n13175), .A2(n13176), .ZN(n13173) );
  XNOR2_X1 U13225 ( .A(n13177), .B(n13178), .ZN(n12822) );
  XNOR2_X1 U13226 ( .A(n13179), .B(n13180), .ZN(n13178) );
  XNOR2_X1 U13227 ( .A(n13181), .B(n13182), .ZN(n12814) );
  XOR2_X1 U13228 ( .A(n13183), .B(n13184), .Z(n13182) );
  NAND2_X1 U13229 ( .A1(a_14_), .A2(b_8_), .ZN(n13184) );
  XNOR2_X1 U13230 ( .A(n13185), .B(n13186), .ZN(n12805) );
  XNOR2_X1 U13231 ( .A(n13187), .B(n13188), .ZN(n13185) );
  XNOR2_X1 U13232 ( .A(n13189), .B(n13190), .ZN(n12952) );
  XNOR2_X1 U13233 ( .A(n13191), .B(n13192), .ZN(n13190) );
  XNOR2_X1 U13234 ( .A(n13193), .B(n13194), .ZN(n12794) );
  XNOR2_X1 U13235 ( .A(n13195), .B(n13196), .ZN(n13193) );
  XNOR2_X1 U13236 ( .A(n13197), .B(n13198), .ZN(n12956) );
  XNOR2_X1 U13237 ( .A(n13199), .B(n13200), .ZN(n13198) );
  XNOR2_X1 U13238 ( .A(n13201), .B(n13202), .ZN(n12960) );
  XOR2_X1 U13239 ( .A(n13203), .B(n13204), .Z(n13202) );
  XNOR2_X1 U13240 ( .A(n13205), .B(n13206), .ZN(n12964) );
  XNOR2_X1 U13241 ( .A(n13207), .B(n13208), .ZN(n13206) );
  XNOR2_X1 U13242 ( .A(n13209), .B(n13210), .ZN(n12968) );
  XNOR2_X1 U13243 ( .A(n13211), .B(n13212), .ZN(n13210) );
  XOR2_X1 U13244 ( .A(n13213), .B(n13214), .Z(n12972) );
  XOR2_X1 U13245 ( .A(n13215), .B(n13216), .Z(n13213) );
  NOR2_X1 U13246 ( .A1(n12909), .A2(n7455), .ZN(n13216) );
  XNOR2_X1 U13247 ( .A(n13217), .B(n13218), .ZN(n12975) );
  XOR2_X1 U13248 ( .A(n13219), .B(n13220), .Z(n13218) );
  NAND2_X1 U13249 ( .A1(a_4_), .A2(b_8_), .ZN(n13220) );
  XOR2_X1 U13250 ( .A(n13221), .B(n13222), .Z(n12979) );
  XOR2_X1 U13251 ( .A(n13223), .B(n13224), .Z(n13221) );
  NOR2_X1 U13252 ( .A1(n12909), .A2(n7464), .ZN(n13224) );
  XOR2_X1 U13253 ( .A(n13225), .B(n13226), .Z(n12984) );
  XOR2_X1 U13254 ( .A(n13227), .B(n13228), .Z(n13225) );
  NOR2_X1 U13255 ( .A1(n12909), .A2(n7469), .ZN(n13228) );
  XOR2_X1 U13256 ( .A(n13229), .B(n13230), .Z(n12988) );
  XOR2_X1 U13257 ( .A(n13231), .B(n13232), .Z(n13229) );
  NOR2_X1 U13258 ( .A1(n12909), .A2(n7669), .ZN(n13232) );
  XOR2_X1 U13259 ( .A(n13233), .B(n12754), .Z(n12994) );
  INV_X1 U13260 ( .A(n13234), .ZN(n12754) );
  INV_X1 U13261 ( .A(n12753), .ZN(n13233) );
  XOR2_X1 U13262 ( .A(n13235), .B(n13236), .Z(n12753) );
  NOR2_X1 U13263 ( .A1(n7478), .A2(n12909), .ZN(n13236) );
  NAND2_X1 U13264 ( .A1(n13237), .A2(n13238), .ZN(n7320) );
  OR2_X1 U13265 ( .A1(n13238), .A2(n13237), .ZN(n7319) );
  NAND2_X1 U13266 ( .A1(n13239), .A2(n13240), .ZN(n13237) );
  NAND2_X1 U13267 ( .A1(n13241), .A2(n13242), .ZN(n13240) );
  XOR2_X1 U13268 ( .A(n13243), .B(n13244), .Z(n13242) );
  INV_X1 U13269 ( .A(n13245), .ZN(n13241) );
  OR2_X1 U13270 ( .A1(n12993), .A2(n12992), .ZN(n13238) );
  AND2_X1 U13271 ( .A1(n13246), .A2(n13247), .ZN(n12992) );
  NAND2_X1 U13272 ( .A1(n13248), .A2(b_8_), .ZN(n13247) );
  NOR2_X1 U13273 ( .A1(n13249), .A2(n7478), .ZN(n13248) );
  NOR2_X1 U13274 ( .A1(n13234), .A2(n13235), .ZN(n13249) );
  NAND2_X1 U13275 ( .A1(n13234), .A2(n13235), .ZN(n13246) );
  NAND2_X1 U13276 ( .A1(n13250), .A2(n13251), .ZN(n13235) );
  NAND2_X1 U13277 ( .A1(n13252), .A2(a_1_), .ZN(n13251) );
  NOR2_X1 U13278 ( .A1(n13253), .A2(n12909), .ZN(n13252) );
  NOR2_X1 U13279 ( .A1(n13230), .A2(n13231), .ZN(n13253) );
  NAND2_X1 U13280 ( .A1(n13230), .A2(n13231), .ZN(n13250) );
  NAND2_X1 U13281 ( .A1(n13254), .A2(n13255), .ZN(n13231) );
  NAND2_X1 U13282 ( .A1(n13256), .A2(a_2_), .ZN(n13255) );
  NOR2_X1 U13283 ( .A1(n13257), .A2(n12909), .ZN(n13256) );
  NOR2_X1 U13284 ( .A1(n13226), .A2(n13227), .ZN(n13257) );
  NAND2_X1 U13285 ( .A1(n13226), .A2(n13227), .ZN(n13254) );
  NAND2_X1 U13286 ( .A1(n13258), .A2(n13259), .ZN(n13227) );
  NAND2_X1 U13287 ( .A1(n13260), .A2(a_3_), .ZN(n13259) );
  NOR2_X1 U13288 ( .A1(n13261), .A2(n12909), .ZN(n13260) );
  NOR2_X1 U13289 ( .A1(n13222), .A2(n13223), .ZN(n13261) );
  NAND2_X1 U13290 ( .A1(n13222), .A2(n13223), .ZN(n13258) );
  NAND2_X1 U13291 ( .A1(n13262), .A2(n13263), .ZN(n13223) );
  NAND2_X1 U13292 ( .A1(n13264), .A2(a_4_), .ZN(n13263) );
  NOR2_X1 U13293 ( .A1(n13265), .A2(n12909), .ZN(n13264) );
  NOR2_X1 U13294 ( .A1(n13217), .A2(n13219), .ZN(n13265) );
  NAND2_X1 U13295 ( .A1(n13217), .A2(n13219), .ZN(n13262) );
  NAND2_X1 U13296 ( .A1(n13266), .A2(n13267), .ZN(n13219) );
  NAND2_X1 U13297 ( .A1(n13268), .A2(a_5_), .ZN(n13267) );
  NOR2_X1 U13298 ( .A1(n13269), .A2(n12909), .ZN(n13268) );
  NOR2_X1 U13299 ( .A1(n13214), .A2(n13215), .ZN(n13269) );
  NAND2_X1 U13300 ( .A1(n13214), .A2(n13215), .ZN(n13266) );
  NAND2_X1 U13301 ( .A1(n13270), .A2(n13271), .ZN(n13215) );
  NAND2_X1 U13302 ( .A1(n13212), .A2(n13272), .ZN(n13271) );
  OR2_X1 U13303 ( .A1(n13211), .A2(n13209), .ZN(n13272) );
  NOR2_X1 U13304 ( .A1(n7450), .A2(n12909), .ZN(n13212) );
  NAND2_X1 U13305 ( .A1(n13209), .A2(n13211), .ZN(n13270) );
  NAND2_X1 U13306 ( .A1(n13273), .A2(n13274), .ZN(n13211) );
  NAND2_X1 U13307 ( .A1(n13208), .A2(n13275), .ZN(n13274) );
  NAND2_X1 U13308 ( .A1(n13205), .A2(n13207), .ZN(n13275) );
  NOR2_X1 U13309 ( .A1(n7445), .A2(n12909), .ZN(n13208) );
  OR2_X1 U13310 ( .A1(n13205), .A2(n13207), .ZN(n13273) );
  NAND2_X1 U13311 ( .A1(n13276), .A2(n13277), .ZN(n13207) );
  NAND2_X1 U13312 ( .A1(n13278), .A2(n13204), .ZN(n13277) );
  NAND2_X1 U13313 ( .A1(n13201), .A2(n13203), .ZN(n13278) );
  OR2_X1 U13314 ( .A1(n13203), .A2(n13201), .ZN(n13276) );
  XOR2_X1 U13315 ( .A(n13279), .B(n13280), .Z(n13201) );
  XOR2_X1 U13316 ( .A(n13281), .B(n13282), .Z(n13279) );
  NOR2_X1 U13317 ( .A1(n13127), .A2(n7704), .ZN(n13282) );
  NAND2_X1 U13318 ( .A1(n13283), .A2(n13284), .ZN(n13203) );
  NAND2_X1 U13319 ( .A1(n13200), .A2(n13285), .ZN(n13284) );
  OR2_X1 U13320 ( .A1(n13199), .A2(n13197), .ZN(n13285) );
  NOR2_X1 U13321 ( .A1(n7704), .A2(n12909), .ZN(n13200) );
  NAND2_X1 U13322 ( .A1(n13197), .A2(n13199), .ZN(n13283) );
  NAND2_X1 U13323 ( .A1(n13286), .A2(n13287), .ZN(n13199) );
  NAND2_X1 U13324 ( .A1(n13036), .A2(n13288), .ZN(n13287) );
  OR2_X1 U13325 ( .A1(n13035), .A2(n13033), .ZN(n13288) );
  NOR2_X1 U13326 ( .A1(n7709), .A2(n12909), .ZN(n13036) );
  NAND2_X1 U13327 ( .A1(n13033), .A2(n13035), .ZN(n13286) );
  NAND2_X1 U13328 ( .A1(n13289), .A2(n13290), .ZN(n13035) );
  NAND2_X1 U13329 ( .A1(n13196), .A2(n13291), .ZN(n13290) );
  NAND2_X1 U13330 ( .A1(n13195), .A2(n13194), .ZN(n13291) );
  NOR2_X1 U13331 ( .A1(n12909), .A2(n7424), .ZN(n13196) );
  OR2_X1 U13332 ( .A1(n13194), .A2(n13195), .ZN(n13289) );
  AND2_X1 U13333 ( .A1(n13292), .A2(n13293), .ZN(n13195) );
  NAND2_X1 U13334 ( .A1(n13192), .A2(n13294), .ZN(n13293) );
  OR2_X1 U13335 ( .A1(n13189), .A2(n13191), .ZN(n13294) );
  NOR2_X1 U13336 ( .A1(n7718), .A2(n12909), .ZN(n13192) );
  NAND2_X1 U13337 ( .A1(n13189), .A2(n13191), .ZN(n13292) );
  NAND2_X1 U13338 ( .A1(n13295), .A2(n13296), .ZN(n13191) );
  NAND2_X1 U13339 ( .A1(n13188), .A2(n13297), .ZN(n13296) );
  NAND2_X1 U13340 ( .A1(n13187), .A2(n13186), .ZN(n13297) );
  NOR2_X1 U13341 ( .A1(n7415), .A2(n12909), .ZN(n13188) );
  OR2_X1 U13342 ( .A1(n13186), .A2(n13187), .ZN(n13295) );
  AND2_X1 U13343 ( .A1(n13298), .A2(n13299), .ZN(n13187) );
  NAND2_X1 U13344 ( .A1(n13300), .A2(a_14_), .ZN(n13299) );
  NOR2_X1 U13345 ( .A1(n13301), .A2(n12909), .ZN(n13300) );
  NOR2_X1 U13346 ( .A1(n13183), .A2(n13181), .ZN(n13301) );
  NAND2_X1 U13347 ( .A1(n13181), .A2(n13183), .ZN(n13298) );
  NAND2_X1 U13348 ( .A1(n13302), .A2(n13303), .ZN(n13183) );
  NAND2_X1 U13349 ( .A1(n13180), .A2(n13304), .ZN(n13303) );
  OR2_X1 U13350 ( .A1(n13179), .A2(n13177), .ZN(n13304) );
  NOR2_X1 U13351 ( .A1(n7406), .A2(n12909), .ZN(n13180) );
  NAND2_X1 U13352 ( .A1(n13177), .A2(n13179), .ZN(n13302) );
  NAND2_X1 U13353 ( .A1(n13175), .A2(n13305), .ZN(n13179) );
  NAND2_X1 U13354 ( .A1(n13174), .A2(n13176), .ZN(n13305) );
  NAND2_X1 U13355 ( .A1(n13306), .A2(n13307), .ZN(n13176) );
  NAND2_X1 U13356 ( .A1(a_16_), .A2(b_8_), .ZN(n13307) );
  INV_X1 U13357 ( .A(n13308), .ZN(n13306) );
  XNOR2_X1 U13358 ( .A(n13309), .B(n13310), .ZN(n13174) );
  XOR2_X1 U13359 ( .A(n13311), .B(n13312), .Z(n13310) );
  NAND2_X1 U13360 ( .A1(a_17_), .A2(b_7_), .ZN(n13312) );
  NAND2_X1 U13361 ( .A1(a_16_), .A2(n13308), .ZN(n13175) );
  NAND2_X1 U13362 ( .A1(n13171), .A2(n13313), .ZN(n13308) );
  NAND2_X1 U13363 ( .A1(n13170), .A2(n13172), .ZN(n13313) );
  NAND2_X1 U13364 ( .A1(n13314), .A2(n13315), .ZN(n13172) );
  NAND2_X1 U13365 ( .A1(a_17_), .A2(b_8_), .ZN(n13315) );
  INV_X1 U13366 ( .A(n13316), .ZN(n13314) );
  XNOR2_X1 U13367 ( .A(n13317), .B(n13318), .ZN(n13170) );
  XOR2_X1 U13368 ( .A(n13319), .B(n13320), .Z(n13318) );
  NAND2_X1 U13369 ( .A1(a_18_), .A2(b_7_), .ZN(n13320) );
  NAND2_X1 U13370 ( .A1(a_17_), .A2(n13316), .ZN(n13171) );
  NAND2_X1 U13371 ( .A1(n13321), .A2(n13322), .ZN(n13316) );
  NAND2_X1 U13372 ( .A1(n13323), .A2(a_18_), .ZN(n13322) );
  NOR2_X1 U13373 ( .A1(n13324), .A2(n12909), .ZN(n13323) );
  NOR2_X1 U13374 ( .A1(n13167), .A2(n13166), .ZN(n13324) );
  NAND2_X1 U13375 ( .A1(n13166), .A2(n13167), .ZN(n13321) );
  NAND2_X1 U13376 ( .A1(n13325), .A2(n13326), .ZN(n13167) );
  NAND2_X1 U13377 ( .A1(n13164), .A2(n13327), .ZN(n13326) );
  OR2_X1 U13378 ( .A1(n13162), .A2(n13163), .ZN(n13327) );
  NOR2_X1 U13379 ( .A1(n7750), .A2(n12909), .ZN(n13164) );
  NAND2_X1 U13380 ( .A1(n13162), .A2(n13163), .ZN(n13325) );
  NAND2_X1 U13381 ( .A1(n13328), .A2(n13329), .ZN(n13163) );
  NAND2_X1 U13382 ( .A1(n13159), .A2(n13330), .ZN(n13329) );
  NAND2_X1 U13383 ( .A1(n13160), .A2(n13158), .ZN(n13330) );
  NOR2_X1 U13384 ( .A1(n12909), .A2(n7755), .ZN(n13159) );
  OR2_X1 U13385 ( .A1(n13158), .A2(n13160), .ZN(n13328) );
  AND2_X1 U13386 ( .A1(n13331), .A2(n13332), .ZN(n13160) );
  NAND2_X1 U13387 ( .A1(n13156), .A2(n13333), .ZN(n13332) );
  NAND2_X1 U13388 ( .A1(n13155), .A2(n13154), .ZN(n13333) );
  NOR2_X1 U13389 ( .A1(n12909), .A2(n7760), .ZN(n13156) );
  OR2_X1 U13390 ( .A1(n13154), .A2(n13155), .ZN(n13331) );
  AND2_X1 U13391 ( .A1(n13334), .A2(n13335), .ZN(n13155) );
  NAND2_X1 U13392 ( .A1(n13152), .A2(n13336), .ZN(n13335) );
  NAND2_X1 U13393 ( .A1(n13151), .A2(n13150), .ZN(n13336) );
  NOR2_X1 U13394 ( .A1(n7765), .A2(n12909), .ZN(n13152) );
  OR2_X1 U13395 ( .A1(n13150), .A2(n13151), .ZN(n13334) );
  AND2_X1 U13396 ( .A1(n13337), .A2(n13338), .ZN(n13151) );
  NAND2_X1 U13397 ( .A1(n13339), .A2(b_8_), .ZN(n13338) );
  NOR2_X1 U13398 ( .A1(n13340), .A2(n8014), .ZN(n13339) );
  NOR2_X1 U13399 ( .A1(n13146), .A2(n13147), .ZN(n13340) );
  NAND2_X1 U13400 ( .A1(n13146), .A2(n13147), .ZN(n13337) );
  NAND2_X1 U13401 ( .A1(n13341), .A2(n13342), .ZN(n13147) );
  NAND2_X1 U13402 ( .A1(n13343), .A2(a_24_), .ZN(n13342) );
  NOR2_X1 U13403 ( .A1(n13344), .A2(n12909), .ZN(n13343) );
  NOR2_X1 U13404 ( .A1(n13142), .A2(n13143), .ZN(n13344) );
  NAND2_X1 U13405 ( .A1(n13142), .A2(n13143), .ZN(n13341) );
  NAND2_X1 U13406 ( .A1(n13345), .A2(n13346), .ZN(n13143) );
  NAND2_X1 U13407 ( .A1(n13140), .A2(n13347), .ZN(n13346) );
  OR2_X1 U13408 ( .A1(n13138), .A2(n13139), .ZN(n13347) );
  NOR2_X1 U13409 ( .A1(n12909), .A2(n8022), .ZN(n13140) );
  NAND2_X1 U13410 ( .A1(n13138), .A2(n13139), .ZN(n13345) );
  NAND2_X1 U13411 ( .A1(n13135), .A2(n13348), .ZN(n13139) );
  NAND2_X1 U13412 ( .A1(n13134), .A2(n13136), .ZN(n13348) );
  NAND2_X1 U13413 ( .A1(n13349), .A2(n13350), .ZN(n13136) );
  NAND2_X1 U13414 ( .A1(a_26_), .A2(b_8_), .ZN(n13350) );
  INV_X1 U13415 ( .A(n13351), .ZN(n13349) );
  XNOR2_X1 U13416 ( .A(n13352), .B(n13353), .ZN(n13134) );
  NAND2_X1 U13417 ( .A1(n13354), .A2(n13355), .ZN(n13352) );
  NAND2_X1 U13418 ( .A1(a_26_), .A2(n13351), .ZN(n13135) );
  NAND2_X1 U13419 ( .A1(n13104), .A2(n13356), .ZN(n13351) );
  NAND2_X1 U13420 ( .A1(n13103), .A2(n13105), .ZN(n13356) );
  NAND2_X1 U13421 ( .A1(n13357), .A2(n13358), .ZN(n13105) );
  NAND2_X1 U13422 ( .A1(a_27_), .A2(b_8_), .ZN(n13358) );
  INV_X1 U13423 ( .A(n13359), .ZN(n13357) );
  XNOR2_X1 U13424 ( .A(n13360), .B(n13361), .ZN(n13103) );
  XOR2_X1 U13425 ( .A(n13362), .B(n13363), .Z(n13361) );
  NAND2_X1 U13426 ( .A1(b_7_), .A2(a_28_), .ZN(n13363) );
  NAND2_X1 U13427 ( .A1(a_27_), .A2(n13359), .ZN(n13104) );
  NAND2_X1 U13428 ( .A1(n13364), .A2(n13365), .ZN(n13359) );
  NAND2_X1 U13429 ( .A1(n13366), .A2(a_28_), .ZN(n13365) );
  NOR2_X1 U13430 ( .A1(n13367), .A2(n12909), .ZN(n13366) );
  NOR2_X1 U13431 ( .A1(n13110), .A2(n13112), .ZN(n13367) );
  NAND2_X1 U13432 ( .A1(n13110), .A2(n13112), .ZN(n13364) );
  NAND2_X1 U13433 ( .A1(n13368), .A2(n13369), .ZN(n13112) );
  NAND2_X1 U13434 ( .A1(n13130), .A2(n13370), .ZN(n13369) );
  NAND2_X1 U13435 ( .A1(n13132), .A2(n13131), .ZN(n13370) );
  NOR2_X1 U13436 ( .A1(n12909), .A2(n7337), .ZN(n13130) );
  OR2_X1 U13437 ( .A1(n13131), .A2(n13132), .ZN(n13368) );
  AND2_X1 U13438 ( .A1(n13371), .A2(n13372), .ZN(n13132) );
  NAND2_X1 U13439 ( .A1(n13373), .A2(b_6_), .ZN(n13372) );
  NOR2_X1 U13440 ( .A1(n13374), .A2(n7817), .ZN(n13373) );
  NOR2_X1 U13441 ( .A1(n7816), .A2(n13127), .ZN(n13374) );
  NAND2_X1 U13442 ( .A1(n13375), .A2(b_7_), .ZN(n13371) );
  NOR2_X1 U13443 ( .A1(n13376), .A2(n8052), .ZN(n13375) );
  NOR2_X1 U13444 ( .A1(n7810), .A2(n13377), .ZN(n13376) );
  NAND2_X1 U13445 ( .A1(n13378), .A2(b_7_), .ZN(n13131) );
  NOR2_X1 U13446 ( .A1(n8055), .A2(n12909), .ZN(n13378) );
  XOR2_X1 U13447 ( .A(n13379), .B(n13380), .Z(n13110) );
  XOR2_X1 U13448 ( .A(n13381), .B(n13382), .Z(n13379) );
  XNOR2_X1 U13449 ( .A(n13383), .B(n13384), .ZN(n13138) );
  NAND2_X1 U13450 ( .A1(n13385), .A2(n13386), .ZN(n13383) );
  XOR2_X1 U13451 ( .A(n13387), .B(n13388), .Z(n13142) );
  XOR2_X1 U13452 ( .A(n13389), .B(n13390), .Z(n13387) );
  XOR2_X1 U13453 ( .A(n13391), .B(n13392), .Z(n13146) );
  XOR2_X1 U13454 ( .A(n13393), .B(n13394), .Z(n13391) );
  XNOR2_X1 U13455 ( .A(n13395), .B(n13396), .ZN(n13150) );
  XOR2_X1 U13456 ( .A(n13397), .B(n13398), .Z(n13395) );
  NOR2_X1 U13457 ( .A1(n8014), .A2(n13127), .ZN(n13398) );
  XOR2_X1 U13458 ( .A(n13399), .B(n13400), .Z(n13154) );
  NAND2_X1 U13459 ( .A1(n13401), .A2(n13402), .ZN(n13399) );
  XNOR2_X1 U13460 ( .A(n13403), .B(n13404), .ZN(n13158) );
  XOR2_X1 U13461 ( .A(n13405), .B(n13406), .Z(n13403) );
  NOR2_X1 U13462 ( .A1(n7760), .A2(n13127), .ZN(n13406) );
  XNOR2_X1 U13463 ( .A(n13407), .B(n13408), .ZN(n13162) );
  XOR2_X1 U13464 ( .A(n13409), .B(n13410), .Z(n13408) );
  NAND2_X1 U13465 ( .A1(b_7_), .A2(a_20_), .ZN(n13410) );
  XNOR2_X1 U13466 ( .A(n13411), .B(n13412), .ZN(n13166) );
  XOR2_X1 U13467 ( .A(n13413), .B(n13414), .Z(n13412) );
  NAND2_X1 U13468 ( .A1(a_19_), .A2(b_7_), .ZN(n13414) );
  XOR2_X1 U13469 ( .A(n13415), .B(n13416), .Z(n13177) );
  XOR2_X1 U13470 ( .A(n13417), .B(n13418), .Z(n13415) );
  NOR2_X1 U13471 ( .A1(n13127), .A2(n7736), .ZN(n13418) );
  XOR2_X1 U13472 ( .A(n13419), .B(n13420), .Z(n13181) );
  XOR2_X1 U13473 ( .A(n13421), .B(n13422), .Z(n13419) );
  NOR2_X1 U13474 ( .A1(n13127), .A2(n7406), .ZN(n13422) );
  XNOR2_X1 U13475 ( .A(n13423), .B(n13424), .ZN(n13186) );
  XOR2_X1 U13476 ( .A(n13425), .B(n13426), .Z(n13423) );
  NOR2_X1 U13477 ( .A1(n13127), .A2(n7727), .ZN(n13426) );
  XOR2_X1 U13478 ( .A(n13427), .B(n13428), .Z(n13189) );
  XOR2_X1 U13479 ( .A(n13429), .B(n13430), .Z(n13427) );
  NOR2_X1 U13480 ( .A1(n13127), .A2(n7415), .ZN(n13430) );
  XNOR2_X1 U13481 ( .A(n13431), .B(n13432), .ZN(n13194) );
  XOR2_X1 U13482 ( .A(n13433), .B(n13434), .Z(n13431) );
  NOR2_X1 U13483 ( .A1(n13127), .A2(n7718), .ZN(n13434) );
  XOR2_X1 U13484 ( .A(n13435), .B(n13436), .Z(n13033) );
  XOR2_X1 U13485 ( .A(n13437), .B(n13438), .Z(n13435) );
  NOR2_X1 U13486 ( .A1(n7424), .A2(n13127), .ZN(n13438) );
  XOR2_X1 U13487 ( .A(n13439), .B(n13440), .Z(n13197) );
  XOR2_X1 U13488 ( .A(n13441), .B(n13442), .Z(n13439) );
  NOR2_X1 U13489 ( .A1(n13127), .A2(n7709), .ZN(n13442) );
  XNOR2_X1 U13490 ( .A(n13443), .B(n13444), .ZN(n13205) );
  XOR2_X1 U13491 ( .A(n13445), .B(n13446), .Z(n13443) );
  NOR2_X1 U13492 ( .A1(n13127), .A2(n7699), .ZN(n13446) );
  XOR2_X1 U13493 ( .A(n13447), .B(n13448), .Z(n13209) );
  XOR2_X1 U13494 ( .A(n13449), .B(n13450), .Z(n13447) );
  XOR2_X1 U13495 ( .A(n13451), .B(n13452), .Z(n13214) );
  XNOR2_X1 U13496 ( .A(n13453), .B(n13454), .ZN(n13451) );
  NAND2_X1 U13497 ( .A1(a_6_), .A2(b_7_), .ZN(n13453) );
  XOR2_X1 U13498 ( .A(n13455), .B(n13456), .Z(n13217) );
  XOR2_X1 U13499 ( .A(n13457), .B(n13458), .Z(n13455) );
  NOR2_X1 U13500 ( .A1(n13127), .A2(n7455), .ZN(n13458) );
  XOR2_X1 U13501 ( .A(n13459), .B(n13460), .Z(n13222) );
  XOR2_X1 U13502 ( .A(n13461), .B(n13462), .Z(n13459) );
  NOR2_X1 U13503 ( .A1(n13127), .A2(n7682), .ZN(n13462) );
  XOR2_X1 U13504 ( .A(n13463), .B(n13464), .Z(n13226) );
  XOR2_X1 U13505 ( .A(n13465), .B(n13466), .Z(n13463) );
  NOR2_X1 U13506 ( .A1(n13127), .A2(n7464), .ZN(n13466) );
  XOR2_X1 U13507 ( .A(n13467), .B(n13468), .Z(n13230) );
  XOR2_X1 U13508 ( .A(n13469), .B(n13470), .Z(n13467) );
  NOR2_X1 U13509 ( .A1(n13127), .A2(n7469), .ZN(n13470) );
  XNOR2_X1 U13510 ( .A(n13471), .B(n13472), .ZN(n13234) );
  XOR2_X1 U13511 ( .A(n13473), .B(n13474), .Z(n13472) );
  NAND2_X1 U13512 ( .A1(a_1_), .A2(b_7_), .ZN(n13474) );
  XOR2_X1 U13513 ( .A(n13475), .B(n13476), .Z(n12993) );
  XNOR2_X1 U13514 ( .A(n13477), .B(n13478), .ZN(n13476) );
  NAND2_X1 U13515 ( .A1(n13479), .A2(n13239), .ZN(n7323) );
  OR2_X1 U13516 ( .A1(n13239), .A2(n13479), .ZN(n7324) );
  XNOR2_X1 U13517 ( .A(n13480), .B(n13481), .ZN(n13479) );
  NAND2_X1 U13518 ( .A1(n13482), .A2(n13245), .ZN(n13239) );
  NAND2_X1 U13519 ( .A1(n13483), .A2(n13484), .ZN(n13245) );
  NAND2_X1 U13520 ( .A1(n13478), .A2(n13485), .ZN(n13484) );
  OR2_X1 U13521 ( .A1(n13475), .A2(n13477), .ZN(n13485) );
  NOR2_X1 U13522 ( .A1(n13127), .A2(n7478), .ZN(n13478) );
  NAND2_X1 U13523 ( .A1(n13475), .A2(n13477), .ZN(n13483) );
  NAND2_X1 U13524 ( .A1(n13486), .A2(n13487), .ZN(n13477) );
  NAND2_X1 U13525 ( .A1(n13488), .A2(a_1_), .ZN(n13487) );
  NOR2_X1 U13526 ( .A1(n13489), .A2(n13127), .ZN(n13488) );
  NOR2_X1 U13527 ( .A1(n13473), .A2(n13471), .ZN(n13489) );
  NAND2_X1 U13528 ( .A1(n13471), .A2(n13473), .ZN(n13486) );
  NAND2_X1 U13529 ( .A1(n13490), .A2(n13491), .ZN(n13473) );
  NAND2_X1 U13530 ( .A1(n13492), .A2(a_2_), .ZN(n13491) );
  NOR2_X1 U13531 ( .A1(n13493), .A2(n13127), .ZN(n13492) );
  NOR2_X1 U13532 ( .A1(n13469), .A2(n13468), .ZN(n13493) );
  NAND2_X1 U13533 ( .A1(n13468), .A2(n13469), .ZN(n13490) );
  NAND2_X1 U13534 ( .A1(n13494), .A2(n13495), .ZN(n13469) );
  NAND2_X1 U13535 ( .A1(n13496), .A2(a_3_), .ZN(n13495) );
  NOR2_X1 U13536 ( .A1(n13497), .A2(n13127), .ZN(n13496) );
  NOR2_X1 U13537 ( .A1(n13465), .A2(n13464), .ZN(n13497) );
  NAND2_X1 U13538 ( .A1(n13464), .A2(n13465), .ZN(n13494) );
  NAND2_X1 U13539 ( .A1(n13498), .A2(n13499), .ZN(n13465) );
  NAND2_X1 U13540 ( .A1(n13500), .A2(a_4_), .ZN(n13499) );
  NOR2_X1 U13541 ( .A1(n13501), .A2(n13127), .ZN(n13500) );
  NOR2_X1 U13542 ( .A1(n13461), .A2(n13460), .ZN(n13501) );
  NAND2_X1 U13543 ( .A1(n13460), .A2(n13461), .ZN(n13498) );
  NAND2_X1 U13544 ( .A1(n13502), .A2(n13503), .ZN(n13461) );
  NAND2_X1 U13545 ( .A1(n13504), .A2(a_5_), .ZN(n13503) );
  NOR2_X1 U13546 ( .A1(n13505), .A2(n13127), .ZN(n13504) );
  NOR2_X1 U13547 ( .A1(n13457), .A2(n13456), .ZN(n13505) );
  NAND2_X1 U13548 ( .A1(n13456), .A2(n13457), .ZN(n13502) );
  NAND2_X1 U13549 ( .A1(n13506), .A2(n13507), .ZN(n13457) );
  NAND2_X1 U13550 ( .A1(n13508), .A2(a_6_), .ZN(n13507) );
  NOR2_X1 U13551 ( .A1(n13509), .A2(n13127), .ZN(n13508) );
  NOR2_X1 U13552 ( .A1(n13454), .A2(n13452), .ZN(n13509) );
  NAND2_X1 U13553 ( .A1(n13452), .A2(n13454), .ZN(n13506) );
  NAND2_X1 U13554 ( .A1(n13510), .A2(n13511), .ZN(n13454) );
  NAND2_X1 U13555 ( .A1(n13448), .A2(n13512), .ZN(n13511) );
  OR2_X1 U13556 ( .A1(n13449), .A2(n13450), .ZN(n13512) );
  XOR2_X1 U13557 ( .A(n13513), .B(n13514), .Z(n13448) );
  XOR2_X1 U13558 ( .A(n13515), .B(n13516), .Z(n13513) );
  NOR2_X1 U13559 ( .A1(n13377), .A2(n7699), .ZN(n13516) );
  NAND2_X1 U13560 ( .A1(n13450), .A2(n13449), .ZN(n13510) );
  NAND2_X1 U13561 ( .A1(n13517), .A2(n13518), .ZN(n13449) );
  NAND2_X1 U13562 ( .A1(n13519), .A2(a_8_), .ZN(n13518) );
  NOR2_X1 U13563 ( .A1(n13520), .A2(n13127), .ZN(n13519) );
  NOR2_X1 U13564 ( .A1(n13445), .A2(n13444), .ZN(n13520) );
  NAND2_X1 U13565 ( .A1(n13444), .A2(n13445), .ZN(n13517) );
  NAND2_X1 U13566 ( .A1(n13521), .A2(n13522), .ZN(n13445) );
  NAND2_X1 U13567 ( .A1(n13523), .A2(a_9_), .ZN(n13522) );
  NOR2_X1 U13568 ( .A1(n13524), .A2(n13127), .ZN(n13523) );
  NOR2_X1 U13569 ( .A1(n13281), .A2(n13280), .ZN(n13524) );
  NAND2_X1 U13570 ( .A1(n13280), .A2(n13281), .ZN(n13521) );
  NAND2_X1 U13571 ( .A1(n13525), .A2(n13526), .ZN(n13281) );
  NAND2_X1 U13572 ( .A1(n13527), .A2(a_10_), .ZN(n13526) );
  NOR2_X1 U13573 ( .A1(n13528), .A2(n13127), .ZN(n13527) );
  NOR2_X1 U13574 ( .A1(n13441), .A2(n13440), .ZN(n13528) );
  NAND2_X1 U13575 ( .A1(n13440), .A2(n13441), .ZN(n13525) );
  NAND2_X1 U13576 ( .A1(n13529), .A2(n13530), .ZN(n13441) );
  NAND2_X1 U13577 ( .A1(n13531), .A2(b_7_), .ZN(n13530) );
  NOR2_X1 U13578 ( .A1(n13532), .A2(n7424), .ZN(n13531) );
  NOR2_X1 U13579 ( .A1(n13437), .A2(n13436), .ZN(n13532) );
  NAND2_X1 U13580 ( .A1(n13436), .A2(n13437), .ZN(n13529) );
  NAND2_X1 U13581 ( .A1(n13533), .A2(n13534), .ZN(n13437) );
  NAND2_X1 U13582 ( .A1(n13535), .A2(a_12_), .ZN(n13534) );
  NOR2_X1 U13583 ( .A1(n13536), .A2(n13127), .ZN(n13535) );
  NOR2_X1 U13584 ( .A1(n13433), .A2(n13432), .ZN(n13536) );
  NAND2_X1 U13585 ( .A1(n13432), .A2(n13433), .ZN(n13533) );
  NAND2_X1 U13586 ( .A1(n13537), .A2(n13538), .ZN(n13433) );
  NAND2_X1 U13587 ( .A1(n13539), .A2(a_13_), .ZN(n13538) );
  NOR2_X1 U13588 ( .A1(n13540), .A2(n13127), .ZN(n13539) );
  NOR2_X1 U13589 ( .A1(n13428), .A2(n13429), .ZN(n13540) );
  NAND2_X1 U13590 ( .A1(n13428), .A2(n13429), .ZN(n13537) );
  NAND2_X1 U13591 ( .A1(n13541), .A2(n13542), .ZN(n13429) );
  NAND2_X1 U13592 ( .A1(n13543), .A2(a_14_), .ZN(n13542) );
  NOR2_X1 U13593 ( .A1(n13544), .A2(n13127), .ZN(n13543) );
  NOR2_X1 U13594 ( .A1(n13425), .A2(n13424), .ZN(n13544) );
  NAND2_X1 U13595 ( .A1(n13424), .A2(n13425), .ZN(n13541) );
  NAND2_X1 U13596 ( .A1(n13545), .A2(n13546), .ZN(n13425) );
  NAND2_X1 U13597 ( .A1(n13547), .A2(a_15_), .ZN(n13546) );
  NOR2_X1 U13598 ( .A1(n13548), .A2(n13127), .ZN(n13547) );
  NOR2_X1 U13599 ( .A1(n13420), .A2(n13421), .ZN(n13548) );
  NAND2_X1 U13600 ( .A1(n13420), .A2(n13421), .ZN(n13545) );
  NAND2_X1 U13601 ( .A1(n13549), .A2(n13550), .ZN(n13421) );
  NAND2_X1 U13602 ( .A1(n13551), .A2(a_16_), .ZN(n13550) );
  NOR2_X1 U13603 ( .A1(n13552), .A2(n13127), .ZN(n13551) );
  NOR2_X1 U13604 ( .A1(n13417), .A2(n13416), .ZN(n13552) );
  NAND2_X1 U13605 ( .A1(n13416), .A2(n13417), .ZN(n13549) );
  NAND2_X1 U13606 ( .A1(n13553), .A2(n13554), .ZN(n13417) );
  NAND2_X1 U13607 ( .A1(n13555), .A2(a_17_), .ZN(n13554) );
  NOR2_X1 U13608 ( .A1(n13556), .A2(n13127), .ZN(n13555) );
  NOR2_X1 U13609 ( .A1(n13309), .A2(n13311), .ZN(n13556) );
  NAND2_X1 U13610 ( .A1(n13309), .A2(n13311), .ZN(n13553) );
  NAND2_X1 U13611 ( .A1(n13557), .A2(n13558), .ZN(n13311) );
  NAND2_X1 U13612 ( .A1(n13559), .A2(a_18_), .ZN(n13558) );
  NOR2_X1 U13613 ( .A1(n13560), .A2(n13127), .ZN(n13559) );
  NOR2_X1 U13614 ( .A1(n13319), .A2(n13317), .ZN(n13560) );
  NAND2_X1 U13615 ( .A1(n13317), .A2(n13319), .ZN(n13557) );
  NAND2_X1 U13616 ( .A1(n13561), .A2(n13562), .ZN(n13319) );
  NAND2_X1 U13617 ( .A1(n13563), .A2(a_19_), .ZN(n13562) );
  NOR2_X1 U13618 ( .A1(n13564), .A2(n13127), .ZN(n13563) );
  NOR2_X1 U13619 ( .A1(n13411), .A2(n13413), .ZN(n13564) );
  NAND2_X1 U13620 ( .A1(n13411), .A2(n13413), .ZN(n13561) );
  NAND2_X1 U13621 ( .A1(n13565), .A2(n13566), .ZN(n13413) );
  NAND2_X1 U13622 ( .A1(n13567), .A2(b_7_), .ZN(n13566) );
  NOR2_X1 U13623 ( .A1(n13568), .A2(n7755), .ZN(n13567) );
  NOR2_X1 U13624 ( .A1(n13407), .A2(n13409), .ZN(n13568) );
  NAND2_X1 U13625 ( .A1(n13407), .A2(n13409), .ZN(n13565) );
  NAND2_X1 U13626 ( .A1(n13569), .A2(n13570), .ZN(n13409) );
  NAND2_X1 U13627 ( .A1(n13571), .A2(b_7_), .ZN(n13570) );
  NOR2_X1 U13628 ( .A1(n13572), .A2(n7760), .ZN(n13571) );
  NOR2_X1 U13629 ( .A1(n13405), .A2(n13404), .ZN(n13572) );
  NAND2_X1 U13630 ( .A1(n13404), .A2(n13405), .ZN(n13569) );
  NAND2_X1 U13631 ( .A1(n13401), .A2(n13573), .ZN(n13405) );
  NAND2_X1 U13632 ( .A1(n13400), .A2(n13402), .ZN(n13573) );
  NAND2_X1 U13633 ( .A1(n13574), .A2(n13575), .ZN(n13402) );
  NAND2_X1 U13634 ( .A1(a_22_), .A2(b_7_), .ZN(n13575) );
  INV_X1 U13635 ( .A(n13576), .ZN(n13574) );
  XOR2_X1 U13636 ( .A(n13577), .B(n13578), .Z(n13400) );
  XOR2_X1 U13637 ( .A(n13579), .B(n13580), .Z(n13577) );
  NOR2_X1 U13638 ( .A1(n8014), .A2(n13377), .ZN(n13580) );
  NAND2_X1 U13639 ( .A1(a_22_), .A2(n13576), .ZN(n13401) );
  NAND2_X1 U13640 ( .A1(n13581), .A2(n13582), .ZN(n13576) );
  NAND2_X1 U13641 ( .A1(n13583), .A2(b_7_), .ZN(n13582) );
  NOR2_X1 U13642 ( .A1(n13584), .A2(n8014), .ZN(n13583) );
  NOR2_X1 U13643 ( .A1(n13397), .A2(n13396), .ZN(n13584) );
  NAND2_X1 U13644 ( .A1(n13396), .A2(n13397), .ZN(n13581) );
  NAND2_X1 U13645 ( .A1(n13585), .A2(n13586), .ZN(n13397) );
  NAND2_X1 U13646 ( .A1(n13394), .A2(n13587), .ZN(n13586) );
  OR2_X1 U13647 ( .A1(n13392), .A2(n13393), .ZN(n13587) );
  NOR2_X1 U13648 ( .A1(n7774), .A2(n13127), .ZN(n13394) );
  NAND2_X1 U13649 ( .A1(n13392), .A2(n13393), .ZN(n13585) );
  NAND2_X1 U13650 ( .A1(n13588), .A2(n13589), .ZN(n13393) );
  NAND2_X1 U13651 ( .A1(n13390), .A2(n13590), .ZN(n13589) );
  OR2_X1 U13652 ( .A1(n13388), .A2(n13389), .ZN(n13590) );
  NOR2_X1 U13653 ( .A1(n13127), .A2(n8022), .ZN(n13390) );
  NAND2_X1 U13654 ( .A1(n13388), .A2(n13389), .ZN(n13588) );
  NAND2_X1 U13655 ( .A1(n13385), .A2(n13591), .ZN(n13389) );
  NAND2_X1 U13656 ( .A1(n13384), .A2(n13386), .ZN(n13591) );
  NAND2_X1 U13657 ( .A1(n13592), .A2(n13593), .ZN(n13386) );
  NAND2_X1 U13658 ( .A1(a_26_), .A2(b_7_), .ZN(n13593) );
  INV_X1 U13659 ( .A(n13594), .ZN(n13592) );
  XNOR2_X1 U13660 ( .A(n13595), .B(n13596), .ZN(n13384) );
  NAND2_X1 U13661 ( .A1(n13597), .A2(n13598), .ZN(n13595) );
  NAND2_X1 U13662 ( .A1(a_26_), .A2(n13594), .ZN(n13385) );
  NAND2_X1 U13663 ( .A1(n13354), .A2(n13599), .ZN(n13594) );
  NAND2_X1 U13664 ( .A1(n13353), .A2(n13355), .ZN(n13599) );
  NAND2_X1 U13665 ( .A1(n13600), .A2(n13601), .ZN(n13355) );
  NAND2_X1 U13666 ( .A1(b_7_), .A2(a_27_), .ZN(n13601) );
  INV_X1 U13667 ( .A(n13602), .ZN(n13600) );
  XNOR2_X1 U13668 ( .A(n13603), .B(n13604), .ZN(n13353) );
  XOR2_X1 U13669 ( .A(n13605), .B(n13606), .Z(n13604) );
  NAND2_X1 U13670 ( .A1(b_6_), .A2(a_28_), .ZN(n13606) );
  NAND2_X1 U13671 ( .A1(a_27_), .A2(n13602), .ZN(n13354) );
  NAND2_X1 U13672 ( .A1(n13607), .A2(n13608), .ZN(n13602) );
  NAND2_X1 U13673 ( .A1(n13609), .A2(b_7_), .ZN(n13608) );
  NOR2_X1 U13674 ( .A1(n13610), .A2(n7803), .ZN(n13609) );
  NOR2_X1 U13675 ( .A1(n13360), .A2(n13362), .ZN(n13610) );
  NAND2_X1 U13676 ( .A1(n13360), .A2(n13362), .ZN(n13607) );
  NAND2_X1 U13677 ( .A1(n13611), .A2(n13612), .ZN(n13362) );
  NAND2_X1 U13678 ( .A1(n13380), .A2(n13613), .ZN(n13612) );
  NAND2_X1 U13679 ( .A1(n13382), .A2(n13381), .ZN(n13613) );
  NOR2_X1 U13680 ( .A1(n13127), .A2(n7337), .ZN(n13380) );
  OR2_X1 U13681 ( .A1(n13381), .A2(n13382), .ZN(n13611) );
  AND2_X1 U13682 ( .A1(n13614), .A2(n13615), .ZN(n13382) );
  NAND2_X1 U13683 ( .A1(n13616), .A2(b_5_), .ZN(n13615) );
  NOR2_X1 U13684 ( .A1(n13617), .A2(n7817), .ZN(n13616) );
  NOR2_X1 U13685 ( .A1(n7816), .A2(n13377), .ZN(n13617) );
  NAND2_X1 U13686 ( .A1(n13618), .A2(b_6_), .ZN(n13614) );
  NOR2_X1 U13687 ( .A1(n13619), .A2(n8052), .ZN(n13618) );
  NOR2_X1 U13688 ( .A1(n7810), .A2(n13620), .ZN(n13619) );
  NAND2_X1 U13689 ( .A1(n13621), .A2(b_6_), .ZN(n13381) );
  NOR2_X1 U13690 ( .A1(n8055), .A2(n13127), .ZN(n13621) );
  XOR2_X1 U13691 ( .A(n13622), .B(n13623), .Z(n13360) );
  XOR2_X1 U13692 ( .A(n13624), .B(n13625), .Z(n13622) );
  XNOR2_X1 U13693 ( .A(n13626), .B(n13627), .ZN(n13388) );
  NAND2_X1 U13694 ( .A1(n13628), .A2(n13629), .ZN(n13626) );
  XNOR2_X1 U13695 ( .A(n13630), .B(n13631), .ZN(n13392) );
  NAND2_X1 U13696 ( .A1(n13632), .A2(n13633), .ZN(n13630) );
  XNOR2_X1 U13697 ( .A(n13634), .B(n13635), .ZN(n13396) );
  XNOR2_X1 U13698 ( .A(n13636), .B(n13637), .ZN(n13635) );
  XNOR2_X1 U13699 ( .A(n13638), .B(n13639), .ZN(n13404) );
  NAND2_X1 U13700 ( .A1(n13640), .A2(n13641), .ZN(n13638) );
  XNOR2_X1 U13701 ( .A(n13642), .B(n13643), .ZN(n13407) );
  XNOR2_X1 U13702 ( .A(n13644), .B(n13645), .ZN(n13643) );
  XNOR2_X1 U13703 ( .A(n13646), .B(n13647), .ZN(n13411) );
  XOR2_X1 U13704 ( .A(n13648), .B(n13649), .Z(n13647) );
  NAND2_X1 U13705 ( .A1(b_6_), .A2(a_20_), .ZN(n13649) );
  XNOR2_X1 U13706 ( .A(n13650), .B(n13651), .ZN(n13317) );
  XNOR2_X1 U13707 ( .A(n13652), .B(n13653), .ZN(n13650) );
  XOR2_X1 U13708 ( .A(n13654), .B(n13655), .Z(n13309) );
  XOR2_X1 U13709 ( .A(n13656), .B(n13657), .Z(n13654) );
  XNOR2_X1 U13710 ( .A(n13658), .B(n13659), .ZN(n13416) );
  XNOR2_X1 U13711 ( .A(n13660), .B(n13661), .ZN(n13658) );
  XNOR2_X1 U13712 ( .A(n13662), .B(n13663), .ZN(n13420) );
  XNOR2_X1 U13713 ( .A(n13664), .B(n13665), .ZN(n13663) );
  XNOR2_X1 U13714 ( .A(n13666), .B(n13667), .ZN(n13424) );
  XNOR2_X1 U13715 ( .A(n13668), .B(n13669), .ZN(n13667) );
  XNOR2_X1 U13716 ( .A(n13670), .B(n13671), .ZN(n13428) );
  XNOR2_X1 U13717 ( .A(n13672), .B(n13673), .ZN(n13671) );
  XNOR2_X1 U13718 ( .A(n13674), .B(n13675), .ZN(n13432) );
  XNOR2_X1 U13719 ( .A(n13676), .B(n13677), .ZN(n13675) );
  XNOR2_X1 U13720 ( .A(n13678), .B(n13679), .ZN(n13436) );
  XNOR2_X1 U13721 ( .A(n13680), .B(n13681), .ZN(n13679) );
  XNOR2_X1 U13722 ( .A(n13682), .B(n13683), .ZN(n13440) );
  XNOR2_X1 U13723 ( .A(n13684), .B(n13685), .ZN(n13683) );
  XNOR2_X1 U13724 ( .A(n13686), .B(n13687), .ZN(n13280) );
  XNOR2_X1 U13725 ( .A(n13688), .B(n13689), .ZN(n13687) );
  XNOR2_X1 U13726 ( .A(n13690), .B(n13691), .ZN(n13444) );
  XOR2_X1 U13727 ( .A(n13692), .B(n13693), .Z(n13691) );
  NAND2_X1 U13728 ( .A1(a_9_), .A2(b_6_), .ZN(n13693) );
  XOR2_X1 U13729 ( .A(n13694), .B(n13695), .Z(n13452) );
  XOR2_X1 U13730 ( .A(n13696), .B(n13697), .Z(n13694) );
  NOR2_X1 U13731 ( .A1(n13377), .A2(n7445), .ZN(n13697) );
  XNOR2_X1 U13732 ( .A(n13698), .B(n13699), .ZN(n13456) );
  XNOR2_X1 U13733 ( .A(n13700), .B(n13701), .ZN(n13698) );
  XNOR2_X1 U13734 ( .A(n13702), .B(n13703), .ZN(n13460) );
  XOR2_X1 U13735 ( .A(n13704), .B(n13705), .Z(n13703) );
  NAND2_X1 U13736 ( .A1(a_5_), .A2(b_6_), .ZN(n13705) );
  XOR2_X1 U13737 ( .A(n13706), .B(n13707), .Z(n13464) );
  XOR2_X1 U13738 ( .A(n13708), .B(n13709), .Z(n13706) );
  NOR2_X1 U13739 ( .A1(n13377), .A2(n7682), .ZN(n13709) );
  XOR2_X1 U13740 ( .A(n13710), .B(n13711), .Z(n13468) );
  XOR2_X1 U13741 ( .A(n13712), .B(n13713), .Z(n13710) );
  NOR2_X1 U13742 ( .A1(n13377), .A2(n7464), .ZN(n13713) );
  XNOR2_X1 U13743 ( .A(n13714), .B(n13715), .ZN(n13471) );
  XOR2_X1 U13744 ( .A(n13716), .B(n13717), .Z(n13715) );
  NAND2_X1 U13745 ( .A1(a_2_), .A2(b_6_), .ZN(n13717) );
  XOR2_X1 U13746 ( .A(n13718), .B(n13719), .Z(n13475) );
  XOR2_X1 U13747 ( .A(n13720), .B(n13721), .Z(n13718) );
  NOR2_X1 U13748 ( .A1(n13377), .A2(n7669), .ZN(n13721) );
  XNOR2_X1 U13749 ( .A(n13243), .B(n13244), .ZN(n13482) );
  XNOR2_X1 U13750 ( .A(n13722), .B(n13723), .ZN(n13243) );
  NOR2_X1 U13751 ( .A1(n7478), .A2(n13377), .ZN(n13723) );
  NAND2_X1 U13752 ( .A1(n13724), .A2(n13725), .ZN(n7347) );
  OR2_X1 U13753 ( .A1(n13725), .A2(n13724), .ZN(n7346) );
  NAND2_X1 U13754 ( .A1(n13726), .A2(n13727), .ZN(n13724) );
  NAND2_X1 U13755 ( .A1(n13728), .A2(n13729), .ZN(n13727) );
  XOR2_X1 U13756 ( .A(n13730), .B(n13731), .Z(n13729) );
  INV_X1 U13757 ( .A(n13732), .ZN(n13728) );
  NAND2_X1 U13758 ( .A1(n13481), .A2(n13480), .ZN(n13725) );
  NAND2_X1 U13759 ( .A1(n13733), .A2(n13734), .ZN(n13480) );
  NAND2_X1 U13760 ( .A1(n13735), .A2(b_6_), .ZN(n13734) );
  NOR2_X1 U13761 ( .A1(n13736), .A2(n7478), .ZN(n13735) );
  NOR2_X1 U13762 ( .A1(n13722), .A2(n13244), .ZN(n13736) );
  NAND2_X1 U13763 ( .A1(n13244), .A2(n13722), .ZN(n13733) );
  NAND2_X1 U13764 ( .A1(n13737), .A2(n13738), .ZN(n13722) );
  NAND2_X1 U13765 ( .A1(n13739), .A2(a_1_), .ZN(n13738) );
  NOR2_X1 U13766 ( .A1(n13740), .A2(n13377), .ZN(n13739) );
  NOR2_X1 U13767 ( .A1(n13719), .A2(n13720), .ZN(n13740) );
  NAND2_X1 U13768 ( .A1(n13719), .A2(n13720), .ZN(n13737) );
  NAND2_X1 U13769 ( .A1(n13741), .A2(n13742), .ZN(n13720) );
  NAND2_X1 U13770 ( .A1(n13743), .A2(a_2_), .ZN(n13742) );
  NOR2_X1 U13771 ( .A1(n13744), .A2(n13377), .ZN(n13743) );
  NOR2_X1 U13772 ( .A1(n13714), .A2(n13716), .ZN(n13744) );
  NAND2_X1 U13773 ( .A1(n13714), .A2(n13716), .ZN(n13741) );
  NAND2_X1 U13774 ( .A1(n13745), .A2(n13746), .ZN(n13716) );
  NAND2_X1 U13775 ( .A1(n13747), .A2(a_3_), .ZN(n13746) );
  NOR2_X1 U13776 ( .A1(n13748), .A2(n13377), .ZN(n13747) );
  NOR2_X1 U13777 ( .A1(n13711), .A2(n13712), .ZN(n13748) );
  NAND2_X1 U13778 ( .A1(n13711), .A2(n13712), .ZN(n13745) );
  NAND2_X1 U13779 ( .A1(n13749), .A2(n13750), .ZN(n13712) );
  NAND2_X1 U13780 ( .A1(n13751), .A2(a_4_), .ZN(n13750) );
  NOR2_X1 U13781 ( .A1(n13752), .A2(n13377), .ZN(n13751) );
  NOR2_X1 U13782 ( .A1(n13707), .A2(n13708), .ZN(n13752) );
  NAND2_X1 U13783 ( .A1(n13707), .A2(n13708), .ZN(n13749) );
  NAND2_X1 U13784 ( .A1(n13753), .A2(n13754), .ZN(n13708) );
  NAND2_X1 U13785 ( .A1(n13755), .A2(a_5_), .ZN(n13754) );
  NOR2_X1 U13786 ( .A1(n13756), .A2(n13377), .ZN(n13755) );
  NOR2_X1 U13787 ( .A1(n13702), .A2(n13704), .ZN(n13756) );
  NAND2_X1 U13788 ( .A1(n13702), .A2(n13704), .ZN(n13753) );
  NAND2_X1 U13789 ( .A1(n13757), .A2(n13758), .ZN(n13704) );
  NAND2_X1 U13790 ( .A1(n13701), .A2(n13759), .ZN(n13758) );
  NAND2_X1 U13791 ( .A1(n13700), .A2(n13699), .ZN(n13759) );
  OR2_X1 U13792 ( .A1(n13699), .A2(n13700), .ZN(n13757) );
  AND2_X1 U13793 ( .A1(n13760), .A2(n13761), .ZN(n13700) );
  NAND2_X1 U13794 ( .A1(n13762), .A2(a_7_), .ZN(n13761) );
  NOR2_X1 U13795 ( .A1(n13763), .A2(n13377), .ZN(n13762) );
  NOR2_X1 U13796 ( .A1(n13695), .A2(n13696), .ZN(n13763) );
  NAND2_X1 U13797 ( .A1(n13695), .A2(n13696), .ZN(n13760) );
  NAND2_X1 U13798 ( .A1(n13764), .A2(n13765), .ZN(n13696) );
  NAND2_X1 U13799 ( .A1(n13766), .A2(a_8_), .ZN(n13765) );
  NOR2_X1 U13800 ( .A1(n13767), .A2(n13377), .ZN(n13766) );
  NOR2_X1 U13801 ( .A1(n13514), .A2(n13515), .ZN(n13767) );
  NAND2_X1 U13802 ( .A1(n13514), .A2(n13515), .ZN(n13764) );
  NAND2_X1 U13803 ( .A1(n13768), .A2(n13769), .ZN(n13515) );
  NAND2_X1 U13804 ( .A1(n13770), .A2(a_9_), .ZN(n13769) );
  NOR2_X1 U13805 ( .A1(n13771), .A2(n13377), .ZN(n13770) );
  NOR2_X1 U13806 ( .A1(n13690), .A2(n13692), .ZN(n13771) );
  NAND2_X1 U13807 ( .A1(n13690), .A2(n13692), .ZN(n13768) );
  NAND2_X1 U13808 ( .A1(n13772), .A2(n13773), .ZN(n13692) );
  NAND2_X1 U13809 ( .A1(n13689), .A2(n13774), .ZN(n13773) );
  OR2_X1 U13810 ( .A1(n13688), .A2(n13686), .ZN(n13774) );
  NOR2_X1 U13811 ( .A1(n7709), .A2(n13377), .ZN(n13689) );
  NAND2_X1 U13812 ( .A1(n13686), .A2(n13688), .ZN(n13772) );
  NAND2_X1 U13813 ( .A1(n13775), .A2(n13776), .ZN(n13688) );
  NAND2_X1 U13814 ( .A1(n13685), .A2(n13777), .ZN(n13776) );
  OR2_X1 U13815 ( .A1(n13684), .A2(n13682), .ZN(n13777) );
  NOR2_X1 U13816 ( .A1(n13377), .A2(n7424), .ZN(n13685) );
  NAND2_X1 U13817 ( .A1(n13682), .A2(n13684), .ZN(n13775) );
  NAND2_X1 U13818 ( .A1(n13778), .A2(n13779), .ZN(n13684) );
  NAND2_X1 U13819 ( .A1(n13681), .A2(n13780), .ZN(n13779) );
  OR2_X1 U13820 ( .A1(n13680), .A2(n13678), .ZN(n13780) );
  NOR2_X1 U13821 ( .A1(n7718), .A2(n13377), .ZN(n13681) );
  NAND2_X1 U13822 ( .A1(n13678), .A2(n13680), .ZN(n13778) );
  NAND2_X1 U13823 ( .A1(n13781), .A2(n13782), .ZN(n13680) );
  NAND2_X1 U13824 ( .A1(n13677), .A2(n13783), .ZN(n13782) );
  OR2_X1 U13825 ( .A1(n13676), .A2(n13674), .ZN(n13783) );
  NOR2_X1 U13826 ( .A1(n7415), .A2(n13377), .ZN(n13677) );
  NAND2_X1 U13827 ( .A1(n13674), .A2(n13676), .ZN(n13781) );
  NAND2_X1 U13828 ( .A1(n13784), .A2(n13785), .ZN(n13676) );
  NAND2_X1 U13829 ( .A1(n13673), .A2(n13786), .ZN(n13785) );
  OR2_X1 U13830 ( .A1(n13670), .A2(n13672), .ZN(n13786) );
  NOR2_X1 U13831 ( .A1(n7727), .A2(n13377), .ZN(n13673) );
  NAND2_X1 U13832 ( .A1(n13670), .A2(n13672), .ZN(n13784) );
  NAND2_X1 U13833 ( .A1(n13787), .A2(n13788), .ZN(n13672) );
  NAND2_X1 U13834 ( .A1(n13669), .A2(n13789), .ZN(n13788) );
  OR2_X1 U13835 ( .A1(n13668), .A2(n13666), .ZN(n13789) );
  NOR2_X1 U13836 ( .A1(n7406), .A2(n13377), .ZN(n13669) );
  NAND2_X1 U13837 ( .A1(n13666), .A2(n13668), .ZN(n13787) );
  NAND2_X1 U13838 ( .A1(n13790), .A2(n13791), .ZN(n13668) );
  NAND2_X1 U13839 ( .A1(n13665), .A2(n13792), .ZN(n13791) );
  OR2_X1 U13840 ( .A1(n13662), .A2(n13664), .ZN(n13792) );
  NOR2_X1 U13841 ( .A1(n7736), .A2(n13377), .ZN(n13665) );
  NAND2_X1 U13842 ( .A1(n13662), .A2(n13664), .ZN(n13790) );
  NAND2_X1 U13843 ( .A1(n13793), .A2(n13794), .ZN(n13664) );
  NAND2_X1 U13844 ( .A1(n13661), .A2(n13795), .ZN(n13794) );
  NAND2_X1 U13845 ( .A1(n13660), .A2(n13659), .ZN(n13795) );
  NOR2_X1 U13846 ( .A1(n7397), .A2(n13377), .ZN(n13661) );
  OR2_X1 U13847 ( .A1(n13659), .A2(n13660), .ZN(n13793) );
  AND2_X1 U13848 ( .A1(n13796), .A2(n13797), .ZN(n13660) );
  NAND2_X1 U13849 ( .A1(n13657), .A2(n13798), .ZN(n13797) );
  OR2_X1 U13850 ( .A1(n13655), .A2(n13656), .ZN(n13798) );
  NOR2_X1 U13851 ( .A1(n7745), .A2(n13377), .ZN(n13657) );
  NAND2_X1 U13852 ( .A1(n13655), .A2(n13656), .ZN(n13796) );
  NAND2_X1 U13853 ( .A1(n13799), .A2(n13800), .ZN(n13656) );
  NAND2_X1 U13854 ( .A1(n13652), .A2(n13801), .ZN(n13800) );
  NAND2_X1 U13855 ( .A1(n13653), .A2(n13651), .ZN(n13801) );
  NOR2_X1 U13856 ( .A1(n7750), .A2(n13377), .ZN(n13652) );
  OR2_X1 U13857 ( .A1(n13651), .A2(n13653), .ZN(n13799) );
  AND2_X1 U13858 ( .A1(n13802), .A2(n13803), .ZN(n13653) );
  NAND2_X1 U13859 ( .A1(n13804), .A2(b_6_), .ZN(n13803) );
  NOR2_X1 U13860 ( .A1(n13805), .A2(n7755), .ZN(n13804) );
  NOR2_X1 U13861 ( .A1(n13648), .A2(n13646), .ZN(n13805) );
  NAND2_X1 U13862 ( .A1(n13646), .A2(n13648), .ZN(n13802) );
  NAND2_X1 U13863 ( .A1(n13806), .A2(n13807), .ZN(n13648) );
  NAND2_X1 U13864 ( .A1(n13645), .A2(n13808), .ZN(n13807) );
  OR2_X1 U13865 ( .A1(n13642), .A2(n13644), .ZN(n13808) );
  NOR2_X1 U13866 ( .A1(n13377), .A2(n7760), .ZN(n13645) );
  NAND2_X1 U13867 ( .A1(n13642), .A2(n13644), .ZN(n13806) );
  NAND2_X1 U13868 ( .A1(n13640), .A2(n13809), .ZN(n13644) );
  NAND2_X1 U13869 ( .A1(n13639), .A2(n13641), .ZN(n13809) );
  NAND2_X1 U13870 ( .A1(n13810), .A2(n13811), .ZN(n13641) );
  NAND2_X1 U13871 ( .A1(a_22_), .A2(b_6_), .ZN(n13811) );
  INV_X1 U13872 ( .A(n13812), .ZN(n13810) );
  XOR2_X1 U13873 ( .A(n13813), .B(n13814), .Z(n13639) );
  XOR2_X1 U13874 ( .A(n13815), .B(n13816), .Z(n13813) );
  NOR2_X1 U13875 ( .A1(n8014), .A2(n13620), .ZN(n13816) );
  NAND2_X1 U13876 ( .A1(a_22_), .A2(n13812), .ZN(n13640) );
  NAND2_X1 U13877 ( .A1(n13817), .A2(n13818), .ZN(n13812) );
  NAND2_X1 U13878 ( .A1(n13819), .A2(b_6_), .ZN(n13818) );
  NOR2_X1 U13879 ( .A1(n13820), .A2(n8014), .ZN(n13819) );
  NOR2_X1 U13880 ( .A1(n13579), .A2(n13578), .ZN(n13820) );
  NAND2_X1 U13881 ( .A1(n13578), .A2(n13579), .ZN(n13817) );
  NAND2_X1 U13882 ( .A1(n13821), .A2(n13822), .ZN(n13579) );
  NAND2_X1 U13883 ( .A1(n13637), .A2(n13823), .ZN(n13822) );
  OR2_X1 U13884 ( .A1(n13636), .A2(n13634), .ZN(n13823) );
  NOR2_X1 U13885 ( .A1(n7774), .A2(n13377), .ZN(n13637) );
  NAND2_X1 U13886 ( .A1(n13634), .A2(n13636), .ZN(n13821) );
  NAND2_X1 U13887 ( .A1(n13632), .A2(n13824), .ZN(n13636) );
  NAND2_X1 U13888 ( .A1(n13631), .A2(n13633), .ZN(n13824) );
  NAND2_X1 U13889 ( .A1(n13825), .A2(n13826), .ZN(n13633) );
  NAND2_X1 U13890 ( .A1(b_6_), .A2(a_25_), .ZN(n13826) );
  INV_X1 U13891 ( .A(n13827), .ZN(n13825) );
  XNOR2_X1 U13892 ( .A(n13828), .B(n13829), .ZN(n13631) );
  NAND2_X1 U13893 ( .A1(n13830), .A2(n13831), .ZN(n13828) );
  NAND2_X1 U13894 ( .A1(a_25_), .A2(n13827), .ZN(n13632) );
  NAND2_X1 U13895 ( .A1(n13628), .A2(n13832), .ZN(n13827) );
  NAND2_X1 U13896 ( .A1(n13627), .A2(n13629), .ZN(n13832) );
  NAND2_X1 U13897 ( .A1(n13833), .A2(n13834), .ZN(n13629) );
  NAND2_X1 U13898 ( .A1(b_6_), .A2(a_26_), .ZN(n13834) );
  INV_X1 U13899 ( .A(n13835), .ZN(n13833) );
  XNOR2_X1 U13900 ( .A(n13836), .B(n13837), .ZN(n13627) );
  NAND2_X1 U13901 ( .A1(n13838), .A2(n13839), .ZN(n13836) );
  NAND2_X1 U13902 ( .A1(a_26_), .A2(n13835), .ZN(n13628) );
  NAND2_X1 U13903 ( .A1(n13597), .A2(n13840), .ZN(n13835) );
  NAND2_X1 U13904 ( .A1(n13596), .A2(n13598), .ZN(n13840) );
  NAND2_X1 U13905 ( .A1(n13841), .A2(n13842), .ZN(n13598) );
  NAND2_X1 U13906 ( .A1(b_6_), .A2(a_27_), .ZN(n13842) );
  INV_X1 U13907 ( .A(n13843), .ZN(n13841) );
  XNOR2_X1 U13908 ( .A(n13844), .B(n13845), .ZN(n13596) );
  XOR2_X1 U13909 ( .A(n13846), .B(n13847), .Z(n13845) );
  NAND2_X1 U13910 ( .A1(b_5_), .A2(a_28_), .ZN(n13847) );
  NAND2_X1 U13911 ( .A1(a_27_), .A2(n13843), .ZN(n13597) );
  NAND2_X1 U13912 ( .A1(n13848), .A2(n13849), .ZN(n13843) );
  NAND2_X1 U13913 ( .A1(n13850), .A2(b_6_), .ZN(n13849) );
  NOR2_X1 U13914 ( .A1(n13851), .A2(n7803), .ZN(n13850) );
  NOR2_X1 U13915 ( .A1(n13603), .A2(n13605), .ZN(n13851) );
  NAND2_X1 U13916 ( .A1(n13603), .A2(n13605), .ZN(n13848) );
  NAND2_X1 U13917 ( .A1(n13852), .A2(n13853), .ZN(n13605) );
  NAND2_X1 U13918 ( .A1(n13623), .A2(n13854), .ZN(n13853) );
  NAND2_X1 U13919 ( .A1(n13625), .A2(n13624), .ZN(n13854) );
  NOR2_X1 U13920 ( .A1(n13377), .A2(n7337), .ZN(n13623) );
  OR2_X1 U13921 ( .A1(n13624), .A2(n13625), .ZN(n13852) );
  AND2_X1 U13922 ( .A1(n13855), .A2(n13856), .ZN(n13625) );
  NAND2_X1 U13923 ( .A1(n13857), .A2(b_4_), .ZN(n13856) );
  NOR2_X1 U13924 ( .A1(n13858), .A2(n7817), .ZN(n13857) );
  NOR2_X1 U13925 ( .A1(n7816), .A2(n13620), .ZN(n13858) );
  NAND2_X1 U13926 ( .A1(n13859), .A2(b_5_), .ZN(n13855) );
  NOR2_X1 U13927 ( .A1(n13860), .A2(n8052), .ZN(n13859) );
  NOR2_X1 U13928 ( .A1(n7810), .A2(n13861), .ZN(n13860) );
  NAND2_X1 U13929 ( .A1(n13862), .A2(b_5_), .ZN(n13624) );
  NOR2_X1 U13930 ( .A1(n8055), .A2(n13377), .ZN(n13862) );
  XOR2_X1 U13931 ( .A(n13863), .B(n13864), .Z(n13603) );
  XOR2_X1 U13932 ( .A(n13865), .B(n13866), .Z(n13863) );
  XNOR2_X1 U13933 ( .A(n13867), .B(n13868), .ZN(n13634) );
  NAND2_X1 U13934 ( .A1(n13869), .A2(n13870), .ZN(n13867) );
  XNOR2_X1 U13935 ( .A(n13871), .B(n13872), .ZN(n13578) );
  XOR2_X1 U13936 ( .A(n13873), .B(n13874), .Z(n13872) );
  NAND2_X1 U13937 ( .A1(a_24_), .A2(b_5_), .ZN(n13874) );
  XOR2_X1 U13938 ( .A(n13875), .B(n13876), .Z(n13642) );
  XOR2_X1 U13939 ( .A(n13877), .B(n13878), .Z(n13875) );
  NOR2_X1 U13940 ( .A1(n13620), .A2(n7765), .ZN(n13878) );
  XOR2_X1 U13941 ( .A(n13879), .B(n13880), .Z(n13646) );
  XOR2_X1 U13942 ( .A(n13881), .B(n13882), .Z(n13879) );
  NOR2_X1 U13943 ( .A1(n7760), .A2(n13620), .ZN(n13882) );
  XNOR2_X1 U13944 ( .A(n13883), .B(n13884), .ZN(n13651) );
  XOR2_X1 U13945 ( .A(n13885), .B(n13886), .Z(n13883) );
  NOR2_X1 U13946 ( .A1(n7755), .A2(n13620), .ZN(n13886) );
  XOR2_X1 U13947 ( .A(n13887), .B(n13888), .Z(n13655) );
  XOR2_X1 U13948 ( .A(n13889), .B(n13890), .Z(n13887) );
  NOR2_X1 U13949 ( .A1(n13620), .A2(n7750), .ZN(n13890) );
  XNOR2_X1 U13950 ( .A(n13891), .B(n13892), .ZN(n13659) );
  XOR2_X1 U13951 ( .A(n13893), .B(n13894), .Z(n13891) );
  NOR2_X1 U13952 ( .A1(n13620), .A2(n7745), .ZN(n13894) );
  XOR2_X1 U13953 ( .A(n13895), .B(n13896), .Z(n13662) );
  XOR2_X1 U13954 ( .A(n13897), .B(n13898), .Z(n13895) );
  NOR2_X1 U13955 ( .A1(n13620), .A2(n7397), .ZN(n13898) );
  XOR2_X1 U13956 ( .A(n13899), .B(n13900), .Z(n13666) );
  XOR2_X1 U13957 ( .A(n13901), .B(n13902), .Z(n13899) );
  NOR2_X1 U13958 ( .A1(n13620), .A2(n7736), .ZN(n13902) );
  XOR2_X1 U13959 ( .A(n13903), .B(n13904), .Z(n13670) );
  XOR2_X1 U13960 ( .A(n13905), .B(n13906), .Z(n13903) );
  NOR2_X1 U13961 ( .A1(n13620), .A2(n7406), .ZN(n13906) );
  XOR2_X1 U13962 ( .A(n13907), .B(n13908), .Z(n13674) );
  XOR2_X1 U13963 ( .A(n13909), .B(n13910), .Z(n13907) );
  NOR2_X1 U13964 ( .A1(n13620), .A2(n7727), .ZN(n13910) );
  XOR2_X1 U13965 ( .A(n13911), .B(n13912), .Z(n13678) );
  XOR2_X1 U13966 ( .A(n13913), .B(n13914), .Z(n13911) );
  NOR2_X1 U13967 ( .A1(n13620), .A2(n7415), .ZN(n13914) );
  XOR2_X1 U13968 ( .A(n13915), .B(n13916), .Z(n13682) );
  XOR2_X1 U13969 ( .A(n13917), .B(n13918), .Z(n13915) );
  NOR2_X1 U13970 ( .A1(n13620), .A2(n7718), .ZN(n13918) );
  XOR2_X1 U13971 ( .A(n13919), .B(n13920), .Z(n13686) );
  XOR2_X1 U13972 ( .A(n13921), .B(n13922), .Z(n13919) );
  NOR2_X1 U13973 ( .A1(n7424), .A2(n13620), .ZN(n13922) );
  XOR2_X1 U13974 ( .A(n13923), .B(n13924), .Z(n13690) );
  XOR2_X1 U13975 ( .A(n13925), .B(n13926), .Z(n13923) );
  NOR2_X1 U13976 ( .A1(n13620), .A2(n7709), .ZN(n13926) );
  XOR2_X1 U13977 ( .A(n13927), .B(n13928), .Z(n13514) );
  XOR2_X1 U13978 ( .A(n13929), .B(n13930), .Z(n13927) );
  NOR2_X1 U13979 ( .A1(n13620), .A2(n7704), .ZN(n13930) );
  XOR2_X1 U13980 ( .A(n13931), .B(n13932), .Z(n13695) );
  XOR2_X1 U13981 ( .A(n13933), .B(n13934), .Z(n13931) );
  NOR2_X1 U13982 ( .A1(n13620), .A2(n7699), .ZN(n13934) );
  XNOR2_X1 U13983 ( .A(n13935), .B(n13936), .ZN(n13699) );
  XOR2_X1 U13984 ( .A(n13937), .B(n13938), .Z(n13935) );
  NOR2_X1 U13985 ( .A1(n13620), .A2(n7445), .ZN(n13938) );
  XOR2_X1 U13986 ( .A(n13939), .B(n13940), .Z(n13702) );
  XOR2_X1 U13987 ( .A(n13941), .B(n13942), .Z(n13939) );
  NOR2_X1 U13988 ( .A1(n13620), .A2(n7450), .ZN(n13942) );
  XOR2_X1 U13989 ( .A(n13943), .B(n13944), .Z(n13707) );
  XOR2_X1 U13990 ( .A(n13945), .B(n13946), .Z(n13943) );
  XOR2_X1 U13991 ( .A(n13947), .B(n13948), .Z(n13711) );
  XNOR2_X1 U13992 ( .A(n13949), .B(n13950), .ZN(n13947) );
  NAND2_X1 U13993 ( .A1(a_4_), .A2(b_5_), .ZN(n13949) );
  XOR2_X1 U13994 ( .A(n13951), .B(n13952), .Z(n13714) );
  XOR2_X1 U13995 ( .A(n13953), .B(n13954), .Z(n13951) );
  NOR2_X1 U13996 ( .A1(n13620), .A2(n7464), .ZN(n13954) );
  XOR2_X1 U13997 ( .A(n13955), .B(n13956), .Z(n13719) );
  XOR2_X1 U13998 ( .A(n13957), .B(n13958), .Z(n13955) );
  NOR2_X1 U13999 ( .A1(n13620), .A2(n7469), .ZN(n13958) );
  XOR2_X1 U14000 ( .A(n13959), .B(n13960), .Z(n13244) );
  XOR2_X1 U14001 ( .A(n13961), .B(n13962), .Z(n13959) );
  NOR2_X1 U14002 ( .A1(n13620), .A2(n7669), .ZN(n13962) );
  XOR2_X1 U14003 ( .A(n13963), .B(n13964), .Z(n13481) );
  XOR2_X1 U14004 ( .A(n13965), .B(n13966), .Z(n13963) );
  NAND2_X1 U14005 ( .A1(n13967), .A2(n13726), .ZN(n7391) );
  OR2_X1 U14006 ( .A1(n13726), .A2(n13967), .ZN(n7392) );
  XNOR2_X1 U14007 ( .A(n13968), .B(n13969), .ZN(n13967) );
  NAND2_X1 U14008 ( .A1(n13970), .A2(n13732), .ZN(n13726) );
  NAND2_X1 U14009 ( .A1(n13971), .A2(n13972), .ZN(n13732) );
  NAND2_X1 U14010 ( .A1(n13966), .A2(n13973), .ZN(n13972) );
  OR2_X1 U14011 ( .A1(n13964), .A2(n13965), .ZN(n13973) );
  NOR2_X1 U14012 ( .A1(n13620), .A2(n7478), .ZN(n13966) );
  NAND2_X1 U14013 ( .A1(n13964), .A2(n13965), .ZN(n13971) );
  NAND2_X1 U14014 ( .A1(n13974), .A2(n13975), .ZN(n13965) );
  NAND2_X1 U14015 ( .A1(n13976), .A2(a_1_), .ZN(n13975) );
  NOR2_X1 U14016 ( .A1(n13977), .A2(n13620), .ZN(n13976) );
  NOR2_X1 U14017 ( .A1(n13960), .A2(n13961), .ZN(n13977) );
  NAND2_X1 U14018 ( .A1(n13960), .A2(n13961), .ZN(n13974) );
  NAND2_X1 U14019 ( .A1(n13978), .A2(n13979), .ZN(n13961) );
  NAND2_X1 U14020 ( .A1(n13980), .A2(a_2_), .ZN(n13979) );
  NOR2_X1 U14021 ( .A1(n13981), .A2(n13620), .ZN(n13980) );
  NOR2_X1 U14022 ( .A1(n13957), .A2(n13956), .ZN(n13981) );
  NAND2_X1 U14023 ( .A1(n13956), .A2(n13957), .ZN(n13978) );
  NAND2_X1 U14024 ( .A1(n13982), .A2(n13983), .ZN(n13957) );
  NAND2_X1 U14025 ( .A1(n13984), .A2(a_3_), .ZN(n13983) );
  NOR2_X1 U14026 ( .A1(n13985), .A2(n13620), .ZN(n13984) );
  NOR2_X1 U14027 ( .A1(n13953), .A2(n13952), .ZN(n13985) );
  NAND2_X1 U14028 ( .A1(n13952), .A2(n13953), .ZN(n13982) );
  NAND2_X1 U14029 ( .A1(n13986), .A2(n13987), .ZN(n13953) );
  NAND2_X1 U14030 ( .A1(n13988), .A2(a_4_), .ZN(n13987) );
  NOR2_X1 U14031 ( .A1(n13989), .A2(n13620), .ZN(n13988) );
  NOR2_X1 U14032 ( .A1(n13950), .A2(n13948), .ZN(n13989) );
  NAND2_X1 U14033 ( .A1(n13948), .A2(n13950), .ZN(n13986) );
  NAND2_X1 U14034 ( .A1(n13990), .A2(n13991), .ZN(n13950) );
  NAND2_X1 U14035 ( .A1(n13944), .A2(n13992), .ZN(n13991) );
  OR2_X1 U14036 ( .A1(n13945), .A2(n13946), .ZN(n13992) );
  XOR2_X1 U14037 ( .A(n13993), .B(n13994), .Z(n13944) );
  XOR2_X1 U14038 ( .A(n13995), .B(n13996), .Z(n13993) );
  NOR2_X1 U14039 ( .A1(n13861), .A2(n7450), .ZN(n13996) );
  NAND2_X1 U14040 ( .A1(n13946), .A2(n13945), .ZN(n13990) );
  NAND2_X1 U14041 ( .A1(n13997), .A2(n13998), .ZN(n13945) );
  NAND2_X1 U14042 ( .A1(n13999), .A2(a_6_), .ZN(n13998) );
  NOR2_X1 U14043 ( .A1(n14000), .A2(n13620), .ZN(n13999) );
  NOR2_X1 U14044 ( .A1(n13941), .A2(n13940), .ZN(n14000) );
  NAND2_X1 U14045 ( .A1(n13940), .A2(n13941), .ZN(n13997) );
  NAND2_X1 U14046 ( .A1(n14001), .A2(n14002), .ZN(n13941) );
  NAND2_X1 U14047 ( .A1(n14003), .A2(a_7_), .ZN(n14002) );
  NOR2_X1 U14048 ( .A1(n14004), .A2(n13620), .ZN(n14003) );
  NOR2_X1 U14049 ( .A1(n13937), .A2(n13936), .ZN(n14004) );
  NAND2_X1 U14050 ( .A1(n13936), .A2(n13937), .ZN(n14001) );
  NAND2_X1 U14051 ( .A1(n14005), .A2(n14006), .ZN(n13937) );
  NAND2_X1 U14052 ( .A1(n14007), .A2(a_8_), .ZN(n14006) );
  NOR2_X1 U14053 ( .A1(n14008), .A2(n13620), .ZN(n14007) );
  NOR2_X1 U14054 ( .A1(n13933), .A2(n13932), .ZN(n14008) );
  NAND2_X1 U14055 ( .A1(n13932), .A2(n13933), .ZN(n14005) );
  NAND2_X1 U14056 ( .A1(n14009), .A2(n14010), .ZN(n13933) );
  NAND2_X1 U14057 ( .A1(n14011), .A2(a_9_), .ZN(n14010) );
  NOR2_X1 U14058 ( .A1(n14012), .A2(n13620), .ZN(n14011) );
  NOR2_X1 U14059 ( .A1(n13929), .A2(n13928), .ZN(n14012) );
  NAND2_X1 U14060 ( .A1(n13928), .A2(n13929), .ZN(n14009) );
  NAND2_X1 U14061 ( .A1(n14013), .A2(n14014), .ZN(n13929) );
  NAND2_X1 U14062 ( .A1(n14015), .A2(a_10_), .ZN(n14014) );
  NOR2_X1 U14063 ( .A1(n14016), .A2(n13620), .ZN(n14015) );
  NOR2_X1 U14064 ( .A1(n13925), .A2(n13924), .ZN(n14016) );
  NAND2_X1 U14065 ( .A1(n13924), .A2(n13925), .ZN(n14013) );
  NAND2_X1 U14066 ( .A1(n14017), .A2(n14018), .ZN(n13925) );
  NAND2_X1 U14067 ( .A1(n14019), .A2(b_5_), .ZN(n14018) );
  NOR2_X1 U14068 ( .A1(n14020), .A2(n7424), .ZN(n14019) );
  NOR2_X1 U14069 ( .A1(n13921), .A2(n13920), .ZN(n14020) );
  NAND2_X1 U14070 ( .A1(n13920), .A2(n13921), .ZN(n14017) );
  NAND2_X1 U14071 ( .A1(n14021), .A2(n14022), .ZN(n13921) );
  NAND2_X1 U14072 ( .A1(n14023), .A2(a_12_), .ZN(n14022) );
  NOR2_X1 U14073 ( .A1(n14024), .A2(n13620), .ZN(n14023) );
  NOR2_X1 U14074 ( .A1(n13917), .A2(n13916), .ZN(n14024) );
  NAND2_X1 U14075 ( .A1(n13916), .A2(n13917), .ZN(n14021) );
  NAND2_X1 U14076 ( .A1(n14025), .A2(n14026), .ZN(n13917) );
  NAND2_X1 U14077 ( .A1(n14027), .A2(a_13_), .ZN(n14026) );
  NOR2_X1 U14078 ( .A1(n14028), .A2(n13620), .ZN(n14027) );
  NOR2_X1 U14079 ( .A1(n13913), .A2(n13912), .ZN(n14028) );
  NAND2_X1 U14080 ( .A1(n13912), .A2(n13913), .ZN(n14025) );
  NAND2_X1 U14081 ( .A1(n14029), .A2(n14030), .ZN(n13913) );
  NAND2_X1 U14082 ( .A1(n14031), .A2(a_14_), .ZN(n14030) );
  NOR2_X1 U14083 ( .A1(n14032), .A2(n13620), .ZN(n14031) );
  NOR2_X1 U14084 ( .A1(n13909), .A2(n13908), .ZN(n14032) );
  NAND2_X1 U14085 ( .A1(n13908), .A2(n13909), .ZN(n14029) );
  NAND2_X1 U14086 ( .A1(n14033), .A2(n14034), .ZN(n13909) );
  NAND2_X1 U14087 ( .A1(n14035), .A2(a_15_), .ZN(n14034) );
  NOR2_X1 U14088 ( .A1(n14036), .A2(n13620), .ZN(n14035) );
  NOR2_X1 U14089 ( .A1(n13904), .A2(n13905), .ZN(n14036) );
  NAND2_X1 U14090 ( .A1(n13904), .A2(n13905), .ZN(n14033) );
  NAND2_X1 U14091 ( .A1(n14037), .A2(n14038), .ZN(n13905) );
  NAND2_X1 U14092 ( .A1(n14039), .A2(a_16_), .ZN(n14038) );
  NOR2_X1 U14093 ( .A1(n14040), .A2(n13620), .ZN(n14039) );
  NOR2_X1 U14094 ( .A1(n13901), .A2(n13900), .ZN(n14040) );
  NAND2_X1 U14095 ( .A1(n13900), .A2(n13901), .ZN(n14037) );
  NAND2_X1 U14096 ( .A1(n14041), .A2(n14042), .ZN(n13901) );
  NAND2_X1 U14097 ( .A1(n14043), .A2(a_17_), .ZN(n14042) );
  NOR2_X1 U14098 ( .A1(n14044), .A2(n13620), .ZN(n14043) );
  NOR2_X1 U14099 ( .A1(n13896), .A2(n13897), .ZN(n14044) );
  NAND2_X1 U14100 ( .A1(n13896), .A2(n13897), .ZN(n14041) );
  NAND2_X1 U14101 ( .A1(n14045), .A2(n14046), .ZN(n13897) );
  NAND2_X1 U14102 ( .A1(n14047), .A2(a_18_), .ZN(n14046) );
  NOR2_X1 U14103 ( .A1(n14048), .A2(n13620), .ZN(n14047) );
  NOR2_X1 U14104 ( .A1(n13893), .A2(n13892), .ZN(n14048) );
  NAND2_X1 U14105 ( .A1(n13892), .A2(n13893), .ZN(n14045) );
  NAND2_X1 U14106 ( .A1(n14049), .A2(n14050), .ZN(n13893) );
  NAND2_X1 U14107 ( .A1(n14051), .A2(a_19_), .ZN(n14050) );
  NOR2_X1 U14108 ( .A1(n14052), .A2(n13620), .ZN(n14051) );
  NOR2_X1 U14109 ( .A1(n13888), .A2(n13889), .ZN(n14052) );
  NAND2_X1 U14110 ( .A1(n13888), .A2(n13889), .ZN(n14049) );
  NAND2_X1 U14111 ( .A1(n14053), .A2(n14054), .ZN(n13889) );
  NAND2_X1 U14112 ( .A1(n14055), .A2(b_5_), .ZN(n14054) );
  NOR2_X1 U14113 ( .A1(n14056), .A2(n7755), .ZN(n14055) );
  NOR2_X1 U14114 ( .A1(n13885), .A2(n13884), .ZN(n14056) );
  NAND2_X1 U14115 ( .A1(n13884), .A2(n13885), .ZN(n14053) );
  NAND2_X1 U14116 ( .A1(n14057), .A2(n14058), .ZN(n13885) );
  NAND2_X1 U14117 ( .A1(n14059), .A2(b_5_), .ZN(n14058) );
  NOR2_X1 U14118 ( .A1(n14060), .A2(n7760), .ZN(n14059) );
  NOR2_X1 U14119 ( .A1(n13880), .A2(n13881), .ZN(n14060) );
  NAND2_X1 U14120 ( .A1(n13880), .A2(n13881), .ZN(n14057) );
  NAND2_X1 U14121 ( .A1(n14061), .A2(n14062), .ZN(n13881) );
  NAND2_X1 U14122 ( .A1(n14063), .A2(a_22_), .ZN(n14062) );
  NOR2_X1 U14123 ( .A1(n14064), .A2(n13620), .ZN(n14063) );
  NOR2_X1 U14124 ( .A1(n13876), .A2(n13877), .ZN(n14064) );
  NAND2_X1 U14125 ( .A1(n13876), .A2(n13877), .ZN(n14061) );
  NAND2_X1 U14126 ( .A1(n14065), .A2(n14066), .ZN(n13877) );
  NAND2_X1 U14127 ( .A1(n14067), .A2(b_5_), .ZN(n14066) );
  NOR2_X1 U14128 ( .A1(n14068), .A2(n8014), .ZN(n14067) );
  NOR2_X1 U14129 ( .A1(n13814), .A2(n13815), .ZN(n14068) );
  NAND2_X1 U14130 ( .A1(n13814), .A2(n13815), .ZN(n14065) );
  NAND2_X1 U14131 ( .A1(n14069), .A2(n14070), .ZN(n13815) );
  NAND2_X1 U14132 ( .A1(n14071), .A2(a_24_), .ZN(n14070) );
  NOR2_X1 U14133 ( .A1(n14072), .A2(n13620), .ZN(n14071) );
  NOR2_X1 U14134 ( .A1(n13871), .A2(n13873), .ZN(n14072) );
  NAND2_X1 U14135 ( .A1(n13871), .A2(n13873), .ZN(n14069) );
  NAND2_X1 U14136 ( .A1(n13869), .A2(n14073), .ZN(n13873) );
  NAND2_X1 U14137 ( .A1(n13868), .A2(n13870), .ZN(n14073) );
  NAND2_X1 U14138 ( .A1(n14074), .A2(n14075), .ZN(n13870) );
  NAND2_X1 U14139 ( .A1(b_5_), .A2(a_25_), .ZN(n14075) );
  INV_X1 U14140 ( .A(n14076), .ZN(n14074) );
  XNOR2_X1 U14141 ( .A(n14077), .B(n14078), .ZN(n13868) );
  NAND2_X1 U14142 ( .A1(n14079), .A2(n14080), .ZN(n14077) );
  NAND2_X1 U14143 ( .A1(a_25_), .A2(n14076), .ZN(n13869) );
  NAND2_X1 U14144 ( .A1(n13830), .A2(n14081), .ZN(n14076) );
  NAND2_X1 U14145 ( .A1(n13829), .A2(n13831), .ZN(n14081) );
  NAND2_X1 U14146 ( .A1(n14082), .A2(n14083), .ZN(n13831) );
  NAND2_X1 U14147 ( .A1(b_5_), .A2(a_26_), .ZN(n14083) );
  INV_X1 U14148 ( .A(n14084), .ZN(n14082) );
  XNOR2_X1 U14149 ( .A(n14085), .B(n14086), .ZN(n13829) );
  NAND2_X1 U14150 ( .A1(n14087), .A2(n14088), .ZN(n14085) );
  NAND2_X1 U14151 ( .A1(a_26_), .A2(n14084), .ZN(n13830) );
  NAND2_X1 U14152 ( .A1(n13838), .A2(n14089), .ZN(n14084) );
  NAND2_X1 U14153 ( .A1(n13837), .A2(n13839), .ZN(n14089) );
  NAND2_X1 U14154 ( .A1(n14090), .A2(n14091), .ZN(n13839) );
  NAND2_X1 U14155 ( .A1(b_5_), .A2(a_27_), .ZN(n14091) );
  INV_X1 U14156 ( .A(n14092), .ZN(n14090) );
  XNOR2_X1 U14157 ( .A(n14093), .B(n14094), .ZN(n13837) );
  XOR2_X1 U14158 ( .A(n14095), .B(n14096), .Z(n14094) );
  NAND2_X1 U14159 ( .A1(b_4_), .A2(a_28_), .ZN(n14096) );
  NAND2_X1 U14160 ( .A1(a_27_), .A2(n14092), .ZN(n13838) );
  NAND2_X1 U14161 ( .A1(n14097), .A2(n14098), .ZN(n14092) );
  NAND2_X1 U14162 ( .A1(n14099), .A2(b_5_), .ZN(n14098) );
  NOR2_X1 U14163 ( .A1(n14100), .A2(n7803), .ZN(n14099) );
  NOR2_X1 U14164 ( .A1(n13844), .A2(n13846), .ZN(n14100) );
  NAND2_X1 U14165 ( .A1(n13844), .A2(n13846), .ZN(n14097) );
  NAND2_X1 U14166 ( .A1(n14101), .A2(n14102), .ZN(n13846) );
  NAND2_X1 U14167 ( .A1(n13864), .A2(n14103), .ZN(n14102) );
  NAND2_X1 U14168 ( .A1(n13866), .A2(n13865), .ZN(n14103) );
  NOR2_X1 U14169 ( .A1(n13620), .A2(n7337), .ZN(n13864) );
  OR2_X1 U14170 ( .A1(n13865), .A2(n13866), .ZN(n14101) );
  AND2_X1 U14171 ( .A1(n14104), .A2(n14105), .ZN(n13866) );
  NAND2_X1 U14172 ( .A1(n14106), .A2(b_3_), .ZN(n14105) );
  NOR2_X1 U14173 ( .A1(n14107), .A2(n7817), .ZN(n14106) );
  NOR2_X1 U14174 ( .A1(n7816), .A2(n13861), .ZN(n14107) );
  NAND2_X1 U14175 ( .A1(n14108), .A2(b_4_), .ZN(n14104) );
  NOR2_X1 U14176 ( .A1(n14109), .A2(n8052), .ZN(n14108) );
  NOR2_X1 U14177 ( .A1(n7810), .A2(n14110), .ZN(n14109) );
  NAND2_X1 U14178 ( .A1(n14111), .A2(b_4_), .ZN(n13865) );
  NOR2_X1 U14179 ( .A1(n8055), .A2(n13620), .ZN(n14111) );
  XOR2_X1 U14180 ( .A(n14112), .B(n14113), .Z(n13844) );
  XOR2_X1 U14181 ( .A(n14114), .B(n14115), .Z(n14112) );
  XOR2_X1 U14182 ( .A(n14116), .B(n14117), .Z(n13871) );
  XOR2_X1 U14183 ( .A(n14118), .B(n14119), .Z(n14116) );
  XOR2_X1 U14184 ( .A(n14120), .B(n14121), .Z(n13814) );
  XOR2_X1 U14185 ( .A(n14122), .B(n14123), .Z(n14120) );
  XOR2_X1 U14186 ( .A(n14124), .B(n14125), .Z(n13876) );
  XOR2_X1 U14187 ( .A(n14126), .B(n14127), .Z(n14124) );
  XOR2_X1 U14188 ( .A(n14128), .B(n14129), .Z(n13880) );
  XOR2_X1 U14189 ( .A(n14130), .B(n14131), .Z(n14128) );
  XNOR2_X1 U14190 ( .A(n14132), .B(n14133), .ZN(n13884) );
  XNOR2_X1 U14191 ( .A(n14134), .B(n14135), .ZN(n14132) );
  XNOR2_X1 U14192 ( .A(n14136), .B(n14137), .ZN(n13888) );
  XNOR2_X1 U14193 ( .A(n14138), .B(n14139), .ZN(n14137) );
  XNOR2_X1 U14194 ( .A(n14140), .B(n14141), .ZN(n13892) );
  XNOR2_X1 U14195 ( .A(n14142), .B(n14143), .ZN(n14140) );
  XOR2_X1 U14196 ( .A(n14144), .B(n14145), .Z(n13896) );
  XOR2_X1 U14197 ( .A(n14146), .B(n14147), .Z(n14144) );
  XNOR2_X1 U14198 ( .A(n14148), .B(n14149), .ZN(n13900) );
  XNOR2_X1 U14199 ( .A(n14150), .B(n14151), .ZN(n14148) );
  XNOR2_X1 U14200 ( .A(n14152), .B(n14153), .ZN(n13904) );
  XNOR2_X1 U14201 ( .A(n14154), .B(n14155), .ZN(n14153) );
  XNOR2_X1 U14202 ( .A(n14156), .B(n14157), .ZN(n13908) );
  XNOR2_X1 U14203 ( .A(n14158), .B(n14159), .ZN(n14156) );
  XNOR2_X1 U14204 ( .A(n14160), .B(n14161), .ZN(n13912) );
  XNOR2_X1 U14205 ( .A(n14162), .B(n14163), .ZN(n14161) );
  XOR2_X1 U14206 ( .A(n14164), .B(n14165), .Z(n13916) );
  XOR2_X1 U14207 ( .A(n14166), .B(n14167), .Z(n14164) );
  NOR2_X1 U14208 ( .A1(n13861), .A2(n7415), .ZN(n14167) );
  XOR2_X1 U14209 ( .A(n14168), .B(n14169), .Z(n13920) );
  XOR2_X1 U14210 ( .A(n14170), .B(n14171), .Z(n14168) );
  NOR2_X1 U14211 ( .A1(n13861), .A2(n7718), .ZN(n14171) );
  XNOR2_X1 U14212 ( .A(n14172), .B(n14173), .ZN(n13924) );
  XOR2_X1 U14213 ( .A(n14174), .B(n14175), .Z(n14173) );
  NAND2_X1 U14214 ( .A1(b_4_), .A2(a_11_), .ZN(n14175) );
  XNOR2_X1 U14215 ( .A(n14176), .B(n14177), .ZN(n13928) );
  XOR2_X1 U14216 ( .A(n14178), .B(n14179), .Z(n14177) );
  NAND2_X1 U14217 ( .A1(a_10_), .A2(b_4_), .ZN(n14179) );
  XNOR2_X1 U14218 ( .A(n14180), .B(n14181), .ZN(n13932) );
  XOR2_X1 U14219 ( .A(n14182), .B(n14183), .Z(n14181) );
  NAND2_X1 U14220 ( .A1(a_9_), .A2(b_4_), .ZN(n14183) );
  XOR2_X1 U14221 ( .A(n14184), .B(n14185), .Z(n13936) );
  XOR2_X1 U14222 ( .A(n14186), .B(n14187), .Z(n14184) );
  NOR2_X1 U14223 ( .A1(n13861), .A2(n7699), .ZN(n14187) );
  XOR2_X1 U14224 ( .A(n14188), .B(n14189), .Z(n13940) );
  XOR2_X1 U14225 ( .A(n14190), .B(n14191), .Z(n14188) );
  NOR2_X1 U14226 ( .A1(n13861), .A2(n7445), .ZN(n14191) );
  XOR2_X1 U14227 ( .A(n14192), .B(n14193), .Z(n13948) );
  XOR2_X1 U14228 ( .A(n14194), .B(n14195), .Z(n14192) );
  NOR2_X1 U14229 ( .A1(n13861), .A2(n7455), .ZN(n14195) );
  XNOR2_X1 U14230 ( .A(n14196), .B(n14197), .ZN(n13952) );
  XNOR2_X1 U14231 ( .A(n14198), .B(n14199), .ZN(n14196) );
  XOR2_X1 U14232 ( .A(n14200), .B(n14201), .Z(n13956) );
  XNOR2_X1 U14233 ( .A(n14202), .B(n14203), .ZN(n14200) );
  NAND2_X1 U14234 ( .A1(a_3_), .A2(b_4_), .ZN(n14202) );
  XOR2_X1 U14235 ( .A(n14204), .B(n14205), .Z(n13960) );
  XOR2_X1 U14236 ( .A(n14206), .B(n14207), .Z(n14204) );
  NOR2_X1 U14237 ( .A1(n13861), .A2(n7469), .ZN(n14207) );
  XOR2_X1 U14238 ( .A(n14208), .B(n14209), .Z(n13964) );
  XOR2_X1 U14239 ( .A(n14210), .B(n14211), .Z(n14208) );
  NOR2_X1 U14240 ( .A1(n13861), .A2(n7669), .ZN(n14211) );
  XNOR2_X1 U14241 ( .A(n13730), .B(n13731), .ZN(n13970) );
  XNOR2_X1 U14242 ( .A(n14212), .B(n14213), .ZN(n13730) );
  NOR2_X1 U14243 ( .A1(n7478), .A2(n13861), .ZN(n14213) );
  NAND2_X1 U14244 ( .A1(n14214), .A2(n14215), .ZN(n7440) );
  OR2_X1 U14245 ( .A1(n14215), .A2(n14214), .ZN(n7439) );
  NAND2_X1 U14246 ( .A1(n14216), .A2(n14217), .ZN(n14214) );
  NAND2_X1 U14247 ( .A1(n14218), .A2(n14219), .ZN(n14217) );
  INV_X1 U14248 ( .A(n14220), .ZN(n14219) );
  XNOR2_X1 U14249 ( .A(n14221), .B(n14222), .ZN(n14218) );
  NAND2_X1 U14250 ( .A1(n13969), .A2(n13968), .ZN(n14215) );
  NAND2_X1 U14251 ( .A1(n14223), .A2(n14224), .ZN(n13968) );
  NAND2_X1 U14252 ( .A1(n14225), .A2(b_4_), .ZN(n14224) );
  NOR2_X1 U14253 ( .A1(n14226), .A2(n7478), .ZN(n14225) );
  NOR2_X1 U14254 ( .A1(n14212), .A2(n13731), .ZN(n14226) );
  NAND2_X1 U14255 ( .A1(n13731), .A2(n14212), .ZN(n14223) );
  NAND2_X1 U14256 ( .A1(n14227), .A2(n14228), .ZN(n14212) );
  NAND2_X1 U14257 ( .A1(n14229), .A2(a_1_), .ZN(n14228) );
  NOR2_X1 U14258 ( .A1(n14230), .A2(n13861), .ZN(n14229) );
  NOR2_X1 U14259 ( .A1(n14209), .A2(n14210), .ZN(n14230) );
  NAND2_X1 U14260 ( .A1(n14209), .A2(n14210), .ZN(n14227) );
  NAND2_X1 U14261 ( .A1(n14231), .A2(n14232), .ZN(n14210) );
  NAND2_X1 U14262 ( .A1(n14233), .A2(a_2_), .ZN(n14232) );
  NOR2_X1 U14263 ( .A1(n14234), .A2(n13861), .ZN(n14233) );
  NOR2_X1 U14264 ( .A1(n14206), .A2(n14205), .ZN(n14234) );
  NAND2_X1 U14265 ( .A1(n14205), .A2(n14206), .ZN(n14231) );
  NAND2_X1 U14266 ( .A1(n14235), .A2(n14236), .ZN(n14206) );
  NAND2_X1 U14267 ( .A1(n14237), .A2(a_3_), .ZN(n14236) );
  NOR2_X1 U14268 ( .A1(n14238), .A2(n13861), .ZN(n14237) );
  NOR2_X1 U14269 ( .A1(n14201), .A2(n14203), .ZN(n14238) );
  NAND2_X1 U14270 ( .A1(n14201), .A2(n14203), .ZN(n14235) );
  NAND2_X1 U14271 ( .A1(n14239), .A2(n14240), .ZN(n14203) );
  NAND2_X1 U14272 ( .A1(n14199), .A2(n14241), .ZN(n14240) );
  NAND2_X1 U14273 ( .A1(n14198), .A2(n14197), .ZN(n14241) );
  OR2_X1 U14274 ( .A1(n14197), .A2(n14198), .ZN(n14239) );
  AND2_X1 U14275 ( .A1(n14242), .A2(n14243), .ZN(n14198) );
  NAND2_X1 U14276 ( .A1(n14244), .A2(a_5_), .ZN(n14243) );
  NOR2_X1 U14277 ( .A1(n14245), .A2(n13861), .ZN(n14244) );
  NOR2_X1 U14278 ( .A1(n14193), .A2(n14194), .ZN(n14245) );
  NAND2_X1 U14279 ( .A1(n14193), .A2(n14194), .ZN(n14242) );
  NAND2_X1 U14280 ( .A1(n14246), .A2(n14247), .ZN(n14194) );
  NAND2_X1 U14281 ( .A1(n14248), .A2(a_6_), .ZN(n14247) );
  NOR2_X1 U14282 ( .A1(n14249), .A2(n13861), .ZN(n14248) );
  NOR2_X1 U14283 ( .A1(n13994), .A2(n13995), .ZN(n14249) );
  NAND2_X1 U14284 ( .A1(n13994), .A2(n13995), .ZN(n14246) );
  NAND2_X1 U14285 ( .A1(n14250), .A2(n14251), .ZN(n13995) );
  NAND2_X1 U14286 ( .A1(n14252), .A2(a_7_), .ZN(n14251) );
  NOR2_X1 U14287 ( .A1(n14253), .A2(n13861), .ZN(n14252) );
  NOR2_X1 U14288 ( .A1(n14189), .A2(n14190), .ZN(n14253) );
  NAND2_X1 U14289 ( .A1(n14189), .A2(n14190), .ZN(n14250) );
  NAND2_X1 U14290 ( .A1(n14254), .A2(n14255), .ZN(n14190) );
  NAND2_X1 U14291 ( .A1(n14256), .A2(a_8_), .ZN(n14255) );
  NOR2_X1 U14292 ( .A1(n14257), .A2(n13861), .ZN(n14256) );
  NOR2_X1 U14293 ( .A1(n14185), .A2(n14186), .ZN(n14257) );
  NAND2_X1 U14294 ( .A1(n14185), .A2(n14186), .ZN(n14254) );
  NAND2_X1 U14295 ( .A1(n14258), .A2(n14259), .ZN(n14186) );
  NAND2_X1 U14296 ( .A1(n14260), .A2(a_9_), .ZN(n14259) );
  NOR2_X1 U14297 ( .A1(n14261), .A2(n13861), .ZN(n14260) );
  NOR2_X1 U14298 ( .A1(n14180), .A2(n14182), .ZN(n14261) );
  NAND2_X1 U14299 ( .A1(n14180), .A2(n14182), .ZN(n14258) );
  NAND2_X1 U14300 ( .A1(n14262), .A2(n14263), .ZN(n14182) );
  NAND2_X1 U14301 ( .A1(n14264), .A2(a_10_), .ZN(n14263) );
  NOR2_X1 U14302 ( .A1(n14265), .A2(n13861), .ZN(n14264) );
  NOR2_X1 U14303 ( .A1(n14176), .A2(n14178), .ZN(n14265) );
  NAND2_X1 U14304 ( .A1(n14176), .A2(n14178), .ZN(n14262) );
  NAND2_X1 U14305 ( .A1(n14266), .A2(n14267), .ZN(n14178) );
  NAND2_X1 U14306 ( .A1(n14268), .A2(b_4_), .ZN(n14267) );
  NOR2_X1 U14307 ( .A1(n14269), .A2(n7424), .ZN(n14268) );
  NOR2_X1 U14308 ( .A1(n14172), .A2(n14174), .ZN(n14269) );
  NAND2_X1 U14309 ( .A1(n14172), .A2(n14174), .ZN(n14266) );
  NAND2_X1 U14310 ( .A1(n14270), .A2(n14271), .ZN(n14174) );
  NAND2_X1 U14311 ( .A1(n14272), .A2(a_12_), .ZN(n14271) );
  NOR2_X1 U14312 ( .A1(n14273), .A2(n13861), .ZN(n14272) );
  NOR2_X1 U14313 ( .A1(n14169), .A2(n14170), .ZN(n14273) );
  NAND2_X1 U14314 ( .A1(n14169), .A2(n14170), .ZN(n14270) );
  NAND2_X1 U14315 ( .A1(n14274), .A2(n14275), .ZN(n14170) );
  NAND2_X1 U14316 ( .A1(n14276), .A2(a_13_), .ZN(n14275) );
  NOR2_X1 U14317 ( .A1(n14277), .A2(n13861), .ZN(n14276) );
  NOR2_X1 U14318 ( .A1(n14165), .A2(n14166), .ZN(n14277) );
  NAND2_X1 U14319 ( .A1(n14165), .A2(n14166), .ZN(n14274) );
  NAND2_X1 U14320 ( .A1(n14278), .A2(n14279), .ZN(n14166) );
  NAND2_X1 U14321 ( .A1(n14163), .A2(n14280), .ZN(n14279) );
  OR2_X1 U14322 ( .A1(n14162), .A2(n14160), .ZN(n14280) );
  NOR2_X1 U14323 ( .A1(n7727), .A2(n13861), .ZN(n14163) );
  NAND2_X1 U14324 ( .A1(n14160), .A2(n14162), .ZN(n14278) );
  NAND2_X1 U14325 ( .A1(n14281), .A2(n14282), .ZN(n14162) );
  NAND2_X1 U14326 ( .A1(n14159), .A2(n14283), .ZN(n14282) );
  NAND2_X1 U14327 ( .A1(n14158), .A2(n14157), .ZN(n14283) );
  NOR2_X1 U14328 ( .A1(n7406), .A2(n13861), .ZN(n14159) );
  OR2_X1 U14329 ( .A1(n14157), .A2(n14158), .ZN(n14281) );
  AND2_X1 U14330 ( .A1(n14284), .A2(n14285), .ZN(n14158) );
  NAND2_X1 U14331 ( .A1(n14155), .A2(n14286), .ZN(n14285) );
  OR2_X1 U14332 ( .A1(n14152), .A2(n14154), .ZN(n14286) );
  NOR2_X1 U14333 ( .A1(n7736), .A2(n13861), .ZN(n14155) );
  NAND2_X1 U14334 ( .A1(n14152), .A2(n14154), .ZN(n14284) );
  NAND2_X1 U14335 ( .A1(n14287), .A2(n14288), .ZN(n14154) );
  NAND2_X1 U14336 ( .A1(n14151), .A2(n14289), .ZN(n14288) );
  NAND2_X1 U14337 ( .A1(n14150), .A2(n14149), .ZN(n14289) );
  NOR2_X1 U14338 ( .A1(n7397), .A2(n13861), .ZN(n14151) );
  OR2_X1 U14339 ( .A1(n14149), .A2(n14150), .ZN(n14287) );
  AND2_X1 U14340 ( .A1(n14290), .A2(n14291), .ZN(n14150) );
  NAND2_X1 U14341 ( .A1(n14147), .A2(n14292), .ZN(n14291) );
  OR2_X1 U14342 ( .A1(n14145), .A2(n14146), .ZN(n14292) );
  NOR2_X1 U14343 ( .A1(n7745), .A2(n13861), .ZN(n14147) );
  NAND2_X1 U14344 ( .A1(n14145), .A2(n14146), .ZN(n14290) );
  NAND2_X1 U14345 ( .A1(n14293), .A2(n14294), .ZN(n14146) );
  NAND2_X1 U14346 ( .A1(n14143), .A2(n14295), .ZN(n14294) );
  NAND2_X1 U14347 ( .A1(n14142), .A2(n14141), .ZN(n14295) );
  NOR2_X1 U14348 ( .A1(n7750), .A2(n13861), .ZN(n14143) );
  OR2_X1 U14349 ( .A1(n14141), .A2(n14142), .ZN(n14293) );
  AND2_X1 U14350 ( .A1(n14296), .A2(n14297), .ZN(n14142) );
  NAND2_X1 U14351 ( .A1(n14139), .A2(n14298), .ZN(n14297) );
  OR2_X1 U14352 ( .A1(n14136), .A2(n14138), .ZN(n14298) );
  NOR2_X1 U14353 ( .A1(n13861), .A2(n7755), .ZN(n14139) );
  NAND2_X1 U14354 ( .A1(n14136), .A2(n14138), .ZN(n14296) );
  NAND2_X1 U14355 ( .A1(n14299), .A2(n14300), .ZN(n14138) );
  NAND2_X1 U14356 ( .A1(n14135), .A2(n14301), .ZN(n14300) );
  NAND2_X1 U14357 ( .A1(n14134), .A2(n14133), .ZN(n14301) );
  NOR2_X1 U14358 ( .A1(n13861), .A2(n7760), .ZN(n14135) );
  OR2_X1 U14359 ( .A1(n14133), .A2(n14134), .ZN(n14299) );
  AND2_X1 U14360 ( .A1(n14302), .A2(n14303), .ZN(n14134) );
  NAND2_X1 U14361 ( .A1(n14131), .A2(n14304), .ZN(n14303) );
  OR2_X1 U14362 ( .A1(n14129), .A2(n14130), .ZN(n14304) );
  NOR2_X1 U14363 ( .A1(n7765), .A2(n13861), .ZN(n14131) );
  NAND2_X1 U14364 ( .A1(n14129), .A2(n14130), .ZN(n14302) );
  NAND2_X1 U14365 ( .A1(n14305), .A2(n14306), .ZN(n14130) );
  NAND2_X1 U14366 ( .A1(n14127), .A2(n14307), .ZN(n14306) );
  OR2_X1 U14367 ( .A1(n14125), .A2(n14126), .ZN(n14307) );
  NOR2_X1 U14368 ( .A1(n13861), .A2(n8014), .ZN(n14127) );
  NAND2_X1 U14369 ( .A1(n14125), .A2(n14126), .ZN(n14305) );
  NAND2_X1 U14370 ( .A1(n14308), .A2(n14309), .ZN(n14126) );
  NAND2_X1 U14371 ( .A1(n14123), .A2(n14310), .ZN(n14309) );
  OR2_X1 U14372 ( .A1(n14121), .A2(n14122), .ZN(n14310) );
  NOR2_X1 U14373 ( .A1(n7774), .A2(n13861), .ZN(n14123) );
  NAND2_X1 U14374 ( .A1(n14121), .A2(n14122), .ZN(n14308) );
  NAND2_X1 U14375 ( .A1(n14311), .A2(n14312), .ZN(n14122) );
  NAND2_X1 U14376 ( .A1(n14119), .A2(n14313), .ZN(n14312) );
  OR2_X1 U14377 ( .A1(n14117), .A2(n14118), .ZN(n14313) );
  NOR2_X1 U14378 ( .A1(n13861), .A2(n8022), .ZN(n14119) );
  NAND2_X1 U14379 ( .A1(n14117), .A2(n14118), .ZN(n14311) );
  NAND2_X1 U14380 ( .A1(n14079), .A2(n14314), .ZN(n14118) );
  NAND2_X1 U14381 ( .A1(n14078), .A2(n14080), .ZN(n14314) );
  NAND2_X1 U14382 ( .A1(n14315), .A2(n14316), .ZN(n14080) );
  NAND2_X1 U14383 ( .A1(b_4_), .A2(a_26_), .ZN(n14316) );
  INV_X1 U14384 ( .A(n14317), .ZN(n14315) );
  XNOR2_X1 U14385 ( .A(n14318), .B(n14319), .ZN(n14078) );
  NAND2_X1 U14386 ( .A1(n14320), .A2(n14321), .ZN(n14318) );
  NAND2_X1 U14387 ( .A1(a_26_), .A2(n14317), .ZN(n14079) );
  NAND2_X1 U14388 ( .A1(n14087), .A2(n14322), .ZN(n14317) );
  NAND2_X1 U14389 ( .A1(n14086), .A2(n14088), .ZN(n14322) );
  NAND2_X1 U14390 ( .A1(n14323), .A2(n14324), .ZN(n14088) );
  NAND2_X1 U14391 ( .A1(b_4_), .A2(a_27_), .ZN(n14324) );
  INV_X1 U14392 ( .A(n14325), .ZN(n14323) );
  XNOR2_X1 U14393 ( .A(n14326), .B(n14327), .ZN(n14086) );
  XOR2_X1 U14394 ( .A(n14328), .B(n14329), .Z(n14327) );
  NAND2_X1 U14395 ( .A1(b_3_), .A2(a_28_), .ZN(n14329) );
  NAND2_X1 U14396 ( .A1(a_27_), .A2(n14325), .ZN(n14087) );
  NAND2_X1 U14397 ( .A1(n14330), .A2(n14331), .ZN(n14325) );
  NAND2_X1 U14398 ( .A1(n14332), .A2(b_4_), .ZN(n14331) );
  NOR2_X1 U14399 ( .A1(n14333), .A2(n7803), .ZN(n14332) );
  NOR2_X1 U14400 ( .A1(n14093), .A2(n14095), .ZN(n14333) );
  NAND2_X1 U14401 ( .A1(n14093), .A2(n14095), .ZN(n14330) );
  NAND2_X1 U14402 ( .A1(n14334), .A2(n14335), .ZN(n14095) );
  NAND2_X1 U14403 ( .A1(n14113), .A2(n14336), .ZN(n14335) );
  NAND2_X1 U14404 ( .A1(n14115), .A2(n14114), .ZN(n14336) );
  NOR2_X1 U14405 ( .A1(n13861), .A2(n7337), .ZN(n14113) );
  OR2_X1 U14406 ( .A1(n14114), .A2(n14115), .ZN(n14334) );
  AND2_X1 U14407 ( .A1(n14337), .A2(n14338), .ZN(n14115) );
  NAND2_X1 U14408 ( .A1(n14339), .A2(b_2_), .ZN(n14338) );
  NOR2_X1 U14409 ( .A1(n14340), .A2(n7817), .ZN(n14339) );
  NOR2_X1 U14410 ( .A1(n7816), .A2(n14110), .ZN(n14340) );
  NAND2_X1 U14411 ( .A1(n14341), .A2(b_3_), .ZN(n14337) );
  NOR2_X1 U14412 ( .A1(n14342), .A2(n8052), .ZN(n14341) );
  NOR2_X1 U14413 ( .A1(n7810), .A2(n14343), .ZN(n14342) );
  NAND2_X1 U14414 ( .A1(n14344), .A2(b_3_), .ZN(n14114) );
  NOR2_X1 U14415 ( .A1(n8055), .A2(n13861), .ZN(n14344) );
  XOR2_X1 U14416 ( .A(n14345), .B(n14346), .Z(n14093) );
  XOR2_X1 U14417 ( .A(n14347), .B(n14348), .Z(n14345) );
  XNOR2_X1 U14418 ( .A(n14349), .B(n14350), .ZN(n14117) );
  NAND2_X1 U14419 ( .A1(n14351), .A2(n14352), .ZN(n14349) );
  XNOR2_X1 U14420 ( .A(n14353), .B(n14354), .ZN(n14121) );
  NAND2_X1 U14421 ( .A1(n14355), .A2(n14356), .ZN(n14353) );
  XOR2_X1 U14422 ( .A(n14357), .B(n14358), .Z(n14125) );
  XOR2_X1 U14423 ( .A(n14359), .B(n14360), .Z(n14357) );
  NOR2_X1 U14424 ( .A1(n7774), .A2(n14110), .ZN(n14360) );
  XNOR2_X1 U14425 ( .A(n14361), .B(n14362), .ZN(n14129) );
  NAND2_X1 U14426 ( .A1(n14363), .A2(n14364), .ZN(n14361) );
  XNOR2_X1 U14427 ( .A(n14365), .B(n14366), .ZN(n14133) );
  XOR2_X1 U14428 ( .A(n14367), .B(n14368), .Z(n14365) );
  NOR2_X1 U14429 ( .A1(n14110), .A2(n7765), .ZN(n14368) );
  XNOR2_X1 U14430 ( .A(n14369), .B(n14370), .ZN(n14136) );
  NAND2_X1 U14431 ( .A1(n14371), .A2(n14372), .ZN(n14369) );
  XNOR2_X1 U14432 ( .A(n14373), .B(n14374), .ZN(n14141) );
  XNOR2_X1 U14433 ( .A(n14375), .B(n14376), .ZN(n14373) );
  NAND2_X1 U14434 ( .A1(b_3_), .A2(a_20_), .ZN(n14375) );
  XNOR2_X1 U14435 ( .A(n14377), .B(n14378), .ZN(n14145) );
  NAND2_X1 U14436 ( .A1(n14379), .A2(n14380), .ZN(n14377) );
  XNOR2_X1 U14437 ( .A(n14381), .B(n14382), .ZN(n14149) );
  XOR2_X1 U14438 ( .A(n14383), .B(n14384), .Z(n14381) );
  NOR2_X1 U14439 ( .A1(n14110), .A2(n7745), .ZN(n14384) );
  XNOR2_X1 U14440 ( .A(n14385), .B(n14386), .ZN(n14152) );
  NAND2_X1 U14441 ( .A1(n14387), .A2(n14388), .ZN(n14385) );
  XNOR2_X1 U14442 ( .A(n14389), .B(n14390), .ZN(n14157) );
  XOR2_X1 U14443 ( .A(n14391), .B(n14392), .Z(n14389) );
  NOR2_X1 U14444 ( .A1(n14110), .A2(n7736), .ZN(n14392) );
  XNOR2_X1 U14445 ( .A(n14393), .B(n14394), .ZN(n14160) );
  NAND2_X1 U14446 ( .A1(n14395), .A2(n14396), .ZN(n14393) );
  XOR2_X1 U14447 ( .A(n14397), .B(n14398), .Z(n14165) );
  XOR2_X1 U14448 ( .A(n14399), .B(n14400), .Z(n14397) );
  NOR2_X1 U14449 ( .A1(n14110), .A2(n7727), .ZN(n14400) );
  XNOR2_X1 U14450 ( .A(n14401), .B(n14402), .ZN(n14169) );
  NAND2_X1 U14451 ( .A1(n14403), .A2(n14404), .ZN(n14401) );
  XOR2_X1 U14452 ( .A(n14405), .B(n14406), .Z(n14172) );
  XOR2_X1 U14453 ( .A(n14407), .B(n14408), .Z(n14405) );
  NOR2_X1 U14454 ( .A1(n14110), .A2(n7718), .ZN(n14408) );
  XNOR2_X1 U14455 ( .A(n14409), .B(n14410), .ZN(n14176) );
  NAND2_X1 U14456 ( .A1(n14411), .A2(n14412), .ZN(n14409) );
  XOR2_X1 U14457 ( .A(n14413), .B(n14414), .Z(n14180) );
  XOR2_X1 U14458 ( .A(n14415), .B(n14416), .Z(n14413) );
  NOR2_X1 U14459 ( .A1(n14110), .A2(n7709), .ZN(n14416) );
  XNOR2_X1 U14460 ( .A(n14417), .B(n14418), .ZN(n14185) );
  NAND2_X1 U14461 ( .A1(n14419), .A2(n14420), .ZN(n14417) );
  XOR2_X1 U14462 ( .A(n14421), .B(n14422), .Z(n14189) );
  XOR2_X1 U14463 ( .A(n14423), .B(n14424), .Z(n14421) );
  NOR2_X1 U14464 ( .A1(n14110), .A2(n7699), .ZN(n14424) );
  XNOR2_X1 U14465 ( .A(n14425), .B(n14426), .ZN(n13994) );
  NAND2_X1 U14466 ( .A1(n14427), .A2(n14428), .ZN(n14425) );
  XOR2_X1 U14467 ( .A(n14429), .B(n14430), .Z(n14193) );
  XOR2_X1 U14468 ( .A(n14431), .B(n14432), .Z(n14429) );
  NOR2_X1 U14469 ( .A1(n14110), .A2(n7450), .ZN(n14432) );
  XOR2_X1 U14470 ( .A(n14433), .B(n14434), .Z(n14197) );
  NAND2_X1 U14471 ( .A1(n14435), .A2(n14436), .ZN(n14433) );
  XOR2_X1 U14472 ( .A(n14437), .B(n14438), .Z(n14201) );
  XOR2_X1 U14473 ( .A(n14439), .B(n14440), .Z(n14437) );
  NOR2_X1 U14474 ( .A1(n14110), .A2(n7682), .ZN(n14440) );
  XOR2_X1 U14475 ( .A(n14441), .B(n14442), .Z(n14205) );
  XOR2_X1 U14476 ( .A(n14443), .B(n14444), .Z(n14441) );
  XOR2_X1 U14477 ( .A(n14445), .B(n14446), .Z(n14209) );
  XOR2_X1 U14478 ( .A(n14447), .B(n14448), .Z(n14445) );
  NOR2_X1 U14479 ( .A1(n14110), .A2(n7469), .ZN(n14448) );
  XNOR2_X1 U14480 ( .A(n14449), .B(n14450), .ZN(n13731) );
  NAND2_X1 U14481 ( .A1(n14451), .A2(n14452), .ZN(n14449) );
  XOR2_X1 U14482 ( .A(n14453), .B(n14454), .Z(n13969) );
  XOR2_X1 U14483 ( .A(n14455), .B(n14456), .Z(n14453) );
  NAND2_X1 U14484 ( .A1(n14457), .A2(n14216), .ZN(n7487) );
  XNOR2_X1 U14485 ( .A(n14458), .B(n14459), .ZN(n14457) );
  OR2_X1 U14486 ( .A1(n14460), .A2(n14216), .ZN(n7488) );
  NAND2_X1 U14487 ( .A1(n14461), .A2(n14220), .ZN(n14216) );
  NAND2_X1 U14488 ( .A1(n14462), .A2(n14463), .ZN(n14220) );
  NAND2_X1 U14489 ( .A1(n14456), .A2(n14464), .ZN(n14463) );
  OR2_X1 U14490 ( .A1(n14454), .A2(n14455), .ZN(n14464) );
  NOR2_X1 U14491 ( .A1(n14110), .A2(n7478), .ZN(n14456) );
  NAND2_X1 U14492 ( .A1(n14454), .A2(n14455), .ZN(n14462) );
  NAND2_X1 U14493 ( .A1(n14451), .A2(n14465), .ZN(n14455) );
  NAND2_X1 U14494 ( .A1(n14450), .A2(n14452), .ZN(n14465) );
  NAND2_X1 U14495 ( .A1(n14466), .A2(n14467), .ZN(n14452) );
  NAND2_X1 U14496 ( .A1(a_1_), .A2(b_3_), .ZN(n14467) );
  INV_X1 U14497 ( .A(n14468), .ZN(n14466) );
  XNOR2_X1 U14498 ( .A(n14469), .B(n14470), .ZN(n14450) );
  XNOR2_X1 U14499 ( .A(n14471), .B(n14472), .ZN(n14469) );
  NAND2_X1 U14500 ( .A1(a_1_), .A2(n14468), .ZN(n14451) );
  NAND2_X1 U14501 ( .A1(n14473), .A2(n14474), .ZN(n14468) );
  NAND2_X1 U14502 ( .A1(n14475), .A2(a_2_), .ZN(n14474) );
  NOR2_X1 U14503 ( .A1(n14476), .A2(n14110), .ZN(n14475) );
  NOR2_X1 U14504 ( .A1(n14447), .A2(n14446), .ZN(n14476) );
  NAND2_X1 U14505 ( .A1(n14446), .A2(n14447), .ZN(n14473) );
  NAND2_X1 U14506 ( .A1(n14477), .A2(n14478), .ZN(n14447) );
  NAND2_X1 U14507 ( .A1(n14442), .A2(n14479), .ZN(n14478) );
  OR2_X1 U14508 ( .A1(n14443), .A2(n14444), .ZN(n14479) );
  XNOR2_X1 U14509 ( .A(n14480), .B(n14481), .ZN(n14442) );
  NAND2_X1 U14510 ( .A1(n14482), .A2(n14483), .ZN(n14480) );
  NAND2_X1 U14511 ( .A1(n14444), .A2(n14443), .ZN(n14477) );
  NAND2_X1 U14512 ( .A1(n14484), .A2(n14485), .ZN(n14443) );
  NAND2_X1 U14513 ( .A1(n14486), .A2(a_4_), .ZN(n14485) );
  NOR2_X1 U14514 ( .A1(n14487), .A2(n14110), .ZN(n14486) );
  NOR2_X1 U14515 ( .A1(n14439), .A2(n14438), .ZN(n14487) );
  NAND2_X1 U14516 ( .A1(n14438), .A2(n14439), .ZN(n14484) );
  NAND2_X1 U14517 ( .A1(n14435), .A2(n14488), .ZN(n14439) );
  NAND2_X1 U14518 ( .A1(n14434), .A2(n14436), .ZN(n14488) );
  NAND2_X1 U14519 ( .A1(n14489), .A2(n14490), .ZN(n14436) );
  NAND2_X1 U14520 ( .A1(a_5_), .A2(b_3_), .ZN(n14490) );
  INV_X1 U14521 ( .A(n14491), .ZN(n14489) );
  XNOR2_X1 U14522 ( .A(n14492), .B(n14493), .ZN(n14434) );
  NAND2_X1 U14523 ( .A1(n14494), .A2(n14495), .ZN(n14492) );
  NAND2_X1 U14524 ( .A1(a_5_), .A2(n14491), .ZN(n14435) );
  NAND2_X1 U14525 ( .A1(n14496), .A2(n14497), .ZN(n14491) );
  NAND2_X1 U14526 ( .A1(n14498), .A2(a_6_), .ZN(n14497) );
  NOR2_X1 U14527 ( .A1(n14499), .A2(n14110), .ZN(n14498) );
  NOR2_X1 U14528 ( .A1(n14431), .A2(n14430), .ZN(n14499) );
  NAND2_X1 U14529 ( .A1(n14430), .A2(n14431), .ZN(n14496) );
  NAND2_X1 U14530 ( .A1(n14427), .A2(n14500), .ZN(n14431) );
  NAND2_X1 U14531 ( .A1(n14426), .A2(n14428), .ZN(n14500) );
  NAND2_X1 U14532 ( .A1(n14501), .A2(n14502), .ZN(n14428) );
  NAND2_X1 U14533 ( .A1(a_7_), .A2(b_3_), .ZN(n14502) );
  INV_X1 U14534 ( .A(n14503), .ZN(n14501) );
  XNOR2_X1 U14535 ( .A(n14504), .B(n14505), .ZN(n14426) );
  NAND2_X1 U14536 ( .A1(n14506), .A2(n14507), .ZN(n14504) );
  NAND2_X1 U14537 ( .A1(a_7_), .A2(n14503), .ZN(n14427) );
  NAND2_X1 U14538 ( .A1(n14508), .A2(n14509), .ZN(n14503) );
  NAND2_X1 U14539 ( .A1(n14510), .A2(a_8_), .ZN(n14509) );
  NOR2_X1 U14540 ( .A1(n14511), .A2(n14110), .ZN(n14510) );
  NOR2_X1 U14541 ( .A1(n14423), .A2(n14422), .ZN(n14511) );
  NAND2_X1 U14542 ( .A1(n14422), .A2(n14423), .ZN(n14508) );
  NAND2_X1 U14543 ( .A1(n14419), .A2(n14512), .ZN(n14423) );
  NAND2_X1 U14544 ( .A1(n14418), .A2(n14420), .ZN(n14512) );
  NAND2_X1 U14545 ( .A1(n14513), .A2(n14514), .ZN(n14420) );
  NAND2_X1 U14546 ( .A1(a_9_), .A2(b_3_), .ZN(n14514) );
  INV_X1 U14547 ( .A(n14515), .ZN(n14513) );
  XNOR2_X1 U14548 ( .A(n14516), .B(n14517), .ZN(n14418) );
  NAND2_X1 U14549 ( .A1(n14518), .A2(n14519), .ZN(n14516) );
  NAND2_X1 U14550 ( .A1(a_9_), .A2(n14515), .ZN(n14419) );
  NAND2_X1 U14551 ( .A1(n14520), .A2(n14521), .ZN(n14515) );
  NAND2_X1 U14552 ( .A1(n14522), .A2(a_10_), .ZN(n14521) );
  NOR2_X1 U14553 ( .A1(n14523), .A2(n14110), .ZN(n14522) );
  NOR2_X1 U14554 ( .A1(n14415), .A2(n14414), .ZN(n14523) );
  NAND2_X1 U14555 ( .A1(n14414), .A2(n14415), .ZN(n14520) );
  NAND2_X1 U14556 ( .A1(n14411), .A2(n14524), .ZN(n14415) );
  NAND2_X1 U14557 ( .A1(n14410), .A2(n14412), .ZN(n14524) );
  NAND2_X1 U14558 ( .A1(n14525), .A2(n14526), .ZN(n14412) );
  NAND2_X1 U14559 ( .A1(b_3_), .A2(a_11_), .ZN(n14526) );
  INV_X1 U14560 ( .A(n14527), .ZN(n14525) );
  XNOR2_X1 U14561 ( .A(n14528), .B(n14529), .ZN(n14410) );
  NAND2_X1 U14562 ( .A1(n14530), .A2(n14531), .ZN(n14528) );
  NAND2_X1 U14563 ( .A1(a_11_), .A2(n14527), .ZN(n14411) );
  NAND2_X1 U14564 ( .A1(n14532), .A2(n14533), .ZN(n14527) );
  NAND2_X1 U14565 ( .A1(n14534), .A2(a_12_), .ZN(n14533) );
  NOR2_X1 U14566 ( .A1(n14535), .A2(n14110), .ZN(n14534) );
  NOR2_X1 U14567 ( .A1(n14407), .A2(n14406), .ZN(n14535) );
  NAND2_X1 U14568 ( .A1(n14406), .A2(n14407), .ZN(n14532) );
  NAND2_X1 U14569 ( .A1(n14403), .A2(n14536), .ZN(n14407) );
  NAND2_X1 U14570 ( .A1(n14402), .A2(n14404), .ZN(n14536) );
  NAND2_X1 U14571 ( .A1(n14537), .A2(n14538), .ZN(n14404) );
  NAND2_X1 U14572 ( .A1(a_13_), .A2(b_3_), .ZN(n14538) );
  INV_X1 U14573 ( .A(n14539), .ZN(n14537) );
  XNOR2_X1 U14574 ( .A(n14540), .B(n14541), .ZN(n14402) );
  NAND2_X1 U14575 ( .A1(n14542), .A2(n14543), .ZN(n14540) );
  NAND2_X1 U14576 ( .A1(a_13_), .A2(n14539), .ZN(n14403) );
  NAND2_X1 U14577 ( .A1(n14544), .A2(n14545), .ZN(n14539) );
  NAND2_X1 U14578 ( .A1(n14546), .A2(a_14_), .ZN(n14545) );
  NOR2_X1 U14579 ( .A1(n14547), .A2(n14110), .ZN(n14546) );
  NOR2_X1 U14580 ( .A1(n14399), .A2(n14398), .ZN(n14547) );
  NAND2_X1 U14581 ( .A1(n14398), .A2(n14399), .ZN(n14544) );
  NAND2_X1 U14582 ( .A1(n14395), .A2(n14548), .ZN(n14399) );
  NAND2_X1 U14583 ( .A1(n14394), .A2(n14396), .ZN(n14548) );
  NAND2_X1 U14584 ( .A1(n14549), .A2(n14550), .ZN(n14396) );
  NAND2_X1 U14585 ( .A1(a_15_), .A2(b_3_), .ZN(n14550) );
  INV_X1 U14586 ( .A(n14551), .ZN(n14549) );
  XNOR2_X1 U14587 ( .A(n14552), .B(n14553), .ZN(n14394) );
  NAND2_X1 U14588 ( .A1(n14554), .A2(n14555), .ZN(n14552) );
  NAND2_X1 U14589 ( .A1(a_15_), .A2(n14551), .ZN(n14395) );
  NAND2_X1 U14590 ( .A1(n14556), .A2(n14557), .ZN(n14551) );
  NAND2_X1 U14591 ( .A1(n14558), .A2(a_16_), .ZN(n14557) );
  NOR2_X1 U14592 ( .A1(n14559), .A2(n14110), .ZN(n14558) );
  NOR2_X1 U14593 ( .A1(n14391), .A2(n14390), .ZN(n14559) );
  NAND2_X1 U14594 ( .A1(n14390), .A2(n14391), .ZN(n14556) );
  NAND2_X1 U14595 ( .A1(n14387), .A2(n14560), .ZN(n14391) );
  NAND2_X1 U14596 ( .A1(n14386), .A2(n14388), .ZN(n14560) );
  NAND2_X1 U14597 ( .A1(n14561), .A2(n14562), .ZN(n14388) );
  NAND2_X1 U14598 ( .A1(a_17_), .A2(b_3_), .ZN(n14562) );
  INV_X1 U14599 ( .A(n14563), .ZN(n14561) );
  XNOR2_X1 U14600 ( .A(n14564), .B(n14565), .ZN(n14386) );
  XNOR2_X1 U14601 ( .A(n14566), .B(n14567), .ZN(n14564) );
  NAND2_X1 U14602 ( .A1(a_17_), .A2(n14563), .ZN(n14387) );
  NAND2_X1 U14603 ( .A1(n14568), .A2(n14569), .ZN(n14563) );
  NAND2_X1 U14604 ( .A1(n14570), .A2(a_18_), .ZN(n14569) );
  NOR2_X1 U14605 ( .A1(n14571), .A2(n14110), .ZN(n14570) );
  NOR2_X1 U14606 ( .A1(n14383), .A2(n14382), .ZN(n14571) );
  NAND2_X1 U14607 ( .A1(n14382), .A2(n14383), .ZN(n14568) );
  NAND2_X1 U14608 ( .A1(n14379), .A2(n14572), .ZN(n14383) );
  NAND2_X1 U14609 ( .A1(n14378), .A2(n14380), .ZN(n14572) );
  NAND2_X1 U14610 ( .A1(n14573), .A2(n14574), .ZN(n14380) );
  NAND2_X1 U14611 ( .A1(a_19_), .A2(b_3_), .ZN(n14574) );
  INV_X1 U14612 ( .A(n14575), .ZN(n14573) );
  XNOR2_X1 U14613 ( .A(n14576), .B(n14577), .ZN(n14378) );
  XNOR2_X1 U14614 ( .A(n14578), .B(n14579), .ZN(n14576) );
  NAND2_X1 U14615 ( .A1(a_19_), .A2(n14575), .ZN(n14379) );
  NAND2_X1 U14616 ( .A1(n14580), .A2(n14581), .ZN(n14575) );
  NAND2_X1 U14617 ( .A1(n14582), .A2(b_3_), .ZN(n14581) );
  NOR2_X1 U14618 ( .A1(n14583), .A2(n7755), .ZN(n14582) );
  NOR2_X1 U14619 ( .A1(n14376), .A2(n14374), .ZN(n14583) );
  NAND2_X1 U14620 ( .A1(n14374), .A2(n14376), .ZN(n14580) );
  NAND2_X1 U14621 ( .A1(n14371), .A2(n14584), .ZN(n14376) );
  NAND2_X1 U14622 ( .A1(n14370), .A2(n14372), .ZN(n14584) );
  NAND2_X1 U14623 ( .A1(n14585), .A2(n14586), .ZN(n14372) );
  NAND2_X1 U14624 ( .A1(b_3_), .A2(a_21_), .ZN(n14586) );
  INV_X1 U14625 ( .A(n14587), .ZN(n14585) );
  XNOR2_X1 U14626 ( .A(n14588), .B(n14589), .ZN(n14370) );
  XNOR2_X1 U14627 ( .A(n14590), .B(n14591), .ZN(n14589) );
  NAND2_X1 U14628 ( .A1(a_21_), .A2(n14587), .ZN(n14371) );
  NAND2_X1 U14629 ( .A1(n14592), .A2(n14593), .ZN(n14587) );
  NAND2_X1 U14630 ( .A1(n14594), .A2(a_22_), .ZN(n14593) );
  NOR2_X1 U14631 ( .A1(n14595), .A2(n14110), .ZN(n14594) );
  NOR2_X1 U14632 ( .A1(n14367), .A2(n14366), .ZN(n14595) );
  NAND2_X1 U14633 ( .A1(n14366), .A2(n14367), .ZN(n14592) );
  NAND2_X1 U14634 ( .A1(n14363), .A2(n14596), .ZN(n14367) );
  NAND2_X1 U14635 ( .A1(n14362), .A2(n14364), .ZN(n14596) );
  NAND2_X1 U14636 ( .A1(n14597), .A2(n14598), .ZN(n14364) );
  NAND2_X1 U14637 ( .A1(b_3_), .A2(a_23_), .ZN(n14598) );
  INV_X1 U14638 ( .A(n14599), .ZN(n14597) );
  XNOR2_X1 U14639 ( .A(n14600), .B(n14601), .ZN(n14362) );
  XNOR2_X1 U14640 ( .A(n14602), .B(n14603), .ZN(n14601) );
  NAND2_X1 U14641 ( .A1(a_23_), .A2(n14599), .ZN(n14363) );
  NAND2_X1 U14642 ( .A1(n14604), .A2(n14605), .ZN(n14599) );
  NAND2_X1 U14643 ( .A1(n14606), .A2(b_3_), .ZN(n14605) );
  NOR2_X1 U14644 ( .A1(n14607), .A2(n7774), .ZN(n14606) );
  NOR2_X1 U14645 ( .A1(n14358), .A2(n14359), .ZN(n14607) );
  NAND2_X1 U14646 ( .A1(n14358), .A2(n14359), .ZN(n14604) );
  NAND2_X1 U14647 ( .A1(n14355), .A2(n14608), .ZN(n14359) );
  NAND2_X1 U14648 ( .A1(n14354), .A2(n14356), .ZN(n14608) );
  NAND2_X1 U14649 ( .A1(n14609), .A2(n14610), .ZN(n14356) );
  NAND2_X1 U14650 ( .A1(b_3_), .A2(a_25_), .ZN(n14610) );
  INV_X1 U14651 ( .A(n14611), .ZN(n14609) );
  XNOR2_X1 U14652 ( .A(n14612), .B(n14613), .ZN(n14354) );
  XOR2_X1 U14653 ( .A(n14614), .B(n14615), .Z(n14613) );
  NAND2_X1 U14654 ( .A1(b_2_), .A2(a_26_), .ZN(n14615) );
  NAND2_X1 U14655 ( .A1(a_25_), .A2(n14611), .ZN(n14355) );
  NAND2_X1 U14656 ( .A1(n14351), .A2(n14616), .ZN(n14611) );
  NAND2_X1 U14657 ( .A1(n14350), .A2(n14352), .ZN(n14616) );
  NAND2_X1 U14658 ( .A1(n14617), .A2(n14618), .ZN(n14352) );
  NAND2_X1 U14659 ( .A1(b_3_), .A2(a_26_), .ZN(n14618) );
  INV_X1 U14660 ( .A(n14619), .ZN(n14617) );
  XNOR2_X1 U14661 ( .A(n14620), .B(n14621), .ZN(n14350) );
  XNOR2_X1 U14662 ( .A(n14622), .B(n14623), .ZN(n14620) );
  NAND2_X1 U14663 ( .A1(a_26_), .A2(n14619), .ZN(n14351) );
  NAND2_X1 U14664 ( .A1(n14320), .A2(n14624), .ZN(n14619) );
  NAND2_X1 U14665 ( .A1(n14319), .A2(n14321), .ZN(n14624) );
  NAND2_X1 U14666 ( .A1(n14625), .A2(n14626), .ZN(n14321) );
  NAND2_X1 U14667 ( .A1(b_3_), .A2(a_27_), .ZN(n14626) );
  INV_X1 U14668 ( .A(n14627), .ZN(n14625) );
  XOR2_X1 U14669 ( .A(n14628), .B(n14629), .Z(n14319) );
  XNOR2_X1 U14670 ( .A(n14630), .B(n14631), .ZN(n14628) );
  NAND2_X1 U14671 ( .A1(b_2_), .A2(a_28_), .ZN(n14630) );
  NAND2_X1 U14672 ( .A1(a_27_), .A2(n14627), .ZN(n14320) );
  NAND2_X1 U14673 ( .A1(n14632), .A2(n14633), .ZN(n14627) );
  NAND2_X1 U14674 ( .A1(n14634), .A2(b_3_), .ZN(n14633) );
  NOR2_X1 U14675 ( .A1(n14635), .A2(n7803), .ZN(n14634) );
  NOR2_X1 U14676 ( .A1(n14326), .A2(n14328), .ZN(n14635) );
  NAND2_X1 U14677 ( .A1(n14326), .A2(n14328), .ZN(n14632) );
  NAND2_X1 U14678 ( .A1(n14636), .A2(n14637), .ZN(n14328) );
  NAND2_X1 U14679 ( .A1(n14346), .A2(n14638), .ZN(n14637) );
  NAND2_X1 U14680 ( .A1(n14348), .A2(n14347), .ZN(n14638) );
  NOR2_X1 U14681 ( .A1(n14110), .A2(n7337), .ZN(n14346) );
  OR2_X1 U14682 ( .A1(n14347), .A2(n14348), .ZN(n14636) );
  AND2_X1 U14683 ( .A1(n14639), .A2(n14640), .ZN(n14348) );
  NAND2_X1 U14684 ( .A1(n14641), .A2(b_1_), .ZN(n14640) );
  NOR2_X1 U14685 ( .A1(n14642), .A2(n7817), .ZN(n14641) );
  NOR2_X1 U14686 ( .A1(n7816), .A2(n14343), .ZN(n14642) );
  NAND2_X1 U14687 ( .A1(n14643), .A2(b_2_), .ZN(n14639) );
  NOR2_X1 U14688 ( .A1(n14644), .A2(n8052), .ZN(n14643) );
  NOR2_X1 U14689 ( .A1(n7810), .A2(n14645), .ZN(n14644) );
  NAND2_X1 U14690 ( .A1(n14646), .A2(b_2_), .ZN(n14347) );
  NOR2_X1 U14691 ( .A1(n8055), .A2(n14110), .ZN(n14646) );
  XOR2_X1 U14692 ( .A(n14647), .B(n14648), .Z(n14326) );
  NOR2_X1 U14693 ( .A1(n7337), .A2(n14343), .ZN(n14648) );
  XOR2_X1 U14694 ( .A(n14649), .B(n14650), .Z(n14647) );
  XNOR2_X1 U14695 ( .A(n14651), .B(n14652), .ZN(n14358) );
  NAND2_X1 U14696 ( .A1(n14653), .A2(n14654), .ZN(n14651) );
  XNOR2_X1 U14697 ( .A(n14655), .B(n14656), .ZN(n14366) );
  XOR2_X1 U14698 ( .A(n14657), .B(n14658), .Z(n14656) );
  NAND2_X1 U14699 ( .A1(b_2_), .A2(a_23_), .ZN(n14658) );
  XOR2_X1 U14700 ( .A(n14659), .B(n14660), .Z(n14374) );
  XOR2_X1 U14701 ( .A(n14661), .B(n14662), .Z(n14659) );
  NOR2_X1 U14702 ( .A1(n7760), .A2(n14343), .ZN(n14662) );
  XOR2_X1 U14703 ( .A(n14663), .B(n14664), .Z(n14382) );
  XOR2_X1 U14704 ( .A(n14665), .B(n14666), .Z(n14663) );
  NOR2_X1 U14705 ( .A1(n14343), .A2(n7750), .ZN(n14666) );
  XNOR2_X1 U14706 ( .A(n14667), .B(n14668), .ZN(n14390) );
  XNOR2_X1 U14707 ( .A(n14669), .B(n14670), .ZN(n14667) );
  XNOR2_X1 U14708 ( .A(n14671), .B(n14672), .ZN(n14398) );
  XNOR2_X1 U14709 ( .A(n14673), .B(n14674), .ZN(n14671) );
  XNOR2_X1 U14710 ( .A(n14675), .B(n14676), .ZN(n14406) );
  XNOR2_X1 U14711 ( .A(n14677), .B(n14678), .ZN(n14675) );
  XNOR2_X1 U14712 ( .A(n14679), .B(n14680), .ZN(n14414) );
  XNOR2_X1 U14713 ( .A(n14681), .B(n14682), .ZN(n14679) );
  XNOR2_X1 U14714 ( .A(n14683), .B(n14684), .ZN(n14422) );
  XNOR2_X1 U14715 ( .A(n14685), .B(n14686), .ZN(n14683) );
  XNOR2_X1 U14716 ( .A(n14687), .B(n14688), .ZN(n14430) );
  XNOR2_X1 U14717 ( .A(n14689), .B(n14690), .ZN(n14687) );
  XNOR2_X1 U14718 ( .A(n14691), .B(n14692), .ZN(n14438) );
  XNOR2_X1 U14719 ( .A(n14693), .B(n14694), .ZN(n14691) );
  XNOR2_X1 U14720 ( .A(n14695), .B(n14696), .ZN(n14446) );
  XNOR2_X1 U14721 ( .A(n14697), .B(n14698), .ZN(n14695) );
  XOR2_X1 U14722 ( .A(n14699), .B(n14700), .Z(n14454) );
  XOR2_X1 U14723 ( .A(n14701), .B(n14702), .Z(n14699) );
  XOR2_X1 U14724 ( .A(n14221), .B(n14222), .Z(n14461) );
  XOR2_X1 U14725 ( .A(n14703), .B(n14704), .Z(n14221) );
  OR2_X1 U14726 ( .A1(n14705), .A2(n14706), .ZN(n14460) );
  NOR2_X1 U14727 ( .A1(n14459), .A2(n14458), .ZN(n14706) );
  NAND2_X1 U14728 ( .A1(n14707), .A2(n14708), .ZN(n7532) );
  XOR2_X1 U14729 ( .A(n14709), .B(n14710), .Z(n14707) );
  NOR2_X1 U14730 ( .A1(n7531), .A2(n14711), .ZN(n7573) );
  AND2_X1 U14731 ( .A1(n14712), .A2(n14705), .ZN(n7531) );
  INV_X1 U14732 ( .A(n14708), .ZN(n14705) );
  NAND2_X1 U14733 ( .A1(n14459), .A2(n14458), .ZN(n14708) );
  NAND2_X1 U14734 ( .A1(n14713), .A2(n14714), .ZN(n14458) );
  NAND2_X1 U14735 ( .A1(n14703), .A2(n14715), .ZN(n14714) );
  OR2_X1 U14736 ( .A1(n14704), .A2(n14222), .ZN(n14715) );
  NOR2_X1 U14737 ( .A1(n14343), .A2(n7478), .ZN(n14703) );
  NAND2_X1 U14738 ( .A1(n14222), .A2(n14704), .ZN(n14713) );
  NAND2_X1 U14739 ( .A1(n14716), .A2(n14717), .ZN(n14704) );
  NAND2_X1 U14740 ( .A1(n14702), .A2(n14718), .ZN(n14717) );
  OR2_X1 U14741 ( .A1(n14701), .A2(n14700), .ZN(n14718) );
  NOR2_X1 U14742 ( .A1(n7669), .A2(n14343), .ZN(n14702) );
  NAND2_X1 U14743 ( .A1(n14700), .A2(n14701), .ZN(n14716) );
  NAND2_X1 U14744 ( .A1(n14719), .A2(n14720), .ZN(n14701) );
  NAND2_X1 U14745 ( .A1(n14471), .A2(n14721), .ZN(n14720) );
  NAND2_X1 U14746 ( .A1(n14472), .A2(n14470), .ZN(n14721) );
  OR2_X1 U14747 ( .A1(n14470), .A2(n14472), .ZN(n14719) );
  AND2_X1 U14748 ( .A1(n14722), .A2(n14723), .ZN(n14472) );
  NAND2_X1 U14749 ( .A1(n14698), .A2(n14724), .ZN(n14723) );
  NAND2_X1 U14750 ( .A1(n14697), .A2(n14696), .ZN(n14724) );
  NOR2_X1 U14751 ( .A1(n7464), .A2(n14343), .ZN(n14698) );
  OR2_X1 U14752 ( .A1(n14696), .A2(n14697), .ZN(n14722) );
  AND2_X1 U14753 ( .A1(n14482), .A2(n14725), .ZN(n14697) );
  NAND2_X1 U14754 ( .A1(n14481), .A2(n14483), .ZN(n14725) );
  NAND2_X1 U14755 ( .A1(n14726), .A2(n14727), .ZN(n14483) );
  NAND2_X1 U14756 ( .A1(a_4_), .A2(b_2_), .ZN(n14727) );
  INV_X1 U14757 ( .A(n14728), .ZN(n14726) );
  XOR2_X1 U14758 ( .A(n14729), .B(n14730), .Z(n14481) );
  NOR2_X1 U14759 ( .A1(n14645), .A2(n7455), .ZN(n14730) );
  XOR2_X1 U14760 ( .A(n14731), .B(n14732), .Z(n14729) );
  NAND2_X1 U14761 ( .A1(a_4_), .A2(n14728), .ZN(n14482) );
  NAND2_X1 U14762 ( .A1(n14733), .A2(n14734), .ZN(n14728) );
  NAND2_X1 U14763 ( .A1(n14694), .A2(n14735), .ZN(n14734) );
  NAND2_X1 U14764 ( .A1(n14693), .A2(n14692), .ZN(n14735) );
  NOR2_X1 U14765 ( .A1(n7455), .A2(n14343), .ZN(n14694) );
  OR2_X1 U14766 ( .A1(n14692), .A2(n14693), .ZN(n14733) );
  AND2_X1 U14767 ( .A1(n14494), .A2(n14736), .ZN(n14693) );
  NAND2_X1 U14768 ( .A1(n14493), .A2(n14495), .ZN(n14736) );
  NAND2_X1 U14769 ( .A1(n14737), .A2(n14738), .ZN(n14495) );
  NAND2_X1 U14770 ( .A1(a_6_), .A2(b_2_), .ZN(n14738) );
  INV_X1 U14771 ( .A(n14739), .ZN(n14737) );
  XOR2_X1 U14772 ( .A(n14740), .B(n14741), .Z(n14493) );
  NOR2_X1 U14773 ( .A1(n14645), .A2(n7445), .ZN(n14741) );
  XOR2_X1 U14774 ( .A(n14742), .B(n14743), .Z(n14740) );
  NAND2_X1 U14775 ( .A1(a_6_), .A2(n14739), .ZN(n14494) );
  NAND2_X1 U14776 ( .A1(n14744), .A2(n14745), .ZN(n14739) );
  NAND2_X1 U14777 ( .A1(n14690), .A2(n14746), .ZN(n14745) );
  NAND2_X1 U14778 ( .A1(n14689), .A2(n14688), .ZN(n14746) );
  NOR2_X1 U14779 ( .A1(n7445), .A2(n14343), .ZN(n14690) );
  OR2_X1 U14780 ( .A1(n14688), .A2(n14689), .ZN(n14744) );
  AND2_X1 U14781 ( .A1(n14506), .A2(n14747), .ZN(n14689) );
  NAND2_X1 U14782 ( .A1(n14505), .A2(n14507), .ZN(n14747) );
  NAND2_X1 U14783 ( .A1(n14748), .A2(n14749), .ZN(n14507) );
  NAND2_X1 U14784 ( .A1(a_8_), .A2(b_2_), .ZN(n14749) );
  INV_X1 U14785 ( .A(n14750), .ZN(n14748) );
  XOR2_X1 U14786 ( .A(n14751), .B(n14752), .Z(n14505) );
  NOR2_X1 U14787 ( .A1(n14645), .A2(n7704), .ZN(n14752) );
  XOR2_X1 U14788 ( .A(n14753), .B(n14754), .Z(n14751) );
  NAND2_X1 U14789 ( .A1(a_8_), .A2(n14750), .ZN(n14506) );
  NAND2_X1 U14790 ( .A1(n14755), .A2(n14756), .ZN(n14750) );
  NAND2_X1 U14791 ( .A1(n14686), .A2(n14757), .ZN(n14756) );
  NAND2_X1 U14792 ( .A1(n14685), .A2(n14684), .ZN(n14757) );
  NOR2_X1 U14793 ( .A1(n7704), .A2(n14343), .ZN(n14686) );
  OR2_X1 U14794 ( .A1(n14684), .A2(n14685), .ZN(n14755) );
  AND2_X1 U14795 ( .A1(n14518), .A2(n14758), .ZN(n14685) );
  NAND2_X1 U14796 ( .A1(n14517), .A2(n14519), .ZN(n14758) );
  NAND2_X1 U14797 ( .A1(n14759), .A2(n14760), .ZN(n14519) );
  NAND2_X1 U14798 ( .A1(a_10_), .A2(b_2_), .ZN(n14760) );
  INV_X1 U14799 ( .A(n14761), .ZN(n14759) );
  XOR2_X1 U14800 ( .A(n14762), .B(n14763), .Z(n14517) );
  NOR2_X1 U14801 ( .A1(n7424), .A2(n14645), .ZN(n14763) );
  XOR2_X1 U14802 ( .A(n14764), .B(n14765), .Z(n14762) );
  NAND2_X1 U14803 ( .A1(a_10_), .A2(n14761), .ZN(n14518) );
  NAND2_X1 U14804 ( .A1(n14766), .A2(n14767), .ZN(n14761) );
  NAND2_X1 U14805 ( .A1(n14682), .A2(n14768), .ZN(n14767) );
  NAND2_X1 U14806 ( .A1(n14681), .A2(n14680), .ZN(n14768) );
  NOR2_X1 U14807 ( .A1(n14343), .A2(n7424), .ZN(n14682) );
  OR2_X1 U14808 ( .A1(n14680), .A2(n14681), .ZN(n14766) );
  AND2_X1 U14809 ( .A1(n14530), .A2(n14769), .ZN(n14681) );
  NAND2_X1 U14810 ( .A1(n14529), .A2(n14531), .ZN(n14769) );
  NAND2_X1 U14811 ( .A1(n14770), .A2(n14771), .ZN(n14531) );
  NAND2_X1 U14812 ( .A1(a_12_), .A2(b_2_), .ZN(n14771) );
  INV_X1 U14813 ( .A(n14772), .ZN(n14770) );
  XOR2_X1 U14814 ( .A(n14773), .B(n14774), .Z(n14529) );
  NOR2_X1 U14815 ( .A1(n14645), .A2(n7415), .ZN(n14774) );
  XOR2_X1 U14816 ( .A(n14775), .B(n14776), .Z(n14773) );
  NAND2_X1 U14817 ( .A1(a_12_), .A2(n14772), .ZN(n14530) );
  NAND2_X1 U14818 ( .A1(n14777), .A2(n14778), .ZN(n14772) );
  NAND2_X1 U14819 ( .A1(n14678), .A2(n14779), .ZN(n14778) );
  NAND2_X1 U14820 ( .A1(n14677), .A2(n14676), .ZN(n14779) );
  NOR2_X1 U14821 ( .A1(n7415), .A2(n14343), .ZN(n14678) );
  OR2_X1 U14822 ( .A1(n14676), .A2(n14677), .ZN(n14777) );
  AND2_X1 U14823 ( .A1(n14542), .A2(n14780), .ZN(n14677) );
  NAND2_X1 U14824 ( .A1(n14541), .A2(n14543), .ZN(n14780) );
  NAND2_X1 U14825 ( .A1(n14781), .A2(n14782), .ZN(n14543) );
  NAND2_X1 U14826 ( .A1(a_14_), .A2(b_2_), .ZN(n14782) );
  INV_X1 U14827 ( .A(n14783), .ZN(n14781) );
  XOR2_X1 U14828 ( .A(n14784), .B(n14785), .Z(n14541) );
  NOR2_X1 U14829 ( .A1(n14645), .A2(n7406), .ZN(n14785) );
  XOR2_X1 U14830 ( .A(n14786), .B(n14787), .Z(n14784) );
  NAND2_X1 U14831 ( .A1(a_14_), .A2(n14783), .ZN(n14542) );
  NAND2_X1 U14832 ( .A1(n14788), .A2(n14789), .ZN(n14783) );
  NAND2_X1 U14833 ( .A1(n14674), .A2(n14790), .ZN(n14789) );
  NAND2_X1 U14834 ( .A1(n14673), .A2(n14672), .ZN(n14790) );
  NOR2_X1 U14835 ( .A1(n7406), .A2(n14343), .ZN(n14674) );
  OR2_X1 U14836 ( .A1(n14672), .A2(n14673), .ZN(n14788) );
  AND2_X1 U14837 ( .A1(n14554), .A2(n14791), .ZN(n14673) );
  NAND2_X1 U14838 ( .A1(n14553), .A2(n14555), .ZN(n14791) );
  NAND2_X1 U14839 ( .A1(n14792), .A2(n14793), .ZN(n14555) );
  NAND2_X1 U14840 ( .A1(a_16_), .A2(b_2_), .ZN(n14793) );
  INV_X1 U14841 ( .A(n14794), .ZN(n14792) );
  XOR2_X1 U14842 ( .A(n14795), .B(n14796), .Z(n14553) );
  NOR2_X1 U14843 ( .A1(n14645), .A2(n7397), .ZN(n14796) );
  XOR2_X1 U14844 ( .A(n14797), .B(n14798), .Z(n14795) );
  NAND2_X1 U14845 ( .A1(a_16_), .A2(n14794), .ZN(n14554) );
  NAND2_X1 U14846 ( .A1(n14799), .A2(n14800), .ZN(n14794) );
  NAND2_X1 U14847 ( .A1(n14670), .A2(n14801), .ZN(n14800) );
  NAND2_X1 U14848 ( .A1(n14669), .A2(n14668), .ZN(n14801) );
  NOR2_X1 U14849 ( .A1(n7397), .A2(n14343), .ZN(n14670) );
  OR2_X1 U14850 ( .A1(n14668), .A2(n14669), .ZN(n14799) );
  AND2_X1 U14851 ( .A1(n14802), .A2(n14803), .ZN(n14669) );
  NAND2_X1 U14852 ( .A1(n14567), .A2(n14804), .ZN(n14803) );
  NAND2_X1 U14853 ( .A1(n14566), .A2(n14565), .ZN(n14804) );
  NOR2_X1 U14854 ( .A1(n7745), .A2(n14343), .ZN(n14567) );
  OR2_X1 U14855 ( .A1(n14565), .A2(n14566), .ZN(n14802) );
  AND2_X1 U14856 ( .A1(n14805), .A2(n14806), .ZN(n14566) );
  NAND2_X1 U14857 ( .A1(n14807), .A2(a_19_), .ZN(n14806) );
  NOR2_X1 U14858 ( .A1(n14808), .A2(n14343), .ZN(n14807) );
  NOR2_X1 U14859 ( .A1(n14664), .A2(n14665), .ZN(n14808) );
  NAND2_X1 U14860 ( .A1(n14664), .A2(n14665), .ZN(n14805) );
  NAND2_X1 U14861 ( .A1(n14809), .A2(n14810), .ZN(n14665) );
  NAND2_X1 U14862 ( .A1(n14579), .A2(n14811), .ZN(n14810) );
  NAND2_X1 U14863 ( .A1(n14578), .A2(n14577), .ZN(n14811) );
  NOR2_X1 U14864 ( .A1(n14343), .A2(n7755), .ZN(n14579) );
  OR2_X1 U14865 ( .A1(n14577), .A2(n14578), .ZN(n14809) );
  AND2_X1 U14866 ( .A1(n14812), .A2(n14813), .ZN(n14578) );
  NAND2_X1 U14867 ( .A1(n14814), .A2(b_2_), .ZN(n14813) );
  NOR2_X1 U14868 ( .A1(n14815), .A2(n7760), .ZN(n14814) );
  NOR2_X1 U14869 ( .A1(n14660), .A2(n14661), .ZN(n14815) );
  NAND2_X1 U14870 ( .A1(n14660), .A2(n14661), .ZN(n14812) );
  NAND2_X1 U14871 ( .A1(n14816), .A2(n14817), .ZN(n14661) );
  NAND2_X1 U14872 ( .A1(n14591), .A2(n14818), .ZN(n14817) );
  OR2_X1 U14873 ( .A1(n14590), .A2(n14588), .ZN(n14818) );
  NOR2_X1 U14874 ( .A1(n7765), .A2(n14343), .ZN(n14591) );
  NAND2_X1 U14875 ( .A1(n14588), .A2(n14590), .ZN(n14816) );
  NAND2_X1 U14876 ( .A1(n14819), .A2(n14820), .ZN(n14590) );
  NAND2_X1 U14877 ( .A1(n14821), .A2(b_2_), .ZN(n14820) );
  NOR2_X1 U14878 ( .A1(n14822), .A2(n8014), .ZN(n14821) );
  NOR2_X1 U14879 ( .A1(n14655), .A2(n14657), .ZN(n14822) );
  NAND2_X1 U14880 ( .A1(n14655), .A2(n14657), .ZN(n14819) );
  NAND2_X1 U14881 ( .A1(n14823), .A2(n14824), .ZN(n14657) );
  NAND2_X1 U14882 ( .A1(n14603), .A2(n14825), .ZN(n14824) );
  OR2_X1 U14883 ( .A1(n14602), .A2(n14600), .ZN(n14825) );
  NOR2_X1 U14884 ( .A1(n14343), .A2(n7774), .ZN(n14603) );
  NAND2_X1 U14885 ( .A1(n14600), .A2(n14602), .ZN(n14823) );
  NAND2_X1 U14886 ( .A1(n14653), .A2(n14826), .ZN(n14602) );
  NAND2_X1 U14887 ( .A1(n14652), .A2(n14654), .ZN(n14826) );
  NAND2_X1 U14888 ( .A1(n14827), .A2(n14828), .ZN(n14654) );
  NAND2_X1 U14889 ( .A1(b_2_), .A2(a_25_), .ZN(n14828) );
  INV_X1 U14890 ( .A(n14829), .ZN(n14827) );
  XOR2_X1 U14891 ( .A(n14830), .B(n14831), .Z(n14652) );
  NOR2_X1 U14892 ( .A1(n14832), .A2(n14833), .ZN(n14831) );
  INV_X1 U14893 ( .A(n14834), .ZN(n14833) );
  NOR2_X1 U14894 ( .A1(n14835), .A2(n14836), .ZN(n14832) );
  NAND2_X1 U14895 ( .A1(a_25_), .A2(n14829), .ZN(n14653) );
  NAND2_X1 U14896 ( .A1(n14837), .A2(n14838), .ZN(n14829) );
  NAND2_X1 U14897 ( .A1(n14839), .A2(b_2_), .ZN(n14838) );
  NOR2_X1 U14898 ( .A1(n14840), .A2(n7356), .ZN(n14839) );
  NOR2_X1 U14899 ( .A1(n14612), .A2(n14614), .ZN(n14840) );
  NAND2_X1 U14900 ( .A1(n14612), .A2(n14614), .ZN(n14837) );
  NAND2_X1 U14901 ( .A1(n14841), .A2(n14842), .ZN(n14614) );
  NAND2_X1 U14902 ( .A1(n14622), .A2(n14843), .ZN(n14842) );
  NAND2_X1 U14903 ( .A1(n14623), .A2(n14621), .ZN(n14843) );
  NOR2_X1 U14904 ( .A1(n14343), .A2(n14844), .ZN(n14622) );
  OR2_X1 U14905 ( .A1(n14621), .A2(n14623), .ZN(n14841) );
  AND2_X1 U14906 ( .A1(n14845), .A2(n14846), .ZN(n14623) );
  NAND2_X1 U14907 ( .A1(n14847), .A2(b_2_), .ZN(n14846) );
  NOR2_X1 U14908 ( .A1(n14848), .A2(n7803), .ZN(n14847) );
  NOR2_X1 U14909 ( .A1(n14631), .A2(n14629), .ZN(n14848) );
  NAND2_X1 U14910 ( .A1(n14629), .A2(n14631), .ZN(n14845) );
  NAND2_X1 U14911 ( .A1(n14849), .A2(n14850), .ZN(n14631) );
  NAND2_X1 U14912 ( .A1(n14851), .A2(b_2_), .ZN(n14850) );
  NOR2_X1 U14913 ( .A1(n14852), .A2(n7337), .ZN(n14851) );
  NOR2_X1 U14914 ( .A1(n14649), .A2(n14650), .ZN(n14852) );
  NAND2_X1 U14915 ( .A1(n14649), .A2(n14650), .ZN(n14849) );
  NAND2_X1 U14916 ( .A1(n14853), .A2(n14854), .ZN(n14650) );
  NAND2_X1 U14917 ( .A1(n14855), .A2(b_0_), .ZN(n14854) );
  NOR2_X1 U14918 ( .A1(n14856), .A2(n7817), .ZN(n14855) );
  NOR2_X1 U14919 ( .A1(n7816), .A2(n14645), .ZN(n14856) );
  NAND2_X1 U14920 ( .A1(a_31_), .A2(n8052), .ZN(n7328) );
  NAND2_X1 U14921 ( .A1(n14857), .A2(b_1_), .ZN(n14853) );
  NOR2_X1 U14922 ( .A1(n14858), .A2(n8052), .ZN(n14857) );
  NOR2_X1 U14923 ( .A1(n7810), .A2(n14859), .ZN(n14858) );
  NAND2_X1 U14924 ( .A1(a_30_), .A2(n7817), .ZN(n7332) );
  AND2_X1 U14925 ( .A1(n14860), .A2(b_1_), .ZN(n14649) );
  NOR2_X1 U14926 ( .A1(n8055), .A2(n14343), .ZN(n14860) );
  XNOR2_X1 U14927 ( .A(n14861), .B(n14862), .ZN(n14629) );
  XNOR2_X1 U14928 ( .A(n14863), .B(n14864), .ZN(n14862) );
  NAND2_X1 U14929 ( .A1(b_0_), .A2(a_30_), .ZN(n14861) );
  XNOR2_X1 U14930 ( .A(n14865), .B(n14866), .ZN(n14621) );
  NOR2_X1 U14931 ( .A1(n7337), .A2(n14859), .ZN(n14866) );
  XOR2_X1 U14932 ( .A(n14867), .B(n14868), .Z(n14865) );
  XOR2_X1 U14933 ( .A(n14869), .B(n14870), .Z(n14612) );
  NOR2_X1 U14934 ( .A1(n7803), .A2(n14859), .ZN(n14870) );
  XOR2_X1 U14935 ( .A(n14871), .B(n14872), .Z(n14869) );
  XOR2_X1 U14936 ( .A(n14873), .B(n14874), .Z(n14600) );
  NOR2_X1 U14937 ( .A1(n7356), .A2(n14859), .ZN(n14874) );
  XOR2_X1 U14938 ( .A(n14875), .B(n14876), .Z(n14873) );
  XOR2_X1 U14939 ( .A(n14877), .B(n14878), .Z(n14655) );
  NOR2_X1 U14940 ( .A1(n14879), .A2(n14880), .ZN(n14878) );
  INV_X1 U14941 ( .A(n14881), .ZN(n14880) );
  NOR2_X1 U14942 ( .A1(n14882), .A2(n14883), .ZN(n14879) );
  XOR2_X1 U14943 ( .A(n14884), .B(n14885), .Z(n14588) );
  NOR2_X1 U14944 ( .A1(n7774), .A2(n14859), .ZN(n14885) );
  XOR2_X1 U14945 ( .A(n14886), .B(n14887), .Z(n14884) );
  XOR2_X1 U14946 ( .A(n14888), .B(n14889), .Z(n14660) );
  NOR2_X1 U14947 ( .A1(n14890), .A2(n14891), .ZN(n14889) );
  INV_X1 U14948 ( .A(n14892), .ZN(n14891) );
  NOR2_X1 U14949 ( .A1(n14893), .A2(n14894), .ZN(n14890) );
  XNOR2_X1 U14950 ( .A(n14895), .B(n14896), .ZN(n14577) );
  NOR2_X1 U14951 ( .A1(n7765), .A2(n14859), .ZN(n14896) );
  XOR2_X1 U14952 ( .A(n14897), .B(n14898), .Z(n14895) );
  XOR2_X1 U14953 ( .A(n14899), .B(n14900), .Z(n14664) );
  NOR2_X1 U14954 ( .A1(n14901), .A2(n14902), .ZN(n14900) );
  INV_X1 U14955 ( .A(n14903), .ZN(n14902) );
  NOR2_X1 U14956 ( .A1(n14904), .A2(n14905), .ZN(n14901) );
  XNOR2_X1 U14957 ( .A(n14906), .B(n14907), .ZN(n14565) );
  NOR2_X1 U14958 ( .A1(n7755), .A2(n14859), .ZN(n14907) );
  XOR2_X1 U14959 ( .A(n14908), .B(n14909), .Z(n14906) );
  XNOR2_X1 U14960 ( .A(n14910), .B(n14911), .ZN(n14668) );
  NOR2_X1 U14961 ( .A1(n14912), .A2(n14913), .ZN(n14911) );
  INV_X1 U14962 ( .A(n14914), .ZN(n14913) );
  NOR2_X1 U14963 ( .A1(n14915), .A2(n14916), .ZN(n14912) );
  XNOR2_X1 U14964 ( .A(n14917), .B(n14918), .ZN(n14672) );
  NOR2_X1 U14965 ( .A1(n14919), .A2(n14920), .ZN(n14918) );
  INV_X1 U14966 ( .A(n14921), .ZN(n14920) );
  NOR2_X1 U14967 ( .A1(n14922), .A2(n14923), .ZN(n14919) );
  XNOR2_X1 U14968 ( .A(n14924), .B(n14925), .ZN(n14676) );
  NOR2_X1 U14969 ( .A1(n14926), .A2(n14927), .ZN(n14925) );
  INV_X1 U14970 ( .A(n14928), .ZN(n14927) );
  NOR2_X1 U14971 ( .A1(n14929), .A2(n14930), .ZN(n14926) );
  XNOR2_X1 U14972 ( .A(n14931), .B(n14932), .ZN(n14680) );
  NOR2_X1 U14973 ( .A1(n14933), .A2(n14934), .ZN(n14932) );
  INV_X1 U14974 ( .A(n14935), .ZN(n14934) );
  NOR2_X1 U14975 ( .A1(n14936), .A2(n14937), .ZN(n14933) );
  XNOR2_X1 U14976 ( .A(n14938), .B(n14939), .ZN(n14684) );
  NOR2_X1 U14977 ( .A1(n14940), .A2(n14941), .ZN(n14939) );
  INV_X1 U14978 ( .A(n14942), .ZN(n14941) );
  NOR2_X1 U14979 ( .A1(n14943), .A2(n14944), .ZN(n14940) );
  XNOR2_X1 U14980 ( .A(n14945), .B(n14946), .ZN(n14688) );
  NOR2_X1 U14981 ( .A1(n14947), .A2(n14948), .ZN(n14946) );
  INV_X1 U14982 ( .A(n14949), .ZN(n14948) );
  NOR2_X1 U14983 ( .A1(n14950), .A2(n14951), .ZN(n14947) );
  XNOR2_X1 U14984 ( .A(n14952), .B(n14953), .ZN(n14692) );
  NOR2_X1 U14985 ( .A1(n14954), .A2(n14955), .ZN(n14953) );
  INV_X1 U14986 ( .A(n14956), .ZN(n14955) );
  NOR2_X1 U14987 ( .A1(n14957), .A2(n14958), .ZN(n14954) );
  XNOR2_X1 U14988 ( .A(n14959), .B(n14960), .ZN(n14696) );
  NOR2_X1 U14989 ( .A1(n14961), .A2(n14962), .ZN(n14960) );
  INV_X1 U14990 ( .A(n14963), .ZN(n14962) );
  NOR2_X1 U14991 ( .A1(n14964), .A2(n14965), .ZN(n14961) );
  XNOR2_X1 U14992 ( .A(n14966), .B(n14967), .ZN(n14470) );
  NOR2_X1 U14993 ( .A1(n14645), .A2(n7464), .ZN(n14967) );
  XOR2_X1 U14994 ( .A(n14968), .B(n14969), .Z(n14966) );
  XOR2_X1 U14995 ( .A(n14970), .B(n14971), .Z(n14700) );
  NOR2_X1 U14996 ( .A1(n14972), .A2(n14973), .ZN(n14971) );
  INV_X1 U14997 ( .A(n14974), .ZN(n14973) );
  NOR2_X1 U14998 ( .A1(n14975), .A2(n14976), .ZN(n14972) );
  XOR2_X1 U14999 ( .A(n14977), .B(n14978), .Z(n14222) );
  NOR2_X1 U15000 ( .A1(n14859), .A2(n7469), .ZN(n14978) );
  XOR2_X1 U15001 ( .A(n14979), .B(n14980), .Z(n14977) );
  XOR2_X1 U15002 ( .A(n14981), .B(n14982), .Z(n14459) );
  NOR2_X1 U15003 ( .A1(n14983), .A2(n14984), .ZN(n14982) );
  INV_X1 U15004 ( .A(n14985), .ZN(n14984) );
  NOR2_X1 U15005 ( .A1(n14986), .A2(n14987), .ZN(n14983) );
  NOR2_X1 U15006 ( .A1(n14711), .A2(n14709), .ZN(n14712) );
  AND2_X1 U15007 ( .A1(a_0_), .A2(n14710), .ZN(n14711) );
  NAND2_X1 U15008 ( .A1(n14985), .A2(n14988), .ZN(n14710) );
  NAND2_X1 U15009 ( .A1(n14989), .A2(n14981), .ZN(n14988) );
  NAND2_X1 U15010 ( .A1(n14990), .A2(n14991), .ZN(n14981) );
  NAND2_X1 U15011 ( .A1(n14992), .A2(a_2_), .ZN(n14991) );
  NOR2_X1 U15012 ( .A1(n14993), .A2(n14859), .ZN(n14992) );
  NOR2_X1 U15013 ( .A1(n14980), .A2(n14979), .ZN(n14993) );
  NAND2_X1 U15014 ( .A1(n14980), .A2(n14979), .ZN(n14990) );
  NAND2_X1 U15015 ( .A1(n14974), .A2(n14994), .ZN(n14979) );
  NAND2_X1 U15016 ( .A1(n14995), .A2(n14970), .ZN(n14994) );
  NAND2_X1 U15017 ( .A1(n14996), .A2(n14997), .ZN(n14970) );
  NAND2_X1 U15018 ( .A1(n14998), .A2(a_3_), .ZN(n14997) );
  NOR2_X1 U15019 ( .A1(n14999), .A2(n14645), .ZN(n14998) );
  NOR2_X1 U15020 ( .A1(n14969), .A2(n14968), .ZN(n14999) );
  NAND2_X1 U15021 ( .A1(n14969), .A2(n14968), .ZN(n14996) );
  NAND2_X1 U15022 ( .A1(n14963), .A2(n15000), .ZN(n14968) );
  NAND2_X1 U15023 ( .A1(n15001), .A2(n14959), .ZN(n15000) );
  NAND2_X1 U15024 ( .A1(n15002), .A2(n15003), .ZN(n14959) );
  NAND2_X1 U15025 ( .A1(n15004), .A2(a_5_), .ZN(n15003) );
  NOR2_X1 U15026 ( .A1(n15005), .A2(n14645), .ZN(n15004) );
  NOR2_X1 U15027 ( .A1(n14732), .A2(n14731), .ZN(n15005) );
  NAND2_X1 U15028 ( .A1(n14732), .A2(n14731), .ZN(n15002) );
  NAND2_X1 U15029 ( .A1(n14956), .A2(n15006), .ZN(n14731) );
  NAND2_X1 U15030 ( .A1(n15007), .A2(n14952), .ZN(n15006) );
  NAND2_X1 U15031 ( .A1(n15008), .A2(n15009), .ZN(n14952) );
  NAND2_X1 U15032 ( .A1(n15010), .A2(a_7_), .ZN(n15009) );
  NOR2_X1 U15033 ( .A1(n15011), .A2(n14645), .ZN(n15010) );
  NOR2_X1 U15034 ( .A1(n14743), .A2(n14742), .ZN(n15011) );
  NAND2_X1 U15035 ( .A1(n14743), .A2(n14742), .ZN(n15008) );
  NAND2_X1 U15036 ( .A1(n14949), .A2(n15012), .ZN(n14742) );
  NAND2_X1 U15037 ( .A1(n15013), .A2(n14945), .ZN(n15012) );
  NAND2_X1 U15038 ( .A1(n15014), .A2(n15015), .ZN(n14945) );
  NAND2_X1 U15039 ( .A1(n15016), .A2(a_9_), .ZN(n15015) );
  NOR2_X1 U15040 ( .A1(n15017), .A2(n14645), .ZN(n15016) );
  NOR2_X1 U15041 ( .A1(n14754), .A2(n14753), .ZN(n15017) );
  NAND2_X1 U15042 ( .A1(n14754), .A2(n14753), .ZN(n15014) );
  NAND2_X1 U15043 ( .A1(n14942), .A2(n15018), .ZN(n14753) );
  NAND2_X1 U15044 ( .A1(n15019), .A2(n14938), .ZN(n15018) );
  NAND2_X1 U15045 ( .A1(n15020), .A2(n15021), .ZN(n14938) );
  NAND2_X1 U15046 ( .A1(n15022), .A2(b_1_), .ZN(n15021) );
  NOR2_X1 U15047 ( .A1(n15023), .A2(n7424), .ZN(n15022) );
  NOR2_X1 U15048 ( .A1(n14765), .A2(n14764), .ZN(n15023) );
  NAND2_X1 U15049 ( .A1(n14765), .A2(n14764), .ZN(n15020) );
  NAND2_X1 U15050 ( .A1(n14935), .A2(n15024), .ZN(n14764) );
  NAND2_X1 U15051 ( .A1(n15025), .A2(n14931), .ZN(n15024) );
  NAND2_X1 U15052 ( .A1(n15026), .A2(n15027), .ZN(n14931) );
  NAND2_X1 U15053 ( .A1(n15028), .A2(a_13_), .ZN(n15027) );
  NOR2_X1 U15054 ( .A1(n15029), .A2(n14645), .ZN(n15028) );
  NOR2_X1 U15055 ( .A1(n14776), .A2(n14775), .ZN(n15029) );
  NAND2_X1 U15056 ( .A1(n14776), .A2(n14775), .ZN(n15026) );
  NAND2_X1 U15057 ( .A1(n14928), .A2(n15030), .ZN(n14775) );
  NAND2_X1 U15058 ( .A1(n15031), .A2(n14924), .ZN(n15030) );
  NAND2_X1 U15059 ( .A1(n15032), .A2(n15033), .ZN(n14924) );
  NAND2_X1 U15060 ( .A1(n15034), .A2(a_15_), .ZN(n15033) );
  NOR2_X1 U15061 ( .A1(n15035), .A2(n14645), .ZN(n15034) );
  NOR2_X1 U15062 ( .A1(n14787), .A2(n14786), .ZN(n15035) );
  NAND2_X1 U15063 ( .A1(n14787), .A2(n14786), .ZN(n15032) );
  NAND2_X1 U15064 ( .A1(n14921), .A2(n15036), .ZN(n14786) );
  NAND2_X1 U15065 ( .A1(n15037), .A2(n14917), .ZN(n15036) );
  NAND2_X1 U15066 ( .A1(n15038), .A2(n15039), .ZN(n14917) );
  NAND2_X1 U15067 ( .A1(n15040), .A2(a_17_), .ZN(n15039) );
  NOR2_X1 U15068 ( .A1(n15041), .A2(n14645), .ZN(n15040) );
  NOR2_X1 U15069 ( .A1(n14798), .A2(n14797), .ZN(n15041) );
  NAND2_X1 U15070 ( .A1(n14798), .A2(n14797), .ZN(n15038) );
  NAND2_X1 U15071 ( .A1(n14914), .A2(n15042), .ZN(n14797) );
  NAND2_X1 U15072 ( .A1(n15043), .A2(n14910), .ZN(n15042) );
  NAND2_X1 U15073 ( .A1(n15044), .A2(n15045), .ZN(n14910) );
  NAND2_X1 U15074 ( .A1(n15046), .A2(b_0_), .ZN(n15045) );
  NOR2_X1 U15075 ( .A1(n15047), .A2(n7755), .ZN(n15046) );
  NOR2_X1 U15076 ( .A1(n14909), .A2(n14908), .ZN(n15047) );
  NAND2_X1 U15077 ( .A1(n14909), .A2(n14908), .ZN(n15044) );
  NAND2_X1 U15078 ( .A1(n14903), .A2(n15048), .ZN(n14908) );
  NAND2_X1 U15079 ( .A1(n15049), .A2(n14899), .ZN(n15048) );
  NAND2_X1 U15080 ( .A1(n15050), .A2(n15051), .ZN(n14899) );
  NAND2_X1 U15081 ( .A1(n15052), .A2(b_0_), .ZN(n15051) );
  NOR2_X1 U15082 ( .A1(n15053), .A2(n7765), .ZN(n15052) );
  NOR2_X1 U15083 ( .A1(n14898), .A2(n14897), .ZN(n15053) );
  NAND2_X1 U15084 ( .A1(n14898), .A2(n14897), .ZN(n15050) );
  NAND2_X1 U15085 ( .A1(n14892), .A2(n15054), .ZN(n14897) );
  NAND2_X1 U15086 ( .A1(n15055), .A2(n14888), .ZN(n15054) );
  NAND2_X1 U15087 ( .A1(n15056), .A2(n15057), .ZN(n14888) );
  NAND2_X1 U15088 ( .A1(n15058), .A2(b_0_), .ZN(n15057) );
  NOR2_X1 U15089 ( .A1(n15059), .A2(n7774), .ZN(n15058) );
  NOR2_X1 U15090 ( .A1(n14887), .A2(n14886), .ZN(n15059) );
  NAND2_X1 U15091 ( .A1(n14887), .A2(n14886), .ZN(n15056) );
  NAND2_X1 U15092 ( .A1(n14881), .A2(n15060), .ZN(n14886) );
  NAND2_X1 U15093 ( .A1(n15061), .A2(n14877), .ZN(n15060) );
  NAND2_X1 U15094 ( .A1(n15062), .A2(n15063), .ZN(n14877) );
  NAND2_X1 U15095 ( .A1(n15064), .A2(b_0_), .ZN(n15063) );
  NOR2_X1 U15096 ( .A1(n15065), .A2(n7356), .ZN(n15064) );
  NOR2_X1 U15097 ( .A1(n14876), .A2(n14875), .ZN(n15065) );
  NAND2_X1 U15098 ( .A1(n14876), .A2(n14875), .ZN(n15062) );
  NAND2_X1 U15099 ( .A1(n14834), .A2(n15066), .ZN(n14875) );
  NAND2_X1 U15100 ( .A1(n15067), .A2(n14830), .ZN(n15066) );
  NAND2_X1 U15101 ( .A1(n15068), .A2(n15069), .ZN(n14830) );
  NAND2_X1 U15102 ( .A1(n15070), .A2(b_0_), .ZN(n15069) );
  NOR2_X1 U15103 ( .A1(n15071), .A2(n7803), .ZN(n15070) );
  NOR2_X1 U15104 ( .A1(n14872), .A2(n14871), .ZN(n15071) );
  NAND2_X1 U15105 ( .A1(n14872), .A2(n14871), .ZN(n15068) );
  NAND2_X1 U15106 ( .A1(n15072), .A2(n15073), .ZN(n14871) );
  NAND2_X1 U15107 ( .A1(n15074), .A2(b_0_), .ZN(n15073) );
  NOR2_X1 U15108 ( .A1(n15075), .A2(n7337), .ZN(n15074) );
  NOR2_X1 U15109 ( .A1(n14868), .A2(n14867), .ZN(n15075) );
  NAND2_X1 U15110 ( .A1(n14868), .A2(n14867), .ZN(n15072) );
  NAND2_X1 U15111 ( .A1(n14864), .A2(n15076), .ZN(n14867) );
  NAND2_X1 U15112 ( .A1(n15077), .A2(n14863), .ZN(n15076) );
  NOR2_X1 U15113 ( .A1(n14645), .A2(n7337), .ZN(n14863) );
  NOR2_X1 U15114 ( .A1(n8052), .A2(n14859), .ZN(n15077) );
  NAND2_X1 U15115 ( .A1(n15078), .A2(b_0_), .ZN(n14864) );
  NOR2_X1 U15116 ( .A1(n8055), .A2(n14645), .ZN(n15078) );
  NOR2_X1 U15117 ( .A1(n14645), .A2(n7803), .ZN(n14868) );
  NOR2_X1 U15118 ( .A1(n14645), .A2(n14844), .ZN(n14872) );
  OR2_X1 U15119 ( .A1(n14835), .A2(a_27_), .ZN(n15067) );
  NAND2_X1 U15120 ( .A1(n14836), .A2(n14835), .ZN(n14834) );
  NOR2_X1 U15121 ( .A1(n14645), .A2(n7356), .ZN(n14835) );
  NOR2_X1 U15122 ( .A1(n14844), .A2(n14859), .ZN(n14836) );
  NOR2_X1 U15123 ( .A1(n14645), .A2(n8022), .ZN(n14876) );
  OR2_X1 U15124 ( .A1(n14882), .A2(a_25_), .ZN(n15061) );
  NAND2_X1 U15125 ( .A1(n14883), .A2(n14882), .ZN(n14881) );
  NOR2_X1 U15126 ( .A1(n14645), .A2(n7774), .ZN(n14882) );
  NOR2_X1 U15127 ( .A1(n8022), .A2(n14859), .ZN(n14883) );
  NOR2_X1 U15128 ( .A1(n14645), .A2(n8014), .ZN(n14887) );
  OR2_X1 U15129 ( .A1(n14893), .A2(a_23_), .ZN(n15055) );
  NAND2_X1 U15130 ( .A1(n14894), .A2(n14893), .ZN(n14892) );
  NOR2_X1 U15131 ( .A1(n14645), .A2(n7765), .ZN(n14893) );
  NOR2_X1 U15132 ( .A1(n8014), .A2(n14859), .ZN(n14894) );
  NOR2_X1 U15133 ( .A1(n14645), .A2(n7760), .ZN(n14898) );
  OR2_X1 U15134 ( .A1(n14904), .A2(a_21_), .ZN(n15049) );
  NAND2_X1 U15135 ( .A1(n14905), .A2(n14904), .ZN(n14903) );
  NOR2_X1 U15136 ( .A1(n14645), .A2(n7755), .ZN(n14904) );
  NOR2_X1 U15137 ( .A1(n7760), .A2(n14859), .ZN(n14905) );
  NOR2_X1 U15138 ( .A1(n7750), .A2(n14645), .ZN(n14909) );
  OR2_X1 U15139 ( .A1(n14915), .A2(a_19_), .ZN(n15043) );
  NAND2_X1 U15140 ( .A1(n14916), .A2(n14915), .ZN(n14914) );
  NOR2_X1 U15141 ( .A1(n7745), .A2(n14645), .ZN(n14915) );
  NOR2_X1 U15142 ( .A1(n14859), .A2(n7750), .ZN(n14916) );
  NOR2_X1 U15143 ( .A1(n7745), .A2(n14859), .ZN(n14798) );
  OR2_X1 U15144 ( .A1(n14922), .A2(a_16_), .ZN(n15037) );
  NAND2_X1 U15145 ( .A1(n14923), .A2(n14922), .ZN(n14921) );
  NOR2_X1 U15146 ( .A1(n7397), .A2(n14859), .ZN(n14922) );
  NOR2_X1 U15147 ( .A1(n14645), .A2(n7736), .ZN(n14923) );
  NOR2_X1 U15148 ( .A1(n7736), .A2(n14859), .ZN(n14787) );
  OR2_X1 U15149 ( .A1(n14929), .A2(a_14_), .ZN(n15031) );
  NAND2_X1 U15150 ( .A1(n14930), .A2(n14929), .ZN(n14928) );
  NOR2_X1 U15151 ( .A1(n7406), .A2(n14859), .ZN(n14929) );
  NOR2_X1 U15152 ( .A1(n14645), .A2(n7727), .ZN(n14930) );
  NOR2_X1 U15153 ( .A1(n7727), .A2(n14859), .ZN(n14776) );
  OR2_X1 U15154 ( .A1(n14936), .A2(a_12_), .ZN(n15025) );
  NAND2_X1 U15155 ( .A1(n14937), .A2(n14936), .ZN(n14935) );
  NOR2_X1 U15156 ( .A1(n7415), .A2(n14859), .ZN(n14936) );
  NOR2_X1 U15157 ( .A1(n14645), .A2(n7718), .ZN(n14937) );
  NOR2_X1 U15158 ( .A1(n7718), .A2(n14859), .ZN(n14765) );
  OR2_X1 U15159 ( .A1(n14943), .A2(a_10_), .ZN(n15019) );
  NAND2_X1 U15160 ( .A1(n14944), .A2(n14943), .ZN(n14942) );
  NOR2_X1 U15161 ( .A1(n14859), .A2(n7424), .ZN(n14943) );
  NOR2_X1 U15162 ( .A1(n14645), .A2(n7709), .ZN(n14944) );
  NOR2_X1 U15163 ( .A1(n7709), .A2(n14859), .ZN(n14754) );
  OR2_X1 U15164 ( .A1(n14950), .A2(a_8_), .ZN(n15013) );
  NAND2_X1 U15165 ( .A1(n14951), .A2(n14950), .ZN(n14949) );
  NOR2_X1 U15166 ( .A1(n7704), .A2(n14859), .ZN(n14950) );
  NOR2_X1 U15167 ( .A1(n14645), .A2(n7699), .ZN(n14951) );
  NOR2_X1 U15168 ( .A1(n7699), .A2(n14859), .ZN(n14743) );
  OR2_X1 U15169 ( .A1(n14957), .A2(a_6_), .ZN(n15007) );
  NAND2_X1 U15170 ( .A1(n14958), .A2(n14957), .ZN(n14956) );
  NOR2_X1 U15171 ( .A1(n7445), .A2(n14859), .ZN(n14957) );
  NOR2_X1 U15172 ( .A1(n14645), .A2(n7450), .ZN(n14958) );
  NOR2_X1 U15173 ( .A1(n7450), .A2(n14859), .ZN(n14732) );
  OR2_X1 U15174 ( .A1(n14964), .A2(a_4_), .ZN(n15001) );
  NAND2_X1 U15175 ( .A1(n14965), .A2(n14964), .ZN(n14963) );
  NOR2_X1 U15176 ( .A1(n7455), .A2(n14859), .ZN(n14964) );
  NOR2_X1 U15177 ( .A1(n14645), .A2(n7682), .ZN(n14965) );
  NOR2_X1 U15178 ( .A1(n7682), .A2(n14859), .ZN(n14969) );
  OR2_X1 U15179 ( .A1(n14975), .A2(a_2_), .ZN(n14995) );
  NAND2_X1 U15180 ( .A1(n14976), .A2(n14975), .ZN(n14974) );
  NOR2_X1 U15181 ( .A1(n7464), .A2(n14859), .ZN(n14975) );
  NOR2_X1 U15182 ( .A1(n14645), .A2(n7469), .ZN(n14976) );
  OR2_X1 U15183 ( .A1(n14986), .A2(a_0_), .ZN(n14989) );
  NAND2_X1 U15184 ( .A1(n14987), .A2(n14986), .ZN(n14985) );
  NOR2_X1 U15185 ( .A1(n7669), .A2(n14859), .ZN(n14986) );
  NOR2_X1 U15186 ( .A1(n7478), .A2(n14645), .ZN(n14987) );
  NAND2_X1 U15187 ( .A1(n15079), .A2(n15080), .ZN(Result_add_9_) );
  NAND2_X1 U15188 ( .A1(n12788), .A2(n15081), .ZN(n15080) );
  INV_X1 U15189 ( .A(n15082), .ZN(n12788) );
  NOR2_X1 U15190 ( .A1(n15083), .A2(n15084), .ZN(n15079) );
  NOR2_X1 U15191 ( .A1(b_9_), .A2(n15085), .ZN(n15084) );
  XOR2_X1 U15192 ( .A(n7704), .B(n15081), .Z(n15085) );
  NOR2_X1 U15193 ( .A1(n12638), .A2(n15086), .ZN(n15083) );
  OR2_X1 U15194 ( .A1(n15081), .A2(a_9_), .ZN(n15086) );
  XOR2_X1 U15195 ( .A(n15087), .B(n15088), .Z(Result_add_8_) );
  AND2_X1 U15196 ( .A1(n15089), .A2(n13204), .ZN(n15088) );
  NAND2_X1 U15197 ( .A1(n15090), .A2(n15091), .ZN(Result_add_7_) );
  NAND2_X1 U15198 ( .A1(n13450), .A2(n15092), .ZN(n15091) );
  INV_X1 U15199 ( .A(n15093), .ZN(n13450) );
  NOR2_X1 U15200 ( .A1(n15094), .A2(n15095), .ZN(n15090) );
  NOR2_X1 U15201 ( .A1(b_7_), .A2(n15096), .ZN(n15095) );
  XOR2_X1 U15202 ( .A(n7445), .B(n15092), .Z(n15096) );
  NOR2_X1 U15203 ( .A1(n13127), .A2(n15097), .ZN(n15094) );
  OR2_X1 U15204 ( .A1(n15092), .A2(a_7_), .ZN(n15097) );
  XNOR2_X1 U15205 ( .A(n15098), .B(n15099), .ZN(Result_add_6_) );
  NOR2_X1 U15206 ( .A1(n15100), .A2(n13701), .ZN(n15099) );
  NAND2_X1 U15207 ( .A1(n15101), .A2(n15102), .ZN(Result_add_5_) );
  NAND2_X1 U15208 ( .A1(n13946), .A2(n15103), .ZN(n15102) );
  INV_X1 U15209 ( .A(n15104), .ZN(n13946) );
  NOR2_X1 U15210 ( .A1(n15105), .A2(n15106), .ZN(n15101) );
  NOR2_X1 U15211 ( .A1(b_5_), .A2(n15107), .ZN(n15106) );
  XOR2_X1 U15212 ( .A(n7455), .B(n15103), .Z(n15107) );
  NOR2_X1 U15213 ( .A1(n13620), .A2(n15108), .ZN(n15105) );
  NAND2_X1 U15214 ( .A1(n15109), .A2(n7455), .ZN(n15108) );
  XNOR2_X1 U15215 ( .A(n15110), .B(n15111), .ZN(Result_add_4_) );
  NOR2_X1 U15216 ( .A1(n15112), .A2(n14199), .ZN(n15111) );
  NAND2_X1 U15217 ( .A1(n15113), .A2(n15114), .ZN(Result_add_3_) );
  NAND2_X1 U15218 ( .A1(n14444), .A2(n15115), .ZN(n15114) );
  INV_X1 U15219 ( .A(n15116), .ZN(n14444) );
  NOR2_X1 U15220 ( .A1(n15117), .A2(n15118), .ZN(n15113) );
  NOR2_X1 U15221 ( .A1(b_3_), .A2(n15119), .ZN(n15118) );
  XOR2_X1 U15222 ( .A(n7464), .B(n15115), .Z(n15119) );
  NOR2_X1 U15223 ( .A1(n14110), .A2(n15120), .ZN(n15117) );
  NAND2_X1 U15224 ( .A1(n15121), .A2(n7464), .ZN(n15120) );
  XOR2_X1 U15225 ( .A(b_31_), .B(a_31_), .Z(Result_add_31_) );
  NAND2_X1 U15226 ( .A1(n15122), .A2(n15123), .ZN(Result_add_30_) );
  INV_X1 U15227 ( .A(n7338), .ZN(n15123) );
  NOR2_X1 U15228 ( .A1(n7818), .A2(n15124), .ZN(n7338) );
  NOR2_X1 U15229 ( .A1(n15125), .A2(n15126), .ZN(n15122) );
  NOR2_X1 U15230 ( .A1(n7334), .A2(n15127), .ZN(n15126) );
  NAND2_X1 U15231 ( .A1(n15124), .A2(n8052), .ZN(n15127) );
  NOR2_X1 U15232 ( .A1(b_30_), .A2(n15128), .ZN(n15125) );
  XOR2_X1 U15233 ( .A(n15124), .B(a_30_), .Z(n15128) );
  XNOR2_X1 U15234 ( .A(n15129), .B(n15130), .ZN(Result_add_2_) );
  NOR2_X1 U15235 ( .A1(n15131), .A2(n14471), .ZN(n15130) );
  NAND2_X1 U15236 ( .A1(n15132), .A2(n15133), .ZN(Result_add_29_) );
  NAND2_X1 U15237 ( .A1(n8057), .A2(n15134), .ZN(n15133) );
  INV_X1 U15238 ( .A(n15135), .ZN(n8057) );
  NOR2_X1 U15239 ( .A1(n15136), .A2(n15137), .ZN(n15132) );
  NOR2_X1 U15240 ( .A1(b_29_), .A2(n15138), .ZN(n15137) );
  XOR2_X1 U15241 ( .A(a_29_), .B(n15139), .Z(n15138) );
  NOR2_X1 U15242 ( .A1(n7814), .A2(n15140), .ZN(n15136) );
  NAND2_X1 U15243 ( .A1(n15139), .A2(n7337), .ZN(n15140) );
  INV_X1 U15244 ( .A(n15134), .ZN(n15139) );
  XNOR2_X1 U15245 ( .A(n15141), .B(n15142), .ZN(Result_add_28_) );
  NAND2_X1 U15246 ( .A1(n8278), .A2(n15143), .ZN(n15141) );
  NAND2_X1 U15247 ( .A1(n15144), .A2(n15145), .ZN(Result_add_27_) );
  NAND2_X1 U15248 ( .A1(n8513), .A2(n15146), .ZN(n15145) );
  INV_X1 U15249 ( .A(n15147), .ZN(n8513) );
  NOR2_X1 U15250 ( .A1(n15148), .A2(n15149), .ZN(n15144) );
  NOR2_X1 U15251 ( .A1(b_27_), .A2(n15150), .ZN(n15149) );
  XOR2_X1 U15252 ( .A(n14844), .B(n15146), .Z(n15150) );
  NOR2_X1 U15253 ( .A1(n8292), .A2(n15151), .ZN(n15148) );
  OR2_X1 U15254 ( .A1(n15146), .A2(a_27_), .ZN(n15151) );
  XOR2_X1 U15255 ( .A(n15152), .B(n15153), .Z(Result_add_26_) );
  AND2_X1 U15256 ( .A1(n15154), .A2(n8985), .ZN(n15153) );
  NAND2_X1 U15257 ( .A1(n15155), .A2(n15156), .ZN(Result_add_25_) );
  NAND2_X1 U15258 ( .A1(n9024), .A2(n15157), .ZN(n15156) );
  INV_X1 U15259 ( .A(n15158), .ZN(n9024) );
  NOR2_X1 U15260 ( .A1(n15159), .A2(n15160), .ZN(n15155) );
  NOR2_X1 U15261 ( .A1(b_25_), .A2(n15161), .ZN(n15160) );
  XOR2_X1 U15262 ( .A(n8022), .B(n15157), .Z(n15161) );
  NOR2_X1 U15263 ( .A1(n8775), .A2(n15162), .ZN(n15159) );
  OR2_X1 U15264 ( .A1(n15157), .A2(a_25_), .ZN(n15162) );
  XNOR2_X1 U15265 ( .A(n15163), .B(n15164), .ZN(Result_add_24_) );
  NOR2_X1 U15266 ( .A1(n15165), .A2(n9272), .ZN(n15164) );
  NAND2_X1 U15267 ( .A1(n15166), .A2(n15167), .ZN(Result_add_23_) );
  NAND2_X1 U15268 ( .A1(n9521), .A2(n15168), .ZN(n15167) );
  INV_X1 U15269 ( .A(n15169), .ZN(n9521) );
  NOR2_X1 U15270 ( .A1(n15170), .A2(n15171), .ZN(n15166) );
  NOR2_X1 U15271 ( .A1(b_23_), .A2(n15172), .ZN(n15171) );
  XOR2_X1 U15272 ( .A(n8014), .B(n15168), .Z(n15172) );
  NOR2_X1 U15273 ( .A1(n9256), .A2(n15173), .ZN(n15170) );
  NAND2_X1 U15274 ( .A1(n15174), .A2(n8014), .ZN(n15173) );
  XNOR2_X1 U15275 ( .A(n15175), .B(n15176), .ZN(Result_add_22_) );
  NOR2_X1 U15276 ( .A1(n15177), .A2(n9758), .ZN(n15176) );
  NAND2_X1 U15277 ( .A1(n15178), .A2(n15179), .ZN(Result_add_21_) );
  NAND2_X1 U15278 ( .A1(n9995), .A2(n15180), .ZN(n15179) );
  INV_X1 U15279 ( .A(n15181), .ZN(n9995) );
  NOR2_X1 U15280 ( .A1(n15182), .A2(n15183), .ZN(n15178) );
  NOR2_X1 U15281 ( .A1(b_21_), .A2(n15184), .ZN(n15183) );
  XOR2_X1 U15282 ( .A(n7760), .B(n15180), .Z(n15184) );
  NOR2_X1 U15283 ( .A1(n9734), .A2(n15185), .ZN(n15182) );
  NAND2_X1 U15284 ( .A1(n15186), .A2(n7760), .ZN(n15185) );
  XOR2_X1 U15285 ( .A(n15187), .B(n15188), .Z(Result_add_20_) );
  AND2_X1 U15286 ( .A1(n15189), .A2(n10412), .ZN(n15188) );
  NAND2_X1 U15287 ( .A1(n15190), .A2(n15191), .ZN(Result_add_1_) );
  NAND2_X1 U15288 ( .A1(n15192), .A2(n15193), .ZN(n15191) );
  OR2_X1 U15289 ( .A1(n14980), .A2(n15194), .ZN(n15192) );
  NAND2_X1 U15290 ( .A1(n15195), .A2(n15196), .ZN(n15190) );
  XOR2_X1 U15291 ( .A(b_1_), .B(a_1_), .Z(n15195) );
  NAND2_X1 U15292 ( .A1(n15197), .A2(n15198), .ZN(Result_add_19_) );
  NAND2_X1 U15293 ( .A1(n10496), .A2(n15199), .ZN(n15198) );
  INV_X1 U15294 ( .A(n15200), .ZN(n10496) );
  NOR2_X1 U15295 ( .A1(n15201), .A2(n15202), .ZN(n15197) );
  NOR2_X1 U15296 ( .A1(b_19_), .A2(n15203), .ZN(n15202) );
  XOR2_X1 U15297 ( .A(n7750), .B(n15199), .Z(n15203) );
  NOR2_X1 U15298 ( .A1(n10207), .A2(n15204), .ZN(n15201) );
  OR2_X1 U15299 ( .A1(n15199), .A2(a_19_), .ZN(n15204) );
  XNOR2_X1 U15300 ( .A(n15205), .B(n15206), .ZN(Result_add_18_) );
  NOR2_X1 U15301 ( .A1(n15207), .A2(n10733), .ZN(n15206) );
  NAND2_X1 U15302 ( .A1(n15208), .A2(n15209), .ZN(Result_add_17_) );
  NAND2_X1 U15303 ( .A1(n11005), .A2(n15210), .ZN(n15209) );
  NOR2_X1 U15304 ( .A1(n15211), .A2(n15212), .ZN(n15208) );
  NOR2_X1 U15305 ( .A1(b_17_), .A2(n15213), .ZN(n15212) );
  XOR2_X1 U15306 ( .A(n7397), .B(n15210), .Z(n15213) );
  NOR2_X1 U15307 ( .A1(n10693), .A2(n15214), .ZN(n15211) );
  NAND2_X1 U15308 ( .A1(n15215), .A2(n7397), .ZN(n15214) );
  XNOR2_X1 U15309 ( .A(n15216), .B(n15217), .ZN(Result_add_16_) );
  NOR2_X1 U15310 ( .A1(n15218), .A2(n11223), .ZN(n15217) );
  NAND2_X1 U15311 ( .A1(n15219), .A2(n15220), .ZN(Result_add_15_) );
  NAND2_X1 U15312 ( .A1(n11479), .A2(n15221), .ZN(n15220) );
  INV_X1 U15313 ( .A(n15222), .ZN(n11479) );
  NOR2_X1 U15314 ( .A1(n15223), .A2(n15224), .ZN(n15219) );
  NOR2_X1 U15315 ( .A1(b_15_), .A2(n15225), .ZN(n15224) );
  XOR2_X1 U15316 ( .A(n7406), .B(n15221), .Z(n15225) );
  NOR2_X1 U15317 ( .A1(n11175), .A2(n15226), .ZN(n15223) );
  NAND2_X1 U15318 ( .A1(n15227), .A2(n7406), .ZN(n15226) );
  XOR2_X1 U15319 ( .A(n15228), .B(n15229), .Z(Result_add_14_) );
  AND2_X1 U15320 ( .A1(n15230), .A2(n11717), .ZN(n15229) );
  NAND2_X1 U15321 ( .A1(n15231), .A2(n15232), .ZN(Result_add_13_) );
  NAND2_X1 U15322 ( .A1(n11862), .A2(n15233), .ZN(n15232) );
  INV_X1 U15323 ( .A(n15234), .ZN(n11862) );
  NOR2_X1 U15324 ( .A1(n15235), .A2(n15236), .ZN(n15231) );
  NOR2_X1 U15325 ( .A1(b_13_), .A2(n15237), .ZN(n15236) );
  XOR2_X1 U15326 ( .A(n7415), .B(n15233), .Z(n15237) );
  NOR2_X1 U15327 ( .A1(n11664), .A2(n15238), .ZN(n15235) );
  OR2_X1 U15328 ( .A1(n15233), .A2(a_13_), .ZN(n15238) );
  XOR2_X1 U15329 ( .A(n15239), .B(n15240), .Z(Result_add_12_) );
  AND2_X1 U15330 ( .A1(n15241), .A2(n12340), .ZN(n15240) );
  NAND2_X1 U15331 ( .A1(n15242), .A2(n15243), .ZN(Result_add_11_) );
  NAND2_X1 U15332 ( .A1(n12481), .A2(n15244), .ZN(n15243) );
  INV_X1 U15333 ( .A(n15245), .ZN(n12481) );
  NOR2_X1 U15334 ( .A1(n15246), .A2(n15247), .ZN(n15242) );
  NOR2_X1 U15335 ( .A1(b_11_), .A2(n15248), .ZN(n15247) );
  XOR2_X1 U15336 ( .A(n7424), .B(n15244), .Z(n15248) );
  NOR2_X1 U15337 ( .A1(n12145), .A2(n15249), .ZN(n15246) );
  OR2_X1 U15338 ( .A1(n15244), .A2(a_11_), .ZN(n15249) );
  XOR2_X1 U15339 ( .A(n15250), .B(n15251), .Z(Result_add_10_) );
  AND2_X1 U15340 ( .A1(n15252), .A2(n12800), .ZN(n15251) );
  XOR2_X1 U15341 ( .A(n15253), .B(n15254), .Z(Result_add_0_) );
  NOR2_X1 U15342 ( .A1(n15255), .A2(n15256), .ZN(n15254) );
  INV_X1 U15343 ( .A(n14709), .ZN(n15256) );
  NAND2_X1 U15344 ( .A1(b_0_), .A2(a_0_), .ZN(n14709) );
  NOR2_X1 U15345 ( .A1(b_0_), .A2(a_0_), .ZN(n15255) );
  NOR2_X1 U15346 ( .A1(n15194), .A2(n15257), .ZN(n15253) );
  NOR2_X1 U15347 ( .A1(n14980), .A2(n15193), .ZN(n15257) );
  INV_X1 U15348 ( .A(n15196), .ZN(n15193) );
  NOR2_X1 U15349 ( .A1(n14471), .A2(n15258), .ZN(n15196) );
  NOR2_X1 U15350 ( .A1(n15131), .A2(n15129), .ZN(n15258) );
  AND2_X1 U15351 ( .A1(n15116), .A2(n15259), .ZN(n15129) );
  NAND2_X1 U15352 ( .A1(n15260), .A2(n15115), .ZN(n15259) );
  INV_X1 U15353 ( .A(n15121), .ZN(n15115) );
  NOR2_X1 U15354 ( .A1(n14199), .A2(n15261), .ZN(n15121) );
  NOR2_X1 U15355 ( .A1(n15112), .A2(n15110), .ZN(n15261) );
  AND2_X1 U15356 ( .A1(n15104), .A2(n15262), .ZN(n15110) );
  NAND2_X1 U15357 ( .A1(n15263), .A2(n15103), .ZN(n15262) );
  INV_X1 U15358 ( .A(n15109), .ZN(n15103) );
  NOR2_X1 U15359 ( .A1(n13701), .A2(n15264), .ZN(n15109) );
  NOR2_X1 U15360 ( .A1(n15100), .A2(n15098), .ZN(n15264) );
  AND2_X1 U15361 ( .A1(n15093), .A2(n15265), .ZN(n15098) );
  NAND2_X1 U15362 ( .A1(n15266), .A2(n15092), .ZN(n15265) );
  NAND2_X1 U15363 ( .A1(n13204), .A2(n15267), .ZN(n15092) );
  NAND2_X1 U15364 ( .A1(n15089), .A2(n15087), .ZN(n15267) );
  NAND2_X1 U15365 ( .A1(n15082), .A2(n15268), .ZN(n15087) );
  NAND2_X1 U15366 ( .A1(n15269), .A2(n15081), .ZN(n15268) );
  NAND2_X1 U15367 ( .A1(n12800), .A2(n15270), .ZN(n15081) );
  NAND2_X1 U15368 ( .A1(n15252), .A2(n15250), .ZN(n15270) );
  NAND2_X1 U15369 ( .A1(n15245), .A2(n15271), .ZN(n15250) );
  NAND2_X1 U15370 ( .A1(n15272), .A2(n15244), .ZN(n15271) );
  NAND2_X1 U15371 ( .A1(n12340), .A2(n15273), .ZN(n15244) );
  NAND2_X1 U15372 ( .A1(n15241), .A2(n15239), .ZN(n15273) );
  NAND2_X1 U15373 ( .A1(n15234), .A2(n15274), .ZN(n15239) );
  NAND2_X1 U15374 ( .A1(n15275), .A2(n15233), .ZN(n15274) );
  NAND2_X1 U15375 ( .A1(n11717), .A2(n15276), .ZN(n15233) );
  NAND2_X1 U15376 ( .A1(n15230), .A2(n15228), .ZN(n15276) );
  NAND2_X1 U15377 ( .A1(n15222), .A2(n15277), .ZN(n15228) );
  NAND2_X1 U15378 ( .A1(n15278), .A2(n15221), .ZN(n15277) );
  INV_X1 U15379 ( .A(n15227), .ZN(n15221) );
  NOR2_X1 U15380 ( .A1(n11223), .A2(n15279), .ZN(n15227) );
  NOR2_X1 U15381 ( .A1(n15218), .A2(n15216), .ZN(n15279) );
  NOR2_X1 U15382 ( .A1(n11005), .A2(n15280), .ZN(n15216) );
  AND2_X1 U15383 ( .A1(n15281), .A2(n15210), .ZN(n15280) );
  INV_X1 U15384 ( .A(n15215), .ZN(n15210) );
  NOR2_X1 U15385 ( .A1(n10733), .A2(n15282), .ZN(n15215) );
  NOR2_X1 U15386 ( .A1(n15207), .A2(n15205), .ZN(n15282) );
  AND2_X1 U15387 ( .A1(n15200), .A2(n15283), .ZN(n15205) );
  NAND2_X1 U15388 ( .A1(n15284), .A2(n15199), .ZN(n15283) );
  NAND2_X1 U15389 ( .A1(n10412), .A2(n15285), .ZN(n15199) );
  NAND2_X1 U15390 ( .A1(n15189), .A2(n15187), .ZN(n15285) );
  NAND2_X1 U15391 ( .A1(n15181), .A2(n15286), .ZN(n15187) );
  NAND2_X1 U15392 ( .A1(n15287), .A2(n15180), .ZN(n15286) );
  INV_X1 U15393 ( .A(n15186), .ZN(n15180) );
  NOR2_X1 U15394 ( .A1(n9758), .A2(n15288), .ZN(n15186) );
  NOR2_X1 U15395 ( .A1(n15177), .A2(n15175), .ZN(n15288) );
  AND2_X1 U15396 ( .A1(n15169), .A2(n15289), .ZN(n15175) );
  NAND2_X1 U15397 ( .A1(n15290), .A2(n15168), .ZN(n15289) );
  INV_X1 U15398 ( .A(n15174), .ZN(n15168) );
  NOR2_X1 U15399 ( .A1(n9272), .A2(n15291), .ZN(n15174) );
  NOR2_X1 U15400 ( .A1(n15165), .A2(n15163), .ZN(n15291) );
  AND2_X1 U15401 ( .A1(n15158), .A2(n15292), .ZN(n15163) );
  NAND2_X1 U15402 ( .A1(n15293), .A2(n15157), .ZN(n15292) );
  NAND2_X1 U15403 ( .A1(n8985), .A2(n15294), .ZN(n15157) );
  NAND2_X1 U15404 ( .A1(n15154), .A2(n15152), .ZN(n15294) );
  NAND2_X1 U15405 ( .A1(n15147), .A2(n15295), .ZN(n15152) );
  NAND2_X1 U15406 ( .A1(n15296), .A2(n15146), .ZN(n15295) );
  NAND2_X1 U15407 ( .A1(n8278), .A2(n15297), .ZN(n15146) );
  NAND2_X1 U15408 ( .A1(n15143), .A2(n15142), .ZN(n15297) );
  NAND2_X1 U15409 ( .A1(n15135), .A2(n15298), .ZN(n15142) );
  NAND2_X1 U15410 ( .A1(n15299), .A2(n15134), .ZN(n15298) );
  NAND2_X1 U15411 ( .A1(n7818), .A2(n15300), .ZN(n15134) );
  NAND2_X1 U15412 ( .A1(Result_mul_63_), .A2(n15301), .ZN(n15300) );
  NAND2_X1 U15413 ( .A1(n7334), .A2(n8052), .ZN(n15301) );
  INV_X1 U15414 ( .A(b_30_), .ZN(n7334) );
  INV_X1 U15415 ( .A(n15124), .ZN(Result_mul_63_) );
  NAND2_X1 U15416 ( .A1(b_31_), .A2(a_31_), .ZN(n15124) );
  NAND2_X1 U15417 ( .A1(b_30_), .A2(a_30_), .ZN(n7818) );
  NAND2_X1 U15418 ( .A1(n7814), .A2(n7337), .ZN(n15299) );
  INV_X1 U15419 ( .A(b_29_), .ZN(n7814) );
  NAND2_X1 U15420 ( .A1(b_29_), .A2(a_29_), .ZN(n15135) );
  NAND2_X1 U15421 ( .A1(n8053), .A2(n7803), .ZN(n15143) );
  INV_X1 U15422 ( .A(b_28_), .ZN(n8053) );
  NAND2_X1 U15423 ( .A1(b_28_), .A2(a_28_), .ZN(n8278) );
  NAND2_X1 U15424 ( .A1(n8292), .A2(n14844), .ZN(n15296) );
  INV_X1 U15425 ( .A(a_27_), .ZN(n14844) );
  NAND2_X1 U15426 ( .A1(b_27_), .A2(a_27_), .ZN(n15147) );
  NAND2_X1 U15427 ( .A1(n8535), .A2(n7356), .ZN(n15154) );
  INV_X1 U15428 ( .A(a_26_), .ZN(n7356) );
  INV_X1 U15429 ( .A(b_26_), .ZN(n8535) );
  NAND2_X1 U15430 ( .A1(b_26_), .A2(a_26_), .ZN(n8985) );
  NAND2_X1 U15431 ( .A1(n8775), .A2(n8022), .ZN(n15293) );
  INV_X1 U15432 ( .A(b_25_), .ZN(n8775) );
  NAND2_X1 U15433 ( .A1(b_25_), .A2(a_25_), .ZN(n15158) );
  NOR2_X1 U15434 ( .A1(b_24_), .A2(a_24_), .ZN(n15165) );
  NOR2_X1 U15435 ( .A1(n9007), .A2(n7774), .ZN(n9272) );
  INV_X1 U15436 ( .A(b_24_), .ZN(n9007) );
  NAND2_X1 U15437 ( .A1(n9256), .A2(n8014), .ZN(n15290) );
  INV_X1 U15438 ( .A(b_23_), .ZN(n9256) );
  NAND2_X1 U15439 ( .A1(b_23_), .A2(a_23_), .ZN(n15169) );
  NOR2_X1 U15440 ( .A1(b_22_), .A2(a_22_), .ZN(n15177) );
  NOR2_X1 U15441 ( .A1(n9500), .A2(n7765), .ZN(n9758) );
  INV_X1 U15442 ( .A(b_22_), .ZN(n9500) );
  NAND2_X1 U15443 ( .A1(n9734), .A2(n7760), .ZN(n15287) );
  NAND2_X1 U15444 ( .A1(b_21_), .A2(a_21_), .ZN(n15181) );
  NAND2_X1 U15445 ( .A1(n9966), .A2(n7755), .ZN(n15189) );
  INV_X1 U15446 ( .A(b_20_), .ZN(n9966) );
  NAND2_X1 U15447 ( .A1(b_20_), .A2(a_20_), .ZN(n10412) );
  NAND2_X1 U15448 ( .A1(n10207), .A2(n7750), .ZN(n15284) );
  NAND2_X1 U15449 ( .A1(b_19_), .A2(a_19_), .ZN(n15200) );
  NOR2_X1 U15450 ( .A1(b_18_), .A2(a_18_), .ZN(n15207) );
  NOR2_X1 U15451 ( .A1(n10459), .A2(n7745), .ZN(n10733) );
  INV_X1 U15452 ( .A(b_18_), .ZN(n10459) );
  NAND2_X1 U15453 ( .A1(n10693), .A2(n7397), .ZN(n15281) );
  NOR2_X1 U15454 ( .A1(n10693), .A2(n7397), .ZN(n11005) );
  NOR2_X1 U15455 ( .A1(b_16_), .A2(a_16_), .ZN(n15218) );
  NOR2_X1 U15456 ( .A1(n10964), .A2(n7736), .ZN(n11223) );
  INV_X1 U15457 ( .A(b_16_), .ZN(n10964) );
  NAND2_X1 U15458 ( .A1(n11175), .A2(n7406), .ZN(n15278) );
  INV_X1 U15459 ( .A(b_15_), .ZN(n11175) );
  NAND2_X1 U15460 ( .A1(b_15_), .A2(a_15_), .ZN(n15222) );
  NAND2_X1 U15461 ( .A1(n11426), .A2(n7727), .ZN(n15230) );
  INV_X1 U15462 ( .A(b_14_), .ZN(n11426) );
  NAND2_X1 U15463 ( .A1(b_14_), .A2(a_14_), .ZN(n11717) );
  NAND2_X1 U15464 ( .A1(n11664), .A2(n7415), .ZN(n15275) );
  INV_X1 U15465 ( .A(b_13_), .ZN(n11664) );
  NAND2_X1 U15466 ( .A1(b_13_), .A2(a_13_), .ZN(n15234) );
  NAND2_X1 U15467 ( .A1(n11945), .A2(n7718), .ZN(n15241) );
  INV_X1 U15468 ( .A(b_12_), .ZN(n11945) );
  NAND2_X1 U15469 ( .A1(b_12_), .A2(a_12_), .ZN(n12340) );
  NAND2_X1 U15470 ( .A1(n12145), .A2(n7424), .ZN(n15272) );
  NAND2_X1 U15471 ( .A1(a_11_), .A2(b_11_), .ZN(n15245) );
  NAND2_X1 U15472 ( .A1(n12422), .A2(n7709), .ZN(n15252) );
  NAND2_X1 U15473 ( .A1(a_10_), .A2(b_10_), .ZN(n12800) );
  NAND2_X1 U15474 ( .A1(n12638), .A2(n7704), .ZN(n15269) );
  NAND2_X1 U15475 ( .A1(a_9_), .A2(b_9_), .ZN(n15082) );
  NAND2_X1 U15476 ( .A1(n12909), .A2(n7699), .ZN(n15089) );
  NAND2_X1 U15477 ( .A1(a_8_), .A2(b_8_), .ZN(n13204) );
  NAND2_X1 U15478 ( .A1(n13127), .A2(n7445), .ZN(n15266) );
  NAND2_X1 U15479 ( .A1(a_7_), .A2(b_7_), .ZN(n15093) );
  NOR2_X1 U15480 ( .A1(b_6_), .A2(a_6_), .ZN(n15100) );
  NOR2_X1 U15481 ( .A1(n7450), .A2(n13377), .ZN(n13701) );
  NAND2_X1 U15482 ( .A1(n13620), .A2(n7455), .ZN(n15263) );
  NAND2_X1 U15483 ( .A1(a_5_), .A2(b_5_), .ZN(n15104) );
  NOR2_X1 U15484 ( .A1(b_4_), .A2(a_4_), .ZN(n15112) );
  NOR2_X1 U15485 ( .A1(n7682), .A2(n13861), .ZN(n14199) );
  NAND2_X1 U15486 ( .A1(n14110), .A2(n7464), .ZN(n15260) );
  NAND2_X1 U15487 ( .A1(a_3_), .A2(b_3_), .ZN(n15116) );
  NOR2_X1 U15488 ( .A1(b_2_), .A2(a_2_), .ZN(n15131) );
  NOR2_X1 U15489 ( .A1(n7469), .A2(n14343), .ZN(n14471) );
  INV_X1 U15490 ( .A(b_2_), .ZN(n14343) );
  NOR2_X1 U15491 ( .A1(n7669), .A2(n14645), .ZN(n14980) );
  NOR2_X1 U15492 ( .A1(b_1_), .A2(a_1_), .ZN(n15194) );
endmodule

