module add_mul_sub_32_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, 
        a_18_, a_19_, a_20_, a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, 
        a_28_, a_29_, a_30_, a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, 
        b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, 
        b_17_, b_18_, b_19_, b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, 
        b_27_, b_28_, b_29_, b_30_, b_31_, operation_0_, operation_1_, 
        Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_, 
        Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_, 
        Result_12_, Result_13_, Result_14_, Result_15_, Result_16_, Result_17_, 
        Result_18_, Result_19_, Result_20_, Result_21_, Result_22_, Result_23_, 
        Result_24_, Result_25_, Result_26_, Result_27_, Result_28_, Result_29_, 
        Result_30_, Result_31_, Result_32_, Result_33_, Result_34_, Result_35_, 
        Result_36_, Result_37_, Result_38_, Result_39_, Result_40_, Result_41_, 
        Result_42_, Result_43_, Result_44_, Result_45_, Result_46_, Result_47_, 
        Result_48_, Result_49_, Result_50_, Result_51_, Result_52_, Result_53_, 
        Result_54_, Result_55_, Result_56_, Result_57_, Result_58_, Result_59_, 
        Result_60_, Result_61_, Result_62_, Result_63_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, a_19_, a_20_,
         a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, a_29_, a_30_,
         a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_,
         b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, b_18_, b_19_,
         b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, b_28_, b_29_,
         b_30_, b_31_, operation_0_, operation_1_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_,
         Result_32_, Result_33_, Result_34_, Result_35_, Result_36_,
         Result_37_, Result_38_, Result_39_, Result_40_, Result_41_,
         Result_42_, Result_43_, Result_44_, Result_45_, Result_46_,
         Result_47_, Result_48_, Result_49_, Result_50_, Result_51_,
         Result_52_, Result_53_, Result_54_, Result_55_, Result_56_,
         Result_57_, Result_58_, Result_59_, Result_60_, Result_61_,
         Result_62_, Result_63_;
  wire   n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626,
         n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
         n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
         n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,
         n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
         n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666,
         n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674,
         n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
         n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
         n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706,
         n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
         n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,
         n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
         n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,
         n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746,
         n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
         n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,
         n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770,
         n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778,
         n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786,
         n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794,
         n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802,
         n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810,
         n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818,
         n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826,
         n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834,
         n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842,
         n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850,
         n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858,
         n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866,
         n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874,
         n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882,
         n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890,
         n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898,
         n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906,
         n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914,
         n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922,
         n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930,
         n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938,
         n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946,
         n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954,
         n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962,
         n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970,
         n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978,
         n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986,
         n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994,
         n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002,
         n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010,
         n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
         n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,
         n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034,
         n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,
         n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050,
         n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058,
         n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066,
         n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
         n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082,
         n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,
         n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,
         n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106,
         n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114,
         n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122,
         n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130,
         n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
         n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146,
         n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154,
         n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,
         n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170,
         n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178,
         n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186,
         n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194,
         n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202,
         n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
         n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218,
         n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226,
         n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
         n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242,
         n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250,
         n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258,
         n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266,
         n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274,
         n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282,
         n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290,
         n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298,
         n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
         n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314,
         n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322,
         n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330,
         n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
         n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346,
         n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354,
         n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,
         n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370,
         n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
         n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386,
         n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394,
         n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402,
         n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
         n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,
         n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,
         n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,
         n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442,
         n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
         n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458,
         n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466,
         n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,
         n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
         n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490,
         n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
         n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
         n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
         n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
         n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538,
         n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546,
         n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
         n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562,
         n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,
         n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
         n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,
         n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
         n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602,
         n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610,
         n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618,
         n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626,
         n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634,
         n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642,
         n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650,
         n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658,
         n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
         n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674,
         n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682,
         n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690,
         n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
         n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706,
         n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714,
         n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722,
         n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730,
         n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,
         n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746,
         n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754,
         n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762,
         n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770,
         n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778,
         n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786,
         n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794,
         n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802,
         n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,
         n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818,
         n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826,
         n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834,
         n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842,
         n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850,
         n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858,
         n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866,
         n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874,
         n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,
         n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890,
         n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898,
         n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906,
         n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914,
         n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922,
         n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930,
         n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938,
         n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946,
         n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,
         n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962,
         n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970,
         n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978,
         n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986,
         n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994,
         n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002,
         n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010,
         n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018,
         n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
         n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034,
         n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042,
         n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050,
         n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058,
         n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
         n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074,
         n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082,
         n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090,
         n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
         n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106,
         n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114,
         n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122,
         n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130,
         n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,
         n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,
         n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
         n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
         n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
         n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178,
         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,
         n18187, n18188, n18189, n18190;

  INV_X2 U9088 ( .A(b_1_), .ZN(n9982) );
  INV_X2 U9089 ( .A(b_21_), .ZN(n10052) );
  INV_X2 U9090 ( .A(b_27_), .ZN(n11041) );
  INV_X2 U9091 ( .A(b_25_), .ZN(n9245) );
  INV_X2 U9092 ( .A(n18016), .ZN(n9030) );
  INV_X2 U9093 ( .A(n9064), .ZN(n9091) );
  NAND2_X2 U9094 ( .A1(n9979), .A2(n9980), .ZN(n9064) );
  INV_X1 U9095 ( .A(n10045), .ZN(n9024) );
  INV_X2 U9096 ( .A(n9024), .ZN(n9025) );
  NAND2_X4 U9097 ( .A1(operation_0_), .A2(n9979), .ZN(n9092) );
  INV_X4 U9098 ( .A(a_29_), .ZN(n9121) );
  INV_X1 U9099 ( .A(n9032), .ZN(n9026) );
  INV_X4 U9100 ( .A(n9026), .ZN(n9027) );
  INV_X1 U9101 ( .A(n9066), .ZN(n9028) );
  INV_X4 U9102 ( .A(n9028), .ZN(n9029) );
  INV_X2 U9103 ( .A(b_31_), .ZN(n9077) );
  INV_X2 U9104 ( .A(a_6_), .ZN(n10081) );
  INV_X2 U9105 ( .A(a_14_), .ZN(n10065) );
  INV_X2 U9106 ( .A(a_12_), .ZN(n10070) );
  INV_X2 U9107 ( .A(a_5_), .ZN(n10083) );
  INV_X2 U9108 ( .A(a_9_), .ZN(n10076) );
  INV_X2 U9109 ( .A(a_19_), .ZN(n9415) );
  INV_X2 U9110 ( .A(n9081), .ZN(n10486) );
  INV_X2 U9111 ( .A(a_0_), .ZN(n10093) );
  INV_X2 U9112 ( .A(a_1_), .ZN(n9983) );
  INV_X2 U9113 ( .A(a_15_), .ZN(n9534) );
  INV_X2 U9114 ( .A(b_5_), .ZN(n10082) );
  INV_X2 U9115 ( .A(b_28_), .ZN(n10786) );
  INV_X2 U9116 ( .A(b_26_), .ZN(n9217) );
  INV_X2 U9117 ( .A(b_30_), .ZN(n9080) );
  INV_X2 U9118 ( .A(b_23_), .ZN(n9302) );
  NAND2_X2 U9119 ( .A1(a_30_), .A2(n10044), .ZN(n10489) );
  INV_X2 U9120 ( .A(b_8_), .ZN(n10078) );
  INV_X2 U9121 ( .A(b_24_), .ZN(n10049) );
  INV_X2 U9122 ( .A(a_10_), .ZN(n10073) );
  INV_X2 U9123 ( .A(a_18_), .ZN(n10058) );
  INV_X2 U9124 ( .A(a_11_), .ZN(n9649) );
  INV_X2 U9125 ( .A(b_4_), .ZN(n10084) );
  INV_X2 U9126 ( .A(b_2_), .ZN(n10087) );
  INV_X2 U9127 ( .A(b_0_), .ZN(n10094) );
  INV_X2 U9128 ( .A(a_25_), .ZN(n10048) );
  INV_X2 U9129 ( .A(a_26_), .ZN(n10047) );
  INV_X2 U9130 ( .A(a_20_), .ZN(n10054) );
  INV_X2 U9131 ( .A(b_17_), .ZN(n10059) );
  INV_X2 U9132 ( .A(a_28_), .ZN(n9136) );
  INV_X2 U9133 ( .A(b_11_), .ZN(n10071) );
  INV_X2 U9134 ( .A(a_23_), .ZN(n10051) );
  NAND2_X1 U9135 ( .A1(n9030), .A2(n9031), .ZN(Result_9_) );
  NAND2_X1 U9136 ( .A1(n9027), .A2(n9033), .ZN(n9031) );
  XOR2_X1 U9137 ( .A(n9034), .B(n9035), .Z(n9033) );
  NOR2_X1 U9138 ( .A1(n9036), .A2(n9037), .ZN(n9035) );
  INV_X1 U9139 ( .A(n9038), .ZN(n9037) );
  NOR2_X1 U9140 ( .A1(n9039), .A2(n9040), .ZN(n9036) );
  NAND2_X1 U9141 ( .A1(n9030), .A2(n9041), .ZN(Result_8_) );
  NAND2_X1 U9142 ( .A1(n9027), .A2(n9042), .ZN(n9041) );
  XOR2_X1 U9143 ( .A(n9043), .B(n9044), .Z(n9042) );
  NAND2_X1 U9144 ( .A1(n9030), .A2(n9045), .ZN(Result_7_) );
  NAND2_X1 U9145 ( .A1(n9027), .A2(n9046), .ZN(n9045) );
  XOR2_X1 U9146 ( .A(n9047), .B(n9048), .Z(n9046) );
  NOR2_X1 U9147 ( .A1(n9049), .A2(n9050), .ZN(n9048) );
  INV_X1 U9148 ( .A(n9051), .ZN(n9050) );
  NOR2_X1 U9149 ( .A1(n9052), .A2(n9053), .ZN(n9049) );
  NAND2_X1 U9150 ( .A1(n9030), .A2(n9054), .ZN(Result_6_) );
  NAND2_X1 U9151 ( .A1(n9027), .A2(n9055), .ZN(n9054) );
  XOR2_X1 U9152 ( .A(n9056), .B(n9057), .Z(n9055) );
  NAND2_X1 U9153 ( .A1(n9058), .A2(n9059), .ZN(Result_63_) );
  NAND2_X1 U9154 ( .A1(n9060), .A2(n9027), .ZN(n9059) );
  NAND2_X1 U9155 ( .A1(n9061), .A2(n9062), .ZN(n9058) );
  NAND2_X1 U9156 ( .A1(n9063), .A2(n9064), .ZN(n9062) );
  NOR2_X1 U9157 ( .A1(n9065), .A2(n9029), .ZN(n9063) );
  NAND2_X1 U9158 ( .A1(n9067), .A2(n9068), .ZN(n9061) );
  NAND2_X1 U9159 ( .A1(n9069), .A2(n9070), .ZN(Result_62_) );
  NAND2_X1 U9160 ( .A1(n9027), .A2(n9071), .ZN(n9070) );
  NAND2_X1 U9161 ( .A1(n9072), .A2(n9073), .ZN(n9071) );
  NAND2_X1 U9162 ( .A1(n9074), .A2(a_30_), .ZN(n9073) );
  NOR2_X1 U9163 ( .A1(n9075), .A2(n9076), .ZN(n9072) );
  NOR2_X1 U9164 ( .A1(n9077), .A2(n9078), .ZN(n9076) );
  NOR2_X1 U9165 ( .A1(n9079), .A2(n9080), .ZN(n9075) );
  NOR2_X1 U9166 ( .A1(n9081), .A2(n9082), .ZN(n9079) );
  NOR2_X1 U9167 ( .A1(n9083), .A2(n9084), .ZN(n9069) );
  NOR2_X1 U9168 ( .A1(n9085), .A2(n9086), .ZN(n9084) );
  NOR2_X1 U9169 ( .A1(n9087), .A2(n9088), .ZN(n9085) );
  NAND2_X1 U9170 ( .A1(n9089), .A2(n9090), .ZN(n9088) );
  NAND2_X1 U9171 ( .A1(n9091), .A2(n9060), .ZN(n9090) );
  NAND2_X1 U9172 ( .A1(n9074), .A2(n9029), .ZN(n9089) );
  NOR2_X1 U9173 ( .A1(n9067), .A2(n9092), .ZN(n9087) );
  INV_X1 U9174 ( .A(n9082), .ZN(n9067) );
  NOR2_X1 U9175 ( .A1(n9093), .A2(n9094), .ZN(n9083) );
  NOR2_X1 U9176 ( .A1(n9095), .A2(n9096), .ZN(n9094) );
  NAND2_X1 U9177 ( .A1(n9097), .A2(n9098), .ZN(n9096) );
  NAND2_X1 U9178 ( .A1(n9091), .A2(n9099), .ZN(n9098) );
  NAND2_X1 U9179 ( .A1(n9029), .A2(n9068), .ZN(n9097) );
  NOR2_X1 U9180 ( .A1(n9082), .A2(n9092), .ZN(n9095) );
  INV_X1 U9181 ( .A(n9086), .ZN(n9093) );
  NAND2_X1 U9182 ( .A1(n9100), .A2(n9078), .ZN(n9086) );
  NAND2_X1 U9183 ( .A1(n9101), .A2(n9102), .ZN(Result_61_) );
  NAND2_X1 U9184 ( .A1(n9103), .A2(n9027), .ZN(n9102) );
  XNOR2_X1 U9185 ( .A(n9104), .B(n9105), .ZN(n9103) );
  XOR2_X1 U9186 ( .A(n9106), .B(n9107), .Z(n9105) );
  NOR2_X1 U9187 ( .A1(n9108), .A2(n9109), .ZN(n9101) );
  NOR2_X1 U9188 ( .A1(n9110), .A2(n9111), .ZN(n9109) );
  NOR2_X1 U9189 ( .A1(n9112), .A2(n9113), .ZN(n9110) );
  NAND2_X1 U9190 ( .A1(n9114), .A2(n9115), .ZN(n9113) );
  NAND2_X1 U9191 ( .A1(n9091), .A2(n9116), .ZN(n9115) );
  NAND2_X1 U9192 ( .A1(n9029), .A2(n9117), .ZN(n9114) );
  NOR2_X1 U9193 ( .A1(n9118), .A2(n9092), .ZN(n9112) );
  NOR2_X1 U9194 ( .A1(n9119), .A2(n9120), .ZN(n9108) );
  INV_X1 U9195 ( .A(n9111), .ZN(n9120) );
  XNOR2_X1 U9196 ( .A(b_29_), .B(n9121), .ZN(n9111) );
  NOR2_X1 U9197 ( .A1(n9122), .A2(n9123), .ZN(n9119) );
  NAND2_X1 U9198 ( .A1(n9124), .A2(n9125), .ZN(n9123) );
  INV_X1 U9199 ( .A(n9126), .ZN(n9125) );
  NOR2_X1 U9200 ( .A1(n9116), .A2(n9064), .ZN(n9126) );
  NAND2_X1 U9201 ( .A1(n9029), .A2(n9127), .ZN(n9124) );
  NOR2_X1 U9202 ( .A1(n9128), .A2(n9092), .ZN(n9122) );
  NAND2_X1 U9203 ( .A1(n9129), .A2(n9130), .ZN(Result_60_) );
  NAND2_X1 U9204 ( .A1(n9131), .A2(n9027), .ZN(n9130) );
  XNOR2_X1 U9205 ( .A(n9132), .B(n9133), .ZN(n9131) );
  XNOR2_X1 U9206 ( .A(n9134), .B(n9135), .ZN(n9132) );
  NOR2_X1 U9207 ( .A1(n9136), .A2(n9077), .ZN(n9135) );
  NOR2_X1 U9208 ( .A1(n9137), .A2(n9138), .ZN(n9129) );
  NOR2_X1 U9209 ( .A1(n9139), .A2(n9140), .ZN(n9138) );
  NOR2_X1 U9210 ( .A1(n9141), .A2(n9142), .ZN(n9139) );
  NAND2_X1 U9211 ( .A1(n9143), .A2(n9144), .ZN(n9142) );
  NAND2_X1 U9212 ( .A1(n9091), .A2(n9145), .ZN(n9144) );
  NAND2_X1 U9213 ( .A1(n9029), .A2(n9146), .ZN(n9143) );
  NOR2_X1 U9214 ( .A1(n9092), .A2(n9147), .ZN(n9141) );
  NOR2_X1 U9215 ( .A1(n9148), .A2(n9149), .ZN(n9137) );
  NOR2_X1 U9216 ( .A1(n9150), .A2(n9151), .ZN(n9149) );
  NAND2_X1 U9217 ( .A1(n9152), .A2(n9153), .ZN(n9151) );
  NAND2_X1 U9218 ( .A1(n9154), .A2(n9091), .ZN(n9153) );
  NAND2_X1 U9219 ( .A1(n9029), .A2(n9155), .ZN(n9152) );
  INV_X1 U9220 ( .A(n9156), .ZN(n9150) );
  NAND2_X1 U9221 ( .A1(n9147), .A2(n9065), .ZN(n9156) );
  INV_X1 U9222 ( .A(n9140), .ZN(n9148) );
  NAND2_X1 U9223 ( .A1(n9157), .A2(n9158), .ZN(n9140) );
  NAND2_X1 U9224 ( .A1(n9030), .A2(n9159), .ZN(Result_5_) );
  NAND2_X1 U9225 ( .A1(n9027), .A2(n9160), .ZN(n9159) );
  XOR2_X1 U9226 ( .A(n9161), .B(n9162), .Z(n9160) );
  NOR2_X1 U9227 ( .A1(n9163), .A2(n9164), .ZN(n9162) );
  INV_X1 U9228 ( .A(n9165), .ZN(n9164) );
  NOR2_X1 U9229 ( .A1(n9166), .A2(n9167), .ZN(n9163) );
  NAND2_X1 U9230 ( .A1(n9168), .A2(n9169), .ZN(Result_59_) );
  NAND2_X1 U9231 ( .A1(n9170), .A2(n9027), .ZN(n9169) );
  XNOR2_X1 U9232 ( .A(n9171), .B(n9172), .ZN(n9170) );
  XOR2_X1 U9233 ( .A(n9173), .B(n9174), .Z(n9172) );
  NOR2_X1 U9234 ( .A1(n9175), .A2(n9176), .ZN(n9168) );
  NOR2_X1 U9235 ( .A1(n9177), .A2(n9178), .ZN(n9176) );
  NOR2_X1 U9236 ( .A1(n9179), .A2(n9180), .ZN(n9177) );
  NAND2_X1 U9237 ( .A1(n9181), .A2(n9182), .ZN(n9180) );
  INV_X1 U9238 ( .A(n9183), .ZN(n9182) );
  NOR2_X1 U9239 ( .A1(n9064), .A2(n9184), .ZN(n9183) );
  NAND2_X1 U9240 ( .A1(n9029), .A2(n9185), .ZN(n9181) );
  NOR2_X1 U9241 ( .A1(n9092), .A2(n9186), .ZN(n9179) );
  NOR2_X1 U9242 ( .A1(n9187), .A2(n9188), .ZN(n9175) );
  NOR2_X1 U9243 ( .A1(n9189), .A2(n9190), .ZN(n9188) );
  NAND2_X1 U9244 ( .A1(n9191), .A2(n9192), .ZN(n9190) );
  NAND2_X1 U9245 ( .A1(n9184), .A2(n9091), .ZN(n9192) );
  NAND2_X1 U9246 ( .A1(n9193), .A2(n9029), .ZN(n9191) );
  INV_X1 U9247 ( .A(n9185), .ZN(n9193) );
  INV_X1 U9248 ( .A(n9194), .ZN(n9189) );
  NAND2_X1 U9249 ( .A1(n9186), .A2(n9065), .ZN(n9194) );
  INV_X1 U9250 ( .A(n9178), .ZN(n9187) );
  NAND2_X1 U9251 ( .A1(n9195), .A2(n9196), .ZN(n9178) );
  NAND2_X1 U9252 ( .A1(n9197), .A2(n9198), .ZN(Result_58_) );
  NAND2_X1 U9253 ( .A1(n9199), .A2(n9027), .ZN(n9198) );
  XNOR2_X1 U9254 ( .A(n9200), .B(n9201), .ZN(n9199) );
  XNOR2_X1 U9255 ( .A(n9202), .B(n9203), .ZN(n9200) );
  NOR2_X1 U9256 ( .A1(n9204), .A2(n9205), .ZN(n9197) );
  NOR2_X1 U9257 ( .A1(n9206), .A2(n9207), .ZN(n9205) );
  NOR2_X1 U9258 ( .A1(n9208), .A2(n9209), .ZN(n9206) );
  NAND2_X1 U9259 ( .A1(n9210), .A2(n9211), .ZN(n9209) );
  NAND2_X1 U9260 ( .A1(n9091), .A2(n9212), .ZN(n9211) );
  NAND2_X1 U9261 ( .A1(n9029), .A2(n9213), .ZN(n9210) );
  NOR2_X1 U9262 ( .A1(n9214), .A2(n9092), .ZN(n9208) );
  NOR2_X1 U9263 ( .A1(n9215), .A2(n9216), .ZN(n9204) );
  INV_X1 U9264 ( .A(n9207), .ZN(n9216) );
  XNOR2_X1 U9265 ( .A(a_26_), .B(n9217), .ZN(n9207) );
  NOR2_X1 U9266 ( .A1(n9218), .A2(n9219), .ZN(n9215) );
  NAND2_X1 U9267 ( .A1(n9220), .A2(n9221), .ZN(n9219) );
  NAND2_X1 U9268 ( .A1(n9222), .A2(n9091), .ZN(n9221) );
  NAND2_X1 U9269 ( .A1(n9029), .A2(n9223), .ZN(n9220) );
  NOR2_X1 U9270 ( .A1(n9224), .A2(n9092), .ZN(n9218) );
  NAND2_X1 U9271 ( .A1(n9225), .A2(n9226), .ZN(Result_57_) );
  NAND2_X1 U9272 ( .A1(n9227), .A2(n9027), .ZN(n9226) );
  XNOR2_X1 U9273 ( .A(n9228), .B(n9229), .ZN(n9227) );
  NAND2_X1 U9274 ( .A1(n9230), .A2(n9231), .ZN(n9228) );
  NOR2_X1 U9275 ( .A1(n9232), .A2(n9233), .ZN(n9225) );
  NOR2_X1 U9276 ( .A1(n9234), .A2(n9235), .ZN(n9233) );
  NOR2_X1 U9277 ( .A1(n9236), .A2(n9237), .ZN(n9234) );
  NAND2_X1 U9278 ( .A1(n9238), .A2(n9239), .ZN(n9237) );
  NAND2_X1 U9279 ( .A1(n9091), .A2(n9240), .ZN(n9239) );
  NAND2_X1 U9280 ( .A1(n9029), .A2(n9241), .ZN(n9238) );
  NOR2_X1 U9281 ( .A1(n9242), .A2(n9092), .ZN(n9236) );
  NOR2_X1 U9282 ( .A1(n9243), .A2(n9244), .ZN(n9232) );
  INV_X1 U9283 ( .A(n9235), .ZN(n9244) );
  XNOR2_X1 U9284 ( .A(a_25_), .B(n9245), .ZN(n9235) );
  NOR2_X1 U9285 ( .A1(n9246), .A2(n9247), .ZN(n9243) );
  NAND2_X1 U9286 ( .A1(n9248), .A2(n9249), .ZN(n9247) );
  INV_X1 U9287 ( .A(n9250), .ZN(n9249) );
  NOR2_X1 U9288 ( .A1(n9240), .A2(n9064), .ZN(n9250) );
  NAND2_X1 U9289 ( .A1(n9029), .A2(n9251), .ZN(n9248) );
  NOR2_X1 U9290 ( .A1(n9252), .A2(n9092), .ZN(n9246) );
  NAND2_X1 U9291 ( .A1(n9253), .A2(n9254), .ZN(Result_56_) );
  NAND2_X1 U9292 ( .A1(n9027), .A2(n9255), .ZN(n9254) );
  XOR2_X1 U9293 ( .A(n9256), .B(n9257), .Z(n9255) );
  XOR2_X1 U9294 ( .A(n9258), .B(n9259), .Z(n9257) );
  NOR2_X1 U9295 ( .A1(n9260), .A2(n9261), .ZN(n9253) );
  NOR2_X1 U9296 ( .A1(n9262), .A2(n9263), .ZN(n9261) );
  NOR2_X1 U9297 ( .A1(n9264), .A2(n9265), .ZN(n9262) );
  NAND2_X1 U9298 ( .A1(n9266), .A2(n9267), .ZN(n9265) );
  NAND2_X1 U9299 ( .A1(n9091), .A2(n9268), .ZN(n9267) );
  NAND2_X1 U9300 ( .A1(n9029), .A2(n9269), .ZN(n9266) );
  INV_X1 U9301 ( .A(n9270), .ZN(n9264) );
  NAND2_X1 U9302 ( .A1(n9271), .A2(n9065), .ZN(n9270) );
  NOR2_X1 U9303 ( .A1(n9272), .A2(n9273), .ZN(n9260) );
  NOR2_X1 U9304 ( .A1(n9274), .A2(n9275), .ZN(n9273) );
  NAND2_X1 U9305 ( .A1(n9276), .A2(n9277), .ZN(n9275) );
  INV_X1 U9306 ( .A(n9278), .ZN(n9277) );
  NOR2_X1 U9307 ( .A1(n9268), .A2(n9064), .ZN(n9278) );
  NAND2_X1 U9308 ( .A1(n9029), .A2(n9279), .ZN(n9276) );
  NOR2_X1 U9309 ( .A1(n9092), .A2(n9271), .ZN(n9274) );
  INV_X1 U9310 ( .A(n9263), .ZN(n9272) );
  NAND2_X1 U9311 ( .A1(n9280), .A2(n9281), .ZN(n9263) );
  NAND2_X1 U9312 ( .A1(n9282), .A2(n9283), .ZN(Result_55_) );
  NAND2_X1 U9313 ( .A1(n9027), .A2(n9284), .ZN(n9283) );
  XOR2_X1 U9314 ( .A(n9285), .B(n9286), .Z(n9284) );
  XOR2_X1 U9315 ( .A(n9287), .B(n9288), .Z(n9286) );
  NOR2_X1 U9316 ( .A1(n9289), .A2(n9290), .ZN(n9282) );
  NOR2_X1 U9317 ( .A1(n9291), .A2(n9292), .ZN(n9290) );
  NOR2_X1 U9318 ( .A1(n9293), .A2(n9294), .ZN(n9291) );
  NAND2_X1 U9319 ( .A1(n9295), .A2(n9296), .ZN(n9294) );
  NAND2_X1 U9320 ( .A1(n9091), .A2(n9297), .ZN(n9296) );
  NAND2_X1 U9321 ( .A1(n9029), .A2(n9298), .ZN(n9295) );
  NOR2_X1 U9322 ( .A1(n9299), .A2(n9092), .ZN(n9293) );
  NOR2_X1 U9323 ( .A1(n9300), .A2(n9301), .ZN(n9289) );
  INV_X1 U9324 ( .A(n9292), .ZN(n9301) );
  XNOR2_X1 U9325 ( .A(a_23_), .B(n9302), .ZN(n9292) );
  NOR2_X1 U9326 ( .A1(n9303), .A2(n9304), .ZN(n9300) );
  NAND2_X1 U9327 ( .A1(n9305), .A2(n9306), .ZN(n9304) );
  INV_X1 U9328 ( .A(n9307), .ZN(n9306) );
  NOR2_X1 U9329 ( .A1(n9297), .A2(n9064), .ZN(n9307) );
  NAND2_X1 U9330 ( .A1(n9029), .A2(n9308), .ZN(n9305) );
  NOR2_X1 U9331 ( .A1(n9309), .A2(n9092), .ZN(n9303) );
  NAND2_X1 U9332 ( .A1(n9310), .A2(n9311), .ZN(Result_54_) );
  NAND2_X1 U9333 ( .A1(n9027), .A2(n9312), .ZN(n9311) );
  XNOR2_X1 U9334 ( .A(n9313), .B(n9314), .ZN(n9312) );
  XOR2_X1 U9335 ( .A(n9315), .B(n9316), .Z(n9314) );
  NOR2_X1 U9336 ( .A1(n9317), .A2(n9318), .ZN(n9310) );
  NOR2_X1 U9337 ( .A1(n9319), .A2(n9320), .ZN(n9318) );
  NOR2_X1 U9338 ( .A1(n9321), .A2(n9322), .ZN(n9319) );
  NAND2_X1 U9339 ( .A1(n9323), .A2(n9324), .ZN(n9322) );
  NAND2_X1 U9340 ( .A1(n9091), .A2(n9325), .ZN(n9324) );
  NAND2_X1 U9341 ( .A1(n9029), .A2(n9326), .ZN(n9323) );
  NOR2_X1 U9342 ( .A1(n9327), .A2(n9092), .ZN(n9321) );
  NOR2_X1 U9343 ( .A1(n9328), .A2(n9329), .ZN(n9317) );
  INV_X1 U9344 ( .A(n9320), .ZN(n9329) );
  XNOR2_X1 U9345 ( .A(b_22_), .B(n9330), .ZN(n9320) );
  NOR2_X1 U9346 ( .A1(n9331), .A2(n9332), .ZN(n9328) );
  NAND2_X1 U9347 ( .A1(n9333), .A2(n9334), .ZN(n9332) );
  NAND2_X1 U9348 ( .A1(n9335), .A2(n9091), .ZN(n9334) );
  NAND2_X1 U9349 ( .A1(n9029), .A2(n9336), .ZN(n9333) );
  NOR2_X1 U9350 ( .A1(n9337), .A2(n9092), .ZN(n9331) );
  NAND2_X1 U9351 ( .A1(n9338), .A2(n9339), .ZN(Result_53_) );
  NAND2_X1 U9352 ( .A1(n9027), .A2(n9340), .ZN(n9339) );
  XNOR2_X1 U9353 ( .A(n9341), .B(n9342), .ZN(n9340) );
  NAND2_X1 U9354 ( .A1(n9343), .A2(n9344), .ZN(n9341) );
  NOR2_X1 U9355 ( .A1(n9345), .A2(n9346), .ZN(n9338) );
  NOR2_X1 U9356 ( .A1(n9347), .A2(n9348), .ZN(n9346) );
  NOR2_X1 U9357 ( .A1(n9349), .A2(n9350), .ZN(n9347) );
  NAND2_X1 U9358 ( .A1(n9351), .A2(n9352), .ZN(n9350) );
  NAND2_X1 U9359 ( .A1(n9091), .A2(n9353), .ZN(n9352) );
  NAND2_X1 U9360 ( .A1(n9029), .A2(n9354), .ZN(n9351) );
  NOR2_X1 U9361 ( .A1(n9355), .A2(n9092), .ZN(n9349) );
  NOR2_X1 U9362 ( .A1(n9356), .A2(n9357), .ZN(n9345) );
  INV_X1 U9363 ( .A(n9348), .ZN(n9357) );
  XNOR2_X1 U9364 ( .A(b_21_), .B(n9358), .ZN(n9348) );
  NOR2_X1 U9365 ( .A1(n9359), .A2(n9360), .ZN(n9356) );
  NAND2_X1 U9366 ( .A1(n9361), .A2(n9362), .ZN(n9360) );
  NAND2_X1 U9367 ( .A1(n9363), .A2(n9091), .ZN(n9362) );
  NAND2_X1 U9368 ( .A1(n9029), .A2(n9364), .ZN(n9361) );
  NOR2_X1 U9369 ( .A1(n9365), .A2(n9092), .ZN(n9359) );
  NAND2_X1 U9370 ( .A1(n9366), .A2(n9367), .ZN(Result_52_) );
  NAND2_X1 U9371 ( .A1(n9027), .A2(n9368), .ZN(n9367) );
  XOR2_X1 U9372 ( .A(n9369), .B(n9370), .Z(n9368) );
  XOR2_X1 U9373 ( .A(n9371), .B(n9372), .Z(n9370) );
  NOR2_X1 U9374 ( .A1(n9373), .A2(n9374), .ZN(n9366) );
  NOR2_X1 U9375 ( .A1(n9375), .A2(n9376), .ZN(n9374) );
  NOR2_X1 U9376 ( .A1(n9377), .A2(n9378), .ZN(n9375) );
  NAND2_X1 U9377 ( .A1(n9379), .A2(n9380), .ZN(n9378) );
  INV_X1 U9378 ( .A(n9381), .ZN(n9380) );
  NOR2_X1 U9379 ( .A1(n9382), .A2(n9064), .ZN(n9381) );
  NAND2_X1 U9380 ( .A1(n9029), .A2(n9383), .ZN(n9379) );
  NOR2_X1 U9381 ( .A1(n9384), .A2(n9092), .ZN(n9377) );
  NOR2_X1 U9382 ( .A1(n9385), .A2(n9386), .ZN(n9373) );
  NOR2_X1 U9383 ( .A1(n9387), .A2(n9388), .ZN(n9386) );
  NAND2_X1 U9384 ( .A1(n9389), .A2(n9390), .ZN(n9388) );
  NAND2_X1 U9385 ( .A1(n9091), .A2(n9382), .ZN(n9390) );
  NAND2_X1 U9386 ( .A1(n9029), .A2(n9391), .ZN(n9389) );
  NOR2_X1 U9387 ( .A1(n9392), .A2(n9092), .ZN(n9387) );
  INV_X1 U9388 ( .A(n9376), .ZN(n9385) );
  NAND2_X1 U9389 ( .A1(n9393), .A2(n9394), .ZN(n9376) );
  NAND2_X1 U9390 ( .A1(n9395), .A2(n9396), .ZN(Result_51_) );
  NAND2_X1 U9391 ( .A1(n9397), .A2(n9027), .ZN(n9396) );
  XNOR2_X1 U9392 ( .A(n9398), .B(n9399), .ZN(n9397) );
  XNOR2_X1 U9393 ( .A(n9400), .B(n9401), .ZN(n9398) );
  NOR2_X1 U9394 ( .A1(n9402), .A2(n9403), .ZN(n9395) );
  NOR2_X1 U9395 ( .A1(n9404), .A2(n9405), .ZN(n9403) );
  NOR2_X1 U9396 ( .A1(n9406), .A2(n9407), .ZN(n9404) );
  NAND2_X1 U9397 ( .A1(n9408), .A2(n9409), .ZN(n9407) );
  NAND2_X1 U9398 ( .A1(n9091), .A2(n9410), .ZN(n9409) );
  NAND2_X1 U9399 ( .A1(n9029), .A2(n9411), .ZN(n9408) );
  NOR2_X1 U9400 ( .A1(n9412), .A2(n9092), .ZN(n9406) );
  NOR2_X1 U9401 ( .A1(n9413), .A2(n9414), .ZN(n9402) );
  INV_X1 U9402 ( .A(n9405), .ZN(n9414) );
  XNOR2_X1 U9403 ( .A(b_19_), .B(n9415), .ZN(n9405) );
  NOR2_X1 U9404 ( .A1(n9416), .A2(n9417), .ZN(n9413) );
  NAND2_X1 U9405 ( .A1(n9418), .A2(n9419), .ZN(n9417) );
  INV_X1 U9406 ( .A(n9420), .ZN(n9419) );
  NOR2_X1 U9407 ( .A1(n9410), .A2(n9064), .ZN(n9420) );
  NAND2_X1 U9408 ( .A1(n9029), .A2(n9421), .ZN(n9418) );
  NOR2_X1 U9409 ( .A1(n9422), .A2(n9092), .ZN(n9416) );
  NAND2_X1 U9410 ( .A1(n9423), .A2(n9424), .ZN(Result_50_) );
  NAND2_X1 U9411 ( .A1(n9425), .A2(n9027), .ZN(n9424) );
  XOR2_X1 U9412 ( .A(n9426), .B(n9427), .Z(n9425) );
  XOR2_X1 U9413 ( .A(n9428), .B(n9429), .Z(n9426) );
  NOR2_X1 U9414 ( .A1(n9430), .A2(n9431), .ZN(n9423) );
  NOR2_X1 U9415 ( .A1(n9432), .A2(n9433), .ZN(n9431) );
  NOR2_X1 U9416 ( .A1(n9434), .A2(n9435), .ZN(n9432) );
  NAND2_X1 U9417 ( .A1(n9436), .A2(n9437), .ZN(n9435) );
  INV_X1 U9418 ( .A(n9438), .ZN(n9437) );
  NOR2_X1 U9419 ( .A1(n9439), .A2(n9064), .ZN(n9438) );
  NAND2_X1 U9420 ( .A1(n9029), .A2(n9440), .ZN(n9436) );
  NOR2_X1 U9421 ( .A1(n9441), .A2(n9092), .ZN(n9434) );
  NOR2_X1 U9422 ( .A1(n9442), .A2(n9443), .ZN(n9430) );
  NOR2_X1 U9423 ( .A1(n9444), .A2(n9445), .ZN(n9443) );
  NAND2_X1 U9424 ( .A1(n9446), .A2(n9447), .ZN(n9445) );
  NAND2_X1 U9425 ( .A1(n9091), .A2(n9439), .ZN(n9447) );
  NAND2_X1 U9426 ( .A1(n9029), .A2(n9448), .ZN(n9446) );
  NOR2_X1 U9427 ( .A1(n9449), .A2(n9092), .ZN(n9444) );
  INV_X1 U9428 ( .A(n9433), .ZN(n9442) );
  NAND2_X1 U9429 ( .A1(n9450), .A2(n9451), .ZN(n9433) );
  NAND2_X1 U9430 ( .A1(n9030), .A2(n9452), .ZN(Result_4_) );
  NAND2_X1 U9431 ( .A1(n9453), .A2(n9027), .ZN(n9452) );
  XOR2_X1 U9432 ( .A(n9454), .B(n9455), .Z(n9453) );
  NAND2_X1 U9433 ( .A1(n9456), .A2(n9457), .ZN(Result_49_) );
  NAND2_X1 U9434 ( .A1(n9027), .A2(n9458), .ZN(n9457) );
  XOR2_X1 U9435 ( .A(n9459), .B(n9460), .Z(n9458) );
  XNOR2_X1 U9436 ( .A(n9461), .B(n9462), .ZN(n9460) );
  NAND2_X1 U9437 ( .A1(a_17_), .A2(b_31_), .ZN(n9462) );
  NOR2_X1 U9438 ( .A1(n9463), .A2(n9464), .ZN(n9456) );
  NOR2_X1 U9439 ( .A1(n9465), .A2(n9466), .ZN(n9464) );
  NOR2_X1 U9440 ( .A1(n9467), .A2(n9468), .ZN(n9465) );
  NAND2_X1 U9441 ( .A1(n9469), .A2(n9470), .ZN(n9468) );
  INV_X1 U9442 ( .A(n9471), .ZN(n9470) );
  NOR2_X1 U9443 ( .A1(n9472), .A2(n9064), .ZN(n9471) );
  NAND2_X1 U9444 ( .A1(n9029), .A2(n9473), .ZN(n9469) );
  NOR2_X1 U9445 ( .A1(n9474), .A2(n9092), .ZN(n9467) );
  NOR2_X1 U9446 ( .A1(n9475), .A2(n9476), .ZN(n9463) );
  NOR2_X1 U9447 ( .A1(n9477), .A2(n9478), .ZN(n9476) );
  NAND2_X1 U9448 ( .A1(n9479), .A2(n9480), .ZN(n9478) );
  NAND2_X1 U9449 ( .A1(n9091), .A2(n9472), .ZN(n9480) );
  NAND2_X1 U9450 ( .A1(n9029), .A2(n9481), .ZN(n9479) );
  NOR2_X1 U9451 ( .A1(n9482), .A2(n9092), .ZN(n9477) );
  INV_X1 U9452 ( .A(n9466), .ZN(n9475) );
  NAND2_X1 U9453 ( .A1(n9483), .A2(n9484), .ZN(n9466) );
  NAND2_X1 U9454 ( .A1(n9485), .A2(n9486), .ZN(Result_48_) );
  NAND2_X1 U9455 ( .A1(n9487), .A2(n9027), .ZN(n9486) );
  XNOR2_X1 U9456 ( .A(n9488), .B(n9489), .ZN(n9487) );
  XOR2_X1 U9457 ( .A(n9490), .B(n9491), .Z(n9489) );
  NAND2_X1 U9458 ( .A1(a_16_), .A2(b_31_), .ZN(n9491) );
  NOR2_X1 U9459 ( .A1(n9492), .A2(n9493), .ZN(n9485) );
  NOR2_X1 U9460 ( .A1(n9494), .A2(n9495), .ZN(n9493) );
  NOR2_X1 U9461 ( .A1(n9496), .A2(n9497), .ZN(n9494) );
  NAND2_X1 U9462 ( .A1(n9498), .A2(n9499), .ZN(n9497) );
  INV_X1 U9463 ( .A(n9500), .ZN(n9499) );
  NOR2_X1 U9464 ( .A1(n9501), .A2(n9064), .ZN(n9500) );
  NAND2_X1 U9465 ( .A1(n9029), .A2(n9502), .ZN(n9498) );
  NOR2_X1 U9466 ( .A1(n9503), .A2(n9092), .ZN(n9496) );
  NOR2_X1 U9467 ( .A1(n9504), .A2(n9505), .ZN(n9492) );
  NOR2_X1 U9468 ( .A1(n9506), .A2(n9507), .ZN(n9505) );
  NAND2_X1 U9469 ( .A1(n9508), .A2(n9509), .ZN(n9507) );
  NAND2_X1 U9470 ( .A1(n9091), .A2(n9501), .ZN(n9509) );
  NAND2_X1 U9471 ( .A1(n9029), .A2(n9510), .ZN(n9508) );
  NOR2_X1 U9472 ( .A1(n9511), .A2(n9092), .ZN(n9506) );
  INV_X1 U9473 ( .A(n9495), .ZN(n9504) );
  NAND2_X1 U9474 ( .A1(n9512), .A2(n9513), .ZN(n9495) );
  NAND2_X1 U9475 ( .A1(n9514), .A2(n9515), .ZN(Result_47_) );
  NAND2_X1 U9476 ( .A1(n9516), .A2(n9027), .ZN(n9515) );
  XNOR2_X1 U9477 ( .A(n9517), .B(n9518), .ZN(n9516) );
  XOR2_X1 U9478 ( .A(n9519), .B(n9520), .Z(n9518) );
  NAND2_X1 U9479 ( .A1(a_15_), .A2(b_31_), .ZN(n9520) );
  NOR2_X1 U9480 ( .A1(n9521), .A2(n9522), .ZN(n9514) );
  NOR2_X1 U9481 ( .A1(n9523), .A2(n9524), .ZN(n9522) );
  NOR2_X1 U9482 ( .A1(n9525), .A2(n9526), .ZN(n9523) );
  NAND2_X1 U9483 ( .A1(n9527), .A2(n9528), .ZN(n9526) );
  NAND2_X1 U9484 ( .A1(n9091), .A2(n9529), .ZN(n9528) );
  NAND2_X1 U9485 ( .A1(n9029), .A2(n9530), .ZN(n9527) );
  NOR2_X1 U9486 ( .A1(n9531), .A2(n9092), .ZN(n9525) );
  NOR2_X1 U9487 ( .A1(n9532), .A2(n9533), .ZN(n9521) );
  INV_X1 U9488 ( .A(n9524), .ZN(n9533) );
  XNOR2_X1 U9489 ( .A(b_15_), .B(n9534), .ZN(n9524) );
  NOR2_X1 U9490 ( .A1(n9535), .A2(n9536), .ZN(n9532) );
  NAND2_X1 U9491 ( .A1(n9537), .A2(n9538), .ZN(n9536) );
  INV_X1 U9492 ( .A(n9539), .ZN(n9538) );
  NOR2_X1 U9493 ( .A1(n9529), .A2(n9064), .ZN(n9539) );
  NAND2_X1 U9494 ( .A1(n9029), .A2(n9540), .ZN(n9537) );
  NOR2_X1 U9495 ( .A1(n9541), .A2(n9092), .ZN(n9535) );
  NAND2_X1 U9496 ( .A1(n9542), .A2(n9543), .ZN(Result_46_) );
  NAND2_X1 U9497 ( .A1(n9027), .A2(n9544), .ZN(n9543) );
  XNOR2_X1 U9498 ( .A(n9545), .B(n9546), .ZN(n9544) );
  XOR2_X1 U9499 ( .A(n9547), .B(n9548), .Z(n9546) );
  NAND2_X1 U9500 ( .A1(a_14_), .A2(b_31_), .ZN(n9548) );
  NOR2_X1 U9501 ( .A1(n9549), .A2(n9550), .ZN(n9542) );
  NOR2_X1 U9502 ( .A1(n9551), .A2(n9552), .ZN(n9550) );
  NOR2_X1 U9503 ( .A1(n9553), .A2(n9554), .ZN(n9551) );
  NAND2_X1 U9504 ( .A1(n9555), .A2(n9556), .ZN(n9554) );
  INV_X1 U9505 ( .A(n9557), .ZN(n9556) );
  NOR2_X1 U9506 ( .A1(n9558), .A2(n9064), .ZN(n9557) );
  NAND2_X1 U9507 ( .A1(n9029), .A2(n9559), .ZN(n9555) );
  NOR2_X1 U9508 ( .A1(n9560), .A2(n9092), .ZN(n9553) );
  NOR2_X1 U9509 ( .A1(n9561), .A2(n9562), .ZN(n9549) );
  NOR2_X1 U9510 ( .A1(n9563), .A2(n9564), .ZN(n9562) );
  NAND2_X1 U9511 ( .A1(n9565), .A2(n9566), .ZN(n9564) );
  NAND2_X1 U9512 ( .A1(n9091), .A2(n9558), .ZN(n9566) );
  NAND2_X1 U9513 ( .A1(n9029), .A2(n9567), .ZN(n9565) );
  NOR2_X1 U9514 ( .A1(n9568), .A2(n9092), .ZN(n9563) );
  INV_X1 U9515 ( .A(n9552), .ZN(n9561) );
  NAND2_X1 U9516 ( .A1(n9569), .A2(n9570), .ZN(n9552) );
  NAND2_X1 U9517 ( .A1(n9571), .A2(n9572), .ZN(Result_45_) );
  NAND2_X1 U9518 ( .A1(n9027), .A2(n9573), .ZN(n9572) );
  XNOR2_X1 U9519 ( .A(n9574), .B(n9575), .ZN(n9573) );
  XOR2_X1 U9520 ( .A(n9576), .B(n9577), .Z(n9575) );
  NAND2_X1 U9521 ( .A1(a_13_), .A2(b_31_), .ZN(n9577) );
  NOR2_X1 U9522 ( .A1(n9578), .A2(n9579), .ZN(n9571) );
  NOR2_X1 U9523 ( .A1(n9580), .A2(n9581), .ZN(n9579) );
  NOR2_X1 U9524 ( .A1(n9582), .A2(n9583), .ZN(n9580) );
  NAND2_X1 U9525 ( .A1(n9584), .A2(n9585), .ZN(n9583) );
  INV_X1 U9526 ( .A(n9586), .ZN(n9585) );
  NOR2_X1 U9527 ( .A1(n9587), .A2(n9064), .ZN(n9586) );
  NAND2_X1 U9528 ( .A1(n9029), .A2(n9588), .ZN(n9584) );
  NOR2_X1 U9529 ( .A1(n9589), .A2(n9092), .ZN(n9582) );
  NOR2_X1 U9530 ( .A1(n9590), .A2(n9591), .ZN(n9578) );
  NOR2_X1 U9531 ( .A1(n9592), .A2(n9593), .ZN(n9591) );
  NAND2_X1 U9532 ( .A1(n9594), .A2(n9595), .ZN(n9593) );
  NAND2_X1 U9533 ( .A1(n9091), .A2(n9587), .ZN(n9595) );
  NAND2_X1 U9534 ( .A1(n9029), .A2(n9596), .ZN(n9594) );
  NOR2_X1 U9535 ( .A1(n9597), .A2(n9092), .ZN(n9592) );
  INV_X1 U9536 ( .A(n9581), .ZN(n9590) );
  NAND2_X1 U9537 ( .A1(n9598), .A2(n9599), .ZN(n9581) );
  NAND2_X1 U9538 ( .A1(n9600), .A2(n9601), .ZN(Result_44_) );
  NAND2_X1 U9539 ( .A1(n9027), .A2(n9602), .ZN(n9601) );
  XNOR2_X1 U9540 ( .A(n9603), .B(n9604), .ZN(n9602) );
  XOR2_X1 U9541 ( .A(n9605), .B(n9606), .Z(n9604) );
  NAND2_X1 U9542 ( .A1(a_12_), .A2(b_31_), .ZN(n9606) );
  NOR2_X1 U9543 ( .A1(n9607), .A2(n9608), .ZN(n9600) );
  NOR2_X1 U9544 ( .A1(n9609), .A2(n9610), .ZN(n9608) );
  NOR2_X1 U9545 ( .A1(n9611), .A2(n9612), .ZN(n9609) );
  NAND2_X1 U9546 ( .A1(n9613), .A2(n9614), .ZN(n9612) );
  INV_X1 U9547 ( .A(n9615), .ZN(n9614) );
  NOR2_X1 U9548 ( .A1(n9616), .A2(n9064), .ZN(n9615) );
  NAND2_X1 U9549 ( .A1(n9029), .A2(n9617), .ZN(n9613) );
  NOR2_X1 U9550 ( .A1(n9618), .A2(n9092), .ZN(n9611) );
  NOR2_X1 U9551 ( .A1(n9619), .A2(n9620), .ZN(n9607) );
  NOR2_X1 U9552 ( .A1(n9621), .A2(n9622), .ZN(n9620) );
  NAND2_X1 U9553 ( .A1(n9623), .A2(n9624), .ZN(n9622) );
  NAND2_X1 U9554 ( .A1(n9091), .A2(n9616), .ZN(n9624) );
  NAND2_X1 U9555 ( .A1(n9029), .A2(n9625), .ZN(n9623) );
  NOR2_X1 U9556 ( .A1(n9626), .A2(n9092), .ZN(n9621) );
  INV_X1 U9557 ( .A(n9610), .ZN(n9619) );
  NAND2_X1 U9558 ( .A1(n9627), .A2(n9628), .ZN(n9610) );
  NAND2_X1 U9559 ( .A1(n9629), .A2(n9630), .ZN(Result_43_) );
  NAND2_X1 U9560 ( .A1(n9027), .A2(n9631), .ZN(n9630) );
  XNOR2_X1 U9561 ( .A(n9632), .B(n9633), .ZN(n9631) );
  XOR2_X1 U9562 ( .A(n9634), .B(n9635), .Z(n9633) );
  NAND2_X1 U9563 ( .A1(a_11_), .A2(b_31_), .ZN(n9635) );
  NOR2_X1 U9564 ( .A1(n9636), .A2(n9637), .ZN(n9629) );
  NOR2_X1 U9565 ( .A1(n9638), .A2(n9639), .ZN(n9637) );
  NOR2_X1 U9566 ( .A1(n9640), .A2(n9641), .ZN(n9638) );
  NAND2_X1 U9567 ( .A1(n9642), .A2(n9643), .ZN(n9641) );
  NAND2_X1 U9568 ( .A1(n9091), .A2(n9644), .ZN(n9643) );
  NAND2_X1 U9569 ( .A1(n9029), .A2(n9645), .ZN(n9642) );
  NOR2_X1 U9570 ( .A1(n9646), .A2(n9092), .ZN(n9640) );
  NOR2_X1 U9571 ( .A1(n9647), .A2(n9648), .ZN(n9636) );
  INV_X1 U9572 ( .A(n9639), .ZN(n9648) );
  XNOR2_X1 U9573 ( .A(b_11_), .B(n9649), .ZN(n9639) );
  NOR2_X1 U9574 ( .A1(n9650), .A2(n9651), .ZN(n9647) );
  NAND2_X1 U9575 ( .A1(n9652), .A2(n9653), .ZN(n9651) );
  INV_X1 U9576 ( .A(n9654), .ZN(n9653) );
  NOR2_X1 U9577 ( .A1(n9644), .A2(n9064), .ZN(n9654) );
  NAND2_X1 U9578 ( .A1(n9029), .A2(n9655), .ZN(n9652) );
  NOR2_X1 U9579 ( .A1(n9656), .A2(n9092), .ZN(n9650) );
  NAND2_X1 U9580 ( .A1(n9657), .A2(n9658), .ZN(Result_42_) );
  NAND2_X1 U9581 ( .A1(n9659), .A2(n9027), .ZN(n9658) );
  XNOR2_X1 U9582 ( .A(n9660), .B(n9661), .ZN(n9659) );
  XOR2_X1 U9583 ( .A(n9662), .B(n9663), .Z(n9661) );
  NAND2_X1 U9584 ( .A1(a_10_), .A2(b_31_), .ZN(n9663) );
  NOR2_X1 U9585 ( .A1(n9664), .A2(n9665), .ZN(n9657) );
  NOR2_X1 U9586 ( .A1(n9666), .A2(n9667), .ZN(n9665) );
  NOR2_X1 U9587 ( .A1(n9668), .A2(n9669), .ZN(n9666) );
  NAND2_X1 U9588 ( .A1(n9670), .A2(n9671), .ZN(n9669) );
  INV_X1 U9589 ( .A(n9672), .ZN(n9671) );
  NOR2_X1 U9590 ( .A1(n9673), .A2(n9064), .ZN(n9672) );
  NAND2_X1 U9591 ( .A1(n9029), .A2(n9674), .ZN(n9670) );
  NOR2_X1 U9592 ( .A1(n9675), .A2(n9092), .ZN(n9668) );
  NOR2_X1 U9593 ( .A1(n9676), .A2(n9677), .ZN(n9664) );
  NOR2_X1 U9594 ( .A1(n9678), .A2(n9679), .ZN(n9677) );
  NAND2_X1 U9595 ( .A1(n9680), .A2(n9681), .ZN(n9679) );
  NAND2_X1 U9596 ( .A1(n9091), .A2(n9673), .ZN(n9681) );
  NAND2_X1 U9597 ( .A1(n9029), .A2(n9682), .ZN(n9680) );
  NOR2_X1 U9598 ( .A1(n9683), .A2(n9092), .ZN(n9678) );
  INV_X1 U9599 ( .A(n9667), .ZN(n9676) );
  NAND2_X1 U9600 ( .A1(n9684), .A2(n9685), .ZN(n9667) );
  NAND2_X1 U9601 ( .A1(n9686), .A2(n9687), .ZN(Result_41_) );
  NAND2_X1 U9602 ( .A1(n9688), .A2(n9027), .ZN(n9687) );
  XNOR2_X1 U9603 ( .A(n9689), .B(n9690), .ZN(n9688) );
  XOR2_X1 U9604 ( .A(n9691), .B(n9692), .Z(n9690) );
  NAND2_X1 U9605 ( .A1(a_9_), .A2(b_31_), .ZN(n9692) );
  NOR2_X1 U9606 ( .A1(n9693), .A2(n9694), .ZN(n9686) );
  NOR2_X1 U9607 ( .A1(n9695), .A2(n9696), .ZN(n9694) );
  NOR2_X1 U9608 ( .A1(n9697), .A2(n9698), .ZN(n9695) );
  NAND2_X1 U9609 ( .A1(n9699), .A2(n9700), .ZN(n9698) );
  INV_X1 U9610 ( .A(n9701), .ZN(n9700) );
  NOR2_X1 U9611 ( .A1(n9702), .A2(n9064), .ZN(n9701) );
  NAND2_X1 U9612 ( .A1(n9029), .A2(n9703), .ZN(n9699) );
  NOR2_X1 U9613 ( .A1(n9704), .A2(n9092), .ZN(n9697) );
  NOR2_X1 U9614 ( .A1(n9705), .A2(n9706), .ZN(n9693) );
  NOR2_X1 U9615 ( .A1(n9707), .A2(n9708), .ZN(n9706) );
  NAND2_X1 U9616 ( .A1(n9709), .A2(n9710), .ZN(n9708) );
  NAND2_X1 U9617 ( .A1(n9091), .A2(n9702), .ZN(n9710) );
  NAND2_X1 U9618 ( .A1(n9029), .A2(n9711), .ZN(n9709) );
  NOR2_X1 U9619 ( .A1(n9712), .A2(n9092), .ZN(n9707) );
  INV_X1 U9620 ( .A(n9696), .ZN(n9705) );
  NAND2_X1 U9621 ( .A1(n9713), .A2(n9714), .ZN(n9696) );
  NAND2_X1 U9622 ( .A1(n9715), .A2(n9716), .ZN(Result_40_) );
  NAND2_X1 U9623 ( .A1(n9027), .A2(n9717), .ZN(n9716) );
  XNOR2_X1 U9624 ( .A(n9718), .B(n9719), .ZN(n9717) );
  XOR2_X1 U9625 ( .A(n9720), .B(n9721), .Z(n9719) );
  NAND2_X1 U9626 ( .A1(a_8_), .A2(b_31_), .ZN(n9721) );
  NOR2_X1 U9627 ( .A1(n9722), .A2(n9723), .ZN(n9715) );
  NOR2_X1 U9628 ( .A1(n9724), .A2(n9725), .ZN(n9723) );
  NOR2_X1 U9629 ( .A1(n9726), .A2(n9727), .ZN(n9724) );
  NAND2_X1 U9630 ( .A1(n9728), .A2(n9729), .ZN(n9727) );
  INV_X1 U9631 ( .A(n9730), .ZN(n9729) );
  NOR2_X1 U9632 ( .A1(n9731), .A2(n9064), .ZN(n9730) );
  NAND2_X1 U9633 ( .A1(n9029), .A2(n9732), .ZN(n9728) );
  NOR2_X1 U9634 ( .A1(n9733), .A2(n9092), .ZN(n9726) );
  NOR2_X1 U9635 ( .A1(n9734), .A2(n9735), .ZN(n9722) );
  NOR2_X1 U9636 ( .A1(n9736), .A2(n9737), .ZN(n9735) );
  NAND2_X1 U9637 ( .A1(n9738), .A2(n9739), .ZN(n9737) );
  NAND2_X1 U9638 ( .A1(n9091), .A2(n9731), .ZN(n9739) );
  NAND2_X1 U9639 ( .A1(n9029), .A2(n9740), .ZN(n9738) );
  NOR2_X1 U9640 ( .A1(n9741), .A2(n9092), .ZN(n9736) );
  INV_X1 U9641 ( .A(n9725), .ZN(n9734) );
  NAND2_X1 U9642 ( .A1(n9742), .A2(n9743), .ZN(n9725) );
  NAND2_X1 U9643 ( .A1(n9030), .A2(n9744), .ZN(Result_3_) );
  NAND2_X1 U9644 ( .A1(n9027), .A2(n9745), .ZN(n9744) );
  XOR2_X1 U9645 ( .A(n9746), .B(n9747), .Z(n9745) );
  NOR2_X1 U9646 ( .A1(n9748), .A2(n9749), .ZN(n9747) );
  INV_X1 U9647 ( .A(n9750), .ZN(n9749) );
  NOR2_X1 U9648 ( .A1(n9751), .A2(n9752), .ZN(n9748) );
  NAND2_X1 U9649 ( .A1(n9753), .A2(n9754), .ZN(Result_39_) );
  NAND2_X1 U9650 ( .A1(n9027), .A2(n9755), .ZN(n9754) );
  XNOR2_X1 U9651 ( .A(n9756), .B(n9757), .ZN(n9755) );
  XOR2_X1 U9652 ( .A(n9758), .B(n9759), .Z(n9757) );
  NAND2_X1 U9653 ( .A1(a_7_), .A2(b_31_), .ZN(n9759) );
  NOR2_X1 U9654 ( .A1(n9760), .A2(n9761), .ZN(n9753) );
  NOR2_X1 U9655 ( .A1(n9762), .A2(n9763), .ZN(n9761) );
  NOR2_X1 U9656 ( .A1(n9764), .A2(n9765), .ZN(n9762) );
  NAND2_X1 U9657 ( .A1(n9766), .A2(n9767), .ZN(n9765) );
  NAND2_X1 U9658 ( .A1(n9091), .A2(n9768), .ZN(n9767) );
  NAND2_X1 U9659 ( .A1(n9029), .A2(n9769), .ZN(n9766) );
  NOR2_X1 U9660 ( .A1(n9770), .A2(n9092), .ZN(n9764) );
  NOR2_X1 U9661 ( .A1(n9771), .A2(n9772), .ZN(n9760) );
  INV_X1 U9662 ( .A(n9763), .ZN(n9772) );
  XNOR2_X1 U9663 ( .A(b_7_), .B(n9773), .ZN(n9763) );
  NOR2_X1 U9664 ( .A1(n9774), .A2(n9775), .ZN(n9771) );
  NAND2_X1 U9665 ( .A1(n9776), .A2(n9777), .ZN(n9775) );
  NAND2_X1 U9666 ( .A1(n9778), .A2(n9091), .ZN(n9777) );
  NAND2_X1 U9667 ( .A1(n9029), .A2(n9779), .ZN(n9776) );
  NOR2_X1 U9668 ( .A1(n9780), .A2(n9092), .ZN(n9774) );
  NAND2_X1 U9669 ( .A1(n9781), .A2(n9782), .ZN(Result_38_) );
  NAND2_X1 U9670 ( .A1(n9027), .A2(n9783), .ZN(n9782) );
  XNOR2_X1 U9671 ( .A(n9784), .B(n9785), .ZN(n9783) );
  XOR2_X1 U9672 ( .A(n9786), .B(n9787), .Z(n9785) );
  NAND2_X1 U9673 ( .A1(a_6_), .A2(b_31_), .ZN(n9787) );
  NOR2_X1 U9674 ( .A1(n9788), .A2(n9789), .ZN(n9781) );
  NOR2_X1 U9675 ( .A1(n9790), .A2(n9791), .ZN(n9789) );
  NOR2_X1 U9676 ( .A1(n9792), .A2(n9793), .ZN(n9790) );
  NAND2_X1 U9677 ( .A1(n9794), .A2(n9795), .ZN(n9793) );
  NAND2_X1 U9678 ( .A1(n9796), .A2(n9091), .ZN(n9795) );
  NAND2_X1 U9679 ( .A1(n9029), .A2(n9797), .ZN(n9794) );
  NOR2_X1 U9680 ( .A1(n9798), .A2(n9092), .ZN(n9792) );
  NOR2_X1 U9681 ( .A1(n9799), .A2(n9800), .ZN(n9788) );
  NOR2_X1 U9682 ( .A1(n9801), .A2(n9802), .ZN(n9800) );
  NAND2_X1 U9683 ( .A1(n9803), .A2(n9804), .ZN(n9802) );
  NAND2_X1 U9684 ( .A1(n9091), .A2(n9805), .ZN(n9804) );
  NAND2_X1 U9685 ( .A1(n9029), .A2(n9806), .ZN(n9803) );
  NOR2_X1 U9686 ( .A1(n9807), .A2(n9092), .ZN(n9801) );
  INV_X1 U9687 ( .A(n9791), .ZN(n9799) );
  NAND2_X1 U9688 ( .A1(n9808), .A2(n9809), .ZN(n9791) );
  NAND2_X1 U9689 ( .A1(n9810), .A2(n9811), .ZN(Result_37_) );
  NAND2_X1 U9690 ( .A1(n9027), .A2(n9812), .ZN(n9811) );
  XNOR2_X1 U9691 ( .A(n9813), .B(n9814), .ZN(n9812) );
  XOR2_X1 U9692 ( .A(n9815), .B(n9816), .Z(n9814) );
  NAND2_X1 U9693 ( .A1(a_5_), .A2(b_31_), .ZN(n9816) );
  NOR2_X1 U9694 ( .A1(n9817), .A2(n9818), .ZN(n9810) );
  NOR2_X1 U9695 ( .A1(n9819), .A2(n9820), .ZN(n9818) );
  NOR2_X1 U9696 ( .A1(n9821), .A2(n9822), .ZN(n9819) );
  NAND2_X1 U9697 ( .A1(n9823), .A2(n9824), .ZN(n9822) );
  INV_X1 U9698 ( .A(n9825), .ZN(n9824) );
  NOR2_X1 U9699 ( .A1(n9826), .A2(n9064), .ZN(n9825) );
  NAND2_X1 U9700 ( .A1(n9029), .A2(n9827), .ZN(n9823) );
  NOR2_X1 U9701 ( .A1(n9828), .A2(n9092), .ZN(n9821) );
  NOR2_X1 U9702 ( .A1(n9829), .A2(n9830), .ZN(n9817) );
  NOR2_X1 U9703 ( .A1(n9831), .A2(n9832), .ZN(n9830) );
  NAND2_X1 U9704 ( .A1(n9833), .A2(n9834), .ZN(n9832) );
  NAND2_X1 U9705 ( .A1(n9091), .A2(n9826), .ZN(n9834) );
  NAND2_X1 U9706 ( .A1(n9029), .A2(n9835), .ZN(n9833) );
  NOR2_X1 U9707 ( .A1(n9836), .A2(n9092), .ZN(n9831) );
  INV_X1 U9708 ( .A(n9820), .ZN(n9829) );
  NAND2_X1 U9709 ( .A1(n9837), .A2(n9838), .ZN(n9820) );
  NAND2_X1 U9710 ( .A1(n9839), .A2(n9840), .ZN(Result_36_) );
  NAND2_X1 U9711 ( .A1(n9027), .A2(n9841), .ZN(n9840) );
  XNOR2_X1 U9712 ( .A(n9842), .B(n9843), .ZN(n9841) );
  XOR2_X1 U9713 ( .A(n9844), .B(n9845), .Z(n9843) );
  NAND2_X1 U9714 ( .A1(a_4_), .A2(b_31_), .ZN(n9845) );
  NOR2_X1 U9715 ( .A1(n9846), .A2(n9847), .ZN(n9839) );
  NOR2_X1 U9716 ( .A1(n9848), .A2(n9849), .ZN(n9847) );
  NOR2_X1 U9717 ( .A1(n9850), .A2(n9851), .ZN(n9848) );
  NAND2_X1 U9718 ( .A1(n9852), .A2(n9853), .ZN(n9851) );
  INV_X1 U9719 ( .A(n9854), .ZN(n9853) );
  NOR2_X1 U9720 ( .A1(n9855), .A2(n9064), .ZN(n9854) );
  NAND2_X1 U9721 ( .A1(n9029), .A2(n9856), .ZN(n9852) );
  NOR2_X1 U9722 ( .A1(n9857), .A2(n9092), .ZN(n9850) );
  NOR2_X1 U9723 ( .A1(n9858), .A2(n9859), .ZN(n9846) );
  NOR2_X1 U9724 ( .A1(n9860), .A2(n9861), .ZN(n9859) );
  NAND2_X1 U9725 ( .A1(n9862), .A2(n9863), .ZN(n9861) );
  NAND2_X1 U9726 ( .A1(n9091), .A2(n9855), .ZN(n9863) );
  NAND2_X1 U9727 ( .A1(n9029), .A2(n9864), .ZN(n9862) );
  NOR2_X1 U9728 ( .A1(n9865), .A2(n9092), .ZN(n9860) );
  INV_X1 U9729 ( .A(n9849), .ZN(n9858) );
  NAND2_X1 U9730 ( .A1(n9866), .A2(n9867), .ZN(n9849) );
  NAND2_X1 U9731 ( .A1(n9868), .A2(n9869), .ZN(Result_35_) );
  NAND2_X1 U9732 ( .A1(n9870), .A2(n9027), .ZN(n9869) );
  XNOR2_X1 U9733 ( .A(n9871), .B(n9872), .ZN(n9870) );
  XOR2_X1 U9734 ( .A(n9873), .B(n9874), .Z(n9872) );
  NAND2_X1 U9735 ( .A1(a_3_), .A2(b_31_), .ZN(n9874) );
  NOR2_X1 U9736 ( .A1(n9875), .A2(n9876), .ZN(n9868) );
  NOR2_X1 U9737 ( .A1(n9877), .A2(n9878), .ZN(n9876) );
  NOR2_X1 U9738 ( .A1(n9879), .A2(n9880), .ZN(n9877) );
  NAND2_X1 U9739 ( .A1(n9881), .A2(n9882), .ZN(n9880) );
  NAND2_X1 U9740 ( .A1(n9091), .A2(n9883), .ZN(n9882) );
  NAND2_X1 U9741 ( .A1(n9029), .A2(n9884), .ZN(n9881) );
  NOR2_X1 U9742 ( .A1(n9885), .A2(n9092), .ZN(n9879) );
  NOR2_X1 U9743 ( .A1(n9886), .A2(n9887), .ZN(n9875) );
  INV_X1 U9744 ( .A(n9878), .ZN(n9887) );
  XNOR2_X1 U9745 ( .A(a_3_), .B(n9888), .ZN(n9878) );
  NOR2_X1 U9746 ( .A1(n9889), .A2(n9890), .ZN(n9886) );
  NAND2_X1 U9747 ( .A1(n9891), .A2(n9892), .ZN(n9890) );
  INV_X1 U9748 ( .A(n9893), .ZN(n9892) );
  NOR2_X1 U9749 ( .A1(n9883), .A2(n9064), .ZN(n9893) );
  NAND2_X1 U9750 ( .A1(n9029), .A2(n9894), .ZN(n9891) );
  NOR2_X1 U9751 ( .A1(n9895), .A2(n9092), .ZN(n9889) );
  NAND2_X1 U9752 ( .A1(n9896), .A2(n9897), .ZN(Result_34_) );
  NAND2_X1 U9753 ( .A1(n9027), .A2(n9898), .ZN(n9897) );
  XNOR2_X1 U9754 ( .A(n9899), .B(n9900), .ZN(n9898) );
  XOR2_X1 U9755 ( .A(n9901), .B(n9902), .Z(n9900) );
  NAND2_X1 U9756 ( .A1(a_2_), .A2(b_31_), .ZN(n9902) );
  NOR2_X1 U9757 ( .A1(n9903), .A2(n9904), .ZN(n9896) );
  NOR2_X1 U9758 ( .A1(n9905), .A2(n9906), .ZN(n9904) );
  NOR2_X1 U9759 ( .A1(n9907), .A2(n9908), .ZN(n9905) );
  NAND2_X1 U9760 ( .A1(n9909), .A2(n9910), .ZN(n9908) );
  INV_X1 U9761 ( .A(n9911), .ZN(n9910) );
  NOR2_X1 U9762 ( .A1(n9912), .A2(n9064), .ZN(n9911) );
  NAND2_X1 U9763 ( .A1(n9029), .A2(n9913), .ZN(n9909) );
  NOR2_X1 U9764 ( .A1(n9914), .A2(n9092), .ZN(n9907) );
  NOR2_X1 U9765 ( .A1(n9915), .A2(n9916), .ZN(n9903) );
  NOR2_X1 U9766 ( .A1(n9917), .A2(n9918), .ZN(n9916) );
  NAND2_X1 U9767 ( .A1(n9919), .A2(n9920), .ZN(n9918) );
  NAND2_X1 U9768 ( .A1(n9091), .A2(n9912), .ZN(n9920) );
  NAND2_X1 U9769 ( .A1(n9029), .A2(n9921), .ZN(n9919) );
  NOR2_X1 U9770 ( .A1(n9922), .A2(n9092), .ZN(n9917) );
  INV_X1 U9771 ( .A(n9906), .ZN(n9915) );
  NAND2_X1 U9772 ( .A1(n9923), .A2(n9924), .ZN(n9906) );
  NAND2_X1 U9773 ( .A1(n9925), .A2(n9926), .ZN(Result_33_) );
  NAND2_X1 U9774 ( .A1(n9927), .A2(n9027), .ZN(n9926) );
  XNOR2_X1 U9775 ( .A(n9928), .B(n9929), .ZN(n9927) );
  XOR2_X1 U9776 ( .A(n9930), .B(n9931), .Z(n9929) );
  NAND2_X1 U9777 ( .A1(a_1_), .A2(b_31_), .ZN(n9931) );
  NOR2_X1 U9778 ( .A1(n9932), .A2(n9933), .ZN(n9925) );
  NOR2_X1 U9779 ( .A1(n9934), .A2(n9935), .ZN(n9933) );
  NOR2_X1 U9780 ( .A1(n9936), .A2(n9937), .ZN(n9934) );
  NAND2_X1 U9781 ( .A1(n9938), .A2(n9939), .ZN(n9937) );
  NAND2_X1 U9782 ( .A1(n9940), .A2(n9091), .ZN(n9939) );
  NAND2_X1 U9783 ( .A1(n9029), .A2(n9941), .ZN(n9938) );
  NOR2_X1 U9784 ( .A1(n9942), .A2(n9092), .ZN(n9936) );
  NOR2_X1 U9785 ( .A1(n9943), .A2(n9944), .ZN(n9932) );
  NOR2_X1 U9786 ( .A1(n9945), .A2(n9946), .ZN(n9944) );
  NAND2_X1 U9787 ( .A1(n9947), .A2(n9948), .ZN(n9946) );
  NAND2_X1 U9788 ( .A1(n9091), .A2(n9949), .ZN(n9948) );
  NAND2_X1 U9789 ( .A1(n9029), .A2(n9950), .ZN(n9947) );
  NOR2_X1 U9790 ( .A1(n9951), .A2(n9092), .ZN(n9945) );
  INV_X1 U9791 ( .A(n9935), .ZN(n9943) );
  NAND2_X1 U9792 ( .A1(n9952), .A2(n9953), .ZN(n9935) );
  NAND2_X1 U9793 ( .A1(n9954), .A2(n9955), .ZN(Result_32_) );
  NAND2_X1 U9794 ( .A1(n9956), .A2(n9027), .ZN(n9955) );
  XNOR2_X1 U9795 ( .A(n9957), .B(n9958), .ZN(n9956) );
  XOR2_X1 U9796 ( .A(n9959), .B(n9960), .Z(n9958) );
  NAND2_X1 U9797 ( .A1(a_0_), .A2(b_31_), .ZN(n9960) );
  NOR2_X1 U9798 ( .A1(n9961), .A2(n9962), .ZN(n9954) );
  NOR2_X1 U9799 ( .A1(n9963), .A2(n9964), .ZN(n9962) );
  NOR2_X1 U9800 ( .A1(n9965), .A2(n9966), .ZN(n9963) );
  NAND2_X1 U9801 ( .A1(n9967), .A2(n9968), .ZN(n9966) );
  NAND2_X1 U9802 ( .A1(n9091), .A2(n9969), .ZN(n9968) );
  NAND2_X1 U9803 ( .A1(n9029), .A2(n9970), .ZN(n9967) );
  NOR2_X1 U9804 ( .A1(n9971), .A2(n9092), .ZN(n9965) );
  NOR2_X1 U9805 ( .A1(n9972), .A2(n9973), .ZN(n9961) );
  NOR2_X1 U9806 ( .A1(n9974), .A2(n9975), .ZN(n9973) );
  NAND2_X1 U9807 ( .A1(n9976), .A2(n9977), .ZN(n9975) );
  INV_X1 U9808 ( .A(n9978), .ZN(n9977) );
  NOR2_X1 U9809 ( .A1(n9969), .A2(n9064), .ZN(n9978) );
  NAND2_X1 U9810 ( .A1(n9981), .A2(n9953), .ZN(n9969) );
  NAND2_X1 U9811 ( .A1(n9982), .A2(n9983), .ZN(n9953) );
  NAND2_X1 U9812 ( .A1(n9940), .A2(n9952), .ZN(n9981) );
  INV_X1 U9813 ( .A(n9949), .ZN(n9940) );
  NAND2_X1 U9814 ( .A1(n9923), .A2(n9984), .ZN(n9949) );
  NAND2_X1 U9815 ( .A1(n9924), .A2(n9912), .ZN(n9984) );
  NAND2_X1 U9816 ( .A1(n9985), .A2(n9986), .ZN(n9912) );
  NAND2_X1 U9817 ( .A1(n9987), .A2(n9883), .ZN(n9986) );
  NAND2_X1 U9818 ( .A1(n9866), .A2(n9988), .ZN(n9883) );
  NAND2_X1 U9819 ( .A1(n9867), .A2(n9855), .ZN(n9988) );
  NAND2_X1 U9820 ( .A1(n9837), .A2(n9989), .ZN(n9855) );
  NAND2_X1 U9821 ( .A1(n9838), .A2(n9826), .ZN(n9989) );
  NAND2_X1 U9822 ( .A1(n9808), .A2(n9990), .ZN(n9826) );
  NAND2_X1 U9823 ( .A1(n9809), .A2(n9805), .ZN(n9990) );
  INV_X1 U9824 ( .A(n9796), .ZN(n9805) );
  NOR2_X1 U9825 ( .A1(n9991), .A2(n9992), .ZN(n9796) );
  NOR2_X1 U9826 ( .A1(n9993), .A2(n9778), .ZN(n9992) );
  INV_X1 U9827 ( .A(n9768), .ZN(n9778) );
  NAND2_X1 U9828 ( .A1(n9742), .A2(n9994), .ZN(n9768) );
  NAND2_X1 U9829 ( .A1(n9743), .A2(n9731), .ZN(n9994) );
  NAND2_X1 U9830 ( .A1(n9713), .A2(n9995), .ZN(n9731) );
  NAND2_X1 U9831 ( .A1(n9714), .A2(n9702), .ZN(n9995) );
  NAND2_X1 U9832 ( .A1(n9684), .A2(n9996), .ZN(n9702) );
  NAND2_X1 U9833 ( .A1(n9685), .A2(n9673), .ZN(n9996) );
  NAND2_X1 U9834 ( .A1(n9997), .A2(n9998), .ZN(n9673) );
  NAND2_X1 U9835 ( .A1(n9999), .A2(n9644), .ZN(n9998) );
  NAND2_X1 U9836 ( .A1(n9627), .A2(n10000), .ZN(n9644) );
  NAND2_X1 U9837 ( .A1(n9628), .A2(n9616), .ZN(n10000) );
  NAND2_X1 U9838 ( .A1(n9598), .A2(n10001), .ZN(n9616) );
  NAND2_X1 U9839 ( .A1(n9599), .A2(n9587), .ZN(n10001) );
  NAND2_X1 U9840 ( .A1(n9569), .A2(n10002), .ZN(n9587) );
  NAND2_X1 U9841 ( .A1(n9570), .A2(n9558), .ZN(n10002) );
  NAND2_X1 U9842 ( .A1(n10003), .A2(n10004), .ZN(n9558) );
  NAND2_X1 U9843 ( .A1(n10005), .A2(n9529), .ZN(n10004) );
  NAND2_X1 U9844 ( .A1(n9512), .A2(n10006), .ZN(n9529) );
  NAND2_X1 U9845 ( .A1(n9513), .A2(n9501), .ZN(n10006) );
  NAND2_X1 U9846 ( .A1(n9483), .A2(n10007), .ZN(n9501) );
  NAND2_X1 U9847 ( .A1(n9484), .A2(n9472), .ZN(n10007) );
  NAND2_X1 U9848 ( .A1(n9450), .A2(n10008), .ZN(n9472) );
  NAND2_X1 U9849 ( .A1(n9451), .A2(n9439), .ZN(n10008) );
  NAND2_X1 U9850 ( .A1(n10009), .A2(n10010), .ZN(n9439) );
  NAND2_X1 U9851 ( .A1(n10011), .A2(n9410), .ZN(n10010) );
  NAND2_X1 U9852 ( .A1(n9393), .A2(n10012), .ZN(n9410) );
  NAND2_X1 U9853 ( .A1(n9394), .A2(n9382), .ZN(n10012) );
  NAND2_X1 U9854 ( .A1(n10013), .A2(n10014), .ZN(n9382) );
  NAND2_X1 U9855 ( .A1(n10015), .A2(n9353), .ZN(n10014) );
  INV_X1 U9856 ( .A(n9363), .ZN(n9353) );
  NOR2_X1 U9857 ( .A1(n10016), .A2(n10017), .ZN(n9363) );
  NOR2_X1 U9858 ( .A1(n10018), .A2(n9335), .ZN(n10017) );
  INV_X1 U9859 ( .A(n9325), .ZN(n9335) );
  NAND2_X1 U9860 ( .A1(n10019), .A2(n10020), .ZN(n9325) );
  NAND2_X1 U9861 ( .A1(n10021), .A2(n9297), .ZN(n10020) );
  NAND2_X1 U9862 ( .A1(n10022), .A2(n10023), .ZN(n9297) );
  NAND2_X1 U9863 ( .A1(n10024), .A2(n9268), .ZN(n10023) );
  NAND2_X1 U9864 ( .A1(n10025), .A2(n10026), .ZN(n9268) );
  NAND2_X1 U9865 ( .A1(n10027), .A2(n9240), .ZN(n10026) );
  NAND2_X1 U9866 ( .A1(n10028), .A2(n10029), .ZN(n9240) );
  NAND2_X1 U9867 ( .A1(n10030), .A2(n9212), .ZN(n10029) );
  INV_X1 U9868 ( .A(n9222), .ZN(n9212) );
  NOR2_X1 U9869 ( .A1(n10031), .A2(n10032), .ZN(n9222) );
  NOR2_X1 U9870 ( .A1(n10033), .A2(n9184), .ZN(n10032) );
  NOR2_X1 U9871 ( .A1(n10034), .A2(n10035), .ZN(n9184) );
  NOR2_X1 U9872 ( .A1(n10036), .A2(n9154), .ZN(n10035) );
  INV_X1 U9873 ( .A(n9145), .ZN(n9154) );
  NAND2_X1 U9874 ( .A1(n10037), .A2(n10038), .ZN(n9145) );
  NAND2_X1 U9875 ( .A1(n10039), .A2(n9116), .ZN(n10038) );
  NAND2_X1 U9876 ( .A1(n10040), .A2(n10041), .ZN(n9116) );
  NAND2_X1 U9877 ( .A1(b_30_), .A2(n10042), .ZN(n10041) );
  NAND2_X1 U9878 ( .A1(n10043), .A2(n9099), .ZN(n10042) );
  INV_X1 U9879 ( .A(n9060), .ZN(n9099) );
  NOR2_X1 U9880 ( .A1(n10044), .A2(n9077), .ZN(n9060) );
  NAND2_X1 U9881 ( .A1(n9025), .A2(b_31_), .ZN(n10040) );
  NAND2_X1 U9882 ( .A1(n10046), .A2(n9121), .ZN(n10039) );
  NOR2_X1 U9883 ( .A1(b_28_), .A2(a_28_), .ZN(n10036) );
  NOR2_X1 U9884 ( .A1(b_27_), .A2(a_27_), .ZN(n10033) );
  NAND2_X1 U9885 ( .A1(n9217), .A2(n10047), .ZN(n10030) );
  NAND2_X1 U9886 ( .A1(n9245), .A2(n10048), .ZN(n10027) );
  NAND2_X1 U9887 ( .A1(n10049), .A2(n10050), .ZN(n10024) );
  NAND2_X1 U9888 ( .A1(n9302), .A2(n10051), .ZN(n10021) );
  NOR2_X1 U9889 ( .A1(b_22_), .A2(a_22_), .ZN(n10018) );
  NAND2_X1 U9890 ( .A1(n10052), .A2(n9358), .ZN(n10015) );
  NAND2_X1 U9891 ( .A1(n10053), .A2(n10054), .ZN(n9394) );
  INV_X1 U9892 ( .A(n10055), .ZN(n9393) );
  NAND2_X1 U9893 ( .A1(n10056), .A2(n9415), .ZN(n10011) );
  NAND2_X1 U9894 ( .A1(n10057), .A2(n10058), .ZN(n9451) );
  NAND2_X1 U9895 ( .A1(n10059), .A2(n10060), .ZN(n9484) );
  NAND2_X1 U9896 ( .A1(n10061), .A2(n10062), .ZN(n9513) );
  NAND2_X1 U9897 ( .A1(n10063), .A2(n9534), .ZN(n10005) );
  NAND2_X1 U9898 ( .A1(n10064), .A2(n10065), .ZN(n9570) );
  NAND2_X1 U9899 ( .A1(n10066), .A2(n10067), .ZN(n9599) );
  INV_X1 U9900 ( .A(n10068), .ZN(n9598) );
  NAND2_X1 U9901 ( .A1(n10069), .A2(n10070), .ZN(n9628) );
  NAND2_X1 U9902 ( .A1(n10071), .A2(n9649), .ZN(n9999) );
  NAND2_X1 U9903 ( .A1(n10072), .A2(n10073), .ZN(n9685) );
  INV_X1 U9904 ( .A(n10074), .ZN(n9684) );
  NAND2_X1 U9905 ( .A1(n10075), .A2(n10076), .ZN(n9714) );
  INV_X1 U9906 ( .A(n10077), .ZN(n9713) );
  NAND2_X1 U9907 ( .A1(n10078), .A2(n10079), .ZN(n9743) );
  NOR2_X1 U9908 ( .A1(b_7_), .A2(a_7_), .ZN(n9993) );
  NAND2_X1 U9909 ( .A1(n10080), .A2(n10081), .ZN(n9809) );
  NAND2_X1 U9910 ( .A1(n10082), .A2(n10083), .ZN(n9838) );
  NAND2_X1 U9911 ( .A1(n10084), .A2(n10085), .ZN(n9867) );
  NAND2_X1 U9912 ( .A1(n9888), .A2(n10086), .ZN(n9987) );
  NAND2_X1 U9913 ( .A1(n10087), .A2(n10088), .ZN(n9924) );
  NAND2_X1 U9914 ( .A1(n9029), .A2(n10089), .ZN(n9976) );
  NOR2_X1 U9915 ( .A1(n10090), .A2(n9092), .ZN(n9974) );
  INV_X1 U9916 ( .A(n9964), .ZN(n9972) );
  NAND2_X1 U9917 ( .A1(n10091), .A2(n10092), .ZN(n9964) );
  NAND2_X1 U9918 ( .A1(n10093), .A2(n10094), .ZN(n10092) );
  NAND2_X1 U9919 ( .A1(n9030), .A2(n10095), .ZN(Result_31_) );
  NAND2_X1 U9920 ( .A1(n10096), .A2(n9027), .ZN(n10095) );
  XNOR2_X1 U9921 ( .A(n10097), .B(n10098), .ZN(n10096) );
  NAND2_X1 U9922 ( .A1(n9030), .A2(n10099), .ZN(Result_30_) );
  NAND2_X1 U9923 ( .A1(n10100), .A2(n9027), .ZN(n10099) );
  NOR2_X1 U9924 ( .A1(n10101), .A2(n10102), .ZN(n10100) );
  NOR2_X1 U9925 ( .A1(n10103), .A2(n10104), .ZN(n10102) );
  NOR2_X1 U9926 ( .A1(n10105), .A2(n10098), .ZN(n10103) );
  INV_X1 U9927 ( .A(n10097), .ZN(n10105) );
  NAND2_X1 U9928 ( .A1(n9030), .A2(n10106), .ZN(Result_2_) );
  NAND2_X1 U9929 ( .A1(n10107), .A2(n9027), .ZN(n10106) );
  XOR2_X1 U9930 ( .A(n10108), .B(n10109), .Z(n10107) );
  NAND2_X1 U9931 ( .A1(n9030), .A2(n10110), .ZN(Result_29_) );
  NAND2_X1 U9932 ( .A1(n9027), .A2(n10111), .ZN(n10110) );
  XNOR2_X1 U9933 ( .A(n10101), .B(n10112), .ZN(n10111) );
  NAND2_X1 U9934 ( .A1(n10113), .A2(n10114), .ZN(n10112) );
  NAND2_X1 U9935 ( .A1(n9030), .A2(n10115), .ZN(Result_28_) );
  NAND2_X1 U9936 ( .A1(n10116), .A2(n9027), .ZN(n10115) );
  XNOR2_X1 U9937 ( .A(n10117), .B(n10118), .ZN(n10116) );
  NAND2_X1 U9938 ( .A1(n10119), .A2(n10120), .ZN(n10118) );
  NAND2_X1 U9939 ( .A1(n9030), .A2(n10121), .ZN(Result_27_) );
  NAND2_X1 U9940 ( .A1(n10122), .A2(n9027), .ZN(n10121) );
  XNOR2_X1 U9941 ( .A(n10123), .B(n10124), .ZN(n10122) );
  NAND2_X1 U9942 ( .A1(n10125), .A2(n10126), .ZN(n10124) );
  NAND2_X1 U9943 ( .A1(n9030), .A2(n10127), .ZN(Result_26_) );
  NAND2_X1 U9944 ( .A1(n10128), .A2(n9027), .ZN(n10127) );
  XNOR2_X1 U9945 ( .A(n10129), .B(n10130), .ZN(n10128) );
  NAND2_X1 U9946 ( .A1(n10131), .A2(n10132), .ZN(n10130) );
  NAND2_X1 U9947 ( .A1(n9030), .A2(n10133), .ZN(Result_25_) );
  NAND2_X1 U9948 ( .A1(n10134), .A2(n9027), .ZN(n10133) );
  XOR2_X1 U9949 ( .A(n10135), .B(n10136), .Z(n10134) );
  NOR2_X1 U9950 ( .A1(n10137), .A2(n10138), .ZN(n10136) );
  NOR2_X1 U9951 ( .A1(n10139), .A2(n10140), .ZN(n10138) );
  INV_X1 U9952 ( .A(n10141), .ZN(n10137) );
  NAND2_X1 U9953 ( .A1(n9030), .A2(n10142), .ZN(Result_24_) );
  NAND2_X1 U9954 ( .A1(n10143), .A2(n9027), .ZN(n10142) );
  XNOR2_X1 U9955 ( .A(n10144), .B(n10145), .ZN(n10143) );
  NAND2_X1 U9956 ( .A1(n10146), .A2(n10147), .ZN(n10145) );
  NAND2_X1 U9957 ( .A1(n9030), .A2(n10148), .ZN(Result_23_) );
  NAND2_X1 U9958 ( .A1(n10149), .A2(n9027), .ZN(n10148) );
  XNOR2_X1 U9959 ( .A(n10150), .B(n10151), .ZN(n10149) );
  NAND2_X1 U9960 ( .A1(n10152), .A2(n10153), .ZN(n10151) );
  NAND2_X1 U9961 ( .A1(n9030), .A2(n10154), .ZN(Result_22_) );
  NAND2_X1 U9962 ( .A1(n10155), .A2(n9027), .ZN(n10154) );
  XNOR2_X1 U9963 ( .A(n10156), .B(n10157), .ZN(n10155) );
  NAND2_X1 U9964 ( .A1(n10158), .A2(n10159), .ZN(n10157) );
  NAND2_X1 U9965 ( .A1(n9030), .A2(n10160), .ZN(Result_21_) );
  NAND2_X1 U9966 ( .A1(n10161), .A2(n9027), .ZN(n10160) );
  XNOR2_X1 U9967 ( .A(n10162), .B(n10163), .ZN(n10161) );
  NAND2_X1 U9968 ( .A1(n10164), .A2(n10165), .ZN(n10163) );
  NAND2_X1 U9969 ( .A1(n9030), .A2(n10166), .ZN(Result_20_) );
  NAND2_X1 U9970 ( .A1(n10167), .A2(n9027), .ZN(n10166) );
  XNOR2_X1 U9971 ( .A(n10168), .B(n10169), .ZN(n10167) );
  NAND2_X1 U9972 ( .A1(n10170), .A2(n10171), .ZN(n10169) );
  NAND2_X1 U9973 ( .A1(n9030), .A2(n10172), .ZN(Result_1_) );
  NAND2_X1 U9974 ( .A1(n9027), .A2(n10173), .ZN(n10172) );
  XNOR2_X1 U9975 ( .A(n10174), .B(n10175), .ZN(n10173) );
  NOR2_X1 U9976 ( .A1(n10176), .A2(n10177), .ZN(n10175) );
  NAND2_X1 U9977 ( .A1(n9030), .A2(n10178), .ZN(Result_19_) );
  NAND2_X1 U9978 ( .A1(n10179), .A2(n9027), .ZN(n10178) );
  XNOR2_X1 U9979 ( .A(n10180), .B(n10181), .ZN(n10179) );
  NAND2_X1 U9980 ( .A1(n10182), .A2(n10183), .ZN(n10181) );
  NAND2_X1 U9981 ( .A1(n9030), .A2(n10184), .ZN(Result_18_) );
  NAND2_X1 U9982 ( .A1(n10185), .A2(n9027), .ZN(n10184) );
  XNOR2_X1 U9983 ( .A(n10186), .B(n10187), .ZN(n10185) );
  NAND2_X1 U9984 ( .A1(n10188), .A2(n10189), .ZN(n10187) );
  NAND2_X1 U9985 ( .A1(n9030), .A2(n10190), .ZN(Result_17_) );
  NAND2_X1 U9986 ( .A1(n10191), .A2(n9027), .ZN(n10190) );
  XOR2_X1 U9987 ( .A(n10192), .B(n10193), .Z(n10191) );
  NOR2_X1 U9988 ( .A1(n10194), .A2(n10195), .ZN(n10193) );
  INV_X1 U9989 ( .A(n10196), .ZN(n10195) );
  NOR2_X1 U9990 ( .A1(n10197), .A2(n10198), .ZN(n10194) );
  NAND2_X1 U9991 ( .A1(n9030), .A2(n10199), .ZN(Result_16_) );
  NAND2_X1 U9992 ( .A1(n10200), .A2(n9027), .ZN(n10199) );
  XNOR2_X1 U9993 ( .A(n10201), .B(n10202), .ZN(n10200) );
  NAND2_X1 U9994 ( .A1(n10203), .A2(n10204), .ZN(n10202) );
  NAND2_X1 U9995 ( .A1(n9030), .A2(n10205), .ZN(Result_15_) );
  NAND2_X1 U9996 ( .A1(n10206), .A2(n9027), .ZN(n10205) );
  XOR2_X1 U9997 ( .A(n10207), .B(n10208), .Z(n10206) );
  NOR2_X1 U9998 ( .A1(n10209), .A2(n10210), .ZN(n10208) );
  INV_X1 U9999 ( .A(n10211), .ZN(n10210) );
  NOR2_X1 U10000 ( .A1(n10212), .A2(n10213), .ZN(n10209) );
  NAND2_X1 U10001 ( .A1(n9030), .A2(n10214), .ZN(Result_14_) );
  NAND2_X1 U10002 ( .A1(n10215), .A2(n9027), .ZN(n10214) );
  XOR2_X1 U10003 ( .A(n10216), .B(n10217), .Z(n10215) );
  NAND2_X1 U10004 ( .A1(n9030), .A2(n10218), .ZN(Result_13_) );
  NAND2_X1 U10005 ( .A1(n9027), .A2(n10219), .ZN(n10218) );
  XOR2_X1 U10006 ( .A(n10220), .B(n10221), .Z(n10219) );
  NOR2_X1 U10007 ( .A1(n10222), .A2(n10223), .ZN(n10221) );
  INV_X1 U10008 ( .A(n10224), .ZN(n10223) );
  NOR2_X1 U10009 ( .A1(n10225), .A2(n10226), .ZN(n10222) );
  NAND2_X1 U10010 ( .A1(n9030), .A2(n10227), .ZN(Result_12_) );
  NAND2_X1 U10011 ( .A1(n9027), .A2(n10228), .ZN(n10227) );
  XOR2_X1 U10012 ( .A(n10229), .B(n10230), .Z(n10228) );
  NAND2_X1 U10013 ( .A1(n9030), .A2(n10231), .ZN(Result_11_) );
  NAND2_X1 U10014 ( .A1(n9027), .A2(n10232), .ZN(n10231) );
  XOR2_X1 U10015 ( .A(n10233), .B(n10234), .Z(n10232) );
  NOR2_X1 U10016 ( .A1(n10235), .A2(n10236), .ZN(n10234) );
  INV_X1 U10017 ( .A(n10237), .ZN(n10236) );
  NOR2_X1 U10018 ( .A1(n10238), .A2(n10239), .ZN(n10235) );
  NAND2_X1 U10019 ( .A1(n9030), .A2(n10240), .ZN(Result_10_) );
  NAND2_X1 U10020 ( .A1(n10241), .A2(n9027), .ZN(n10240) );
  XOR2_X1 U10021 ( .A(n10242), .B(n10243), .Z(n10241) );
  NAND2_X1 U10022 ( .A1(n9030), .A2(n10244), .ZN(Result_0_) );
  NAND2_X1 U10023 ( .A1(n9027), .A2(n10245), .ZN(n10244) );
  NAND2_X1 U10024 ( .A1(n10246), .A2(n10247), .ZN(n10245) );
  NAND2_X1 U10025 ( .A1(a_0_), .A2(n10248), .ZN(n10247) );
  NOR2_X1 U10026 ( .A1(n10177), .A2(n10249), .ZN(n10246) );
  NOR2_X1 U10027 ( .A1(n10176), .A2(n10174), .ZN(n10249) );
  INV_X1 U10028 ( .A(n10250), .ZN(n10174) );
  NOR2_X1 U10029 ( .A1(n10108), .A2(n10109), .ZN(n10250) );
  NOR2_X1 U10030 ( .A1(n10251), .A2(n10252), .ZN(n10109) );
  NAND2_X1 U10031 ( .A1(n9750), .A2(n10253), .ZN(n10251) );
  NAND2_X1 U10032 ( .A1(n9746), .A2(n9751), .ZN(n10253) );
  NOR2_X1 U10033 ( .A1(n9454), .A2(n9455), .ZN(n9746) );
  NOR2_X1 U10034 ( .A1(n10254), .A2(n10255), .ZN(n9455) );
  NAND2_X1 U10035 ( .A1(n9165), .A2(n10256), .ZN(n10254) );
  NAND2_X1 U10036 ( .A1(n9161), .A2(n9166), .ZN(n10256) );
  NOR2_X1 U10037 ( .A1(n9057), .A2(n9056), .ZN(n9161) );
  NOR2_X1 U10038 ( .A1(n10257), .A2(n10258), .ZN(n9056) );
  NAND2_X1 U10039 ( .A1(n9051), .A2(n10259), .ZN(n10257) );
  NAND2_X1 U10040 ( .A1(n9047), .A2(n9052), .ZN(n10259) );
  NOR2_X1 U10041 ( .A1(n9044), .A2(n9043), .ZN(n9047) );
  NOR2_X1 U10042 ( .A1(n10260), .A2(n10261), .ZN(n9043) );
  NAND2_X1 U10043 ( .A1(n9038), .A2(n10262), .ZN(n10260) );
  NAND2_X1 U10044 ( .A1(n9034), .A2(n9039), .ZN(n10262) );
  NOR2_X1 U10045 ( .A1(n10242), .A2(n10243), .ZN(n9034) );
  NOR2_X1 U10046 ( .A1(n10263), .A2(n10264), .ZN(n10243) );
  NAND2_X1 U10047 ( .A1(n10237), .A2(n10265), .ZN(n10264) );
  NAND2_X1 U10048 ( .A1(n10238), .A2(n10233), .ZN(n10265) );
  NOR2_X1 U10049 ( .A1(n10230), .A2(n10229), .ZN(n10233) );
  NOR2_X1 U10050 ( .A1(n10266), .A2(n10267), .ZN(n10229) );
  NAND2_X1 U10051 ( .A1(n10224), .A2(n10268), .ZN(n10267) );
  NAND2_X1 U10052 ( .A1(n10225), .A2(n10220), .ZN(n10268) );
  NOR2_X1 U10053 ( .A1(n10216), .A2(n10217), .ZN(n10220) );
  NOR2_X1 U10054 ( .A1(n10269), .A2(n10270), .ZN(n10217) );
  NAND2_X1 U10055 ( .A1(n10211), .A2(n10271), .ZN(n10270) );
  NAND2_X1 U10056 ( .A1(n10212), .A2(n10207), .ZN(n10271) );
  NAND2_X1 U10057 ( .A1(n10272), .A2(n10203), .ZN(n10207) );
  NAND2_X1 U10058 ( .A1(n10273), .A2(n10274), .ZN(n10203) );
  NAND2_X1 U10059 ( .A1(n10204), .A2(n10201), .ZN(n10272) );
  NAND2_X1 U10060 ( .A1(n10196), .A2(n10275), .ZN(n10201) );
  NAND2_X1 U10061 ( .A1(n10197), .A2(n10192), .ZN(n10275) );
  NAND2_X1 U10062 ( .A1(n10276), .A2(n10188), .ZN(n10192) );
  NAND2_X1 U10063 ( .A1(n10277), .A2(n10278), .ZN(n10188) );
  NAND2_X1 U10064 ( .A1(n10186), .A2(n10189), .ZN(n10276) );
  INV_X1 U10065 ( .A(n10279), .ZN(n10189) );
  NOR2_X1 U10066 ( .A1(n10277), .A2(n10278), .ZN(n10279) );
  XOR2_X1 U10067 ( .A(n10280), .B(n10281), .Z(n10277) );
  NAND2_X1 U10068 ( .A1(n10183), .A2(n10282), .ZN(n10186) );
  NAND2_X1 U10069 ( .A1(n10180), .A2(n10182), .ZN(n10282) );
  NAND2_X1 U10070 ( .A1(n10283), .A2(n10284), .ZN(n10182) );
  NAND2_X1 U10071 ( .A1(n10170), .A2(n10285), .ZN(n10180) );
  NAND2_X1 U10072 ( .A1(n10168), .A2(n10171), .ZN(n10285) );
  NAND2_X1 U10073 ( .A1(n10286), .A2(n10287), .ZN(n10171) );
  XNOR2_X1 U10074 ( .A(n10288), .B(n10289), .ZN(n10286) );
  NAND2_X1 U10075 ( .A1(n10164), .A2(n10290), .ZN(n10168) );
  NAND2_X1 U10076 ( .A1(n10165), .A2(n10162), .ZN(n10290) );
  NAND2_X1 U10077 ( .A1(n10159), .A2(n10291), .ZN(n10162) );
  NAND2_X1 U10078 ( .A1(n10156), .A2(n10158), .ZN(n10291) );
  NAND2_X1 U10079 ( .A1(n10292), .A2(n10293), .ZN(n10158) );
  XNOR2_X1 U10080 ( .A(n10294), .B(n10295), .ZN(n10292) );
  NAND2_X1 U10081 ( .A1(n10153), .A2(n10296), .ZN(n10156) );
  NAND2_X1 U10082 ( .A1(n10150), .A2(n10152), .ZN(n10296) );
  NAND2_X1 U10083 ( .A1(n10297), .A2(n10298), .ZN(n10152) );
  NAND2_X1 U10084 ( .A1(n10146), .A2(n10299), .ZN(n10150) );
  NAND2_X1 U10085 ( .A1(n10144), .A2(n10147), .ZN(n10299) );
  NAND2_X1 U10086 ( .A1(n10300), .A2(n10301), .ZN(n10147) );
  XNOR2_X1 U10087 ( .A(n10302), .B(n10303), .ZN(n10300) );
  NAND2_X1 U10088 ( .A1(n10141), .A2(n10304), .ZN(n10144) );
  NAND2_X1 U10089 ( .A1(n10140), .A2(n10135), .ZN(n10304) );
  NAND2_X1 U10090 ( .A1(n10305), .A2(n10131), .ZN(n10135) );
  NAND2_X1 U10091 ( .A1(n10306), .A2(n10307), .ZN(n10131) );
  INV_X1 U10092 ( .A(n10308), .ZN(n10307) );
  NAND2_X1 U10093 ( .A1(n10129), .A2(n10132), .ZN(n10305) );
  NAND2_X1 U10094 ( .A1(n10309), .A2(n10308), .ZN(n10132) );
  INV_X1 U10095 ( .A(n10306), .ZN(n10309) );
  XOR2_X1 U10096 ( .A(n10310), .B(n10311), .Z(n10306) );
  NAND2_X1 U10097 ( .A1(n10125), .A2(n10312), .ZN(n10129) );
  NAND2_X1 U10098 ( .A1(n10123), .A2(n10126), .ZN(n10312) );
  NAND2_X1 U10099 ( .A1(n10313), .A2(n10314), .ZN(n10126) );
  NAND2_X1 U10100 ( .A1(n10120), .A2(n10315), .ZN(n10123) );
  NAND2_X1 U10101 ( .A1(n10117), .A2(n10119), .ZN(n10315) );
  NAND2_X1 U10102 ( .A1(n10316), .A2(n10317), .ZN(n10119) );
  NAND2_X1 U10103 ( .A1(n10113), .A2(n10318), .ZN(n10117) );
  NAND2_X1 U10104 ( .A1(n10101), .A2(n10114), .ZN(n10318) );
  NAND2_X1 U10105 ( .A1(n10319), .A2(n10320), .ZN(n10114) );
  NOR2_X1 U10106 ( .A1(n10321), .A2(n10098), .ZN(n10101) );
  XNOR2_X1 U10107 ( .A(n10322), .B(n10323), .ZN(n10098) );
  XOR2_X1 U10108 ( .A(n10324), .B(n10325), .Z(n10322) );
  NOR2_X1 U10109 ( .A1(n9080), .A2(n10093), .ZN(n10325) );
  NAND2_X1 U10110 ( .A1(n10097), .A2(n10104), .ZN(n10321) );
  XOR2_X1 U10111 ( .A(n10326), .B(n10327), .Z(n10104) );
  NAND2_X1 U10112 ( .A1(n10328), .A2(n10329), .ZN(n10097) );
  NAND2_X1 U10113 ( .A1(n10330), .A2(a_0_), .ZN(n10329) );
  NOR2_X1 U10114 ( .A1(n10331), .A2(n9077), .ZN(n10330) );
  NOR2_X1 U10115 ( .A1(n9957), .A2(n9959), .ZN(n10331) );
  NAND2_X1 U10116 ( .A1(n9957), .A2(n9959), .ZN(n10328) );
  NAND2_X1 U10117 ( .A1(n10332), .A2(n10333), .ZN(n9959) );
  NAND2_X1 U10118 ( .A1(n10334), .A2(a_1_), .ZN(n10333) );
  NOR2_X1 U10119 ( .A1(n10335), .A2(n9077), .ZN(n10334) );
  NOR2_X1 U10120 ( .A1(n9928), .A2(n9930), .ZN(n10335) );
  NAND2_X1 U10121 ( .A1(n9928), .A2(n9930), .ZN(n10332) );
  NAND2_X1 U10122 ( .A1(n10336), .A2(n10337), .ZN(n9930) );
  NAND2_X1 U10123 ( .A1(n10338), .A2(a_2_), .ZN(n10337) );
  NOR2_X1 U10124 ( .A1(n10339), .A2(n9077), .ZN(n10338) );
  NOR2_X1 U10125 ( .A1(n9899), .A2(n9901), .ZN(n10339) );
  NAND2_X1 U10126 ( .A1(n9899), .A2(n9901), .ZN(n10336) );
  NAND2_X1 U10127 ( .A1(n10340), .A2(n10341), .ZN(n9901) );
  NAND2_X1 U10128 ( .A1(n10342), .A2(a_3_), .ZN(n10341) );
  NOR2_X1 U10129 ( .A1(n10343), .A2(n9077), .ZN(n10342) );
  NOR2_X1 U10130 ( .A1(n9871), .A2(n9873), .ZN(n10343) );
  NAND2_X1 U10131 ( .A1(n9871), .A2(n9873), .ZN(n10340) );
  NAND2_X1 U10132 ( .A1(n10344), .A2(n10345), .ZN(n9873) );
  NAND2_X1 U10133 ( .A1(n10346), .A2(a_4_), .ZN(n10345) );
  NOR2_X1 U10134 ( .A1(n10347), .A2(n9077), .ZN(n10346) );
  NOR2_X1 U10135 ( .A1(n9842), .A2(n9844), .ZN(n10347) );
  NAND2_X1 U10136 ( .A1(n9842), .A2(n9844), .ZN(n10344) );
  NAND2_X1 U10137 ( .A1(n10348), .A2(n10349), .ZN(n9844) );
  NAND2_X1 U10138 ( .A1(n10350), .A2(a_5_), .ZN(n10349) );
  NOR2_X1 U10139 ( .A1(n10351), .A2(n9077), .ZN(n10350) );
  NOR2_X1 U10140 ( .A1(n9813), .A2(n9815), .ZN(n10351) );
  NAND2_X1 U10141 ( .A1(n9813), .A2(n9815), .ZN(n10348) );
  NAND2_X1 U10142 ( .A1(n10352), .A2(n10353), .ZN(n9815) );
  NAND2_X1 U10143 ( .A1(n10354), .A2(a_6_), .ZN(n10353) );
  NOR2_X1 U10144 ( .A1(n10355), .A2(n9077), .ZN(n10354) );
  NOR2_X1 U10145 ( .A1(n9784), .A2(n9786), .ZN(n10355) );
  NAND2_X1 U10146 ( .A1(n9784), .A2(n9786), .ZN(n10352) );
  NAND2_X1 U10147 ( .A1(n10356), .A2(n10357), .ZN(n9786) );
  NAND2_X1 U10148 ( .A1(n10358), .A2(a_7_), .ZN(n10357) );
  NOR2_X1 U10149 ( .A1(n10359), .A2(n9077), .ZN(n10358) );
  NOR2_X1 U10150 ( .A1(n9756), .A2(n9758), .ZN(n10359) );
  NAND2_X1 U10151 ( .A1(n9756), .A2(n9758), .ZN(n10356) );
  NAND2_X1 U10152 ( .A1(n10360), .A2(n10361), .ZN(n9758) );
  NAND2_X1 U10153 ( .A1(n10362), .A2(a_8_), .ZN(n10361) );
  NOR2_X1 U10154 ( .A1(n10363), .A2(n9077), .ZN(n10362) );
  NOR2_X1 U10155 ( .A1(n9718), .A2(n9720), .ZN(n10363) );
  NAND2_X1 U10156 ( .A1(n9718), .A2(n9720), .ZN(n10360) );
  NAND2_X1 U10157 ( .A1(n10364), .A2(n10365), .ZN(n9720) );
  NAND2_X1 U10158 ( .A1(n10366), .A2(a_9_), .ZN(n10365) );
  NOR2_X1 U10159 ( .A1(n10367), .A2(n9077), .ZN(n10366) );
  NOR2_X1 U10160 ( .A1(n9689), .A2(n9691), .ZN(n10367) );
  NAND2_X1 U10161 ( .A1(n9689), .A2(n9691), .ZN(n10364) );
  NAND2_X1 U10162 ( .A1(n10368), .A2(n10369), .ZN(n9691) );
  NAND2_X1 U10163 ( .A1(n10370), .A2(a_10_), .ZN(n10369) );
  NOR2_X1 U10164 ( .A1(n10371), .A2(n9077), .ZN(n10370) );
  NOR2_X1 U10165 ( .A1(n9660), .A2(n9662), .ZN(n10371) );
  NAND2_X1 U10166 ( .A1(n9660), .A2(n9662), .ZN(n10368) );
  NAND2_X1 U10167 ( .A1(n10372), .A2(n10373), .ZN(n9662) );
  NAND2_X1 U10168 ( .A1(n10374), .A2(a_11_), .ZN(n10373) );
  NOR2_X1 U10169 ( .A1(n10375), .A2(n9077), .ZN(n10374) );
  NOR2_X1 U10170 ( .A1(n9632), .A2(n9634), .ZN(n10375) );
  NAND2_X1 U10171 ( .A1(n9632), .A2(n9634), .ZN(n10372) );
  NAND2_X1 U10172 ( .A1(n10376), .A2(n10377), .ZN(n9634) );
  NAND2_X1 U10173 ( .A1(n10378), .A2(a_12_), .ZN(n10377) );
  NOR2_X1 U10174 ( .A1(n10379), .A2(n9077), .ZN(n10378) );
  NOR2_X1 U10175 ( .A1(n9603), .A2(n9605), .ZN(n10379) );
  NAND2_X1 U10176 ( .A1(n9603), .A2(n9605), .ZN(n10376) );
  NAND2_X1 U10177 ( .A1(n10380), .A2(n10381), .ZN(n9605) );
  NAND2_X1 U10178 ( .A1(n10382), .A2(a_13_), .ZN(n10381) );
  NOR2_X1 U10179 ( .A1(n10383), .A2(n9077), .ZN(n10382) );
  NOR2_X1 U10180 ( .A1(n9574), .A2(n9576), .ZN(n10383) );
  NAND2_X1 U10181 ( .A1(n9574), .A2(n9576), .ZN(n10380) );
  NAND2_X1 U10182 ( .A1(n10384), .A2(n10385), .ZN(n9576) );
  NAND2_X1 U10183 ( .A1(n10386), .A2(a_14_), .ZN(n10385) );
  NOR2_X1 U10184 ( .A1(n10387), .A2(n9077), .ZN(n10386) );
  NOR2_X1 U10185 ( .A1(n9545), .A2(n9547), .ZN(n10387) );
  NAND2_X1 U10186 ( .A1(n9545), .A2(n9547), .ZN(n10384) );
  NAND2_X1 U10187 ( .A1(n10388), .A2(n10389), .ZN(n9547) );
  NAND2_X1 U10188 ( .A1(n10390), .A2(a_15_), .ZN(n10389) );
  NOR2_X1 U10189 ( .A1(n10391), .A2(n9077), .ZN(n10390) );
  NOR2_X1 U10190 ( .A1(n9517), .A2(n9519), .ZN(n10391) );
  NAND2_X1 U10191 ( .A1(n9517), .A2(n9519), .ZN(n10388) );
  NAND2_X1 U10192 ( .A1(n10392), .A2(n10393), .ZN(n9519) );
  NAND2_X1 U10193 ( .A1(n10394), .A2(a_16_), .ZN(n10393) );
  NOR2_X1 U10194 ( .A1(n10395), .A2(n9077), .ZN(n10394) );
  NOR2_X1 U10195 ( .A1(n9488), .A2(n9490), .ZN(n10395) );
  NAND2_X1 U10196 ( .A1(n9488), .A2(n9490), .ZN(n10392) );
  NAND2_X1 U10197 ( .A1(n10396), .A2(n10397), .ZN(n9490) );
  NAND2_X1 U10198 ( .A1(n10398), .A2(a_17_), .ZN(n10397) );
  NOR2_X1 U10199 ( .A1(n10399), .A2(n9077), .ZN(n10398) );
  NOR2_X1 U10200 ( .A1(n9461), .A2(n9459), .ZN(n10399) );
  NAND2_X1 U10201 ( .A1(n9461), .A2(n9459), .ZN(n10396) );
  XNOR2_X1 U10202 ( .A(n10400), .B(n10401), .ZN(n9459) );
  NAND2_X1 U10203 ( .A1(n10402), .A2(n10403), .ZN(n10400) );
  NOR2_X1 U10204 ( .A1(n10404), .A2(n10405), .ZN(n9461) );
  NOR2_X1 U10205 ( .A1(n9427), .A2(n10406), .ZN(n10405) );
  NOR2_X1 U10206 ( .A1(n9428), .A2(n9429), .ZN(n10406) );
  XNOR2_X1 U10207 ( .A(n10407), .B(n10408), .ZN(n9427) );
  XNOR2_X1 U10208 ( .A(n10409), .B(n10410), .ZN(n10407) );
  NOR2_X1 U10209 ( .A1(n9080), .A2(n9415), .ZN(n10410) );
  INV_X1 U10210 ( .A(n10411), .ZN(n10404) );
  NAND2_X1 U10211 ( .A1(n9429), .A2(n9428), .ZN(n10411) );
  NAND2_X1 U10212 ( .A1(a_18_), .A2(b_31_), .ZN(n9428) );
  NOR2_X1 U10213 ( .A1(n10412), .A2(n10413), .ZN(n9429) );
  INV_X1 U10214 ( .A(n10414), .ZN(n10413) );
  NAND2_X1 U10215 ( .A1(n9400), .A2(n10415), .ZN(n10414) );
  NAND2_X1 U10216 ( .A1(n9401), .A2(n9399), .ZN(n10415) );
  NOR2_X1 U10217 ( .A1(n9415), .A2(n9077), .ZN(n9400) );
  NOR2_X1 U10218 ( .A1(n9399), .A2(n9401), .ZN(n10412) );
  NOR2_X1 U10219 ( .A1(n10416), .A2(n10417), .ZN(n9401) );
  INV_X1 U10220 ( .A(n10418), .ZN(n10417) );
  NAND2_X1 U10221 ( .A1(n9371), .A2(n10419), .ZN(n10418) );
  NAND2_X1 U10222 ( .A1(n9372), .A2(n9369), .ZN(n10419) );
  NOR2_X1 U10223 ( .A1(n10054), .A2(n9077), .ZN(n9371) );
  NOR2_X1 U10224 ( .A1(n9369), .A2(n9372), .ZN(n10416) );
  INV_X1 U10225 ( .A(n10420), .ZN(n9372) );
  NAND2_X1 U10226 ( .A1(n9343), .A2(n10421), .ZN(n10420) );
  NAND2_X1 U10227 ( .A1(n9342), .A2(n9344), .ZN(n10421) );
  NAND2_X1 U10228 ( .A1(n10422), .A2(n10423), .ZN(n9344) );
  NAND2_X1 U10229 ( .A1(a_21_), .A2(b_31_), .ZN(n10422) );
  XNOR2_X1 U10230 ( .A(n10424), .B(n10425), .ZN(n9342) );
  XNOR2_X1 U10231 ( .A(n10426), .B(n10427), .ZN(n10424) );
  INV_X1 U10232 ( .A(n10428), .ZN(n9343) );
  NOR2_X1 U10233 ( .A1(n10423), .A2(n9358), .ZN(n10428) );
  NAND2_X1 U10234 ( .A1(n10429), .A2(n10430), .ZN(n10423) );
  NAND2_X1 U10235 ( .A1(n10431), .A2(n9315), .ZN(n10430) );
  NAND2_X1 U10236 ( .A1(a_22_), .A2(b_31_), .ZN(n9315) );
  NAND2_X1 U10237 ( .A1(n9313), .A2(n9316), .ZN(n10431) );
  INV_X1 U10238 ( .A(n10432), .ZN(n10429) );
  NOR2_X1 U10239 ( .A1(n9316), .A2(n9313), .ZN(n10432) );
  XOR2_X1 U10240 ( .A(n10433), .B(n10434), .Z(n9313) );
  XOR2_X1 U10241 ( .A(n10435), .B(n10436), .Z(n10433) );
  NOR2_X1 U10242 ( .A1(n9080), .A2(n10051), .ZN(n10436) );
  NAND2_X1 U10243 ( .A1(n10437), .A2(n10438), .ZN(n9316) );
  NAND2_X1 U10244 ( .A1(n9287), .A2(n10439), .ZN(n10438) );
  INV_X1 U10245 ( .A(n10440), .ZN(n10439) );
  NOR2_X1 U10246 ( .A1(n9288), .A2(n9285), .ZN(n10440) );
  NOR2_X1 U10247 ( .A1(n10051), .A2(n9077), .ZN(n9287) );
  NAND2_X1 U10248 ( .A1(n9285), .A2(n9288), .ZN(n10437) );
  NAND2_X1 U10249 ( .A1(n10441), .A2(n10442), .ZN(n9288) );
  NAND2_X1 U10250 ( .A1(n9259), .A2(n10443), .ZN(n10442) );
  INV_X1 U10251 ( .A(n10444), .ZN(n10443) );
  NOR2_X1 U10252 ( .A1(n9258), .A2(n9256), .ZN(n10444) );
  NOR2_X1 U10253 ( .A1(n10050), .A2(n9077), .ZN(n9259) );
  NAND2_X1 U10254 ( .A1(n9256), .A2(n9258), .ZN(n10441) );
  NAND2_X1 U10255 ( .A1(n9230), .A2(n10445), .ZN(n9258) );
  NAND2_X1 U10256 ( .A1(n9229), .A2(n9231), .ZN(n10445) );
  NAND2_X1 U10257 ( .A1(n10446), .A2(n10447), .ZN(n9231) );
  NAND2_X1 U10258 ( .A1(a_25_), .A2(b_31_), .ZN(n10447) );
  INV_X1 U10259 ( .A(n10448), .ZN(n10446) );
  XOR2_X1 U10260 ( .A(n10449), .B(n10450), .Z(n9229) );
  XNOR2_X1 U10261 ( .A(n10451), .B(n10452), .ZN(n10450) );
  NAND2_X1 U10262 ( .A1(a_25_), .A2(n10448), .ZN(n9230) );
  NAND2_X1 U10263 ( .A1(n10453), .A2(n10454), .ZN(n10448) );
  NAND2_X1 U10264 ( .A1(n9201), .A2(n10455), .ZN(n10454) );
  INV_X1 U10265 ( .A(n10456), .ZN(n10455) );
  NOR2_X1 U10266 ( .A1(n9203), .A2(n9202), .ZN(n10456) );
  XNOR2_X1 U10267 ( .A(n10457), .B(n10458), .ZN(n9201) );
  NAND2_X1 U10268 ( .A1(n10459), .A2(n10460), .ZN(n10457) );
  NAND2_X1 U10269 ( .A1(n9203), .A2(n9202), .ZN(n10453) );
  NOR2_X1 U10270 ( .A1(n10047), .A2(n9077), .ZN(n9202) );
  NOR2_X1 U10271 ( .A1(n10461), .A2(n10462), .ZN(n9203) );
  INV_X1 U10272 ( .A(n10463), .ZN(n10462) );
  NAND2_X1 U10273 ( .A1(n10464), .A2(n9173), .ZN(n10463) );
  NAND2_X1 U10274 ( .A1(b_31_), .A2(a_27_), .ZN(n9173) );
  NAND2_X1 U10275 ( .A1(n9171), .A2(n9174), .ZN(n10464) );
  NOR2_X1 U10276 ( .A1(n9174), .A2(n9171), .ZN(n10461) );
  XNOR2_X1 U10277 ( .A(n10465), .B(n10466), .ZN(n9171) );
  XOR2_X1 U10278 ( .A(n10467), .B(n10468), .Z(n10466) );
  NAND2_X1 U10279 ( .A1(b_30_), .A2(a_28_), .ZN(n10468) );
  NAND2_X1 U10280 ( .A1(n10469), .A2(n10470), .ZN(n9174) );
  NAND2_X1 U10281 ( .A1(n10471), .A2(b_31_), .ZN(n10470) );
  NOR2_X1 U10282 ( .A1(n10472), .A2(n9136), .ZN(n10471) );
  NOR2_X1 U10283 ( .A1(n9134), .A2(n9133), .ZN(n10472) );
  NAND2_X1 U10284 ( .A1(n9134), .A2(n9133), .ZN(n10469) );
  XOR2_X1 U10285 ( .A(n10473), .B(n10474), .Z(n9133) );
  NOR2_X1 U10286 ( .A1(n9080), .A2(n9121), .ZN(n10474) );
  XNOR2_X1 U10287 ( .A(n10475), .B(n10476), .ZN(n10473) );
  NOR2_X1 U10288 ( .A1(n10477), .A2(n10478), .ZN(n9134) );
  INV_X1 U10289 ( .A(n10479), .ZN(n10478) );
  NAND2_X1 U10290 ( .A1(n10480), .A2(n9106), .ZN(n10479) );
  NAND2_X1 U10291 ( .A1(a_29_), .A2(b_31_), .ZN(n9106) );
  NAND2_X1 U10292 ( .A1(n9104), .A2(n9107), .ZN(n10480) );
  NOR2_X1 U10293 ( .A1(n9107), .A2(n9104), .ZN(n10477) );
  INV_X1 U10294 ( .A(n10481), .ZN(n9104) );
  NAND2_X1 U10295 ( .A1(n10482), .A2(n9025), .ZN(n10481) );
  NOR2_X1 U10296 ( .A1(n9077), .A2(n9080), .ZN(n10482) );
  NAND2_X1 U10297 ( .A1(n10483), .A2(n10484), .ZN(n9107) );
  NAND2_X1 U10298 ( .A1(b_29_), .A2(n10485), .ZN(n10484) );
  NAND2_X1 U10299 ( .A1(n10486), .A2(n10487), .ZN(n10485) );
  NAND2_X1 U10300 ( .A1(a_31_), .A2(n9080), .ZN(n10487) );
  NAND2_X1 U10301 ( .A1(b_30_), .A2(n10488), .ZN(n10483) );
  NAND2_X1 U10302 ( .A1(n10489), .A2(n10490), .ZN(n10488) );
  NAND2_X1 U10303 ( .A1(a_30_), .A2(n10046), .ZN(n10490) );
  XOR2_X1 U10304 ( .A(n10491), .B(n10492), .Z(n9256) );
  XOR2_X1 U10305 ( .A(n10493), .B(n10494), .Z(n10492) );
  XOR2_X1 U10306 ( .A(n10495), .B(n10496), .Z(n9285) );
  XOR2_X1 U10307 ( .A(n10497), .B(n10498), .Z(n10495) );
  XOR2_X1 U10308 ( .A(n10499), .B(n10500), .Z(n9369) );
  NAND2_X1 U10309 ( .A1(n10501), .A2(n10502), .ZN(n10499) );
  XNOR2_X1 U10310 ( .A(n10503), .B(n10504), .ZN(n9399) );
  XNOR2_X1 U10311 ( .A(n10505), .B(n10506), .ZN(n10504) );
  XNOR2_X1 U10312 ( .A(n10507), .B(n10508), .ZN(n9488) );
  NAND2_X1 U10313 ( .A1(n10509), .A2(n10510), .ZN(n10507) );
  XNOR2_X1 U10314 ( .A(n10511), .B(n10512), .ZN(n9517) );
  NAND2_X1 U10315 ( .A1(n10513), .A2(n10514), .ZN(n10511) );
  XOR2_X1 U10316 ( .A(n10515), .B(n10516), .Z(n9545) );
  XOR2_X1 U10317 ( .A(n10517), .B(n10518), .Z(n10515) );
  NOR2_X1 U10318 ( .A1(n9080), .A2(n9534), .ZN(n10518) );
  XNOR2_X1 U10319 ( .A(n10519), .B(n10520), .ZN(n9574) );
  NAND2_X1 U10320 ( .A1(n10521), .A2(n10522), .ZN(n10519) );
  XNOR2_X1 U10321 ( .A(n10523), .B(n10524), .ZN(n9603) );
  NAND2_X1 U10322 ( .A1(n10525), .A2(n10526), .ZN(n10523) );
  XNOR2_X1 U10323 ( .A(n10527), .B(n10528), .ZN(n9632) );
  NAND2_X1 U10324 ( .A1(n10529), .A2(n10530), .ZN(n10527) );
  XOR2_X1 U10325 ( .A(n10531), .B(n10532), .Z(n9660) );
  XOR2_X1 U10326 ( .A(n10533), .B(n10534), .Z(n10531) );
  NOR2_X1 U10327 ( .A1(n9080), .A2(n9649), .ZN(n10534) );
  XOR2_X1 U10328 ( .A(n10535), .B(n10536), .Z(n9689) );
  XNOR2_X1 U10329 ( .A(n10537), .B(n10538), .ZN(n10536) );
  XNOR2_X1 U10330 ( .A(n10539), .B(n10540), .ZN(n9718) );
  XNOR2_X1 U10331 ( .A(n10541), .B(n10542), .ZN(n10539) );
  NOR2_X1 U10332 ( .A1(n9080), .A2(n10076), .ZN(n10542) );
  XNOR2_X1 U10333 ( .A(n10543), .B(n10544), .ZN(n9756) );
  NAND2_X1 U10334 ( .A1(n10545), .A2(n10546), .ZN(n10543) );
  XNOR2_X1 U10335 ( .A(n10547), .B(n10548), .ZN(n9784) );
  NAND2_X1 U10336 ( .A1(n10549), .A2(n10550), .ZN(n10547) );
  XNOR2_X1 U10337 ( .A(n10551), .B(n10552), .ZN(n9813) );
  NAND2_X1 U10338 ( .A1(n10553), .A2(n10554), .ZN(n10551) );
  XOR2_X1 U10339 ( .A(n10555), .B(n10556), .Z(n9842) );
  XOR2_X1 U10340 ( .A(n10557), .B(n10558), .Z(n10555) );
  NOR2_X1 U10341 ( .A1(n9080), .A2(n10083), .ZN(n10558) );
  XNOR2_X1 U10342 ( .A(n10559), .B(n10560), .ZN(n9871) );
  NAND2_X1 U10343 ( .A1(n10561), .A2(n10562), .ZN(n10559) );
  XNOR2_X1 U10344 ( .A(n10563), .B(n10564), .ZN(n9899) );
  NAND2_X1 U10345 ( .A1(n10565), .A2(n10566), .ZN(n10563) );
  XOR2_X1 U10346 ( .A(n10567), .B(n10568), .Z(n9928) );
  XNOR2_X1 U10347 ( .A(n10569), .B(n10570), .ZN(n10568) );
  XNOR2_X1 U10348 ( .A(n10571), .B(n10572), .ZN(n9957) );
  XNOR2_X1 U10349 ( .A(n10573), .B(n10574), .ZN(n10571) );
  INV_X1 U10350 ( .A(n10575), .ZN(n10113) );
  NOR2_X1 U10351 ( .A1(n10320), .A2(n10319), .ZN(n10575) );
  XNOR2_X1 U10352 ( .A(n10576), .B(n10577), .ZN(n10319) );
  NAND2_X1 U10353 ( .A1(n10327), .A2(n10326), .ZN(n10320) );
  NAND2_X1 U10354 ( .A1(n10578), .A2(n10579), .ZN(n10326) );
  NAND2_X1 U10355 ( .A1(n10580), .A2(a_0_), .ZN(n10579) );
  NOR2_X1 U10356 ( .A1(n10581), .A2(n9080), .ZN(n10580) );
  NOR2_X1 U10357 ( .A1(n10323), .A2(n10324), .ZN(n10581) );
  NAND2_X1 U10358 ( .A1(n10323), .A2(n10324), .ZN(n10578) );
  NAND2_X1 U10359 ( .A1(n10582), .A2(n10583), .ZN(n10324) );
  NAND2_X1 U10360 ( .A1(n10574), .A2(n10584), .ZN(n10583) );
  INV_X1 U10361 ( .A(n10585), .ZN(n10584) );
  NOR2_X1 U10362 ( .A1(n10572), .A2(n10573), .ZN(n10585) );
  NOR2_X1 U10363 ( .A1(n9983), .A2(n9080), .ZN(n10574) );
  NAND2_X1 U10364 ( .A1(n10573), .A2(n10572), .ZN(n10582) );
  XNOR2_X1 U10365 ( .A(n10586), .B(n10587), .ZN(n10572) );
  XNOR2_X1 U10366 ( .A(n10588), .B(n10589), .ZN(n10586) );
  NOR2_X1 U10367 ( .A1(n10590), .A2(n10591), .ZN(n10573) );
  INV_X1 U10368 ( .A(n10592), .ZN(n10591) );
  NAND2_X1 U10369 ( .A1(n10567), .A2(n10593), .ZN(n10592) );
  NAND2_X1 U10370 ( .A1(n10570), .A2(n10569), .ZN(n10593) );
  XOR2_X1 U10371 ( .A(n10594), .B(n10595), .Z(n10567) );
  NAND2_X1 U10372 ( .A1(n10596), .A2(n10597), .ZN(n10594) );
  NOR2_X1 U10373 ( .A1(n10569), .A2(n10570), .ZN(n10590) );
  NOR2_X1 U10374 ( .A1(n10088), .A2(n9080), .ZN(n10570) );
  NAND2_X1 U10375 ( .A1(n10565), .A2(n10598), .ZN(n10569) );
  NAND2_X1 U10376 ( .A1(n10564), .A2(n10566), .ZN(n10598) );
  NAND2_X1 U10377 ( .A1(n10599), .A2(n10600), .ZN(n10566) );
  NAND2_X1 U10378 ( .A1(a_3_), .A2(b_30_), .ZN(n10600) );
  INV_X1 U10379 ( .A(n10601), .ZN(n10599) );
  XOR2_X1 U10380 ( .A(n10602), .B(n10603), .Z(n10564) );
  XNOR2_X1 U10381 ( .A(n10604), .B(n10605), .ZN(n10603) );
  NAND2_X1 U10382 ( .A1(a_3_), .A2(n10601), .ZN(n10565) );
  NAND2_X1 U10383 ( .A1(n10561), .A2(n10606), .ZN(n10601) );
  NAND2_X1 U10384 ( .A1(n10560), .A2(n10562), .ZN(n10606) );
  NAND2_X1 U10385 ( .A1(n10607), .A2(n10608), .ZN(n10562) );
  NAND2_X1 U10386 ( .A1(a_4_), .A2(b_30_), .ZN(n10608) );
  INV_X1 U10387 ( .A(n10609), .ZN(n10607) );
  XOR2_X1 U10388 ( .A(n10610), .B(n10611), .Z(n10560) );
  XOR2_X1 U10389 ( .A(n10612), .B(n10613), .Z(n10610) );
  NOR2_X1 U10390 ( .A1(n10083), .A2(n10046), .ZN(n10613) );
  NAND2_X1 U10391 ( .A1(a_4_), .A2(n10609), .ZN(n10561) );
  NAND2_X1 U10392 ( .A1(n10614), .A2(n10615), .ZN(n10609) );
  NAND2_X1 U10393 ( .A1(n10616), .A2(a_5_), .ZN(n10615) );
  NOR2_X1 U10394 ( .A1(n10617), .A2(n9080), .ZN(n10616) );
  NOR2_X1 U10395 ( .A1(n10557), .A2(n10556), .ZN(n10617) );
  NAND2_X1 U10396 ( .A1(n10556), .A2(n10557), .ZN(n10614) );
  NAND2_X1 U10397 ( .A1(n10553), .A2(n10618), .ZN(n10557) );
  NAND2_X1 U10398 ( .A1(n10552), .A2(n10554), .ZN(n10618) );
  NAND2_X1 U10399 ( .A1(n10619), .A2(n10620), .ZN(n10554) );
  NAND2_X1 U10400 ( .A1(a_6_), .A2(b_30_), .ZN(n10620) );
  INV_X1 U10401 ( .A(n10621), .ZN(n10619) );
  XNOR2_X1 U10402 ( .A(n10622), .B(n10623), .ZN(n10552) );
  NAND2_X1 U10403 ( .A1(n10624), .A2(n10625), .ZN(n10622) );
  NAND2_X1 U10404 ( .A1(a_6_), .A2(n10621), .ZN(n10553) );
  NAND2_X1 U10405 ( .A1(n10549), .A2(n10626), .ZN(n10621) );
  NAND2_X1 U10406 ( .A1(n10548), .A2(n10550), .ZN(n10626) );
  NAND2_X1 U10407 ( .A1(n10627), .A2(n10628), .ZN(n10550) );
  NAND2_X1 U10408 ( .A1(a_7_), .A2(b_30_), .ZN(n10628) );
  INV_X1 U10409 ( .A(n10629), .ZN(n10627) );
  XNOR2_X1 U10410 ( .A(n10630), .B(n10631), .ZN(n10548) );
  NAND2_X1 U10411 ( .A1(n10632), .A2(n10633), .ZN(n10630) );
  NAND2_X1 U10412 ( .A1(a_7_), .A2(n10629), .ZN(n10549) );
  NAND2_X1 U10413 ( .A1(n10545), .A2(n10634), .ZN(n10629) );
  NAND2_X1 U10414 ( .A1(n10544), .A2(n10546), .ZN(n10634) );
  NAND2_X1 U10415 ( .A1(n10635), .A2(n10636), .ZN(n10546) );
  NAND2_X1 U10416 ( .A1(a_8_), .A2(b_30_), .ZN(n10636) );
  INV_X1 U10417 ( .A(n10637), .ZN(n10635) );
  XNOR2_X1 U10418 ( .A(n10638), .B(n10639), .ZN(n10544) );
  XNOR2_X1 U10419 ( .A(n10640), .B(n10641), .ZN(n10638) );
  NOR2_X1 U10420 ( .A1(n10076), .A2(n10046), .ZN(n10641) );
  NAND2_X1 U10421 ( .A1(a_8_), .A2(n10637), .ZN(n10545) );
  NAND2_X1 U10422 ( .A1(n10642), .A2(n10643), .ZN(n10637) );
  NAND2_X1 U10423 ( .A1(n10644), .A2(a_9_), .ZN(n10643) );
  NOR2_X1 U10424 ( .A1(n10645), .A2(n9080), .ZN(n10644) );
  NOR2_X1 U10425 ( .A1(n10541), .A2(n10540), .ZN(n10645) );
  NAND2_X1 U10426 ( .A1(n10540), .A2(n10541), .ZN(n10642) );
  NOR2_X1 U10427 ( .A1(n10646), .A2(n10647), .ZN(n10541) );
  INV_X1 U10428 ( .A(n10648), .ZN(n10647) );
  NAND2_X1 U10429 ( .A1(n10535), .A2(n10649), .ZN(n10648) );
  NAND2_X1 U10430 ( .A1(n10538), .A2(n10537), .ZN(n10649) );
  XNOR2_X1 U10431 ( .A(n10650), .B(n10651), .ZN(n10535) );
  XOR2_X1 U10432 ( .A(n10652), .B(n10653), .Z(n10650) );
  NOR2_X1 U10433 ( .A1(n9649), .A2(n10046), .ZN(n10653) );
  NOR2_X1 U10434 ( .A1(n10537), .A2(n10538), .ZN(n10646) );
  NOR2_X1 U10435 ( .A1(n10073), .A2(n9080), .ZN(n10538) );
  NAND2_X1 U10436 ( .A1(n10654), .A2(n10655), .ZN(n10537) );
  NAND2_X1 U10437 ( .A1(n10656), .A2(a_11_), .ZN(n10655) );
  NOR2_X1 U10438 ( .A1(n10657), .A2(n9080), .ZN(n10656) );
  NOR2_X1 U10439 ( .A1(n10532), .A2(n10533), .ZN(n10657) );
  NAND2_X1 U10440 ( .A1(n10532), .A2(n10533), .ZN(n10654) );
  NAND2_X1 U10441 ( .A1(n10529), .A2(n10658), .ZN(n10533) );
  NAND2_X1 U10442 ( .A1(n10528), .A2(n10530), .ZN(n10658) );
  NAND2_X1 U10443 ( .A1(n10659), .A2(n10660), .ZN(n10530) );
  NAND2_X1 U10444 ( .A1(a_12_), .A2(b_30_), .ZN(n10660) );
  INV_X1 U10445 ( .A(n10661), .ZN(n10659) );
  XNOR2_X1 U10446 ( .A(n10662), .B(n10663), .ZN(n10528) );
  NAND2_X1 U10447 ( .A1(n10664), .A2(n10665), .ZN(n10662) );
  NAND2_X1 U10448 ( .A1(a_12_), .A2(n10661), .ZN(n10529) );
  NAND2_X1 U10449 ( .A1(n10525), .A2(n10666), .ZN(n10661) );
  NAND2_X1 U10450 ( .A1(n10524), .A2(n10526), .ZN(n10666) );
  NAND2_X1 U10451 ( .A1(n10667), .A2(n10668), .ZN(n10526) );
  NAND2_X1 U10452 ( .A1(a_13_), .A2(b_30_), .ZN(n10668) );
  INV_X1 U10453 ( .A(n10669), .ZN(n10667) );
  XNOR2_X1 U10454 ( .A(n10670), .B(n10671), .ZN(n10524) );
  NAND2_X1 U10455 ( .A1(n10672), .A2(n10673), .ZN(n10670) );
  NAND2_X1 U10456 ( .A1(a_13_), .A2(n10669), .ZN(n10525) );
  NAND2_X1 U10457 ( .A1(n10521), .A2(n10674), .ZN(n10669) );
  NAND2_X1 U10458 ( .A1(n10520), .A2(n10522), .ZN(n10674) );
  NAND2_X1 U10459 ( .A1(n10675), .A2(n10676), .ZN(n10522) );
  NAND2_X1 U10460 ( .A1(a_14_), .A2(b_30_), .ZN(n10676) );
  INV_X1 U10461 ( .A(n10677), .ZN(n10675) );
  XOR2_X1 U10462 ( .A(n10678), .B(n10679), .Z(n10520) );
  XOR2_X1 U10463 ( .A(n10680), .B(n10681), .Z(n10678) );
  NOR2_X1 U10464 ( .A1(n9534), .A2(n10046), .ZN(n10681) );
  NAND2_X1 U10465 ( .A1(a_14_), .A2(n10677), .ZN(n10521) );
  NAND2_X1 U10466 ( .A1(n10682), .A2(n10683), .ZN(n10677) );
  NAND2_X1 U10467 ( .A1(n10684), .A2(a_15_), .ZN(n10683) );
  NOR2_X1 U10468 ( .A1(n10685), .A2(n9080), .ZN(n10684) );
  NOR2_X1 U10469 ( .A1(n10517), .A2(n10516), .ZN(n10685) );
  NAND2_X1 U10470 ( .A1(n10516), .A2(n10517), .ZN(n10682) );
  NAND2_X1 U10471 ( .A1(n10513), .A2(n10686), .ZN(n10517) );
  NAND2_X1 U10472 ( .A1(n10512), .A2(n10514), .ZN(n10686) );
  NAND2_X1 U10473 ( .A1(n10687), .A2(n10688), .ZN(n10514) );
  NAND2_X1 U10474 ( .A1(a_16_), .A2(b_30_), .ZN(n10688) );
  INV_X1 U10475 ( .A(n10689), .ZN(n10687) );
  XNOR2_X1 U10476 ( .A(n10690), .B(n10691), .ZN(n10512) );
  NAND2_X1 U10477 ( .A1(n10692), .A2(n10693), .ZN(n10690) );
  NAND2_X1 U10478 ( .A1(a_16_), .A2(n10689), .ZN(n10513) );
  NAND2_X1 U10479 ( .A1(n10509), .A2(n10694), .ZN(n10689) );
  NAND2_X1 U10480 ( .A1(n10508), .A2(n10510), .ZN(n10694) );
  NAND2_X1 U10481 ( .A1(n10695), .A2(n10696), .ZN(n10510) );
  NAND2_X1 U10482 ( .A1(a_17_), .A2(b_30_), .ZN(n10696) );
  INV_X1 U10483 ( .A(n10697), .ZN(n10695) );
  XNOR2_X1 U10484 ( .A(n10698), .B(n10699), .ZN(n10508) );
  NAND2_X1 U10485 ( .A1(n10700), .A2(n10701), .ZN(n10698) );
  NAND2_X1 U10486 ( .A1(a_17_), .A2(n10697), .ZN(n10509) );
  NAND2_X1 U10487 ( .A1(n10402), .A2(n10702), .ZN(n10697) );
  NAND2_X1 U10488 ( .A1(n10401), .A2(n10403), .ZN(n10702) );
  NAND2_X1 U10489 ( .A1(n10703), .A2(n10704), .ZN(n10403) );
  NAND2_X1 U10490 ( .A1(a_18_), .A2(b_30_), .ZN(n10704) );
  INV_X1 U10491 ( .A(n10705), .ZN(n10703) );
  XNOR2_X1 U10492 ( .A(n10706), .B(n10707), .ZN(n10401) );
  XOR2_X1 U10493 ( .A(n10708), .B(n10709), .Z(n10707) );
  NAND2_X1 U10494 ( .A1(b_29_), .A2(a_19_), .ZN(n10709) );
  NAND2_X1 U10495 ( .A1(a_18_), .A2(n10705), .ZN(n10402) );
  NAND2_X1 U10496 ( .A1(n10710), .A2(n10711), .ZN(n10705) );
  NAND2_X1 U10497 ( .A1(n10712), .A2(a_19_), .ZN(n10711) );
  NOR2_X1 U10498 ( .A1(n10713), .A2(n9080), .ZN(n10712) );
  NOR2_X1 U10499 ( .A1(n10409), .A2(n10408), .ZN(n10713) );
  NAND2_X1 U10500 ( .A1(n10409), .A2(n10408), .ZN(n10710) );
  XNOR2_X1 U10501 ( .A(n10714), .B(n10715), .ZN(n10408) );
  NAND2_X1 U10502 ( .A1(n10716), .A2(n10717), .ZN(n10714) );
  NOR2_X1 U10503 ( .A1(n10718), .A2(n10719), .ZN(n10409) );
  INV_X1 U10504 ( .A(n10720), .ZN(n10719) );
  NAND2_X1 U10505 ( .A1(n10503), .A2(n10721), .ZN(n10720) );
  NAND2_X1 U10506 ( .A1(n10506), .A2(n10505), .ZN(n10721) );
  XOR2_X1 U10507 ( .A(n10722), .B(n10723), .Z(n10503) );
  NAND2_X1 U10508 ( .A1(n10724), .A2(n10725), .ZN(n10722) );
  NOR2_X1 U10509 ( .A1(n10505), .A2(n10506), .ZN(n10718) );
  NOR2_X1 U10510 ( .A1(n10054), .A2(n9080), .ZN(n10506) );
  NAND2_X1 U10511 ( .A1(n10501), .A2(n10726), .ZN(n10505) );
  NAND2_X1 U10512 ( .A1(n10500), .A2(n10502), .ZN(n10726) );
  NAND2_X1 U10513 ( .A1(n10727), .A2(n10728), .ZN(n10502) );
  NAND2_X1 U10514 ( .A1(a_21_), .A2(b_30_), .ZN(n10727) );
  XNOR2_X1 U10515 ( .A(n10729), .B(n10730), .ZN(n10500) );
  NAND2_X1 U10516 ( .A1(n10731), .A2(n10732), .ZN(n10729) );
  INV_X1 U10517 ( .A(n10733), .ZN(n10501) );
  NOR2_X1 U10518 ( .A1(n10728), .A2(n9358), .ZN(n10733) );
  NAND2_X1 U10519 ( .A1(n10734), .A2(n10735), .ZN(n10728) );
  NAND2_X1 U10520 ( .A1(n10425), .A2(n10736), .ZN(n10735) );
  NAND2_X1 U10521 ( .A1(n10426), .A2(n10737), .ZN(n10736) );
  XNOR2_X1 U10522 ( .A(n10738), .B(n10739), .ZN(n10425) );
  XOR2_X1 U10523 ( .A(n10740), .B(n10741), .Z(n10738) );
  NOR2_X1 U10524 ( .A1(n10051), .A2(n10046), .ZN(n10741) );
  NAND2_X1 U10525 ( .A1(n10427), .A2(n10742), .ZN(n10734) );
  INV_X1 U10526 ( .A(n10426), .ZN(n10742) );
  NOR2_X1 U10527 ( .A1(n9330), .A2(n9080), .ZN(n10426) );
  INV_X1 U10528 ( .A(n10737), .ZN(n10427) );
  NAND2_X1 U10529 ( .A1(n10743), .A2(n10744), .ZN(n10737) );
  NAND2_X1 U10530 ( .A1(n10745), .A2(a_23_), .ZN(n10744) );
  NOR2_X1 U10531 ( .A1(n10746), .A2(n9080), .ZN(n10745) );
  NOR2_X1 U10532 ( .A1(n10435), .A2(n10434), .ZN(n10746) );
  NAND2_X1 U10533 ( .A1(n10434), .A2(n10435), .ZN(n10743) );
  NAND2_X1 U10534 ( .A1(n10747), .A2(n10748), .ZN(n10435) );
  NAND2_X1 U10535 ( .A1(n10498), .A2(n10749), .ZN(n10748) );
  INV_X1 U10536 ( .A(n10750), .ZN(n10749) );
  NOR2_X1 U10537 ( .A1(n10496), .A2(n10497), .ZN(n10750) );
  NOR2_X1 U10538 ( .A1(n10050), .A2(n9080), .ZN(n10498) );
  NAND2_X1 U10539 ( .A1(n10496), .A2(n10497), .ZN(n10747) );
  NAND2_X1 U10540 ( .A1(n10751), .A2(n10752), .ZN(n10497) );
  NAND2_X1 U10541 ( .A1(n10494), .A2(n10753), .ZN(n10752) );
  INV_X1 U10542 ( .A(n10754), .ZN(n10753) );
  NOR2_X1 U10543 ( .A1(n10491), .A2(n10493), .ZN(n10754) );
  NOR2_X1 U10544 ( .A1(n10048), .A2(n9080), .ZN(n10494) );
  NAND2_X1 U10545 ( .A1(n10491), .A2(n10493), .ZN(n10751) );
  NOR2_X1 U10546 ( .A1(n10755), .A2(n10756), .ZN(n10493) );
  INV_X1 U10547 ( .A(n10757), .ZN(n10756) );
  NAND2_X1 U10548 ( .A1(n10449), .A2(n10758), .ZN(n10757) );
  NAND2_X1 U10549 ( .A1(n10452), .A2(n10451), .ZN(n10758) );
  XOR2_X1 U10550 ( .A(n10759), .B(n10760), .Z(n10449) );
  NAND2_X1 U10551 ( .A1(n10761), .A2(n10762), .ZN(n10759) );
  NOR2_X1 U10552 ( .A1(n10451), .A2(n10452), .ZN(n10755) );
  NOR2_X1 U10553 ( .A1(n10047), .A2(n9080), .ZN(n10452) );
  NAND2_X1 U10554 ( .A1(n10459), .A2(n10763), .ZN(n10451) );
  NAND2_X1 U10555 ( .A1(n10458), .A2(n10460), .ZN(n10763) );
  NAND2_X1 U10556 ( .A1(n10764), .A2(n10765), .ZN(n10460) );
  NAND2_X1 U10557 ( .A1(b_30_), .A2(a_27_), .ZN(n10765) );
  INV_X1 U10558 ( .A(n10766), .ZN(n10764) );
  XNOR2_X1 U10559 ( .A(n10767), .B(n10768), .ZN(n10458) );
  XNOR2_X1 U10560 ( .A(n10769), .B(n10770), .ZN(n10767) );
  NOR2_X1 U10561 ( .A1(n9136), .A2(n10046), .ZN(n10770) );
  NAND2_X1 U10562 ( .A1(a_27_), .A2(n10766), .ZN(n10459) );
  NAND2_X1 U10563 ( .A1(n10771), .A2(n10772), .ZN(n10766) );
  NAND2_X1 U10564 ( .A1(n10773), .A2(b_30_), .ZN(n10772) );
  NOR2_X1 U10565 ( .A1(n10774), .A2(n9136), .ZN(n10773) );
  NOR2_X1 U10566 ( .A1(n10465), .A2(n10467), .ZN(n10774) );
  NAND2_X1 U10567 ( .A1(n10465), .A2(n10467), .ZN(n10771) );
  NAND2_X1 U10568 ( .A1(n10775), .A2(n10776), .ZN(n10467) );
  NAND2_X1 U10569 ( .A1(n10777), .A2(a_29_), .ZN(n10776) );
  NOR2_X1 U10570 ( .A1(n10778), .A2(n9080), .ZN(n10777) );
  NOR2_X1 U10571 ( .A1(n10779), .A2(n10475), .ZN(n10778) );
  NAND2_X1 U10572 ( .A1(n10779), .A2(n10475), .ZN(n10775) );
  NAND2_X1 U10573 ( .A1(n10780), .A2(n10781), .ZN(n10475) );
  NAND2_X1 U10574 ( .A1(b_28_), .A2(n10782), .ZN(n10781) );
  NAND2_X1 U10575 ( .A1(n10486), .A2(n10783), .ZN(n10782) );
  NAND2_X1 U10576 ( .A1(a_31_), .A2(n10046), .ZN(n10783) );
  NAND2_X1 U10577 ( .A1(b_29_), .A2(n10784), .ZN(n10780) );
  NAND2_X1 U10578 ( .A1(n10489), .A2(n10785), .ZN(n10784) );
  NAND2_X1 U10579 ( .A1(a_30_), .A2(n10786), .ZN(n10785) );
  INV_X1 U10580 ( .A(n10476), .ZN(n10779) );
  NAND2_X1 U10581 ( .A1(n10787), .A2(n9025), .ZN(n10476) );
  NOR2_X1 U10582 ( .A1(n9080), .A2(n10046), .ZN(n10787) );
  XNOR2_X1 U10583 ( .A(n10788), .B(n10037), .ZN(n10465) );
  INV_X1 U10584 ( .A(n10789), .ZN(n10037) );
  XNOR2_X1 U10585 ( .A(n10790), .B(n10791), .ZN(n10788) );
  XOR2_X1 U10586 ( .A(n10792), .B(n10793), .Z(n10491) );
  XNOR2_X1 U10587 ( .A(n10794), .B(n10795), .ZN(n10793) );
  XNOR2_X1 U10588 ( .A(n10796), .B(n10797), .ZN(n10496) );
  XNOR2_X1 U10589 ( .A(n10798), .B(n10799), .ZN(n10797) );
  XNOR2_X1 U10590 ( .A(n10800), .B(n10801), .ZN(n10434) );
  XNOR2_X1 U10591 ( .A(n10802), .B(n10803), .ZN(n10800) );
  XNOR2_X1 U10592 ( .A(n10804), .B(n10805), .ZN(n10516) );
  NAND2_X1 U10593 ( .A1(n10806), .A2(n10807), .ZN(n10804) );
  XNOR2_X1 U10594 ( .A(n10808), .B(n10809), .ZN(n10532) );
  NAND2_X1 U10595 ( .A1(n10810), .A2(n10811), .ZN(n10808) );
  XOR2_X1 U10596 ( .A(n10812), .B(n10813), .Z(n10540) );
  XNOR2_X1 U10597 ( .A(n10814), .B(n10815), .ZN(n10813) );
  XNOR2_X1 U10598 ( .A(n10816), .B(n10817), .ZN(n10556) );
  NAND2_X1 U10599 ( .A1(n10818), .A2(n10819), .ZN(n10816) );
  XNOR2_X1 U10600 ( .A(n10820), .B(n10821), .ZN(n10323) );
  XNOR2_X1 U10601 ( .A(n10822), .B(n10823), .ZN(n10820) );
  XNOR2_X1 U10602 ( .A(n10824), .B(n10825), .ZN(n10327) );
  NAND2_X1 U10603 ( .A1(n10826), .A2(n10827), .ZN(n10824) );
  INV_X1 U10604 ( .A(n10828), .ZN(n10120) );
  NOR2_X1 U10605 ( .A1(n10317), .A2(n10316), .ZN(n10828) );
  XNOR2_X1 U10606 ( .A(n10829), .B(n10830), .ZN(n10316) );
  NAND2_X1 U10607 ( .A1(n10577), .A2(n10576), .ZN(n10317) );
  NAND2_X1 U10608 ( .A1(n10826), .A2(n10831), .ZN(n10576) );
  NAND2_X1 U10609 ( .A1(n10825), .A2(n10827), .ZN(n10831) );
  NAND2_X1 U10610 ( .A1(n10832), .A2(n10833), .ZN(n10827) );
  NAND2_X1 U10611 ( .A1(b_29_), .A2(a_0_), .ZN(n10833) );
  XOR2_X1 U10612 ( .A(n10834), .B(n10835), .Z(n10825) );
  XOR2_X1 U10613 ( .A(n10836), .B(n10837), .Z(n10834) );
  NAND2_X1 U10614 ( .A1(a_0_), .A2(n10838), .ZN(n10826) );
  INV_X1 U10615 ( .A(n10832), .ZN(n10838) );
  NOR2_X1 U10616 ( .A1(n10839), .A2(n10840), .ZN(n10832) );
  INV_X1 U10617 ( .A(n10841), .ZN(n10840) );
  NAND2_X1 U10618 ( .A1(n10823), .A2(n10842), .ZN(n10841) );
  NAND2_X1 U10619 ( .A1(n10822), .A2(n10821), .ZN(n10842) );
  NOR2_X1 U10620 ( .A1(n10046), .A2(n9983), .ZN(n10823) );
  NOR2_X1 U10621 ( .A1(n10821), .A2(n10822), .ZN(n10839) );
  NOR2_X1 U10622 ( .A1(n10843), .A2(n10844), .ZN(n10822) );
  INV_X1 U10623 ( .A(n10845), .ZN(n10844) );
  NAND2_X1 U10624 ( .A1(n10588), .A2(n10846), .ZN(n10845) );
  NAND2_X1 U10625 ( .A1(n10587), .A2(n10589), .ZN(n10846) );
  NAND2_X1 U10626 ( .A1(n10596), .A2(n10847), .ZN(n10588) );
  NAND2_X1 U10627 ( .A1(n10595), .A2(n10597), .ZN(n10847) );
  NAND2_X1 U10628 ( .A1(n10848), .A2(n10849), .ZN(n10597) );
  NAND2_X1 U10629 ( .A1(b_29_), .A2(a_3_), .ZN(n10848) );
  XNOR2_X1 U10630 ( .A(n10850), .B(n10851), .ZN(n10595) );
  XOR2_X1 U10631 ( .A(n10852), .B(n10853), .Z(n10851) );
  NAND2_X1 U10632 ( .A1(a_4_), .A2(b_28_), .ZN(n10853) );
  NAND2_X1 U10633 ( .A1(n10854), .A2(a_3_), .ZN(n10596) );
  INV_X1 U10634 ( .A(n10849), .ZN(n10854) );
  NAND2_X1 U10635 ( .A1(n10855), .A2(n10856), .ZN(n10849) );
  NAND2_X1 U10636 ( .A1(n10602), .A2(n10857), .ZN(n10856) );
  NAND2_X1 U10637 ( .A1(n10605), .A2(n10604), .ZN(n10857) );
  XNOR2_X1 U10638 ( .A(n10858), .B(n10859), .ZN(n10602) );
  XNOR2_X1 U10639 ( .A(n10860), .B(n10861), .ZN(n10859) );
  NAND2_X1 U10640 ( .A1(a_5_), .A2(b_28_), .ZN(n10861) );
  INV_X1 U10641 ( .A(n10862), .ZN(n10855) );
  NOR2_X1 U10642 ( .A1(n10604), .A2(n10605), .ZN(n10862) );
  NOR2_X1 U10643 ( .A1(n10046), .A2(n10085), .ZN(n10605) );
  NAND2_X1 U10644 ( .A1(n10863), .A2(n10864), .ZN(n10604) );
  NAND2_X1 U10645 ( .A1(n10865), .A2(b_29_), .ZN(n10864) );
  NOR2_X1 U10646 ( .A1(n10866), .A2(n10083), .ZN(n10865) );
  NOR2_X1 U10647 ( .A1(n10611), .A2(n10612), .ZN(n10866) );
  NAND2_X1 U10648 ( .A1(n10611), .A2(n10612), .ZN(n10863) );
  NAND2_X1 U10649 ( .A1(n10818), .A2(n10867), .ZN(n10612) );
  NAND2_X1 U10650 ( .A1(n10817), .A2(n10819), .ZN(n10867) );
  NAND2_X1 U10651 ( .A1(n10868), .A2(n10869), .ZN(n10819) );
  NAND2_X1 U10652 ( .A1(b_29_), .A2(a_6_), .ZN(n10869) );
  INV_X1 U10653 ( .A(n10870), .ZN(n10868) );
  XNOR2_X1 U10654 ( .A(n10871), .B(n10872), .ZN(n10817) );
  NAND2_X1 U10655 ( .A1(n10873), .A2(n10874), .ZN(n10871) );
  NAND2_X1 U10656 ( .A1(a_6_), .A2(n10870), .ZN(n10818) );
  NAND2_X1 U10657 ( .A1(n10624), .A2(n10875), .ZN(n10870) );
  NAND2_X1 U10658 ( .A1(n10623), .A2(n10625), .ZN(n10875) );
  NAND2_X1 U10659 ( .A1(n10876), .A2(n10877), .ZN(n10625) );
  NAND2_X1 U10660 ( .A1(b_29_), .A2(a_7_), .ZN(n10877) );
  INV_X1 U10661 ( .A(n10878), .ZN(n10876) );
  XNOR2_X1 U10662 ( .A(n10879), .B(n10880), .ZN(n10623) );
  NAND2_X1 U10663 ( .A1(n10881), .A2(n10882), .ZN(n10879) );
  NAND2_X1 U10664 ( .A1(a_7_), .A2(n10878), .ZN(n10624) );
  NAND2_X1 U10665 ( .A1(n10632), .A2(n10883), .ZN(n10878) );
  NAND2_X1 U10666 ( .A1(n10631), .A2(n10633), .ZN(n10883) );
  NAND2_X1 U10667 ( .A1(n10884), .A2(n10885), .ZN(n10633) );
  NAND2_X1 U10668 ( .A1(b_29_), .A2(a_8_), .ZN(n10885) );
  INV_X1 U10669 ( .A(n10886), .ZN(n10884) );
  XNOR2_X1 U10670 ( .A(n10887), .B(n10888), .ZN(n10631) );
  XNOR2_X1 U10671 ( .A(n10889), .B(n10890), .ZN(n10887) );
  NOR2_X1 U10672 ( .A1(n10786), .A2(n10076), .ZN(n10890) );
  NAND2_X1 U10673 ( .A1(a_8_), .A2(n10886), .ZN(n10632) );
  NAND2_X1 U10674 ( .A1(n10891), .A2(n10892), .ZN(n10886) );
  NAND2_X1 U10675 ( .A1(n10893), .A2(b_29_), .ZN(n10892) );
  NOR2_X1 U10676 ( .A1(n10894), .A2(n10076), .ZN(n10893) );
  NOR2_X1 U10677 ( .A1(n10640), .A2(n10639), .ZN(n10894) );
  NAND2_X1 U10678 ( .A1(n10640), .A2(n10639), .ZN(n10891) );
  XOR2_X1 U10679 ( .A(n10895), .B(n10896), .Z(n10639) );
  XNOR2_X1 U10680 ( .A(n10897), .B(n10898), .ZN(n10896) );
  NOR2_X1 U10681 ( .A1(n10899), .A2(n10900), .ZN(n10640) );
  INV_X1 U10682 ( .A(n10901), .ZN(n10900) );
  NAND2_X1 U10683 ( .A1(n10812), .A2(n10902), .ZN(n10901) );
  NAND2_X1 U10684 ( .A1(n10815), .A2(n10814), .ZN(n10902) );
  XNOR2_X1 U10685 ( .A(n10903), .B(n10904), .ZN(n10812) );
  XOR2_X1 U10686 ( .A(n10905), .B(n10906), .Z(n10903) );
  NOR2_X1 U10687 ( .A1(n10786), .A2(n9649), .ZN(n10906) );
  NOR2_X1 U10688 ( .A1(n10814), .A2(n10815), .ZN(n10899) );
  NOR2_X1 U10689 ( .A1(n10046), .A2(n10073), .ZN(n10815) );
  NAND2_X1 U10690 ( .A1(n10907), .A2(n10908), .ZN(n10814) );
  NAND2_X1 U10691 ( .A1(n10909), .A2(b_29_), .ZN(n10908) );
  NOR2_X1 U10692 ( .A1(n10910), .A2(n9649), .ZN(n10909) );
  NOR2_X1 U10693 ( .A1(n10651), .A2(n10652), .ZN(n10910) );
  NAND2_X1 U10694 ( .A1(n10651), .A2(n10652), .ZN(n10907) );
  NAND2_X1 U10695 ( .A1(n10810), .A2(n10911), .ZN(n10652) );
  NAND2_X1 U10696 ( .A1(n10809), .A2(n10811), .ZN(n10911) );
  NAND2_X1 U10697 ( .A1(n10912), .A2(n10913), .ZN(n10811) );
  NAND2_X1 U10698 ( .A1(b_29_), .A2(a_12_), .ZN(n10913) );
  INV_X1 U10699 ( .A(n10914), .ZN(n10912) );
  XNOR2_X1 U10700 ( .A(n10915), .B(n10916), .ZN(n10809) );
  NAND2_X1 U10701 ( .A1(n10917), .A2(n10918), .ZN(n10915) );
  NAND2_X1 U10702 ( .A1(a_12_), .A2(n10914), .ZN(n10810) );
  NAND2_X1 U10703 ( .A1(n10664), .A2(n10919), .ZN(n10914) );
  NAND2_X1 U10704 ( .A1(n10663), .A2(n10665), .ZN(n10919) );
  NAND2_X1 U10705 ( .A1(n10920), .A2(n10921), .ZN(n10665) );
  NAND2_X1 U10706 ( .A1(b_29_), .A2(a_13_), .ZN(n10921) );
  INV_X1 U10707 ( .A(n10922), .ZN(n10920) );
  XNOR2_X1 U10708 ( .A(n10923), .B(n10924), .ZN(n10663) );
  NAND2_X1 U10709 ( .A1(n10925), .A2(n10926), .ZN(n10923) );
  NAND2_X1 U10710 ( .A1(a_13_), .A2(n10922), .ZN(n10664) );
  NAND2_X1 U10711 ( .A1(n10672), .A2(n10927), .ZN(n10922) );
  NAND2_X1 U10712 ( .A1(n10671), .A2(n10673), .ZN(n10927) );
  NAND2_X1 U10713 ( .A1(n10928), .A2(n10929), .ZN(n10673) );
  NAND2_X1 U10714 ( .A1(b_29_), .A2(a_14_), .ZN(n10929) );
  INV_X1 U10715 ( .A(n10930), .ZN(n10928) );
  XOR2_X1 U10716 ( .A(n10931), .B(n10932), .Z(n10671) );
  XOR2_X1 U10717 ( .A(n10933), .B(n10934), .Z(n10931) );
  NOR2_X1 U10718 ( .A1(n10786), .A2(n9534), .ZN(n10934) );
  NAND2_X1 U10719 ( .A1(a_14_), .A2(n10930), .ZN(n10672) );
  NAND2_X1 U10720 ( .A1(n10935), .A2(n10936), .ZN(n10930) );
  NAND2_X1 U10721 ( .A1(n10937), .A2(b_29_), .ZN(n10936) );
  NOR2_X1 U10722 ( .A1(n10938), .A2(n9534), .ZN(n10937) );
  NOR2_X1 U10723 ( .A1(n10679), .A2(n10680), .ZN(n10938) );
  NAND2_X1 U10724 ( .A1(n10679), .A2(n10680), .ZN(n10935) );
  NAND2_X1 U10725 ( .A1(n10806), .A2(n10939), .ZN(n10680) );
  NAND2_X1 U10726 ( .A1(n10805), .A2(n10807), .ZN(n10939) );
  NAND2_X1 U10727 ( .A1(n10940), .A2(n10941), .ZN(n10807) );
  NAND2_X1 U10728 ( .A1(b_29_), .A2(a_16_), .ZN(n10941) );
  INV_X1 U10729 ( .A(n10942), .ZN(n10940) );
  XNOR2_X1 U10730 ( .A(n10943), .B(n10944), .ZN(n10805) );
  NAND2_X1 U10731 ( .A1(n10945), .A2(n10946), .ZN(n10943) );
  NAND2_X1 U10732 ( .A1(a_16_), .A2(n10942), .ZN(n10806) );
  NAND2_X1 U10733 ( .A1(n10692), .A2(n10947), .ZN(n10942) );
  NAND2_X1 U10734 ( .A1(n10691), .A2(n10693), .ZN(n10947) );
  NAND2_X1 U10735 ( .A1(n10948), .A2(n10949), .ZN(n10693) );
  NAND2_X1 U10736 ( .A1(b_29_), .A2(a_17_), .ZN(n10949) );
  INV_X1 U10737 ( .A(n10950), .ZN(n10948) );
  XNOR2_X1 U10738 ( .A(n10951), .B(n10952), .ZN(n10691) );
  NAND2_X1 U10739 ( .A1(n10953), .A2(n10954), .ZN(n10951) );
  NAND2_X1 U10740 ( .A1(a_17_), .A2(n10950), .ZN(n10692) );
  NAND2_X1 U10741 ( .A1(n10700), .A2(n10955), .ZN(n10950) );
  NAND2_X1 U10742 ( .A1(n10699), .A2(n10701), .ZN(n10955) );
  NAND2_X1 U10743 ( .A1(n10956), .A2(n10957), .ZN(n10701) );
  NAND2_X1 U10744 ( .A1(b_29_), .A2(a_18_), .ZN(n10957) );
  INV_X1 U10745 ( .A(n10958), .ZN(n10956) );
  XNOR2_X1 U10746 ( .A(n10959), .B(n10960), .ZN(n10699) );
  XOR2_X1 U10747 ( .A(n10961), .B(n10962), .Z(n10960) );
  NAND2_X1 U10748 ( .A1(a_19_), .A2(b_28_), .ZN(n10962) );
  NAND2_X1 U10749 ( .A1(a_18_), .A2(n10958), .ZN(n10700) );
  NAND2_X1 U10750 ( .A1(n10963), .A2(n10964), .ZN(n10958) );
  NAND2_X1 U10751 ( .A1(n10965), .A2(b_29_), .ZN(n10964) );
  NOR2_X1 U10752 ( .A1(n10966), .A2(n9415), .ZN(n10965) );
  NOR2_X1 U10753 ( .A1(n10706), .A2(n10708), .ZN(n10966) );
  NAND2_X1 U10754 ( .A1(n10706), .A2(n10708), .ZN(n10963) );
  NAND2_X1 U10755 ( .A1(n10716), .A2(n10967), .ZN(n10708) );
  NAND2_X1 U10756 ( .A1(n10715), .A2(n10717), .ZN(n10967) );
  NAND2_X1 U10757 ( .A1(n10968), .A2(n10969), .ZN(n10717) );
  NAND2_X1 U10758 ( .A1(b_29_), .A2(a_20_), .ZN(n10969) );
  INV_X1 U10759 ( .A(n10970), .ZN(n10968) );
  XNOR2_X1 U10760 ( .A(n10971), .B(n10972), .ZN(n10715) );
  NAND2_X1 U10761 ( .A1(n10973), .A2(n10974), .ZN(n10971) );
  NAND2_X1 U10762 ( .A1(a_20_), .A2(n10970), .ZN(n10716) );
  NAND2_X1 U10763 ( .A1(n10724), .A2(n10975), .ZN(n10970) );
  NAND2_X1 U10764 ( .A1(n10723), .A2(n10725), .ZN(n10975) );
  NAND2_X1 U10765 ( .A1(n10976), .A2(n10977), .ZN(n10725) );
  NAND2_X1 U10766 ( .A1(b_29_), .A2(a_21_), .ZN(n10977) );
  INV_X1 U10767 ( .A(n10978), .ZN(n10976) );
  XNOR2_X1 U10768 ( .A(n10979), .B(n10980), .ZN(n10723) );
  NAND2_X1 U10769 ( .A1(n10981), .A2(n10982), .ZN(n10979) );
  NAND2_X1 U10770 ( .A1(a_21_), .A2(n10978), .ZN(n10724) );
  NAND2_X1 U10771 ( .A1(n10731), .A2(n10983), .ZN(n10978) );
  NAND2_X1 U10772 ( .A1(n10730), .A2(n10732), .ZN(n10983) );
  NAND2_X1 U10773 ( .A1(n10984), .A2(n10985), .ZN(n10732) );
  NAND2_X1 U10774 ( .A1(b_29_), .A2(a_22_), .ZN(n10985) );
  INV_X1 U10775 ( .A(n10986), .ZN(n10984) );
  XOR2_X1 U10776 ( .A(n10987), .B(n10988), .Z(n10730) );
  XOR2_X1 U10777 ( .A(n10989), .B(n10990), .Z(n10987) );
  NOR2_X1 U10778 ( .A1(n10786), .A2(n10051), .ZN(n10990) );
  NAND2_X1 U10779 ( .A1(a_22_), .A2(n10986), .ZN(n10731) );
  NAND2_X1 U10780 ( .A1(n10991), .A2(n10992), .ZN(n10986) );
  NAND2_X1 U10781 ( .A1(n10993), .A2(b_29_), .ZN(n10992) );
  NOR2_X1 U10782 ( .A1(n10994), .A2(n10051), .ZN(n10993) );
  NOR2_X1 U10783 ( .A1(n10739), .A2(n10740), .ZN(n10994) );
  NAND2_X1 U10784 ( .A1(n10739), .A2(n10740), .ZN(n10991) );
  NAND2_X1 U10785 ( .A1(n10995), .A2(n10996), .ZN(n10740) );
  NAND2_X1 U10786 ( .A1(n10803), .A2(n10997), .ZN(n10996) );
  NAND2_X1 U10787 ( .A1(n10802), .A2(n10801), .ZN(n10997) );
  NOR2_X1 U10788 ( .A1(n10046), .A2(n10050), .ZN(n10803) );
  INV_X1 U10789 ( .A(n10998), .ZN(n10995) );
  NOR2_X1 U10790 ( .A1(n10801), .A2(n10802), .ZN(n10998) );
  NOR2_X1 U10791 ( .A1(n10999), .A2(n11000), .ZN(n10802) );
  INV_X1 U10792 ( .A(n11001), .ZN(n11000) );
  NAND2_X1 U10793 ( .A1(n10799), .A2(n11002), .ZN(n11001) );
  NAND2_X1 U10794 ( .A1(n10796), .A2(n10798), .ZN(n11002) );
  NOR2_X1 U10795 ( .A1(n10046), .A2(n10048), .ZN(n10799) );
  NOR2_X1 U10796 ( .A1(n10798), .A2(n10796), .ZN(n10999) );
  XNOR2_X1 U10797 ( .A(n11003), .B(n11004), .ZN(n10796) );
  XNOR2_X1 U10798 ( .A(n11005), .B(n11006), .ZN(n11004) );
  NAND2_X1 U10799 ( .A1(n11007), .A2(n11008), .ZN(n10798) );
  NAND2_X1 U10800 ( .A1(n10792), .A2(n11009), .ZN(n11008) );
  NAND2_X1 U10801 ( .A1(n10795), .A2(n10794), .ZN(n11009) );
  XOR2_X1 U10802 ( .A(n11010), .B(n11011), .Z(n10792) );
  XNOR2_X1 U10803 ( .A(n11012), .B(n11013), .ZN(n11010) );
  INV_X1 U10804 ( .A(n11014), .ZN(n11007) );
  NOR2_X1 U10805 ( .A1(n10794), .A2(n10795), .ZN(n11014) );
  NOR2_X1 U10806 ( .A1(n10046), .A2(n10047), .ZN(n10795) );
  NAND2_X1 U10807 ( .A1(n10761), .A2(n11015), .ZN(n10794) );
  NAND2_X1 U10808 ( .A1(n10760), .A2(n10762), .ZN(n11015) );
  NAND2_X1 U10809 ( .A1(n11016), .A2(n11017), .ZN(n10762) );
  NAND2_X1 U10810 ( .A1(b_29_), .A2(a_27_), .ZN(n11017) );
  INV_X1 U10811 ( .A(n11018), .ZN(n11016) );
  XOR2_X1 U10812 ( .A(n11019), .B(n11020), .Z(n10760) );
  XNOR2_X1 U10813 ( .A(n11021), .B(n10034), .ZN(n11020) );
  NAND2_X1 U10814 ( .A1(a_27_), .A2(n11018), .ZN(n10761) );
  NAND2_X1 U10815 ( .A1(n11022), .A2(n11023), .ZN(n11018) );
  NAND2_X1 U10816 ( .A1(n11024), .A2(b_29_), .ZN(n11023) );
  NOR2_X1 U10817 ( .A1(n11025), .A2(n9136), .ZN(n11024) );
  NOR2_X1 U10818 ( .A1(n10769), .A2(n10768), .ZN(n11025) );
  NAND2_X1 U10819 ( .A1(n10769), .A2(n10768), .ZN(n11022) );
  XOR2_X1 U10820 ( .A(n11026), .B(n11027), .Z(n10768) );
  NOR2_X1 U10821 ( .A1(n9121), .A2(n10786), .ZN(n11027) );
  XNOR2_X1 U10822 ( .A(n11028), .B(n11029), .ZN(n11026) );
  NOR2_X1 U10823 ( .A1(n11030), .A2(n11031), .ZN(n10769) );
  INV_X1 U10824 ( .A(n11032), .ZN(n11031) );
  NAND2_X1 U10825 ( .A1(n11033), .A2(n10791), .ZN(n11032) );
  NAND2_X1 U10826 ( .A1(n11034), .A2(n9025), .ZN(n10791) );
  NOR2_X1 U10827 ( .A1(n10786), .A2(n10046), .ZN(n11034) );
  NAND2_X1 U10828 ( .A1(n10789), .A2(n10790), .ZN(n11033) );
  NOR2_X1 U10829 ( .A1(n10790), .A2(n10789), .ZN(n11030) );
  NOR2_X1 U10830 ( .A1(n10046), .A2(n9121), .ZN(n10789) );
  NAND2_X1 U10831 ( .A1(n11035), .A2(n11036), .ZN(n10790) );
  NAND2_X1 U10832 ( .A1(b_27_), .A2(n11037), .ZN(n11036) );
  NAND2_X1 U10833 ( .A1(n10486), .A2(n11038), .ZN(n11037) );
  NAND2_X1 U10834 ( .A1(a_31_), .A2(n10786), .ZN(n11038) );
  NAND2_X1 U10835 ( .A1(b_28_), .A2(n11039), .ZN(n11035) );
  NAND2_X1 U10836 ( .A1(n10489), .A2(n11040), .ZN(n11039) );
  NAND2_X1 U10837 ( .A1(a_30_), .A2(n11041), .ZN(n11040) );
  XNOR2_X1 U10838 ( .A(n11042), .B(n11043), .ZN(n10801) );
  XOR2_X1 U10839 ( .A(n11044), .B(n11045), .Z(n11043) );
  XNOR2_X1 U10840 ( .A(n11046), .B(n11047), .ZN(n10739) );
  XNOR2_X1 U10841 ( .A(n11048), .B(n11049), .ZN(n11047) );
  XNOR2_X1 U10842 ( .A(n11050), .B(n11051), .ZN(n10706) );
  NAND2_X1 U10843 ( .A1(n11052), .A2(n11053), .ZN(n11050) );
  XNOR2_X1 U10844 ( .A(n11054), .B(n11055), .ZN(n10679) );
  NAND2_X1 U10845 ( .A1(n11056), .A2(n11057), .ZN(n11054) );
  XNOR2_X1 U10846 ( .A(n11058), .B(n11059), .ZN(n10651) );
  NAND2_X1 U10847 ( .A1(n11060), .A2(n11061), .ZN(n11058) );
  XOR2_X1 U10848 ( .A(n11062), .B(n11063), .Z(n10611) );
  XNOR2_X1 U10849 ( .A(n11064), .B(n11065), .ZN(n11063) );
  NOR2_X1 U10850 ( .A1(n10589), .A2(n10587), .ZN(n10843) );
  XOR2_X1 U10851 ( .A(n11066), .B(n11067), .Z(n10587) );
  XOR2_X1 U10852 ( .A(n11068), .B(n11069), .Z(n11067) );
  NAND2_X1 U10853 ( .A1(a_3_), .A2(b_28_), .ZN(n11069) );
  NAND2_X1 U10854 ( .A1(b_29_), .A2(a_2_), .ZN(n10589) );
  XNOR2_X1 U10855 ( .A(n11070), .B(n11071), .ZN(n10821) );
  XOR2_X1 U10856 ( .A(n11072), .B(n11073), .Z(n11070) );
  XOR2_X1 U10857 ( .A(n11074), .B(n11075), .Z(n10577) );
  XOR2_X1 U10858 ( .A(n11076), .B(n11077), .Z(n11074) );
  INV_X1 U10859 ( .A(n11078), .ZN(n10125) );
  NOR2_X1 U10860 ( .A1(n10313), .A2(n10314), .ZN(n11078) );
  NAND2_X1 U10861 ( .A1(n11079), .A2(n10308), .ZN(n10314) );
  NAND2_X1 U10862 ( .A1(n11080), .A2(n11081), .ZN(n10308) );
  XOR2_X1 U10863 ( .A(n11082), .B(n11083), .Z(n11080) );
  NAND2_X1 U10864 ( .A1(n11084), .A2(n11085), .ZN(n11079) );
  INV_X1 U10865 ( .A(n11081), .ZN(n11085) );
  NAND2_X1 U10866 ( .A1(n11086), .A2(n11087), .ZN(n11081) );
  NAND2_X1 U10867 ( .A1(n11088), .A2(a_0_), .ZN(n11087) );
  NOR2_X1 U10868 ( .A1(n11089), .A2(n11041), .ZN(n11088) );
  NOR2_X1 U10869 ( .A1(n11090), .A2(n11091), .ZN(n11089) );
  NAND2_X1 U10870 ( .A1(n11090), .A2(n11091), .ZN(n11086) );
  XNOR2_X1 U10871 ( .A(n11083), .B(n11082), .ZN(n11084) );
  XOR2_X1 U10872 ( .A(n11092), .B(n11093), .Z(n11083) );
  NAND2_X1 U10873 ( .A1(n10830), .A2(n10829), .ZN(n10313) );
  NAND2_X1 U10874 ( .A1(n11094), .A2(n11095), .ZN(n10829) );
  NAND2_X1 U10875 ( .A1(n11076), .A2(n11096), .ZN(n11095) );
  INV_X1 U10876 ( .A(n11097), .ZN(n11096) );
  NOR2_X1 U10877 ( .A1(n11077), .A2(n11075), .ZN(n11097) );
  NOR2_X1 U10878 ( .A1(n10093), .A2(n10786), .ZN(n11076) );
  NAND2_X1 U10879 ( .A1(n11075), .A2(n11077), .ZN(n11094) );
  NAND2_X1 U10880 ( .A1(n11098), .A2(n11099), .ZN(n11077) );
  NAND2_X1 U10881 ( .A1(n10837), .A2(n11100), .ZN(n11099) );
  INV_X1 U10882 ( .A(n11101), .ZN(n11100) );
  NOR2_X1 U10883 ( .A1(n10836), .A2(n10835), .ZN(n11101) );
  NOR2_X1 U10884 ( .A1(n9983), .A2(n10786), .ZN(n10837) );
  NAND2_X1 U10885 ( .A1(n10835), .A2(n10836), .ZN(n11098) );
  NAND2_X1 U10886 ( .A1(n11102), .A2(n11103), .ZN(n10836) );
  NAND2_X1 U10887 ( .A1(n11073), .A2(n11104), .ZN(n11103) );
  INV_X1 U10888 ( .A(n11105), .ZN(n11104) );
  NOR2_X1 U10889 ( .A1(n11072), .A2(n11071), .ZN(n11105) );
  NOR2_X1 U10890 ( .A1(n10088), .A2(n10786), .ZN(n11073) );
  NAND2_X1 U10891 ( .A1(n11071), .A2(n11072), .ZN(n11102) );
  NAND2_X1 U10892 ( .A1(n11106), .A2(n11107), .ZN(n11072) );
  NAND2_X1 U10893 ( .A1(n11108), .A2(a_3_), .ZN(n11107) );
  NOR2_X1 U10894 ( .A1(n11109), .A2(n10786), .ZN(n11108) );
  NOR2_X1 U10895 ( .A1(n11066), .A2(n11068), .ZN(n11109) );
  NAND2_X1 U10896 ( .A1(n11066), .A2(n11068), .ZN(n11106) );
  NAND2_X1 U10897 ( .A1(n11110), .A2(n11111), .ZN(n11068) );
  NAND2_X1 U10898 ( .A1(n11112), .A2(a_4_), .ZN(n11111) );
  NOR2_X1 U10899 ( .A1(n11113), .A2(n10786), .ZN(n11112) );
  NOR2_X1 U10900 ( .A1(n10850), .A2(n10852), .ZN(n11113) );
  NAND2_X1 U10901 ( .A1(n10850), .A2(n10852), .ZN(n11110) );
  NAND2_X1 U10902 ( .A1(n11114), .A2(n11115), .ZN(n10852) );
  NAND2_X1 U10903 ( .A1(n11116), .A2(a_5_), .ZN(n11115) );
  NOR2_X1 U10904 ( .A1(n11117), .A2(n10786), .ZN(n11116) );
  NOR2_X1 U10905 ( .A1(n10860), .A2(n10858), .ZN(n11117) );
  NAND2_X1 U10906 ( .A1(n10860), .A2(n10858), .ZN(n11114) );
  XNOR2_X1 U10907 ( .A(n11118), .B(n11119), .ZN(n10858) );
  XNOR2_X1 U10908 ( .A(n11120), .B(n11121), .ZN(n11118) );
  NOR2_X1 U10909 ( .A1(n11122), .A2(n11123), .ZN(n10860) );
  INV_X1 U10910 ( .A(n11124), .ZN(n11123) );
  NAND2_X1 U10911 ( .A1(n11062), .A2(n11125), .ZN(n11124) );
  NAND2_X1 U10912 ( .A1(n11065), .A2(n11064), .ZN(n11125) );
  XOR2_X1 U10913 ( .A(n11126), .B(n11127), .Z(n11062) );
  NAND2_X1 U10914 ( .A1(n11128), .A2(n11129), .ZN(n11126) );
  NOR2_X1 U10915 ( .A1(n11064), .A2(n11065), .ZN(n11122) );
  NOR2_X1 U10916 ( .A1(n10081), .A2(n10786), .ZN(n11065) );
  NAND2_X1 U10917 ( .A1(n10873), .A2(n11130), .ZN(n11064) );
  NAND2_X1 U10918 ( .A1(n10872), .A2(n10874), .ZN(n11130) );
  NAND2_X1 U10919 ( .A1(n11131), .A2(n11132), .ZN(n10874) );
  NAND2_X1 U10920 ( .A1(a_7_), .A2(b_28_), .ZN(n11132) );
  INV_X1 U10921 ( .A(n11133), .ZN(n11131) );
  XNOR2_X1 U10922 ( .A(n11134), .B(n11135), .ZN(n10872) );
  NAND2_X1 U10923 ( .A1(n11136), .A2(n11137), .ZN(n11134) );
  NAND2_X1 U10924 ( .A1(a_7_), .A2(n11133), .ZN(n10873) );
  NAND2_X1 U10925 ( .A1(n10881), .A2(n11138), .ZN(n11133) );
  NAND2_X1 U10926 ( .A1(n10880), .A2(n10882), .ZN(n11138) );
  NAND2_X1 U10927 ( .A1(n11139), .A2(n11140), .ZN(n10882) );
  NAND2_X1 U10928 ( .A1(a_8_), .A2(b_28_), .ZN(n11140) );
  INV_X1 U10929 ( .A(n11141), .ZN(n11139) );
  XNOR2_X1 U10930 ( .A(n11142), .B(n11143), .ZN(n10880) );
  XNOR2_X1 U10931 ( .A(n11144), .B(n11145), .ZN(n11142) );
  NOR2_X1 U10932 ( .A1(n11041), .A2(n10076), .ZN(n11145) );
  NAND2_X1 U10933 ( .A1(a_8_), .A2(n11141), .ZN(n10881) );
  NAND2_X1 U10934 ( .A1(n11146), .A2(n11147), .ZN(n11141) );
  NAND2_X1 U10935 ( .A1(n11148), .A2(a_9_), .ZN(n11147) );
  NOR2_X1 U10936 ( .A1(n11149), .A2(n10786), .ZN(n11148) );
  NOR2_X1 U10937 ( .A1(n10889), .A2(n10888), .ZN(n11149) );
  NAND2_X1 U10938 ( .A1(n10889), .A2(n10888), .ZN(n11146) );
  XOR2_X1 U10939 ( .A(n11150), .B(n11151), .Z(n10888) );
  XNOR2_X1 U10940 ( .A(n11152), .B(n11153), .ZN(n11151) );
  NOR2_X1 U10941 ( .A1(n11154), .A2(n11155), .ZN(n10889) );
  INV_X1 U10942 ( .A(n11156), .ZN(n11155) );
  NAND2_X1 U10943 ( .A1(n10895), .A2(n11157), .ZN(n11156) );
  NAND2_X1 U10944 ( .A1(n10898), .A2(n10897), .ZN(n11157) );
  XNOR2_X1 U10945 ( .A(n11158), .B(n11159), .ZN(n10895) );
  XOR2_X1 U10946 ( .A(n11160), .B(n11161), .Z(n11158) );
  NOR2_X1 U10947 ( .A1(n11041), .A2(n9649), .ZN(n11161) );
  NOR2_X1 U10948 ( .A1(n10897), .A2(n10898), .ZN(n11154) );
  NOR2_X1 U10949 ( .A1(n10073), .A2(n10786), .ZN(n10898) );
  NAND2_X1 U10950 ( .A1(n11162), .A2(n11163), .ZN(n10897) );
  NAND2_X1 U10951 ( .A1(n11164), .A2(a_11_), .ZN(n11163) );
  NOR2_X1 U10952 ( .A1(n11165), .A2(n10786), .ZN(n11164) );
  NOR2_X1 U10953 ( .A1(n10904), .A2(n10905), .ZN(n11165) );
  NAND2_X1 U10954 ( .A1(n10904), .A2(n10905), .ZN(n11162) );
  NAND2_X1 U10955 ( .A1(n11060), .A2(n11166), .ZN(n10905) );
  NAND2_X1 U10956 ( .A1(n11059), .A2(n11061), .ZN(n11166) );
  NAND2_X1 U10957 ( .A1(n11167), .A2(n11168), .ZN(n11061) );
  NAND2_X1 U10958 ( .A1(a_12_), .A2(b_28_), .ZN(n11168) );
  INV_X1 U10959 ( .A(n11169), .ZN(n11167) );
  XNOR2_X1 U10960 ( .A(n11170), .B(n11171), .ZN(n11059) );
  NAND2_X1 U10961 ( .A1(n11172), .A2(n11173), .ZN(n11170) );
  NAND2_X1 U10962 ( .A1(a_12_), .A2(n11169), .ZN(n11060) );
  NAND2_X1 U10963 ( .A1(n10917), .A2(n11174), .ZN(n11169) );
  NAND2_X1 U10964 ( .A1(n10916), .A2(n10918), .ZN(n11174) );
  NAND2_X1 U10965 ( .A1(n11175), .A2(n11176), .ZN(n10918) );
  NAND2_X1 U10966 ( .A1(a_13_), .A2(b_28_), .ZN(n11176) );
  INV_X1 U10967 ( .A(n11177), .ZN(n11175) );
  XNOR2_X1 U10968 ( .A(n11178), .B(n11179), .ZN(n10916) );
  NAND2_X1 U10969 ( .A1(n11180), .A2(n11181), .ZN(n11178) );
  NAND2_X1 U10970 ( .A1(a_13_), .A2(n11177), .ZN(n10917) );
  NAND2_X1 U10971 ( .A1(n10925), .A2(n11182), .ZN(n11177) );
  NAND2_X1 U10972 ( .A1(n10924), .A2(n10926), .ZN(n11182) );
  NAND2_X1 U10973 ( .A1(n11183), .A2(n11184), .ZN(n10926) );
  NAND2_X1 U10974 ( .A1(a_14_), .A2(b_28_), .ZN(n11184) );
  INV_X1 U10975 ( .A(n11185), .ZN(n11183) );
  XOR2_X1 U10976 ( .A(n11186), .B(n11187), .Z(n10924) );
  XOR2_X1 U10977 ( .A(n11188), .B(n11189), .Z(n11186) );
  NOR2_X1 U10978 ( .A1(n11041), .A2(n9534), .ZN(n11189) );
  NAND2_X1 U10979 ( .A1(a_14_), .A2(n11185), .ZN(n10925) );
  NAND2_X1 U10980 ( .A1(n11190), .A2(n11191), .ZN(n11185) );
  NAND2_X1 U10981 ( .A1(n11192), .A2(a_15_), .ZN(n11191) );
  NOR2_X1 U10982 ( .A1(n11193), .A2(n10786), .ZN(n11192) );
  NOR2_X1 U10983 ( .A1(n10932), .A2(n10933), .ZN(n11193) );
  NAND2_X1 U10984 ( .A1(n10932), .A2(n10933), .ZN(n11190) );
  NAND2_X1 U10985 ( .A1(n11056), .A2(n11194), .ZN(n10933) );
  NAND2_X1 U10986 ( .A1(n11055), .A2(n11057), .ZN(n11194) );
  NAND2_X1 U10987 ( .A1(n11195), .A2(n11196), .ZN(n11057) );
  NAND2_X1 U10988 ( .A1(a_16_), .A2(b_28_), .ZN(n11196) );
  INV_X1 U10989 ( .A(n11197), .ZN(n11195) );
  XNOR2_X1 U10990 ( .A(n11198), .B(n11199), .ZN(n11055) );
  NAND2_X1 U10991 ( .A1(n11200), .A2(n11201), .ZN(n11198) );
  NAND2_X1 U10992 ( .A1(a_16_), .A2(n11197), .ZN(n11056) );
  NAND2_X1 U10993 ( .A1(n10945), .A2(n11202), .ZN(n11197) );
  NAND2_X1 U10994 ( .A1(n10944), .A2(n10946), .ZN(n11202) );
  NAND2_X1 U10995 ( .A1(n11203), .A2(n11204), .ZN(n10946) );
  NAND2_X1 U10996 ( .A1(a_17_), .A2(b_28_), .ZN(n11204) );
  INV_X1 U10997 ( .A(n11205), .ZN(n11203) );
  XNOR2_X1 U10998 ( .A(n11206), .B(n11207), .ZN(n10944) );
  NAND2_X1 U10999 ( .A1(n11208), .A2(n11209), .ZN(n11206) );
  NAND2_X1 U11000 ( .A1(a_17_), .A2(n11205), .ZN(n10945) );
  NAND2_X1 U11001 ( .A1(n10953), .A2(n11210), .ZN(n11205) );
  NAND2_X1 U11002 ( .A1(n10952), .A2(n10954), .ZN(n11210) );
  NAND2_X1 U11003 ( .A1(n11211), .A2(n11212), .ZN(n10954) );
  NAND2_X1 U11004 ( .A1(a_18_), .A2(b_28_), .ZN(n11212) );
  INV_X1 U11005 ( .A(n11213), .ZN(n11211) );
  XOR2_X1 U11006 ( .A(n11214), .B(n11215), .Z(n10952) );
  XOR2_X1 U11007 ( .A(n11216), .B(n11217), .Z(n11214) );
  NOR2_X1 U11008 ( .A1(n11041), .A2(n9415), .ZN(n11217) );
  NAND2_X1 U11009 ( .A1(a_18_), .A2(n11213), .ZN(n10953) );
  NAND2_X1 U11010 ( .A1(n11218), .A2(n11219), .ZN(n11213) );
  NAND2_X1 U11011 ( .A1(n11220), .A2(a_19_), .ZN(n11219) );
  NOR2_X1 U11012 ( .A1(n11221), .A2(n10786), .ZN(n11220) );
  NOR2_X1 U11013 ( .A1(n10959), .A2(n10961), .ZN(n11221) );
  NAND2_X1 U11014 ( .A1(n10959), .A2(n10961), .ZN(n11218) );
  NAND2_X1 U11015 ( .A1(n11052), .A2(n11222), .ZN(n10961) );
  NAND2_X1 U11016 ( .A1(n11051), .A2(n11053), .ZN(n11222) );
  NAND2_X1 U11017 ( .A1(n11223), .A2(n11224), .ZN(n11053) );
  NAND2_X1 U11018 ( .A1(a_20_), .A2(b_28_), .ZN(n11224) );
  INV_X1 U11019 ( .A(n11225), .ZN(n11223) );
  XNOR2_X1 U11020 ( .A(n11226), .B(n11227), .ZN(n11051) );
  NAND2_X1 U11021 ( .A1(n11228), .A2(n11229), .ZN(n11226) );
  NAND2_X1 U11022 ( .A1(a_20_), .A2(n11225), .ZN(n11052) );
  NAND2_X1 U11023 ( .A1(n10973), .A2(n11230), .ZN(n11225) );
  NAND2_X1 U11024 ( .A1(n10972), .A2(n10974), .ZN(n11230) );
  NAND2_X1 U11025 ( .A1(n11231), .A2(n11232), .ZN(n10974) );
  NAND2_X1 U11026 ( .A1(a_21_), .A2(b_28_), .ZN(n11232) );
  INV_X1 U11027 ( .A(n11233), .ZN(n11231) );
  XNOR2_X1 U11028 ( .A(n11234), .B(n11235), .ZN(n10972) );
  NAND2_X1 U11029 ( .A1(n11236), .A2(n11237), .ZN(n11234) );
  NAND2_X1 U11030 ( .A1(a_21_), .A2(n11233), .ZN(n10973) );
  NAND2_X1 U11031 ( .A1(n10981), .A2(n11238), .ZN(n11233) );
  NAND2_X1 U11032 ( .A1(n10980), .A2(n10982), .ZN(n11238) );
  NAND2_X1 U11033 ( .A1(n11239), .A2(n11240), .ZN(n10982) );
  NAND2_X1 U11034 ( .A1(a_22_), .A2(b_28_), .ZN(n11240) );
  INV_X1 U11035 ( .A(n11241), .ZN(n11239) );
  XOR2_X1 U11036 ( .A(n11242), .B(n11243), .Z(n10980) );
  XOR2_X1 U11037 ( .A(n11244), .B(n11245), .Z(n11242) );
  NOR2_X1 U11038 ( .A1(n11041), .A2(n10051), .ZN(n11245) );
  NAND2_X1 U11039 ( .A1(a_22_), .A2(n11241), .ZN(n10981) );
  NAND2_X1 U11040 ( .A1(n11246), .A2(n11247), .ZN(n11241) );
  NAND2_X1 U11041 ( .A1(n11248), .A2(a_23_), .ZN(n11247) );
  NOR2_X1 U11042 ( .A1(n11249), .A2(n10786), .ZN(n11248) );
  NOR2_X1 U11043 ( .A1(n10988), .A2(n10989), .ZN(n11249) );
  NAND2_X1 U11044 ( .A1(n10988), .A2(n10989), .ZN(n11246) );
  NAND2_X1 U11045 ( .A1(n11250), .A2(n11251), .ZN(n10989) );
  INV_X1 U11046 ( .A(n11252), .ZN(n11251) );
  NOR2_X1 U11047 ( .A1(n11253), .A2(n11254), .ZN(n11252) );
  NOR2_X1 U11048 ( .A1(n11048), .A2(n11046), .ZN(n11254) );
  INV_X1 U11049 ( .A(n11049), .ZN(n11253) );
  NOR2_X1 U11050 ( .A1(n10050), .A2(n10786), .ZN(n11049) );
  NAND2_X1 U11051 ( .A1(n11046), .A2(n11048), .ZN(n11250) );
  NAND2_X1 U11052 ( .A1(n11255), .A2(n11256), .ZN(n11048) );
  NAND2_X1 U11053 ( .A1(n11045), .A2(n11257), .ZN(n11256) );
  INV_X1 U11054 ( .A(n11258), .ZN(n11257) );
  NOR2_X1 U11055 ( .A1(n11042), .A2(n11044), .ZN(n11258) );
  NOR2_X1 U11056 ( .A1(n10048), .A2(n10786), .ZN(n11045) );
  NAND2_X1 U11057 ( .A1(n11044), .A2(n11042), .ZN(n11255) );
  XOR2_X1 U11058 ( .A(n11259), .B(n11260), .Z(n11042) );
  XOR2_X1 U11059 ( .A(n11261), .B(n11262), .Z(n11259) );
  NOR2_X1 U11060 ( .A1(n11263), .A2(n11264), .ZN(n11044) );
  INV_X1 U11061 ( .A(n11265), .ZN(n11264) );
  NAND2_X1 U11062 ( .A1(n11003), .A2(n11266), .ZN(n11265) );
  NAND2_X1 U11063 ( .A1(n11006), .A2(n11005), .ZN(n11266) );
  XNOR2_X1 U11064 ( .A(n11267), .B(n11268), .ZN(n11003) );
  XNOR2_X1 U11065 ( .A(n10031), .B(n11269), .ZN(n11268) );
  NOR2_X1 U11066 ( .A1(n11005), .A2(n11006), .ZN(n11263) );
  NOR2_X1 U11067 ( .A1(n10047), .A2(n10786), .ZN(n11006) );
  NAND2_X1 U11068 ( .A1(n11270), .A2(n11271), .ZN(n11005) );
  NAND2_X1 U11069 ( .A1(n11013), .A2(n11272), .ZN(n11271) );
  INV_X1 U11070 ( .A(n11273), .ZN(n11272) );
  NOR2_X1 U11071 ( .A1(n11011), .A2(n11012), .ZN(n11273) );
  NOR2_X1 U11072 ( .A1(n10786), .A2(n11274), .ZN(n11013) );
  NAND2_X1 U11073 ( .A1(n11012), .A2(n11011), .ZN(n11270) );
  XNOR2_X1 U11074 ( .A(n11275), .B(n11276), .ZN(n11011) );
  XOR2_X1 U11075 ( .A(n11277), .B(n11278), .Z(n11276) );
  NAND2_X1 U11076 ( .A1(b_27_), .A2(a_28_), .ZN(n11278) );
  NOR2_X1 U11077 ( .A1(n11279), .A2(n11280), .ZN(n11012) );
  INV_X1 U11078 ( .A(n11281), .ZN(n11280) );
  NAND2_X1 U11079 ( .A1(n11019), .A2(n11282), .ZN(n11281) );
  NAND2_X1 U11080 ( .A1(n10034), .A2(n11021), .ZN(n11282) );
  XNOR2_X1 U11081 ( .A(n11283), .B(n11284), .ZN(n11019) );
  NOR2_X1 U11082 ( .A1(n9121), .A2(n11041), .ZN(n11284) );
  XNOR2_X1 U11083 ( .A(n11285), .B(n11286), .ZN(n11283) );
  NOR2_X1 U11084 ( .A1(n11021), .A2(n10034), .ZN(n11279) );
  NOR2_X1 U11085 ( .A1(n10786), .A2(n9136), .ZN(n10034) );
  NAND2_X1 U11086 ( .A1(n11287), .A2(n11288), .ZN(n11021) );
  NAND2_X1 U11087 ( .A1(n11289), .A2(b_28_), .ZN(n11288) );
  NOR2_X1 U11088 ( .A1(n11290), .A2(n9121), .ZN(n11289) );
  NOR2_X1 U11089 ( .A1(n11291), .A2(n11028), .ZN(n11290) );
  NAND2_X1 U11090 ( .A1(n11291), .A2(n11028), .ZN(n11287) );
  NAND2_X1 U11091 ( .A1(n11292), .A2(n11293), .ZN(n11028) );
  NAND2_X1 U11092 ( .A1(b_26_), .A2(n11294), .ZN(n11293) );
  NAND2_X1 U11093 ( .A1(n10486), .A2(n11295), .ZN(n11294) );
  NAND2_X1 U11094 ( .A1(a_31_), .A2(n11041), .ZN(n11295) );
  NAND2_X1 U11095 ( .A1(b_27_), .A2(n11296), .ZN(n11292) );
  NAND2_X1 U11096 ( .A1(n10489), .A2(n11297), .ZN(n11296) );
  NAND2_X1 U11097 ( .A1(a_30_), .A2(n9217), .ZN(n11297) );
  INV_X1 U11098 ( .A(n11029), .ZN(n11291) );
  NAND2_X1 U11099 ( .A1(n11298), .A2(n9025), .ZN(n11029) );
  NOR2_X1 U11100 ( .A1(n10786), .A2(n11041), .ZN(n11298) );
  XNOR2_X1 U11101 ( .A(n11299), .B(n11300), .ZN(n11046) );
  XNOR2_X1 U11102 ( .A(n11301), .B(n11302), .ZN(n11300) );
  XNOR2_X1 U11103 ( .A(n11303), .B(n11304), .ZN(n10988) );
  XNOR2_X1 U11104 ( .A(n11305), .B(n11306), .ZN(n11304) );
  XNOR2_X1 U11105 ( .A(n11307), .B(n11308), .ZN(n10959) );
  NAND2_X1 U11106 ( .A1(n11309), .A2(n11310), .ZN(n11307) );
  XNOR2_X1 U11107 ( .A(n11311), .B(n11312), .ZN(n10932) );
  NAND2_X1 U11108 ( .A1(n11313), .A2(n11314), .ZN(n11311) );
  XNOR2_X1 U11109 ( .A(n11315), .B(n11316), .ZN(n10904) );
  NAND2_X1 U11110 ( .A1(n11317), .A2(n11318), .ZN(n11315) );
  XNOR2_X1 U11111 ( .A(n11319), .B(n11320), .ZN(n10850) );
  XNOR2_X1 U11112 ( .A(n11321), .B(n11322), .ZN(n11319) );
  XNOR2_X1 U11113 ( .A(n11323), .B(n11324), .ZN(n11066) );
  XNOR2_X1 U11114 ( .A(n11325), .B(n11326), .ZN(n11323) );
  XOR2_X1 U11115 ( .A(n11327), .B(n11328), .Z(n11071) );
  XOR2_X1 U11116 ( .A(n11329), .B(n11330), .Z(n11327) );
  NOR2_X1 U11117 ( .A1(n11041), .A2(n10086), .ZN(n11330) );
  XNOR2_X1 U11118 ( .A(n11331), .B(n11332), .ZN(n10835) );
  NAND2_X1 U11119 ( .A1(n11333), .A2(n11334), .ZN(n11331) );
  XOR2_X1 U11120 ( .A(n11335), .B(n11336), .Z(n11075) );
  XOR2_X1 U11121 ( .A(n11337), .B(n11338), .Z(n11335) );
  NOR2_X1 U11122 ( .A1(n11041), .A2(n9983), .ZN(n11338) );
  XNOR2_X1 U11123 ( .A(n11090), .B(n11339), .ZN(n10830) );
  XOR2_X1 U11124 ( .A(n11091), .B(n11340), .Z(n11339) );
  NAND2_X1 U11125 ( .A1(a_0_), .A2(b_27_), .ZN(n11340) );
  NAND2_X1 U11126 ( .A1(n11341), .A2(n11342), .ZN(n11091) );
  NAND2_X1 U11127 ( .A1(n11343), .A2(a_1_), .ZN(n11342) );
  NOR2_X1 U11128 ( .A1(n11344), .A2(n11041), .ZN(n11343) );
  NOR2_X1 U11129 ( .A1(n11336), .A2(n11337), .ZN(n11344) );
  NAND2_X1 U11130 ( .A1(n11336), .A2(n11337), .ZN(n11341) );
  NAND2_X1 U11131 ( .A1(n11333), .A2(n11345), .ZN(n11337) );
  NAND2_X1 U11132 ( .A1(n11332), .A2(n11334), .ZN(n11345) );
  NAND2_X1 U11133 ( .A1(n11346), .A2(n11347), .ZN(n11334) );
  NAND2_X1 U11134 ( .A1(a_2_), .A2(b_27_), .ZN(n11347) );
  INV_X1 U11135 ( .A(n11348), .ZN(n11346) );
  XNOR2_X1 U11136 ( .A(n11349), .B(n11350), .ZN(n11332) );
  XOR2_X1 U11137 ( .A(n11351), .B(n11352), .Z(n11350) );
  NAND2_X1 U11138 ( .A1(a_2_), .A2(n11348), .ZN(n11333) );
  NAND2_X1 U11139 ( .A1(n11353), .A2(n11354), .ZN(n11348) );
  NAND2_X1 U11140 ( .A1(n11355), .A2(a_3_), .ZN(n11354) );
  NOR2_X1 U11141 ( .A1(n11356), .A2(n11041), .ZN(n11355) );
  NOR2_X1 U11142 ( .A1(n11328), .A2(n11329), .ZN(n11356) );
  NAND2_X1 U11143 ( .A1(n11328), .A2(n11329), .ZN(n11353) );
  NAND2_X1 U11144 ( .A1(n11357), .A2(n11358), .ZN(n11329) );
  NAND2_X1 U11145 ( .A1(n11325), .A2(n11359), .ZN(n11358) );
  NAND2_X1 U11146 ( .A1(n11326), .A2(n11324), .ZN(n11359) );
  NOR2_X1 U11147 ( .A1(n10085), .A2(n11041), .ZN(n11325) );
  INV_X1 U11148 ( .A(n11360), .ZN(n11357) );
  NOR2_X1 U11149 ( .A1(n11324), .A2(n11326), .ZN(n11360) );
  NOR2_X1 U11150 ( .A1(n11361), .A2(n11362), .ZN(n11326) );
  INV_X1 U11151 ( .A(n11363), .ZN(n11362) );
  NAND2_X1 U11152 ( .A1(n11322), .A2(n11364), .ZN(n11363) );
  NAND2_X1 U11153 ( .A1(n11321), .A2(n11320), .ZN(n11364) );
  NOR2_X1 U11154 ( .A1(n10083), .A2(n11041), .ZN(n11322) );
  NOR2_X1 U11155 ( .A1(n11320), .A2(n11321), .ZN(n11361) );
  NOR2_X1 U11156 ( .A1(n11365), .A2(n11366), .ZN(n11321) );
  INV_X1 U11157 ( .A(n11367), .ZN(n11366) );
  NAND2_X1 U11158 ( .A1(n11120), .A2(n11368), .ZN(n11367) );
  NAND2_X1 U11159 ( .A1(n11119), .A2(n11121), .ZN(n11368) );
  NAND2_X1 U11160 ( .A1(n11128), .A2(n11369), .ZN(n11120) );
  NAND2_X1 U11161 ( .A1(n11127), .A2(n11129), .ZN(n11369) );
  NAND2_X1 U11162 ( .A1(n11370), .A2(n11371), .ZN(n11129) );
  NAND2_X1 U11163 ( .A1(a_7_), .A2(b_27_), .ZN(n11371) );
  INV_X1 U11164 ( .A(n11372), .ZN(n11370) );
  XNOR2_X1 U11165 ( .A(n11373), .B(n11374), .ZN(n11127) );
  XOR2_X1 U11166 ( .A(n11375), .B(n11376), .Z(n11374) );
  NAND2_X1 U11167 ( .A1(a_8_), .A2(b_26_), .ZN(n11376) );
  NAND2_X1 U11168 ( .A1(a_7_), .A2(n11372), .ZN(n11128) );
  NAND2_X1 U11169 ( .A1(n11136), .A2(n11377), .ZN(n11372) );
  NAND2_X1 U11170 ( .A1(n11135), .A2(n11137), .ZN(n11377) );
  NAND2_X1 U11171 ( .A1(n11378), .A2(n11379), .ZN(n11137) );
  NAND2_X1 U11172 ( .A1(a_8_), .A2(b_27_), .ZN(n11379) );
  INV_X1 U11173 ( .A(n11380), .ZN(n11378) );
  XNOR2_X1 U11174 ( .A(n11381), .B(n11382), .ZN(n11135) );
  XNOR2_X1 U11175 ( .A(n11383), .B(n11384), .ZN(n11381) );
  NOR2_X1 U11176 ( .A1(n9217), .A2(n10076), .ZN(n11384) );
  NAND2_X1 U11177 ( .A1(a_8_), .A2(n11380), .ZN(n11136) );
  NAND2_X1 U11178 ( .A1(n11385), .A2(n11386), .ZN(n11380) );
  NAND2_X1 U11179 ( .A1(n11387), .A2(a_9_), .ZN(n11386) );
  NOR2_X1 U11180 ( .A1(n11388), .A2(n11041), .ZN(n11387) );
  NOR2_X1 U11181 ( .A1(n11144), .A2(n11143), .ZN(n11388) );
  NAND2_X1 U11182 ( .A1(n11144), .A2(n11143), .ZN(n11385) );
  XOR2_X1 U11183 ( .A(n11389), .B(n11390), .Z(n11143) );
  XNOR2_X1 U11184 ( .A(n11391), .B(n11392), .ZN(n11390) );
  NOR2_X1 U11185 ( .A1(n11393), .A2(n11394), .ZN(n11144) );
  INV_X1 U11186 ( .A(n11395), .ZN(n11394) );
  NAND2_X1 U11187 ( .A1(n11150), .A2(n11396), .ZN(n11395) );
  NAND2_X1 U11188 ( .A1(n11153), .A2(n11152), .ZN(n11396) );
  XOR2_X1 U11189 ( .A(n11397), .B(n11398), .Z(n11150) );
  XOR2_X1 U11190 ( .A(n11399), .B(n11400), .Z(n11398) );
  NAND2_X1 U11191 ( .A1(a_11_), .A2(b_26_), .ZN(n11400) );
  NOR2_X1 U11192 ( .A1(n11152), .A2(n11153), .ZN(n11393) );
  NOR2_X1 U11193 ( .A1(n10073), .A2(n11041), .ZN(n11153) );
  NAND2_X1 U11194 ( .A1(n11401), .A2(n11402), .ZN(n11152) );
  NAND2_X1 U11195 ( .A1(n11403), .A2(a_11_), .ZN(n11402) );
  NOR2_X1 U11196 ( .A1(n11404), .A2(n11041), .ZN(n11403) );
  NOR2_X1 U11197 ( .A1(n11159), .A2(n11160), .ZN(n11404) );
  NAND2_X1 U11198 ( .A1(n11159), .A2(n11160), .ZN(n11401) );
  NAND2_X1 U11199 ( .A1(n11317), .A2(n11405), .ZN(n11160) );
  NAND2_X1 U11200 ( .A1(n11316), .A2(n11318), .ZN(n11405) );
  NAND2_X1 U11201 ( .A1(n11406), .A2(n11407), .ZN(n11318) );
  NAND2_X1 U11202 ( .A1(a_12_), .A2(b_27_), .ZN(n11407) );
  INV_X1 U11203 ( .A(n11408), .ZN(n11406) );
  XNOR2_X1 U11204 ( .A(n11409), .B(n11410), .ZN(n11316) );
  NAND2_X1 U11205 ( .A1(n11411), .A2(n11412), .ZN(n11409) );
  NAND2_X1 U11206 ( .A1(a_12_), .A2(n11408), .ZN(n11317) );
  NAND2_X1 U11207 ( .A1(n11172), .A2(n11413), .ZN(n11408) );
  NAND2_X1 U11208 ( .A1(n11171), .A2(n11173), .ZN(n11413) );
  NAND2_X1 U11209 ( .A1(n11414), .A2(n11415), .ZN(n11173) );
  NAND2_X1 U11210 ( .A1(a_13_), .A2(b_27_), .ZN(n11415) );
  INV_X1 U11211 ( .A(n11416), .ZN(n11414) );
  XNOR2_X1 U11212 ( .A(n11417), .B(n11418), .ZN(n11171) );
  NAND2_X1 U11213 ( .A1(n11419), .A2(n11420), .ZN(n11417) );
  NAND2_X1 U11214 ( .A1(a_13_), .A2(n11416), .ZN(n11172) );
  NAND2_X1 U11215 ( .A1(n11180), .A2(n11421), .ZN(n11416) );
  NAND2_X1 U11216 ( .A1(n11179), .A2(n11181), .ZN(n11421) );
  NAND2_X1 U11217 ( .A1(n11422), .A2(n11423), .ZN(n11181) );
  NAND2_X1 U11218 ( .A1(a_14_), .A2(b_27_), .ZN(n11423) );
  INV_X1 U11219 ( .A(n11424), .ZN(n11422) );
  XOR2_X1 U11220 ( .A(n11425), .B(n11426), .Z(n11179) );
  XOR2_X1 U11221 ( .A(n11427), .B(n11428), .Z(n11425) );
  NOR2_X1 U11222 ( .A1(n9217), .A2(n9534), .ZN(n11428) );
  NAND2_X1 U11223 ( .A1(a_14_), .A2(n11424), .ZN(n11180) );
  NAND2_X1 U11224 ( .A1(n11429), .A2(n11430), .ZN(n11424) );
  NAND2_X1 U11225 ( .A1(n11431), .A2(a_15_), .ZN(n11430) );
  NOR2_X1 U11226 ( .A1(n11432), .A2(n11041), .ZN(n11431) );
  NOR2_X1 U11227 ( .A1(n11187), .A2(n11188), .ZN(n11432) );
  NAND2_X1 U11228 ( .A1(n11187), .A2(n11188), .ZN(n11429) );
  NAND2_X1 U11229 ( .A1(n11313), .A2(n11433), .ZN(n11188) );
  NAND2_X1 U11230 ( .A1(n11312), .A2(n11314), .ZN(n11433) );
  NAND2_X1 U11231 ( .A1(n11434), .A2(n11435), .ZN(n11314) );
  NAND2_X1 U11232 ( .A1(a_16_), .A2(b_27_), .ZN(n11435) );
  INV_X1 U11233 ( .A(n11436), .ZN(n11434) );
  XNOR2_X1 U11234 ( .A(n11437), .B(n11438), .ZN(n11312) );
  NAND2_X1 U11235 ( .A1(n11439), .A2(n11440), .ZN(n11437) );
  NAND2_X1 U11236 ( .A1(a_16_), .A2(n11436), .ZN(n11313) );
  NAND2_X1 U11237 ( .A1(n11200), .A2(n11441), .ZN(n11436) );
  NAND2_X1 U11238 ( .A1(n11199), .A2(n11201), .ZN(n11441) );
  NAND2_X1 U11239 ( .A1(n11442), .A2(n11443), .ZN(n11201) );
  NAND2_X1 U11240 ( .A1(a_17_), .A2(b_27_), .ZN(n11443) );
  INV_X1 U11241 ( .A(n11444), .ZN(n11442) );
  XNOR2_X1 U11242 ( .A(n11445), .B(n11446), .ZN(n11199) );
  NAND2_X1 U11243 ( .A1(n11447), .A2(n11448), .ZN(n11445) );
  NAND2_X1 U11244 ( .A1(a_17_), .A2(n11444), .ZN(n11200) );
  NAND2_X1 U11245 ( .A1(n11208), .A2(n11449), .ZN(n11444) );
  NAND2_X1 U11246 ( .A1(n11207), .A2(n11209), .ZN(n11449) );
  NAND2_X1 U11247 ( .A1(n11450), .A2(n11451), .ZN(n11209) );
  NAND2_X1 U11248 ( .A1(a_18_), .A2(b_27_), .ZN(n11451) );
  INV_X1 U11249 ( .A(n11452), .ZN(n11450) );
  XNOR2_X1 U11250 ( .A(n11453), .B(n11454), .ZN(n11207) );
  XOR2_X1 U11251 ( .A(n11455), .B(n11456), .Z(n11454) );
  NAND2_X1 U11252 ( .A1(a_19_), .A2(b_26_), .ZN(n11456) );
  NAND2_X1 U11253 ( .A1(a_18_), .A2(n11452), .ZN(n11208) );
  NAND2_X1 U11254 ( .A1(n11457), .A2(n11458), .ZN(n11452) );
  NAND2_X1 U11255 ( .A1(n11459), .A2(a_19_), .ZN(n11458) );
  NOR2_X1 U11256 ( .A1(n11460), .A2(n11041), .ZN(n11459) );
  NOR2_X1 U11257 ( .A1(n11215), .A2(n11216), .ZN(n11460) );
  NAND2_X1 U11258 ( .A1(n11215), .A2(n11216), .ZN(n11457) );
  NAND2_X1 U11259 ( .A1(n11309), .A2(n11461), .ZN(n11216) );
  NAND2_X1 U11260 ( .A1(n11308), .A2(n11310), .ZN(n11461) );
  NAND2_X1 U11261 ( .A1(n11462), .A2(n11463), .ZN(n11310) );
  NAND2_X1 U11262 ( .A1(a_20_), .A2(b_27_), .ZN(n11463) );
  INV_X1 U11263 ( .A(n11464), .ZN(n11462) );
  XNOR2_X1 U11264 ( .A(n11465), .B(n11466), .ZN(n11308) );
  NAND2_X1 U11265 ( .A1(n11467), .A2(n11468), .ZN(n11465) );
  NAND2_X1 U11266 ( .A1(a_20_), .A2(n11464), .ZN(n11309) );
  NAND2_X1 U11267 ( .A1(n11228), .A2(n11469), .ZN(n11464) );
  NAND2_X1 U11268 ( .A1(n11227), .A2(n11229), .ZN(n11469) );
  NAND2_X1 U11269 ( .A1(n11470), .A2(n11471), .ZN(n11229) );
  NAND2_X1 U11270 ( .A1(a_21_), .A2(b_27_), .ZN(n11471) );
  INV_X1 U11271 ( .A(n11472), .ZN(n11470) );
  XNOR2_X1 U11272 ( .A(n11473), .B(n11474), .ZN(n11227) );
  NAND2_X1 U11273 ( .A1(n11475), .A2(n11476), .ZN(n11473) );
  NAND2_X1 U11274 ( .A1(a_21_), .A2(n11472), .ZN(n11228) );
  NAND2_X1 U11275 ( .A1(n11236), .A2(n11477), .ZN(n11472) );
  NAND2_X1 U11276 ( .A1(n11235), .A2(n11237), .ZN(n11477) );
  NAND2_X1 U11277 ( .A1(n11478), .A2(n11479), .ZN(n11237) );
  NAND2_X1 U11278 ( .A1(a_22_), .A2(b_27_), .ZN(n11479) );
  INV_X1 U11279 ( .A(n11480), .ZN(n11478) );
  XOR2_X1 U11280 ( .A(n11481), .B(n11482), .Z(n11235) );
  XOR2_X1 U11281 ( .A(n11483), .B(n11484), .Z(n11481) );
  NOR2_X1 U11282 ( .A1(n9217), .A2(n10051), .ZN(n11484) );
  NAND2_X1 U11283 ( .A1(a_22_), .A2(n11480), .ZN(n11236) );
  NAND2_X1 U11284 ( .A1(n11485), .A2(n11486), .ZN(n11480) );
  NAND2_X1 U11285 ( .A1(n11487), .A2(a_23_), .ZN(n11486) );
  NOR2_X1 U11286 ( .A1(n11488), .A2(n11041), .ZN(n11487) );
  NOR2_X1 U11287 ( .A1(n11243), .A2(n11244), .ZN(n11488) );
  NAND2_X1 U11288 ( .A1(n11243), .A2(n11244), .ZN(n11485) );
  NAND2_X1 U11289 ( .A1(n11489), .A2(n11490), .ZN(n11244) );
  INV_X1 U11290 ( .A(n11491), .ZN(n11490) );
  NOR2_X1 U11291 ( .A1(n11492), .A2(n11493), .ZN(n11491) );
  NOR2_X1 U11292 ( .A1(n11305), .A2(n11303), .ZN(n11493) );
  INV_X1 U11293 ( .A(n11306), .ZN(n11492) );
  NOR2_X1 U11294 ( .A1(n10050), .A2(n11041), .ZN(n11306) );
  NAND2_X1 U11295 ( .A1(n11303), .A2(n11305), .ZN(n11489) );
  NAND2_X1 U11296 ( .A1(n11494), .A2(n11495), .ZN(n11305) );
  NAND2_X1 U11297 ( .A1(n11302), .A2(n11496), .ZN(n11495) );
  NAND2_X1 U11298 ( .A1(n11299), .A2(n11301), .ZN(n11496) );
  NOR2_X1 U11299 ( .A1(n10048), .A2(n11041), .ZN(n11302) );
  INV_X1 U11300 ( .A(n11497), .ZN(n11494) );
  NOR2_X1 U11301 ( .A1(n11301), .A2(n11299), .ZN(n11497) );
  XNOR2_X1 U11302 ( .A(n11498), .B(n11499), .ZN(n11299) );
  XNOR2_X1 U11303 ( .A(n11500), .B(n11501), .ZN(n11499) );
  NAND2_X1 U11304 ( .A1(n11502), .A2(n11503), .ZN(n11301) );
  INV_X1 U11305 ( .A(n11504), .ZN(n11503) );
  NOR2_X1 U11306 ( .A1(n11260), .A2(n11505), .ZN(n11504) );
  NOR2_X1 U11307 ( .A1(n11261), .A2(n11262), .ZN(n11505) );
  XNOR2_X1 U11308 ( .A(n11506), .B(n11507), .ZN(n11260) );
  NAND2_X1 U11309 ( .A1(n11508), .A2(n11509), .ZN(n11506) );
  NAND2_X1 U11310 ( .A1(n11262), .A2(n11261), .ZN(n11502) );
  NAND2_X1 U11311 ( .A1(a_26_), .A2(b_27_), .ZN(n11261) );
  NOR2_X1 U11312 ( .A1(n11510), .A2(n11511), .ZN(n11262) );
  NOR2_X1 U11313 ( .A1(n11267), .A2(n11512), .ZN(n11511) );
  NOR2_X1 U11314 ( .A1(n11269), .A2(n10031), .ZN(n11512) );
  XOR2_X1 U11315 ( .A(n11513), .B(n11514), .Z(n11267) );
  XOR2_X1 U11316 ( .A(n11515), .B(n11516), .Z(n11514) );
  NAND2_X1 U11317 ( .A1(b_26_), .A2(a_28_), .ZN(n11516) );
  INV_X1 U11318 ( .A(n11517), .ZN(n11510) );
  NAND2_X1 U11319 ( .A1(n10031), .A2(n11269), .ZN(n11517) );
  NAND2_X1 U11320 ( .A1(n11518), .A2(n11519), .ZN(n11269) );
  NAND2_X1 U11321 ( .A1(n11520), .A2(b_27_), .ZN(n11519) );
  NOR2_X1 U11322 ( .A1(n11521), .A2(n9136), .ZN(n11520) );
  NOR2_X1 U11323 ( .A1(n11275), .A2(n11277), .ZN(n11521) );
  NAND2_X1 U11324 ( .A1(n11275), .A2(n11277), .ZN(n11518) );
  NAND2_X1 U11325 ( .A1(n11522), .A2(n11523), .ZN(n11277) );
  NAND2_X1 U11326 ( .A1(n11524), .A2(b_27_), .ZN(n11523) );
  NOR2_X1 U11327 ( .A1(n11525), .A2(n9121), .ZN(n11524) );
  NOR2_X1 U11328 ( .A1(n11526), .A2(n11285), .ZN(n11525) );
  NAND2_X1 U11329 ( .A1(n11526), .A2(n11285), .ZN(n11522) );
  NAND2_X1 U11330 ( .A1(n11527), .A2(n11528), .ZN(n11285) );
  NAND2_X1 U11331 ( .A1(b_25_), .A2(n11529), .ZN(n11528) );
  NAND2_X1 U11332 ( .A1(n10486), .A2(n11530), .ZN(n11529) );
  NAND2_X1 U11333 ( .A1(a_31_), .A2(n9217), .ZN(n11530) );
  NAND2_X1 U11334 ( .A1(b_26_), .A2(n11531), .ZN(n11527) );
  NAND2_X1 U11335 ( .A1(n10489), .A2(n11532), .ZN(n11531) );
  NAND2_X1 U11336 ( .A1(a_30_), .A2(n9245), .ZN(n11532) );
  INV_X1 U11337 ( .A(n11286), .ZN(n11526) );
  NAND2_X1 U11338 ( .A1(n11533), .A2(n9025), .ZN(n11286) );
  NOR2_X1 U11339 ( .A1(n11041), .A2(n9217), .ZN(n11533) );
  XOR2_X1 U11340 ( .A(n11534), .B(n11535), .Z(n11275) );
  NOR2_X1 U11341 ( .A1(n9121), .A2(n9217), .ZN(n11535) );
  XNOR2_X1 U11342 ( .A(n11536), .B(n11537), .ZN(n11534) );
  NOR2_X1 U11343 ( .A1(n11041), .A2(n11274), .ZN(n10031) );
  XNOR2_X1 U11344 ( .A(n11538), .B(n11539), .ZN(n11303) );
  XNOR2_X1 U11345 ( .A(n11540), .B(n11541), .ZN(n11539) );
  XNOR2_X1 U11346 ( .A(n11542), .B(n11543), .ZN(n11243) );
  XNOR2_X1 U11347 ( .A(n11544), .B(n11545), .ZN(n11543) );
  XNOR2_X1 U11348 ( .A(n11546), .B(n11547), .ZN(n11215) );
  NAND2_X1 U11349 ( .A1(n11548), .A2(n11549), .ZN(n11546) );
  XNOR2_X1 U11350 ( .A(n11550), .B(n11551), .ZN(n11187) );
  NAND2_X1 U11351 ( .A1(n11552), .A2(n11553), .ZN(n11550) );
  XNOR2_X1 U11352 ( .A(n11554), .B(n11555), .ZN(n11159) );
  NAND2_X1 U11353 ( .A1(n11556), .A2(n11557), .ZN(n11554) );
  NOR2_X1 U11354 ( .A1(n11121), .A2(n11119), .ZN(n11365) );
  XOR2_X1 U11355 ( .A(n11558), .B(n11559), .Z(n11119) );
  XOR2_X1 U11356 ( .A(n11560), .B(n11561), .Z(n11559) );
  NAND2_X1 U11357 ( .A1(a_7_), .A2(b_26_), .ZN(n11561) );
  NAND2_X1 U11358 ( .A1(a_6_), .A2(b_27_), .ZN(n11121) );
  XOR2_X1 U11359 ( .A(n11562), .B(n11563), .Z(n11320) );
  XNOR2_X1 U11360 ( .A(n11564), .B(n11565), .ZN(n11563) );
  XNOR2_X1 U11361 ( .A(n11566), .B(n11567), .ZN(n11324) );
  XOR2_X1 U11362 ( .A(n11568), .B(n11569), .Z(n11566) );
  NOR2_X1 U11363 ( .A1(n9217), .A2(n10083), .ZN(n11569) );
  XNOR2_X1 U11364 ( .A(n11570), .B(n11571), .ZN(n11328) );
  XOR2_X1 U11365 ( .A(n11572), .B(n11573), .Z(n11571) );
  NAND2_X1 U11366 ( .A1(a_4_), .A2(b_26_), .ZN(n11573) );
  XNOR2_X1 U11367 ( .A(n11574), .B(n11575), .ZN(n11336) );
  XNOR2_X1 U11368 ( .A(n11576), .B(n11577), .ZN(n11574) );
  XNOR2_X1 U11369 ( .A(n11578), .B(n11579), .ZN(n11090) );
  XNOR2_X1 U11370 ( .A(n11580), .B(n11581), .ZN(n11578) );
  NAND2_X1 U11371 ( .A1(n10139), .A2(n10140), .ZN(n10141) );
  INV_X1 U11372 ( .A(n11582), .ZN(n10140) );
  NAND2_X1 U11373 ( .A1(n11583), .A2(n10301), .ZN(n11582) );
  NAND2_X1 U11374 ( .A1(n11584), .A2(n11585), .ZN(n11583) );
  INV_X1 U11375 ( .A(n11586), .ZN(n11585) );
  XOR2_X1 U11376 ( .A(n11587), .B(n11588), .Z(n11584) );
  NOR2_X1 U11377 ( .A1(n10311), .A2(n10310), .ZN(n10139) );
  NOR2_X1 U11378 ( .A1(n11589), .A2(n11590), .ZN(n10310) );
  INV_X1 U11379 ( .A(n11591), .ZN(n11590) );
  NAND2_X1 U11380 ( .A1(n11093), .A2(n11592), .ZN(n11591) );
  NAND2_X1 U11381 ( .A1(n11092), .A2(n11082), .ZN(n11592) );
  NOR2_X1 U11382 ( .A1(n10093), .A2(n9217), .ZN(n11093) );
  NOR2_X1 U11383 ( .A1(n11082), .A2(n11092), .ZN(n11589) );
  NOR2_X1 U11384 ( .A1(n11593), .A2(n11594), .ZN(n11092) );
  INV_X1 U11385 ( .A(n11595), .ZN(n11594) );
  NAND2_X1 U11386 ( .A1(n11581), .A2(n11596), .ZN(n11595) );
  NAND2_X1 U11387 ( .A1(n11579), .A2(n11580), .ZN(n11596) );
  NOR2_X1 U11388 ( .A1(n9983), .A2(n9217), .ZN(n11581) );
  NOR2_X1 U11389 ( .A1(n11579), .A2(n11580), .ZN(n11593) );
  NOR2_X1 U11390 ( .A1(n11597), .A2(n11598), .ZN(n11580) );
  INV_X1 U11391 ( .A(n11599), .ZN(n11598) );
  NAND2_X1 U11392 ( .A1(n11576), .A2(n11600), .ZN(n11599) );
  NAND2_X1 U11393 ( .A1(n11577), .A2(n11575), .ZN(n11600) );
  NOR2_X1 U11394 ( .A1(n10088), .A2(n9217), .ZN(n11576) );
  NOR2_X1 U11395 ( .A1(n11575), .A2(n11577), .ZN(n11597) );
  NOR2_X1 U11396 ( .A1(n11601), .A2(n11602), .ZN(n11577) );
  NOR2_X1 U11397 ( .A1(n11352), .A2(n11603), .ZN(n11602) );
  NOR2_X1 U11398 ( .A1(n11351), .A2(n11349), .ZN(n11603) );
  NAND2_X1 U11399 ( .A1(a_3_), .A2(b_26_), .ZN(n11352) );
  INV_X1 U11400 ( .A(n11604), .ZN(n11601) );
  NAND2_X1 U11401 ( .A1(n11349), .A2(n11351), .ZN(n11604) );
  NAND2_X1 U11402 ( .A1(n11605), .A2(n11606), .ZN(n11351) );
  NAND2_X1 U11403 ( .A1(n11607), .A2(a_4_), .ZN(n11606) );
  NOR2_X1 U11404 ( .A1(n11608), .A2(n9217), .ZN(n11607) );
  NOR2_X1 U11405 ( .A1(n11570), .A2(n11572), .ZN(n11608) );
  NAND2_X1 U11406 ( .A1(n11570), .A2(n11572), .ZN(n11605) );
  NAND2_X1 U11407 ( .A1(n11609), .A2(n11610), .ZN(n11572) );
  NAND2_X1 U11408 ( .A1(n11611), .A2(a_5_), .ZN(n11610) );
  NOR2_X1 U11409 ( .A1(n11612), .A2(n9217), .ZN(n11611) );
  NOR2_X1 U11410 ( .A1(n11568), .A2(n11567), .ZN(n11612) );
  NAND2_X1 U11411 ( .A1(n11567), .A2(n11568), .ZN(n11609) );
  NAND2_X1 U11412 ( .A1(n11613), .A2(n11614), .ZN(n11568) );
  NAND2_X1 U11413 ( .A1(n11564), .A2(n11615), .ZN(n11614) );
  NAND2_X1 U11414 ( .A1(n11616), .A2(n11617), .ZN(n11615) );
  INV_X1 U11415 ( .A(n11565), .ZN(n11617) );
  INV_X1 U11416 ( .A(n11562), .ZN(n11616) );
  NAND2_X1 U11417 ( .A1(n11618), .A2(n11619), .ZN(n11564) );
  NAND2_X1 U11418 ( .A1(n11620), .A2(a_7_), .ZN(n11619) );
  NOR2_X1 U11419 ( .A1(n11621), .A2(n9217), .ZN(n11620) );
  NOR2_X1 U11420 ( .A1(n11560), .A2(n11558), .ZN(n11621) );
  NAND2_X1 U11421 ( .A1(n11558), .A2(n11560), .ZN(n11618) );
  NAND2_X1 U11422 ( .A1(n11622), .A2(n11623), .ZN(n11560) );
  NAND2_X1 U11423 ( .A1(n11624), .A2(a_8_), .ZN(n11623) );
  NOR2_X1 U11424 ( .A1(n11625), .A2(n9217), .ZN(n11624) );
  NOR2_X1 U11425 ( .A1(n11373), .A2(n11375), .ZN(n11625) );
  NAND2_X1 U11426 ( .A1(n11373), .A2(n11375), .ZN(n11622) );
  NAND2_X1 U11427 ( .A1(n11626), .A2(n11627), .ZN(n11375) );
  NAND2_X1 U11428 ( .A1(n11628), .A2(a_9_), .ZN(n11627) );
  NOR2_X1 U11429 ( .A1(n11629), .A2(n9217), .ZN(n11628) );
  NOR2_X1 U11430 ( .A1(n11383), .A2(n11382), .ZN(n11629) );
  NAND2_X1 U11431 ( .A1(n11383), .A2(n11382), .ZN(n11626) );
  XOR2_X1 U11432 ( .A(n11630), .B(n11631), .Z(n11382) );
  XOR2_X1 U11433 ( .A(n11632), .B(n11633), .Z(n11631) );
  NOR2_X1 U11434 ( .A1(n11634), .A2(n11635), .ZN(n11383) );
  INV_X1 U11435 ( .A(n11636), .ZN(n11635) );
  NAND2_X1 U11436 ( .A1(n11389), .A2(n11637), .ZN(n11636) );
  NAND2_X1 U11437 ( .A1(n11392), .A2(n11391), .ZN(n11637) );
  XNOR2_X1 U11438 ( .A(n11638), .B(n11639), .ZN(n11389) );
  XOR2_X1 U11439 ( .A(n11640), .B(n11641), .Z(n11638) );
  NOR2_X1 U11440 ( .A1(n9245), .A2(n9649), .ZN(n11641) );
  NOR2_X1 U11441 ( .A1(n11391), .A2(n11392), .ZN(n11634) );
  NOR2_X1 U11442 ( .A1(n10073), .A2(n9217), .ZN(n11392) );
  NAND2_X1 U11443 ( .A1(n11642), .A2(n11643), .ZN(n11391) );
  NAND2_X1 U11444 ( .A1(n11644), .A2(a_11_), .ZN(n11643) );
  NOR2_X1 U11445 ( .A1(n11645), .A2(n9217), .ZN(n11644) );
  NOR2_X1 U11446 ( .A1(n11397), .A2(n11399), .ZN(n11645) );
  NAND2_X1 U11447 ( .A1(n11397), .A2(n11399), .ZN(n11642) );
  NAND2_X1 U11448 ( .A1(n11556), .A2(n11646), .ZN(n11399) );
  NAND2_X1 U11449 ( .A1(n11555), .A2(n11557), .ZN(n11646) );
  NAND2_X1 U11450 ( .A1(n11647), .A2(n11648), .ZN(n11557) );
  NAND2_X1 U11451 ( .A1(a_12_), .A2(b_26_), .ZN(n11648) );
  INV_X1 U11452 ( .A(n11649), .ZN(n11647) );
  XNOR2_X1 U11453 ( .A(n11650), .B(n11651), .ZN(n11555) );
  NAND2_X1 U11454 ( .A1(n11652), .A2(n11653), .ZN(n11650) );
  NAND2_X1 U11455 ( .A1(a_12_), .A2(n11649), .ZN(n11556) );
  NAND2_X1 U11456 ( .A1(n11411), .A2(n11654), .ZN(n11649) );
  NAND2_X1 U11457 ( .A1(n11410), .A2(n11412), .ZN(n11654) );
  NAND2_X1 U11458 ( .A1(n11655), .A2(n11656), .ZN(n11412) );
  NAND2_X1 U11459 ( .A1(a_13_), .A2(b_26_), .ZN(n11656) );
  INV_X1 U11460 ( .A(n11657), .ZN(n11655) );
  XNOR2_X1 U11461 ( .A(n11658), .B(n11659), .ZN(n11410) );
  NAND2_X1 U11462 ( .A1(n11660), .A2(n11661), .ZN(n11658) );
  NAND2_X1 U11463 ( .A1(a_13_), .A2(n11657), .ZN(n11411) );
  NAND2_X1 U11464 ( .A1(n11419), .A2(n11662), .ZN(n11657) );
  NAND2_X1 U11465 ( .A1(n11418), .A2(n11420), .ZN(n11662) );
  NAND2_X1 U11466 ( .A1(n11663), .A2(n11664), .ZN(n11420) );
  NAND2_X1 U11467 ( .A1(a_14_), .A2(b_26_), .ZN(n11664) );
  INV_X1 U11468 ( .A(n11665), .ZN(n11663) );
  XNOR2_X1 U11469 ( .A(n11666), .B(n11667), .ZN(n11418) );
  XOR2_X1 U11470 ( .A(n11668), .B(n11669), .Z(n11667) );
  NAND2_X1 U11471 ( .A1(a_15_), .A2(b_25_), .ZN(n11669) );
  NAND2_X1 U11472 ( .A1(a_14_), .A2(n11665), .ZN(n11419) );
  NAND2_X1 U11473 ( .A1(n11670), .A2(n11671), .ZN(n11665) );
  NAND2_X1 U11474 ( .A1(n11672), .A2(a_15_), .ZN(n11671) );
  NOR2_X1 U11475 ( .A1(n11673), .A2(n9217), .ZN(n11672) );
  NOR2_X1 U11476 ( .A1(n11426), .A2(n11427), .ZN(n11673) );
  NAND2_X1 U11477 ( .A1(n11426), .A2(n11427), .ZN(n11670) );
  NAND2_X1 U11478 ( .A1(n11552), .A2(n11674), .ZN(n11427) );
  NAND2_X1 U11479 ( .A1(n11551), .A2(n11553), .ZN(n11674) );
  NAND2_X1 U11480 ( .A1(n11675), .A2(n11676), .ZN(n11553) );
  NAND2_X1 U11481 ( .A1(a_16_), .A2(b_26_), .ZN(n11676) );
  INV_X1 U11482 ( .A(n11677), .ZN(n11675) );
  XNOR2_X1 U11483 ( .A(n11678), .B(n11679), .ZN(n11551) );
  NAND2_X1 U11484 ( .A1(n11680), .A2(n11681), .ZN(n11678) );
  NAND2_X1 U11485 ( .A1(a_16_), .A2(n11677), .ZN(n11552) );
  NAND2_X1 U11486 ( .A1(n11439), .A2(n11682), .ZN(n11677) );
  NAND2_X1 U11487 ( .A1(n11438), .A2(n11440), .ZN(n11682) );
  NAND2_X1 U11488 ( .A1(n11683), .A2(n11684), .ZN(n11440) );
  NAND2_X1 U11489 ( .A1(a_17_), .A2(b_26_), .ZN(n11684) );
  INV_X1 U11490 ( .A(n11685), .ZN(n11683) );
  XNOR2_X1 U11491 ( .A(n11686), .B(n11687), .ZN(n11438) );
  XOR2_X1 U11492 ( .A(n11688), .B(n11689), .Z(n11686) );
  NAND2_X1 U11493 ( .A1(a_17_), .A2(n11685), .ZN(n11439) );
  NAND2_X1 U11494 ( .A1(n11447), .A2(n11690), .ZN(n11685) );
  NAND2_X1 U11495 ( .A1(n11446), .A2(n11448), .ZN(n11690) );
  NAND2_X1 U11496 ( .A1(n11691), .A2(n11692), .ZN(n11448) );
  NAND2_X1 U11497 ( .A1(a_18_), .A2(b_26_), .ZN(n11692) );
  INV_X1 U11498 ( .A(n11693), .ZN(n11691) );
  XNOR2_X1 U11499 ( .A(n11694), .B(n11695), .ZN(n11446) );
  XOR2_X1 U11500 ( .A(n11696), .B(n11697), .Z(n11695) );
  NAND2_X1 U11501 ( .A1(a_19_), .A2(b_25_), .ZN(n11697) );
  NAND2_X1 U11502 ( .A1(a_18_), .A2(n11693), .ZN(n11447) );
  NAND2_X1 U11503 ( .A1(n11698), .A2(n11699), .ZN(n11693) );
  NAND2_X1 U11504 ( .A1(n11700), .A2(a_19_), .ZN(n11699) );
  NOR2_X1 U11505 ( .A1(n11701), .A2(n9217), .ZN(n11700) );
  NOR2_X1 U11506 ( .A1(n11453), .A2(n11455), .ZN(n11701) );
  NAND2_X1 U11507 ( .A1(n11453), .A2(n11455), .ZN(n11698) );
  NAND2_X1 U11508 ( .A1(n11548), .A2(n11702), .ZN(n11455) );
  NAND2_X1 U11509 ( .A1(n11547), .A2(n11549), .ZN(n11702) );
  NAND2_X1 U11510 ( .A1(n11703), .A2(n11704), .ZN(n11549) );
  NAND2_X1 U11511 ( .A1(a_20_), .A2(b_26_), .ZN(n11704) );
  INV_X1 U11512 ( .A(n11705), .ZN(n11703) );
  XNOR2_X1 U11513 ( .A(n11706), .B(n11707), .ZN(n11547) );
  NAND2_X1 U11514 ( .A1(n11708), .A2(n11709), .ZN(n11706) );
  NAND2_X1 U11515 ( .A1(a_20_), .A2(n11705), .ZN(n11548) );
  NAND2_X1 U11516 ( .A1(n11467), .A2(n11710), .ZN(n11705) );
  NAND2_X1 U11517 ( .A1(n11466), .A2(n11468), .ZN(n11710) );
  NAND2_X1 U11518 ( .A1(n11711), .A2(n11712), .ZN(n11468) );
  NAND2_X1 U11519 ( .A1(a_21_), .A2(b_26_), .ZN(n11712) );
  INV_X1 U11520 ( .A(n11713), .ZN(n11711) );
  XNOR2_X1 U11521 ( .A(n11714), .B(n11715), .ZN(n11466) );
  NAND2_X1 U11522 ( .A1(n11716), .A2(n11717), .ZN(n11714) );
  NAND2_X1 U11523 ( .A1(a_21_), .A2(n11713), .ZN(n11467) );
  NAND2_X1 U11524 ( .A1(n11475), .A2(n11718), .ZN(n11713) );
  NAND2_X1 U11525 ( .A1(n11474), .A2(n11476), .ZN(n11718) );
  NAND2_X1 U11526 ( .A1(n11719), .A2(n11720), .ZN(n11476) );
  NAND2_X1 U11527 ( .A1(a_22_), .A2(b_26_), .ZN(n11720) );
  INV_X1 U11528 ( .A(n11721), .ZN(n11719) );
  XNOR2_X1 U11529 ( .A(n11722), .B(n11723), .ZN(n11474) );
  XOR2_X1 U11530 ( .A(n11724), .B(n11725), .Z(n11723) );
  NAND2_X1 U11531 ( .A1(a_23_), .A2(b_25_), .ZN(n11725) );
  NAND2_X1 U11532 ( .A1(a_22_), .A2(n11721), .ZN(n11475) );
  NAND2_X1 U11533 ( .A1(n11726), .A2(n11727), .ZN(n11721) );
  NAND2_X1 U11534 ( .A1(n11728), .A2(a_23_), .ZN(n11727) );
  NOR2_X1 U11535 ( .A1(n11729), .A2(n9217), .ZN(n11728) );
  NOR2_X1 U11536 ( .A1(n11482), .A2(n11483), .ZN(n11729) );
  NAND2_X1 U11537 ( .A1(n11482), .A2(n11483), .ZN(n11726) );
  NAND2_X1 U11538 ( .A1(n11730), .A2(n11731), .ZN(n11483) );
  NAND2_X1 U11539 ( .A1(n11545), .A2(n11732), .ZN(n11731) );
  INV_X1 U11540 ( .A(n11733), .ZN(n11732) );
  NOR2_X1 U11541 ( .A1(n11544), .A2(n11542), .ZN(n11733) );
  NOR2_X1 U11542 ( .A1(n10050), .A2(n9217), .ZN(n11545) );
  NAND2_X1 U11543 ( .A1(n11542), .A2(n11544), .ZN(n11730) );
  NAND2_X1 U11544 ( .A1(n11734), .A2(n11735), .ZN(n11544) );
  NAND2_X1 U11545 ( .A1(n11541), .A2(n11736), .ZN(n11735) );
  NAND2_X1 U11546 ( .A1(n11538), .A2(n11540), .ZN(n11736) );
  NOR2_X1 U11547 ( .A1(n10048), .A2(n9217), .ZN(n11541) );
  INV_X1 U11548 ( .A(n11737), .ZN(n11734) );
  NOR2_X1 U11549 ( .A1(n11540), .A2(n11538), .ZN(n11737) );
  XNOR2_X1 U11550 ( .A(n11738), .B(n11739), .ZN(n11538) );
  XNOR2_X1 U11551 ( .A(n11740), .B(n11741), .ZN(n11739) );
  NAND2_X1 U11552 ( .A1(n11742), .A2(n11743), .ZN(n11540) );
  NAND2_X1 U11553 ( .A1(n11498), .A2(n11744), .ZN(n11743) );
  NAND2_X1 U11554 ( .A1(n11501), .A2(n11500), .ZN(n11744) );
  INV_X1 U11555 ( .A(n10028), .ZN(n11501) );
  XOR2_X1 U11556 ( .A(n11745), .B(n11746), .Z(n11498) );
  NAND2_X1 U11557 ( .A1(n11747), .A2(n11748), .ZN(n11745) );
  NAND2_X1 U11558 ( .A1(n11749), .A2(n10028), .ZN(n11742) );
  NAND2_X1 U11559 ( .A1(b_26_), .A2(a_26_), .ZN(n10028) );
  INV_X1 U11560 ( .A(n11500), .ZN(n11749) );
  NAND2_X1 U11561 ( .A1(n11508), .A2(n11750), .ZN(n11500) );
  NAND2_X1 U11562 ( .A1(n11507), .A2(n11509), .ZN(n11750) );
  NAND2_X1 U11563 ( .A1(n11751), .A2(n11752), .ZN(n11509) );
  NAND2_X1 U11564 ( .A1(b_26_), .A2(a_27_), .ZN(n11752) );
  INV_X1 U11565 ( .A(n11753), .ZN(n11751) );
  XNOR2_X1 U11566 ( .A(n11754), .B(n11755), .ZN(n11507) );
  XOR2_X1 U11567 ( .A(n11756), .B(n11757), .Z(n11755) );
  NAND2_X1 U11568 ( .A1(b_25_), .A2(a_28_), .ZN(n11757) );
  NAND2_X1 U11569 ( .A1(a_27_), .A2(n11753), .ZN(n11508) );
  NAND2_X1 U11570 ( .A1(n11758), .A2(n11759), .ZN(n11753) );
  NAND2_X1 U11571 ( .A1(n11760), .A2(b_26_), .ZN(n11759) );
  NOR2_X1 U11572 ( .A1(n11761), .A2(n9136), .ZN(n11760) );
  NOR2_X1 U11573 ( .A1(n11513), .A2(n11515), .ZN(n11761) );
  NAND2_X1 U11574 ( .A1(n11513), .A2(n11515), .ZN(n11758) );
  NAND2_X1 U11575 ( .A1(n11762), .A2(n11763), .ZN(n11515) );
  NAND2_X1 U11576 ( .A1(n11764), .A2(b_26_), .ZN(n11763) );
  NOR2_X1 U11577 ( .A1(n11765), .A2(n9121), .ZN(n11764) );
  NOR2_X1 U11578 ( .A1(n11766), .A2(n11536), .ZN(n11765) );
  NAND2_X1 U11579 ( .A1(n11766), .A2(n11536), .ZN(n11762) );
  NAND2_X1 U11580 ( .A1(n11767), .A2(n11768), .ZN(n11536) );
  NAND2_X1 U11581 ( .A1(b_24_), .A2(n11769), .ZN(n11768) );
  NAND2_X1 U11582 ( .A1(n10486), .A2(n11770), .ZN(n11769) );
  NAND2_X1 U11583 ( .A1(a_31_), .A2(n9245), .ZN(n11770) );
  NAND2_X1 U11584 ( .A1(b_25_), .A2(n11771), .ZN(n11767) );
  NAND2_X1 U11585 ( .A1(n10489), .A2(n11772), .ZN(n11771) );
  NAND2_X1 U11586 ( .A1(a_30_), .A2(n10049), .ZN(n11772) );
  INV_X1 U11587 ( .A(n11537), .ZN(n11766) );
  NAND2_X1 U11588 ( .A1(n11773), .A2(n9025), .ZN(n11537) );
  NOR2_X1 U11589 ( .A1(n9217), .A2(n9245), .ZN(n11773) );
  XOR2_X1 U11590 ( .A(n11774), .B(n11775), .Z(n11513) );
  NOR2_X1 U11591 ( .A1(n9121), .A2(n9245), .ZN(n11775) );
  XNOR2_X1 U11592 ( .A(n11776), .B(n11777), .ZN(n11774) );
  XNOR2_X1 U11593 ( .A(n11778), .B(n11779), .ZN(n11542) );
  XOR2_X1 U11594 ( .A(n11780), .B(n10025), .Z(n11779) );
  XNOR2_X1 U11595 ( .A(n11781), .B(n11782), .ZN(n11482) );
  XNOR2_X1 U11596 ( .A(n11783), .B(n11784), .ZN(n11782) );
  XNOR2_X1 U11597 ( .A(n11785), .B(n11786), .ZN(n11453) );
  NAND2_X1 U11598 ( .A1(n11787), .A2(n11788), .ZN(n11785) );
  XNOR2_X1 U11599 ( .A(n11789), .B(n11790), .ZN(n11426) );
  NAND2_X1 U11600 ( .A1(n11791), .A2(n11792), .ZN(n11789) );
  XNOR2_X1 U11601 ( .A(n11793), .B(n11794), .ZN(n11397) );
  NAND2_X1 U11602 ( .A1(n11795), .A2(n11796), .ZN(n11793) );
  XOR2_X1 U11603 ( .A(n11797), .B(n11798), .Z(n11373) );
  XOR2_X1 U11604 ( .A(n11799), .B(n11800), .Z(n11797) );
  NOR2_X1 U11605 ( .A1(n9245), .A2(n10076), .ZN(n11800) );
  XNOR2_X1 U11606 ( .A(n11801), .B(n11802), .ZN(n11558) );
  XOR2_X1 U11607 ( .A(n11803), .B(n11804), .Z(n11802) );
  NAND2_X1 U11608 ( .A1(a_8_), .A2(b_25_), .ZN(n11804) );
  NAND2_X1 U11609 ( .A1(n11565), .A2(n11562), .ZN(n11613) );
  XNOR2_X1 U11610 ( .A(n11805), .B(n11806), .ZN(n11562) );
  XOR2_X1 U11611 ( .A(n11807), .B(n11808), .Z(n11806) );
  NAND2_X1 U11612 ( .A1(a_7_), .A2(b_25_), .ZN(n11808) );
  NOR2_X1 U11613 ( .A1(n10081), .A2(n9217), .ZN(n11565) );
  XNOR2_X1 U11614 ( .A(n11809), .B(n11810), .ZN(n11567) );
  NAND2_X1 U11615 ( .A1(n11811), .A2(n11812), .ZN(n11809) );
  XOR2_X1 U11616 ( .A(n11813), .B(n11814), .Z(n11570) );
  XOR2_X1 U11617 ( .A(n11815), .B(n11816), .Z(n11813) );
  NOR2_X1 U11618 ( .A1(n9245), .A2(n10083), .ZN(n11816) );
  XNOR2_X1 U11619 ( .A(n11817), .B(n11818), .ZN(n11349) );
  NAND2_X1 U11620 ( .A1(n11819), .A2(n11820), .ZN(n11817) );
  XNOR2_X1 U11621 ( .A(n11821), .B(n11822), .ZN(n11575) );
  XOR2_X1 U11622 ( .A(n11823), .B(n11824), .Z(n11821) );
  NOR2_X1 U11623 ( .A1(n9245), .A2(n10086), .ZN(n11824) );
  XOR2_X1 U11624 ( .A(n11825), .B(n11826), .Z(n11579) );
  XOR2_X1 U11625 ( .A(n11827), .B(n11828), .Z(n11826) );
  NAND2_X1 U11626 ( .A1(a_2_), .A2(b_25_), .ZN(n11828) );
  XOR2_X1 U11627 ( .A(n11829), .B(n11830), .Z(n11082) );
  XOR2_X1 U11628 ( .A(n11831), .B(n11832), .Z(n11830) );
  NAND2_X1 U11629 ( .A1(a_1_), .A2(b_25_), .ZN(n11832) );
  XOR2_X1 U11630 ( .A(n11833), .B(n11834), .Z(n10311) );
  XOR2_X1 U11631 ( .A(n11835), .B(n11836), .Z(n11834) );
  NAND2_X1 U11632 ( .A1(a_0_), .A2(b_25_), .ZN(n11836) );
  INV_X1 U11633 ( .A(n11837), .ZN(n10146) );
  NOR2_X1 U11634 ( .A1(n11838), .A2(n10301), .ZN(n11837) );
  NAND2_X1 U11635 ( .A1(n11839), .A2(n11586), .ZN(n10301) );
  NAND2_X1 U11636 ( .A1(n11840), .A2(n11841), .ZN(n11586) );
  NAND2_X1 U11637 ( .A1(n11842), .A2(a_0_), .ZN(n11841) );
  NOR2_X1 U11638 ( .A1(n11843), .A2(n9245), .ZN(n11842) );
  NOR2_X1 U11639 ( .A1(n11833), .A2(n11835), .ZN(n11843) );
  NAND2_X1 U11640 ( .A1(n11833), .A2(n11835), .ZN(n11840) );
  NAND2_X1 U11641 ( .A1(n11844), .A2(n11845), .ZN(n11835) );
  NAND2_X1 U11642 ( .A1(n11846), .A2(a_1_), .ZN(n11845) );
  NOR2_X1 U11643 ( .A1(n11847), .A2(n9245), .ZN(n11846) );
  NOR2_X1 U11644 ( .A1(n11829), .A2(n11831), .ZN(n11847) );
  NAND2_X1 U11645 ( .A1(n11829), .A2(n11831), .ZN(n11844) );
  NAND2_X1 U11646 ( .A1(n11848), .A2(n11849), .ZN(n11831) );
  NAND2_X1 U11647 ( .A1(n11850), .A2(a_2_), .ZN(n11849) );
  NOR2_X1 U11648 ( .A1(n11851), .A2(n9245), .ZN(n11850) );
  NOR2_X1 U11649 ( .A1(n11825), .A2(n11827), .ZN(n11851) );
  NAND2_X1 U11650 ( .A1(n11825), .A2(n11827), .ZN(n11848) );
  NAND2_X1 U11651 ( .A1(n11852), .A2(n11853), .ZN(n11827) );
  NAND2_X1 U11652 ( .A1(n11854), .A2(a_3_), .ZN(n11853) );
  NOR2_X1 U11653 ( .A1(n11855), .A2(n9245), .ZN(n11854) );
  NOR2_X1 U11654 ( .A1(n11822), .A2(n11823), .ZN(n11855) );
  NAND2_X1 U11655 ( .A1(n11822), .A2(n11823), .ZN(n11852) );
  NAND2_X1 U11656 ( .A1(n11819), .A2(n11856), .ZN(n11823) );
  NAND2_X1 U11657 ( .A1(n11818), .A2(n11820), .ZN(n11856) );
  NAND2_X1 U11658 ( .A1(n11857), .A2(n11858), .ZN(n11820) );
  NAND2_X1 U11659 ( .A1(a_4_), .A2(b_25_), .ZN(n11858) );
  INV_X1 U11660 ( .A(n11859), .ZN(n11857) );
  XOR2_X1 U11661 ( .A(n11860), .B(n11861), .Z(n11818) );
  XOR2_X1 U11662 ( .A(n11862), .B(n11863), .Z(n11860) );
  NAND2_X1 U11663 ( .A1(a_4_), .A2(n11859), .ZN(n11819) );
  NAND2_X1 U11664 ( .A1(n11864), .A2(n11865), .ZN(n11859) );
  NAND2_X1 U11665 ( .A1(n11866), .A2(a_5_), .ZN(n11865) );
  NOR2_X1 U11666 ( .A1(n11867), .A2(n9245), .ZN(n11866) );
  NOR2_X1 U11667 ( .A1(n11814), .A2(n11815), .ZN(n11867) );
  NAND2_X1 U11668 ( .A1(n11814), .A2(n11815), .ZN(n11864) );
  NAND2_X1 U11669 ( .A1(n11811), .A2(n11868), .ZN(n11815) );
  NAND2_X1 U11670 ( .A1(n11810), .A2(n11812), .ZN(n11868) );
  NAND2_X1 U11671 ( .A1(n11869), .A2(n11870), .ZN(n11812) );
  NAND2_X1 U11672 ( .A1(a_6_), .A2(b_25_), .ZN(n11870) );
  INV_X1 U11673 ( .A(n11871), .ZN(n11869) );
  XNOR2_X1 U11674 ( .A(n11872), .B(n11873), .ZN(n11810) );
  NAND2_X1 U11675 ( .A1(n11874), .A2(n11875), .ZN(n11872) );
  NAND2_X1 U11676 ( .A1(a_6_), .A2(n11871), .ZN(n11811) );
  NAND2_X1 U11677 ( .A1(n11876), .A2(n11877), .ZN(n11871) );
  NAND2_X1 U11678 ( .A1(n11878), .A2(a_7_), .ZN(n11877) );
  NOR2_X1 U11679 ( .A1(n11879), .A2(n9245), .ZN(n11878) );
  NOR2_X1 U11680 ( .A1(n11805), .A2(n11807), .ZN(n11879) );
  NAND2_X1 U11681 ( .A1(n11805), .A2(n11807), .ZN(n11876) );
  NAND2_X1 U11682 ( .A1(n11880), .A2(n11881), .ZN(n11807) );
  NAND2_X1 U11683 ( .A1(n11882), .A2(a_8_), .ZN(n11881) );
  NOR2_X1 U11684 ( .A1(n11883), .A2(n9245), .ZN(n11882) );
  NOR2_X1 U11685 ( .A1(n11801), .A2(n11803), .ZN(n11883) );
  NAND2_X1 U11686 ( .A1(n11801), .A2(n11803), .ZN(n11880) );
  NAND2_X1 U11687 ( .A1(n11884), .A2(n11885), .ZN(n11803) );
  NAND2_X1 U11688 ( .A1(n11886), .A2(a_9_), .ZN(n11885) );
  NOR2_X1 U11689 ( .A1(n11887), .A2(n9245), .ZN(n11886) );
  NOR2_X1 U11690 ( .A1(n11798), .A2(n11799), .ZN(n11887) );
  NAND2_X1 U11691 ( .A1(n11798), .A2(n11799), .ZN(n11884) );
  NAND2_X1 U11692 ( .A1(n11888), .A2(n11889), .ZN(n11799) );
  NAND2_X1 U11693 ( .A1(n11632), .A2(n11890), .ZN(n11889) );
  NAND2_X1 U11694 ( .A1(n11630), .A2(n11633), .ZN(n11890) );
  NAND2_X1 U11695 ( .A1(n11891), .A2(n11892), .ZN(n11632) );
  NAND2_X1 U11696 ( .A1(n11893), .A2(a_11_), .ZN(n11892) );
  NOR2_X1 U11697 ( .A1(n11894), .A2(n9245), .ZN(n11893) );
  NOR2_X1 U11698 ( .A1(n11639), .A2(n11640), .ZN(n11894) );
  NAND2_X1 U11699 ( .A1(n11639), .A2(n11640), .ZN(n11891) );
  NAND2_X1 U11700 ( .A1(n11795), .A2(n11895), .ZN(n11640) );
  NAND2_X1 U11701 ( .A1(n11794), .A2(n11796), .ZN(n11895) );
  NAND2_X1 U11702 ( .A1(n11896), .A2(n11897), .ZN(n11796) );
  NAND2_X1 U11703 ( .A1(a_12_), .A2(b_25_), .ZN(n11897) );
  INV_X1 U11704 ( .A(n11898), .ZN(n11896) );
  XNOR2_X1 U11705 ( .A(n11899), .B(n11900), .ZN(n11794) );
  NAND2_X1 U11706 ( .A1(n11901), .A2(n11902), .ZN(n11899) );
  NAND2_X1 U11707 ( .A1(a_12_), .A2(n11898), .ZN(n11795) );
  NAND2_X1 U11708 ( .A1(n11652), .A2(n11903), .ZN(n11898) );
  NAND2_X1 U11709 ( .A1(n11651), .A2(n11653), .ZN(n11903) );
  NAND2_X1 U11710 ( .A1(n11904), .A2(n11905), .ZN(n11653) );
  NAND2_X1 U11711 ( .A1(a_13_), .A2(b_25_), .ZN(n11905) );
  INV_X1 U11712 ( .A(n11906), .ZN(n11904) );
  XOR2_X1 U11713 ( .A(n11907), .B(n11908), .Z(n11651) );
  XNOR2_X1 U11714 ( .A(n11909), .B(n11910), .ZN(n11908) );
  NAND2_X1 U11715 ( .A1(a_13_), .A2(n11906), .ZN(n11652) );
  NAND2_X1 U11716 ( .A1(n11660), .A2(n11911), .ZN(n11906) );
  NAND2_X1 U11717 ( .A1(n11659), .A2(n11661), .ZN(n11911) );
  NAND2_X1 U11718 ( .A1(n11912), .A2(n11913), .ZN(n11661) );
  NAND2_X1 U11719 ( .A1(a_14_), .A2(b_25_), .ZN(n11913) );
  INV_X1 U11720 ( .A(n11914), .ZN(n11912) );
  XOR2_X1 U11721 ( .A(n11915), .B(n11916), .Z(n11659) );
  XNOR2_X1 U11722 ( .A(n11917), .B(n11918), .ZN(n11916) );
  NAND2_X1 U11723 ( .A1(a_15_), .A2(b_24_), .ZN(n11918) );
  NAND2_X1 U11724 ( .A1(a_14_), .A2(n11914), .ZN(n11660) );
  NAND2_X1 U11725 ( .A1(n11919), .A2(n11920), .ZN(n11914) );
  NAND2_X1 U11726 ( .A1(n11921), .A2(a_15_), .ZN(n11920) );
  NOR2_X1 U11727 ( .A1(n11922), .A2(n9245), .ZN(n11921) );
  NOR2_X1 U11728 ( .A1(n11666), .A2(n11668), .ZN(n11922) );
  NAND2_X1 U11729 ( .A1(n11666), .A2(n11668), .ZN(n11919) );
  NAND2_X1 U11730 ( .A1(n11791), .A2(n11923), .ZN(n11668) );
  NAND2_X1 U11731 ( .A1(n11790), .A2(n11792), .ZN(n11923) );
  NAND2_X1 U11732 ( .A1(n11924), .A2(n11925), .ZN(n11792) );
  NAND2_X1 U11733 ( .A1(a_16_), .A2(b_25_), .ZN(n11925) );
  INV_X1 U11734 ( .A(n11926), .ZN(n11924) );
  XNOR2_X1 U11735 ( .A(n11927), .B(n11928), .ZN(n11790) );
  XNOR2_X1 U11736 ( .A(n11929), .B(n11930), .ZN(n11927) );
  NAND2_X1 U11737 ( .A1(a_16_), .A2(n11926), .ZN(n11791) );
  NAND2_X1 U11738 ( .A1(n11680), .A2(n11931), .ZN(n11926) );
  NAND2_X1 U11739 ( .A1(n11679), .A2(n11681), .ZN(n11931) );
  NAND2_X1 U11740 ( .A1(n11932), .A2(n11933), .ZN(n11681) );
  NAND2_X1 U11741 ( .A1(a_17_), .A2(b_25_), .ZN(n11932) );
  XNOR2_X1 U11742 ( .A(n11934), .B(n11935), .ZN(n11679) );
  XOR2_X1 U11743 ( .A(n11936), .B(n11937), .Z(n11934) );
  NAND2_X1 U11744 ( .A1(n11938), .A2(a_17_), .ZN(n11680) );
  INV_X1 U11745 ( .A(n11933), .ZN(n11938) );
  NAND2_X1 U11746 ( .A1(n11939), .A2(n11940), .ZN(n11933) );
  NAND2_X1 U11747 ( .A1(n11687), .A2(n11941), .ZN(n11940) );
  NAND2_X1 U11748 ( .A1(n11689), .A2(n11688), .ZN(n11941) );
  XNOR2_X1 U11749 ( .A(n11942), .B(n11943), .ZN(n11687) );
  XOR2_X1 U11750 ( .A(n11944), .B(n11945), .Z(n11942) );
  INV_X1 U11751 ( .A(n11946), .ZN(n11939) );
  NOR2_X1 U11752 ( .A1(n11688), .A2(n11689), .ZN(n11946) );
  NOR2_X1 U11753 ( .A1(n10058), .A2(n9245), .ZN(n11689) );
  NAND2_X1 U11754 ( .A1(n11947), .A2(n11948), .ZN(n11688) );
  NAND2_X1 U11755 ( .A1(n11949), .A2(a_19_), .ZN(n11948) );
  NOR2_X1 U11756 ( .A1(n11950), .A2(n9245), .ZN(n11949) );
  NOR2_X1 U11757 ( .A1(n11694), .A2(n11696), .ZN(n11950) );
  NAND2_X1 U11758 ( .A1(n11694), .A2(n11696), .ZN(n11947) );
  NAND2_X1 U11759 ( .A1(n11787), .A2(n11951), .ZN(n11696) );
  NAND2_X1 U11760 ( .A1(n11786), .A2(n11788), .ZN(n11951) );
  NAND2_X1 U11761 ( .A1(n11952), .A2(n11953), .ZN(n11788) );
  NAND2_X1 U11762 ( .A1(a_20_), .A2(b_25_), .ZN(n11953) );
  INV_X1 U11763 ( .A(n11954), .ZN(n11952) );
  XNOR2_X1 U11764 ( .A(n11955), .B(n11956), .ZN(n11786) );
  NAND2_X1 U11765 ( .A1(n11957), .A2(n11958), .ZN(n11955) );
  NAND2_X1 U11766 ( .A1(a_20_), .A2(n11954), .ZN(n11787) );
  NAND2_X1 U11767 ( .A1(n11708), .A2(n11959), .ZN(n11954) );
  NAND2_X1 U11768 ( .A1(n11707), .A2(n11709), .ZN(n11959) );
  NAND2_X1 U11769 ( .A1(n11960), .A2(n11961), .ZN(n11709) );
  NAND2_X1 U11770 ( .A1(a_21_), .A2(b_25_), .ZN(n11961) );
  INV_X1 U11771 ( .A(n11962), .ZN(n11960) );
  XNOR2_X1 U11772 ( .A(n11963), .B(n11964), .ZN(n11707) );
  NAND2_X1 U11773 ( .A1(n11965), .A2(n11966), .ZN(n11963) );
  NAND2_X1 U11774 ( .A1(a_21_), .A2(n11962), .ZN(n11708) );
  NAND2_X1 U11775 ( .A1(n11716), .A2(n11967), .ZN(n11962) );
  NAND2_X1 U11776 ( .A1(n11715), .A2(n11717), .ZN(n11967) );
  NAND2_X1 U11777 ( .A1(n11968), .A2(n11969), .ZN(n11717) );
  NAND2_X1 U11778 ( .A1(a_22_), .A2(b_25_), .ZN(n11969) );
  INV_X1 U11779 ( .A(n11970), .ZN(n11968) );
  XOR2_X1 U11780 ( .A(n11971), .B(n11972), .Z(n11715) );
  XOR2_X1 U11781 ( .A(n11973), .B(n11974), .Z(n11971) );
  NOR2_X1 U11782 ( .A1(n10049), .A2(n10051), .ZN(n11974) );
  NAND2_X1 U11783 ( .A1(a_22_), .A2(n11970), .ZN(n11716) );
  NAND2_X1 U11784 ( .A1(n11975), .A2(n11976), .ZN(n11970) );
  NAND2_X1 U11785 ( .A1(n11977), .A2(a_23_), .ZN(n11976) );
  NOR2_X1 U11786 ( .A1(n11978), .A2(n9245), .ZN(n11977) );
  NOR2_X1 U11787 ( .A1(n11722), .A2(n11724), .ZN(n11978) );
  NAND2_X1 U11788 ( .A1(n11722), .A2(n11724), .ZN(n11975) );
  NAND2_X1 U11789 ( .A1(n11979), .A2(n11980), .ZN(n11724) );
  NAND2_X1 U11790 ( .A1(n11784), .A2(n11981), .ZN(n11980) );
  NAND2_X1 U11791 ( .A1(n11781), .A2(n11783), .ZN(n11981) );
  NOR2_X1 U11792 ( .A1(n10050), .A2(n9245), .ZN(n11784) );
  INV_X1 U11793 ( .A(n11982), .ZN(n11979) );
  NOR2_X1 U11794 ( .A1(n11783), .A2(n11781), .ZN(n11982) );
  XNOR2_X1 U11795 ( .A(n11983), .B(n11984), .ZN(n11781) );
  XOR2_X1 U11796 ( .A(n11985), .B(n11986), .Z(n11984) );
  NAND2_X1 U11797 ( .A1(n11987), .A2(n11988), .ZN(n11783) );
  NAND2_X1 U11798 ( .A1(n11778), .A2(n11989), .ZN(n11988) );
  INV_X1 U11799 ( .A(n11990), .ZN(n11989) );
  NOR2_X1 U11800 ( .A1(n11780), .A2(n10025), .ZN(n11990) );
  XNOR2_X1 U11801 ( .A(n11991), .B(n11992), .ZN(n11778) );
  XNOR2_X1 U11802 ( .A(n11993), .B(n11994), .ZN(n11992) );
  NAND2_X1 U11803 ( .A1(n10025), .A2(n11780), .ZN(n11987) );
  NAND2_X1 U11804 ( .A1(n11995), .A2(n11996), .ZN(n11780) );
  NAND2_X1 U11805 ( .A1(n11738), .A2(n11997), .ZN(n11996) );
  NAND2_X1 U11806 ( .A1(n11741), .A2(n11740), .ZN(n11997) );
  XOR2_X1 U11807 ( .A(n11998), .B(n11999), .Z(n11738) );
  NAND2_X1 U11808 ( .A1(n12000), .A2(n12001), .ZN(n11998) );
  INV_X1 U11809 ( .A(n12002), .ZN(n11995) );
  NOR2_X1 U11810 ( .A1(n11740), .A2(n11741), .ZN(n12002) );
  NOR2_X1 U11811 ( .A1(n9245), .A2(n10047), .ZN(n11741) );
  NAND2_X1 U11812 ( .A1(n11747), .A2(n12003), .ZN(n11740) );
  NAND2_X1 U11813 ( .A1(n11746), .A2(n11748), .ZN(n12003) );
  NAND2_X1 U11814 ( .A1(n12004), .A2(n12005), .ZN(n11748) );
  NAND2_X1 U11815 ( .A1(b_25_), .A2(a_27_), .ZN(n12005) );
  INV_X1 U11816 ( .A(n12006), .ZN(n12004) );
  XNOR2_X1 U11817 ( .A(n12007), .B(n12008), .ZN(n11746) );
  XOR2_X1 U11818 ( .A(n12009), .B(n12010), .Z(n12008) );
  NAND2_X1 U11819 ( .A1(a_28_), .A2(b_24_), .ZN(n12010) );
  NAND2_X1 U11820 ( .A1(a_27_), .A2(n12006), .ZN(n11747) );
  NAND2_X1 U11821 ( .A1(n12011), .A2(n12012), .ZN(n12006) );
  NAND2_X1 U11822 ( .A1(n12013), .A2(b_25_), .ZN(n12012) );
  NOR2_X1 U11823 ( .A1(n12014), .A2(n9136), .ZN(n12013) );
  NOR2_X1 U11824 ( .A1(n11754), .A2(n11756), .ZN(n12014) );
  NAND2_X1 U11825 ( .A1(n11754), .A2(n11756), .ZN(n12011) );
  NAND2_X1 U11826 ( .A1(n12015), .A2(n12016), .ZN(n11756) );
  NAND2_X1 U11827 ( .A1(n12017), .A2(b_25_), .ZN(n12016) );
  NOR2_X1 U11828 ( .A1(n12018), .A2(n9121), .ZN(n12017) );
  NOR2_X1 U11829 ( .A1(n12019), .A2(n11776), .ZN(n12018) );
  NAND2_X1 U11830 ( .A1(n12019), .A2(n11776), .ZN(n12015) );
  NAND2_X1 U11831 ( .A1(n12020), .A2(n12021), .ZN(n11776) );
  NAND2_X1 U11832 ( .A1(b_23_), .A2(n12022), .ZN(n12021) );
  NAND2_X1 U11833 ( .A1(n10486), .A2(n12023), .ZN(n12022) );
  NAND2_X1 U11834 ( .A1(a_31_), .A2(n10049), .ZN(n12023) );
  NAND2_X1 U11835 ( .A1(b_24_), .A2(n12024), .ZN(n12020) );
  NAND2_X1 U11836 ( .A1(n10489), .A2(n12025), .ZN(n12024) );
  NAND2_X1 U11837 ( .A1(a_30_), .A2(n9302), .ZN(n12025) );
  INV_X1 U11838 ( .A(n11777), .ZN(n12019) );
  NAND2_X1 U11839 ( .A1(n12026), .A2(n9025), .ZN(n11777) );
  NOR2_X1 U11840 ( .A1(n10049), .A2(n9245), .ZN(n12026) );
  XOR2_X1 U11841 ( .A(n12027), .B(n12028), .Z(n11754) );
  NOR2_X1 U11842 ( .A1(n10049), .A2(n9121), .ZN(n12028) );
  XNOR2_X1 U11843 ( .A(n12029), .B(n12030), .ZN(n12027) );
  NAND2_X1 U11844 ( .A1(b_25_), .A2(a_25_), .ZN(n10025) );
  XNOR2_X1 U11845 ( .A(n12031), .B(n12032), .ZN(n11722) );
  XNOR2_X1 U11846 ( .A(n12033), .B(n12034), .ZN(n12032) );
  XNOR2_X1 U11847 ( .A(n12035), .B(n12036), .ZN(n11694) );
  XOR2_X1 U11848 ( .A(n12037), .B(n12038), .Z(n12035) );
  XNOR2_X1 U11849 ( .A(n12039), .B(n12040), .ZN(n11666) );
  XOR2_X1 U11850 ( .A(n12041), .B(n12042), .Z(n12039) );
  XNOR2_X1 U11851 ( .A(n12043), .B(n12044), .ZN(n11639) );
  XOR2_X1 U11852 ( .A(n12045), .B(n12046), .Z(n12044) );
  NAND2_X1 U11853 ( .A1(a_12_), .A2(b_24_), .ZN(n12046) );
  INV_X1 U11854 ( .A(n12047), .ZN(n11888) );
  NOR2_X1 U11855 ( .A1(n11633), .A2(n11630), .ZN(n12047) );
  XNOR2_X1 U11856 ( .A(n12048), .B(n12049), .ZN(n11630) );
  XOR2_X1 U11857 ( .A(n12050), .B(n12051), .Z(n12048) );
  NOR2_X1 U11858 ( .A1(n10049), .A2(n9649), .ZN(n12051) );
  NAND2_X1 U11859 ( .A1(a_10_), .A2(b_25_), .ZN(n11633) );
  XNOR2_X1 U11860 ( .A(n12052), .B(n12053), .ZN(n11798) );
  NAND2_X1 U11861 ( .A1(n12054), .A2(n12055), .ZN(n12052) );
  XOR2_X1 U11862 ( .A(n12056), .B(n12057), .Z(n11801) );
  XOR2_X1 U11863 ( .A(n12058), .B(n12059), .Z(n12056) );
  NOR2_X1 U11864 ( .A1(n10049), .A2(n10076), .ZN(n12059) );
  XNOR2_X1 U11865 ( .A(n12060), .B(n12061), .ZN(n11805) );
  XOR2_X1 U11866 ( .A(n12062), .B(n12063), .Z(n12061) );
  NAND2_X1 U11867 ( .A1(a_8_), .A2(b_24_), .ZN(n12063) );
  XOR2_X1 U11868 ( .A(n12064), .B(n12065), .Z(n11814) );
  XOR2_X1 U11869 ( .A(n12066), .B(n12067), .Z(n12064) );
  XOR2_X1 U11870 ( .A(n12068), .B(n12069), .Z(n11822) );
  XNOR2_X1 U11871 ( .A(n12070), .B(n12071), .ZN(n12068) );
  NAND2_X1 U11872 ( .A1(a_4_), .A2(b_24_), .ZN(n12070) );
  XNOR2_X1 U11873 ( .A(n12072), .B(n12073), .ZN(n11825) );
  NAND2_X1 U11874 ( .A1(n12074), .A2(n12075), .ZN(n12072) );
  XNOR2_X1 U11875 ( .A(n12076), .B(n12077), .ZN(n11829) );
  NAND2_X1 U11876 ( .A1(n12078), .A2(n12079), .ZN(n12076) );
  XNOR2_X1 U11877 ( .A(n12080), .B(n12081), .ZN(n11833) );
  XOR2_X1 U11878 ( .A(n12082), .B(n12083), .Z(n12081) );
  NAND2_X1 U11879 ( .A1(a_1_), .A2(b_24_), .ZN(n12083) );
  XNOR2_X1 U11880 ( .A(n11587), .B(n11588), .ZN(n11839) );
  NAND2_X1 U11881 ( .A1(n12084), .A2(n12085), .ZN(n11587) );
  NAND2_X1 U11882 ( .A1(n10298), .A2(n12086), .ZN(n11838) );
  INV_X1 U11883 ( .A(n12087), .ZN(n12086) );
  NOR2_X1 U11884 ( .A1(n10303), .A2(n10302), .ZN(n12087) );
  INV_X1 U11885 ( .A(n12088), .ZN(n10153) );
  NOR2_X1 U11886 ( .A1(n10298), .A2(n10297), .ZN(n12088) );
  NAND2_X1 U11887 ( .A1(n10293), .A2(n12089), .ZN(n10297) );
  NAND2_X1 U11888 ( .A1(n12090), .A2(n12091), .ZN(n12089) );
  INV_X1 U11889 ( .A(n12092), .ZN(n12091) );
  XNOR2_X1 U11890 ( .A(n12093), .B(n12094), .ZN(n12090) );
  NAND2_X1 U11891 ( .A1(n10303), .A2(n10302), .ZN(n10298) );
  NAND2_X1 U11892 ( .A1(n12084), .A2(n12095), .ZN(n10302) );
  NAND2_X1 U11893 ( .A1(n11588), .A2(n12085), .ZN(n12095) );
  NAND2_X1 U11894 ( .A1(n12096), .A2(n12097), .ZN(n12085) );
  NAND2_X1 U11895 ( .A1(a_0_), .A2(b_24_), .ZN(n12097) );
  INV_X1 U11896 ( .A(n12098), .ZN(n12096) );
  XOR2_X1 U11897 ( .A(n12099), .B(n12100), .Z(n11588) );
  XOR2_X1 U11898 ( .A(n12101), .B(n12102), .Z(n12099) );
  NOR2_X1 U11899 ( .A1(n9302), .A2(n9983), .ZN(n12102) );
  NAND2_X1 U11900 ( .A1(a_0_), .A2(n12098), .ZN(n12084) );
  NAND2_X1 U11901 ( .A1(n12103), .A2(n12104), .ZN(n12098) );
  NAND2_X1 U11902 ( .A1(n12105), .A2(a_1_), .ZN(n12104) );
  NOR2_X1 U11903 ( .A1(n12106), .A2(n10049), .ZN(n12105) );
  NOR2_X1 U11904 ( .A1(n12080), .A2(n12082), .ZN(n12106) );
  NAND2_X1 U11905 ( .A1(n12080), .A2(n12082), .ZN(n12103) );
  NAND2_X1 U11906 ( .A1(n12078), .A2(n12107), .ZN(n12082) );
  NAND2_X1 U11907 ( .A1(n12077), .A2(n12079), .ZN(n12107) );
  NAND2_X1 U11908 ( .A1(n12108), .A2(n12109), .ZN(n12079) );
  NAND2_X1 U11909 ( .A1(a_2_), .A2(b_24_), .ZN(n12109) );
  INV_X1 U11910 ( .A(n12110), .ZN(n12108) );
  XOR2_X1 U11911 ( .A(n12111), .B(n12112), .Z(n12077) );
  XNOR2_X1 U11912 ( .A(n12113), .B(n12114), .ZN(n12112) );
  NAND2_X1 U11913 ( .A1(a_2_), .A2(n12110), .ZN(n12078) );
  NAND2_X1 U11914 ( .A1(n12074), .A2(n12115), .ZN(n12110) );
  NAND2_X1 U11915 ( .A1(n12073), .A2(n12075), .ZN(n12115) );
  NAND2_X1 U11916 ( .A1(n12116), .A2(n12117), .ZN(n12075) );
  NAND2_X1 U11917 ( .A1(a_3_), .A2(b_24_), .ZN(n12117) );
  INV_X1 U11918 ( .A(n12118), .ZN(n12116) );
  XOR2_X1 U11919 ( .A(n12119), .B(n12120), .Z(n12073) );
  XOR2_X1 U11920 ( .A(n12121), .B(n12122), .Z(n12119) );
  NOR2_X1 U11921 ( .A1(n9302), .A2(n10085), .ZN(n12122) );
  NAND2_X1 U11922 ( .A1(a_3_), .A2(n12118), .ZN(n12074) );
  NAND2_X1 U11923 ( .A1(n12123), .A2(n12124), .ZN(n12118) );
  NAND2_X1 U11924 ( .A1(n12125), .A2(a_4_), .ZN(n12124) );
  NOR2_X1 U11925 ( .A1(n12126), .A2(n10049), .ZN(n12125) );
  NOR2_X1 U11926 ( .A1(n12069), .A2(n12071), .ZN(n12126) );
  NAND2_X1 U11927 ( .A1(n12069), .A2(n12071), .ZN(n12123) );
  NAND2_X1 U11928 ( .A1(n12127), .A2(n12128), .ZN(n12071) );
  NAND2_X1 U11929 ( .A1(n11863), .A2(n12129), .ZN(n12128) );
  INV_X1 U11930 ( .A(n12130), .ZN(n12129) );
  NOR2_X1 U11931 ( .A1(n11862), .A2(n11861), .ZN(n12130) );
  NOR2_X1 U11932 ( .A1(n10083), .A2(n10049), .ZN(n11863) );
  NAND2_X1 U11933 ( .A1(n11861), .A2(n11862), .ZN(n12127) );
  NAND2_X1 U11934 ( .A1(n12131), .A2(n12132), .ZN(n11862) );
  NAND2_X1 U11935 ( .A1(n12067), .A2(n12133), .ZN(n12132) );
  INV_X1 U11936 ( .A(n12134), .ZN(n12133) );
  NOR2_X1 U11937 ( .A1(n12066), .A2(n12065), .ZN(n12134) );
  NOR2_X1 U11938 ( .A1(n10081), .A2(n10049), .ZN(n12067) );
  NAND2_X1 U11939 ( .A1(n12065), .A2(n12066), .ZN(n12131) );
  NAND2_X1 U11940 ( .A1(n11874), .A2(n12135), .ZN(n12066) );
  NAND2_X1 U11941 ( .A1(n11873), .A2(n11875), .ZN(n12135) );
  NAND2_X1 U11942 ( .A1(n12136), .A2(n12137), .ZN(n11875) );
  NAND2_X1 U11943 ( .A1(a_7_), .A2(b_24_), .ZN(n12137) );
  INV_X1 U11944 ( .A(n12138), .ZN(n12136) );
  XNOR2_X1 U11945 ( .A(n12139), .B(n12140), .ZN(n11873) );
  XNOR2_X1 U11946 ( .A(n12141), .B(n12142), .ZN(n12140) );
  NAND2_X1 U11947 ( .A1(a_7_), .A2(n12138), .ZN(n11874) );
  NAND2_X1 U11948 ( .A1(n12143), .A2(n12144), .ZN(n12138) );
  NAND2_X1 U11949 ( .A1(n12145), .A2(a_8_), .ZN(n12144) );
  NOR2_X1 U11950 ( .A1(n12146), .A2(n10049), .ZN(n12145) );
  NOR2_X1 U11951 ( .A1(n12060), .A2(n12062), .ZN(n12146) );
  NAND2_X1 U11952 ( .A1(n12060), .A2(n12062), .ZN(n12143) );
  NAND2_X1 U11953 ( .A1(n12147), .A2(n12148), .ZN(n12062) );
  NAND2_X1 U11954 ( .A1(n12149), .A2(a_9_), .ZN(n12148) );
  NOR2_X1 U11955 ( .A1(n12150), .A2(n10049), .ZN(n12149) );
  NOR2_X1 U11956 ( .A1(n12057), .A2(n12058), .ZN(n12150) );
  NAND2_X1 U11957 ( .A1(n12057), .A2(n12058), .ZN(n12147) );
  NAND2_X1 U11958 ( .A1(n12054), .A2(n12151), .ZN(n12058) );
  NAND2_X1 U11959 ( .A1(n12053), .A2(n12055), .ZN(n12151) );
  NAND2_X1 U11960 ( .A1(n12152), .A2(n12153), .ZN(n12055) );
  NAND2_X1 U11961 ( .A1(a_10_), .A2(b_24_), .ZN(n12153) );
  INV_X1 U11962 ( .A(n12154), .ZN(n12152) );
  XOR2_X1 U11963 ( .A(n12155), .B(n12156), .Z(n12053) );
  XOR2_X1 U11964 ( .A(n12157), .B(n12158), .Z(n12155) );
  NOR2_X1 U11965 ( .A1(n9302), .A2(n9649), .ZN(n12158) );
  NAND2_X1 U11966 ( .A1(a_10_), .A2(n12154), .ZN(n12054) );
  NAND2_X1 U11967 ( .A1(n12159), .A2(n12160), .ZN(n12154) );
  NAND2_X1 U11968 ( .A1(n12161), .A2(a_11_), .ZN(n12160) );
  NOR2_X1 U11969 ( .A1(n12162), .A2(n10049), .ZN(n12161) );
  NOR2_X1 U11970 ( .A1(n12049), .A2(n12050), .ZN(n12162) );
  NAND2_X1 U11971 ( .A1(n12049), .A2(n12050), .ZN(n12159) );
  NAND2_X1 U11972 ( .A1(n12163), .A2(n12164), .ZN(n12050) );
  NAND2_X1 U11973 ( .A1(n12165), .A2(a_12_), .ZN(n12164) );
  NOR2_X1 U11974 ( .A1(n12166), .A2(n10049), .ZN(n12165) );
  NOR2_X1 U11975 ( .A1(n12043), .A2(n12045), .ZN(n12166) );
  NAND2_X1 U11976 ( .A1(n12043), .A2(n12045), .ZN(n12163) );
  NAND2_X1 U11977 ( .A1(n11901), .A2(n12167), .ZN(n12045) );
  NAND2_X1 U11978 ( .A1(n11900), .A2(n11902), .ZN(n12167) );
  NAND2_X1 U11979 ( .A1(n12168), .A2(n12169), .ZN(n11902) );
  NAND2_X1 U11980 ( .A1(a_13_), .A2(b_24_), .ZN(n12168) );
  XNOR2_X1 U11981 ( .A(n12170), .B(n12171), .ZN(n11900) );
  NAND2_X1 U11982 ( .A1(n12172), .A2(n12173), .ZN(n12170) );
  NAND2_X1 U11983 ( .A1(n12174), .A2(a_13_), .ZN(n11901) );
  INV_X1 U11984 ( .A(n12169), .ZN(n12174) );
  NAND2_X1 U11985 ( .A1(n12175), .A2(n12176), .ZN(n12169) );
  NAND2_X1 U11986 ( .A1(n11907), .A2(n12177), .ZN(n12176) );
  NAND2_X1 U11987 ( .A1(n11910), .A2(n11909), .ZN(n12177) );
  XNOR2_X1 U11988 ( .A(n12178), .B(n12179), .ZN(n11907) );
  XOR2_X1 U11989 ( .A(n12180), .B(n12181), .Z(n12178) );
  NOR2_X1 U11990 ( .A1(n9302), .A2(n9534), .ZN(n12181) );
  INV_X1 U11991 ( .A(n12182), .ZN(n12175) );
  NOR2_X1 U11992 ( .A1(n11909), .A2(n11910), .ZN(n12182) );
  NOR2_X1 U11993 ( .A1(n10065), .A2(n10049), .ZN(n11910) );
  NAND2_X1 U11994 ( .A1(n12183), .A2(n12184), .ZN(n11909) );
  NAND2_X1 U11995 ( .A1(n12185), .A2(a_15_), .ZN(n12184) );
  NOR2_X1 U11996 ( .A1(n12186), .A2(n10049), .ZN(n12185) );
  NOR2_X1 U11997 ( .A1(n11917), .A2(n11915), .ZN(n12186) );
  NAND2_X1 U11998 ( .A1(n11917), .A2(n11915), .ZN(n12183) );
  XNOR2_X1 U11999 ( .A(n12187), .B(n12188), .ZN(n11915) );
  NAND2_X1 U12000 ( .A1(n12189), .A2(n12190), .ZN(n12187) );
  NOR2_X1 U12001 ( .A1(n12191), .A2(n12192), .ZN(n11917) );
  INV_X1 U12002 ( .A(n12193), .ZN(n12192) );
  NAND2_X1 U12003 ( .A1(n12040), .A2(n12194), .ZN(n12193) );
  NAND2_X1 U12004 ( .A1(n12042), .A2(n12041), .ZN(n12194) );
  XOR2_X1 U12005 ( .A(n12195), .B(n12196), .Z(n12040) );
  NAND2_X1 U12006 ( .A1(n12197), .A2(n12198), .ZN(n12195) );
  NOR2_X1 U12007 ( .A1(n12041), .A2(n12042), .ZN(n12191) );
  NOR2_X1 U12008 ( .A1(n10062), .A2(n10049), .ZN(n12042) );
  NAND2_X1 U12009 ( .A1(n12199), .A2(n12200), .ZN(n12041) );
  NAND2_X1 U12010 ( .A1(n11930), .A2(n12201), .ZN(n12200) );
  INV_X1 U12011 ( .A(n12202), .ZN(n12201) );
  NOR2_X1 U12012 ( .A1(n11928), .A2(n11929), .ZN(n12202) );
  NOR2_X1 U12013 ( .A1(n10060), .A2(n10049), .ZN(n11930) );
  NAND2_X1 U12014 ( .A1(n11929), .A2(n11928), .ZN(n12199) );
  XNOR2_X1 U12015 ( .A(n12203), .B(n12204), .ZN(n11928) );
  NAND2_X1 U12016 ( .A1(n12205), .A2(n12206), .ZN(n12203) );
  NOR2_X1 U12017 ( .A1(n12207), .A2(n12208), .ZN(n11929) );
  INV_X1 U12018 ( .A(n12209), .ZN(n12208) );
  NAND2_X1 U12019 ( .A1(n11935), .A2(n12210), .ZN(n12209) );
  NAND2_X1 U12020 ( .A1(n11937), .A2(n11936), .ZN(n12210) );
  XOR2_X1 U12021 ( .A(n12211), .B(n12212), .Z(n11935) );
  XOR2_X1 U12022 ( .A(n12213), .B(n12214), .Z(n12212) );
  NAND2_X1 U12023 ( .A1(a_19_), .A2(b_23_), .ZN(n12214) );
  NOR2_X1 U12024 ( .A1(n11936), .A2(n11937), .ZN(n12207) );
  NOR2_X1 U12025 ( .A1(n10058), .A2(n10049), .ZN(n11937) );
  NAND2_X1 U12026 ( .A1(n12215), .A2(n12216), .ZN(n11936) );
  NAND2_X1 U12027 ( .A1(n11945), .A2(n12217), .ZN(n12216) );
  NAND2_X1 U12028 ( .A1(n11943), .A2(n11944), .ZN(n12217) );
  NOR2_X1 U12029 ( .A1(n9415), .A2(n10049), .ZN(n11945) );
  INV_X1 U12030 ( .A(n12218), .ZN(n12215) );
  NOR2_X1 U12031 ( .A1(n11944), .A2(n11943), .ZN(n12218) );
  XOR2_X1 U12032 ( .A(n12219), .B(n12220), .Z(n11943) );
  NAND2_X1 U12033 ( .A1(n12221), .A2(n12222), .ZN(n12219) );
  NAND2_X1 U12034 ( .A1(n12223), .A2(n12224), .ZN(n11944) );
  NAND2_X1 U12035 ( .A1(n12036), .A2(n12225), .ZN(n12224) );
  NAND2_X1 U12036 ( .A1(n12038), .A2(n12037), .ZN(n12225) );
  XOR2_X1 U12037 ( .A(n12226), .B(n12227), .Z(n12036) );
  NAND2_X1 U12038 ( .A1(n12228), .A2(n12229), .ZN(n12226) );
  INV_X1 U12039 ( .A(n12230), .ZN(n12223) );
  NOR2_X1 U12040 ( .A1(n12037), .A2(n12038), .ZN(n12230) );
  NOR2_X1 U12041 ( .A1(n10054), .A2(n10049), .ZN(n12038) );
  NAND2_X1 U12042 ( .A1(n11957), .A2(n12231), .ZN(n12037) );
  NAND2_X1 U12043 ( .A1(n11956), .A2(n11958), .ZN(n12231) );
  NAND2_X1 U12044 ( .A1(n12232), .A2(n12233), .ZN(n11958) );
  NAND2_X1 U12045 ( .A1(a_21_), .A2(b_24_), .ZN(n12233) );
  INV_X1 U12046 ( .A(n12234), .ZN(n12232) );
  XNOR2_X1 U12047 ( .A(n12235), .B(n12236), .ZN(n11956) );
  NAND2_X1 U12048 ( .A1(n12237), .A2(n12238), .ZN(n12235) );
  NAND2_X1 U12049 ( .A1(a_21_), .A2(n12234), .ZN(n11957) );
  NAND2_X1 U12050 ( .A1(n11965), .A2(n12239), .ZN(n12234) );
  NAND2_X1 U12051 ( .A1(n11964), .A2(n11966), .ZN(n12239) );
  NAND2_X1 U12052 ( .A1(n12240), .A2(n12241), .ZN(n11966) );
  NAND2_X1 U12053 ( .A1(a_22_), .A2(b_24_), .ZN(n12241) );
  INV_X1 U12054 ( .A(n12242), .ZN(n12240) );
  XNOR2_X1 U12055 ( .A(n12243), .B(n12244), .ZN(n11964) );
  XNOR2_X1 U12056 ( .A(n12245), .B(n12246), .ZN(n12243) );
  NAND2_X1 U12057 ( .A1(a_22_), .A2(n12242), .ZN(n11965) );
  NAND2_X1 U12058 ( .A1(n12247), .A2(n12248), .ZN(n12242) );
  NAND2_X1 U12059 ( .A1(n12249), .A2(a_23_), .ZN(n12248) );
  NOR2_X1 U12060 ( .A1(n12250), .A2(n10049), .ZN(n12249) );
  NOR2_X1 U12061 ( .A1(n11972), .A2(n11973), .ZN(n12250) );
  NAND2_X1 U12062 ( .A1(n11972), .A2(n11973), .ZN(n12247) );
  NAND2_X1 U12063 ( .A1(n12251), .A2(n12252), .ZN(n11973) );
  INV_X1 U12064 ( .A(n12253), .ZN(n12252) );
  NOR2_X1 U12065 ( .A1(n10022), .A2(n12254), .ZN(n12253) );
  NOR2_X1 U12066 ( .A1(n12033), .A2(n12031), .ZN(n12254) );
  INV_X1 U12067 ( .A(n12034), .ZN(n10022) );
  NOR2_X1 U12068 ( .A1(n10050), .A2(n10049), .ZN(n12034) );
  NAND2_X1 U12069 ( .A1(n12031), .A2(n12033), .ZN(n12251) );
  NAND2_X1 U12070 ( .A1(n12255), .A2(n12256), .ZN(n12033) );
  NAND2_X1 U12071 ( .A1(n11986), .A2(n12257), .ZN(n12256) );
  INV_X1 U12072 ( .A(n12258), .ZN(n12257) );
  NOR2_X1 U12073 ( .A1(n11983), .A2(n11985), .ZN(n12258) );
  NOR2_X1 U12074 ( .A1(n10048), .A2(n10049), .ZN(n11986) );
  NAND2_X1 U12075 ( .A1(n11985), .A2(n11983), .ZN(n12255) );
  XOR2_X1 U12076 ( .A(n12259), .B(n12260), .Z(n11983) );
  XNOR2_X1 U12077 ( .A(n12261), .B(n12262), .ZN(n12260) );
  NOR2_X1 U12078 ( .A1(n12263), .A2(n12264), .ZN(n11985) );
  INV_X1 U12079 ( .A(n12265), .ZN(n12264) );
  NAND2_X1 U12080 ( .A1(n11991), .A2(n12266), .ZN(n12265) );
  NAND2_X1 U12081 ( .A1(n11994), .A2(n11993), .ZN(n12266) );
  XOR2_X1 U12082 ( .A(n12267), .B(n12268), .Z(n11991) );
  NAND2_X1 U12083 ( .A1(n12269), .A2(n12270), .ZN(n12267) );
  NOR2_X1 U12084 ( .A1(n11993), .A2(n11994), .ZN(n12263) );
  NOR2_X1 U12085 ( .A1(n10047), .A2(n10049), .ZN(n11994) );
  NAND2_X1 U12086 ( .A1(n12000), .A2(n12271), .ZN(n11993) );
  NAND2_X1 U12087 ( .A1(n11999), .A2(n12001), .ZN(n12271) );
  NAND2_X1 U12088 ( .A1(n12272), .A2(n12273), .ZN(n12001) );
  NAND2_X1 U12089 ( .A1(a_27_), .A2(b_24_), .ZN(n12273) );
  INV_X1 U12090 ( .A(n12274), .ZN(n12272) );
  XNOR2_X1 U12091 ( .A(n12275), .B(n12276), .ZN(n11999) );
  XOR2_X1 U12092 ( .A(n12277), .B(n12278), .Z(n12276) );
  NAND2_X1 U12093 ( .A1(b_23_), .A2(a_28_), .ZN(n12278) );
  NAND2_X1 U12094 ( .A1(a_27_), .A2(n12274), .ZN(n12000) );
  NAND2_X1 U12095 ( .A1(n12279), .A2(n12280), .ZN(n12274) );
  NAND2_X1 U12096 ( .A1(n12281), .A2(a_28_), .ZN(n12280) );
  NOR2_X1 U12097 ( .A1(n12282), .A2(n10049), .ZN(n12281) );
  NOR2_X1 U12098 ( .A1(n12007), .A2(n12009), .ZN(n12282) );
  NAND2_X1 U12099 ( .A1(n12007), .A2(n12009), .ZN(n12279) );
  NAND2_X1 U12100 ( .A1(n12283), .A2(n12284), .ZN(n12009) );
  NAND2_X1 U12101 ( .A1(n12285), .A2(a_29_), .ZN(n12284) );
  NOR2_X1 U12102 ( .A1(n12286), .A2(n10049), .ZN(n12285) );
  NOR2_X1 U12103 ( .A1(n12287), .A2(n12029), .ZN(n12286) );
  NAND2_X1 U12104 ( .A1(n12287), .A2(n12029), .ZN(n12283) );
  NAND2_X1 U12105 ( .A1(n12288), .A2(n12289), .ZN(n12029) );
  NAND2_X1 U12106 ( .A1(b_22_), .A2(n12290), .ZN(n12289) );
  NAND2_X1 U12107 ( .A1(n10486), .A2(n12291), .ZN(n12290) );
  NAND2_X1 U12108 ( .A1(a_31_), .A2(n9302), .ZN(n12291) );
  NAND2_X1 U12109 ( .A1(b_23_), .A2(n12292), .ZN(n12288) );
  NAND2_X1 U12110 ( .A1(n10489), .A2(n12293), .ZN(n12292) );
  NAND2_X1 U12111 ( .A1(a_30_), .A2(n12294), .ZN(n12293) );
  INV_X1 U12112 ( .A(n12030), .ZN(n12287) );
  NAND2_X1 U12113 ( .A1(n12295), .A2(n9025), .ZN(n12030) );
  NOR2_X1 U12114 ( .A1(n10049), .A2(n9302), .ZN(n12295) );
  XOR2_X1 U12115 ( .A(n12296), .B(n12297), .Z(n12007) );
  NOR2_X1 U12116 ( .A1(n9121), .A2(n9302), .ZN(n12297) );
  XNOR2_X1 U12117 ( .A(n12298), .B(n12299), .ZN(n12296) );
  XOR2_X1 U12118 ( .A(n12300), .B(n12301), .Z(n12031) );
  XOR2_X1 U12119 ( .A(n12302), .B(n12303), .Z(n12301) );
  XNOR2_X1 U12120 ( .A(n12304), .B(n12305), .ZN(n11972) );
  XOR2_X1 U12121 ( .A(n12306), .B(n12307), .Z(n12305) );
  XOR2_X1 U12122 ( .A(n12308), .B(n12309), .Z(n12043) );
  XOR2_X1 U12123 ( .A(n12310), .B(n12311), .Z(n12308) );
  NOR2_X1 U12124 ( .A1(n9302), .A2(n10067), .ZN(n12311) );
  XNOR2_X1 U12125 ( .A(n12312), .B(n12313), .ZN(n12049) );
  NAND2_X1 U12126 ( .A1(n12314), .A2(n12315), .ZN(n12312) );
  XNOR2_X1 U12127 ( .A(n12316), .B(n12317), .ZN(n12057) );
  XNOR2_X1 U12128 ( .A(n12318), .B(n12319), .ZN(n12316) );
  XNOR2_X1 U12129 ( .A(n12320), .B(n12321), .ZN(n12060) );
  XNOR2_X1 U12130 ( .A(n12322), .B(n12323), .ZN(n12320) );
  XOR2_X1 U12131 ( .A(n12324), .B(n12325), .Z(n12065) );
  XNOR2_X1 U12132 ( .A(n12326), .B(n12327), .ZN(n12324) );
  NAND2_X1 U12133 ( .A1(a_7_), .A2(b_23_), .ZN(n12326) );
  XNOR2_X1 U12134 ( .A(n12328), .B(n12329), .ZN(n11861) );
  NAND2_X1 U12135 ( .A1(n12330), .A2(n12331), .ZN(n12328) );
  XOR2_X1 U12136 ( .A(n12332), .B(n12333), .Z(n12069) );
  XOR2_X1 U12137 ( .A(n12334), .B(n12335), .Z(n12332) );
  NOR2_X1 U12138 ( .A1(n9302), .A2(n10083), .ZN(n12335) );
  XNOR2_X1 U12139 ( .A(n12336), .B(n12337), .ZN(n12080) );
  NAND2_X1 U12140 ( .A1(n12338), .A2(n12339), .ZN(n12336) );
  XOR2_X1 U12141 ( .A(n12340), .B(n12341), .Z(n10303) );
  XNOR2_X1 U12142 ( .A(n12342), .B(n12343), .ZN(n12341) );
  INV_X1 U12143 ( .A(n12344), .ZN(n10159) );
  NOR2_X1 U12144 ( .A1(n12345), .A2(n10293), .ZN(n12344) );
  NAND2_X1 U12145 ( .A1(n12092), .A2(n12346), .ZN(n10293) );
  XNOR2_X1 U12146 ( .A(n12347), .B(n12093), .ZN(n12346) );
  XOR2_X1 U12147 ( .A(n12348), .B(n12349), .Z(n12093) );
  INV_X1 U12148 ( .A(n12094), .ZN(n12347) );
  NOR2_X1 U12149 ( .A1(n12350), .A2(n12351), .ZN(n12092) );
  INV_X1 U12150 ( .A(n12352), .ZN(n12351) );
  NAND2_X1 U12151 ( .A1(n12340), .A2(n12353), .ZN(n12352) );
  NAND2_X1 U12152 ( .A1(n12343), .A2(n12342), .ZN(n12353) );
  XOR2_X1 U12153 ( .A(n12354), .B(n12355), .Z(n12340) );
  NAND2_X1 U12154 ( .A1(n12356), .A2(n12357), .ZN(n12354) );
  NOR2_X1 U12155 ( .A1(n12342), .A2(n12343), .ZN(n12350) );
  NOR2_X1 U12156 ( .A1(n10093), .A2(n9302), .ZN(n12343) );
  NAND2_X1 U12157 ( .A1(n12358), .A2(n12359), .ZN(n12342) );
  NAND2_X1 U12158 ( .A1(n12360), .A2(a_1_), .ZN(n12359) );
  NOR2_X1 U12159 ( .A1(n12361), .A2(n9302), .ZN(n12360) );
  NOR2_X1 U12160 ( .A1(n12100), .A2(n12101), .ZN(n12361) );
  NAND2_X1 U12161 ( .A1(n12100), .A2(n12101), .ZN(n12358) );
  NAND2_X1 U12162 ( .A1(n12338), .A2(n12362), .ZN(n12101) );
  NAND2_X1 U12163 ( .A1(n12337), .A2(n12339), .ZN(n12362) );
  NAND2_X1 U12164 ( .A1(n12363), .A2(n12364), .ZN(n12339) );
  NAND2_X1 U12165 ( .A1(a_2_), .A2(b_23_), .ZN(n12363) );
  XNOR2_X1 U12166 ( .A(n12365), .B(n12366), .ZN(n12337) );
  NAND2_X1 U12167 ( .A1(n12367), .A2(n12368), .ZN(n12365) );
  NAND2_X1 U12168 ( .A1(n12369), .A2(a_2_), .ZN(n12338) );
  INV_X1 U12169 ( .A(n12364), .ZN(n12369) );
  NAND2_X1 U12170 ( .A1(n12370), .A2(n12371), .ZN(n12364) );
  NAND2_X1 U12171 ( .A1(n12111), .A2(n12372), .ZN(n12371) );
  NAND2_X1 U12172 ( .A1(n12114), .A2(n12113), .ZN(n12372) );
  XOR2_X1 U12173 ( .A(n12373), .B(n12374), .Z(n12111) );
  NAND2_X1 U12174 ( .A1(n12375), .A2(n12376), .ZN(n12373) );
  INV_X1 U12175 ( .A(n12377), .ZN(n12370) );
  NOR2_X1 U12176 ( .A1(n12113), .A2(n12114), .ZN(n12377) );
  NOR2_X1 U12177 ( .A1(n10086), .A2(n9302), .ZN(n12114) );
  NAND2_X1 U12178 ( .A1(n12378), .A2(n12379), .ZN(n12113) );
  NAND2_X1 U12179 ( .A1(n12380), .A2(a_4_), .ZN(n12379) );
  NOR2_X1 U12180 ( .A1(n12381), .A2(n9302), .ZN(n12380) );
  NOR2_X1 U12181 ( .A1(n12120), .A2(n12121), .ZN(n12381) );
  NAND2_X1 U12182 ( .A1(n12120), .A2(n12121), .ZN(n12378) );
  NAND2_X1 U12183 ( .A1(n12382), .A2(n12383), .ZN(n12121) );
  NAND2_X1 U12184 ( .A1(n12384), .A2(a_5_), .ZN(n12383) );
  NOR2_X1 U12185 ( .A1(n12385), .A2(n9302), .ZN(n12384) );
  NOR2_X1 U12186 ( .A1(n12333), .A2(n12334), .ZN(n12385) );
  NAND2_X1 U12187 ( .A1(n12333), .A2(n12334), .ZN(n12382) );
  NAND2_X1 U12188 ( .A1(n12330), .A2(n12386), .ZN(n12334) );
  NAND2_X1 U12189 ( .A1(n12329), .A2(n12331), .ZN(n12386) );
  NAND2_X1 U12190 ( .A1(n12387), .A2(n12388), .ZN(n12331) );
  NAND2_X1 U12191 ( .A1(a_6_), .A2(b_23_), .ZN(n12388) );
  INV_X1 U12192 ( .A(n12389), .ZN(n12387) );
  XNOR2_X1 U12193 ( .A(n12390), .B(n12391), .ZN(n12329) );
  NAND2_X1 U12194 ( .A1(n12392), .A2(n12393), .ZN(n12390) );
  NAND2_X1 U12195 ( .A1(a_6_), .A2(n12389), .ZN(n12330) );
  NAND2_X1 U12196 ( .A1(n12394), .A2(n12395), .ZN(n12389) );
  NAND2_X1 U12197 ( .A1(n12396), .A2(a_7_), .ZN(n12395) );
  NOR2_X1 U12198 ( .A1(n12397), .A2(n9302), .ZN(n12396) );
  NOR2_X1 U12199 ( .A1(n12325), .A2(n12327), .ZN(n12397) );
  NAND2_X1 U12200 ( .A1(n12325), .A2(n12327), .ZN(n12394) );
  NAND2_X1 U12201 ( .A1(n12398), .A2(n12399), .ZN(n12327) );
  NAND2_X1 U12202 ( .A1(n12142), .A2(n12400), .ZN(n12399) );
  INV_X1 U12203 ( .A(n12401), .ZN(n12400) );
  NOR2_X1 U12204 ( .A1(n12141), .A2(n12139), .ZN(n12401) );
  NOR2_X1 U12205 ( .A1(n10079), .A2(n9302), .ZN(n12142) );
  NAND2_X1 U12206 ( .A1(n12139), .A2(n12141), .ZN(n12398) );
  NAND2_X1 U12207 ( .A1(n12402), .A2(n12403), .ZN(n12141) );
  NAND2_X1 U12208 ( .A1(n12323), .A2(n12404), .ZN(n12403) );
  NAND2_X1 U12209 ( .A1(n12322), .A2(n12321), .ZN(n12404) );
  NOR2_X1 U12210 ( .A1(n10076), .A2(n9302), .ZN(n12323) );
  INV_X1 U12211 ( .A(n12405), .ZN(n12402) );
  NOR2_X1 U12212 ( .A1(n12321), .A2(n12322), .ZN(n12405) );
  NOR2_X1 U12213 ( .A1(n12406), .A2(n12407), .ZN(n12322) );
  INV_X1 U12214 ( .A(n12408), .ZN(n12407) );
  NAND2_X1 U12215 ( .A1(n12318), .A2(n12409), .ZN(n12408) );
  NAND2_X1 U12216 ( .A1(n12317), .A2(n12319), .ZN(n12409) );
  NAND2_X1 U12217 ( .A1(n12410), .A2(n12411), .ZN(n12318) );
  NAND2_X1 U12218 ( .A1(n12412), .A2(a_11_), .ZN(n12411) );
  NOR2_X1 U12219 ( .A1(n12413), .A2(n9302), .ZN(n12412) );
  NOR2_X1 U12220 ( .A1(n12156), .A2(n12157), .ZN(n12413) );
  NAND2_X1 U12221 ( .A1(n12156), .A2(n12157), .ZN(n12410) );
  NAND2_X1 U12222 ( .A1(n12314), .A2(n12414), .ZN(n12157) );
  NAND2_X1 U12223 ( .A1(n12313), .A2(n12315), .ZN(n12414) );
  NAND2_X1 U12224 ( .A1(n12415), .A2(n12416), .ZN(n12315) );
  NAND2_X1 U12225 ( .A1(a_12_), .A2(b_23_), .ZN(n12416) );
  INV_X1 U12226 ( .A(n12417), .ZN(n12415) );
  XNOR2_X1 U12227 ( .A(n12418), .B(n12419), .ZN(n12313) );
  NAND2_X1 U12228 ( .A1(n12420), .A2(n12421), .ZN(n12418) );
  NAND2_X1 U12229 ( .A1(a_12_), .A2(n12417), .ZN(n12314) );
  NAND2_X1 U12230 ( .A1(n12422), .A2(n12423), .ZN(n12417) );
  NAND2_X1 U12231 ( .A1(n12424), .A2(a_13_), .ZN(n12423) );
  NOR2_X1 U12232 ( .A1(n12425), .A2(n9302), .ZN(n12424) );
  NOR2_X1 U12233 ( .A1(n12309), .A2(n12310), .ZN(n12425) );
  NAND2_X1 U12234 ( .A1(n12309), .A2(n12310), .ZN(n12422) );
  NAND2_X1 U12235 ( .A1(n12172), .A2(n12426), .ZN(n12310) );
  NAND2_X1 U12236 ( .A1(n12171), .A2(n12173), .ZN(n12426) );
  NAND2_X1 U12237 ( .A1(n12427), .A2(n12428), .ZN(n12173) );
  NAND2_X1 U12238 ( .A1(a_14_), .A2(b_23_), .ZN(n12428) );
  INV_X1 U12239 ( .A(n12429), .ZN(n12427) );
  XNOR2_X1 U12240 ( .A(n12430), .B(n12431), .ZN(n12171) );
  XOR2_X1 U12241 ( .A(n12432), .B(n12433), .Z(n12431) );
  NAND2_X1 U12242 ( .A1(a_15_), .A2(b_22_), .ZN(n12433) );
  NAND2_X1 U12243 ( .A1(a_14_), .A2(n12429), .ZN(n12172) );
  NAND2_X1 U12244 ( .A1(n12434), .A2(n12435), .ZN(n12429) );
  NAND2_X1 U12245 ( .A1(n12436), .A2(a_15_), .ZN(n12435) );
  NOR2_X1 U12246 ( .A1(n12437), .A2(n9302), .ZN(n12436) );
  NOR2_X1 U12247 ( .A1(n12179), .A2(n12180), .ZN(n12437) );
  NAND2_X1 U12248 ( .A1(n12179), .A2(n12180), .ZN(n12434) );
  NAND2_X1 U12249 ( .A1(n12189), .A2(n12438), .ZN(n12180) );
  NAND2_X1 U12250 ( .A1(n12188), .A2(n12190), .ZN(n12438) );
  NAND2_X1 U12251 ( .A1(n12439), .A2(n12440), .ZN(n12190) );
  NAND2_X1 U12252 ( .A1(a_16_), .A2(b_23_), .ZN(n12440) );
  INV_X1 U12253 ( .A(n12441), .ZN(n12439) );
  XNOR2_X1 U12254 ( .A(n12442), .B(n12443), .ZN(n12188) );
  NAND2_X1 U12255 ( .A1(n12444), .A2(n12445), .ZN(n12442) );
  NAND2_X1 U12256 ( .A1(a_16_), .A2(n12441), .ZN(n12189) );
  NAND2_X1 U12257 ( .A1(n12197), .A2(n12446), .ZN(n12441) );
  NAND2_X1 U12258 ( .A1(n12196), .A2(n12198), .ZN(n12446) );
  NAND2_X1 U12259 ( .A1(n12447), .A2(n12448), .ZN(n12198) );
  NAND2_X1 U12260 ( .A1(a_17_), .A2(b_23_), .ZN(n12448) );
  INV_X1 U12261 ( .A(n12449), .ZN(n12447) );
  XNOR2_X1 U12262 ( .A(n12450), .B(n12451), .ZN(n12196) );
  NAND2_X1 U12263 ( .A1(n12452), .A2(n12453), .ZN(n12450) );
  NAND2_X1 U12264 ( .A1(a_17_), .A2(n12449), .ZN(n12197) );
  NAND2_X1 U12265 ( .A1(n12205), .A2(n12454), .ZN(n12449) );
  NAND2_X1 U12266 ( .A1(n12204), .A2(n12206), .ZN(n12454) );
  NAND2_X1 U12267 ( .A1(n12455), .A2(n12456), .ZN(n12206) );
  NAND2_X1 U12268 ( .A1(a_18_), .A2(b_23_), .ZN(n12456) );
  INV_X1 U12269 ( .A(n12457), .ZN(n12455) );
  XOR2_X1 U12270 ( .A(n12458), .B(n12459), .Z(n12204) );
  XOR2_X1 U12271 ( .A(n12460), .B(n12461), .Z(n12458) );
  NOR2_X1 U12272 ( .A1(n12294), .A2(n9415), .ZN(n12461) );
  NAND2_X1 U12273 ( .A1(a_18_), .A2(n12457), .ZN(n12205) );
  NAND2_X1 U12274 ( .A1(n12462), .A2(n12463), .ZN(n12457) );
  NAND2_X1 U12275 ( .A1(n12464), .A2(a_19_), .ZN(n12463) );
  NOR2_X1 U12276 ( .A1(n12465), .A2(n9302), .ZN(n12464) );
  NOR2_X1 U12277 ( .A1(n12211), .A2(n12213), .ZN(n12465) );
  NAND2_X1 U12278 ( .A1(n12211), .A2(n12213), .ZN(n12462) );
  NAND2_X1 U12279 ( .A1(n12221), .A2(n12466), .ZN(n12213) );
  NAND2_X1 U12280 ( .A1(n12220), .A2(n12222), .ZN(n12466) );
  NAND2_X1 U12281 ( .A1(n12467), .A2(n12468), .ZN(n12222) );
  NAND2_X1 U12282 ( .A1(a_20_), .A2(b_23_), .ZN(n12468) );
  INV_X1 U12283 ( .A(n12469), .ZN(n12467) );
  XNOR2_X1 U12284 ( .A(n12470), .B(n12471), .ZN(n12220) );
  NAND2_X1 U12285 ( .A1(n12472), .A2(n12473), .ZN(n12470) );
  NAND2_X1 U12286 ( .A1(a_20_), .A2(n12469), .ZN(n12221) );
  NAND2_X1 U12287 ( .A1(n12228), .A2(n12474), .ZN(n12469) );
  NAND2_X1 U12288 ( .A1(n12227), .A2(n12229), .ZN(n12474) );
  NAND2_X1 U12289 ( .A1(n12475), .A2(n12476), .ZN(n12229) );
  NAND2_X1 U12290 ( .A1(a_21_), .A2(b_23_), .ZN(n12476) );
  INV_X1 U12291 ( .A(n12477), .ZN(n12475) );
  XOR2_X1 U12292 ( .A(n12478), .B(n12479), .Z(n12227) );
  XNOR2_X1 U12293 ( .A(n12480), .B(n10016), .ZN(n12479) );
  NAND2_X1 U12294 ( .A1(a_21_), .A2(n12477), .ZN(n12228) );
  NAND2_X1 U12295 ( .A1(n12237), .A2(n12481), .ZN(n12477) );
  NAND2_X1 U12296 ( .A1(n12236), .A2(n12238), .ZN(n12481) );
  NAND2_X1 U12297 ( .A1(n12482), .A2(n12483), .ZN(n12238) );
  NAND2_X1 U12298 ( .A1(a_22_), .A2(b_23_), .ZN(n12482) );
  XOR2_X1 U12299 ( .A(n12484), .B(n12485), .Z(n12236) );
  XOR2_X1 U12300 ( .A(n12486), .B(n12487), .Z(n12484) );
  NOR2_X1 U12301 ( .A1(n10051), .A2(n12294), .ZN(n12487) );
  INV_X1 U12302 ( .A(n12488), .ZN(n12237) );
  NOR2_X1 U12303 ( .A1(n12483), .A2(n9330), .ZN(n12488) );
  NAND2_X1 U12304 ( .A1(n12489), .A2(n12490), .ZN(n12483) );
  NAND2_X1 U12305 ( .A1(n12244), .A2(n12491), .ZN(n12490) );
  NAND2_X1 U12306 ( .A1(n12246), .A2(n12492), .ZN(n12491) );
  INV_X1 U12307 ( .A(n12245), .ZN(n12492) );
  XOR2_X1 U12308 ( .A(n12493), .B(n12494), .Z(n12244) );
  XNOR2_X1 U12309 ( .A(n12495), .B(n12496), .ZN(n12494) );
  NAND2_X1 U12310 ( .A1(n12245), .A2(n10019), .ZN(n12489) );
  INV_X1 U12311 ( .A(n12246), .ZN(n10019) );
  NOR2_X1 U12312 ( .A1(n9302), .A2(n10051), .ZN(n12246) );
  NOR2_X1 U12313 ( .A1(n12497), .A2(n12498), .ZN(n12245) );
  NOR2_X1 U12314 ( .A1(n12307), .A2(n12499), .ZN(n12498) );
  NOR2_X1 U12315 ( .A1(n12306), .A2(n12304), .ZN(n12499) );
  NAND2_X1 U12316 ( .A1(b_23_), .A2(a_24_), .ZN(n12307) );
  INV_X1 U12317 ( .A(n12500), .ZN(n12497) );
  NAND2_X1 U12318 ( .A1(n12304), .A2(n12306), .ZN(n12500) );
  NAND2_X1 U12319 ( .A1(n12501), .A2(n12502), .ZN(n12306) );
  NAND2_X1 U12320 ( .A1(n12303), .A2(n12503), .ZN(n12502) );
  INV_X1 U12321 ( .A(n12504), .ZN(n12503) );
  NOR2_X1 U12322 ( .A1(n12300), .A2(n12302), .ZN(n12504) );
  NOR2_X1 U12323 ( .A1(n9302), .A2(n10048), .ZN(n12303) );
  NAND2_X1 U12324 ( .A1(n12302), .A2(n12300), .ZN(n12501) );
  XOR2_X1 U12325 ( .A(n12505), .B(n12506), .Z(n12300) );
  XNOR2_X1 U12326 ( .A(n12507), .B(n12508), .ZN(n12506) );
  NOR2_X1 U12327 ( .A1(n12509), .A2(n12510), .ZN(n12302) );
  INV_X1 U12328 ( .A(n12511), .ZN(n12510) );
  NAND2_X1 U12329 ( .A1(n12259), .A2(n12512), .ZN(n12511) );
  NAND2_X1 U12330 ( .A1(n12262), .A2(n12261), .ZN(n12512) );
  XOR2_X1 U12331 ( .A(n12513), .B(n12514), .Z(n12259) );
  NAND2_X1 U12332 ( .A1(n12515), .A2(n12516), .ZN(n12513) );
  NOR2_X1 U12333 ( .A1(n12261), .A2(n12262), .ZN(n12509) );
  NOR2_X1 U12334 ( .A1(n9302), .A2(n10047), .ZN(n12262) );
  NAND2_X1 U12335 ( .A1(n12269), .A2(n12517), .ZN(n12261) );
  NAND2_X1 U12336 ( .A1(n12268), .A2(n12270), .ZN(n12517) );
  NAND2_X1 U12337 ( .A1(n12518), .A2(n12519), .ZN(n12270) );
  NAND2_X1 U12338 ( .A1(b_23_), .A2(a_27_), .ZN(n12519) );
  INV_X1 U12339 ( .A(n12520), .ZN(n12518) );
  XNOR2_X1 U12340 ( .A(n12521), .B(n12522), .ZN(n12268) );
  XOR2_X1 U12341 ( .A(n12523), .B(n12524), .Z(n12522) );
  NAND2_X1 U12342 ( .A1(b_22_), .A2(a_28_), .ZN(n12524) );
  NAND2_X1 U12343 ( .A1(a_27_), .A2(n12520), .ZN(n12269) );
  NAND2_X1 U12344 ( .A1(n12525), .A2(n12526), .ZN(n12520) );
  NAND2_X1 U12345 ( .A1(n12527), .A2(b_23_), .ZN(n12526) );
  NOR2_X1 U12346 ( .A1(n12528), .A2(n9136), .ZN(n12527) );
  NOR2_X1 U12347 ( .A1(n12275), .A2(n12277), .ZN(n12528) );
  NAND2_X1 U12348 ( .A1(n12275), .A2(n12277), .ZN(n12525) );
  NAND2_X1 U12349 ( .A1(n12529), .A2(n12530), .ZN(n12277) );
  NAND2_X1 U12350 ( .A1(n12531), .A2(b_23_), .ZN(n12530) );
  NOR2_X1 U12351 ( .A1(n12532), .A2(n9121), .ZN(n12531) );
  NOR2_X1 U12352 ( .A1(n12533), .A2(n12298), .ZN(n12532) );
  NAND2_X1 U12353 ( .A1(n12533), .A2(n12298), .ZN(n12529) );
  NAND2_X1 U12354 ( .A1(n12534), .A2(n12535), .ZN(n12298) );
  NAND2_X1 U12355 ( .A1(b_21_), .A2(n12536), .ZN(n12535) );
  NAND2_X1 U12356 ( .A1(n10486), .A2(n12537), .ZN(n12536) );
  NAND2_X1 U12357 ( .A1(a_31_), .A2(n12294), .ZN(n12537) );
  NAND2_X1 U12358 ( .A1(b_22_), .A2(n12538), .ZN(n12534) );
  NAND2_X1 U12359 ( .A1(n10489), .A2(n12539), .ZN(n12538) );
  NAND2_X1 U12360 ( .A1(a_30_), .A2(n10052), .ZN(n12539) );
  INV_X1 U12361 ( .A(n12299), .ZN(n12533) );
  NAND2_X1 U12362 ( .A1(n12540), .A2(n9025), .ZN(n12299) );
  NOR2_X1 U12363 ( .A1(n9302), .A2(n12294), .ZN(n12540) );
  XOR2_X1 U12364 ( .A(n12541), .B(n12542), .Z(n12275) );
  NOR2_X1 U12365 ( .A1(n9121), .A2(n12294), .ZN(n12542) );
  XNOR2_X1 U12366 ( .A(n12543), .B(n12544), .ZN(n12541) );
  XNOR2_X1 U12367 ( .A(n12545), .B(n12546), .ZN(n12304) );
  XNOR2_X1 U12368 ( .A(n12547), .B(n12548), .ZN(n12546) );
  XNOR2_X1 U12369 ( .A(n12549), .B(n12550), .ZN(n12211) );
  NAND2_X1 U12370 ( .A1(n12551), .A2(n12552), .ZN(n12549) );
  XNOR2_X1 U12371 ( .A(n12553), .B(n12554), .ZN(n12179) );
  NAND2_X1 U12372 ( .A1(n12555), .A2(n12556), .ZN(n12553) );
  XOR2_X1 U12373 ( .A(n12557), .B(n12558), .Z(n12309) );
  XNOR2_X1 U12374 ( .A(n12559), .B(n12560), .ZN(n12558) );
  XOR2_X1 U12375 ( .A(n12561), .B(n12562), .Z(n12156) );
  XOR2_X1 U12376 ( .A(n12563), .B(n12564), .Z(n12561) );
  NOR2_X1 U12377 ( .A1(n12294), .A2(n10070), .ZN(n12564) );
  NOR2_X1 U12378 ( .A1(n12319), .A2(n12317), .ZN(n12406) );
  XOR2_X1 U12379 ( .A(n12565), .B(n12566), .Z(n12317) );
  NAND2_X1 U12380 ( .A1(n12567), .A2(n12568), .ZN(n12565) );
  NAND2_X1 U12381 ( .A1(a_10_), .A2(b_23_), .ZN(n12319) );
  XOR2_X1 U12382 ( .A(n12569), .B(n12570), .Z(n12321) );
  XOR2_X1 U12383 ( .A(n12571), .B(n12572), .Z(n12569) );
  XNOR2_X1 U12384 ( .A(n12573), .B(n12574), .ZN(n12139) );
  NAND2_X1 U12385 ( .A1(n12575), .A2(n12576), .ZN(n12573) );
  XNOR2_X1 U12386 ( .A(n12577), .B(n12578), .ZN(n12325) );
  NAND2_X1 U12387 ( .A1(n12579), .A2(n12580), .ZN(n12577) );
  XOR2_X1 U12388 ( .A(n12581), .B(n12582), .Z(n12333) );
  XOR2_X1 U12389 ( .A(n12583), .B(n12584), .Z(n12581) );
  NOR2_X1 U12390 ( .A1(n12294), .A2(n10081), .ZN(n12584) );
  XNOR2_X1 U12391 ( .A(n12585), .B(n12586), .ZN(n12120) );
  NAND2_X1 U12392 ( .A1(n12587), .A2(n12588), .ZN(n12585) );
  XNOR2_X1 U12393 ( .A(n12589), .B(n12590), .ZN(n12100) );
  NAND2_X1 U12394 ( .A1(n12591), .A2(n12592), .ZN(n12589) );
  NAND2_X1 U12395 ( .A1(n12593), .A2(n12594), .ZN(n12345) );
  INV_X1 U12396 ( .A(n12595), .ZN(n12594) );
  NOR2_X1 U12397 ( .A1(n10295), .A2(n10294), .ZN(n12595) );
  NAND2_X1 U12398 ( .A1(n12596), .A2(n12593), .ZN(n10165) );
  INV_X1 U12399 ( .A(n12597), .ZN(n10164) );
  NOR2_X1 U12400 ( .A1(n12593), .A2(n12596), .ZN(n12597) );
  XNOR2_X1 U12401 ( .A(n12598), .B(n12599), .ZN(n12596) );
  NAND2_X1 U12402 ( .A1(n10295), .A2(n10294), .ZN(n12593) );
  NAND2_X1 U12403 ( .A1(n12600), .A2(n12601), .ZN(n10294) );
  NAND2_X1 U12404 ( .A1(n12349), .A2(n12602), .ZN(n12601) );
  INV_X1 U12405 ( .A(n12603), .ZN(n12602) );
  NOR2_X1 U12406 ( .A1(n12348), .A2(n12094), .ZN(n12603) );
  NOR2_X1 U12407 ( .A1(n10093), .A2(n12294), .ZN(n12349) );
  NAND2_X1 U12408 ( .A1(n12094), .A2(n12348), .ZN(n12600) );
  NAND2_X1 U12409 ( .A1(n12356), .A2(n12604), .ZN(n12348) );
  NAND2_X1 U12410 ( .A1(n12355), .A2(n12357), .ZN(n12604) );
  NAND2_X1 U12411 ( .A1(n12605), .A2(n12606), .ZN(n12357) );
  NAND2_X1 U12412 ( .A1(a_1_), .A2(b_22_), .ZN(n12606) );
  INV_X1 U12413 ( .A(n12607), .ZN(n12605) );
  XOR2_X1 U12414 ( .A(n12608), .B(n12609), .Z(n12355) );
  XNOR2_X1 U12415 ( .A(n12610), .B(n12611), .ZN(n12609) );
  NAND2_X1 U12416 ( .A1(a_1_), .A2(n12607), .ZN(n12356) );
  NAND2_X1 U12417 ( .A1(n12591), .A2(n12612), .ZN(n12607) );
  NAND2_X1 U12418 ( .A1(n12590), .A2(n12592), .ZN(n12612) );
  NAND2_X1 U12419 ( .A1(n12613), .A2(n12614), .ZN(n12592) );
  NAND2_X1 U12420 ( .A1(a_2_), .A2(b_22_), .ZN(n12614) );
  INV_X1 U12421 ( .A(n12615), .ZN(n12613) );
  XNOR2_X1 U12422 ( .A(n12616), .B(n12617), .ZN(n12590) );
  NAND2_X1 U12423 ( .A1(n12618), .A2(n12619), .ZN(n12616) );
  NAND2_X1 U12424 ( .A1(a_2_), .A2(n12615), .ZN(n12591) );
  NAND2_X1 U12425 ( .A1(n12367), .A2(n12620), .ZN(n12615) );
  NAND2_X1 U12426 ( .A1(n12366), .A2(n12368), .ZN(n12620) );
  NAND2_X1 U12427 ( .A1(n12621), .A2(n12622), .ZN(n12368) );
  NAND2_X1 U12428 ( .A1(a_3_), .A2(b_22_), .ZN(n12622) );
  INV_X1 U12429 ( .A(n12623), .ZN(n12621) );
  XOR2_X1 U12430 ( .A(n12624), .B(n12625), .Z(n12366) );
  XNOR2_X1 U12431 ( .A(n12626), .B(n12627), .ZN(n12625) );
  NAND2_X1 U12432 ( .A1(a_3_), .A2(n12623), .ZN(n12367) );
  NAND2_X1 U12433 ( .A1(n12375), .A2(n12628), .ZN(n12623) );
  NAND2_X1 U12434 ( .A1(n12374), .A2(n12376), .ZN(n12628) );
  NAND2_X1 U12435 ( .A1(n12629), .A2(n12630), .ZN(n12376) );
  NAND2_X1 U12436 ( .A1(a_4_), .A2(b_22_), .ZN(n12630) );
  INV_X1 U12437 ( .A(n12631), .ZN(n12629) );
  XNOR2_X1 U12438 ( .A(n12632), .B(n12633), .ZN(n12374) );
  XNOR2_X1 U12439 ( .A(n12634), .B(n12635), .ZN(n12632) );
  NOR2_X1 U12440 ( .A1(n10052), .A2(n10083), .ZN(n12635) );
  NAND2_X1 U12441 ( .A1(a_4_), .A2(n12631), .ZN(n12375) );
  NAND2_X1 U12442 ( .A1(n12587), .A2(n12636), .ZN(n12631) );
  NAND2_X1 U12443 ( .A1(n12586), .A2(n12588), .ZN(n12636) );
  NAND2_X1 U12444 ( .A1(n12637), .A2(n12638), .ZN(n12588) );
  NAND2_X1 U12445 ( .A1(a_5_), .A2(b_22_), .ZN(n12638) );
  INV_X1 U12446 ( .A(n12639), .ZN(n12637) );
  XOR2_X1 U12447 ( .A(n12640), .B(n12641), .Z(n12586) );
  XNOR2_X1 U12448 ( .A(n12642), .B(n12643), .ZN(n12641) );
  NAND2_X1 U12449 ( .A1(a_5_), .A2(n12639), .ZN(n12587) );
  NAND2_X1 U12450 ( .A1(n12644), .A2(n12645), .ZN(n12639) );
  NAND2_X1 U12451 ( .A1(n12646), .A2(a_6_), .ZN(n12645) );
  NOR2_X1 U12452 ( .A1(n12647), .A2(n12294), .ZN(n12646) );
  NOR2_X1 U12453 ( .A1(n12582), .A2(n12583), .ZN(n12647) );
  NAND2_X1 U12454 ( .A1(n12582), .A2(n12583), .ZN(n12644) );
  NAND2_X1 U12455 ( .A1(n12392), .A2(n12648), .ZN(n12583) );
  NAND2_X1 U12456 ( .A1(n12391), .A2(n12393), .ZN(n12648) );
  NAND2_X1 U12457 ( .A1(n12649), .A2(n12650), .ZN(n12393) );
  NAND2_X1 U12458 ( .A1(a_7_), .A2(b_22_), .ZN(n12650) );
  INV_X1 U12459 ( .A(n12651), .ZN(n12649) );
  XNOR2_X1 U12460 ( .A(n12652), .B(n12653), .ZN(n12391) );
  XOR2_X1 U12461 ( .A(n12654), .B(n12655), .Z(n12652) );
  NAND2_X1 U12462 ( .A1(a_7_), .A2(n12651), .ZN(n12392) );
  NAND2_X1 U12463 ( .A1(n12579), .A2(n12656), .ZN(n12651) );
  NAND2_X1 U12464 ( .A1(n12578), .A2(n12580), .ZN(n12656) );
  NAND2_X1 U12465 ( .A1(n12657), .A2(n12658), .ZN(n12580) );
  NAND2_X1 U12466 ( .A1(a_8_), .A2(b_22_), .ZN(n12658) );
  INV_X1 U12467 ( .A(n12659), .ZN(n12657) );
  XNOR2_X1 U12468 ( .A(n12660), .B(n12661), .ZN(n12578) );
  NAND2_X1 U12469 ( .A1(n12662), .A2(n12663), .ZN(n12660) );
  NAND2_X1 U12470 ( .A1(a_8_), .A2(n12659), .ZN(n12579) );
  NAND2_X1 U12471 ( .A1(n12575), .A2(n12664), .ZN(n12659) );
  NAND2_X1 U12472 ( .A1(n12574), .A2(n12576), .ZN(n12664) );
  NAND2_X1 U12473 ( .A1(n12665), .A2(n12666), .ZN(n12576) );
  NAND2_X1 U12474 ( .A1(a_9_), .A2(b_22_), .ZN(n12665) );
  XNOR2_X1 U12475 ( .A(n12667), .B(n12668), .ZN(n12574) );
  XOR2_X1 U12476 ( .A(n12669), .B(n12670), .Z(n12668) );
  NAND2_X1 U12477 ( .A1(a_10_), .A2(b_21_), .ZN(n12670) );
  NAND2_X1 U12478 ( .A1(n12671), .A2(a_9_), .ZN(n12575) );
  INV_X1 U12479 ( .A(n12666), .ZN(n12671) );
  NAND2_X1 U12480 ( .A1(n12672), .A2(n12673), .ZN(n12666) );
  NAND2_X1 U12481 ( .A1(n12570), .A2(n12674), .ZN(n12673) );
  NAND2_X1 U12482 ( .A1(n12572), .A2(n12571), .ZN(n12674) );
  XNOR2_X1 U12483 ( .A(n12675), .B(n12676), .ZN(n12570) );
  XOR2_X1 U12484 ( .A(n12677), .B(n12678), .Z(n12675) );
  NOR2_X1 U12485 ( .A1(n10052), .A2(n9649), .ZN(n12678) );
  INV_X1 U12486 ( .A(n12679), .ZN(n12672) );
  NOR2_X1 U12487 ( .A1(n12571), .A2(n12572), .ZN(n12679) );
  NOR2_X1 U12488 ( .A1(n10073), .A2(n12294), .ZN(n12572) );
  NAND2_X1 U12489 ( .A1(n12567), .A2(n12680), .ZN(n12571) );
  NAND2_X1 U12490 ( .A1(n12566), .A2(n12568), .ZN(n12680) );
  NAND2_X1 U12491 ( .A1(n12681), .A2(n12682), .ZN(n12568) );
  NAND2_X1 U12492 ( .A1(a_11_), .A2(b_22_), .ZN(n12682) );
  INV_X1 U12493 ( .A(n12683), .ZN(n12681) );
  XNOR2_X1 U12494 ( .A(n12684), .B(n12685), .ZN(n12566) );
  NAND2_X1 U12495 ( .A1(n12686), .A2(n12687), .ZN(n12684) );
  NAND2_X1 U12496 ( .A1(a_11_), .A2(n12683), .ZN(n12567) );
  NAND2_X1 U12497 ( .A1(n12688), .A2(n12689), .ZN(n12683) );
  NAND2_X1 U12498 ( .A1(n12690), .A2(a_12_), .ZN(n12689) );
  NOR2_X1 U12499 ( .A1(n12691), .A2(n12294), .ZN(n12690) );
  NOR2_X1 U12500 ( .A1(n12562), .A2(n12563), .ZN(n12691) );
  NAND2_X1 U12501 ( .A1(n12562), .A2(n12563), .ZN(n12688) );
  NAND2_X1 U12502 ( .A1(n12420), .A2(n12692), .ZN(n12563) );
  NAND2_X1 U12503 ( .A1(n12419), .A2(n12421), .ZN(n12692) );
  NAND2_X1 U12504 ( .A1(n12693), .A2(n12694), .ZN(n12421) );
  NAND2_X1 U12505 ( .A1(a_13_), .A2(b_22_), .ZN(n12693) );
  XNOR2_X1 U12506 ( .A(n12695), .B(n12696), .ZN(n12419) );
  XOR2_X1 U12507 ( .A(n12697), .B(n12698), .Z(n12696) );
  NAND2_X1 U12508 ( .A1(a_14_), .A2(b_21_), .ZN(n12698) );
  NAND2_X1 U12509 ( .A1(n12699), .A2(a_13_), .ZN(n12420) );
  INV_X1 U12510 ( .A(n12694), .ZN(n12699) );
  NAND2_X1 U12511 ( .A1(n12700), .A2(n12701), .ZN(n12694) );
  NAND2_X1 U12512 ( .A1(n12557), .A2(n12702), .ZN(n12701) );
  NAND2_X1 U12513 ( .A1(n12560), .A2(n12559), .ZN(n12702) );
  XNOR2_X1 U12514 ( .A(n12703), .B(n12704), .ZN(n12557) );
  XOR2_X1 U12515 ( .A(n12705), .B(n12706), .Z(n12703) );
  NOR2_X1 U12516 ( .A1(n10052), .A2(n9534), .ZN(n12706) );
  INV_X1 U12517 ( .A(n12707), .ZN(n12700) );
  NOR2_X1 U12518 ( .A1(n12559), .A2(n12560), .ZN(n12707) );
  NOR2_X1 U12519 ( .A1(n10065), .A2(n12294), .ZN(n12560) );
  NAND2_X1 U12520 ( .A1(n12708), .A2(n12709), .ZN(n12559) );
  NAND2_X1 U12521 ( .A1(n12710), .A2(a_15_), .ZN(n12709) );
  NOR2_X1 U12522 ( .A1(n12711), .A2(n12294), .ZN(n12710) );
  NOR2_X1 U12523 ( .A1(n12430), .A2(n12432), .ZN(n12711) );
  NAND2_X1 U12524 ( .A1(n12430), .A2(n12432), .ZN(n12708) );
  NAND2_X1 U12525 ( .A1(n12555), .A2(n12712), .ZN(n12432) );
  NAND2_X1 U12526 ( .A1(n12554), .A2(n12556), .ZN(n12712) );
  NAND2_X1 U12527 ( .A1(n12713), .A2(n12714), .ZN(n12556) );
  NAND2_X1 U12528 ( .A1(a_16_), .A2(b_22_), .ZN(n12714) );
  INV_X1 U12529 ( .A(n12715), .ZN(n12713) );
  XNOR2_X1 U12530 ( .A(n12716), .B(n12717), .ZN(n12554) );
  NAND2_X1 U12531 ( .A1(n12718), .A2(n12719), .ZN(n12716) );
  NAND2_X1 U12532 ( .A1(a_16_), .A2(n12715), .ZN(n12555) );
  NAND2_X1 U12533 ( .A1(n12444), .A2(n12720), .ZN(n12715) );
  NAND2_X1 U12534 ( .A1(n12443), .A2(n12445), .ZN(n12720) );
  NAND2_X1 U12535 ( .A1(n12721), .A2(n12722), .ZN(n12445) );
  NAND2_X1 U12536 ( .A1(a_17_), .A2(b_22_), .ZN(n12722) );
  INV_X1 U12537 ( .A(n12723), .ZN(n12721) );
  XNOR2_X1 U12538 ( .A(n12724), .B(n12725), .ZN(n12443) );
  NAND2_X1 U12539 ( .A1(n12726), .A2(n12727), .ZN(n12724) );
  NAND2_X1 U12540 ( .A1(a_17_), .A2(n12723), .ZN(n12444) );
  NAND2_X1 U12541 ( .A1(n12452), .A2(n12728), .ZN(n12723) );
  NAND2_X1 U12542 ( .A1(n12451), .A2(n12453), .ZN(n12728) );
  NAND2_X1 U12543 ( .A1(n12729), .A2(n12730), .ZN(n12453) );
  NAND2_X1 U12544 ( .A1(a_18_), .A2(b_22_), .ZN(n12730) );
  INV_X1 U12545 ( .A(n12731), .ZN(n12729) );
  XOR2_X1 U12546 ( .A(n12732), .B(n12733), .Z(n12451) );
  XNOR2_X1 U12547 ( .A(n12734), .B(n12735), .ZN(n12733) );
  NAND2_X1 U12548 ( .A1(a_19_), .A2(b_21_), .ZN(n12735) );
  NAND2_X1 U12549 ( .A1(a_18_), .A2(n12731), .ZN(n12452) );
  NAND2_X1 U12550 ( .A1(n12736), .A2(n12737), .ZN(n12731) );
  NAND2_X1 U12551 ( .A1(n12738), .A2(a_19_), .ZN(n12737) );
  NOR2_X1 U12552 ( .A1(n12739), .A2(n12294), .ZN(n12738) );
  NOR2_X1 U12553 ( .A1(n12459), .A2(n12460), .ZN(n12739) );
  NAND2_X1 U12554 ( .A1(n12459), .A2(n12460), .ZN(n12736) );
  NAND2_X1 U12555 ( .A1(n12551), .A2(n12740), .ZN(n12460) );
  NAND2_X1 U12556 ( .A1(n12550), .A2(n12552), .ZN(n12740) );
  NAND2_X1 U12557 ( .A1(n12741), .A2(n12742), .ZN(n12552) );
  NAND2_X1 U12558 ( .A1(a_20_), .A2(b_22_), .ZN(n12742) );
  INV_X1 U12559 ( .A(n12743), .ZN(n12741) );
  XNOR2_X1 U12560 ( .A(n12744), .B(n12745), .ZN(n12550) );
  XNOR2_X1 U12561 ( .A(n12746), .B(n12747), .ZN(n12744) );
  NAND2_X1 U12562 ( .A1(a_20_), .A2(n12743), .ZN(n12551) );
  NAND2_X1 U12563 ( .A1(n12472), .A2(n12748), .ZN(n12743) );
  NAND2_X1 U12564 ( .A1(n12471), .A2(n12473), .ZN(n12748) );
  NAND2_X1 U12565 ( .A1(n12749), .A2(n12750), .ZN(n12473) );
  NAND2_X1 U12566 ( .A1(a_21_), .A2(b_22_), .ZN(n12749) );
  XNOR2_X1 U12567 ( .A(n12751), .B(n12752), .ZN(n12471) );
  NAND2_X1 U12568 ( .A1(n12753), .A2(n12754), .ZN(n12751) );
  NAND2_X1 U12569 ( .A1(n12755), .A2(a_21_), .ZN(n12472) );
  INV_X1 U12570 ( .A(n12750), .ZN(n12755) );
  NAND2_X1 U12571 ( .A1(n12756), .A2(n12757), .ZN(n12750) );
  NAND2_X1 U12572 ( .A1(n12478), .A2(n12758), .ZN(n12757) );
  NAND2_X1 U12573 ( .A1(n10016), .A2(n12480), .ZN(n12758) );
  XNOR2_X1 U12574 ( .A(n12759), .B(n12760), .ZN(n12478) );
  XOR2_X1 U12575 ( .A(n12761), .B(n12762), .Z(n12759) );
  NOR2_X1 U12576 ( .A1(n10051), .A2(n10052), .ZN(n12762) );
  INV_X1 U12577 ( .A(n12763), .ZN(n12756) );
  NOR2_X1 U12578 ( .A1(n12480), .A2(n10016), .ZN(n12763) );
  NOR2_X1 U12579 ( .A1(n12294), .A2(n9330), .ZN(n10016) );
  NAND2_X1 U12580 ( .A1(n12764), .A2(n12765), .ZN(n12480) );
  NAND2_X1 U12581 ( .A1(n12766), .A2(b_22_), .ZN(n12765) );
  NOR2_X1 U12582 ( .A1(n12767), .A2(n10051), .ZN(n12766) );
  NOR2_X1 U12583 ( .A1(n12485), .A2(n12486), .ZN(n12767) );
  NAND2_X1 U12584 ( .A1(n12485), .A2(n12486), .ZN(n12764) );
  NAND2_X1 U12585 ( .A1(n12768), .A2(n12769), .ZN(n12486) );
  INV_X1 U12586 ( .A(n12770), .ZN(n12769) );
  NOR2_X1 U12587 ( .A1(n12771), .A2(n12772), .ZN(n12770) );
  NOR2_X1 U12588 ( .A1(n12495), .A2(n12493), .ZN(n12772) );
  INV_X1 U12589 ( .A(n12496), .ZN(n12771) );
  NOR2_X1 U12590 ( .A1(n12294), .A2(n10050), .ZN(n12496) );
  NAND2_X1 U12591 ( .A1(n12493), .A2(n12495), .ZN(n12768) );
  NAND2_X1 U12592 ( .A1(n12773), .A2(n12774), .ZN(n12495) );
  NAND2_X1 U12593 ( .A1(n12548), .A2(n12775), .ZN(n12774) );
  NAND2_X1 U12594 ( .A1(n12545), .A2(n12547), .ZN(n12775) );
  NOR2_X1 U12595 ( .A1(n12294), .A2(n10048), .ZN(n12548) );
  INV_X1 U12596 ( .A(n12776), .ZN(n12773) );
  NOR2_X1 U12597 ( .A1(n12547), .A2(n12545), .ZN(n12776) );
  XNOR2_X1 U12598 ( .A(n12777), .B(n12778), .ZN(n12545) );
  XNOR2_X1 U12599 ( .A(n12779), .B(n12780), .ZN(n12778) );
  NAND2_X1 U12600 ( .A1(n12781), .A2(n12782), .ZN(n12547) );
  NAND2_X1 U12601 ( .A1(n12505), .A2(n12783), .ZN(n12782) );
  NAND2_X1 U12602 ( .A1(n12508), .A2(n12507), .ZN(n12783) );
  XOR2_X1 U12603 ( .A(n12784), .B(n12785), .Z(n12505) );
  NAND2_X1 U12604 ( .A1(n12786), .A2(n12787), .ZN(n12784) );
  INV_X1 U12605 ( .A(n12788), .ZN(n12781) );
  NOR2_X1 U12606 ( .A1(n12507), .A2(n12508), .ZN(n12788) );
  NOR2_X1 U12607 ( .A1(n12294), .A2(n10047), .ZN(n12508) );
  NAND2_X1 U12608 ( .A1(n12515), .A2(n12789), .ZN(n12507) );
  NAND2_X1 U12609 ( .A1(n12514), .A2(n12516), .ZN(n12789) );
  NAND2_X1 U12610 ( .A1(n12790), .A2(n12791), .ZN(n12516) );
  NAND2_X1 U12611 ( .A1(b_22_), .A2(a_27_), .ZN(n12791) );
  INV_X1 U12612 ( .A(n12792), .ZN(n12790) );
  XNOR2_X1 U12613 ( .A(n12793), .B(n12794), .ZN(n12514) );
  XOR2_X1 U12614 ( .A(n12795), .B(n12796), .Z(n12794) );
  NAND2_X1 U12615 ( .A1(b_21_), .A2(a_28_), .ZN(n12796) );
  NAND2_X1 U12616 ( .A1(a_27_), .A2(n12792), .ZN(n12515) );
  NAND2_X1 U12617 ( .A1(n12797), .A2(n12798), .ZN(n12792) );
  NAND2_X1 U12618 ( .A1(n12799), .A2(b_22_), .ZN(n12798) );
  NOR2_X1 U12619 ( .A1(n12800), .A2(n9136), .ZN(n12799) );
  NOR2_X1 U12620 ( .A1(n12521), .A2(n12523), .ZN(n12800) );
  NAND2_X1 U12621 ( .A1(n12521), .A2(n12523), .ZN(n12797) );
  NAND2_X1 U12622 ( .A1(n12801), .A2(n12802), .ZN(n12523) );
  NAND2_X1 U12623 ( .A1(n12803), .A2(b_22_), .ZN(n12802) );
  NOR2_X1 U12624 ( .A1(n12804), .A2(n9121), .ZN(n12803) );
  NOR2_X1 U12625 ( .A1(n12805), .A2(n12543), .ZN(n12804) );
  NAND2_X1 U12626 ( .A1(n12805), .A2(n12543), .ZN(n12801) );
  NAND2_X1 U12627 ( .A1(n12806), .A2(n12807), .ZN(n12543) );
  NAND2_X1 U12628 ( .A1(b_20_), .A2(n12808), .ZN(n12807) );
  NAND2_X1 U12629 ( .A1(n10486), .A2(n12809), .ZN(n12808) );
  NAND2_X1 U12630 ( .A1(a_31_), .A2(n10052), .ZN(n12809) );
  NAND2_X1 U12631 ( .A1(b_21_), .A2(n12810), .ZN(n12806) );
  NAND2_X1 U12632 ( .A1(n10489), .A2(n12811), .ZN(n12810) );
  NAND2_X1 U12633 ( .A1(a_30_), .A2(n10053), .ZN(n12811) );
  INV_X1 U12634 ( .A(n12544), .ZN(n12805) );
  NAND2_X1 U12635 ( .A1(n12812), .A2(n9025), .ZN(n12544) );
  NOR2_X1 U12636 ( .A1(n12294), .A2(n10052), .ZN(n12812) );
  XOR2_X1 U12637 ( .A(n12813), .B(n12814), .Z(n12521) );
  NOR2_X1 U12638 ( .A1(n9121), .A2(n10052), .ZN(n12814) );
  XNOR2_X1 U12639 ( .A(n12815), .B(n12816), .ZN(n12813) );
  XOR2_X1 U12640 ( .A(n12817), .B(n12818), .Z(n12493) );
  XOR2_X1 U12641 ( .A(n12819), .B(n12820), .Z(n12818) );
  XNOR2_X1 U12642 ( .A(n12821), .B(n12822), .ZN(n12485) );
  XNOR2_X1 U12643 ( .A(n12823), .B(n12824), .ZN(n12822) );
  XNOR2_X1 U12644 ( .A(n12825), .B(n12826), .ZN(n12459) );
  XOR2_X1 U12645 ( .A(n12827), .B(n12828), .Z(n12826) );
  XNOR2_X1 U12646 ( .A(n12829), .B(n12830), .ZN(n12430) );
  NAND2_X1 U12647 ( .A1(n12831), .A2(n12832), .ZN(n12829) );
  XNOR2_X1 U12648 ( .A(n12833), .B(n12834), .ZN(n12562) );
  NAND2_X1 U12649 ( .A1(n12835), .A2(n12836), .ZN(n12833) );
  XNOR2_X1 U12650 ( .A(n12837), .B(n12838), .ZN(n12582) );
  XNOR2_X1 U12651 ( .A(n12839), .B(n12840), .ZN(n12837) );
  NOR2_X1 U12652 ( .A1(n10052), .A2(n9773), .ZN(n12840) );
  XNOR2_X1 U12653 ( .A(n12841), .B(n12842), .ZN(n12094) );
  NAND2_X1 U12654 ( .A1(n12843), .A2(n12844), .ZN(n12841) );
  XOR2_X1 U12655 ( .A(n12845), .B(n12846), .Z(n10295) );
  XNOR2_X1 U12656 ( .A(n12847), .B(n12848), .ZN(n12846) );
  INV_X1 U12657 ( .A(n12849), .ZN(n10170) );
  NOR2_X1 U12658 ( .A1(n10287), .A2(n12850), .ZN(n12849) );
  NAND2_X1 U12659 ( .A1(n10284), .A2(n12851), .ZN(n12850) );
  INV_X1 U12660 ( .A(n12852), .ZN(n12851) );
  NOR2_X1 U12661 ( .A1(n10288), .A2(n10289), .ZN(n12852) );
  NAND2_X1 U12662 ( .A1(n12598), .A2(n12599), .ZN(n10287) );
  XNOR2_X1 U12663 ( .A(n12853), .B(n12854), .ZN(n12599) );
  NAND2_X1 U12664 ( .A1(n12855), .A2(n12856), .ZN(n12853) );
  NOR2_X1 U12665 ( .A1(n12857), .A2(n12858), .ZN(n12598) );
  INV_X1 U12666 ( .A(n12859), .ZN(n12858) );
  NAND2_X1 U12667 ( .A1(n12845), .A2(n12860), .ZN(n12859) );
  NAND2_X1 U12668 ( .A1(n12848), .A2(n12847), .ZN(n12860) );
  XOR2_X1 U12669 ( .A(n12861), .B(n12862), .Z(n12845) );
  XOR2_X1 U12670 ( .A(n12863), .B(n12864), .Z(n12861) );
  NOR2_X1 U12671 ( .A1(n12847), .A2(n12848), .ZN(n12857) );
  NOR2_X1 U12672 ( .A1(n10093), .A2(n10052), .ZN(n12848) );
  NAND2_X1 U12673 ( .A1(n12843), .A2(n12865), .ZN(n12847) );
  NAND2_X1 U12674 ( .A1(n12842), .A2(n12844), .ZN(n12865) );
  NAND2_X1 U12675 ( .A1(n12866), .A2(n12867), .ZN(n12844) );
  NAND2_X1 U12676 ( .A1(a_1_), .A2(b_21_), .ZN(n12866) );
  XNOR2_X1 U12677 ( .A(n12868), .B(n12869), .ZN(n12842) );
  NAND2_X1 U12678 ( .A1(n12870), .A2(n12871), .ZN(n12868) );
  NAND2_X1 U12679 ( .A1(n12872), .A2(a_1_), .ZN(n12843) );
  INV_X1 U12680 ( .A(n12867), .ZN(n12872) );
  NAND2_X1 U12681 ( .A1(n12873), .A2(n12874), .ZN(n12867) );
  NAND2_X1 U12682 ( .A1(n12608), .A2(n12875), .ZN(n12874) );
  NAND2_X1 U12683 ( .A1(n12611), .A2(n12610), .ZN(n12875) );
  XOR2_X1 U12684 ( .A(n12876), .B(n12877), .Z(n12608) );
  NAND2_X1 U12685 ( .A1(n12878), .A2(n12879), .ZN(n12876) );
  INV_X1 U12686 ( .A(n12880), .ZN(n12873) );
  NOR2_X1 U12687 ( .A1(n12610), .A2(n12611), .ZN(n12880) );
  NOR2_X1 U12688 ( .A1(n10088), .A2(n10052), .ZN(n12611) );
  NAND2_X1 U12689 ( .A1(n12618), .A2(n12881), .ZN(n12610) );
  NAND2_X1 U12690 ( .A1(n12617), .A2(n12619), .ZN(n12881) );
  NAND2_X1 U12691 ( .A1(n12882), .A2(n12883), .ZN(n12619) );
  NAND2_X1 U12692 ( .A1(a_3_), .A2(b_21_), .ZN(n12882) );
  XNOR2_X1 U12693 ( .A(n12884), .B(n12885), .ZN(n12617) );
  NAND2_X1 U12694 ( .A1(n12886), .A2(n12887), .ZN(n12884) );
  NAND2_X1 U12695 ( .A1(n12888), .A2(a_3_), .ZN(n12618) );
  INV_X1 U12696 ( .A(n12883), .ZN(n12888) );
  NAND2_X1 U12697 ( .A1(n12889), .A2(n12890), .ZN(n12883) );
  NAND2_X1 U12698 ( .A1(n12624), .A2(n12891), .ZN(n12890) );
  NAND2_X1 U12699 ( .A1(n12627), .A2(n12626), .ZN(n12891) );
  XOR2_X1 U12700 ( .A(n12892), .B(n12893), .Z(n12624) );
  NAND2_X1 U12701 ( .A1(n12894), .A2(n12895), .ZN(n12892) );
  INV_X1 U12702 ( .A(n12896), .ZN(n12889) );
  NOR2_X1 U12703 ( .A1(n12626), .A2(n12627), .ZN(n12896) );
  NOR2_X1 U12704 ( .A1(n10085), .A2(n10052), .ZN(n12627) );
  NAND2_X1 U12705 ( .A1(n12897), .A2(n12898), .ZN(n12626) );
  NAND2_X1 U12706 ( .A1(n12899), .A2(a_5_), .ZN(n12898) );
  NOR2_X1 U12707 ( .A1(n12900), .A2(n10052), .ZN(n12899) );
  NOR2_X1 U12708 ( .A1(n12634), .A2(n12633), .ZN(n12900) );
  NAND2_X1 U12709 ( .A1(n12634), .A2(n12633), .ZN(n12897) );
  XNOR2_X1 U12710 ( .A(n12901), .B(n12902), .ZN(n12633) );
  NAND2_X1 U12711 ( .A1(n12903), .A2(n12904), .ZN(n12901) );
  NOR2_X1 U12712 ( .A1(n12905), .A2(n12906), .ZN(n12634) );
  INV_X1 U12713 ( .A(n12907), .ZN(n12906) );
  NAND2_X1 U12714 ( .A1(n12640), .A2(n12908), .ZN(n12907) );
  NAND2_X1 U12715 ( .A1(n12643), .A2(n12642), .ZN(n12908) );
  XNOR2_X1 U12716 ( .A(n12909), .B(n12910), .ZN(n12640) );
  XOR2_X1 U12717 ( .A(n12911), .B(n12912), .Z(n12909) );
  NOR2_X1 U12718 ( .A1(n9773), .A2(n10053), .ZN(n12912) );
  NOR2_X1 U12719 ( .A1(n12642), .A2(n12643), .ZN(n12905) );
  NOR2_X1 U12720 ( .A1(n10081), .A2(n10052), .ZN(n12643) );
  NAND2_X1 U12721 ( .A1(n12913), .A2(n12914), .ZN(n12642) );
  NAND2_X1 U12722 ( .A1(n12915), .A2(a_7_), .ZN(n12914) );
  NOR2_X1 U12723 ( .A1(n12916), .A2(n10052), .ZN(n12915) );
  NOR2_X1 U12724 ( .A1(n12839), .A2(n12838), .ZN(n12916) );
  NAND2_X1 U12725 ( .A1(n12839), .A2(n12838), .ZN(n12913) );
  XNOR2_X1 U12726 ( .A(n12917), .B(n12918), .ZN(n12838) );
  NAND2_X1 U12727 ( .A1(n12919), .A2(n12920), .ZN(n12917) );
  NOR2_X1 U12728 ( .A1(n12921), .A2(n12922), .ZN(n12839) );
  INV_X1 U12729 ( .A(n12923), .ZN(n12922) );
  NAND2_X1 U12730 ( .A1(n12653), .A2(n12924), .ZN(n12923) );
  NAND2_X1 U12731 ( .A1(n12655), .A2(n12654), .ZN(n12924) );
  XOR2_X1 U12732 ( .A(n12925), .B(n12926), .Z(n12653) );
  XOR2_X1 U12733 ( .A(n12927), .B(n12928), .Z(n12926) );
  NAND2_X1 U12734 ( .A1(b_20_), .A2(a_9_), .ZN(n12928) );
  NOR2_X1 U12735 ( .A1(n12654), .A2(n12655), .ZN(n12921) );
  NOR2_X1 U12736 ( .A1(n10079), .A2(n10052), .ZN(n12655) );
  NAND2_X1 U12737 ( .A1(n12662), .A2(n12929), .ZN(n12654) );
  NAND2_X1 U12738 ( .A1(n12661), .A2(n12663), .ZN(n12929) );
  NAND2_X1 U12739 ( .A1(n12930), .A2(n12931), .ZN(n12663) );
  NAND2_X1 U12740 ( .A1(a_9_), .A2(b_21_), .ZN(n12931) );
  INV_X1 U12741 ( .A(n12932), .ZN(n12930) );
  XNOR2_X1 U12742 ( .A(n12933), .B(n12934), .ZN(n12661) );
  XOR2_X1 U12743 ( .A(n12935), .B(n12936), .Z(n12934) );
  NAND2_X1 U12744 ( .A1(b_20_), .A2(a_10_), .ZN(n12936) );
  NAND2_X1 U12745 ( .A1(a_9_), .A2(n12932), .ZN(n12662) );
  NAND2_X1 U12746 ( .A1(n12937), .A2(n12938), .ZN(n12932) );
  NAND2_X1 U12747 ( .A1(n12939), .A2(a_10_), .ZN(n12938) );
  NOR2_X1 U12748 ( .A1(n12940), .A2(n10052), .ZN(n12939) );
  NOR2_X1 U12749 ( .A1(n12667), .A2(n12669), .ZN(n12940) );
  NAND2_X1 U12750 ( .A1(n12667), .A2(n12669), .ZN(n12937) );
  NAND2_X1 U12751 ( .A1(n12941), .A2(n12942), .ZN(n12669) );
  NAND2_X1 U12752 ( .A1(n12943), .A2(a_11_), .ZN(n12942) );
  NOR2_X1 U12753 ( .A1(n12944), .A2(n10052), .ZN(n12943) );
  NOR2_X1 U12754 ( .A1(n12676), .A2(n12677), .ZN(n12944) );
  NAND2_X1 U12755 ( .A1(n12676), .A2(n12677), .ZN(n12941) );
  NAND2_X1 U12756 ( .A1(n12686), .A2(n12945), .ZN(n12677) );
  NAND2_X1 U12757 ( .A1(n12685), .A2(n12687), .ZN(n12945) );
  NAND2_X1 U12758 ( .A1(n12946), .A2(n12947), .ZN(n12687) );
  NAND2_X1 U12759 ( .A1(a_12_), .A2(b_21_), .ZN(n12947) );
  INV_X1 U12760 ( .A(n12948), .ZN(n12946) );
  XNOR2_X1 U12761 ( .A(n12949), .B(n12950), .ZN(n12685) );
  NAND2_X1 U12762 ( .A1(n12951), .A2(n12952), .ZN(n12949) );
  NAND2_X1 U12763 ( .A1(a_12_), .A2(n12948), .ZN(n12686) );
  NAND2_X1 U12764 ( .A1(n12835), .A2(n12953), .ZN(n12948) );
  NAND2_X1 U12765 ( .A1(n12834), .A2(n12836), .ZN(n12953) );
  NAND2_X1 U12766 ( .A1(n12954), .A2(n12955), .ZN(n12836) );
  NAND2_X1 U12767 ( .A1(a_13_), .A2(b_21_), .ZN(n12955) );
  INV_X1 U12768 ( .A(n12956), .ZN(n12954) );
  XOR2_X1 U12769 ( .A(n12957), .B(n12958), .Z(n12834) );
  XNOR2_X1 U12770 ( .A(n12959), .B(n12960), .ZN(n12958) );
  NAND2_X1 U12771 ( .A1(a_13_), .A2(n12956), .ZN(n12835) );
  NAND2_X1 U12772 ( .A1(n12961), .A2(n12962), .ZN(n12956) );
  NAND2_X1 U12773 ( .A1(n12963), .A2(a_14_), .ZN(n12962) );
  NOR2_X1 U12774 ( .A1(n12964), .A2(n10052), .ZN(n12963) );
  NOR2_X1 U12775 ( .A1(n12695), .A2(n12697), .ZN(n12964) );
  NAND2_X1 U12776 ( .A1(n12695), .A2(n12697), .ZN(n12961) );
  NAND2_X1 U12777 ( .A1(n12965), .A2(n12966), .ZN(n12697) );
  NAND2_X1 U12778 ( .A1(n12967), .A2(a_15_), .ZN(n12966) );
  NOR2_X1 U12779 ( .A1(n12968), .A2(n10052), .ZN(n12967) );
  NOR2_X1 U12780 ( .A1(n12704), .A2(n12705), .ZN(n12968) );
  NAND2_X1 U12781 ( .A1(n12704), .A2(n12705), .ZN(n12965) );
  NAND2_X1 U12782 ( .A1(n12831), .A2(n12969), .ZN(n12705) );
  NAND2_X1 U12783 ( .A1(n12830), .A2(n12832), .ZN(n12969) );
  NAND2_X1 U12784 ( .A1(n12970), .A2(n12971), .ZN(n12832) );
  NAND2_X1 U12785 ( .A1(a_16_), .A2(b_21_), .ZN(n12971) );
  INV_X1 U12786 ( .A(n12972), .ZN(n12970) );
  XNOR2_X1 U12787 ( .A(n12973), .B(n12974), .ZN(n12830) );
  NAND2_X1 U12788 ( .A1(n12975), .A2(n12976), .ZN(n12973) );
  NAND2_X1 U12789 ( .A1(a_16_), .A2(n12972), .ZN(n12831) );
  NAND2_X1 U12790 ( .A1(n12718), .A2(n12977), .ZN(n12972) );
  NAND2_X1 U12791 ( .A1(n12717), .A2(n12719), .ZN(n12977) );
  NAND2_X1 U12792 ( .A1(n12978), .A2(n12979), .ZN(n12719) );
  NAND2_X1 U12793 ( .A1(a_17_), .A2(b_21_), .ZN(n12979) );
  INV_X1 U12794 ( .A(n12980), .ZN(n12978) );
  XOR2_X1 U12795 ( .A(n12981), .B(n12982), .Z(n12717) );
  XNOR2_X1 U12796 ( .A(n12983), .B(n12984), .ZN(n12982) );
  NAND2_X1 U12797 ( .A1(a_17_), .A2(n12980), .ZN(n12718) );
  NAND2_X1 U12798 ( .A1(n12726), .A2(n12985), .ZN(n12980) );
  NAND2_X1 U12799 ( .A1(n12725), .A2(n12727), .ZN(n12985) );
  NAND2_X1 U12800 ( .A1(n12986), .A2(n12987), .ZN(n12727) );
  NAND2_X1 U12801 ( .A1(a_18_), .A2(b_21_), .ZN(n12987) );
  INV_X1 U12802 ( .A(n12988), .ZN(n12986) );
  XNOR2_X1 U12803 ( .A(n12989), .B(n12990), .ZN(n12725) );
  XOR2_X1 U12804 ( .A(n12991), .B(n12992), .Z(n12990) );
  NAND2_X1 U12805 ( .A1(b_20_), .A2(a_19_), .ZN(n12992) );
  NAND2_X1 U12806 ( .A1(a_18_), .A2(n12988), .ZN(n12726) );
  NAND2_X1 U12807 ( .A1(n12993), .A2(n12994), .ZN(n12988) );
  NAND2_X1 U12808 ( .A1(n12995), .A2(a_19_), .ZN(n12994) );
  NOR2_X1 U12809 ( .A1(n12996), .A2(n10052), .ZN(n12995) );
  NOR2_X1 U12810 ( .A1(n12734), .A2(n12732), .ZN(n12996) );
  NAND2_X1 U12811 ( .A1(n12734), .A2(n12732), .ZN(n12993) );
  XNOR2_X1 U12812 ( .A(n12997), .B(n12998), .ZN(n12732) );
  XNOR2_X1 U12813 ( .A(n10055), .B(n12999), .ZN(n12998) );
  INV_X1 U12814 ( .A(n13000), .ZN(n12734) );
  NAND2_X1 U12815 ( .A1(n13001), .A2(n13002), .ZN(n13000) );
  NAND2_X1 U12816 ( .A1(n12825), .A2(n13003), .ZN(n13002) );
  INV_X1 U12817 ( .A(n13004), .ZN(n13003) );
  NOR2_X1 U12818 ( .A1(n12827), .A2(n12828), .ZN(n13004) );
  XOR2_X1 U12819 ( .A(n13005), .B(n13006), .Z(n12825) );
  NAND2_X1 U12820 ( .A1(n13007), .A2(n13008), .ZN(n13005) );
  NAND2_X1 U12821 ( .A1(n12828), .A2(n12827), .ZN(n13001) );
  NAND2_X1 U12822 ( .A1(n13009), .A2(n13010), .ZN(n12827) );
  NAND2_X1 U12823 ( .A1(n12745), .A2(n13011), .ZN(n13010) );
  NAND2_X1 U12824 ( .A1(n12747), .A2(n13012), .ZN(n13011) );
  INV_X1 U12825 ( .A(n10013), .ZN(n12747) );
  XOR2_X1 U12826 ( .A(n13013), .B(n13014), .Z(n12745) );
  NAND2_X1 U12827 ( .A1(n13015), .A2(n13016), .ZN(n13013) );
  NAND2_X1 U12828 ( .A1(n12746), .A2(n10013), .ZN(n13009) );
  NAND2_X1 U12829 ( .A1(b_21_), .A2(a_21_), .ZN(n10013) );
  INV_X1 U12830 ( .A(n13012), .ZN(n12746) );
  NAND2_X1 U12831 ( .A1(n12753), .A2(n13017), .ZN(n13012) );
  NAND2_X1 U12832 ( .A1(n12752), .A2(n12754), .ZN(n13017) );
  NAND2_X1 U12833 ( .A1(n13018), .A2(n13019), .ZN(n12754) );
  NAND2_X1 U12834 ( .A1(b_21_), .A2(a_22_), .ZN(n13019) );
  INV_X1 U12835 ( .A(n13020), .ZN(n13018) );
  XOR2_X1 U12836 ( .A(n13021), .B(n13022), .Z(n12752) );
  XOR2_X1 U12837 ( .A(n13023), .B(n13024), .Z(n13021) );
  NOR2_X1 U12838 ( .A1(n10051), .A2(n10053), .ZN(n13024) );
  NAND2_X1 U12839 ( .A1(a_22_), .A2(n13020), .ZN(n12753) );
  NAND2_X1 U12840 ( .A1(n13025), .A2(n13026), .ZN(n13020) );
  NAND2_X1 U12841 ( .A1(n13027), .A2(b_21_), .ZN(n13026) );
  NOR2_X1 U12842 ( .A1(n13028), .A2(n10051), .ZN(n13027) );
  NOR2_X1 U12843 ( .A1(n12760), .A2(n12761), .ZN(n13028) );
  NAND2_X1 U12844 ( .A1(n12760), .A2(n12761), .ZN(n13025) );
  NAND2_X1 U12845 ( .A1(n13029), .A2(n13030), .ZN(n12761) );
  INV_X1 U12846 ( .A(n13031), .ZN(n13030) );
  NOR2_X1 U12847 ( .A1(n13032), .A2(n13033), .ZN(n13031) );
  NOR2_X1 U12848 ( .A1(n12823), .A2(n12821), .ZN(n13033) );
  INV_X1 U12849 ( .A(n12824), .ZN(n13032) );
  NOR2_X1 U12850 ( .A1(n10052), .A2(n10050), .ZN(n12824) );
  NAND2_X1 U12851 ( .A1(n12821), .A2(n12823), .ZN(n13029) );
  NAND2_X1 U12852 ( .A1(n13034), .A2(n13035), .ZN(n12823) );
  NAND2_X1 U12853 ( .A1(n12820), .A2(n13036), .ZN(n13035) );
  INV_X1 U12854 ( .A(n13037), .ZN(n13036) );
  NOR2_X1 U12855 ( .A1(n12817), .A2(n12819), .ZN(n13037) );
  NOR2_X1 U12856 ( .A1(n10052), .A2(n10048), .ZN(n12820) );
  NAND2_X1 U12857 ( .A1(n12819), .A2(n12817), .ZN(n13034) );
  XOR2_X1 U12858 ( .A(n13038), .B(n13039), .Z(n12817) );
  XNOR2_X1 U12859 ( .A(n13040), .B(n13041), .ZN(n13039) );
  NOR2_X1 U12860 ( .A1(n13042), .A2(n13043), .ZN(n12819) );
  INV_X1 U12861 ( .A(n13044), .ZN(n13043) );
  NAND2_X1 U12862 ( .A1(n12777), .A2(n13045), .ZN(n13044) );
  NAND2_X1 U12863 ( .A1(n12780), .A2(n12779), .ZN(n13045) );
  XOR2_X1 U12864 ( .A(n13046), .B(n13047), .Z(n12777) );
  NAND2_X1 U12865 ( .A1(n13048), .A2(n13049), .ZN(n13046) );
  NOR2_X1 U12866 ( .A1(n12779), .A2(n12780), .ZN(n13042) );
  NOR2_X1 U12867 ( .A1(n10052), .A2(n10047), .ZN(n12780) );
  NAND2_X1 U12868 ( .A1(n12786), .A2(n13050), .ZN(n12779) );
  NAND2_X1 U12869 ( .A1(n12785), .A2(n12787), .ZN(n13050) );
  NAND2_X1 U12870 ( .A1(n13051), .A2(n13052), .ZN(n12787) );
  NAND2_X1 U12871 ( .A1(b_21_), .A2(a_27_), .ZN(n13052) );
  INV_X1 U12872 ( .A(n13053), .ZN(n13051) );
  XNOR2_X1 U12873 ( .A(n13054), .B(n13055), .ZN(n12785) );
  XOR2_X1 U12874 ( .A(n13056), .B(n13057), .Z(n13055) );
  NAND2_X1 U12875 ( .A1(b_20_), .A2(a_28_), .ZN(n13057) );
  NAND2_X1 U12876 ( .A1(a_27_), .A2(n13053), .ZN(n12786) );
  NAND2_X1 U12877 ( .A1(n13058), .A2(n13059), .ZN(n13053) );
  NAND2_X1 U12878 ( .A1(n13060), .A2(b_21_), .ZN(n13059) );
  NOR2_X1 U12879 ( .A1(n13061), .A2(n9136), .ZN(n13060) );
  NOR2_X1 U12880 ( .A1(n12793), .A2(n12795), .ZN(n13061) );
  NAND2_X1 U12881 ( .A1(n12793), .A2(n12795), .ZN(n13058) );
  NAND2_X1 U12882 ( .A1(n13062), .A2(n13063), .ZN(n12795) );
  NAND2_X1 U12883 ( .A1(n13064), .A2(b_21_), .ZN(n13063) );
  NOR2_X1 U12884 ( .A1(n13065), .A2(n9121), .ZN(n13064) );
  NOR2_X1 U12885 ( .A1(n13066), .A2(n12815), .ZN(n13065) );
  NAND2_X1 U12886 ( .A1(n13066), .A2(n12815), .ZN(n13062) );
  NAND2_X1 U12887 ( .A1(n13067), .A2(n13068), .ZN(n12815) );
  NAND2_X1 U12888 ( .A1(b_19_), .A2(n13069), .ZN(n13068) );
  NAND2_X1 U12889 ( .A1(n10486), .A2(n13070), .ZN(n13069) );
  NAND2_X1 U12890 ( .A1(a_31_), .A2(n10053), .ZN(n13070) );
  NAND2_X1 U12891 ( .A1(b_20_), .A2(n13071), .ZN(n13067) );
  NAND2_X1 U12892 ( .A1(n10489), .A2(n13072), .ZN(n13071) );
  NAND2_X1 U12893 ( .A1(a_30_), .A2(n10056), .ZN(n13072) );
  INV_X1 U12894 ( .A(n12816), .ZN(n13066) );
  NAND2_X1 U12895 ( .A1(n13073), .A2(n9025), .ZN(n12816) );
  NOR2_X1 U12896 ( .A1(n10052), .A2(n10053), .ZN(n13073) );
  XOR2_X1 U12897 ( .A(n13074), .B(n13075), .Z(n12793) );
  NOR2_X1 U12898 ( .A1(n9121), .A2(n10053), .ZN(n13075) );
  XNOR2_X1 U12899 ( .A(n13076), .B(n13077), .ZN(n13074) );
  XNOR2_X1 U12900 ( .A(n13078), .B(n13079), .ZN(n12821) );
  XNOR2_X1 U12901 ( .A(n13080), .B(n13081), .ZN(n13079) );
  XNOR2_X1 U12902 ( .A(n13082), .B(n13083), .ZN(n12760) );
  XNOR2_X1 U12903 ( .A(n13084), .B(n13085), .ZN(n13083) );
  NAND2_X1 U12904 ( .A1(a_20_), .A2(b_21_), .ZN(n12828) );
  XNOR2_X1 U12905 ( .A(n13086), .B(n13087), .ZN(n12704) );
  NAND2_X1 U12906 ( .A1(n13088), .A2(n13089), .ZN(n13086) );
  XNOR2_X1 U12907 ( .A(n13090), .B(n13091), .ZN(n12695) );
  NAND2_X1 U12908 ( .A1(n13092), .A2(n13093), .ZN(n13090) );
  XOR2_X1 U12909 ( .A(n13094), .B(n13095), .Z(n12676) );
  XOR2_X1 U12910 ( .A(n13096), .B(n13097), .Z(n13094) );
  NOR2_X1 U12911 ( .A1(n10070), .A2(n10053), .ZN(n13097) );
  XNOR2_X1 U12912 ( .A(n13098), .B(n13099), .ZN(n12667) );
  XOR2_X1 U12913 ( .A(n13100), .B(n13101), .Z(n13099) );
  NAND2_X1 U12914 ( .A1(b_20_), .A2(a_11_), .ZN(n13101) );
  INV_X1 U12915 ( .A(n13102), .ZN(n10183) );
  NOR2_X1 U12916 ( .A1(n10284), .A2(n10283), .ZN(n13102) );
  NAND2_X1 U12917 ( .A1(n13103), .A2(n13104), .ZN(n10283) );
  NAND2_X1 U12918 ( .A1(n13105), .A2(n13106), .ZN(n13104) );
  INV_X1 U12919 ( .A(n10278), .ZN(n13103) );
  NOR2_X1 U12920 ( .A1(n13106), .A2(n13105), .ZN(n10278) );
  INV_X1 U12921 ( .A(n13107), .ZN(n13105) );
  NAND2_X1 U12922 ( .A1(n13108), .A2(n13109), .ZN(n13107) );
  NAND2_X1 U12923 ( .A1(n13110), .A2(b_19_), .ZN(n13109) );
  NOR2_X1 U12924 ( .A1(n13111), .A2(n10093), .ZN(n13110) );
  NOR2_X1 U12925 ( .A1(n13112), .A2(n13113), .ZN(n13111) );
  NAND2_X1 U12926 ( .A1(n13112), .A2(n13113), .ZN(n13108) );
  XNOR2_X1 U12927 ( .A(n13114), .B(n13115), .ZN(n13106) );
  XOR2_X1 U12928 ( .A(n13116), .B(n13117), .Z(n13114) );
  NAND2_X1 U12929 ( .A1(n10288), .A2(n10289), .ZN(n10284) );
  NAND2_X1 U12930 ( .A1(n12855), .A2(n13118), .ZN(n10289) );
  NAND2_X1 U12931 ( .A1(n12854), .A2(n12856), .ZN(n13118) );
  NAND2_X1 U12932 ( .A1(n13119), .A2(n13120), .ZN(n12856) );
  NAND2_X1 U12933 ( .A1(b_20_), .A2(a_0_), .ZN(n13119) );
  XOR2_X1 U12934 ( .A(n13121), .B(n13122), .Z(n12854) );
  XNOR2_X1 U12935 ( .A(n13123), .B(n13124), .ZN(n13122) );
  NAND2_X1 U12936 ( .A1(n13125), .A2(a_0_), .ZN(n12855) );
  INV_X1 U12937 ( .A(n13120), .ZN(n13125) );
  NAND2_X1 U12938 ( .A1(n13126), .A2(n13127), .ZN(n13120) );
  NAND2_X1 U12939 ( .A1(n12862), .A2(n13128), .ZN(n13127) );
  NAND2_X1 U12940 ( .A1(n12864), .A2(n12863), .ZN(n13128) );
  XNOR2_X1 U12941 ( .A(n13129), .B(n13130), .ZN(n12862) );
  NOR2_X1 U12942 ( .A1(n13131), .A2(n13132), .ZN(n13130) );
  INV_X1 U12943 ( .A(n13133), .ZN(n13132) );
  NOR2_X1 U12944 ( .A1(n13134), .A2(n13135), .ZN(n13131) );
  NOR2_X1 U12945 ( .A1(n10088), .A2(n10056), .ZN(n13135) );
  INV_X1 U12946 ( .A(n13136), .ZN(n13126) );
  NOR2_X1 U12947 ( .A1(n12863), .A2(n12864), .ZN(n13136) );
  NOR2_X1 U12948 ( .A1(n10053), .A2(n9983), .ZN(n12864) );
  NAND2_X1 U12949 ( .A1(n12870), .A2(n13137), .ZN(n12863) );
  NAND2_X1 U12950 ( .A1(n12869), .A2(n12871), .ZN(n13137) );
  NAND2_X1 U12951 ( .A1(n13138), .A2(n13139), .ZN(n12871) );
  NAND2_X1 U12952 ( .A1(b_20_), .A2(a_2_), .ZN(n13139) );
  INV_X1 U12953 ( .A(n13140), .ZN(n13138) );
  XNOR2_X1 U12954 ( .A(n13141), .B(n13142), .ZN(n12869) );
  XOR2_X1 U12955 ( .A(n13143), .B(n13144), .Z(n13141) );
  NAND2_X1 U12956 ( .A1(a_2_), .A2(n13140), .ZN(n12870) );
  NAND2_X1 U12957 ( .A1(n12878), .A2(n13145), .ZN(n13140) );
  NAND2_X1 U12958 ( .A1(n12877), .A2(n12879), .ZN(n13145) );
  NAND2_X1 U12959 ( .A1(n13146), .A2(n13147), .ZN(n12879) );
  NAND2_X1 U12960 ( .A1(b_20_), .A2(a_3_), .ZN(n13147) );
  INV_X1 U12961 ( .A(n13148), .ZN(n13146) );
  XNOR2_X1 U12962 ( .A(n13149), .B(n13150), .ZN(n12877) );
  NAND2_X1 U12963 ( .A1(n13151), .A2(n13152), .ZN(n13149) );
  NAND2_X1 U12964 ( .A1(a_3_), .A2(n13148), .ZN(n12878) );
  NAND2_X1 U12965 ( .A1(n12886), .A2(n13153), .ZN(n13148) );
  NAND2_X1 U12966 ( .A1(n12885), .A2(n12887), .ZN(n13153) );
  NAND2_X1 U12967 ( .A1(n13154), .A2(n13155), .ZN(n12887) );
  NAND2_X1 U12968 ( .A1(b_20_), .A2(a_4_), .ZN(n13155) );
  INV_X1 U12969 ( .A(n13156), .ZN(n13154) );
  XOR2_X1 U12970 ( .A(n13157), .B(n13158), .Z(n12885) );
  XNOR2_X1 U12971 ( .A(n13159), .B(n13160), .ZN(n13158) );
  NAND2_X1 U12972 ( .A1(a_4_), .A2(n13156), .ZN(n12886) );
  NAND2_X1 U12973 ( .A1(n12894), .A2(n13161), .ZN(n13156) );
  NAND2_X1 U12974 ( .A1(n12893), .A2(n12895), .ZN(n13161) );
  NAND2_X1 U12975 ( .A1(n13162), .A2(n13163), .ZN(n12895) );
  NAND2_X1 U12976 ( .A1(b_20_), .A2(a_5_), .ZN(n13163) );
  INV_X1 U12977 ( .A(n13164), .ZN(n13162) );
  XNOR2_X1 U12978 ( .A(n13165), .B(n13166), .ZN(n12893) );
  NAND2_X1 U12979 ( .A1(n13167), .A2(n13168), .ZN(n13165) );
  NAND2_X1 U12980 ( .A1(a_5_), .A2(n13164), .ZN(n12894) );
  NAND2_X1 U12981 ( .A1(n12903), .A2(n13169), .ZN(n13164) );
  NAND2_X1 U12982 ( .A1(n12902), .A2(n12904), .ZN(n13169) );
  NAND2_X1 U12983 ( .A1(n13170), .A2(n13171), .ZN(n12904) );
  NAND2_X1 U12984 ( .A1(b_20_), .A2(a_6_), .ZN(n13171) );
  INV_X1 U12985 ( .A(n13172), .ZN(n13170) );
  XOR2_X1 U12986 ( .A(n13173), .B(n13174), .Z(n12902) );
  XNOR2_X1 U12987 ( .A(n13175), .B(n13176), .ZN(n13174) );
  NAND2_X1 U12988 ( .A1(a_6_), .A2(n13172), .ZN(n12903) );
  NAND2_X1 U12989 ( .A1(n13177), .A2(n13178), .ZN(n13172) );
  NAND2_X1 U12990 ( .A1(n13179), .A2(b_20_), .ZN(n13178) );
  NOR2_X1 U12991 ( .A1(n13180), .A2(n9773), .ZN(n13179) );
  NOR2_X1 U12992 ( .A1(n12910), .A2(n12911), .ZN(n13180) );
  NAND2_X1 U12993 ( .A1(n12910), .A2(n12911), .ZN(n13177) );
  NAND2_X1 U12994 ( .A1(n12919), .A2(n13181), .ZN(n12911) );
  NAND2_X1 U12995 ( .A1(n12918), .A2(n12920), .ZN(n13181) );
  NAND2_X1 U12996 ( .A1(n13182), .A2(n13183), .ZN(n12920) );
  NAND2_X1 U12997 ( .A1(b_20_), .A2(a_8_), .ZN(n13183) );
  INV_X1 U12998 ( .A(n13184), .ZN(n13182) );
  XOR2_X1 U12999 ( .A(n13185), .B(n13186), .Z(n12918) );
  XNOR2_X1 U13000 ( .A(n13187), .B(n13188), .ZN(n13186) );
  NAND2_X1 U13001 ( .A1(a_8_), .A2(n13184), .ZN(n12919) );
  NAND2_X1 U13002 ( .A1(n13189), .A2(n13190), .ZN(n13184) );
  NAND2_X1 U13003 ( .A1(n13191), .A2(b_20_), .ZN(n13190) );
  NOR2_X1 U13004 ( .A1(n13192), .A2(n10076), .ZN(n13191) );
  NOR2_X1 U13005 ( .A1(n12925), .A2(n12927), .ZN(n13192) );
  NAND2_X1 U13006 ( .A1(n12925), .A2(n12927), .ZN(n13189) );
  NAND2_X1 U13007 ( .A1(n13193), .A2(n13194), .ZN(n12927) );
  NAND2_X1 U13008 ( .A1(n13195), .A2(b_20_), .ZN(n13194) );
  NOR2_X1 U13009 ( .A1(n13196), .A2(n10073), .ZN(n13195) );
  NOR2_X1 U13010 ( .A1(n12933), .A2(n12935), .ZN(n13196) );
  NAND2_X1 U13011 ( .A1(n12933), .A2(n12935), .ZN(n13193) );
  NAND2_X1 U13012 ( .A1(n13197), .A2(n13198), .ZN(n12935) );
  NAND2_X1 U13013 ( .A1(n13199), .A2(b_20_), .ZN(n13198) );
  NOR2_X1 U13014 ( .A1(n13200), .A2(n9649), .ZN(n13199) );
  NOR2_X1 U13015 ( .A1(n13098), .A2(n13100), .ZN(n13200) );
  NAND2_X1 U13016 ( .A1(n13098), .A2(n13100), .ZN(n13197) );
  NAND2_X1 U13017 ( .A1(n13201), .A2(n13202), .ZN(n13100) );
  NAND2_X1 U13018 ( .A1(n13203), .A2(b_20_), .ZN(n13202) );
  NOR2_X1 U13019 ( .A1(n13204), .A2(n10070), .ZN(n13203) );
  NOR2_X1 U13020 ( .A1(n13095), .A2(n13096), .ZN(n13204) );
  NAND2_X1 U13021 ( .A1(n13095), .A2(n13096), .ZN(n13201) );
  NAND2_X1 U13022 ( .A1(n12951), .A2(n13205), .ZN(n13096) );
  NAND2_X1 U13023 ( .A1(n12950), .A2(n12952), .ZN(n13205) );
  NAND2_X1 U13024 ( .A1(n13206), .A2(n13207), .ZN(n12952) );
  NAND2_X1 U13025 ( .A1(b_20_), .A2(a_13_), .ZN(n13206) );
  XOR2_X1 U13026 ( .A(n13208), .B(n13209), .Z(n12950) );
  XOR2_X1 U13027 ( .A(n13210), .B(n13211), .Z(n13208) );
  NOR2_X1 U13028 ( .A1(n10065), .A2(n10056), .ZN(n13211) );
  NAND2_X1 U13029 ( .A1(n13212), .A2(a_13_), .ZN(n12951) );
  INV_X1 U13030 ( .A(n13207), .ZN(n13212) );
  NAND2_X1 U13031 ( .A1(n13213), .A2(n13214), .ZN(n13207) );
  NAND2_X1 U13032 ( .A1(n12957), .A2(n13215), .ZN(n13214) );
  NAND2_X1 U13033 ( .A1(n12960), .A2(n12959), .ZN(n13215) );
  XNOR2_X1 U13034 ( .A(n13216), .B(n13217), .ZN(n12957) );
  XOR2_X1 U13035 ( .A(n13218), .B(n13219), .Z(n13216) );
  NOR2_X1 U13036 ( .A1(n9534), .A2(n10056), .ZN(n13219) );
  INV_X1 U13037 ( .A(n13220), .ZN(n13213) );
  NOR2_X1 U13038 ( .A1(n12959), .A2(n12960), .ZN(n13220) );
  NOR2_X1 U13039 ( .A1(n10053), .A2(n10065), .ZN(n12960) );
  NAND2_X1 U13040 ( .A1(n13092), .A2(n13221), .ZN(n12959) );
  NAND2_X1 U13041 ( .A1(n13091), .A2(n13093), .ZN(n13221) );
  NAND2_X1 U13042 ( .A1(n13222), .A2(n13223), .ZN(n13093) );
  NAND2_X1 U13043 ( .A1(b_20_), .A2(a_15_), .ZN(n13223) );
  INV_X1 U13044 ( .A(n13224), .ZN(n13222) );
  XNOR2_X1 U13045 ( .A(n13225), .B(n13226), .ZN(n13091) );
  NAND2_X1 U13046 ( .A1(n13227), .A2(n13228), .ZN(n13225) );
  NAND2_X1 U13047 ( .A1(a_15_), .A2(n13224), .ZN(n13092) );
  NAND2_X1 U13048 ( .A1(n13088), .A2(n13229), .ZN(n13224) );
  NAND2_X1 U13049 ( .A1(n13087), .A2(n13089), .ZN(n13229) );
  NAND2_X1 U13050 ( .A1(n13230), .A2(n13231), .ZN(n13089) );
  NAND2_X1 U13051 ( .A1(b_20_), .A2(a_16_), .ZN(n13231) );
  INV_X1 U13052 ( .A(n13232), .ZN(n13230) );
  XNOR2_X1 U13053 ( .A(n13233), .B(n13234), .ZN(n13087) );
  NAND2_X1 U13054 ( .A1(n13235), .A2(n13236), .ZN(n13233) );
  NAND2_X1 U13055 ( .A1(a_16_), .A2(n13232), .ZN(n13088) );
  NAND2_X1 U13056 ( .A1(n12975), .A2(n13237), .ZN(n13232) );
  NAND2_X1 U13057 ( .A1(n12974), .A2(n12976), .ZN(n13237) );
  NAND2_X1 U13058 ( .A1(n13238), .A2(n13239), .ZN(n12976) );
  NAND2_X1 U13059 ( .A1(b_20_), .A2(a_17_), .ZN(n13238) );
  XOR2_X1 U13060 ( .A(n13240), .B(n13241), .Z(n12974) );
  XOR2_X1 U13061 ( .A(n13242), .B(n13243), .Z(n13240) );
  NAND2_X1 U13062 ( .A1(n13244), .A2(a_17_), .ZN(n12975) );
  INV_X1 U13063 ( .A(n13239), .ZN(n13244) );
  NAND2_X1 U13064 ( .A1(n13245), .A2(n13246), .ZN(n13239) );
  NAND2_X1 U13065 ( .A1(n12981), .A2(n13247), .ZN(n13246) );
  NAND2_X1 U13066 ( .A1(n12984), .A2(n12983), .ZN(n13247) );
  XOR2_X1 U13067 ( .A(n13248), .B(n13249), .Z(n12981) );
  XOR2_X1 U13068 ( .A(n13250), .B(n10009), .Z(n13249) );
  INV_X1 U13069 ( .A(n13251), .ZN(n13245) );
  NOR2_X1 U13070 ( .A1(n12983), .A2(n12984), .ZN(n13251) );
  NOR2_X1 U13071 ( .A1(n10053), .A2(n10058), .ZN(n12984) );
  NAND2_X1 U13072 ( .A1(n13252), .A2(n13253), .ZN(n12983) );
  NAND2_X1 U13073 ( .A1(n13254), .A2(b_20_), .ZN(n13253) );
  NOR2_X1 U13074 ( .A1(n13255), .A2(n9415), .ZN(n13254) );
  NOR2_X1 U13075 ( .A1(n12989), .A2(n12991), .ZN(n13255) );
  NAND2_X1 U13076 ( .A1(n12989), .A2(n12991), .ZN(n13252) );
  NAND2_X1 U13077 ( .A1(n13256), .A2(n13257), .ZN(n12991) );
  NAND2_X1 U13078 ( .A1(n12997), .A2(n13258), .ZN(n13257) );
  INV_X1 U13079 ( .A(n13259), .ZN(n13258) );
  NOR2_X1 U13080 ( .A1(n12999), .A2(n10055), .ZN(n13259) );
  XNOR2_X1 U13081 ( .A(n13260), .B(n13261), .ZN(n12997) );
  NAND2_X1 U13082 ( .A1(n13262), .A2(n13263), .ZN(n13260) );
  NAND2_X1 U13083 ( .A1(n10055), .A2(n12999), .ZN(n13256) );
  NAND2_X1 U13084 ( .A1(n13007), .A2(n13264), .ZN(n12999) );
  NAND2_X1 U13085 ( .A1(n13006), .A2(n13008), .ZN(n13264) );
  NAND2_X1 U13086 ( .A1(n13265), .A2(n13266), .ZN(n13008) );
  NAND2_X1 U13087 ( .A1(b_20_), .A2(a_21_), .ZN(n13266) );
  INV_X1 U13088 ( .A(n13267), .ZN(n13265) );
  XNOR2_X1 U13089 ( .A(n13268), .B(n13269), .ZN(n13006) );
  NAND2_X1 U13090 ( .A1(n13270), .A2(n13271), .ZN(n13268) );
  NAND2_X1 U13091 ( .A1(a_21_), .A2(n13267), .ZN(n13007) );
  NAND2_X1 U13092 ( .A1(n13015), .A2(n13272), .ZN(n13267) );
  NAND2_X1 U13093 ( .A1(n13014), .A2(n13016), .ZN(n13272) );
  NAND2_X1 U13094 ( .A1(n13273), .A2(n13274), .ZN(n13016) );
  NAND2_X1 U13095 ( .A1(b_20_), .A2(a_22_), .ZN(n13274) );
  INV_X1 U13096 ( .A(n13275), .ZN(n13273) );
  XOR2_X1 U13097 ( .A(n13276), .B(n13277), .Z(n13014) );
  XOR2_X1 U13098 ( .A(n13278), .B(n13279), .Z(n13276) );
  NOR2_X1 U13099 ( .A1(n10051), .A2(n10056), .ZN(n13279) );
  NAND2_X1 U13100 ( .A1(a_22_), .A2(n13275), .ZN(n13015) );
  NAND2_X1 U13101 ( .A1(n13280), .A2(n13281), .ZN(n13275) );
  NAND2_X1 U13102 ( .A1(n13282), .A2(b_20_), .ZN(n13281) );
  NOR2_X1 U13103 ( .A1(n13283), .A2(n10051), .ZN(n13282) );
  NOR2_X1 U13104 ( .A1(n13022), .A2(n13023), .ZN(n13283) );
  NAND2_X1 U13105 ( .A1(n13022), .A2(n13023), .ZN(n13280) );
  NAND2_X1 U13106 ( .A1(n13284), .A2(n13285), .ZN(n13023) );
  INV_X1 U13107 ( .A(n13286), .ZN(n13285) );
  NOR2_X1 U13108 ( .A1(n13287), .A2(n13288), .ZN(n13286) );
  NOR2_X1 U13109 ( .A1(n13084), .A2(n13082), .ZN(n13288) );
  INV_X1 U13110 ( .A(n13085), .ZN(n13287) );
  NOR2_X1 U13111 ( .A1(n10053), .A2(n10050), .ZN(n13085) );
  NAND2_X1 U13112 ( .A1(n13082), .A2(n13084), .ZN(n13284) );
  NAND2_X1 U13113 ( .A1(n13289), .A2(n13290), .ZN(n13084) );
  NAND2_X1 U13114 ( .A1(n13081), .A2(n13291), .ZN(n13290) );
  NAND2_X1 U13115 ( .A1(n13078), .A2(n13080), .ZN(n13291) );
  NOR2_X1 U13116 ( .A1(n10053), .A2(n10048), .ZN(n13081) );
  INV_X1 U13117 ( .A(n13292), .ZN(n13289) );
  NOR2_X1 U13118 ( .A1(n13080), .A2(n13078), .ZN(n13292) );
  XNOR2_X1 U13119 ( .A(n13293), .B(n13294), .ZN(n13078) );
  XNOR2_X1 U13120 ( .A(n13295), .B(n13296), .ZN(n13294) );
  NAND2_X1 U13121 ( .A1(n13297), .A2(n13298), .ZN(n13080) );
  NAND2_X1 U13122 ( .A1(n13038), .A2(n13299), .ZN(n13298) );
  NAND2_X1 U13123 ( .A1(n13041), .A2(n13040), .ZN(n13299) );
  XOR2_X1 U13124 ( .A(n13300), .B(n13301), .Z(n13038) );
  NAND2_X1 U13125 ( .A1(n13302), .A2(n13303), .ZN(n13300) );
  INV_X1 U13126 ( .A(n13304), .ZN(n13297) );
  NOR2_X1 U13127 ( .A1(n13040), .A2(n13041), .ZN(n13304) );
  NOR2_X1 U13128 ( .A1(n10053), .A2(n10047), .ZN(n13041) );
  NAND2_X1 U13129 ( .A1(n13048), .A2(n13305), .ZN(n13040) );
  NAND2_X1 U13130 ( .A1(n13047), .A2(n13049), .ZN(n13305) );
  NAND2_X1 U13131 ( .A1(n13306), .A2(n13307), .ZN(n13049) );
  NAND2_X1 U13132 ( .A1(b_20_), .A2(a_27_), .ZN(n13307) );
  INV_X1 U13133 ( .A(n13308), .ZN(n13306) );
  XNOR2_X1 U13134 ( .A(n13309), .B(n13310), .ZN(n13047) );
  XOR2_X1 U13135 ( .A(n13311), .B(n13312), .Z(n13310) );
  NAND2_X1 U13136 ( .A1(b_19_), .A2(a_28_), .ZN(n13312) );
  NAND2_X1 U13137 ( .A1(a_27_), .A2(n13308), .ZN(n13048) );
  NAND2_X1 U13138 ( .A1(n13313), .A2(n13314), .ZN(n13308) );
  NAND2_X1 U13139 ( .A1(n13315), .A2(b_20_), .ZN(n13314) );
  NOR2_X1 U13140 ( .A1(n13316), .A2(n9136), .ZN(n13315) );
  NOR2_X1 U13141 ( .A1(n13054), .A2(n13056), .ZN(n13316) );
  NAND2_X1 U13142 ( .A1(n13054), .A2(n13056), .ZN(n13313) );
  NAND2_X1 U13143 ( .A1(n13317), .A2(n13318), .ZN(n13056) );
  NAND2_X1 U13144 ( .A1(n13319), .A2(b_20_), .ZN(n13318) );
  NOR2_X1 U13145 ( .A1(n13320), .A2(n9121), .ZN(n13319) );
  NOR2_X1 U13146 ( .A1(n13321), .A2(n13076), .ZN(n13320) );
  NAND2_X1 U13147 ( .A1(n13321), .A2(n13076), .ZN(n13317) );
  NAND2_X1 U13148 ( .A1(n13322), .A2(n13323), .ZN(n13076) );
  NAND2_X1 U13149 ( .A1(b_18_), .A2(n13324), .ZN(n13323) );
  NAND2_X1 U13150 ( .A1(n10486), .A2(n13325), .ZN(n13324) );
  NAND2_X1 U13151 ( .A1(a_31_), .A2(n10056), .ZN(n13325) );
  NAND2_X1 U13152 ( .A1(b_19_), .A2(n13326), .ZN(n13322) );
  NAND2_X1 U13153 ( .A1(n10489), .A2(n13327), .ZN(n13326) );
  NAND2_X1 U13154 ( .A1(a_30_), .A2(n10057), .ZN(n13327) );
  INV_X1 U13155 ( .A(n13077), .ZN(n13321) );
  NAND2_X1 U13156 ( .A1(n13328), .A2(n9025), .ZN(n13077) );
  NOR2_X1 U13157 ( .A1(n10053), .A2(n10056), .ZN(n13328) );
  XOR2_X1 U13158 ( .A(n13329), .B(n13330), .Z(n13054) );
  NOR2_X1 U13159 ( .A1(n9121), .A2(n10056), .ZN(n13330) );
  XNOR2_X1 U13160 ( .A(n13331), .B(n13332), .ZN(n13329) );
  XNOR2_X1 U13161 ( .A(n13333), .B(n13334), .ZN(n13082) );
  XNOR2_X1 U13162 ( .A(n13335), .B(n13336), .ZN(n13334) );
  XNOR2_X1 U13163 ( .A(n13337), .B(n13338), .ZN(n13022) );
  XNOR2_X1 U13164 ( .A(n13339), .B(n13340), .ZN(n13338) );
  NOR2_X1 U13165 ( .A1(n10053), .A2(n10054), .ZN(n10055) );
  XOR2_X1 U13166 ( .A(n13341), .B(n13342), .Z(n12989) );
  XNOR2_X1 U13167 ( .A(n13343), .B(n13344), .ZN(n13342) );
  XNOR2_X1 U13168 ( .A(n13345), .B(n13346), .ZN(n13095) );
  NAND2_X1 U13169 ( .A1(n13347), .A2(n13348), .ZN(n13345) );
  XOR2_X1 U13170 ( .A(n13349), .B(n13350), .Z(n13098) );
  XOR2_X1 U13171 ( .A(n13351), .B(n13352), .Z(n13349) );
  XOR2_X1 U13172 ( .A(n13353), .B(n13354), .Z(n12933) );
  XNOR2_X1 U13173 ( .A(n13355), .B(n13356), .ZN(n13353) );
  XOR2_X1 U13174 ( .A(n13357), .B(n13358), .Z(n12925) );
  XOR2_X1 U13175 ( .A(n13359), .B(n13360), .Z(n13357) );
  NOR2_X1 U13176 ( .A1(n10073), .A2(n10056), .ZN(n13360) );
  XNOR2_X1 U13177 ( .A(n13361), .B(n13362), .ZN(n12910) );
  NAND2_X1 U13178 ( .A1(n13363), .A2(n13364), .ZN(n13361) );
  XOR2_X1 U13179 ( .A(n13113), .B(n13365), .Z(n10288) );
  XNOR2_X1 U13180 ( .A(n13112), .B(n13366), .ZN(n13365) );
  NAND2_X1 U13181 ( .A1(b_19_), .A2(a_0_), .ZN(n13366) );
  NOR2_X1 U13182 ( .A1(n13367), .A2(n13368), .ZN(n13112) );
  INV_X1 U13183 ( .A(n13369), .ZN(n13368) );
  NAND2_X1 U13184 ( .A1(n13121), .A2(n13370), .ZN(n13369) );
  NAND2_X1 U13185 ( .A1(n13124), .A2(n13123), .ZN(n13370) );
  XNOR2_X1 U13186 ( .A(n13371), .B(n13372), .ZN(n13121) );
  XOR2_X1 U13187 ( .A(n13373), .B(n13374), .Z(n13372) );
  NOR2_X1 U13188 ( .A1(n13123), .A2(n13124), .ZN(n13367) );
  NOR2_X1 U13189 ( .A1(n10056), .A2(n9983), .ZN(n13124) );
  NAND2_X1 U13190 ( .A1(n13133), .A2(n13375), .ZN(n13123) );
  NAND2_X1 U13191 ( .A1(n13129), .A2(n13376), .ZN(n13375) );
  NAND2_X1 U13192 ( .A1(n13377), .A2(n13378), .ZN(n13376) );
  NAND2_X1 U13193 ( .A1(b_19_), .A2(a_2_), .ZN(n13378) );
  INV_X1 U13194 ( .A(n13134), .ZN(n13377) );
  XNOR2_X1 U13195 ( .A(n13379), .B(n13380), .ZN(n13129) );
  XOR2_X1 U13196 ( .A(n13381), .B(n13382), .Z(n13379) );
  NAND2_X1 U13197 ( .A1(n13134), .A2(a_2_), .ZN(n13133) );
  NOR2_X1 U13198 ( .A1(n13383), .A2(n13384), .ZN(n13134) );
  INV_X1 U13199 ( .A(n13385), .ZN(n13384) );
  NAND2_X1 U13200 ( .A1(n13142), .A2(n13386), .ZN(n13385) );
  NAND2_X1 U13201 ( .A1(n13144), .A2(n13143), .ZN(n13386) );
  XOR2_X1 U13202 ( .A(n13387), .B(n13388), .Z(n13142) );
  XNOR2_X1 U13203 ( .A(n13389), .B(n13390), .ZN(n13387) );
  NOR2_X1 U13204 ( .A1(n13143), .A2(n13144), .ZN(n13383) );
  NOR2_X1 U13205 ( .A1(n10056), .A2(n10086), .ZN(n13144) );
  NAND2_X1 U13206 ( .A1(n13151), .A2(n13391), .ZN(n13143) );
  NAND2_X1 U13207 ( .A1(n13150), .A2(n13152), .ZN(n13391) );
  NAND2_X1 U13208 ( .A1(n13392), .A2(n13393), .ZN(n13152) );
  NAND2_X1 U13209 ( .A1(b_19_), .A2(a_4_), .ZN(n13392) );
  XNOR2_X1 U13210 ( .A(n13394), .B(n13395), .ZN(n13150) );
  XOR2_X1 U13211 ( .A(n13396), .B(n13397), .Z(n13394) );
  NAND2_X1 U13212 ( .A1(n13398), .A2(a_4_), .ZN(n13151) );
  INV_X1 U13213 ( .A(n13393), .ZN(n13398) );
  NAND2_X1 U13214 ( .A1(n13399), .A2(n13400), .ZN(n13393) );
  NAND2_X1 U13215 ( .A1(n13157), .A2(n13401), .ZN(n13400) );
  NAND2_X1 U13216 ( .A1(n13160), .A2(n13159), .ZN(n13401) );
  XOR2_X1 U13217 ( .A(n13402), .B(n13403), .Z(n13157) );
  XNOR2_X1 U13218 ( .A(n13404), .B(n13405), .ZN(n13403) );
  INV_X1 U13219 ( .A(n13406), .ZN(n13399) );
  NOR2_X1 U13220 ( .A1(n13159), .A2(n13160), .ZN(n13406) );
  NOR2_X1 U13221 ( .A1(n10056), .A2(n10083), .ZN(n13160) );
  NAND2_X1 U13222 ( .A1(n13167), .A2(n13407), .ZN(n13159) );
  NAND2_X1 U13223 ( .A1(n13166), .A2(n13168), .ZN(n13407) );
  NAND2_X1 U13224 ( .A1(n13408), .A2(n13409), .ZN(n13168) );
  NAND2_X1 U13225 ( .A1(b_19_), .A2(a_6_), .ZN(n13408) );
  XOR2_X1 U13226 ( .A(n13410), .B(n13411), .Z(n13166) );
  XNOR2_X1 U13227 ( .A(n13412), .B(n13413), .ZN(n13411) );
  NAND2_X1 U13228 ( .A1(n13414), .A2(a_6_), .ZN(n13167) );
  INV_X1 U13229 ( .A(n13409), .ZN(n13414) );
  NAND2_X1 U13230 ( .A1(n13415), .A2(n13416), .ZN(n13409) );
  NAND2_X1 U13231 ( .A1(n13173), .A2(n13417), .ZN(n13416) );
  NAND2_X1 U13232 ( .A1(n13176), .A2(n13175), .ZN(n13417) );
  XOR2_X1 U13233 ( .A(n13418), .B(n13419), .Z(n13173) );
  XNOR2_X1 U13234 ( .A(n13420), .B(n13421), .ZN(n13419) );
  INV_X1 U13235 ( .A(n13422), .ZN(n13415) );
  NOR2_X1 U13236 ( .A1(n13175), .A2(n13176), .ZN(n13422) );
  NOR2_X1 U13237 ( .A1(n10056), .A2(n9773), .ZN(n13176) );
  NAND2_X1 U13238 ( .A1(n13363), .A2(n13423), .ZN(n13175) );
  NAND2_X1 U13239 ( .A1(n13362), .A2(n13364), .ZN(n13423) );
  NAND2_X1 U13240 ( .A1(n13424), .A2(n13425), .ZN(n13364) );
  NAND2_X1 U13241 ( .A1(b_19_), .A2(a_8_), .ZN(n13424) );
  XNOR2_X1 U13242 ( .A(n13426), .B(n13427), .ZN(n13362) );
  XOR2_X1 U13243 ( .A(n13428), .B(n13429), .Z(n13426) );
  NAND2_X1 U13244 ( .A1(n13430), .A2(a_8_), .ZN(n13363) );
  INV_X1 U13245 ( .A(n13425), .ZN(n13430) );
  NAND2_X1 U13246 ( .A1(n13431), .A2(n13432), .ZN(n13425) );
  NAND2_X1 U13247 ( .A1(n13185), .A2(n13433), .ZN(n13432) );
  NAND2_X1 U13248 ( .A1(n13188), .A2(n13187), .ZN(n13433) );
  XOR2_X1 U13249 ( .A(n13434), .B(n13435), .Z(n13185) );
  XNOR2_X1 U13250 ( .A(n13436), .B(n13437), .ZN(n13434) );
  INV_X1 U13251 ( .A(n13438), .ZN(n13431) );
  NOR2_X1 U13252 ( .A1(n13187), .A2(n13188), .ZN(n13438) );
  NOR2_X1 U13253 ( .A1(n10056), .A2(n10076), .ZN(n13188) );
  NAND2_X1 U13254 ( .A1(n13439), .A2(n13440), .ZN(n13187) );
  NAND2_X1 U13255 ( .A1(n13441), .A2(b_19_), .ZN(n13440) );
  NOR2_X1 U13256 ( .A1(n13442), .A2(n10073), .ZN(n13441) );
  NOR2_X1 U13257 ( .A1(n13358), .A2(n13359), .ZN(n13442) );
  NAND2_X1 U13258 ( .A1(n13358), .A2(n13359), .ZN(n13439) );
  NAND2_X1 U13259 ( .A1(n13443), .A2(n13444), .ZN(n13359) );
  INV_X1 U13260 ( .A(n13445), .ZN(n13444) );
  NOR2_X1 U13261 ( .A1(n13355), .A2(n13446), .ZN(n13445) );
  NOR2_X1 U13262 ( .A1(n13356), .A2(n13354), .ZN(n13446) );
  NAND2_X1 U13263 ( .A1(b_19_), .A2(a_11_), .ZN(n13355) );
  NAND2_X1 U13264 ( .A1(n13354), .A2(n13356), .ZN(n13443) );
  NAND2_X1 U13265 ( .A1(n13447), .A2(n13448), .ZN(n13356) );
  NAND2_X1 U13266 ( .A1(n13352), .A2(n13449), .ZN(n13448) );
  INV_X1 U13267 ( .A(n13450), .ZN(n13449) );
  NOR2_X1 U13268 ( .A1(n13351), .A2(n13350), .ZN(n13450) );
  NOR2_X1 U13269 ( .A1(n10056), .A2(n10070), .ZN(n13352) );
  NAND2_X1 U13270 ( .A1(n13350), .A2(n13351), .ZN(n13447) );
  NAND2_X1 U13271 ( .A1(n13347), .A2(n13451), .ZN(n13351) );
  NAND2_X1 U13272 ( .A1(n13346), .A2(n13348), .ZN(n13451) );
  NAND2_X1 U13273 ( .A1(n13452), .A2(n13453), .ZN(n13348) );
  NAND2_X1 U13274 ( .A1(b_19_), .A2(a_13_), .ZN(n13453) );
  INV_X1 U13275 ( .A(n13454), .ZN(n13452) );
  XNOR2_X1 U13276 ( .A(n13455), .B(n13456), .ZN(n13346) );
  XOR2_X1 U13277 ( .A(n13457), .B(n13458), .Z(n13456) );
  NAND2_X1 U13278 ( .A1(b_18_), .A2(a_14_), .ZN(n13458) );
  NAND2_X1 U13279 ( .A1(a_13_), .A2(n13454), .ZN(n13347) );
  NAND2_X1 U13280 ( .A1(n13459), .A2(n13460), .ZN(n13454) );
  NAND2_X1 U13281 ( .A1(n13461), .A2(b_19_), .ZN(n13460) );
  NOR2_X1 U13282 ( .A1(n13462), .A2(n10065), .ZN(n13461) );
  NOR2_X1 U13283 ( .A1(n13209), .A2(n13210), .ZN(n13462) );
  NAND2_X1 U13284 ( .A1(n13209), .A2(n13210), .ZN(n13459) );
  NAND2_X1 U13285 ( .A1(n13463), .A2(n13464), .ZN(n13210) );
  NAND2_X1 U13286 ( .A1(n13465), .A2(b_19_), .ZN(n13464) );
  NOR2_X1 U13287 ( .A1(n13466), .A2(n9534), .ZN(n13465) );
  NOR2_X1 U13288 ( .A1(n13217), .A2(n13218), .ZN(n13466) );
  NAND2_X1 U13289 ( .A1(n13217), .A2(n13218), .ZN(n13463) );
  NAND2_X1 U13290 ( .A1(n13227), .A2(n13467), .ZN(n13218) );
  NAND2_X1 U13291 ( .A1(n13226), .A2(n13228), .ZN(n13467) );
  NAND2_X1 U13292 ( .A1(n13468), .A2(n13469), .ZN(n13228) );
  NAND2_X1 U13293 ( .A1(b_19_), .A2(a_16_), .ZN(n13469) );
  INV_X1 U13294 ( .A(n13470), .ZN(n13468) );
  XNOR2_X1 U13295 ( .A(n13471), .B(n13472), .ZN(n13226) );
  NAND2_X1 U13296 ( .A1(n13473), .A2(n13474), .ZN(n13471) );
  NAND2_X1 U13297 ( .A1(a_16_), .A2(n13470), .ZN(n13227) );
  NAND2_X1 U13298 ( .A1(n13235), .A2(n13475), .ZN(n13470) );
  NAND2_X1 U13299 ( .A1(n13234), .A2(n13236), .ZN(n13475) );
  NAND2_X1 U13300 ( .A1(n13476), .A2(n13477), .ZN(n13236) );
  NAND2_X1 U13301 ( .A1(b_19_), .A2(a_17_), .ZN(n13477) );
  INV_X1 U13302 ( .A(n13478), .ZN(n13476) );
  XNOR2_X1 U13303 ( .A(n13479), .B(n13480), .ZN(n13234) );
  XNOR2_X1 U13304 ( .A(n13481), .B(n9450), .ZN(n13479) );
  NAND2_X1 U13305 ( .A1(a_17_), .A2(n13478), .ZN(n13235) );
  NAND2_X1 U13306 ( .A1(n13482), .A2(n13483), .ZN(n13478) );
  NAND2_X1 U13307 ( .A1(n13243), .A2(n13484), .ZN(n13483) );
  NAND2_X1 U13308 ( .A1(n13241), .A2(n13242), .ZN(n13484) );
  NOR2_X1 U13309 ( .A1(n10056), .A2(n10058), .ZN(n13243) );
  INV_X1 U13310 ( .A(n13485), .ZN(n13482) );
  NOR2_X1 U13311 ( .A1(n13242), .A2(n13241), .ZN(n13485) );
  XOR2_X1 U13312 ( .A(n13486), .B(n13487), .Z(n13241) );
  NAND2_X1 U13313 ( .A1(n13488), .A2(n13489), .ZN(n13486) );
  NAND2_X1 U13314 ( .A1(n13490), .A2(n13491), .ZN(n13242) );
  NAND2_X1 U13315 ( .A1(n13248), .A2(n13492), .ZN(n13491) );
  INV_X1 U13316 ( .A(n13493), .ZN(n13492) );
  NOR2_X1 U13317 ( .A1(n13250), .A2(n10009), .ZN(n13493) );
  XNOR2_X1 U13318 ( .A(n13494), .B(n13495), .ZN(n13248) );
  XOR2_X1 U13319 ( .A(n13496), .B(n13497), .Z(n13494) );
  NOR2_X1 U13320 ( .A1(n10054), .A2(n10057), .ZN(n13497) );
  NAND2_X1 U13321 ( .A1(n10009), .A2(n13250), .ZN(n13490) );
  NAND2_X1 U13322 ( .A1(n13498), .A2(n13499), .ZN(n13250) );
  NAND2_X1 U13323 ( .A1(n13341), .A2(n13500), .ZN(n13499) );
  NAND2_X1 U13324 ( .A1(n13344), .A2(n13343), .ZN(n13500) );
  XOR2_X1 U13325 ( .A(n13501), .B(n13502), .Z(n13341) );
  NAND2_X1 U13326 ( .A1(n13503), .A2(n13504), .ZN(n13501) );
  INV_X1 U13327 ( .A(n13505), .ZN(n13498) );
  NOR2_X1 U13328 ( .A1(n13343), .A2(n13344), .ZN(n13505) );
  NOR2_X1 U13329 ( .A1(n10056), .A2(n10054), .ZN(n13344) );
  NAND2_X1 U13330 ( .A1(n13262), .A2(n13506), .ZN(n13343) );
  NAND2_X1 U13331 ( .A1(n13261), .A2(n13263), .ZN(n13506) );
  NAND2_X1 U13332 ( .A1(n13507), .A2(n13508), .ZN(n13263) );
  NAND2_X1 U13333 ( .A1(b_19_), .A2(a_21_), .ZN(n13508) );
  INV_X1 U13334 ( .A(n13509), .ZN(n13507) );
  XNOR2_X1 U13335 ( .A(n13510), .B(n13511), .ZN(n13261) );
  NAND2_X1 U13336 ( .A1(n13512), .A2(n13513), .ZN(n13510) );
  NAND2_X1 U13337 ( .A1(a_21_), .A2(n13509), .ZN(n13262) );
  NAND2_X1 U13338 ( .A1(n13270), .A2(n13514), .ZN(n13509) );
  NAND2_X1 U13339 ( .A1(n13269), .A2(n13271), .ZN(n13514) );
  NAND2_X1 U13340 ( .A1(n13515), .A2(n13516), .ZN(n13271) );
  NAND2_X1 U13341 ( .A1(b_19_), .A2(a_22_), .ZN(n13516) );
  INV_X1 U13342 ( .A(n13517), .ZN(n13515) );
  XOR2_X1 U13343 ( .A(n13518), .B(n13519), .Z(n13269) );
  XOR2_X1 U13344 ( .A(n13520), .B(n13521), .Z(n13518) );
  NOR2_X1 U13345 ( .A1(n10051), .A2(n10057), .ZN(n13521) );
  NAND2_X1 U13346 ( .A1(a_22_), .A2(n13517), .ZN(n13270) );
  NAND2_X1 U13347 ( .A1(n13522), .A2(n13523), .ZN(n13517) );
  NAND2_X1 U13348 ( .A1(n13524), .A2(b_19_), .ZN(n13523) );
  NOR2_X1 U13349 ( .A1(n13525), .A2(n10051), .ZN(n13524) );
  NOR2_X1 U13350 ( .A1(n13277), .A2(n13278), .ZN(n13525) );
  NAND2_X1 U13351 ( .A1(n13277), .A2(n13278), .ZN(n13522) );
  NAND2_X1 U13352 ( .A1(n13526), .A2(n13527), .ZN(n13278) );
  INV_X1 U13353 ( .A(n13528), .ZN(n13527) );
  NOR2_X1 U13354 ( .A1(n13529), .A2(n13530), .ZN(n13528) );
  NOR2_X1 U13355 ( .A1(n13339), .A2(n13337), .ZN(n13530) );
  INV_X1 U13356 ( .A(n13340), .ZN(n13529) );
  NOR2_X1 U13357 ( .A1(n10056), .A2(n10050), .ZN(n13340) );
  NAND2_X1 U13358 ( .A1(n13337), .A2(n13339), .ZN(n13526) );
  NAND2_X1 U13359 ( .A1(n13531), .A2(n13532), .ZN(n13339) );
  NAND2_X1 U13360 ( .A1(n13336), .A2(n13533), .ZN(n13532) );
  NAND2_X1 U13361 ( .A1(n13333), .A2(n13335), .ZN(n13533) );
  NOR2_X1 U13362 ( .A1(n10056), .A2(n10048), .ZN(n13336) );
  INV_X1 U13363 ( .A(n13534), .ZN(n13531) );
  NOR2_X1 U13364 ( .A1(n13335), .A2(n13333), .ZN(n13534) );
  XNOR2_X1 U13365 ( .A(n13535), .B(n13536), .ZN(n13333) );
  XNOR2_X1 U13366 ( .A(n13537), .B(n13538), .ZN(n13536) );
  NAND2_X1 U13367 ( .A1(n13539), .A2(n13540), .ZN(n13335) );
  NAND2_X1 U13368 ( .A1(n13293), .A2(n13541), .ZN(n13540) );
  NAND2_X1 U13369 ( .A1(n13296), .A2(n13295), .ZN(n13541) );
  XOR2_X1 U13370 ( .A(n13542), .B(n13543), .Z(n13293) );
  NAND2_X1 U13371 ( .A1(n13544), .A2(n13545), .ZN(n13542) );
  INV_X1 U13372 ( .A(n13546), .ZN(n13539) );
  NOR2_X1 U13373 ( .A1(n13295), .A2(n13296), .ZN(n13546) );
  NOR2_X1 U13374 ( .A1(n10056), .A2(n10047), .ZN(n13296) );
  NAND2_X1 U13375 ( .A1(n13302), .A2(n13547), .ZN(n13295) );
  NAND2_X1 U13376 ( .A1(n13301), .A2(n13303), .ZN(n13547) );
  NAND2_X1 U13377 ( .A1(n13548), .A2(n13549), .ZN(n13303) );
  NAND2_X1 U13378 ( .A1(b_19_), .A2(a_27_), .ZN(n13549) );
  INV_X1 U13379 ( .A(n13550), .ZN(n13548) );
  XNOR2_X1 U13380 ( .A(n13551), .B(n13552), .ZN(n13301) );
  XOR2_X1 U13381 ( .A(n13553), .B(n13554), .Z(n13552) );
  NAND2_X1 U13382 ( .A1(b_18_), .A2(a_28_), .ZN(n13554) );
  NAND2_X1 U13383 ( .A1(a_27_), .A2(n13550), .ZN(n13302) );
  NAND2_X1 U13384 ( .A1(n13555), .A2(n13556), .ZN(n13550) );
  NAND2_X1 U13385 ( .A1(n13557), .A2(b_19_), .ZN(n13556) );
  NOR2_X1 U13386 ( .A1(n13558), .A2(n9136), .ZN(n13557) );
  NOR2_X1 U13387 ( .A1(n13309), .A2(n13311), .ZN(n13558) );
  NAND2_X1 U13388 ( .A1(n13309), .A2(n13311), .ZN(n13555) );
  NAND2_X1 U13389 ( .A1(n13559), .A2(n13560), .ZN(n13311) );
  NAND2_X1 U13390 ( .A1(n13561), .A2(b_19_), .ZN(n13560) );
  NOR2_X1 U13391 ( .A1(n13562), .A2(n9121), .ZN(n13561) );
  NOR2_X1 U13392 ( .A1(n13563), .A2(n13331), .ZN(n13562) );
  NAND2_X1 U13393 ( .A1(n13563), .A2(n13331), .ZN(n13559) );
  NAND2_X1 U13394 ( .A1(n13564), .A2(n13565), .ZN(n13331) );
  NAND2_X1 U13395 ( .A1(b_17_), .A2(n13566), .ZN(n13565) );
  NAND2_X1 U13396 ( .A1(n10486), .A2(n13567), .ZN(n13566) );
  NAND2_X1 U13397 ( .A1(a_31_), .A2(n10057), .ZN(n13567) );
  NAND2_X1 U13398 ( .A1(b_18_), .A2(n13568), .ZN(n13564) );
  NAND2_X1 U13399 ( .A1(n10489), .A2(n13569), .ZN(n13568) );
  NAND2_X1 U13400 ( .A1(a_30_), .A2(n10059), .ZN(n13569) );
  INV_X1 U13401 ( .A(n13332), .ZN(n13563) );
  NAND2_X1 U13402 ( .A1(n13570), .A2(n9025), .ZN(n13332) );
  NOR2_X1 U13403 ( .A1(n10056), .A2(n10057), .ZN(n13570) );
  XOR2_X1 U13404 ( .A(n13571), .B(n13572), .Z(n13309) );
  NOR2_X1 U13405 ( .A1(n9121), .A2(n10057), .ZN(n13572) );
  XNOR2_X1 U13406 ( .A(n13573), .B(n13574), .ZN(n13571) );
  XNOR2_X1 U13407 ( .A(n13575), .B(n13576), .ZN(n13337) );
  XNOR2_X1 U13408 ( .A(n13577), .B(n13578), .ZN(n13576) );
  XNOR2_X1 U13409 ( .A(n13579), .B(n13580), .ZN(n13277) );
  XNOR2_X1 U13410 ( .A(n13581), .B(n13582), .ZN(n13580) );
  NAND2_X1 U13411 ( .A1(b_19_), .A2(a_19_), .ZN(n10009) );
  XNOR2_X1 U13412 ( .A(n13583), .B(n13584), .ZN(n13217) );
  NAND2_X1 U13413 ( .A1(n13585), .A2(n13586), .ZN(n13583) );
  XNOR2_X1 U13414 ( .A(n13587), .B(n13588), .ZN(n13209) );
  XOR2_X1 U13415 ( .A(n13589), .B(n13590), .Z(n13588) );
  NAND2_X1 U13416 ( .A1(b_18_), .A2(a_15_), .ZN(n13590) );
  XNOR2_X1 U13417 ( .A(n13591), .B(n13592), .ZN(n13350) );
  NAND2_X1 U13418 ( .A1(n13593), .A2(n13594), .ZN(n13591) );
  XOR2_X1 U13419 ( .A(n13595), .B(n13596), .Z(n13354) );
  XOR2_X1 U13420 ( .A(n13597), .B(n13598), .Z(n13595) );
  NOR2_X1 U13421 ( .A1(n10070), .A2(n10057), .ZN(n13598) );
  XOR2_X1 U13422 ( .A(n13599), .B(n13600), .Z(n13358) );
  XNOR2_X1 U13423 ( .A(n13601), .B(n13602), .ZN(n13600) );
  XOR2_X1 U13424 ( .A(n13603), .B(n13604), .Z(n13113) );
  XOR2_X1 U13425 ( .A(n13605), .B(n13606), .Z(n13603) );
  NAND2_X1 U13426 ( .A1(n10198), .A2(n10197), .ZN(n10196) );
  NOR2_X1 U13427 ( .A1(n13607), .A2(n10274), .ZN(n10197) );
  NOR2_X1 U13428 ( .A1(n13608), .A2(n13609), .ZN(n13607) );
  XNOR2_X1 U13429 ( .A(n13610), .B(n13611), .ZN(n13609) );
  NOR2_X1 U13430 ( .A1(n10280), .A2(n10281), .ZN(n10198) );
  XNOR2_X1 U13431 ( .A(n13612), .B(n13613), .ZN(n10281) );
  XNOR2_X1 U13432 ( .A(n13614), .B(n13615), .ZN(n13613) );
  NAND2_X1 U13433 ( .A1(a_0_), .A2(b_17_), .ZN(n13615) );
  INV_X1 U13434 ( .A(n13616), .ZN(n10280) );
  NAND2_X1 U13435 ( .A1(n13617), .A2(n13618), .ZN(n13616) );
  NAND2_X1 U13436 ( .A1(n13117), .A2(n13619), .ZN(n13618) );
  INV_X1 U13437 ( .A(n13620), .ZN(n13619) );
  NOR2_X1 U13438 ( .A1(n13115), .A2(n13116), .ZN(n13620) );
  NOR2_X1 U13439 ( .A1(n10057), .A2(n10093), .ZN(n13117) );
  NAND2_X1 U13440 ( .A1(n13115), .A2(n13116), .ZN(n13617) );
  NAND2_X1 U13441 ( .A1(n13621), .A2(n13622), .ZN(n13116) );
  NAND2_X1 U13442 ( .A1(n13606), .A2(n13623), .ZN(n13622) );
  INV_X1 U13443 ( .A(n13624), .ZN(n13623) );
  NOR2_X1 U13444 ( .A1(n13604), .A2(n13605), .ZN(n13624) );
  NOR2_X1 U13445 ( .A1(n10057), .A2(n9983), .ZN(n13606) );
  NAND2_X1 U13446 ( .A1(n13604), .A2(n13605), .ZN(n13621) );
  NAND2_X1 U13447 ( .A1(n13625), .A2(n13626), .ZN(n13605) );
  NAND2_X1 U13448 ( .A1(n13374), .A2(n13627), .ZN(n13626) );
  INV_X1 U13449 ( .A(n13628), .ZN(n13627) );
  NOR2_X1 U13450 ( .A1(n13371), .A2(n13373), .ZN(n13628) );
  NOR2_X1 U13451 ( .A1(n10057), .A2(n10088), .ZN(n13374) );
  NAND2_X1 U13452 ( .A1(n13371), .A2(n13373), .ZN(n13625) );
  NOR2_X1 U13453 ( .A1(n13629), .A2(n13630), .ZN(n13373) );
  INV_X1 U13454 ( .A(n13631), .ZN(n13630) );
  NAND2_X1 U13455 ( .A1(n13380), .A2(n13632), .ZN(n13631) );
  NAND2_X1 U13456 ( .A1(n13382), .A2(n13381), .ZN(n13632) );
  XOR2_X1 U13457 ( .A(n13633), .B(n13634), .Z(n13380) );
  XNOR2_X1 U13458 ( .A(n13635), .B(n13636), .ZN(n13633) );
  NOR2_X1 U13459 ( .A1(n10059), .A2(n10085), .ZN(n13636) );
  NOR2_X1 U13460 ( .A1(n13381), .A2(n13382), .ZN(n13629) );
  NOR2_X1 U13461 ( .A1(n10057), .A2(n10086), .ZN(n13382) );
  NAND2_X1 U13462 ( .A1(n13637), .A2(n13638), .ZN(n13381) );
  NAND2_X1 U13463 ( .A1(n13390), .A2(n13639), .ZN(n13638) );
  INV_X1 U13464 ( .A(n13640), .ZN(n13639) );
  NOR2_X1 U13465 ( .A1(n13388), .A2(n13389), .ZN(n13640) );
  NOR2_X1 U13466 ( .A1(n10057), .A2(n10085), .ZN(n13390) );
  NAND2_X1 U13467 ( .A1(n13389), .A2(n13388), .ZN(n13637) );
  XOR2_X1 U13468 ( .A(n13641), .B(n13642), .Z(n13388) );
  XNOR2_X1 U13469 ( .A(n13643), .B(n13644), .ZN(n13642) );
  NOR2_X1 U13470 ( .A1(n13645), .A2(n13646), .ZN(n13389) );
  INV_X1 U13471 ( .A(n13647), .ZN(n13646) );
  NAND2_X1 U13472 ( .A1(n13395), .A2(n13648), .ZN(n13647) );
  NAND2_X1 U13473 ( .A1(n13397), .A2(n13396), .ZN(n13648) );
  XNOR2_X1 U13474 ( .A(n13649), .B(n13650), .ZN(n13395) );
  XOR2_X1 U13475 ( .A(n13651), .B(n13652), .Z(n13649) );
  NOR2_X1 U13476 ( .A1(n10059), .A2(n10081), .ZN(n13652) );
  NOR2_X1 U13477 ( .A1(n13396), .A2(n13397), .ZN(n13645) );
  NOR2_X1 U13478 ( .A1(n10057), .A2(n10083), .ZN(n13397) );
  NAND2_X1 U13479 ( .A1(n13653), .A2(n13654), .ZN(n13396) );
  NAND2_X1 U13480 ( .A1(n13405), .A2(n13655), .ZN(n13654) );
  NAND2_X1 U13481 ( .A1(n13402), .A2(n13404), .ZN(n13655) );
  NOR2_X1 U13482 ( .A1(n10057), .A2(n10081), .ZN(n13405) );
  INV_X1 U13483 ( .A(n13656), .ZN(n13653) );
  NOR2_X1 U13484 ( .A1(n13404), .A2(n13402), .ZN(n13656) );
  XOR2_X1 U13485 ( .A(n13657), .B(n13658), .Z(n13402) );
  NAND2_X1 U13486 ( .A1(n13659), .A2(n13660), .ZN(n13657) );
  NAND2_X1 U13487 ( .A1(n13661), .A2(n13662), .ZN(n13404) );
  NAND2_X1 U13488 ( .A1(n13410), .A2(n13663), .ZN(n13662) );
  NAND2_X1 U13489 ( .A1(n13413), .A2(n13412), .ZN(n13663) );
  XNOR2_X1 U13490 ( .A(n13664), .B(n13665), .ZN(n13410) );
  XNOR2_X1 U13491 ( .A(n13666), .B(n13667), .ZN(n13665) );
  INV_X1 U13492 ( .A(n13668), .ZN(n13661) );
  NOR2_X1 U13493 ( .A1(n13412), .A2(n13413), .ZN(n13668) );
  NOR2_X1 U13494 ( .A1(n10057), .A2(n9773), .ZN(n13413) );
  NAND2_X1 U13495 ( .A1(n13669), .A2(n13670), .ZN(n13412) );
  NAND2_X1 U13496 ( .A1(n13421), .A2(n13671), .ZN(n13670) );
  NAND2_X1 U13497 ( .A1(n13418), .A2(n13420), .ZN(n13671) );
  NOR2_X1 U13498 ( .A1(n10057), .A2(n10079), .ZN(n13421) );
  INV_X1 U13499 ( .A(n13672), .ZN(n13669) );
  NOR2_X1 U13500 ( .A1(n13420), .A2(n13418), .ZN(n13672) );
  XOR2_X1 U13501 ( .A(n13673), .B(n13674), .Z(n13418) );
  NAND2_X1 U13502 ( .A1(n13675), .A2(n13676), .ZN(n13673) );
  NAND2_X1 U13503 ( .A1(n13677), .A2(n13678), .ZN(n13420) );
  NAND2_X1 U13504 ( .A1(n13427), .A2(n13679), .ZN(n13678) );
  NAND2_X1 U13505 ( .A1(n13429), .A2(n13428), .ZN(n13679) );
  XNOR2_X1 U13506 ( .A(n13680), .B(n13681), .ZN(n13427) );
  XNOR2_X1 U13507 ( .A(n13682), .B(n13683), .ZN(n13681) );
  INV_X1 U13508 ( .A(n13684), .ZN(n13677) );
  NOR2_X1 U13509 ( .A1(n13428), .A2(n13429), .ZN(n13684) );
  NOR2_X1 U13510 ( .A1(n10057), .A2(n10076), .ZN(n13429) );
  NAND2_X1 U13511 ( .A1(n13685), .A2(n13686), .ZN(n13428) );
  NAND2_X1 U13512 ( .A1(n13437), .A2(n13687), .ZN(n13686) );
  INV_X1 U13513 ( .A(n13688), .ZN(n13687) );
  NOR2_X1 U13514 ( .A1(n13435), .A2(n13436), .ZN(n13688) );
  NOR2_X1 U13515 ( .A1(n10057), .A2(n10073), .ZN(n13437) );
  NAND2_X1 U13516 ( .A1(n13436), .A2(n13435), .ZN(n13685) );
  XNOR2_X1 U13517 ( .A(n13689), .B(n13690), .ZN(n13435) );
  XNOR2_X1 U13518 ( .A(n13691), .B(n13692), .ZN(n13689) );
  NOR2_X1 U13519 ( .A1(n10059), .A2(n9649), .ZN(n13692) );
  NOR2_X1 U13520 ( .A1(n13693), .A2(n13694), .ZN(n13436) );
  INV_X1 U13521 ( .A(n13695), .ZN(n13694) );
  NAND2_X1 U13522 ( .A1(n13599), .A2(n13696), .ZN(n13695) );
  NAND2_X1 U13523 ( .A1(n13602), .A2(n13601), .ZN(n13696) );
  XOR2_X1 U13524 ( .A(n13697), .B(n13698), .Z(n13599) );
  XOR2_X1 U13525 ( .A(n13699), .B(n13700), .Z(n13697) );
  NOR2_X1 U13526 ( .A1(n13601), .A2(n13602), .ZN(n13693) );
  NOR2_X1 U13527 ( .A1(n10057), .A2(n9649), .ZN(n13602) );
  NAND2_X1 U13528 ( .A1(n13701), .A2(n13702), .ZN(n13601) );
  NAND2_X1 U13529 ( .A1(n13703), .A2(b_18_), .ZN(n13702) );
  NOR2_X1 U13530 ( .A1(n13704), .A2(n10070), .ZN(n13703) );
  NOR2_X1 U13531 ( .A1(n13596), .A2(n13597), .ZN(n13704) );
  NAND2_X1 U13532 ( .A1(n13596), .A2(n13597), .ZN(n13701) );
  NAND2_X1 U13533 ( .A1(n13593), .A2(n13705), .ZN(n13597) );
  NAND2_X1 U13534 ( .A1(n13592), .A2(n13594), .ZN(n13705) );
  NAND2_X1 U13535 ( .A1(n13706), .A2(n13707), .ZN(n13594) );
  NAND2_X1 U13536 ( .A1(b_18_), .A2(a_13_), .ZN(n13707) );
  INV_X1 U13537 ( .A(n13708), .ZN(n13706) );
  XOR2_X1 U13538 ( .A(n13709), .B(n13710), .Z(n13592) );
  XOR2_X1 U13539 ( .A(n13711), .B(n13712), .Z(n13709) );
  NOR2_X1 U13540 ( .A1(n10059), .A2(n10065), .ZN(n13712) );
  NAND2_X1 U13541 ( .A1(a_13_), .A2(n13708), .ZN(n13593) );
  NAND2_X1 U13542 ( .A1(n13713), .A2(n13714), .ZN(n13708) );
  NAND2_X1 U13543 ( .A1(n13715), .A2(b_18_), .ZN(n13714) );
  NOR2_X1 U13544 ( .A1(n13716), .A2(n10065), .ZN(n13715) );
  NOR2_X1 U13545 ( .A1(n13455), .A2(n13457), .ZN(n13716) );
  NAND2_X1 U13546 ( .A1(n13455), .A2(n13457), .ZN(n13713) );
  NAND2_X1 U13547 ( .A1(n13717), .A2(n13718), .ZN(n13457) );
  NAND2_X1 U13548 ( .A1(n13719), .A2(b_18_), .ZN(n13718) );
  NOR2_X1 U13549 ( .A1(n13720), .A2(n9534), .ZN(n13719) );
  NOR2_X1 U13550 ( .A1(n13587), .A2(n13589), .ZN(n13720) );
  NAND2_X1 U13551 ( .A1(n13587), .A2(n13589), .ZN(n13717) );
  NAND2_X1 U13552 ( .A1(n13585), .A2(n13721), .ZN(n13589) );
  NAND2_X1 U13553 ( .A1(n13584), .A2(n13586), .ZN(n13721) );
  NAND2_X1 U13554 ( .A1(n13722), .A2(n13723), .ZN(n13586) );
  NAND2_X1 U13555 ( .A1(b_18_), .A2(a_16_), .ZN(n13723) );
  INV_X1 U13556 ( .A(n13724), .ZN(n13722) );
  XNOR2_X1 U13557 ( .A(n13725), .B(n13726), .ZN(n13584) );
  XNOR2_X1 U13558 ( .A(n13727), .B(n13728), .ZN(n13725) );
  NAND2_X1 U13559 ( .A1(a_16_), .A2(n13724), .ZN(n13585) );
  NAND2_X1 U13560 ( .A1(n13473), .A2(n13729), .ZN(n13724) );
  NAND2_X1 U13561 ( .A1(n13472), .A2(n13474), .ZN(n13729) );
  NAND2_X1 U13562 ( .A1(n13730), .A2(n13731), .ZN(n13474) );
  NAND2_X1 U13563 ( .A1(b_18_), .A2(a_17_), .ZN(n13730) );
  XOR2_X1 U13564 ( .A(n13732), .B(n13733), .Z(n13472) );
  XOR2_X1 U13565 ( .A(n13734), .B(n13735), .Z(n13732) );
  NOR2_X1 U13566 ( .A1(n10058), .A2(n10059), .ZN(n13735) );
  INV_X1 U13567 ( .A(n13736), .ZN(n13473) );
  NOR2_X1 U13568 ( .A1(n13731), .A2(n10060), .ZN(n13736) );
  NAND2_X1 U13569 ( .A1(n13737), .A2(n13738), .ZN(n13731) );
  NAND2_X1 U13570 ( .A1(n13480), .A2(n13739), .ZN(n13738) );
  NAND2_X1 U13571 ( .A1(n13740), .A2(n13481), .ZN(n13739) );
  XOR2_X1 U13572 ( .A(n13741), .B(n13742), .Z(n13480) );
  XNOR2_X1 U13573 ( .A(n13743), .B(n13744), .ZN(n13742) );
  INV_X1 U13574 ( .A(n13745), .ZN(n13737) );
  NOR2_X1 U13575 ( .A1(n13481), .A2(n13740), .ZN(n13745) );
  INV_X1 U13576 ( .A(n9450), .ZN(n13740) );
  NAND2_X1 U13577 ( .A1(b_18_), .A2(a_18_), .ZN(n9450) );
  NAND2_X1 U13578 ( .A1(n13488), .A2(n13746), .ZN(n13481) );
  NAND2_X1 U13579 ( .A1(n13487), .A2(n13489), .ZN(n13746) );
  NAND2_X1 U13580 ( .A1(n13747), .A2(n13748), .ZN(n13489) );
  NAND2_X1 U13581 ( .A1(b_18_), .A2(a_19_), .ZN(n13748) );
  INV_X1 U13582 ( .A(n13749), .ZN(n13747) );
  XNOR2_X1 U13583 ( .A(n13750), .B(n13751), .ZN(n13487) );
  XOR2_X1 U13584 ( .A(n13752), .B(n13753), .Z(n13750) );
  NAND2_X1 U13585 ( .A1(a_19_), .A2(n13749), .ZN(n13488) );
  NAND2_X1 U13586 ( .A1(n13754), .A2(n13755), .ZN(n13749) );
  NAND2_X1 U13587 ( .A1(n13756), .A2(b_18_), .ZN(n13755) );
  NOR2_X1 U13588 ( .A1(n13757), .A2(n10054), .ZN(n13756) );
  NOR2_X1 U13589 ( .A1(n13495), .A2(n13496), .ZN(n13757) );
  NAND2_X1 U13590 ( .A1(n13495), .A2(n13496), .ZN(n13754) );
  NAND2_X1 U13591 ( .A1(n13503), .A2(n13758), .ZN(n13496) );
  NAND2_X1 U13592 ( .A1(n13502), .A2(n13504), .ZN(n13758) );
  NAND2_X1 U13593 ( .A1(n13759), .A2(n13760), .ZN(n13504) );
  NAND2_X1 U13594 ( .A1(b_18_), .A2(a_21_), .ZN(n13760) );
  INV_X1 U13595 ( .A(n13761), .ZN(n13759) );
  XNOR2_X1 U13596 ( .A(n13762), .B(n13763), .ZN(n13502) );
  XOR2_X1 U13597 ( .A(n13764), .B(n13765), .Z(n13763) );
  NAND2_X1 U13598 ( .A1(b_17_), .A2(a_22_), .ZN(n13765) );
  NAND2_X1 U13599 ( .A1(a_21_), .A2(n13761), .ZN(n13503) );
  NAND2_X1 U13600 ( .A1(n13512), .A2(n13766), .ZN(n13761) );
  NAND2_X1 U13601 ( .A1(n13511), .A2(n13513), .ZN(n13766) );
  NAND2_X1 U13602 ( .A1(n13767), .A2(n13768), .ZN(n13513) );
  NAND2_X1 U13603 ( .A1(b_18_), .A2(a_22_), .ZN(n13768) );
  INV_X1 U13604 ( .A(n13769), .ZN(n13767) );
  XOR2_X1 U13605 ( .A(n13770), .B(n13771), .Z(n13511) );
  XOR2_X1 U13606 ( .A(n13772), .B(n13773), .Z(n13770) );
  NOR2_X1 U13607 ( .A1(n10051), .A2(n10059), .ZN(n13773) );
  NAND2_X1 U13608 ( .A1(a_22_), .A2(n13769), .ZN(n13512) );
  NAND2_X1 U13609 ( .A1(n13774), .A2(n13775), .ZN(n13769) );
  NAND2_X1 U13610 ( .A1(n13776), .A2(b_18_), .ZN(n13775) );
  NOR2_X1 U13611 ( .A1(n13777), .A2(n10051), .ZN(n13776) );
  NOR2_X1 U13612 ( .A1(n13520), .A2(n13519), .ZN(n13777) );
  NAND2_X1 U13613 ( .A1(n13519), .A2(n13520), .ZN(n13774) );
  NAND2_X1 U13614 ( .A1(n13778), .A2(n13779), .ZN(n13520) );
  INV_X1 U13615 ( .A(n13780), .ZN(n13779) );
  NOR2_X1 U13616 ( .A1(n13781), .A2(n13782), .ZN(n13780) );
  NOR2_X1 U13617 ( .A1(n13581), .A2(n13579), .ZN(n13782) );
  INV_X1 U13618 ( .A(n13582), .ZN(n13781) );
  NOR2_X1 U13619 ( .A1(n10057), .A2(n10050), .ZN(n13582) );
  NAND2_X1 U13620 ( .A1(n13579), .A2(n13581), .ZN(n13778) );
  NAND2_X1 U13621 ( .A1(n13783), .A2(n13784), .ZN(n13581) );
  NAND2_X1 U13622 ( .A1(n13578), .A2(n13785), .ZN(n13784) );
  NAND2_X1 U13623 ( .A1(n13575), .A2(n13577), .ZN(n13785) );
  NOR2_X1 U13624 ( .A1(n10057), .A2(n10048), .ZN(n13578) );
  INV_X1 U13625 ( .A(n13786), .ZN(n13783) );
  NOR2_X1 U13626 ( .A1(n13575), .A2(n13577), .ZN(n13786) );
  NAND2_X1 U13627 ( .A1(n13787), .A2(n13788), .ZN(n13577) );
  NAND2_X1 U13628 ( .A1(n13535), .A2(n13789), .ZN(n13788) );
  NAND2_X1 U13629 ( .A1(n13538), .A2(n13537), .ZN(n13789) );
  XOR2_X1 U13630 ( .A(n13790), .B(n13791), .Z(n13535) );
  NAND2_X1 U13631 ( .A1(n13792), .A2(n13793), .ZN(n13790) );
  INV_X1 U13632 ( .A(n13794), .ZN(n13787) );
  NOR2_X1 U13633 ( .A1(n13537), .A2(n13538), .ZN(n13794) );
  NOR2_X1 U13634 ( .A1(n10057), .A2(n10047), .ZN(n13538) );
  NAND2_X1 U13635 ( .A1(n13544), .A2(n13795), .ZN(n13537) );
  NAND2_X1 U13636 ( .A1(n13543), .A2(n13545), .ZN(n13795) );
  NAND2_X1 U13637 ( .A1(n13796), .A2(n13797), .ZN(n13545) );
  NAND2_X1 U13638 ( .A1(b_18_), .A2(a_27_), .ZN(n13797) );
  INV_X1 U13639 ( .A(n13798), .ZN(n13796) );
  XNOR2_X1 U13640 ( .A(n13799), .B(n13800), .ZN(n13543) );
  XOR2_X1 U13641 ( .A(n13801), .B(n13802), .Z(n13800) );
  NAND2_X1 U13642 ( .A1(b_17_), .A2(a_28_), .ZN(n13802) );
  NAND2_X1 U13643 ( .A1(a_27_), .A2(n13798), .ZN(n13544) );
  NAND2_X1 U13644 ( .A1(n13803), .A2(n13804), .ZN(n13798) );
  NAND2_X1 U13645 ( .A1(n13805), .A2(b_18_), .ZN(n13804) );
  NOR2_X1 U13646 ( .A1(n13806), .A2(n9136), .ZN(n13805) );
  NOR2_X1 U13647 ( .A1(n13551), .A2(n13553), .ZN(n13806) );
  NAND2_X1 U13648 ( .A1(n13551), .A2(n13553), .ZN(n13803) );
  NAND2_X1 U13649 ( .A1(n13807), .A2(n13808), .ZN(n13553) );
  NAND2_X1 U13650 ( .A1(n13809), .A2(b_18_), .ZN(n13808) );
  NOR2_X1 U13651 ( .A1(n13810), .A2(n9121), .ZN(n13809) );
  NOR2_X1 U13652 ( .A1(n13811), .A2(n13573), .ZN(n13810) );
  NAND2_X1 U13653 ( .A1(n13811), .A2(n13573), .ZN(n13807) );
  NAND2_X1 U13654 ( .A1(n13812), .A2(n13813), .ZN(n13573) );
  NAND2_X1 U13655 ( .A1(b_16_), .A2(n13814), .ZN(n13813) );
  NAND2_X1 U13656 ( .A1(n10486), .A2(n13815), .ZN(n13814) );
  NAND2_X1 U13657 ( .A1(a_31_), .A2(n10059), .ZN(n13815) );
  NAND2_X1 U13658 ( .A1(b_17_), .A2(n13816), .ZN(n13812) );
  NAND2_X1 U13659 ( .A1(n10489), .A2(n13817), .ZN(n13816) );
  NAND2_X1 U13660 ( .A1(a_30_), .A2(n10061), .ZN(n13817) );
  INV_X1 U13661 ( .A(n13574), .ZN(n13811) );
  NAND2_X1 U13662 ( .A1(n13818), .A2(n9025), .ZN(n13574) );
  NOR2_X1 U13663 ( .A1(n10059), .A2(n10057), .ZN(n13818) );
  XOR2_X1 U13664 ( .A(n13819), .B(n13820), .Z(n13551) );
  NOR2_X1 U13665 ( .A1(n9121), .A2(n10059), .ZN(n13820) );
  XNOR2_X1 U13666 ( .A(n13821), .B(n13822), .ZN(n13819) );
  XNOR2_X1 U13667 ( .A(n13823), .B(n13824), .ZN(n13575) );
  XNOR2_X1 U13668 ( .A(n13825), .B(n13826), .ZN(n13824) );
  XNOR2_X1 U13669 ( .A(n13827), .B(n13828), .ZN(n13579) );
  XNOR2_X1 U13670 ( .A(n13829), .B(n13830), .ZN(n13828) );
  XNOR2_X1 U13671 ( .A(n13831), .B(n13832), .ZN(n13519) );
  XNOR2_X1 U13672 ( .A(n13833), .B(n13834), .ZN(n13832) );
  XNOR2_X1 U13673 ( .A(n13835), .B(n13836), .ZN(n13495) );
  NAND2_X1 U13674 ( .A1(n13837), .A2(n13838), .ZN(n13835) );
  XOR2_X1 U13675 ( .A(n13839), .B(n13840), .Z(n13587) );
  XNOR2_X1 U13676 ( .A(n13841), .B(n13842), .ZN(n13839) );
  XOR2_X1 U13677 ( .A(n13843), .B(n13844), .Z(n13455) );
  XNOR2_X1 U13678 ( .A(n13845), .B(n13846), .ZN(n13844) );
  NAND2_X1 U13679 ( .A1(a_15_), .A2(b_17_), .ZN(n13846) );
  XNOR2_X1 U13680 ( .A(n13847), .B(n13848), .ZN(n13596) );
  NAND2_X1 U13681 ( .A1(n13849), .A2(n13850), .ZN(n13847) );
  XOR2_X1 U13682 ( .A(n13851), .B(n13852), .Z(n13371) );
  XNOR2_X1 U13683 ( .A(n13853), .B(n13854), .ZN(n13852) );
  XNOR2_X1 U13684 ( .A(n13855), .B(n13856), .ZN(n13604) );
  XNOR2_X1 U13685 ( .A(n13857), .B(n13858), .ZN(n13855) );
  NOR2_X1 U13686 ( .A1(n10059), .A2(n10088), .ZN(n13858) );
  XOR2_X1 U13687 ( .A(n13859), .B(n13860), .Z(n13115) );
  XNOR2_X1 U13688 ( .A(n13861), .B(n13862), .ZN(n13860) );
  INV_X1 U13689 ( .A(n13863), .ZN(n10204) );
  NOR2_X1 U13690 ( .A1(n10273), .A2(n10274), .ZN(n13863) );
  NOR2_X1 U13691 ( .A1(n13864), .A2(n13865), .ZN(n10274) );
  INV_X1 U13692 ( .A(n13608), .ZN(n13865) );
  NAND2_X1 U13693 ( .A1(n13866), .A2(n13867), .ZN(n13608) );
  NAND2_X1 U13694 ( .A1(n13868), .A2(a_0_), .ZN(n13867) );
  NOR2_X1 U13695 ( .A1(n13869), .A2(n10059), .ZN(n13868) );
  NOR2_X1 U13696 ( .A1(n13614), .A2(n13612), .ZN(n13869) );
  NAND2_X1 U13697 ( .A1(n13614), .A2(n13612), .ZN(n13866) );
  XNOR2_X1 U13698 ( .A(n13870), .B(n13871), .ZN(n13612) );
  NAND2_X1 U13699 ( .A1(n13872), .A2(n13873), .ZN(n13870) );
  NOR2_X1 U13700 ( .A1(n13874), .A2(n13875), .ZN(n13614) );
  INV_X1 U13701 ( .A(n13876), .ZN(n13875) );
  NAND2_X1 U13702 ( .A1(n13859), .A2(n13877), .ZN(n13876) );
  NAND2_X1 U13703 ( .A1(n13862), .A2(n13861), .ZN(n13877) );
  XOR2_X1 U13704 ( .A(n13878), .B(n13879), .Z(n13859) );
  NAND2_X1 U13705 ( .A1(n13880), .A2(n13881), .ZN(n13878) );
  NOR2_X1 U13706 ( .A1(n13861), .A2(n13862), .ZN(n13874) );
  NOR2_X1 U13707 ( .A1(n9983), .A2(n10059), .ZN(n13862) );
  NAND2_X1 U13708 ( .A1(n13882), .A2(n13883), .ZN(n13861) );
  NAND2_X1 U13709 ( .A1(n13884), .A2(a_2_), .ZN(n13883) );
  NOR2_X1 U13710 ( .A1(n13885), .A2(n10059), .ZN(n13884) );
  NOR2_X1 U13711 ( .A1(n13857), .A2(n13856), .ZN(n13885) );
  NAND2_X1 U13712 ( .A1(n13857), .A2(n13856), .ZN(n13882) );
  XNOR2_X1 U13713 ( .A(n13886), .B(n13887), .ZN(n13856) );
  NAND2_X1 U13714 ( .A1(n13888), .A2(n13889), .ZN(n13886) );
  NOR2_X1 U13715 ( .A1(n13890), .A2(n13891), .ZN(n13857) );
  INV_X1 U13716 ( .A(n13892), .ZN(n13891) );
  NAND2_X1 U13717 ( .A1(n13851), .A2(n13893), .ZN(n13892) );
  NAND2_X1 U13718 ( .A1(n13854), .A2(n13853), .ZN(n13893) );
  XOR2_X1 U13719 ( .A(n13894), .B(n13895), .Z(n13851) );
  NAND2_X1 U13720 ( .A1(n13896), .A2(n13897), .ZN(n13894) );
  NOR2_X1 U13721 ( .A1(n13853), .A2(n13854), .ZN(n13890) );
  NOR2_X1 U13722 ( .A1(n10086), .A2(n10059), .ZN(n13854) );
  NAND2_X1 U13723 ( .A1(n13898), .A2(n13899), .ZN(n13853) );
  NAND2_X1 U13724 ( .A1(n13900), .A2(a_4_), .ZN(n13899) );
  NOR2_X1 U13725 ( .A1(n13901), .A2(n10059), .ZN(n13900) );
  NOR2_X1 U13726 ( .A1(n13635), .A2(n13634), .ZN(n13901) );
  NAND2_X1 U13727 ( .A1(n13635), .A2(n13634), .ZN(n13898) );
  XNOR2_X1 U13728 ( .A(n13902), .B(n13903), .ZN(n13634) );
  NAND2_X1 U13729 ( .A1(n13904), .A2(n13905), .ZN(n13902) );
  NOR2_X1 U13730 ( .A1(n13906), .A2(n13907), .ZN(n13635) );
  INV_X1 U13731 ( .A(n13908), .ZN(n13907) );
  NAND2_X1 U13732 ( .A1(n13641), .A2(n13909), .ZN(n13908) );
  NAND2_X1 U13733 ( .A1(n13644), .A2(n13643), .ZN(n13909) );
  XNOR2_X1 U13734 ( .A(n13910), .B(n13911), .ZN(n13641) );
  XOR2_X1 U13735 ( .A(n13912), .B(n13913), .Z(n13910) );
  NOR2_X1 U13736 ( .A1(n10061), .A2(n10081), .ZN(n13913) );
  NOR2_X1 U13737 ( .A1(n13643), .A2(n13644), .ZN(n13906) );
  NOR2_X1 U13738 ( .A1(n10083), .A2(n10059), .ZN(n13644) );
  NAND2_X1 U13739 ( .A1(n13914), .A2(n13915), .ZN(n13643) );
  NAND2_X1 U13740 ( .A1(n13916), .A2(a_6_), .ZN(n13915) );
  NOR2_X1 U13741 ( .A1(n13917), .A2(n10059), .ZN(n13916) );
  NOR2_X1 U13742 ( .A1(n13650), .A2(n13651), .ZN(n13917) );
  NAND2_X1 U13743 ( .A1(n13650), .A2(n13651), .ZN(n13914) );
  NAND2_X1 U13744 ( .A1(n13659), .A2(n13918), .ZN(n13651) );
  NAND2_X1 U13745 ( .A1(n13658), .A2(n13660), .ZN(n13918) );
  NAND2_X1 U13746 ( .A1(n13919), .A2(n13920), .ZN(n13660) );
  NAND2_X1 U13747 ( .A1(a_7_), .A2(b_17_), .ZN(n13919) );
  XOR2_X1 U13748 ( .A(n13921), .B(n13922), .Z(n13658) );
  XNOR2_X1 U13749 ( .A(n13923), .B(n13924), .ZN(n13922) );
  NAND2_X1 U13750 ( .A1(a_8_), .A2(b_16_), .ZN(n13924) );
  NAND2_X1 U13751 ( .A1(n13925), .A2(a_7_), .ZN(n13659) );
  INV_X1 U13752 ( .A(n13920), .ZN(n13925) );
  NAND2_X1 U13753 ( .A1(n13926), .A2(n13927), .ZN(n13920) );
  NAND2_X1 U13754 ( .A1(n13664), .A2(n13928), .ZN(n13927) );
  NAND2_X1 U13755 ( .A1(n13667), .A2(n13666), .ZN(n13928) );
  XNOR2_X1 U13756 ( .A(n13929), .B(n13930), .ZN(n13664) );
  XNOR2_X1 U13757 ( .A(n13931), .B(n13932), .ZN(n13930) );
  INV_X1 U13758 ( .A(n13933), .ZN(n13926) );
  NOR2_X1 U13759 ( .A1(n13666), .A2(n13667), .ZN(n13933) );
  NOR2_X1 U13760 ( .A1(n10079), .A2(n10059), .ZN(n13667) );
  NAND2_X1 U13761 ( .A1(n13675), .A2(n13934), .ZN(n13666) );
  NAND2_X1 U13762 ( .A1(n13674), .A2(n13676), .ZN(n13934) );
  NAND2_X1 U13763 ( .A1(n13935), .A2(n13936), .ZN(n13676) );
  NAND2_X1 U13764 ( .A1(a_9_), .A2(b_17_), .ZN(n13935) );
  XNOR2_X1 U13765 ( .A(n13937), .B(n13938), .ZN(n13674) );
  NAND2_X1 U13766 ( .A1(n13939), .A2(n13940), .ZN(n13937) );
  NAND2_X1 U13767 ( .A1(n13941), .A2(a_9_), .ZN(n13675) );
  INV_X1 U13768 ( .A(n13936), .ZN(n13941) );
  NAND2_X1 U13769 ( .A1(n13942), .A2(n13943), .ZN(n13936) );
  NAND2_X1 U13770 ( .A1(n13680), .A2(n13944), .ZN(n13943) );
  NAND2_X1 U13771 ( .A1(n13683), .A2(n13682), .ZN(n13944) );
  XOR2_X1 U13772 ( .A(n13945), .B(n13946), .Z(n13680) );
  NAND2_X1 U13773 ( .A1(n13947), .A2(n13948), .ZN(n13945) );
  INV_X1 U13774 ( .A(n13949), .ZN(n13942) );
  NOR2_X1 U13775 ( .A1(n13682), .A2(n13683), .ZN(n13949) );
  NOR2_X1 U13776 ( .A1(n10073), .A2(n10059), .ZN(n13683) );
  NAND2_X1 U13777 ( .A1(n13950), .A2(n13951), .ZN(n13682) );
  NAND2_X1 U13778 ( .A1(n13952), .A2(a_11_), .ZN(n13951) );
  NOR2_X1 U13779 ( .A1(n13953), .A2(n10059), .ZN(n13952) );
  NOR2_X1 U13780 ( .A1(n13691), .A2(n13690), .ZN(n13953) );
  NAND2_X1 U13781 ( .A1(n13691), .A2(n13690), .ZN(n13950) );
  XNOR2_X1 U13782 ( .A(n13954), .B(n13955), .ZN(n13690) );
  NAND2_X1 U13783 ( .A1(n13956), .A2(n13957), .ZN(n13954) );
  NOR2_X1 U13784 ( .A1(n13958), .A2(n13959), .ZN(n13691) );
  INV_X1 U13785 ( .A(n13960), .ZN(n13959) );
  NAND2_X1 U13786 ( .A1(n13698), .A2(n13961), .ZN(n13960) );
  NAND2_X1 U13787 ( .A1(n13700), .A2(n13699), .ZN(n13961) );
  XNOR2_X1 U13788 ( .A(n13962), .B(n13963), .ZN(n13698) );
  XOR2_X1 U13789 ( .A(n13964), .B(n13965), .Z(n13962) );
  NOR2_X1 U13790 ( .A1(n10061), .A2(n10067), .ZN(n13965) );
  NOR2_X1 U13791 ( .A1(n13699), .A2(n13700), .ZN(n13958) );
  NOR2_X1 U13792 ( .A1(n10070), .A2(n10059), .ZN(n13700) );
  NAND2_X1 U13793 ( .A1(n13849), .A2(n13966), .ZN(n13699) );
  NAND2_X1 U13794 ( .A1(n13848), .A2(n13850), .ZN(n13966) );
  NAND2_X1 U13795 ( .A1(n13967), .A2(n13968), .ZN(n13850) );
  NAND2_X1 U13796 ( .A1(a_13_), .A2(b_17_), .ZN(n13968) );
  INV_X1 U13797 ( .A(n13969), .ZN(n13967) );
  XOR2_X1 U13798 ( .A(n13970), .B(n13971), .Z(n13848) );
  XNOR2_X1 U13799 ( .A(n13972), .B(n13973), .ZN(n13970) );
  NAND2_X1 U13800 ( .A1(a_14_), .A2(b_16_), .ZN(n13972) );
  NAND2_X1 U13801 ( .A1(a_13_), .A2(n13969), .ZN(n13849) );
  NAND2_X1 U13802 ( .A1(n13974), .A2(n13975), .ZN(n13969) );
  NAND2_X1 U13803 ( .A1(n13976), .A2(a_14_), .ZN(n13975) );
  NOR2_X1 U13804 ( .A1(n13977), .A2(n10059), .ZN(n13976) );
  NOR2_X1 U13805 ( .A1(n13710), .A2(n13711), .ZN(n13977) );
  NAND2_X1 U13806 ( .A1(n13710), .A2(n13711), .ZN(n13974) );
  NAND2_X1 U13807 ( .A1(n13978), .A2(n13979), .ZN(n13711) );
  NAND2_X1 U13808 ( .A1(n13980), .A2(a_15_), .ZN(n13979) );
  NOR2_X1 U13809 ( .A1(n13981), .A2(n10059), .ZN(n13980) );
  NOR2_X1 U13810 ( .A1(n13845), .A2(n13843), .ZN(n13981) );
  NAND2_X1 U13811 ( .A1(n13845), .A2(n13843), .ZN(n13978) );
  XOR2_X1 U13812 ( .A(n13982), .B(n13983), .Z(n13843) );
  XNOR2_X1 U13813 ( .A(n13984), .B(n9512), .ZN(n13982) );
  NOR2_X1 U13814 ( .A1(n13985), .A2(n13986), .ZN(n13845) );
  INV_X1 U13815 ( .A(n13987), .ZN(n13986) );
  NAND2_X1 U13816 ( .A1(n13840), .A2(n13988), .ZN(n13987) );
  NAND2_X1 U13817 ( .A1(n13841), .A2(n13842), .ZN(n13988) );
  XOR2_X1 U13818 ( .A(n13989), .B(n13990), .Z(n13840) );
  NAND2_X1 U13819 ( .A1(n13991), .A2(n13992), .ZN(n13989) );
  NOR2_X1 U13820 ( .A1(n13842), .A2(n13841), .ZN(n13985) );
  INV_X1 U13821 ( .A(n13993), .ZN(n13841) );
  NAND2_X1 U13822 ( .A1(n13994), .A2(n13995), .ZN(n13993) );
  NAND2_X1 U13823 ( .A1(n13726), .A2(n13996), .ZN(n13995) );
  NAND2_X1 U13824 ( .A1(n13727), .A2(n13997), .ZN(n13996) );
  XNOR2_X1 U13825 ( .A(n13998), .B(n13999), .ZN(n13726) );
  XOR2_X1 U13826 ( .A(n14000), .B(n14001), .Z(n13998) );
  NOR2_X1 U13827 ( .A1(n10058), .A2(n10061), .ZN(n14001) );
  NAND2_X1 U13828 ( .A1(n13728), .A2(n9483), .ZN(n13994) );
  INV_X1 U13829 ( .A(n13727), .ZN(n9483) );
  NOR2_X1 U13830 ( .A1(n10059), .A2(n10060), .ZN(n13727) );
  INV_X1 U13831 ( .A(n13997), .ZN(n13728) );
  NAND2_X1 U13832 ( .A1(n14002), .A2(n14003), .ZN(n13997) );
  NAND2_X1 U13833 ( .A1(n14004), .A2(b_17_), .ZN(n14003) );
  NOR2_X1 U13834 ( .A1(n14005), .A2(n10058), .ZN(n14004) );
  NOR2_X1 U13835 ( .A1(n13733), .A2(n13734), .ZN(n14005) );
  NAND2_X1 U13836 ( .A1(n13733), .A2(n13734), .ZN(n14002) );
  NAND2_X1 U13837 ( .A1(n14006), .A2(n14007), .ZN(n13734) );
  NAND2_X1 U13838 ( .A1(n13744), .A2(n14008), .ZN(n14007) );
  NAND2_X1 U13839 ( .A1(n13741), .A2(n13743), .ZN(n14008) );
  NOR2_X1 U13840 ( .A1(n10059), .A2(n9415), .ZN(n13744) );
  INV_X1 U13841 ( .A(n14009), .ZN(n14006) );
  NOR2_X1 U13842 ( .A1(n13743), .A2(n13741), .ZN(n14009) );
  XOR2_X1 U13843 ( .A(n14010), .B(n14011), .Z(n13741) );
  XNOR2_X1 U13844 ( .A(n14012), .B(n14013), .ZN(n14010) );
  NAND2_X1 U13845 ( .A1(n14014), .A2(n14015), .ZN(n13743) );
  NAND2_X1 U13846 ( .A1(n13751), .A2(n14016), .ZN(n14015) );
  NAND2_X1 U13847 ( .A1(n13753), .A2(n13752), .ZN(n14016) );
  XNOR2_X1 U13848 ( .A(n14017), .B(n14018), .ZN(n13751) );
  XOR2_X1 U13849 ( .A(n14019), .B(n14020), .Z(n14017) );
  INV_X1 U13850 ( .A(n14021), .ZN(n14014) );
  NOR2_X1 U13851 ( .A1(n13752), .A2(n13753), .ZN(n14021) );
  NOR2_X1 U13852 ( .A1(n10059), .A2(n10054), .ZN(n13753) );
  NAND2_X1 U13853 ( .A1(n13837), .A2(n14022), .ZN(n13752) );
  NAND2_X1 U13854 ( .A1(n13836), .A2(n13838), .ZN(n14022) );
  NAND2_X1 U13855 ( .A1(n14023), .A2(n14024), .ZN(n13838) );
  NAND2_X1 U13856 ( .A1(b_17_), .A2(a_21_), .ZN(n14024) );
  INV_X1 U13857 ( .A(n14025), .ZN(n14023) );
  XNOR2_X1 U13858 ( .A(n14026), .B(n14027), .ZN(n13836) );
  NAND2_X1 U13859 ( .A1(n14028), .A2(n14029), .ZN(n14026) );
  NAND2_X1 U13860 ( .A1(a_21_), .A2(n14025), .ZN(n13837) );
  NAND2_X1 U13861 ( .A1(n14030), .A2(n14031), .ZN(n14025) );
  NAND2_X1 U13862 ( .A1(n14032), .A2(b_17_), .ZN(n14031) );
  NOR2_X1 U13863 ( .A1(n14033), .A2(n9330), .ZN(n14032) );
  NOR2_X1 U13864 ( .A1(n13762), .A2(n13764), .ZN(n14033) );
  NAND2_X1 U13865 ( .A1(n13762), .A2(n13764), .ZN(n14030) );
  NAND2_X1 U13866 ( .A1(n14034), .A2(n14035), .ZN(n13764) );
  NAND2_X1 U13867 ( .A1(n14036), .A2(b_17_), .ZN(n14035) );
  NOR2_X1 U13868 ( .A1(n14037), .A2(n10051), .ZN(n14036) );
  NOR2_X1 U13869 ( .A1(n13771), .A2(n13772), .ZN(n14037) );
  NAND2_X1 U13870 ( .A1(n13771), .A2(n13772), .ZN(n14034) );
  NAND2_X1 U13871 ( .A1(n14038), .A2(n14039), .ZN(n13772) );
  INV_X1 U13872 ( .A(n14040), .ZN(n14039) );
  NOR2_X1 U13873 ( .A1(n14041), .A2(n14042), .ZN(n14040) );
  NOR2_X1 U13874 ( .A1(n13833), .A2(n13831), .ZN(n14042) );
  INV_X1 U13875 ( .A(n13834), .ZN(n14041) );
  NOR2_X1 U13876 ( .A1(n10059), .A2(n10050), .ZN(n13834) );
  NAND2_X1 U13877 ( .A1(n13831), .A2(n13833), .ZN(n14038) );
  NAND2_X1 U13878 ( .A1(n14043), .A2(n14044), .ZN(n13833) );
  NAND2_X1 U13879 ( .A1(n13830), .A2(n14045), .ZN(n14044) );
  NAND2_X1 U13880 ( .A1(n13827), .A2(n13829), .ZN(n14045) );
  NOR2_X1 U13881 ( .A1(n10059), .A2(n10048), .ZN(n13830) );
  INV_X1 U13882 ( .A(n14046), .ZN(n14043) );
  NOR2_X1 U13883 ( .A1(n13829), .A2(n13827), .ZN(n14046) );
  XNOR2_X1 U13884 ( .A(n14047), .B(n14048), .ZN(n13827) );
  XNOR2_X1 U13885 ( .A(n14049), .B(n14050), .ZN(n14048) );
  NAND2_X1 U13886 ( .A1(n14051), .A2(n14052), .ZN(n13829) );
  NAND2_X1 U13887 ( .A1(n13823), .A2(n14053), .ZN(n14052) );
  NAND2_X1 U13888 ( .A1(n13826), .A2(n13825), .ZN(n14053) );
  XOR2_X1 U13889 ( .A(n14054), .B(n14055), .Z(n13823) );
  NAND2_X1 U13890 ( .A1(n14056), .A2(n14057), .ZN(n14054) );
  INV_X1 U13891 ( .A(n14058), .ZN(n14051) );
  NOR2_X1 U13892 ( .A1(n13825), .A2(n13826), .ZN(n14058) );
  NOR2_X1 U13893 ( .A1(n10059), .A2(n10047), .ZN(n13826) );
  NAND2_X1 U13894 ( .A1(n13792), .A2(n14059), .ZN(n13825) );
  NAND2_X1 U13895 ( .A1(n13791), .A2(n13793), .ZN(n14059) );
  NAND2_X1 U13896 ( .A1(n14060), .A2(n14061), .ZN(n13793) );
  NAND2_X1 U13897 ( .A1(b_17_), .A2(a_27_), .ZN(n14061) );
  INV_X1 U13898 ( .A(n14062), .ZN(n14060) );
  XNOR2_X1 U13899 ( .A(n14063), .B(n14064), .ZN(n13791) );
  XOR2_X1 U13900 ( .A(n14065), .B(n14066), .Z(n14064) );
  NAND2_X1 U13901 ( .A1(b_16_), .A2(a_28_), .ZN(n14066) );
  NAND2_X1 U13902 ( .A1(a_27_), .A2(n14062), .ZN(n13792) );
  NAND2_X1 U13903 ( .A1(n14067), .A2(n14068), .ZN(n14062) );
  NAND2_X1 U13904 ( .A1(n14069), .A2(b_17_), .ZN(n14068) );
  NOR2_X1 U13905 ( .A1(n14070), .A2(n9136), .ZN(n14069) );
  NOR2_X1 U13906 ( .A1(n13799), .A2(n13801), .ZN(n14070) );
  NAND2_X1 U13907 ( .A1(n13799), .A2(n13801), .ZN(n14067) );
  NAND2_X1 U13908 ( .A1(n14071), .A2(n14072), .ZN(n13801) );
  NAND2_X1 U13909 ( .A1(n14073), .A2(b_17_), .ZN(n14072) );
  NOR2_X1 U13910 ( .A1(n14074), .A2(n9121), .ZN(n14073) );
  NOR2_X1 U13911 ( .A1(n14075), .A2(n13821), .ZN(n14074) );
  NAND2_X1 U13912 ( .A1(n14075), .A2(n13821), .ZN(n14071) );
  NAND2_X1 U13913 ( .A1(n14076), .A2(n14077), .ZN(n13821) );
  NAND2_X1 U13914 ( .A1(b_15_), .A2(n14078), .ZN(n14077) );
  NAND2_X1 U13915 ( .A1(n10486), .A2(n14079), .ZN(n14078) );
  NAND2_X1 U13916 ( .A1(a_31_), .A2(n10061), .ZN(n14079) );
  NAND2_X1 U13917 ( .A1(b_16_), .A2(n14080), .ZN(n14076) );
  NAND2_X1 U13918 ( .A1(n10489), .A2(n14081), .ZN(n14080) );
  NAND2_X1 U13919 ( .A1(a_30_), .A2(n10063), .ZN(n14081) );
  INV_X1 U13920 ( .A(n13822), .ZN(n14075) );
  NAND2_X1 U13921 ( .A1(n14082), .A2(n9025), .ZN(n13822) );
  NOR2_X1 U13922 ( .A1(n10059), .A2(n10061), .ZN(n14082) );
  XOR2_X1 U13923 ( .A(n14083), .B(n14084), .Z(n13799) );
  NOR2_X1 U13924 ( .A1(n9121), .A2(n10061), .ZN(n14084) );
  XNOR2_X1 U13925 ( .A(n14085), .B(n14086), .ZN(n14083) );
  XNOR2_X1 U13926 ( .A(n14087), .B(n14088), .ZN(n13831) );
  XNOR2_X1 U13927 ( .A(n14089), .B(n14090), .ZN(n14088) );
  XNOR2_X1 U13928 ( .A(n14091), .B(n14092), .ZN(n13771) );
  XOR2_X1 U13929 ( .A(n14093), .B(n14094), .Z(n14092) );
  XNOR2_X1 U13930 ( .A(n14095), .B(n14096), .ZN(n13762) );
  NAND2_X1 U13931 ( .A1(n14097), .A2(n14098), .ZN(n14095) );
  XOR2_X1 U13932 ( .A(n14099), .B(n14100), .Z(n13733) );
  XOR2_X1 U13933 ( .A(n14101), .B(n14102), .Z(n14099) );
  NOR2_X1 U13934 ( .A1(n9415), .A2(n10061), .ZN(n14102) );
  NOR2_X1 U13935 ( .A1(n10062), .A2(n10059), .ZN(n13842) );
  XNOR2_X1 U13936 ( .A(n14103), .B(n14104), .ZN(n13710) );
  XOR2_X1 U13937 ( .A(n14105), .B(n14106), .Z(n14104) );
  NAND2_X1 U13938 ( .A1(a_15_), .A2(b_16_), .ZN(n14106) );
  XNOR2_X1 U13939 ( .A(n14107), .B(n14108), .ZN(n13650) );
  NAND2_X1 U13940 ( .A1(n14109), .A2(n14110), .ZN(n14107) );
  XNOR2_X1 U13941 ( .A(n14111), .B(n13611), .ZN(n13864) );
  XNOR2_X1 U13942 ( .A(n14112), .B(n14113), .ZN(n13611) );
  XOR2_X1 U13943 ( .A(n14114), .B(n14115), .Z(n10273) );
  NAND2_X1 U13944 ( .A1(n10213), .A2(n10212), .ZN(n10211) );
  NOR2_X1 U13945 ( .A1(n14116), .A2(n10269), .ZN(n10212) );
  NOR2_X1 U13946 ( .A1(n14117), .A2(n14118), .ZN(n14116) );
  NOR2_X1 U13947 ( .A1(n14114), .A2(n14115), .ZN(n10213) );
  NAND2_X1 U13948 ( .A1(n14119), .A2(n14120), .ZN(n14115) );
  NAND2_X1 U13949 ( .A1(n14111), .A2(n14121), .ZN(n14120) );
  NAND2_X1 U13950 ( .A1(n14113), .A2(n14112), .ZN(n14121) );
  INV_X1 U13951 ( .A(n13610), .ZN(n14111) );
  XOR2_X1 U13952 ( .A(n14122), .B(n14123), .Z(n13610) );
  XOR2_X1 U13953 ( .A(n14124), .B(n14125), .Z(n14122) );
  NOR2_X1 U13954 ( .A1(n9983), .A2(n10063), .ZN(n14125) );
  INV_X1 U13955 ( .A(n14126), .ZN(n14119) );
  NOR2_X1 U13956 ( .A1(n14112), .A2(n14113), .ZN(n14126) );
  NOR2_X1 U13957 ( .A1(n10093), .A2(n10061), .ZN(n14113) );
  NAND2_X1 U13958 ( .A1(n13872), .A2(n14127), .ZN(n14112) );
  NAND2_X1 U13959 ( .A1(n13871), .A2(n13873), .ZN(n14127) );
  NAND2_X1 U13960 ( .A1(n14128), .A2(n14129), .ZN(n13873) );
  NAND2_X1 U13961 ( .A1(a_1_), .A2(b_16_), .ZN(n14129) );
  INV_X1 U13962 ( .A(n14130), .ZN(n14128) );
  XNOR2_X1 U13963 ( .A(n14131), .B(n14132), .ZN(n13871) );
  XOR2_X1 U13964 ( .A(n14133), .B(n14134), .Z(n14132) );
  NAND2_X1 U13965 ( .A1(b_15_), .A2(a_2_), .ZN(n14134) );
  NAND2_X1 U13966 ( .A1(a_1_), .A2(n14130), .ZN(n13872) );
  NAND2_X1 U13967 ( .A1(n13880), .A2(n14135), .ZN(n14130) );
  NAND2_X1 U13968 ( .A1(n13879), .A2(n13881), .ZN(n14135) );
  NAND2_X1 U13969 ( .A1(n14136), .A2(n14137), .ZN(n13881) );
  NAND2_X1 U13970 ( .A1(a_2_), .A2(b_16_), .ZN(n14137) );
  INV_X1 U13971 ( .A(n14138), .ZN(n14136) );
  XNOR2_X1 U13972 ( .A(n14139), .B(n14140), .ZN(n13879) );
  XOR2_X1 U13973 ( .A(n14141), .B(n14142), .Z(n14140) );
  NAND2_X1 U13974 ( .A1(b_15_), .A2(a_3_), .ZN(n14142) );
  NAND2_X1 U13975 ( .A1(a_2_), .A2(n14138), .ZN(n13880) );
  NAND2_X1 U13976 ( .A1(n13888), .A2(n14143), .ZN(n14138) );
  NAND2_X1 U13977 ( .A1(n13887), .A2(n13889), .ZN(n14143) );
  NAND2_X1 U13978 ( .A1(n14144), .A2(n14145), .ZN(n13889) );
  NAND2_X1 U13979 ( .A1(a_3_), .A2(b_16_), .ZN(n14145) );
  INV_X1 U13980 ( .A(n14146), .ZN(n14144) );
  XOR2_X1 U13981 ( .A(n14147), .B(n14148), .Z(n13887) );
  XOR2_X1 U13982 ( .A(n14149), .B(n14150), .Z(n14147) );
  NOR2_X1 U13983 ( .A1(n10085), .A2(n10063), .ZN(n14150) );
  NAND2_X1 U13984 ( .A1(a_3_), .A2(n14146), .ZN(n13888) );
  NAND2_X1 U13985 ( .A1(n13896), .A2(n14151), .ZN(n14146) );
  NAND2_X1 U13986 ( .A1(n13895), .A2(n13897), .ZN(n14151) );
  NAND2_X1 U13987 ( .A1(n14152), .A2(n14153), .ZN(n13897) );
  NAND2_X1 U13988 ( .A1(a_4_), .A2(b_16_), .ZN(n14153) );
  INV_X1 U13989 ( .A(n14154), .ZN(n14152) );
  XNOR2_X1 U13990 ( .A(n14155), .B(n14156), .ZN(n13895) );
  XOR2_X1 U13991 ( .A(n14157), .B(n14158), .Z(n14156) );
  NAND2_X1 U13992 ( .A1(b_15_), .A2(a_5_), .ZN(n14158) );
  NAND2_X1 U13993 ( .A1(a_4_), .A2(n14154), .ZN(n13896) );
  NAND2_X1 U13994 ( .A1(n13904), .A2(n14159), .ZN(n14154) );
  NAND2_X1 U13995 ( .A1(n13903), .A2(n13905), .ZN(n14159) );
  NAND2_X1 U13996 ( .A1(n14160), .A2(n14161), .ZN(n13905) );
  NAND2_X1 U13997 ( .A1(a_5_), .A2(b_16_), .ZN(n14161) );
  INV_X1 U13998 ( .A(n14162), .ZN(n14160) );
  XNOR2_X1 U13999 ( .A(n14163), .B(n14164), .ZN(n13903) );
  XOR2_X1 U14000 ( .A(n14165), .B(n14166), .Z(n14164) );
  NAND2_X1 U14001 ( .A1(b_15_), .A2(a_6_), .ZN(n14166) );
  NAND2_X1 U14002 ( .A1(a_5_), .A2(n14162), .ZN(n13904) );
  NAND2_X1 U14003 ( .A1(n14167), .A2(n14168), .ZN(n14162) );
  NAND2_X1 U14004 ( .A1(n14169), .A2(a_6_), .ZN(n14168) );
  NOR2_X1 U14005 ( .A1(n14170), .A2(n10061), .ZN(n14169) );
  NOR2_X1 U14006 ( .A1(n13912), .A2(n13911), .ZN(n14170) );
  NAND2_X1 U14007 ( .A1(n13911), .A2(n13912), .ZN(n14167) );
  NAND2_X1 U14008 ( .A1(n14109), .A2(n14171), .ZN(n13912) );
  NAND2_X1 U14009 ( .A1(n14108), .A2(n14110), .ZN(n14171) );
  NAND2_X1 U14010 ( .A1(n14172), .A2(n14173), .ZN(n14110) );
  NAND2_X1 U14011 ( .A1(a_7_), .A2(b_16_), .ZN(n14173) );
  INV_X1 U14012 ( .A(n14174), .ZN(n14172) );
  XNOR2_X1 U14013 ( .A(n14175), .B(n14176), .ZN(n14108) );
  XNOR2_X1 U14014 ( .A(n14177), .B(n14178), .ZN(n14175) );
  NAND2_X1 U14015 ( .A1(a_7_), .A2(n14174), .ZN(n14109) );
  NAND2_X1 U14016 ( .A1(n14179), .A2(n14180), .ZN(n14174) );
  NAND2_X1 U14017 ( .A1(n14181), .A2(a_8_), .ZN(n14180) );
  NOR2_X1 U14018 ( .A1(n14182), .A2(n10061), .ZN(n14181) );
  NOR2_X1 U14019 ( .A1(n13923), .A2(n13921), .ZN(n14182) );
  NAND2_X1 U14020 ( .A1(n13923), .A2(n13921), .ZN(n14179) );
  XOR2_X1 U14021 ( .A(n14183), .B(n14184), .Z(n13921) );
  XNOR2_X1 U14022 ( .A(n14185), .B(n14186), .ZN(n14184) );
  NAND2_X1 U14023 ( .A1(b_15_), .A2(a_9_), .ZN(n14186) );
  NOR2_X1 U14024 ( .A1(n14187), .A2(n14188), .ZN(n13923) );
  INV_X1 U14025 ( .A(n14189), .ZN(n14188) );
  NAND2_X1 U14026 ( .A1(n13929), .A2(n14190), .ZN(n14189) );
  NAND2_X1 U14027 ( .A1(n13932), .A2(n13931), .ZN(n14190) );
  XOR2_X1 U14028 ( .A(n14191), .B(n14192), .Z(n13929) );
  XOR2_X1 U14029 ( .A(n14193), .B(n14194), .Z(n14191) );
  NOR2_X1 U14030 ( .A1(n13931), .A2(n13932), .ZN(n14187) );
  NOR2_X1 U14031 ( .A1(n10076), .A2(n10061), .ZN(n13932) );
  NAND2_X1 U14032 ( .A1(n13939), .A2(n14195), .ZN(n13931) );
  NAND2_X1 U14033 ( .A1(n13938), .A2(n13940), .ZN(n14195) );
  NAND2_X1 U14034 ( .A1(n14196), .A2(n14197), .ZN(n13940) );
  NAND2_X1 U14035 ( .A1(a_10_), .A2(b_16_), .ZN(n14197) );
  INV_X1 U14036 ( .A(n14198), .ZN(n14196) );
  XNOR2_X1 U14037 ( .A(n14199), .B(n14200), .ZN(n13938) );
  XOR2_X1 U14038 ( .A(n14201), .B(n14202), .Z(n14200) );
  NAND2_X1 U14039 ( .A1(b_15_), .A2(a_11_), .ZN(n14202) );
  NAND2_X1 U14040 ( .A1(a_10_), .A2(n14198), .ZN(n13939) );
  NAND2_X1 U14041 ( .A1(n13947), .A2(n14203), .ZN(n14198) );
  NAND2_X1 U14042 ( .A1(n13946), .A2(n13948), .ZN(n14203) );
  NAND2_X1 U14043 ( .A1(n14204), .A2(n14205), .ZN(n13948) );
  NAND2_X1 U14044 ( .A1(a_11_), .A2(b_16_), .ZN(n14205) );
  INV_X1 U14045 ( .A(n14206), .ZN(n14204) );
  XNOR2_X1 U14046 ( .A(n14207), .B(n14208), .ZN(n13946) );
  XNOR2_X1 U14047 ( .A(n14209), .B(n14210), .ZN(n14207) );
  NOR2_X1 U14048 ( .A1(n10070), .A2(n10063), .ZN(n14210) );
  NAND2_X1 U14049 ( .A1(a_11_), .A2(n14206), .ZN(n13947) );
  NAND2_X1 U14050 ( .A1(n13956), .A2(n14211), .ZN(n14206) );
  NAND2_X1 U14051 ( .A1(n13955), .A2(n13957), .ZN(n14211) );
  NAND2_X1 U14052 ( .A1(n14212), .A2(n14213), .ZN(n13957) );
  NAND2_X1 U14053 ( .A1(a_12_), .A2(b_16_), .ZN(n14213) );
  INV_X1 U14054 ( .A(n14214), .ZN(n14212) );
  XOR2_X1 U14055 ( .A(n14215), .B(n14216), .Z(n13955) );
  XNOR2_X1 U14056 ( .A(n14217), .B(n14218), .ZN(n14216) );
  NAND2_X1 U14057 ( .A1(a_12_), .A2(n14214), .ZN(n13956) );
  NAND2_X1 U14058 ( .A1(n14219), .A2(n14220), .ZN(n14214) );
  NAND2_X1 U14059 ( .A1(n14221), .A2(a_13_), .ZN(n14220) );
  NOR2_X1 U14060 ( .A1(n14222), .A2(n10061), .ZN(n14221) );
  NOR2_X1 U14061 ( .A1(n13964), .A2(n13963), .ZN(n14222) );
  NAND2_X1 U14062 ( .A1(n13963), .A2(n13964), .ZN(n14219) );
  NAND2_X1 U14063 ( .A1(n14223), .A2(n14224), .ZN(n13964) );
  NAND2_X1 U14064 ( .A1(n14225), .A2(a_14_), .ZN(n14224) );
  NOR2_X1 U14065 ( .A1(n14226), .A2(n10061), .ZN(n14225) );
  NOR2_X1 U14066 ( .A1(n13973), .A2(n13971), .ZN(n14226) );
  NAND2_X1 U14067 ( .A1(n13971), .A2(n13973), .ZN(n14223) );
  NAND2_X1 U14068 ( .A1(n14227), .A2(n14228), .ZN(n13973) );
  NAND2_X1 U14069 ( .A1(n14229), .A2(a_15_), .ZN(n14228) );
  NOR2_X1 U14070 ( .A1(n14230), .A2(n10061), .ZN(n14229) );
  NOR2_X1 U14071 ( .A1(n14105), .A2(n14103), .ZN(n14230) );
  NAND2_X1 U14072 ( .A1(n14103), .A2(n14105), .ZN(n14227) );
  NAND2_X1 U14073 ( .A1(n14231), .A2(n14232), .ZN(n14105) );
  NAND2_X1 U14074 ( .A1(n13983), .A2(n14233), .ZN(n14232) );
  INV_X1 U14075 ( .A(n14234), .ZN(n14233) );
  NOR2_X1 U14076 ( .A1(n13984), .A2(n14235), .ZN(n14234) );
  XNOR2_X1 U14077 ( .A(n14236), .B(n14237), .ZN(n13983) );
  NAND2_X1 U14078 ( .A1(n14238), .A2(n14239), .ZN(n14236) );
  NAND2_X1 U14079 ( .A1(n14235), .A2(n13984), .ZN(n14231) );
  NAND2_X1 U14080 ( .A1(n13991), .A2(n14240), .ZN(n13984) );
  NAND2_X1 U14081 ( .A1(n13990), .A2(n13992), .ZN(n14240) );
  NAND2_X1 U14082 ( .A1(n14241), .A2(n14242), .ZN(n13992) );
  NAND2_X1 U14083 ( .A1(b_16_), .A2(a_17_), .ZN(n14242) );
  INV_X1 U14084 ( .A(n14243), .ZN(n14241) );
  XNOR2_X1 U14085 ( .A(n14244), .B(n14245), .ZN(n13990) );
  XOR2_X1 U14086 ( .A(n14246), .B(n14247), .Z(n14245) );
  NAND2_X1 U14087 ( .A1(b_15_), .A2(a_18_), .ZN(n14247) );
  NAND2_X1 U14088 ( .A1(a_17_), .A2(n14243), .ZN(n13991) );
  NAND2_X1 U14089 ( .A1(n14248), .A2(n14249), .ZN(n14243) );
  NAND2_X1 U14090 ( .A1(n14250), .A2(b_16_), .ZN(n14249) );
  NOR2_X1 U14091 ( .A1(n14251), .A2(n10058), .ZN(n14250) );
  NOR2_X1 U14092 ( .A1(n14000), .A2(n13999), .ZN(n14251) );
  NAND2_X1 U14093 ( .A1(n13999), .A2(n14000), .ZN(n14248) );
  NAND2_X1 U14094 ( .A1(n14252), .A2(n14253), .ZN(n14000) );
  NAND2_X1 U14095 ( .A1(n14254), .A2(b_16_), .ZN(n14253) );
  NOR2_X1 U14096 ( .A1(n14255), .A2(n9415), .ZN(n14254) );
  NOR2_X1 U14097 ( .A1(n14100), .A2(n14101), .ZN(n14255) );
  NAND2_X1 U14098 ( .A1(n14100), .A2(n14101), .ZN(n14252) );
  NAND2_X1 U14099 ( .A1(n14256), .A2(n14257), .ZN(n14101) );
  NAND2_X1 U14100 ( .A1(n14013), .A2(n14258), .ZN(n14257) );
  INV_X1 U14101 ( .A(n14259), .ZN(n14258) );
  NOR2_X1 U14102 ( .A1(n14011), .A2(n14012), .ZN(n14259) );
  NOR2_X1 U14103 ( .A1(n10061), .A2(n10054), .ZN(n14013) );
  NAND2_X1 U14104 ( .A1(n14012), .A2(n14011), .ZN(n14256) );
  XNOR2_X1 U14105 ( .A(n14260), .B(n14261), .ZN(n14011) );
  NAND2_X1 U14106 ( .A1(n14262), .A2(n14263), .ZN(n14260) );
  NOR2_X1 U14107 ( .A1(n14264), .A2(n14265), .ZN(n14012) );
  NOR2_X1 U14108 ( .A1(n14018), .A2(n14266), .ZN(n14265) );
  INV_X1 U14109 ( .A(n14267), .ZN(n14266) );
  NAND2_X1 U14110 ( .A1(n14020), .A2(n14019), .ZN(n14267) );
  XOR2_X1 U14111 ( .A(n14268), .B(n14269), .Z(n14018) );
  XOR2_X1 U14112 ( .A(n14270), .B(n14271), .Z(n14268) );
  NOR2_X1 U14113 ( .A1(n14019), .A2(n14020), .ZN(n14264) );
  NOR2_X1 U14114 ( .A1(n10061), .A2(n9358), .ZN(n14020) );
  NAND2_X1 U14115 ( .A1(n14028), .A2(n14272), .ZN(n14019) );
  NAND2_X1 U14116 ( .A1(n14027), .A2(n14029), .ZN(n14272) );
  NAND2_X1 U14117 ( .A1(n14273), .A2(n14274), .ZN(n14029) );
  NAND2_X1 U14118 ( .A1(b_16_), .A2(a_22_), .ZN(n14274) );
  INV_X1 U14119 ( .A(n14275), .ZN(n14273) );
  XOR2_X1 U14120 ( .A(n14276), .B(n14277), .Z(n14027) );
  XNOR2_X1 U14121 ( .A(n14278), .B(n14279), .ZN(n14276) );
  NAND2_X1 U14122 ( .A1(a_22_), .A2(n14275), .ZN(n14028) );
  NAND2_X1 U14123 ( .A1(n14097), .A2(n14280), .ZN(n14275) );
  NAND2_X1 U14124 ( .A1(n14096), .A2(n14098), .ZN(n14280) );
  NAND2_X1 U14125 ( .A1(n14281), .A2(n14282), .ZN(n14098) );
  NAND2_X1 U14126 ( .A1(b_16_), .A2(a_23_), .ZN(n14282) );
  INV_X1 U14127 ( .A(n14283), .ZN(n14281) );
  XNOR2_X1 U14128 ( .A(n14284), .B(n14285), .ZN(n14096) );
  XOR2_X1 U14129 ( .A(n14286), .B(n14287), .Z(n14285) );
  NAND2_X1 U14130 ( .A1(a_23_), .A2(n14283), .ZN(n14097) );
  NAND2_X1 U14131 ( .A1(n14288), .A2(n14289), .ZN(n14283) );
  INV_X1 U14132 ( .A(n14290), .ZN(n14289) );
  NOR2_X1 U14133 ( .A1(n14094), .A2(n14291), .ZN(n14290) );
  NOR2_X1 U14134 ( .A1(n14093), .A2(n14091), .ZN(n14291) );
  NAND2_X1 U14135 ( .A1(b_16_), .A2(a_24_), .ZN(n14094) );
  NAND2_X1 U14136 ( .A1(n14091), .A2(n14093), .ZN(n14288) );
  NAND2_X1 U14137 ( .A1(n14292), .A2(n14293), .ZN(n14093) );
  NAND2_X1 U14138 ( .A1(n14090), .A2(n14294), .ZN(n14293) );
  NAND2_X1 U14139 ( .A1(n14087), .A2(n14089), .ZN(n14294) );
  NOR2_X1 U14140 ( .A1(n10061), .A2(n10048), .ZN(n14090) );
  INV_X1 U14141 ( .A(n14295), .ZN(n14292) );
  NOR2_X1 U14142 ( .A1(n14087), .A2(n14089), .ZN(n14295) );
  NAND2_X1 U14143 ( .A1(n14296), .A2(n14297), .ZN(n14089) );
  NAND2_X1 U14144 ( .A1(n14047), .A2(n14298), .ZN(n14297) );
  NAND2_X1 U14145 ( .A1(n14050), .A2(n14049), .ZN(n14298) );
  XOR2_X1 U14146 ( .A(n14299), .B(n14300), .Z(n14047) );
  NAND2_X1 U14147 ( .A1(n14301), .A2(n14302), .ZN(n14299) );
  INV_X1 U14148 ( .A(n14303), .ZN(n14296) );
  NOR2_X1 U14149 ( .A1(n14049), .A2(n14050), .ZN(n14303) );
  NOR2_X1 U14150 ( .A1(n10061), .A2(n10047), .ZN(n14050) );
  NAND2_X1 U14151 ( .A1(n14056), .A2(n14304), .ZN(n14049) );
  NAND2_X1 U14152 ( .A1(n14055), .A2(n14057), .ZN(n14304) );
  NAND2_X1 U14153 ( .A1(n14305), .A2(n14306), .ZN(n14057) );
  NAND2_X1 U14154 ( .A1(b_16_), .A2(a_27_), .ZN(n14306) );
  INV_X1 U14155 ( .A(n14307), .ZN(n14305) );
  XNOR2_X1 U14156 ( .A(n14308), .B(n14309), .ZN(n14055) );
  XOR2_X1 U14157 ( .A(n14310), .B(n14311), .Z(n14309) );
  NAND2_X1 U14158 ( .A1(b_15_), .A2(a_28_), .ZN(n14311) );
  NAND2_X1 U14159 ( .A1(a_27_), .A2(n14307), .ZN(n14056) );
  NAND2_X1 U14160 ( .A1(n14312), .A2(n14313), .ZN(n14307) );
  NAND2_X1 U14161 ( .A1(n14314), .A2(b_16_), .ZN(n14313) );
  NOR2_X1 U14162 ( .A1(n14315), .A2(n9136), .ZN(n14314) );
  NOR2_X1 U14163 ( .A1(n14063), .A2(n14065), .ZN(n14315) );
  NAND2_X1 U14164 ( .A1(n14063), .A2(n14065), .ZN(n14312) );
  NAND2_X1 U14165 ( .A1(n14316), .A2(n14317), .ZN(n14065) );
  NAND2_X1 U14166 ( .A1(n14318), .A2(b_16_), .ZN(n14317) );
  NOR2_X1 U14167 ( .A1(n14319), .A2(n9121), .ZN(n14318) );
  NOR2_X1 U14168 ( .A1(n14320), .A2(n14085), .ZN(n14319) );
  NAND2_X1 U14169 ( .A1(n14320), .A2(n14085), .ZN(n14316) );
  NAND2_X1 U14170 ( .A1(n14321), .A2(n14322), .ZN(n14085) );
  NAND2_X1 U14171 ( .A1(b_14_), .A2(n14323), .ZN(n14322) );
  NAND2_X1 U14172 ( .A1(n10486), .A2(n14324), .ZN(n14323) );
  NAND2_X1 U14173 ( .A1(a_31_), .A2(n10063), .ZN(n14324) );
  NAND2_X1 U14174 ( .A1(b_15_), .A2(n14325), .ZN(n14321) );
  NAND2_X1 U14175 ( .A1(n10489), .A2(n14326), .ZN(n14325) );
  NAND2_X1 U14176 ( .A1(a_30_), .A2(n10064), .ZN(n14326) );
  INV_X1 U14177 ( .A(n14086), .ZN(n14320) );
  NAND2_X1 U14178 ( .A1(n14327), .A2(n9025), .ZN(n14086) );
  NOR2_X1 U14179 ( .A1(n10061), .A2(n10063), .ZN(n14327) );
  XOR2_X1 U14180 ( .A(n14328), .B(n14329), .Z(n14063) );
  NOR2_X1 U14181 ( .A1(n9121), .A2(n10063), .ZN(n14329) );
  XNOR2_X1 U14182 ( .A(n14330), .B(n14331), .ZN(n14328) );
  XNOR2_X1 U14183 ( .A(n14332), .B(n14333), .ZN(n14087) );
  XNOR2_X1 U14184 ( .A(n14334), .B(n14335), .ZN(n14333) );
  XNOR2_X1 U14185 ( .A(n14336), .B(n14337), .ZN(n14091) );
  XNOR2_X1 U14186 ( .A(n14338), .B(n14339), .ZN(n14337) );
  XOR2_X1 U14187 ( .A(n14340), .B(n14341), .Z(n14100) );
  XOR2_X1 U14188 ( .A(n14342), .B(n14343), .Z(n14340) );
  NOR2_X1 U14189 ( .A1(n10054), .A2(n10063), .ZN(n14343) );
  XNOR2_X1 U14190 ( .A(n14344), .B(n14345), .ZN(n13999) );
  XOR2_X1 U14191 ( .A(n14346), .B(n14347), .Z(n14345) );
  NAND2_X1 U14192 ( .A1(b_15_), .A2(a_19_), .ZN(n14347) );
  INV_X1 U14193 ( .A(n9512), .ZN(n14235) );
  NAND2_X1 U14194 ( .A1(b_16_), .A2(a_16_), .ZN(n9512) );
  XNOR2_X1 U14195 ( .A(n14348), .B(n14349), .ZN(n14103) );
  XOR2_X1 U14196 ( .A(n14350), .B(n14351), .Z(n14348) );
  XNOR2_X1 U14197 ( .A(n14352), .B(n14353), .ZN(n13971) );
  XOR2_X1 U14198 ( .A(n14354), .B(n10003), .Z(n14353) );
  XNOR2_X1 U14199 ( .A(n14355), .B(n14356), .ZN(n13963) );
  XNOR2_X1 U14200 ( .A(n14357), .B(n14358), .ZN(n14355) );
  NOR2_X1 U14201 ( .A1(n10065), .A2(n10063), .ZN(n14358) );
  XNOR2_X1 U14202 ( .A(n14359), .B(n14360), .ZN(n13911) );
  XNOR2_X1 U14203 ( .A(n14361), .B(n14362), .ZN(n14359) );
  NOR2_X1 U14204 ( .A1(n9773), .A2(n10063), .ZN(n14362) );
  XNOR2_X1 U14205 ( .A(n14363), .B(n14364), .ZN(n14114) );
  XOR2_X1 U14206 ( .A(n14365), .B(n14366), .Z(n14363) );
  NOR2_X1 U14207 ( .A1(n10093), .A2(n10063), .ZN(n14366) );
  INV_X1 U14208 ( .A(n14367), .ZN(n10269) );
  NAND2_X1 U14209 ( .A1(n14117), .A2(n14118), .ZN(n14367) );
  NAND2_X1 U14210 ( .A1(n14368), .A2(n14369), .ZN(n14118) );
  NAND2_X1 U14211 ( .A1(n14370), .A2(b_15_), .ZN(n14369) );
  NOR2_X1 U14212 ( .A1(n14371), .A2(n10093), .ZN(n14370) );
  NOR2_X1 U14213 ( .A1(n14364), .A2(n14365), .ZN(n14371) );
  NAND2_X1 U14214 ( .A1(n14364), .A2(n14365), .ZN(n14368) );
  NAND2_X1 U14215 ( .A1(n14372), .A2(n14373), .ZN(n14365) );
  NAND2_X1 U14216 ( .A1(n14374), .A2(b_15_), .ZN(n14373) );
  NOR2_X1 U14217 ( .A1(n14375), .A2(n9983), .ZN(n14374) );
  NOR2_X1 U14218 ( .A1(n14123), .A2(n14124), .ZN(n14375) );
  NAND2_X1 U14219 ( .A1(n14123), .A2(n14124), .ZN(n14372) );
  NAND2_X1 U14220 ( .A1(n14376), .A2(n14377), .ZN(n14124) );
  NAND2_X1 U14221 ( .A1(n14378), .A2(b_15_), .ZN(n14377) );
  NOR2_X1 U14222 ( .A1(n14379), .A2(n10088), .ZN(n14378) );
  NOR2_X1 U14223 ( .A1(n14131), .A2(n14133), .ZN(n14379) );
  NAND2_X1 U14224 ( .A1(n14131), .A2(n14133), .ZN(n14376) );
  NAND2_X1 U14225 ( .A1(n14380), .A2(n14381), .ZN(n14133) );
  NAND2_X1 U14226 ( .A1(n14382), .A2(b_15_), .ZN(n14381) );
  NOR2_X1 U14227 ( .A1(n14383), .A2(n10086), .ZN(n14382) );
  NOR2_X1 U14228 ( .A1(n14139), .A2(n14141), .ZN(n14383) );
  NAND2_X1 U14229 ( .A1(n14139), .A2(n14141), .ZN(n14380) );
  NAND2_X1 U14230 ( .A1(n14384), .A2(n14385), .ZN(n14141) );
  NAND2_X1 U14231 ( .A1(n14386), .A2(b_15_), .ZN(n14385) );
  NOR2_X1 U14232 ( .A1(n14387), .A2(n10085), .ZN(n14386) );
  NOR2_X1 U14233 ( .A1(n14148), .A2(n14149), .ZN(n14387) );
  NAND2_X1 U14234 ( .A1(n14148), .A2(n14149), .ZN(n14384) );
  NAND2_X1 U14235 ( .A1(n14388), .A2(n14389), .ZN(n14149) );
  NAND2_X1 U14236 ( .A1(n14390), .A2(b_15_), .ZN(n14389) );
  NOR2_X1 U14237 ( .A1(n14391), .A2(n10083), .ZN(n14390) );
  NOR2_X1 U14238 ( .A1(n14155), .A2(n14157), .ZN(n14391) );
  NAND2_X1 U14239 ( .A1(n14155), .A2(n14157), .ZN(n14388) );
  NAND2_X1 U14240 ( .A1(n14392), .A2(n14393), .ZN(n14157) );
  NAND2_X1 U14241 ( .A1(n14394), .A2(b_15_), .ZN(n14393) );
  NOR2_X1 U14242 ( .A1(n14395), .A2(n10081), .ZN(n14394) );
  NOR2_X1 U14243 ( .A1(n14163), .A2(n14165), .ZN(n14395) );
  NAND2_X1 U14244 ( .A1(n14163), .A2(n14165), .ZN(n14392) );
  NAND2_X1 U14245 ( .A1(n14396), .A2(n14397), .ZN(n14165) );
  NAND2_X1 U14246 ( .A1(n14398), .A2(b_15_), .ZN(n14397) );
  NOR2_X1 U14247 ( .A1(n14399), .A2(n9773), .ZN(n14398) );
  NOR2_X1 U14248 ( .A1(n14361), .A2(n14360), .ZN(n14399) );
  NAND2_X1 U14249 ( .A1(n14361), .A2(n14360), .ZN(n14396) );
  XOR2_X1 U14250 ( .A(n14400), .B(n14401), .Z(n14360) );
  XNOR2_X1 U14251 ( .A(n14402), .B(n14403), .ZN(n14401) );
  INV_X1 U14252 ( .A(n14404), .ZN(n14361) );
  NAND2_X1 U14253 ( .A1(n14405), .A2(n14406), .ZN(n14404) );
  NAND2_X1 U14254 ( .A1(n14176), .A2(n14407), .ZN(n14406) );
  NAND2_X1 U14255 ( .A1(n14177), .A2(n14408), .ZN(n14407) );
  XOR2_X1 U14256 ( .A(n14409), .B(n14410), .Z(n14176) );
  XNOR2_X1 U14257 ( .A(n14411), .B(n14412), .ZN(n14410) );
  NAND2_X1 U14258 ( .A1(n14178), .A2(n14413), .ZN(n14405) );
  INV_X1 U14259 ( .A(n14177), .ZN(n14413) );
  NOR2_X1 U14260 ( .A1(n10063), .A2(n10079), .ZN(n14177) );
  INV_X1 U14261 ( .A(n14408), .ZN(n14178) );
  NAND2_X1 U14262 ( .A1(n14414), .A2(n14415), .ZN(n14408) );
  NAND2_X1 U14263 ( .A1(n14416), .A2(b_15_), .ZN(n14415) );
  NOR2_X1 U14264 ( .A1(n14417), .A2(n10076), .ZN(n14416) );
  NOR2_X1 U14265 ( .A1(n14185), .A2(n14183), .ZN(n14417) );
  NAND2_X1 U14266 ( .A1(n14185), .A2(n14183), .ZN(n14414) );
  XNOR2_X1 U14267 ( .A(n14418), .B(n14419), .ZN(n14183) );
  XOR2_X1 U14268 ( .A(n14420), .B(n14421), .Z(n14418) );
  NOR2_X1 U14269 ( .A1(n14422), .A2(n14423), .ZN(n14185) );
  INV_X1 U14270 ( .A(n14424), .ZN(n14423) );
  NAND2_X1 U14271 ( .A1(n14192), .A2(n14425), .ZN(n14424) );
  NAND2_X1 U14272 ( .A1(n14194), .A2(n14193), .ZN(n14425) );
  XOR2_X1 U14273 ( .A(n14426), .B(n14427), .Z(n14192) );
  XNOR2_X1 U14274 ( .A(n14428), .B(n14429), .ZN(n14427) );
  NOR2_X1 U14275 ( .A1(n14193), .A2(n14194), .ZN(n14422) );
  NOR2_X1 U14276 ( .A1(n10063), .A2(n10073), .ZN(n14194) );
  NAND2_X1 U14277 ( .A1(n14430), .A2(n14431), .ZN(n14193) );
  NAND2_X1 U14278 ( .A1(n14432), .A2(b_15_), .ZN(n14431) );
  NOR2_X1 U14279 ( .A1(n14433), .A2(n9649), .ZN(n14432) );
  NOR2_X1 U14280 ( .A1(n14199), .A2(n14201), .ZN(n14433) );
  NAND2_X1 U14281 ( .A1(n14199), .A2(n14201), .ZN(n14430) );
  NAND2_X1 U14282 ( .A1(n14434), .A2(n14435), .ZN(n14201) );
  NAND2_X1 U14283 ( .A1(n14436), .A2(b_15_), .ZN(n14435) );
  NOR2_X1 U14284 ( .A1(n14437), .A2(n10070), .ZN(n14436) );
  NOR2_X1 U14285 ( .A1(n14209), .A2(n14208), .ZN(n14437) );
  NAND2_X1 U14286 ( .A1(n14209), .A2(n14208), .ZN(n14434) );
  XNOR2_X1 U14287 ( .A(n14438), .B(n14439), .ZN(n14208) );
  XNOR2_X1 U14288 ( .A(n14440), .B(n14441), .ZN(n14438) );
  NOR2_X1 U14289 ( .A1(n14442), .A2(n14443), .ZN(n14209) );
  INV_X1 U14290 ( .A(n14444), .ZN(n14443) );
  NAND2_X1 U14291 ( .A1(n14215), .A2(n14445), .ZN(n14444) );
  NAND2_X1 U14292 ( .A1(n14218), .A2(n14217), .ZN(n14445) );
  XOR2_X1 U14293 ( .A(n14446), .B(n14447), .Z(n14215) );
  XNOR2_X1 U14294 ( .A(n14448), .B(n9569), .ZN(n14446) );
  INV_X1 U14295 ( .A(n14449), .ZN(n9569) );
  NOR2_X1 U14296 ( .A1(n14217), .A2(n14218), .ZN(n14442) );
  NOR2_X1 U14297 ( .A1(n10063), .A2(n10067), .ZN(n14218) );
  NAND2_X1 U14298 ( .A1(n14450), .A2(n14451), .ZN(n14217) );
  NAND2_X1 U14299 ( .A1(n14452), .A2(b_15_), .ZN(n14451) );
  NOR2_X1 U14300 ( .A1(n14453), .A2(n10065), .ZN(n14452) );
  NOR2_X1 U14301 ( .A1(n14357), .A2(n14356), .ZN(n14453) );
  NAND2_X1 U14302 ( .A1(n14357), .A2(n14356), .ZN(n14450) );
  XNOR2_X1 U14303 ( .A(n14454), .B(n14455), .ZN(n14356) );
  NAND2_X1 U14304 ( .A1(n14456), .A2(n14457), .ZN(n14454) );
  INV_X1 U14305 ( .A(n14458), .ZN(n14357) );
  NAND2_X1 U14306 ( .A1(n14459), .A2(n14460), .ZN(n14458) );
  NAND2_X1 U14307 ( .A1(n14352), .A2(n14461), .ZN(n14460) );
  INV_X1 U14308 ( .A(n14462), .ZN(n14461) );
  NOR2_X1 U14309 ( .A1(n14354), .A2(n10003), .ZN(n14462) );
  XOR2_X1 U14310 ( .A(n14463), .B(n14464), .Z(n14352) );
  NAND2_X1 U14311 ( .A1(n14465), .A2(n14466), .ZN(n14463) );
  NAND2_X1 U14312 ( .A1(n10003), .A2(n14354), .ZN(n14459) );
  NAND2_X1 U14313 ( .A1(n14467), .A2(n14468), .ZN(n14354) );
  NAND2_X1 U14314 ( .A1(n14349), .A2(n14469), .ZN(n14468) );
  NAND2_X1 U14315 ( .A1(n14351), .A2(n14350), .ZN(n14469) );
  XOR2_X1 U14316 ( .A(n14470), .B(n14471), .Z(n14349) );
  NAND2_X1 U14317 ( .A1(n14472), .A2(n14473), .ZN(n14470) );
  INV_X1 U14318 ( .A(n14474), .ZN(n14467) );
  NOR2_X1 U14319 ( .A1(n14350), .A2(n14351), .ZN(n14474) );
  NOR2_X1 U14320 ( .A1(n10063), .A2(n10062), .ZN(n14351) );
  NAND2_X1 U14321 ( .A1(n14238), .A2(n14475), .ZN(n14350) );
  NAND2_X1 U14322 ( .A1(n14237), .A2(n14239), .ZN(n14475) );
  NAND2_X1 U14323 ( .A1(n14476), .A2(n14477), .ZN(n14239) );
  NAND2_X1 U14324 ( .A1(b_15_), .A2(a_17_), .ZN(n14477) );
  INV_X1 U14325 ( .A(n14478), .ZN(n14476) );
  XNOR2_X1 U14326 ( .A(n14479), .B(n14480), .ZN(n14237) );
  XOR2_X1 U14327 ( .A(n14481), .B(n14482), .Z(n14480) );
  NAND2_X1 U14328 ( .A1(b_14_), .A2(a_18_), .ZN(n14482) );
  NAND2_X1 U14329 ( .A1(a_17_), .A2(n14478), .ZN(n14238) );
  NAND2_X1 U14330 ( .A1(n14483), .A2(n14484), .ZN(n14478) );
  NAND2_X1 U14331 ( .A1(n14485), .A2(b_15_), .ZN(n14484) );
  NOR2_X1 U14332 ( .A1(n14486), .A2(n10058), .ZN(n14485) );
  NOR2_X1 U14333 ( .A1(n14244), .A2(n14246), .ZN(n14486) );
  NAND2_X1 U14334 ( .A1(n14244), .A2(n14246), .ZN(n14483) );
  NAND2_X1 U14335 ( .A1(n14487), .A2(n14488), .ZN(n14246) );
  NAND2_X1 U14336 ( .A1(n14489), .A2(b_15_), .ZN(n14488) );
  NOR2_X1 U14337 ( .A1(n14490), .A2(n9415), .ZN(n14489) );
  NOR2_X1 U14338 ( .A1(n14344), .A2(n14346), .ZN(n14490) );
  NAND2_X1 U14339 ( .A1(n14344), .A2(n14346), .ZN(n14487) );
  NAND2_X1 U14340 ( .A1(n14491), .A2(n14492), .ZN(n14346) );
  NAND2_X1 U14341 ( .A1(n14493), .A2(b_15_), .ZN(n14492) );
  NOR2_X1 U14342 ( .A1(n14494), .A2(n10054), .ZN(n14493) );
  NOR2_X1 U14343 ( .A1(n14341), .A2(n14342), .ZN(n14494) );
  NAND2_X1 U14344 ( .A1(n14341), .A2(n14342), .ZN(n14491) );
  NAND2_X1 U14345 ( .A1(n14262), .A2(n14495), .ZN(n14342) );
  NAND2_X1 U14346 ( .A1(n14261), .A2(n14263), .ZN(n14495) );
  NAND2_X1 U14347 ( .A1(n14496), .A2(n14497), .ZN(n14263) );
  NAND2_X1 U14348 ( .A1(b_15_), .A2(a_21_), .ZN(n14497) );
  INV_X1 U14349 ( .A(n14498), .ZN(n14496) );
  XNOR2_X1 U14350 ( .A(n14499), .B(n14500), .ZN(n14261) );
  XNOR2_X1 U14351 ( .A(n14501), .B(n14502), .ZN(n14499) );
  NAND2_X1 U14352 ( .A1(a_21_), .A2(n14498), .ZN(n14262) );
  NAND2_X1 U14353 ( .A1(n14503), .A2(n14504), .ZN(n14498) );
  NAND2_X1 U14354 ( .A1(n14271), .A2(n14505), .ZN(n14504) );
  INV_X1 U14355 ( .A(n14506), .ZN(n14505) );
  NOR2_X1 U14356 ( .A1(n14270), .A2(n14269), .ZN(n14506) );
  NOR2_X1 U14357 ( .A1(n10063), .A2(n9330), .ZN(n14271) );
  NAND2_X1 U14358 ( .A1(n14269), .A2(n14270), .ZN(n14503) );
  NAND2_X1 U14359 ( .A1(n14507), .A2(n14508), .ZN(n14270) );
  NAND2_X1 U14360 ( .A1(n14279), .A2(n14509), .ZN(n14508) );
  NAND2_X1 U14361 ( .A1(n14278), .A2(n14510), .ZN(n14509) );
  INV_X1 U14362 ( .A(n14277), .ZN(n14510) );
  NOR2_X1 U14363 ( .A1(n10063), .A2(n10051), .ZN(n14279) );
  NAND2_X1 U14364 ( .A1(n14277), .A2(n14511), .ZN(n14507) );
  INV_X1 U14365 ( .A(n14278), .ZN(n14511) );
  NOR2_X1 U14366 ( .A1(n14512), .A2(n14513), .ZN(n14278) );
  NOR2_X1 U14367 ( .A1(n14287), .A2(n14514), .ZN(n14513) );
  NOR2_X1 U14368 ( .A1(n14286), .A2(n14284), .ZN(n14514) );
  NAND2_X1 U14369 ( .A1(b_15_), .A2(a_24_), .ZN(n14287) );
  INV_X1 U14370 ( .A(n14515), .ZN(n14512) );
  NAND2_X1 U14371 ( .A1(n14284), .A2(n14286), .ZN(n14515) );
  NAND2_X1 U14372 ( .A1(n14516), .A2(n14517), .ZN(n14286) );
  NAND2_X1 U14373 ( .A1(n14339), .A2(n14518), .ZN(n14517) );
  NAND2_X1 U14374 ( .A1(n14336), .A2(n14338), .ZN(n14518) );
  NOR2_X1 U14375 ( .A1(n10063), .A2(n10048), .ZN(n14339) );
  INV_X1 U14376 ( .A(n14519), .ZN(n14516) );
  NOR2_X1 U14377 ( .A1(n14338), .A2(n14336), .ZN(n14519) );
  XNOR2_X1 U14378 ( .A(n14520), .B(n14521), .ZN(n14336) );
  XNOR2_X1 U14379 ( .A(n14522), .B(n14523), .ZN(n14521) );
  NAND2_X1 U14380 ( .A1(n14524), .A2(n14525), .ZN(n14338) );
  NAND2_X1 U14381 ( .A1(n14332), .A2(n14526), .ZN(n14525) );
  NAND2_X1 U14382 ( .A1(n14335), .A2(n14334), .ZN(n14526) );
  XOR2_X1 U14383 ( .A(n14527), .B(n14528), .Z(n14332) );
  NAND2_X1 U14384 ( .A1(n14529), .A2(n14530), .ZN(n14527) );
  INV_X1 U14385 ( .A(n14531), .ZN(n14524) );
  NOR2_X1 U14386 ( .A1(n14334), .A2(n14335), .ZN(n14531) );
  NOR2_X1 U14387 ( .A1(n10063), .A2(n10047), .ZN(n14335) );
  NAND2_X1 U14388 ( .A1(n14301), .A2(n14532), .ZN(n14334) );
  NAND2_X1 U14389 ( .A1(n14300), .A2(n14302), .ZN(n14532) );
  NAND2_X1 U14390 ( .A1(n14533), .A2(n14534), .ZN(n14302) );
  NAND2_X1 U14391 ( .A1(b_15_), .A2(a_27_), .ZN(n14534) );
  INV_X1 U14392 ( .A(n14535), .ZN(n14533) );
  XNOR2_X1 U14393 ( .A(n14536), .B(n14537), .ZN(n14300) );
  XOR2_X1 U14394 ( .A(n14538), .B(n14539), .Z(n14537) );
  NAND2_X1 U14395 ( .A1(b_14_), .A2(a_28_), .ZN(n14539) );
  NAND2_X1 U14396 ( .A1(a_27_), .A2(n14535), .ZN(n14301) );
  NAND2_X1 U14397 ( .A1(n14540), .A2(n14541), .ZN(n14535) );
  NAND2_X1 U14398 ( .A1(n14542), .A2(b_15_), .ZN(n14541) );
  NOR2_X1 U14399 ( .A1(n14543), .A2(n9136), .ZN(n14542) );
  NOR2_X1 U14400 ( .A1(n14308), .A2(n14310), .ZN(n14543) );
  NAND2_X1 U14401 ( .A1(n14308), .A2(n14310), .ZN(n14540) );
  NAND2_X1 U14402 ( .A1(n14544), .A2(n14545), .ZN(n14310) );
  NAND2_X1 U14403 ( .A1(n14546), .A2(b_15_), .ZN(n14545) );
  NOR2_X1 U14404 ( .A1(n14547), .A2(n9121), .ZN(n14546) );
  NOR2_X1 U14405 ( .A1(n14548), .A2(n14330), .ZN(n14547) );
  NAND2_X1 U14406 ( .A1(n14548), .A2(n14330), .ZN(n14544) );
  NAND2_X1 U14407 ( .A1(n14549), .A2(n14550), .ZN(n14330) );
  NAND2_X1 U14408 ( .A1(b_13_), .A2(n14551), .ZN(n14550) );
  NAND2_X1 U14409 ( .A1(n10486), .A2(n14552), .ZN(n14551) );
  NAND2_X1 U14410 ( .A1(a_31_), .A2(n10064), .ZN(n14552) );
  NAND2_X1 U14411 ( .A1(b_14_), .A2(n14553), .ZN(n14549) );
  NAND2_X1 U14412 ( .A1(n10489), .A2(n14554), .ZN(n14553) );
  NAND2_X1 U14413 ( .A1(a_30_), .A2(n10066), .ZN(n14554) );
  INV_X1 U14414 ( .A(n14331), .ZN(n14548) );
  NAND2_X1 U14415 ( .A1(n14555), .A2(n9025), .ZN(n14331) );
  NOR2_X1 U14416 ( .A1(n10063), .A2(n10064), .ZN(n14555) );
  XOR2_X1 U14417 ( .A(n14556), .B(n14557), .Z(n14308) );
  NOR2_X1 U14418 ( .A1(n9121), .A2(n10064), .ZN(n14557) );
  XNOR2_X1 U14419 ( .A(n14558), .B(n14559), .ZN(n14556) );
  XNOR2_X1 U14420 ( .A(n14560), .B(n14561), .ZN(n14284) );
  XNOR2_X1 U14421 ( .A(n14562), .B(n14563), .ZN(n14561) );
  XOR2_X1 U14422 ( .A(n14564), .B(n14565), .Z(n14277) );
  XNOR2_X1 U14423 ( .A(n14566), .B(n14567), .ZN(n14565) );
  XNOR2_X1 U14424 ( .A(n14568), .B(n14569), .ZN(n14269) );
  XNOR2_X1 U14425 ( .A(n14570), .B(n14571), .ZN(n14568) );
  XNOR2_X1 U14426 ( .A(n14572), .B(n14573), .ZN(n14341) );
  NAND2_X1 U14427 ( .A1(n14574), .A2(n14575), .ZN(n14572) );
  XOR2_X1 U14428 ( .A(n14576), .B(n14577), .Z(n14344) );
  XOR2_X1 U14429 ( .A(n14578), .B(n14579), .Z(n14576) );
  NOR2_X1 U14430 ( .A1(n10054), .A2(n10064), .ZN(n14579) );
  XNOR2_X1 U14431 ( .A(n14580), .B(n14581), .ZN(n14244) );
  XOR2_X1 U14432 ( .A(n14582), .B(n14583), .Z(n14581) );
  NAND2_X1 U14433 ( .A1(b_14_), .A2(a_19_), .ZN(n14583) );
  NAND2_X1 U14434 ( .A1(b_15_), .A2(a_15_), .ZN(n10003) );
  XNOR2_X1 U14435 ( .A(n14584), .B(n14585), .ZN(n14199) );
  XOR2_X1 U14436 ( .A(n14586), .B(n14587), .Z(n14584) );
  XNOR2_X1 U14437 ( .A(n14588), .B(n14589), .ZN(n14163) );
  NAND2_X1 U14438 ( .A1(n14590), .A2(n14591), .ZN(n14588) );
  XNOR2_X1 U14439 ( .A(n14592), .B(n14593), .ZN(n14155) );
  XOR2_X1 U14440 ( .A(n14594), .B(n14595), .Z(n14593) );
  NAND2_X1 U14441 ( .A1(b_14_), .A2(a_6_), .ZN(n14595) );
  XNOR2_X1 U14442 ( .A(n14596), .B(n14597), .ZN(n14148) );
  NAND2_X1 U14443 ( .A1(n14598), .A2(n14599), .ZN(n14596) );
  XNOR2_X1 U14444 ( .A(n14600), .B(n14601), .ZN(n14139) );
  NAND2_X1 U14445 ( .A1(n14602), .A2(n14603), .ZN(n14600) );
  XNOR2_X1 U14446 ( .A(n14604), .B(n14605), .ZN(n14131) );
  NAND2_X1 U14447 ( .A1(n14606), .A2(n14607), .ZN(n14604) );
  XNOR2_X1 U14448 ( .A(n14608), .B(n14609), .ZN(n14123) );
  NAND2_X1 U14449 ( .A1(n14610), .A2(n14611), .ZN(n14608) );
  XNOR2_X1 U14450 ( .A(n14612), .B(n14613), .ZN(n14364) );
  NAND2_X1 U14451 ( .A1(n14614), .A2(n14615), .ZN(n14612) );
  XOR2_X1 U14452 ( .A(n14616), .B(n14617), .Z(n14117) );
  XNOR2_X1 U14453 ( .A(n14618), .B(n14619), .ZN(n14617) );
  XNOR2_X1 U14454 ( .A(n14620), .B(n14621), .ZN(n10216) );
  NAND2_X1 U14455 ( .A1(n10226), .A2(n10225), .ZN(n10224) );
  NOR2_X1 U14456 ( .A1(n14622), .A2(n10266), .ZN(n10225) );
  NOR2_X1 U14457 ( .A1(n14623), .A2(n14624), .ZN(n14622) );
  NOR2_X1 U14458 ( .A1(n14621), .A2(n14620), .ZN(n10226) );
  XNOR2_X1 U14459 ( .A(n14625), .B(n14626), .ZN(n14620) );
  XOR2_X1 U14460 ( .A(n14627), .B(n14628), .Z(n14625) );
  NOR2_X1 U14461 ( .A1(n10093), .A2(n10066), .ZN(n14628) );
  NAND2_X1 U14462 ( .A1(n14629), .A2(n14630), .ZN(n14621) );
  NAND2_X1 U14463 ( .A1(n14616), .A2(n14631), .ZN(n14630) );
  NAND2_X1 U14464 ( .A1(n14619), .A2(n14618), .ZN(n14631) );
  XNOR2_X1 U14465 ( .A(n14632), .B(n14633), .ZN(n14616) );
  XOR2_X1 U14466 ( .A(n14634), .B(n14635), .Z(n14632) );
  NOR2_X1 U14467 ( .A1(n9983), .A2(n10066), .ZN(n14635) );
  INV_X1 U14468 ( .A(n14636), .ZN(n14629) );
  NOR2_X1 U14469 ( .A1(n14618), .A2(n14619), .ZN(n14636) );
  NOR2_X1 U14470 ( .A1(n10064), .A2(n10093), .ZN(n14619) );
  NAND2_X1 U14471 ( .A1(n14614), .A2(n14637), .ZN(n14618) );
  NAND2_X1 U14472 ( .A1(n14613), .A2(n14615), .ZN(n14637) );
  NAND2_X1 U14473 ( .A1(n14638), .A2(n14639), .ZN(n14615) );
  NAND2_X1 U14474 ( .A1(b_14_), .A2(a_1_), .ZN(n14639) );
  INV_X1 U14475 ( .A(n14640), .ZN(n14638) );
  XOR2_X1 U14476 ( .A(n14641), .B(n14642), .Z(n14613) );
  XOR2_X1 U14477 ( .A(n14643), .B(n14644), .Z(n14641) );
  NOR2_X1 U14478 ( .A1(n10088), .A2(n10066), .ZN(n14644) );
  NAND2_X1 U14479 ( .A1(a_1_), .A2(n14640), .ZN(n14614) );
  NAND2_X1 U14480 ( .A1(n14610), .A2(n14645), .ZN(n14640) );
  NAND2_X1 U14481 ( .A1(n14609), .A2(n14611), .ZN(n14645) );
  NAND2_X1 U14482 ( .A1(n14646), .A2(n14647), .ZN(n14611) );
  NAND2_X1 U14483 ( .A1(b_14_), .A2(a_2_), .ZN(n14647) );
  INV_X1 U14484 ( .A(n14648), .ZN(n14646) );
  XOR2_X1 U14485 ( .A(n14649), .B(n14650), .Z(n14609) );
  XOR2_X1 U14486 ( .A(n14651), .B(n14652), .Z(n14649) );
  NOR2_X1 U14487 ( .A1(n10086), .A2(n10066), .ZN(n14652) );
  NAND2_X1 U14488 ( .A1(a_2_), .A2(n14648), .ZN(n14610) );
  NAND2_X1 U14489 ( .A1(n14606), .A2(n14653), .ZN(n14648) );
  NAND2_X1 U14490 ( .A1(n14605), .A2(n14607), .ZN(n14653) );
  NAND2_X1 U14491 ( .A1(n14654), .A2(n14655), .ZN(n14607) );
  NAND2_X1 U14492 ( .A1(b_14_), .A2(a_3_), .ZN(n14655) );
  INV_X1 U14493 ( .A(n14656), .ZN(n14654) );
  XOR2_X1 U14494 ( .A(n14657), .B(n14658), .Z(n14605) );
  XOR2_X1 U14495 ( .A(n14659), .B(n14660), .Z(n14657) );
  NOR2_X1 U14496 ( .A1(n10085), .A2(n10066), .ZN(n14660) );
  NAND2_X1 U14497 ( .A1(a_3_), .A2(n14656), .ZN(n14606) );
  NAND2_X1 U14498 ( .A1(n14602), .A2(n14661), .ZN(n14656) );
  NAND2_X1 U14499 ( .A1(n14601), .A2(n14603), .ZN(n14661) );
  NAND2_X1 U14500 ( .A1(n14662), .A2(n14663), .ZN(n14603) );
  NAND2_X1 U14501 ( .A1(b_14_), .A2(a_4_), .ZN(n14663) );
  INV_X1 U14502 ( .A(n14664), .ZN(n14662) );
  XNOR2_X1 U14503 ( .A(n14665), .B(n14666), .ZN(n14601) );
  XOR2_X1 U14504 ( .A(n14667), .B(n14668), .Z(n14666) );
  NAND2_X1 U14505 ( .A1(b_13_), .A2(a_5_), .ZN(n14668) );
  NAND2_X1 U14506 ( .A1(a_4_), .A2(n14664), .ZN(n14602) );
  NAND2_X1 U14507 ( .A1(n14598), .A2(n14669), .ZN(n14664) );
  NAND2_X1 U14508 ( .A1(n14597), .A2(n14599), .ZN(n14669) );
  NAND2_X1 U14509 ( .A1(n14670), .A2(n14671), .ZN(n14599) );
  NAND2_X1 U14510 ( .A1(b_14_), .A2(a_5_), .ZN(n14671) );
  INV_X1 U14511 ( .A(n14672), .ZN(n14670) );
  XNOR2_X1 U14512 ( .A(n14673), .B(n14674), .ZN(n14597) );
  XOR2_X1 U14513 ( .A(n14675), .B(n14676), .Z(n14674) );
  NAND2_X1 U14514 ( .A1(b_13_), .A2(a_6_), .ZN(n14676) );
  NAND2_X1 U14515 ( .A1(a_5_), .A2(n14672), .ZN(n14598) );
  NAND2_X1 U14516 ( .A1(n14677), .A2(n14678), .ZN(n14672) );
  NAND2_X1 U14517 ( .A1(n14679), .A2(b_14_), .ZN(n14678) );
  NOR2_X1 U14518 ( .A1(n14680), .A2(n10081), .ZN(n14679) );
  NOR2_X1 U14519 ( .A1(n14594), .A2(n14592), .ZN(n14680) );
  NAND2_X1 U14520 ( .A1(n14592), .A2(n14594), .ZN(n14677) );
  NAND2_X1 U14521 ( .A1(n14590), .A2(n14681), .ZN(n14594) );
  NAND2_X1 U14522 ( .A1(n14589), .A2(n14591), .ZN(n14681) );
  NAND2_X1 U14523 ( .A1(n14682), .A2(n14683), .ZN(n14591) );
  NAND2_X1 U14524 ( .A1(b_14_), .A2(a_7_), .ZN(n14682) );
  XNOR2_X1 U14525 ( .A(n14684), .B(n14685), .ZN(n14589) );
  XOR2_X1 U14526 ( .A(n14686), .B(n14687), .Z(n14684) );
  NAND2_X1 U14527 ( .A1(n14688), .A2(a_7_), .ZN(n14590) );
  INV_X1 U14528 ( .A(n14683), .ZN(n14688) );
  NAND2_X1 U14529 ( .A1(n14689), .A2(n14690), .ZN(n14683) );
  NAND2_X1 U14530 ( .A1(n14400), .A2(n14691), .ZN(n14690) );
  NAND2_X1 U14531 ( .A1(n14403), .A2(n14402), .ZN(n14691) );
  XNOR2_X1 U14532 ( .A(n14692), .B(n14693), .ZN(n14400) );
  XOR2_X1 U14533 ( .A(n14694), .B(n14695), .Z(n14692) );
  NOR2_X1 U14534 ( .A1(n10076), .A2(n10066), .ZN(n14695) );
  INV_X1 U14535 ( .A(n14696), .ZN(n14689) );
  NOR2_X1 U14536 ( .A1(n14402), .A2(n14403), .ZN(n14696) );
  NOR2_X1 U14537 ( .A1(n10064), .A2(n10079), .ZN(n14403) );
  NAND2_X1 U14538 ( .A1(n14697), .A2(n14698), .ZN(n14402) );
  NAND2_X1 U14539 ( .A1(n14412), .A2(n14699), .ZN(n14698) );
  NAND2_X1 U14540 ( .A1(n14409), .A2(n14411), .ZN(n14699) );
  NOR2_X1 U14541 ( .A1(n10064), .A2(n10076), .ZN(n14412) );
  INV_X1 U14542 ( .A(n14700), .ZN(n14697) );
  NOR2_X1 U14543 ( .A1(n14411), .A2(n14409), .ZN(n14700) );
  XNOR2_X1 U14544 ( .A(n14701), .B(n14702), .ZN(n14409) );
  XOR2_X1 U14545 ( .A(n14703), .B(n14704), .Z(n14701) );
  NOR2_X1 U14546 ( .A1(n10073), .A2(n10066), .ZN(n14704) );
  NAND2_X1 U14547 ( .A1(n14705), .A2(n14706), .ZN(n14411) );
  NAND2_X1 U14548 ( .A1(n14419), .A2(n14707), .ZN(n14706) );
  NAND2_X1 U14549 ( .A1(n14421), .A2(n14420), .ZN(n14707) );
  XNOR2_X1 U14550 ( .A(n14708), .B(n14709), .ZN(n14419) );
  XNOR2_X1 U14551 ( .A(n14710), .B(n14711), .ZN(n14708) );
  NAND2_X1 U14552 ( .A1(b_13_), .A2(a_11_), .ZN(n14710) );
  INV_X1 U14553 ( .A(n14712), .ZN(n14705) );
  NOR2_X1 U14554 ( .A1(n14420), .A2(n14421), .ZN(n14712) );
  NOR2_X1 U14555 ( .A1(n10064), .A2(n10073), .ZN(n14421) );
  NAND2_X1 U14556 ( .A1(n14713), .A2(n14714), .ZN(n14420) );
  NAND2_X1 U14557 ( .A1(n14429), .A2(n14715), .ZN(n14714) );
  NAND2_X1 U14558 ( .A1(n14426), .A2(n14428), .ZN(n14715) );
  NOR2_X1 U14559 ( .A1(n10064), .A2(n9649), .ZN(n14429) );
  INV_X1 U14560 ( .A(n14716), .ZN(n14713) );
  NOR2_X1 U14561 ( .A1(n14428), .A2(n14426), .ZN(n14716) );
  XNOR2_X1 U14562 ( .A(n14717), .B(n14718), .ZN(n14426) );
  XNOR2_X1 U14563 ( .A(n14719), .B(n14720), .ZN(n14718) );
  NAND2_X1 U14564 ( .A1(b_13_), .A2(a_12_), .ZN(n14720) );
  NAND2_X1 U14565 ( .A1(n14721), .A2(n14722), .ZN(n14428) );
  NAND2_X1 U14566 ( .A1(n14585), .A2(n14723), .ZN(n14722) );
  NAND2_X1 U14567 ( .A1(n14587), .A2(n14586), .ZN(n14723) );
  XNOR2_X1 U14568 ( .A(n14724), .B(n14725), .ZN(n14585) );
  XNOR2_X1 U14569 ( .A(n14726), .B(n10068), .ZN(n14725) );
  INV_X1 U14570 ( .A(n14727), .ZN(n14721) );
  NOR2_X1 U14571 ( .A1(n14586), .A2(n14587), .ZN(n14727) );
  NOR2_X1 U14572 ( .A1(n10064), .A2(n10070), .ZN(n14587) );
  NAND2_X1 U14573 ( .A1(n14728), .A2(n14729), .ZN(n14586) );
  NAND2_X1 U14574 ( .A1(n14441), .A2(n14730), .ZN(n14729) );
  INV_X1 U14575 ( .A(n14731), .ZN(n14730) );
  NOR2_X1 U14576 ( .A1(n14439), .A2(n14440), .ZN(n14731) );
  NOR2_X1 U14577 ( .A1(n10064), .A2(n10067), .ZN(n14441) );
  NAND2_X1 U14578 ( .A1(n14440), .A2(n14439), .ZN(n14728) );
  XNOR2_X1 U14579 ( .A(n14732), .B(n14733), .ZN(n14439) );
  XOR2_X1 U14580 ( .A(n14734), .B(n14735), .Z(n14733) );
  NAND2_X1 U14581 ( .A1(b_13_), .A2(a_14_), .ZN(n14735) );
  NOR2_X1 U14582 ( .A1(n14736), .A2(n14737), .ZN(n14440) );
  INV_X1 U14583 ( .A(n14738), .ZN(n14737) );
  NAND2_X1 U14584 ( .A1(n14447), .A2(n14739), .ZN(n14738) );
  NAND2_X1 U14585 ( .A1(n14449), .A2(n14448), .ZN(n14739) );
  XOR2_X1 U14586 ( .A(n14740), .B(n14741), .Z(n14447) );
  XNOR2_X1 U14587 ( .A(n14742), .B(n14743), .ZN(n14740) );
  NOR2_X1 U14588 ( .A1(n9534), .A2(n10066), .ZN(n14743) );
  NOR2_X1 U14589 ( .A1(n14448), .A2(n14449), .ZN(n14736) );
  NOR2_X1 U14590 ( .A1(n10064), .A2(n10065), .ZN(n14449) );
  NAND2_X1 U14591 ( .A1(n14456), .A2(n14744), .ZN(n14448) );
  NAND2_X1 U14592 ( .A1(n14455), .A2(n14457), .ZN(n14744) );
  NAND2_X1 U14593 ( .A1(n14745), .A2(n14746), .ZN(n14457) );
  NAND2_X1 U14594 ( .A1(b_14_), .A2(a_15_), .ZN(n14746) );
  INV_X1 U14595 ( .A(n14747), .ZN(n14745) );
  XNOR2_X1 U14596 ( .A(n14748), .B(n14749), .ZN(n14455) );
  XOR2_X1 U14597 ( .A(n14750), .B(n14751), .Z(n14748) );
  NAND2_X1 U14598 ( .A1(a_15_), .A2(n14747), .ZN(n14456) );
  NAND2_X1 U14599 ( .A1(n14465), .A2(n14752), .ZN(n14747) );
  NAND2_X1 U14600 ( .A1(n14464), .A2(n14466), .ZN(n14752) );
  NAND2_X1 U14601 ( .A1(n14753), .A2(n14754), .ZN(n14466) );
  NAND2_X1 U14602 ( .A1(b_14_), .A2(a_16_), .ZN(n14754) );
  INV_X1 U14603 ( .A(n14755), .ZN(n14753) );
  XNOR2_X1 U14604 ( .A(n14756), .B(n14757), .ZN(n14464) );
  NAND2_X1 U14605 ( .A1(n14758), .A2(n14759), .ZN(n14756) );
  NAND2_X1 U14606 ( .A1(a_16_), .A2(n14755), .ZN(n14465) );
  NAND2_X1 U14607 ( .A1(n14472), .A2(n14760), .ZN(n14755) );
  NAND2_X1 U14608 ( .A1(n14471), .A2(n14473), .ZN(n14760) );
  NAND2_X1 U14609 ( .A1(n14761), .A2(n14762), .ZN(n14473) );
  NAND2_X1 U14610 ( .A1(b_14_), .A2(a_17_), .ZN(n14762) );
  INV_X1 U14611 ( .A(n14763), .ZN(n14761) );
  XNOR2_X1 U14612 ( .A(n14764), .B(n14765), .ZN(n14471) );
  XOR2_X1 U14613 ( .A(n14766), .B(n14767), .Z(n14765) );
  NAND2_X1 U14614 ( .A1(b_13_), .A2(a_18_), .ZN(n14767) );
  NAND2_X1 U14615 ( .A1(a_17_), .A2(n14763), .ZN(n14472) );
  NAND2_X1 U14616 ( .A1(n14768), .A2(n14769), .ZN(n14763) );
  NAND2_X1 U14617 ( .A1(n14770), .A2(b_14_), .ZN(n14769) );
  NOR2_X1 U14618 ( .A1(n14771), .A2(n10058), .ZN(n14770) );
  NOR2_X1 U14619 ( .A1(n14479), .A2(n14481), .ZN(n14771) );
  NAND2_X1 U14620 ( .A1(n14479), .A2(n14481), .ZN(n14768) );
  NAND2_X1 U14621 ( .A1(n14772), .A2(n14773), .ZN(n14481) );
  NAND2_X1 U14622 ( .A1(n14774), .A2(b_14_), .ZN(n14773) );
  NOR2_X1 U14623 ( .A1(n14775), .A2(n9415), .ZN(n14774) );
  NOR2_X1 U14624 ( .A1(n14580), .A2(n14582), .ZN(n14775) );
  NAND2_X1 U14625 ( .A1(n14580), .A2(n14582), .ZN(n14772) );
  NAND2_X1 U14626 ( .A1(n14776), .A2(n14777), .ZN(n14582) );
  NAND2_X1 U14627 ( .A1(n14778), .A2(b_14_), .ZN(n14777) );
  NOR2_X1 U14628 ( .A1(n14779), .A2(n10054), .ZN(n14778) );
  NOR2_X1 U14629 ( .A1(n14578), .A2(n14577), .ZN(n14779) );
  NAND2_X1 U14630 ( .A1(n14577), .A2(n14578), .ZN(n14776) );
  NAND2_X1 U14631 ( .A1(n14574), .A2(n14780), .ZN(n14578) );
  NAND2_X1 U14632 ( .A1(n14573), .A2(n14575), .ZN(n14780) );
  NAND2_X1 U14633 ( .A1(n14781), .A2(n14782), .ZN(n14575) );
  NAND2_X1 U14634 ( .A1(b_14_), .A2(a_21_), .ZN(n14782) );
  INV_X1 U14635 ( .A(n14783), .ZN(n14781) );
  XNOR2_X1 U14636 ( .A(n14784), .B(n14785), .ZN(n14573) );
  XOR2_X1 U14637 ( .A(n14786), .B(n14787), .Z(n14785) );
  NAND2_X1 U14638 ( .A1(a_21_), .A2(n14783), .ZN(n14574) );
  NAND2_X1 U14639 ( .A1(n14788), .A2(n14789), .ZN(n14783) );
  NAND2_X1 U14640 ( .A1(n14502), .A2(n14790), .ZN(n14789) );
  NAND2_X1 U14641 ( .A1(n14501), .A2(n14500), .ZN(n14790) );
  NOR2_X1 U14642 ( .A1(n10064), .A2(n9330), .ZN(n14502) );
  INV_X1 U14643 ( .A(n14791), .ZN(n14788) );
  NOR2_X1 U14644 ( .A1(n14500), .A2(n14501), .ZN(n14791) );
  NOR2_X1 U14645 ( .A1(n14792), .A2(n14793), .ZN(n14501) );
  INV_X1 U14646 ( .A(n14794), .ZN(n14793) );
  NAND2_X1 U14647 ( .A1(n14571), .A2(n14795), .ZN(n14794) );
  NAND2_X1 U14648 ( .A1(n14569), .A2(n14570), .ZN(n14795) );
  NOR2_X1 U14649 ( .A1(n10064), .A2(n10051), .ZN(n14571) );
  NOR2_X1 U14650 ( .A1(n14569), .A2(n14570), .ZN(n14792) );
  NOR2_X1 U14651 ( .A1(n14796), .A2(n14797), .ZN(n14570) );
  NOR2_X1 U14652 ( .A1(n14567), .A2(n14798), .ZN(n14797) );
  NOR2_X1 U14653 ( .A1(n14799), .A2(n14800), .ZN(n14798) );
  INV_X1 U14654 ( .A(n14564), .ZN(n14800) );
  INV_X1 U14655 ( .A(n14566), .ZN(n14799) );
  NAND2_X1 U14656 ( .A1(b_14_), .A2(a_24_), .ZN(n14567) );
  NOR2_X1 U14657 ( .A1(n14564), .A2(n14566), .ZN(n14796) );
  NOR2_X1 U14658 ( .A1(n14801), .A2(n14802), .ZN(n14566) );
  INV_X1 U14659 ( .A(n14803), .ZN(n14802) );
  NAND2_X1 U14660 ( .A1(n14563), .A2(n14804), .ZN(n14803) );
  NAND2_X1 U14661 ( .A1(n14560), .A2(n14562), .ZN(n14804) );
  NOR2_X1 U14662 ( .A1(n10064), .A2(n10048), .ZN(n14563) );
  NOR2_X1 U14663 ( .A1(n14560), .A2(n14562), .ZN(n14801) );
  NAND2_X1 U14664 ( .A1(n14805), .A2(n14806), .ZN(n14562) );
  NAND2_X1 U14665 ( .A1(n14520), .A2(n14807), .ZN(n14806) );
  NAND2_X1 U14666 ( .A1(n14523), .A2(n14522), .ZN(n14807) );
  XOR2_X1 U14667 ( .A(n14808), .B(n14809), .Z(n14520) );
  NAND2_X1 U14668 ( .A1(n14810), .A2(n14811), .ZN(n14808) );
  INV_X1 U14669 ( .A(n14812), .ZN(n14805) );
  NOR2_X1 U14670 ( .A1(n14522), .A2(n14523), .ZN(n14812) );
  NOR2_X1 U14671 ( .A1(n10064), .A2(n10047), .ZN(n14523) );
  NAND2_X1 U14672 ( .A1(n14529), .A2(n14813), .ZN(n14522) );
  NAND2_X1 U14673 ( .A1(n14528), .A2(n14530), .ZN(n14813) );
  NAND2_X1 U14674 ( .A1(n14814), .A2(n14815), .ZN(n14530) );
  NAND2_X1 U14675 ( .A1(b_14_), .A2(a_27_), .ZN(n14815) );
  INV_X1 U14676 ( .A(n14816), .ZN(n14814) );
  XNOR2_X1 U14677 ( .A(n14817), .B(n14818), .ZN(n14528) );
  XOR2_X1 U14678 ( .A(n14819), .B(n14820), .Z(n14818) );
  NAND2_X1 U14679 ( .A1(b_13_), .A2(a_28_), .ZN(n14820) );
  NAND2_X1 U14680 ( .A1(a_27_), .A2(n14816), .ZN(n14529) );
  NAND2_X1 U14681 ( .A1(n14821), .A2(n14822), .ZN(n14816) );
  NAND2_X1 U14682 ( .A1(n14823), .A2(b_14_), .ZN(n14822) );
  NOR2_X1 U14683 ( .A1(n14824), .A2(n9136), .ZN(n14823) );
  NOR2_X1 U14684 ( .A1(n14536), .A2(n14538), .ZN(n14824) );
  NAND2_X1 U14685 ( .A1(n14536), .A2(n14538), .ZN(n14821) );
  NAND2_X1 U14686 ( .A1(n14825), .A2(n14826), .ZN(n14538) );
  NAND2_X1 U14687 ( .A1(n14827), .A2(b_14_), .ZN(n14826) );
  NOR2_X1 U14688 ( .A1(n14828), .A2(n9121), .ZN(n14827) );
  NOR2_X1 U14689 ( .A1(n14829), .A2(n14558), .ZN(n14828) );
  NAND2_X1 U14690 ( .A1(n14829), .A2(n14558), .ZN(n14825) );
  NAND2_X1 U14691 ( .A1(n14830), .A2(n14831), .ZN(n14558) );
  NAND2_X1 U14692 ( .A1(b_12_), .A2(n14832), .ZN(n14831) );
  NAND2_X1 U14693 ( .A1(n10486), .A2(n14833), .ZN(n14832) );
  NAND2_X1 U14694 ( .A1(a_31_), .A2(n10066), .ZN(n14833) );
  NAND2_X1 U14695 ( .A1(b_13_), .A2(n14834), .ZN(n14830) );
  NAND2_X1 U14696 ( .A1(n10489), .A2(n14835), .ZN(n14834) );
  NAND2_X1 U14697 ( .A1(a_30_), .A2(n10069), .ZN(n14835) );
  INV_X1 U14698 ( .A(n14559), .ZN(n14829) );
  NAND2_X1 U14699 ( .A1(n14836), .A2(n9025), .ZN(n14559) );
  NOR2_X1 U14700 ( .A1(n10064), .A2(n10066), .ZN(n14836) );
  XOR2_X1 U14701 ( .A(n14837), .B(n14838), .Z(n14536) );
  NOR2_X1 U14702 ( .A1(n9121), .A2(n10066), .ZN(n14838) );
  XNOR2_X1 U14703 ( .A(n14839), .B(n14840), .ZN(n14837) );
  XNOR2_X1 U14704 ( .A(n14841), .B(n14842), .ZN(n14560) );
  XNOR2_X1 U14705 ( .A(n14843), .B(n14844), .ZN(n14842) );
  XNOR2_X1 U14706 ( .A(n14845), .B(n14846), .ZN(n14564) );
  XOR2_X1 U14707 ( .A(n14847), .B(n14848), .Z(n14846) );
  XOR2_X1 U14708 ( .A(n14849), .B(n14850), .Z(n14569) );
  XOR2_X1 U14709 ( .A(n14851), .B(n14852), .Z(n14850) );
  XNOR2_X1 U14710 ( .A(n14853), .B(n14854), .ZN(n14500) );
  XOR2_X1 U14711 ( .A(n14855), .B(n14856), .Z(n14853) );
  XNOR2_X1 U14712 ( .A(n14857), .B(n14858), .ZN(n14577) );
  NAND2_X1 U14713 ( .A1(n14859), .A2(n14860), .ZN(n14857) );
  XOR2_X1 U14714 ( .A(n14861), .B(n14862), .Z(n14580) );
  XOR2_X1 U14715 ( .A(n14863), .B(n14864), .Z(n14861) );
  NOR2_X1 U14716 ( .A1(n10054), .A2(n10066), .ZN(n14864) );
  XNOR2_X1 U14717 ( .A(n14865), .B(n14866), .ZN(n14479) );
  XOR2_X1 U14718 ( .A(n14867), .B(n14868), .Z(n14866) );
  NAND2_X1 U14719 ( .A1(b_13_), .A2(a_19_), .ZN(n14868) );
  XOR2_X1 U14720 ( .A(n14869), .B(n14870), .Z(n14592) );
  XNOR2_X1 U14721 ( .A(n14871), .B(n14872), .ZN(n14870) );
  NAND2_X1 U14722 ( .A1(b_13_), .A2(a_7_), .ZN(n14872) );
  INV_X1 U14723 ( .A(n14873), .ZN(n10266) );
  NAND2_X1 U14724 ( .A1(n14623), .A2(n14624), .ZN(n14873) );
  NAND2_X1 U14725 ( .A1(n14874), .A2(n14875), .ZN(n14624) );
  NAND2_X1 U14726 ( .A1(n14876), .A2(b_13_), .ZN(n14875) );
  NOR2_X1 U14727 ( .A1(n14877), .A2(n10093), .ZN(n14876) );
  NOR2_X1 U14728 ( .A1(n14626), .A2(n14627), .ZN(n14877) );
  NAND2_X1 U14729 ( .A1(n14626), .A2(n14627), .ZN(n14874) );
  NAND2_X1 U14730 ( .A1(n14878), .A2(n14879), .ZN(n14627) );
  NAND2_X1 U14731 ( .A1(n14880), .A2(b_13_), .ZN(n14879) );
  NOR2_X1 U14732 ( .A1(n14881), .A2(n9983), .ZN(n14880) );
  NOR2_X1 U14733 ( .A1(n14633), .A2(n14634), .ZN(n14881) );
  NAND2_X1 U14734 ( .A1(n14633), .A2(n14634), .ZN(n14878) );
  NAND2_X1 U14735 ( .A1(n14882), .A2(n14883), .ZN(n14634) );
  NAND2_X1 U14736 ( .A1(n14884), .A2(b_13_), .ZN(n14883) );
  NOR2_X1 U14737 ( .A1(n14885), .A2(n10088), .ZN(n14884) );
  NOR2_X1 U14738 ( .A1(n14642), .A2(n14643), .ZN(n14885) );
  NAND2_X1 U14739 ( .A1(n14642), .A2(n14643), .ZN(n14882) );
  NAND2_X1 U14740 ( .A1(n14886), .A2(n14887), .ZN(n14643) );
  NAND2_X1 U14741 ( .A1(n14888), .A2(b_13_), .ZN(n14887) );
  NOR2_X1 U14742 ( .A1(n14889), .A2(n10086), .ZN(n14888) );
  NOR2_X1 U14743 ( .A1(n14650), .A2(n14651), .ZN(n14889) );
  NAND2_X1 U14744 ( .A1(n14650), .A2(n14651), .ZN(n14886) );
  NAND2_X1 U14745 ( .A1(n14890), .A2(n14891), .ZN(n14651) );
  NAND2_X1 U14746 ( .A1(n14892), .A2(b_13_), .ZN(n14891) );
  NOR2_X1 U14747 ( .A1(n14893), .A2(n10085), .ZN(n14892) );
  NOR2_X1 U14748 ( .A1(n14658), .A2(n14659), .ZN(n14893) );
  NAND2_X1 U14749 ( .A1(n14658), .A2(n14659), .ZN(n14890) );
  NAND2_X1 U14750 ( .A1(n14894), .A2(n14895), .ZN(n14659) );
  NAND2_X1 U14751 ( .A1(n14896), .A2(b_13_), .ZN(n14895) );
  NOR2_X1 U14752 ( .A1(n14897), .A2(n10083), .ZN(n14896) );
  NOR2_X1 U14753 ( .A1(n14665), .A2(n14667), .ZN(n14897) );
  NAND2_X1 U14754 ( .A1(n14665), .A2(n14667), .ZN(n14894) );
  NAND2_X1 U14755 ( .A1(n14898), .A2(n14899), .ZN(n14667) );
  NAND2_X1 U14756 ( .A1(n14900), .A2(b_13_), .ZN(n14899) );
  NOR2_X1 U14757 ( .A1(n14901), .A2(n10081), .ZN(n14900) );
  NOR2_X1 U14758 ( .A1(n14673), .A2(n14675), .ZN(n14901) );
  NAND2_X1 U14759 ( .A1(n14673), .A2(n14675), .ZN(n14898) );
  NAND2_X1 U14760 ( .A1(n14902), .A2(n14903), .ZN(n14675) );
  NAND2_X1 U14761 ( .A1(n14904), .A2(b_13_), .ZN(n14903) );
  NOR2_X1 U14762 ( .A1(n14905), .A2(n9773), .ZN(n14904) );
  NOR2_X1 U14763 ( .A1(n14871), .A2(n14869), .ZN(n14905) );
  NAND2_X1 U14764 ( .A1(n14871), .A2(n14869), .ZN(n14902) );
  XNOR2_X1 U14765 ( .A(n14906), .B(n14907), .ZN(n14869) );
  NAND2_X1 U14766 ( .A1(n14908), .A2(n14909), .ZN(n14906) );
  NOR2_X1 U14767 ( .A1(n14910), .A2(n14911), .ZN(n14871) );
  INV_X1 U14768 ( .A(n14912), .ZN(n14911) );
  NAND2_X1 U14769 ( .A1(n14685), .A2(n14913), .ZN(n14912) );
  NAND2_X1 U14770 ( .A1(n14687), .A2(n14686), .ZN(n14913) );
  XOR2_X1 U14771 ( .A(n14914), .B(n14915), .Z(n14685) );
  NAND2_X1 U14772 ( .A1(n14916), .A2(n14917), .ZN(n14914) );
  NOR2_X1 U14773 ( .A1(n14686), .A2(n14687), .ZN(n14910) );
  NOR2_X1 U14774 ( .A1(n10066), .A2(n10079), .ZN(n14687) );
  NAND2_X1 U14775 ( .A1(n14918), .A2(n14919), .ZN(n14686) );
  NAND2_X1 U14776 ( .A1(n14920), .A2(b_13_), .ZN(n14919) );
  NOR2_X1 U14777 ( .A1(n14921), .A2(n10076), .ZN(n14920) );
  NOR2_X1 U14778 ( .A1(n14693), .A2(n14694), .ZN(n14921) );
  NAND2_X1 U14779 ( .A1(n14693), .A2(n14694), .ZN(n14918) );
  NAND2_X1 U14780 ( .A1(n14922), .A2(n14923), .ZN(n14694) );
  NAND2_X1 U14781 ( .A1(n14924), .A2(b_13_), .ZN(n14923) );
  NOR2_X1 U14782 ( .A1(n14925), .A2(n10073), .ZN(n14924) );
  NOR2_X1 U14783 ( .A1(n14702), .A2(n14703), .ZN(n14925) );
  NAND2_X1 U14784 ( .A1(n14702), .A2(n14703), .ZN(n14922) );
  NAND2_X1 U14785 ( .A1(n14926), .A2(n14927), .ZN(n14703) );
  NAND2_X1 U14786 ( .A1(n14928), .A2(b_13_), .ZN(n14927) );
  NOR2_X1 U14787 ( .A1(n14929), .A2(n9649), .ZN(n14928) );
  NOR2_X1 U14788 ( .A1(n14709), .A2(n14711), .ZN(n14929) );
  NAND2_X1 U14789 ( .A1(n14709), .A2(n14711), .ZN(n14926) );
  NAND2_X1 U14790 ( .A1(n14930), .A2(n14931), .ZN(n14711) );
  NAND2_X1 U14791 ( .A1(n14932), .A2(b_13_), .ZN(n14931) );
  NOR2_X1 U14792 ( .A1(n14933), .A2(n10070), .ZN(n14932) );
  NOR2_X1 U14793 ( .A1(n14719), .A2(n14717), .ZN(n14933) );
  NAND2_X1 U14794 ( .A1(n14719), .A2(n14717), .ZN(n14930) );
  XOR2_X1 U14795 ( .A(n14934), .B(n14935), .Z(n14717) );
  XNOR2_X1 U14796 ( .A(n14936), .B(n14937), .ZN(n14935) );
  NOR2_X1 U14797 ( .A1(n14938), .A2(n14939), .ZN(n14719) );
  INV_X1 U14798 ( .A(n14940), .ZN(n14939) );
  NAND2_X1 U14799 ( .A1(n14724), .A2(n14941), .ZN(n14940) );
  NAND2_X1 U14800 ( .A1(n10068), .A2(n14726), .ZN(n14941) );
  XOR2_X1 U14801 ( .A(n14942), .B(n14943), .Z(n14724) );
  NAND2_X1 U14802 ( .A1(n14944), .A2(n14945), .ZN(n14942) );
  NOR2_X1 U14803 ( .A1(n14726), .A2(n10068), .ZN(n14938) );
  NOR2_X1 U14804 ( .A1(n10066), .A2(n10067), .ZN(n10068) );
  NAND2_X1 U14805 ( .A1(n14946), .A2(n14947), .ZN(n14726) );
  NAND2_X1 U14806 ( .A1(n14948), .A2(b_13_), .ZN(n14947) );
  NOR2_X1 U14807 ( .A1(n14949), .A2(n10065), .ZN(n14948) );
  NOR2_X1 U14808 ( .A1(n14732), .A2(n14734), .ZN(n14949) );
  NAND2_X1 U14809 ( .A1(n14732), .A2(n14734), .ZN(n14946) );
  NAND2_X1 U14810 ( .A1(n14950), .A2(n14951), .ZN(n14734) );
  NAND2_X1 U14811 ( .A1(n14952), .A2(b_13_), .ZN(n14951) );
  NOR2_X1 U14812 ( .A1(n14953), .A2(n9534), .ZN(n14952) );
  NOR2_X1 U14813 ( .A1(n14742), .A2(n14741), .ZN(n14953) );
  NAND2_X1 U14814 ( .A1(n14742), .A2(n14741), .ZN(n14950) );
  XNOR2_X1 U14815 ( .A(n14954), .B(n14955), .ZN(n14741) );
  NAND2_X1 U14816 ( .A1(n14956), .A2(n14957), .ZN(n14954) );
  NOR2_X1 U14817 ( .A1(n14958), .A2(n14959), .ZN(n14742) );
  INV_X1 U14818 ( .A(n14960), .ZN(n14959) );
  NAND2_X1 U14819 ( .A1(n14749), .A2(n14961), .ZN(n14960) );
  NAND2_X1 U14820 ( .A1(n14751), .A2(n14750), .ZN(n14961) );
  XOR2_X1 U14821 ( .A(n14962), .B(n14963), .Z(n14749) );
  XOR2_X1 U14822 ( .A(n14964), .B(n14965), .Z(n14963) );
  NAND2_X1 U14823 ( .A1(b_12_), .A2(a_17_), .ZN(n14965) );
  NOR2_X1 U14824 ( .A1(n14750), .A2(n14751), .ZN(n14958) );
  NOR2_X1 U14825 ( .A1(n10066), .A2(n10062), .ZN(n14751) );
  NAND2_X1 U14826 ( .A1(n14758), .A2(n14966), .ZN(n14750) );
  NAND2_X1 U14827 ( .A1(n14757), .A2(n14759), .ZN(n14966) );
  NAND2_X1 U14828 ( .A1(n14967), .A2(n14968), .ZN(n14759) );
  NAND2_X1 U14829 ( .A1(b_13_), .A2(a_17_), .ZN(n14968) );
  INV_X1 U14830 ( .A(n14969), .ZN(n14967) );
  XNOR2_X1 U14831 ( .A(n14970), .B(n14971), .ZN(n14757) );
  XOR2_X1 U14832 ( .A(n14972), .B(n14973), .Z(n14971) );
  NAND2_X1 U14833 ( .A1(b_12_), .A2(a_18_), .ZN(n14973) );
  NAND2_X1 U14834 ( .A1(a_17_), .A2(n14969), .ZN(n14758) );
  NAND2_X1 U14835 ( .A1(n14974), .A2(n14975), .ZN(n14969) );
  NAND2_X1 U14836 ( .A1(n14976), .A2(b_13_), .ZN(n14975) );
  NOR2_X1 U14837 ( .A1(n14977), .A2(n10058), .ZN(n14976) );
  NOR2_X1 U14838 ( .A1(n14764), .A2(n14766), .ZN(n14977) );
  NAND2_X1 U14839 ( .A1(n14764), .A2(n14766), .ZN(n14974) );
  NAND2_X1 U14840 ( .A1(n14978), .A2(n14979), .ZN(n14766) );
  NAND2_X1 U14841 ( .A1(n14980), .A2(b_13_), .ZN(n14979) );
  NOR2_X1 U14842 ( .A1(n14981), .A2(n9415), .ZN(n14980) );
  NOR2_X1 U14843 ( .A1(n14865), .A2(n14867), .ZN(n14981) );
  NAND2_X1 U14844 ( .A1(n14865), .A2(n14867), .ZN(n14978) );
  NAND2_X1 U14845 ( .A1(n14982), .A2(n14983), .ZN(n14867) );
  NAND2_X1 U14846 ( .A1(n14984), .A2(b_13_), .ZN(n14983) );
  NOR2_X1 U14847 ( .A1(n14985), .A2(n10054), .ZN(n14984) );
  NOR2_X1 U14848 ( .A1(n14862), .A2(n14863), .ZN(n14985) );
  NAND2_X1 U14849 ( .A1(n14862), .A2(n14863), .ZN(n14982) );
  NAND2_X1 U14850 ( .A1(n14859), .A2(n14986), .ZN(n14863) );
  NAND2_X1 U14851 ( .A1(n14858), .A2(n14860), .ZN(n14986) );
  NAND2_X1 U14852 ( .A1(n14987), .A2(n14988), .ZN(n14860) );
  NAND2_X1 U14853 ( .A1(b_13_), .A2(a_21_), .ZN(n14988) );
  INV_X1 U14854 ( .A(n14989), .ZN(n14987) );
  XOR2_X1 U14855 ( .A(n14990), .B(n14991), .Z(n14858) );
  XOR2_X1 U14856 ( .A(n14992), .B(n14993), .Z(n14990) );
  NAND2_X1 U14857 ( .A1(a_21_), .A2(n14989), .ZN(n14859) );
  NAND2_X1 U14858 ( .A1(n14994), .A2(n14995), .ZN(n14989) );
  INV_X1 U14859 ( .A(n14996), .ZN(n14995) );
  NOR2_X1 U14860 ( .A1(n14787), .A2(n14997), .ZN(n14996) );
  NOR2_X1 U14861 ( .A1(n14786), .A2(n14784), .ZN(n14997) );
  NAND2_X1 U14862 ( .A1(b_13_), .A2(a_22_), .ZN(n14787) );
  NAND2_X1 U14863 ( .A1(n14784), .A2(n14786), .ZN(n14994) );
  NAND2_X1 U14864 ( .A1(n14998), .A2(n14999), .ZN(n14786) );
  NAND2_X1 U14865 ( .A1(n14856), .A2(n15000), .ZN(n14999) );
  INV_X1 U14866 ( .A(n15001), .ZN(n15000) );
  NOR2_X1 U14867 ( .A1(n14855), .A2(n14854), .ZN(n15001) );
  NOR2_X1 U14868 ( .A1(n10066), .A2(n10051), .ZN(n14856) );
  NAND2_X1 U14869 ( .A1(n14854), .A2(n14855), .ZN(n14998) );
  NAND2_X1 U14870 ( .A1(n15002), .A2(n15003), .ZN(n14855) );
  INV_X1 U14871 ( .A(n15004), .ZN(n15003) );
  NOR2_X1 U14872 ( .A1(n14852), .A2(n15005), .ZN(n15004) );
  NOR2_X1 U14873 ( .A1(n14851), .A2(n14849), .ZN(n15005) );
  NAND2_X1 U14874 ( .A1(b_13_), .A2(a_24_), .ZN(n14852) );
  NAND2_X1 U14875 ( .A1(n14849), .A2(n14851), .ZN(n15002) );
  NAND2_X1 U14876 ( .A1(n15006), .A2(n15007), .ZN(n14851) );
  NAND2_X1 U14877 ( .A1(n14848), .A2(n15008), .ZN(n15007) );
  INV_X1 U14878 ( .A(n15009), .ZN(n15008) );
  NOR2_X1 U14879 ( .A1(n14845), .A2(n14847), .ZN(n15009) );
  NOR2_X1 U14880 ( .A1(n10066), .A2(n10048), .ZN(n14848) );
  NAND2_X1 U14881 ( .A1(n14847), .A2(n14845), .ZN(n15006) );
  XOR2_X1 U14882 ( .A(n15010), .B(n15011), .Z(n14845) );
  XNOR2_X1 U14883 ( .A(n15012), .B(n15013), .ZN(n15011) );
  NOR2_X1 U14884 ( .A1(n15014), .A2(n15015), .ZN(n14847) );
  INV_X1 U14885 ( .A(n15016), .ZN(n15015) );
  NAND2_X1 U14886 ( .A1(n14841), .A2(n15017), .ZN(n15016) );
  NAND2_X1 U14887 ( .A1(n14844), .A2(n14843), .ZN(n15017) );
  XOR2_X1 U14888 ( .A(n15018), .B(n15019), .Z(n14841) );
  NAND2_X1 U14889 ( .A1(n15020), .A2(n15021), .ZN(n15018) );
  NOR2_X1 U14890 ( .A1(n14843), .A2(n14844), .ZN(n15014) );
  NOR2_X1 U14891 ( .A1(n10066), .A2(n10047), .ZN(n14844) );
  NAND2_X1 U14892 ( .A1(n14810), .A2(n15022), .ZN(n14843) );
  NAND2_X1 U14893 ( .A1(n14809), .A2(n14811), .ZN(n15022) );
  NAND2_X1 U14894 ( .A1(n15023), .A2(n15024), .ZN(n14811) );
  NAND2_X1 U14895 ( .A1(b_13_), .A2(a_27_), .ZN(n15024) );
  INV_X1 U14896 ( .A(n15025), .ZN(n15023) );
  XNOR2_X1 U14897 ( .A(n15026), .B(n15027), .ZN(n14809) );
  XOR2_X1 U14898 ( .A(n15028), .B(n15029), .Z(n15027) );
  NAND2_X1 U14899 ( .A1(b_12_), .A2(a_28_), .ZN(n15029) );
  NAND2_X1 U14900 ( .A1(a_27_), .A2(n15025), .ZN(n14810) );
  NAND2_X1 U14901 ( .A1(n15030), .A2(n15031), .ZN(n15025) );
  NAND2_X1 U14902 ( .A1(n15032), .A2(b_13_), .ZN(n15031) );
  NOR2_X1 U14903 ( .A1(n15033), .A2(n9136), .ZN(n15032) );
  NOR2_X1 U14904 ( .A1(n14817), .A2(n14819), .ZN(n15033) );
  NAND2_X1 U14905 ( .A1(n14817), .A2(n14819), .ZN(n15030) );
  NAND2_X1 U14906 ( .A1(n15034), .A2(n15035), .ZN(n14819) );
  NAND2_X1 U14907 ( .A1(n15036), .A2(b_13_), .ZN(n15035) );
  NOR2_X1 U14908 ( .A1(n15037), .A2(n9121), .ZN(n15036) );
  NOR2_X1 U14909 ( .A1(n15038), .A2(n14839), .ZN(n15037) );
  NAND2_X1 U14910 ( .A1(n15038), .A2(n14839), .ZN(n15034) );
  NAND2_X1 U14911 ( .A1(n15039), .A2(n15040), .ZN(n14839) );
  NAND2_X1 U14912 ( .A1(b_11_), .A2(n15041), .ZN(n15040) );
  NAND2_X1 U14913 ( .A1(n10486), .A2(n15042), .ZN(n15041) );
  NAND2_X1 U14914 ( .A1(a_31_), .A2(n10069), .ZN(n15042) );
  NAND2_X1 U14915 ( .A1(b_12_), .A2(n15043), .ZN(n15039) );
  NAND2_X1 U14916 ( .A1(n10489), .A2(n15044), .ZN(n15043) );
  NAND2_X1 U14917 ( .A1(a_30_), .A2(n10071), .ZN(n15044) );
  INV_X1 U14918 ( .A(n14840), .ZN(n15038) );
  NAND2_X1 U14919 ( .A1(n15045), .A2(n9025), .ZN(n14840) );
  NOR2_X1 U14920 ( .A1(n10066), .A2(n10069), .ZN(n15045) );
  XOR2_X1 U14921 ( .A(n15046), .B(n15047), .Z(n14817) );
  NOR2_X1 U14922 ( .A1(n9121), .A2(n10069), .ZN(n15047) );
  XNOR2_X1 U14923 ( .A(n15048), .B(n15049), .ZN(n15046) );
  XOR2_X1 U14924 ( .A(n15050), .B(n15051), .Z(n14849) );
  XOR2_X1 U14925 ( .A(n15052), .B(n15053), .Z(n15051) );
  XNOR2_X1 U14926 ( .A(n15054), .B(n15055), .ZN(n14854) );
  XOR2_X1 U14927 ( .A(n15056), .B(n15057), .Z(n15055) );
  XOR2_X1 U14928 ( .A(n15058), .B(n15059), .Z(n14784) );
  XOR2_X1 U14929 ( .A(n15060), .B(n15061), .Z(n15058) );
  XNOR2_X1 U14930 ( .A(n15062), .B(n15063), .ZN(n14862) );
  NAND2_X1 U14931 ( .A1(n15064), .A2(n15065), .ZN(n15062) );
  XOR2_X1 U14932 ( .A(n15066), .B(n15067), .Z(n14865) );
  XOR2_X1 U14933 ( .A(n15068), .B(n15069), .Z(n15066) );
  NOR2_X1 U14934 ( .A1(n10054), .A2(n10069), .ZN(n15069) );
  XNOR2_X1 U14935 ( .A(n15070), .B(n15071), .ZN(n14764) );
  XOR2_X1 U14936 ( .A(n15072), .B(n15073), .Z(n15071) );
  NAND2_X1 U14937 ( .A1(b_12_), .A2(a_19_), .ZN(n15073) );
  XOR2_X1 U14938 ( .A(n15074), .B(n15075), .Z(n14732) );
  XOR2_X1 U14939 ( .A(n15076), .B(n15077), .Z(n15074) );
  NOR2_X1 U14940 ( .A1(n9534), .A2(n10069), .ZN(n15077) );
  XNOR2_X1 U14941 ( .A(n15078), .B(n15079), .ZN(n14709) );
  XOR2_X1 U14942 ( .A(n15080), .B(n9627), .Z(n15079) );
  XOR2_X1 U14943 ( .A(n15081), .B(n15082), .Z(n14702) );
  XOR2_X1 U14944 ( .A(n15083), .B(n15084), .Z(n15082) );
  XNOR2_X1 U14945 ( .A(n15085), .B(n15086), .ZN(n14693) );
  NAND2_X1 U14946 ( .A1(n15087), .A2(n15088), .ZN(n15085) );
  XNOR2_X1 U14947 ( .A(n15089), .B(n15090), .ZN(n14673) );
  NAND2_X1 U14948 ( .A1(n15091), .A2(n15092), .ZN(n15089) );
  XNOR2_X1 U14949 ( .A(n15093), .B(n15094), .ZN(n14665) );
  NAND2_X1 U14950 ( .A1(n15095), .A2(n15096), .ZN(n15093) );
  XNOR2_X1 U14951 ( .A(n15097), .B(n15098), .ZN(n14658) );
  NAND2_X1 U14952 ( .A1(n15099), .A2(n15100), .ZN(n15097) );
  XNOR2_X1 U14953 ( .A(n15101), .B(n15102), .ZN(n14650) );
  NAND2_X1 U14954 ( .A1(n15103), .A2(n15104), .ZN(n15101) );
  XNOR2_X1 U14955 ( .A(n15105), .B(n15106), .ZN(n14642) );
  NAND2_X1 U14956 ( .A1(n15107), .A2(n15108), .ZN(n15105) );
  XNOR2_X1 U14957 ( .A(n15109), .B(n15110), .ZN(n14633) );
  NAND2_X1 U14958 ( .A1(n15111), .A2(n15112), .ZN(n15109) );
  XOR2_X1 U14959 ( .A(n15113), .B(n15114), .Z(n14626) );
  XNOR2_X1 U14960 ( .A(n15115), .B(n15116), .ZN(n15114) );
  XNOR2_X1 U14961 ( .A(n15117), .B(n15118), .ZN(n14623) );
  XNOR2_X1 U14962 ( .A(n15119), .B(n15120), .ZN(n15118) );
  XNOR2_X1 U14963 ( .A(n15121), .B(n15122), .ZN(n10230) );
  NAND2_X1 U14964 ( .A1(n10239), .A2(n10238), .ZN(n10237) );
  NOR2_X1 U14965 ( .A1(n15123), .A2(n10263), .ZN(n10238) );
  NOR2_X1 U14966 ( .A1(n15124), .A2(n15125), .ZN(n15123) );
  INV_X1 U14967 ( .A(n15126), .ZN(n10239) );
  NAND2_X1 U14968 ( .A1(n15122), .A2(n15121), .ZN(n15126) );
  NAND2_X1 U14969 ( .A1(n15127), .A2(n15128), .ZN(n15121) );
  NAND2_X1 U14970 ( .A1(n15120), .A2(n15129), .ZN(n15128) );
  NAND2_X1 U14971 ( .A1(n15117), .A2(n15119), .ZN(n15129) );
  NOR2_X1 U14972 ( .A1(n10069), .A2(n10093), .ZN(n15120) );
  INV_X1 U14973 ( .A(n15130), .ZN(n15127) );
  NOR2_X1 U14974 ( .A1(n15119), .A2(n15117), .ZN(n15130) );
  XNOR2_X1 U14975 ( .A(n15131), .B(n15132), .ZN(n15117) );
  XOR2_X1 U14976 ( .A(n15133), .B(n15134), .Z(n15131) );
  NOR2_X1 U14977 ( .A1(n10071), .A2(n9983), .ZN(n15134) );
  NAND2_X1 U14978 ( .A1(n15135), .A2(n15136), .ZN(n15119) );
  NAND2_X1 U14979 ( .A1(n15113), .A2(n15137), .ZN(n15136) );
  NAND2_X1 U14980 ( .A1(n15116), .A2(n15115), .ZN(n15137) );
  XNOR2_X1 U14981 ( .A(n15138), .B(n15139), .ZN(n15113) );
  XOR2_X1 U14982 ( .A(n15140), .B(n15141), .Z(n15138) );
  NOR2_X1 U14983 ( .A1(n10071), .A2(n10088), .ZN(n15141) );
  INV_X1 U14984 ( .A(n15142), .ZN(n15135) );
  NOR2_X1 U14985 ( .A1(n15115), .A2(n15116), .ZN(n15142) );
  NOR2_X1 U14986 ( .A1(n10069), .A2(n9983), .ZN(n15116) );
  NAND2_X1 U14987 ( .A1(n15111), .A2(n15143), .ZN(n15115) );
  NAND2_X1 U14988 ( .A1(n15110), .A2(n15112), .ZN(n15143) );
  NAND2_X1 U14989 ( .A1(n15144), .A2(n15145), .ZN(n15112) );
  NAND2_X1 U14990 ( .A1(b_12_), .A2(a_2_), .ZN(n15145) );
  INV_X1 U14991 ( .A(n15146), .ZN(n15144) );
  XOR2_X1 U14992 ( .A(n15147), .B(n15148), .Z(n15110) );
  XOR2_X1 U14993 ( .A(n15149), .B(n15150), .Z(n15147) );
  NOR2_X1 U14994 ( .A1(n10071), .A2(n10086), .ZN(n15150) );
  NAND2_X1 U14995 ( .A1(a_2_), .A2(n15146), .ZN(n15111) );
  NAND2_X1 U14996 ( .A1(n15107), .A2(n15151), .ZN(n15146) );
  NAND2_X1 U14997 ( .A1(n15106), .A2(n15108), .ZN(n15151) );
  NAND2_X1 U14998 ( .A1(n15152), .A2(n15153), .ZN(n15108) );
  NAND2_X1 U14999 ( .A1(b_12_), .A2(a_3_), .ZN(n15153) );
  INV_X1 U15000 ( .A(n15154), .ZN(n15152) );
  XOR2_X1 U15001 ( .A(n15155), .B(n15156), .Z(n15106) );
  XOR2_X1 U15002 ( .A(n15157), .B(n15158), .Z(n15155) );
  NOR2_X1 U15003 ( .A1(n10071), .A2(n10085), .ZN(n15158) );
  NAND2_X1 U15004 ( .A1(a_3_), .A2(n15154), .ZN(n15107) );
  NAND2_X1 U15005 ( .A1(n15103), .A2(n15159), .ZN(n15154) );
  NAND2_X1 U15006 ( .A1(n15102), .A2(n15104), .ZN(n15159) );
  NAND2_X1 U15007 ( .A1(n15160), .A2(n15161), .ZN(n15104) );
  NAND2_X1 U15008 ( .A1(b_12_), .A2(a_4_), .ZN(n15161) );
  INV_X1 U15009 ( .A(n15162), .ZN(n15160) );
  XOR2_X1 U15010 ( .A(n15163), .B(n15164), .Z(n15102) );
  XOR2_X1 U15011 ( .A(n15165), .B(n15166), .Z(n15163) );
  NOR2_X1 U15012 ( .A1(n10071), .A2(n10083), .ZN(n15166) );
  NAND2_X1 U15013 ( .A1(a_4_), .A2(n15162), .ZN(n15103) );
  NAND2_X1 U15014 ( .A1(n15099), .A2(n15167), .ZN(n15162) );
  NAND2_X1 U15015 ( .A1(n15098), .A2(n15100), .ZN(n15167) );
  NAND2_X1 U15016 ( .A1(n15168), .A2(n15169), .ZN(n15100) );
  NAND2_X1 U15017 ( .A1(b_12_), .A2(a_5_), .ZN(n15169) );
  INV_X1 U15018 ( .A(n15170), .ZN(n15168) );
  XOR2_X1 U15019 ( .A(n15171), .B(n15172), .Z(n15098) );
  XOR2_X1 U15020 ( .A(n15173), .B(n15174), .Z(n15171) );
  NOR2_X1 U15021 ( .A1(n10071), .A2(n10081), .ZN(n15174) );
  NAND2_X1 U15022 ( .A1(a_5_), .A2(n15170), .ZN(n15099) );
  NAND2_X1 U15023 ( .A1(n15095), .A2(n15175), .ZN(n15170) );
  NAND2_X1 U15024 ( .A1(n15094), .A2(n15096), .ZN(n15175) );
  NAND2_X1 U15025 ( .A1(n15176), .A2(n15177), .ZN(n15096) );
  NAND2_X1 U15026 ( .A1(b_12_), .A2(a_6_), .ZN(n15177) );
  INV_X1 U15027 ( .A(n15178), .ZN(n15176) );
  XOR2_X1 U15028 ( .A(n15179), .B(n15180), .Z(n15094) );
  XOR2_X1 U15029 ( .A(n15181), .B(n15182), .Z(n15179) );
  NOR2_X1 U15030 ( .A1(n10071), .A2(n9773), .ZN(n15182) );
  NAND2_X1 U15031 ( .A1(a_6_), .A2(n15178), .ZN(n15095) );
  NAND2_X1 U15032 ( .A1(n15091), .A2(n15183), .ZN(n15178) );
  NAND2_X1 U15033 ( .A1(n15090), .A2(n15092), .ZN(n15183) );
  NAND2_X1 U15034 ( .A1(n15184), .A2(n15185), .ZN(n15092) );
  NAND2_X1 U15035 ( .A1(b_12_), .A2(a_7_), .ZN(n15185) );
  INV_X1 U15036 ( .A(n15186), .ZN(n15184) );
  XOR2_X1 U15037 ( .A(n15187), .B(n15188), .Z(n15090) );
  XOR2_X1 U15038 ( .A(n15189), .B(n15190), .Z(n15187) );
  NOR2_X1 U15039 ( .A1(n10071), .A2(n10079), .ZN(n15190) );
  NAND2_X1 U15040 ( .A1(a_7_), .A2(n15186), .ZN(n15091) );
  NAND2_X1 U15041 ( .A1(n14908), .A2(n15191), .ZN(n15186) );
  NAND2_X1 U15042 ( .A1(n14907), .A2(n14909), .ZN(n15191) );
  NAND2_X1 U15043 ( .A1(n15192), .A2(n15193), .ZN(n14909) );
  NAND2_X1 U15044 ( .A1(b_12_), .A2(a_8_), .ZN(n15193) );
  INV_X1 U15045 ( .A(n15194), .ZN(n15192) );
  XOR2_X1 U15046 ( .A(n15195), .B(n15196), .Z(n14907) );
  XNOR2_X1 U15047 ( .A(n15197), .B(n15198), .ZN(n15195) );
  NAND2_X1 U15048 ( .A1(a_9_), .A2(b_11_), .ZN(n15197) );
  NAND2_X1 U15049 ( .A1(a_8_), .A2(n15194), .ZN(n14908) );
  NAND2_X1 U15050 ( .A1(n14916), .A2(n15199), .ZN(n15194) );
  NAND2_X1 U15051 ( .A1(n14915), .A2(n14917), .ZN(n15199) );
  NAND2_X1 U15052 ( .A1(n15200), .A2(n15201), .ZN(n14917) );
  NAND2_X1 U15053 ( .A1(b_12_), .A2(a_9_), .ZN(n15201) );
  INV_X1 U15054 ( .A(n15202), .ZN(n15200) );
  XOR2_X1 U15055 ( .A(n15203), .B(n15204), .Z(n14915) );
  XNOR2_X1 U15056 ( .A(n15205), .B(n15206), .ZN(n15204) );
  NAND2_X1 U15057 ( .A1(a_10_), .A2(b_11_), .ZN(n15206) );
  NAND2_X1 U15058 ( .A1(a_9_), .A2(n15202), .ZN(n14916) );
  NAND2_X1 U15059 ( .A1(n15087), .A2(n15207), .ZN(n15202) );
  NAND2_X1 U15060 ( .A1(n15086), .A2(n15088), .ZN(n15207) );
  NAND2_X1 U15061 ( .A1(n15208), .A2(n15209), .ZN(n15088) );
  NAND2_X1 U15062 ( .A1(b_12_), .A2(a_10_), .ZN(n15208) );
  XNOR2_X1 U15063 ( .A(n15210), .B(n15211), .ZN(n15086) );
  XNOR2_X1 U15064 ( .A(n15212), .B(n9997), .ZN(n15210) );
  INV_X1 U15065 ( .A(n15213), .ZN(n9997) );
  INV_X1 U15066 ( .A(n15214), .ZN(n15087) );
  NOR2_X1 U15067 ( .A1(n15209), .A2(n10073), .ZN(n15214) );
  NAND2_X1 U15068 ( .A1(n15215), .A2(n15216), .ZN(n15209) );
  INV_X1 U15069 ( .A(n15217), .ZN(n15216) );
  NOR2_X1 U15070 ( .A1(n15081), .A2(n15218), .ZN(n15217) );
  NOR2_X1 U15071 ( .A1(n15084), .A2(n15083), .ZN(n15218) );
  XOR2_X1 U15072 ( .A(n15219), .B(n15220), .Z(n15081) );
  XOR2_X1 U15073 ( .A(n15221), .B(n15222), .Z(n15219) );
  NOR2_X1 U15074 ( .A1(n10070), .A2(n10071), .ZN(n15222) );
  NAND2_X1 U15075 ( .A1(n15084), .A2(n15083), .ZN(n15215) );
  NAND2_X1 U15076 ( .A1(n15223), .A2(n15224), .ZN(n15083) );
  NAND2_X1 U15077 ( .A1(n15078), .A2(n15225), .ZN(n15224) );
  INV_X1 U15078 ( .A(n15226), .ZN(n15225) );
  NOR2_X1 U15079 ( .A1(n9627), .A2(n15080), .ZN(n15226) );
  XOR2_X1 U15080 ( .A(n15227), .B(n15228), .Z(n15078) );
  XOR2_X1 U15081 ( .A(n15229), .B(n15230), .Z(n15228) );
  NAND2_X1 U15082 ( .A1(b_11_), .A2(a_13_), .ZN(n15230) );
  NAND2_X1 U15083 ( .A1(n9627), .A2(n15080), .ZN(n15223) );
  NAND2_X1 U15084 ( .A1(n15231), .A2(n15232), .ZN(n15080) );
  NAND2_X1 U15085 ( .A1(n14934), .A2(n15233), .ZN(n15232) );
  NAND2_X1 U15086 ( .A1(n14937), .A2(n14936), .ZN(n15233) );
  XOR2_X1 U15087 ( .A(n15234), .B(n15235), .Z(n14934) );
  XOR2_X1 U15088 ( .A(n15236), .B(n15237), .Z(n15235) );
  NAND2_X1 U15089 ( .A1(b_11_), .A2(a_14_), .ZN(n15237) );
  INV_X1 U15090 ( .A(n15238), .ZN(n15231) );
  NOR2_X1 U15091 ( .A1(n14936), .A2(n14937), .ZN(n15238) );
  NOR2_X1 U15092 ( .A1(n10069), .A2(n10067), .ZN(n14937) );
  NAND2_X1 U15093 ( .A1(n14944), .A2(n15239), .ZN(n14936) );
  NAND2_X1 U15094 ( .A1(n14943), .A2(n14945), .ZN(n15239) );
  NAND2_X1 U15095 ( .A1(n15240), .A2(n15241), .ZN(n14945) );
  NAND2_X1 U15096 ( .A1(b_12_), .A2(a_14_), .ZN(n15241) );
  INV_X1 U15097 ( .A(n15242), .ZN(n15240) );
  XNOR2_X1 U15098 ( .A(n15243), .B(n15244), .ZN(n14943) );
  XOR2_X1 U15099 ( .A(n15245), .B(n15246), .Z(n15244) );
  NAND2_X1 U15100 ( .A1(b_11_), .A2(a_15_), .ZN(n15246) );
  NAND2_X1 U15101 ( .A1(a_14_), .A2(n15242), .ZN(n14944) );
  NAND2_X1 U15102 ( .A1(n15247), .A2(n15248), .ZN(n15242) );
  NAND2_X1 U15103 ( .A1(n15249), .A2(b_12_), .ZN(n15248) );
  NOR2_X1 U15104 ( .A1(n15250), .A2(n9534), .ZN(n15249) );
  NOR2_X1 U15105 ( .A1(n15076), .A2(n15075), .ZN(n15250) );
  NAND2_X1 U15106 ( .A1(n15075), .A2(n15076), .ZN(n15247) );
  NAND2_X1 U15107 ( .A1(n14956), .A2(n15251), .ZN(n15076) );
  NAND2_X1 U15108 ( .A1(n14955), .A2(n14957), .ZN(n15251) );
  NAND2_X1 U15109 ( .A1(n15252), .A2(n15253), .ZN(n14957) );
  NAND2_X1 U15110 ( .A1(b_12_), .A2(a_16_), .ZN(n15253) );
  INV_X1 U15111 ( .A(n15254), .ZN(n15252) );
  XOR2_X1 U15112 ( .A(n15255), .B(n15256), .Z(n14955) );
  XNOR2_X1 U15113 ( .A(n15257), .B(n15258), .ZN(n15256) );
  NAND2_X1 U15114 ( .A1(a_16_), .A2(n15254), .ZN(n14956) );
  NAND2_X1 U15115 ( .A1(n15259), .A2(n15260), .ZN(n15254) );
  NAND2_X1 U15116 ( .A1(n15261), .A2(b_12_), .ZN(n15260) );
  NOR2_X1 U15117 ( .A1(n15262), .A2(n10060), .ZN(n15261) );
  NOR2_X1 U15118 ( .A1(n14964), .A2(n14962), .ZN(n15262) );
  NAND2_X1 U15119 ( .A1(n14962), .A2(n14964), .ZN(n15259) );
  NAND2_X1 U15120 ( .A1(n15263), .A2(n15264), .ZN(n14964) );
  NAND2_X1 U15121 ( .A1(n15265), .A2(b_12_), .ZN(n15264) );
  NOR2_X1 U15122 ( .A1(n15266), .A2(n10058), .ZN(n15265) );
  NOR2_X1 U15123 ( .A1(n14970), .A2(n14972), .ZN(n15266) );
  NAND2_X1 U15124 ( .A1(n14970), .A2(n14972), .ZN(n15263) );
  NAND2_X1 U15125 ( .A1(n15267), .A2(n15268), .ZN(n14972) );
  NAND2_X1 U15126 ( .A1(n15269), .A2(b_12_), .ZN(n15268) );
  NOR2_X1 U15127 ( .A1(n15270), .A2(n9415), .ZN(n15269) );
  NOR2_X1 U15128 ( .A1(n15070), .A2(n15072), .ZN(n15270) );
  NAND2_X1 U15129 ( .A1(n15070), .A2(n15072), .ZN(n15267) );
  NAND2_X1 U15130 ( .A1(n15271), .A2(n15272), .ZN(n15072) );
  NAND2_X1 U15131 ( .A1(n15273), .A2(b_12_), .ZN(n15272) );
  NOR2_X1 U15132 ( .A1(n15274), .A2(n10054), .ZN(n15273) );
  NOR2_X1 U15133 ( .A1(n15067), .A2(n15068), .ZN(n15274) );
  NAND2_X1 U15134 ( .A1(n15067), .A2(n15068), .ZN(n15271) );
  NAND2_X1 U15135 ( .A1(n15064), .A2(n15275), .ZN(n15068) );
  NAND2_X1 U15136 ( .A1(n15063), .A2(n15065), .ZN(n15275) );
  NAND2_X1 U15137 ( .A1(n15276), .A2(n15277), .ZN(n15065) );
  NAND2_X1 U15138 ( .A1(b_12_), .A2(a_21_), .ZN(n15277) );
  INV_X1 U15139 ( .A(n15278), .ZN(n15276) );
  XOR2_X1 U15140 ( .A(n15279), .B(n15280), .Z(n15063) );
  XOR2_X1 U15141 ( .A(n15281), .B(n15282), .Z(n15279) );
  NAND2_X1 U15142 ( .A1(a_21_), .A2(n15278), .ZN(n15064) );
  NAND2_X1 U15143 ( .A1(n15283), .A2(n15284), .ZN(n15278) );
  NAND2_X1 U15144 ( .A1(n14993), .A2(n15285), .ZN(n15284) );
  INV_X1 U15145 ( .A(n15286), .ZN(n15285) );
  NOR2_X1 U15146 ( .A1(n14992), .A2(n14991), .ZN(n15286) );
  NOR2_X1 U15147 ( .A1(n10069), .A2(n9330), .ZN(n14993) );
  NAND2_X1 U15148 ( .A1(n14991), .A2(n14992), .ZN(n15283) );
  NAND2_X1 U15149 ( .A1(n15287), .A2(n15288), .ZN(n14992) );
  NAND2_X1 U15150 ( .A1(n15061), .A2(n15289), .ZN(n15288) );
  INV_X1 U15151 ( .A(n15290), .ZN(n15289) );
  NOR2_X1 U15152 ( .A1(n15059), .A2(n15060), .ZN(n15290) );
  NOR2_X1 U15153 ( .A1(n10069), .A2(n10051), .ZN(n15061) );
  NAND2_X1 U15154 ( .A1(n15059), .A2(n15060), .ZN(n15287) );
  NAND2_X1 U15155 ( .A1(n15291), .A2(n15292), .ZN(n15060) );
  INV_X1 U15156 ( .A(n15293), .ZN(n15292) );
  NOR2_X1 U15157 ( .A1(n15057), .A2(n15294), .ZN(n15293) );
  NOR2_X1 U15158 ( .A1(n15056), .A2(n15054), .ZN(n15294) );
  NAND2_X1 U15159 ( .A1(b_12_), .A2(a_24_), .ZN(n15057) );
  NAND2_X1 U15160 ( .A1(n15054), .A2(n15056), .ZN(n15291) );
  NAND2_X1 U15161 ( .A1(n15295), .A2(n15296), .ZN(n15056) );
  NAND2_X1 U15162 ( .A1(n15053), .A2(n15297), .ZN(n15296) );
  INV_X1 U15163 ( .A(n15298), .ZN(n15297) );
  NOR2_X1 U15164 ( .A1(n15050), .A2(n15052), .ZN(n15298) );
  NOR2_X1 U15165 ( .A1(n10069), .A2(n10048), .ZN(n15053) );
  NAND2_X1 U15166 ( .A1(n15050), .A2(n15052), .ZN(n15295) );
  NOR2_X1 U15167 ( .A1(n15299), .A2(n15300), .ZN(n15052) );
  INV_X1 U15168 ( .A(n15301), .ZN(n15300) );
  NAND2_X1 U15169 ( .A1(n15010), .A2(n15302), .ZN(n15301) );
  NAND2_X1 U15170 ( .A1(n15013), .A2(n15012), .ZN(n15302) );
  XOR2_X1 U15171 ( .A(n15303), .B(n15304), .Z(n15010) );
  NAND2_X1 U15172 ( .A1(n15305), .A2(n15306), .ZN(n15303) );
  NOR2_X1 U15173 ( .A1(n15012), .A2(n15013), .ZN(n15299) );
  NOR2_X1 U15174 ( .A1(n10069), .A2(n10047), .ZN(n15013) );
  NAND2_X1 U15175 ( .A1(n15020), .A2(n15307), .ZN(n15012) );
  NAND2_X1 U15176 ( .A1(n15019), .A2(n15021), .ZN(n15307) );
  NAND2_X1 U15177 ( .A1(n15308), .A2(n15309), .ZN(n15021) );
  NAND2_X1 U15178 ( .A1(b_12_), .A2(a_27_), .ZN(n15309) );
  INV_X1 U15179 ( .A(n15310), .ZN(n15308) );
  XNOR2_X1 U15180 ( .A(n15311), .B(n15312), .ZN(n15019) );
  XOR2_X1 U15181 ( .A(n15313), .B(n15314), .Z(n15312) );
  NAND2_X1 U15182 ( .A1(b_11_), .A2(a_28_), .ZN(n15314) );
  NAND2_X1 U15183 ( .A1(a_27_), .A2(n15310), .ZN(n15020) );
  NAND2_X1 U15184 ( .A1(n15315), .A2(n15316), .ZN(n15310) );
  NAND2_X1 U15185 ( .A1(n15317), .A2(b_12_), .ZN(n15316) );
  NOR2_X1 U15186 ( .A1(n15318), .A2(n9136), .ZN(n15317) );
  NOR2_X1 U15187 ( .A1(n15026), .A2(n15028), .ZN(n15318) );
  NAND2_X1 U15188 ( .A1(n15026), .A2(n15028), .ZN(n15315) );
  NAND2_X1 U15189 ( .A1(n15319), .A2(n15320), .ZN(n15028) );
  NAND2_X1 U15190 ( .A1(n15321), .A2(b_12_), .ZN(n15320) );
  NOR2_X1 U15191 ( .A1(n15322), .A2(n9121), .ZN(n15321) );
  NOR2_X1 U15192 ( .A1(n15323), .A2(n15048), .ZN(n15322) );
  NAND2_X1 U15193 ( .A1(n15323), .A2(n15048), .ZN(n15319) );
  NAND2_X1 U15194 ( .A1(n15324), .A2(n15325), .ZN(n15048) );
  NAND2_X1 U15195 ( .A1(b_10_), .A2(n15326), .ZN(n15325) );
  NAND2_X1 U15196 ( .A1(n10486), .A2(n15327), .ZN(n15326) );
  NAND2_X1 U15197 ( .A1(a_31_), .A2(n10071), .ZN(n15327) );
  NAND2_X1 U15198 ( .A1(b_11_), .A2(n15328), .ZN(n15324) );
  NAND2_X1 U15199 ( .A1(n10489), .A2(n15329), .ZN(n15328) );
  NAND2_X1 U15200 ( .A1(a_30_), .A2(n10072), .ZN(n15329) );
  INV_X1 U15201 ( .A(n15049), .ZN(n15323) );
  NAND2_X1 U15202 ( .A1(n15330), .A2(n9025), .ZN(n15049) );
  NOR2_X1 U15203 ( .A1(n10071), .A2(n10069), .ZN(n15330) );
  XOR2_X1 U15204 ( .A(n15331), .B(n15332), .Z(n15026) );
  NOR2_X1 U15205 ( .A1(n9121), .A2(n10071), .ZN(n15332) );
  XNOR2_X1 U15206 ( .A(n15333), .B(n15334), .ZN(n15331) );
  XOR2_X1 U15207 ( .A(n15335), .B(n15336), .Z(n15050) );
  XNOR2_X1 U15208 ( .A(n15337), .B(n15338), .ZN(n15336) );
  XOR2_X1 U15209 ( .A(n15339), .B(n15340), .Z(n15054) );
  XOR2_X1 U15210 ( .A(n15341), .B(n15342), .Z(n15340) );
  XNOR2_X1 U15211 ( .A(n15343), .B(n15344), .ZN(n15059) );
  XOR2_X1 U15212 ( .A(n15345), .B(n15346), .Z(n15344) );
  XOR2_X1 U15213 ( .A(n15347), .B(n15348), .Z(n14991) );
  XOR2_X1 U15214 ( .A(n15349), .B(n15350), .Z(n15347) );
  XNOR2_X1 U15215 ( .A(n15351), .B(n15352), .ZN(n15067) );
  XNOR2_X1 U15216 ( .A(n15353), .B(n15354), .ZN(n15352) );
  XNOR2_X1 U15217 ( .A(n15355), .B(n15356), .ZN(n15070) );
  XOR2_X1 U15218 ( .A(n15357), .B(n15358), .Z(n15356) );
  XNOR2_X1 U15219 ( .A(n15359), .B(n15360), .ZN(n14970) );
  XNOR2_X1 U15220 ( .A(n15361), .B(n15362), .ZN(n15359) );
  XOR2_X1 U15221 ( .A(n15363), .B(n15364), .Z(n14962) );
  XOR2_X1 U15222 ( .A(n15365), .B(n15366), .Z(n15363) );
  NOR2_X1 U15223 ( .A1(n10058), .A2(n10071), .ZN(n15366) );
  XNOR2_X1 U15224 ( .A(n15367), .B(n15368), .ZN(n15075) );
  XNOR2_X1 U15225 ( .A(n15369), .B(n15370), .ZN(n15367) );
  NOR2_X1 U15226 ( .A1(n10062), .A2(n10071), .ZN(n15370) );
  NAND2_X1 U15227 ( .A1(b_12_), .A2(a_12_), .ZN(n9627) );
  NAND2_X1 U15228 ( .A1(b_12_), .A2(a_11_), .ZN(n15084) );
  XNOR2_X1 U15229 ( .A(n15371), .B(n15372), .ZN(n15122) );
  XOR2_X1 U15230 ( .A(n15373), .B(n15374), .Z(n15372) );
  NAND2_X1 U15231 ( .A1(a_0_), .A2(b_11_), .ZN(n15374) );
  INV_X1 U15232 ( .A(n15375), .ZN(n10263) );
  NAND2_X1 U15233 ( .A1(n15125), .A2(n15124), .ZN(n15375) );
  NAND2_X1 U15234 ( .A1(n15376), .A2(n15377), .ZN(n15124) );
  NAND2_X1 U15235 ( .A1(n15378), .A2(a_0_), .ZN(n15377) );
  NOR2_X1 U15236 ( .A1(n15379), .A2(n10071), .ZN(n15378) );
  NOR2_X1 U15237 ( .A1(n15371), .A2(n15373), .ZN(n15379) );
  NAND2_X1 U15238 ( .A1(n15371), .A2(n15373), .ZN(n15376) );
  NAND2_X1 U15239 ( .A1(n15380), .A2(n15381), .ZN(n15373) );
  NAND2_X1 U15240 ( .A1(n15382), .A2(a_1_), .ZN(n15381) );
  NOR2_X1 U15241 ( .A1(n15383), .A2(n10071), .ZN(n15382) );
  NOR2_X1 U15242 ( .A1(n15132), .A2(n15133), .ZN(n15383) );
  NAND2_X1 U15243 ( .A1(n15132), .A2(n15133), .ZN(n15380) );
  NAND2_X1 U15244 ( .A1(n15384), .A2(n15385), .ZN(n15133) );
  NAND2_X1 U15245 ( .A1(n15386), .A2(a_2_), .ZN(n15385) );
  NOR2_X1 U15246 ( .A1(n15387), .A2(n10071), .ZN(n15386) );
  NOR2_X1 U15247 ( .A1(n15139), .A2(n15140), .ZN(n15387) );
  NAND2_X1 U15248 ( .A1(n15139), .A2(n15140), .ZN(n15384) );
  NAND2_X1 U15249 ( .A1(n15388), .A2(n15389), .ZN(n15140) );
  NAND2_X1 U15250 ( .A1(n15390), .A2(a_3_), .ZN(n15389) );
  NOR2_X1 U15251 ( .A1(n15391), .A2(n10071), .ZN(n15390) );
  NOR2_X1 U15252 ( .A1(n15148), .A2(n15149), .ZN(n15391) );
  NAND2_X1 U15253 ( .A1(n15148), .A2(n15149), .ZN(n15388) );
  NAND2_X1 U15254 ( .A1(n15392), .A2(n15393), .ZN(n15149) );
  NAND2_X1 U15255 ( .A1(n15394), .A2(a_4_), .ZN(n15393) );
  NOR2_X1 U15256 ( .A1(n15395), .A2(n10071), .ZN(n15394) );
  NOR2_X1 U15257 ( .A1(n15156), .A2(n15157), .ZN(n15395) );
  NAND2_X1 U15258 ( .A1(n15156), .A2(n15157), .ZN(n15392) );
  NAND2_X1 U15259 ( .A1(n15396), .A2(n15397), .ZN(n15157) );
  NAND2_X1 U15260 ( .A1(n15398), .A2(a_5_), .ZN(n15397) );
  NOR2_X1 U15261 ( .A1(n15399), .A2(n10071), .ZN(n15398) );
  NOR2_X1 U15262 ( .A1(n15164), .A2(n15165), .ZN(n15399) );
  NAND2_X1 U15263 ( .A1(n15164), .A2(n15165), .ZN(n15396) );
  NAND2_X1 U15264 ( .A1(n15400), .A2(n15401), .ZN(n15165) );
  NAND2_X1 U15265 ( .A1(n15402), .A2(a_6_), .ZN(n15401) );
  NOR2_X1 U15266 ( .A1(n15403), .A2(n10071), .ZN(n15402) );
  NOR2_X1 U15267 ( .A1(n15172), .A2(n15173), .ZN(n15403) );
  NAND2_X1 U15268 ( .A1(n15172), .A2(n15173), .ZN(n15400) );
  NAND2_X1 U15269 ( .A1(n15404), .A2(n15405), .ZN(n15173) );
  NAND2_X1 U15270 ( .A1(n15406), .A2(a_7_), .ZN(n15405) );
  NOR2_X1 U15271 ( .A1(n15407), .A2(n10071), .ZN(n15406) );
  NOR2_X1 U15272 ( .A1(n15180), .A2(n15181), .ZN(n15407) );
  NAND2_X1 U15273 ( .A1(n15180), .A2(n15181), .ZN(n15404) );
  NAND2_X1 U15274 ( .A1(n15408), .A2(n15409), .ZN(n15181) );
  NAND2_X1 U15275 ( .A1(n15410), .A2(a_8_), .ZN(n15409) );
  NOR2_X1 U15276 ( .A1(n15411), .A2(n10071), .ZN(n15410) );
  NOR2_X1 U15277 ( .A1(n15188), .A2(n15189), .ZN(n15411) );
  NAND2_X1 U15278 ( .A1(n15188), .A2(n15189), .ZN(n15408) );
  NAND2_X1 U15279 ( .A1(n15412), .A2(n15413), .ZN(n15189) );
  NAND2_X1 U15280 ( .A1(n15414), .A2(a_9_), .ZN(n15413) );
  NOR2_X1 U15281 ( .A1(n15415), .A2(n10071), .ZN(n15414) );
  NOR2_X1 U15282 ( .A1(n15196), .A2(n15198), .ZN(n15415) );
  NAND2_X1 U15283 ( .A1(n15196), .A2(n15198), .ZN(n15412) );
  NAND2_X1 U15284 ( .A1(n15416), .A2(n15417), .ZN(n15198) );
  NAND2_X1 U15285 ( .A1(n15418), .A2(a_10_), .ZN(n15417) );
  NOR2_X1 U15286 ( .A1(n15419), .A2(n10071), .ZN(n15418) );
  NOR2_X1 U15287 ( .A1(n15205), .A2(n15203), .ZN(n15419) );
  NAND2_X1 U15288 ( .A1(n15205), .A2(n15203), .ZN(n15416) );
  XNOR2_X1 U15289 ( .A(n15420), .B(n15421), .ZN(n15203) );
  NAND2_X1 U15290 ( .A1(n15422), .A2(n15423), .ZN(n15420) );
  NOR2_X1 U15291 ( .A1(n15424), .A2(n15425), .ZN(n15205) );
  INV_X1 U15292 ( .A(n15426), .ZN(n15425) );
  NAND2_X1 U15293 ( .A1(n15211), .A2(n15427), .ZN(n15426) );
  NAND2_X1 U15294 ( .A1(n15213), .A2(n15212), .ZN(n15427) );
  XOR2_X1 U15295 ( .A(n15428), .B(n15429), .Z(n15211) );
  NAND2_X1 U15296 ( .A1(n15430), .A2(n15431), .ZN(n15428) );
  NOR2_X1 U15297 ( .A1(n15212), .A2(n15213), .ZN(n15424) );
  NOR2_X1 U15298 ( .A1(n10071), .A2(n9649), .ZN(n15213) );
  NAND2_X1 U15299 ( .A1(n15432), .A2(n15433), .ZN(n15212) );
  NAND2_X1 U15300 ( .A1(n15434), .A2(b_11_), .ZN(n15433) );
  NOR2_X1 U15301 ( .A1(n15435), .A2(n10070), .ZN(n15434) );
  NOR2_X1 U15302 ( .A1(n15220), .A2(n15221), .ZN(n15435) );
  NAND2_X1 U15303 ( .A1(n15220), .A2(n15221), .ZN(n15432) );
  NAND2_X1 U15304 ( .A1(n15436), .A2(n15437), .ZN(n15221) );
  NAND2_X1 U15305 ( .A1(n15438), .A2(b_11_), .ZN(n15437) );
  NOR2_X1 U15306 ( .A1(n15439), .A2(n10067), .ZN(n15438) );
  NOR2_X1 U15307 ( .A1(n15227), .A2(n15229), .ZN(n15439) );
  NAND2_X1 U15308 ( .A1(n15227), .A2(n15229), .ZN(n15436) );
  NAND2_X1 U15309 ( .A1(n15440), .A2(n15441), .ZN(n15229) );
  NAND2_X1 U15310 ( .A1(n15442), .A2(b_11_), .ZN(n15441) );
  NOR2_X1 U15311 ( .A1(n15443), .A2(n10065), .ZN(n15442) );
  NOR2_X1 U15312 ( .A1(n15234), .A2(n15236), .ZN(n15443) );
  NAND2_X1 U15313 ( .A1(n15234), .A2(n15236), .ZN(n15440) );
  NAND2_X1 U15314 ( .A1(n15444), .A2(n15445), .ZN(n15236) );
  NAND2_X1 U15315 ( .A1(n15446), .A2(b_11_), .ZN(n15445) );
  NOR2_X1 U15316 ( .A1(n15447), .A2(n9534), .ZN(n15446) );
  NOR2_X1 U15317 ( .A1(n15243), .A2(n15245), .ZN(n15447) );
  NAND2_X1 U15318 ( .A1(n15243), .A2(n15245), .ZN(n15444) );
  NAND2_X1 U15319 ( .A1(n15448), .A2(n15449), .ZN(n15245) );
  NAND2_X1 U15320 ( .A1(n15450), .A2(b_11_), .ZN(n15449) );
  NOR2_X1 U15321 ( .A1(n15451), .A2(n10062), .ZN(n15450) );
  NOR2_X1 U15322 ( .A1(n15369), .A2(n15368), .ZN(n15451) );
  NAND2_X1 U15323 ( .A1(n15369), .A2(n15368), .ZN(n15448) );
  XNOR2_X1 U15324 ( .A(n15452), .B(n15453), .ZN(n15368) );
  NAND2_X1 U15325 ( .A1(n15454), .A2(n15455), .ZN(n15452) );
  NOR2_X1 U15326 ( .A1(n15456), .A2(n15457), .ZN(n15369) );
  INV_X1 U15327 ( .A(n15458), .ZN(n15457) );
  NAND2_X1 U15328 ( .A1(n15255), .A2(n15459), .ZN(n15458) );
  NAND2_X1 U15329 ( .A1(n15258), .A2(n15257), .ZN(n15459) );
  XOR2_X1 U15330 ( .A(n15460), .B(n15461), .Z(n15255) );
  XNOR2_X1 U15331 ( .A(n15462), .B(n15463), .ZN(n15460) );
  NOR2_X1 U15332 ( .A1(n10058), .A2(n10072), .ZN(n15463) );
  NOR2_X1 U15333 ( .A1(n15257), .A2(n15258), .ZN(n15456) );
  NOR2_X1 U15334 ( .A1(n10071), .A2(n10060), .ZN(n15258) );
  NAND2_X1 U15335 ( .A1(n15464), .A2(n15465), .ZN(n15257) );
  NAND2_X1 U15336 ( .A1(n15466), .A2(b_11_), .ZN(n15465) );
  NOR2_X1 U15337 ( .A1(n15467), .A2(n10058), .ZN(n15466) );
  NOR2_X1 U15338 ( .A1(n15364), .A2(n15365), .ZN(n15467) );
  NAND2_X1 U15339 ( .A1(n15364), .A2(n15365), .ZN(n15464) );
  NAND2_X1 U15340 ( .A1(n15468), .A2(n15469), .ZN(n15365) );
  NAND2_X1 U15341 ( .A1(n15361), .A2(n15470), .ZN(n15469) );
  NAND2_X1 U15342 ( .A1(n15362), .A2(n15360), .ZN(n15470) );
  NOR2_X1 U15343 ( .A1(n10071), .A2(n9415), .ZN(n15361) );
  INV_X1 U15344 ( .A(n15471), .ZN(n15468) );
  NOR2_X1 U15345 ( .A1(n15360), .A2(n15362), .ZN(n15471) );
  NOR2_X1 U15346 ( .A1(n15472), .A2(n15473), .ZN(n15362) );
  NOR2_X1 U15347 ( .A1(n15358), .A2(n15474), .ZN(n15473) );
  NOR2_X1 U15348 ( .A1(n15357), .A2(n15355), .ZN(n15474) );
  NAND2_X1 U15349 ( .A1(b_11_), .A2(a_20_), .ZN(n15358) );
  INV_X1 U15350 ( .A(n15475), .ZN(n15472) );
  NAND2_X1 U15351 ( .A1(n15355), .A2(n15357), .ZN(n15475) );
  NAND2_X1 U15352 ( .A1(n15476), .A2(n15477), .ZN(n15357) );
  NAND2_X1 U15353 ( .A1(n15354), .A2(n15478), .ZN(n15477) );
  INV_X1 U15354 ( .A(n15479), .ZN(n15478) );
  NOR2_X1 U15355 ( .A1(n15353), .A2(n15351), .ZN(n15479) );
  NOR2_X1 U15356 ( .A1(n10071), .A2(n9358), .ZN(n15354) );
  NAND2_X1 U15357 ( .A1(n15351), .A2(n15353), .ZN(n15476) );
  NAND2_X1 U15358 ( .A1(n15480), .A2(n15481), .ZN(n15353) );
  NAND2_X1 U15359 ( .A1(n15282), .A2(n15482), .ZN(n15481) );
  INV_X1 U15360 ( .A(n15483), .ZN(n15482) );
  NOR2_X1 U15361 ( .A1(n15281), .A2(n15280), .ZN(n15483) );
  NOR2_X1 U15362 ( .A1(n10071), .A2(n9330), .ZN(n15282) );
  NAND2_X1 U15363 ( .A1(n15280), .A2(n15281), .ZN(n15480) );
  NAND2_X1 U15364 ( .A1(n15484), .A2(n15485), .ZN(n15281) );
  NAND2_X1 U15365 ( .A1(n15350), .A2(n15486), .ZN(n15485) );
  INV_X1 U15366 ( .A(n15487), .ZN(n15486) );
  NOR2_X1 U15367 ( .A1(n15349), .A2(n15348), .ZN(n15487) );
  NOR2_X1 U15368 ( .A1(n10071), .A2(n10051), .ZN(n15350) );
  NAND2_X1 U15369 ( .A1(n15348), .A2(n15349), .ZN(n15484) );
  NAND2_X1 U15370 ( .A1(n15488), .A2(n15489), .ZN(n15349) );
  INV_X1 U15371 ( .A(n15490), .ZN(n15489) );
  NOR2_X1 U15372 ( .A1(n15346), .A2(n15491), .ZN(n15490) );
  NOR2_X1 U15373 ( .A1(n15345), .A2(n15343), .ZN(n15491) );
  NAND2_X1 U15374 ( .A1(b_11_), .A2(a_24_), .ZN(n15346) );
  NAND2_X1 U15375 ( .A1(n15343), .A2(n15345), .ZN(n15488) );
  NAND2_X1 U15376 ( .A1(n15492), .A2(n15493), .ZN(n15345) );
  NAND2_X1 U15377 ( .A1(n15342), .A2(n15494), .ZN(n15493) );
  INV_X1 U15378 ( .A(n15495), .ZN(n15494) );
  NOR2_X1 U15379 ( .A1(n15339), .A2(n15341), .ZN(n15495) );
  NOR2_X1 U15380 ( .A1(n10071), .A2(n10048), .ZN(n15342) );
  NAND2_X1 U15381 ( .A1(n15341), .A2(n15339), .ZN(n15492) );
  XOR2_X1 U15382 ( .A(n15496), .B(n15497), .Z(n15339) );
  XNOR2_X1 U15383 ( .A(n15498), .B(n15499), .ZN(n15497) );
  NOR2_X1 U15384 ( .A1(n15500), .A2(n15501), .ZN(n15341) );
  INV_X1 U15385 ( .A(n15502), .ZN(n15501) );
  NAND2_X1 U15386 ( .A1(n15335), .A2(n15503), .ZN(n15502) );
  NAND2_X1 U15387 ( .A1(n15338), .A2(n15337), .ZN(n15503) );
  XOR2_X1 U15388 ( .A(n15504), .B(n15505), .Z(n15335) );
  NAND2_X1 U15389 ( .A1(n15506), .A2(n15507), .ZN(n15504) );
  NOR2_X1 U15390 ( .A1(n15337), .A2(n15338), .ZN(n15500) );
  NOR2_X1 U15391 ( .A1(n10071), .A2(n10047), .ZN(n15338) );
  NAND2_X1 U15392 ( .A1(n15305), .A2(n15508), .ZN(n15337) );
  NAND2_X1 U15393 ( .A1(n15304), .A2(n15306), .ZN(n15508) );
  NAND2_X1 U15394 ( .A1(n15509), .A2(n15510), .ZN(n15306) );
  NAND2_X1 U15395 ( .A1(b_11_), .A2(a_27_), .ZN(n15510) );
  INV_X1 U15396 ( .A(n15511), .ZN(n15509) );
  XNOR2_X1 U15397 ( .A(n15512), .B(n15513), .ZN(n15304) );
  XOR2_X1 U15398 ( .A(n15514), .B(n15515), .Z(n15513) );
  NAND2_X1 U15399 ( .A1(b_10_), .A2(a_28_), .ZN(n15515) );
  NAND2_X1 U15400 ( .A1(a_27_), .A2(n15511), .ZN(n15305) );
  NAND2_X1 U15401 ( .A1(n15516), .A2(n15517), .ZN(n15511) );
  NAND2_X1 U15402 ( .A1(n15518), .A2(b_11_), .ZN(n15517) );
  NOR2_X1 U15403 ( .A1(n15519), .A2(n9136), .ZN(n15518) );
  NOR2_X1 U15404 ( .A1(n15311), .A2(n15313), .ZN(n15519) );
  NAND2_X1 U15405 ( .A1(n15311), .A2(n15313), .ZN(n15516) );
  NAND2_X1 U15406 ( .A1(n15520), .A2(n15521), .ZN(n15313) );
  NAND2_X1 U15407 ( .A1(n15522), .A2(b_11_), .ZN(n15521) );
  NOR2_X1 U15408 ( .A1(n15523), .A2(n9121), .ZN(n15522) );
  NOR2_X1 U15409 ( .A1(n15524), .A2(n15333), .ZN(n15523) );
  NAND2_X1 U15410 ( .A1(n15524), .A2(n15333), .ZN(n15520) );
  NAND2_X1 U15411 ( .A1(n15525), .A2(n15526), .ZN(n15333) );
  NAND2_X1 U15412 ( .A1(b_10_), .A2(n15527), .ZN(n15526) );
  NAND2_X1 U15413 ( .A1(n10489), .A2(n15528), .ZN(n15527) );
  NAND2_X1 U15414 ( .A1(a_30_), .A2(n10075), .ZN(n15528) );
  NAND2_X1 U15415 ( .A1(b_9_), .A2(n15529), .ZN(n15525) );
  NAND2_X1 U15416 ( .A1(n10486), .A2(n15530), .ZN(n15529) );
  NAND2_X1 U15417 ( .A1(a_31_), .A2(n10072), .ZN(n15530) );
  INV_X1 U15418 ( .A(n15334), .ZN(n15524) );
  NAND2_X1 U15419 ( .A1(n15531), .A2(n9025), .ZN(n15334) );
  NOR2_X1 U15420 ( .A1(n10071), .A2(n10072), .ZN(n15531) );
  XOR2_X1 U15421 ( .A(n15532), .B(n15533), .Z(n15311) );
  NOR2_X1 U15422 ( .A1(n9121), .A2(n10072), .ZN(n15533) );
  XNOR2_X1 U15423 ( .A(n15534), .B(n15535), .ZN(n15532) );
  XOR2_X1 U15424 ( .A(n15536), .B(n15537), .Z(n15343) );
  XOR2_X1 U15425 ( .A(n15538), .B(n15539), .Z(n15537) );
  XNOR2_X1 U15426 ( .A(n15540), .B(n15541), .ZN(n15348) );
  XOR2_X1 U15427 ( .A(n15542), .B(n15543), .Z(n15541) );
  XOR2_X1 U15428 ( .A(n15544), .B(n15545), .Z(n15280) );
  XOR2_X1 U15429 ( .A(n15546), .B(n15547), .Z(n15544) );
  XOR2_X1 U15430 ( .A(n15548), .B(n15549), .Z(n15351) );
  XOR2_X1 U15431 ( .A(n15550), .B(n15551), .Z(n15548) );
  XNOR2_X1 U15432 ( .A(n15552), .B(n15553), .ZN(n15355) );
  NAND2_X1 U15433 ( .A1(n15554), .A2(n15555), .ZN(n15552) );
  XNOR2_X1 U15434 ( .A(n15556), .B(n15557), .ZN(n15360) );
  XOR2_X1 U15435 ( .A(n15558), .B(n15559), .Z(n15556) );
  NOR2_X1 U15436 ( .A1(n10054), .A2(n10072), .ZN(n15559) );
  XOR2_X1 U15437 ( .A(n15560), .B(n15561), .Z(n15364) );
  XNOR2_X1 U15438 ( .A(n15562), .B(n15563), .ZN(n15561) );
  XNOR2_X1 U15439 ( .A(n15564), .B(n15565), .ZN(n15243) );
  NAND2_X1 U15440 ( .A1(n15566), .A2(n15567), .ZN(n15564) );
  XNOR2_X1 U15441 ( .A(n15568), .B(n15569), .ZN(n15234) );
  NAND2_X1 U15442 ( .A1(n15570), .A2(n15571), .ZN(n15568) );
  XNOR2_X1 U15443 ( .A(n15572), .B(n15573), .ZN(n15227) );
  NAND2_X1 U15444 ( .A1(n15574), .A2(n15575), .ZN(n15572) );
  XNOR2_X1 U15445 ( .A(n15576), .B(n15577), .ZN(n15220) );
  NAND2_X1 U15446 ( .A1(n15578), .A2(n15579), .ZN(n15576) );
  XOR2_X1 U15447 ( .A(n15580), .B(n15581), .Z(n15196) );
  XNOR2_X1 U15448 ( .A(n10074), .B(n15582), .ZN(n15581) );
  XNOR2_X1 U15449 ( .A(n15583), .B(n15584), .ZN(n15188) );
  NAND2_X1 U15450 ( .A1(n15585), .A2(n15586), .ZN(n15583) );
  XOR2_X1 U15451 ( .A(n15587), .B(n15588), .Z(n15180) );
  XNOR2_X1 U15452 ( .A(n15589), .B(n15590), .ZN(n15588) );
  XNOR2_X1 U15453 ( .A(n15591), .B(n15592), .ZN(n15172) );
  XNOR2_X1 U15454 ( .A(n15593), .B(n15594), .ZN(n15592) );
  XOR2_X1 U15455 ( .A(n15595), .B(n15596), .Z(n15164) );
  XOR2_X1 U15456 ( .A(n15597), .B(n15598), .Z(n15595) );
  XOR2_X1 U15457 ( .A(n15599), .B(n15600), .Z(n15156) );
  XOR2_X1 U15458 ( .A(n15601), .B(n15602), .Z(n15599) );
  XNOR2_X1 U15459 ( .A(n15603), .B(n15604), .ZN(n15148) );
  XOR2_X1 U15460 ( .A(n15605), .B(n15606), .Z(n15604) );
  XNOR2_X1 U15461 ( .A(n15607), .B(n15608), .ZN(n15139) );
  XNOR2_X1 U15462 ( .A(n15609), .B(n15610), .ZN(n15608) );
  XOR2_X1 U15463 ( .A(n15611), .B(n15612), .Z(n15132) );
  XOR2_X1 U15464 ( .A(n15613), .B(n15614), .Z(n15611) );
  XOR2_X1 U15465 ( .A(n15615), .B(n15616), .Z(n15371) );
  XOR2_X1 U15466 ( .A(n15617), .B(n15618), .Z(n15615) );
  XNOR2_X1 U15467 ( .A(n15619), .B(n15620), .ZN(n15125) );
  XNOR2_X1 U15468 ( .A(n15621), .B(n15622), .ZN(n15620) );
  XOR2_X1 U15469 ( .A(n15623), .B(n15624), .Z(n10242) );
  NAND2_X1 U15470 ( .A1(n9039), .A2(n9040), .ZN(n9038) );
  NOR2_X1 U15471 ( .A1(n15624), .A2(n15625), .ZN(n9040) );
  INV_X1 U15472 ( .A(n15623), .ZN(n15625) );
  NAND2_X1 U15473 ( .A1(n15626), .A2(n15627), .ZN(n15623) );
  NAND2_X1 U15474 ( .A1(n15622), .A2(n15628), .ZN(n15627) );
  INV_X1 U15475 ( .A(n15629), .ZN(n15628) );
  NOR2_X1 U15476 ( .A1(n15619), .A2(n15621), .ZN(n15629) );
  NOR2_X1 U15477 ( .A1(n10072), .A2(n10093), .ZN(n15622) );
  NAND2_X1 U15478 ( .A1(n15619), .A2(n15621), .ZN(n15626) );
  NAND2_X1 U15479 ( .A1(n15630), .A2(n15631), .ZN(n15621) );
  NAND2_X1 U15480 ( .A1(n15618), .A2(n15632), .ZN(n15631) );
  INV_X1 U15481 ( .A(n15633), .ZN(n15632) );
  NOR2_X1 U15482 ( .A1(n15616), .A2(n15617), .ZN(n15633) );
  NOR2_X1 U15483 ( .A1(n10072), .A2(n9983), .ZN(n15618) );
  NAND2_X1 U15484 ( .A1(n15616), .A2(n15617), .ZN(n15630) );
  NAND2_X1 U15485 ( .A1(n15634), .A2(n15635), .ZN(n15617) );
  NAND2_X1 U15486 ( .A1(n15614), .A2(n15636), .ZN(n15635) );
  INV_X1 U15487 ( .A(n15637), .ZN(n15636) );
  NOR2_X1 U15488 ( .A1(n15612), .A2(n15613), .ZN(n15637) );
  NOR2_X1 U15489 ( .A1(n10072), .A2(n10088), .ZN(n15614) );
  NAND2_X1 U15490 ( .A1(n15612), .A2(n15613), .ZN(n15634) );
  NAND2_X1 U15491 ( .A1(n15638), .A2(n15639), .ZN(n15613) );
  NAND2_X1 U15492 ( .A1(n15610), .A2(n15640), .ZN(n15639) );
  INV_X1 U15493 ( .A(n15641), .ZN(n15640) );
  NOR2_X1 U15494 ( .A1(n15607), .A2(n15609), .ZN(n15641) );
  NOR2_X1 U15495 ( .A1(n10072), .A2(n10086), .ZN(n15610) );
  NAND2_X1 U15496 ( .A1(n15607), .A2(n15609), .ZN(n15638) );
  NAND2_X1 U15497 ( .A1(n15642), .A2(n15643), .ZN(n15609) );
  INV_X1 U15498 ( .A(n15644), .ZN(n15643) );
  NOR2_X1 U15499 ( .A1(n15606), .A2(n15645), .ZN(n15644) );
  NOR2_X1 U15500 ( .A1(n15603), .A2(n15605), .ZN(n15645) );
  NAND2_X1 U15501 ( .A1(b_10_), .A2(a_4_), .ZN(n15606) );
  NAND2_X1 U15502 ( .A1(n15603), .A2(n15605), .ZN(n15642) );
  NAND2_X1 U15503 ( .A1(n15646), .A2(n15647), .ZN(n15605) );
  NAND2_X1 U15504 ( .A1(n15602), .A2(n15648), .ZN(n15647) );
  INV_X1 U15505 ( .A(n15649), .ZN(n15648) );
  NOR2_X1 U15506 ( .A1(n15600), .A2(n15601), .ZN(n15649) );
  NOR2_X1 U15507 ( .A1(n10072), .A2(n10083), .ZN(n15602) );
  NAND2_X1 U15508 ( .A1(n15600), .A2(n15601), .ZN(n15646) );
  NAND2_X1 U15509 ( .A1(n15650), .A2(n15651), .ZN(n15601) );
  NAND2_X1 U15510 ( .A1(n15598), .A2(n15652), .ZN(n15651) );
  INV_X1 U15511 ( .A(n15653), .ZN(n15652) );
  NOR2_X1 U15512 ( .A1(n15596), .A2(n15597), .ZN(n15653) );
  NOR2_X1 U15513 ( .A1(n10072), .A2(n10081), .ZN(n15598) );
  NAND2_X1 U15514 ( .A1(n15596), .A2(n15597), .ZN(n15650) );
  NAND2_X1 U15515 ( .A1(n15654), .A2(n15655), .ZN(n15597) );
  NAND2_X1 U15516 ( .A1(n15594), .A2(n15656), .ZN(n15655) );
  NAND2_X1 U15517 ( .A1(n15591), .A2(n15593), .ZN(n15656) );
  NOR2_X1 U15518 ( .A1(n10072), .A2(n9773), .ZN(n15594) );
  INV_X1 U15519 ( .A(n15657), .ZN(n15654) );
  NOR2_X1 U15520 ( .A1(n15593), .A2(n15591), .ZN(n15657) );
  XNOR2_X1 U15521 ( .A(n15658), .B(n15659), .ZN(n15591) );
  XNOR2_X1 U15522 ( .A(n15660), .B(n15661), .ZN(n15659) );
  NAND2_X1 U15523 ( .A1(b_9_), .A2(a_8_), .ZN(n15661) );
  NAND2_X1 U15524 ( .A1(n15662), .A2(n15663), .ZN(n15593) );
  NAND2_X1 U15525 ( .A1(n15587), .A2(n15664), .ZN(n15663) );
  NAND2_X1 U15526 ( .A1(n15590), .A2(n15589), .ZN(n15664) );
  XNOR2_X1 U15527 ( .A(n15665), .B(n15666), .ZN(n15587) );
  XNOR2_X1 U15528 ( .A(n15667), .B(n10077), .ZN(n15666) );
  INV_X1 U15529 ( .A(n15668), .ZN(n15662) );
  NOR2_X1 U15530 ( .A1(n15589), .A2(n15590), .ZN(n15668) );
  NOR2_X1 U15531 ( .A1(n10072), .A2(n10079), .ZN(n15590) );
  NAND2_X1 U15532 ( .A1(n15585), .A2(n15669), .ZN(n15589) );
  NAND2_X1 U15533 ( .A1(n15584), .A2(n15586), .ZN(n15669) );
  NAND2_X1 U15534 ( .A1(n15670), .A2(n15671), .ZN(n15586) );
  NAND2_X1 U15535 ( .A1(b_10_), .A2(a_9_), .ZN(n15671) );
  INV_X1 U15536 ( .A(n15672), .ZN(n15670) );
  XNOR2_X1 U15537 ( .A(n15673), .B(n15674), .ZN(n15584) );
  XOR2_X1 U15538 ( .A(n15675), .B(n15676), .Z(n15674) );
  NAND2_X1 U15539 ( .A1(b_9_), .A2(a_10_), .ZN(n15676) );
  NAND2_X1 U15540 ( .A1(a_9_), .A2(n15672), .ZN(n15585) );
  NAND2_X1 U15541 ( .A1(n15677), .A2(n15678), .ZN(n15672) );
  INV_X1 U15542 ( .A(n15679), .ZN(n15678) );
  NOR2_X1 U15543 ( .A1(n15580), .A2(n15680), .ZN(n15679) );
  NOR2_X1 U15544 ( .A1(n15582), .A2(n10074), .ZN(n15680) );
  XNOR2_X1 U15545 ( .A(n15681), .B(n15682), .ZN(n15580) );
  XOR2_X1 U15546 ( .A(n15683), .B(n15684), .Z(n15681) );
  NOR2_X1 U15547 ( .A1(n9649), .A2(n10075), .ZN(n15684) );
  NAND2_X1 U15548 ( .A1(n10074), .A2(n15582), .ZN(n15677) );
  NAND2_X1 U15549 ( .A1(n15422), .A2(n15685), .ZN(n15582) );
  NAND2_X1 U15550 ( .A1(n15421), .A2(n15423), .ZN(n15685) );
  NAND2_X1 U15551 ( .A1(n15686), .A2(n15687), .ZN(n15423) );
  NAND2_X1 U15552 ( .A1(b_10_), .A2(a_11_), .ZN(n15687) );
  INV_X1 U15553 ( .A(n15688), .ZN(n15686) );
  XNOR2_X1 U15554 ( .A(n15689), .B(n15690), .ZN(n15421) );
  XOR2_X1 U15555 ( .A(n15691), .B(n15692), .Z(n15690) );
  NAND2_X1 U15556 ( .A1(b_9_), .A2(a_12_), .ZN(n15692) );
  NAND2_X1 U15557 ( .A1(a_11_), .A2(n15688), .ZN(n15422) );
  NAND2_X1 U15558 ( .A1(n15430), .A2(n15693), .ZN(n15688) );
  NAND2_X1 U15559 ( .A1(n15429), .A2(n15431), .ZN(n15693) );
  NAND2_X1 U15560 ( .A1(n15694), .A2(n15695), .ZN(n15431) );
  NAND2_X1 U15561 ( .A1(b_10_), .A2(a_12_), .ZN(n15695) );
  INV_X1 U15562 ( .A(n15696), .ZN(n15694) );
  XOR2_X1 U15563 ( .A(n15697), .B(n15698), .Z(n15429) );
  XNOR2_X1 U15564 ( .A(n15699), .B(n15700), .ZN(n15698) );
  NAND2_X1 U15565 ( .A1(b_9_), .A2(a_13_), .ZN(n15700) );
  NAND2_X1 U15566 ( .A1(a_12_), .A2(n15696), .ZN(n15430) );
  NAND2_X1 U15567 ( .A1(n15578), .A2(n15701), .ZN(n15696) );
  NAND2_X1 U15568 ( .A1(n15577), .A2(n15579), .ZN(n15701) );
  NAND2_X1 U15569 ( .A1(n15702), .A2(n15703), .ZN(n15579) );
  NAND2_X1 U15570 ( .A1(b_10_), .A2(a_13_), .ZN(n15703) );
  INV_X1 U15571 ( .A(n15704), .ZN(n15702) );
  XNOR2_X1 U15572 ( .A(n15705), .B(n15706), .ZN(n15577) );
  XOR2_X1 U15573 ( .A(n15707), .B(n15708), .Z(n15705) );
  NAND2_X1 U15574 ( .A1(a_13_), .A2(n15704), .ZN(n15578) );
  NAND2_X1 U15575 ( .A1(n15574), .A2(n15709), .ZN(n15704) );
  NAND2_X1 U15576 ( .A1(n15573), .A2(n15575), .ZN(n15709) );
  NAND2_X1 U15577 ( .A1(n15710), .A2(n15711), .ZN(n15575) );
  NAND2_X1 U15578 ( .A1(b_10_), .A2(a_14_), .ZN(n15711) );
  INV_X1 U15579 ( .A(n15712), .ZN(n15710) );
  XNOR2_X1 U15580 ( .A(n15713), .B(n15714), .ZN(n15573) );
  XOR2_X1 U15581 ( .A(n15715), .B(n15716), .Z(n15714) );
  NAND2_X1 U15582 ( .A1(b_9_), .A2(a_15_), .ZN(n15716) );
  NAND2_X1 U15583 ( .A1(a_14_), .A2(n15712), .ZN(n15574) );
  NAND2_X1 U15584 ( .A1(n15570), .A2(n15717), .ZN(n15712) );
  NAND2_X1 U15585 ( .A1(n15569), .A2(n15571), .ZN(n15717) );
  NAND2_X1 U15586 ( .A1(n15718), .A2(n15719), .ZN(n15571) );
  NAND2_X1 U15587 ( .A1(b_10_), .A2(a_15_), .ZN(n15719) );
  INV_X1 U15588 ( .A(n15720), .ZN(n15718) );
  XNOR2_X1 U15589 ( .A(n15721), .B(n15722), .ZN(n15569) );
  XOR2_X1 U15590 ( .A(n15723), .B(n15724), .Z(n15722) );
  NAND2_X1 U15591 ( .A1(b_9_), .A2(a_16_), .ZN(n15724) );
  NAND2_X1 U15592 ( .A1(a_15_), .A2(n15720), .ZN(n15570) );
  NAND2_X1 U15593 ( .A1(n15566), .A2(n15725), .ZN(n15720) );
  NAND2_X1 U15594 ( .A1(n15565), .A2(n15567), .ZN(n15725) );
  NAND2_X1 U15595 ( .A1(n15726), .A2(n15727), .ZN(n15567) );
  NAND2_X1 U15596 ( .A1(b_10_), .A2(a_16_), .ZN(n15727) );
  INV_X1 U15597 ( .A(n15728), .ZN(n15726) );
  XOR2_X1 U15598 ( .A(n15729), .B(n15730), .Z(n15565) );
  XOR2_X1 U15599 ( .A(n15731), .B(n15732), .Z(n15729) );
  NOR2_X1 U15600 ( .A1(n10060), .A2(n10075), .ZN(n15732) );
  NAND2_X1 U15601 ( .A1(a_16_), .A2(n15728), .ZN(n15566) );
  NAND2_X1 U15602 ( .A1(n15454), .A2(n15733), .ZN(n15728) );
  NAND2_X1 U15603 ( .A1(n15453), .A2(n15455), .ZN(n15733) );
  NAND2_X1 U15604 ( .A1(n15734), .A2(n15735), .ZN(n15455) );
  NAND2_X1 U15605 ( .A1(b_10_), .A2(a_17_), .ZN(n15735) );
  INV_X1 U15606 ( .A(n15736), .ZN(n15734) );
  XOR2_X1 U15607 ( .A(n15737), .B(n15738), .Z(n15453) );
  XOR2_X1 U15608 ( .A(n15739), .B(n15740), .Z(n15737) );
  NOR2_X1 U15609 ( .A1(n10058), .A2(n10075), .ZN(n15740) );
  NAND2_X1 U15610 ( .A1(a_17_), .A2(n15736), .ZN(n15454) );
  NAND2_X1 U15611 ( .A1(n15741), .A2(n15742), .ZN(n15736) );
  NAND2_X1 U15612 ( .A1(n15743), .A2(b_10_), .ZN(n15742) );
  NOR2_X1 U15613 ( .A1(n15744), .A2(n10058), .ZN(n15743) );
  NOR2_X1 U15614 ( .A1(n15462), .A2(n15461), .ZN(n15744) );
  NAND2_X1 U15615 ( .A1(n15461), .A2(n15462), .ZN(n15741) );
  NOR2_X1 U15616 ( .A1(n15745), .A2(n15746), .ZN(n15462) );
  INV_X1 U15617 ( .A(n15747), .ZN(n15746) );
  NAND2_X1 U15618 ( .A1(n15560), .A2(n15748), .ZN(n15747) );
  NAND2_X1 U15619 ( .A1(n15563), .A2(n15562), .ZN(n15748) );
  XNOR2_X1 U15620 ( .A(n15749), .B(n15750), .ZN(n15560) );
  XOR2_X1 U15621 ( .A(n15751), .B(n15752), .Z(n15749) );
  NOR2_X1 U15622 ( .A1(n10054), .A2(n10075), .ZN(n15752) );
  NOR2_X1 U15623 ( .A1(n15562), .A2(n15563), .ZN(n15745) );
  NOR2_X1 U15624 ( .A1(n10072), .A2(n9415), .ZN(n15563) );
  NAND2_X1 U15625 ( .A1(n15753), .A2(n15754), .ZN(n15562) );
  NAND2_X1 U15626 ( .A1(n15755), .A2(b_10_), .ZN(n15754) );
  NOR2_X1 U15627 ( .A1(n15756), .A2(n10054), .ZN(n15755) );
  NOR2_X1 U15628 ( .A1(n15557), .A2(n15558), .ZN(n15756) );
  NAND2_X1 U15629 ( .A1(n15557), .A2(n15558), .ZN(n15753) );
  NAND2_X1 U15630 ( .A1(n15554), .A2(n15757), .ZN(n15558) );
  NAND2_X1 U15631 ( .A1(n15553), .A2(n15555), .ZN(n15757) );
  NAND2_X1 U15632 ( .A1(n15758), .A2(n15759), .ZN(n15555) );
  NAND2_X1 U15633 ( .A1(b_10_), .A2(a_21_), .ZN(n15759) );
  INV_X1 U15634 ( .A(n15760), .ZN(n15758) );
  XOR2_X1 U15635 ( .A(n15761), .B(n15762), .Z(n15553) );
  XOR2_X1 U15636 ( .A(n15763), .B(n15764), .Z(n15761) );
  NAND2_X1 U15637 ( .A1(a_21_), .A2(n15760), .ZN(n15554) );
  NAND2_X1 U15638 ( .A1(n15765), .A2(n15766), .ZN(n15760) );
  NAND2_X1 U15639 ( .A1(n15551), .A2(n15767), .ZN(n15766) );
  INV_X1 U15640 ( .A(n15768), .ZN(n15767) );
  NOR2_X1 U15641 ( .A1(n15550), .A2(n15549), .ZN(n15768) );
  NOR2_X1 U15642 ( .A1(n10072), .A2(n9330), .ZN(n15551) );
  NAND2_X1 U15643 ( .A1(n15549), .A2(n15550), .ZN(n15765) );
  NAND2_X1 U15644 ( .A1(n15769), .A2(n15770), .ZN(n15550) );
  NAND2_X1 U15645 ( .A1(n15547), .A2(n15771), .ZN(n15770) );
  INV_X1 U15646 ( .A(n15772), .ZN(n15771) );
  NOR2_X1 U15647 ( .A1(n15545), .A2(n15546), .ZN(n15772) );
  NOR2_X1 U15648 ( .A1(n10072), .A2(n10051), .ZN(n15547) );
  NAND2_X1 U15649 ( .A1(n15545), .A2(n15546), .ZN(n15769) );
  NAND2_X1 U15650 ( .A1(n15773), .A2(n15774), .ZN(n15546) );
  INV_X1 U15651 ( .A(n15775), .ZN(n15774) );
  NOR2_X1 U15652 ( .A1(n15543), .A2(n15776), .ZN(n15775) );
  NOR2_X1 U15653 ( .A1(n15542), .A2(n15540), .ZN(n15776) );
  NAND2_X1 U15654 ( .A1(b_10_), .A2(a_24_), .ZN(n15543) );
  NAND2_X1 U15655 ( .A1(n15540), .A2(n15542), .ZN(n15773) );
  NAND2_X1 U15656 ( .A1(n15777), .A2(n15778), .ZN(n15542) );
  NAND2_X1 U15657 ( .A1(n15539), .A2(n15779), .ZN(n15778) );
  INV_X1 U15658 ( .A(n15780), .ZN(n15779) );
  NOR2_X1 U15659 ( .A1(n15536), .A2(n15538), .ZN(n15780) );
  NOR2_X1 U15660 ( .A1(n10072), .A2(n10048), .ZN(n15539) );
  NAND2_X1 U15661 ( .A1(n15536), .A2(n15538), .ZN(n15777) );
  NOR2_X1 U15662 ( .A1(n15781), .A2(n15782), .ZN(n15538) );
  INV_X1 U15663 ( .A(n15783), .ZN(n15782) );
  NAND2_X1 U15664 ( .A1(n15496), .A2(n15784), .ZN(n15783) );
  NAND2_X1 U15665 ( .A1(n15499), .A2(n15498), .ZN(n15784) );
  XOR2_X1 U15666 ( .A(n15785), .B(n15786), .Z(n15496) );
  NAND2_X1 U15667 ( .A1(n15787), .A2(n15788), .ZN(n15785) );
  NOR2_X1 U15668 ( .A1(n15498), .A2(n15499), .ZN(n15781) );
  NOR2_X1 U15669 ( .A1(n10072), .A2(n10047), .ZN(n15499) );
  NAND2_X1 U15670 ( .A1(n15506), .A2(n15789), .ZN(n15498) );
  NAND2_X1 U15671 ( .A1(n15505), .A2(n15507), .ZN(n15789) );
  NAND2_X1 U15672 ( .A1(n15790), .A2(n15791), .ZN(n15507) );
  NAND2_X1 U15673 ( .A1(b_10_), .A2(a_27_), .ZN(n15791) );
  INV_X1 U15674 ( .A(n15792), .ZN(n15790) );
  XNOR2_X1 U15675 ( .A(n15793), .B(n15794), .ZN(n15505) );
  XOR2_X1 U15676 ( .A(n15795), .B(n15796), .Z(n15794) );
  NAND2_X1 U15677 ( .A1(b_9_), .A2(a_28_), .ZN(n15796) );
  NAND2_X1 U15678 ( .A1(a_27_), .A2(n15792), .ZN(n15506) );
  NAND2_X1 U15679 ( .A1(n15797), .A2(n15798), .ZN(n15792) );
  NAND2_X1 U15680 ( .A1(n15799), .A2(b_10_), .ZN(n15798) );
  NOR2_X1 U15681 ( .A1(n15800), .A2(n9136), .ZN(n15799) );
  NOR2_X1 U15682 ( .A1(n15512), .A2(n15514), .ZN(n15800) );
  NAND2_X1 U15683 ( .A1(n15512), .A2(n15514), .ZN(n15797) );
  NAND2_X1 U15684 ( .A1(n15801), .A2(n15802), .ZN(n15514) );
  NAND2_X1 U15685 ( .A1(n15803), .A2(b_10_), .ZN(n15802) );
  NOR2_X1 U15686 ( .A1(n15804), .A2(n9121), .ZN(n15803) );
  NOR2_X1 U15687 ( .A1(n15805), .A2(n15534), .ZN(n15804) );
  NAND2_X1 U15688 ( .A1(n15805), .A2(n15534), .ZN(n15801) );
  NAND2_X1 U15689 ( .A1(n15806), .A2(n15807), .ZN(n15534) );
  NAND2_X1 U15690 ( .A1(b_8_), .A2(n15808), .ZN(n15807) );
  NAND2_X1 U15691 ( .A1(n10486), .A2(n15809), .ZN(n15808) );
  NAND2_X1 U15692 ( .A1(a_31_), .A2(n10075), .ZN(n15809) );
  NAND2_X1 U15693 ( .A1(b_9_), .A2(n15810), .ZN(n15806) );
  NAND2_X1 U15694 ( .A1(n10489), .A2(n15811), .ZN(n15810) );
  NAND2_X1 U15695 ( .A1(a_30_), .A2(n10078), .ZN(n15811) );
  INV_X1 U15696 ( .A(n15535), .ZN(n15805) );
  NAND2_X1 U15697 ( .A1(n15812), .A2(n9025), .ZN(n15535) );
  NOR2_X1 U15698 ( .A1(n10072), .A2(n10075), .ZN(n15812) );
  XOR2_X1 U15699 ( .A(n15813), .B(n15814), .Z(n15512) );
  NOR2_X1 U15700 ( .A1(n9121), .A2(n10075), .ZN(n15814) );
  XNOR2_X1 U15701 ( .A(n15815), .B(n15816), .ZN(n15813) );
  XOR2_X1 U15702 ( .A(n15817), .B(n15818), .Z(n15536) );
  XNOR2_X1 U15703 ( .A(n15819), .B(n15820), .ZN(n15818) );
  XOR2_X1 U15704 ( .A(n15821), .B(n15822), .Z(n15540) );
  XOR2_X1 U15705 ( .A(n15823), .B(n15824), .Z(n15822) );
  XNOR2_X1 U15706 ( .A(n15825), .B(n15826), .ZN(n15545) );
  XOR2_X1 U15707 ( .A(n15827), .B(n15828), .Z(n15826) );
  XOR2_X1 U15708 ( .A(n15829), .B(n15830), .Z(n15549) );
  XOR2_X1 U15709 ( .A(n15831), .B(n15832), .Z(n15829) );
  XNOR2_X1 U15710 ( .A(n15833), .B(n15834), .ZN(n15557) );
  NAND2_X1 U15711 ( .A1(n15835), .A2(n15836), .ZN(n15833) );
  XNOR2_X1 U15712 ( .A(n15837), .B(n15838), .ZN(n15461) );
  XOR2_X1 U15713 ( .A(n15839), .B(n15840), .Z(n15838) );
  NAND2_X1 U15714 ( .A1(b_9_), .A2(a_19_), .ZN(n15840) );
  NOR2_X1 U15715 ( .A1(n10072), .A2(n10073), .ZN(n10074) );
  XNOR2_X1 U15716 ( .A(n15841), .B(n15842), .ZN(n15596) );
  XOR2_X1 U15717 ( .A(n15843), .B(n15844), .Z(n15842) );
  NAND2_X1 U15718 ( .A1(b_9_), .A2(a_7_), .ZN(n15844) );
  XNOR2_X1 U15719 ( .A(n15845), .B(n15846), .ZN(n15600) );
  XOR2_X1 U15720 ( .A(n15847), .B(n15848), .Z(n15846) );
  NAND2_X1 U15721 ( .A1(b_9_), .A2(a_6_), .ZN(n15848) );
  XOR2_X1 U15722 ( .A(n15849), .B(n15850), .Z(n15603) );
  XOR2_X1 U15723 ( .A(n15851), .B(n15852), .Z(n15849) );
  NOR2_X1 U15724 ( .A1(n10083), .A2(n10075), .ZN(n15852) );
  XOR2_X1 U15725 ( .A(n15853), .B(n15854), .Z(n15607) );
  XOR2_X1 U15726 ( .A(n15855), .B(n15856), .Z(n15853) );
  NOR2_X1 U15727 ( .A1(n10085), .A2(n10075), .ZN(n15856) );
  XNOR2_X1 U15728 ( .A(n15857), .B(n15858), .ZN(n15612) );
  XOR2_X1 U15729 ( .A(n15859), .B(n15860), .Z(n15858) );
  NAND2_X1 U15730 ( .A1(b_9_), .A2(a_3_), .ZN(n15860) );
  XOR2_X1 U15731 ( .A(n15861), .B(n15862), .Z(n15616) );
  XOR2_X1 U15732 ( .A(n15863), .B(n15864), .Z(n15861) );
  NOR2_X1 U15733 ( .A1(n10088), .A2(n10075), .ZN(n15864) );
  XOR2_X1 U15734 ( .A(n15865), .B(n15866), .Z(n15619) );
  XOR2_X1 U15735 ( .A(n15867), .B(n15868), .Z(n15865) );
  NOR2_X1 U15736 ( .A1(n9983), .A2(n10075), .ZN(n15868) );
  XNOR2_X1 U15737 ( .A(n15869), .B(n15870), .ZN(n15624) );
  XOR2_X1 U15738 ( .A(n15871), .B(n15872), .Z(n15869) );
  NOR2_X1 U15739 ( .A1(n10093), .A2(n10075), .ZN(n15872) );
  NOR2_X1 U15740 ( .A1(n15873), .A2(n10261), .ZN(n9039) );
  INV_X1 U15741 ( .A(n15874), .ZN(n10261) );
  NAND2_X1 U15742 ( .A1(n15875), .A2(n15876), .ZN(n15874) );
  NOR2_X1 U15743 ( .A1(n15876), .A2(n15875), .ZN(n15873) );
  XNOR2_X1 U15744 ( .A(n15877), .B(n15878), .ZN(n15875) );
  XNOR2_X1 U15745 ( .A(n15879), .B(n15880), .ZN(n15878) );
  NAND2_X1 U15746 ( .A1(n15881), .A2(n15882), .ZN(n15876) );
  NAND2_X1 U15747 ( .A1(n15883), .A2(b_9_), .ZN(n15882) );
  NOR2_X1 U15748 ( .A1(n15884), .A2(n10093), .ZN(n15883) );
  NOR2_X1 U15749 ( .A1(n15871), .A2(n15870), .ZN(n15884) );
  NAND2_X1 U15750 ( .A1(n15870), .A2(n15871), .ZN(n15881) );
  NAND2_X1 U15751 ( .A1(n15885), .A2(n15886), .ZN(n15871) );
  NAND2_X1 U15752 ( .A1(n15887), .A2(b_9_), .ZN(n15886) );
  NOR2_X1 U15753 ( .A1(n15888), .A2(n9983), .ZN(n15887) );
  NOR2_X1 U15754 ( .A1(n15866), .A2(n15867), .ZN(n15888) );
  NAND2_X1 U15755 ( .A1(n15866), .A2(n15867), .ZN(n15885) );
  NAND2_X1 U15756 ( .A1(n15889), .A2(n15890), .ZN(n15867) );
  NAND2_X1 U15757 ( .A1(n15891), .A2(b_9_), .ZN(n15890) );
  NOR2_X1 U15758 ( .A1(n15892), .A2(n10088), .ZN(n15891) );
  NOR2_X1 U15759 ( .A1(n15862), .A2(n15863), .ZN(n15892) );
  NAND2_X1 U15760 ( .A1(n15862), .A2(n15863), .ZN(n15889) );
  NAND2_X1 U15761 ( .A1(n15893), .A2(n15894), .ZN(n15863) );
  NAND2_X1 U15762 ( .A1(n15895), .A2(b_9_), .ZN(n15894) );
  NOR2_X1 U15763 ( .A1(n15896), .A2(n10086), .ZN(n15895) );
  NOR2_X1 U15764 ( .A1(n15857), .A2(n15859), .ZN(n15896) );
  NAND2_X1 U15765 ( .A1(n15857), .A2(n15859), .ZN(n15893) );
  NAND2_X1 U15766 ( .A1(n15897), .A2(n15898), .ZN(n15859) );
  NAND2_X1 U15767 ( .A1(n15899), .A2(b_9_), .ZN(n15898) );
  NOR2_X1 U15768 ( .A1(n15900), .A2(n10085), .ZN(n15899) );
  NOR2_X1 U15769 ( .A1(n15854), .A2(n15855), .ZN(n15900) );
  NAND2_X1 U15770 ( .A1(n15854), .A2(n15855), .ZN(n15897) );
  NAND2_X1 U15771 ( .A1(n15901), .A2(n15902), .ZN(n15855) );
  NAND2_X1 U15772 ( .A1(n15903), .A2(b_9_), .ZN(n15902) );
  NOR2_X1 U15773 ( .A1(n15904), .A2(n10083), .ZN(n15903) );
  NOR2_X1 U15774 ( .A1(n15850), .A2(n15851), .ZN(n15904) );
  NAND2_X1 U15775 ( .A1(n15850), .A2(n15851), .ZN(n15901) );
  NAND2_X1 U15776 ( .A1(n15905), .A2(n15906), .ZN(n15851) );
  NAND2_X1 U15777 ( .A1(n15907), .A2(b_9_), .ZN(n15906) );
  NOR2_X1 U15778 ( .A1(n15908), .A2(n10081), .ZN(n15907) );
  NOR2_X1 U15779 ( .A1(n15845), .A2(n15847), .ZN(n15908) );
  NAND2_X1 U15780 ( .A1(n15845), .A2(n15847), .ZN(n15905) );
  NAND2_X1 U15781 ( .A1(n15909), .A2(n15910), .ZN(n15847) );
  NAND2_X1 U15782 ( .A1(n15911), .A2(b_9_), .ZN(n15910) );
  NOR2_X1 U15783 ( .A1(n15912), .A2(n9773), .ZN(n15911) );
  NOR2_X1 U15784 ( .A1(n15841), .A2(n15843), .ZN(n15912) );
  NAND2_X1 U15785 ( .A1(n15841), .A2(n15843), .ZN(n15909) );
  NAND2_X1 U15786 ( .A1(n15913), .A2(n15914), .ZN(n15843) );
  NAND2_X1 U15787 ( .A1(n15915), .A2(b_9_), .ZN(n15914) );
  NOR2_X1 U15788 ( .A1(n15916), .A2(n10079), .ZN(n15915) );
  NOR2_X1 U15789 ( .A1(n15660), .A2(n15658), .ZN(n15916) );
  NAND2_X1 U15790 ( .A1(n15660), .A2(n15658), .ZN(n15913) );
  XOR2_X1 U15791 ( .A(n15917), .B(n15918), .Z(n15658) );
  XNOR2_X1 U15792 ( .A(n15919), .B(n15920), .ZN(n15918) );
  NOR2_X1 U15793 ( .A1(n15921), .A2(n15922), .ZN(n15660) );
  INV_X1 U15794 ( .A(n15923), .ZN(n15922) );
  NAND2_X1 U15795 ( .A1(n15665), .A2(n15924), .ZN(n15923) );
  NAND2_X1 U15796 ( .A1(n10077), .A2(n15667), .ZN(n15924) );
  XOR2_X1 U15797 ( .A(n15925), .B(n15926), .Z(n15665) );
  XOR2_X1 U15798 ( .A(n15927), .B(n15928), .Z(n15926) );
  NOR2_X1 U15799 ( .A1(n15667), .A2(n10077), .ZN(n15921) );
  NOR2_X1 U15800 ( .A1(n10075), .A2(n10076), .ZN(n10077) );
  NAND2_X1 U15801 ( .A1(n15929), .A2(n15930), .ZN(n15667) );
  NAND2_X1 U15802 ( .A1(n15931), .A2(b_9_), .ZN(n15930) );
  NOR2_X1 U15803 ( .A1(n15932), .A2(n10073), .ZN(n15931) );
  NOR2_X1 U15804 ( .A1(n15675), .A2(n15673), .ZN(n15932) );
  NAND2_X1 U15805 ( .A1(n15673), .A2(n15675), .ZN(n15929) );
  NAND2_X1 U15806 ( .A1(n15933), .A2(n15934), .ZN(n15675) );
  NAND2_X1 U15807 ( .A1(n15935), .A2(b_9_), .ZN(n15934) );
  NOR2_X1 U15808 ( .A1(n15936), .A2(n9649), .ZN(n15935) );
  NOR2_X1 U15809 ( .A1(n15682), .A2(n15683), .ZN(n15936) );
  NAND2_X1 U15810 ( .A1(n15682), .A2(n15683), .ZN(n15933) );
  NAND2_X1 U15811 ( .A1(n15937), .A2(n15938), .ZN(n15683) );
  NAND2_X1 U15812 ( .A1(n15939), .A2(b_9_), .ZN(n15938) );
  NOR2_X1 U15813 ( .A1(n15940), .A2(n10070), .ZN(n15939) );
  NOR2_X1 U15814 ( .A1(n15689), .A2(n15691), .ZN(n15940) );
  NAND2_X1 U15815 ( .A1(n15689), .A2(n15691), .ZN(n15937) );
  NAND2_X1 U15816 ( .A1(n15941), .A2(n15942), .ZN(n15691) );
  NAND2_X1 U15817 ( .A1(n15943), .A2(b_9_), .ZN(n15942) );
  NOR2_X1 U15818 ( .A1(n15944), .A2(n10067), .ZN(n15943) );
  NOR2_X1 U15819 ( .A1(n15699), .A2(n15697), .ZN(n15944) );
  NAND2_X1 U15820 ( .A1(n15697), .A2(n15699), .ZN(n15941) );
  NOR2_X1 U15821 ( .A1(n15945), .A2(n15946), .ZN(n15699) );
  INV_X1 U15822 ( .A(n15947), .ZN(n15946) );
  NAND2_X1 U15823 ( .A1(n15706), .A2(n15948), .ZN(n15947) );
  NAND2_X1 U15824 ( .A1(n15708), .A2(n15707), .ZN(n15948) );
  XOR2_X1 U15825 ( .A(n15949), .B(n15950), .Z(n15706) );
  XNOR2_X1 U15826 ( .A(n15951), .B(n15952), .ZN(n15950) );
  NOR2_X1 U15827 ( .A1(n15707), .A2(n15708), .ZN(n15945) );
  NOR2_X1 U15828 ( .A1(n10075), .A2(n10065), .ZN(n15708) );
  NAND2_X1 U15829 ( .A1(n15953), .A2(n15954), .ZN(n15707) );
  NAND2_X1 U15830 ( .A1(n15955), .A2(b_9_), .ZN(n15954) );
  NOR2_X1 U15831 ( .A1(n15956), .A2(n9534), .ZN(n15955) );
  NOR2_X1 U15832 ( .A1(n15715), .A2(n15713), .ZN(n15956) );
  NAND2_X1 U15833 ( .A1(n15713), .A2(n15715), .ZN(n15953) );
  NAND2_X1 U15834 ( .A1(n15957), .A2(n15958), .ZN(n15715) );
  NAND2_X1 U15835 ( .A1(n15959), .A2(b_9_), .ZN(n15958) );
  NOR2_X1 U15836 ( .A1(n15960), .A2(n10062), .ZN(n15959) );
  NOR2_X1 U15837 ( .A1(n15721), .A2(n15723), .ZN(n15960) );
  NAND2_X1 U15838 ( .A1(n15721), .A2(n15723), .ZN(n15957) );
  NAND2_X1 U15839 ( .A1(n15961), .A2(n15962), .ZN(n15723) );
  NAND2_X1 U15840 ( .A1(n15963), .A2(b_9_), .ZN(n15962) );
  NOR2_X1 U15841 ( .A1(n15964), .A2(n10060), .ZN(n15963) );
  NOR2_X1 U15842 ( .A1(n15730), .A2(n15731), .ZN(n15964) );
  NAND2_X1 U15843 ( .A1(n15730), .A2(n15731), .ZN(n15961) );
  NAND2_X1 U15844 ( .A1(n15965), .A2(n15966), .ZN(n15731) );
  NAND2_X1 U15845 ( .A1(n15967), .A2(b_9_), .ZN(n15966) );
  NOR2_X1 U15846 ( .A1(n15968), .A2(n10058), .ZN(n15967) );
  NOR2_X1 U15847 ( .A1(n15738), .A2(n15739), .ZN(n15968) );
  NAND2_X1 U15848 ( .A1(n15738), .A2(n15739), .ZN(n15965) );
  NAND2_X1 U15849 ( .A1(n15969), .A2(n15970), .ZN(n15739) );
  NAND2_X1 U15850 ( .A1(n15971), .A2(b_9_), .ZN(n15970) );
  NOR2_X1 U15851 ( .A1(n15972), .A2(n9415), .ZN(n15971) );
  NOR2_X1 U15852 ( .A1(n15839), .A2(n15837), .ZN(n15972) );
  NAND2_X1 U15853 ( .A1(n15837), .A2(n15839), .ZN(n15969) );
  NAND2_X1 U15854 ( .A1(n15973), .A2(n15974), .ZN(n15839) );
  NAND2_X1 U15855 ( .A1(n15975), .A2(b_9_), .ZN(n15974) );
  NOR2_X1 U15856 ( .A1(n15976), .A2(n10054), .ZN(n15975) );
  NOR2_X1 U15857 ( .A1(n15750), .A2(n15751), .ZN(n15976) );
  NAND2_X1 U15858 ( .A1(n15750), .A2(n15751), .ZN(n15973) );
  NAND2_X1 U15859 ( .A1(n15835), .A2(n15977), .ZN(n15751) );
  NAND2_X1 U15860 ( .A1(n15834), .A2(n15836), .ZN(n15977) );
  NAND2_X1 U15861 ( .A1(n15978), .A2(n15979), .ZN(n15836) );
  NAND2_X1 U15862 ( .A1(b_9_), .A2(a_21_), .ZN(n15979) );
  INV_X1 U15863 ( .A(n15980), .ZN(n15978) );
  XOR2_X1 U15864 ( .A(n15981), .B(n15982), .Z(n15834) );
  XOR2_X1 U15865 ( .A(n15983), .B(n15984), .Z(n15981) );
  NAND2_X1 U15866 ( .A1(a_21_), .A2(n15980), .ZN(n15835) );
  NAND2_X1 U15867 ( .A1(n15985), .A2(n15986), .ZN(n15980) );
  NAND2_X1 U15868 ( .A1(n15764), .A2(n15987), .ZN(n15986) );
  INV_X1 U15869 ( .A(n15988), .ZN(n15987) );
  NOR2_X1 U15870 ( .A1(n15763), .A2(n15762), .ZN(n15988) );
  NOR2_X1 U15871 ( .A1(n10075), .A2(n9330), .ZN(n15764) );
  NAND2_X1 U15872 ( .A1(n15762), .A2(n15763), .ZN(n15985) );
  NAND2_X1 U15873 ( .A1(n15989), .A2(n15990), .ZN(n15763) );
  NAND2_X1 U15874 ( .A1(n15832), .A2(n15991), .ZN(n15990) );
  INV_X1 U15875 ( .A(n15992), .ZN(n15991) );
  NOR2_X1 U15876 ( .A1(n15830), .A2(n15831), .ZN(n15992) );
  NOR2_X1 U15877 ( .A1(n10075), .A2(n10051), .ZN(n15832) );
  NAND2_X1 U15878 ( .A1(n15830), .A2(n15831), .ZN(n15989) );
  NAND2_X1 U15879 ( .A1(n15993), .A2(n15994), .ZN(n15831) );
  INV_X1 U15880 ( .A(n15995), .ZN(n15994) );
  NOR2_X1 U15881 ( .A1(n15828), .A2(n15996), .ZN(n15995) );
  NOR2_X1 U15882 ( .A1(n15827), .A2(n15825), .ZN(n15996) );
  NAND2_X1 U15883 ( .A1(b_9_), .A2(a_24_), .ZN(n15828) );
  NAND2_X1 U15884 ( .A1(n15825), .A2(n15827), .ZN(n15993) );
  NAND2_X1 U15885 ( .A1(n15997), .A2(n15998), .ZN(n15827) );
  NAND2_X1 U15886 ( .A1(n15824), .A2(n15999), .ZN(n15998) );
  INV_X1 U15887 ( .A(n16000), .ZN(n15999) );
  NOR2_X1 U15888 ( .A1(n15821), .A2(n15823), .ZN(n16000) );
  NOR2_X1 U15889 ( .A1(n10075), .A2(n10048), .ZN(n15824) );
  NAND2_X1 U15890 ( .A1(n15821), .A2(n15823), .ZN(n15997) );
  NOR2_X1 U15891 ( .A1(n16001), .A2(n16002), .ZN(n15823) );
  INV_X1 U15892 ( .A(n16003), .ZN(n16002) );
  NAND2_X1 U15893 ( .A1(n15817), .A2(n16004), .ZN(n16003) );
  NAND2_X1 U15894 ( .A1(n15820), .A2(n15819), .ZN(n16004) );
  XOR2_X1 U15895 ( .A(n16005), .B(n16006), .Z(n15817) );
  NAND2_X1 U15896 ( .A1(n16007), .A2(n16008), .ZN(n16005) );
  NOR2_X1 U15897 ( .A1(n15819), .A2(n15820), .ZN(n16001) );
  NOR2_X1 U15898 ( .A1(n10075), .A2(n10047), .ZN(n15820) );
  NAND2_X1 U15899 ( .A1(n15787), .A2(n16009), .ZN(n15819) );
  NAND2_X1 U15900 ( .A1(n15786), .A2(n15788), .ZN(n16009) );
  NAND2_X1 U15901 ( .A1(n16010), .A2(n16011), .ZN(n15788) );
  NAND2_X1 U15902 ( .A1(b_9_), .A2(a_27_), .ZN(n16011) );
  INV_X1 U15903 ( .A(n16012), .ZN(n16010) );
  XNOR2_X1 U15904 ( .A(n16013), .B(n16014), .ZN(n15786) );
  XOR2_X1 U15905 ( .A(n16015), .B(n16016), .Z(n16014) );
  NAND2_X1 U15906 ( .A1(b_8_), .A2(a_28_), .ZN(n16016) );
  NAND2_X1 U15907 ( .A1(a_27_), .A2(n16012), .ZN(n15787) );
  NAND2_X1 U15908 ( .A1(n16017), .A2(n16018), .ZN(n16012) );
  NAND2_X1 U15909 ( .A1(n16019), .A2(b_9_), .ZN(n16018) );
  NOR2_X1 U15910 ( .A1(n16020), .A2(n9136), .ZN(n16019) );
  NOR2_X1 U15911 ( .A1(n15793), .A2(n15795), .ZN(n16020) );
  NAND2_X1 U15912 ( .A1(n15793), .A2(n15795), .ZN(n16017) );
  NAND2_X1 U15913 ( .A1(n16021), .A2(n16022), .ZN(n15795) );
  NAND2_X1 U15914 ( .A1(n16023), .A2(b_9_), .ZN(n16022) );
  NOR2_X1 U15915 ( .A1(n16024), .A2(n9121), .ZN(n16023) );
  NOR2_X1 U15916 ( .A1(n16025), .A2(n15815), .ZN(n16024) );
  NAND2_X1 U15917 ( .A1(n16025), .A2(n15815), .ZN(n16021) );
  NAND2_X1 U15918 ( .A1(n16026), .A2(n16027), .ZN(n15815) );
  NAND2_X1 U15919 ( .A1(b_7_), .A2(n16028), .ZN(n16027) );
  NAND2_X1 U15920 ( .A1(n10486), .A2(n16029), .ZN(n16028) );
  NAND2_X1 U15921 ( .A1(a_31_), .A2(n10078), .ZN(n16029) );
  NAND2_X1 U15922 ( .A1(b_8_), .A2(n16030), .ZN(n16026) );
  NAND2_X1 U15923 ( .A1(n10489), .A2(n16031), .ZN(n16030) );
  NAND2_X1 U15924 ( .A1(a_30_), .A2(n16032), .ZN(n16031) );
  INV_X1 U15925 ( .A(n15816), .ZN(n16025) );
  NAND2_X1 U15926 ( .A1(n16033), .A2(n9025), .ZN(n15816) );
  NOR2_X1 U15927 ( .A1(n10075), .A2(n10078), .ZN(n16033) );
  XOR2_X1 U15928 ( .A(n16034), .B(n16035), .Z(n15793) );
  NOR2_X1 U15929 ( .A1(n9121), .A2(n10078), .ZN(n16035) );
  XNOR2_X1 U15930 ( .A(n16036), .B(n16037), .ZN(n16034) );
  XOR2_X1 U15931 ( .A(n16038), .B(n16039), .Z(n15821) );
  XNOR2_X1 U15932 ( .A(n16040), .B(n16041), .ZN(n16039) );
  XOR2_X1 U15933 ( .A(n16042), .B(n16043), .Z(n15825) );
  XOR2_X1 U15934 ( .A(n16044), .B(n16045), .Z(n16043) );
  XNOR2_X1 U15935 ( .A(n16046), .B(n16047), .ZN(n15830) );
  XOR2_X1 U15936 ( .A(n16048), .B(n16049), .Z(n16047) );
  XOR2_X1 U15937 ( .A(n16050), .B(n16051), .Z(n15762) );
  XOR2_X1 U15938 ( .A(n16052), .B(n16053), .Z(n16050) );
  XNOR2_X1 U15939 ( .A(n16054), .B(n16055), .ZN(n15750) );
  XOR2_X1 U15940 ( .A(n16056), .B(n16057), .Z(n16055) );
  XNOR2_X1 U15941 ( .A(n16058), .B(n16059), .ZN(n15837) );
  XNOR2_X1 U15942 ( .A(n16060), .B(n16061), .ZN(n16058) );
  XNOR2_X1 U15943 ( .A(n16062), .B(n16063), .ZN(n15738) );
  XNOR2_X1 U15944 ( .A(n16064), .B(n16065), .ZN(n16062) );
  XNOR2_X1 U15945 ( .A(n16066), .B(n16067), .ZN(n15730) );
  XOR2_X1 U15946 ( .A(n16068), .B(n16069), .Z(n16066) );
  XOR2_X1 U15947 ( .A(n16070), .B(n16071), .Z(n15721) );
  XOR2_X1 U15948 ( .A(n16072), .B(n16073), .Z(n16071) );
  XNOR2_X1 U15949 ( .A(n16074), .B(n16075), .ZN(n15713) );
  XOR2_X1 U15950 ( .A(n16076), .B(n16077), .Z(n16074) );
  XOR2_X1 U15951 ( .A(n16078), .B(n16079), .Z(n15697) );
  XNOR2_X1 U15952 ( .A(n16080), .B(n16081), .ZN(n16079) );
  XOR2_X1 U15953 ( .A(n16082), .B(n16083), .Z(n15689) );
  XOR2_X1 U15954 ( .A(n16084), .B(n16085), .Z(n16083) );
  XNOR2_X1 U15955 ( .A(n16086), .B(n16087), .ZN(n15682) );
  XOR2_X1 U15956 ( .A(n16088), .B(n16089), .Z(n16087) );
  XNOR2_X1 U15957 ( .A(n16090), .B(n16091), .ZN(n15673) );
  XNOR2_X1 U15958 ( .A(n16092), .B(n16093), .ZN(n16091) );
  XNOR2_X1 U15959 ( .A(n16094), .B(n16095), .ZN(n15841) );
  XNOR2_X1 U15960 ( .A(n16096), .B(n9742), .ZN(n16094) );
  INV_X1 U15961 ( .A(n16097), .ZN(n9742) );
  XNOR2_X1 U15962 ( .A(n16098), .B(n16099), .ZN(n15845) );
  XNOR2_X1 U15963 ( .A(n16100), .B(n16101), .ZN(n16099) );
  XOR2_X1 U15964 ( .A(n16102), .B(n16103), .Z(n15850) );
  XOR2_X1 U15965 ( .A(n16104), .B(n16105), .Z(n16102) );
  XOR2_X1 U15966 ( .A(n16106), .B(n16107), .Z(n15854) );
  XOR2_X1 U15967 ( .A(n16108), .B(n16109), .Z(n16106) );
  XOR2_X1 U15968 ( .A(n16110), .B(n16111), .Z(n15857) );
  XOR2_X1 U15969 ( .A(n16112), .B(n16113), .Z(n16110) );
  XNOR2_X1 U15970 ( .A(n16114), .B(n16115), .ZN(n15862) );
  XNOR2_X1 U15971 ( .A(n16116), .B(n16117), .ZN(n16115) );
  XNOR2_X1 U15972 ( .A(n16118), .B(n16119), .ZN(n15866) );
  XNOR2_X1 U15973 ( .A(n16120), .B(n16121), .ZN(n16118) );
  XNOR2_X1 U15974 ( .A(n16122), .B(n16123), .ZN(n15870) );
  XNOR2_X1 U15975 ( .A(n16124), .B(n16125), .ZN(n16122) );
  XNOR2_X1 U15976 ( .A(n16126), .B(n16127), .ZN(n9044) );
  NAND2_X1 U15977 ( .A1(n9052), .A2(n9053), .ZN(n9051) );
  INV_X1 U15978 ( .A(n16128), .ZN(n9053) );
  NAND2_X1 U15979 ( .A1(n16127), .A2(n16126), .ZN(n16128) );
  NAND2_X1 U15980 ( .A1(n16129), .A2(n16130), .ZN(n16126) );
  NAND2_X1 U15981 ( .A1(n15880), .A2(n16131), .ZN(n16130) );
  INV_X1 U15982 ( .A(n16132), .ZN(n16131) );
  NOR2_X1 U15983 ( .A1(n15877), .A2(n15879), .ZN(n16132) );
  NOR2_X1 U15984 ( .A1(n10078), .A2(n10093), .ZN(n15880) );
  NAND2_X1 U15985 ( .A1(n15877), .A2(n15879), .ZN(n16129) );
  NAND2_X1 U15986 ( .A1(n16133), .A2(n16134), .ZN(n15879) );
  NAND2_X1 U15987 ( .A1(n16125), .A2(n16135), .ZN(n16134) );
  NAND2_X1 U15988 ( .A1(n16124), .A2(n16123), .ZN(n16135) );
  NOR2_X1 U15989 ( .A1(n10078), .A2(n9983), .ZN(n16125) );
  INV_X1 U15990 ( .A(n16136), .ZN(n16133) );
  NOR2_X1 U15991 ( .A1(n16123), .A2(n16124), .ZN(n16136) );
  NOR2_X1 U15992 ( .A1(n16137), .A2(n16138), .ZN(n16124) );
  INV_X1 U15993 ( .A(n16139), .ZN(n16138) );
  NAND2_X1 U15994 ( .A1(n16120), .A2(n16140), .ZN(n16139) );
  NAND2_X1 U15995 ( .A1(n16119), .A2(n16121), .ZN(n16140) );
  NOR2_X1 U15996 ( .A1(n10078), .A2(n10088), .ZN(n16120) );
  NOR2_X1 U15997 ( .A1(n16119), .A2(n16121), .ZN(n16137) );
  INV_X1 U15998 ( .A(n16141), .ZN(n16121) );
  NAND2_X1 U15999 ( .A1(n16142), .A2(n16143), .ZN(n16141) );
  NAND2_X1 U16000 ( .A1(n16117), .A2(n16144), .ZN(n16143) );
  INV_X1 U16001 ( .A(n16145), .ZN(n16144) );
  NOR2_X1 U16002 ( .A1(n16114), .A2(n16116), .ZN(n16145) );
  NOR2_X1 U16003 ( .A1(n10078), .A2(n10086), .ZN(n16117) );
  NAND2_X1 U16004 ( .A1(n16114), .A2(n16116), .ZN(n16142) );
  NAND2_X1 U16005 ( .A1(n16146), .A2(n16147), .ZN(n16116) );
  NAND2_X1 U16006 ( .A1(n16113), .A2(n16148), .ZN(n16147) );
  INV_X1 U16007 ( .A(n16149), .ZN(n16148) );
  NOR2_X1 U16008 ( .A1(n16111), .A2(n16112), .ZN(n16149) );
  NOR2_X1 U16009 ( .A1(n10078), .A2(n10085), .ZN(n16113) );
  NAND2_X1 U16010 ( .A1(n16111), .A2(n16112), .ZN(n16146) );
  NAND2_X1 U16011 ( .A1(n16150), .A2(n16151), .ZN(n16112) );
  NAND2_X1 U16012 ( .A1(n16109), .A2(n16152), .ZN(n16151) );
  INV_X1 U16013 ( .A(n16153), .ZN(n16152) );
  NOR2_X1 U16014 ( .A1(n16107), .A2(n16108), .ZN(n16153) );
  NOR2_X1 U16015 ( .A1(n10078), .A2(n10083), .ZN(n16109) );
  NAND2_X1 U16016 ( .A1(n16107), .A2(n16108), .ZN(n16150) );
  NAND2_X1 U16017 ( .A1(n16154), .A2(n16155), .ZN(n16108) );
  NAND2_X1 U16018 ( .A1(n16105), .A2(n16156), .ZN(n16155) );
  INV_X1 U16019 ( .A(n16157), .ZN(n16156) );
  NOR2_X1 U16020 ( .A1(n16103), .A2(n16104), .ZN(n16157) );
  NOR2_X1 U16021 ( .A1(n10078), .A2(n10081), .ZN(n16105) );
  NAND2_X1 U16022 ( .A1(n16103), .A2(n16104), .ZN(n16154) );
  NAND2_X1 U16023 ( .A1(n16158), .A2(n16159), .ZN(n16104) );
  NAND2_X1 U16024 ( .A1(n16101), .A2(n16160), .ZN(n16159) );
  NAND2_X1 U16025 ( .A1(n16098), .A2(n16100), .ZN(n16160) );
  NOR2_X1 U16026 ( .A1(n10078), .A2(n9773), .ZN(n16101) );
  INV_X1 U16027 ( .A(n16161), .ZN(n16158) );
  NOR2_X1 U16028 ( .A1(n16098), .A2(n16100), .ZN(n16161) );
  NAND2_X1 U16029 ( .A1(n16162), .A2(n16163), .ZN(n16100) );
  NAND2_X1 U16030 ( .A1(n16095), .A2(n16164), .ZN(n16163) );
  NAND2_X1 U16031 ( .A1(n16097), .A2(n16096), .ZN(n16164) );
  XOR2_X1 U16032 ( .A(n16165), .B(n16166), .Z(n16095) );
  XOR2_X1 U16033 ( .A(n16167), .B(n16168), .Z(n16166) );
  NAND2_X1 U16034 ( .A1(b_7_), .A2(a_9_), .ZN(n16168) );
  INV_X1 U16035 ( .A(n16169), .ZN(n16162) );
  NOR2_X1 U16036 ( .A1(n16096), .A2(n16097), .ZN(n16169) );
  NOR2_X1 U16037 ( .A1(n10078), .A2(n10079), .ZN(n16097) );
  NAND2_X1 U16038 ( .A1(n16170), .A2(n16171), .ZN(n16096) );
  NAND2_X1 U16039 ( .A1(n15920), .A2(n16172), .ZN(n16171) );
  NAND2_X1 U16040 ( .A1(n16173), .A2(n15917), .ZN(n16172) );
  INV_X1 U16041 ( .A(n15919), .ZN(n16173) );
  NOR2_X1 U16042 ( .A1(n10078), .A2(n10076), .ZN(n15920) );
  NAND2_X1 U16043 ( .A1(n16174), .A2(n15919), .ZN(n16170) );
  NAND2_X1 U16044 ( .A1(n16175), .A2(n16176), .ZN(n15919) );
  INV_X1 U16045 ( .A(n16177), .ZN(n16176) );
  NOR2_X1 U16046 ( .A1(n15928), .A2(n16178), .ZN(n16177) );
  NOR2_X1 U16047 ( .A1(n15927), .A2(n15925), .ZN(n16178) );
  NAND2_X1 U16048 ( .A1(b_8_), .A2(a_10_), .ZN(n15928) );
  NAND2_X1 U16049 ( .A1(n15925), .A2(n15927), .ZN(n16175) );
  NAND2_X1 U16050 ( .A1(n16179), .A2(n16180), .ZN(n15927) );
  NAND2_X1 U16051 ( .A1(n16093), .A2(n16181), .ZN(n16180) );
  INV_X1 U16052 ( .A(n16182), .ZN(n16181) );
  NOR2_X1 U16053 ( .A1(n16092), .A2(n16090), .ZN(n16182) );
  NOR2_X1 U16054 ( .A1(n10078), .A2(n9649), .ZN(n16093) );
  NAND2_X1 U16055 ( .A1(n16090), .A2(n16092), .ZN(n16179) );
  NAND2_X1 U16056 ( .A1(n16183), .A2(n16184), .ZN(n16092) );
  INV_X1 U16057 ( .A(n16185), .ZN(n16184) );
  NOR2_X1 U16058 ( .A1(n16089), .A2(n16186), .ZN(n16185) );
  NOR2_X1 U16059 ( .A1(n16086), .A2(n16088), .ZN(n16186) );
  NAND2_X1 U16060 ( .A1(b_8_), .A2(a_12_), .ZN(n16089) );
  NAND2_X1 U16061 ( .A1(n16086), .A2(n16088), .ZN(n16183) );
  NAND2_X1 U16062 ( .A1(n16187), .A2(n16188), .ZN(n16088) );
  NAND2_X1 U16063 ( .A1(n16085), .A2(n16189), .ZN(n16188) );
  INV_X1 U16064 ( .A(n16190), .ZN(n16189) );
  NOR2_X1 U16065 ( .A1(n16082), .A2(n16084), .ZN(n16190) );
  NOR2_X1 U16066 ( .A1(n10078), .A2(n10067), .ZN(n16085) );
  NAND2_X1 U16067 ( .A1(n16082), .A2(n16084), .ZN(n16187) );
  NOR2_X1 U16068 ( .A1(n16191), .A2(n16192), .ZN(n16084) );
  INV_X1 U16069 ( .A(n16193), .ZN(n16192) );
  NAND2_X1 U16070 ( .A1(n16078), .A2(n16194), .ZN(n16193) );
  NAND2_X1 U16071 ( .A1(n16081), .A2(n16080), .ZN(n16194) );
  XNOR2_X1 U16072 ( .A(n16195), .B(n16196), .ZN(n16078) );
  XOR2_X1 U16073 ( .A(n16197), .B(n16198), .Z(n16195) );
  NOR2_X1 U16074 ( .A1(n9534), .A2(n16032), .ZN(n16198) );
  NOR2_X1 U16075 ( .A1(n16080), .A2(n16081), .ZN(n16191) );
  NOR2_X1 U16076 ( .A1(n10078), .A2(n10065), .ZN(n16081) );
  NAND2_X1 U16077 ( .A1(n16199), .A2(n16200), .ZN(n16080) );
  NAND2_X1 U16078 ( .A1(n15952), .A2(n16201), .ZN(n16200) );
  NAND2_X1 U16079 ( .A1(n15949), .A2(n15951), .ZN(n16201) );
  NOR2_X1 U16080 ( .A1(n10078), .A2(n9534), .ZN(n15952) );
  INV_X1 U16081 ( .A(n16202), .ZN(n16199) );
  NOR2_X1 U16082 ( .A1(n15949), .A2(n15951), .ZN(n16202) );
  NAND2_X1 U16083 ( .A1(n16203), .A2(n16204), .ZN(n15951) );
  NAND2_X1 U16084 ( .A1(n16075), .A2(n16205), .ZN(n16204) );
  NAND2_X1 U16085 ( .A1(n16077), .A2(n16076), .ZN(n16205) );
  XOR2_X1 U16086 ( .A(n16206), .B(n16207), .Z(n16075) );
  XOR2_X1 U16087 ( .A(n16208), .B(n16209), .Z(n16207) );
  NAND2_X1 U16088 ( .A1(b_7_), .A2(a_17_), .ZN(n16209) );
  INV_X1 U16089 ( .A(n16210), .ZN(n16203) );
  NOR2_X1 U16090 ( .A1(n16076), .A2(n16077), .ZN(n16210) );
  NOR2_X1 U16091 ( .A1(n10078), .A2(n10062), .ZN(n16077) );
  NAND2_X1 U16092 ( .A1(n16211), .A2(n16212), .ZN(n16076) );
  NAND2_X1 U16093 ( .A1(n16073), .A2(n16213), .ZN(n16212) );
  INV_X1 U16094 ( .A(n16214), .ZN(n16213) );
  NOR2_X1 U16095 ( .A1(n16070), .A2(n16072), .ZN(n16214) );
  NOR2_X1 U16096 ( .A1(n10078), .A2(n10060), .ZN(n16073) );
  NAND2_X1 U16097 ( .A1(n16070), .A2(n16072), .ZN(n16211) );
  NOR2_X1 U16098 ( .A1(n16215), .A2(n16216), .ZN(n16072) );
  INV_X1 U16099 ( .A(n16217), .ZN(n16216) );
  NAND2_X1 U16100 ( .A1(n16067), .A2(n16218), .ZN(n16217) );
  NAND2_X1 U16101 ( .A1(n16069), .A2(n16068), .ZN(n16218) );
  XOR2_X1 U16102 ( .A(n16219), .B(n16220), .Z(n16067) );
  XOR2_X1 U16103 ( .A(n16221), .B(n16222), .Z(n16220) );
  NAND2_X1 U16104 ( .A1(b_7_), .A2(a_19_), .ZN(n16222) );
  NOR2_X1 U16105 ( .A1(n16068), .A2(n16069), .ZN(n16215) );
  NOR2_X1 U16106 ( .A1(n10078), .A2(n10058), .ZN(n16069) );
  NAND2_X1 U16107 ( .A1(n16223), .A2(n16224), .ZN(n16068) );
  NAND2_X1 U16108 ( .A1(n16064), .A2(n16225), .ZN(n16224) );
  NAND2_X1 U16109 ( .A1(n16063), .A2(n16065), .ZN(n16225) );
  NOR2_X1 U16110 ( .A1(n10078), .A2(n9415), .ZN(n16064) );
  INV_X1 U16111 ( .A(n16226), .ZN(n16223) );
  NOR2_X1 U16112 ( .A1(n16063), .A2(n16065), .ZN(n16226) );
  NOR2_X1 U16113 ( .A1(n16227), .A2(n16228), .ZN(n16065) );
  INV_X1 U16114 ( .A(n16229), .ZN(n16228) );
  NAND2_X1 U16115 ( .A1(n16061), .A2(n16230), .ZN(n16229) );
  NAND2_X1 U16116 ( .A1(n16060), .A2(n16059), .ZN(n16230) );
  NOR2_X1 U16117 ( .A1(n10078), .A2(n10054), .ZN(n16061) );
  NOR2_X1 U16118 ( .A1(n16059), .A2(n16060), .ZN(n16227) );
  NOR2_X1 U16119 ( .A1(n16231), .A2(n16232), .ZN(n16060) );
  NOR2_X1 U16120 ( .A1(n16057), .A2(n16233), .ZN(n16232) );
  NOR2_X1 U16121 ( .A1(n16054), .A2(n16056), .ZN(n16233) );
  NAND2_X1 U16122 ( .A1(b_8_), .A2(a_21_), .ZN(n16057) );
  INV_X1 U16123 ( .A(n16234), .ZN(n16231) );
  NAND2_X1 U16124 ( .A1(n16054), .A2(n16056), .ZN(n16234) );
  NAND2_X1 U16125 ( .A1(n16235), .A2(n16236), .ZN(n16056) );
  NAND2_X1 U16126 ( .A1(n15984), .A2(n16237), .ZN(n16236) );
  INV_X1 U16127 ( .A(n16238), .ZN(n16237) );
  NOR2_X1 U16128 ( .A1(n15982), .A2(n15983), .ZN(n16238) );
  NOR2_X1 U16129 ( .A1(n10078), .A2(n9330), .ZN(n15984) );
  NAND2_X1 U16130 ( .A1(n15982), .A2(n15983), .ZN(n16235) );
  NAND2_X1 U16131 ( .A1(n16239), .A2(n16240), .ZN(n15983) );
  NAND2_X1 U16132 ( .A1(n16053), .A2(n16241), .ZN(n16240) );
  INV_X1 U16133 ( .A(n16242), .ZN(n16241) );
  NOR2_X1 U16134 ( .A1(n16051), .A2(n16052), .ZN(n16242) );
  NOR2_X1 U16135 ( .A1(n10078), .A2(n10051), .ZN(n16053) );
  NAND2_X1 U16136 ( .A1(n16051), .A2(n16052), .ZN(n16239) );
  NAND2_X1 U16137 ( .A1(n16243), .A2(n16244), .ZN(n16052) );
  INV_X1 U16138 ( .A(n16245), .ZN(n16244) );
  NOR2_X1 U16139 ( .A1(n16049), .A2(n16246), .ZN(n16245) );
  NOR2_X1 U16140 ( .A1(n16048), .A2(n16046), .ZN(n16246) );
  NAND2_X1 U16141 ( .A1(b_8_), .A2(a_24_), .ZN(n16049) );
  NAND2_X1 U16142 ( .A1(n16046), .A2(n16048), .ZN(n16243) );
  NAND2_X1 U16143 ( .A1(n16247), .A2(n16248), .ZN(n16048) );
  NAND2_X1 U16144 ( .A1(n16045), .A2(n16249), .ZN(n16248) );
  INV_X1 U16145 ( .A(n16250), .ZN(n16249) );
  NOR2_X1 U16146 ( .A1(n16042), .A2(n16044), .ZN(n16250) );
  NOR2_X1 U16147 ( .A1(n10078), .A2(n10048), .ZN(n16045) );
  NAND2_X1 U16148 ( .A1(n16042), .A2(n16044), .ZN(n16247) );
  NOR2_X1 U16149 ( .A1(n16251), .A2(n16252), .ZN(n16044) );
  INV_X1 U16150 ( .A(n16253), .ZN(n16252) );
  NAND2_X1 U16151 ( .A1(n16038), .A2(n16254), .ZN(n16253) );
  NAND2_X1 U16152 ( .A1(n16041), .A2(n16040), .ZN(n16254) );
  XOR2_X1 U16153 ( .A(n16255), .B(n16256), .Z(n16038) );
  NAND2_X1 U16154 ( .A1(n16257), .A2(n16258), .ZN(n16255) );
  NOR2_X1 U16155 ( .A1(n16040), .A2(n16041), .ZN(n16251) );
  NOR2_X1 U16156 ( .A1(n10078), .A2(n10047), .ZN(n16041) );
  NAND2_X1 U16157 ( .A1(n16007), .A2(n16259), .ZN(n16040) );
  NAND2_X1 U16158 ( .A1(n16006), .A2(n16008), .ZN(n16259) );
  NAND2_X1 U16159 ( .A1(n16260), .A2(n16261), .ZN(n16008) );
  NAND2_X1 U16160 ( .A1(b_8_), .A2(a_27_), .ZN(n16261) );
  INV_X1 U16161 ( .A(n16262), .ZN(n16260) );
  XNOR2_X1 U16162 ( .A(n16263), .B(n16264), .ZN(n16006) );
  XOR2_X1 U16163 ( .A(n16265), .B(n16266), .Z(n16264) );
  NAND2_X1 U16164 ( .A1(b_7_), .A2(a_28_), .ZN(n16266) );
  NAND2_X1 U16165 ( .A1(a_27_), .A2(n16262), .ZN(n16007) );
  NAND2_X1 U16166 ( .A1(n16267), .A2(n16268), .ZN(n16262) );
  NAND2_X1 U16167 ( .A1(n16269), .A2(b_8_), .ZN(n16268) );
  NOR2_X1 U16168 ( .A1(n16270), .A2(n9136), .ZN(n16269) );
  NOR2_X1 U16169 ( .A1(n16013), .A2(n16015), .ZN(n16270) );
  NAND2_X1 U16170 ( .A1(n16013), .A2(n16015), .ZN(n16267) );
  NAND2_X1 U16171 ( .A1(n16271), .A2(n16272), .ZN(n16015) );
  NAND2_X1 U16172 ( .A1(n16273), .A2(b_8_), .ZN(n16272) );
  NOR2_X1 U16173 ( .A1(n16274), .A2(n9121), .ZN(n16273) );
  NOR2_X1 U16174 ( .A1(n16275), .A2(n16036), .ZN(n16274) );
  NAND2_X1 U16175 ( .A1(n16275), .A2(n16036), .ZN(n16271) );
  NAND2_X1 U16176 ( .A1(n16276), .A2(n16277), .ZN(n16036) );
  NAND2_X1 U16177 ( .A1(b_6_), .A2(n16278), .ZN(n16277) );
  NAND2_X1 U16178 ( .A1(n10486), .A2(n16279), .ZN(n16278) );
  NAND2_X1 U16179 ( .A1(a_31_), .A2(n16032), .ZN(n16279) );
  NAND2_X1 U16180 ( .A1(b_7_), .A2(n16280), .ZN(n16276) );
  NAND2_X1 U16181 ( .A1(n10489), .A2(n16281), .ZN(n16280) );
  NAND2_X1 U16182 ( .A1(a_30_), .A2(n10080), .ZN(n16281) );
  INV_X1 U16183 ( .A(n16037), .ZN(n16275) );
  NAND2_X1 U16184 ( .A1(n16282), .A2(n9025), .ZN(n16037) );
  NOR2_X1 U16185 ( .A1(n16032), .A2(n10078), .ZN(n16282) );
  XOR2_X1 U16186 ( .A(n16283), .B(n16284), .Z(n16013) );
  NOR2_X1 U16187 ( .A1(n9121), .A2(n16032), .ZN(n16284) );
  XNOR2_X1 U16188 ( .A(n16285), .B(n16286), .ZN(n16283) );
  XOR2_X1 U16189 ( .A(n16287), .B(n16288), .Z(n16042) );
  XNOR2_X1 U16190 ( .A(n16289), .B(n16290), .ZN(n16288) );
  XOR2_X1 U16191 ( .A(n16291), .B(n16292), .Z(n16046) );
  XOR2_X1 U16192 ( .A(n16293), .B(n16294), .Z(n16292) );
  XNOR2_X1 U16193 ( .A(n16295), .B(n16296), .ZN(n16051) );
  XOR2_X1 U16194 ( .A(n16297), .B(n16298), .Z(n16296) );
  XNOR2_X1 U16195 ( .A(n16299), .B(n16300), .ZN(n15982) );
  XNOR2_X1 U16196 ( .A(n16301), .B(n16302), .ZN(n16299) );
  XNOR2_X1 U16197 ( .A(n16303), .B(n16304), .ZN(n16054) );
  NAND2_X1 U16198 ( .A1(n16305), .A2(n16306), .ZN(n16303) );
  XOR2_X1 U16199 ( .A(n16307), .B(n16308), .Z(n16059) );
  XOR2_X1 U16200 ( .A(n16309), .B(n16310), .Z(n16307) );
  XNOR2_X1 U16201 ( .A(n16311), .B(n16312), .ZN(n16063) );
  XNOR2_X1 U16202 ( .A(n16313), .B(n16314), .ZN(n16312) );
  NAND2_X1 U16203 ( .A1(b_7_), .A2(a_20_), .ZN(n16314) );
  XNOR2_X1 U16204 ( .A(n16315), .B(n16316), .ZN(n16070) );
  XOR2_X1 U16205 ( .A(n16317), .B(n16318), .Z(n16316) );
  NAND2_X1 U16206 ( .A1(b_7_), .A2(a_18_), .ZN(n16318) );
  XNOR2_X1 U16207 ( .A(n16319), .B(n16320), .ZN(n15949) );
  XOR2_X1 U16208 ( .A(n16321), .B(n16322), .Z(n16319) );
  NOR2_X1 U16209 ( .A1(n10062), .A2(n16032), .ZN(n16322) );
  XNOR2_X1 U16210 ( .A(n16323), .B(n16324), .ZN(n16082) );
  XOR2_X1 U16211 ( .A(n16325), .B(n16326), .Z(n16324) );
  NAND2_X1 U16212 ( .A1(b_7_), .A2(a_14_), .ZN(n16326) );
  XOR2_X1 U16213 ( .A(n16327), .B(n16328), .Z(n16086) );
  XOR2_X1 U16214 ( .A(n16329), .B(n16330), .Z(n16327) );
  NOR2_X1 U16215 ( .A1(n10067), .A2(n16032), .ZN(n16330) );
  XNOR2_X1 U16216 ( .A(n16331), .B(n16332), .ZN(n16090) );
  XOR2_X1 U16217 ( .A(n16333), .B(n16334), .Z(n16332) );
  NAND2_X1 U16218 ( .A1(b_7_), .A2(a_12_), .ZN(n16334) );
  XOR2_X1 U16219 ( .A(n16335), .B(n16336), .Z(n15925) );
  XOR2_X1 U16220 ( .A(n16337), .B(n16338), .Z(n16335) );
  NOR2_X1 U16221 ( .A1(n9649), .A2(n16032), .ZN(n16338) );
  INV_X1 U16222 ( .A(n15917), .ZN(n16174) );
  XOR2_X1 U16223 ( .A(n16339), .B(n16340), .Z(n15917) );
  XOR2_X1 U16224 ( .A(n16341), .B(n16342), .Z(n16340) );
  NAND2_X1 U16225 ( .A1(b_7_), .A2(a_10_), .ZN(n16342) );
  XOR2_X1 U16226 ( .A(n16343), .B(n16344), .Z(n16098) );
  XOR2_X1 U16227 ( .A(n16345), .B(n16346), .Z(n16344) );
  NAND2_X1 U16228 ( .A1(b_7_), .A2(a_8_), .ZN(n16346) );
  XOR2_X1 U16229 ( .A(n16347), .B(n16348), .Z(n16103) );
  XNOR2_X1 U16230 ( .A(n16349), .B(n9991), .ZN(n16348) );
  XNOR2_X1 U16231 ( .A(n16350), .B(n16351), .ZN(n16107) );
  XNOR2_X1 U16232 ( .A(n16352), .B(n16353), .ZN(n16351) );
  XNOR2_X1 U16233 ( .A(n16354), .B(n16355), .ZN(n16111) );
  XNOR2_X1 U16234 ( .A(n16356), .B(n16357), .ZN(n16354) );
  XNOR2_X1 U16235 ( .A(n16358), .B(n16359), .ZN(n16114) );
  XNOR2_X1 U16236 ( .A(n16360), .B(n16361), .ZN(n16358) );
  XOR2_X1 U16237 ( .A(n16362), .B(n16363), .Z(n16119) );
  XNOR2_X1 U16238 ( .A(n16364), .B(n16365), .ZN(n16362) );
  XOR2_X1 U16239 ( .A(n16366), .B(n16367), .Z(n16123) );
  XNOR2_X1 U16240 ( .A(n16368), .B(n16369), .ZN(n16366) );
  XNOR2_X1 U16241 ( .A(n16370), .B(n16371), .ZN(n15877) );
  XNOR2_X1 U16242 ( .A(n16372), .B(n16373), .ZN(n16370) );
  XNOR2_X1 U16243 ( .A(n16374), .B(n16375), .ZN(n16127) );
  XNOR2_X1 U16244 ( .A(n16376), .B(n16377), .ZN(n16375) );
  NOR2_X1 U16245 ( .A1(n16378), .A2(n10258), .ZN(n9052) );
  INV_X1 U16246 ( .A(n16379), .ZN(n10258) );
  NAND2_X1 U16247 ( .A1(n16380), .A2(n16381), .ZN(n16379) );
  NOR2_X1 U16248 ( .A1(n16381), .A2(n16380), .ZN(n16378) );
  XNOR2_X1 U16249 ( .A(n16382), .B(n16383), .ZN(n16380) );
  XNOR2_X1 U16250 ( .A(n16384), .B(n16385), .ZN(n16383) );
  NAND2_X1 U16251 ( .A1(n16386), .A2(n16387), .ZN(n16381) );
  NAND2_X1 U16252 ( .A1(n16377), .A2(n16388), .ZN(n16387) );
  NAND2_X1 U16253 ( .A1(n16389), .A2(n16390), .ZN(n16388) );
  NOR2_X1 U16254 ( .A1(n10093), .A2(n16032), .ZN(n16377) );
  NAND2_X1 U16255 ( .A1(n16374), .A2(n16376), .ZN(n16386) );
  INV_X1 U16256 ( .A(n16389), .ZN(n16376) );
  NOR2_X1 U16257 ( .A1(n16391), .A2(n16392), .ZN(n16389) );
  INV_X1 U16258 ( .A(n16393), .ZN(n16392) );
  NAND2_X1 U16259 ( .A1(n16373), .A2(n16394), .ZN(n16393) );
  NAND2_X1 U16260 ( .A1(n16372), .A2(n16371), .ZN(n16394) );
  NOR2_X1 U16261 ( .A1(n9983), .A2(n16032), .ZN(n16373) );
  NOR2_X1 U16262 ( .A1(n16371), .A2(n16372), .ZN(n16391) );
  NOR2_X1 U16263 ( .A1(n16395), .A2(n16396), .ZN(n16372) );
  INV_X1 U16264 ( .A(n16397), .ZN(n16396) );
  NAND2_X1 U16265 ( .A1(n16368), .A2(n16398), .ZN(n16397) );
  NAND2_X1 U16266 ( .A1(n16367), .A2(n16369), .ZN(n16398) );
  NOR2_X1 U16267 ( .A1(n10088), .A2(n16032), .ZN(n16368) );
  NOR2_X1 U16268 ( .A1(n16367), .A2(n16369), .ZN(n16395) );
  NOR2_X1 U16269 ( .A1(n16399), .A2(n16400), .ZN(n16369) );
  INV_X1 U16270 ( .A(n16401), .ZN(n16400) );
  NAND2_X1 U16271 ( .A1(n16365), .A2(n16402), .ZN(n16401) );
  NAND2_X1 U16272 ( .A1(n16364), .A2(n16363), .ZN(n16402) );
  NOR2_X1 U16273 ( .A1(n10086), .A2(n16032), .ZN(n16365) );
  NOR2_X1 U16274 ( .A1(n16363), .A2(n16364), .ZN(n16399) );
  NOR2_X1 U16275 ( .A1(n16403), .A2(n16404), .ZN(n16364) );
  INV_X1 U16276 ( .A(n16405), .ZN(n16404) );
  NAND2_X1 U16277 ( .A1(n16360), .A2(n16406), .ZN(n16405) );
  NAND2_X1 U16278 ( .A1(n16361), .A2(n16359), .ZN(n16406) );
  NOR2_X1 U16279 ( .A1(n10085), .A2(n16032), .ZN(n16360) );
  NOR2_X1 U16280 ( .A1(n16359), .A2(n16361), .ZN(n16403) );
  NOR2_X1 U16281 ( .A1(n16407), .A2(n16408), .ZN(n16361) );
  INV_X1 U16282 ( .A(n16409), .ZN(n16408) );
  NAND2_X1 U16283 ( .A1(n16357), .A2(n16410), .ZN(n16409) );
  NAND2_X1 U16284 ( .A1(n16356), .A2(n16355), .ZN(n16410) );
  NOR2_X1 U16285 ( .A1(n10083), .A2(n16032), .ZN(n16357) );
  NOR2_X1 U16286 ( .A1(n16355), .A2(n16356), .ZN(n16407) );
  NOR2_X1 U16287 ( .A1(n16411), .A2(n16412), .ZN(n16356) );
  INV_X1 U16288 ( .A(n16413), .ZN(n16412) );
  NAND2_X1 U16289 ( .A1(n16353), .A2(n16414), .ZN(n16413) );
  NAND2_X1 U16290 ( .A1(n16350), .A2(n16352), .ZN(n16414) );
  NOR2_X1 U16291 ( .A1(n10081), .A2(n16032), .ZN(n16353) );
  NOR2_X1 U16292 ( .A1(n16352), .A2(n16350), .ZN(n16411) );
  XOR2_X1 U16293 ( .A(n16415), .B(n16416), .Z(n16350) );
  XOR2_X1 U16294 ( .A(n16417), .B(n16418), .Z(n16416) );
  NAND2_X1 U16295 ( .A1(n16419), .A2(n16420), .ZN(n16352) );
  NAND2_X1 U16296 ( .A1(n16347), .A2(n16421), .ZN(n16420) );
  NAND2_X1 U16297 ( .A1(n9991), .A2(n16349), .ZN(n16421) );
  XOR2_X1 U16298 ( .A(n16422), .B(n16423), .Z(n16347) );
  XNOR2_X1 U16299 ( .A(n16424), .B(n16425), .ZN(n16423) );
  INV_X1 U16300 ( .A(n16426), .ZN(n16419) );
  NOR2_X1 U16301 ( .A1(n16349), .A2(n9991), .ZN(n16426) );
  NOR2_X1 U16302 ( .A1(n16032), .A2(n9773), .ZN(n9991) );
  NAND2_X1 U16303 ( .A1(n16427), .A2(n16428), .ZN(n16349) );
  NAND2_X1 U16304 ( .A1(n16429), .A2(b_7_), .ZN(n16428) );
  NOR2_X1 U16305 ( .A1(n16430), .A2(n10079), .ZN(n16429) );
  NOR2_X1 U16306 ( .A1(n16345), .A2(n16343), .ZN(n16430) );
  NAND2_X1 U16307 ( .A1(n16343), .A2(n16345), .ZN(n16427) );
  NAND2_X1 U16308 ( .A1(n16431), .A2(n16432), .ZN(n16345) );
  NAND2_X1 U16309 ( .A1(n16433), .A2(b_7_), .ZN(n16432) );
  NOR2_X1 U16310 ( .A1(n16434), .A2(n10076), .ZN(n16433) );
  NOR2_X1 U16311 ( .A1(n16165), .A2(n16167), .ZN(n16434) );
  NAND2_X1 U16312 ( .A1(n16165), .A2(n16167), .ZN(n16431) );
  NAND2_X1 U16313 ( .A1(n16435), .A2(n16436), .ZN(n16167) );
  NAND2_X1 U16314 ( .A1(n16437), .A2(b_7_), .ZN(n16436) );
  NOR2_X1 U16315 ( .A1(n16438), .A2(n10073), .ZN(n16437) );
  NOR2_X1 U16316 ( .A1(n16341), .A2(n16339), .ZN(n16438) );
  NAND2_X1 U16317 ( .A1(n16339), .A2(n16341), .ZN(n16435) );
  NAND2_X1 U16318 ( .A1(n16439), .A2(n16440), .ZN(n16341) );
  NAND2_X1 U16319 ( .A1(n16441), .A2(b_7_), .ZN(n16440) );
  NOR2_X1 U16320 ( .A1(n16442), .A2(n9649), .ZN(n16441) );
  NOR2_X1 U16321 ( .A1(n16337), .A2(n16336), .ZN(n16442) );
  NAND2_X1 U16322 ( .A1(n16336), .A2(n16337), .ZN(n16439) );
  NAND2_X1 U16323 ( .A1(n16443), .A2(n16444), .ZN(n16337) );
  NAND2_X1 U16324 ( .A1(n16445), .A2(b_7_), .ZN(n16444) );
  NOR2_X1 U16325 ( .A1(n16446), .A2(n10070), .ZN(n16445) );
  NOR2_X1 U16326 ( .A1(n16333), .A2(n16331), .ZN(n16446) );
  NAND2_X1 U16327 ( .A1(n16331), .A2(n16333), .ZN(n16443) );
  NAND2_X1 U16328 ( .A1(n16447), .A2(n16448), .ZN(n16333) );
  NAND2_X1 U16329 ( .A1(n16449), .A2(b_7_), .ZN(n16448) );
  NOR2_X1 U16330 ( .A1(n16450), .A2(n10067), .ZN(n16449) );
  NOR2_X1 U16331 ( .A1(n16328), .A2(n16329), .ZN(n16450) );
  NAND2_X1 U16332 ( .A1(n16328), .A2(n16329), .ZN(n16447) );
  NAND2_X1 U16333 ( .A1(n16451), .A2(n16452), .ZN(n16329) );
  NAND2_X1 U16334 ( .A1(n16453), .A2(b_7_), .ZN(n16452) );
  NOR2_X1 U16335 ( .A1(n16454), .A2(n10065), .ZN(n16453) );
  NOR2_X1 U16336 ( .A1(n16325), .A2(n16323), .ZN(n16454) );
  NAND2_X1 U16337 ( .A1(n16323), .A2(n16325), .ZN(n16451) );
  NAND2_X1 U16338 ( .A1(n16455), .A2(n16456), .ZN(n16325) );
  NAND2_X1 U16339 ( .A1(n16457), .A2(b_7_), .ZN(n16456) );
  NOR2_X1 U16340 ( .A1(n16458), .A2(n9534), .ZN(n16457) );
  NOR2_X1 U16341 ( .A1(n16196), .A2(n16197), .ZN(n16458) );
  NAND2_X1 U16342 ( .A1(n16196), .A2(n16197), .ZN(n16455) );
  NAND2_X1 U16343 ( .A1(n16459), .A2(n16460), .ZN(n16197) );
  NAND2_X1 U16344 ( .A1(n16461), .A2(b_7_), .ZN(n16460) );
  NOR2_X1 U16345 ( .A1(n16462), .A2(n10062), .ZN(n16461) );
  NOR2_X1 U16346 ( .A1(n16321), .A2(n16320), .ZN(n16462) );
  NAND2_X1 U16347 ( .A1(n16320), .A2(n16321), .ZN(n16459) );
  NAND2_X1 U16348 ( .A1(n16463), .A2(n16464), .ZN(n16321) );
  NAND2_X1 U16349 ( .A1(n16465), .A2(b_7_), .ZN(n16464) );
  NOR2_X1 U16350 ( .A1(n16466), .A2(n10060), .ZN(n16465) );
  NOR2_X1 U16351 ( .A1(n16208), .A2(n16206), .ZN(n16466) );
  NAND2_X1 U16352 ( .A1(n16206), .A2(n16208), .ZN(n16463) );
  NAND2_X1 U16353 ( .A1(n16467), .A2(n16468), .ZN(n16208) );
  NAND2_X1 U16354 ( .A1(n16469), .A2(b_7_), .ZN(n16468) );
  NOR2_X1 U16355 ( .A1(n16470), .A2(n10058), .ZN(n16469) );
  NOR2_X1 U16356 ( .A1(n16317), .A2(n16315), .ZN(n16470) );
  NAND2_X1 U16357 ( .A1(n16315), .A2(n16317), .ZN(n16467) );
  NAND2_X1 U16358 ( .A1(n16471), .A2(n16472), .ZN(n16317) );
  NAND2_X1 U16359 ( .A1(n16473), .A2(b_7_), .ZN(n16472) );
  NOR2_X1 U16360 ( .A1(n16474), .A2(n9415), .ZN(n16473) );
  NOR2_X1 U16361 ( .A1(n16219), .A2(n16221), .ZN(n16474) );
  NAND2_X1 U16362 ( .A1(n16219), .A2(n16221), .ZN(n16471) );
  NAND2_X1 U16363 ( .A1(n16475), .A2(n16476), .ZN(n16221) );
  NAND2_X1 U16364 ( .A1(n16477), .A2(b_7_), .ZN(n16476) );
  NOR2_X1 U16365 ( .A1(n16478), .A2(n10054), .ZN(n16477) );
  NOR2_X1 U16366 ( .A1(n16313), .A2(n16311), .ZN(n16478) );
  NAND2_X1 U16367 ( .A1(n16313), .A2(n16311), .ZN(n16475) );
  XNOR2_X1 U16368 ( .A(n16479), .B(n16480), .ZN(n16311) );
  NAND2_X1 U16369 ( .A1(n16481), .A2(n16482), .ZN(n16479) );
  NOR2_X1 U16370 ( .A1(n16483), .A2(n16484), .ZN(n16313) );
  INV_X1 U16371 ( .A(n16485), .ZN(n16484) );
  NAND2_X1 U16372 ( .A1(n16308), .A2(n16486), .ZN(n16485) );
  NAND2_X1 U16373 ( .A1(n16310), .A2(n16309), .ZN(n16486) );
  XOR2_X1 U16374 ( .A(n16487), .B(n16488), .Z(n16308) );
  NAND2_X1 U16375 ( .A1(n16489), .A2(n16490), .ZN(n16487) );
  NOR2_X1 U16376 ( .A1(n16309), .A2(n16310), .ZN(n16483) );
  NOR2_X1 U16377 ( .A1(n16032), .A2(n9358), .ZN(n16310) );
  NAND2_X1 U16378 ( .A1(n16305), .A2(n16491), .ZN(n16309) );
  NAND2_X1 U16379 ( .A1(n16304), .A2(n16306), .ZN(n16491) );
  NAND2_X1 U16380 ( .A1(n16492), .A2(n16493), .ZN(n16306) );
  NAND2_X1 U16381 ( .A1(b_7_), .A2(a_22_), .ZN(n16493) );
  INV_X1 U16382 ( .A(n16494), .ZN(n16492) );
  XNOR2_X1 U16383 ( .A(n16495), .B(n16496), .ZN(n16304) );
  XOR2_X1 U16384 ( .A(n16497), .B(n16498), .Z(n16496) );
  NAND2_X1 U16385 ( .A1(b_6_), .A2(a_23_), .ZN(n16498) );
  NAND2_X1 U16386 ( .A1(a_22_), .A2(n16494), .ZN(n16305) );
  NAND2_X1 U16387 ( .A1(n16499), .A2(n16500), .ZN(n16494) );
  NAND2_X1 U16388 ( .A1(n16302), .A2(n16501), .ZN(n16500) );
  NAND2_X1 U16389 ( .A1(n16301), .A2(n16300), .ZN(n16501) );
  NOR2_X1 U16390 ( .A1(n16032), .A2(n10051), .ZN(n16302) );
  INV_X1 U16391 ( .A(n16502), .ZN(n16499) );
  NOR2_X1 U16392 ( .A1(n16300), .A2(n16301), .ZN(n16502) );
  NOR2_X1 U16393 ( .A1(n16503), .A2(n16504), .ZN(n16301) );
  NOR2_X1 U16394 ( .A1(n16298), .A2(n16505), .ZN(n16504) );
  NOR2_X1 U16395 ( .A1(n16297), .A2(n16295), .ZN(n16505) );
  NAND2_X1 U16396 ( .A1(b_7_), .A2(a_24_), .ZN(n16298) );
  INV_X1 U16397 ( .A(n16506), .ZN(n16503) );
  NAND2_X1 U16398 ( .A1(n16295), .A2(n16297), .ZN(n16506) );
  NAND2_X1 U16399 ( .A1(n16507), .A2(n16508), .ZN(n16297) );
  NAND2_X1 U16400 ( .A1(n16294), .A2(n16509), .ZN(n16508) );
  INV_X1 U16401 ( .A(n16510), .ZN(n16509) );
  NOR2_X1 U16402 ( .A1(n16291), .A2(n16293), .ZN(n16510) );
  NOR2_X1 U16403 ( .A1(n16032), .A2(n10048), .ZN(n16294) );
  NAND2_X1 U16404 ( .A1(n16291), .A2(n16293), .ZN(n16507) );
  NOR2_X1 U16405 ( .A1(n16511), .A2(n16512), .ZN(n16293) );
  INV_X1 U16406 ( .A(n16513), .ZN(n16512) );
  NAND2_X1 U16407 ( .A1(n16287), .A2(n16514), .ZN(n16513) );
  NAND2_X1 U16408 ( .A1(n16290), .A2(n16289), .ZN(n16514) );
  XOR2_X1 U16409 ( .A(n16515), .B(n16516), .Z(n16287) );
  NAND2_X1 U16410 ( .A1(n16517), .A2(n16518), .ZN(n16515) );
  NOR2_X1 U16411 ( .A1(n16289), .A2(n16290), .ZN(n16511) );
  NOR2_X1 U16412 ( .A1(n16032), .A2(n10047), .ZN(n16290) );
  NAND2_X1 U16413 ( .A1(n16257), .A2(n16519), .ZN(n16289) );
  NAND2_X1 U16414 ( .A1(n16256), .A2(n16258), .ZN(n16519) );
  NAND2_X1 U16415 ( .A1(n16520), .A2(n16521), .ZN(n16258) );
  NAND2_X1 U16416 ( .A1(b_7_), .A2(a_27_), .ZN(n16521) );
  INV_X1 U16417 ( .A(n16522), .ZN(n16520) );
  XNOR2_X1 U16418 ( .A(n16523), .B(n16524), .ZN(n16256) );
  XOR2_X1 U16419 ( .A(n16525), .B(n16526), .Z(n16524) );
  NAND2_X1 U16420 ( .A1(b_6_), .A2(a_28_), .ZN(n16526) );
  NAND2_X1 U16421 ( .A1(a_27_), .A2(n16522), .ZN(n16257) );
  NAND2_X1 U16422 ( .A1(n16527), .A2(n16528), .ZN(n16522) );
  NAND2_X1 U16423 ( .A1(n16529), .A2(b_7_), .ZN(n16528) );
  NOR2_X1 U16424 ( .A1(n16530), .A2(n9136), .ZN(n16529) );
  NOR2_X1 U16425 ( .A1(n16263), .A2(n16265), .ZN(n16530) );
  NAND2_X1 U16426 ( .A1(n16263), .A2(n16265), .ZN(n16527) );
  NAND2_X1 U16427 ( .A1(n16531), .A2(n16532), .ZN(n16265) );
  NAND2_X1 U16428 ( .A1(n16533), .A2(b_7_), .ZN(n16532) );
  NOR2_X1 U16429 ( .A1(n16534), .A2(n9121), .ZN(n16533) );
  NOR2_X1 U16430 ( .A1(n16535), .A2(n16285), .ZN(n16534) );
  NAND2_X1 U16431 ( .A1(n16535), .A2(n16285), .ZN(n16531) );
  NAND2_X1 U16432 ( .A1(n16536), .A2(n16537), .ZN(n16285) );
  NAND2_X1 U16433 ( .A1(b_5_), .A2(n16538), .ZN(n16537) );
  NAND2_X1 U16434 ( .A1(n10486), .A2(n16539), .ZN(n16538) );
  NAND2_X1 U16435 ( .A1(a_31_), .A2(n10080), .ZN(n16539) );
  NAND2_X1 U16436 ( .A1(b_6_), .A2(n16540), .ZN(n16536) );
  NAND2_X1 U16437 ( .A1(n10489), .A2(n16541), .ZN(n16540) );
  NAND2_X1 U16438 ( .A1(a_30_), .A2(n10082), .ZN(n16541) );
  INV_X1 U16439 ( .A(n16286), .ZN(n16535) );
  NAND2_X1 U16440 ( .A1(n16542), .A2(n9025), .ZN(n16286) );
  NOR2_X1 U16441 ( .A1(n16032), .A2(n10080), .ZN(n16542) );
  XOR2_X1 U16442 ( .A(n16543), .B(n16544), .Z(n16263) );
  NOR2_X1 U16443 ( .A1(n9121), .A2(n10080), .ZN(n16544) );
  XNOR2_X1 U16444 ( .A(n16545), .B(n16546), .ZN(n16543) );
  XOR2_X1 U16445 ( .A(n16547), .B(n16548), .Z(n16291) );
  XNOR2_X1 U16446 ( .A(n16549), .B(n16550), .ZN(n16548) );
  XOR2_X1 U16447 ( .A(n16551), .B(n16552), .Z(n16295) );
  XOR2_X1 U16448 ( .A(n16553), .B(n16554), .Z(n16552) );
  XOR2_X1 U16449 ( .A(n16555), .B(n16556), .Z(n16300) );
  XOR2_X1 U16450 ( .A(n16557), .B(n16558), .Z(n16556) );
  NAND2_X1 U16451 ( .A1(b_6_), .A2(a_24_), .ZN(n16558) );
  XNOR2_X1 U16452 ( .A(n16559), .B(n16560), .ZN(n16219) );
  NAND2_X1 U16453 ( .A1(n16561), .A2(n16562), .ZN(n16559) );
  XOR2_X1 U16454 ( .A(n16563), .B(n16564), .Z(n16315) );
  XNOR2_X1 U16455 ( .A(n16565), .B(n16566), .ZN(n16564) );
  XNOR2_X1 U16456 ( .A(n16567), .B(n16568), .ZN(n16206) );
  XNOR2_X1 U16457 ( .A(n16569), .B(n16570), .ZN(n16568) );
  XNOR2_X1 U16458 ( .A(n16571), .B(n16572), .ZN(n16320) );
  XOR2_X1 U16459 ( .A(n16573), .B(n16574), .Z(n16572) );
  XNOR2_X1 U16460 ( .A(n16575), .B(n16576), .ZN(n16196) );
  XNOR2_X1 U16461 ( .A(n16577), .B(n16578), .ZN(n16576) );
  XNOR2_X1 U16462 ( .A(n16579), .B(n16580), .ZN(n16323) );
  XOR2_X1 U16463 ( .A(n16581), .B(n16582), .Z(n16580) );
  XNOR2_X1 U16464 ( .A(n16583), .B(n16584), .ZN(n16328) );
  XNOR2_X1 U16465 ( .A(n16585), .B(n16586), .ZN(n16584) );
  XNOR2_X1 U16466 ( .A(n16587), .B(n16588), .ZN(n16331) );
  XOR2_X1 U16467 ( .A(n16589), .B(n16590), .Z(n16588) );
  XOR2_X1 U16468 ( .A(n16591), .B(n16592), .Z(n16336) );
  XOR2_X1 U16469 ( .A(n16593), .B(n16594), .Z(n16592) );
  XNOR2_X1 U16470 ( .A(n16595), .B(n16596), .ZN(n16339) );
  XOR2_X1 U16471 ( .A(n16597), .B(n16598), .Z(n16596) );
  XNOR2_X1 U16472 ( .A(n16599), .B(n16600), .ZN(n16165) );
  XNOR2_X1 U16473 ( .A(n16601), .B(n16602), .ZN(n16600) );
  XNOR2_X1 U16474 ( .A(n16603), .B(n16604), .ZN(n16343) );
  XOR2_X1 U16475 ( .A(n16605), .B(n16606), .Z(n16604) );
  XNOR2_X1 U16476 ( .A(n16607), .B(n16608), .ZN(n16355) );
  XNOR2_X1 U16477 ( .A(n16609), .B(n9808), .ZN(n16608) );
  XOR2_X1 U16478 ( .A(n16610), .B(n16611), .Z(n16359) );
  XNOR2_X1 U16479 ( .A(n16612), .B(n16613), .ZN(n16611) );
  XOR2_X1 U16480 ( .A(n16614), .B(n16615), .Z(n16363) );
  XNOR2_X1 U16481 ( .A(n16616), .B(n16617), .ZN(n16615) );
  XNOR2_X1 U16482 ( .A(n16618), .B(n16619), .ZN(n16367) );
  XOR2_X1 U16483 ( .A(n16620), .B(n16621), .Z(n16618) );
  XNOR2_X1 U16484 ( .A(n16622), .B(n16623), .ZN(n16371) );
  XOR2_X1 U16485 ( .A(n16624), .B(n16625), .Z(n16622) );
  INV_X1 U16486 ( .A(n16390), .ZN(n16374) );
  XOR2_X1 U16487 ( .A(n16626), .B(n16627), .Z(n16390) );
  XNOR2_X1 U16488 ( .A(n16628), .B(n16629), .ZN(n16627) );
  XOR2_X1 U16489 ( .A(n16630), .B(n16631), .Z(n9057) );
  NAND2_X1 U16490 ( .A1(n9166), .A2(n9167), .ZN(n9165) );
  NOR2_X1 U16491 ( .A1(n16630), .A2(n16632), .ZN(n9167) );
  INV_X1 U16492 ( .A(n16631), .ZN(n16632) );
  NAND2_X1 U16493 ( .A1(n16633), .A2(n16634), .ZN(n16631) );
  NAND2_X1 U16494 ( .A1(n16385), .A2(n16635), .ZN(n16634) );
  INV_X1 U16495 ( .A(n16636), .ZN(n16635) );
  NOR2_X1 U16496 ( .A1(n16384), .A2(n16382), .ZN(n16636) );
  NOR2_X1 U16497 ( .A1(n10080), .A2(n10093), .ZN(n16385) );
  NAND2_X1 U16498 ( .A1(n16382), .A2(n16384), .ZN(n16633) );
  NAND2_X1 U16499 ( .A1(n16637), .A2(n16638), .ZN(n16384) );
  NAND2_X1 U16500 ( .A1(n16629), .A2(n16639), .ZN(n16638) );
  INV_X1 U16501 ( .A(n16640), .ZN(n16639) );
  NOR2_X1 U16502 ( .A1(n16626), .A2(n16628), .ZN(n16640) );
  NOR2_X1 U16503 ( .A1(n10080), .A2(n9983), .ZN(n16629) );
  NAND2_X1 U16504 ( .A1(n16626), .A2(n16628), .ZN(n16637) );
  NAND2_X1 U16505 ( .A1(n16641), .A2(n16642), .ZN(n16628) );
  NAND2_X1 U16506 ( .A1(n16624), .A2(n16643), .ZN(n16642) );
  INV_X1 U16507 ( .A(n16644), .ZN(n16643) );
  NOR2_X1 U16508 ( .A1(n16623), .A2(n16625), .ZN(n16644) );
  NOR2_X1 U16509 ( .A1(n10080), .A2(n10088), .ZN(n16624) );
  NAND2_X1 U16510 ( .A1(n16623), .A2(n16625), .ZN(n16641) );
  NAND2_X1 U16511 ( .A1(n16645), .A2(n16646), .ZN(n16625) );
  NAND2_X1 U16512 ( .A1(n16621), .A2(n16647), .ZN(n16646) );
  INV_X1 U16513 ( .A(n16648), .ZN(n16647) );
  NOR2_X1 U16514 ( .A1(n16620), .A2(n16619), .ZN(n16648) );
  NOR2_X1 U16515 ( .A1(n10080), .A2(n10086), .ZN(n16621) );
  NAND2_X1 U16516 ( .A1(n16619), .A2(n16620), .ZN(n16645) );
  NAND2_X1 U16517 ( .A1(n16649), .A2(n16650), .ZN(n16620) );
  NAND2_X1 U16518 ( .A1(n16617), .A2(n16651), .ZN(n16650) );
  INV_X1 U16519 ( .A(n16652), .ZN(n16651) );
  NOR2_X1 U16520 ( .A1(n16614), .A2(n16616), .ZN(n16652) );
  NOR2_X1 U16521 ( .A1(n10080), .A2(n10085), .ZN(n16617) );
  NAND2_X1 U16522 ( .A1(n16614), .A2(n16616), .ZN(n16649) );
  NAND2_X1 U16523 ( .A1(n16653), .A2(n16654), .ZN(n16616) );
  NAND2_X1 U16524 ( .A1(n16613), .A2(n16655), .ZN(n16654) );
  NAND2_X1 U16525 ( .A1(n16610), .A2(n16612), .ZN(n16655) );
  NOR2_X1 U16526 ( .A1(n10080), .A2(n10083), .ZN(n16613) );
  INV_X1 U16527 ( .A(n16656), .ZN(n16653) );
  NOR2_X1 U16528 ( .A1(n16610), .A2(n16612), .ZN(n16656) );
  NAND2_X1 U16529 ( .A1(n16657), .A2(n16658), .ZN(n16612) );
  NAND2_X1 U16530 ( .A1(n16607), .A2(n16659), .ZN(n16658) );
  INV_X1 U16531 ( .A(n16660), .ZN(n16659) );
  NOR2_X1 U16532 ( .A1(n9808), .A2(n16609), .ZN(n16660) );
  XNOR2_X1 U16533 ( .A(n16661), .B(n16662), .ZN(n16607) );
  XOR2_X1 U16534 ( .A(n16663), .B(n16664), .Z(n16661) );
  NOR2_X1 U16535 ( .A1(n9773), .A2(n10082), .ZN(n16664) );
  NAND2_X1 U16536 ( .A1(n16609), .A2(n9808), .ZN(n16657) );
  NAND2_X1 U16537 ( .A1(b_6_), .A2(a_6_), .ZN(n9808) );
  NOR2_X1 U16538 ( .A1(n16665), .A2(n16666), .ZN(n16609) );
  NOR2_X1 U16539 ( .A1(n16418), .A2(n16667), .ZN(n16666) );
  NOR2_X1 U16540 ( .A1(n16417), .A2(n16415), .ZN(n16667) );
  NAND2_X1 U16541 ( .A1(b_6_), .A2(a_7_), .ZN(n16418) );
  INV_X1 U16542 ( .A(n16668), .ZN(n16665) );
  NAND2_X1 U16543 ( .A1(n16415), .A2(n16417), .ZN(n16668) );
  NAND2_X1 U16544 ( .A1(n16669), .A2(n16670), .ZN(n16417) );
  NAND2_X1 U16545 ( .A1(n16425), .A2(n16671), .ZN(n16670) );
  NAND2_X1 U16546 ( .A1(n16672), .A2(n16673), .ZN(n16671) );
  INV_X1 U16547 ( .A(n16424), .ZN(n16673) );
  INV_X1 U16548 ( .A(n16422), .ZN(n16672) );
  NOR2_X1 U16549 ( .A1(n10080), .A2(n10079), .ZN(n16425) );
  NAND2_X1 U16550 ( .A1(n16422), .A2(n16424), .ZN(n16669) );
  NAND2_X1 U16551 ( .A1(n16674), .A2(n16675), .ZN(n16424) );
  INV_X1 U16552 ( .A(n16676), .ZN(n16675) );
  NOR2_X1 U16553 ( .A1(n16606), .A2(n16677), .ZN(n16676) );
  NOR2_X1 U16554 ( .A1(n16605), .A2(n16603), .ZN(n16677) );
  NAND2_X1 U16555 ( .A1(b_6_), .A2(a_9_), .ZN(n16606) );
  NAND2_X1 U16556 ( .A1(n16603), .A2(n16605), .ZN(n16674) );
  NAND2_X1 U16557 ( .A1(n16678), .A2(n16679), .ZN(n16605) );
  NAND2_X1 U16558 ( .A1(n16602), .A2(n16680), .ZN(n16679) );
  NAND2_X1 U16559 ( .A1(n16681), .A2(n16682), .ZN(n16680) );
  INV_X1 U16560 ( .A(n16601), .ZN(n16682) );
  INV_X1 U16561 ( .A(n16599), .ZN(n16681) );
  NOR2_X1 U16562 ( .A1(n10080), .A2(n10073), .ZN(n16602) );
  NAND2_X1 U16563 ( .A1(n16599), .A2(n16601), .ZN(n16678) );
  NAND2_X1 U16564 ( .A1(n16683), .A2(n16684), .ZN(n16601) );
  INV_X1 U16565 ( .A(n16685), .ZN(n16684) );
  NOR2_X1 U16566 ( .A1(n16598), .A2(n16686), .ZN(n16685) );
  NOR2_X1 U16567 ( .A1(n16597), .A2(n16595), .ZN(n16686) );
  NAND2_X1 U16568 ( .A1(b_6_), .A2(a_11_), .ZN(n16598) );
  NAND2_X1 U16569 ( .A1(n16595), .A2(n16597), .ZN(n16683) );
  NAND2_X1 U16570 ( .A1(n16687), .A2(n16688), .ZN(n16597) );
  NAND2_X1 U16571 ( .A1(n16594), .A2(n16689), .ZN(n16688) );
  NAND2_X1 U16572 ( .A1(n16593), .A2(n16591), .ZN(n16689) );
  NOR2_X1 U16573 ( .A1(n10080), .A2(n10070), .ZN(n16594) );
  INV_X1 U16574 ( .A(n16690), .ZN(n16687) );
  NOR2_X1 U16575 ( .A1(n16591), .A2(n16593), .ZN(n16690) );
  NOR2_X1 U16576 ( .A1(n16691), .A2(n16692), .ZN(n16593) );
  NOR2_X1 U16577 ( .A1(n16590), .A2(n16693), .ZN(n16692) );
  NOR2_X1 U16578 ( .A1(n16589), .A2(n16587), .ZN(n16693) );
  NAND2_X1 U16579 ( .A1(b_6_), .A2(a_13_), .ZN(n16590) );
  INV_X1 U16580 ( .A(n16694), .ZN(n16691) );
  NAND2_X1 U16581 ( .A1(n16587), .A2(n16589), .ZN(n16694) );
  NAND2_X1 U16582 ( .A1(n16695), .A2(n16696), .ZN(n16589) );
  NAND2_X1 U16583 ( .A1(n16586), .A2(n16697), .ZN(n16696) );
  INV_X1 U16584 ( .A(n16698), .ZN(n16697) );
  NOR2_X1 U16585 ( .A1(n16583), .A2(n16585), .ZN(n16698) );
  NOR2_X1 U16586 ( .A1(n10080), .A2(n10065), .ZN(n16586) );
  NAND2_X1 U16587 ( .A1(n16583), .A2(n16585), .ZN(n16695) );
  NAND2_X1 U16588 ( .A1(n16699), .A2(n16700), .ZN(n16585) );
  INV_X1 U16589 ( .A(n16701), .ZN(n16700) );
  NOR2_X1 U16590 ( .A1(n16582), .A2(n16702), .ZN(n16701) );
  NOR2_X1 U16591 ( .A1(n16581), .A2(n16579), .ZN(n16702) );
  NAND2_X1 U16592 ( .A1(b_6_), .A2(a_15_), .ZN(n16582) );
  NAND2_X1 U16593 ( .A1(n16579), .A2(n16581), .ZN(n16699) );
  NAND2_X1 U16594 ( .A1(n16703), .A2(n16704), .ZN(n16581) );
  NAND2_X1 U16595 ( .A1(n16578), .A2(n16705), .ZN(n16704) );
  INV_X1 U16596 ( .A(n16706), .ZN(n16705) );
  NOR2_X1 U16597 ( .A1(n16575), .A2(n16577), .ZN(n16706) );
  NOR2_X1 U16598 ( .A1(n10080), .A2(n10062), .ZN(n16578) );
  NAND2_X1 U16599 ( .A1(n16575), .A2(n16577), .ZN(n16703) );
  NAND2_X1 U16600 ( .A1(n16707), .A2(n16708), .ZN(n16577) );
  INV_X1 U16601 ( .A(n16709), .ZN(n16708) );
  NOR2_X1 U16602 ( .A1(n16574), .A2(n16710), .ZN(n16709) );
  NOR2_X1 U16603 ( .A1(n16573), .A2(n16571), .ZN(n16710) );
  NAND2_X1 U16604 ( .A1(b_6_), .A2(a_17_), .ZN(n16574) );
  NAND2_X1 U16605 ( .A1(n16571), .A2(n16573), .ZN(n16707) );
  NAND2_X1 U16606 ( .A1(n16711), .A2(n16712), .ZN(n16573) );
  NAND2_X1 U16607 ( .A1(n16570), .A2(n16713), .ZN(n16712) );
  NAND2_X1 U16608 ( .A1(n16567), .A2(n16569), .ZN(n16713) );
  NOR2_X1 U16609 ( .A1(n10080), .A2(n10058), .ZN(n16570) );
  INV_X1 U16610 ( .A(n16714), .ZN(n16711) );
  NOR2_X1 U16611 ( .A1(n16569), .A2(n16567), .ZN(n16714) );
  XNOR2_X1 U16612 ( .A(n16715), .B(n16716), .ZN(n16567) );
  XOR2_X1 U16613 ( .A(n16717), .B(n16718), .Z(n16715) );
  NOR2_X1 U16614 ( .A1(n9415), .A2(n10082), .ZN(n16718) );
  NAND2_X1 U16615 ( .A1(n16719), .A2(n16720), .ZN(n16569) );
  NAND2_X1 U16616 ( .A1(n16563), .A2(n16721), .ZN(n16720) );
  NAND2_X1 U16617 ( .A1(n16566), .A2(n16565), .ZN(n16721) );
  XNOR2_X1 U16618 ( .A(n16722), .B(n16723), .ZN(n16563) );
  XOR2_X1 U16619 ( .A(n16724), .B(n16725), .Z(n16722) );
  NOR2_X1 U16620 ( .A1(n10054), .A2(n10082), .ZN(n16725) );
  INV_X1 U16621 ( .A(n16726), .ZN(n16719) );
  NOR2_X1 U16622 ( .A1(n16565), .A2(n16566), .ZN(n16726) );
  NOR2_X1 U16623 ( .A1(n10080), .A2(n9415), .ZN(n16566) );
  NAND2_X1 U16624 ( .A1(n16561), .A2(n16727), .ZN(n16565) );
  NAND2_X1 U16625 ( .A1(n16560), .A2(n16562), .ZN(n16727) );
  NAND2_X1 U16626 ( .A1(n16728), .A2(n16729), .ZN(n16562) );
  NAND2_X1 U16627 ( .A1(b_6_), .A2(a_20_), .ZN(n16729) );
  INV_X1 U16628 ( .A(n16730), .ZN(n16728) );
  XNOR2_X1 U16629 ( .A(n16731), .B(n16732), .ZN(n16560) );
  XOR2_X1 U16630 ( .A(n16733), .B(n16734), .Z(n16732) );
  NAND2_X1 U16631 ( .A1(b_5_), .A2(a_21_), .ZN(n16734) );
  NAND2_X1 U16632 ( .A1(a_20_), .A2(n16730), .ZN(n16561) );
  NAND2_X1 U16633 ( .A1(n16481), .A2(n16735), .ZN(n16730) );
  NAND2_X1 U16634 ( .A1(n16480), .A2(n16482), .ZN(n16735) );
  NAND2_X1 U16635 ( .A1(n16736), .A2(n16737), .ZN(n16482) );
  NAND2_X1 U16636 ( .A1(b_6_), .A2(a_21_), .ZN(n16737) );
  INV_X1 U16637 ( .A(n16738), .ZN(n16736) );
  XNOR2_X1 U16638 ( .A(n16739), .B(n16740), .ZN(n16480) );
  XOR2_X1 U16639 ( .A(n16741), .B(n16742), .Z(n16740) );
  NAND2_X1 U16640 ( .A1(b_5_), .A2(a_22_), .ZN(n16742) );
  NAND2_X1 U16641 ( .A1(a_21_), .A2(n16738), .ZN(n16481) );
  NAND2_X1 U16642 ( .A1(n16489), .A2(n16743), .ZN(n16738) );
  NAND2_X1 U16643 ( .A1(n16488), .A2(n16490), .ZN(n16743) );
  NAND2_X1 U16644 ( .A1(n16744), .A2(n16745), .ZN(n16490) );
  NAND2_X1 U16645 ( .A1(b_6_), .A2(a_22_), .ZN(n16745) );
  INV_X1 U16646 ( .A(n16746), .ZN(n16744) );
  XNOR2_X1 U16647 ( .A(n16747), .B(n16748), .ZN(n16488) );
  XOR2_X1 U16648 ( .A(n16749), .B(n16750), .Z(n16748) );
  NAND2_X1 U16649 ( .A1(b_5_), .A2(a_23_), .ZN(n16750) );
  NAND2_X1 U16650 ( .A1(a_22_), .A2(n16746), .ZN(n16489) );
  NAND2_X1 U16651 ( .A1(n16751), .A2(n16752), .ZN(n16746) );
  NAND2_X1 U16652 ( .A1(n16753), .A2(b_6_), .ZN(n16752) );
  NOR2_X1 U16653 ( .A1(n16754), .A2(n10051), .ZN(n16753) );
  NOR2_X1 U16654 ( .A1(n16495), .A2(n16497), .ZN(n16754) );
  NAND2_X1 U16655 ( .A1(n16495), .A2(n16497), .ZN(n16751) );
  NAND2_X1 U16656 ( .A1(n16755), .A2(n16756), .ZN(n16497) );
  NAND2_X1 U16657 ( .A1(n16757), .A2(b_6_), .ZN(n16756) );
  NOR2_X1 U16658 ( .A1(n16758), .A2(n10050), .ZN(n16757) );
  NOR2_X1 U16659 ( .A1(n16557), .A2(n16555), .ZN(n16758) );
  NAND2_X1 U16660 ( .A1(n16555), .A2(n16557), .ZN(n16755) );
  NAND2_X1 U16661 ( .A1(n16759), .A2(n16760), .ZN(n16557) );
  NAND2_X1 U16662 ( .A1(n16554), .A2(n16761), .ZN(n16760) );
  INV_X1 U16663 ( .A(n16762), .ZN(n16761) );
  NOR2_X1 U16664 ( .A1(n16551), .A2(n16553), .ZN(n16762) );
  NOR2_X1 U16665 ( .A1(n10080), .A2(n10048), .ZN(n16554) );
  NAND2_X1 U16666 ( .A1(n16551), .A2(n16553), .ZN(n16759) );
  NOR2_X1 U16667 ( .A1(n16763), .A2(n16764), .ZN(n16553) );
  INV_X1 U16668 ( .A(n16765), .ZN(n16764) );
  NAND2_X1 U16669 ( .A1(n16547), .A2(n16766), .ZN(n16765) );
  NAND2_X1 U16670 ( .A1(n16550), .A2(n16549), .ZN(n16766) );
  XOR2_X1 U16671 ( .A(n16767), .B(n16768), .Z(n16547) );
  NAND2_X1 U16672 ( .A1(n16769), .A2(n16770), .ZN(n16767) );
  NOR2_X1 U16673 ( .A1(n16549), .A2(n16550), .ZN(n16763) );
  NOR2_X1 U16674 ( .A1(n10080), .A2(n10047), .ZN(n16550) );
  NAND2_X1 U16675 ( .A1(n16517), .A2(n16771), .ZN(n16549) );
  NAND2_X1 U16676 ( .A1(n16516), .A2(n16518), .ZN(n16771) );
  NAND2_X1 U16677 ( .A1(n16772), .A2(n16773), .ZN(n16518) );
  NAND2_X1 U16678 ( .A1(b_6_), .A2(a_27_), .ZN(n16773) );
  INV_X1 U16679 ( .A(n16774), .ZN(n16772) );
  XNOR2_X1 U16680 ( .A(n16775), .B(n16776), .ZN(n16516) );
  XOR2_X1 U16681 ( .A(n16777), .B(n16778), .Z(n16776) );
  NAND2_X1 U16682 ( .A1(b_5_), .A2(a_28_), .ZN(n16778) );
  NAND2_X1 U16683 ( .A1(a_27_), .A2(n16774), .ZN(n16517) );
  NAND2_X1 U16684 ( .A1(n16779), .A2(n16780), .ZN(n16774) );
  NAND2_X1 U16685 ( .A1(n16781), .A2(b_6_), .ZN(n16780) );
  NOR2_X1 U16686 ( .A1(n16782), .A2(n9136), .ZN(n16781) );
  NOR2_X1 U16687 ( .A1(n16523), .A2(n16525), .ZN(n16782) );
  NAND2_X1 U16688 ( .A1(n16523), .A2(n16525), .ZN(n16779) );
  NAND2_X1 U16689 ( .A1(n16783), .A2(n16784), .ZN(n16525) );
  NAND2_X1 U16690 ( .A1(n16785), .A2(b_6_), .ZN(n16784) );
  NOR2_X1 U16691 ( .A1(n16786), .A2(n9121), .ZN(n16785) );
  NOR2_X1 U16692 ( .A1(n16787), .A2(n16545), .ZN(n16786) );
  NAND2_X1 U16693 ( .A1(n16787), .A2(n16545), .ZN(n16783) );
  NAND2_X1 U16694 ( .A1(n16788), .A2(n16789), .ZN(n16545) );
  NAND2_X1 U16695 ( .A1(b_4_), .A2(n16790), .ZN(n16789) );
  NAND2_X1 U16696 ( .A1(n10486), .A2(n16791), .ZN(n16790) );
  NAND2_X1 U16697 ( .A1(a_31_), .A2(n10082), .ZN(n16791) );
  NAND2_X1 U16698 ( .A1(b_5_), .A2(n16792), .ZN(n16788) );
  NAND2_X1 U16699 ( .A1(n10489), .A2(n16793), .ZN(n16792) );
  NAND2_X1 U16700 ( .A1(a_30_), .A2(n10084), .ZN(n16793) );
  INV_X1 U16701 ( .A(n16546), .ZN(n16787) );
  NAND2_X1 U16702 ( .A1(n16794), .A2(n9025), .ZN(n16546) );
  NOR2_X1 U16703 ( .A1(n10080), .A2(n10082), .ZN(n16794) );
  XOR2_X1 U16704 ( .A(n16795), .B(n16796), .Z(n16523) );
  NOR2_X1 U16705 ( .A1(n9121), .A2(n10082), .ZN(n16796) );
  XNOR2_X1 U16706 ( .A(n16797), .B(n16798), .ZN(n16795) );
  XOR2_X1 U16707 ( .A(n16799), .B(n16800), .Z(n16551) );
  XNOR2_X1 U16708 ( .A(n16801), .B(n16802), .ZN(n16800) );
  XNOR2_X1 U16709 ( .A(n16803), .B(n16804), .ZN(n16555) );
  XNOR2_X1 U16710 ( .A(n16805), .B(n16806), .ZN(n16804) );
  XNOR2_X1 U16711 ( .A(n16807), .B(n16808), .ZN(n16495) );
  XOR2_X1 U16712 ( .A(n16809), .B(n16810), .Z(n16808) );
  NAND2_X1 U16713 ( .A1(b_5_), .A2(a_24_), .ZN(n16810) );
  XOR2_X1 U16714 ( .A(n16811), .B(n16812), .Z(n16571) );
  XOR2_X1 U16715 ( .A(n16813), .B(n16814), .Z(n16811) );
  NOR2_X1 U16716 ( .A1(n10058), .A2(n10082), .ZN(n16814) );
  XOR2_X1 U16717 ( .A(n16815), .B(n16816), .Z(n16575) );
  XOR2_X1 U16718 ( .A(n16817), .B(n16818), .Z(n16815) );
  NOR2_X1 U16719 ( .A1(n10060), .A2(n10082), .ZN(n16818) );
  XOR2_X1 U16720 ( .A(n16819), .B(n16820), .Z(n16579) );
  XOR2_X1 U16721 ( .A(n16821), .B(n16822), .Z(n16819) );
  NOR2_X1 U16722 ( .A1(n10062), .A2(n10082), .ZN(n16822) );
  XOR2_X1 U16723 ( .A(n16823), .B(n16824), .Z(n16583) );
  XOR2_X1 U16724 ( .A(n16825), .B(n16826), .Z(n16823) );
  NOR2_X1 U16725 ( .A1(n9534), .A2(n10082), .ZN(n16826) );
  XOR2_X1 U16726 ( .A(n16827), .B(n16828), .Z(n16587) );
  XOR2_X1 U16727 ( .A(n16829), .B(n16830), .Z(n16827) );
  NOR2_X1 U16728 ( .A1(n10065), .A2(n10082), .ZN(n16830) );
  XNOR2_X1 U16729 ( .A(n16831), .B(n16832), .ZN(n16591) );
  XOR2_X1 U16730 ( .A(n16833), .B(n16834), .Z(n16831) );
  NOR2_X1 U16731 ( .A1(n10067), .A2(n10082), .ZN(n16834) );
  XOR2_X1 U16732 ( .A(n16835), .B(n16836), .Z(n16595) );
  XOR2_X1 U16733 ( .A(n16837), .B(n16838), .Z(n16835) );
  NOR2_X1 U16734 ( .A1(n10070), .A2(n10082), .ZN(n16838) );
  XOR2_X1 U16735 ( .A(n16839), .B(n16840), .Z(n16599) );
  XOR2_X1 U16736 ( .A(n16841), .B(n16842), .Z(n16839) );
  NOR2_X1 U16737 ( .A1(n9649), .A2(n10082), .ZN(n16842) );
  XOR2_X1 U16738 ( .A(n16843), .B(n16844), .Z(n16603) );
  XOR2_X1 U16739 ( .A(n16845), .B(n16846), .Z(n16843) );
  NOR2_X1 U16740 ( .A1(n10073), .A2(n10082), .ZN(n16846) );
  XOR2_X1 U16741 ( .A(n16847), .B(n16848), .Z(n16422) );
  XOR2_X1 U16742 ( .A(n16849), .B(n16850), .Z(n16847) );
  NOR2_X1 U16743 ( .A1(n10076), .A2(n10082), .ZN(n16850) );
  XOR2_X1 U16744 ( .A(n16851), .B(n16852), .Z(n16415) );
  XOR2_X1 U16745 ( .A(n16853), .B(n16854), .Z(n16851) );
  NOR2_X1 U16746 ( .A1(n10079), .A2(n10082), .ZN(n16854) );
  XNOR2_X1 U16747 ( .A(n16855), .B(n16856), .ZN(n16610) );
  XOR2_X1 U16748 ( .A(n16857), .B(n16858), .Z(n16855) );
  NOR2_X1 U16749 ( .A1(n10081), .A2(n10082), .ZN(n16858) );
  XOR2_X1 U16750 ( .A(n16859), .B(n16860), .Z(n16614) );
  XNOR2_X1 U16751 ( .A(n16861), .B(n9837), .ZN(n16859) );
  XOR2_X1 U16752 ( .A(n16862), .B(n16863), .Z(n16619) );
  XNOR2_X1 U16753 ( .A(n16864), .B(n16865), .ZN(n16862) );
  NAND2_X1 U16754 ( .A1(b_5_), .A2(a_4_), .ZN(n16864) );
  XOR2_X1 U16755 ( .A(n16866), .B(n16867), .Z(n16623) );
  XOR2_X1 U16756 ( .A(n16868), .B(n16869), .Z(n16866) );
  NOR2_X1 U16757 ( .A1(n10086), .A2(n10082), .ZN(n16869) );
  XOR2_X1 U16758 ( .A(n16870), .B(n16871), .Z(n16626) );
  XOR2_X1 U16759 ( .A(n16872), .B(n16873), .Z(n16870) );
  NOR2_X1 U16760 ( .A1(n10088), .A2(n10082), .ZN(n16873) );
  XOR2_X1 U16761 ( .A(n16874), .B(n16875), .Z(n16382) );
  XOR2_X1 U16762 ( .A(n16876), .B(n16877), .Z(n16874) );
  NOR2_X1 U16763 ( .A1(n9983), .A2(n10082), .ZN(n16877) );
  XNOR2_X1 U16764 ( .A(n16878), .B(n16879), .ZN(n16630) );
  XOR2_X1 U16765 ( .A(n16880), .B(n16881), .Z(n16878) );
  NOR2_X1 U16766 ( .A1(n10093), .A2(n10082), .ZN(n16881) );
  NOR2_X1 U16767 ( .A1(n16882), .A2(n10255), .ZN(n9166) );
  INV_X1 U16768 ( .A(n16883), .ZN(n10255) );
  NAND2_X1 U16769 ( .A1(n16884), .A2(n16885), .ZN(n16883) );
  NOR2_X1 U16770 ( .A1(n16885), .A2(n16884), .ZN(n16882) );
  XNOR2_X1 U16771 ( .A(n16886), .B(n16887), .ZN(n16884) );
  XNOR2_X1 U16772 ( .A(n16888), .B(n16889), .ZN(n16886) );
  NAND2_X1 U16773 ( .A1(n16890), .A2(n16891), .ZN(n16885) );
  NAND2_X1 U16774 ( .A1(n16892), .A2(b_5_), .ZN(n16891) );
  NOR2_X1 U16775 ( .A1(n16893), .A2(n10093), .ZN(n16892) );
  NOR2_X1 U16776 ( .A1(n16879), .A2(n16880), .ZN(n16893) );
  NAND2_X1 U16777 ( .A1(n16879), .A2(n16880), .ZN(n16890) );
  NAND2_X1 U16778 ( .A1(n16894), .A2(n16895), .ZN(n16880) );
  NAND2_X1 U16779 ( .A1(n16896), .A2(b_5_), .ZN(n16895) );
  NOR2_X1 U16780 ( .A1(n16897), .A2(n9983), .ZN(n16896) );
  NOR2_X1 U16781 ( .A1(n16876), .A2(n16875), .ZN(n16897) );
  NAND2_X1 U16782 ( .A1(n16875), .A2(n16876), .ZN(n16894) );
  NAND2_X1 U16783 ( .A1(n16898), .A2(n16899), .ZN(n16876) );
  NAND2_X1 U16784 ( .A1(n16900), .A2(b_5_), .ZN(n16899) );
  NOR2_X1 U16785 ( .A1(n16901), .A2(n10088), .ZN(n16900) );
  NOR2_X1 U16786 ( .A1(n16871), .A2(n16872), .ZN(n16901) );
  NAND2_X1 U16787 ( .A1(n16871), .A2(n16872), .ZN(n16898) );
  NAND2_X1 U16788 ( .A1(n16902), .A2(n16903), .ZN(n16872) );
  NAND2_X1 U16789 ( .A1(n16904), .A2(b_5_), .ZN(n16903) );
  NOR2_X1 U16790 ( .A1(n16905), .A2(n10086), .ZN(n16904) );
  NOR2_X1 U16791 ( .A1(n16867), .A2(n16868), .ZN(n16905) );
  NAND2_X1 U16792 ( .A1(n16867), .A2(n16868), .ZN(n16902) );
  NAND2_X1 U16793 ( .A1(n16906), .A2(n16907), .ZN(n16868) );
  NAND2_X1 U16794 ( .A1(n16908), .A2(b_5_), .ZN(n16907) );
  NOR2_X1 U16795 ( .A1(n16909), .A2(n10085), .ZN(n16908) );
  NOR2_X1 U16796 ( .A1(n16865), .A2(n16863), .ZN(n16909) );
  NAND2_X1 U16797 ( .A1(n16863), .A2(n16865), .ZN(n16906) );
  NAND2_X1 U16798 ( .A1(n16910), .A2(n16911), .ZN(n16865) );
  NAND2_X1 U16799 ( .A1(n16860), .A2(n16912), .ZN(n16911) );
  NAND2_X1 U16800 ( .A1(n16913), .A2(n9837), .ZN(n16912) );
  INV_X1 U16801 ( .A(n16861), .ZN(n16913) );
  XNOR2_X1 U16802 ( .A(n16914), .B(n16915), .ZN(n16860) );
  XNOR2_X1 U16803 ( .A(n16916), .B(n16917), .ZN(n16915) );
  NAND2_X1 U16804 ( .A1(n16918), .A2(n16861), .ZN(n16910) );
  NAND2_X1 U16805 ( .A1(n16919), .A2(n16920), .ZN(n16861) );
  NAND2_X1 U16806 ( .A1(n16921), .A2(b_5_), .ZN(n16920) );
  NOR2_X1 U16807 ( .A1(n16922), .A2(n10081), .ZN(n16921) );
  NOR2_X1 U16808 ( .A1(n16857), .A2(n16856), .ZN(n16922) );
  NAND2_X1 U16809 ( .A1(n16856), .A2(n16857), .ZN(n16919) );
  NAND2_X1 U16810 ( .A1(n16923), .A2(n16924), .ZN(n16857) );
  NAND2_X1 U16811 ( .A1(n16925), .A2(b_5_), .ZN(n16924) );
  NOR2_X1 U16812 ( .A1(n16926), .A2(n9773), .ZN(n16925) );
  NOR2_X1 U16813 ( .A1(n16662), .A2(n16663), .ZN(n16926) );
  NAND2_X1 U16814 ( .A1(n16662), .A2(n16663), .ZN(n16923) );
  NAND2_X1 U16815 ( .A1(n16927), .A2(n16928), .ZN(n16663) );
  NAND2_X1 U16816 ( .A1(n16929), .A2(b_5_), .ZN(n16928) );
  NOR2_X1 U16817 ( .A1(n16930), .A2(n10079), .ZN(n16929) );
  NOR2_X1 U16818 ( .A1(n16853), .A2(n16852), .ZN(n16930) );
  NAND2_X1 U16819 ( .A1(n16852), .A2(n16853), .ZN(n16927) );
  NAND2_X1 U16820 ( .A1(n16931), .A2(n16932), .ZN(n16853) );
  NAND2_X1 U16821 ( .A1(n16933), .A2(b_5_), .ZN(n16932) );
  NOR2_X1 U16822 ( .A1(n16934), .A2(n10076), .ZN(n16933) );
  NOR2_X1 U16823 ( .A1(n16848), .A2(n16849), .ZN(n16934) );
  NAND2_X1 U16824 ( .A1(n16848), .A2(n16849), .ZN(n16931) );
  NAND2_X1 U16825 ( .A1(n16935), .A2(n16936), .ZN(n16849) );
  NAND2_X1 U16826 ( .A1(n16937), .A2(b_5_), .ZN(n16936) );
  NOR2_X1 U16827 ( .A1(n16938), .A2(n10073), .ZN(n16937) );
  NOR2_X1 U16828 ( .A1(n16845), .A2(n16844), .ZN(n16938) );
  NAND2_X1 U16829 ( .A1(n16844), .A2(n16845), .ZN(n16935) );
  NAND2_X1 U16830 ( .A1(n16939), .A2(n16940), .ZN(n16845) );
  NAND2_X1 U16831 ( .A1(n16941), .A2(b_5_), .ZN(n16940) );
  NOR2_X1 U16832 ( .A1(n16942), .A2(n9649), .ZN(n16941) );
  NOR2_X1 U16833 ( .A1(n16840), .A2(n16841), .ZN(n16942) );
  NAND2_X1 U16834 ( .A1(n16840), .A2(n16841), .ZN(n16939) );
  NAND2_X1 U16835 ( .A1(n16943), .A2(n16944), .ZN(n16841) );
  NAND2_X1 U16836 ( .A1(n16945), .A2(b_5_), .ZN(n16944) );
  NOR2_X1 U16837 ( .A1(n16946), .A2(n10070), .ZN(n16945) );
  NOR2_X1 U16838 ( .A1(n16837), .A2(n16836), .ZN(n16946) );
  NAND2_X1 U16839 ( .A1(n16836), .A2(n16837), .ZN(n16943) );
  NAND2_X1 U16840 ( .A1(n16947), .A2(n16948), .ZN(n16837) );
  NAND2_X1 U16841 ( .A1(n16949), .A2(b_5_), .ZN(n16948) );
  NOR2_X1 U16842 ( .A1(n16950), .A2(n10067), .ZN(n16949) );
  NOR2_X1 U16843 ( .A1(n16833), .A2(n16832), .ZN(n16950) );
  NAND2_X1 U16844 ( .A1(n16832), .A2(n16833), .ZN(n16947) );
  NAND2_X1 U16845 ( .A1(n16951), .A2(n16952), .ZN(n16833) );
  NAND2_X1 U16846 ( .A1(n16953), .A2(b_5_), .ZN(n16952) );
  NOR2_X1 U16847 ( .A1(n16954), .A2(n10065), .ZN(n16953) );
  NOR2_X1 U16848 ( .A1(n16829), .A2(n16828), .ZN(n16954) );
  NAND2_X1 U16849 ( .A1(n16828), .A2(n16829), .ZN(n16951) );
  NAND2_X1 U16850 ( .A1(n16955), .A2(n16956), .ZN(n16829) );
  NAND2_X1 U16851 ( .A1(n16957), .A2(b_5_), .ZN(n16956) );
  NOR2_X1 U16852 ( .A1(n16958), .A2(n9534), .ZN(n16957) );
  NOR2_X1 U16853 ( .A1(n16824), .A2(n16825), .ZN(n16958) );
  NAND2_X1 U16854 ( .A1(n16824), .A2(n16825), .ZN(n16955) );
  NAND2_X1 U16855 ( .A1(n16959), .A2(n16960), .ZN(n16825) );
  NAND2_X1 U16856 ( .A1(n16961), .A2(b_5_), .ZN(n16960) );
  NOR2_X1 U16857 ( .A1(n16962), .A2(n10062), .ZN(n16961) );
  NOR2_X1 U16858 ( .A1(n16821), .A2(n16820), .ZN(n16962) );
  NAND2_X1 U16859 ( .A1(n16820), .A2(n16821), .ZN(n16959) );
  NAND2_X1 U16860 ( .A1(n16963), .A2(n16964), .ZN(n16821) );
  NAND2_X1 U16861 ( .A1(n16965), .A2(b_5_), .ZN(n16964) );
  NOR2_X1 U16862 ( .A1(n16966), .A2(n10060), .ZN(n16965) );
  NOR2_X1 U16863 ( .A1(n16816), .A2(n16817), .ZN(n16966) );
  NAND2_X1 U16864 ( .A1(n16816), .A2(n16817), .ZN(n16963) );
  NAND2_X1 U16865 ( .A1(n16967), .A2(n16968), .ZN(n16817) );
  NAND2_X1 U16866 ( .A1(n16969), .A2(b_5_), .ZN(n16968) );
  NOR2_X1 U16867 ( .A1(n16970), .A2(n10058), .ZN(n16969) );
  NOR2_X1 U16868 ( .A1(n16813), .A2(n16812), .ZN(n16970) );
  NAND2_X1 U16869 ( .A1(n16812), .A2(n16813), .ZN(n16967) );
  NAND2_X1 U16870 ( .A1(n16971), .A2(n16972), .ZN(n16813) );
  NAND2_X1 U16871 ( .A1(n16973), .A2(b_5_), .ZN(n16972) );
  NOR2_X1 U16872 ( .A1(n16974), .A2(n9415), .ZN(n16973) );
  NOR2_X1 U16873 ( .A1(n16716), .A2(n16717), .ZN(n16974) );
  NAND2_X1 U16874 ( .A1(n16716), .A2(n16717), .ZN(n16971) );
  NAND2_X1 U16875 ( .A1(n16975), .A2(n16976), .ZN(n16717) );
  NAND2_X1 U16876 ( .A1(n16977), .A2(b_5_), .ZN(n16976) );
  NOR2_X1 U16877 ( .A1(n16978), .A2(n10054), .ZN(n16977) );
  NOR2_X1 U16878 ( .A1(n16724), .A2(n16723), .ZN(n16978) );
  NAND2_X1 U16879 ( .A1(n16723), .A2(n16724), .ZN(n16975) );
  NAND2_X1 U16880 ( .A1(n16979), .A2(n16980), .ZN(n16724) );
  NAND2_X1 U16881 ( .A1(n16981), .A2(b_5_), .ZN(n16980) );
  NOR2_X1 U16882 ( .A1(n16982), .A2(n9358), .ZN(n16981) );
  NOR2_X1 U16883 ( .A1(n16733), .A2(n16731), .ZN(n16982) );
  NAND2_X1 U16884 ( .A1(n16731), .A2(n16733), .ZN(n16979) );
  NAND2_X1 U16885 ( .A1(n16983), .A2(n16984), .ZN(n16733) );
  NAND2_X1 U16886 ( .A1(n16985), .A2(b_5_), .ZN(n16984) );
  NOR2_X1 U16887 ( .A1(n16986), .A2(n9330), .ZN(n16985) );
  NOR2_X1 U16888 ( .A1(n16739), .A2(n16741), .ZN(n16986) );
  NAND2_X1 U16889 ( .A1(n16739), .A2(n16741), .ZN(n16983) );
  NAND2_X1 U16890 ( .A1(n16987), .A2(n16988), .ZN(n16741) );
  NAND2_X1 U16891 ( .A1(n16989), .A2(b_5_), .ZN(n16988) );
  NOR2_X1 U16892 ( .A1(n16990), .A2(n10051), .ZN(n16989) );
  NOR2_X1 U16893 ( .A1(n16747), .A2(n16749), .ZN(n16990) );
  NAND2_X1 U16894 ( .A1(n16747), .A2(n16749), .ZN(n16987) );
  NAND2_X1 U16895 ( .A1(n16991), .A2(n16992), .ZN(n16749) );
  NAND2_X1 U16896 ( .A1(n16993), .A2(b_5_), .ZN(n16992) );
  NOR2_X1 U16897 ( .A1(n16994), .A2(n10050), .ZN(n16993) );
  NOR2_X1 U16898 ( .A1(n16809), .A2(n16807), .ZN(n16994) );
  NAND2_X1 U16899 ( .A1(n16807), .A2(n16809), .ZN(n16991) );
  NAND2_X1 U16900 ( .A1(n16995), .A2(n16996), .ZN(n16809) );
  NAND2_X1 U16901 ( .A1(n16806), .A2(n16997), .ZN(n16996) );
  NAND2_X1 U16902 ( .A1(n16803), .A2(n16805), .ZN(n16997) );
  NOR2_X1 U16903 ( .A1(n10082), .A2(n10048), .ZN(n16806) );
  INV_X1 U16904 ( .A(n16998), .ZN(n16995) );
  NOR2_X1 U16905 ( .A1(n16805), .A2(n16803), .ZN(n16998) );
  XNOR2_X1 U16906 ( .A(n16999), .B(n17000), .ZN(n16803) );
  XNOR2_X1 U16907 ( .A(n17001), .B(n17002), .ZN(n17000) );
  NAND2_X1 U16908 ( .A1(n17003), .A2(n17004), .ZN(n16805) );
  NAND2_X1 U16909 ( .A1(n16799), .A2(n17005), .ZN(n17004) );
  NAND2_X1 U16910 ( .A1(n16802), .A2(n16801), .ZN(n17005) );
  XOR2_X1 U16911 ( .A(n17006), .B(n17007), .Z(n16799) );
  NAND2_X1 U16912 ( .A1(n17008), .A2(n17009), .ZN(n17006) );
  INV_X1 U16913 ( .A(n17010), .ZN(n17003) );
  NOR2_X1 U16914 ( .A1(n16801), .A2(n16802), .ZN(n17010) );
  NOR2_X1 U16915 ( .A1(n10082), .A2(n10047), .ZN(n16802) );
  NAND2_X1 U16916 ( .A1(n16769), .A2(n17011), .ZN(n16801) );
  NAND2_X1 U16917 ( .A1(n16768), .A2(n16770), .ZN(n17011) );
  NAND2_X1 U16918 ( .A1(n17012), .A2(n17013), .ZN(n16770) );
  NAND2_X1 U16919 ( .A1(b_5_), .A2(a_27_), .ZN(n17013) );
  INV_X1 U16920 ( .A(n17014), .ZN(n17012) );
  XNOR2_X1 U16921 ( .A(n17015), .B(n17016), .ZN(n16768) );
  XOR2_X1 U16922 ( .A(n17017), .B(n17018), .Z(n17016) );
  NAND2_X1 U16923 ( .A1(b_4_), .A2(a_28_), .ZN(n17018) );
  NAND2_X1 U16924 ( .A1(a_27_), .A2(n17014), .ZN(n16769) );
  NAND2_X1 U16925 ( .A1(n17019), .A2(n17020), .ZN(n17014) );
  NAND2_X1 U16926 ( .A1(n17021), .A2(b_5_), .ZN(n17020) );
  NOR2_X1 U16927 ( .A1(n17022), .A2(n9136), .ZN(n17021) );
  NOR2_X1 U16928 ( .A1(n16775), .A2(n16777), .ZN(n17022) );
  NAND2_X1 U16929 ( .A1(n16775), .A2(n16777), .ZN(n17019) );
  NAND2_X1 U16930 ( .A1(n17023), .A2(n17024), .ZN(n16777) );
  NAND2_X1 U16931 ( .A1(n17025), .A2(b_5_), .ZN(n17024) );
  NOR2_X1 U16932 ( .A1(n17026), .A2(n9121), .ZN(n17025) );
  NOR2_X1 U16933 ( .A1(n17027), .A2(n16797), .ZN(n17026) );
  NAND2_X1 U16934 ( .A1(n17027), .A2(n16797), .ZN(n17023) );
  NAND2_X1 U16935 ( .A1(n17028), .A2(n17029), .ZN(n16797) );
  NAND2_X1 U16936 ( .A1(b_3_), .A2(n17030), .ZN(n17029) );
  NAND2_X1 U16937 ( .A1(n10486), .A2(n17031), .ZN(n17030) );
  NAND2_X1 U16938 ( .A1(a_31_), .A2(n10084), .ZN(n17031) );
  NAND2_X1 U16939 ( .A1(b_4_), .A2(n17032), .ZN(n17028) );
  NAND2_X1 U16940 ( .A1(n10489), .A2(n17033), .ZN(n17032) );
  NAND2_X1 U16941 ( .A1(a_30_), .A2(n9888), .ZN(n17033) );
  INV_X1 U16942 ( .A(n16798), .ZN(n17027) );
  NAND2_X1 U16943 ( .A1(n17034), .A2(n9025), .ZN(n16798) );
  NOR2_X1 U16944 ( .A1(n10082), .A2(n10084), .ZN(n17034) );
  XOR2_X1 U16945 ( .A(n17035), .B(n17036), .Z(n16775) );
  NOR2_X1 U16946 ( .A1(n9121), .A2(n10084), .ZN(n17036) );
  XNOR2_X1 U16947 ( .A(n17037), .B(n17038), .ZN(n17035) );
  XNOR2_X1 U16948 ( .A(n17039), .B(n17040), .ZN(n16807) );
  XNOR2_X1 U16949 ( .A(n17041), .B(n17042), .ZN(n17040) );
  XNOR2_X1 U16950 ( .A(n17043), .B(n17044), .ZN(n16747) );
  XOR2_X1 U16951 ( .A(n17045), .B(n17046), .Z(n17044) );
  XOR2_X1 U16952 ( .A(n17047), .B(n17048), .Z(n16739) );
  XNOR2_X1 U16953 ( .A(n17049), .B(n17050), .ZN(n17047) );
  XNOR2_X1 U16954 ( .A(n17051), .B(n17052), .ZN(n16731) );
  XNOR2_X1 U16955 ( .A(n17053), .B(n17054), .ZN(n17051) );
  XNOR2_X1 U16956 ( .A(n17055), .B(n17056), .ZN(n16723) );
  XNOR2_X1 U16957 ( .A(n17057), .B(n17058), .ZN(n17055) );
  XNOR2_X1 U16958 ( .A(n17059), .B(n17060), .ZN(n16716) );
  XNOR2_X1 U16959 ( .A(n17061), .B(n17062), .ZN(n17059) );
  XOR2_X1 U16960 ( .A(n17063), .B(n17064), .Z(n16812) );
  XOR2_X1 U16961 ( .A(n17065), .B(n17066), .Z(n17063) );
  XNOR2_X1 U16962 ( .A(n17067), .B(n17068), .ZN(n16816) );
  XNOR2_X1 U16963 ( .A(n17069), .B(n17070), .ZN(n17068) );
  XOR2_X1 U16964 ( .A(n17071), .B(n17072), .Z(n16820) );
  XOR2_X1 U16965 ( .A(n17073), .B(n17074), .Z(n17071) );
  XNOR2_X1 U16966 ( .A(n17075), .B(n17076), .ZN(n16824) );
  XNOR2_X1 U16967 ( .A(n17077), .B(n17078), .ZN(n17076) );
  XOR2_X1 U16968 ( .A(n17079), .B(n17080), .Z(n16828) );
  XOR2_X1 U16969 ( .A(n17081), .B(n17082), .Z(n17079) );
  XNOR2_X1 U16970 ( .A(n17083), .B(n17084), .ZN(n16832) );
  XNOR2_X1 U16971 ( .A(n17085), .B(n17086), .ZN(n17084) );
  XNOR2_X1 U16972 ( .A(n17087), .B(n17088), .ZN(n16836) );
  XOR2_X1 U16973 ( .A(n17089), .B(n17090), .Z(n17088) );
  XNOR2_X1 U16974 ( .A(n17091), .B(n17092), .ZN(n16840) );
  XNOR2_X1 U16975 ( .A(n17093), .B(n17094), .ZN(n17092) );
  XOR2_X1 U16976 ( .A(n17095), .B(n17096), .Z(n16844) );
  XOR2_X1 U16977 ( .A(n17097), .B(n17098), .Z(n17095) );
  XNOR2_X1 U16978 ( .A(n17099), .B(n17100), .ZN(n16848) );
  XNOR2_X1 U16979 ( .A(n17101), .B(n17102), .ZN(n17100) );
  XOR2_X1 U16980 ( .A(n17103), .B(n17104), .Z(n16852) );
  XOR2_X1 U16981 ( .A(n17105), .B(n17106), .Z(n17103) );
  XNOR2_X1 U16982 ( .A(n17107), .B(n17108), .ZN(n16662) );
  XNOR2_X1 U16983 ( .A(n17109), .B(n17110), .ZN(n17108) );
  XOR2_X1 U16984 ( .A(n17111), .B(n17112), .Z(n16856) );
  XOR2_X1 U16985 ( .A(n17113), .B(n17114), .Z(n17111) );
  INV_X1 U16986 ( .A(n9837), .ZN(n16918) );
  NAND2_X1 U16987 ( .A1(b_5_), .A2(a_5_), .ZN(n9837) );
  XNOR2_X1 U16988 ( .A(n17115), .B(n17116), .ZN(n16863) );
  XNOR2_X1 U16989 ( .A(n17117), .B(n17118), .ZN(n17115) );
  XOR2_X1 U16990 ( .A(n17119), .B(n17120), .Z(n16867) );
  XNOR2_X1 U16991 ( .A(n17121), .B(n9866), .ZN(n17120) );
  XNOR2_X1 U16992 ( .A(n17122), .B(n17123), .ZN(n16871) );
  XNOR2_X1 U16993 ( .A(n17124), .B(n17125), .ZN(n17123) );
  XNOR2_X1 U16994 ( .A(n17126), .B(n17127), .ZN(n16875) );
  XNOR2_X1 U16995 ( .A(n17128), .B(n17129), .ZN(n17127) );
  XNOR2_X1 U16996 ( .A(n17130), .B(n17131), .ZN(n16879) );
  XNOR2_X1 U16997 ( .A(n17132), .B(n17133), .ZN(n17131) );
  XOR2_X1 U16998 ( .A(n17134), .B(n17135), .Z(n9454) );
  NAND2_X1 U16999 ( .A1(n9751), .A2(n9752), .ZN(n9750) );
  NOR2_X1 U17000 ( .A1(n17135), .A2(n17136), .ZN(n9752) );
  INV_X1 U17001 ( .A(n17134), .ZN(n17136) );
  NAND2_X1 U17002 ( .A1(n17137), .A2(n17138), .ZN(n17134) );
  NAND2_X1 U17003 ( .A1(n16889), .A2(n17139), .ZN(n17138) );
  INV_X1 U17004 ( .A(n17140), .ZN(n17139) );
  NOR2_X1 U17005 ( .A1(n16887), .A2(n16888), .ZN(n17140) );
  NOR2_X1 U17006 ( .A1(n10084), .A2(n10093), .ZN(n16889) );
  NAND2_X1 U17007 ( .A1(n16887), .A2(n16888), .ZN(n17137) );
  NAND2_X1 U17008 ( .A1(n17141), .A2(n17142), .ZN(n16888) );
  NAND2_X1 U17009 ( .A1(n17133), .A2(n17143), .ZN(n17142) );
  INV_X1 U17010 ( .A(n17144), .ZN(n17143) );
  NOR2_X1 U17011 ( .A1(n17130), .A2(n17132), .ZN(n17144) );
  NOR2_X1 U17012 ( .A1(n10084), .A2(n9983), .ZN(n17133) );
  NAND2_X1 U17013 ( .A1(n17130), .A2(n17132), .ZN(n17141) );
  NAND2_X1 U17014 ( .A1(n17145), .A2(n17146), .ZN(n17132) );
  NAND2_X1 U17015 ( .A1(n17129), .A2(n17147), .ZN(n17146) );
  NAND2_X1 U17016 ( .A1(n17148), .A2(n17149), .ZN(n17147) );
  NOR2_X1 U17017 ( .A1(n10084), .A2(n10088), .ZN(n17129) );
  NAND2_X1 U17018 ( .A1(n17126), .A2(n17128), .ZN(n17145) );
  INV_X1 U17019 ( .A(n17148), .ZN(n17128) );
  NOR2_X1 U17020 ( .A1(n17150), .A2(n17151), .ZN(n17148) );
  INV_X1 U17021 ( .A(n17152), .ZN(n17151) );
  NAND2_X1 U17022 ( .A1(n17125), .A2(n17153), .ZN(n17152) );
  NAND2_X1 U17023 ( .A1(n17122), .A2(n17124), .ZN(n17153) );
  NOR2_X1 U17024 ( .A1(n10084), .A2(n10086), .ZN(n17125) );
  NOR2_X1 U17025 ( .A1(n17122), .A2(n17124), .ZN(n17150) );
  NAND2_X1 U17026 ( .A1(n17154), .A2(n17155), .ZN(n17124) );
  NAND2_X1 U17027 ( .A1(n17119), .A2(n17156), .ZN(n17155) );
  INV_X1 U17028 ( .A(n17157), .ZN(n17156) );
  NOR2_X1 U17029 ( .A1(n9866), .A2(n17121), .ZN(n17157) );
  XOR2_X1 U17030 ( .A(n17158), .B(n17159), .Z(n17119) );
  NAND2_X1 U17031 ( .A1(n17160), .A2(n17161), .ZN(n17158) );
  NAND2_X1 U17032 ( .A1(n17121), .A2(n9866), .ZN(n17154) );
  NAND2_X1 U17033 ( .A1(b_4_), .A2(a_4_), .ZN(n9866) );
  NOR2_X1 U17034 ( .A1(n17162), .A2(n17163), .ZN(n17121) );
  INV_X1 U17035 ( .A(n17164), .ZN(n17163) );
  NAND2_X1 U17036 ( .A1(n17118), .A2(n17165), .ZN(n17164) );
  NAND2_X1 U17037 ( .A1(n17117), .A2(n17116), .ZN(n17165) );
  NOR2_X1 U17038 ( .A1(n10084), .A2(n10083), .ZN(n17118) );
  NOR2_X1 U17039 ( .A1(n17116), .A2(n17117), .ZN(n17162) );
  INV_X1 U17040 ( .A(n17166), .ZN(n17117) );
  NAND2_X1 U17041 ( .A1(n17167), .A2(n17168), .ZN(n17166) );
  NAND2_X1 U17042 ( .A1(n16917), .A2(n17169), .ZN(n17168) );
  INV_X1 U17043 ( .A(n17170), .ZN(n17169) );
  NOR2_X1 U17044 ( .A1(n16914), .A2(n16916), .ZN(n17170) );
  NOR2_X1 U17045 ( .A1(n10084), .A2(n10081), .ZN(n16917) );
  NAND2_X1 U17046 ( .A1(n16914), .A2(n16916), .ZN(n17167) );
  NAND2_X1 U17047 ( .A1(n17171), .A2(n17172), .ZN(n16916) );
  NAND2_X1 U17048 ( .A1(n17114), .A2(n17173), .ZN(n17172) );
  INV_X1 U17049 ( .A(n17174), .ZN(n17173) );
  NOR2_X1 U17050 ( .A1(n17113), .A2(n17112), .ZN(n17174) );
  NOR2_X1 U17051 ( .A1(n10084), .A2(n9773), .ZN(n17114) );
  NAND2_X1 U17052 ( .A1(n17112), .A2(n17113), .ZN(n17171) );
  NAND2_X1 U17053 ( .A1(n17175), .A2(n17176), .ZN(n17113) );
  NAND2_X1 U17054 ( .A1(n17110), .A2(n17177), .ZN(n17176) );
  INV_X1 U17055 ( .A(n17178), .ZN(n17177) );
  NOR2_X1 U17056 ( .A1(n17107), .A2(n17109), .ZN(n17178) );
  NOR2_X1 U17057 ( .A1(n10084), .A2(n10079), .ZN(n17110) );
  NAND2_X1 U17058 ( .A1(n17107), .A2(n17109), .ZN(n17175) );
  NAND2_X1 U17059 ( .A1(n17179), .A2(n17180), .ZN(n17109) );
  NAND2_X1 U17060 ( .A1(n17106), .A2(n17181), .ZN(n17180) );
  INV_X1 U17061 ( .A(n17182), .ZN(n17181) );
  NOR2_X1 U17062 ( .A1(n17105), .A2(n17104), .ZN(n17182) );
  NOR2_X1 U17063 ( .A1(n10084), .A2(n10076), .ZN(n17106) );
  NAND2_X1 U17064 ( .A1(n17104), .A2(n17105), .ZN(n17179) );
  NAND2_X1 U17065 ( .A1(n17183), .A2(n17184), .ZN(n17105) );
  NAND2_X1 U17066 ( .A1(n17102), .A2(n17185), .ZN(n17184) );
  INV_X1 U17067 ( .A(n17186), .ZN(n17185) );
  NOR2_X1 U17068 ( .A1(n17099), .A2(n17101), .ZN(n17186) );
  NOR2_X1 U17069 ( .A1(n10084), .A2(n10073), .ZN(n17102) );
  NAND2_X1 U17070 ( .A1(n17099), .A2(n17101), .ZN(n17183) );
  NAND2_X1 U17071 ( .A1(n17187), .A2(n17188), .ZN(n17101) );
  NAND2_X1 U17072 ( .A1(n17098), .A2(n17189), .ZN(n17188) );
  INV_X1 U17073 ( .A(n17190), .ZN(n17189) );
  NOR2_X1 U17074 ( .A1(n17097), .A2(n17096), .ZN(n17190) );
  NOR2_X1 U17075 ( .A1(n10084), .A2(n9649), .ZN(n17098) );
  NAND2_X1 U17076 ( .A1(n17096), .A2(n17097), .ZN(n17187) );
  NAND2_X1 U17077 ( .A1(n17191), .A2(n17192), .ZN(n17097) );
  NAND2_X1 U17078 ( .A1(n17094), .A2(n17193), .ZN(n17192) );
  INV_X1 U17079 ( .A(n17194), .ZN(n17193) );
  NOR2_X1 U17080 ( .A1(n17091), .A2(n17093), .ZN(n17194) );
  NOR2_X1 U17081 ( .A1(n10084), .A2(n10070), .ZN(n17094) );
  NAND2_X1 U17082 ( .A1(n17091), .A2(n17093), .ZN(n17191) );
  NAND2_X1 U17083 ( .A1(n17195), .A2(n17196), .ZN(n17093) );
  INV_X1 U17084 ( .A(n17197), .ZN(n17196) );
  NOR2_X1 U17085 ( .A1(n17090), .A2(n17198), .ZN(n17197) );
  NOR2_X1 U17086 ( .A1(n17089), .A2(n17087), .ZN(n17198) );
  NAND2_X1 U17087 ( .A1(b_4_), .A2(a_13_), .ZN(n17090) );
  NAND2_X1 U17088 ( .A1(n17087), .A2(n17089), .ZN(n17195) );
  NAND2_X1 U17089 ( .A1(n17199), .A2(n17200), .ZN(n17089) );
  NAND2_X1 U17090 ( .A1(n17086), .A2(n17201), .ZN(n17200) );
  INV_X1 U17091 ( .A(n17202), .ZN(n17201) );
  NOR2_X1 U17092 ( .A1(n17085), .A2(n17083), .ZN(n17202) );
  NOR2_X1 U17093 ( .A1(n10084), .A2(n10065), .ZN(n17086) );
  NAND2_X1 U17094 ( .A1(n17083), .A2(n17085), .ZN(n17199) );
  NAND2_X1 U17095 ( .A1(n17203), .A2(n17204), .ZN(n17085) );
  NAND2_X1 U17096 ( .A1(n17082), .A2(n17205), .ZN(n17204) );
  INV_X1 U17097 ( .A(n17206), .ZN(n17205) );
  NOR2_X1 U17098 ( .A1(n17081), .A2(n17080), .ZN(n17206) );
  NOR2_X1 U17099 ( .A1(n10084), .A2(n9534), .ZN(n17082) );
  NAND2_X1 U17100 ( .A1(n17080), .A2(n17081), .ZN(n17203) );
  NAND2_X1 U17101 ( .A1(n17207), .A2(n17208), .ZN(n17081) );
  NAND2_X1 U17102 ( .A1(n17078), .A2(n17209), .ZN(n17208) );
  INV_X1 U17103 ( .A(n17210), .ZN(n17209) );
  NOR2_X1 U17104 ( .A1(n17075), .A2(n17077), .ZN(n17210) );
  NOR2_X1 U17105 ( .A1(n10084), .A2(n10062), .ZN(n17078) );
  NAND2_X1 U17106 ( .A1(n17075), .A2(n17077), .ZN(n17207) );
  NAND2_X1 U17107 ( .A1(n17211), .A2(n17212), .ZN(n17077) );
  NAND2_X1 U17108 ( .A1(n17074), .A2(n17213), .ZN(n17212) );
  INV_X1 U17109 ( .A(n17214), .ZN(n17213) );
  NOR2_X1 U17110 ( .A1(n17073), .A2(n17072), .ZN(n17214) );
  NOR2_X1 U17111 ( .A1(n10084), .A2(n10060), .ZN(n17074) );
  NAND2_X1 U17112 ( .A1(n17072), .A2(n17073), .ZN(n17211) );
  NAND2_X1 U17113 ( .A1(n17215), .A2(n17216), .ZN(n17073) );
  NAND2_X1 U17114 ( .A1(n17070), .A2(n17217), .ZN(n17216) );
  INV_X1 U17115 ( .A(n17218), .ZN(n17217) );
  NOR2_X1 U17116 ( .A1(n17067), .A2(n17069), .ZN(n17218) );
  NOR2_X1 U17117 ( .A1(n10084), .A2(n10058), .ZN(n17070) );
  NAND2_X1 U17118 ( .A1(n17067), .A2(n17069), .ZN(n17215) );
  NAND2_X1 U17119 ( .A1(n17219), .A2(n17220), .ZN(n17069) );
  NAND2_X1 U17120 ( .A1(n17066), .A2(n17221), .ZN(n17220) );
  INV_X1 U17121 ( .A(n17222), .ZN(n17221) );
  NOR2_X1 U17122 ( .A1(n17065), .A2(n17064), .ZN(n17222) );
  NOR2_X1 U17123 ( .A1(n10084), .A2(n9415), .ZN(n17066) );
  NAND2_X1 U17124 ( .A1(n17064), .A2(n17065), .ZN(n17219) );
  NAND2_X1 U17125 ( .A1(n17223), .A2(n17224), .ZN(n17065) );
  NAND2_X1 U17126 ( .A1(n17062), .A2(n17225), .ZN(n17224) );
  NAND2_X1 U17127 ( .A1(n17060), .A2(n17061), .ZN(n17225) );
  NOR2_X1 U17128 ( .A1(n10084), .A2(n10054), .ZN(n17062) );
  NAND2_X1 U17129 ( .A1(n17226), .A2(n17227), .ZN(n17223) );
  INV_X1 U17130 ( .A(n17061), .ZN(n17227) );
  NOR2_X1 U17131 ( .A1(n17228), .A2(n17229), .ZN(n17061) );
  INV_X1 U17132 ( .A(n17230), .ZN(n17229) );
  NAND2_X1 U17133 ( .A1(n17058), .A2(n17231), .ZN(n17230) );
  NAND2_X1 U17134 ( .A1(n17057), .A2(n17056), .ZN(n17231) );
  NOR2_X1 U17135 ( .A1(n10084), .A2(n9358), .ZN(n17058) );
  NOR2_X1 U17136 ( .A1(n17056), .A2(n17057), .ZN(n17228) );
  NOR2_X1 U17137 ( .A1(n17232), .A2(n17233), .ZN(n17057) );
  INV_X1 U17138 ( .A(n17234), .ZN(n17233) );
  NAND2_X1 U17139 ( .A1(n17054), .A2(n17235), .ZN(n17234) );
  NAND2_X1 U17140 ( .A1(n17053), .A2(n17052), .ZN(n17235) );
  NOR2_X1 U17141 ( .A1(n10084), .A2(n9330), .ZN(n17054) );
  NOR2_X1 U17142 ( .A1(n17052), .A2(n17053), .ZN(n17232) );
  INV_X1 U17143 ( .A(n17236), .ZN(n17053) );
  NAND2_X1 U17144 ( .A1(n17237), .A2(n17238), .ZN(n17236) );
  NAND2_X1 U17145 ( .A1(n17050), .A2(n17239), .ZN(n17238) );
  NAND2_X1 U17146 ( .A1(n17240), .A2(n17049), .ZN(n17239) );
  INV_X1 U17147 ( .A(n17048), .ZN(n17240) );
  NOR2_X1 U17148 ( .A1(n10084), .A2(n10051), .ZN(n17050) );
  NAND2_X1 U17149 ( .A1(n17048), .A2(n17241), .ZN(n17237) );
  INV_X1 U17150 ( .A(n17049), .ZN(n17241) );
  NOR2_X1 U17151 ( .A1(n17242), .A2(n17243), .ZN(n17049) );
  NOR2_X1 U17152 ( .A1(n17046), .A2(n17244), .ZN(n17243) );
  NOR2_X1 U17153 ( .A1(n17043), .A2(n17045), .ZN(n17244) );
  NAND2_X1 U17154 ( .A1(b_4_), .A2(a_24_), .ZN(n17046) );
  INV_X1 U17155 ( .A(n17245), .ZN(n17242) );
  NAND2_X1 U17156 ( .A1(n17043), .A2(n17045), .ZN(n17245) );
  NAND2_X1 U17157 ( .A1(n17246), .A2(n17247), .ZN(n17045) );
  NAND2_X1 U17158 ( .A1(n17042), .A2(n17248), .ZN(n17247) );
  NAND2_X1 U17159 ( .A1(n17039), .A2(n17041), .ZN(n17248) );
  NOR2_X1 U17160 ( .A1(n10084), .A2(n10048), .ZN(n17042) );
  INV_X1 U17161 ( .A(n17249), .ZN(n17246) );
  NOR2_X1 U17162 ( .A1(n17041), .A2(n17039), .ZN(n17249) );
  XNOR2_X1 U17163 ( .A(n17250), .B(n17251), .ZN(n17039) );
  XNOR2_X1 U17164 ( .A(n17252), .B(n17253), .ZN(n17251) );
  NAND2_X1 U17165 ( .A1(n17254), .A2(n17255), .ZN(n17041) );
  NAND2_X1 U17166 ( .A1(n16999), .A2(n17256), .ZN(n17255) );
  NAND2_X1 U17167 ( .A1(n17002), .A2(n17001), .ZN(n17256) );
  XOR2_X1 U17168 ( .A(n17257), .B(n17258), .Z(n16999) );
  NAND2_X1 U17169 ( .A1(n17259), .A2(n17260), .ZN(n17257) );
  INV_X1 U17170 ( .A(n17261), .ZN(n17254) );
  NOR2_X1 U17171 ( .A1(n17001), .A2(n17002), .ZN(n17261) );
  NOR2_X1 U17172 ( .A1(n10084), .A2(n10047), .ZN(n17002) );
  NAND2_X1 U17173 ( .A1(n17008), .A2(n17262), .ZN(n17001) );
  NAND2_X1 U17174 ( .A1(n17007), .A2(n17009), .ZN(n17262) );
  NAND2_X1 U17175 ( .A1(n17263), .A2(n17264), .ZN(n17009) );
  NAND2_X1 U17176 ( .A1(b_4_), .A2(a_27_), .ZN(n17264) );
  INV_X1 U17177 ( .A(n17265), .ZN(n17263) );
  XNOR2_X1 U17178 ( .A(n17266), .B(n17267), .ZN(n17007) );
  XOR2_X1 U17179 ( .A(n17268), .B(n17269), .Z(n17267) );
  NAND2_X1 U17180 ( .A1(b_3_), .A2(a_28_), .ZN(n17269) );
  NAND2_X1 U17181 ( .A1(a_27_), .A2(n17265), .ZN(n17008) );
  NAND2_X1 U17182 ( .A1(n17270), .A2(n17271), .ZN(n17265) );
  NAND2_X1 U17183 ( .A1(n17272), .A2(b_4_), .ZN(n17271) );
  NOR2_X1 U17184 ( .A1(n17273), .A2(n9136), .ZN(n17272) );
  NOR2_X1 U17185 ( .A1(n17015), .A2(n17017), .ZN(n17273) );
  NAND2_X1 U17186 ( .A1(n17015), .A2(n17017), .ZN(n17270) );
  NAND2_X1 U17187 ( .A1(n17274), .A2(n17275), .ZN(n17017) );
  NAND2_X1 U17188 ( .A1(n17276), .A2(b_4_), .ZN(n17275) );
  NOR2_X1 U17189 ( .A1(n17277), .A2(n9121), .ZN(n17276) );
  NOR2_X1 U17190 ( .A1(n17278), .A2(n17037), .ZN(n17277) );
  NAND2_X1 U17191 ( .A1(n17278), .A2(n17037), .ZN(n17274) );
  NAND2_X1 U17192 ( .A1(n17279), .A2(n17280), .ZN(n17037) );
  NAND2_X1 U17193 ( .A1(b_2_), .A2(n17281), .ZN(n17280) );
  NAND2_X1 U17194 ( .A1(n10486), .A2(n17282), .ZN(n17281) );
  NAND2_X1 U17195 ( .A1(a_31_), .A2(n9888), .ZN(n17282) );
  NAND2_X1 U17196 ( .A1(b_3_), .A2(n17283), .ZN(n17279) );
  NAND2_X1 U17197 ( .A1(n10489), .A2(n17284), .ZN(n17283) );
  NAND2_X1 U17198 ( .A1(a_30_), .A2(n10087), .ZN(n17284) );
  INV_X1 U17199 ( .A(n17038), .ZN(n17278) );
  NAND2_X1 U17200 ( .A1(n17285), .A2(n9025), .ZN(n17038) );
  NOR2_X1 U17201 ( .A1(n9888), .A2(n10084), .ZN(n17285) );
  XOR2_X1 U17202 ( .A(n17286), .B(n17287), .Z(n17015) );
  NOR2_X1 U17203 ( .A1(n9121), .A2(n9888), .ZN(n17287) );
  XNOR2_X1 U17204 ( .A(n17288), .B(n17289), .ZN(n17286) );
  XNOR2_X1 U17205 ( .A(n17290), .B(n17291), .ZN(n17043) );
  XNOR2_X1 U17206 ( .A(n17292), .B(n17293), .ZN(n17291) );
  XOR2_X1 U17207 ( .A(n17294), .B(n17295), .Z(n17048) );
  XNOR2_X1 U17208 ( .A(n17296), .B(n17297), .ZN(n17295) );
  XOR2_X1 U17209 ( .A(n17298), .B(n17299), .Z(n17052) );
  NAND2_X1 U17210 ( .A1(n17300), .A2(n17301), .ZN(n17298) );
  XNOR2_X1 U17211 ( .A(n17302), .B(n17303), .ZN(n17056) );
  XOR2_X1 U17212 ( .A(n17304), .B(n17305), .Z(n17302) );
  NOR2_X1 U17213 ( .A1(n9330), .A2(n9888), .ZN(n17305) );
  INV_X1 U17214 ( .A(n17060), .ZN(n17226) );
  XOR2_X1 U17215 ( .A(n17306), .B(n17307), .Z(n17060) );
  NAND2_X1 U17216 ( .A1(n17308), .A2(n17309), .ZN(n17306) );
  XOR2_X1 U17217 ( .A(n17310), .B(n17311), .Z(n17064) );
  XOR2_X1 U17218 ( .A(n17312), .B(n17313), .Z(n17310) );
  NOR2_X1 U17219 ( .A1(n10054), .A2(n9888), .ZN(n17313) );
  XNOR2_X1 U17220 ( .A(n17314), .B(n17315), .ZN(n17067) );
  NAND2_X1 U17221 ( .A1(n17316), .A2(n17317), .ZN(n17314) );
  XOR2_X1 U17222 ( .A(n17318), .B(n17319), .Z(n17072) );
  XOR2_X1 U17223 ( .A(n17320), .B(n17321), .Z(n17318) );
  NOR2_X1 U17224 ( .A1(n10058), .A2(n9888), .ZN(n17321) );
  XNOR2_X1 U17225 ( .A(n17322), .B(n17323), .ZN(n17075) );
  NAND2_X1 U17226 ( .A1(n17324), .A2(n17325), .ZN(n17322) );
  XOR2_X1 U17227 ( .A(n17326), .B(n17327), .Z(n17080) );
  XOR2_X1 U17228 ( .A(n17328), .B(n17329), .Z(n17326) );
  NOR2_X1 U17229 ( .A1(n10062), .A2(n9888), .ZN(n17329) );
  XNOR2_X1 U17230 ( .A(n17330), .B(n17331), .ZN(n17083) );
  NAND2_X1 U17231 ( .A1(n17332), .A2(n17333), .ZN(n17330) );
  XOR2_X1 U17232 ( .A(n17334), .B(n17335), .Z(n17087) );
  XOR2_X1 U17233 ( .A(n17336), .B(n17337), .Z(n17334) );
  NOR2_X1 U17234 ( .A1(n10065), .A2(n9888), .ZN(n17337) );
  XNOR2_X1 U17235 ( .A(n17338), .B(n17339), .ZN(n17091) );
  NAND2_X1 U17236 ( .A1(n17340), .A2(n17341), .ZN(n17338) );
  XOR2_X1 U17237 ( .A(n17342), .B(n17343), .Z(n17096) );
  XOR2_X1 U17238 ( .A(n17344), .B(n17345), .Z(n17342) );
  NOR2_X1 U17239 ( .A1(n10070), .A2(n9888), .ZN(n17345) );
  XNOR2_X1 U17240 ( .A(n17346), .B(n17347), .ZN(n17099) );
  NAND2_X1 U17241 ( .A1(n17348), .A2(n17349), .ZN(n17346) );
  XOR2_X1 U17242 ( .A(n17350), .B(n17351), .Z(n17104) );
  XOR2_X1 U17243 ( .A(n17352), .B(n17353), .Z(n17350) );
  NOR2_X1 U17244 ( .A1(n10073), .A2(n9888), .ZN(n17353) );
  XNOR2_X1 U17245 ( .A(n17354), .B(n17355), .ZN(n17107) );
  NAND2_X1 U17246 ( .A1(n17356), .A2(n17357), .ZN(n17354) );
  XOR2_X1 U17247 ( .A(n17358), .B(n17359), .Z(n17112) );
  XOR2_X1 U17248 ( .A(n17360), .B(n17361), .Z(n17358) );
  NOR2_X1 U17249 ( .A1(n10079), .A2(n9888), .ZN(n17361) );
  XNOR2_X1 U17250 ( .A(n17362), .B(n17363), .ZN(n16914) );
  NAND2_X1 U17251 ( .A1(n17364), .A2(n17365), .ZN(n17362) );
  XNOR2_X1 U17252 ( .A(n17366), .B(n17367), .ZN(n17116) );
  XOR2_X1 U17253 ( .A(n17368), .B(n17369), .Z(n17366) );
  NOR2_X1 U17254 ( .A1(n10081), .A2(n9888), .ZN(n17369) );
  XNOR2_X1 U17255 ( .A(n17370), .B(n17371), .ZN(n17122) );
  XOR2_X1 U17256 ( .A(n17372), .B(n17373), .Z(n17370) );
  NOR2_X1 U17257 ( .A1(n10085), .A2(n9888), .ZN(n17373) );
  INV_X1 U17258 ( .A(n17149), .ZN(n17126) );
  XOR2_X1 U17259 ( .A(n17374), .B(n17375), .Z(n17149) );
  XNOR2_X1 U17260 ( .A(n17376), .B(n9985), .ZN(n17374) );
  INV_X1 U17261 ( .A(n17377), .ZN(n9985) );
  XOR2_X1 U17262 ( .A(n17378), .B(n17379), .Z(n17130) );
  XNOR2_X1 U17263 ( .A(n17380), .B(n17381), .ZN(n17379) );
  NAND2_X1 U17264 ( .A1(a_2_), .A2(b_3_), .ZN(n17381) );
  XNOR2_X1 U17265 ( .A(n17382), .B(n17383), .ZN(n16887) );
  NAND2_X1 U17266 ( .A1(n17384), .A2(n17385), .ZN(n17382) );
  XNOR2_X1 U17267 ( .A(n17386), .B(n17387), .ZN(n17135) );
  XOR2_X1 U17268 ( .A(n17388), .B(n17389), .Z(n17386) );
  NOR2_X1 U17269 ( .A1(n9888), .A2(n10093), .ZN(n17389) );
  NOR2_X1 U17270 ( .A1(n17390), .A2(n10252), .ZN(n9751) );
  INV_X1 U17271 ( .A(n17391), .ZN(n10252) );
  NAND2_X1 U17272 ( .A1(n17392), .A2(n17393), .ZN(n17391) );
  NOR2_X1 U17273 ( .A1(n17392), .A2(n17393), .ZN(n17390) );
  NAND2_X1 U17274 ( .A1(n17394), .A2(n17395), .ZN(n17393) );
  NAND2_X1 U17275 ( .A1(n17396), .A2(a_0_), .ZN(n17395) );
  NOR2_X1 U17276 ( .A1(n17397), .A2(n9888), .ZN(n17396) );
  NOR2_X1 U17277 ( .A1(n17388), .A2(n17387), .ZN(n17397) );
  NAND2_X1 U17278 ( .A1(n17387), .A2(n17388), .ZN(n17394) );
  NAND2_X1 U17279 ( .A1(n17384), .A2(n17398), .ZN(n17388) );
  NAND2_X1 U17280 ( .A1(n17383), .A2(n17385), .ZN(n17398) );
  NAND2_X1 U17281 ( .A1(n17399), .A2(n17400), .ZN(n17385) );
  NAND2_X1 U17282 ( .A1(a_1_), .A2(b_3_), .ZN(n17400) );
  INV_X1 U17283 ( .A(n17401), .ZN(n17399) );
  XNOR2_X1 U17284 ( .A(n17402), .B(n17403), .ZN(n17383) );
  XOR2_X1 U17285 ( .A(n17404), .B(n9923), .Z(n17402) );
  NAND2_X1 U17286 ( .A1(a_1_), .A2(n17401), .ZN(n17384) );
  NAND2_X1 U17287 ( .A1(n17405), .A2(n17406), .ZN(n17401) );
  NAND2_X1 U17288 ( .A1(n17407), .A2(a_2_), .ZN(n17406) );
  NOR2_X1 U17289 ( .A1(n17408), .A2(n9888), .ZN(n17407) );
  NOR2_X1 U17290 ( .A1(n17380), .A2(n17378), .ZN(n17408) );
  NAND2_X1 U17291 ( .A1(n17380), .A2(n17378), .ZN(n17405) );
  XNOR2_X1 U17292 ( .A(n17409), .B(n17410), .ZN(n17378) );
  XNOR2_X1 U17293 ( .A(n17411), .B(n17412), .ZN(n17409) );
  NOR2_X1 U17294 ( .A1(n17413), .A2(n17414), .ZN(n17380) );
  INV_X1 U17295 ( .A(n17415), .ZN(n17414) );
  NAND2_X1 U17296 ( .A1(n17375), .A2(n17416), .ZN(n17415) );
  NAND2_X1 U17297 ( .A1(n17377), .A2(n17376), .ZN(n17416) );
  XOR2_X1 U17298 ( .A(n17417), .B(n17418), .Z(n17375) );
  XNOR2_X1 U17299 ( .A(n17419), .B(n17420), .ZN(n17417) );
  NOR2_X1 U17300 ( .A1(n17376), .A2(n17377), .ZN(n17413) );
  NOR2_X1 U17301 ( .A1(n9888), .A2(n10086), .ZN(n17377) );
  NAND2_X1 U17302 ( .A1(n17421), .A2(n17422), .ZN(n17376) );
  NAND2_X1 U17303 ( .A1(n17423), .A2(b_3_), .ZN(n17422) );
  NOR2_X1 U17304 ( .A1(n17424), .A2(n10085), .ZN(n17423) );
  NOR2_X1 U17305 ( .A1(n17372), .A2(n17371), .ZN(n17424) );
  NAND2_X1 U17306 ( .A1(n17371), .A2(n17372), .ZN(n17421) );
  NAND2_X1 U17307 ( .A1(n17160), .A2(n17425), .ZN(n17372) );
  NAND2_X1 U17308 ( .A1(n17159), .A2(n17161), .ZN(n17425) );
  NAND2_X1 U17309 ( .A1(n17426), .A2(n17427), .ZN(n17161) );
  NAND2_X1 U17310 ( .A1(b_3_), .A2(a_5_), .ZN(n17427) );
  INV_X1 U17311 ( .A(n17428), .ZN(n17426) );
  XNOR2_X1 U17312 ( .A(n17429), .B(n17430), .ZN(n17159) );
  XNOR2_X1 U17313 ( .A(n17431), .B(n17432), .ZN(n17429) );
  NAND2_X1 U17314 ( .A1(a_5_), .A2(n17428), .ZN(n17160) );
  NAND2_X1 U17315 ( .A1(n17433), .A2(n17434), .ZN(n17428) );
  NAND2_X1 U17316 ( .A1(n17435), .A2(b_3_), .ZN(n17434) );
  NOR2_X1 U17317 ( .A1(n17436), .A2(n10081), .ZN(n17435) );
  NOR2_X1 U17318 ( .A1(n17368), .A2(n17367), .ZN(n17436) );
  NAND2_X1 U17319 ( .A1(n17367), .A2(n17368), .ZN(n17433) );
  NAND2_X1 U17320 ( .A1(n17364), .A2(n17437), .ZN(n17368) );
  NAND2_X1 U17321 ( .A1(n17363), .A2(n17365), .ZN(n17437) );
  NAND2_X1 U17322 ( .A1(n17438), .A2(n17439), .ZN(n17365) );
  NAND2_X1 U17323 ( .A1(b_3_), .A2(a_7_), .ZN(n17439) );
  INV_X1 U17324 ( .A(n17440), .ZN(n17438) );
  XNOR2_X1 U17325 ( .A(n17441), .B(n17442), .ZN(n17363) );
  XNOR2_X1 U17326 ( .A(n17443), .B(n17444), .ZN(n17441) );
  NAND2_X1 U17327 ( .A1(a_7_), .A2(n17440), .ZN(n17364) );
  NAND2_X1 U17328 ( .A1(n17445), .A2(n17446), .ZN(n17440) );
  NAND2_X1 U17329 ( .A1(n17447), .A2(b_3_), .ZN(n17446) );
  NOR2_X1 U17330 ( .A1(n17448), .A2(n10079), .ZN(n17447) );
  NOR2_X1 U17331 ( .A1(n17360), .A2(n17359), .ZN(n17448) );
  NAND2_X1 U17332 ( .A1(n17359), .A2(n17360), .ZN(n17445) );
  NAND2_X1 U17333 ( .A1(n17356), .A2(n17449), .ZN(n17360) );
  NAND2_X1 U17334 ( .A1(n17355), .A2(n17357), .ZN(n17449) );
  NAND2_X1 U17335 ( .A1(n17450), .A2(n17451), .ZN(n17357) );
  NAND2_X1 U17336 ( .A1(b_3_), .A2(a_9_), .ZN(n17451) );
  INV_X1 U17337 ( .A(n17452), .ZN(n17450) );
  XNOR2_X1 U17338 ( .A(n17453), .B(n17454), .ZN(n17355) );
  XNOR2_X1 U17339 ( .A(n17455), .B(n17456), .ZN(n17453) );
  NAND2_X1 U17340 ( .A1(a_9_), .A2(n17452), .ZN(n17356) );
  NAND2_X1 U17341 ( .A1(n17457), .A2(n17458), .ZN(n17452) );
  NAND2_X1 U17342 ( .A1(n17459), .A2(b_3_), .ZN(n17458) );
  NOR2_X1 U17343 ( .A1(n17460), .A2(n10073), .ZN(n17459) );
  NOR2_X1 U17344 ( .A1(n17352), .A2(n17351), .ZN(n17460) );
  NAND2_X1 U17345 ( .A1(n17351), .A2(n17352), .ZN(n17457) );
  NAND2_X1 U17346 ( .A1(n17348), .A2(n17461), .ZN(n17352) );
  NAND2_X1 U17347 ( .A1(n17347), .A2(n17349), .ZN(n17461) );
  NAND2_X1 U17348 ( .A1(n17462), .A2(n17463), .ZN(n17349) );
  NAND2_X1 U17349 ( .A1(b_3_), .A2(a_11_), .ZN(n17463) );
  INV_X1 U17350 ( .A(n17464), .ZN(n17462) );
  XNOR2_X1 U17351 ( .A(n17465), .B(n17466), .ZN(n17347) );
  XNOR2_X1 U17352 ( .A(n17467), .B(n17468), .ZN(n17465) );
  NAND2_X1 U17353 ( .A1(a_11_), .A2(n17464), .ZN(n17348) );
  NAND2_X1 U17354 ( .A1(n17469), .A2(n17470), .ZN(n17464) );
  NAND2_X1 U17355 ( .A1(n17471), .A2(b_3_), .ZN(n17470) );
  NOR2_X1 U17356 ( .A1(n17472), .A2(n10070), .ZN(n17471) );
  NOR2_X1 U17357 ( .A1(n17344), .A2(n17343), .ZN(n17472) );
  NAND2_X1 U17358 ( .A1(n17343), .A2(n17344), .ZN(n17469) );
  NAND2_X1 U17359 ( .A1(n17340), .A2(n17473), .ZN(n17344) );
  NAND2_X1 U17360 ( .A1(n17339), .A2(n17341), .ZN(n17473) );
  NAND2_X1 U17361 ( .A1(n17474), .A2(n17475), .ZN(n17341) );
  NAND2_X1 U17362 ( .A1(b_3_), .A2(a_13_), .ZN(n17475) );
  INV_X1 U17363 ( .A(n17476), .ZN(n17474) );
  XNOR2_X1 U17364 ( .A(n17477), .B(n17478), .ZN(n17339) );
  XNOR2_X1 U17365 ( .A(n17479), .B(n17480), .ZN(n17477) );
  NAND2_X1 U17366 ( .A1(a_13_), .A2(n17476), .ZN(n17340) );
  NAND2_X1 U17367 ( .A1(n17481), .A2(n17482), .ZN(n17476) );
  NAND2_X1 U17368 ( .A1(n17483), .A2(b_3_), .ZN(n17482) );
  NOR2_X1 U17369 ( .A1(n17484), .A2(n10065), .ZN(n17483) );
  NOR2_X1 U17370 ( .A1(n17336), .A2(n17335), .ZN(n17484) );
  NAND2_X1 U17371 ( .A1(n17335), .A2(n17336), .ZN(n17481) );
  NAND2_X1 U17372 ( .A1(n17332), .A2(n17485), .ZN(n17336) );
  NAND2_X1 U17373 ( .A1(n17331), .A2(n17333), .ZN(n17485) );
  NAND2_X1 U17374 ( .A1(n17486), .A2(n17487), .ZN(n17333) );
  NAND2_X1 U17375 ( .A1(b_3_), .A2(a_15_), .ZN(n17487) );
  INV_X1 U17376 ( .A(n17488), .ZN(n17486) );
  XNOR2_X1 U17377 ( .A(n17489), .B(n17490), .ZN(n17331) );
  XNOR2_X1 U17378 ( .A(n17491), .B(n17492), .ZN(n17489) );
  NAND2_X1 U17379 ( .A1(a_15_), .A2(n17488), .ZN(n17332) );
  NAND2_X1 U17380 ( .A1(n17493), .A2(n17494), .ZN(n17488) );
  NAND2_X1 U17381 ( .A1(n17495), .A2(b_3_), .ZN(n17494) );
  NOR2_X1 U17382 ( .A1(n17496), .A2(n10062), .ZN(n17495) );
  NOR2_X1 U17383 ( .A1(n17328), .A2(n17327), .ZN(n17496) );
  NAND2_X1 U17384 ( .A1(n17327), .A2(n17328), .ZN(n17493) );
  NAND2_X1 U17385 ( .A1(n17324), .A2(n17497), .ZN(n17328) );
  NAND2_X1 U17386 ( .A1(n17323), .A2(n17325), .ZN(n17497) );
  NAND2_X1 U17387 ( .A1(n17498), .A2(n17499), .ZN(n17325) );
  NAND2_X1 U17388 ( .A1(b_3_), .A2(a_17_), .ZN(n17499) );
  INV_X1 U17389 ( .A(n17500), .ZN(n17498) );
  XNOR2_X1 U17390 ( .A(n17501), .B(n17502), .ZN(n17323) );
  XNOR2_X1 U17391 ( .A(n17503), .B(n17504), .ZN(n17501) );
  NAND2_X1 U17392 ( .A1(a_17_), .A2(n17500), .ZN(n17324) );
  NAND2_X1 U17393 ( .A1(n17505), .A2(n17506), .ZN(n17500) );
  NAND2_X1 U17394 ( .A1(n17507), .A2(b_3_), .ZN(n17506) );
  NOR2_X1 U17395 ( .A1(n17508), .A2(n10058), .ZN(n17507) );
  NOR2_X1 U17396 ( .A1(n17320), .A2(n17319), .ZN(n17508) );
  NAND2_X1 U17397 ( .A1(n17319), .A2(n17320), .ZN(n17505) );
  NAND2_X1 U17398 ( .A1(n17316), .A2(n17509), .ZN(n17320) );
  NAND2_X1 U17399 ( .A1(n17315), .A2(n17317), .ZN(n17509) );
  NAND2_X1 U17400 ( .A1(n17510), .A2(n17511), .ZN(n17317) );
  NAND2_X1 U17401 ( .A1(b_3_), .A2(a_19_), .ZN(n17511) );
  INV_X1 U17402 ( .A(n17512), .ZN(n17510) );
  XNOR2_X1 U17403 ( .A(n17513), .B(n17514), .ZN(n17315) );
  XNOR2_X1 U17404 ( .A(n17515), .B(n17516), .ZN(n17513) );
  NAND2_X1 U17405 ( .A1(a_19_), .A2(n17512), .ZN(n17316) );
  NAND2_X1 U17406 ( .A1(n17517), .A2(n17518), .ZN(n17512) );
  NAND2_X1 U17407 ( .A1(n17519), .A2(b_3_), .ZN(n17518) );
  NOR2_X1 U17408 ( .A1(n17520), .A2(n10054), .ZN(n17519) );
  NOR2_X1 U17409 ( .A1(n17312), .A2(n17311), .ZN(n17520) );
  NAND2_X1 U17410 ( .A1(n17311), .A2(n17312), .ZN(n17517) );
  NAND2_X1 U17411 ( .A1(n17308), .A2(n17521), .ZN(n17312) );
  NAND2_X1 U17412 ( .A1(n17307), .A2(n17309), .ZN(n17521) );
  NAND2_X1 U17413 ( .A1(n17522), .A2(n17523), .ZN(n17309) );
  NAND2_X1 U17414 ( .A1(b_3_), .A2(a_21_), .ZN(n17523) );
  INV_X1 U17415 ( .A(n17524), .ZN(n17522) );
  XNOR2_X1 U17416 ( .A(n17525), .B(n17526), .ZN(n17307) );
  XNOR2_X1 U17417 ( .A(n17527), .B(n17528), .ZN(n17525) );
  NAND2_X1 U17418 ( .A1(a_21_), .A2(n17524), .ZN(n17308) );
  NAND2_X1 U17419 ( .A1(n17529), .A2(n17530), .ZN(n17524) );
  NAND2_X1 U17420 ( .A1(n17531), .A2(b_3_), .ZN(n17530) );
  NOR2_X1 U17421 ( .A1(n17532), .A2(n9330), .ZN(n17531) );
  NOR2_X1 U17422 ( .A1(n17304), .A2(n17303), .ZN(n17532) );
  NAND2_X1 U17423 ( .A1(n17303), .A2(n17304), .ZN(n17529) );
  NAND2_X1 U17424 ( .A1(n17300), .A2(n17533), .ZN(n17304) );
  NAND2_X1 U17425 ( .A1(n17299), .A2(n17301), .ZN(n17533) );
  NAND2_X1 U17426 ( .A1(n17534), .A2(n17535), .ZN(n17301) );
  NAND2_X1 U17427 ( .A1(b_3_), .A2(a_23_), .ZN(n17535) );
  XNOR2_X1 U17428 ( .A(n17536), .B(n17537), .ZN(n17299) );
  NAND2_X1 U17429 ( .A1(n17538), .A2(n17539), .ZN(n17536) );
  INV_X1 U17430 ( .A(n17540), .ZN(n17300) );
  NOR2_X1 U17431 ( .A1(n10051), .A2(n17534), .ZN(n17540) );
  NOR2_X1 U17432 ( .A1(n17541), .A2(n17542), .ZN(n17534) );
  NOR2_X1 U17433 ( .A1(n17297), .A2(n17543), .ZN(n17542) );
  NOR2_X1 U17434 ( .A1(n17544), .A2(n17545), .ZN(n17543) );
  INV_X1 U17435 ( .A(n17294), .ZN(n17545) );
  INV_X1 U17436 ( .A(n17296), .ZN(n17544) );
  NAND2_X1 U17437 ( .A1(b_3_), .A2(a_24_), .ZN(n17297) );
  NOR2_X1 U17438 ( .A1(n17294), .A2(n17296), .ZN(n17541) );
  NOR2_X1 U17439 ( .A1(n17546), .A2(n17547), .ZN(n17296) );
  INV_X1 U17440 ( .A(n17548), .ZN(n17547) );
  NAND2_X1 U17441 ( .A1(n17293), .A2(n17549), .ZN(n17548) );
  NAND2_X1 U17442 ( .A1(n17290), .A2(n17292), .ZN(n17549) );
  NOR2_X1 U17443 ( .A1(n9888), .A2(n10048), .ZN(n17293) );
  NOR2_X1 U17444 ( .A1(n17292), .A2(n17290), .ZN(n17546) );
  XOR2_X1 U17445 ( .A(n17550), .B(n17551), .Z(n17290) );
  XNOR2_X1 U17446 ( .A(n17552), .B(n17553), .ZN(n17551) );
  NOR2_X1 U17447 ( .A1(n10047), .A2(n10087), .ZN(n17553) );
  NAND2_X1 U17448 ( .A1(n17554), .A2(n17555), .ZN(n17292) );
  NAND2_X1 U17449 ( .A1(n17250), .A2(n17556), .ZN(n17555) );
  NAND2_X1 U17450 ( .A1(n17253), .A2(n17252), .ZN(n17556) );
  XOR2_X1 U17451 ( .A(n17557), .B(n17558), .Z(n17250) );
  NAND2_X1 U17452 ( .A1(n17559), .A2(n17560), .ZN(n17557) );
  INV_X1 U17453 ( .A(n17561), .ZN(n17554) );
  NOR2_X1 U17454 ( .A1(n17252), .A2(n17253), .ZN(n17561) );
  NOR2_X1 U17455 ( .A1(n9888), .A2(n10047), .ZN(n17253) );
  NAND2_X1 U17456 ( .A1(n17259), .A2(n17562), .ZN(n17252) );
  NAND2_X1 U17457 ( .A1(n17258), .A2(n17260), .ZN(n17562) );
  NAND2_X1 U17458 ( .A1(n17563), .A2(n17564), .ZN(n17260) );
  NAND2_X1 U17459 ( .A1(b_3_), .A2(a_27_), .ZN(n17564) );
  INV_X1 U17460 ( .A(n17565), .ZN(n17563) );
  XNOR2_X1 U17461 ( .A(n17566), .B(n17567), .ZN(n17258) );
  XOR2_X1 U17462 ( .A(n17568), .B(n17569), .Z(n17567) );
  NAND2_X1 U17463 ( .A1(b_2_), .A2(a_28_), .ZN(n17569) );
  NAND2_X1 U17464 ( .A1(a_27_), .A2(n17565), .ZN(n17259) );
  NAND2_X1 U17465 ( .A1(n17570), .A2(n17571), .ZN(n17565) );
  NAND2_X1 U17466 ( .A1(n17572), .A2(b_3_), .ZN(n17571) );
  NOR2_X1 U17467 ( .A1(n17573), .A2(n9136), .ZN(n17572) );
  NOR2_X1 U17468 ( .A1(n17266), .A2(n17268), .ZN(n17573) );
  NAND2_X1 U17469 ( .A1(n17266), .A2(n17268), .ZN(n17570) );
  NAND2_X1 U17470 ( .A1(n17574), .A2(n17575), .ZN(n17268) );
  NAND2_X1 U17471 ( .A1(n17576), .A2(b_3_), .ZN(n17575) );
  NOR2_X1 U17472 ( .A1(n17577), .A2(n9121), .ZN(n17576) );
  NOR2_X1 U17473 ( .A1(n17578), .A2(n17288), .ZN(n17577) );
  NAND2_X1 U17474 ( .A1(n17578), .A2(n17288), .ZN(n17574) );
  NAND2_X1 U17475 ( .A1(n17579), .A2(n17580), .ZN(n17288) );
  NAND2_X1 U17476 ( .A1(b_1_), .A2(n17581), .ZN(n17580) );
  NAND2_X1 U17477 ( .A1(n10486), .A2(n17582), .ZN(n17581) );
  NAND2_X1 U17478 ( .A1(a_31_), .A2(n10087), .ZN(n17582) );
  NAND2_X1 U17479 ( .A1(b_2_), .A2(n17583), .ZN(n17579) );
  NAND2_X1 U17480 ( .A1(n10489), .A2(n17584), .ZN(n17583) );
  NAND2_X1 U17481 ( .A1(a_30_), .A2(n9982), .ZN(n17584) );
  INV_X1 U17482 ( .A(n17289), .ZN(n17578) );
  NAND2_X1 U17483 ( .A1(n17585), .A2(n9025), .ZN(n17289) );
  NOR2_X1 U17484 ( .A1(n9888), .A2(n10087), .ZN(n17585) );
  XOR2_X1 U17485 ( .A(n17586), .B(n17587), .Z(n17266) );
  NOR2_X1 U17486 ( .A1(n9121), .A2(n10087), .ZN(n17587) );
  XNOR2_X1 U17487 ( .A(n17588), .B(n17589), .ZN(n17586) );
  XOR2_X1 U17488 ( .A(n17590), .B(n17591), .Z(n17294) );
  NAND2_X1 U17489 ( .A1(n17592), .A2(n17593), .ZN(n17590) );
  XNOR2_X1 U17490 ( .A(n17594), .B(n17595), .ZN(n17303) );
  XNOR2_X1 U17491 ( .A(n17596), .B(n17597), .ZN(n17594) );
  XNOR2_X1 U17492 ( .A(n17598), .B(n17599), .ZN(n17311) );
  XNOR2_X1 U17493 ( .A(n17600), .B(n17601), .ZN(n17598) );
  XNOR2_X1 U17494 ( .A(n17602), .B(n17603), .ZN(n17319) );
  XNOR2_X1 U17495 ( .A(n17604), .B(n17605), .ZN(n17602) );
  XNOR2_X1 U17496 ( .A(n17606), .B(n17607), .ZN(n17327) );
  XNOR2_X1 U17497 ( .A(n17608), .B(n17609), .ZN(n17606) );
  XNOR2_X1 U17498 ( .A(n17610), .B(n17611), .ZN(n17335) );
  XNOR2_X1 U17499 ( .A(n17612), .B(n17613), .ZN(n17610) );
  XNOR2_X1 U17500 ( .A(n17614), .B(n17615), .ZN(n17343) );
  XNOR2_X1 U17501 ( .A(n17616), .B(n17617), .ZN(n17614) );
  XNOR2_X1 U17502 ( .A(n17618), .B(n17619), .ZN(n17351) );
  XNOR2_X1 U17503 ( .A(n17620), .B(n17621), .ZN(n17618) );
  XNOR2_X1 U17504 ( .A(n17622), .B(n17623), .ZN(n17359) );
  XNOR2_X1 U17505 ( .A(n17624), .B(n17625), .ZN(n17622) );
  XNOR2_X1 U17506 ( .A(n17626), .B(n17627), .ZN(n17367) );
  XNOR2_X1 U17507 ( .A(n17628), .B(n17629), .ZN(n17626) );
  XNOR2_X1 U17508 ( .A(n17630), .B(n17631), .ZN(n17371) );
  XNOR2_X1 U17509 ( .A(n17632), .B(n17633), .ZN(n17630) );
  XNOR2_X1 U17510 ( .A(n17634), .B(n17635), .ZN(n17387) );
  XNOR2_X1 U17511 ( .A(n17636), .B(n17637), .ZN(n17634) );
  XNOR2_X1 U17512 ( .A(n17638), .B(n17639), .ZN(n17392) );
  XNOR2_X1 U17513 ( .A(n17640), .B(n17641), .ZN(n17639) );
  XNOR2_X1 U17514 ( .A(n17642), .B(n17643), .ZN(n10108) );
  NOR2_X1 U17515 ( .A1(n17644), .A2(n17645), .ZN(n10176) );
  INV_X1 U17516 ( .A(n17646), .ZN(n17645) );
  XNOR2_X1 U17517 ( .A(n10248), .B(n10091), .ZN(n17644) );
  NOR2_X1 U17518 ( .A1(n17647), .A2(n17646), .ZN(n10177) );
  NAND2_X1 U17519 ( .A1(n17643), .A2(n17642), .ZN(n17646) );
  NAND2_X1 U17520 ( .A1(n17648), .A2(n17649), .ZN(n17642) );
  NAND2_X1 U17521 ( .A1(n17641), .A2(n17650), .ZN(n17649) );
  INV_X1 U17522 ( .A(n17651), .ZN(n17650) );
  NOR2_X1 U17523 ( .A1(n17640), .A2(n17638), .ZN(n17651) );
  NOR2_X1 U17524 ( .A1(n10087), .A2(n10093), .ZN(n17641) );
  NAND2_X1 U17525 ( .A1(n17638), .A2(n17640), .ZN(n17648) );
  NAND2_X1 U17526 ( .A1(n17652), .A2(n17653), .ZN(n17640) );
  NAND2_X1 U17527 ( .A1(n17637), .A2(n17654), .ZN(n17653) );
  NAND2_X1 U17528 ( .A1(n17636), .A2(n17635), .ZN(n17654) );
  NOR2_X1 U17529 ( .A1(n10087), .A2(n9983), .ZN(n17637) );
  INV_X1 U17530 ( .A(n17655), .ZN(n17652) );
  NOR2_X1 U17531 ( .A1(n17635), .A2(n17636), .ZN(n17655) );
  NOR2_X1 U17532 ( .A1(n17656), .A2(n17657), .ZN(n17636) );
  NOR2_X1 U17533 ( .A1(n9923), .A2(n17658), .ZN(n17657) );
  INV_X1 U17534 ( .A(n17659), .ZN(n17658) );
  NAND2_X1 U17535 ( .A1(n17404), .A2(n17403), .ZN(n17659) );
  NAND2_X1 U17536 ( .A1(b_2_), .A2(a_2_), .ZN(n9923) );
  NOR2_X1 U17537 ( .A1(n17403), .A2(n17404), .ZN(n17656) );
  NOR2_X1 U17538 ( .A1(n17660), .A2(n17661), .ZN(n17404) );
  INV_X1 U17539 ( .A(n17662), .ZN(n17661) );
  NAND2_X1 U17540 ( .A1(n17412), .A2(n17663), .ZN(n17662) );
  NAND2_X1 U17541 ( .A1(n17411), .A2(n17410), .ZN(n17663) );
  NOR2_X1 U17542 ( .A1(n10087), .A2(n10086), .ZN(n17412) );
  NOR2_X1 U17543 ( .A1(n17410), .A2(n17411), .ZN(n17660) );
  NOR2_X1 U17544 ( .A1(n17664), .A2(n17665), .ZN(n17411) );
  INV_X1 U17545 ( .A(n17666), .ZN(n17665) );
  NAND2_X1 U17546 ( .A1(n17420), .A2(n17667), .ZN(n17666) );
  NAND2_X1 U17547 ( .A1(n17419), .A2(n17418), .ZN(n17667) );
  NOR2_X1 U17548 ( .A1(n10087), .A2(n10085), .ZN(n17420) );
  NOR2_X1 U17549 ( .A1(n17418), .A2(n17419), .ZN(n17664) );
  NOR2_X1 U17550 ( .A1(n17668), .A2(n17669), .ZN(n17419) );
  INV_X1 U17551 ( .A(n17670), .ZN(n17669) );
  NAND2_X1 U17552 ( .A1(n17633), .A2(n17671), .ZN(n17670) );
  NAND2_X1 U17553 ( .A1(n17632), .A2(n17631), .ZN(n17671) );
  NOR2_X1 U17554 ( .A1(n10087), .A2(n10083), .ZN(n17633) );
  NOR2_X1 U17555 ( .A1(n17631), .A2(n17632), .ZN(n17668) );
  NOR2_X1 U17556 ( .A1(n17672), .A2(n17673), .ZN(n17632) );
  INV_X1 U17557 ( .A(n17674), .ZN(n17673) );
  NAND2_X1 U17558 ( .A1(n17432), .A2(n17675), .ZN(n17674) );
  NAND2_X1 U17559 ( .A1(n17431), .A2(n17430), .ZN(n17675) );
  NOR2_X1 U17560 ( .A1(n10087), .A2(n10081), .ZN(n17432) );
  NOR2_X1 U17561 ( .A1(n17430), .A2(n17431), .ZN(n17672) );
  NOR2_X1 U17562 ( .A1(n17676), .A2(n17677), .ZN(n17431) );
  INV_X1 U17563 ( .A(n17678), .ZN(n17677) );
  NAND2_X1 U17564 ( .A1(n17629), .A2(n17679), .ZN(n17678) );
  NAND2_X1 U17565 ( .A1(n17628), .A2(n17627), .ZN(n17679) );
  NOR2_X1 U17566 ( .A1(n10087), .A2(n9773), .ZN(n17629) );
  NOR2_X1 U17567 ( .A1(n17627), .A2(n17628), .ZN(n17676) );
  NOR2_X1 U17568 ( .A1(n17680), .A2(n17681), .ZN(n17628) );
  INV_X1 U17569 ( .A(n17682), .ZN(n17681) );
  NAND2_X1 U17570 ( .A1(n17444), .A2(n17683), .ZN(n17682) );
  NAND2_X1 U17571 ( .A1(n17443), .A2(n17442), .ZN(n17683) );
  NOR2_X1 U17572 ( .A1(n10087), .A2(n10079), .ZN(n17444) );
  NOR2_X1 U17573 ( .A1(n17442), .A2(n17443), .ZN(n17680) );
  NOR2_X1 U17574 ( .A1(n17684), .A2(n17685), .ZN(n17443) );
  INV_X1 U17575 ( .A(n17686), .ZN(n17685) );
  NAND2_X1 U17576 ( .A1(n17625), .A2(n17687), .ZN(n17686) );
  NAND2_X1 U17577 ( .A1(n17624), .A2(n17623), .ZN(n17687) );
  NOR2_X1 U17578 ( .A1(n10087), .A2(n10076), .ZN(n17625) );
  NOR2_X1 U17579 ( .A1(n17623), .A2(n17624), .ZN(n17684) );
  NOR2_X1 U17580 ( .A1(n17688), .A2(n17689), .ZN(n17624) );
  INV_X1 U17581 ( .A(n17690), .ZN(n17689) );
  NAND2_X1 U17582 ( .A1(n17456), .A2(n17691), .ZN(n17690) );
  NAND2_X1 U17583 ( .A1(n17455), .A2(n17454), .ZN(n17691) );
  NOR2_X1 U17584 ( .A1(n10087), .A2(n10073), .ZN(n17456) );
  NOR2_X1 U17585 ( .A1(n17454), .A2(n17455), .ZN(n17688) );
  NOR2_X1 U17586 ( .A1(n17692), .A2(n17693), .ZN(n17455) );
  INV_X1 U17587 ( .A(n17694), .ZN(n17693) );
  NAND2_X1 U17588 ( .A1(n17621), .A2(n17695), .ZN(n17694) );
  NAND2_X1 U17589 ( .A1(n17620), .A2(n17619), .ZN(n17695) );
  NOR2_X1 U17590 ( .A1(n10087), .A2(n9649), .ZN(n17621) );
  NOR2_X1 U17591 ( .A1(n17619), .A2(n17620), .ZN(n17692) );
  NOR2_X1 U17592 ( .A1(n17696), .A2(n17697), .ZN(n17620) );
  INV_X1 U17593 ( .A(n17698), .ZN(n17697) );
  NAND2_X1 U17594 ( .A1(n17468), .A2(n17699), .ZN(n17698) );
  NAND2_X1 U17595 ( .A1(n17467), .A2(n17466), .ZN(n17699) );
  NOR2_X1 U17596 ( .A1(n10087), .A2(n10070), .ZN(n17468) );
  NOR2_X1 U17597 ( .A1(n17466), .A2(n17467), .ZN(n17696) );
  NOR2_X1 U17598 ( .A1(n17700), .A2(n17701), .ZN(n17467) );
  INV_X1 U17599 ( .A(n17702), .ZN(n17701) );
  NAND2_X1 U17600 ( .A1(n17617), .A2(n17703), .ZN(n17702) );
  NAND2_X1 U17601 ( .A1(n17616), .A2(n17615), .ZN(n17703) );
  NOR2_X1 U17602 ( .A1(n10087), .A2(n10067), .ZN(n17617) );
  NOR2_X1 U17603 ( .A1(n17615), .A2(n17616), .ZN(n17700) );
  NOR2_X1 U17604 ( .A1(n17704), .A2(n17705), .ZN(n17616) );
  INV_X1 U17605 ( .A(n17706), .ZN(n17705) );
  NAND2_X1 U17606 ( .A1(n17480), .A2(n17707), .ZN(n17706) );
  NAND2_X1 U17607 ( .A1(n17479), .A2(n17478), .ZN(n17707) );
  NOR2_X1 U17608 ( .A1(n10087), .A2(n10065), .ZN(n17480) );
  NOR2_X1 U17609 ( .A1(n17478), .A2(n17479), .ZN(n17704) );
  NOR2_X1 U17610 ( .A1(n17708), .A2(n17709), .ZN(n17479) );
  INV_X1 U17611 ( .A(n17710), .ZN(n17709) );
  NAND2_X1 U17612 ( .A1(n17613), .A2(n17711), .ZN(n17710) );
  NAND2_X1 U17613 ( .A1(n17612), .A2(n17611), .ZN(n17711) );
  NOR2_X1 U17614 ( .A1(n10087), .A2(n9534), .ZN(n17613) );
  NOR2_X1 U17615 ( .A1(n17611), .A2(n17612), .ZN(n17708) );
  NOR2_X1 U17616 ( .A1(n17712), .A2(n17713), .ZN(n17612) );
  INV_X1 U17617 ( .A(n17714), .ZN(n17713) );
  NAND2_X1 U17618 ( .A1(n17491), .A2(n17715), .ZN(n17714) );
  NAND2_X1 U17619 ( .A1(n17490), .A2(n17492), .ZN(n17715) );
  NOR2_X1 U17620 ( .A1(n10087), .A2(n10062), .ZN(n17491) );
  NOR2_X1 U17621 ( .A1(n17490), .A2(n17492), .ZN(n17712) );
  NOR2_X1 U17622 ( .A1(n17716), .A2(n17717), .ZN(n17492) );
  INV_X1 U17623 ( .A(n17718), .ZN(n17717) );
  NAND2_X1 U17624 ( .A1(n17609), .A2(n17719), .ZN(n17718) );
  NAND2_X1 U17625 ( .A1(n17608), .A2(n17607), .ZN(n17719) );
  NOR2_X1 U17626 ( .A1(n10087), .A2(n10060), .ZN(n17609) );
  NOR2_X1 U17627 ( .A1(n17607), .A2(n17608), .ZN(n17716) );
  NOR2_X1 U17628 ( .A1(n17720), .A2(n17721), .ZN(n17608) );
  INV_X1 U17629 ( .A(n17722), .ZN(n17721) );
  NAND2_X1 U17630 ( .A1(n17504), .A2(n17723), .ZN(n17722) );
  NAND2_X1 U17631 ( .A1(n17503), .A2(n17502), .ZN(n17723) );
  NOR2_X1 U17632 ( .A1(n10087), .A2(n10058), .ZN(n17504) );
  NOR2_X1 U17633 ( .A1(n17502), .A2(n17503), .ZN(n17720) );
  NOR2_X1 U17634 ( .A1(n17724), .A2(n17725), .ZN(n17503) );
  INV_X1 U17635 ( .A(n17726), .ZN(n17725) );
  NAND2_X1 U17636 ( .A1(n17605), .A2(n17727), .ZN(n17726) );
  NAND2_X1 U17637 ( .A1(n17604), .A2(n17603), .ZN(n17727) );
  NOR2_X1 U17638 ( .A1(n10087), .A2(n9415), .ZN(n17605) );
  NOR2_X1 U17639 ( .A1(n17603), .A2(n17604), .ZN(n17724) );
  NOR2_X1 U17640 ( .A1(n17728), .A2(n17729), .ZN(n17604) );
  INV_X1 U17641 ( .A(n17730), .ZN(n17729) );
  NAND2_X1 U17642 ( .A1(n17516), .A2(n17731), .ZN(n17730) );
  NAND2_X1 U17643 ( .A1(n17515), .A2(n17514), .ZN(n17731) );
  NOR2_X1 U17644 ( .A1(n10087), .A2(n10054), .ZN(n17516) );
  NOR2_X1 U17645 ( .A1(n17514), .A2(n17515), .ZN(n17728) );
  NOR2_X1 U17646 ( .A1(n17732), .A2(n17733), .ZN(n17515) );
  INV_X1 U17647 ( .A(n17734), .ZN(n17733) );
  NAND2_X1 U17648 ( .A1(n17601), .A2(n17735), .ZN(n17734) );
  NAND2_X1 U17649 ( .A1(n17600), .A2(n17599), .ZN(n17735) );
  NOR2_X1 U17650 ( .A1(n10087), .A2(n9358), .ZN(n17601) );
  NOR2_X1 U17651 ( .A1(n17599), .A2(n17600), .ZN(n17732) );
  NOR2_X1 U17652 ( .A1(n17736), .A2(n17737), .ZN(n17600) );
  INV_X1 U17653 ( .A(n17738), .ZN(n17737) );
  NAND2_X1 U17654 ( .A1(n17528), .A2(n17739), .ZN(n17738) );
  NAND2_X1 U17655 ( .A1(n17527), .A2(n17526), .ZN(n17739) );
  NOR2_X1 U17656 ( .A1(n10087), .A2(n9330), .ZN(n17528) );
  NOR2_X1 U17657 ( .A1(n17526), .A2(n17527), .ZN(n17736) );
  NOR2_X1 U17658 ( .A1(n17740), .A2(n17741), .ZN(n17527) );
  INV_X1 U17659 ( .A(n17742), .ZN(n17741) );
  NAND2_X1 U17660 ( .A1(n17597), .A2(n17743), .ZN(n17742) );
  NAND2_X1 U17661 ( .A1(n17596), .A2(n17595), .ZN(n17743) );
  NOR2_X1 U17662 ( .A1(n10087), .A2(n10051), .ZN(n17597) );
  NOR2_X1 U17663 ( .A1(n17595), .A2(n17596), .ZN(n17740) );
  INV_X1 U17664 ( .A(n17744), .ZN(n17596) );
  NAND2_X1 U17665 ( .A1(n17538), .A2(n17745), .ZN(n17744) );
  NAND2_X1 U17666 ( .A1(n17537), .A2(n17539), .ZN(n17745) );
  NAND2_X1 U17667 ( .A1(n17746), .A2(n17747), .ZN(n17539) );
  NAND2_X1 U17668 ( .A1(b_2_), .A2(a_24_), .ZN(n17747) );
  INV_X1 U17669 ( .A(n17748), .ZN(n17746) );
  XOR2_X1 U17670 ( .A(n17749), .B(n17750), .Z(n17537) );
  XNOR2_X1 U17671 ( .A(n17751), .B(n17752), .ZN(n17750) );
  NAND2_X1 U17672 ( .A1(b_1_), .A2(a_25_), .ZN(n17749) );
  NAND2_X1 U17673 ( .A1(a_24_), .A2(n17748), .ZN(n17538) );
  NAND2_X1 U17674 ( .A1(n17592), .A2(n17753), .ZN(n17748) );
  NAND2_X1 U17675 ( .A1(n17591), .A2(n17593), .ZN(n17753) );
  NAND2_X1 U17676 ( .A1(n17754), .A2(n17755), .ZN(n17593) );
  NAND2_X1 U17677 ( .A1(b_2_), .A2(a_25_), .ZN(n17755) );
  INV_X1 U17678 ( .A(n17756), .ZN(n17754) );
  XOR2_X1 U17679 ( .A(n17757), .B(n17758), .Z(n17591) );
  XNOR2_X1 U17680 ( .A(n17759), .B(n17760), .ZN(n17758) );
  NAND2_X1 U17681 ( .A1(b_1_), .A2(a_26_), .ZN(n17757) );
  NAND2_X1 U17682 ( .A1(a_25_), .A2(n17756), .ZN(n17592) );
  NAND2_X1 U17683 ( .A1(n17761), .A2(n17762), .ZN(n17756) );
  NAND2_X1 U17684 ( .A1(n17763), .A2(b_2_), .ZN(n17762) );
  NOR2_X1 U17685 ( .A1(n17764), .A2(n10047), .ZN(n17763) );
  NOR2_X1 U17686 ( .A1(n17550), .A2(n17552), .ZN(n17764) );
  NAND2_X1 U17687 ( .A1(n17550), .A2(n17552), .ZN(n17761) );
  NAND2_X1 U17688 ( .A1(n17559), .A2(n17765), .ZN(n17552) );
  NAND2_X1 U17689 ( .A1(n17558), .A2(n17560), .ZN(n17765) );
  NAND2_X1 U17690 ( .A1(n17766), .A2(n17767), .ZN(n17560) );
  NAND2_X1 U17691 ( .A1(b_2_), .A2(a_27_), .ZN(n17767) );
  INV_X1 U17692 ( .A(n17768), .ZN(n17766) );
  XOR2_X1 U17693 ( .A(n17769), .B(n17770), .Z(n17558) );
  NOR2_X1 U17694 ( .A1(n9136), .A2(n9982), .ZN(n17770) );
  XOR2_X1 U17695 ( .A(n17771), .B(n17772), .Z(n17769) );
  NAND2_X1 U17696 ( .A1(a_27_), .A2(n17768), .ZN(n17559) );
  NAND2_X1 U17697 ( .A1(n17773), .A2(n17774), .ZN(n17768) );
  NAND2_X1 U17698 ( .A1(n17775), .A2(b_2_), .ZN(n17774) );
  NOR2_X1 U17699 ( .A1(n17776), .A2(n9136), .ZN(n17775) );
  NOR2_X1 U17700 ( .A1(n17568), .A2(n17566), .ZN(n17776) );
  NAND2_X1 U17701 ( .A1(n17566), .A2(n17568), .ZN(n17773) );
  NAND2_X1 U17702 ( .A1(n17777), .A2(n17778), .ZN(n17568) );
  NAND2_X1 U17703 ( .A1(n17779), .A2(b_2_), .ZN(n17778) );
  NOR2_X1 U17704 ( .A1(n17780), .A2(n9121), .ZN(n17779) );
  NOR2_X1 U17705 ( .A1(n17781), .A2(n17588), .ZN(n17780) );
  NAND2_X1 U17706 ( .A1(n17781), .A2(n17588), .ZN(n17777) );
  NAND2_X1 U17707 ( .A1(n17782), .A2(n17783), .ZN(n17588) );
  NAND2_X1 U17708 ( .A1(b_0_), .A2(n17784), .ZN(n17783) );
  NAND2_X1 U17709 ( .A1(n10486), .A2(n17785), .ZN(n17784) );
  NAND2_X1 U17710 ( .A1(a_31_), .A2(n9982), .ZN(n17785) );
  NOR2_X1 U17711 ( .A1(n10044), .A2(a_30_), .ZN(n9081) );
  NAND2_X1 U17712 ( .A1(b_1_), .A2(n17786), .ZN(n17782) );
  NAND2_X1 U17713 ( .A1(n10489), .A2(n17787), .ZN(n17786) );
  NAND2_X1 U17714 ( .A1(a_30_), .A2(n10094), .ZN(n17787) );
  INV_X1 U17715 ( .A(n17589), .ZN(n17781) );
  NAND2_X1 U17716 ( .A1(n17788), .A2(n9025), .ZN(n17589) );
  NOR2_X1 U17717 ( .A1(n10087), .A2(n9982), .ZN(n17788) );
  XNOR2_X1 U17718 ( .A(n17789), .B(n17790), .ZN(n17566) );
  XOR2_X1 U17719 ( .A(n17791), .B(n17792), .Z(n17789) );
  XOR2_X1 U17720 ( .A(n17793), .B(n17794), .Z(n17550) );
  XNOR2_X1 U17721 ( .A(n17795), .B(n17796), .ZN(n17794) );
  NAND2_X1 U17722 ( .A1(b_1_), .A2(a_27_), .ZN(n17793) );
  XNOR2_X1 U17723 ( .A(n17797), .B(n17798), .ZN(n17595) );
  XNOR2_X1 U17724 ( .A(n17799), .B(n17800), .ZN(n17798) );
  NAND2_X1 U17725 ( .A1(b_1_), .A2(a_24_), .ZN(n17797) );
  XNOR2_X1 U17726 ( .A(n17801), .B(n17802), .ZN(n17526) );
  XNOR2_X1 U17727 ( .A(n17803), .B(n17804), .ZN(n17802) );
  NAND2_X1 U17728 ( .A1(b_1_), .A2(a_23_), .ZN(n17801) );
  XNOR2_X1 U17729 ( .A(n17805), .B(n17806), .ZN(n17599) );
  XNOR2_X1 U17730 ( .A(n17807), .B(n17808), .ZN(n17806) );
  NAND2_X1 U17731 ( .A1(b_1_), .A2(a_22_), .ZN(n17805) );
  XNOR2_X1 U17732 ( .A(n17809), .B(n17810), .ZN(n17514) );
  XNOR2_X1 U17733 ( .A(n17811), .B(n17812), .ZN(n17810) );
  NAND2_X1 U17734 ( .A1(b_1_), .A2(a_21_), .ZN(n17809) );
  XNOR2_X1 U17735 ( .A(n17813), .B(n17814), .ZN(n17603) );
  XNOR2_X1 U17736 ( .A(n17815), .B(n17816), .ZN(n17814) );
  NAND2_X1 U17737 ( .A1(b_1_), .A2(a_20_), .ZN(n17813) );
  XNOR2_X1 U17738 ( .A(n17817), .B(n17818), .ZN(n17502) );
  XNOR2_X1 U17739 ( .A(n17819), .B(n17820), .ZN(n17818) );
  NAND2_X1 U17740 ( .A1(b_1_), .A2(a_19_), .ZN(n17817) );
  XOR2_X1 U17741 ( .A(n17821), .B(n17822), .Z(n17607) );
  XOR2_X1 U17742 ( .A(n17823), .B(n17824), .Z(n17822) );
  XNOR2_X1 U17743 ( .A(n17825), .B(n17826), .ZN(n17490) );
  XOR2_X1 U17744 ( .A(n17827), .B(n17828), .Z(n17826) );
  XOR2_X1 U17745 ( .A(n17829), .B(n17830), .Z(n17611) );
  XNOR2_X1 U17746 ( .A(n17831), .B(n17832), .ZN(n17830) );
  XNOR2_X1 U17747 ( .A(n17833), .B(n17834), .ZN(n17478) );
  XOR2_X1 U17748 ( .A(n17835), .B(n17836), .Z(n17833) );
  XNOR2_X1 U17749 ( .A(n17837), .B(n17838), .ZN(n17615) );
  XOR2_X1 U17750 ( .A(n17839), .B(n17840), .Z(n17837) );
  XNOR2_X1 U17751 ( .A(n17841), .B(n17842), .ZN(n17466) );
  XOR2_X1 U17752 ( .A(n17843), .B(n17844), .Z(n17841) );
  XNOR2_X1 U17753 ( .A(n17845), .B(n17846), .ZN(n17619) );
  XOR2_X1 U17754 ( .A(n17847), .B(n17848), .Z(n17845) );
  XNOR2_X1 U17755 ( .A(n17849), .B(n17850), .ZN(n17454) );
  XOR2_X1 U17756 ( .A(n17851), .B(n17852), .Z(n17849) );
  XNOR2_X1 U17757 ( .A(n17853), .B(n17854), .ZN(n17623) );
  XOR2_X1 U17758 ( .A(n17855), .B(n17856), .Z(n17853) );
  XNOR2_X1 U17759 ( .A(n17857), .B(n17858), .ZN(n17442) );
  XOR2_X1 U17760 ( .A(n17859), .B(n17860), .Z(n17857) );
  XNOR2_X1 U17761 ( .A(n17861), .B(n17862), .ZN(n17627) );
  XOR2_X1 U17762 ( .A(n17863), .B(n17864), .Z(n17861) );
  XNOR2_X1 U17763 ( .A(n17865), .B(n17866), .ZN(n17430) );
  XOR2_X1 U17764 ( .A(n17867), .B(n17868), .Z(n17865) );
  XNOR2_X1 U17765 ( .A(n17869), .B(n17870), .ZN(n17631) );
  XOR2_X1 U17766 ( .A(n17871), .B(n17872), .Z(n17869) );
  XNOR2_X1 U17767 ( .A(n17873), .B(n17874), .ZN(n17418) );
  XOR2_X1 U17768 ( .A(n17875), .B(n17876), .Z(n17873) );
  XNOR2_X1 U17769 ( .A(n17877), .B(n17878), .ZN(n17410) );
  XOR2_X1 U17770 ( .A(n17879), .B(n17880), .Z(n17877) );
  XNOR2_X1 U17771 ( .A(n17881), .B(n17882), .ZN(n17403) );
  XOR2_X1 U17772 ( .A(n17883), .B(n17884), .Z(n17881) );
  XNOR2_X1 U17773 ( .A(n17885), .B(n17886), .ZN(n17635) );
  XOR2_X1 U17774 ( .A(n17887), .B(n17888), .Z(n17885) );
  XOR2_X1 U17775 ( .A(n17889), .B(n17890), .Z(n17638) );
  XNOR2_X1 U17776 ( .A(n17891), .B(n9952), .ZN(n17889) );
  XOR2_X1 U17777 ( .A(n17892), .B(n17893), .Z(n17643) );
  XOR2_X1 U17778 ( .A(n17894), .B(n17895), .Z(n17892) );
  INV_X1 U17779 ( .A(n17896), .ZN(n17647) );
  NOR2_X1 U17780 ( .A1(n10248), .A2(n10091), .ZN(n17896) );
  NAND2_X1 U17781 ( .A1(b_0_), .A2(a_0_), .ZN(n10091) );
  NAND2_X1 U17782 ( .A1(n17897), .A2(n17898), .ZN(n10248) );
  NAND2_X1 U17783 ( .A1(n17893), .A2(n17899), .ZN(n17898) );
  INV_X1 U17784 ( .A(n17900), .ZN(n17899) );
  NOR2_X1 U17785 ( .A1(n17894), .A2(n17895), .ZN(n17900) );
  NOR2_X1 U17786 ( .A1(n10094), .A2(n9983), .ZN(n17893) );
  NAND2_X1 U17787 ( .A1(n17895), .A2(n17894), .ZN(n17897) );
  NAND2_X1 U17788 ( .A1(n17901), .A2(n17902), .ZN(n17894) );
  NAND2_X1 U17789 ( .A1(n17890), .A2(n17903), .ZN(n17902) );
  NAND2_X1 U17790 ( .A1(n17904), .A2(n9952), .ZN(n17903) );
  INV_X1 U17791 ( .A(n17891), .ZN(n17904) );
  NOR2_X1 U17792 ( .A1(n10094), .A2(n10088), .ZN(n17890) );
  NAND2_X1 U17793 ( .A1(n17905), .A2(n17891), .ZN(n17901) );
  NAND2_X1 U17794 ( .A1(n17906), .A2(n17907), .ZN(n17891) );
  NAND2_X1 U17795 ( .A1(n17886), .A2(n17908), .ZN(n17907) );
  INV_X1 U17796 ( .A(n17909), .ZN(n17908) );
  NOR2_X1 U17797 ( .A1(n17887), .A2(n17888), .ZN(n17909) );
  NOR2_X1 U17798 ( .A1(n9982), .A2(n10088), .ZN(n17886) );
  NAND2_X1 U17799 ( .A1(n17888), .A2(n17887), .ZN(n17906) );
  NAND2_X1 U17800 ( .A1(n17910), .A2(n17911), .ZN(n17887) );
  NAND2_X1 U17801 ( .A1(n17882), .A2(n17912), .ZN(n17911) );
  INV_X1 U17802 ( .A(n17913), .ZN(n17912) );
  NOR2_X1 U17803 ( .A1(n17883), .A2(n17884), .ZN(n17913) );
  NOR2_X1 U17804 ( .A1(n9982), .A2(n10086), .ZN(n17882) );
  NAND2_X1 U17805 ( .A1(n17884), .A2(n17883), .ZN(n17910) );
  NAND2_X1 U17806 ( .A1(n17914), .A2(n17915), .ZN(n17883) );
  NAND2_X1 U17807 ( .A1(n17878), .A2(n17916), .ZN(n17915) );
  INV_X1 U17808 ( .A(n17917), .ZN(n17916) );
  NOR2_X1 U17809 ( .A1(n17879), .A2(n17880), .ZN(n17917) );
  NOR2_X1 U17810 ( .A1(n9982), .A2(n10085), .ZN(n17878) );
  NAND2_X1 U17811 ( .A1(n17880), .A2(n17879), .ZN(n17914) );
  NAND2_X1 U17812 ( .A1(n17918), .A2(n17919), .ZN(n17879) );
  NAND2_X1 U17813 ( .A1(n17874), .A2(n17920), .ZN(n17919) );
  INV_X1 U17814 ( .A(n17921), .ZN(n17920) );
  NOR2_X1 U17815 ( .A1(n17875), .A2(n17876), .ZN(n17921) );
  NOR2_X1 U17816 ( .A1(n9982), .A2(n10083), .ZN(n17874) );
  NAND2_X1 U17817 ( .A1(n17876), .A2(n17875), .ZN(n17918) );
  NAND2_X1 U17818 ( .A1(n17922), .A2(n17923), .ZN(n17875) );
  NAND2_X1 U17819 ( .A1(n17870), .A2(n17924), .ZN(n17923) );
  INV_X1 U17820 ( .A(n17925), .ZN(n17924) );
  NOR2_X1 U17821 ( .A1(n17871), .A2(n17872), .ZN(n17925) );
  NOR2_X1 U17822 ( .A1(n9982), .A2(n10081), .ZN(n17870) );
  NAND2_X1 U17823 ( .A1(n17872), .A2(n17871), .ZN(n17922) );
  NAND2_X1 U17824 ( .A1(n17926), .A2(n17927), .ZN(n17871) );
  NAND2_X1 U17825 ( .A1(n17866), .A2(n17928), .ZN(n17927) );
  INV_X1 U17826 ( .A(n17929), .ZN(n17928) );
  NOR2_X1 U17827 ( .A1(n17867), .A2(n17868), .ZN(n17929) );
  NOR2_X1 U17828 ( .A1(n9982), .A2(n9773), .ZN(n17866) );
  NAND2_X1 U17829 ( .A1(n17868), .A2(n17867), .ZN(n17926) );
  NAND2_X1 U17830 ( .A1(n17930), .A2(n17931), .ZN(n17867) );
  NAND2_X1 U17831 ( .A1(n17862), .A2(n17932), .ZN(n17931) );
  INV_X1 U17832 ( .A(n17933), .ZN(n17932) );
  NOR2_X1 U17833 ( .A1(n17863), .A2(n17864), .ZN(n17933) );
  NOR2_X1 U17834 ( .A1(n9982), .A2(n10079), .ZN(n17862) );
  NAND2_X1 U17835 ( .A1(n17864), .A2(n17863), .ZN(n17930) );
  NAND2_X1 U17836 ( .A1(n17934), .A2(n17935), .ZN(n17863) );
  NAND2_X1 U17837 ( .A1(n17858), .A2(n17936), .ZN(n17935) );
  INV_X1 U17838 ( .A(n17937), .ZN(n17936) );
  NOR2_X1 U17839 ( .A1(n17859), .A2(n17860), .ZN(n17937) );
  NOR2_X1 U17840 ( .A1(n9982), .A2(n10076), .ZN(n17858) );
  NAND2_X1 U17841 ( .A1(n17860), .A2(n17859), .ZN(n17934) );
  NAND2_X1 U17842 ( .A1(n17938), .A2(n17939), .ZN(n17859) );
  NAND2_X1 U17843 ( .A1(n17854), .A2(n17940), .ZN(n17939) );
  INV_X1 U17844 ( .A(n17941), .ZN(n17940) );
  NOR2_X1 U17845 ( .A1(n17855), .A2(n17856), .ZN(n17941) );
  NOR2_X1 U17846 ( .A1(n9982), .A2(n10073), .ZN(n17854) );
  NAND2_X1 U17847 ( .A1(n17856), .A2(n17855), .ZN(n17938) );
  NAND2_X1 U17848 ( .A1(n17942), .A2(n17943), .ZN(n17855) );
  NAND2_X1 U17849 ( .A1(n17850), .A2(n17944), .ZN(n17943) );
  INV_X1 U17850 ( .A(n17945), .ZN(n17944) );
  NOR2_X1 U17851 ( .A1(n17851), .A2(n17852), .ZN(n17945) );
  NOR2_X1 U17852 ( .A1(n9982), .A2(n9649), .ZN(n17850) );
  NAND2_X1 U17853 ( .A1(n17852), .A2(n17851), .ZN(n17942) );
  NAND2_X1 U17854 ( .A1(n17946), .A2(n17947), .ZN(n17851) );
  NAND2_X1 U17855 ( .A1(n17846), .A2(n17948), .ZN(n17947) );
  INV_X1 U17856 ( .A(n17949), .ZN(n17948) );
  NOR2_X1 U17857 ( .A1(n17847), .A2(n17848), .ZN(n17949) );
  NOR2_X1 U17858 ( .A1(n9982), .A2(n10070), .ZN(n17846) );
  NAND2_X1 U17859 ( .A1(n17848), .A2(n17847), .ZN(n17946) );
  NAND2_X1 U17860 ( .A1(n17950), .A2(n17951), .ZN(n17847) );
  NAND2_X1 U17861 ( .A1(n17842), .A2(n17952), .ZN(n17951) );
  INV_X1 U17862 ( .A(n17953), .ZN(n17952) );
  NOR2_X1 U17863 ( .A1(n17843), .A2(n17844), .ZN(n17953) );
  NOR2_X1 U17864 ( .A1(n9982), .A2(n10067), .ZN(n17842) );
  NAND2_X1 U17865 ( .A1(n17844), .A2(n17843), .ZN(n17950) );
  NAND2_X1 U17866 ( .A1(n17954), .A2(n17955), .ZN(n17843) );
  NAND2_X1 U17867 ( .A1(n17838), .A2(n17956), .ZN(n17955) );
  INV_X1 U17868 ( .A(n17957), .ZN(n17956) );
  NOR2_X1 U17869 ( .A1(n17839), .A2(n17840), .ZN(n17957) );
  NOR2_X1 U17870 ( .A1(n9982), .A2(n10065), .ZN(n17838) );
  NAND2_X1 U17871 ( .A1(n17840), .A2(n17839), .ZN(n17954) );
  NAND2_X1 U17872 ( .A1(n17958), .A2(n17959), .ZN(n17839) );
  NAND2_X1 U17873 ( .A1(n17834), .A2(n17960), .ZN(n17959) );
  INV_X1 U17874 ( .A(n17961), .ZN(n17960) );
  NOR2_X1 U17875 ( .A1(n17835), .A2(n17836), .ZN(n17961) );
  NOR2_X1 U17876 ( .A1(n9982), .A2(n9534), .ZN(n17834) );
  NAND2_X1 U17877 ( .A1(n17836), .A2(n17835), .ZN(n17958) );
  NAND2_X1 U17878 ( .A1(n17962), .A2(n17963), .ZN(n17835) );
  NAND2_X1 U17879 ( .A1(n17829), .A2(n17964), .ZN(n17963) );
  NAND2_X1 U17880 ( .A1(n17831), .A2(n17832), .ZN(n17964) );
  NOR2_X1 U17881 ( .A1(n9982), .A2(n10062), .ZN(n17829) );
  INV_X1 U17882 ( .A(n17965), .ZN(n17962) );
  NOR2_X1 U17883 ( .A1(n17832), .A2(n17831), .ZN(n17965) );
  NOR2_X1 U17884 ( .A1(n17966), .A2(n17967), .ZN(n17831) );
  INV_X1 U17885 ( .A(n17968), .ZN(n17967) );
  NAND2_X1 U17886 ( .A1(n17825), .A2(n17969), .ZN(n17968) );
  NAND2_X1 U17887 ( .A1(n17828), .A2(n17827), .ZN(n17969) );
  NOR2_X1 U17888 ( .A1(n9982), .A2(n10060), .ZN(n17825) );
  NOR2_X1 U17889 ( .A1(n17828), .A2(n17827), .ZN(n17966) );
  NAND2_X1 U17890 ( .A1(b_0_), .A2(a_18_), .ZN(n17827) );
  NAND2_X1 U17891 ( .A1(n17970), .A2(n17971), .ZN(n17828) );
  NAND2_X1 U17892 ( .A1(n17972), .A2(n17823), .ZN(n17971) );
  NAND2_X1 U17893 ( .A1(b_0_), .A2(a_19_), .ZN(n17823) );
  NAND2_X1 U17894 ( .A1(n17821), .A2(n17824), .ZN(n17972) );
  INV_X1 U17895 ( .A(n17973), .ZN(n17970) );
  NOR2_X1 U17896 ( .A1(n17824), .A2(n17821), .ZN(n17973) );
  NOR2_X1 U17897 ( .A1(n9982), .A2(n10058), .ZN(n17821) );
  NAND2_X1 U17898 ( .A1(n17974), .A2(n17975), .ZN(n17824) );
  NAND2_X1 U17899 ( .A1(n17976), .A2(b_1_), .ZN(n17975) );
  NOR2_X1 U17900 ( .A1(n17977), .A2(n9415), .ZN(n17976) );
  NOR2_X1 U17901 ( .A1(n17819), .A2(n17820), .ZN(n17977) );
  NAND2_X1 U17902 ( .A1(n17819), .A2(n17820), .ZN(n17974) );
  NAND2_X1 U17903 ( .A1(n17978), .A2(n17979), .ZN(n17820) );
  NAND2_X1 U17904 ( .A1(n17980), .A2(b_1_), .ZN(n17979) );
  NOR2_X1 U17905 ( .A1(n17981), .A2(n10054), .ZN(n17980) );
  NOR2_X1 U17906 ( .A1(n17815), .A2(n17816), .ZN(n17981) );
  NAND2_X1 U17907 ( .A1(n17815), .A2(n17816), .ZN(n17978) );
  NAND2_X1 U17908 ( .A1(n17982), .A2(n17983), .ZN(n17816) );
  NAND2_X1 U17909 ( .A1(n17984), .A2(b_1_), .ZN(n17983) );
  NOR2_X1 U17910 ( .A1(n17985), .A2(n9358), .ZN(n17984) );
  NOR2_X1 U17911 ( .A1(n17811), .A2(n17812), .ZN(n17985) );
  NAND2_X1 U17912 ( .A1(n17811), .A2(n17812), .ZN(n17982) );
  NAND2_X1 U17913 ( .A1(n17986), .A2(n17987), .ZN(n17812) );
  NAND2_X1 U17914 ( .A1(n17988), .A2(b_1_), .ZN(n17987) );
  NOR2_X1 U17915 ( .A1(n17989), .A2(n9330), .ZN(n17988) );
  NOR2_X1 U17916 ( .A1(n17807), .A2(n17808), .ZN(n17989) );
  NAND2_X1 U17917 ( .A1(n17807), .A2(n17808), .ZN(n17986) );
  NAND2_X1 U17918 ( .A1(n17990), .A2(n17991), .ZN(n17808) );
  NAND2_X1 U17919 ( .A1(n17992), .A2(b_1_), .ZN(n17991) );
  NOR2_X1 U17920 ( .A1(n17993), .A2(n10051), .ZN(n17992) );
  NOR2_X1 U17921 ( .A1(n17803), .A2(n17804), .ZN(n17993) );
  NAND2_X1 U17922 ( .A1(n17803), .A2(n17804), .ZN(n17990) );
  NAND2_X1 U17923 ( .A1(n17994), .A2(n17995), .ZN(n17804) );
  NAND2_X1 U17924 ( .A1(n17996), .A2(b_1_), .ZN(n17995) );
  NOR2_X1 U17925 ( .A1(n17997), .A2(n10050), .ZN(n17996) );
  NOR2_X1 U17926 ( .A1(n17799), .A2(n17800), .ZN(n17997) );
  NAND2_X1 U17927 ( .A1(n17799), .A2(n17800), .ZN(n17994) );
  NAND2_X1 U17928 ( .A1(n17998), .A2(n17999), .ZN(n17800) );
  NAND2_X1 U17929 ( .A1(n18000), .A2(b_1_), .ZN(n17999) );
  NOR2_X1 U17930 ( .A1(n18001), .A2(n10048), .ZN(n18000) );
  NOR2_X1 U17931 ( .A1(n17751), .A2(n17752), .ZN(n18001) );
  NAND2_X1 U17932 ( .A1(n17751), .A2(n17752), .ZN(n17998) );
  NAND2_X1 U17933 ( .A1(n18002), .A2(n18003), .ZN(n17752) );
  NAND2_X1 U17934 ( .A1(n18004), .A2(b_1_), .ZN(n18003) );
  NOR2_X1 U17935 ( .A1(n18005), .A2(n10047), .ZN(n18004) );
  NOR2_X1 U17936 ( .A1(n17759), .A2(n17760), .ZN(n18005) );
  NAND2_X1 U17937 ( .A1(n17759), .A2(n17760), .ZN(n18002) );
  NAND2_X1 U17938 ( .A1(n18006), .A2(n18007), .ZN(n17760) );
  NAND2_X1 U17939 ( .A1(n18008), .A2(b_1_), .ZN(n18007) );
  NOR2_X1 U17940 ( .A1(n18009), .A2(n11274), .ZN(n18008) );
  NOR2_X1 U17941 ( .A1(n17795), .A2(n17796), .ZN(n18009) );
  NAND2_X1 U17942 ( .A1(n17795), .A2(n17796), .ZN(n18006) );
  NAND2_X1 U17943 ( .A1(n18010), .A2(n18011), .ZN(n17796) );
  NAND2_X1 U17944 ( .A1(n18012), .A2(b_1_), .ZN(n18011) );
  NOR2_X1 U17945 ( .A1(n18013), .A2(n9136), .ZN(n18012) );
  NOR2_X1 U17946 ( .A1(n17771), .A2(n17772), .ZN(n18013) );
  NAND2_X1 U17947 ( .A1(n17771), .A2(n17772), .ZN(n18010) );
  NAND2_X1 U17948 ( .A1(n17792), .A2(n18014), .ZN(n17772) );
  NAND2_X1 U17949 ( .A1(n17790), .A2(n17791), .ZN(n18014) );
  NOR2_X1 U17950 ( .A1(n9982), .A2(n9121), .ZN(n17791) );
  NOR2_X1 U17951 ( .A1(n10043), .A2(n10094), .ZN(n17790) );
  NAND2_X1 U17952 ( .A1(n18015), .A2(n9025), .ZN(n17792) );
  NOR2_X1 U17953 ( .A1(n10044), .A2(n10043), .ZN(n10045) );
  NOR2_X1 U17954 ( .A1(n10094), .A2(n9982), .ZN(n18015) );
  NOR2_X1 U17955 ( .A1(n10094), .A2(n9121), .ZN(n17771) );
  NOR2_X1 U17956 ( .A1(n10094), .A2(n9136), .ZN(n17795) );
  NOR2_X1 U17957 ( .A1(n10094), .A2(n11274), .ZN(n17759) );
  NOR2_X1 U17958 ( .A1(n10094), .A2(n10047), .ZN(n17751) );
  NOR2_X1 U17959 ( .A1(n10094), .A2(n10048), .ZN(n17799) );
  NOR2_X1 U17960 ( .A1(n10094), .A2(n10050), .ZN(n17803) );
  NOR2_X1 U17961 ( .A1(n10094), .A2(n10051), .ZN(n17807) );
  NOR2_X1 U17962 ( .A1(n10094), .A2(n9330), .ZN(n17811) );
  NOR2_X1 U17963 ( .A1(n10094), .A2(n9358), .ZN(n17815) );
  NOR2_X1 U17964 ( .A1(n10094), .A2(n10054), .ZN(n17819) );
  NAND2_X1 U17965 ( .A1(b_0_), .A2(a_17_), .ZN(n17832) );
  NOR2_X1 U17966 ( .A1(n10094), .A2(n10062), .ZN(n17836) );
  NOR2_X1 U17967 ( .A1(n10094), .A2(n9534), .ZN(n17840) );
  NOR2_X1 U17968 ( .A1(n10094), .A2(n10065), .ZN(n17844) );
  NOR2_X1 U17969 ( .A1(n10094), .A2(n10067), .ZN(n17848) );
  NOR2_X1 U17970 ( .A1(n10094), .A2(n10070), .ZN(n17852) );
  NOR2_X1 U17971 ( .A1(n10094), .A2(n9649), .ZN(n17856) );
  NOR2_X1 U17972 ( .A1(n10094), .A2(n10073), .ZN(n17860) );
  NOR2_X1 U17973 ( .A1(n10094), .A2(n10076), .ZN(n17864) );
  NOR2_X1 U17974 ( .A1(n10094), .A2(n10079), .ZN(n17868) );
  NOR2_X1 U17975 ( .A1(n10094), .A2(n9773), .ZN(n17872) );
  NOR2_X1 U17976 ( .A1(n10094), .A2(n10081), .ZN(n17876) );
  NOR2_X1 U17977 ( .A1(n10094), .A2(n10083), .ZN(n17880) );
  NOR2_X1 U17978 ( .A1(n10094), .A2(n10085), .ZN(n17884) );
  NOR2_X1 U17979 ( .A1(n10094), .A2(n10086), .ZN(n17888) );
  INV_X1 U17980 ( .A(n9952), .ZN(n17905) );
  NAND2_X1 U17981 ( .A1(b_1_), .A2(a_1_), .ZN(n9952) );
  NOR2_X1 U17982 ( .A1(n9982), .A2(n10093), .ZN(n17895) );
  NOR2_X1 U17983 ( .A1(n9980), .A2(n9979), .ZN(n9032) );
  INV_X1 U17984 ( .A(operation_0_), .ZN(n9980) );
  NAND2_X1 U17985 ( .A1(n18017), .A2(n18018), .ZN(n18016) );
  NAND2_X1 U17986 ( .A1(n9029), .A2(n18019), .ZN(n18018) );
  NAND2_X1 U17987 ( .A1(n18020), .A2(n18021), .ZN(n18019) );
  NAND2_X1 U17988 ( .A1(b_0_), .A2(n18022), .ZN(n18021) );
  NAND2_X1 U17989 ( .A1(a_0_), .A2(n9970), .ZN(n18022) );
  NAND2_X1 U17990 ( .A1(n10089), .A2(n10093), .ZN(n18020) );
  INV_X1 U17991 ( .A(n9970), .ZN(n10089) );
  NAND2_X1 U17992 ( .A1(n18023), .A2(n18024), .ZN(n9970) );
  NAND2_X1 U17993 ( .A1(n18025), .A2(n9982), .ZN(n18024) );
  NAND2_X1 U17994 ( .A1(n9950), .A2(n9983), .ZN(n18025) );
  INV_X1 U17995 ( .A(n9941), .ZN(n9950) );
  NAND2_X1 U17996 ( .A1(a_1_), .A2(n9941), .ZN(n18023) );
  NAND2_X1 U17997 ( .A1(n18026), .A2(n18027), .ZN(n9941) );
  NAND2_X1 U17998 ( .A1(n18028), .A2(n10087), .ZN(n18027) );
  NAND2_X1 U17999 ( .A1(n10088), .A2(n9921), .ZN(n18028) );
  NAND2_X1 U18000 ( .A1(a_2_), .A2(n9913), .ZN(n18026) );
  INV_X1 U18001 ( .A(n9921), .ZN(n9913) );
  NAND2_X1 U18002 ( .A1(n18029), .A2(n18030), .ZN(n9921) );
  NAND2_X1 U18003 ( .A1(b_3_), .A2(n18031), .ZN(n18030) );
  NAND2_X1 U18004 ( .A1(a_3_), .A2(n9894), .ZN(n18031) );
  NAND2_X1 U18005 ( .A1(n9884), .A2(n10086), .ZN(n18029) );
  INV_X1 U18006 ( .A(n9894), .ZN(n9884) );
  NAND2_X1 U18007 ( .A1(n18032), .A2(n18033), .ZN(n9894) );
  NAND2_X1 U18008 ( .A1(n18034), .A2(n10084), .ZN(n18033) );
  NAND2_X1 U18009 ( .A1(n9864), .A2(n10085), .ZN(n18034) );
  INV_X1 U18010 ( .A(n9856), .ZN(n9864) );
  NAND2_X1 U18011 ( .A1(a_4_), .A2(n9856), .ZN(n18032) );
  NAND2_X1 U18012 ( .A1(n18035), .A2(n18036), .ZN(n9856) );
  NAND2_X1 U18013 ( .A1(n18037), .A2(n10082), .ZN(n18036) );
  NAND2_X1 U18014 ( .A1(n9835), .A2(n10083), .ZN(n18037) );
  INV_X1 U18015 ( .A(n9827), .ZN(n9835) );
  NAND2_X1 U18016 ( .A1(a_5_), .A2(n9827), .ZN(n18035) );
  NAND2_X1 U18017 ( .A1(n18038), .A2(n18039), .ZN(n9827) );
  NAND2_X1 U18018 ( .A1(n18040), .A2(n10080), .ZN(n18039) );
  INV_X1 U18019 ( .A(b_6_), .ZN(n10080) );
  NAND2_X1 U18020 ( .A1(n10081), .A2(n9806), .ZN(n18040) );
  NAND2_X1 U18021 ( .A1(a_6_), .A2(n9797), .ZN(n18038) );
  INV_X1 U18022 ( .A(n9806), .ZN(n9797) );
  NAND2_X1 U18023 ( .A1(n18041), .A2(n18042), .ZN(n9806) );
  NAND2_X1 U18024 ( .A1(b_7_), .A2(n18043), .ZN(n18042) );
  NAND2_X1 U18025 ( .A1(a_7_), .A2(n9779), .ZN(n18043) );
  NAND2_X1 U18026 ( .A1(n9769), .A2(n9773), .ZN(n18041) );
  INV_X1 U18027 ( .A(n9779), .ZN(n9769) );
  NAND2_X1 U18028 ( .A1(n18044), .A2(n18045), .ZN(n9779) );
  NAND2_X1 U18029 ( .A1(n18046), .A2(n10078), .ZN(n18045) );
  NAND2_X1 U18030 ( .A1(n9740), .A2(n10079), .ZN(n18046) );
  INV_X1 U18031 ( .A(n9732), .ZN(n9740) );
  NAND2_X1 U18032 ( .A1(a_8_), .A2(n9732), .ZN(n18044) );
  NAND2_X1 U18033 ( .A1(n18047), .A2(n18048), .ZN(n9732) );
  NAND2_X1 U18034 ( .A1(n18049), .A2(n10075), .ZN(n18048) );
  INV_X1 U18035 ( .A(b_9_), .ZN(n10075) );
  NAND2_X1 U18036 ( .A1(n9711), .A2(n10076), .ZN(n18049) );
  INV_X1 U18037 ( .A(n9703), .ZN(n9711) );
  NAND2_X1 U18038 ( .A1(a_9_), .A2(n9703), .ZN(n18047) );
  NAND2_X1 U18039 ( .A1(n18050), .A2(n18051), .ZN(n9703) );
  NAND2_X1 U18040 ( .A1(n18052), .A2(n10072), .ZN(n18051) );
  INV_X1 U18041 ( .A(b_10_), .ZN(n10072) );
  NAND2_X1 U18042 ( .A1(n10073), .A2(n9682), .ZN(n18052) );
  NAND2_X1 U18043 ( .A1(a_10_), .A2(n9674), .ZN(n18050) );
  INV_X1 U18044 ( .A(n9682), .ZN(n9674) );
  NAND2_X1 U18045 ( .A1(n18053), .A2(n18054), .ZN(n9682) );
  NAND2_X1 U18046 ( .A1(b_11_), .A2(n18055), .ZN(n18054) );
  NAND2_X1 U18047 ( .A1(a_11_), .A2(n9655), .ZN(n18055) );
  NAND2_X1 U18048 ( .A1(n9645), .A2(n9649), .ZN(n18053) );
  INV_X1 U18049 ( .A(n9655), .ZN(n9645) );
  NAND2_X1 U18050 ( .A1(n18056), .A2(n18057), .ZN(n9655) );
  NAND2_X1 U18051 ( .A1(n18058), .A2(n10069), .ZN(n18057) );
  INV_X1 U18052 ( .A(b_12_), .ZN(n10069) );
  NAND2_X1 U18053 ( .A1(n9625), .A2(n10070), .ZN(n18058) );
  INV_X1 U18054 ( .A(n9617), .ZN(n9625) );
  NAND2_X1 U18055 ( .A1(a_12_), .A2(n9617), .ZN(n18056) );
  NAND2_X1 U18056 ( .A1(n18059), .A2(n18060), .ZN(n9617) );
  NAND2_X1 U18057 ( .A1(n18061), .A2(n10066), .ZN(n18060) );
  INV_X1 U18058 ( .A(b_13_), .ZN(n10066) );
  NAND2_X1 U18059 ( .A1(n9596), .A2(n10067), .ZN(n18061) );
  INV_X1 U18060 ( .A(n9588), .ZN(n9596) );
  NAND2_X1 U18061 ( .A1(a_13_), .A2(n9588), .ZN(n18059) );
  NAND2_X1 U18062 ( .A1(n18062), .A2(n18063), .ZN(n9588) );
  NAND2_X1 U18063 ( .A1(n18064), .A2(n10064), .ZN(n18063) );
  INV_X1 U18064 ( .A(b_14_), .ZN(n10064) );
  NAND2_X1 U18065 ( .A1(n9567), .A2(n10065), .ZN(n18064) );
  INV_X1 U18066 ( .A(n9559), .ZN(n9567) );
  NAND2_X1 U18067 ( .A1(a_14_), .A2(n9559), .ZN(n18062) );
  NAND2_X1 U18068 ( .A1(n18065), .A2(n18066), .ZN(n9559) );
  NAND2_X1 U18069 ( .A1(n18067), .A2(n10063), .ZN(n18066) );
  INV_X1 U18070 ( .A(b_15_), .ZN(n10063) );
  NAND2_X1 U18071 ( .A1(n9534), .A2(n9530), .ZN(n18067) );
  NAND2_X1 U18072 ( .A1(a_15_), .A2(n9540), .ZN(n18065) );
  INV_X1 U18073 ( .A(n9530), .ZN(n9540) );
  NAND2_X1 U18074 ( .A1(n18068), .A2(n18069), .ZN(n9530) );
  NAND2_X1 U18075 ( .A1(b_16_), .A2(n18070), .ZN(n18069) );
  NAND2_X1 U18076 ( .A1(a_16_), .A2(n9502), .ZN(n18070) );
  INV_X1 U18077 ( .A(n9510), .ZN(n9502) );
  NAND2_X1 U18078 ( .A1(n9510), .A2(n10062), .ZN(n18068) );
  NAND2_X1 U18079 ( .A1(n18071), .A2(n18072), .ZN(n9510) );
  NAND2_X1 U18080 ( .A1(b_17_), .A2(n18073), .ZN(n18072) );
  NAND2_X1 U18081 ( .A1(a_17_), .A2(n9473), .ZN(n18073) );
  NAND2_X1 U18082 ( .A1(n9481), .A2(n10060), .ZN(n18071) );
  INV_X1 U18083 ( .A(n9473), .ZN(n9481) );
  NAND2_X1 U18084 ( .A1(n18074), .A2(n18075), .ZN(n9473) );
  NAND2_X1 U18085 ( .A1(n18076), .A2(n10057), .ZN(n18075) );
  INV_X1 U18086 ( .A(b_18_), .ZN(n10057) );
  NAND2_X1 U18087 ( .A1(n9448), .A2(n10058), .ZN(n18076) );
  INV_X1 U18088 ( .A(n9440), .ZN(n9448) );
  NAND2_X1 U18089 ( .A1(a_18_), .A2(n9440), .ZN(n18074) );
  NAND2_X1 U18090 ( .A1(n18077), .A2(n18078), .ZN(n9440) );
  NAND2_X1 U18091 ( .A1(n18079), .A2(n10056), .ZN(n18078) );
  INV_X1 U18092 ( .A(b_19_), .ZN(n10056) );
  NAND2_X1 U18093 ( .A1(n9411), .A2(n9415), .ZN(n18079) );
  INV_X1 U18094 ( .A(n9421), .ZN(n9411) );
  NAND2_X1 U18095 ( .A1(a_19_), .A2(n9421), .ZN(n18077) );
  NAND2_X1 U18096 ( .A1(n18080), .A2(n18081), .ZN(n9421) );
  NAND2_X1 U18097 ( .A1(n18082), .A2(n10053), .ZN(n18081) );
  INV_X1 U18098 ( .A(b_20_), .ZN(n10053) );
  NAND2_X1 U18099 ( .A1(n10054), .A2(n9391), .ZN(n18082) );
  NAND2_X1 U18100 ( .A1(a_20_), .A2(n9383), .ZN(n18080) );
  INV_X1 U18101 ( .A(n9391), .ZN(n9383) );
  NAND2_X1 U18102 ( .A1(n18083), .A2(n18084), .ZN(n9391) );
  NAND2_X1 U18103 ( .A1(b_21_), .A2(n18085), .ZN(n18084) );
  NAND2_X1 U18104 ( .A1(a_21_), .A2(n9364), .ZN(n18085) );
  INV_X1 U18105 ( .A(n9354), .ZN(n9364) );
  NAND2_X1 U18106 ( .A1(n9354), .A2(n9358), .ZN(n18083) );
  NAND2_X1 U18107 ( .A1(n18086), .A2(n18087), .ZN(n9354) );
  NAND2_X1 U18108 ( .A1(b_22_), .A2(n18088), .ZN(n18087) );
  NAND2_X1 U18109 ( .A1(a_22_), .A2(n9336), .ZN(n18088) );
  INV_X1 U18110 ( .A(n9326), .ZN(n9336) );
  NAND2_X1 U18111 ( .A1(n9326), .A2(n9330), .ZN(n18086) );
  NAND2_X1 U18112 ( .A1(n18089), .A2(n18090), .ZN(n9326) );
  NAND2_X1 U18113 ( .A1(b_23_), .A2(n18091), .ZN(n18090) );
  NAND2_X1 U18114 ( .A1(a_23_), .A2(n9308), .ZN(n18091) );
  NAND2_X1 U18115 ( .A1(n9298), .A2(n10051), .ZN(n18089) );
  INV_X1 U18116 ( .A(n9308), .ZN(n9298) );
  NAND2_X1 U18117 ( .A1(n9281), .A2(n18092), .ZN(n9308) );
  NAND2_X1 U18118 ( .A1(n9279), .A2(n9280), .ZN(n18092) );
  INV_X1 U18119 ( .A(n9269), .ZN(n9279) );
  NAND2_X1 U18120 ( .A1(n18093), .A2(n18094), .ZN(n9269) );
  NAND2_X1 U18121 ( .A1(b_25_), .A2(n18095), .ZN(n18094) );
  NAND2_X1 U18122 ( .A1(a_25_), .A2(n9251), .ZN(n18095) );
  INV_X1 U18123 ( .A(n9241), .ZN(n9251) );
  NAND2_X1 U18124 ( .A1(n9241), .A2(n10048), .ZN(n18093) );
  NAND2_X1 U18125 ( .A1(n18096), .A2(n18097), .ZN(n9241) );
  NAND2_X1 U18126 ( .A1(b_26_), .A2(n18098), .ZN(n18097) );
  NAND2_X1 U18127 ( .A1(a_26_), .A2(n9223), .ZN(n18098) );
  INV_X1 U18128 ( .A(n9213), .ZN(n9223) );
  NAND2_X1 U18129 ( .A1(n9213), .A2(n10047), .ZN(n18096) );
  NAND2_X1 U18130 ( .A1(n9196), .A2(n18099), .ZN(n9213) );
  NAND2_X1 U18131 ( .A1(n9185), .A2(n9195), .ZN(n18099) );
  NAND2_X1 U18132 ( .A1(n9158), .A2(n18100), .ZN(n9185) );
  NAND2_X1 U18133 ( .A1(n9146), .A2(n9157), .ZN(n18100) );
  INV_X1 U18134 ( .A(n9155), .ZN(n9146) );
  NAND2_X1 U18135 ( .A1(n18101), .A2(n18102), .ZN(n9155) );
  NAND2_X1 U18136 ( .A1(n18103), .A2(n10046), .ZN(n18102) );
  INV_X1 U18137 ( .A(b_29_), .ZN(n10046) );
  NAND2_X1 U18138 ( .A1(n9117), .A2(n9121), .ZN(n18103) );
  INV_X1 U18139 ( .A(n9127), .ZN(n9117) );
  NAND2_X1 U18140 ( .A1(a_29_), .A2(n9127), .ZN(n18101) );
  NAND2_X1 U18141 ( .A1(n9078), .A2(n18104), .ZN(n9127) );
  NAND2_X1 U18142 ( .A1(n9100), .A2(n9068), .ZN(n18104) );
  INV_X1 U18143 ( .A(n9074), .ZN(n9068) );
  NOR2_X1 U18144 ( .A1(n9077), .A2(a_31_), .ZN(n9074) );
  NOR2_X1 U18145 ( .A1(n9979), .A2(operation_0_), .ZN(n9066) );
  NAND2_X1 U18146 ( .A1(n9065), .A2(n18105), .ZN(n18017) );
  NAND2_X1 U18147 ( .A1(n18106), .A2(n18107), .ZN(n18105) );
  NAND2_X1 U18148 ( .A1(n18108), .A2(n10094), .ZN(n18107) );
  NAND2_X1 U18149 ( .A1(n10093), .A2(n10090), .ZN(n18108) );
  NAND2_X1 U18150 ( .A1(n9971), .A2(a_0_), .ZN(n18106) );
  INV_X1 U18151 ( .A(n10090), .ZN(n9971) );
  NAND2_X1 U18152 ( .A1(n18109), .A2(n18110), .ZN(n10090) );
  NAND2_X1 U18153 ( .A1(b_1_), .A2(n18111), .ZN(n18110) );
  NAND2_X1 U18154 ( .A1(n9942), .A2(a_1_), .ZN(n18111) );
  INV_X1 U18155 ( .A(n9951), .ZN(n9942) );
  NAND2_X1 U18156 ( .A1(n9951), .A2(n9983), .ZN(n18109) );
  NAND2_X1 U18157 ( .A1(n18112), .A2(n18113), .ZN(n9951) );
  NAND2_X1 U18158 ( .A1(b_2_), .A2(n18114), .ZN(n18113) );
  NAND2_X1 U18159 ( .A1(a_2_), .A2(n9914), .ZN(n18114) );
  NAND2_X1 U18160 ( .A1(n9922), .A2(n10088), .ZN(n18112) );
  INV_X1 U18161 ( .A(a_2_), .ZN(n10088) );
  INV_X1 U18162 ( .A(n9914), .ZN(n9922) );
  NAND2_X1 U18163 ( .A1(n18115), .A2(n18116), .ZN(n9914) );
  NAND2_X1 U18164 ( .A1(n18117), .A2(n9888), .ZN(n18116) );
  INV_X1 U18165 ( .A(b_3_), .ZN(n9888) );
  NAND2_X1 U18166 ( .A1(n10086), .A2(n9885), .ZN(n18117) );
  INV_X1 U18167 ( .A(a_3_), .ZN(n10086) );
  NAND2_X1 U18168 ( .A1(n9895), .A2(a_3_), .ZN(n18115) );
  INV_X1 U18169 ( .A(n9885), .ZN(n9895) );
  NAND2_X1 U18170 ( .A1(n18118), .A2(n18119), .ZN(n9885) );
  NAND2_X1 U18171 ( .A1(b_4_), .A2(n18120), .ZN(n18119) );
  NAND2_X1 U18172 ( .A1(n9857), .A2(a_4_), .ZN(n18120) );
  INV_X1 U18173 ( .A(n9865), .ZN(n9857) );
  NAND2_X1 U18174 ( .A1(n9865), .A2(n10085), .ZN(n18118) );
  INV_X1 U18175 ( .A(a_4_), .ZN(n10085) );
  NAND2_X1 U18176 ( .A1(n18121), .A2(n18122), .ZN(n9865) );
  NAND2_X1 U18177 ( .A1(b_5_), .A2(n18123), .ZN(n18122) );
  NAND2_X1 U18178 ( .A1(n9828), .A2(a_5_), .ZN(n18123) );
  INV_X1 U18179 ( .A(n9836), .ZN(n9828) );
  NAND2_X1 U18180 ( .A1(n9836), .A2(n10083), .ZN(n18121) );
  NAND2_X1 U18181 ( .A1(n18124), .A2(n18125), .ZN(n9836) );
  NAND2_X1 U18182 ( .A1(b_6_), .A2(n18126), .ZN(n18125) );
  NAND2_X1 U18183 ( .A1(a_6_), .A2(n9798), .ZN(n18126) );
  NAND2_X1 U18184 ( .A1(n9807), .A2(n10081), .ZN(n18124) );
  INV_X1 U18185 ( .A(n9798), .ZN(n9807) );
  NAND2_X1 U18186 ( .A1(n18127), .A2(n18128), .ZN(n9798) );
  NAND2_X1 U18187 ( .A1(n18129), .A2(n16032), .ZN(n18128) );
  INV_X1 U18188 ( .A(b_7_), .ZN(n16032) );
  NAND2_X1 U18189 ( .A1(n9773), .A2(n9770), .ZN(n18129) );
  INV_X1 U18190 ( .A(a_7_), .ZN(n9773) );
  NAND2_X1 U18191 ( .A1(n9780), .A2(a_7_), .ZN(n18127) );
  INV_X1 U18192 ( .A(n9770), .ZN(n9780) );
  NAND2_X1 U18193 ( .A1(n18130), .A2(n18131), .ZN(n9770) );
  NAND2_X1 U18194 ( .A1(b_8_), .A2(n18132), .ZN(n18131) );
  NAND2_X1 U18195 ( .A1(n9733), .A2(a_8_), .ZN(n18132) );
  INV_X1 U18196 ( .A(n9741), .ZN(n9733) );
  NAND2_X1 U18197 ( .A1(n9741), .A2(n10079), .ZN(n18130) );
  INV_X1 U18198 ( .A(a_8_), .ZN(n10079) );
  NAND2_X1 U18199 ( .A1(n18133), .A2(n18134), .ZN(n9741) );
  NAND2_X1 U18200 ( .A1(b_9_), .A2(n18135), .ZN(n18134) );
  NAND2_X1 U18201 ( .A1(n9704), .A2(a_9_), .ZN(n18135) );
  INV_X1 U18202 ( .A(n9712), .ZN(n9704) );
  NAND2_X1 U18203 ( .A1(n9712), .A2(n10076), .ZN(n18133) );
  NAND2_X1 U18204 ( .A1(n18136), .A2(n18137), .ZN(n9712) );
  NAND2_X1 U18205 ( .A1(b_10_), .A2(n18138), .ZN(n18137) );
  NAND2_X1 U18206 ( .A1(a_10_), .A2(n9675), .ZN(n18138) );
  NAND2_X1 U18207 ( .A1(n9683), .A2(n10073), .ZN(n18136) );
  INV_X1 U18208 ( .A(n9675), .ZN(n9683) );
  NAND2_X1 U18209 ( .A1(n18139), .A2(n18140), .ZN(n9675) );
  NAND2_X1 U18210 ( .A1(n18141), .A2(n10071), .ZN(n18140) );
  NAND2_X1 U18211 ( .A1(n9649), .A2(n9646), .ZN(n18141) );
  NAND2_X1 U18212 ( .A1(n9656), .A2(a_11_), .ZN(n18139) );
  INV_X1 U18213 ( .A(n9646), .ZN(n9656) );
  NAND2_X1 U18214 ( .A1(n18142), .A2(n18143), .ZN(n9646) );
  NAND2_X1 U18215 ( .A1(b_12_), .A2(n18144), .ZN(n18143) );
  NAND2_X1 U18216 ( .A1(n9618), .A2(a_12_), .ZN(n18144) );
  INV_X1 U18217 ( .A(n9626), .ZN(n9618) );
  NAND2_X1 U18218 ( .A1(n9626), .A2(n10070), .ZN(n18142) );
  NAND2_X1 U18219 ( .A1(n18145), .A2(n18146), .ZN(n9626) );
  NAND2_X1 U18220 ( .A1(b_13_), .A2(n18147), .ZN(n18146) );
  NAND2_X1 U18221 ( .A1(n9589), .A2(a_13_), .ZN(n18147) );
  INV_X1 U18222 ( .A(n9597), .ZN(n9589) );
  NAND2_X1 U18223 ( .A1(n9597), .A2(n10067), .ZN(n18145) );
  INV_X1 U18224 ( .A(a_13_), .ZN(n10067) );
  NAND2_X1 U18225 ( .A1(n18148), .A2(n18149), .ZN(n9597) );
  NAND2_X1 U18226 ( .A1(b_14_), .A2(n18150), .ZN(n18149) );
  NAND2_X1 U18227 ( .A1(n9560), .A2(a_14_), .ZN(n18150) );
  INV_X1 U18228 ( .A(n9568), .ZN(n9560) );
  NAND2_X1 U18229 ( .A1(n9568), .A2(n10065), .ZN(n18148) );
  NAND2_X1 U18230 ( .A1(n18151), .A2(n18152), .ZN(n9568) );
  NAND2_X1 U18231 ( .A1(b_15_), .A2(n18153), .ZN(n18152) );
  NAND2_X1 U18232 ( .A1(a_15_), .A2(n9541), .ZN(n18153) );
  NAND2_X1 U18233 ( .A1(n9531), .A2(n9534), .ZN(n18151) );
  INV_X1 U18234 ( .A(n9541), .ZN(n9531) );
  NAND2_X1 U18235 ( .A1(n18154), .A2(n18155), .ZN(n9541) );
  NAND2_X1 U18236 ( .A1(n18156), .A2(n10061), .ZN(n18155) );
  INV_X1 U18237 ( .A(b_16_), .ZN(n10061) );
  NAND2_X1 U18238 ( .A1(n9511), .A2(n10062), .ZN(n18156) );
  INV_X1 U18239 ( .A(a_16_), .ZN(n10062) );
  INV_X1 U18240 ( .A(n9503), .ZN(n9511) );
  NAND2_X1 U18241 ( .A1(a_16_), .A2(n9503), .ZN(n18154) );
  NAND2_X1 U18242 ( .A1(n18157), .A2(n18158), .ZN(n9503) );
  NAND2_X1 U18243 ( .A1(n18159), .A2(n10059), .ZN(n18158) );
  NAND2_X1 U18244 ( .A1(n10060), .A2(n9482), .ZN(n18159) );
  INV_X1 U18245 ( .A(a_17_), .ZN(n10060) );
  NAND2_X1 U18246 ( .A1(n9474), .A2(a_17_), .ZN(n18157) );
  INV_X1 U18247 ( .A(n9482), .ZN(n9474) );
  NAND2_X1 U18248 ( .A1(n18160), .A2(n18161), .ZN(n9482) );
  NAND2_X1 U18249 ( .A1(b_18_), .A2(n18162), .ZN(n18161) );
  NAND2_X1 U18250 ( .A1(n9441), .A2(a_18_), .ZN(n18162) );
  INV_X1 U18251 ( .A(n9449), .ZN(n9441) );
  NAND2_X1 U18252 ( .A1(n9449), .A2(n10058), .ZN(n18160) );
  NAND2_X1 U18253 ( .A1(n18163), .A2(n18164), .ZN(n9449) );
  NAND2_X1 U18254 ( .A1(b_19_), .A2(n18165), .ZN(n18164) );
  NAND2_X1 U18255 ( .A1(n9422), .A2(a_19_), .ZN(n18165) );
  INV_X1 U18256 ( .A(n9412), .ZN(n9422) );
  NAND2_X1 U18257 ( .A1(n9412), .A2(n9415), .ZN(n18163) );
  NAND2_X1 U18258 ( .A1(n18166), .A2(n18167), .ZN(n9412) );
  NAND2_X1 U18259 ( .A1(b_20_), .A2(n18168), .ZN(n18167) );
  NAND2_X1 U18260 ( .A1(a_20_), .A2(n9384), .ZN(n18168) );
  NAND2_X1 U18261 ( .A1(n9392), .A2(n10054), .ZN(n18166) );
  INV_X1 U18262 ( .A(n9384), .ZN(n9392) );
  NAND2_X1 U18263 ( .A1(n18169), .A2(n18170), .ZN(n9384) );
  NAND2_X1 U18264 ( .A1(n18171), .A2(n10052), .ZN(n18170) );
  NAND2_X1 U18265 ( .A1(n9355), .A2(n9358), .ZN(n18171) );
  INV_X1 U18266 ( .A(a_21_), .ZN(n9358) );
  INV_X1 U18267 ( .A(n9365), .ZN(n9355) );
  NAND2_X1 U18268 ( .A1(a_21_), .A2(n9365), .ZN(n18169) );
  NAND2_X1 U18269 ( .A1(n18172), .A2(n18173), .ZN(n9365) );
  NAND2_X1 U18270 ( .A1(n18174), .A2(n12294), .ZN(n18173) );
  INV_X1 U18271 ( .A(b_22_), .ZN(n12294) );
  NAND2_X1 U18272 ( .A1(n9327), .A2(n9330), .ZN(n18174) );
  INV_X1 U18273 ( .A(a_22_), .ZN(n9330) );
  INV_X1 U18274 ( .A(n9337), .ZN(n9327) );
  NAND2_X1 U18275 ( .A1(a_22_), .A2(n9337), .ZN(n18172) );
  NAND2_X1 U18276 ( .A1(n18175), .A2(n18176), .ZN(n9337) );
  NAND2_X1 U18277 ( .A1(n18177), .A2(n9302), .ZN(n18176) );
  NAND2_X1 U18278 ( .A1(n9299), .A2(n10051), .ZN(n18177) );
  INV_X1 U18279 ( .A(n9309), .ZN(n9299) );
  NAND2_X1 U18280 ( .A1(a_23_), .A2(n9309), .ZN(n18175) );
  NAND2_X1 U18281 ( .A1(n9281), .A2(n18178), .ZN(n9309) );
  NAND2_X1 U18282 ( .A1(n9280), .A2(n9271), .ZN(n18178) );
  NAND2_X1 U18283 ( .A1(n18179), .A2(n18180), .ZN(n9271) );
  NAND2_X1 U18284 ( .A1(n18181), .A2(n9245), .ZN(n18180) );
  NAND2_X1 U18285 ( .A1(n9242), .A2(n10048), .ZN(n18181) );
  INV_X1 U18286 ( .A(n9252), .ZN(n9242) );
  NAND2_X1 U18287 ( .A1(a_25_), .A2(n9252), .ZN(n18179) );
  NAND2_X1 U18288 ( .A1(n18182), .A2(n18183), .ZN(n9252) );
  NAND2_X1 U18289 ( .A1(n18184), .A2(n9217), .ZN(n18183) );
  NAND2_X1 U18290 ( .A1(n10047), .A2(n9214), .ZN(n18184) );
  NAND2_X1 U18291 ( .A1(n9224), .A2(a_26_), .ZN(n18182) );
  INV_X1 U18292 ( .A(n9214), .ZN(n9224) );
  NAND2_X1 U18293 ( .A1(n9196), .A2(n18185), .ZN(n9214) );
  NAND2_X1 U18294 ( .A1(n9195), .A2(n9186), .ZN(n18185) );
  NAND2_X1 U18295 ( .A1(n9158), .A2(n18186), .ZN(n9186) );
  NAND2_X1 U18296 ( .A1(n9157), .A2(n9147), .ZN(n18186) );
  NAND2_X1 U18297 ( .A1(n18187), .A2(n18188), .ZN(n9147) );
  NAND2_X1 U18298 ( .A1(b_29_), .A2(n18189), .ZN(n18188) );
  NAND2_X1 U18299 ( .A1(a_29_), .A2(n9128), .ZN(n18189) );
  NAND2_X1 U18300 ( .A1(n9118), .A2(n9121), .ZN(n18187) );
  INV_X1 U18301 ( .A(n9128), .ZN(n9118) );
  NAND2_X1 U18302 ( .A1(n9078), .A2(n18190), .ZN(n9128) );
  NAND2_X1 U18303 ( .A1(n9082), .A2(n9100), .ZN(n18190) );
  NAND2_X1 U18304 ( .A1(b_30_), .A2(n10043), .ZN(n9100) );
  INV_X1 U18305 ( .A(a_30_), .ZN(n10043) );
  NOR2_X1 U18306 ( .A1(n10044), .A2(b_31_), .ZN(n9082) );
  INV_X1 U18307 ( .A(a_31_), .ZN(n10044) );
  NAND2_X1 U18308 ( .A1(a_30_), .A2(n9080), .ZN(n9078) );
  NAND2_X1 U18309 ( .A1(a_28_), .A2(n10786), .ZN(n9157) );
  NAND2_X1 U18310 ( .A1(b_28_), .A2(n9136), .ZN(n9158) );
  NAND2_X1 U18311 ( .A1(a_27_), .A2(n11041), .ZN(n9195) );
  NAND2_X1 U18312 ( .A1(b_27_), .A2(n11274), .ZN(n9196) );
  INV_X1 U18313 ( .A(a_27_), .ZN(n11274) );
  NAND2_X1 U18314 ( .A1(b_24_), .A2(n10050), .ZN(n9280) );
  INV_X1 U18315 ( .A(a_24_), .ZN(n10050) );
  NAND2_X1 U18316 ( .A1(a_24_), .A2(n10049), .ZN(n9281) );
  INV_X1 U18317 ( .A(n9092), .ZN(n9065) );
  INV_X1 U18318 ( .A(operation_1_), .ZN(n9979) );
endmodule

