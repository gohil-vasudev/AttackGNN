module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n445_, new_n236_, new_n238_, new_n479_, new_n250_, new_n288_, new_n421_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n186_, new_n365_, new_n339_, new_n197_, new_n386_, new_n401_, new_n389_, new_n246_, new_n170_, new_n266_, new_n367_, new_n173_, new_n220_, new_n419_, new_n214_, new_n451_, new_n489_, new_n114_, new_n188_, new_n240_, new_n413_, new_n211_, new_n123_, new_n127_, new_n342_, new_n462_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n427_, new_n234_, new_n393_, new_n418_, new_n292_, new_n215_, new_n152_, new_n157_, new_n153_, new_n133_, new_n257_, new_n212_, new_n364_, new_n449_, new_n484_, new_n272_, new_n282_, new_n201_, new_n192_, new_n414_, new_n110_, new_n315_, new_n124_, new_n326_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n248_, new_n350_, new_n117_, new_n167_, new_n385_, new_n461_, new_n297_, new_n361_, new_n150_, new_n108_, new_n137_, new_n183_, new_n463_, new_n303_, new_n351_, new_n325_, new_n180_, new_n318_, new_n321_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n423_, new_n205_, new_n498_, new_n141_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n256_, new_n381_, new_n388_, new_n194_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n314_, new_n118_, new_n363_, new_n165_, new_n441_, new_n477_, new_n216_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n395_, new_n383_, new_n343_, new_n210_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n187_, new_n311_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n349_, new_n244_, new_n172_, new_n488_, new_n277_, new_n402_, new_n286_, new_n335_, new_n347_, new_n346_, new_n198_, new_n438_, new_n208_, new_n179_, new_n436_, new_n397_, new_n399_, new_n233_, new_n469_, new_n391_, new_n178_, new_n295_, new_n359_, new_n132_, new_n166_, new_n162_, new_n457_, new_n161_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n155_, new_n410_, new_n113_, new_n371_, new_n202_, new_n296_, new_n308_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n291_, new_n261_, new_n309_, new_n323_, new_n259_, new_n362_, new_n227_, new_n416_, new_n222_, new_n400_, new_n328_, new_n460_, new_n130_, new_n471_, new_n268_, new_n374_, new_n376_, new_n380_, new_n138_, new_n310_, new_n144_, new_n275_, new_n352_, new_n126_, new_n177_, new_n493_, new_n264_, new_n379_, new_n273_, new_n224_, new_n270_, new_n143_, new_n125_, new_n145_, new_n253_, new_n403_, new_n475_, new_n237_, new_n149_, new_n260_, new_n251_, new_n189_, new_n300_, new_n106_, new_n411_, new_n107_, new_n182_, new_n407_, new_n480_, new_n151_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n428_, new_n199_, new_n146_, new_n302_, new_n191_, new_n225_, new_n387_, new_n476_, new_n112_, new_n121_, new_n415_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n154_, new_n131_, new_n255_, new_n459_, new_n174_, new_n468_, new_n354_, new_n392_, new_n340_, new_n147_, new_n285_, new_n502_, new_n209_, new_n337_, new_n203_, new_n316_, new_n417_, new_n332_, new_n453_, new_n163_, new_n148_, new_n122_, new_n111_, new_n252_, new_n160_, new_n312_, new_n242_, new_n115_, new_n307_, new_n190_, new_n408_, new_n213_, new_n134_, new_n433_, new_n435_, new_n109_, new_n265_, new_n370_, new_n278_, new_n304_, new_n217_, new_n269_, new_n129_, new_n412_, new_n327_, new_n495_, new_n431_, new_n196_, new_n319_, new_n338_, new_n336_, new_n377_, new_n247_, new_n330_, new_n375_, new_n294_, new_n195_, new_n357_, new_n320_, new_n245_, new_n467_, new_n404_, new_n193_, new_n128_, new_n358_, new_n348_, new_n159_, new_n322_, new_n228_, new_n289_, new_n425_, new_n175_, new_n226_, new_n185_, new_n373_, new_n171_, new_n434_, new_n200_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n168_, new_n279_, new_n455_, new_n120_, new_n406_, new_n356_, new_n229_, new_n464_, new_n204_, new_n181_, new_n135_, new_n405_;

not g000 ( new_n106_, N1 );
xnor g001 ( new_n107_, N89, N93 );
xnor g002 ( new_n108_, N81, N85 );
xor g003 ( new_n109_, new_n107_, new_n108_ );
xnor g004 ( new_n110_, N73, N77 );
xor g005 ( new_n111_, N65, N69 );
xnor g006 ( new_n112_, new_n111_, new_n110_ );
nand g007 ( new_n113_, new_n109_, new_n112_ );
xnor g008 ( new_n114_, new_n107_, new_n108_ );
xnor g009 ( new_n115_, N65, N69 );
xnor g010 ( new_n116_, new_n110_, new_n115_ );
nand g011 ( new_n117_, new_n114_, new_n116_ );
nand g012 ( new_n118_, new_n113_, new_n117_ );
nand g013 ( new_n119_, new_n118_, N129, N137 );
nand g014 ( new_n120_, N129, N137 );
nand g015 ( new_n121_, new_n113_, new_n117_, new_n120_ );
nand g016 ( new_n122_, new_n119_, new_n121_ );
xnor g017 ( new_n123_, N1, N17 );
xnor g018 ( new_n124_, N33, N49 );
xnor g019 ( new_n125_, new_n123_, new_n124_ );
xnor g020 ( new_n126_, new_n122_, new_n125_ );
not g021 ( new_n127_, keyIn_0_13 );
not g022 ( new_n128_, keyIn_0_11 );
not g023 ( new_n129_, keyIn_0_9 );
not g024 ( new_n130_, keyIn_0_2 );
not g025 ( new_n131_, N37 );
nand g026 ( new_n132_, new_n131_, N33 );
not g027 ( new_n133_, N33 );
nand g028 ( new_n134_, new_n133_, N37 );
nand g029 ( new_n135_, new_n132_, new_n134_ );
nand g030 ( new_n136_, new_n135_, new_n130_ );
nand g031 ( new_n137_, new_n132_, new_n134_, keyIn_0_2 );
not g032 ( new_n138_, keyIn_0_3 );
not g033 ( new_n139_, N45 );
nand g034 ( new_n140_, new_n139_, N41 );
not g035 ( new_n141_, N41 );
nand g036 ( new_n142_, new_n141_, N45 );
nand g037 ( new_n143_, new_n140_, new_n142_ );
nand g038 ( new_n144_, new_n143_, new_n138_ );
nand g039 ( new_n145_, new_n140_, new_n142_, keyIn_0_3 );
nand g040 ( new_n146_, new_n136_, new_n144_, new_n137_, new_n145_ );
nand g041 ( new_n147_, new_n136_, new_n137_ );
nand g042 ( new_n148_, new_n144_, new_n145_ );
nand g043 ( new_n149_, new_n147_, new_n148_ );
nand g044 ( new_n150_, new_n149_, new_n146_ );
nand g045 ( new_n151_, new_n150_, keyIn_0_7 );
not g046 ( new_n152_, keyIn_0_7 );
nand g047 ( new_n153_, new_n149_, new_n152_, new_n146_ );
not g048 ( new_n154_, keyIn_0_8 );
not g049 ( new_n155_, N53 );
nand g050 ( new_n156_, new_n155_, N49 );
not g051 ( new_n157_, N49 );
nand g052 ( new_n158_, new_n157_, N53 );
nand g053 ( new_n159_, new_n156_, new_n158_ );
nand g054 ( new_n160_, new_n159_, keyIn_0_4 );
not g055 ( new_n161_, keyIn_0_4 );
nand g056 ( new_n162_, new_n156_, new_n158_, new_n161_ );
not g057 ( new_n163_, keyIn_0_5 );
not g058 ( new_n164_, N61 );
nand g059 ( new_n165_, new_n164_, N57 );
not g060 ( new_n166_, N57 );
nand g061 ( new_n167_, new_n166_, N61 );
nand g062 ( new_n168_, new_n165_, new_n167_ );
nand g063 ( new_n169_, new_n168_, new_n163_ );
nand g064 ( new_n170_, new_n165_, new_n167_, keyIn_0_5 );
nand g065 ( new_n171_, new_n160_, new_n169_, new_n162_, new_n170_ );
nand g066 ( new_n172_, new_n160_, new_n162_ );
nand g067 ( new_n173_, new_n169_, new_n170_ );
nand g068 ( new_n174_, new_n172_, new_n173_ );
nand g069 ( new_n175_, new_n174_, new_n154_, new_n171_ );
nand g070 ( new_n176_, new_n174_, new_n171_ );
nand g071 ( new_n177_, new_n176_, keyIn_0_8 );
nand g072 ( new_n178_, new_n177_, new_n175_ );
nand g073 ( new_n179_, new_n178_, new_n151_, new_n153_ );
nand g074 ( new_n180_, new_n151_, new_n153_ );
nand g075 ( new_n181_, new_n180_, new_n175_, new_n177_ );
nand g076 ( new_n182_, new_n179_, new_n181_ );
nand g077 ( new_n183_, new_n182_, new_n129_ );
nand g078 ( new_n184_, new_n179_, new_n181_, keyIn_0_9 );
nand g079 ( new_n185_, new_n183_, new_n184_ );
nand g080 ( new_n186_, N134, N137 );
nand g081 ( new_n187_, new_n185_, new_n186_ );
nand g082 ( new_n188_, new_n183_, N134, N137, new_n184_ );
nand g083 ( new_n189_, new_n187_, new_n188_ );
nand g084 ( new_n190_, new_n189_, new_n128_ );
nand g085 ( new_n191_, new_n187_, keyIn_0_11, new_n188_ );
nand g086 ( new_n192_, new_n190_, new_n191_ );
xnor g087 ( new_n193_, N69, N85 );
xnor g088 ( new_n194_, N101, N117 );
xnor g089 ( new_n195_, new_n193_, new_n194_ );
nand g090 ( new_n196_, new_n192_, new_n195_ );
not g091 ( new_n197_, new_n195_ );
nand g092 ( new_n198_, new_n190_, new_n191_, new_n197_ );
nand g093 ( new_n199_, new_n196_, new_n198_ );
nand g094 ( new_n200_, new_n199_, new_n127_ );
nand g095 ( new_n201_, new_n196_, keyIn_0_13, new_n198_ );
nand g096 ( new_n202_, new_n200_, keyIn_0_15, new_n201_ );
not g097 ( new_n203_, keyIn_0_15 );
nand g098 ( new_n204_, new_n200_, new_n201_ );
nand g099 ( new_n205_, new_n204_, new_n203_ );
nand g100 ( new_n206_, new_n205_, new_n202_ );
not g101 ( new_n207_, keyIn_0_14 );
not g102 ( new_n208_, keyIn_0_10 );
not g103 ( new_n209_, keyIn_0_0 );
not g104 ( new_n210_, N5 );
nand g105 ( new_n211_, new_n210_, N1 );
nand g106 ( new_n212_, new_n106_, N5 );
nand g107 ( new_n213_, new_n211_, new_n212_ );
nand g108 ( new_n214_, new_n213_, new_n209_ );
nand g109 ( new_n215_, new_n211_, new_n212_, keyIn_0_0 );
not g110 ( new_n216_, N13 );
nand g111 ( new_n217_, new_n216_, N9 );
not g112 ( new_n218_, N9 );
nand g113 ( new_n219_, new_n218_, N13 );
nand g114 ( new_n220_, new_n217_, new_n219_ );
nand g115 ( new_n221_, new_n220_, keyIn_0_1 );
not g116 ( new_n222_, keyIn_0_1 );
nand g117 ( new_n223_, new_n217_, new_n219_, new_n222_ );
nand g118 ( new_n224_, new_n214_, new_n221_, new_n215_, new_n223_ );
nand g119 ( new_n225_, new_n214_, new_n215_ );
nand g120 ( new_n226_, new_n221_, new_n223_ );
nand g121 ( new_n227_, new_n225_, new_n226_ );
nand g122 ( new_n228_, new_n227_, keyIn_0_6, new_n224_ );
not g123 ( new_n229_, keyIn_0_6 );
nand g124 ( new_n230_, new_n227_, new_n224_ );
nand g125 ( new_n231_, new_n230_, new_n229_ );
nand g126 ( new_n232_, new_n231_, new_n228_ );
nand g127 ( new_n233_, new_n232_, new_n151_, new_n153_ );
nand g128 ( new_n234_, new_n180_, new_n228_, new_n231_ );
nand g129 ( new_n235_, new_n233_, new_n234_ );
nand g130 ( new_n236_, new_n235_, new_n208_ );
nand g131 ( new_n237_, new_n233_, new_n234_, keyIn_0_10 );
nand g132 ( new_n238_, new_n236_, new_n237_ );
nand g133 ( new_n239_, N135, N137 );
not g134 ( new_n240_, new_n239_ );
nand g135 ( new_n241_, new_n238_, new_n240_ );
nand g136 ( new_n242_, new_n236_, new_n237_, new_n239_ );
nand g137 ( new_n243_, new_n241_, keyIn_0_12, new_n242_ );
not g138 ( new_n244_, keyIn_0_12 );
nand g139 ( new_n245_, new_n241_, new_n242_ );
nand g140 ( new_n246_, new_n245_, new_n244_ );
nand g141 ( new_n247_, new_n246_, new_n243_ );
xnor g142 ( new_n248_, N73, N89 );
xnor g143 ( new_n249_, N105, N121 );
xnor g144 ( new_n250_, new_n248_, new_n249_ );
nand g145 ( new_n251_, new_n247_, new_n250_ );
not g146 ( new_n252_, new_n250_ );
nand g147 ( new_n253_, new_n246_, new_n243_, new_n252_ );
nand g148 ( new_n254_, new_n251_, new_n207_, new_n253_ );
nand g149 ( new_n255_, new_n251_, new_n253_ );
nand g150 ( new_n256_, new_n255_, keyIn_0_14 );
nand g151 ( new_n257_, new_n256_, new_n254_ );
not g152 ( new_n258_, new_n125_ );
xnor g153 ( new_n259_, new_n122_, new_n258_ );
xnor g154 ( new_n260_, N97, N101 );
xnor g155 ( new_n261_, N105, N109 );
xor g156 ( new_n262_, new_n260_, new_n261_ );
xnor g157 ( new_n263_, N121, N125 );
xnor g158 ( new_n264_, N113, N117 );
xor g159 ( new_n265_, new_n263_, new_n264_ );
nand g160 ( new_n266_, new_n262_, new_n265_ );
xnor g161 ( new_n267_, new_n260_, new_n261_ );
xnor g162 ( new_n268_, new_n263_, new_n264_ );
nand g163 ( new_n269_, new_n267_, new_n268_ );
nand g164 ( new_n270_, N130, N137 );
nand g165 ( new_n271_, new_n266_, new_n269_, new_n270_ );
nand g166 ( new_n272_, new_n266_, new_n269_ );
nand g167 ( new_n273_, new_n272_, N130, N137 );
nand g168 ( new_n274_, new_n273_, new_n271_ );
xnor g169 ( new_n275_, N5, N21 );
xnor g170 ( new_n276_, N37, N53 );
xnor g171 ( new_n277_, new_n275_, new_n276_ );
xnor g172 ( new_n278_, new_n274_, new_n277_ );
nand g173 ( new_n279_, new_n262_, new_n112_ );
nand g174 ( new_n280_, new_n116_, new_n267_ );
nand g175 ( new_n281_, N131, N137 );
nand g176 ( new_n282_, new_n279_, new_n280_, new_n281_ );
nand g177 ( new_n283_, new_n279_, new_n280_ );
nand g178 ( new_n284_, new_n283_, N131, N137 );
nand g179 ( new_n285_, new_n284_, new_n282_ );
xnor g180 ( new_n286_, N9, N25 );
xnor g181 ( new_n287_, N41, N57 );
xnor g182 ( new_n288_, new_n286_, new_n287_ );
not g183 ( new_n289_, new_n288_ );
xnor g184 ( new_n290_, new_n285_, new_n289_ );
nand g185 ( new_n291_, new_n278_, new_n259_, new_n290_ );
not g186 ( new_n292_, new_n277_ );
xnor g187 ( new_n293_, new_n274_, new_n292_ );
nand g188 ( new_n294_, new_n293_, new_n290_, new_n126_ );
nand g189 ( new_n295_, new_n291_, new_n294_ );
xnor g190 ( new_n296_, new_n265_, new_n114_ );
nand g191 ( new_n297_, N132, N137 );
nand g192 ( new_n298_, new_n296_, new_n297_ );
xnor g193 ( new_n299_, new_n114_, new_n268_ );
nand g194 ( new_n300_, new_n299_, N132, N137 );
nand g195 ( new_n301_, new_n298_, new_n300_ );
xnor g196 ( new_n302_, N13, N29 );
xnor g197 ( new_n303_, N45, N61 );
xnor g198 ( new_n304_, new_n302_, new_n303_ );
not g199 ( new_n305_, new_n304_ );
xnor g200 ( new_n306_, new_n301_, new_n305_ );
nand g201 ( new_n307_, new_n295_, new_n306_ );
nand g202 ( new_n308_, new_n298_, new_n300_, new_n305_ );
nand g203 ( new_n309_, new_n301_, new_n304_ );
nand g204 ( new_n310_, new_n309_, new_n308_ );
nand g205 ( new_n311_, new_n290_, new_n310_ );
xnor g206 ( new_n312_, new_n285_, new_n288_ );
nand g207 ( new_n313_, new_n306_, new_n312_ );
nand g208 ( new_n314_, new_n313_, new_n311_ );
nand g209 ( new_n315_, new_n293_, new_n259_ );
not g210 ( new_n316_, new_n315_ );
nand g211 ( new_n317_, new_n314_, new_n316_ );
nand g212 ( new_n318_, new_n307_, new_n317_ );
nand g213 ( new_n319_, new_n318_, keyIn_0_17 );
not g214 ( new_n320_, keyIn_0_17 );
nand g215 ( new_n321_, new_n307_, new_n317_, new_n320_ );
nand g216 ( new_n322_, new_n319_, new_n321_ );
xnor g217 ( new_n323_, N17, N21 );
xnor g218 ( new_n324_, N25, N29 );
xnor g219 ( new_n325_, new_n323_, new_n324_ );
xor g220 ( new_n326_, new_n178_, new_n325_ );
nand g221 ( new_n327_, N136, N137 );
xnor g222 ( new_n328_, new_n326_, new_n327_ );
xnor g223 ( new_n329_, N77, N93 );
xnor g224 ( new_n330_, N109, N125 );
xnor g225 ( new_n331_, new_n329_, new_n330_ );
xor g226 ( new_n332_, new_n328_, new_n331_ );
nand g227 ( new_n333_, new_n322_, new_n332_ );
not g228 ( new_n334_, new_n333_ );
xor g229 ( new_n335_, new_n232_, new_n325_ );
nand g230 ( new_n336_, N133, N137 );
xnor g231 ( new_n337_, new_n335_, new_n336_ );
xnor g232 ( new_n338_, N65, N81 );
xnor g233 ( new_n339_, N97, N113 );
xnor g234 ( new_n340_, new_n338_, new_n339_ );
xnor g235 ( new_n341_, new_n337_, new_n340_ );
nand g236 ( new_n342_, new_n257_, new_n334_, new_n341_ );
not g237 ( new_n343_, new_n342_ );
nand g238 ( new_n344_, new_n343_, new_n206_ );
nand g239 ( new_n345_, new_n344_, keyIn_0_18 );
not g240 ( new_n346_, keyIn_0_18 );
nand g241 ( new_n347_, new_n343_, new_n206_, new_n346_ );
nand g242 ( new_n348_, new_n345_, new_n347_ );
nand g243 ( new_n349_, new_n348_, new_n126_ );
nand g244 ( new_n350_, new_n349_, keyIn_0_20 );
not g245 ( new_n351_, keyIn_0_20 );
nand g246 ( new_n352_, new_n348_, new_n351_, new_n126_ );
nand g247 ( new_n353_, new_n350_, new_n352_ );
nand g248 ( new_n354_, new_n353_, new_n106_ );
nand g249 ( new_n355_, new_n350_, N1, new_n352_ );
nand g250 ( new_n356_, new_n354_, keyIn_0_26, new_n355_ );
not g251 ( new_n357_, keyIn_0_26 );
nand g252 ( new_n358_, new_n354_, new_n355_ );
nand g253 ( new_n359_, new_n358_, new_n357_ );
nand g254 ( N724, new_n359_, new_n356_ );
nand g255 ( new_n361_, new_n348_, new_n278_ );
nand g256 ( new_n362_, new_n361_, keyIn_0_21 );
not g257 ( new_n363_, keyIn_0_21 );
nand g258 ( new_n364_, new_n348_, new_n363_, new_n278_ );
nand g259 ( new_n365_, new_n362_, new_n364_ );
nand g260 ( new_n366_, new_n365_, N5 );
nand g261 ( new_n367_, new_n362_, new_n210_, new_n364_ );
nand g262 ( new_n368_, new_n366_, keyIn_0_27, new_n367_ );
not g263 ( new_n369_, keyIn_0_27 );
nand g264 ( new_n370_, new_n366_, new_n367_ );
nand g265 ( new_n371_, new_n370_, new_n369_ );
nand g266 ( N725, new_n371_, new_n368_ );
not g267 ( new_n373_, keyIn_0_28 );
nand g268 ( new_n374_, new_n348_, new_n312_ );
nand g269 ( new_n375_, new_n374_, keyIn_0_22 );
not g270 ( new_n376_, keyIn_0_22 );
nand g271 ( new_n377_, new_n348_, new_n376_, new_n312_ );
nand g272 ( new_n378_, new_n375_, new_n377_ );
nand g273 ( new_n379_, new_n378_, new_n218_ );
nand g274 ( new_n380_, new_n375_, N9, new_n377_ );
nand g275 ( new_n381_, new_n379_, new_n373_, new_n380_ );
nand g276 ( new_n382_, new_n379_, new_n380_ );
nand g277 ( new_n383_, new_n382_, keyIn_0_28 );
nand g278 ( N726, new_n383_, new_n381_ );
nand g279 ( new_n385_, new_n348_, new_n310_ );
nand g280 ( new_n386_, new_n385_, keyIn_0_23 );
not g281 ( new_n387_, keyIn_0_23 );
nand g282 ( new_n388_, new_n348_, new_n387_, new_n310_ );
nand g283 ( new_n389_, new_n386_, new_n388_ );
nand g284 ( new_n390_, new_n389_, new_n216_ );
nand g285 ( new_n391_, new_n386_, N13, new_n388_ );
nand g286 ( new_n392_, new_n390_, keyIn_0_29, new_n391_ );
not g287 ( new_n393_, keyIn_0_29 );
nand g288 ( new_n394_, new_n390_, new_n391_ );
nand g289 ( new_n395_, new_n394_, new_n393_ );
nand g290 ( N727, new_n395_, new_n392_ );
not g291 ( new_n397_, new_n257_ );
nand g292 ( new_n398_, new_n204_, new_n341_ );
not g293 ( new_n399_, new_n398_ );
not g294 ( new_n400_, new_n332_ );
nand g295 ( new_n401_, new_n322_, new_n400_ );
not g296 ( new_n402_, new_n401_ );
nand g297 ( new_n403_, new_n399_, keyIn_0_19, new_n397_, new_n402_ );
not g298 ( new_n404_, keyIn_0_19 );
nand g299 ( new_n405_, new_n399_, new_n397_, new_n402_ );
nand g300 ( new_n406_, new_n405_, new_n404_ );
nand g301 ( new_n407_, new_n406_, new_n403_ );
nand g302 ( new_n408_, new_n407_, new_n126_ );
xnor g303 ( N728, new_n408_, N17 );
not g304 ( new_n410_, N21 );
nand g305 ( new_n411_, new_n407_, new_n278_ );
nand g306 ( new_n412_, new_n411_, keyIn_0_24 );
not g307 ( new_n413_, keyIn_0_24 );
nand g308 ( new_n414_, new_n407_, new_n413_, new_n278_ );
nand g309 ( new_n415_, new_n412_, new_n410_, new_n414_ );
nand g310 ( new_n416_, new_n412_, new_n414_ );
nand g311 ( new_n417_, new_n416_, N21 );
nand g312 ( new_n418_, new_n417_, keyIn_0_30, new_n415_ );
not g313 ( new_n419_, keyIn_0_30 );
nand g314 ( new_n420_, new_n417_, new_n415_ );
nand g315 ( new_n421_, new_n420_, new_n419_ );
nand g316 ( N729, new_n421_, new_n418_ );
nand g317 ( new_n423_, new_n407_, new_n312_ );
xnor g318 ( N730, new_n423_, N25 );
not g319 ( new_n425_, keyIn_0_25 );
nand g320 ( new_n426_, new_n407_, new_n310_ );
nand g321 ( new_n427_, new_n426_, new_n425_ );
nand g322 ( new_n428_, new_n407_, keyIn_0_25, new_n310_ );
nand g323 ( new_n429_, new_n427_, N29, new_n428_ );
not g324 ( new_n430_, N29 );
nand g325 ( new_n431_, new_n427_, new_n428_ );
nand g326 ( new_n432_, new_n431_, new_n430_ );
nand g327 ( new_n433_, new_n432_, keyIn_0_31, new_n429_ );
not g328 ( new_n434_, keyIn_0_31 );
nand g329 ( new_n435_, new_n432_, new_n429_ );
nand g330 ( new_n436_, new_n435_, new_n434_ );
nand g331 ( N731, new_n436_, new_n433_ );
nor g332 ( new_n438_, new_n397_, new_n204_, new_n333_, new_n341_ );
nand g333 ( new_n439_, new_n438_, new_n126_ );
xnor g334 ( N732, new_n439_, N33 );
nand g335 ( new_n441_, new_n438_, new_n278_ );
xnor g336 ( N733, new_n441_, N37 );
nand g337 ( new_n443_, new_n438_, new_n312_ );
xnor g338 ( N734, new_n443_, N41 );
nand g339 ( new_n445_, new_n438_, new_n310_ );
xnor g340 ( N735, new_n445_, N45 );
not g341 ( new_n447_, new_n204_ );
not g342 ( new_n448_, new_n341_ );
nand g343 ( new_n449_, new_n447_, new_n397_, new_n448_ );
nor g344 ( new_n450_, new_n449_, new_n401_ );
nand g345 ( new_n451_, new_n450_, new_n126_ );
xnor g346 ( N736, new_n451_, N49 );
nand g347 ( new_n453_, new_n450_, new_n278_ );
xnor g348 ( N737, new_n453_, N53 );
nand g349 ( new_n455_, new_n450_, new_n312_ );
xnor g350 ( N738, new_n455_, N57 );
nand g351 ( new_n457_, new_n450_, new_n310_ );
xnor g352 ( N739, new_n457_, N61 );
not g353 ( new_n459_, keyIn_0_16 );
nand g354 ( new_n460_, new_n397_, new_n459_ );
nand g355 ( new_n461_, new_n257_, keyIn_0_16 );
nand g356 ( new_n462_, new_n399_, new_n460_, new_n461_ );
nand g357 ( new_n463_, new_n462_, new_n449_ );
nand g358 ( new_n464_, new_n463_, new_n332_ );
xnor g359 ( new_n465_, new_n257_, new_n332_ );
nand g360 ( new_n466_, new_n465_, new_n204_, new_n448_ );
nand g361 ( new_n467_, new_n464_, new_n466_ );
nor g362 ( new_n468_, new_n313_, new_n259_, new_n278_ );
nand g363 ( new_n469_, new_n467_, new_n341_, new_n468_ );
xnor g364 ( N740, new_n469_, N65 );
nand g365 ( new_n471_, new_n467_, new_n447_, new_n468_ );
xnor g366 ( N741, new_n471_, N69 );
nand g367 ( new_n473_, new_n467_, new_n257_, new_n468_ );
xnor g368 ( N742, new_n473_, N73 );
not g369 ( new_n475_, new_n467_ );
nor g370 ( new_n476_, new_n475_, new_n332_ );
nand g371 ( new_n477_, new_n476_, new_n468_ );
xnor g372 ( N743, new_n477_, N77 );
nor g373 ( new_n479_, new_n294_, new_n306_ );
nand g374 ( new_n480_, new_n467_, new_n341_, new_n479_ );
xnor g375 ( N744, new_n480_, N81 );
nand g376 ( new_n482_, new_n467_, new_n447_, new_n479_ );
xnor g377 ( N745, new_n482_, N85 );
nand g378 ( new_n484_, new_n467_, new_n257_, new_n479_ );
xnor g379 ( N746, new_n484_, N89 );
nand g380 ( new_n486_, new_n476_, new_n479_ );
xnor g381 ( N747, new_n486_, N93 );
nor g382 ( new_n488_, new_n313_, new_n126_, new_n293_ );
nand g383 ( new_n489_, new_n467_, new_n341_, new_n488_ );
xnor g384 ( N748, new_n489_, N97 );
nand g385 ( new_n491_, new_n467_, new_n447_, new_n488_ );
xnor g386 ( N749, new_n491_, N101 );
nand g387 ( new_n493_, new_n467_, new_n257_, new_n488_ );
xnor g388 ( N750, new_n493_, N105 );
nand g389 ( new_n495_, new_n476_, new_n488_ );
xnor g390 ( N751, new_n495_, N109 );
nor g391 ( new_n497_, new_n291_, new_n306_ );
nand g392 ( new_n498_, new_n467_, new_n341_, new_n497_ );
xnor g393 ( N752, new_n498_, N113 );
nand g394 ( new_n500_, new_n467_, new_n447_, new_n497_ );
xnor g395 ( N753, new_n500_, N117 );
nand g396 ( new_n502_, new_n467_, new_n257_, new_n497_ );
xnor g397 ( N754, new_n502_, N121 );
nand g398 ( new_n504_, new_n476_, new_n497_ );
xnor g399 ( N755, new_n504_, N125 );
endmodule