module add_mul_combine_8_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, Result_mul_0_, 
        Result_mul_1_, Result_mul_2_, Result_mul_3_, Result_mul_4_, 
        Result_mul_5_, Result_mul_6_, Result_mul_7_, Result_mul_8_, 
        Result_mul_9_, Result_mul_10_, Result_mul_11_, Result_mul_12_, 
        Result_mul_13_, Result_mul_14_, Result_mul_15_, Result_add_0_, 
        Result_add_1_, Result_add_2_, Result_add_3_, Result_add_4_, 
        Result_add_5_, Result_add_6_, Result_add_7_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_,
         b_4_, b_5_, b_6_, b_7_;
  output Result_mul_0_, Result_mul_1_, Result_mul_2_, Result_mul_3_,
         Result_mul_4_, Result_mul_5_, Result_mul_6_, Result_mul_7_,
         Result_mul_8_, Result_mul_9_, Result_mul_10_, Result_mul_11_,
         Result_mul_12_, Result_mul_13_, Result_mul_14_, Result_mul_15_,
         Result_add_0_, Result_add_1_, Result_add_2_, Result_add_3_,
         Result_add_4_, Result_add_5_, Result_add_6_, Result_add_7_;
  wire   n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594;

  OR2_X1 U827 ( .A1(n803), .A2(n804), .ZN(Result_mul_9_) );
  AND2_X1 U828 ( .A1(n805), .A2(n806), .ZN(n804) );
  INV_X1 U829 ( .A(n807), .ZN(n803) );
  OR2_X1 U830 ( .A1(n806), .A2(n805), .ZN(n807) );
  OR2_X1 U831 ( .A1(n808), .A2(n809), .ZN(n805) );
  AND2_X1 U832 ( .A1(n810), .A2(n811), .ZN(n809) );
  AND2_X1 U833 ( .A1(n812), .A2(n813), .ZN(n808) );
  INV_X1 U834 ( .A(n811), .ZN(n812) );
  OR2_X1 U835 ( .A1(n814), .A2(n815), .ZN(Result_mul_8_) );
  AND2_X1 U836 ( .A1(n816), .A2(n817), .ZN(n815) );
  INV_X1 U837 ( .A(n818), .ZN(n814) );
  OR2_X1 U838 ( .A1(n817), .A2(n816), .ZN(n818) );
  OR2_X1 U839 ( .A1(n819), .A2(n820), .ZN(n816) );
  AND2_X1 U840 ( .A1(n821), .A2(n822), .ZN(n820) );
  AND2_X1 U841 ( .A1(n823), .A2(n824), .ZN(n819) );
  INV_X1 U842 ( .A(n822), .ZN(n823) );
  AND2_X1 U843 ( .A1(n825), .A2(n826), .ZN(Result_mul_7_) );
  OR2_X1 U844 ( .A1(n827), .A2(n828), .ZN(n826) );
  INV_X1 U845 ( .A(n829), .ZN(n828) );
  OR2_X1 U846 ( .A1(n830), .A2(n829), .ZN(n825) );
  AND2_X1 U847 ( .A1(n831), .A2(n832), .ZN(Result_mul_6_) );
  INV_X1 U848 ( .A(n833), .ZN(n832) );
  OR2_X1 U849 ( .A1(n834), .A2(n835), .ZN(n831) );
  AND2_X1 U850 ( .A1(n830), .A2(n829), .ZN(n834) );
  OR2_X1 U851 ( .A1(n836), .A2(n837), .ZN(Result_mul_5_) );
  INV_X1 U852 ( .A(n838), .ZN(n837) );
  OR2_X1 U853 ( .A1(n839), .A2(n833), .ZN(n838) );
  AND2_X1 U854 ( .A1(n833), .A2(n839), .ZN(n836) );
  OR2_X1 U855 ( .A1(n840), .A2(n841), .ZN(n839) );
  AND2_X1 U856 ( .A1(n842), .A2(n843), .ZN(n840) );
  AND2_X1 U857 ( .A1(n844), .A2(n845), .ZN(Result_mul_4_) );
  INV_X1 U858 ( .A(n846), .ZN(n844) );
  AND2_X1 U859 ( .A1(n847), .A2(n848), .ZN(n846) );
  OR2_X1 U860 ( .A1(n849), .A2(n850), .ZN(Result_mul_3_) );
  INV_X1 U861 ( .A(n851), .ZN(n850) );
  OR2_X1 U862 ( .A1(n852), .A2(n853), .ZN(n851) );
  AND2_X1 U863 ( .A1(n853), .A2(n852), .ZN(n849) );
  OR2_X1 U864 ( .A1(n854), .A2(n855), .ZN(n852) );
  AND2_X1 U865 ( .A1(n856), .A2(n857), .ZN(n854) );
  OR2_X1 U866 ( .A1(n858), .A2(n859), .ZN(Result_mul_2_) );
  AND2_X1 U867 ( .A1(n860), .A2(n861), .ZN(n859) );
  OR2_X1 U868 ( .A1(n862), .A2(n863), .ZN(n860) );
  AND2_X1 U869 ( .A1(n864), .A2(n865), .ZN(n863) );
  INV_X1 U870 ( .A(n866), .ZN(n864) );
  AND2_X1 U871 ( .A1(n867), .A2(n866), .ZN(n862) );
  AND2_X1 U872 ( .A1(n868), .A2(n866), .ZN(n858) );
  OR2_X1 U873 ( .A1(n869), .A2(n870), .ZN(Result_mul_1_) );
  INV_X1 U874 ( .A(n871), .ZN(n870) );
  OR2_X1 U875 ( .A1(n872), .A2(n873), .ZN(n871) );
  AND2_X1 U876 ( .A1(n873), .A2(n872), .ZN(n869) );
  OR2_X1 U877 ( .A1(n874), .A2(n875), .ZN(n872) );
  AND2_X1 U878 ( .A1(n876), .A2(n877), .ZN(n874) );
  INV_X1 U879 ( .A(n878), .ZN(n876) );
  OR2_X1 U880 ( .A1(n879), .A2(n880), .ZN(Result_mul_14_) );
  AND2_X1 U881 ( .A1(n881), .A2(n882), .ZN(n880) );
  INV_X1 U882 ( .A(n883), .ZN(n879) );
  OR2_X1 U883 ( .A1(n882), .A2(n881), .ZN(n883) );
  AND2_X1 U884 ( .A1(a_6_), .A2(b_7_), .ZN(n881) );
  OR2_X1 U885 ( .A1(n884), .A2(n885), .ZN(n882) );
  OR2_X1 U886 ( .A1(n886), .A2(n887), .ZN(Result_mul_13_) );
  AND2_X1 U887 ( .A1(n888), .A2(n889), .ZN(n887) );
  INV_X1 U888 ( .A(n890), .ZN(n886) );
  OR2_X1 U889 ( .A1(n889), .A2(n888), .ZN(n890) );
  OR2_X1 U890 ( .A1(n891), .A2(n892), .ZN(n888) );
  AND2_X1 U891 ( .A1(n893), .A2(n894), .ZN(n892) );
  INV_X1 U892 ( .A(n895), .ZN(n893) );
  AND2_X1 U893 ( .A1(n896), .A2(n895), .ZN(n891) );
  OR2_X1 U894 ( .A1(n897), .A2(n898), .ZN(Result_mul_12_) );
  AND2_X1 U895 ( .A1(n899), .A2(n900), .ZN(n898) );
  INV_X1 U896 ( .A(n901), .ZN(n897) );
  OR2_X1 U897 ( .A1(n900), .A2(n899), .ZN(n901) );
  OR2_X1 U898 ( .A1(n902), .A2(n903), .ZN(n899) );
  AND2_X1 U899 ( .A1(n904), .A2(n905), .ZN(n903) );
  AND2_X1 U900 ( .A1(n906), .A2(n907), .ZN(n902) );
  INV_X1 U901 ( .A(n905), .ZN(n906) );
  AND2_X1 U902 ( .A1(n908), .A2(n909), .ZN(Result_mul_11_) );
  INV_X1 U903 ( .A(n910), .ZN(n909) );
  AND2_X1 U904 ( .A1(n911), .A2(n912), .ZN(n910) );
  OR2_X1 U905 ( .A1(n912), .A2(n911), .ZN(n908) );
  AND2_X1 U906 ( .A1(n913), .A2(n914), .ZN(n911) );
  INV_X1 U907 ( .A(n915), .ZN(n914) );
  AND2_X1 U908 ( .A1(n916), .A2(n917), .ZN(n915) );
  OR2_X1 U909 ( .A1(n917), .A2(n916), .ZN(n913) );
  INV_X1 U910 ( .A(n918), .ZN(n916) );
  OR2_X1 U911 ( .A1(n919), .A2(n920), .ZN(Result_mul_10_) );
  AND2_X1 U912 ( .A1(n921), .A2(n922), .ZN(n920) );
  INV_X1 U913 ( .A(n923), .ZN(n919) );
  OR2_X1 U914 ( .A1(n922), .A2(n921), .ZN(n923) );
  OR2_X1 U915 ( .A1(n924), .A2(n925), .ZN(n921) );
  AND2_X1 U916 ( .A1(n926), .A2(n927), .ZN(n925) );
  INV_X1 U917 ( .A(n928), .ZN(n924) );
  OR2_X1 U918 ( .A1(n927), .A2(n926), .ZN(n928) );
  INV_X1 U919 ( .A(n929), .ZN(n926) );
  OR3_X1 U920 ( .A1(n875), .A2(n930), .A3(n931), .ZN(Result_mul_0_) );
  AND2_X1 U921 ( .A1(n932), .A2(a_0_), .ZN(n931) );
  INV_X1 U922 ( .A(n933), .ZN(n932) );
  AND2_X1 U923 ( .A1(n873), .A2(n878), .ZN(n930) );
  INV_X1 U924 ( .A(n934), .ZN(n873) );
  OR2_X1 U925 ( .A1(n935), .A2(n866), .ZN(n934) );
  OR2_X1 U926 ( .A1(n936), .A2(n937), .ZN(n866) );
  AND2_X1 U927 ( .A1(n938), .A2(n939), .ZN(n936) );
  AND2_X1 U928 ( .A1(n861), .A2(n865), .ZN(n935) );
  INV_X1 U929 ( .A(n868), .ZN(n861) );
  OR2_X1 U930 ( .A1(n940), .A2(n855), .ZN(n868) );
  AND2_X1 U931 ( .A1(n941), .A2(n942), .ZN(n855) );
  AND2_X1 U932 ( .A1(n853), .A2(n942), .ZN(n940) );
  INV_X1 U933 ( .A(n857), .ZN(n942) );
  OR2_X1 U934 ( .A1(n867), .A2(n943), .ZN(n857) );
  AND3_X1 U935 ( .A1(n944), .A2(n945), .A3(n946), .ZN(n943) );
  INV_X1 U936 ( .A(n865), .ZN(n867) );
  OR2_X1 U937 ( .A1(n947), .A2(n946), .ZN(n865) );
  OR2_X1 U938 ( .A1(n948), .A2(n949), .ZN(n946) );
  AND2_X1 U939 ( .A1(n950), .A2(n951), .ZN(n949) );
  AND2_X1 U940 ( .A1(n952), .A2(n953), .ZN(n948) );
  OR2_X1 U941 ( .A1(n951), .A2(n950), .ZN(n953) );
  AND2_X1 U942 ( .A1(n944), .A2(n945), .ZN(n947) );
  OR2_X1 U943 ( .A1(n954), .A2(n955), .ZN(n945) );
  INV_X1 U944 ( .A(n956), .ZN(n954) );
  OR2_X1 U945 ( .A1(n957), .A2(n956), .ZN(n944) );
  AND2_X1 U946 ( .A1(n958), .A2(n959), .ZN(n956) );
  INV_X1 U947 ( .A(n960), .ZN(n959) );
  AND2_X1 U948 ( .A1(n961), .A2(n962), .ZN(n960) );
  OR2_X1 U949 ( .A1(n962), .A2(n961), .ZN(n958) );
  INV_X1 U950 ( .A(n963), .ZN(n961) );
  INV_X1 U951 ( .A(n955), .ZN(n957) );
  INV_X1 U952 ( .A(n845), .ZN(n853) );
  OR2_X1 U953 ( .A1(n848), .A2(n847), .ZN(n845) );
  OR2_X1 U954 ( .A1(n964), .A2(n941), .ZN(n847) );
  INV_X1 U955 ( .A(n856), .ZN(n941) );
  OR2_X1 U956 ( .A1(n965), .A2(n966), .ZN(n856) );
  AND2_X1 U957 ( .A1(n965), .A2(n966), .ZN(n964) );
  OR2_X1 U958 ( .A1(n967), .A2(n968), .ZN(n966) );
  AND2_X1 U959 ( .A1(n969), .A2(n970), .ZN(n968) );
  AND2_X1 U960 ( .A1(n971), .A2(n972), .ZN(n967) );
  OR2_X1 U961 ( .A1(n970), .A2(n969), .ZN(n972) );
  INV_X1 U962 ( .A(n973), .ZN(n969) );
  AND2_X1 U963 ( .A1(n974), .A2(n975), .ZN(n965) );
  INV_X1 U964 ( .A(n976), .ZN(n975) );
  AND2_X1 U965 ( .A1(n977), .A2(n952), .ZN(n976) );
  OR2_X1 U966 ( .A1(n952), .A2(n977), .ZN(n974) );
  OR2_X1 U967 ( .A1(n978), .A2(n979), .ZN(n977) );
  AND2_X1 U968 ( .A1(n980), .A2(n951), .ZN(n979) );
  INV_X1 U969 ( .A(n981), .ZN(n951) );
  INV_X1 U970 ( .A(n950), .ZN(n980) );
  AND2_X1 U971 ( .A1(n981), .A2(n950), .ZN(n978) );
  OR2_X1 U972 ( .A1(n982), .A2(n983), .ZN(n950) );
  AND2_X1 U973 ( .A1(n984), .A2(n985), .ZN(n983) );
  AND2_X1 U974 ( .A1(n986), .A2(n987), .ZN(n982) );
  OR2_X1 U975 ( .A1(n985), .A2(n984), .ZN(n987) );
  AND2_X1 U976 ( .A1(b_3_), .A2(a_0_), .ZN(n981) );
  AND2_X1 U977 ( .A1(n988), .A2(n989), .ZN(n952) );
  INV_X1 U978 ( .A(n990), .ZN(n989) );
  AND2_X1 U979 ( .A1(n991), .A2(n992), .ZN(n990) );
  OR2_X1 U980 ( .A1(n992), .A2(n991), .ZN(n988) );
  OR2_X1 U981 ( .A1(n993), .A2(n994), .ZN(n991) );
  INV_X1 U982 ( .A(n995), .ZN(n994) );
  OR2_X1 U983 ( .A1(n996), .A2(n997), .ZN(n995) );
  AND2_X1 U984 ( .A1(n997), .A2(n996), .ZN(n993) );
  INV_X1 U985 ( .A(n998), .ZN(n997) );
  AND2_X1 U986 ( .A1(n999), .A2(n1000), .ZN(n848) );
  INV_X1 U987 ( .A(n1001), .ZN(n999) );
  OR2_X1 U988 ( .A1(n1002), .A2(n841), .ZN(n1001) );
  AND3_X1 U989 ( .A1(n1003), .A2(n1004), .A3(n1005), .ZN(n841) );
  AND2_X1 U990 ( .A1(n833), .A2(n1005), .ZN(n1002) );
  INV_X1 U991 ( .A(n843), .ZN(n1005) );
  OR2_X1 U992 ( .A1(n1006), .A2(n1007), .ZN(n843) );
  AND3_X1 U993 ( .A1(n1008), .A2(n1009), .A3(n1010), .ZN(n1007) );
  INV_X1 U994 ( .A(n1000), .ZN(n1006) );
  OR2_X1 U995 ( .A1(n1011), .A2(n1010), .ZN(n1000) );
  OR2_X1 U996 ( .A1(n1012), .A2(n1013), .ZN(n1010) );
  AND2_X1 U997 ( .A1(n1014), .A2(n1015), .ZN(n1013) );
  AND2_X1 U998 ( .A1(n1016), .A2(n1017), .ZN(n1012) );
  OR2_X1 U999 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  INV_X1 U1000 ( .A(n1018), .ZN(n1015) );
  AND2_X1 U1001 ( .A1(n1008), .A2(n1009), .ZN(n1011) );
  OR2_X1 U1002 ( .A1(n1019), .A2(n971), .ZN(n1009) );
  OR2_X1 U1003 ( .A1(n1020), .A2(n1021), .ZN(n1008) );
  INV_X1 U1004 ( .A(n1019), .ZN(n1021) );
  OR2_X1 U1005 ( .A1(n1022), .A2(n1023), .ZN(n1019) );
  AND2_X1 U1006 ( .A1(n973), .A2(n970), .ZN(n1023) );
  INV_X1 U1007 ( .A(n1024), .ZN(n1022) );
  OR2_X1 U1008 ( .A1(n970), .A2(n973), .ZN(n1024) );
  AND2_X1 U1009 ( .A1(b_4_), .A2(a_0_), .ZN(n973) );
  OR2_X1 U1010 ( .A1(n1025), .A2(n1026), .ZN(n970) );
  AND2_X1 U1011 ( .A1(n1027), .A2(n1028), .ZN(n1026) );
  AND2_X1 U1012 ( .A1(n1029), .A2(n1030), .ZN(n1025) );
  OR2_X1 U1013 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  INV_X1 U1014 ( .A(n1031), .ZN(n1028) );
  INV_X1 U1015 ( .A(n971), .ZN(n1020) );
  AND2_X1 U1016 ( .A1(n1032), .A2(n1033), .ZN(n971) );
  INV_X1 U1017 ( .A(n1034), .ZN(n1033) );
  AND2_X1 U1018 ( .A1(n1035), .A2(n986), .ZN(n1034) );
  OR2_X1 U1019 ( .A1(n986), .A2(n1035), .ZN(n1032) );
  OR2_X1 U1020 ( .A1(n1036), .A2(n1037), .ZN(n1035) );
  AND2_X1 U1021 ( .A1(n1038), .A2(n985), .ZN(n1037) );
  INV_X1 U1022 ( .A(n1039), .ZN(n985) );
  INV_X1 U1023 ( .A(n984), .ZN(n1038) );
  AND2_X1 U1024 ( .A1(n1039), .A2(n984), .ZN(n1036) );
  OR2_X1 U1025 ( .A1(n1040), .A2(n1041), .ZN(n984) );
  AND2_X1 U1026 ( .A1(n1042), .A2(n1043), .ZN(n1041) );
  AND2_X1 U1027 ( .A1(n1044), .A2(n1045), .ZN(n1040) );
  OR2_X1 U1028 ( .A1(n1043), .A2(n1042), .ZN(n1045) );
  INV_X1 U1029 ( .A(n1046), .ZN(n1042) );
  AND2_X1 U1030 ( .A1(b_3_), .A2(a_1_), .ZN(n1039) );
  AND2_X1 U1031 ( .A1(n1047), .A2(n1048), .ZN(n986) );
  INV_X1 U1032 ( .A(n1049), .ZN(n1048) );
  AND2_X1 U1033 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
  OR2_X1 U1034 ( .A1(n1051), .A2(n1050), .ZN(n1047) );
  OR2_X1 U1035 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
  INV_X1 U1036 ( .A(n1054), .ZN(n1053) );
  OR2_X1 U1037 ( .A1(n1055), .A2(n1056), .ZN(n1054) );
  AND2_X1 U1038 ( .A1(n1056), .A2(n1055), .ZN(n1052) );
  AND3_X1 U1039 ( .A1(n830), .A2(n829), .A3(n835), .ZN(n833) );
  AND2_X1 U1040 ( .A1(n842), .A2(n1057), .ZN(n835) );
  OR2_X1 U1041 ( .A1(n1004), .A2(n1003), .ZN(n1057) );
  INV_X1 U1042 ( .A(n1058), .ZN(n1003) );
  OR2_X1 U1043 ( .A1(n1059), .A2(n1058), .ZN(n842) );
  OR2_X1 U1044 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
  AND2_X1 U1045 ( .A1(n1062), .A2(n1063), .ZN(n1061) );
  AND2_X1 U1046 ( .A1(n1064), .A2(n1065), .ZN(n1060) );
  OR2_X1 U1047 ( .A1(n1063), .A2(n1062), .ZN(n1065) );
  INV_X1 U1048 ( .A(n1066), .ZN(n1062) );
  INV_X1 U1049 ( .A(n1004), .ZN(n1059) );
  AND2_X1 U1050 ( .A1(n1067), .A2(n1068), .ZN(n1004) );
  OR2_X1 U1051 ( .A1(n1069), .A2(n1014), .ZN(n1068) );
  INV_X1 U1052 ( .A(n1070), .ZN(n1067) );
  AND2_X1 U1053 ( .A1(n1014), .A2(n1069), .ZN(n1070) );
  AND2_X1 U1054 ( .A1(n1071), .A2(n1072), .ZN(n1069) );
  INV_X1 U1055 ( .A(n1073), .ZN(n1072) );
  AND2_X1 U1056 ( .A1(n1018), .A2(n1017), .ZN(n1073) );
  OR2_X1 U1057 ( .A1(n1017), .A2(n1018), .ZN(n1071) );
  AND2_X1 U1058 ( .A1(b_5_), .A2(a_0_), .ZN(n1018) );
  OR2_X1 U1059 ( .A1(n1074), .A2(n1075), .ZN(n1017) );
  AND2_X1 U1060 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
  AND2_X1 U1061 ( .A1(n1078), .A2(n1079), .ZN(n1074) );
  OR2_X1 U1062 ( .A1(n1077), .A2(n1076), .ZN(n1079) );
  INV_X1 U1063 ( .A(n1080), .ZN(n1076) );
  OR2_X1 U1064 ( .A1(n1081), .A2(n1082), .ZN(n1014) );
  INV_X1 U1065 ( .A(n1083), .ZN(n1082) );
  OR2_X1 U1066 ( .A1(n1084), .A2(n1027), .ZN(n1083) );
  AND2_X1 U1067 ( .A1(n1027), .A2(n1084), .ZN(n1081) );
  AND2_X1 U1068 ( .A1(n1085), .A2(n1086), .ZN(n1084) );
  INV_X1 U1069 ( .A(n1087), .ZN(n1086) );
  AND2_X1 U1070 ( .A1(n1031), .A2(n1030), .ZN(n1087) );
  OR2_X1 U1071 ( .A1(n1030), .A2(n1031), .ZN(n1085) );
  AND2_X1 U1072 ( .A1(b_4_), .A2(a_1_), .ZN(n1031) );
  OR2_X1 U1073 ( .A1(n1088), .A2(n1089), .ZN(n1030) );
  AND2_X1 U1074 ( .A1(n1090), .A2(n1091), .ZN(n1089) );
  AND2_X1 U1075 ( .A1(n1092), .A2(n1093), .ZN(n1088) );
  OR2_X1 U1076 ( .A1(n1091), .A2(n1090), .ZN(n1093) );
  INV_X1 U1077 ( .A(n1094), .ZN(n1090) );
  OR2_X1 U1078 ( .A1(n1095), .A2(n1096), .ZN(n1027) );
  INV_X1 U1079 ( .A(n1097), .ZN(n1096) );
  OR2_X1 U1080 ( .A1(n1098), .A2(n1044), .ZN(n1097) );
  AND2_X1 U1081 ( .A1(n1044), .A2(n1098), .ZN(n1095) );
  AND2_X1 U1082 ( .A1(n1099), .A2(n1100), .ZN(n1098) );
  INV_X1 U1083 ( .A(n1101), .ZN(n1100) );
  AND2_X1 U1084 ( .A1(n1046), .A2(n1043), .ZN(n1101) );
  OR2_X1 U1085 ( .A1(n1043), .A2(n1046), .ZN(n1099) );
  AND2_X1 U1086 ( .A1(b_3_), .A2(a_2_), .ZN(n1046) );
  OR2_X1 U1087 ( .A1(n1102), .A2(n1103), .ZN(n1043) );
  AND2_X1 U1088 ( .A1(n1104), .A2(n1105), .ZN(n1103) );
  AND2_X1 U1089 ( .A1(n1106), .A2(n1107), .ZN(n1102) );
  OR2_X1 U1090 ( .A1(n1105), .A2(n1104), .ZN(n1106) );
  OR2_X1 U1091 ( .A1(n1108), .A2(n1109), .ZN(n1044) );
  INV_X1 U1092 ( .A(n1110), .ZN(n1109) );
  OR2_X1 U1093 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
  AND2_X1 U1094 ( .A1(n1112), .A2(n1111), .ZN(n1108) );
  AND2_X1 U1095 ( .A1(n1113), .A2(n1114), .ZN(n1111) );
  INV_X1 U1096 ( .A(n1115), .ZN(n1114) );
  AND2_X1 U1097 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
  OR2_X1 U1098 ( .A1(n1117), .A2(n1116), .ZN(n1113) );
  AND2_X1 U1099 ( .A1(n1118), .A2(n1119), .ZN(n829) );
  OR2_X1 U1100 ( .A1(n1120), .A2(n1064), .ZN(n1119) );
  INV_X1 U1101 ( .A(n1121), .ZN(n1118) );
  AND2_X1 U1102 ( .A1(n1064), .A2(n1120), .ZN(n1121) );
  AND2_X1 U1103 ( .A1(n1122), .A2(n1123), .ZN(n1120) );
  INV_X1 U1104 ( .A(n1124), .ZN(n1123) );
  AND2_X1 U1105 ( .A1(n1066), .A2(n1063), .ZN(n1124) );
  OR2_X1 U1106 ( .A1(n1063), .A2(n1066), .ZN(n1122) );
  AND2_X1 U1107 ( .A1(b_6_), .A2(a_0_), .ZN(n1066) );
  OR2_X1 U1108 ( .A1(n1125), .A2(n1126), .ZN(n1063) );
  AND2_X1 U1109 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
  AND2_X1 U1110 ( .A1(n1129), .A2(n1130), .ZN(n1125) );
  OR2_X1 U1111 ( .A1(n1128), .A2(n1127), .ZN(n1130) );
  OR2_X1 U1112 ( .A1(n1131), .A2(n1132), .ZN(n1064) );
  INV_X1 U1113 ( .A(n1133), .ZN(n1132) );
  OR2_X1 U1114 ( .A1(n1134), .A2(n1078), .ZN(n1133) );
  AND2_X1 U1115 ( .A1(n1078), .A2(n1134), .ZN(n1131) );
  AND2_X1 U1116 ( .A1(n1135), .A2(n1136), .ZN(n1134) );
  INV_X1 U1117 ( .A(n1137), .ZN(n1136) );
  AND2_X1 U1118 ( .A1(n1080), .A2(n1077), .ZN(n1137) );
  OR2_X1 U1119 ( .A1(n1077), .A2(n1080), .ZN(n1135) );
  AND2_X1 U1120 ( .A1(b_5_), .A2(a_1_), .ZN(n1080) );
  OR2_X1 U1121 ( .A1(n1138), .A2(n1139), .ZN(n1077) );
  AND2_X1 U1122 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
  AND2_X1 U1123 ( .A1(n1142), .A2(n1143), .ZN(n1138) );
  OR2_X1 U1124 ( .A1(n1141), .A2(n1140), .ZN(n1143) );
  OR2_X1 U1125 ( .A1(n1144), .A2(n1145), .ZN(n1078) );
  INV_X1 U1126 ( .A(n1146), .ZN(n1145) );
  OR2_X1 U1127 ( .A1(n1147), .A2(n1092), .ZN(n1146) );
  AND2_X1 U1128 ( .A1(n1092), .A2(n1147), .ZN(n1144) );
  AND2_X1 U1129 ( .A1(n1148), .A2(n1149), .ZN(n1147) );
  INV_X1 U1130 ( .A(n1150), .ZN(n1149) );
  AND2_X1 U1131 ( .A1(n1094), .A2(n1091), .ZN(n1150) );
  OR2_X1 U1132 ( .A1(n1091), .A2(n1094), .ZN(n1148) );
  AND2_X1 U1133 ( .A1(b_4_), .A2(a_2_), .ZN(n1094) );
  OR2_X1 U1134 ( .A1(n1151), .A2(n1152), .ZN(n1091) );
  AND2_X1 U1135 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
  AND2_X1 U1136 ( .A1(n1155), .A2(n1156), .ZN(n1151) );
  OR2_X1 U1137 ( .A1(n1154), .A2(n1153), .ZN(n1156) );
  INV_X1 U1138 ( .A(n1157), .ZN(n1153) );
  OR2_X1 U1139 ( .A1(n1158), .A2(n1159), .ZN(n1092) );
  INV_X1 U1140 ( .A(n1160), .ZN(n1159) );
  OR2_X1 U1141 ( .A1(n1161), .A2(n1104), .ZN(n1160) );
  AND2_X1 U1142 ( .A1(n1104), .A2(n1161), .ZN(n1158) );
  AND2_X1 U1143 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
  OR2_X1 U1144 ( .A1(n1105), .A2(n1164), .ZN(n1163) );
  INV_X1 U1145 ( .A(n1165), .ZN(n1162) );
  AND2_X1 U1146 ( .A1(n1164), .A2(n1105), .ZN(n1165) );
  OR2_X1 U1147 ( .A1(n1166), .A2(n1167), .ZN(n1105) );
  AND2_X1 U1148 ( .A1(n1168), .A2(n1169), .ZN(n1167) );
  AND2_X1 U1149 ( .A1(n1170), .A2(n1171), .ZN(n1166) );
  OR2_X1 U1150 ( .A1(n1169), .A2(n1168), .ZN(n1171) );
  OR2_X1 U1151 ( .A1(n1172), .A2(n1173), .ZN(n1104) );
  INV_X1 U1152 ( .A(n1174), .ZN(n1173) );
  OR2_X1 U1153 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
  AND2_X1 U1154 ( .A1(n1176), .A2(n1175), .ZN(n1172) );
  AND2_X1 U1155 ( .A1(n1177), .A2(n1178), .ZN(n1175) );
  INV_X1 U1156 ( .A(n1179), .ZN(n1178) );
  AND2_X1 U1157 ( .A1(n1180), .A2(n1181), .ZN(n1179) );
  OR2_X1 U1158 ( .A1(n1181), .A2(n1180), .ZN(n1177) );
  INV_X1 U1159 ( .A(n1182), .ZN(n1180) );
  INV_X1 U1160 ( .A(n827), .ZN(n830) );
  OR2_X1 U1161 ( .A1(n1183), .A2(n1184), .ZN(n827) );
  AND2_X1 U1162 ( .A1(n824), .A2(n822), .ZN(n1184) );
  AND2_X1 U1163 ( .A1(n817), .A2(n1185), .ZN(n1183) );
  OR2_X1 U1164 ( .A1(n822), .A2(n824), .ZN(n1185) );
  INV_X1 U1165 ( .A(n821), .ZN(n824) );
  AND2_X1 U1166 ( .A1(b_7_), .A2(a_0_), .ZN(n821) );
  OR2_X1 U1167 ( .A1(n1186), .A2(n1187), .ZN(n822) );
  AND2_X1 U1168 ( .A1(n813), .A2(n811), .ZN(n1187) );
  AND2_X1 U1169 ( .A1(n806), .A2(n1188), .ZN(n1186) );
  OR2_X1 U1170 ( .A1(n811), .A2(n813), .ZN(n1188) );
  INV_X1 U1171 ( .A(n810), .ZN(n813) );
  AND2_X1 U1172 ( .A1(b_7_), .A2(a_1_), .ZN(n810) );
  OR2_X1 U1173 ( .A1(n1189), .A2(n1190), .ZN(n811) );
  AND2_X1 U1174 ( .A1(n929), .A2(n927), .ZN(n1190) );
  AND2_X1 U1175 ( .A1(n922), .A2(n1191), .ZN(n1189) );
  OR2_X1 U1176 ( .A1(n929), .A2(n927), .ZN(n1191) );
  OR2_X1 U1177 ( .A1(n1192), .A2(n1193), .ZN(n927) );
  OR2_X1 U1178 ( .A1(n1194), .A2(n1195), .ZN(n929) );
  AND2_X1 U1179 ( .A1(n918), .A2(n917), .ZN(n1195) );
  AND2_X1 U1180 ( .A1(n912), .A2(n1196), .ZN(n1194) );
  OR2_X1 U1181 ( .A1(n918), .A2(n917), .ZN(n1196) );
  OR2_X1 U1182 ( .A1(n1197), .A2(n1198), .ZN(n917) );
  AND2_X1 U1183 ( .A1(n907), .A2(n905), .ZN(n1198) );
  AND2_X1 U1184 ( .A1(n900), .A2(n1199), .ZN(n1197) );
  OR2_X1 U1185 ( .A1(n907), .A2(n905), .ZN(n1199) );
  OR2_X1 U1186 ( .A1(n1200), .A2(n1201), .ZN(n905) );
  AND2_X1 U1187 ( .A1(n895), .A2(n894), .ZN(n1201) );
  AND2_X1 U1188 ( .A1(n889), .A2(n1202), .ZN(n1200) );
  OR2_X1 U1189 ( .A1(n895), .A2(n894), .ZN(n1202) );
  INV_X1 U1190 ( .A(n896), .ZN(n894) );
  OR2_X1 U1191 ( .A1(n1203), .A2(n1193), .ZN(n895) );
  AND2_X1 U1192 ( .A1(n1204), .A2(n1205), .ZN(n889) );
  OR2_X1 U1193 ( .A1(n1206), .A2(n1207), .ZN(n1205) );
  OR2_X1 U1194 ( .A1(n1208), .A2(n1209), .ZN(n1204) );
  INV_X1 U1195 ( .A(n904), .ZN(n907) );
  AND2_X1 U1196 ( .A1(a_4_), .A2(b_7_), .ZN(n904) );
  AND2_X1 U1197 ( .A1(n1210), .A2(n1211), .ZN(n900) );
  INV_X1 U1198 ( .A(n1212), .ZN(n1211) );
  AND2_X1 U1199 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
  OR2_X1 U1200 ( .A1(n1214), .A2(n1213), .ZN(n1210) );
  OR2_X1 U1201 ( .A1(n1215), .A2(n1216), .ZN(n1213) );
  AND2_X1 U1202 ( .A1(n1217), .A2(n1218), .ZN(n1216) );
  INV_X1 U1203 ( .A(n1219), .ZN(n1215) );
  OR2_X1 U1204 ( .A1(n1218), .A2(n1217), .ZN(n1219) );
  OR2_X1 U1205 ( .A1(n1220), .A2(n1193), .ZN(n918) );
  OR2_X1 U1206 ( .A1(n1221), .A2(n1222), .ZN(n912) );
  INV_X1 U1207 ( .A(n1223), .ZN(n1222) );
  OR2_X1 U1208 ( .A1(n1224), .A2(n1225), .ZN(n1223) );
  AND2_X1 U1209 ( .A1(n1225), .A2(n1224), .ZN(n1221) );
  AND2_X1 U1210 ( .A1(n1226), .A2(n1227), .ZN(n1224) );
  INV_X1 U1211 ( .A(n1228), .ZN(n1227) );
  AND2_X1 U1212 ( .A1(n1229), .A2(n1230), .ZN(n1228) );
  OR2_X1 U1213 ( .A1(n1230), .A2(n1229), .ZN(n1226) );
  INV_X1 U1214 ( .A(n1231), .ZN(n1229) );
  AND2_X1 U1215 ( .A1(n1232), .A2(n1233), .ZN(n922) );
  INV_X1 U1216 ( .A(n1234), .ZN(n1233) );
  AND2_X1 U1217 ( .A1(n1235), .A2(n1236), .ZN(n1234) );
  OR2_X1 U1218 ( .A1(n1236), .A2(n1235), .ZN(n1232) );
  OR2_X1 U1219 ( .A1(n1237), .A2(n1238), .ZN(n1235) );
  INV_X1 U1220 ( .A(n1239), .ZN(n1238) );
  OR2_X1 U1221 ( .A1(n1240), .A2(n1241), .ZN(n1239) );
  AND2_X1 U1222 ( .A1(n1241), .A2(n1240), .ZN(n1237) );
  INV_X1 U1223 ( .A(n1242), .ZN(n1241) );
  AND2_X1 U1224 ( .A1(n1243), .A2(n1244), .ZN(n806) );
  INV_X1 U1225 ( .A(n1245), .ZN(n1244) );
  AND2_X1 U1226 ( .A1(n1246), .A2(n1247), .ZN(n1245) );
  OR2_X1 U1227 ( .A1(n1247), .A2(n1246), .ZN(n1243) );
  OR2_X1 U1228 ( .A1(n1248), .A2(n1249), .ZN(n1246) );
  INV_X1 U1229 ( .A(n1250), .ZN(n1249) );
  OR2_X1 U1230 ( .A1(n1251), .A2(n1252), .ZN(n1250) );
  AND2_X1 U1231 ( .A1(n1252), .A2(n1251), .ZN(n1248) );
  INV_X1 U1232 ( .A(n1253), .ZN(n1252) );
  AND2_X1 U1233 ( .A1(n1254), .A2(n1255), .ZN(n817) );
  INV_X1 U1234 ( .A(n1256), .ZN(n1255) );
  AND2_X1 U1235 ( .A1(n1257), .A2(n1129), .ZN(n1256) );
  OR2_X1 U1236 ( .A1(n1129), .A2(n1257), .ZN(n1254) );
  OR2_X1 U1237 ( .A1(n1258), .A2(n1259), .ZN(n1257) );
  INV_X1 U1238 ( .A(n1260), .ZN(n1259) );
  OR2_X1 U1239 ( .A1(n1127), .A2(n1261), .ZN(n1260) );
  AND2_X1 U1240 ( .A1(n1261), .A2(n1127), .ZN(n1258) );
  OR2_X1 U1241 ( .A1(n885), .A2(n1262), .ZN(n1127) );
  INV_X1 U1242 ( .A(n1128), .ZN(n1261) );
  OR2_X1 U1243 ( .A1(n1263), .A2(n1264), .ZN(n1128) );
  AND2_X1 U1244 ( .A1(n1251), .A2(n1253), .ZN(n1264) );
  AND2_X1 U1245 ( .A1(n1247), .A2(n1265), .ZN(n1263) );
  OR2_X1 U1246 ( .A1(n1253), .A2(n1251), .ZN(n1265) );
  OR2_X1 U1247 ( .A1(n885), .A2(n1192), .ZN(n1251) );
  OR2_X1 U1248 ( .A1(n1266), .A2(n1267), .ZN(n1253) );
  AND2_X1 U1249 ( .A1(n1240), .A2(n1242), .ZN(n1267) );
  AND2_X1 U1250 ( .A1(n1236), .A2(n1268), .ZN(n1266) );
  OR2_X1 U1251 ( .A1(n1240), .A2(n1242), .ZN(n1268) );
  OR2_X1 U1252 ( .A1(n1269), .A2(n1270), .ZN(n1242) );
  AND2_X1 U1253 ( .A1(n1231), .A2(n1230), .ZN(n1270) );
  AND2_X1 U1254 ( .A1(n1225), .A2(n1271), .ZN(n1269) );
  OR2_X1 U1255 ( .A1(n1231), .A2(n1230), .ZN(n1271) );
  OR2_X1 U1256 ( .A1(n1272), .A2(n1273), .ZN(n1230) );
  AND2_X1 U1257 ( .A1(n1274), .A2(n1218), .ZN(n1273) );
  AND2_X1 U1258 ( .A1(n1214), .A2(n1275), .ZN(n1272) );
  OR2_X1 U1259 ( .A1(n1274), .A2(n1218), .ZN(n1275) );
  OR2_X1 U1260 ( .A1(n1206), .A2(n1208), .ZN(n1218) );
  INV_X1 U1261 ( .A(n1207), .ZN(n1208) );
  INV_X1 U1262 ( .A(n1209), .ZN(n1206) );
  AND2_X1 U1263 ( .A1(a_7_), .A2(b_5_), .ZN(n1209) );
  INV_X1 U1264 ( .A(n1217), .ZN(n1274) );
  AND2_X1 U1265 ( .A1(a_5_), .A2(b_6_), .ZN(n1217) );
  AND2_X1 U1266 ( .A1(n1276), .A2(n1277), .ZN(n1214) );
  OR3_X1 U1267 ( .A1(n1278), .A2(n1279), .A3(n1280), .ZN(n1277) );
  OR2_X1 U1268 ( .A1(n1281), .A2(n1282), .ZN(n1276) );
  AND2_X1 U1269 ( .A1(a_6_), .A2(b_5_), .ZN(n1282) );
  OR2_X1 U1270 ( .A1(n1283), .A2(n885), .ZN(n1231) );
  OR2_X1 U1271 ( .A1(n1284), .A2(n1285), .ZN(n1225) );
  AND2_X1 U1272 ( .A1(n1286), .A2(n1287), .ZN(n1285) );
  INV_X1 U1273 ( .A(n1288), .ZN(n1284) );
  OR2_X1 U1274 ( .A1(n1286), .A2(n1287), .ZN(n1288) );
  OR2_X1 U1275 ( .A1(n1289), .A2(n1290), .ZN(n1286) );
  AND2_X1 U1276 ( .A1(n1291), .A2(n1292), .ZN(n1290) );
  AND2_X1 U1277 ( .A1(n1293), .A2(n1294), .ZN(n1289) );
  OR2_X1 U1278 ( .A1(n1220), .A2(n885), .ZN(n1240) );
  AND2_X1 U1279 ( .A1(n1295), .A2(n1296), .ZN(n1236) );
  INV_X1 U1280 ( .A(n1297), .ZN(n1296) );
  AND2_X1 U1281 ( .A1(n1298), .A2(n1299), .ZN(n1297) );
  OR2_X1 U1282 ( .A1(n1299), .A2(n1298), .ZN(n1295) );
  OR2_X1 U1283 ( .A1(n1300), .A2(n1301), .ZN(n1298) );
  AND2_X1 U1284 ( .A1(n1302), .A2(n1303), .ZN(n1301) );
  INV_X1 U1285 ( .A(n1304), .ZN(n1302) );
  AND2_X1 U1286 ( .A1(n1305), .A2(n1304), .ZN(n1300) );
  INV_X1 U1287 ( .A(n1303), .ZN(n1305) );
  AND2_X1 U1288 ( .A1(n1306), .A2(n1307), .ZN(n1247) );
  INV_X1 U1289 ( .A(n1308), .ZN(n1307) );
  AND2_X1 U1290 ( .A1(n1309), .A2(n1310), .ZN(n1308) );
  OR2_X1 U1291 ( .A1(n1310), .A2(n1309), .ZN(n1306) );
  OR2_X1 U1292 ( .A1(n1311), .A2(n1312), .ZN(n1309) );
  INV_X1 U1293 ( .A(n1313), .ZN(n1312) );
  OR2_X1 U1294 ( .A1(n1314), .A2(n1315), .ZN(n1313) );
  AND2_X1 U1295 ( .A1(n1315), .A2(n1314), .ZN(n1311) );
  INV_X1 U1296 ( .A(n1316), .ZN(n1315) );
  AND2_X1 U1297 ( .A1(n1317), .A2(n1318), .ZN(n1129) );
  INV_X1 U1298 ( .A(n1319), .ZN(n1318) );
  AND2_X1 U1299 ( .A1(n1320), .A2(n1142), .ZN(n1319) );
  OR2_X1 U1300 ( .A1(n1142), .A2(n1320), .ZN(n1317) );
  OR2_X1 U1301 ( .A1(n1321), .A2(n1322), .ZN(n1320) );
  INV_X1 U1302 ( .A(n1323), .ZN(n1322) );
  OR2_X1 U1303 ( .A1(n1140), .A2(n1324), .ZN(n1323) );
  AND2_X1 U1304 ( .A1(n1324), .A2(n1140), .ZN(n1321) );
  OR2_X1 U1305 ( .A1(n1278), .A2(n1192), .ZN(n1140) );
  INV_X1 U1306 ( .A(n1141), .ZN(n1324) );
  OR2_X1 U1307 ( .A1(n1325), .A2(n1326), .ZN(n1141) );
  AND2_X1 U1308 ( .A1(n1314), .A2(n1316), .ZN(n1326) );
  AND2_X1 U1309 ( .A1(n1310), .A2(n1327), .ZN(n1325) );
  OR2_X1 U1310 ( .A1(n1316), .A2(n1314), .ZN(n1327) );
  OR2_X1 U1311 ( .A1(n1278), .A2(n1220), .ZN(n1314) );
  OR2_X1 U1312 ( .A1(n1328), .A2(n1329), .ZN(n1316) );
  AND2_X1 U1313 ( .A1(n1304), .A2(n1303), .ZN(n1329) );
  AND2_X1 U1314 ( .A1(n1299), .A2(n1330), .ZN(n1328) );
  OR2_X1 U1315 ( .A1(n1304), .A2(n1303), .ZN(n1330) );
  OR2_X1 U1316 ( .A1(n1331), .A2(n1332), .ZN(n1303) );
  AND2_X1 U1317 ( .A1(n1293), .A2(n1287), .ZN(n1332) );
  AND2_X1 U1318 ( .A1(n1333), .A2(n1294), .ZN(n1331) );
  OR2_X1 U1319 ( .A1(n1293), .A2(n1287), .ZN(n1333) );
  OR3_X1 U1320 ( .A1(n1279), .A2(n1281), .A3(n1278), .ZN(n1287) );
  INV_X1 U1321 ( .A(n1280), .ZN(n1281) );
  INV_X1 U1322 ( .A(n1292), .ZN(n1293) );
  OR2_X1 U1323 ( .A1(n1334), .A2(n1335), .ZN(n1292) );
  AND3_X1 U1324 ( .A1(a_7_), .A2(n1336), .A3(b_3_), .ZN(n1335) );
  INV_X1 U1325 ( .A(n1337), .ZN(n1336) );
  AND2_X1 U1326 ( .A1(a_6_), .A2(b_4_), .ZN(n1337) );
  AND3_X1 U1327 ( .A1(a_6_), .A2(n1338), .A3(b_4_), .ZN(n1334) );
  OR2_X1 U1328 ( .A1(n884), .A2(n1339), .ZN(n1338) );
  OR2_X1 U1329 ( .A1(n1283), .A2(n1278), .ZN(n1304) );
  AND2_X1 U1330 ( .A1(n1340), .A2(n1341), .ZN(n1299) );
  INV_X1 U1331 ( .A(n1342), .ZN(n1341) );
  AND2_X1 U1332 ( .A1(n1343), .A2(n1344), .ZN(n1342) );
  OR2_X1 U1333 ( .A1(n1344), .A2(n1343), .ZN(n1340) );
  OR2_X1 U1334 ( .A1(n1345), .A2(n1346), .ZN(n1343) );
  AND2_X1 U1335 ( .A1(n1347), .A2(n1348), .ZN(n1346) );
  AND2_X1 U1336 ( .A1(n1349), .A2(n1350), .ZN(n1345) );
  AND2_X1 U1337 ( .A1(n1351), .A2(n1352), .ZN(n1310) );
  INV_X1 U1338 ( .A(n1353), .ZN(n1352) );
  AND2_X1 U1339 ( .A1(n1354), .A2(n1355), .ZN(n1353) );
  OR2_X1 U1340 ( .A1(n1355), .A2(n1354), .ZN(n1351) );
  OR2_X1 U1341 ( .A1(n1356), .A2(n1357), .ZN(n1354) );
  INV_X1 U1342 ( .A(n1358), .ZN(n1357) );
  OR2_X1 U1343 ( .A1(n1359), .A2(n1360), .ZN(n1358) );
  AND2_X1 U1344 ( .A1(n1360), .A2(n1359), .ZN(n1356) );
  AND2_X1 U1345 ( .A1(n1361), .A2(n1362), .ZN(n1142) );
  INV_X1 U1346 ( .A(n1363), .ZN(n1362) );
  AND2_X1 U1347 ( .A1(n1364), .A2(n1155), .ZN(n1363) );
  OR2_X1 U1348 ( .A1(n1155), .A2(n1364), .ZN(n1361) );
  OR2_X1 U1349 ( .A1(n1365), .A2(n1366), .ZN(n1364) );
  AND2_X1 U1350 ( .A1(n1157), .A2(n1154), .ZN(n1366) );
  INV_X1 U1351 ( .A(n1367), .ZN(n1365) );
  OR2_X1 U1352 ( .A1(n1154), .A2(n1157), .ZN(n1367) );
  AND2_X1 U1353 ( .A1(b_4_), .A2(a_3_), .ZN(n1157) );
  OR2_X1 U1354 ( .A1(n1368), .A2(n1369), .ZN(n1154) );
  AND2_X1 U1355 ( .A1(n1355), .A2(n1359), .ZN(n1369) );
  AND2_X1 U1356 ( .A1(n1370), .A2(n1371), .ZN(n1368) );
  OR2_X1 U1357 ( .A1(n1355), .A2(n1359), .ZN(n1370) );
  OR2_X1 U1358 ( .A1(n1372), .A2(n1373), .ZN(n1359) );
  AND2_X1 U1359 ( .A1(n1350), .A2(n1348), .ZN(n1373) );
  AND2_X1 U1360 ( .A1(n1344), .A2(n1374), .ZN(n1372) );
  OR2_X1 U1361 ( .A1(n1350), .A2(n1348), .ZN(n1374) );
  INV_X1 U1362 ( .A(n1349), .ZN(n1348) );
  AND2_X1 U1363 ( .A1(n1375), .A2(n1280), .ZN(n1349) );
  AND2_X1 U1364 ( .A1(a_7_), .A2(b_4_), .ZN(n1280) );
  INV_X1 U1365 ( .A(n1347), .ZN(n1350) );
  AND2_X1 U1366 ( .A1(a_5_), .A2(b_4_), .ZN(n1347) );
  AND2_X1 U1367 ( .A1(n1376), .A2(n1377), .ZN(n1344) );
  OR3_X1 U1368 ( .A1(n884), .A2(n1378), .A3(n1375), .ZN(n1377) );
  INV_X1 U1369 ( .A(n1379), .ZN(n1376) );
  AND2_X1 U1370 ( .A1(n1375), .A2(n1380), .ZN(n1379) );
  OR2_X1 U1371 ( .A1(n1378), .A2(n884), .ZN(n1380) );
  AND2_X1 U1372 ( .A1(n1381), .A2(n1382), .ZN(n1355) );
  INV_X1 U1373 ( .A(n1383), .ZN(n1382) );
  AND2_X1 U1374 ( .A1(n1384), .A2(n1385), .ZN(n1383) );
  OR2_X1 U1375 ( .A1(n1385), .A2(n1384), .ZN(n1381) );
  OR2_X1 U1376 ( .A1(n1386), .A2(n1387), .ZN(n1384) );
  AND2_X1 U1377 ( .A1(n1388), .A2(n1389), .ZN(n1387) );
  AND2_X1 U1378 ( .A1(n1390), .A2(n1391), .ZN(n1386) );
  AND2_X1 U1379 ( .A1(n1392), .A2(n1393), .ZN(n1155) );
  INV_X1 U1380 ( .A(n1394), .ZN(n1393) );
  AND2_X1 U1381 ( .A1(n1395), .A2(n1170), .ZN(n1394) );
  OR2_X1 U1382 ( .A1(n1170), .A2(n1395), .ZN(n1392) );
  OR2_X1 U1383 ( .A1(n1396), .A2(n1397), .ZN(n1395) );
  AND2_X1 U1384 ( .A1(n1398), .A2(n1169), .ZN(n1397) );
  INV_X1 U1385 ( .A(n1399), .ZN(n1169) );
  INV_X1 U1386 ( .A(n1168), .ZN(n1398) );
  AND2_X1 U1387 ( .A1(n1399), .A2(n1168), .ZN(n1396) );
  OR2_X1 U1388 ( .A1(n1400), .A2(n1401), .ZN(n1168) );
  AND2_X1 U1389 ( .A1(n1391), .A2(n1389), .ZN(n1401) );
  AND2_X1 U1390 ( .A1(n1385), .A2(n1402), .ZN(n1400) );
  OR2_X1 U1391 ( .A1(n1389), .A2(n1391), .ZN(n1402) );
  INV_X1 U1392 ( .A(n1388), .ZN(n1391) );
  AND3_X1 U1393 ( .A1(b_2_), .A2(a_7_), .A3(n1375), .ZN(n1388) );
  AND2_X1 U1394 ( .A1(a_6_), .A2(b_3_), .ZN(n1375) );
  INV_X1 U1395 ( .A(n1390), .ZN(n1389) );
  AND2_X1 U1396 ( .A1(a_5_), .A2(b_3_), .ZN(n1390) );
  AND2_X1 U1397 ( .A1(n1403), .A2(n1404), .ZN(n1385) );
  INV_X1 U1398 ( .A(n1405), .ZN(n1404) );
  AND2_X1 U1399 ( .A1(n1406), .A2(n1407), .ZN(n1405) );
  OR2_X1 U1400 ( .A1(n1407), .A2(n1406), .ZN(n1403) );
  AND2_X1 U1401 ( .A1(b_3_), .A2(a_4_), .ZN(n1399) );
  AND2_X1 U1402 ( .A1(n1408), .A2(n1409), .ZN(n1170) );
  INV_X1 U1403 ( .A(n1410), .ZN(n1409) );
  AND2_X1 U1404 ( .A1(n1411), .A2(n1412), .ZN(n1410) );
  OR2_X1 U1405 ( .A1(n1412), .A2(n1411), .ZN(n1408) );
  OR2_X1 U1406 ( .A1(n1413), .A2(n1414), .ZN(n1411) );
  AND2_X1 U1407 ( .A1(n1415), .A2(n1416), .ZN(n1414) );
  INV_X1 U1408 ( .A(n1417), .ZN(n1415) );
  AND2_X1 U1409 ( .A1(n1418), .A2(n1417), .ZN(n1413) );
  INV_X1 U1410 ( .A(n1416), .ZN(n1418) );
  AND2_X1 U1411 ( .A1(n878), .A2(n937), .ZN(n875) );
  INV_X1 U1412 ( .A(n877), .ZN(n937) );
  OR2_X1 U1413 ( .A1(n938), .A2(n939), .ZN(n877) );
  OR2_X1 U1414 ( .A1(n1419), .A2(n1420), .ZN(n939) );
  AND2_X1 U1415 ( .A1(n963), .A2(n962), .ZN(n1420) );
  AND2_X1 U1416 ( .A1(n955), .A2(n1421), .ZN(n1419) );
  OR2_X1 U1417 ( .A1(n962), .A2(n963), .ZN(n1421) );
  OR2_X1 U1418 ( .A1(n1378), .A2(n1422), .ZN(n963) );
  OR2_X1 U1419 ( .A1(n1423), .A2(n1424), .ZN(n962) );
  AND2_X1 U1420 ( .A1(n996), .A2(n998), .ZN(n1424) );
  AND2_X1 U1421 ( .A1(n992), .A2(n1425), .ZN(n1423) );
  OR2_X1 U1422 ( .A1(n998), .A2(n996), .ZN(n1425) );
  OR2_X1 U1423 ( .A1(n1378), .A2(n1262), .ZN(n996) );
  OR2_X1 U1424 ( .A1(n1426), .A2(n1427), .ZN(n998) );
  AND2_X1 U1425 ( .A1(n1051), .A2(n1055), .ZN(n1427) );
  AND2_X1 U1426 ( .A1(n1428), .A2(n1429), .ZN(n1426) );
  OR2_X1 U1427 ( .A1(n1051), .A2(n1055), .ZN(n1428) );
  OR2_X1 U1428 ( .A1(n1430), .A2(n1431), .ZN(n1055) );
  AND2_X1 U1429 ( .A1(n1432), .A2(n1117), .ZN(n1431) );
  AND2_X1 U1430 ( .A1(n1112), .A2(n1433), .ZN(n1430) );
  OR2_X1 U1431 ( .A1(n1117), .A2(n1432), .ZN(n1433) );
  INV_X1 U1432 ( .A(n1116), .ZN(n1432) );
  AND2_X1 U1433 ( .A1(b_2_), .A2(a_3_), .ZN(n1116) );
  OR2_X1 U1434 ( .A1(n1434), .A2(n1435), .ZN(n1117) );
  AND2_X1 U1435 ( .A1(n1182), .A2(n1181), .ZN(n1435) );
  AND2_X1 U1436 ( .A1(n1176), .A2(n1436), .ZN(n1434) );
  OR2_X1 U1437 ( .A1(n1181), .A2(n1182), .ZN(n1436) );
  OR2_X1 U1438 ( .A1(n1378), .A2(n1283), .ZN(n1182) );
  OR2_X1 U1439 ( .A1(n1437), .A2(n1438), .ZN(n1181) );
  AND2_X1 U1440 ( .A1(n1417), .A2(n1416), .ZN(n1438) );
  AND2_X1 U1441 ( .A1(n1412), .A2(n1439), .ZN(n1437) );
  OR2_X1 U1442 ( .A1(n1416), .A2(n1417), .ZN(n1439) );
  OR2_X1 U1443 ( .A1(n1378), .A2(n1203), .ZN(n1417) );
  OR2_X1 U1444 ( .A1(n1407), .A2(n1440), .ZN(n1416) );
  INV_X1 U1445 ( .A(n1406), .ZN(n1440) );
  OR2_X1 U1446 ( .A1(n1279), .A2(n1378), .ZN(n1407) );
  AND2_X1 U1447 ( .A1(n1441), .A2(n1442), .ZN(n1412) );
  OR2_X1 U1448 ( .A1(n1443), .A2(n1444), .ZN(n1442) );
  INV_X1 U1449 ( .A(n1445), .ZN(n1441) );
  AND2_X1 U1450 ( .A1(n1444), .A2(n1443), .ZN(n1445) );
  OR2_X1 U1451 ( .A1(n884), .A2(n1446), .ZN(n1443) );
  OR2_X1 U1452 ( .A1(n1447), .A2(n1448), .ZN(n1176) );
  INV_X1 U1453 ( .A(n1449), .ZN(n1448) );
  OR2_X1 U1454 ( .A1(n1450), .A2(n1451), .ZN(n1449) );
  AND2_X1 U1455 ( .A1(n1451), .A2(n1450), .ZN(n1447) );
  OR2_X1 U1456 ( .A1(n1452), .A2(n1453), .ZN(n1450) );
  AND3_X1 U1457 ( .A1(a_6_), .A2(n1454), .A3(b_0_), .ZN(n1453) );
  OR2_X1 U1458 ( .A1(n1455), .A2(n1203), .ZN(n1454) );
  AND3_X1 U1459 ( .A1(b_1_), .A2(n1456), .A3(a_5_), .ZN(n1452) );
  OR2_X1 U1460 ( .A1(n1279), .A2(n1446), .ZN(n1456) );
  OR2_X1 U1461 ( .A1(n1457), .A2(n1458), .ZN(n1112) );
  AND2_X1 U1462 ( .A1(n1459), .A2(n1460), .ZN(n1458) );
  INV_X1 U1463 ( .A(n1461), .ZN(n1457) );
  OR2_X1 U1464 ( .A1(n1459), .A2(n1460), .ZN(n1461) );
  OR2_X1 U1465 ( .A1(n1462), .A2(n1463), .ZN(n1459) );
  AND2_X1 U1466 ( .A1(n1464), .A2(n1465), .ZN(n1463) );
  AND2_X1 U1467 ( .A1(n1466), .A2(n1467), .ZN(n1462) );
  AND2_X1 U1468 ( .A1(n1468), .A2(n1469), .ZN(n1051) );
  INV_X1 U1469 ( .A(n1470), .ZN(n1469) );
  AND2_X1 U1470 ( .A1(n1471), .A2(n1472), .ZN(n1470) );
  OR2_X1 U1471 ( .A1(n1471), .A2(n1472), .ZN(n1468) );
  OR2_X1 U1472 ( .A1(n1473), .A2(n1474), .ZN(n1471) );
  INV_X1 U1473 ( .A(n1475), .ZN(n1474) );
  OR2_X1 U1474 ( .A1(n1476), .A2(n1477), .ZN(n1475) );
  AND2_X1 U1475 ( .A1(n1477), .A2(n1476), .ZN(n1473) );
  INV_X1 U1476 ( .A(n1478), .ZN(n1477) );
  AND2_X1 U1477 ( .A1(n1479), .A2(n1480), .ZN(n992) );
  INV_X1 U1478 ( .A(n1481), .ZN(n1480) );
  AND2_X1 U1479 ( .A1(n1482), .A2(n1483), .ZN(n1481) );
  OR2_X1 U1480 ( .A1(n1482), .A2(n1483), .ZN(n1479) );
  OR2_X1 U1481 ( .A1(n1484), .A2(n1485), .ZN(n1482) );
  AND2_X1 U1482 ( .A1(n1486), .A2(n1487), .ZN(n1485) );
  INV_X1 U1483 ( .A(n1488), .ZN(n1486) );
  AND2_X1 U1484 ( .A1(n1489), .A2(n1488), .ZN(n1484) );
  INV_X1 U1485 ( .A(n1487), .ZN(n1489) );
  AND2_X1 U1486 ( .A1(n1490), .A2(n1491), .ZN(n955) );
  INV_X1 U1487 ( .A(n1492), .ZN(n1491) );
  AND2_X1 U1488 ( .A1(n1493), .A2(n1494), .ZN(n1492) );
  OR2_X1 U1489 ( .A1(n1493), .A2(n1494), .ZN(n1490) );
  OR2_X1 U1490 ( .A1(n1495), .A2(n1496), .ZN(n1493) );
  AND2_X1 U1491 ( .A1(n1497), .A2(n1498), .ZN(n1496) );
  INV_X1 U1492 ( .A(n1499), .ZN(n1495) );
  OR2_X1 U1493 ( .A1(n1498), .A2(n1497), .ZN(n1499) );
  AND2_X1 U1494 ( .A1(n1500), .A2(n1501), .ZN(n938) );
  INV_X1 U1495 ( .A(n1502), .ZN(n1501) );
  AND2_X1 U1496 ( .A1(n1503), .A2(n1504), .ZN(n1502) );
  OR2_X1 U1497 ( .A1(n1503), .A2(n1504), .ZN(n1500) );
  OR2_X1 U1498 ( .A1(n1505), .A2(n1506), .ZN(n1503) );
  INV_X1 U1499 ( .A(n1507), .ZN(n1506) );
  OR2_X1 U1500 ( .A1(n1508), .A2(n1509), .ZN(n1507) );
  AND2_X1 U1501 ( .A1(n1509), .A2(n1508), .ZN(n1505) );
  INV_X1 U1502 ( .A(n1510), .ZN(n1509) );
  OR2_X1 U1503 ( .A1(n1511), .A2(n1512), .ZN(n878) );
  AND2_X1 U1504 ( .A1(n1513), .A2(n933), .ZN(n1512) );
  INV_X1 U1505 ( .A(n1514), .ZN(n1511) );
  OR2_X1 U1506 ( .A1(n933), .A2(n1513), .ZN(n1514) );
  AND2_X1 U1507 ( .A1(b_0_), .A2(a_0_), .ZN(n1513) );
  OR2_X1 U1508 ( .A1(n1515), .A2(n1516), .ZN(n933) );
  AND2_X1 U1509 ( .A1(n1504), .A2(n1510), .ZN(n1516) );
  AND2_X1 U1510 ( .A1(n1517), .A2(n1508), .ZN(n1515) );
  OR2_X1 U1511 ( .A1(n1455), .A2(n1422), .ZN(n1508) );
  OR2_X1 U1512 ( .A1(n1510), .A2(n1504), .ZN(n1517) );
  OR2_X1 U1513 ( .A1(n1262), .A2(n1446), .ZN(n1504) );
  OR2_X1 U1514 ( .A1(n1518), .A2(n1519), .ZN(n1510) );
  AND2_X1 U1515 ( .A1(n1494), .A2(n1498), .ZN(n1519) );
  AND2_X1 U1516 ( .A1(n1520), .A2(n1521), .ZN(n1518) );
  OR2_X1 U1517 ( .A1(n1498), .A2(n1494), .ZN(n1520) );
  OR2_X1 U1518 ( .A1(n1192), .A2(n1446), .ZN(n1494) );
  OR2_X1 U1519 ( .A1(n1522), .A2(n1523), .ZN(n1498) );
  AND2_X1 U1520 ( .A1(n1483), .A2(n1488), .ZN(n1523) );
  AND2_X1 U1521 ( .A1(n1524), .A2(n1487), .ZN(n1522) );
  OR2_X1 U1522 ( .A1(n1220), .A2(n1446), .ZN(n1487) );
  OR2_X1 U1523 ( .A1(n1488), .A2(n1483), .ZN(n1524) );
  OR2_X1 U1524 ( .A1(n1455), .A2(n1192), .ZN(n1483) );
  OR2_X1 U1525 ( .A1(n1525), .A2(n1526), .ZN(n1488) );
  AND2_X1 U1526 ( .A1(n1472), .A2(n1478), .ZN(n1526) );
  AND2_X1 U1527 ( .A1(n1527), .A2(n1476), .ZN(n1525) );
  OR2_X1 U1528 ( .A1(n1455), .A2(n1220), .ZN(n1476) );
  OR2_X1 U1529 ( .A1(n1478), .A2(n1472), .ZN(n1527) );
  OR2_X1 U1530 ( .A1(n1283), .A2(n1446), .ZN(n1472) );
  OR2_X1 U1531 ( .A1(n1528), .A2(n1529), .ZN(n1478) );
  AND2_X1 U1532 ( .A1(n1460), .A2(n1465), .ZN(n1529) );
  AND2_X1 U1533 ( .A1(n1464), .A2(n1530), .ZN(n1528) );
  OR2_X1 U1534 ( .A1(n1465), .A2(n1460), .ZN(n1530) );
  OR2_X1 U1535 ( .A1(n1455), .A2(n1283), .ZN(n1460) );
  INV_X1 U1536 ( .A(a_4_), .ZN(n1283) );
  INV_X1 U1537 ( .A(n1466), .ZN(n1465) );
  INV_X1 U1538 ( .A(n1467), .ZN(n1464) );
  OR2_X1 U1539 ( .A1(n1531), .A2(n1451), .ZN(n1467) );
  AND3_X1 U1540 ( .A1(a_6_), .A2(n1406), .A3(b_0_), .ZN(n1451) );
  AND2_X1 U1541 ( .A1(a_7_), .A2(b_1_), .ZN(n1406) );
  AND2_X1 U1542 ( .A1(n1466), .A2(n1444), .ZN(n1531) );
  AND2_X1 U1543 ( .A1(a_6_), .A2(b_1_), .ZN(n1444) );
  AND2_X1 U1544 ( .A1(a_5_), .A2(b_0_), .ZN(n1466) );
  OR2_X1 U1545 ( .A1(n1532), .A2(n1533), .ZN(Result_add_7_) );
  AND2_X1 U1546 ( .A1(a_7_), .A2(n1193), .ZN(n1533) );
  AND2_X1 U1547 ( .A1(b_7_), .A2(n884), .ZN(n1532) );
  OR3_X1 U1548 ( .A1(n1534), .A2(n1535), .A3(n896), .ZN(Result_add_6_) );
  AND2_X1 U1549 ( .A1(n1207), .A2(Result_mul_15_), .ZN(n896) );
  AND3_X1 U1550 ( .A1(n1536), .A2(n1279), .A3(b_6_), .ZN(n1535) );
  AND2_X1 U1551 ( .A1(n1537), .A2(n885), .ZN(n1534) );
  INV_X1 U1552 ( .A(b_6_), .ZN(n885) );
  OR2_X1 U1553 ( .A1(n1538), .A2(n1539), .ZN(n1537) );
  AND2_X1 U1554 ( .A1(Result_mul_15_), .A2(n1279), .ZN(n1539) );
  INV_X1 U1555 ( .A(a_6_), .ZN(n1279) );
  AND2_X1 U1556 ( .A1(a_6_), .A2(n1536), .ZN(n1538) );
  OR2_X1 U1557 ( .A1(n1540), .A2(n1541), .ZN(Result_add_5_) );
  AND2_X1 U1558 ( .A1(n1542), .A2(n1543), .ZN(n1541) );
  OR2_X1 U1559 ( .A1(n1544), .A2(n1545), .ZN(n1542) );
  AND2_X1 U1560 ( .A1(a_5_), .A2(n1278), .ZN(n1545) );
  AND2_X1 U1561 ( .A1(b_5_), .A2(n1203), .ZN(n1544) );
  AND2_X1 U1562 ( .A1(n1546), .A2(n1547), .ZN(n1540) );
  OR2_X1 U1563 ( .A1(n1291), .A2(n1548), .ZN(n1546) );
  OR2_X1 U1564 ( .A1(n1549), .A2(n1550), .ZN(Result_add_4_) );
  AND2_X1 U1565 ( .A1(n1551), .A2(n1552), .ZN(n1550) );
  AND2_X1 U1566 ( .A1(n1553), .A2(n1554), .ZN(n1549) );
  OR2_X1 U1567 ( .A1(n1555), .A2(n1360), .ZN(n1554) );
  INV_X1 U1568 ( .A(n1556), .ZN(n1553) );
  OR3_X1 U1569 ( .A1(n1557), .A2(n1558), .A3(n1559), .ZN(Result_add_3_) );
  AND2_X1 U1570 ( .A1(n1560), .A2(n1164), .ZN(n1559) );
  AND2_X1 U1571 ( .A1(n1561), .A2(n1339), .ZN(n1558) );
  OR2_X1 U1572 ( .A1(n1562), .A2(n1563), .ZN(n1561) );
  AND2_X1 U1573 ( .A1(n1560), .A2(n1220), .ZN(n1563) );
  INV_X1 U1574 ( .A(n1564), .ZN(n1560) );
  AND2_X1 U1575 ( .A1(a_3_), .A2(n1564), .ZN(n1562) );
  AND3_X1 U1576 ( .A1(n1564), .A2(n1220), .A3(b_3_), .ZN(n1557) );
  OR2_X1 U1577 ( .A1(n1565), .A2(n1566), .ZN(Result_add_2_) );
  INV_X1 U1578 ( .A(n1567), .ZN(n1566) );
  OR2_X1 U1579 ( .A1(n1568), .A2(n1569), .ZN(n1567) );
  AND2_X1 U1580 ( .A1(n1569), .A2(n1568), .ZN(n1565) );
  OR2_X1 U1581 ( .A1(n1570), .A2(n1056), .ZN(n1568) );
  INV_X1 U1582 ( .A(n1571), .ZN(n1569) );
  OR3_X1 U1583 ( .A1(n1572), .A2(n1573), .A3(n1574), .ZN(Result_add_1_) );
  AND2_X1 U1584 ( .A1(n1575), .A2(n1497), .ZN(n1574) );
  AND2_X1 U1585 ( .A1(n1576), .A2(n1455), .ZN(n1573) );
  OR2_X1 U1586 ( .A1(n1577), .A2(n1578), .ZN(n1576) );
  AND2_X1 U1587 ( .A1(n1575), .A2(n1262), .ZN(n1578) );
  INV_X1 U1588 ( .A(n1579), .ZN(n1575) );
  AND2_X1 U1589 ( .A1(a_1_), .A2(n1579), .ZN(n1577) );
  AND3_X1 U1590 ( .A1(n1579), .A2(n1262), .A3(b_1_), .ZN(n1572) );
  OR2_X1 U1591 ( .A1(n1580), .A2(n1581), .ZN(Result_add_0_) );
  AND2_X1 U1592 ( .A1(n1582), .A2(n1583), .ZN(n1581) );
  INV_X1 U1593 ( .A(n1584), .ZN(n1580) );
  OR2_X1 U1594 ( .A1(n1583), .A2(n1582), .ZN(n1584) );
  OR2_X1 U1595 ( .A1(n1585), .A2(n1586), .ZN(n1582) );
  AND2_X1 U1596 ( .A1(a_0_), .A2(n1446), .ZN(n1586) );
  INV_X1 U1597 ( .A(b_0_), .ZN(n1446) );
  AND2_X1 U1598 ( .A1(b_0_), .A2(n1422), .ZN(n1585) );
  INV_X1 U1599 ( .A(a_0_), .ZN(n1422) );
  OR2_X1 U1600 ( .A1(n1587), .A2(n1588), .ZN(n1583) );
  AND2_X1 U1601 ( .A1(n1262), .A2(n1455), .ZN(n1588) );
  INV_X1 U1602 ( .A(b_1_), .ZN(n1455) );
  INV_X1 U1603 ( .A(a_1_), .ZN(n1262) );
  AND2_X1 U1604 ( .A1(n1579), .A2(n1521), .ZN(n1587) );
  INV_X1 U1605 ( .A(n1497), .ZN(n1521) );
  AND2_X1 U1606 ( .A1(b_1_), .A2(a_1_), .ZN(n1497) );
  OR2_X1 U1607 ( .A1(n1589), .A2(n1570), .ZN(n1579) );
  AND2_X1 U1608 ( .A1(n1192), .A2(n1378), .ZN(n1570) );
  INV_X1 U1609 ( .A(b_2_), .ZN(n1378) );
  INV_X1 U1610 ( .A(a_2_), .ZN(n1192) );
  AND2_X1 U1611 ( .A1(n1571), .A2(n1429), .ZN(n1589) );
  INV_X1 U1612 ( .A(n1056), .ZN(n1429) );
  AND2_X1 U1613 ( .A1(b_2_), .A2(a_2_), .ZN(n1056) );
  OR2_X1 U1614 ( .A1(n1590), .A2(n1591), .ZN(n1571) );
  AND2_X1 U1615 ( .A1(n1220), .A2(n1339), .ZN(n1591) );
  INV_X1 U1616 ( .A(b_3_), .ZN(n1339) );
  INV_X1 U1617 ( .A(a_3_), .ZN(n1220) );
  AND2_X1 U1618 ( .A1(n1107), .A2(n1564), .ZN(n1590) );
  OR2_X1 U1619 ( .A1(n1555), .A2(n1551), .ZN(n1564) );
  AND2_X1 U1620 ( .A1(n1371), .A2(n1556), .ZN(n1551) );
  OR2_X1 U1621 ( .A1(n1548), .A2(n1592), .ZN(n1556) );
  AND2_X1 U1622 ( .A1(n1543), .A2(n1294), .ZN(n1592) );
  INV_X1 U1623 ( .A(n1291), .ZN(n1294) );
  AND2_X1 U1624 ( .A1(a_5_), .A2(b_5_), .ZN(n1291) );
  INV_X1 U1625 ( .A(n1547), .ZN(n1543) );
  OR2_X1 U1626 ( .A1(n1593), .A2(n1207), .ZN(n1547) );
  AND2_X1 U1627 ( .A1(a_6_), .A2(b_6_), .ZN(n1207) );
  AND2_X1 U1628 ( .A1(Result_mul_15_), .A2(n1594), .ZN(n1593) );
  OR2_X1 U1629 ( .A1(a_6_), .A2(b_6_), .ZN(n1594) );
  INV_X1 U1630 ( .A(n1536), .ZN(Result_mul_15_) );
  OR2_X1 U1631 ( .A1(n884), .A2(n1193), .ZN(n1536) );
  INV_X1 U1632 ( .A(b_7_), .ZN(n1193) );
  INV_X1 U1633 ( .A(a_7_), .ZN(n884) );
  AND2_X1 U1634 ( .A1(n1203), .A2(n1278), .ZN(n1548) );
  INV_X1 U1635 ( .A(b_5_), .ZN(n1278) );
  INV_X1 U1636 ( .A(a_5_), .ZN(n1203) );
  INV_X1 U1637 ( .A(n1360), .ZN(n1371) );
  AND2_X1 U1638 ( .A1(a_4_), .A2(b_4_), .ZN(n1360) );
  INV_X1 U1639 ( .A(n1552), .ZN(n1555) );
  OR2_X1 U1640 ( .A1(a_4_), .A2(b_4_), .ZN(n1552) );
  INV_X1 U1641 ( .A(n1164), .ZN(n1107) );
  AND2_X1 U1642 ( .A1(b_3_), .A2(a_3_), .ZN(n1164) );
endmodule

