module s38417 ( CK, g1249, g16297, g16355, g16399, g16437, g16496, g1943, 
        g24734, g25420, g25435, g25442, g25489, g26104, g26135, g26149, g2637, 
        g27380, g3212, g3213, g3214, g3215, g3216, g3217, g3218, g3219, g3220, 
        g3221, g3222, g3223, g3224, g3225, g3226, g3227, g3228, g3229, g3230, 
        g3231, g3232, g3233, g3234, g3993, g4088, g4090, g4200, g4321, g4323, 
        g4450, g4590, g51, g5388, g5437, g5472, g5511, g5549, g5555, g5595, 
        g5612, g5629, g563, g5637, g5648, g5657, g5686, g5695, g5738, g5747, 
        g5796, g6225, g6231, g6313, g6368, g6442, g6447, g6485, g6518, g6573, 
        g6642, g6677, g6712, g6750, g6782, g6837, g6895, g6911, g6944, g6979, 
        g7014, g7052, g7084, g7161, g7194, g7229, g7264, g7302, g7334, g7357, 
        g7390, g7425, g7487, g7519, g7909, g7956, g7961, g8007, g8012, g8021, 
        g8023, g8030, g8082, g8087, g8096, g8106, g8167, g8175, g8249, g8251, 
        g8258, g8259, g8260, g8261, g8262, g8263, g8264, g8265, g8266, g8267, 
        g8268, g8269, g8270, g8271, g8272, g8273, g8274, g8275, test_se, 
        test_si1, test_so1, test_si2, test_so2, test_si3, test_so3, test_si4, 
        test_so4, test_si5, test_so5, test_si6, test_so6, test_si7, test_so7, 
        test_si8, test_so8, test_si9, test_so9, test_si10, test_so10, 
        test_si11, test_so11, test_si12, test_so12, test_si13, test_so13, 
        test_si14, test_so14, test_si15, test_so15, test_si16, test_so16, 
        test_si17, test_so17, test_si18, test_so18, test_si19, test_so19, 
        test_si20, test_so20, test_si21, test_so21, test_si22, test_so22, 
        test_si23, test_so23, test_si24, test_so24, test_si25, test_so25, 
        test_si26, test_so26, test_si27, test_so27, test_si28, test_so28, 
        test_si29, test_so29, test_si30, test_so30, test_si31, test_so31, 
        test_si32, test_so32, test_si33, test_so33, test_si34, test_so34, 
        test_si35, test_so35, test_si36, test_so36, test_si37, test_so37, 
        test_si38, test_so38, test_si39, test_so39, test_si40, test_so40, 
        test_si41, test_so41, test_si42, test_so42, test_si43, test_so43, 
        test_si44, test_so44, test_si45, test_so45, test_si46, test_so46, 
        test_si47, test_so47, test_si48, test_so48, test_si49, test_so49, 
        test_si50, test_so50, test_si51, test_so51, test_si52, test_so52, 
        test_si53, test_so53, test_si54, test_so54, test_si55, test_so55, 
        test_si56, test_so56, test_si57, test_so57, test_si58, test_so58, 
        test_si59, test_so59, test_si60, test_so60, test_si61, test_so61, 
        test_si62, test_so62, test_si63, test_so63, test_si64, test_so64, 
        test_si65, test_so65, test_si66, test_so66, test_si67, test_so67, 
        test_si68, test_so68, test_si69, test_so69, test_si70, test_so70, 
        test_si71, test_so71, test_si72, test_so72, test_si73, test_so73, 
        test_si74, test_so74, test_si75, test_so75, test_si76, test_so76, 
        test_si77, test_so77, test_si78, test_so78, test_si79, test_so79, 
        test_si80, test_so80, test_si81, test_so81, test_si82, test_so82, 
        test_si83, test_so83, test_si84, test_so84, test_si85, test_so85, 
        test_si86, test_so86, test_si87, test_so87, test_si88, test_so88, 
        test_si89, test_so89, test_si90, test_so90, test_si91, test_so91, 
        test_si92, test_so92, test_si93, test_so93, test_si94, test_so94, 
        test_si95, test_so95, test_si96, test_so96, test_si97, test_so97, 
        test_si98, test_so98, test_si99, test_so99, test_si100, test_so100 );
  input CK, g1249, g1943, g2637, g3212, g3213, g3214, g3215, g3216, g3217,
         g3218, g3219, g3220, g3221, g3222, g3223, g3224, g3225, g3226, g3227,
         g3228, g3229, g3230, g3231, g3232, g3233, g3234, g51, g563, test_se,
         test_si1, test_si2, test_si3, test_si4, test_si5, test_si6, test_si7,
         test_si8, test_si9, test_si10, test_si11, test_si12, test_si13,
         test_si14, test_si15, test_si16, test_si17, test_si18, test_si19,
         test_si20, test_si21, test_si22, test_si23, test_si24, test_si25,
         test_si26, test_si27, test_si28, test_si29, test_si30, test_si31,
         test_si32, test_si33, test_si34, test_si35, test_si36, test_si37,
         test_si38, test_si39, test_si40, test_si41, test_si42, test_si43,
         test_si44, test_si45, test_si46, test_si47, test_si48, test_si49,
         test_si50, test_si51, test_si52, test_si53, test_si54, test_si55,
         test_si56, test_si57, test_si58, test_si59, test_si60, test_si61,
         test_si62, test_si63, test_si64, test_si65, test_si66, test_si67,
         test_si68, test_si69, test_si70, test_si71, test_si72, test_si73,
         test_si74, test_si75, test_si76, test_si77, test_si78, test_si79,
         test_si80, test_si81, test_si82, test_si83, test_si84, test_si85,
         test_si86, test_si87, test_si88, test_si89, test_si90, test_si91,
         test_si92, test_si93, test_si94, test_si95, test_si96, test_si97,
         test_si98, test_si99, test_si100;
  output g16297, g16355, g16399, g16437, g16496, g24734, g25420, g25435,
         g25442, g25489, g26104, g26135, g26149, g27380, g3993, g4088, g4090,
         g4200, g4321, g4323, g4450, g4590, g5388, g5437, g5472, g5511, g5549,
         g5555, g5595, g5612, g5629, g5637, g5648, g5657, g5686, g5695, g5738,
         g5747, g5796, g6225, g6231, g6313, g6368, g6442, g6447, g6485, g6518,
         g6573, g6642, g6677, g6712, g6750, g6782, g6837, g6895, g6911, g6944,
         g6979, g7014, g7052, g7084, g7161, g7194, g7229, g7264, g7302, g7334,
         g7357, g7390, g7425, g7487, g7519, g7909, g7956, g7961, g8007, g8012,
         g8021, g8023, g8030, g8082, g8087, g8096, g8106, g8167, g8175, g8249,
         g8251, g8258, g8259, g8260, g8261, g8262, g8263, g8264, g8265, g8266,
         g8267, g8268, g8269, g8270, g8271, g8272, g8273, g8274, g8275,
         test_so1, test_so2, test_so3, test_so4, test_so5, test_so6, test_so7,
         test_so8, test_so9, test_so10, test_so11, test_so12, test_so13,
         test_so14, test_so15, test_so16, test_so17, test_so18, test_so19,
         test_so20, test_so21, test_so22, test_so23, test_so24, test_so25,
         test_so26, test_so27, test_so28, test_so29, test_so30, test_so31,
         test_so32, test_so33, test_so34, test_so35, test_so36, test_so37,
         test_so38, test_so39, test_so40, test_so41, test_so42, test_so43,
         test_so44, test_so45, test_so46, test_so47, test_so48, test_so49,
         test_so50, test_so51, test_so52, test_so53, test_so54, test_so55,
         test_so56, test_so57, test_so58, test_so59, test_so60, test_so61,
         test_so62, test_so63, test_so64, test_so65, test_so66, test_so67,
         test_so68, test_so69, test_so70, test_so71, test_so72, test_so73,
         test_so74, test_so75, test_so76, test_so77, test_so78, test_so79,
         test_so80, test_so81, test_so82, test_so83, test_so84, test_so85,
         test_so86, test_so87, test_so88, test_so89, test_so90, test_so91,
         test_so92, test_so93, test_so94, test_so95, test_so96, test_so97,
         test_so98, test_so99, test_so100;
  wire   test_so3, test_so4, test_so5, test_so23, test_so57, test_so63,
         test_so73, test_so99, test_so100, n2230, n2217, n2231, n2374, n2361,
         n2375, DFF_2_n1, n4264, n2445, n2446, n2440, n2426, n2670, n2671,
         n2669, n2685, n2686, n2684, n2718, n2719, n2717, n2982, g2124, n2981,
         n2985, g1430, n2984, n2988, g744, n2987, n2991, g56, n2990, n3742,
         n3741, n8104, g16802, n8103, DFF_1_n1, g16823, n8102, g2950, n4423,
         n4274, g2883, n4330, g22026, g2888, g23358, g2896, n4431, g24473,
         g2892, g25201, g2903, n4305, g26037, g2900, n4291, g26798, g2908,
         n4355, n4273, g2912, n4482, g23357, g2917, n4479, g24476, g2924,
         n4349, g25199, g2920, n4280, DFF_15_n1, n4281, n8099, DFF_16_n1,
         n8098, DFF_18_n1, n4279, g2879, n4351, g2934, g2935, g2938, g2941,
         g2944, g2947, g2953, g2956, g2959, g2962, g2963, g2969, g2972, g2975,
         g2978, g2981, g2874, g18754, g1506, n4288, g18781, g1501, n4565,
         g18803, g1496, n4557, g18821, g1491, n4326, g18835, g1486, n4390,
         g18852, g1481, n4320, g18866, g1476, n4374, g18883, g1471, n4378,
         g21880, g2877, g19154, g813, n4289, g19163, g809, n4567, g19173, g805,
         n4559, g19184, g801, n4327, g20310, g797, n4391, g20343, g793, n4321,
         g20376, g789, n4375, g20417, g785, n4379, g21878, g2873, g19153, g125,
         n4290, g19162, g121, n4569, g19172, g117, n4561, g19144, g113, n4328,
         g19149, g109, n4392, g19157, g105, n4322, g19167, g101, n4376, g19178,
         g97, n4380, g20874, g2857, g18885, g2200, n4287, g18975, g2195, n4563,
         g18968, g2190, n4555, g18942, g2185, n4325, g18906, g2180, n4389,
         g18867, g2175, n4319, g18836, g2170, n4373, g18957, g2165, n4377,
         g21882, g2878, n4598, n4382, n4383, g3109, n4494, g18669, g18719,
         g3211, g18782, g3084, n4445, g17222, g3085, g17225, g3086, g17234,
         g3087, n4344, g17224, g3091, n4448, g17228, g3092, n4451, g17246,
         g3093, g17226, g3094, g17235, g3095, g17269, g3096, g25450, g3097,
         g25451, g3098, g25452, g3099, n4443, g28420, g3100, n4342, g28421,
         g28425, g3102, n4343, g29936, g3103, n4447, g29939, g3104, n4452,
         g29941, g3105, g30796, g3106, n4438, g30798, g3107, g30801, g3108,
         n4334, g17229, g3155, g17247, g3158, g17302, g3161, n4444, g17236,
         g3164, g17270, g3167, g17340, g3170, n4441, g17248, g3173, n4338,
         g17303, g3176, n4450, g17383, g17271, g3182, g17341, g3185, g17429,
         g3088, n8090, DFF_131_n1, n8089, DFF_132_n1, g3197, n8088, DFF_134_n1,
         g3201, n4406, g3204, g3207, n4329, g3188, n4405, g3133, n8087,
         DFF_140_n1, g3128, n8086, n8084, DFF_144_n1, g3124, n8083, DFF_146_n1,
         n8082, n8081, n8080, DFF_149_n1, g3112, g3110, g3111, n8079, n8078,
         n8077, DFF_155_n1, n8076, DFF_156_n1, g3151, n4424, g3142, n4301,
         g185, n4318, n4512, g165, n4369, g22100, g130, g22122, g131, g22141,
         g129, g22123, g133, g22142, g134, g22161, g132, g22025, g142, g22027,
         g143, g22030, g141, g22028, g145, g22031, g146, g22037, g22032, g148,
         g22038, g149, g22047, g147, g22039, g151, g22048, g152, g22063, g150,
         g22049, g154, g22064, g155, g22079, g153, g22065, g157, g22080, g158,
         g22101, g156, g22081, g160, g22102, g161, g22124, g159, g22103,
         g22125, g164, g22143, g162, g25204, g169, g25206, g170, g25211, g168,
         g25207, g172, g25212, g173, g25218, g171, g25213, g175, g25219, g176,
         g25228, g174, g25220, g178, g25229, g179, g25239, g177, g30261, g186,
         g30267, g30275, g192, g30637, g231, g30640, g234, g30645, g237,
         g30668, g195, g30674, g198, g30680, g201, g30641, g240, g30646, g243,
         g30653, g246, g30276, g204, g30284, g207, g30292, g210, g30254, g249,
         g30257, g252, g30262, g30245, g213, g30246, g216, g30248, g219,
         g30258, g258, g30263, g261, g30268, g264, g30635, g222, g30636, g225,
         g30639, g228, g30661, g267, g30669, g270, g30675, g273, g25027, g92,
         g25932, g88, g26529, g83, g27120, g27594, g74, g28145, g70, g28634,
         g65, g29109, g61, g29353, g29579, g52, g180, g181, n4506, g309, n4388,
         g27253, g354, g27255, g343, g27258, g27256, g369, g27259, g358,
         g27265, g361, g27260, g384, g27266, g373, g27277, g376, g27267, g398,
         g27278, g388, g27293, g391, g28732, g408, g28735, g411, g28744, g414,
         g29194, g417, g29197, g420, g29201, g423, g28736, g28745, g428,
         g28754, g426, g26803, g429, g26804, g432, g26807, g435, g26805, g438,
         g26808, g441, g26812, g444, g27759, g448, g27760, g449, g27762, g447,
         g29606, g312, g29608, g313, g29611, g314, g30699, g315, g30700,
         g30702, g317, g30455, g318, g30468, g319, g30482, g320, g29167, g322,
         g29169, g323, g29172, g321, g26655, g403, g26659, g404, g26664, g402,
         g450, n8066, DFF_299_n1, g452, n8065, DFF_301_n1, g454, DFF_303_n1,
         g280, n8062, DFF_305_n1, g282, n8061, DFF_307_n1, g284, n8060,
         DFF_309_n1, g286, n8059, DFF_311_n1, g288, n8058, DFF_313_n1, g290,
         n8057, n4485, n4282, n8056, g21346, g305, n4278, n8055, DFF_328_n1,
         g349, g350, g351, g352, g353, g357, g364, g365, g366, g367, g368,
         g372, g379, g380, g381, g383, g387, g394, g395, g396, g397, g324,
         g337, n4298, n4372, g550, n4313, g554, g18678, g557, n4360, g18726,
         g513, g523, g524, g455, g564, g569, g458, g570, g571, g461, g572,
         g573, g465, g574, g565, g566, g567, g471, g568, g489, n4461, g485,
         n4466, g23067, g486, g23093, g487, g23117, g488, g23385, g23399,
         g24174, g24178, g477, g24207, g478, g24216, g479, g23092, g480,
         g23000, g484, g23022, g464, g24206, g24215, g24228, g528, g535, g542,
         g13149, g543, g544, g21851, g548, g13111, g549, g499, n4541, g13160,
         g558, g559, g27261, g576, g27268, g577, g27279, g575, g27269, g579,
         g27280, g27294, g578, g27281, g582, g27295, g583, g27311, g581,
         g27296, g585, g27312, g586, g27327, g584, g24491, g587, g24498, g590,
         g24507, g593, g24499, g596, g24508, g599, g24519, g602, g28345, g614,
         g28349, g617, g28353, g28342, g605, g28344, g608, g28348, g611,
         g26541, g490, g26545, g493, g26553, g496, g506, n4570, g22578, n4571,
         g525, n8047, DFF_444_n1, n8046, DFF_445_n1, n8045, DFF_446_n1, n8044,
         DFF_447_n1, n8043, DFF_448_n1, DFF_449_n1, g536, g537, g24059, g538,
         n4492, n8040, n4359, g629, n4295, g16654, g630, g20314, g659, n4429,
         g20682, g640, n4404, g633, n4478, g23324, g653, n4422, g24426, g646,
         n4414, g25185, g660, n4403, g672, n4413, g26776, g27672, g679, n4477,
         g28199, g686, n4396, g28668, g692, n4418, g20875, g699, g20879, g700,
         g20891, g698, g20880, g702, g20892, g703, g20901, g701, g20893, g705,
         g20902, g706, g20921, g704, g20903, g708, g20922, g709, g20944, g707,
         g20923, g20945, g712, g20966, g710, g20946, g714, g20967, g715,
         g20989, g713, g20968, g717, g20990, g718, g21009, g716, g20991, g720,
         g21010, g721, g21031, g719, g21011, g723, g21032, g724, g21051, g722,
         g20876, g726, g20881, g20894, g725, g20924, g729, g20947, g730,
         g20969, g728, g20948, g732, g20970, g733, g20992, g731, g25260, g735,
         g25262, g736, g25266, g734, g22218, g738, g739, g22242, g737, n4323,
         n4312, g22126, g818, g22145, g819, g22162, g817, g22146, g821, g22163,
         g822, g22177, g820, g22029, g830, g22033, g831, g22040, g829, g22034,
         g833, g22041, g834, g22054, g832, g22042, g836, g22055, g837, g22066,
         g835, g22056, g22067, g840, g22087, g838, g22068, g842, g22088, g843,
         g22104, g841, g22089, g845, g22105, g846, g22127, g844, g22106, g848,
         g22128, g849, g22147, g847, g22129, g851, g22148, g852, g22164, g850,
         g25209, g857, g25214, g25221, g856, g25215, g860, g25222, g861,
         g25230, g859, g25223, g863, g25231, g864, g25240, g862, g25232, g866,
         g25241, g867, g25248, g865, g30269, g873, g30277, g876, g30285, g879,
         g30643, g918, g30648, g921, g30654, g30676, g882, g30681, g885,
         g30687, g888, g30649, g927, g30655, g930, g30662, g933, g30286, g891,
         g30293, g894, g30298, g897, g30259, g936, g30264, g939, g30270, g942,
         g30247, g900, g30249, g903, g30251, g906, g30265, g30271, g948,
         g30278, g951, g30638, g909, g30642, g912, g30647, g915, g30670, g954,
         g30677, g957, g30682, g960, g25042, g780, g25935, g776, g26530, g771,
         g27123, g767, g27603, g762, g28146, g758, g28635, g753, g29110,
         g29354, g29580, g740, g868, g869, n4363, n4364, g1088, n4381, g996,
         n4387, g27257, g1041, g27262, g1030, g27270, g1033, g27263, g1056,
         g27271, g1045, g27282, g1048, g27272, g27283, g1060, g27297, g1063,
         g27284, g1085, g27298, g1075, g27313, g1078, g28738, g1095, g28746,
         g1098, g28758, g1101, g29198, g1104, g29204, g1107, g29209, g1110,
         g28747, g1114, g28759, g1115, g28767, g1113, g26806, g1116, g26809,
         g26813, g1122, g26810, g1125, g26814, g1128, g26818, g1131, g27761,
         g1135, g27763, g1136, g27765, g1134, g29609, g999, g29612, g1000,
         g29616, g1001, g30701, g1002, g30703, g1003, g30705, g1004, g30470,
         g1005, g30485, g1006, g30500, g29170, g1009, g29173, g1010, g29179,
         g1008, g26661, g1090, g26665, g1091, g26669, g1089, g1137, n8027,
         DFF_649_n1, g1139, n8026, DFF_651_n1, g1141, n8025, DFF_653_n1, g967,
         n8024, DFF_655_n1, g969, DFF_657_n1, g971, n8021, DFF_659_n1, g973,
         n8020, DFF_661_n1, g975, n8019, DFF_663_n1, g977, n8018, n4486, n4283,
         g986, n4432, g992, n4277, n8017, g1029, g1036, g1037, g1038, g1040,
         g1044, g1051, g1052, g1053, g1054, g1055, g1059, g1066, g1067, g1068,
         g1069, g1070, g1074, g1081, g1083, g1084, g1011, g1024, n4371, n4316,
         g1236, n4300, g1240, g18707, g1243, n4353, g18763, g1196, n4304,
         g1199, g1209, g1210, g1142, g1255, g1145, g1256, g1257, g1148, g1258,
         g1259, g1152, g1260, g1251, g1155, g1252, g1253, g1158, g1254, g1176,
         n4460, n4459, g1172, n4465, g23081, g1173, g23111, g23126, g1175,
         g23392, g23406, g24179, g24181, g1164, g24213, g1165, g24223, g1166,
         g23110, g1167, g23014, g1171, g23039, g1151, g24212, g24222, g24235,
         g1214, g1221, g13155, g1229, n4549, n4361, g13124, g1235, g1186,
         n4548, g13171, g1244, g1245, g27273, g1262, g27285, g1263, g27299,
         g1261, g27286, g1265, g27300, g1266, g27314, g1264, g27301, g1268,
         g27315, g1269, g27328, g27316, g1271, g27329, g1272, g27339, g1270,
         g24501, g1273, g24510, g1276, g24521, g1279, g24511, g1282, g24522,
         g1285, g24532, g1288, g28351, g1300, g28355, g1303, g28360, g1306,
         g28346, g1291, g28350, g1294, g28354, g1297, g26547, g26557, g1180,
         g26569, g1183, g1192, n4454, g22615, n8009, DFF_783_n1, DFF_792_n1,
         g1211, n8008, DFF_794_n1, n8007, DFF_795_n1, n8006, DFF_796_n1, n8005,
         DFF_797_n1, n8004, DFF_798_n1, n8003, DFF_799_n1, g1222, g1223,
         g24072, g1224, n4489, n4358, g1315, n4294, g16671, g1316, g20333,
         g1345, n4428, g20717, g1326, n4402, g1319, n4476, g23329, g1339,
         n4421, g24430, g1332, n4412, g25189, g1346, n4401, g1358, n4411,
         g26781, g1352, n4469, g27678, g1365, n4475, g27718, g1372, n4395,
         g28321, g1378, n4417, g20882, g20896, g1386, g20910, g1384, g20897,
         g1388, g20911, g1389, g20925, g1387, g20912, g1391, g20926, g1392,
         g20949, g1390, g20927, g1394, g20950, g1395, g20972, g1393, g20951,
         g1397, g20973, g1398, g20993, g1396, g20974, g1400, g20994, g21015,
         g1399, g20995, g1403, g21016, g1404, g21033, g1402, g21017, g1406,
         g21034, g1407, g21052, g1405, g21035, g1409, g21053, g1410, g21070,
         g1408, g20883, g1412, g20898, g1413, g20913, g1411, g20952, g1415,
         g20975, g1416, g20996, g20976, g1418, g20997, g1419, g21018, g1417,
         g25263, g1421, g25267, g1422, g25270, g1420, g22234, g1424, g1425,
         g22263, g1423, n4317, n4515, g1547, n4368, g22149, g1512, g22166,
         g1513, g22178, g1511, g22167, g22179, g1516, g22191, g1514, g22035,
         g1524, g22043, g1525, g22057, g1523, g22044, g1527, g22058, g1528,
         g22073, g1526, g22059, g1530, g22074, g1531, g22090, g1529, g22075,
         g1533, g22091, g1534, g22112, g1532, g22092, g1536, g22113, g22130,
         g1535, g22114, g1539, g22131, g1540, g22150, g1538, g22132, g1542,
         g22151, g1543, g22168, g1541, g22152, g1545, g22169, g1546, g22180,
         g1544, g25217, g1551, g25224, g1552, g25233, g1550, g25225, g1554,
         g25234, g1555, g25242, g25235, g1557, g25243, g1558, g25249, g1556,
         g25244, g1560, g25250, g1561, g25255, g1559, g30279, g1567, g30287,
         g1570, g30294, g1573, g30651, g1612, g30657, g1615, g30663, g1618,
         g30683, g1576, g30688, g1579, g30692, g1582, g30658, g30664, g1624,
         g30671, g1627, g30295, g1585, g30299, g1588, g30302, g1591, g30266,
         g1630, g30272, g1633, g30280, g1636, g30250, g1594, g30252, g1597,
         g30255, g1600, g30273, g1639, g30281, g1642, g30288, g1645, g30644,
         g1603, g30650, g30656, g1609, g30678, g1648, g30684, g1651, g30689,
         g1654, g25056, g1466, g25938, g1462, g26531, g1457, g27129, g1453,
         g27612, g1448, g28147, g1444, g28636, g1439, g29111, g1435, g29355,
         g29581, g1426, g1562, g1563, n4518, g1690, n4386, g27264, g1735,
         g27274, g1724, g27287, g1727, g27275, g1750, g27288, g1739, g27302,
         g1742, g27289, g1765, g27303, g1754, g27317, g1757, g27304, g1779,
         g27318, g27330, g1772, g28749, g1789, g28760, g1792, g28771, g1795,
         g29205, g1798, g29212, g1801, g29218, g1804, g28761, g1808, g28772,
         g1809, g28778, g1807, g26811, g1810, g26815, g1813, g26820, g1816,
         g26816, g1819, g26821, g1822, g26824, g27764, g1829, g27766, g1830,
         g27768, g1828, g29613, g1693, g29617, g1694, g29620, g1695, g30704,
         g1696, g30706, g1697, g30708, g1698, g30487, g1699, g30503, g1700,
         g30338, g1701, g29178, g1703, g29181, g1704, g29184, g1702, g26667,
         g26670, g1785, g26675, g1783, g1831, n7988, DFF_999_n1, g1833, n7987,
         DFF_1001_n1, g1835, n7986, DFF_1003_n1, g1661, n7985, DFF_1005_n1,
         g1663, n7984, DFF_1007_n1, g1665, n7983, DFF_1009_n1, g1667,
         DFF_1011_n1, g1669, n7980, DFF_1013_n1, g1671, n7979, n4484, n4284,
         g1680, n4488, g1686, n4276, n7978, g1723, g1730, g1731, g1732, g1733,
         g1734, g1738, g1745, g1747, g1748, g1749, g1753, g1760, g1761, g1762,
         g1763, g1764, g1768, g1775, g1776, g1777, g1778, g1705, g1718, n4296,
         n4315, g1930, n4366, g1934, g18743, g1937, n4311, g18794, g1890,
         n4297, g1893, g1903, g1904, g1836, g1944, g1949, g1950, g1951, g1842,
         g1953, g1846, g1954, g1945, g1849, g1946, g1947, g1852, g1948, g1870,
         n4458, n4457, g1866, n4464, g23097, g1867, g23124, g1868, g23137,
         g1869, g23400, g23413, g24182, g24208, g1858, g24219, g1859, g24231,
         g1860, g23123, g1861, g23030, g1865, g23058, g1845, g24218, g24230,
         g24243, g1908, g1915, g1922, g13164, g1923, DFF_1099_n1, n7971,
         g13135, g1929, g1880, n4545, g13182, g1938, g1939, g27290, g1956,
         g27305, g1957, g27319, g1955, g27306, g1959, g27320, g1960, g27331,
         g1958, g27321, g1962, g27332, g1963, g27340, g1961, g27333, g27341,
         g1966, g27346, g1964, g24513, g1967, g24524, g1970, g24534, g1973,
         g24525, g1976, g24535, g1979, g24545, g1982, g28357, g1994, g28362,
         g1997, g28366, g2000, g28352, g1985, g28356, g1988, g28361, g1991,
         g26559, g26573, g1874, g26592, g1877, g1886, n4493, g22651, n7968,
         DFF_1133_n1, DFF_1142_n1, g1905, n7967, DFF_1144_n1, n7966,
         DFF_1145_n1, n7965, DFF_1146_n1, n7964, DFF_1147_n1, n7963,
         DFF_1148_n1, n7962, DFF_1149_n1, g1916, g1917, g24083, n7960, n4357,
         g2009, n4293, g16692, g2010, g20353, g2039, n4427, g20752, g2020,
         n4400, g2013, n4474, g23339, g2033, n4420, g24434, g2026, n4410,
         g25194, g2040, n4399, g2052, n4409, g26789, g2046, n4468, g27682,
         g2059, n4473, g27722, g28325, g2072, n4416, g20899, g2079, g20915,
         g2080, g20934, g2078, g20916, g2082, g20935, g2083, g20953, g2081,
         g20936, g2085, g20954, g2086, g20977, g2084, g20955, g2088, g20978,
         g2089, g20999, g2087, g20979, g2091, g21000, g21019, g2090, g21001,
         g2094, g21020, g2095, g21039, g2093, g21021, g2097, g21040, g2098,
         g21054, g2096, g21041, g2100, g21055, g2101, g21071, g2099, g21056,
         g2103, g21072, g2104, g21080, g2102, g20900, g2106, g20917, g20937,
         g2105, g20980, g2109, g21002, g2110, g21022, g2108, g21003, g2112,
         g21023, g2113, g21042, g2111, g25268, g2115, g25271, g2116, g25279,
         g2114, g22249, g2118, g2119, g22280, g2117, n4324, g2241, n4367,
         g22170, g2206, g22182, g2207, g22192, g2205, g22183, g2209, g22193,
         g2210, g22200, g2208, g22045, g2218, g22060, g2219, g22076, g2217,
         g22061, g2221, g22077, g2222, g22097, g2220, g22078, g2224, g22098,
         g22115, g2223, g22099, g2227, g22116, g2228, g22138, g2226, g22117,
         g2230, g22139, g2231, g22153, g2229, g22140, g2233, g22154, g2234,
         g22171, g2232, g22155, g2236, g22172, g2237, g22184, g2235, g22173,
         g2239, g22185, g22194, g2238, g25227, g2245, g25236, g2246, g25245,
         g2244, g25237, g2248, g25246, g2249, g25251, g2247, g25247, g2251,
         g25252, g2252, g25256, g2250, g25253, g2254, g25257, g2255, g25259,
         g2253, g30289, g2261, g30296, g30300, g2267, g30660, g2306, g30666,
         g2309, g30672, g2312, g30690, g2270, g30693, g2273, g30695, g2276,
         g30667, g2315, g30673, g2318, g30679, g2321, g30301, g2279, g30303,
         g2282, g30304, g2285, g30274, g2324, g30282, g30290, g2330, g30253,
         g2288, g30256, g2291, g30260, g2294, g30283, g2333, g30291, g2336,
         g30297, g2339, g30652, g2297, g30659, g2300, g30665, g2303, g30686,
         g2342, g30691, g2345, g30694, g2348, g25067, g2160, g25940, g26532,
         g2151, g27131, g2147, g27621, g2142, g28148, g2138, g28637, g2133,
         g29112, g2129, g29357, g29582, g2120, g2256, g2257, n4516, g27276,
         g2429, g27291, g2418, g27307, g2421, g27292, g2444, g27308, g2433,
         g27322, g2436, g27309, g2459, g27323, g2448, g27334, g2451, g27324,
         g2473, g27335, g2463, g27342, g2466, g28763, g2483, g28773, g2486,
         g28782, g29213, g2492, g29221, g2495, g29226, g2498, g28774, g2502,
         g28783, g2503, g28788, g2501, g26817, g2504, g26822, g2507, g26825,
         g2510, g26823, g2513, g26826, g2516, g26827, g2519, g27767, g2523,
         g27769, g2524, g27771, g29618, g2387, g29621, g2388, g29623, g2389,
         g30707, g2390, g30709, g2391, g30566, g2392, g30505, g2393, g30341,
         g2394, g30356, g2395, g29182, g2397, g29185, g2398, g29187, g2396,
         g26672, g2478, g26676, g2479, g26025, g2525, n7946, DFF_1349_n1,
         g2527, n7945, DFF_1351_n1, g2529, n7944, DFF_1353_n1, g2355, n7943,
         DFF_1355_n1, g2357, n7942, DFF_1357_n1, g2359, n7941, DFF_1359_n1,
         g2361, n7940, DFF_1361_n1, n7938, DFF_1363_n1, g2365, n7937, n4483,
         n4285, g2374, n4487, g30055, g2380, n4275, n7936, DFF_1378_n1, g2417,
         g2424, g2425, g2426, g2427, g2428, g2432, g2439, g2441, g2442, g2443,
         g2447, g2454, g2455, g2456, g2457, g2458, g2462, g2469, g2470, g2471,
         g2472, g2412, n4314, n4370, g2624, n4299, g2628, g18780, g2631, n4352,
         g18820, g2584, n4303, g2587, g2597, g2598, g2530, g2638, g2643, g2533,
         g2645, g2536, g2646, g2647, g2540, g2648, g2639, g2543, g2640, g2641,
         g2546, g2642, g2564, n4456, n4455, g2560, n4463, g23114, g2561,
         g23133, g2562, g21970, g23407, g23418, g24209, g24214, g2552, g24226,
         g2553, g24238, g2554, g23132, g2555, g23047, g2559, g23076, g2539,
         g24225, g24237, g24250, g2602, g2609, g13175, g2617, n7930, g30072,
         n7929, g13143, g2623, g2574, n4543, g13194, g2632, g2633, g27310,
         g2650, g27325, g2651, g27336, g2649, g27326, g2653, g27337, g2654,
         g27343, g2652, g27338, g2656, g27344, g27347, g2655, g27345, g2659,
         g27348, g2660, g27354, g2658, g24527, g2661, g24537, g2664, g24547,
         g2667, g24538, g2670, g24548, g2673, g24557, g2676, g28364, g2688,
         g28368, g2691, g28371, g2694, g28358, g2679, g28363, g28367, g2685,
         g26575, g2565, g26596, g2568, g26616, g2571, g2580, g22687, n7926,
         g30061, g2599, n7925, DFF_1494_n1, n7924, DFF_1495_n1, n7923,
         DFF_1496_n1, n7922, DFF_1497_n1, n7921, DFF_1498_n1, n7920,
         DFF_1499_n1, g2611, g24092, g2612, n4490, n7918, g2703, n4292, g16718,
         g2704, g20375, g2733, n4426, g20789, g2714, n4398, g2707, n4472,
         g23348, g2727, n4419, g24438, g2720, n4408, g25197, g2734, n4397,
         g2746, n4407, g26795, g27243, g2753, n4471, g27724, g2760, n4393,
         g28328, g2766, n4415, g20918, g2773, g20939, g2774, g20962, g2772,
         g20940, g2776, g20963, g2777, g20981, g2775, g20964, g2779, g20982,
         g2780, g21004, g2778, g20983, g2782, g21005, g2783, g21025, g21006,
         g2785, g21026, g2786, g21043, g2784, g21027, g2788, g21044, g2789,
         g21060, g2787, g21045, g2791, g21061, g2792, g21073, g2790, g21062,
         g2794, g21074, g2795, g21081, g2793, g21075, g2797, g21082, g2798,
         g21094, g20919, g2800, g20941, g2801, g20965, g2799, g21007, g2803,
         g21028, g2804, g21046, g2802, g21029, g2806, g21047, g2807, g21063,
         g2805, g25272, g2809, g25280, g2810, g25288, g2808, g22269, g2812,
         g22284, g2813, g22299, g20877, n7913, DFF_1561_n1, g20884, n7912,
         DFF_1562_n1, n4263_Tj_Payload, n4269, g3043, n4268, g3044, n4267,
         g3045, n4266, g3046, n4265, g3047, n4272, g3048, n4271, g3049, n4270,
         g3050, n4259, g3051, n4236, g3052, n4239, g3053, n4237, n4234, g3056,
         n4233, g3057, n4238, g3058, n4235, g3059, n4240, g3060, n4232, g3061,
         n4245, g3062, n4248, g3063, n4246, g3064, n4243, g3065, n4242, g3066,
         n4247, g3067, n4244, g3068, n4249, g3069, n4241, n4254, g3071, n4257,
         g3072, n4255, g3073, n4252, g3074, n4251, g3075, n4256, g3076, n4253,
         g3077, n4258, g3078, n4250, g2997, g25265, g2993, g26048, n7909,
         g3006, g24445, g3002, g25191, g3013, g26031, g26786, g3024, n4262,
         g3018, n4481, g3028, n4350, g24446, g3036, n4480, g25202, g3032,
         n7907, DFF_1612_n1, g2987, n4365, g16824, g16844, g16853, g16860,
         g16803, g16835, g16851, g16857, g16866, g3083, n4261, N995, n4577,
         g16845, g16854, g16861, g16880, g18755, g18804, g18837, g18868,
         g18907, g2990, N690, n4578, n4260, n4309, n4308, n4307, n4306, n4524,
         n4525, n4511, n4509, n4499, n4520, n3683, n3887, n3686, n3890, n3692,
         n3896, n4513, n3897, n3424, n3427, n3433, n4529, n4530, n4522, n4523,
         n4521, n3171, n3159, n3163, n3893, n3690, n3689, n3431, n3430, n3168,
         n3160, n3164, n3172, n4527, n4528, n4526, n3167, n3894, n3888, n3891,
         n2302, n2289, n2303, n2275, n4066, n4065, n4606, n4618, n4640, n2351,
         n2430, n2792, n2632, n3936, n3252, n3254, n3038, n3070, n3102, n3130,
         n3036, n3068, n3128, n2800, n2798, n2616, n2594, n3940, n3705, n3933,
         n3939, n3016, n3000, n3008, n3023, n3700, n4058, n4101, n3938, n4182,
         n4073, n4057, n4122, n4263, Tj_OUT1, Tj_OUT2, Tj_OUT3, Tj_OUT4,
         Tj_OUT1234, Tj_OUT5, Tj_OUT6, Tj_OUT7, Tj_OUT8, Tj_OUT5678,
         Tj_Trigger, n10, n15, n102, n123, n155, n162, n163, n184, n223, n263,
         n285, n289, n298, n328, n456, n457, n472, n494, n516, n517, n518,
         n531, n532, n533, n534, n539, n586, n615, n616, n672, n819, n833,
         n837, n883, n912, n913, n971, n1122, n1145, n1149, n1194, n1222,
         n1223, n1269, n1396, n1406, n1427, n1431, n1506, n1507, n1542, n1544,
         n1547, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7418,
         n7441, n7442, n7443, n7444, n7445, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7627, n7629, n7630, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7717, n7718, n7719, n7720,
         n7721, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7908, n7910, n7911, n7914, n7915, n7916, n7917, n7919,
         n7927, n7928, n7931, n7932, n7933, n7934, n7935, n7939, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7961, n7969, n7970, n7972, n7973, n7974, n7975, n7976, n7977,
         n7981, n7982, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8010, n8012, n8013, n8014,
         n8015, n8016, n8022, n8023, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8041, n8042, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8063, n8064, n8067, n8069, n8070, n8071,
         n8072, n8073, n8075, n8085, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8100, n8101, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, U3772_n1, U3776_n1, U3777_n1, U3778_n1, U3779_n1,
         U3780_n1, U3781_n1, U3782_n1, U3783_n1, U3784_n1, U3785_n1, U3786_n1,
         U3787_n1, U3901_n1, U3902_n1, U4467_n1, U4904_n1, U4930_n1, U5128_n1,
         U5141_n1, U5749_n1, U5750_n1, U5751_n1, U5752_n1, U5753_n1, U5754_n1,
         U5755_n1, U5756_n1, U5757_n1, U5758_n1, U5759_n1, U5760_n1, U5761_n1,
         U5762_n1, U5763_n1, U5764_n1, U5882_n1, U5939_n1, U5940_n1, U5941_n1,
         U5942_n1, U6140_n1, U6460_n1, U6470_n1, U6562_n1, U6563_n1, U6718_n1,
         U7116_n1, U7118_n1, U7293_n1;
  assign g8251 = test_so3;
  assign g7519 = test_so4;
  assign g4450 = test_so5;
  assign g7909 = test_so23;
  assign g5612 = test_so57;
  assign g5695 = test_so63;
  assign g7084 = test_so73;
  assign g8270 = test_so99;
  assign g8258 = test_so100;

  SDFFX1 DFF_0_Q_reg ( .D(g51), .SI(test_si1), .SE(n8144), .CLK(n8331), .Q(
        n8104), .QN(n14383) );
  SDFFX1 DFF_1_Q_reg ( .D(g16802), .SI(n8104), .SE(n8144), .CLK(n8331), .Q(
        n8103), .QN(DFF_1_n1) );
  SDFFX1 DFF_2_Q_reg ( .D(g16823), .SI(n8103), .SE(n8144), .CLK(n8331), .Q(
        n8102), .QN(DFF_2_n1) );
  SDFFX1 DFF_3_Q_reg ( .D(n4264), .SI(n8102), .SE(n8144), .CLK(n8331), .Q(
        g2950), .QN(n4423) );
  SDFFX1 DFF_4_Q_reg ( .D(n4274), .SI(g2950), .SE(n8145), .CLK(n8332), .Q(
        g2883), .QN(n4330) );
  SDFFX1 DFF_5_Q_reg ( .D(g22026), .SI(g2883), .SE(n8145), .CLK(n8332), .Q(
        g2888), .QN(n8037) );
  SDFFX1 DFF_6_Q_reg ( .D(g23358), .SI(g2888), .SE(n8145), .CLK(n8332), .Q(
        g2896), .QN(n4431) );
  SDFFX1 DFF_7_Q_reg ( .D(g24473), .SI(g2896), .SE(n8145), .CLK(n8332), .Q(
        g2892), .QN(n7764) );
  SDFFX1 DFF_8_Q_reg ( .D(g25201), .SI(g2892), .SE(n8145), .CLK(n8332), .Q(
        g2903), .QN(n4305) );
  SDFFX1 DFF_9_Q_reg ( .D(g26037), .SI(g2903), .SE(n8145), .CLK(n8332), .Q(
        g2900), .QN(n4291) );
  SDFFX1 DFF_10_Q_reg ( .D(g26798), .SI(g2900), .SE(n8145), .CLK(n8332), .Q(
        g2908), .QN(n4355) );
  SDFFX1 DFF_11_Q_reg ( .D(n4273), .SI(g2908), .SE(n8145), .CLK(n8332), .Q(
        g2912), .QN(n4482) );
  SDFFX1 DFF_12_Q_reg ( .D(g23357), .SI(g2912), .SE(n8145), .CLK(n8332), .Q(
        g2917), .QN(n4479) );
  SDFFX1 DFF_13_Q_reg ( .D(g24476), .SI(g2917), .SE(n8145), .CLK(n8332), .Q(
        g2924), .QN(n4349) );
  SDFFX1 DFF_14_Q_reg ( .D(g25199), .SI(g2924), .SE(n8145), .CLK(n8332), .Q(
        g2920), .QN(n7715) );
  SDFFX1 DFF_15_Q_reg ( .D(n4280), .SI(g2920), .SE(n8145), .CLK(n8332), .Q(
        test_so1), .QN(DFF_15_n1) );
  SDFFX1 DFF_16_Q_reg ( .D(n4281), .SI(test_si2), .SE(n8142), .CLK(n8329), .Q(
        n8099), .QN(DFF_16_n1) );
  SDFFX1 DFF_17_Q_reg ( .D(g51), .SI(n8099), .SE(n8142), .CLK(n8329), .Q(g8021) );
  SDFFX1 DFF_18_Q_reg ( .D(g8021), .SI(g8021), .SE(n8142), .CLK(n8329), .Q(
        n8098), .QN(DFF_18_n1) );
  SDFFX1 DFF_19_Q_reg ( .D(n4279), .SI(n8098), .SE(n8142), .CLK(n8329), .Q(
        g2879), .QN(n4351) );
  SDFFX1 DFF_20_Q_reg ( .D(g3212), .SI(g2879), .SE(n8142), .CLK(n8329), .Q(
        g2934), .QN(n8035) );
  SDFFX1 DFF_21_Q_reg ( .D(g3228), .SI(g2934), .SE(n8142), .CLK(n8329), .Q(
        g2935), .QN(n8000) );
  SDFFX1 DFF_22_Q_reg ( .D(g3227), .SI(g2935), .SE(n8143), .CLK(n8330), .Q(
        g2938), .QN(n8001) );
  SDFFX1 DFF_23_Q_reg ( .D(g3226), .SI(g2938), .SE(n8143), .CLK(n8330), .Q(
        g2941), .QN(n7998) );
  SDFFX1 DFF_24_Q_reg ( .D(g3225), .SI(g2941), .SE(n8143), .CLK(n8330), .Q(
        g2944) );
  SDFFX1 DFF_25_Q_reg ( .D(g3224), .SI(g2944), .SE(n8143), .CLK(n8330), .Q(
        g2947), .QN(n8002) );
  SDFFX1 DFF_26_Q_reg ( .D(g3223), .SI(g2947), .SE(n8143), .CLK(n8330), .Q(
        g2953), .QN(n8010) );
  SDFFX1 DFF_27_Q_reg ( .D(g3222), .SI(g2953), .SE(n8143), .CLK(n8330), .Q(
        g2956), .QN(n8012) );
  SDFFX1 DFF_28_Q_reg ( .D(g3221), .SI(g2956), .SE(n8143), .CLK(n8330), .Q(
        g2959), .QN(n7999) );
  SDFFX1 DFF_29_Q_reg ( .D(g3232), .SI(g2959), .SE(n8143), .CLK(n8330), .Q(
        g2962), .QN(n8033) );
  SDFFX1 DFF_30_Q_reg ( .D(g3220), .SI(g2962), .SE(n8143), .CLK(n8330), .Q(
        g2963), .QN(n8015) );
  SDFFX1 DFF_31_Q_reg ( .D(g3219), .SI(g2963), .SE(n8143), .CLK(n8330), .Q(
        test_so2) );
  SDFFX1 DFF_32_Q_reg ( .D(g3218), .SI(test_si3), .SE(n8142), .CLK(n8329), .Q(
        g2969), .QN(n8023) );
  SDFFX1 DFF_33_Q_reg ( .D(g3217), .SI(g2969), .SE(n8142), .CLK(n8329), .Q(
        g2972), .QN(n8016) );
  SDFFX1 DFF_34_Q_reg ( .D(g3216), .SI(g2972), .SE(n8142), .CLK(n8329), .Q(
        g2975), .QN(n8022) );
  SDFFX1 DFF_35_Q_reg ( .D(g3215), .SI(g2975), .SE(n8142), .CLK(n8329), .Q(
        g2978), .QN(n8013) );
  SDFFX1 DFF_36_Q_reg ( .D(g3214), .SI(g2978), .SE(n8142), .CLK(n8329), .Q(
        g2981) );
  SDFFX1 DFF_37_Q_reg ( .D(g3213), .SI(g2981), .SE(n8142), .CLK(n8329), .Q(
        g2874), .QN(n8014) );
  SDFFX1 DFF_38_Q_reg ( .D(g18754), .SI(g2874), .SE(n8143), .CLK(n8330), .Q(
        g1506), .QN(n4288) );
  SDFFX1 DFF_39_Q_reg ( .D(g18781), .SI(g1506), .SE(n8143), .CLK(n8330), .Q(
        g1501), .QN(n4565) );
  SDFFX1 DFF_40_Q_reg ( .D(g18803), .SI(g1501), .SE(n8144), .CLK(n8331), .Q(
        g1496), .QN(n4557) );
  SDFFX1 DFF_41_Q_reg ( .D(g18821), .SI(g1496), .SE(n8144), .CLK(n8331), .Q(
        g1491), .QN(n4326) );
  SDFFX1 DFF_42_Q_reg ( .D(g18835), .SI(g1491), .SE(n8144), .CLK(n8331), .Q(
        g1486), .QN(n4390) );
  SDFFX1 DFF_43_Q_reg ( .D(g18852), .SI(g1486), .SE(n8144), .CLK(n8331), .Q(
        g1481), .QN(n4320) );
  SDFFX1 DFF_44_Q_reg ( .D(g18866), .SI(g1481), .SE(n8144), .CLK(n8331), .Q(
        g1476), .QN(n4374) );
  SDFFX1 DFF_45_Q_reg ( .D(g18883), .SI(g1476), .SE(n8144), .CLK(n8331), .Q(
        g1471), .QN(n4378) );
  SDFFX1 DFF_46_Q_reg ( .D(g21880), .SI(g1471), .SE(n8149), .CLK(n8336), .Q(
        g2877) );
  SDFFX1 DFF_47_Q_reg ( .D(g19154), .SI(g2877), .SE(n8149), .CLK(n8336), .Q(
        test_so3) );
  SDFFX1 DFF_48_Q_reg ( .D(test_so3), .SI(test_si4), .SE(n8149), .CLK(n8336), 
        .Q(g813), .QN(n4289) );
  SDFFX1 DFF_49_Q_reg ( .D(g19163), .SI(g813), .SE(n8149), .CLK(n8336), .Q(
        g4090) );
  SDFFX1 DFF_50_Q_reg ( .D(g4090), .SI(g4090), .SE(n8149), .CLK(n8336), .Q(
        g809), .QN(n4567) );
  SDFFX1 DFF_51_Q_reg ( .D(g19173), .SI(g809), .SE(n8149), .CLK(n8336), .Q(
        g4323) );
  SDFFX1 DFF_52_Q_reg ( .D(g4323), .SI(g4323), .SE(n8149), .CLK(n8336), .Q(
        g805), .QN(n4559) );
  SDFFX1 DFF_53_Q_reg ( .D(g19184), .SI(g805), .SE(n8149), .CLK(n8336), .Q(
        g4590) );
  SDFFX1 DFF_54_Q_reg ( .D(g4590), .SI(g4590), .SE(n8150), .CLK(n8337), .Q(
        g801), .QN(n4327) );
  SDFFX1 DFF_55_Q_reg ( .D(g20310), .SI(g801), .SE(n8150), .CLK(n8337), .Q(
        g6225) );
  SDFFX1 DFF_56_Q_reg ( .D(g6225), .SI(g6225), .SE(n8150), .CLK(n8337), .Q(
        g797), .QN(n4391) );
  SDFFX1 DFF_57_Q_reg ( .D(g20343), .SI(g797), .SE(n8150), .CLK(n8337), .Q(
        g6442) );
  SDFFX1 DFF_58_Q_reg ( .D(g6442), .SI(g6442), .SE(n8150), .CLK(n8337), .Q(
        g793), .QN(n4321) );
  SDFFX1 DFF_59_Q_reg ( .D(g20376), .SI(g793), .SE(n8150), .CLK(n8337), .Q(
        g6895) );
  SDFFX1 DFF_60_Q_reg ( .D(g6895), .SI(g6895), .SE(n8150), .CLK(n8337), .Q(
        g789), .QN(n4375) );
  SDFFX1 DFF_61_Q_reg ( .D(g20417), .SI(g789), .SE(n8150), .CLK(n8337), .Q(
        g7334) );
  SDFFX1 DFF_62_Q_reg ( .D(g7334), .SI(g7334), .SE(n8150), .CLK(n8337), .Q(
        g785), .QN(n4379) );
  SDFFX1 DFF_63_Q_reg ( .D(g21878), .SI(g785), .SE(n8151), .CLK(n8338), .Q(
        test_so4) );
  SDFFX1 DFF_64_Q_reg ( .D(test_so4), .SI(test_si5), .SE(n8151), .CLK(n8338), 
        .Q(g2873) );
  SDFFX1 DFF_65_Q_reg ( .D(g19153), .SI(g2873), .SE(n8151), .CLK(n8338), .Q(
        g8249) );
  SDFFX1 DFF_66_Q_reg ( .D(g8249), .SI(g8249), .SE(n8151), .CLK(n8338), .Q(
        g125), .QN(n4290) );
  SDFFX1 DFF_67_Q_reg ( .D(g19162), .SI(g125), .SE(n8151), .CLK(n8338), .Q(
        g4088) );
  SDFFX1 DFF_68_Q_reg ( .D(g4088), .SI(g4088), .SE(n8151), .CLK(n8338), .Q(
        g121), .QN(n4569) );
  SDFFX1 DFF_69_Q_reg ( .D(g19172), .SI(g121), .SE(n8151), .CLK(n8338), .Q(
        g4321) );
  SDFFX1 DFF_70_Q_reg ( .D(g4321), .SI(g4321), .SE(n8152), .CLK(n8339), .Q(
        g117), .QN(n4561) );
  SDFFX1 DFF_71_Q_reg ( .D(g19144), .SI(g117), .SE(n8152), .CLK(n8339), .Q(
        g8023) );
  SDFFX1 DFF_72_Q_reg ( .D(g8023), .SI(g8023), .SE(n8152), .CLK(n8339), .Q(
        g113), .QN(n4328) );
  SDFFX1 DFF_73_Q_reg ( .D(g19149), .SI(g113), .SE(n8152), .CLK(n8339), .Q(
        g8175) );
  SDFFX1 DFF_74_Q_reg ( .D(g8175), .SI(g8175), .SE(n8152), .CLK(n8339), .Q(
        g109), .QN(n4392) );
  SDFFX1 DFF_75_Q_reg ( .D(g19157), .SI(g109), .SE(n8152), .CLK(n8339), .Q(
        g3993) );
  SDFFX1 DFF_76_Q_reg ( .D(g3993), .SI(g3993), .SE(n8152), .CLK(n8339), .Q(
        g105), .QN(n4322) );
  SDFFX1 DFF_77_Q_reg ( .D(g19167), .SI(g105), .SE(n8152), .CLK(n8339), .Q(
        g4200) );
  SDFFX1 DFF_78_Q_reg ( .D(g4200), .SI(g4200), .SE(n8152), .CLK(n8339), .Q(
        g101), .QN(n4376) );
  SDFFX1 DFF_79_Q_reg ( .D(g19178), .SI(g101), .SE(n8152), .CLK(n8339), .Q(
        test_so5) );
  SDFFX1 DFF_80_Q_reg ( .D(test_so5), .SI(test_si6), .SE(n8152), .CLK(n8339), 
        .Q(g97), .QN(n4380) );
  SDFFX1 DFF_81_Q_reg ( .D(g20874), .SI(g97), .SE(n8152), .CLK(n8339), .Q(
        g8096) );
  SDFFX1 DFF_82_Q_reg ( .D(g8096), .SI(g8096), .SE(n8153), .CLK(n8340), .Q(
        g2857) );
  SDFFX1 DFF_83_Q_reg ( .D(g18885), .SI(g2857), .SE(n8153), .CLK(n8340), .Q(
        g2200), .QN(n4287) );
  SDFFX1 DFF_84_Q_reg ( .D(g18975), .SI(g2200), .SE(n8153), .CLK(n8340), .Q(
        g2195), .QN(n4563) );
  SDFFX1 DFF_85_Q_reg ( .D(g18968), .SI(g2195), .SE(n8153), .CLK(n8340), .Q(
        g2190), .QN(n4555) );
  SDFFX1 DFF_86_Q_reg ( .D(g18942), .SI(g2190), .SE(n8153), .CLK(n8340), .Q(
        g2185), .QN(n4325) );
  SDFFX1 DFF_87_Q_reg ( .D(g18906), .SI(g2185), .SE(n8153), .CLK(n8340), .Q(
        g2180), .QN(n4389) );
  SDFFX1 DFF_88_Q_reg ( .D(g18867), .SI(g2180), .SE(n8153), .CLK(n8340), .Q(
        g2175), .QN(n4319) );
  SDFFX1 DFF_89_Q_reg ( .D(g18836), .SI(g2175), .SE(n8153), .CLK(n8340), .Q(
        g2170), .QN(n4373) );
  SDFFX1 DFF_90_Q_reg ( .D(g18957), .SI(g2170), .SE(n8153), .CLK(n8340), .Q(
        g2165), .QN(n4377) );
  SDFFX1 DFF_91_Q_reg ( .D(g21882), .SI(g2165), .SE(n8170), .CLK(n8357), .Q(
        g2878) );
  SDFFX1 DFF_92_Q_reg ( .D(n4598), .SI(g2878), .SE(n8268), .CLK(n8455), .Q(
        g8106), .QN(n4382) );
  SDFFX1 DFF_93_Q_reg ( .D(g8106), .SI(g8106), .SE(n8268), .CLK(n8455), .Q(
        g8030), .QN(n4383) );
  SDFFX1 DFF_94_Q_reg ( .D(g8030), .SI(g8030), .SE(n8268), .CLK(n8455), .Q(
        g3109), .QN(n4494) );
  SDFFX1 DFF_95_Q_reg ( .D(g18669), .SI(g3109), .SE(n8269), .CLK(n8456), .Q(
        test_so6) );
  SDFFX1 DFF_96_Q_reg ( .D(g18719), .SI(test_si7), .SE(n8269), .CLK(n8456), 
        .Q(g3211) );
  SDFFX1 DFF_97_Q_reg ( .D(g18782), .SI(g3211), .SE(n8269), .CLK(n8456), .Q(
        g3084), .QN(n4445) );
  SDFFX1 DFF_98_Q_reg ( .D(g17222), .SI(g3084), .SE(n8271), .CLK(n8458), .Q(
        g3085) );
  SDFFX1 DFF_99_Q_reg ( .D(g17225), .SI(g3085), .SE(n8271), .CLK(n8458), .Q(
        g3086) );
  SDFFX1 DFF_100_Q_reg ( .D(g17234), .SI(g3086), .SE(n8271), .CLK(n8458), .Q(
        g3087), .QN(n4344) );
  SDFFX1 DFF_101_Q_reg ( .D(g17224), .SI(g3087), .SE(n8271), .CLK(n8458), .Q(
        g3091), .QN(n4448) );
  SDFFX1 DFF_102_Q_reg ( .D(g17228), .SI(g3091), .SE(n8271), .CLK(n8458), .Q(
        g3092), .QN(n4451) );
  SDFFX1 DFF_103_Q_reg ( .D(g17246), .SI(g3092), .SE(n8271), .CLK(n8458), .Q(
        g3093) );
  SDFFX1 DFF_104_Q_reg ( .D(g17226), .SI(g3093), .SE(n8271), .CLK(n8458), .Q(
        g3094) );
  SDFFX1 DFF_105_Q_reg ( .D(g17235), .SI(g3094), .SE(n8271), .CLK(n8458), .Q(
        g3095) );
  SDFFX1 DFF_106_Q_reg ( .D(g17269), .SI(g3095), .SE(n8146), .CLK(n8333), .Q(
        g3096) );
  SDFFX1 DFF_107_Q_reg ( .D(g25450), .SI(g3096), .SE(n8269), .CLK(n8456), .Q(
        g3097) );
  SDFFX1 DFF_108_Q_reg ( .D(g25451), .SI(g3097), .SE(n8269), .CLK(n8456), .Q(
        g3098) );
  SDFFX1 DFF_109_Q_reg ( .D(g25452), .SI(g3098), .SE(n8269), .CLK(n8456), .Q(
        g3099), .QN(n4443) );
  SDFFX1 DFF_110_Q_reg ( .D(g28420), .SI(g3099), .SE(n8269), .CLK(n8456), .Q(
        g3100), .QN(n4342) );
  SDFFX1 DFF_111_Q_reg ( .D(g28421), .SI(g3100), .SE(n8270), .CLK(n8457), .Q(
        test_so7) );
  SDFFX1 DFF_112_Q_reg ( .D(g28425), .SI(test_si8), .SE(n8269), .CLK(n8456), 
        .Q(g3102), .QN(n4343) );
  SDFFX1 DFF_113_Q_reg ( .D(g29936), .SI(g3102), .SE(n8270), .CLK(n8457), .Q(
        g3103), .QN(n4447) );
  SDFFX1 DFF_114_Q_reg ( .D(g29939), .SI(g3103), .SE(n8270), .CLK(n8457), .Q(
        g3104), .QN(n4452) );
  SDFFX1 DFF_115_Q_reg ( .D(g29941), .SI(g3104), .SE(n8270), .CLK(n8457), .Q(
        g3105) );
  SDFFX1 DFF_116_Q_reg ( .D(g30796), .SI(g3105), .SE(n8270), .CLK(n8457), .Q(
        g3106), .QN(n4438) );
  SDFFX1 DFF_117_Q_reg ( .D(g30798), .SI(g3106), .SE(n8270), .CLK(n8457), .Q(
        g3107) );
  SDFFX1 DFF_118_Q_reg ( .D(g30801), .SI(g3107), .SE(n8270), .CLK(n8457), .Q(
        g3108), .QN(n4334) );
  SDFFX1 DFF_119_Q_reg ( .D(g17229), .SI(g3108), .SE(n8270), .CLK(n8457), .Q(
        g3155) );
  SDFFX1 DFF_120_Q_reg ( .D(g17247), .SI(g3155), .SE(n8270), .CLK(n8457), .Q(
        g3158) );
  SDFFX1 DFF_121_Q_reg ( .D(g17302), .SI(g3158), .SE(n8270), .CLK(n8457), .Q(
        g3161), .QN(n4444) );
  SDFFX1 DFF_122_Q_reg ( .D(g17236), .SI(g3161), .SE(n8270), .CLK(n8457), .Q(
        g3164) );
  SDFFX1 DFF_123_Q_reg ( .D(g17270), .SI(g3164), .SE(n8270), .CLK(n8457), .Q(
        g3167) );
  SDFFX1 DFF_124_Q_reg ( .D(g17340), .SI(g3167), .SE(n8271), .CLK(n8458), .Q(
        g3170), .QN(n4441) );
  SDFFX1 DFF_125_Q_reg ( .D(g17248), .SI(g3170), .SE(n8271), .CLK(n8458), .Q(
        g3173), .QN(n4338) );
  SDFFX1 DFF_126_Q_reg ( .D(g17303), .SI(g3173), .SE(n8271), .CLK(n8458), .Q(
        g3176), .QN(n4450) );
  SDFFX1 DFF_127_Q_reg ( .D(g17383), .SI(g3176), .SE(n8271), .CLK(n8458), .Q(
        test_so8) );
  SDFFX1 DFF_128_Q_reg ( .D(g17271), .SI(test_si9), .SE(n8269), .CLK(n8456), 
        .Q(g3182) );
  SDFFX1 DFF_129_Q_reg ( .D(g17341), .SI(g3182), .SE(n8269), .CLK(n8456), .Q(
        g3185) );
  SDFFX1 DFF_130_Q_reg ( .D(g17429), .SI(g3185), .SE(n8269), .CLK(n8456), .Q(
        g3088) );
  SDFFX1 DFF_131_Q_reg ( .D(g24734), .SI(g3088), .SE(n8269), .CLK(n8456), .Q(
        n8090), .QN(DFF_131_n1) );
  SDFFX1 DFF_132_Q_reg ( .D(g25442), .SI(n8090), .SE(n8147), .CLK(n8334), .Q(
        n8089), .QN(DFF_132_n1) );
  SDFFX1 DFF_133_Q_reg ( .D(g25435), .SI(n8089), .SE(n8272), .CLK(n8459), .Q(
        g3197) );
  SDFFX1 DFF_134_Q_reg ( .D(g25420), .SI(g3197), .SE(n8272), .CLK(n8459), .Q(
        n8088), .QN(DFF_134_n1) );
  SDFFX1 DFF_135_Q_reg ( .D(g26149), .SI(n8088), .SE(n8146), .CLK(n8333), .Q(
        g3201), .QN(n4406) );
  SDFFX1 DFF_136_Q_reg ( .D(g26135), .SI(g3201), .SE(n8146), .CLK(n8333), .Q(
        g3204), .QN(n8036) );
  SDFFX1 DFF_137_Q_reg ( .D(g26104), .SI(g3204), .SE(n8146), .CLK(n8333), .Q(
        g3207), .QN(n4329) );
  SDFFX1 DFF_138_Q_reg ( .D(g27380), .SI(g3207), .SE(n8147), .CLK(n8334), .Q(
        g3188), .QN(n4405) );
  SDFFX1 DFF_139_Q_reg ( .D(n102), .SI(g3188), .SE(n8147), .CLK(n8334), .Q(
        g3133), .QN(n7442) );
  SDFFX1 DFF_140_Q_reg ( .D(g26104), .SI(g3133), .SE(n8147), .CLK(n8334), .Q(
        n8087), .QN(DFF_140_n1) );
  SDFFX1 DFF_141_Q_reg ( .D(n263), .SI(n8087), .SE(n8147), .CLK(n8334), .Q(
        g3128) );
  SDFFX1 DFF_142_Q_reg ( .D(g26149), .SI(g3128), .SE(n8147), .CLK(n8334), .Q(
        n8086) );
  SDFFX1 DFF_143_Q_reg ( .D(g25420), .SI(n8086), .SE(n8148), .CLK(n8335), .Q(
        test_so9) );
  SDFFX1 DFF_144_Q_reg ( .D(n289), .SI(test_si10), .SE(n8147), .CLK(n8334), 
        .Q(n8084), .QN(DFF_144_n1) );
  SDFFX1 DFF_145_Q_reg ( .D(g25442), .SI(n8084), .SE(n8147), .CLK(n8334), .Q(
        g3124) );
  SDFFX1 DFF_146_Q_reg ( .D(n298), .SI(g3124), .SE(n8147), .CLK(n8334), .Q(
        n8083), .QN(DFF_146_n1) );
  SDFFX1 DFF_147_Q_reg ( .D(g26104), .SI(n8083), .SE(n8147), .CLK(n8334), .Q(
        n8082), .QN(n14382) );
  SDFFX1 DFF_148_Q_reg ( .D(g26135), .SI(n8082), .SE(n8148), .CLK(n8335), .Q(
        n8081), .QN(n14384) );
  SDFFX1 DFF_149_Q_reg ( .D(g26149), .SI(n8081), .SE(n8148), .CLK(n8335), .Q(
        n8080), .QN(DFF_149_n1) );
  SDFFX1 DFF_150_Q_reg ( .D(g25420), .SI(n8080), .SE(n8148), .CLK(n8335), .Q(
        g3112) );
  SDFFX1 DFF_151_Q_reg ( .D(g25435), .SI(g3112), .SE(n8148), .CLK(n8335), .Q(
        g3110) );
  SDFFX1 DFF_152_Q_reg ( .D(g25442), .SI(g3110), .SE(n8148), .CLK(n8335), .Q(
        g3111) );
  SDFFX1 DFF_153_Q_reg ( .D(g27380), .SI(g3111), .SE(n8148), .CLK(n8335), .Q(
        n8079), .QN(n14385) );
  SDFFX1 DFF_154_Q_reg ( .D(g26104), .SI(n8079), .SE(n8148), .CLK(n8335), .Q(
        n8078), .QN(n14386) );
  SDFFX1 DFF_155_Q_reg ( .D(g26135), .SI(n8078), .SE(n8148), .CLK(n8335), .Q(
        n8077), .QN(DFF_155_n1) );
  SDFFX1 DFF_156_Q_reg ( .D(g26149), .SI(n8077), .SE(n8148), .CLK(n8335), .Q(
        n8076), .QN(DFF_156_n1) );
  SDFFX1 DFF_157_Q_reg ( .D(g27380), .SI(n8076), .SE(n8148), .CLK(n8335), .Q(
        g3151), .QN(n4424) );
  SDFFX1 DFF_158_Q_reg ( .D(g26104), .SI(g3151), .SE(n8148), .CLK(n8335), .Q(
        g3142), .QN(n4301) );
  SDFFX1 DFF_159_Q_reg ( .D(g26135), .SI(g3142), .SE(n8149), .CLK(n8336), .Q(
        test_so10), .QN(n8112) );
  SDFFX1 DFF_160_Q_reg ( .D(n102), .SI(test_si11), .SE(n8146), .CLK(n8333), 
        .Q(g185) );
  SDFFX1 DFF_161_Q_reg ( .D(g2950), .SI(g185), .SE(n8146), .CLK(n8333), .Q(
        g6231), .QN(n4318) );
  SDFFX1 DFF_162_Q_reg ( .D(g6231), .SI(g6231), .SE(n8147), .CLK(n8334), .Q(
        g6313), .QN(n4512) );
  SDFFX1 DFF_163_Q_reg ( .D(g6313), .SI(g6313), .SE(n8147), .CLK(n8334), .Q(
        g165), .QN(n4369) );
  SDFFX1 DFF_164_Q_reg ( .D(g22100), .SI(g165), .SE(n8160), .CLK(n8347), .Q(
        g130), .QN(n7973) );
  SDFFX1 DFF_165_Q_reg ( .D(g22122), .SI(g130), .SE(n8160), .CLK(n8347), .Q(
        g131), .QN(n7972) );
  SDFFX1 DFF_166_Q_reg ( .D(g22141), .SI(g131), .SE(n8160), .CLK(n8347), .Q(
        g129), .QN(n7566) );
  SDFFX1 DFF_167_Q_reg ( .D(g22123), .SI(g129), .SE(n8160), .CLK(n8347), .Q(
        g133), .QN(n7970) );
  SDFFX1 DFF_168_Q_reg ( .D(g22142), .SI(g133), .SE(n8160), .CLK(n8347), .Q(
        g134), .QN(n7969) );
  SDFFX1 DFF_169_Q_reg ( .D(g22161), .SI(g134), .SE(n8160), .CLK(n8347), .Q(
        g132), .QN(n7565) );
  SDFFX1 DFF_170_Q_reg ( .D(g22025), .SI(g132), .SE(n8160), .CLK(n8347), .Q(
        g142), .QN(n7961) );
  SDFFX1 DFF_171_Q_reg ( .D(g22027), .SI(g142), .SE(n8161), .CLK(n8348), .Q(
        g143), .QN(n7959) );
  SDFFX1 DFF_172_Q_reg ( .D(g22030), .SI(g143), .SE(n8161), .CLK(n8348), .Q(
        g141), .QN(n7564) );
  SDFFX1 DFF_173_Q_reg ( .D(g22028), .SI(g141), .SE(n8161), .CLK(n8348), .Q(
        g145), .QN(n7958) );
  SDFFX1 DFF_174_Q_reg ( .D(g22031), .SI(g145), .SE(n8161), .CLK(n8348), .Q(
        g146), .QN(n7957) );
  SDFFX1 DFF_175_Q_reg ( .D(g22037), .SI(g146), .SE(n8161), .CLK(n8348), .Q(
        test_so11), .QN(n8127) );
  SDFFX1 DFF_176_Q_reg ( .D(g22032), .SI(test_si12), .SE(n8159), .CLK(n8346), 
        .Q(g148), .QN(n7956) );
  SDFFX1 DFF_177_Q_reg ( .D(g22038), .SI(g148), .SE(n8159), .CLK(n8346), .Q(
        g149), .QN(n7955) );
  SDFFX1 DFF_178_Q_reg ( .D(g22047), .SI(g149), .SE(n8159), .CLK(n8346), .Q(
        g147), .QN(n7563) );
  SDFFX1 DFF_179_Q_reg ( .D(g22039), .SI(g147), .SE(n8159), .CLK(n8346), .Q(
        g151), .QN(n7954) );
  SDFFX1 DFF_180_Q_reg ( .D(g22048), .SI(g151), .SE(n8159), .CLK(n8346), .Q(
        g152), .QN(n7953) );
  SDFFX1 DFF_181_Q_reg ( .D(g22063), .SI(g152), .SE(n8159), .CLK(n8346), .Q(
        g150), .QN(n7562) );
  SDFFX1 DFF_182_Q_reg ( .D(g22049), .SI(g150), .SE(n8159), .CLK(n8346), .Q(
        g154), .QN(n7952) );
  SDFFX1 DFF_183_Q_reg ( .D(g22064), .SI(g154), .SE(n8159), .CLK(n8346), .Q(
        g155), .QN(n7951) );
  SDFFX1 DFF_184_Q_reg ( .D(g22079), .SI(g155), .SE(n8160), .CLK(n8347), .Q(
        g153), .QN(n7561) );
  SDFFX1 DFF_185_Q_reg ( .D(g22065), .SI(g153), .SE(n8156), .CLK(n8343), .Q(
        g157), .QN(n7950) );
  SDFFX1 DFF_186_Q_reg ( .D(g22080), .SI(g157), .SE(n8158), .CLK(n8345), .Q(
        g158), .QN(n7949) );
  SDFFX1 DFF_187_Q_reg ( .D(g22101), .SI(g158), .SE(n8158), .CLK(n8345), .Q(
        g156), .QN(n7560) );
  SDFFX1 DFF_188_Q_reg ( .D(g22081), .SI(g156), .SE(n8160), .CLK(n8347), .Q(
        g160), .QN(n7522) );
  SDFFX1 DFF_189_Q_reg ( .D(g22102), .SI(g160), .SE(n8160), .CLK(n8347), .Q(
        g161), .QN(n7521) );
  SDFFX1 DFF_190_Q_reg ( .D(g22124), .SI(g161), .SE(n8160), .CLK(n8347), .Q(
        g159), .QN(n7520) );
  SDFFX1 DFF_191_Q_reg ( .D(g22103), .SI(g159), .SE(n8160), .CLK(n8347), .Q(
        test_so12), .QN(n8126) );
  SDFFX1 DFF_192_Q_reg ( .D(g22125), .SI(test_si13), .SE(n8158), .CLK(n8345), 
        .Q(g164), .QN(n7559) );
  SDFFX1 DFF_193_Q_reg ( .D(g22143), .SI(g164), .SE(n8158), .CLK(n8345), .Q(
        g162), .QN(n7558) );
  SDFFX1 DFF_194_Q_reg ( .D(g25204), .SI(g162), .SE(n8158), .CLK(n8345), .Q(
        g169), .QN(n7624) );
  SDFFX1 DFF_195_Q_reg ( .D(g25206), .SI(g169), .SE(n8158), .CLK(n8345), .Q(
        g170), .QN(n7623) );
  SDFFX1 DFF_196_Q_reg ( .D(g25211), .SI(g170), .SE(n8158), .CLK(n8345), .Q(
        g168), .QN(n7622) );
  SDFFX1 DFF_197_Q_reg ( .D(g25207), .SI(g168), .SE(n8158), .CLK(n8345), .Q(
        g172), .QN(n7621) );
  SDFFX1 DFF_198_Q_reg ( .D(g25212), .SI(g172), .SE(n8158), .CLK(n8345), .Q(
        g173), .QN(n7620) );
  SDFFX1 DFF_199_Q_reg ( .D(g25218), .SI(g173), .SE(n8158), .CLK(n8345), .Q(
        g171), .QN(n7619) );
  SDFFX1 DFF_200_Q_reg ( .D(g25213), .SI(g171), .SE(n8158), .CLK(n8345), .Q(
        g175), .QN(n7618) );
  SDFFX1 DFF_201_Q_reg ( .D(g25219), .SI(g175), .SE(n8158), .CLK(n8345), .Q(
        g176), .QN(n7617) );
  SDFFX1 DFF_202_Q_reg ( .D(g25228), .SI(g176), .SE(n8159), .CLK(n8346), .Q(
        g174), .QN(n7616) );
  SDFFX1 DFF_203_Q_reg ( .D(g25220), .SI(g174), .SE(n8159), .CLK(n8346), .Q(
        g178), .QN(n7615) );
  SDFFX1 DFF_204_Q_reg ( .D(g25229), .SI(g178), .SE(n8159), .CLK(n8346), .Q(
        g179), .QN(n7614) );
  SDFFX1 DFF_205_Q_reg ( .D(g25239), .SI(g179), .SE(n8159), .CLK(n8346), .Q(
        g177), .QN(n7613) );
  SDFFX1 DFF_206_Q_reg ( .D(g30261), .SI(g177), .SE(n8163), .CLK(n8350), .Q(
        g186) );
  SDFFX1 DFF_207_Q_reg ( .D(g30267), .SI(g186), .SE(n8163), .CLK(n8350), .Q(
        test_so13) );
  SDFFX1 DFF_208_Q_reg ( .D(g30275), .SI(test_si14), .SE(n8163), .CLK(n8350), 
        .Q(g192) );
  SDFFX1 DFF_209_Q_reg ( .D(g30637), .SI(g192), .SE(n8163), .CLK(n8350), .Q(
        g231) );
  SDFFX1 DFF_210_Q_reg ( .D(g30640), .SI(g231), .SE(n8163), .CLK(n8350), .Q(
        g234) );
  SDFFX1 DFF_211_Q_reg ( .D(g30645), .SI(g234), .SE(n8163), .CLK(n8350), .Q(
        g237) );
  SDFFX1 DFF_212_Q_reg ( .D(g30668), .SI(g237), .SE(n8163), .CLK(n8350), .Q(
        g195) );
  SDFFX1 DFF_213_Q_reg ( .D(g30674), .SI(g195), .SE(n8164), .CLK(n8351), .Q(
        g198) );
  SDFFX1 DFF_214_Q_reg ( .D(g30680), .SI(g198), .SE(n8156), .CLK(n8343), .Q(
        g201) );
  SDFFX1 DFF_215_Q_reg ( .D(g30641), .SI(g201), .SE(n8161), .CLK(n8348), .Q(
        g240) );
  SDFFX1 DFF_216_Q_reg ( .D(g30646), .SI(g240), .SE(n8161), .CLK(n8348), .Q(
        g243) );
  SDFFX1 DFF_217_Q_reg ( .D(g30653), .SI(g243), .SE(n8161), .CLK(n8348), .Q(
        g246) );
  SDFFX1 DFF_218_Q_reg ( .D(g30276), .SI(g246), .SE(n8161), .CLK(n8348), .Q(
        g204) );
  SDFFX1 DFF_219_Q_reg ( .D(g30284), .SI(g204), .SE(n8161), .CLK(n8348), .Q(
        g207) );
  SDFFX1 DFF_220_Q_reg ( .D(g30292), .SI(g207), .SE(n8161), .CLK(n8348), .Q(
        g210) );
  SDFFX1 DFF_221_Q_reg ( .D(g30254), .SI(g210), .SE(n8161), .CLK(n8348), .Q(
        g249) );
  SDFFX1 DFF_222_Q_reg ( .D(g30257), .SI(g249), .SE(n8162), .CLK(n8349), .Q(
        g252) );
  SDFFX1 DFF_223_Q_reg ( .D(g30262), .SI(g252), .SE(n8162), .CLK(n8349), .Q(
        test_so14) );
  SDFFX1 DFF_224_Q_reg ( .D(g30245), .SI(test_si15), .SE(n8162), .CLK(n8349), 
        .Q(g213) );
  SDFFX1 DFF_225_Q_reg ( .D(g30246), .SI(g213), .SE(n8162), .CLK(n8349), .Q(
        g216) );
  SDFFX1 DFF_226_Q_reg ( .D(g30248), .SI(g216), .SE(n8162), .CLK(n8349), .Q(
        g219) );
  SDFFX1 DFF_227_Q_reg ( .D(g30258), .SI(g219), .SE(n8162), .CLK(n8349), .Q(
        g258) );
  SDFFX1 DFF_228_Q_reg ( .D(g30263), .SI(g258), .SE(n8162), .CLK(n8349), .Q(
        g261) );
  SDFFX1 DFF_229_Q_reg ( .D(g30268), .SI(g261), .SE(n8162), .CLK(n8349), .Q(
        g264) );
  SDFFX1 DFF_230_Q_reg ( .D(g30635), .SI(g264), .SE(n8162), .CLK(n8349), .Q(
        g222) );
  SDFFX1 DFF_231_Q_reg ( .D(g30636), .SI(g222), .SE(n8162), .CLK(n8349), .Q(
        g225) );
  SDFFX1 DFF_232_Q_reg ( .D(g30639), .SI(g225), .SE(n8162), .CLK(n8349), .Q(
        g228) );
  SDFFX1 DFF_233_Q_reg ( .D(g30661), .SI(g228), .SE(n8162), .CLK(n8349), .Q(
        g267) );
  SDFFX1 DFF_234_Q_reg ( .D(g30669), .SI(g267), .SE(n8163), .CLK(n8350), .Q(
        g270) );
  SDFFX1 DFF_235_Q_reg ( .D(g30675), .SI(g270), .SE(n8156), .CLK(n8343), .Q(
        g273) );
  SDFFX1 DFF_236_Q_reg ( .D(g25027), .SI(g273), .SE(n8156), .CLK(n8343), .Q(
        g92), .QN(n7714) );
  SDFFX1 DFF_237_Q_reg ( .D(g25932), .SI(g92), .SE(n8156), .CLK(n8343), .Q(g88) );
  SDFFX1 DFF_238_Q_reg ( .D(g26529), .SI(g88), .SE(n8156), .CLK(n8343), .Q(g83), .QN(n7713) );
  SDFFX1 DFF_239_Q_reg ( .D(g27120), .SI(g83), .SE(n8156), .CLK(n8343), .Q(
        test_so15) );
  SDFFX1 DFF_240_Q_reg ( .D(g27594), .SI(test_si16), .SE(n8156), .CLK(n8343), 
        .Q(g74), .QN(n7712) );
  SDFFX1 DFF_241_Q_reg ( .D(g28145), .SI(g74), .SE(n8157), .CLK(n8344), .Q(g70), .QN(n8093) );
  SDFFX1 DFF_242_Q_reg ( .D(g28634), .SI(g70), .SE(n8157), .CLK(n8344), .Q(g65), .QN(n7711) );
  SDFFX1 DFF_243_Q_reg ( .D(g29109), .SI(g65), .SE(n8157), .CLK(n8344), .Q(g61), .QN(n8070) );
  SDFFX1 DFF_244_Q_reg ( .D(g29353), .SI(g61), .SE(n8157), .CLK(n8344), .Q(g56), .QN(n7337) );
  SDFFX1 DFF_245_Q_reg ( .D(g29579), .SI(g56), .SE(n8157), .CLK(n8344), .Q(g52), .QN(n7176) );
  SDFFX1 DFF_246_Q_reg ( .D(n15), .SI(g52), .SE(n8157), .CLK(n8344), .Q(g180)
         );
  SDFFX1 DFF_247_Q_reg ( .D(g180), .SI(g180), .SE(n8157), .CLK(n8344), .Q(
        g5549) );
  SDFFX1 DFF_248_Q_reg ( .D(g5549), .SI(g5549), .SE(n8157), .CLK(n8344), .Q(
        g181), .QN(n7721) );
  SDFFX1 DFF_251_Q_reg ( .D(g6447), .SI(g6447), .SE(n8157), .CLK(n8344), .Q(
        n4640), .QN(n4506) );
  SDFFX1 DFF_252_Q_reg ( .D(g5549), .SI(n4640), .SE(n8157), .CLK(n8344), .Q(
        g309), .QN(n4388) );
  SDFFX1 DFF_253_Q_reg ( .D(g27253), .SI(g309), .SE(n8166), .CLK(n8353), .Q(
        g354), .QN(n7665) );
  SDFFX1 DFF_254_Q_reg ( .D(g27255), .SI(g354), .SE(n8166), .CLK(n8353), .Q(
        g343), .QN(n7664) );
  SDFFX1 DFF_255_Q_reg ( .D(g27258), .SI(g343), .SE(n8166), .CLK(n8353), .Q(
        test_so16), .QN(n8115) );
  SDFFX1 DFF_256_Q_reg ( .D(g27256), .SI(test_si17), .SE(n8167), .CLK(n8354), 
        .Q(g369), .QN(n7643) );
  SDFFX1 DFF_257_Q_reg ( .D(g27259), .SI(g369), .SE(n8167), .CLK(n8354), .Q(
        g358), .QN(n7642) );
  SDFFX1 DFF_258_Q_reg ( .D(g27265), .SI(g358), .SE(n8167), .CLK(n8354), .Q(
        g361), .QN(n7641) );
  SDFFX1 DFF_259_Q_reg ( .D(g27260), .SI(g361), .SE(n8167), .CLK(n8354), .Q(
        g384), .QN(n7391) );
  SDFFX1 DFF_260_Q_reg ( .D(g27266), .SI(g384), .SE(n8167), .CLK(n8354), .Q(
        g373), .QN(n7393) );
  SDFFX1 DFF_261_Q_reg ( .D(g27277), .SI(g373), .SE(n8166), .CLK(n8353), .Q(
        g376), .QN(n7392) );
  SDFFX1 DFF_262_Q_reg ( .D(g27267), .SI(g376), .SE(n8167), .CLK(n8354), .Q(
        g398), .QN(n7654) );
  SDFFX1 DFF_263_Q_reg ( .D(g27278), .SI(g398), .SE(n8167), .CLK(n8354), .Q(
        g388), .QN(n7653) );
  SDFFX1 DFF_264_Q_reg ( .D(g27293), .SI(g388), .SE(n8164), .CLK(n8351), .Q(
        g391), .QN(n7652) );
  SDFFX1 DFF_265_Q_reg ( .D(g28732), .SI(g391), .SE(n8164), .CLK(n8351), .Q(
        g408) );
  SDFFX1 DFF_266_Q_reg ( .D(g28735), .SI(g408), .SE(n8166), .CLK(n8353), .Q(
        g411) );
  SDFFX1 DFF_267_Q_reg ( .D(g28744), .SI(g411), .SE(n8166), .CLK(n8353), .Q(
        g414) );
  SDFFX1 DFF_268_Q_reg ( .D(g29194), .SI(g414), .SE(n8166), .CLK(n8353), .Q(
        g417) );
  SDFFX1 DFF_269_Q_reg ( .D(g29197), .SI(g417), .SE(n8166), .CLK(n8353), .Q(
        g420) );
  SDFFX1 DFF_270_Q_reg ( .D(g29201), .SI(g420), .SE(n8165), .CLK(n8352), .Q(
        g423) );
  SDFFX1 DFF_271_Q_reg ( .D(g28736), .SI(g423), .SE(n8165), .CLK(n8352), .Q(
        test_so17), .QN(n8118) );
  SDFFX1 DFF_272_Q_reg ( .D(g28745), .SI(test_si18), .SE(n8165), .CLK(n8352), 
        .Q(g428), .QN(n7697) );
  SDFFX1 DFF_273_Q_reg ( .D(g28754), .SI(g428), .SE(n8165), .CLK(n8352), .Q(
        g426), .QN(n7696) );
  SDFFX1 DFF_274_Q_reg ( .D(g26803), .SI(g426), .SE(n8165), .CLK(n8352), .Q(
        g429) );
  SDFFX1 DFF_275_Q_reg ( .D(g26804), .SI(g429), .SE(n8165), .CLK(n8352), .Q(
        g432) );
  SDFFX1 DFF_276_Q_reg ( .D(g26807), .SI(g432), .SE(n8165), .CLK(n8352), .Q(
        g435) );
  SDFFX1 DFF_277_Q_reg ( .D(g26805), .SI(g435), .SE(n8165), .CLK(n8352), .Q(
        g438) );
  SDFFX1 DFF_278_Q_reg ( .D(g26808), .SI(g438), .SE(n8165), .CLK(n8352), .Q(
        g441) );
  SDFFX1 DFF_279_Q_reg ( .D(g26812), .SI(g441), .SE(n8166), .CLK(n8353), .Q(
        g444) );
  SDFFX1 DFF_280_Q_reg ( .D(g27759), .SI(g444), .SE(n8166), .CLK(n8353), .Q(
        g448), .QN(n7695) );
  SDFFX1 DFF_281_Q_reg ( .D(g27760), .SI(g448), .SE(n8166), .CLK(n8353), .Q(
        g449), .QN(n7694) );
  SDFFX1 DFF_282_Q_reg ( .D(g27762), .SI(g449), .SE(n8165), .CLK(n8352), .Q(
        g447), .QN(n7693) );
  SDFFX1 DFF_283_Q_reg ( .D(g29606), .SI(g447), .SE(n8165), .CLK(n8352), .Q(
        g312), .QN(n7301) );
  SDFFX1 DFF_284_Q_reg ( .D(g29608), .SI(g312), .SE(n8165), .CLK(n8352), .Q(
        g313), .QN(n7300) );
  SDFFX1 DFF_285_Q_reg ( .D(g29611), .SI(g313), .SE(n8164), .CLK(n8351), .Q(
        g314), .QN(n7299) );
  SDFFX1 DFF_286_Q_reg ( .D(g30699), .SI(g314), .SE(n8164), .CLK(n8351), .Q(
        g315), .QN(n7298) );
  SDFFX1 DFF_287_Q_reg ( .D(g30700), .SI(g315), .SE(n8164), .CLK(n8351), .Q(
        test_so18), .QN(n8140) );
  SDFFX1 DFF_288_Q_reg ( .D(g30702), .SI(test_si19), .SE(n8163), .CLK(n8350), 
        .Q(g317), .QN(n7297) );
  SDFFX1 DFF_289_Q_reg ( .D(g30455), .SI(g317), .SE(n8163), .CLK(n8350), .Q(
        g318), .QN(n7296) );
  SDFFX1 DFF_290_Q_reg ( .D(g30468), .SI(g318), .SE(n8163), .CLK(n8350), .Q(
        g319), .QN(n7295) );
  SDFFX1 DFF_291_Q_reg ( .D(g30482), .SI(g319), .SE(n8163), .CLK(n8350), .Q(
        g320), .QN(n7294) );
  SDFFX1 DFF_292_Q_reg ( .D(g29167), .SI(g320), .SE(n8164), .CLK(n8351), .Q(
        g322), .QN(n7333) );
  SDFFX1 DFF_293_Q_reg ( .D(g29169), .SI(g322), .SE(n8164), .CLK(n8351), .Q(
        g323), .QN(n7332) );
  SDFFX1 DFF_294_Q_reg ( .D(g29172), .SI(g323), .SE(n8164), .CLK(n8351), .Q(
        g321), .QN(n7331) );
  SDFFX1 DFF_295_Q_reg ( .D(g26655), .SI(g321), .SE(n8164), .CLK(n8351), .Q(
        g403), .QN(n7692) );
  SDFFX1 DFF_296_Q_reg ( .D(g26659), .SI(g403), .SE(n8164), .CLK(n8351), .Q(
        g404), .QN(n7691) );
  SDFFX1 DFF_297_Q_reg ( .D(g26664), .SI(g404), .SE(n8164), .CLK(n8351), .Q(
        g402), .QN(n7690) );
  SDFFX1 DFF_298_Q_reg ( .D(n4290), .SI(g402), .SE(n8169), .CLK(n8356), .Q(
        g450) );
  SDFFX1 DFF_299_Q_reg ( .D(g450), .SI(g450), .SE(n8170), .CLK(n8357), .Q(
        n8066), .QN(DFF_299_n1) );
  SDFFX1 DFF_300_Q_reg ( .D(n4569), .SI(n8066), .SE(n8170), .CLK(n8357), .Q(
        g452) );
  SDFFX1 DFF_301_Q_reg ( .D(g452), .SI(g452), .SE(n8170), .CLK(n8357), .Q(
        n8065), .QN(DFF_301_n1) );
  SDFFX1 DFF_302_Q_reg ( .D(n4561), .SI(n8065), .SE(n8170), .CLK(n8357), .Q(
        g454) );
  SDFFX1 DFF_303_Q_reg ( .D(g454), .SI(g454), .SE(n8170), .CLK(n8357), .Q(
        test_so19), .QN(DFF_303_n1) );
  SDFFX1 DFF_304_Q_reg ( .D(n4328), .SI(test_si20), .SE(n8155), .CLK(n8342), 
        .Q(g280) );
  SDFFX1 DFF_305_Q_reg ( .D(g280), .SI(g280), .SE(n8155), .CLK(n8342), .Q(
        n8062), .QN(DFF_305_n1) );
  SDFFX1 DFF_306_Q_reg ( .D(n4392), .SI(n8062), .SE(n8155), .CLK(n8342), .Q(
        g282) );
  SDFFX1 DFF_307_Q_reg ( .D(g282), .SI(g282), .SE(n8155), .CLK(n8342), .Q(
        n8061), .QN(DFF_307_n1) );
  SDFFX1 DFF_308_Q_reg ( .D(n4322), .SI(n8061), .SE(n8155), .CLK(n8342), .Q(
        g284) );
  SDFFX1 DFF_309_Q_reg ( .D(g284), .SI(g284), .SE(n8155), .CLK(n8342), .Q(
        n8060), .QN(DFF_309_n1) );
  SDFFX1 DFF_310_Q_reg ( .D(n4376), .SI(n8060), .SE(n8155), .CLK(n8342), .Q(
        g286) );
  SDFFX1 DFF_311_Q_reg ( .D(g286), .SI(g286), .SE(n8155), .CLK(n8342), .Q(
        n8059), .QN(DFF_311_n1) );
  SDFFX1 DFF_312_Q_reg ( .D(n4380), .SI(n8059), .SE(n8155), .CLK(n8342), .Q(
        g288) );
  SDFFX1 DFF_313_Q_reg ( .D(g288), .SI(g288), .SE(n8155), .CLK(n8342), .Q(
        n8058), .QN(DFF_313_n1) );
  SDFFX1 DFF_314_Q_reg ( .D(g2857), .SI(n8058), .SE(n8156), .CLK(n8343), .Q(
        g290) );
  SDFFX1 DFF_315_Q_reg ( .D(g290), .SI(g290), .SE(n8156), .CLK(n8343), .Q(
        n8057), .QN(n4485) );
  SDFFX1 DFF_316_Q_reg ( .D(n4282), .SI(n8057), .SE(n8166), .CLK(n8353), .Q(
        n8056), .QN(n14388) );
  SDFFX1 DFF_317_Q_reg ( .D(g21346), .SI(n8056), .SE(n8169), .CLK(n8356), .Q(
        g305), .QN(n7445) );
  SDFFX1 DFF_328_Q_reg ( .D(n4278), .SI(g305), .SE(n8167), .CLK(n8354), .Q(
        n8055), .QN(DFF_328_n1) );
  SDFFX1 DFF_329_Q_reg ( .D(g354), .SI(n8055), .SE(n8167), .CLK(n8354), .Q(
        test_so20) );
  SDFFX1 DFF_330_Q_reg ( .D(test_so20), .SI(test_si21), .SE(n8167), .CLK(n8354), .Q(g349) );
  SDFFX1 DFF_331_Q_reg ( .D(g343), .SI(g349), .SE(n8167), .CLK(n8354), .Q(g350) );
  SDFFX1 DFF_332_Q_reg ( .D(g350), .SI(g350), .SE(n8167), .CLK(n8354), .Q(g351) );
  SDFFX1 DFF_333_Q_reg ( .D(test_so16), .SI(g351), .SE(n8168), .CLK(n8355), 
        .Q(g352) );
  SDFFX1 DFF_334_Q_reg ( .D(g352), .SI(g352), .SE(n8168), .CLK(n8355), .Q(g353) );
  SDFFX1 DFF_335_Q_reg ( .D(g369), .SI(g353), .SE(n8168), .CLK(n8355), .Q(g357) );
  SDFFX1 DFF_336_Q_reg ( .D(g357), .SI(g357), .SE(n8168), .CLK(n8355), .Q(g364) );
  SDFFX1 DFF_337_Q_reg ( .D(g358), .SI(g364), .SE(n8168), .CLK(n8355), .Q(g365) );
  SDFFX1 DFF_338_Q_reg ( .D(g365), .SI(g365), .SE(n8168), .CLK(n8355), .Q(g366) );
  SDFFX1 DFF_339_Q_reg ( .D(g361), .SI(g366), .SE(n8168), .CLK(n8355), .Q(g367) );
  SDFFX1 DFF_340_Q_reg ( .D(g367), .SI(g367), .SE(n8168), .CLK(n8355), .Q(g368) );
  SDFFX1 DFF_341_Q_reg ( .D(g384), .SI(g368), .SE(n8168), .CLK(n8355), .Q(g372) );
  SDFFX1 DFF_342_Q_reg ( .D(g372), .SI(g372), .SE(n8168), .CLK(n8355), .Q(g379) );
  SDFFX1 DFF_343_Q_reg ( .D(g373), .SI(g379), .SE(n8168), .CLK(n8355), .Q(g380) );
  SDFFX1 DFF_344_Q_reg ( .D(g380), .SI(g380), .SE(n8168), .CLK(n8355), .Q(g381) );
  SDFFX1 DFF_345_Q_reg ( .D(g376), .SI(g381), .SE(n8169), .CLK(n8356), .Q(
        test_so21) );
  SDFFX1 DFF_346_Q_reg ( .D(test_so21), .SI(test_si22), .SE(n8169), .CLK(n8356), .Q(g383) );
  SDFFX1 DFF_347_Q_reg ( .D(g398), .SI(g383), .SE(n8169), .CLK(n8356), .Q(g387) );
  SDFFX1 DFF_348_Q_reg ( .D(g387), .SI(g387), .SE(n8169), .CLK(n8356), .Q(g394) );
  SDFFX1 DFF_349_Q_reg ( .D(g388), .SI(g394), .SE(n8169), .CLK(n8356), .Q(g395) );
  SDFFX1 DFF_350_Q_reg ( .D(g395), .SI(g395), .SE(n8169), .CLK(n8356), .Q(g396) );
  SDFFX1 DFF_351_Q_reg ( .D(g391), .SI(g396), .SE(n8169), .CLK(n8356), .Q(g397) );
  SDFFX1 DFF_352_Q_reg ( .D(g397), .SI(g397), .SE(n8169), .CLK(n8356), .Q(g324) );
  SDFFX1 DFF_353_Q_reg ( .D(n4598), .SI(g324), .SE(n8173), .CLK(n8360), .Q(
        g5629) );
  SDFFX1 DFF_354_Q_reg ( .D(g5629), .SI(g5629), .SE(n8173), .CLK(n8360), .Q(
        g5648) );
  SDFFX1 DFF_355_Q_reg ( .D(g5648), .SI(g5648), .SE(n8173), .CLK(n8360), .Q(
        g337) );
  SDFFX1 DFF_356_Q_reg ( .D(n4598), .SI(g337), .SE(n8173), .CLK(n8360), .Q(
        g6485), .QN(n4298) );
  SDFFX1 DFF_357_Q_reg ( .D(g6485), .SI(g6485), .SE(n8173), .CLK(n8360), .Q(
        g6642), .QN(n4372) );
  SDFFX1 DFF_358_Q_reg ( .D(g6642), .SI(g6642), .SE(n8173), .CLK(n8360), .Q(
        g550), .QN(n4313) );
  SDFFX1 DFF_359_Q_reg ( .D(n539), .SI(g550), .SE(n8173), .CLK(n8360), .Q(g554), .QN(n7993) );
  SDFFX1 DFF_360_Q_reg ( .D(g18678), .SI(g554), .SE(n8173), .CLK(n8360), .Q(
        g557), .QN(n4360) );
  SDFFX1 DFF_361_Q_reg ( .D(g18726), .SI(g557), .SE(n8173), .CLK(n8360), .Q(
        test_so22), .QN(n8108) );
  SDFFX1 DFF_362_Q_reg ( .D(n534), .SI(test_si23), .SE(n8173), .CLK(n8360), 
        .Q(g513) );
  SDFFX1 DFF_363_Q_reg ( .D(g513), .SI(g513), .SE(n8174), .CLK(n8361), .Q(g523) );
  SDFFX1 DFF_364_Q_reg ( .D(g523), .SI(g523), .SE(n8174), .CLK(n8361), .Q(g524) );
  SDFFX1 DFF_365_Q_reg ( .D(g455), .SI(g524), .SE(n8174), .CLK(n8361), .Q(g564) );
  SDFFX1 DFF_366_Q_reg ( .D(g564), .SI(g564), .SE(n8174), .CLK(n8361), .Q(g569) );
  SDFFX1 DFF_367_Q_reg ( .D(g458), .SI(g569), .SE(n8174), .CLK(n8361), .Q(g570) );
  SDFFX1 DFF_368_Q_reg ( .D(g570), .SI(g570), .SE(n8174), .CLK(n8361), .Q(g571) );
  SDFFX1 DFF_369_Q_reg ( .D(g461), .SI(g571), .SE(n8174), .CLK(n8361), .Q(g572) );
  SDFFX1 DFF_370_Q_reg ( .D(g572), .SI(g572), .SE(n8174), .CLK(n8361), .Q(g573) );
  SDFFX1 DFF_371_Q_reg ( .D(g465), .SI(g573), .SE(n8174), .CLK(n8361), .Q(g574) );
  SDFFX1 DFF_372_Q_reg ( .D(g574), .SI(g574), .SE(n8174), .CLK(n8361), .Q(g565) );
  SDFFX1 DFF_373_Q_reg ( .D(test_so24), .SI(g565), .SE(n8174), .CLK(n8361), 
        .Q(g566) );
  SDFFX1 DFF_374_Q_reg ( .D(g566), .SI(g566), .SE(n8174), .CLK(n8361), .Q(g567) );
  SDFFX1 DFF_375_Q_reg ( .D(g471), .SI(g567), .SE(n8175), .CLK(n8362), .Q(g568) );
  SDFFX1 DFF_376_Q_reg ( .D(g568), .SI(g568), .SE(n8175), .CLK(n8362), .Q(g489) );
  SDFFX1 DFF_377_Q_reg ( .D(g2950), .SI(g489), .SE(n8175), .CLK(n8362), .Q(
        test_so23), .QN(n8100) );
  SDFFX1 DFF_378_Q_reg ( .D(test_so23), .SI(test_si24), .SE(n8175), .CLK(n8362), .Q(g7956), .QN(n4461) );
  SDFFX1 DFF_379_Q_reg ( .D(g7956), .SI(g7956), .SE(n8175), .CLK(n8362), .Q(
        g485), .QN(n4466) );
  SDFFX1 DFF_380_Q_reg ( .D(g23067), .SI(g485), .SE(n8175), .CLK(n8362), .Q(
        g486) );
  SDFFX1 DFF_381_Q_reg ( .D(g23093), .SI(g486), .SE(n8175), .CLK(n8362), .Q(
        g487) );
  SDFFX1 DFF_382_Q_reg ( .D(g23117), .SI(g487), .SE(n8175), .CLK(n8362), .Q(
        g488) );
  SDFFX1 DFF_383_Q_reg ( .D(g23385), .SI(g488), .SE(n8175), .CLK(n8362), .Q(
        g455) );
  SDFFX1 DFF_384_Q_reg ( .D(g23399), .SI(g455), .SE(n8175), .CLK(n8362), .Q(
        g458) );
  SDFFX1 DFF_385_Q_reg ( .D(g24174), .SI(g458), .SE(n8175), .CLK(n8362), .Q(
        g461) );
  SDFFX1 DFF_386_Q_reg ( .D(g24178), .SI(g461), .SE(n8176), .CLK(n8363), .Q(
        g477) );
  SDFFX1 DFF_387_Q_reg ( .D(g24207), .SI(g477), .SE(n8176), .CLK(n8363), .Q(
        g478) );
  SDFFX1 DFF_388_Q_reg ( .D(g24216), .SI(g478), .SE(n8176), .CLK(n8363), .Q(
        g479) );
  SDFFX1 DFF_389_Q_reg ( .D(g23092), .SI(g479), .SE(n8176), .CLK(n8363), .Q(
        g480) );
  SDFFX1 DFF_390_Q_reg ( .D(g23000), .SI(g480), .SE(n8176), .CLK(n8363), .Q(
        g484) );
  SDFFX1 DFF_391_Q_reg ( .D(g23022), .SI(g484), .SE(n8176), .CLK(n8363), .Q(
        g464) );
  SDFFX1 DFF_392_Q_reg ( .D(g24206), .SI(g464), .SE(n8176), .CLK(n8363), .Q(
        g465) );
  SDFFX1 DFF_393_Q_reg ( .D(g24215), .SI(g465), .SE(n8176), .CLK(n8363), .Q(
        test_so24) );
  SDFFX1 DFF_394_Q_reg ( .D(g24228), .SI(test_si25), .SE(n8175), .CLK(n8362), 
        .Q(g471) );
  SDFFX1 DFF_395_Q_reg ( .D(n518), .SI(g471), .SE(n8176), .CLK(n8363), .Q(g528) );
  SDFFX1 DFF_396_Q_reg ( .D(g528), .SI(g528), .SE(n8176), .CLK(n8363), .Q(g535) );
  SDFFX1 DFF_397_Q_reg ( .D(g535), .SI(g535), .SE(n8176), .CLK(n8363), .Q(g542) );
  SDFFX1 DFF_398_Q_reg ( .D(g13149), .SI(g542), .SE(n8176), .CLK(n8363), .Q(
        g543) );
  SDFFX1 DFF_399_Q_reg ( .D(g543), .SI(g543), .SE(n8177), .CLK(n8364), .Q(g544) );
  SDFFX1 DFF_400_Q_reg ( .D(g21851), .SI(g544), .SE(n8177), .CLK(n8364), .Q(
        g548) );
  SDFFX1 DFF_401_Q_reg ( .D(g13111), .SI(g548), .SE(n8177), .CLK(n8364), .Q(
        g549) );
  SDFFX1 DFF_402_Q_reg ( .D(g549), .SI(g549), .SE(n8177), .CLK(n8364), .Q(g499), .QN(n4541) );
  SDFFX1 DFF_403_Q_reg ( .D(g13160), .SI(g499), .SE(n8177), .CLK(n8364), .Q(
        g558) );
  SDFFX1 DFF_404_Q_reg ( .D(g558), .SI(g558), .SE(n8177), .CLK(n8364), .Q(g559), .QN(n7756) );
  SDFFX1 DFF_405_Q_reg ( .D(g27261), .SI(g559), .SE(n8184), .CLK(n8371), .Q(
        g576), .QN(n7347) );
  SDFFX1 DFF_406_Q_reg ( .D(g27268), .SI(g576), .SE(n8185), .CLK(n8372), .Q(
        g577), .QN(n7349) );
  SDFFX1 DFF_407_Q_reg ( .D(g27279), .SI(g577), .SE(n8185), .CLK(n8372), .Q(
        g575), .QN(n7348) );
  SDFFX1 DFF_408_Q_reg ( .D(g27269), .SI(g575), .SE(n8185), .CLK(n8372), .Q(
        g579), .QN(n7359) );
  SDFFX1 DFF_409_Q_reg ( .D(g27280), .SI(g579), .SE(n8185), .CLK(n8372), .Q(
        test_so25), .QN(n8121) );
  SDFFX1 DFF_410_Q_reg ( .D(g27294), .SI(test_si26), .SE(n8185), .CLK(n8372), 
        .Q(g578), .QN(n7360) );
  SDFFX1 DFF_411_Q_reg ( .D(g27281), .SI(g578), .SE(n8185), .CLK(n8372), .Q(
        g582), .QN(n7184) );
  SDFFX1 DFF_412_Q_reg ( .D(g27295), .SI(g582), .SE(n8185), .CLK(n8372), .Q(
        g583), .QN(n7186) );
  SDFFX1 DFF_413_Q_reg ( .D(g27311), .SI(g583), .SE(n8185), .CLK(n8372), .Q(
        g581), .QN(n7185) );
  SDFFX1 DFF_414_Q_reg ( .D(g27296), .SI(g581), .SE(n8184), .CLK(n8371), .Q(
        g585), .QN(n7369) );
  SDFFX1 DFF_415_Q_reg ( .D(g27312), .SI(g585), .SE(n8185), .CLK(n8372), .Q(
        g586), .QN(n7371) );
  SDFFX1 DFF_416_Q_reg ( .D(g27327), .SI(g586), .SE(n8185), .CLK(n8372), .Q(
        g584), .QN(n7370) );
  SDFFX1 DFF_417_Q_reg ( .D(g24491), .SI(g584), .SE(n8185), .CLK(n8372), .Q(
        g587) );
  SDFFX1 DFF_418_Q_reg ( .D(g24498), .SI(g587), .SE(n8185), .CLK(n8372), .Q(
        g590) );
  SDFFX1 DFF_419_Q_reg ( .D(g24507), .SI(g590), .SE(n8186), .CLK(n8373), .Q(
        g593) );
  SDFFX1 DFF_420_Q_reg ( .D(g24499), .SI(g593), .SE(n8186), .CLK(n8373), .Q(
        g596) );
  SDFFX1 DFF_421_Q_reg ( .D(g24508), .SI(g596), .SE(n8186), .CLK(n8373), .Q(
        g599) );
  SDFFX1 DFF_422_Q_reg ( .D(g24519), .SI(g599), .SE(n8186), .CLK(n8373), .Q(
        g602) );
  SDFFX1 DFF_423_Q_reg ( .D(g28345), .SI(g602), .SE(n8186), .CLK(n8373), .Q(
        g614) );
  SDFFX1 DFF_424_Q_reg ( .D(g28349), .SI(g614), .SE(n8186), .CLK(n8373), .Q(
        g617) );
  SDFFX1 DFF_425_Q_reg ( .D(g28353), .SI(g617), .SE(n8186), .CLK(n8373), .Q(
        test_so26) );
  SDFFX1 DFF_426_Q_reg ( .D(g28342), .SI(test_si27), .SE(n8186), .CLK(n8373), 
        .Q(g605) );
  SDFFX1 DFF_427_Q_reg ( .D(g28344), .SI(g605), .SE(n8186), .CLK(n8373), .Q(
        g608) );
  SDFFX1 DFF_428_Q_reg ( .D(g28348), .SI(g608), .SE(n8186), .CLK(n8373), .Q(
        g611) );
  SDFFX1 DFF_429_Q_reg ( .D(g26541), .SI(g611), .SE(n8186), .CLK(n8373), .Q(
        g490) );
  SDFFX1 DFF_430_Q_reg ( .D(g26545), .SI(g490), .SE(n8186), .CLK(n8373), .Q(
        g493) );
  SDFFX1 DFF_431_Q_reg ( .D(g26553), .SI(g493), .SE(n8187), .CLK(n8374), .Q(
        g496) );
  SDFFX1 DFF_432_Q_reg ( .D(g499), .SI(g496), .SE(n8187), .CLK(n8374), .Q(g506), .QN(n4570) );
  SDFFX1 DFF_433_Q_reg ( .D(g22578), .SI(g506), .SE(n8187), .CLK(n8374), .Q(
        n4571), .QN(n7418) );
  SDFFX1 DFF_442_Q_reg ( .D(n533), .SI(n4571), .SE(n8187), .CLK(n8374), .Q(
        g16297), .QN(n8048) );
  SDFFX1 DFF_443_Q_reg ( .D(g16297), .SI(g16297), .SE(n8187), .CLK(n8374), .Q(
        g525), .QN(n8054) );
  SDFFX1 DFF_444_Q_reg ( .D(DFF_299_n1), .SI(g525), .SE(n8187), .CLK(n8374), 
        .Q(n8047), .QN(DFF_444_n1) );
  SDFFX1 DFF_445_Q_reg ( .D(DFF_301_n1), .SI(n8047), .SE(n8187), .CLK(n8374), 
        .Q(n8046), .QN(DFF_445_n1) );
  SDFFX1 DFF_446_Q_reg ( .D(DFF_303_n1), .SI(n8046), .SE(n8187), .CLK(n8374), 
        .Q(n8045), .QN(DFF_446_n1) );
  SDFFX1 DFF_447_Q_reg ( .D(DFF_305_n1), .SI(n8045), .SE(n8187), .CLK(n8374), 
        .Q(n8044), .QN(DFF_447_n1) );
  SDFFX1 DFF_448_Q_reg ( .D(DFF_307_n1), .SI(n8044), .SE(n8187), .CLK(n8374), 
        .Q(n8043), .QN(DFF_448_n1) );
  SDFFX1 DFF_449_Q_reg ( .D(DFF_309_n1), .SI(n8043), .SE(n8187), .CLK(n8374), 
        .Q(test_so27), .QN(DFF_449_n1) );
  SDFFX1 DFF_450_Q_reg ( .D(DFF_311_n1), .SI(test_si28), .SE(n8156), .CLK(
        n8343), .Q(g536), .QN(n7155) );
  SDFFX1 DFF_451_Q_reg ( .D(DFF_313_n1), .SI(g536), .SE(n8156), .CLK(n8343), 
        .Q(g537), .QN(n7154) );
  SDFFX1 DFF_452_Q_reg ( .D(g24059), .SI(g537), .SE(n8169), .CLK(n8356), .Q(
        g538), .QN(n4492) );
  SDFFX1 DFF_453_Q_reg ( .D(n4485), .SI(g538), .SE(n8169), .CLK(n8356), .Q(
        n8040), .QN(n14378) );
  SDFFX1 DFF_455_Q_reg ( .D(g6677), .SI(g6677), .SE(n8172), .CLK(n8359), .Q(
        g6911), .QN(n4359) );
  SDFFX1 DFF_456_Q_reg ( .D(g6911), .SI(g6911), .SE(n8173), .CLK(n8360), .Q(
        g629), .QN(n4295) );
  SDFFX1 DFF_457_Q_reg ( .D(g16654), .SI(g629), .SE(n8173), .CLK(n8360), .Q(
        g630), .QN(n7760) );
  SDFFX1 DFF_458_Q_reg ( .D(g20314), .SI(g630), .SE(n8180), .CLK(n8367), .Q(
        g659), .QN(n4429) );
  SDFFX1 DFF_459_Q_reg ( .D(g20682), .SI(g659), .SE(n8180), .CLK(n8367), .Q(
        g640), .QN(n4404) );
  SDFFX1 DFF_460_Q_reg ( .D(n615), .SI(g640), .SE(n8180), .CLK(n8367), .Q(g633), .QN(n4478) );
  SDFFX1 DFF_461_Q_reg ( .D(g23324), .SI(g633), .SE(n8180), .CLK(n8367), .Q(
        g653), .QN(n4422) );
  SDFFX1 DFF_462_Q_reg ( .D(g24426), .SI(g653), .SE(n8180), .CLK(n8367), .Q(
        g646), .QN(n4414) );
  SDFFX1 DFF_463_Q_reg ( .D(g25185), .SI(g646), .SE(n8180), .CLK(n8367), .Q(
        g660), .QN(n4403) );
  SDFFX1 DFF_464_Q_reg ( .D(n616), .SI(g660), .SE(n8180), .CLK(n8367), .Q(g672), .QN(n4413) );
  SDFFX1 DFF_465_Q_reg ( .D(g26776), .SI(g672), .SE(n8180), .CLK(n8367), .Q(
        test_so28), .QN(n8105) );
  SDFFX1 DFF_466_Q_reg ( .D(g27672), .SI(test_si29), .SE(n8180), .CLK(n8367), 
        .Q(g679), .QN(n4477) );
  SDFFX1 DFF_467_Q_reg ( .D(g28199), .SI(g679), .SE(n8180), .CLK(n8367), .Q(
        g686), .QN(n4396) );
  SDFFX1 DFF_468_Q_reg ( .D(g28668), .SI(g686), .SE(n8180), .CLK(n8367), .Q(
        g692), .QN(n4418) );
  SDFFX1 DFF_469_Q_reg ( .D(g20875), .SI(g692), .SE(n8187), .CLK(n8374), .Q(
        g699), .QN(n7838) );
  SDFFX1 DFF_470_Q_reg ( .D(g20879), .SI(g699), .SE(n8188), .CLK(n8375), .Q(
        g700), .QN(n7837) );
  SDFFX1 DFF_471_Q_reg ( .D(g20891), .SI(g700), .SE(n8188), .CLK(n8375), .Q(
        g698), .QN(n7876) );
  SDFFX1 DFF_472_Q_reg ( .D(g20880), .SI(g698), .SE(n8188), .CLK(n8375), .Q(
        g702), .QN(n7836) );
  SDFFX1 DFF_473_Q_reg ( .D(g20892), .SI(g702), .SE(n8188), .CLK(n8375), .Q(
        g703), .QN(n7835) );
  SDFFX1 DFF_474_Q_reg ( .D(g20901), .SI(g703), .SE(n8189), .CLK(n8376), .Q(
        g701), .QN(n7875) );
  SDFFX1 DFF_475_Q_reg ( .D(g20893), .SI(g701), .SE(n8189), .CLK(n8376), .Q(
        g705), .QN(n7834) );
  SDFFX1 DFF_476_Q_reg ( .D(g20902), .SI(g705), .SE(n8189), .CLK(n8376), .Q(
        g706), .QN(n7833) );
  SDFFX1 DFF_477_Q_reg ( .D(g20921), .SI(g706), .SE(n8189), .CLK(n8376), .Q(
        g704), .QN(n7874) );
  SDFFX1 DFF_478_Q_reg ( .D(g20903), .SI(g704), .SE(n8189), .CLK(n8376), .Q(
        g708), .QN(n7832) );
  SDFFX1 DFF_479_Q_reg ( .D(g20922), .SI(g708), .SE(n8189), .CLK(n8376), .Q(
        g709), .QN(n7831) );
  SDFFX1 DFF_480_Q_reg ( .D(g20944), .SI(g709), .SE(n8189), .CLK(n8376), .Q(
        g707), .QN(n7873) );
  SDFFX1 DFF_481_Q_reg ( .D(g20923), .SI(g707), .SE(n8189), .CLK(n8376), .Q(
        test_so29), .QN(n8137) );
  SDFFX1 DFF_482_Q_reg ( .D(g20945), .SI(test_si30), .SE(n8188), .CLK(n8375), 
        .Q(g712), .QN(n7830) );
  SDFFX1 DFF_483_Q_reg ( .D(g20966), .SI(g712), .SE(n8189), .CLK(n8376), .Q(
        g710), .QN(n7872) );
  SDFFX1 DFF_484_Q_reg ( .D(g20946), .SI(g710), .SE(n8189), .CLK(n8376), .Q(
        g714), .QN(n7829) );
  SDFFX1 DFF_485_Q_reg ( .D(g20967), .SI(g714), .SE(n8189), .CLK(n8376), .Q(
        g715), .QN(n7828) );
  SDFFX1 DFF_486_Q_reg ( .D(g20989), .SI(g715), .SE(n8189), .CLK(n8376), .Q(
        g713), .QN(n7871) );
  SDFFX1 DFF_487_Q_reg ( .D(g20968), .SI(g713), .SE(n8190), .CLK(n8377), .Q(
        g717), .QN(n7827) );
  SDFFX1 DFF_488_Q_reg ( .D(g20990), .SI(g717), .SE(n8190), .CLK(n8377), .Q(
        g718), .QN(n7826) );
  SDFFX1 DFF_489_Q_reg ( .D(g21009), .SI(g718), .SE(n8190), .CLK(n8377), .Q(
        g716), .QN(n7870) );
  SDFFX1 DFF_490_Q_reg ( .D(g20991), .SI(g716), .SE(n8190), .CLK(n8377), .Q(
        g720), .QN(n7825) );
  SDFFX1 DFF_491_Q_reg ( .D(g21010), .SI(g720), .SE(n8190), .CLK(n8377), .Q(
        g721), .QN(n7824) );
  SDFFX1 DFF_492_Q_reg ( .D(g21031), .SI(g721), .SE(n8190), .CLK(n8377), .Q(
        g719), .QN(n7869) );
  SDFFX1 DFF_493_Q_reg ( .D(g21011), .SI(g719), .SE(n8190), .CLK(n8377), .Q(
        g723), .QN(n7823) );
  SDFFX1 DFF_494_Q_reg ( .D(g21032), .SI(g723), .SE(n8190), .CLK(n8377), .Q(
        g724), .QN(n7822) );
  SDFFX1 DFF_495_Q_reg ( .D(g21051), .SI(g724), .SE(n8190), .CLK(n8377), .Q(
        g722), .QN(n7868) );
  SDFFX1 DFF_496_Q_reg ( .D(g20876), .SI(g722), .SE(n8190), .CLK(n8377), .Q(
        g726), .QN(n7821) );
  SDFFX1 DFF_497_Q_reg ( .D(g20881), .SI(g726), .SE(n8190), .CLK(n8377), .Q(
        test_so30), .QN(n8138) );
  SDFFX1 DFF_498_Q_reg ( .D(g20894), .SI(test_si31), .SE(n8188), .CLK(n8375), 
        .Q(g725), .QN(n7867) );
  SDFFX1 DFF_499_Q_reg ( .D(g20924), .SI(g725), .SE(n8188), .CLK(n8375), .Q(
        g729), .QN(n8038) );
  SDFFX1 DFF_500_Q_reg ( .D(g20947), .SI(g729), .SE(n8188), .CLK(n8375), .Q(
        g730), .QN(n7574) );
  SDFFX1 DFF_501_Q_reg ( .D(g20969), .SI(g730), .SE(n8188), .CLK(n8375), .Q(
        g728) );
  SDFFX1 DFF_502_Q_reg ( .D(g20948), .SI(g728), .SE(n8188), .CLK(n8375), .Q(
        g732), .QN(n7578) );
  SDFFX1 DFF_503_Q_reg ( .D(g20970), .SI(g732), .SE(n8188), .CLK(n8375), .Q(
        g733), .QN(n7573) );
  SDFFX1 DFF_504_Q_reg ( .D(g20992), .SI(g733), .SE(n8188), .CLK(n8375), .Q(
        g731), .QN(n7630) );
  SDFFX1 DFF_505_Q_reg ( .D(g25260), .SI(g731), .SE(n8190), .CLK(n8377), .Q(
        g735), .QN(n7509) );
  SDFFX1 DFF_506_Q_reg ( .D(g25262), .SI(g735), .SE(n8191), .CLK(n8378), .Q(
        g736), .QN(n7508) );
  SDFFX1 DFF_507_Q_reg ( .D(g25266), .SI(g736), .SE(n8191), .CLK(n8378), .Q(
        g734), .QN(n7513) );
  SDFFX1 DFF_508_Q_reg ( .D(g22218), .SI(g734), .SE(n8191), .CLK(n8378), .Q(
        g738), .QN(n7880) );
  SDFFX1 DFF_509_Q_reg ( .D(n586), .SI(g738), .SE(n8191), .CLK(n8378), .Q(g739), .QN(n7977) );
  SDFFX1 DFF_510_Q_reg ( .D(g22242), .SI(g739), .SE(n8191), .CLK(n8378), .Q(
        g737), .QN(n7989) );
  SDFFX1 DFF_511_Q_reg ( .D(g2950), .SI(g737), .SE(n8191), .CLK(n8378), .Q(
        g6368), .QN(n4323) );
  SDFFX1 DFF_512_Q_reg ( .D(g6368), .SI(g6368), .SE(n8191), .CLK(n8378), .Q(
        g6518), .QN(n4312) );
  SDFFX1 DFF_513_Q_reg ( .D(g6518), .SI(g6518), .SE(n8191), .CLK(n8378), .Q(
        test_so31), .QN(n8096) );
  SDFFX1 DFF_514_Q_reg ( .D(g22126), .SI(test_si32), .SE(n8192), .CLK(n8379), 
        .Q(g818), .QN(n7948) );
  SDFFX1 DFF_515_Q_reg ( .D(g22145), .SI(g818), .SE(n8195), .CLK(n8382), .Q(
        g819), .QN(n7947) );
  SDFFX1 DFF_516_Q_reg ( .D(g22162), .SI(g819), .SE(n8196), .CLK(n8383), .Q(
        g817), .QN(n7557) );
  SDFFX1 DFF_517_Q_reg ( .D(g22146), .SI(g817), .SE(n8192), .CLK(n8379), .Q(
        g821), .QN(n7939) );
  SDFFX1 DFF_518_Q_reg ( .D(g22163), .SI(g821), .SE(n8196), .CLK(n8383), .Q(
        g822), .QN(n7935) );
  SDFFX1 DFF_519_Q_reg ( .D(g22177), .SI(g822), .SE(n8196), .CLK(n8383), .Q(
        g820), .QN(n7556) );
  SDFFX1 DFF_520_Q_reg ( .D(g22029), .SI(g820), .SE(n8196), .CLK(n8383), .Q(
        g830), .QN(n7934) );
  SDFFX1 DFF_521_Q_reg ( .D(g22033), .SI(g830), .SE(n8196), .CLK(n8383), .Q(
        g831), .QN(n7933) );
  SDFFX1 DFF_522_Q_reg ( .D(g22040), .SI(g831), .SE(n8196), .CLK(n8383), .Q(
        g829), .QN(n7555) );
  SDFFX1 DFF_523_Q_reg ( .D(g22034), .SI(g829), .SE(n8196), .CLK(n8383), .Q(
        g833), .QN(n7932) );
  SDFFX1 DFF_524_Q_reg ( .D(g22041), .SI(g833), .SE(n8196), .CLK(n8383), .Q(
        g834), .QN(n7931) );
  SDFFX1 DFF_525_Q_reg ( .D(g22054), .SI(g834), .SE(n8197), .CLK(n8384), .Q(
        g832), .QN(n7554) );
  SDFFX1 DFF_526_Q_reg ( .D(g22042), .SI(g832), .SE(n8197), .CLK(n8384), .Q(
        g836), .QN(n7928) );
  SDFFX1 DFF_527_Q_reg ( .D(g22055), .SI(g836), .SE(n8197), .CLK(n8384), .Q(
        g837), .QN(n7927) );
  SDFFX1 DFF_528_Q_reg ( .D(g22066), .SI(g837), .SE(n8197), .CLK(n8384), .Q(
        g835), .QN(n7553) );
  SDFFX1 DFF_529_Q_reg ( .D(g22056), .SI(g835), .SE(n8197), .CLK(n8384), .Q(
        test_so32), .QN(n8125) );
  SDFFX1 DFF_530_Q_reg ( .D(g22067), .SI(test_si33), .SE(n8194), .CLK(n8381), 
        .Q(g840), .QN(n7919) );
  SDFFX1 DFF_531_Q_reg ( .D(g22087), .SI(g840), .SE(n8195), .CLK(n8382), .Q(
        g838), .QN(n7552) );
  SDFFX1 DFF_532_Q_reg ( .D(g22068), .SI(g838), .SE(n8195), .CLK(n8382), .Q(
        g842), .QN(n7917) );
  SDFFX1 DFF_533_Q_reg ( .D(g22088), .SI(g842), .SE(n8195), .CLK(n8382), .Q(
        g843), .QN(n7916) );
  SDFFX1 DFF_534_Q_reg ( .D(g22104), .SI(g843), .SE(n8195), .CLK(n8382), .Q(
        g841), .QN(n7551) );
  SDFFX1 DFF_535_Q_reg ( .D(g22089), .SI(g841), .SE(n8195), .CLK(n8382), .Q(
        g845), .QN(n7915) );
  SDFFX1 DFF_536_Q_reg ( .D(g22105), .SI(g845), .SE(n8195), .CLK(n8382), .Q(
        g846), .QN(n7914) );
  SDFFX1 DFF_537_Q_reg ( .D(g22127), .SI(g846), .SE(n8195), .CLK(n8382), .Q(
        g844), .QN(n7550) );
  SDFFX1 DFF_538_Q_reg ( .D(g22106), .SI(g844), .SE(n8195), .CLK(n8382), .Q(
        g848), .QN(n7549) );
  SDFFX1 DFF_539_Q_reg ( .D(g22128), .SI(g848), .SE(n8195), .CLK(n8382), .Q(
        g849), .QN(n7548) );
  SDFFX1 DFF_540_Q_reg ( .D(g22147), .SI(g849), .SE(n8195), .CLK(n8382), .Q(
        g847), .QN(n7547) );
  SDFFX1 DFF_541_Q_reg ( .D(g22129), .SI(g847), .SE(n8195), .CLK(n8382), .Q(
        g851), .QN(n7546) );
  SDFFX1 DFF_542_Q_reg ( .D(g22148), .SI(g851), .SE(n8196), .CLK(n8383), .Q(
        g852), .QN(n7545) );
  SDFFX1 DFF_543_Q_reg ( .D(g22164), .SI(g852), .SE(n8196), .CLK(n8383), .Q(
        g850), .QN(n7544) );
  SDFFX1 DFF_544_Q_reg ( .D(g25209), .SI(g850), .SE(n8196), .CLK(n8383), .Q(
        g857), .QN(n7612) );
  SDFFX1 DFF_545_Q_reg ( .D(g25214), .SI(g857), .SE(n8196), .CLK(n8383), .Q(
        test_so33), .QN(n8117) );
  SDFFX1 DFF_546_Q_reg ( .D(g25221), .SI(test_si34), .SE(n8191), .CLK(n8378), 
        .Q(g856), .QN(n7611) );
  SDFFX1 DFF_547_Q_reg ( .D(g25215), .SI(g856), .SE(n8191), .CLK(n8378), .Q(
        g860), .QN(n7610) );
  SDFFX1 DFF_548_Q_reg ( .D(g25222), .SI(g860), .SE(n8191), .CLK(n8378), .Q(
        g861), .QN(n7609) );
  SDFFX1 DFF_549_Q_reg ( .D(g25230), .SI(g861), .SE(n8191), .CLK(n8378), .Q(
        g859), .QN(n7608) );
  SDFFX1 DFF_550_Q_reg ( .D(g25223), .SI(g859), .SE(n8192), .CLK(n8379), .Q(
        g863), .QN(n7607) );
  SDFFX1 DFF_551_Q_reg ( .D(g25231), .SI(g863), .SE(n8192), .CLK(n8379), .Q(
        g864), .QN(n7606) );
  SDFFX1 DFF_552_Q_reg ( .D(g25240), .SI(g864), .SE(n8192), .CLK(n8379), .Q(
        g862), .QN(n7605) );
  SDFFX1 DFF_553_Q_reg ( .D(g25232), .SI(g862), .SE(n8192), .CLK(n8379), .Q(
        g866), .QN(n7604) );
  SDFFX1 DFF_554_Q_reg ( .D(g25241), .SI(g866), .SE(n8192), .CLK(n8379), .Q(
        g867), .QN(n7603) );
  SDFFX1 DFF_555_Q_reg ( .D(g25248), .SI(g867), .SE(n8192), .CLK(n8379), .Q(
        g865), .QN(n7602) );
  SDFFX1 DFF_556_Q_reg ( .D(g30269), .SI(g865), .SE(n8203), .CLK(n8390), .Q(
        g873) );
  SDFFX1 DFF_557_Q_reg ( .D(g30277), .SI(g873), .SE(n8203), .CLK(n8390), .Q(
        g876) );
  SDFFX1 DFF_558_Q_reg ( .D(g30285), .SI(g876), .SE(n8203), .CLK(n8390), .Q(
        g879) );
  SDFFX1 DFF_559_Q_reg ( .D(g30643), .SI(g879), .SE(n8203), .CLK(n8390), .Q(
        g918) );
  SDFFX1 DFF_560_Q_reg ( .D(g30648), .SI(g918), .SE(n8203), .CLK(n8390), .Q(
        g921) );
  SDFFX1 DFF_561_Q_reg ( .D(g30654), .SI(g921), .SE(n8199), .CLK(n8386), .Q(
        test_so34) );
  SDFFX1 DFF_562_Q_reg ( .D(g30676), .SI(test_si35), .SE(n8192), .CLK(n8379), 
        .Q(g882) );
  SDFFX1 DFF_563_Q_reg ( .D(g30681), .SI(g882), .SE(n8192), .CLK(n8379), .Q(
        g885) );
  SDFFX1 DFF_564_Q_reg ( .D(g30687), .SI(g885), .SE(n8193), .CLK(n8380), .Q(
        g888) );
  SDFFX1 DFF_565_Q_reg ( .D(g30649), .SI(g888), .SE(n8197), .CLK(n8384), .Q(
        g927) );
  SDFFX1 DFF_566_Q_reg ( .D(g30655), .SI(g927), .SE(n8197), .CLK(n8384), .Q(
        g930) );
  SDFFX1 DFF_567_Q_reg ( .D(g30662), .SI(g930), .SE(n8197), .CLK(n8384), .Q(
        g933) );
  SDFFX1 DFF_568_Q_reg ( .D(g30286), .SI(g933), .SE(n8197), .CLK(n8384), .Q(
        g891) );
  SDFFX1 DFF_569_Q_reg ( .D(g30293), .SI(g891), .SE(n8197), .CLK(n8384), .Q(
        g894) );
  SDFFX1 DFF_570_Q_reg ( .D(g30298), .SI(g894), .SE(n8197), .CLK(n8384), .Q(
        g897) );
  SDFFX1 DFF_571_Q_reg ( .D(g30259), .SI(g897), .SE(n8197), .CLK(n8384), .Q(
        g936) );
  SDFFX1 DFF_572_Q_reg ( .D(g30264), .SI(g936), .SE(n8198), .CLK(n8385), .Q(
        g939) );
  SDFFX1 DFF_573_Q_reg ( .D(g30270), .SI(g939), .SE(n8198), .CLK(n8385), .Q(
        g942) );
  SDFFX1 DFF_574_Q_reg ( .D(g30247), .SI(g942), .SE(n8198), .CLK(n8385), .Q(
        g900) );
  SDFFX1 DFF_575_Q_reg ( .D(g30249), .SI(g900), .SE(n8198), .CLK(n8385), .Q(
        g903) );
  SDFFX1 DFF_576_Q_reg ( .D(g30251), .SI(g903), .SE(n8198), .CLK(n8385), .Q(
        g906) );
  SDFFX1 DFF_577_Q_reg ( .D(g30265), .SI(g906), .SE(n8198), .CLK(n8385), .Q(
        test_so35) );
  SDFFX1 DFF_578_Q_reg ( .D(g30271), .SI(test_si36), .SE(n8198), .CLK(n8385), 
        .Q(g948) );
  SDFFX1 DFF_579_Q_reg ( .D(g30278), .SI(g948), .SE(n8198), .CLK(n8385), .Q(
        g951) );
  SDFFX1 DFF_580_Q_reg ( .D(g30638), .SI(g951), .SE(n8198), .CLK(n8385), .Q(
        g909) );
  SDFFX1 DFF_581_Q_reg ( .D(g30642), .SI(g909), .SE(n8199), .CLK(n8386), .Q(
        g912) );
  SDFFX1 DFF_582_Q_reg ( .D(g30647), .SI(g912), .SE(n8198), .CLK(n8385), .Q(
        g915) );
  SDFFX1 DFF_583_Q_reg ( .D(g30670), .SI(g915), .SE(n8198), .CLK(n8385), .Q(
        g954) );
  SDFFX1 DFF_584_Q_reg ( .D(g30677), .SI(g954), .SE(n8198), .CLK(n8385), .Q(
        g957) );
  SDFFX1 DFF_585_Q_reg ( .D(g30682), .SI(g957), .SE(n8193), .CLK(n8380), .Q(
        g960) );
  SDFFX1 DFF_586_Q_reg ( .D(g25042), .SI(g960), .SE(n8193), .CLK(n8380), .Q(
        g780), .QN(n7710) );
  SDFFX1 DFF_587_Q_reg ( .D(g25935), .SI(g780), .SE(n8193), .CLK(n8380), .Q(
        g776), .QN(n8085) );
  SDFFX1 DFF_588_Q_reg ( .D(g26530), .SI(g776), .SE(n8193), .CLK(n8380), .Q(
        g771), .QN(n7709) );
  SDFFX1 DFF_589_Q_reg ( .D(g27123), .SI(g771), .SE(n8193), .CLK(n8380), .Q(
        g767), .QN(n8091) );
  SDFFX1 DFF_590_Q_reg ( .D(g27603), .SI(g767), .SE(n8193), .CLK(n8380), .Q(
        g762), .QN(n7708) );
  SDFFX1 DFF_591_Q_reg ( .D(g28146), .SI(g762), .SE(n8193), .CLK(n8380), .Q(
        g758), .QN(n8092) );
  SDFFX1 DFF_592_Q_reg ( .D(g28635), .SI(g758), .SE(n8193), .CLK(n8380), .Q(
        g753), .QN(n7707) );
  SDFFX1 DFF_593_Q_reg ( .D(g29110), .SI(g753), .SE(n8193), .CLK(n8380), .Q(
        test_so36) );
  SDFFX1 DFF_594_Q_reg ( .D(g29354), .SI(test_si37), .SE(n8193), .CLK(n8380), 
        .Q(g744), .QN(n7336) );
  SDFFX1 DFF_595_Q_reg ( .D(g29580), .SI(g744), .SE(n8193), .CLK(n8380), .Q(
        g740), .QN(n7175) );
  SDFFX1 DFF_596_Q_reg ( .D(n15), .SI(g740), .SE(n8194), .CLK(n8381), .Q(g868)
         );
  SDFFX1 DFF_597_Q_reg ( .D(g868), .SI(g868), .SE(n8194), .CLK(n8381), .Q(
        g5595) );
  SDFFX1 DFF_598_Q_reg ( .D(g5595), .SI(g5595), .SE(n8194), .CLK(n8381), .Q(
        g869), .QN(n7720) );
  SDFFX1 DFF_599_Q_reg ( .D(g2950), .SI(g869), .SE(n8194), .CLK(n8381), .Q(
        g5472), .QN(n4363) );
  SDFFX1 DFF_600_Q_reg ( .D(g5472), .SI(g5472), .SE(n8194), .CLK(n8381), .Q(
        g6712), .QN(n4364) );
  SDFFX1 DFF_601_Q_reg ( .D(g6712), .SI(g6712), .SE(n8194), .CLK(n8381), .Q(
        g1088), .QN(n4381) );
  SDFFX1 DFF_602_Q_reg ( .D(g5595), .SI(g1088), .SE(n8194), .CLK(n8381), .Q(
        g996), .QN(n4387) );
  SDFFX1 DFF_603_Q_reg ( .D(g27257), .SI(g996), .SE(n8202), .CLK(n8389), .Q(
        g1041), .QN(n7663) );
  SDFFX1 DFF_604_Q_reg ( .D(g27262), .SI(g1041), .SE(n8202), .CLK(n8389), .Q(
        g1030), .QN(n7662) );
  SDFFX1 DFF_605_Q_reg ( .D(g27270), .SI(g1030), .SE(n8202), .CLK(n8389), .Q(
        g1033), .QN(n7661) );
  SDFFX1 DFF_606_Q_reg ( .D(g27263), .SI(g1033), .SE(n8202), .CLK(n8389), .Q(
        g1056), .QN(n7640) );
  SDFFX1 DFF_607_Q_reg ( .D(g27271), .SI(g1056), .SE(n8202), .CLK(n8389), .Q(
        g1045), .QN(n7639) );
  SDFFX1 DFF_608_Q_reg ( .D(g27282), .SI(g1045), .SE(n8202), .CLK(n8389), .Q(
        g1048), .QN(n7638) );
  SDFFX1 DFF_609_Q_reg ( .D(g27272), .SI(g1048), .SE(n8202), .CLK(n8389), .Q(
        test_so37), .QN(n8114) );
  SDFFX1 DFF_610_Q_reg ( .D(g27283), .SI(test_si38), .SE(n8202), .CLK(n8389), 
        .Q(g1060), .QN(n7389) );
  SDFFX1 DFF_611_Q_reg ( .D(g27297), .SI(g1060), .SE(n8202), .CLK(n8389), .Q(
        g1063), .QN(n7390) );
  SDFFX1 DFF_612_Q_reg ( .D(g27284), .SI(g1063), .SE(n8203), .CLK(n8390), .Q(
        g1085), .QN(n7651) );
  SDFFX1 DFF_613_Q_reg ( .D(g27298), .SI(g1085), .SE(n8203), .CLK(n8390), .Q(
        g1075), .QN(n7650) );
  SDFFX1 DFF_614_Q_reg ( .D(g27313), .SI(g1075), .SE(n8200), .CLK(n8387), .Q(
        g1078), .QN(n7649) );
  SDFFX1 DFF_615_Q_reg ( .D(g28738), .SI(g1078), .SE(n8200), .CLK(n8387), .Q(
        g1095) );
  SDFFX1 DFF_616_Q_reg ( .D(g28746), .SI(g1095), .SE(n8201), .CLK(n8388), .Q(
        g1098) );
  SDFFX1 DFF_617_Q_reg ( .D(g28758), .SI(g1098), .SE(n8201), .CLK(n8388), .Q(
        g1101) );
  SDFFX1 DFF_618_Q_reg ( .D(g29198), .SI(g1101), .SE(n8202), .CLK(n8389), .Q(
        g1104) );
  SDFFX1 DFF_619_Q_reg ( .D(g29204), .SI(g1104), .SE(n8202), .CLK(n8389), .Q(
        g1107) );
  SDFFX1 DFF_620_Q_reg ( .D(g29209), .SI(g1107), .SE(n8200), .CLK(n8387), .Q(
        g1110) );
  SDFFX1 DFF_621_Q_reg ( .D(g28747), .SI(g1110), .SE(n8200), .CLK(n8387), .Q(
        g1114), .QN(n7689) );
  SDFFX1 DFF_622_Q_reg ( .D(g28759), .SI(g1114), .SE(n8200), .CLK(n8387), .Q(
        g1115), .QN(n7674) );
  SDFFX1 DFF_623_Q_reg ( .D(g28767), .SI(g1115), .SE(n8200), .CLK(n8387), .Q(
        g1113), .QN(n7688) );
  SDFFX1 DFF_624_Q_reg ( .D(g26806), .SI(g1113), .SE(n8200), .CLK(n8387), .Q(
        g1116) );
  SDFFX1 DFF_625_Q_reg ( .D(g26809), .SI(g1116), .SE(n8201), .CLK(n8388), .Q(
        test_so38) );
  SDFFX1 DFF_626_Q_reg ( .D(g26813), .SI(test_si39), .SE(n8201), .CLK(n8388), 
        .Q(g1122) );
  SDFFX1 DFF_627_Q_reg ( .D(g26810), .SI(g1122), .SE(n8201), .CLK(n8388), .Q(
        g1125) );
  SDFFX1 DFF_628_Q_reg ( .D(g26814), .SI(g1125), .SE(n8201), .CLK(n8388), .Q(
        g1128) );
  SDFFX1 DFF_629_Q_reg ( .D(g26818), .SI(g1128), .SE(n8201), .CLK(n8388), .Q(
        g1131) );
  SDFFX1 DFF_630_Q_reg ( .D(g27761), .SI(g1131), .SE(n8201), .CLK(n8388), .Q(
        g1135), .QN(n7687) );
  SDFFX1 DFF_631_Q_reg ( .D(g27763), .SI(g1135), .SE(n8201), .CLK(n8388), .Q(
        g1136), .QN(n7673) );
  SDFFX1 DFF_632_Q_reg ( .D(g27765), .SI(g1136), .SE(n8201), .CLK(n8388), .Q(
        g1134), .QN(n7686) );
  SDFFX1 DFF_633_Q_reg ( .D(g29609), .SI(g1134), .SE(n8201), .CLK(n8388), .Q(
        g999), .QN(n7293) );
  SDFFX1 DFF_634_Q_reg ( .D(g29612), .SI(g999), .SE(n8201), .CLK(n8388), .Q(
        g1000), .QN(n7276) );
  SDFFX1 DFF_635_Q_reg ( .D(g29616), .SI(g1000), .SE(n8200), .CLK(n8387), .Q(
        g1001), .QN(n7292) );
  SDFFX1 DFF_636_Q_reg ( .D(g30701), .SI(g1001), .SE(n8192), .CLK(n8379), .Q(
        g1002), .QN(n7291) );
  SDFFX1 DFF_637_Q_reg ( .D(g30703), .SI(g1002), .SE(n8194), .CLK(n8381), .Q(
        g1003), .QN(n7275) );
  SDFFX1 DFF_638_Q_reg ( .D(g30705), .SI(g1003), .SE(n8194), .CLK(n8381), .Q(
        g1004), .QN(n7290) );
  SDFFX1 DFF_639_Q_reg ( .D(g30470), .SI(g1004), .SE(n8192), .CLK(n8379), .Q(
        g1005), .QN(n7289) );
  SDFFX1 DFF_640_Q_reg ( .D(g30485), .SI(g1005), .SE(n8194), .CLK(n8381), .Q(
        g1006), .QN(n7274) );
  SDFFX1 DFF_641_Q_reg ( .D(g30500), .SI(g1006), .SE(n8194), .CLK(n8381), .Q(
        test_so39), .QN(n8139) );
  SDFFX1 DFF_642_Q_reg ( .D(g29170), .SI(test_si40), .SE(n8203), .CLK(n8390), 
        .Q(g1009), .QN(n7330) );
  SDFFX1 DFF_643_Q_reg ( .D(g29173), .SI(g1009), .SE(n8203), .CLK(n8390), .Q(
        g1010), .QN(n7324) );
  SDFFX1 DFF_644_Q_reg ( .D(g29179), .SI(g1010), .SE(n8199), .CLK(n8386), .Q(
        g1008), .QN(n7329) );
  SDFFX1 DFF_645_Q_reg ( .D(g26661), .SI(g1008), .SE(n8199), .CLK(n8386), .Q(
        g1090), .QN(n7685) );
  SDFFX1 DFF_646_Q_reg ( .D(g26665), .SI(g1090), .SE(n8199), .CLK(n8386), .Q(
        g1091), .QN(n7672) );
  SDFFX1 DFF_647_Q_reg ( .D(g26669), .SI(g1091), .SE(n8199), .CLK(n8386), .Q(
        g1089), .QN(n7684) );
  SDFFX1 DFF_648_Q_reg ( .D(n4289), .SI(g1089), .SE(n8199), .CLK(n8386), .Q(
        g1137) );
  SDFFX1 DFF_649_Q_reg ( .D(g1137), .SI(g1137), .SE(n8199), .CLK(n8386), .Q(
        n8027), .QN(DFF_649_n1) );
  SDFFX1 DFF_650_Q_reg ( .D(n4567), .SI(n8027), .SE(n8199), .CLK(n8386), .Q(
        g1139) );
  SDFFX1 DFF_651_Q_reg ( .D(g1139), .SI(g1139), .SE(n8199), .CLK(n8386), .Q(
        n8026), .QN(DFF_651_n1) );
  SDFFX1 DFF_652_Q_reg ( .D(n4559), .SI(n8026), .SE(n8199), .CLK(n8386), .Q(
        g1141) );
  SDFFX1 DFF_653_Q_reg ( .D(g1141), .SI(g1141), .SE(n8199), .CLK(n8386), .Q(
        n8025), .QN(DFF_653_n1) );
  SDFFX1 DFF_654_Q_reg ( .D(n4327), .SI(n8025), .SE(n8200), .CLK(n8387), .Q(
        g967) );
  SDFFX1 DFF_655_Q_reg ( .D(g967), .SI(g967), .SE(n8200), .CLK(n8387), .Q(
        n8024), .QN(DFF_655_n1) );
  SDFFX1 DFF_656_Q_reg ( .D(n4391), .SI(n8024), .SE(n8200), .CLK(n8387), .Q(
        g969) );
  SDFFX1 DFF_657_Q_reg ( .D(g969), .SI(g969), .SE(n8200), .CLK(n8387), .Q(
        test_so40), .QN(DFF_657_n1) );
  SDFFX1 DFF_658_Q_reg ( .D(n4321), .SI(test_si41), .SE(n8150), .CLK(n8337), 
        .Q(g971) );
  SDFFX1 DFF_659_Q_reg ( .D(g971), .SI(g971), .SE(n8150), .CLK(n8337), .Q(
        n8021), .QN(DFF_659_n1) );
  SDFFX1 DFF_660_Q_reg ( .D(n4375), .SI(n8021), .SE(n8150), .CLK(n8337), .Q(
        g973) );
  SDFFX1 DFF_661_Q_reg ( .D(g973), .SI(g973), .SE(n8151), .CLK(n8338), .Q(
        n8020), .QN(DFF_661_n1) );
  SDFFX1 DFF_662_Q_reg ( .D(n4379), .SI(n8020), .SE(n8151), .CLK(n8338), .Q(
        g975) );
  SDFFX1 DFF_663_Q_reg ( .D(g975), .SI(g975), .SE(n8151), .CLK(n8338), .Q(
        n8019), .QN(DFF_663_n1) );
  SDFFX1 DFF_664_Q_reg ( .D(g2873), .SI(n8019), .SE(n8151), .CLK(n8338), .Q(
        g977) );
  SDFFX1 DFF_665_Q_reg ( .D(g977), .SI(g977), .SE(n8151), .CLK(n8338), .Q(
        n8018), .QN(n4486) );
  SDFFX1 DFF_666_Q_reg ( .D(n4283), .SI(n8018), .SE(n8202), .CLK(n8389), .Q(
        g986), .QN(n4432) );
  SDFFX1 DFF_667_Q_reg ( .D(n457), .SI(g986), .SE(n8203), .CLK(n8390), .Q(g992), .QN(n7717) );
  SDFFX1 DFF_678_Q_reg ( .D(n4277), .SI(g992), .SE(n8203), .CLK(n8390), .Q(
        n8017) );
  SDFFX1 DFF_679_Q_reg ( .D(g1041), .SI(n8017), .SE(n8203), .CLK(n8390), .Q(
        g1029) );
  SDFFX1 DFF_680_Q_reg ( .D(g1029), .SI(g1029), .SE(n8204), .CLK(n8391), .Q(
        g1036) );
  SDFFX1 DFF_681_Q_reg ( .D(g1030), .SI(g1036), .SE(n8204), .CLK(n8391), .Q(
        g1037) );
  SDFFX1 DFF_682_Q_reg ( .D(g1037), .SI(g1037), .SE(n8204), .CLK(n8391), .Q(
        g1038) );
  SDFFX1 DFF_683_Q_reg ( .D(g1033), .SI(g1038), .SE(n8204), .CLK(n8391), .Q(
        test_so41) );
  SDFFX1 DFF_684_Q_reg ( .D(test_so41), .SI(test_si42), .SE(n8204), .CLK(n8391), .Q(g1040) );
  SDFFX1 DFF_685_Q_reg ( .D(g1056), .SI(g1040), .SE(n8204), .CLK(n8391), .Q(
        g1044) );
  SDFFX1 DFF_686_Q_reg ( .D(g1044), .SI(g1044), .SE(n8204), .CLK(n8391), .Q(
        g1051) );
  SDFFX1 DFF_687_Q_reg ( .D(g1045), .SI(g1051), .SE(n8204), .CLK(n8391), .Q(
        g1052) );
  SDFFX1 DFF_688_Q_reg ( .D(g1052), .SI(g1052), .SE(n8204), .CLK(n8391), .Q(
        g1053) );
  SDFFX1 DFF_689_Q_reg ( .D(g1048), .SI(g1053), .SE(n8204), .CLK(n8391), .Q(
        g1054) );
  SDFFX1 DFF_690_Q_reg ( .D(g1054), .SI(g1054), .SE(n8204), .CLK(n8391), .Q(
        g1055) );
  SDFFX1 DFF_691_Q_reg ( .D(test_so37), .SI(g1055), .SE(n8204), .CLK(n8391), 
        .Q(g1059) );
  SDFFX1 DFF_692_Q_reg ( .D(g1059), .SI(g1059), .SE(n8205), .CLK(n8392), .Q(
        g1066) );
  SDFFX1 DFF_693_Q_reg ( .D(g1060), .SI(g1066), .SE(n8205), .CLK(n8392), .Q(
        g1067) );
  SDFFX1 DFF_694_Q_reg ( .D(g1067), .SI(g1067), .SE(n8205), .CLK(n8392), .Q(
        g1068) );
  SDFFX1 DFF_695_Q_reg ( .D(g1063), .SI(g1068), .SE(n8205), .CLK(n8392), .Q(
        g1069) );
  SDFFX1 DFF_696_Q_reg ( .D(g1069), .SI(g1069), .SE(n8205), .CLK(n8392), .Q(
        g1070) );
  SDFFX1 DFF_697_Q_reg ( .D(g1085), .SI(g1070), .SE(n8205), .CLK(n8392), .Q(
        g1074) );
  SDFFX1 DFF_698_Q_reg ( .D(g1074), .SI(g1074), .SE(n8205), .CLK(n8392), .Q(
        g1081) );
  SDFFX1 DFF_699_Q_reg ( .D(g1075), .SI(g1081), .SE(n8205), .CLK(n8392), .Q(
        test_so42) );
  SDFFX1 DFF_700_Q_reg ( .D(test_so42), .SI(test_si43), .SE(n8205), .CLK(n8392), .Q(g1083) );
  SDFFX1 DFF_701_Q_reg ( .D(g1078), .SI(g1083), .SE(n8205), .CLK(n8392), .Q(
        g1084) );
  SDFFX1 DFF_702_Q_reg ( .D(g1084), .SI(g1084), .SE(n8205), .CLK(n8392), .Q(
        g1011) );
  SDFFX1 DFF_703_Q_reg ( .D(n4598), .SI(g1011), .SE(n8205), .CLK(n8392), .Q(
        g5657) );
  SDFFX1 DFF_704_Q_reg ( .D(g5657), .SI(g5657), .SE(n8206), .CLK(n8393), .Q(
        g5686) );
  SDFFX1 DFF_705_Q_reg ( .D(g5686), .SI(g5686), .SE(n8206), .CLK(n8393), .Q(
        g1024) );
  SDFFX1 DFF_706_Q_reg ( .D(n4598), .SI(g1024), .SE(n8206), .CLK(n8393), .Q(
        g6750), .QN(n4371) );
  SDFFX1 DFF_707_Q_reg ( .D(g6750), .SI(g6750), .SE(n8206), .CLK(n8393), .Q(
        g6944), .QN(n4316) );
  SDFFX1 DFF_708_Q_reg ( .D(g6944), .SI(g6944), .SE(n8206), .CLK(n8393), .Q(
        g1236), .QN(n4300) );
  SDFFX1 DFF_709_Q_reg ( .D(n837), .SI(g1236), .SE(n8206), .CLK(n8393), .Q(
        g1240), .QN(n7992) );
  SDFFX1 DFF_710_Q_reg ( .D(g18707), .SI(g1240), .SE(n8206), .CLK(n8393), .Q(
        g1243), .QN(n4353) );
  SDFFX1 DFF_711_Q_reg ( .D(g18763), .SI(g1243), .SE(n8206), .CLK(n8393), .Q(
        g1196), .QN(n4304) );
  SDFFX1 DFF_712_Q_reg ( .D(n819), .SI(g1196), .SE(n8207), .CLK(n8394), .Q(
        g1199) );
  SDFFX1 DFF_713_Q_reg ( .D(g1199), .SI(g1199), .SE(n8207), .CLK(n8394), .Q(
        g1209) );
  SDFFX1 DFF_714_Q_reg ( .D(g1209), .SI(g1209), .SE(n8207), .CLK(n8394), .Q(
        g1210) );
  SDFFX1 DFF_715_Q_reg ( .D(g1142), .SI(g1210), .SE(n8207), .CLK(n8394), .Q(
        test_so43) );
  SDFFX1 DFF_716_Q_reg ( .D(test_so43), .SI(test_si44), .SE(n8208), .CLK(n8395), .Q(g1255) );
  SDFFX1 DFF_717_Q_reg ( .D(g1145), .SI(g1255), .SE(n8208), .CLK(n8395), .Q(
        g1256) );
  SDFFX1 DFF_718_Q_reg ( .D(g1256), .SI(g1256), .SE(n8208), .CLK(n8395), .Q(
        g1257) );
  SDFFX1 DFF_719_Q_reg ( .D(g1148), .SI(g1257), .SE(n8208), .CLK(n8395), .Q(
        g1258) );
  SDFFX1 DFF_720_Q_reg ( .D(g1258), .SI(g1258), .SE(n8208), .CLK(n8395), .Q(
        g1259) );
  SDFFX1 DFF_721_Q_reg ( .D(g1152), .SI(g1259), .SE(n8208), .CLK(n8395), .Q(
        g1260) );
  SDFFX1 DFF_722_Q_reg ( .D(g1260), .SI(g1260), .SE(n8208), .CLK(n8395), .Q(
        g1251) );
  SDFFX1 DFF_723_Q_reg ( .D(g1155), .SI(g1251), .SE(n8208), .CLK(n8395), .Q(
        g1252) );
  SDFFX1 DFF_724_Q_reg ( .D(g1252), .SI(g1252), .SE(n8208), .CLK(n8395), .Q(
        g1253) );
  SDFFX1 DFF_725_Q_reg ( .D(g1158), .SI(g1253), .SE(n8208), .CLK(n8395), .Q(
        g1254) );
  SDFFX1 DFF_726_Q_reg ( .D(g1254), .SI(g1254), .SE(n8208), .CLK(n8395), .Q(
        g1176) );
  SDFFX1 DFF_727_Q_reg ( .D(g2950), .SI(g1176), .SE(n8208), .CLK(n8395), .Q(
        g7961), .QN(n4460) );
  SDFFX1 DFF_728_Q_reg ( .D(g7961), .SI(g7961), .SE(n8209), .CLK(n8396), .Q(
        g8007), .QN(n4459) );
  SDFFX1 DFF_729_Q_reg ( .D(g8007), .SI(g8007), .SE(n8209), .CLK(n8396), .Q(
        g1172), .QN(n4465) );
  SDFFX1 DFF_730_Q_reg ( .D(g23081), .SI(g1172), .SE(n8209), .CLK(n8396), .Q(
        g1173) );
  SDFFX1 DFF_731_Q_reg ( .D(g23111), .SI(g1173), .SE(n8209), .CLK(n8396), .Q(
        test_so44) );
  SDFFX1 DFF_732_Q_reg ( .D(g23126), .SI(test_si45), .SE(n8209), .CLK(n8396), 
        .Q(g1175) );
  SDFFX1 DFF_733_Q_reg ( .D(g23392), .SI(g1175), .SE(n8209), .CLK(n8396), .Q(
        g1142) );
  SDFFX1 DFF_734_Q_reg ( .D(g23406), .SI(g1142), .SE(n8209), .CLK(n8396), .Q(
        g1145) );
  SDFFX1 DFF_735_Q_reg ( .D(g24179), .SI(g1145), .SE(n8209), .CLK(n8396), .Q(
        g1148) );
  SDFFX1 DFF_736_Q_reg ( .D(g24181), .SI(g1148), .SE(n8209), .CLK(n8396), .Q(
        g1164) );
  SDFFX1 DFF_737_Q_reg ( .D(g24213), .SI(g1164), .SE(n8209), .CLK(n8396), .Q(
        g1165) );
  SDFFX1 DFF_738_Q_reg ( .D(g24223), .SI(g1165), .SE(n8209), .CLK(n8396), .Q(
        g1166) );
  SDFFX1 DFF_739_Q_reg ( .D(g23110), .SI(g1166), .SE(n8209), .CLK(n8396), .Q(
        g1167) );
  SDFFX1 DFF_740_Q_reg ( .D(g23014), .SI(g1167), .SE(n8210), .CLK(n8397), .Q(
        g1171) );
  SDFFX1 DFF_741_Q_reg ( .D(g23039), .SI(g1171), .SE(n8210), .CLK(n8397), .Q(
        g1151) );
  SDFFX1 DFF_742_Q_reg ( .D(g24212), .SI(g1151), .SE(n8210), .CLK(n8397), .Q(
        g1152) );
  SDFFX1 DFF_743_Q_reg ( .D(g24222), .SI(g1152), .SE(n8210), .CLK(n8397), .Q(
        g1155) );
  SDFFX1 DFF_744_Q_reg ( .D(g24235), .SI(g1155), .SE(n8210), .CLK(n8397), .Q(
        g1158) );
  SDFFX1 DFF_745_Q_reg ( .D(n833), .SI(g1158), .SE(n8210), .CLK(n8397), .Q(
        g1214) );
  SDFFX1 DFF_746_Q_reg ( .D(g1214), .SI(g1214), .SE(n8210), .CLK(n8397), .Q(
        g1221) );
  SDFFX1 DFF_747_Q_reg ( .D(g1221), .SI(g1221), .SE(n8210), .CLK(n8397), .Q(
        test_so45) );
  SDFFX1 DFF_748_Q_reg ( .D(g13155), .SI(test_si46), .SE(n8210), .CLK(n8397), 
        .Q(g1229) );
  SDFFX1 DFF_749_Q_reg ( .D(g1229), .SI(g1229), .SE(n8210), .CLK(n8397), .Q(
        n4549), .QN(n7153) );
  SDFFX1 DFF_750_Q_reg ( .D(n517), .SI(n4549), .SE(n8211), .CLK(n8398), .Q(
        n4361) );
  SDFFX1 DFF_751_Q_reg ( .D(g13124), .SI(n4361), .SE(n8210), .CLK(n8397), .Q(
        g1235) );
  SDFFX1 DFF_752_Q_reg ( .D(g1235), .SI(g1235), .SE(n8210), .CLK(n8397), .Q(
        g1186), .QN(n4548) );
  SDFFX1 DFF_753_Q_reg ( .D(g13171), .SI(g1186), .SE(n8211), .CLK(n8398), .Q(
        g1244) );
  SDFFX1 DFF_754_Q_reg ( .D(g1244), .SI(g1244), .SE(n8211), .CLK(n8398), .Q(
        g1245), .QN(n7763) );
  SDFFX1 DFF_755_Q_reg ( .D(g27273), .SI(g1245), .SE(n8212), .CLK(n8399), .Q(
        g1262), .QN(n7344) );
  SDFFX1 DFF_756_Q_reg ( .D(g27285), .SI(g1262), .SE(n8212), .CLK(n8399), .Q(
        g1263), .QN(n7346) );
  SDFFX1 DFF_757_Q_reg ( .D(g27299), .SI(g1263), .SE(n8212), .CLK(n8399), .Q(
        g1261), .QN(n7345) );
  SDFFX1 DFF_758_Q_reg ( .D(g27286), .SI(g1261), .SE(n8212), .CLK(n8399), .Q(
        g1265), .QN(n7356) );
  SDFFX1 DFF_759_Q_reg ( .D(g27300), .SI(g1265), .SE(n8212), .CLK(n8399), .Q(
        g1266), .QN(n7358) );
  SDFFX1 DFF_760_Q_reg ( .D(g27314), .SI(g1266), .SE(n8212), .CLK(n8399), .Q(
        g1264), .QN(n7357) );
  SDFFX1 DFF_761_Q_reg ( .D(g27301), .SI(g1264), .SE(n8212), .CLK(n8399), .Q(
        g1268), .QN(n7182) );
  SDFFX1 DFF_762_Q_reg ( .D(g27315), .SI(g1268), .SE(n8212), .CLK(n8399), .Q(
        g1269), .QN(n7183) );
  SDFFX1 DFF_763_Q_reg ( .D(g27328), .SI(g1269), .SE(n8212), .CLK(n8399), .Q(
        test_so46), .QN(n8120) );
  SDFFX1 DFF_764_Q_reg ( .D(g27316), .SI(test_si47), .SE(n8212), .CLK(n8399), 
        .Q(g1271), .QN(n7366) );
  SDFFX1 DFF_765_Q_reg ( .D(g27329), .SI(g1271), .SE(n8212), .CLK(n8399), .Q(
        g1272), .QN(n7368) );
  SDFFX1 DFF_766_Q_reg ( .D(g27339), .SI(g1272), .SE(n8212), .CLK(n8399), .Q(
        g1270), .QN(n7367) );
  SDFFX1 DFF_767_Q_reg ( .D(g24501), .SI(g1270), .SE(n8213), .CLK(n8400), .Q(
        g1273) );
  SDFFX1 DFF_768_Q_reg ( .D(g24510), .SI(g1273), .SE(n8213), .CLK(n8400), .Q(
        g1276) );
  SDFFX1 DFF_769_Q_reg ( .D(g24521), .SI(g1276), .SE(n8213), .CLK(n8400), .Q(
        g1279) );
  SDFFX1 DFF_770_Q_reg ( .D(g24511), .SI(g1279), .SE(n8213), .CLK(n8400), .Q(
        g1282) );
  SDFFX1 DFF_771_Q_reg ( .D(g24522), .SI(g1282), .SE(n8213), .CLK(n8400), .Q(
        g1285) );
  SDFFX1 DFF_772_Q_reg ( .D(g24532), .SI(g1285), .SE(n8213), .CLK(n8400), .Q(
        g1288) );
  SDFFX1 DFF_773_Q_reg ( .D(g28351), .SI(g1288), .SE(n8213), .CLK(n8400), .Q(
        g1300) );
  SDFFX1 DFF_774_Q_reg ( .D(g28355), .SI(g1300), .SE(n8213), .CLK(n8400), .Q(
        g1303) );
  SDFFX1 DFF_775_Q_reg ( .D(g28360), .SI(g1303), .SE(n8213), .CLK(n8400), .Q(
        g1306) );
  SDFFX1 DFF_776_Q_reg ( .D(g28346), .SI(g1306), .SE(n8213), .CLK(n8400), .Q(
        g1291) );
  SDFFX1 DFF_777_Q_reg ( .D(g28350), .SI(g1291), .SE(n8214), .CLK(n8401), .Q(
        g1294) );
  SDFFX1 DFF_778_Q_reg ( .D(g28354), .SI(g1294), .SE(n8214), .CLK(n8401), .Q(
        g1297) );
  SDFFX1 DFF_779_Q_reg ( .D(g26547), .SI(g1297), .SE(n8214), .CLK(n8401), .Q(
        test_so47) );
  SDFFX1 DFF_780_Q_reg ( .D(g26557), .SI(test_si48), .SE(n8214), .CLK(n8401), 
        .Q(g1180) );
  SDFFX1 DFF_781_Q_reg ( .D(g26569), .SI(g1180), .SE(n8214), .CLK(n8401), .Q(
        g1183) );
  SDFFX1 DFF_782_Q_reg ( .D(g1186), .SI(g1183), .SE(n8214), .CLK(n8401), .Q(
        g1192), .QN(n4454) );
  SDFFX1 DFF_783_Q_reg ( .D(g22615), .SI(g1192), .SE(n8214), .CLK(n8401), .Q(
        n8009), .QN(DFF_783_n1) );
  SDFFX1 DFF_792_Q_reg ( .D(n532), .SI(n8009), .SE(n8214), .CLK(n8401), .Q(
        g16355), .QN(DFF_792_n1) );
  SDFFX1 DFF_793_Q_reg ( .D(g16355), .SI(g16355), .SE(n8214), .CLK(n8401), .Q(
        g1211), .QN(n8063) );
  SDFFX1 DFF_794_Q_reg ( .D(DFF_649_n1), .SI(g1211), .SE(n8214), .CLK(n8401), 
        .Q(n8008), .QN(DFF_794_n1) );
  SDFFX1 DFF_795_Q_reg ( .D(DFF_651_n1), .SI(n8008), .SE(n8214), .CLK(n8401), 
        .Q(n8007), .QN(DFF_795_n1) );
  SDFFX1 DFF_796_Q_reg ( .D(DFF_653_n1), .SI(n8007), .SE(n8215), .CLK(n8402), 
        .Q(n8006), .QN(DFF_796_n1) );
  SDFFX1 DFF_797_Q_reg ( .D(DFF_655_n1), .SI(n8006), .SE(n8215), .CLK(n8402), 
        .Q(n8005), .QN(DFF_797_n1) );
  SDFFX1 DFF_798_Q_reg ( .D(DFF_657_n1), .SI(n8005), .SE(n8215), .CLK(n8402), 
        .Q(n8004), .QN(DFF_798_n1) );
  SDFFX1 DFF_799_Q_reg ( .D(DFF_659_n1), .SI(n8004), .SE(n8215), .CLK(n8402), 
        .Q(n8003), .QN(DFF_799_n1) );
  SDFFX1 DFF_800_Q_reg ( .D(DFF_661_n1), .SI(n8003), .SE(n8215), .CLK(n8402), 
        .Q(g1222), .QN(n7161) );
  SDFFX1 DFF_801_Q_reg ( .D(DFF_663_n1), .SI(g1222), .SE(n8215), .CLK(n8402), 
        .Q(g1223), .QN(n7160) );
  SDFFX1 DFF_802_Q_reg ( .D(g24072), .SI(g1223), .SE(n8215), .CLK(n8402), .Q(
        g1224), .QN(n4489) );
  SDFFX1 DFF_803_Q_reg ( .D(n4486), .SI(g1224), .SE(n8215), .CLK(n8402), .Q(
        test_so48), .QN(n14381) );
  SDFFX1 DFF_805_Q_reg ( .D(g6979), .SI(g6979), .SE(n8172), .CLK(n8359), .Q(
        g7161), .QN(n4358) );
  SDFFX1 DFF_806_Q_reg ( .D(g7161), .SI(g7161), .SE(n8172), .CLK(n8359), .Q(
        g1315), .QN(n4294) );
  SDFFX1 DFF_807_Q_reg ( .D(g16671), .SI(g1315), .SE(n8206), .CLK(n8393), .Q(
        g1316), .QN(n7759) );
  SDFFX1 DFF_808_Q_reg ( .D(g20333), .SI(g1316), .SE(n8206), .CLK(n8393), .Q(
        g1345), .QN(n4428) );
  SDFFX1 DFF_809_Q_reg ( .D(g20717), .SI(g1345), .SE(n8206), .CLK(n8393), .Q(
        g1326), .QN(n4402) );
  SDFFX1 DFF_810_Q_reg ( .D(n912), .SI(g1326), .SE(n8206), .CLK(n8393), .Q(
        g1319), .QN(n4476) );
  SDFFX1 DFF_811_Q_reg ( .D(g23329), .SI(g1319), .SE(n8207), .CLK(n8394), .Q(
        g1339), .QN(n4421) );
  SDFFX1 DFF_812_Q_reg ( .D(g24430), .SI(g1339), .SE(n8207), .CLK(n8394), .Q(
        g1332), .QN(n4412) );
  SDFFX1 DFF_813_Q_reg ( .D(g25189), .SI(g1332), .SE(n8207), .CLK(n8394), .Q(
        g1346), .QN(n4401) );
  SDFFX1 DFF_814_Q_reg ( .D(n913), .SI(g1346), .SE(n8207), .CLK(n8394), .Q(
        g1358), .QN(n4411) );
  SDFFX1 DFF_815_Q_reg ( .D(g26781), .SI(g1358), .SE(n8207), .CLK(n8394), .Q(
        g1352), .QN(n4469) );
  SDFFX1 DFF_816_Q_reg ( .D(g27678), .SI(g1352), .SE(n8207), .CLK(n8394), .Q(
        g1365), .QN(n4475) );
  SDFFX1 DFF_817_Q_reg ( .D(g27718), .SI(g1365), .SE(n8207), .CLK(n8394), .Q(
        g1372), .QN(n4395) );
  SDFFX1 DFF_818_Q_reg ( .D(g28321), .SI(g1372), .SE(n8207), .CLK(n8394), .Q(
        g1378), .QN(n4417) );
  SDFFX1 DFF_819_Q_reg ( .D(g20882), .SI(g1378), .SE(n8215), .CLK(n8402), .Q(
        test_so49), .QN(n8136) );
  SDFFX1 DFF_820_Q_reg ( .D(g20896), .SI(test_si50), .SE(n8215), .CLK(n8402), 
        .Q(g1386), .QN(n7820) );
  SDFFX1 DFF_821_Q_reg ( .D(g20910), .SI(g1386), .SE(n8215), .CLK(n8402), .Q(
        g1384), .QN(n7866) );
  SDFFX1 DFF_822_Q_reg ( .D(g20897), .SI(g1384), .SE(n8215), .CLK(n8402), .Q(
        g1388), .QN(n7819) );
  SDFFX1 DFF_823_Q_reg ( .D(g20911), .SI(g1388), .SE(n8216), .CLK(n8403), .Q(
        g1389), .QN(n7818) );
  SDFFX1 DFF_824_Q_reg ( .D(g20925), .SI(g1389), .SE(n8216), .CLK(n8403), .Q(
        g1387), .QN(n7865) );
  SDFFX1 DFF_825_Q_reg ( .D(g20912), .SI(g1387), .SE(n8216), .CLK(n8403), .Q(
        g1391), .QN(n7817) );
  SDFFX1 DFF_826_Q_reg ( .D(g20926), .SI(g1391), .SE(n8216), .CLK(n8403), .Q(
        g1392), .QN(n7816) );
  SDFFX1 DFF_827_Q_reg ( .D(g20949), .SI(g1392), .SE(n8216), .CLK(n8403), .Q(
        g1390), .QN(n7864) );
  SDFFX1 DFF_828_Q_reg ( .D(g20927), .SI(g1390), .SE(n8216), .CLK(n8403), .Q(
        g1394), .QN(n7815) );
  SDFFX1 DFF_829_Q_reg ( .D(g20950), .SI(g1394), .SE(n8216), .CLK(n8403), .Q(
        g1395), .QN(n7814) );
  SDFFX1 DFF_830_Q_reg ( .D(g20972), .SI(g1395), .SE(n8216), .CLK(n8403), .Q(
        g1393), .QN(n7863) );
  SDFFX1 DFF_831_Q_reg ( .D(g20951), .SI(g1393), .SE(n8216), .CLK(n8403), .Q(
        g1397), .QN(n7813) );
  SDFFX1 DFF_832_Q_reg ( .D(g20973), .SI(g1397), .SE(n8216), .CLK(n8403), .Q(
        g1398), .QN(n7812) );
  SDFFX1 DFF_833_Q_reg ( .D(g20993), .SI(g1398), .SE(n8216), .CLK(n8403), .Q(
        g1396), .QN(n7862) );
  SDFFX1 DFF_834_Q_reg ( .D(g20974), .SI(g1396), .SE(n8216), .CLK(n8403), .Q(
        g1400), .QN(n7811) );
  SDFFX1 DFF_835_Q_reg ( .D(g20994), .SI(g1400), .SE(n8217), .CLK(n8404), .Q(
        test_so50), .QN(n8135) );
  SDFFX1 DFF_836_Q_reg ( .D(g21015), .SI(test_si51), .SE(n8217), .CLK(n8404), 
        .Q(g1399), .QN(n7861) );
  SDFFX1 DFF_837_Q_reg ( .D(g20995), .SI(g1399), .SE(n8217), .CLK(n8404), .Q(
        g1403), .QN(n7810) );
  SDFFX1 DFF_838_Q_reg ( .D(g21016), .SI(g1403), .SE(n8217), .CLK(n8404), .Q(
        g1404), .QN(n7809) );
  SDFFX1 DFF_839_Q_reg ( .D(g21033), .SI(g1404), .SE(n8217), .CLK(n8404), .Q(
        g1402), .QN(n7860) );
  SDFFX1 DFF_840_Q_reg ( .D(g21017), .SI(g1402), .SE(n8217), .CLK(n8404), .Q(
        g1406), .QN(n7808) );
  SDFFX1 DFF_841_Q_reg ( .D(g21034), .SI(g1406), .SE(n8217), .CLK(n8404), .Q(
        g1407), .QN(n7807) );
  SDFFX1 DFF_842_Q_reg ( .D(g21052), .SI(g1407), .SE(n8217), .CLK(n8404), .Q(
        g1405), .QN(n7859) );
  SDFFX1 DFF_843_Q_reg ( .D(g21035), .SI(g1405), .SE(n8217), .CLK(n8404), .Q(
        g1409), .QN(n7806) );
  SDFFX1 DFF_844_Q_reg ( .D(g21053), .SI(g1409), .SE(n8217), .CLK(n8404), .Q(
        g1410), .QN(n7805) );
  SDFFX1 DFF_845_Q_reg ( .D(g21070), .SI(g1410), .SE(n8217), .CLK(n8404), .Q(
        g1408), .QN(n7858) );
  SDFFX1 DFF_846_Q_reg ( .D(g20883), .SI(g1408), .SE(n8217), .CLK(n8404), .Q(
        g1412), .QN(n7804) );
  SDFFX1 DFF_847_Q_reg ( .D(g20898), .SI(g1412), .SE(n8218), .CLK(n8405), .Q(
        g1413), .QN(n7803) );
  SDFFX1 DFF_848_Q_reg ( .D(g20913), .SI(g1413), .SE(n8218), .CLK(n8405), .Q(
        g1411), .QN(n7857) );
  SDFFX1 DFF_849_Q_reg ( .D(g20952), .SI(g1411), .SE(n8218), .CLK(n8405), .Q(
        g1415), .QN(n8039) );
  SDFFX1 DFF_850_Q_reg ( .D(g20975), .SI(g1415), .SE(n8218), .CLK(n8405), .Q(
        g1416), .QN(n7572) );
  SDFFX1 DFF_851_Q_reg ( .D(g20996), .SI(g1416), .SE(n8218), .CLK(n8405), .Q(
        test_so51) );
  SDFFX1 DFF_852_Q_reg ( .D(g20976), .SI(test_si52), .SE(n8213), .CLK(n8400), 
        .Q(g1418), .QN(n7577) );
  SDFFX1 DFF_853_Q_reg ( .D(g20997), .SI(g1418), .SE(n8213), .CLK(n8400), .Q(
        g1419), .QN(n7571) );
  SDFFX1 DFF_854_Q_reg ( .D(g21018), .SI(g1419), .SE(n8214), .CLK(n8401), .Q(
        g1417), .QN(n7629) );
  SDFFX1 DFF_855_Q_reg ( .D(g25263), .SI(g1417), .SE(n8218), .CLK(n8405), .Q(
        g1421), .QN(n7507) );
  SDFFX1 DFF_856_Q_reg ( .D(g25267), .SI(g1421), .SE(n8218), .CLK(n8405), .Q(
        g1422), .QN(n7506) );
  SDFFX1 DFF_857_Q_reg ( .D(g25270), .SI(g1422), .SE(n8218), .CLK(n8405), .Q(
        g1420), .QN(n7512) );
  SDFFX1 DFF_858_Q_reg ( .D(g22234), .SI(g1420), .SE(n8218), .CLK(n8405), .Q(
        g1424), .QN(n7879) );
  SDFFX1 DFF_859_Q_reg ( .D(n883), .SI(g1424), .SE(n8218), .CLK(n8405), .Q(
        g1425), .QN(n7976) );
  SDFFX1 DFF_860_Q_reg ( .D(g22263), .SI(g1425), .SE(n8218), .CLK(n8405), .Q(
        g1423), .QN(n7982) );
  SDFFX1 DFF_861_Q_reg ( .D(g2950), .SI(g1423), .SE(n8218), .CLK(n8405), .Q(
        g6573), .QN(n4317) );
  SDFFX1 DFF_862_Q_reg ( .D(g6573), .SI(g6573), .SE(n8219), .CLK(n8406), .Q(
        g6782), .QN(n4515) );
  SDFFX1 DFF_863_Q_reg ( .D(g6782), .SI(g6782), .SE(n8219), .CLK(n8406), .Q(
        g1547), .QN(n4368) );
  SDFFX1 DFF_864_Q_reg ( .D(g22149), .SI(g1547), .SE(n8219), .CLK(n8406), .Q(
        g1512), .QN(n7911) );
  SDFFX1 DFF_865_Q_reg ( .D(g22166), .SI(g1512), .SE(n8223), .CLK(n8410), .Q(
        g1513), .QN(n7910) );
  SDFFX1 DFF_866_Q_reg ( .D(g22178), .SI(g1513), .SE(n8223), .CLK(n8410), .Q(
        g1511), .QN(n7543) );
  SDFFX1 DFF_867_Q_reg ( .D(g22167), .SI(g1511), .SE(n8219), .CLK(n8406), .Q(
        test_so52), .QN(n8110) );
  SDFFX1 DFF_868_Q_reg ( .D(g22179), .SI(test_si53), .SE(n8223), .CLK(n8410), 
        .Q(g1516), .QN(n7908) );
  SDFFX1 DFF_869_Q_reg ( .D(g22191), .SI(g1516), .SE(n8224), .CLK(n8411), .Q(
        g1514), .QN(n7542) );
  SDFFX1 DFF_870_Q_reg ( .D(g22035), .SI(g1514), .SE(n8224), .CLK(n8411), .Q(
        g1524), .QN(n7906) );
  SDFFX1 DFF_871_Q_reg ( .D(g22043), .SI(g1524), .SE(n8224), .CLK(n8411), .Q(
        g1525), .QN(n7905) );
  SDFFX1 DFF_872_Q_reg ( .D(g22057), .SI(g1525), .SE(n8224), .CLK(n8411), .Q(
        g1523), .QN(n7541) );
  SDFFX1 DFF_873_Q_reg ( .D(g22044), .SI(g1523), .SE(n8224), .CLK(n8411), .Q(
        g1527), .QN(n7904) );
  SDFFX1 DFF_874_Q_reg ( .D(g22058), .SI(g1527), .SE(n8224), .CLK(n8411), .Q(
        g1528), .QN(n7903) );
  SDFFX1 DFF_875_Q_reg ( .D(g22073), .SI(g1528), .SE(n8224), .CLK(n8411), .Q(
        g1526), .QN(n7540) );
  SDFFX1 DFF_876_Q_reg ( .D(g22059), .SI(g1526), .SE(n8224), .CLK(n8411), .Q(
        g1530), .QN(n7902) );
  SDFFX1 DFF_877_Q_reg ( .D(g22074), .SI(g1530), .SE(n8224), .CLK(n8411), .Q(
        g1531), .QN(n7901) );
  SDFFX1 DFF_878_Q_reg ( .D(g22090), .SI(g1531), .SE(n8224), .CLK(n8411), .Q(
        g1529), .QN(n7539) );
  SDFFX1 DFF_879_Q_reg ( .D(g22075), .SI(g1529), .SE(n8224), .CLK(n8411), .Q(
        g1533), .QN(n7900) );
  SDFFX1 DFF_880_Q_reg ( .D(g22091), .SI(g1533), .SE(n8224), .CLK(n8411), .Q(
        g1534), .QN(n7899) );
  SDFFX1 DFF_881_Q_reg ( .D(g22112), .SI(g1534), .SE(n8225), .CLK(n8412), .Q(
        g1532), .QN(n7538) );
  SDFFX1 DFF_882_Q_reg ( .D(g22092), .SI(g1532), .SE(n8225), .CLK(n8412), .Q(
        g1536), .QN(n7898) );
  SDFFX1 DFF_883_Q_reg ( .D(g22113), .SI(g1536), .SE(n8225), .CLK(n8412), .Q(
        test_so53), .QN(n8124) );
  SDFFX1 DFF_884_Q_reg ( .D(g22130), .SI(test_si54), .SE(n8222), .CLK(n8409), 
        .Q(g1535), .QN(n7537) );
  SDFFX1 DFF_885_Q_reg ( .D(g22114), .SI(g1535), .SE(n8222), .CLK(n8409), .Q(
        g1539), .QN(n7897) );
  SDFFX1 DFF_886_Q_reg ( .D(g22131), .SI(g1539), .SE(n8222), .CLK(n8409), .Q(
        g1540), .QN(n7896) );
  SDFFX1 DFF_887_Q_reg ( .D(g22150), .SI(g1540), .SE(n8222), .CLK(n8409), .Q(
        g1538), .QN(n7536) );
  SDFFX1 DFF_888_Q_reg ( .D(g22132), .SI(g1538), .SE(n8222), .CLK(n8409), .Q(
        g1542), .QN(n7519) );
  SDFFX1 DFF_889_Q_reg ( .D(g22151), .SI(g1542), .SE(n8222), .CLK(n8409), .Q(
        g1543), .QN(n7518) );
  SDFFX1 DFF_890_Q_reg ( .D(g22168), .SI(g1543), .SE(n8222), .CLK(n8409), .Q(
        g1541), .QN(n7517) );
  SDFFX1 DFF_891_Q_reg ( .D(g22152), .SI(g1541), .SE(n8223), .CLK(n8410), .Q(
        g1545), .QN(n7535) );
  SDFFX1 DFF_892_Q_reg ( .D(g22169), .SI(g1545), .SE(n8223), .CLK(n8410), .Q(
        g1546), .QN(n7534) );
  SDFFX1 DFF_893_Q_reg ( .D(g22180), .SI(g1546), .SE(n8223), .CLK(n8410), .Q(
        g1544), .QN(n7533) );
  SDFFX1 DFF_894_Q_reg ( .D(g25217), .SI(g1544), .SE(n8223), .CLK(n8410), .Q(
        g1551), .QN(n7601) );
  SDFFX1 DFF_895_Q_reg ( .D(g25224), .SI(g1551), .SE(n8223), .CLK(n8410), .Q(
        g1552), .QN(n7600) );
  SDFFX1 DFF_896_Q_reg ( .D(g25233), .SI(g1552), .SE(n8223), .CLK(n8410), .Q(
        g1550), .QN(n7599) );
  SDFFX1 DFF_897_Q_reg ( .D(g25225), .SI(g1550), .SE(n8223), .CLK(n8410), .Q(
        g1554), .QN(n7598) );
  SDFFX1 DFF_898_Q_reg ( .D(g25234), .SI(g1554), .SE(n8223), .CLK(n8410), .Q(
        g1555), .QN(n7597) );
  SDFFX1 DFF_899_Q_reg ( .D(g25242), .SI(g1555), .SE(n8223), .CLK(n8410), .Q(
        test_so54), .QN(n8141) );
  SDFFX1 DFF_900_Q_reg ( .D(g25235), .SI(test_si55), .SE(n8219), .CLK(n8406), 
        .Q(g1557), .QN(n7596) );
  SDFFX1 DFF_901_Q_reg ( .D(g25243), .SI(g1557), .SE(n8219), .CLK(n8406), .Q(
        g1558), .QN(n7595) );
  SDFFX1 DFF_902_Q_reg ( .D(g25249), .SI(g1558), .SE(n8219), .CLK(n8406), .Q(
        g1556), .QN(n7594) );
  SDFFX1 DFF_903_Q_reg ( .D(g25244), .SI(g1556), .SE(n8219), .CLK(n8406), .Q(
        g1560), .QN(n7593) );
  SDFFX1 DFF_904_Q_reg ( .D(g25250), .SI(g1560), .SE(n8219), .CLK(n8406), .Q(
        g1561), .QN(n7592) );
  SDFFX1 DFF_905_Q_reg ( .D(g25255), .SI(g1561), .SE(n8219), .CLK(n8406), .Q(
        g1559), .QN(n7591) );
  SDFFX1 DFF_906_Q_reg ( .D(g30279), .SI(g1559), .SE(n8226), .CLK(n8413), .Q(
        g1567) );
  SDFFX1 DFF_907_Q_reg ( .D(g30287), .SI(g1567), .SE(n8226), .CLK(n8413), .Q(
        g1570) );
  SDFFX1 DFF_908_Q_reg ( .D(g30294), .SI(g1570), .SE(n8226), .CLK(n8413), .Q(
        g1573) );
  SDFFX1 DFF_909_Q_reg ( .D(g30651), .SI(g1573), .SE(n8226), .CLK(n8413), .Q(
        g1612) );
  SDFFX1 DFF_910_Q_reg ( .D(g30657), .SI(g1612), .SE(n8226), .CLK(n8413), .Q(
        g1615) );
  SDFFX1 DFF_911_Q_reg ( .D(g30663), .SI(g1615), .SE(n8225), .CLK(n8412), .Q(
        g1618) );
  SDFFX1 DFF_912_Q_reg ( .D(g30683), .SI(g1618), .SE(n8226), .CLK(n8413), .Q(
        g1576) );
  SDFFX1 DFF_913_Q_reg ( .D(g30688), .SI(g1576), .SE(n8226), .CLK(n8413), .Q(
        g1579) );
  SDFFX1 DFF_914_Q_reg ( .D(g30692), .SI(g1579), .SE(n8219), .CLK(n8406), .Q(
        g1582) );
  SDFFX1 DFF_915_Q_reg ( .D(g30658), .SI(g1582), .SE(n8219), .CLK(n8406), .Q(
        test_so55) );
  SDFFX1 DFF_916_Q_reg ( .D(g30664), .SI(test_si56), .SE(n8220), .CLK(n8407), 
        .Q(g1624) );
  SDFFX1 DFF_917_Q_reg ( .D(g30671), .SI(g1624), .SE(n8220), .CLK(n8407), .Q(
        g1627) );
  SDFFX1 DFF_918_Q_reg ( .D(g30295), .SI(g1627), .SE(n8220), .CLK(n8407), .Q(
        g1585) );
  SDFFX1 DFF_919_Q_reg ( .D(g30299), .SI(g1585), .SE(n8220), .CLK(n8407), .Q(
        g1588) );
  SDFFX1 DFF_920_Q_reg ( .D(g30302), .SI(g1588), .SE(n8220), .CLK(n8407), .Q(
        g1591) );
  SDFFX1 DFF_921_Q_reg ( .D(g30266), .SI(g1591), .SE(n8220), .CLK(n8407), .Q(
        g1630) );
  SDFFX1 DFF_922_Q_reg ( .D(g30272), .SI(g1630), .SE(n8220), .CLK(n8407), .Q(
        g1633) );
  SDFFX1 DFF_923_Q_reg ( .D(g30280), .SI(g1633), .SE(n8220), .CLK(n8407), .Q(
        g1636) );
  SDFFX1 DFF_924_Q_reg ( .D(g30250), .SI(g1636), .SE(n8225), .CLK(n8412), .Q(
        g1594) );
  SDFFX1 DFF_925_Q_reg ( .D(g30252), .SI(g1594), .SE(n8225), .CLK(n8412), .Q(
        g1597) );
  SDFFX1 DFF_926_Q_reg ( .D(g30255), .SI(g1597), .SE(n8225), .CLK(n8412), .Q(
        g1600) );
  SDFFX1 DFF_927_Q_reg ( .D(g30273), .SI(g1600), .SE(n8225), .CLK(n8412), .Q(
        g1639) );
  SDFFX1 DFF_928_Q_reg ( .D(g30281), .SI(g1639), .SE(n8225), .CLK(n8412), .Q(
        g1642) );
  SDFFX1 DFF_929_Q_reg ( .D(g30288), .SI(g1642), .SE(n8225), .CLK(n8412), .Q(
        g1645) );
  SDFFX1 DFF_930_Q_reg ( .D(g30644), .SI(g1645), .SE(n8225), .CLK(n8412), .Q(
        g1603) );
  SDFFX1 DFF_931_Q_reg ( .D(g30650), .SI(g1603), .SE(n8225), .CLK(n8412), .Q(
        test_so56) );
  SDFFX1 DFF_932_Q_reg ( .D(g30656), .SI(test_si57), .SE(n8220), .CLK(n8407), 
        .Q(g1609) );
  SDFFX1 DFF_933_Q_reg ( .D(g30678), .SI(g1609), .SE(n8220), .CLK(n8407), .Q(
        g1648) );
  SDFFX1 DFF_934_Q_reg ( .D(g30684), .SI(g1648), .SE(n8220), .CLK(n8407), .Q(
        g1651) );
  SDFFX1 DFF_935_Q_reg ( .D(g30689), .SI(g1651), .SE(n8220), .CLK(n8407), .Q(
        g1654) );
  SDFFX1 DFF_936_Q_reg ( .D(g25056), .SI(g1654), .SE(n8221), .CLK(n8408), .Q(
        g1466), .QN(n7706) );
  SDFFX1 DFF_937_Q_reg ( .D(g25938), .SI(g1466), .SE(n8221), .CLK(n8408), .Q(
        g1462), .QN(n8069) );
  SDFFX1 DFF_938_Q_reg ( .D(g26531), .SI(g1462), .SE(n8221), .CLK(n8408), .Q(
        g1457), .QN(n7705) );
  SDFFX1 DFF_939_Q_reg ( .D(g27129), .SI(g1457), .SE(n8221), .CLK(n8408), .Q(
        g1453) );
  SDFFX1 DFF_940_Q_reg ( .D(g27612), .SI(g1453), .SE(n8221), .CLK(n8408), .Q(
        g1448), .QN(n7704) );
  SDFFX1 DFF_941_Q_reg ( .D(g28147), .SI(g1448), .SE(n8221), .CLK(n8408), .Q(
        g1444), .QN(n8094) );
  SDFFX1 DFF_942_Q_reg ( .D(g28636), .SI(g1444), .SE(n8221), .CLK(n8408), .Q(
        g1439), .QN(n7703) );
  SDFFX1 DFF_943_Q_reg ( .D(g29111), .SI(g1439), .SE(n8221), .CLK(n8408), .Q(
        g1435), .QN(n8071) );
  SDFFX1 DFF_944_Q_reg ( .D(g29355), .SI(g1435), .SE(n8221), .CLK(n8408), .Q(
        g1430), .QN(n7335) );
  SDFFX1 DFF_945_Q_reg ( .D(g29581), .SI(g1430), .SE(n8221), .CLK(n8408), .Q(
        g1426), .QN(n7174) );
  SDFFX1 DFF_946_Q_reg ( .D(n15), .SI(g1426), .SE(n8221), .CLK(n8408), .Q(
        g1562) );
  SDFFX1 DFF_947_Q_reg ( .D(g1562), .SI(g1562), .SE(n8221), .CLK(n8408), .Q(
        test_so57) );
  SDFFX1 DFF_948_Q_reg ( .D(test_so57), .SI(test_si58), .SE(n8222), .CLK(n8409), .Q(g1563), .QN(n7719) );
  SDFFX1 DFF_949_Q_reg ( .D(g2950), .SI(g1563), .SE(n8222), .CLK(n8409), .Q(
        g5511), .QN(n4518) );
  SDFFX1 DFF_952_Q_reg ( .D(test_so57), .SI(n4618), .SE(n8222), .CLK(n8409), 
        .Q(g1690), .QN(n4386) );
  SDFFX1 DFF_953_Q_reg ( .D(g27264), .SI(g1690), .SE(n8230), .CLK(n8417), .Q(
        g1735), .QN(n7660) );
  SDFFX1 DFF_954_Q_reg ( .D(g27274), .SI(g1735), .SE(n8230), .CLK(n8417), .Q(
        g1724), .QN(n7659) );
  SDFFX1 DFF_955_Q_reg ( .D(g27287), .SI(g1724), .SE(n8230), .CLK(n8417), .Q(
        g1727), .QN(n7658) );
  SDFFX1 DFF_956_Q_reg ( .D(g27275), .SI(g1727), .SE(n8231), .CLK(n8418), .Q(
        g1750), .QN(n7637) );
  SDFFX1 DFF_957_Q_reg ( .D(g27288), .SI(g1750), .SE(n8231), .CLK(n8418), .Q(
        g1739), .QN(n7636) );
  SDFFX1 DFF_958_Q_reg ( .D(g27302), .SI(g1739), .SE(n8231), .CLK(n8418), .Q(
        g1742), .QN(n7635) );
  SDFFX1 DFF_959_Q_reg ( .D(g27289), .SI(g1742), .SE(n8231), .CLK(n8418), .Q(
        g1765), .QN(n7386) );
  SDFFX1 DFF_960_Q_reg ( .D(g27303), .SI(g1765), .SE(n8231), .CLK(n8418), .Q(
        g1754), .QN(n7388) );
  SDFFX1 DFF_961_Q_reg ( .D(g27317), .SI(g1754), .SE(n8230), .CLK(n8417), .Q(
        g1757), .QN(n7387) );
  SDFFX1 DFF_962_Q_reg ( .D(g27304), .SI(g1757), .SE(n8231), .CLK(n8418), .Q(
        g1779), .QN(n7648) );
  SDFFX1 DFF_963_Q_reg ( .D(g27318), .SI(g1779), .SE(n8231), .CLK(n8418), .Q(
        test_so58), .QN(n8113) );
  SDFFX1 DFF_964_Q_reg ( .D(g27330), .SI(test_si59), .SE(n8228), .CLK(n8415), 
        .Q(g1772), .QN(n7647) );
  SDFFX1 DFF_965_Q_reg ( .D(g28749), .SI(g1772), .SE(n8228), .CLK(n8415), .Q(
        g1789) );
  SDFFX1 DFF_966_Q_reg ( .D(g28760), .SI(g1789), .SE(n8230), .CLK(n8417), .Q(
        g1792) );
  SDFFX1 DFF_967_Q_reg ( .D(g28771), .SI(g1792), .SE(n8230), .CLK(n8417), .Q(
        g1795) );
  SDFFX1 DFF_968_Q_reg ( .D(g29205), .SI(g1795), .SE(n8230), .CLK(n8417), .Q(
        g1798) );
  SDFFX1 DFF_969_Q_reg ( .D(g29212), .SI(g1798), .SE(n8230), .CLK(n8417), .Q(
        g1801) );
  SDFFX1 DFF_970_Q_reg ( .D(g29218), .SI(g1801), .SE(n8229), .CLK(n8416), .Q(
        g1804) );
  SDFFX1 DFF_971_Q_reg ( .D(g28761), .SI(g1804), .SE(n8229), .CLK(n8416), .Q(
        g1808), .QN(n7683) );
  SDFFX1 DFF_972_Q_reg ( .D(g28772), .SI(g1808), .SE(n8229), .CLK(n8416), .Q(
        g1809), .QN(n7671) );
  SDFFX1 DFF_973_Q_reg ( .D(g28778), .SI(g1809), .SE(n8229), .CLK(n8416), .Q(
        g1807), .QN(n7682) );
  SDFFX1 DFF_974_Q_reg ( .D(g26811), .SI(g1807), .SE(n8229), .CLK(n8416), .Q(
        g1810) );
  SDFFX1 DFF_975_Q_reg ( .D(g26815), .SI(g1810), .SE(n8229), .CLK(n8416), .Q(
        g1813) );
  SDFFX1 DFF_976_Q_reg ( .D(g26820), .SI(g1813), .SE(n8229), .CLK(n8416), .Q(
        g1816) );
  SDFFX1 DFF_977_Q_reg ( .D(g26816), .SI(g1816), .SE(n8229), .CLK(n8416), .Q(
        g1819) );
  SDFFX1 DFF_978_Q_reg ( .D(g26821), .SI(g1819), .SE(n8229), .CLK(n8416), .Q(
        g1822) );
  SDFFX1 DFF_979_Q_reg ( .D(g26824), .SI(g1822), .SE(n8230), .CLK(n8417), .Q(
        test_so59) );
  SDFFX1 DFF_980_Q_reg ( .D(g27764), .SI(test_si60), .SE(n8230), .CLK(n8417), 
        .Q(g1829), .QN(n7681) );
  SDFFX1 DFF_981_Q_reg ( .D(g27766), .SI(g1829), .SE(n8230), .CLK(n8417), .Q(
        g1830), .QN(n7670) );
  SDFFX1 DFF_982_Q_reg ( .D(g27768), .SI(g1830), .SE(n8229), .CLK(n8416), .Q(
        g1828), .QN(n7680) );
  SDFFX1 DFF_983_Q_reg ( .D(g29613), .SI(g1828), .SE(n8229), .CLK(n8416), .Q(
        g1693), .QN(n7288) );
  SDFFX1 DFF_984_Q_reg ( .D(g29617), .SI(g1693), .SE(n8229), .CLK(n8416), .Q(
        g1694), .QN(n7273) );
  SDFFX1 DFF_985_Q_reg ( .D(g29620), .SI(g1694), .SE(n8226), .CLK(n8413), .Q(
        g1695), .QN(n7287) );
  SDFFX1 DFF_986_Q_reg ( .D(g30704), .SI(g1695), .SE(n8227), .CLK(n8414), .Q(
        g1696), .QN(n7286) );
  SDFFX1 DFF_987_Q_reg ( .D(g30706), .SI(g1696), .SE(n8227), .CLK(n8414), .Q(
        g1697), .QN(n7272) );
  SDFFX1 DFF_988_Q_reg ( .D(g30708), .SI(g1697), .SE(n8226), .CLK(n8413), .Q(
        g1698), .QN(n7285) );
  SDFFX1 DFF_989_Q_reg ( .D(g30487), .SI(g1698), .SE(n8226), .CLK(n8413), .Q(
        g1699), .QN(n7284) );
  SDFFX1 DFF_990_Q_reg ( .D(g30503), .SI(g1699), .SE(n8226), .CLK(n8413), .Q(
        g1700), .QN(n7271) );
  SDFFX1 DFF_991_Q_reg ( .D(g30338), .SI(g1700), .SE(n8226), .CLK(n8413), .Q(
        g1701), .QN(n7283) );
  SDFFX1 DFF_992_Q_reg ( .D(g29178), .SI(g1701), .SE(n8227), .CLK(n8414), .Q(
        g1703), .QN(n7328) );
  SDFFX1 DFF_993_Q_reg ( .D(g29181), .SI(g1703), .SE(n8227), .CLK(n8414), .Q(
        g1704), .QN(n7323) );
  SDFFX1 DFF_994_Q_reg ( .D(g29184), .SI(g1704), .SE(n8227), .CLK(n8414), .Q(
        g1702), .QN(n7327) );
  SDFFX1 DFF_995_Q_reg ( .D(g26667), .SI(g1702), .SE(n8227), .CLK(n8414), .Q(
        test_so60), .QN(n8123) );
  SDFFX1 DFF_996_Q_reg ( .D(g26670), .SI(test_si61), .SE(n8227), .CLK(n8414), 
        .Q(g1785), .QN(n7669) );
  SDFFX1 DFF_997_Q_reg ( .D(g26675), .SI(g1785), .SE(n8227), .CLK(n8414), .Q(
        g1783), .QN(n7679) );
  SDFFX1 DFF_998_Q_reg ( .D(n4288), .SI(g1783), .SE(n8227), .CLK(n8414), .Q(
        g1831) );
  SDFFX1 DFF_999_Q_reg ( .D(g1831), .SI(g1831), .SE(n8227), .CLK(n8414), .Q(
        n7988), .QN(DFF_999_n1) );
  SDFFX1 DFF_1000_Q_reg ( .D(n4565), .SI(n7988), .SE(n8227), .CLK(n8414), .Q(
        g1833) );
  SDFFX1 DFF_1001_Q_reg ( .D(g1833), .SI(g1833), .SE(n8227), .CLK(n8414), .Q(
        n7987), .QN(DFF_1001_n1) );
  SDFFX1 DFF_1002_Q_reg ( .D(n4557), .SI(n7987), .SE(n8228), .CLK(n8415), .Q(
        g1835) );
  SDFFX1 DFF_1003_Q_reg ( .D(g1835), .SI(g1835), .SE(n8228), .CLK(n8415), .Q(
        n7986), .QN(DFF_1003_n1) );
  SDFFX1 DFF_1004_Q_reg ( .D(n4326), .SI(n7986), .SE(n8228), .CLK(n8415), .Q(
        g1661) );
  SDFFX1 DFF_1005_Q_reg ( .D(g1661), .SI(g1661), .SE(n8228), .CLK(n8415), .Q(
        n7985), .QN(DFF_1005_n1) );
  SDFFX1 DFF_1006_Q_reg ( .D(n4390), .SI(n7985), .SE(n8228), .CLK(n8415), .Q(
        g1663) );
  SDFFX1 DFF_1007_Q_reg ( .D(g1663), .SI(g1663), .SE(n8228), .CLK(n8415), .Q(
        n7984), .QN(DFF_1007_n1) );
  SDFFX1 DFF_1008_Q_reg ( .D(n4320), .SI(n7984), .SE(n8228), .CLK(n8415), .Q(
        g1665) );
  SDFFX1 DFF_1009_Q_reg ( .D(g1665), .SI(g1665), .SE(n8228), .CLK(n8415), .Q(
        n7983), .QN(DFF_1009_n1) );
  SDFFX1 DFF_1010_Q_reg ( .D(n4374), .SI(n7983), .SE(n8228), .CLK(n8415), .Q(
        g1667) );
  SDFFX1 DFF_1011_Q_reg ( .D(g1667), .SI(g1667), .SE(n8228), .CLK(n8415), .Q(
        test_so61), .QN(DFF_1011_n1) );
  SDFFX1 DFF_1012_Q_reg ( .D(n4378), .SI(test_si62), .SE(n8144), .CLK(n8331), 
        .Q(g1669) );
  SDFFX1 DFF_1013_Q_reg ( .D(g1669), .SI(g1669), .SE(n8144), .CLK(n8331), .Q(
        n7980), .QN(DFF_1013_n1) );
  SDFFX1 DFF_1014_Q_reg ( .D(g2877), .SI(n7980), .SE(n8149), .CLK(n8336), .Q(
        g1671) );
  SDFFX1 DFF_1015_Q_reg ( .D(g1671), .SI(g1671), .SE(n8149), .CLK(n8336), .Q(
        n7979), .QN(n4484) );
  SDFFX1 DFF_1016_Q_reg ( .D(n4284), .SI(n7979), .SE(n8230), .CLK(n8417), .Q(
        g1680), .QN(n4488) );
  SDFFX1 DFF_1017_Q_reg ( .D(n456), .SI(g1680), .SE(n8231), .CLK(n8418), .Q(
        g1686) );
  SDFFX1 DFF_1028_Q_reg ( .D(n4276), .SI(g1686), .SE(n8231), .CLK(n8418), .Q(
        n7978) );
  SDFFX1 DFF_1029_Q_reg ( .D(g1735), .SI(n7978), .SE(n8231), .CLK(n8418), .Q(
        g1723) );
  SDFFX1 DFF_1030_Q_reg ( .D(g1723), .SI(g1723), .SE(n8231), .CLK(n8418), .Q(
        g1730) );
  SDFFX1 DFF_1031_Q_reg ( .D(g1724), .SI(g1730), .SE(n8231), .CLK(n8418), .Q(
        g1731) );
  SDFFX1 DFF_1032_Q_reg ( .D(g1731), .SI(g1731), .SE(n8232), .CLK(n8419), .Q(
        g1732) );
  SDFFX1 DFF_1033_Q_reg ( .D(g1727), .SI(g1732), .SE(n8232), .CLK(n8419), .Q(
        g1733) );
  SDFFX1 DFF_1034_Q_reg ( .D(g1733), .SI(g1733), .SE(n8232), .CLK(n8419), .Q(
        g1734) );
  SDFFX1 DFF_1035_Q_reg ( .D(g1750), .SI(g1734), .SE(n8232), .CLK(n8419), .Q(
        g1738) );
  SDFFX1 DFF_1036_Q_reg ( .D(g1738), .SI(g1738), .SE(n8232), .CLK(n8419), .Q(
        g1745) );
  SDFFX1 DFF_1037_Q_reg ( .D(g1739), .SI(g1745), .SE(n8232), .CLK(n8419), .Q(
        test_so62) );
  SDFFX1 DFF_1038_Q_reg ( .D(test_so62), .SI(test_si63), .SE(n8232), .CLK(
        n8419), .Q(g1747) );
  SDFFX1 DFF_1039_Q_reg ( .D(g1742), .SI(g1747), .SE(n8232), .CLK(n8419), .Q(
        g1748) );
  SDFFX1 DFF_1040_Q_reg ( .D(g1748), .SI(g1748), .SE(n8232), .CLK(n8419), .Q(
        g1749) );
  SDFFX1 DFF_1041_Q_reg ( .D(g1765), .SI(g1749), .SE(n8232), .CLK(n8419), .Q(
        g1753) );
  SDFFX1 DFF_1042_Q_reg ( .D(g1753), .SI(g1753), .SE(n8232), .CLK(n8419), .Q(
        g1760) );
  SDFFX1 DFF_1043_Q_reg ( .D(g1754), .SI(g1760), .SE(n8232), .CLK(n8419), .Q(
        g1761) );
  SDFFX1 DFF_1044_Q_reg ( .D(g1761), .SI(g1761), .SE(n8233), .CLK(n8420), .Q(
        g1762) );
  SDFFX1 DFF_1045_Q_reg ( .D(g1757), .SI(g1762), .SE(n8233), .CLK(n8420), .Q(
        g1763) );
  SDFFX1 DFF_1046_Q_reg ( .D(g1763), .SI(g1763), .SE(n8233), .CLK(n8420), .Q(
        g1764) );
  SDFFX1 DFF_1047_Q_reg ( .D(g1779), .SI(g1764), .SE(n8233), .CLK(n8420), .Q(
        g1768) );
  SDFFX1 DFF_1048_Q_reg ( .D(g1768), .SI(g1768), .SE(n8233), .CLK(n8420), .Q(
        g1775) );
  SDFFX1 DFF_1049_Q_reg ( .D(test_so58), .SI(g1775), .SE(n8233), .CLK(n8420), 
        .Q(g1776) );
  SDFFX1 DFF_1050_Q_reg ( .D(g1776), .SI(g1776), .SE(n8233), .CLK(n8420), .Q(
        g1777) );
  SDFFX1 DFF_1051_Q_reg ( .D(g1772), .SI(g1777), .SE(n8233), .CLK(n8420), .Q(
        g1778) );
  SDFFX1 DFF_1052_Q_reg ( .D(g1778), .SI(g1778), .SE(n8233), .CLK(n8420), .Q(
        g1705) );
  SDFFX1 DFF_1053_Q_reg ( .D(n4598), .SI(g1705), .SE(n8233), .CLK(n8420), .Q(
        test_so63) );
  SDFFX1 DFF_1054_Q_reg ( .D(test_so63), .SI(test_si64), .SE(n8233), .CLK(
        n8420), .Q(g5738) );
  SDFFX1 DFF_1055_Q_reg ( .D(g5738), .SI(g5738), .SE(n8233), .CLK(n8420), .Q(
        g1718) );
  SDFFX1 DFF_1056_Q_reg ( .D(n4598), .SI(g1718), .SE(n8234), .CLK(n8421), .Q(
        g7052), .QN(n4296) );
  SDFFX1 DFF_1057_Q_reg ( .D(g7052), .SI(g7052), .SE(n8234), .CLK(n8421), .Q(
        g7194), .QN(n4315) );
  SDFFX1 DFF_1058_Q_reg ( .D(g7194), .SI(g7194), .SE(n8234), .CLK(n8421), .Q(
        g1930), .QN(n4366) );
  SDFFX1 DFF_1059_Q_reg ( .D(n1149), .SI(g1930), .SE(n8234), .CLK(n8421), .Q(
        g1934), .QN(n7991) );
  SDFFX1 DFF_1060_Q_reg ( .D(g18743), .SI(g1934), .SE(n8234), .CLK(n8421), .Q(
        g1937), .QN(n4311) );
  SDFFX1 DFF_1061_Q_reg ( .D(g18794), .SI(g1937), .SE(n8234), .CLK(n8421), .Q(
        g1890), .QN(n4297) );
  SDFFX1 DFF_1062_Q_reg ( .D(n1145), .SI(g1890), .SE(n8235), .CLK(n8422), .Q(
        g1893) );
  SDFFX1 DFF_1063_Q_reg ( .D(g1893), .SI(g1893), .SE(n8235), .CLK(n8422), .Q(
        g1903) );
  SDFFX1 DFF_1064_Q_reg ( .D(g1903), .SI(g1903), .SE(n8235), .CLK(n8422), .Q(
        g1904) );
  SDFFX1 DFF_1065_Q_reg ( .D(g1836), .SI(g1904), .SE(n8235), .CLK(n8422), .Q(
        g1944) );
  SDFFX1 DFF_1066_Q_reg ( .D(g1944), .SI(g1944), .SE(n8235), .CLK(n8422), .Q(
        g1949) );
  SDFFX1 DFF_1067_Q_reg ( .D(test_so65), .SI(g1949), .SE(n8235), .CLK(n8422), 
        .Q(g1950) );
  SDFFX1 DFF_1068_Q_reg ( .D(g1950), .SI(g1950), .SE(n8236), .CLK(n8423), .Q(
        g1951) );
  SDFFX1 DFF_1069_Q_reg ( .D(g1842), .SI(g1951), .SE(n8236), .CLK(n8423), .Q(
        test_so64) );
  SDFFX1 DFF_1070_Q_reg ( .D(test_so64), .SI(test_si65), .SE(n8236), .CLK(
        n8423), .Q(g1953) );
  SDFFX1 DFF_1071_Q_reg ( .D(g1846), .SI(g1953), .SE(n8236), .CLK(n8423), .Q(
        g1954) );
  SDFFX1 DFF_1072_Q_reg ( .D(g1954), .SI(g1954), .SE(n8236), .CLK(n8423), .Q(
        g1945) );
  SDFFX1 DFF_1073_Q_reg ( .D(g1849), .SI(g1945), .SE(n8236), .CLK(n8423), .Q(
        g1946) );
  SDFFX1 DFF_1074_Q_reg ( .D(g1946), .SI(g1946), .SE(n8236), .CLK(n8423), .Q(
        g1947) );
  SDFFX1 DFF_1075_Q_reg ( .D(g1852), .SI(g1947), .SE(n8236), .CLK(n8423), .Q(
        g1948) );
  SDFFX1 DFF_1076_Q_reg ( .D(g1948), .SI(g1948), .SE(n8236), .CLK(n8423), .Q(
        g1870) );
  SDFFX1 DFF_1077_Q_reg ( .D(g2950), .SI(g1870), .SE(n8236), .CLK(n8423), .Q(
        g8012), .QN(n4458) );
  SDFFX1 DFF_1078_Q_reg ( .D(g8012), .SI(g8012), .SE(n8236), .CLK(n8423), .Q(
        g8082), .QN(n4457) );
  SDFFX1 DFF_1079_Q_reg ( .D(g8082), .SI(g8082), .SE(n8236), .CLK(n8423), .Q(
        g1866), .QN(n4464) );
  SDFFX1 DFF_1080_Q_reg ( .D(g23097), .SI(g1866), .SE(n8237), .CLK(n8424), .Q(
        g1867) );
  SDFFX1 DFF_1081_Q_reg ( .D(g23124), .SI(g1867), .SE(n8237), .CLK(n8424), .Q(
        g1868) );
  SDFFX1 DFF_1082_Q_reg ( .D(g23137), .SI(g1868), .SE(n8237), .CLK(n8424), .Q(
        g1869) );
  SDFFX1 DFF_1083_Q_reg ( .D(g23400), .SI(g1869), .SE(n8237), .CLK(n8424), .Q(
        g1836) );
  SDFFX1 DFF_1084_Q_reg ( .D(g23413), .SI(g1836), .SE(n8237), .CLK(n8424), .Q(
        test_so65) );
  SDFFX1 DFF_1085_Q_reg ( .D(g24182), .SI(test_si66), .SE(n8237), .CLK(n8424), 
        .Q(g1842) );
  SDFFX1 DFF_1086_Q_reg ( .D(g24208), .SI(g1842), .SE(n8237), .CLK(n8424), .Q(
        g1858) );
  SDFFX1 DFF_1087_Q_reg ( .D(g24219), .SI(g1858), .SE(n8237), .CLK(n8424), .Q(
        g1859) );
  SDFFX1 DFF_1088_Q_reg ( .D(g24231), .SI(g1859), .SE(n8237), .CLK(n8424), .Q(
        g1860) );
  SDFFX1 DFF_1089_Q_reg ( .D(g23123), .SI(g1860), .SE(n8237), .CLK(n8424), .Q(
        g1861) );
  SDFFX1 DFF_1090_Q_reg ( .D(g23030), .SI(g1861), .SE(n8237), .CLK(n8424), .Q(
        g1865) );
  SDFFX1 DFF_1091_Q_reg ( .D(g23058), .SI(g1865), .SE(n8237), .CLK(n8424), .Q(
        g1845) );
  SDFFX1 DFF_1092_Q_reg ( .D(g24218), .SI(g1845), .SE(n8238), .CLK(n8425), .Q(
        g1846) );
  SDFFX1 DFF_1093_Q_reg ( .D(g24230), .SI(g1846), .SE(n8238), .CLK(n8425), .Q(
        g1849) );
  SDFFX1 DFF_1094_Q_reg ( .D(g24243), .SI(g1849), .SE(n8238), .CLK(n8425), .Q(
        g1852) );
  SDFFX1 DFF_1095_Q_reg ( .D(n1122), .SI(g1852), .SE(n8238), .CLK(n8425), .Q(
        g1908) );
  SDFFX1 DFF_1096_Q_reg ( .D(g1908), .SI(g1908), .SE(n8238), .CLK(n8425), .Q(
        g1915) );
  SDFFX1 DFF_1097_Q_reg ( .D(g1915), .SI(g1915), .SE(n8238), .CLK(n8425), .Q(
        g1922) );
  SDFFX1 DFF_1098_Q_reg ( .D(g13164), .SI(g1922), .SE(n8238), .CLK(n8425), .Q(
        g1923) );
  SDFFX1 DFF_1099_Q_reg ( .D(g1923), .SI(g1923), .SE(n8238), .CLK(n8425), .Q(
        test_so66), .QN(DFF_1099_n1) );
  SDFFX1 DFF_1100_Q_reg ( .D(n516), .SI(test_si67), .SE(n8239), .CLK(n8426), 
        .Q(n7971) );
  SDFFX1 DFF_1101_Q_reg ( .D(g13135), .SI(n7971), .SE(n8238), .CLK(n8425), .Q(
        g1929) );
  SDFFX1 DFF_1102_Q_reg ( .D(g1929), .SI(g1929), .SE(n8238), .CLK(n8425), .Q(
        g1880), .QN(n4545) );
  SDFFX1 DFF_1103_Q_reg ( .D(g13182), .SI(g1880), .SE(n8238), .CLK(n8425), .Q(
        g1938) );
  SDFFX1 DFF_1104_Q_reg ( .D(g1938), .SI(g1938), .SE(n8238), .CLK(n8425), .Q(
        g1939), .QN(n7762) );
  SDFFX1 DFF_1105_Q_reg ( .D(g27290), .SI(g1939), .SE(n8240), .CLK(n8427), .Q(
        g1956), .QN(n7341) );
  SDFFX1 DFF_1106_Q_reg ( .D(g27305), .SI(g1956), .SE(n8240), .CLK(n8427), .Q(
        g1957), .QN(n7343) );
  SDFFX1 DFF_1107_Q_reg ( .D(g27319), .SI(g1957), .SE(n8240), .CLK(n8427), .Q(
        g1955), .QN(n7342) );
  SDFFX1 DFF_1108_Q_reg ( .D(g27306), .SI(g1955), .SE(n8240), .CLK(n8427), .Q(
        g1959), .QN(n7353) );
  SDFFX1 DFF_1109_Q_reg ( .D(g27320), .SI(g1959), .SE(n8240), .CLK(n8427), .Q(
        g1960), .QN(n7355) );
  SDFFX1 DFF_1110_Q_reg ( .D(g27331), .SI(g1960), .SE(n8240), .CLK(n8427), .Q(
        g1958), .QN(n7354) );
  SDFFX1 DFF_1111_Q_reg ( .D(g27321), .SI(g1958), .SE(n8241), .CLK(n8428), .Q(
        g1962), .QN(n7179) );
  SDFFX1 DFF_1112_Q_reg ( .D(g27332), .SI(g1962), .SE(n8241), .CLK(n8428), .Q(
        g1963), .QN(n7181) );
  SDFFX1 DFF_1113_Q_reg ( .D(g27340), .SI(g1963), .SE(n8240), .CLK(n8427), .Q(
        g1961), .QN(n7180) );
  SDFFX1 DFF_1114_Q_reg ( .D(g27333), .SI(g1961), .SE(n8241), .CLK(n8428), .Q(
        test_so67), .QN(n8109) );
  SDFFX1 DFF_1115_Q_reg ( .D(g27341), .SI(test_si68), .SE(n8241), .CLK(n8428), 
        .Q(g1966), .QN(n7365) );
  SDFFX1 DFF_1116_Q_reg ( .D(g27346), .SI(g1966), .SE(n8239), .CLK(n8426), .Q(
        g1964), .QN(n7364) );
  SDFFX1 DFF_1117_Q_reg ( .D(g24513), .SI(g1964), .SE(n8239), .CLK(n8426), .Q(
        g1967) );
  SDFFX1 DFF_1118_Q_reg ( .D(g24524), .SI(g1967), .SE(n8240), .CLK(n8427), .Q(
        g1970) );
  SDFFX1 DFF_1119_Q_reg ( .D(g24534), .SI(g1970), .SE(n8240), .CLK(n8427), .Q(
        g1973) );
  SDFFX1 DFF_1120_Q_reg ( .D(g24525), .SI(g1973), .SE(n8240), .CLK(n8427), .Q(
        g1976) );
  SDFFX1 DFF_1121_Q_reg ( .D(g24535), .SI(g1976), .SE(n8240), .CLK(n8427), .Q(
        g1979) );
  SDFFX1 DFF_1122_Q_reg ( .D(g24545), .SI(g1979), .SE(n8240), .CLK(n8427), .Q(
        g1982) );
  SDFFX1 DFF_1123_Q_reg ( .D(g28357), .SI(g1982), .SE(n8241), .CLK(n8428), .Q(
        g1994) );
  SDFFX1 DFF_1124_Q_reg ( .D(g28362), .SI(g1994), .SE(n8241), .CLK(n8428), .Q(
        g1997) );
  SDFFX1 DFF_1125_Q_reg ( .D(g28366), .SI(g1997), .SE(n8241), .CLK(n8428), .Q(
        g2000) );
  SDFFX1 DFF_1126_Q_reg ( .D(g28352), .SI(g2000), .SE(n8241), .CLK(n8428), .Q(
        g1985) );
  SDFFX1 DFF_1127_Q_reg ( .D(g28356), .SI(g1985), .SE(n8241), .CLK(n8428), .Q(
        g1988) );
  SDFFX1 DFF_1128_Q_reg ( .D(g28361), .SI(g1988), .SE(n8241), .CLK(n8428), .Q(
        g1991) );
  SDFFX1 DFF_1129_Q_reg ( .D(g26559), .SI(g1991), .SE(n8241), .CLK(n8428), .Q(
        test_so68) );
  SDFFX1 DFF_1130_Q_reg ( .D(g26573), .SI(test_si69), .SE(n8241), .CLK(n8428), 
        .Q(g1874) );
  SDFFX1 DFF_1131_Q_reg ( .D(g26592), .SI(g1874), .SE(n8242), .CLK(n8429), .Q(
        g1877) );
  SDFFX1 DFF_1132_Q_reg ( .D(g1880), .SI(g1877), .SE(n8242), .CLK(n8429), .Q(
        g1886), .QN(n4493) );
  SDFFX1 DFF_1133_Q_reg ( .D(g22651), .SI(g1886), .SE(n8242), .CLK(n8429), .Q(
        n7968), .QN(DFF_1133_n1) );
  SDFFX1 DFF_1142_Q_reg ( .D(n531), .SI(n7968), .SE(n8242), .CLK(n8429), .Q(
        g16399), .QN(DFF_1142_n1) );
  SDFFX1 DFF_1143_Q_reg ( .D(g16399), .SI(g16399), .SE(n8242), .CLK(n8429), 
        .Q(g1905), .QN(n8064) );
  SDFFX1 DFF_1144_Q_reg ( .D(DFF_999_n1), .SI(g1905), .SE(n8242), .CLK(n8429), 
        .Q(n7967), .QN(DFF_1144_n1) );
  SDFFX1 DFF_1145_Q_reg ( .D(DFF_1001_n1), .SI(n7967), .SE(n8242), .CLK(n8429), 
        .Q(n7966), .QN(DFF_1145_n1) );
  SDFFX1 DFF_1146_Q_reg ( .D(DFF_1003_n1), .SI(n7966), .SE(n8242), .CLK(n8429), 
        .Q(n7965), .QN(DFF_1146_n1) );
  SDFFX1 DFF_1147_Q_reg ( .D(DFF_1005_n1), .SI(n7965), .SE(n8242), .CLK(n8429), 
        .Q(n7964), .QN(DFF_1147_n1) );
  SDFFX1 DFF_1148_Q_reg ( .D(DFF_1007_n1), .SI(n7964), .SE(n8242), .CLK(n8429), 
        .Q(n7963), .QN(DFF_1148_n1) );
  SDFFX1 DFF_1149_Q_reg ( .D(DFF_1009_n1), .SI(n7963), .SE(n8242), .CLK(n8429), 
        .Q(n7962), .QN(DFF_1149_n1) );
  SDFFX1 DFF_1150_Q_reg ( .D(DFF_1011_n1), .SI(n7962), .SE(n8242), .CLK(n8429), 
        .Q(g1916), .QN(n7159) );
  SDFFX1 DFF_1151_Q_reg ( .D(DFF_1013_n1), .SI(g1916), .SE(n8243), .CLK(n8430), 
        .Q(g1917), .QN(n7158) );
  SDFFX1 DFF_1152_Q_reg ( .D(g24083), .SI(g1917), .SE(n8243), .CLK(n8430), .Q(
        test_so69), .QN(n8111) );
  SDFFX1 DFF_1153_Q_reg ( .D(n4484), .SI(test_si70), .SE(n8149), .CLK(n8336), 
        .Q(n7960), .QN(n14380) );
  SDFFX1 DFF_1155_Q_reg ( .D(g7229), .SI(g7229), .SE(n8172), .CLK(n8359), .Q(
        g7357), .QN(n4357) );
  SDFFX1 DFF_1156_Q_reg ( .D(g7357), .SI(g7357), .SE(n8172), .CLK(n8359), .Q(
        g2009), .QN(n4293) );
  SDFFX1 DFF_1157_Q_reg ( .D(g16692), .SI(g2009), .SE(n8234), .CLK(n8421), .Q(
        g2010), .QN(n7758) );
  SDFFX1 DFF_1158_Q_reg ( .D(g20353), .SI(g2010), .SE(n8234), .CLK(n8421), .Q(
        g2039), .QN(n4427) );
  SDFFX1 DFF_1159_Q_reg ( .D(g20752), .SI(g2039), .SE(n8234), .CLK(n8421), .Q(
        g2020), .QN(n4400) );
  SDFFX1 DFF_1160_Q_reg ( .D(n1222), .SI(g2020), .SE(n8234), .CLK(n8421), .Q(
        g2013), .QN(n4474) );
  SDFFX1 DFF_1161_Q_reg ( .D(g23339), .SI(g2013), .SE(n8234), .CLK(n8421), .Q(
        g2033), .QN(n4420) );
  SDFFX1 DFF_1162_Q_reg ( .D(g24434), .SI(g2033), .SE(n8234), .CLK(n8421), .Q(
        g2026), .QN(n4410) );
  SDFFX1 DFF_1163_Q_reg ( .D(g25194), .SI(g2026), .SE(n8235), .CLK(n8422), .Q(
        g2040), .QN(n4399) );
  SDFFX1 DFF_1164_Q_reg ( .D(n1223), .SI(g2040), .SE(n8235), .CLK(n8422), .Q(
        g2052), .QN(n4409) );
  SDFFX1 DFF_1165_Q_reg ( .D(g26789), .SI(g2052), .SE(n8235), .CLK(n8422), .Q(
        g2046), .QN(n4468) );
  SDFFX1 DFF_1166_Q_reg ( .D(g27682), .SI(g2046), .SE(n8235), .CLK(n8422), .Q(
        g2059), .QN(n4473) );
  SDFFX1 DFF_1167_Q_reg ( .D(g27722), .SI(g2059), .SE(n8235), .CLK(n8422), .Q(
        test_so70), .QN(n8106) );
  SDFFX1 DFF_1168_Q_reg ( .D(g28325), .SI(test_si71), .SE(n8235), .CLK(n8422), 
        .Q(g2072), .QN(n4416) );
  SDFFX1 DFF_1169_Q_reg ( .D(g20899), .SI(g2072), .SE(n8243), .CLK(n8430), .Q(
        g2079), .QN(n7802) );
  SDFFX1 DFF_1170_Q_reg ( .D(g20915), .SI(g2079), .SE(n8243), .CLK(n8430), .Q(
        g2080), .QN(n7801) );
  SDFFX1 DFF_1171_Q_reg ( .D(g20934), .SI(g2080), .SE(n8243), .CLK(n8430), .Q(
        g2078), .QN(n7856) );
  SDFFX1 DFF_1172_Q_reg ( .D(g20916), .SI(g2078), .SE(n8243), .CLK(n8430), .Q(
        g2082), .QN(n7800) );
  SDFFX1 DFF_1173_Q_reg ( .D(g20935), .SI(g2082), .SE(n8243), .CLK(n8430), .Q(
        g2083), .QN(n7799) );
  SDFFX1 DFF_1174_Q_reg ( .D(g20953), .SI(g2083), .SE(n8244), .CLK(n8431), .Q(
        g2081), .QN(n7855) );
  SDFFX1 DFF_1175_Q_reg ( .D(g20936), .SI(g2081), .SE(n8244), .CLK(n8431), .Q(
        g2085), .QN(n7798) );
  SDFFX1 DFF_1176_Q_reg ( .D(g20954), .SI(g2085), .SE(n8244), .CLK(n8431), .Q(
        g2086), .QN(n7797) );
  SDFFX1 DFF_1177_Q_reg ( .D(g20977), .SI(g2086), .SE(n8244), .CLK(n8431), .Q(
        g2084), .QN(n7854) );
  SDFFX1 DFF_1178_Q_reg ( .D(g20955), .SI(g2084), .SE(n8244), .CLK(n8431), .Q(
        g2088), .QN(n7796) );
  SDFFX1 DFF_1179_Q_reg ( .D(g20978), .SI(g2088), .SE(n8244), .CLK(n8431), .Q(
        g2089), .QN(n7795) );
  SDFFX1 DFF_1180_Q_reg ( .D(g20999), .SI(g2089), .SE(n8244), .CLK(n8431), .Q(
        g2087), .QN(n7853) );
  SDFFX1 DFF_1181_Q_reg ( .D(g20979), .SI(g2087), .SE(n8244), .CLK(n8431), .Q(
        g2091), .QN(n7794) );
  SDFFX1 DFF_1182_Q_reg ( .D(g21000), .SI(g2091), .SE(n8244), .CLK(n8431), .Q(
        test_so71), .QN(n8133) );
  SDFFX1 DFF_1183_Q_reg ( .D(g21019), .SI(test_si72), .SE(n8244), .CLK(n8431), 
        .Q(g2090), .QN(n7852) );
  SDFFX1 DFF_1184_Q_reg ( .D(g21001), .SI(g2090), .SE(n8245), .CLK(n8432), .Q(
        g2094), .QN(n7793) );
  SDFFX1 DFF_1185_Q_reg ( .D(g21020), .SI(g2094), .SE(n8245), .CLK(n8432), .Q(
        g2095), .QN(n7792) );
  SDFFX1 DFF_1186_Q_reg ( .D(g21039), .SI(g2095), .SE(n8245), .CLK(n8432), .Q(
        g2093), .QN(n7851) );
  SDFFX1 DFF_1187_Q_reg ( .D(g21021), .SI(g2093), .SE(n8245), .CLK(n8432), .Q(
        g2097), .QN(n7791) );
  SDFFX1 DFF_1188_Q_reg ( .D(g21040), .SI(g2097), .SE(n8245), .CLK(n8432), .Q(
        g2098), .QN(n7790) );
  SDFFX1 DFF_1189_Q_reg ( .D(g21054), .SI(g2098), .SE(n8245), .CLK(n8432), .Q(
        g2096), .QN(n7850) );
  SDFFX1 DFF_1190_Q_reg ( .D(g21041), .SI(g2096), .SE(n8245), .CLK(n8432), .Q(
        g2100), .QN(n7789) );
  SDFFX1 DFF_1191_Q_reg ( .D(g21055), .SI(g2100), .SE(n8245), .CLK(n8432), .Q(
        g2101), .QN(n7788) );
  SDFFX1 DFF_1192_Q_reg ( .D(g21071), .SI(g2101), .SE(n8245), .CLK(n8432), .Q(
        g2099), .QN(n7849) );
  SDFFX1 DFF_1193_Q_reg ( .D(g21056), .SI(g2099), .SE(n8245), .CLK(n8432), .Q(
        g2103), .QN(n7787) );
  SDFFX1 DFF_1194_Q_reg ( .D(g21072), .SI(g2103), .SE(n8245), .CLK(n8432), .Q(
        g2104), .QN(n7786) );
  SDFFX1 DFF_1195_Q_reg ( .D(g21080), .SI(g2104), .SE(n8245), .CLK(n8432), .Q(
        g2102), .QN(n7848) );
  SDFFX1 DFF_1196_Q_reg ( .D(g20900), .SI(g2102), .SE(n8246), .CLK(n8433), .Q(
        g2106), .QN(n7785) );
  SDFFX1 DFF_1197_Q_reg ( .D(g20917), .SI(g2106), .SE(n8246), .CLK(n8433), .Q(
        test_so72), .QN(n8134) );
  SDFFX1 DFF_1198_Q_reg ( .D(g20937), .SI(test_si73), .SE(n8243), .CLK(n8430), 
        .Q(g2105), .QN(n7847) );
  SDFFX1 DFF_1199_Q_reg ( .D(g20980), .SI(g2105), .SE(n8243), .CLK(n8430), .Q(
        g2109), .QN(n8041) );
  SDFFX1 DFF_1200_Q_reg ( .D(g21002), .SI(g2109), .SE(n8243), .CLK(n8430), .Q(
        g2110), .QN(n7570) );
  SDFFX1 DFF_1201_Q_reg ( .D(g21022), .SI(g2110), .SE(n8243), .CLK(n8430), .Q(
        g2108) );
  SDFFX1 DFF_1202_Q_reg ( .D(g21003), .SI(g2108), .SE(n8243), .CLK(n8430), .Q(
        g2112), .QN(n7576) );
  SDFFX1 DFF_1203_Q_reg ( .D(g21023), .SI(g2112), .SE(n8244), .CLK(n8431), .Q(
        g2113), .QN(n7569) );
  SDFFX1 DFF_1204_Q_reg ( .D(g21042), .SI(g2113), .SE(n8244), .CLK(n8431), .Q(
        g2111), .QN(n7627) );
  SDFFX1 DFF_1205_Q_reg ( .D(g25268), .SI(g2111), .SE(n8246), .CLK(n8433), .Q(
        g2115), .QN(n7505) );
  SDFFX1 DFF_1206_Q_reg ( .D(g25271), .SI(g2115), .SE(n8246), .CLK(n8433), .Q(
        g2116), .QN(n7504) );
  SDFFX1 DFF_1207_Q_reg ( .D(g25279), .SI(g2116), .SE(n8246), .CLK(n8433), .Q(
        g2114), .QN(n7511) );
  SDFFX1 DFF_1208_Q_reg ( .D(g22249), .SI(g2114), .SE(n8246), .CLK(n8433), .Q(
        g2118), .QN(n7878) );
  SDFFX1 DFF_1209_Q_reg ( .D(n1194), .SI(g2118), .SE(n8246), .CLK(n8433), .Q(
        g2119), .QN(n7975) );
  SDFFX1 DFF_1210_Q_reg ( .D(g22280), .SI(g2119), .SE(n8246), .CLK(n8433), .Q(
        g2117), .QN(n7981) );
  SDFFX1 DFF_1211_Q_reg ( .D(g2950), .SI(g2117), .SE(n8246), .CLK(n8433), .Q(
        g6837), .QN(n4324) );
  SDFFX1 DFF_1212_Q_reg ( .D(g6837), .SI(g6837), .SE(n8246), .CLK(n8433), .Q(
        test_so73), .QN(n8097) );
  SDFFX1 DFF_1213_Q_reg ( .D(test_so73), .SI(test_si74), .SE(n8246), .CLK(
        n8433), .Q(g2241), .QN(n4367) );
  SDFFX1 DFF_1214_Q_reg ( .D(g22170), .SI(g2241), .SE(n8246), .CLK(n8433), .Q(
        g2206), .QN(n7895) );
  SDFFX1 DFF_1215_Q_reg ( .D(g22182), .SI(g2206), .SE(n8251), .CLK(n8438), .Q(
        g2207), .QN(n7894) );
  SDFFX1 DFF_1216_Q_reg ( .D(g22192), .SI(g2207), .SE(n8251), .CLK(n8438), .Q(
        g2205), .QN(n7532) );
  SDFFX1 DFF_1217_Q_reg ( .D(g22183), .SI(g2205), .SE(n8247), .CLK(n8434), .Q(
        g2209), .QN(n7893) );
  SDFFX1 DFF_1218_Q_reg ( .D(g22193), .SI(g2209), .SE(n8251), .CLK(n8438), .Q(
        g2210), .QN(n7892) );
  SDFFX1 DFF_1219_Q_reg ( .D(g22200), .SI(g2210), .SE(n8251), .CLK(n8438), .Q(
        g2208), .QN(n7531) );
  SDFFX1 DFF_1220_Q_reg ( .D(g22045), .SI(g2208), .SE(n8251), .CLK(n8438), .Q(
        g2218), .QN(n7891) );
  SDFFX1 DFF_1221_Q_reg ( .D(g22060), .SI(g2218), .SE(n8251), .CLK(n8438), .Q(
        g2219), .QN(n7890) );
  SDFFX1 DFF_1222_Q_reg ( .D(g22076), .SI(g2219), .SE(n8251), .CLK(n8438), .Q(
        g2217), .QN(n7530) );
  SDFFX1 DFF_1223_Q_reg ( .D(g22061), .SI(g2217), .SE(n8251), .CLK(n8438), .Q(
        g2221), .QN(n7889) );
  SDFFX1 DFF_1224_Q_reg ( .D(g22077), .SI(g2221), .SE(n8251), .CLK(n8438), .Q(
        g2222), .QN(n7888) );
  SDFFX1 DFF_1225_Q_reg ( .D(g22097), .SI(g2222), .SE(n8252), .CLK(n8439), .Q(
        g2220), .QN(n7529) );
  SDFFX1 DFF_1226_Q_reg ( .D(g22078), .SI(g2220), .SE(n8252), .CLK(n8439), .Q(
        g2224), .QN(n7887) );
  SDFFX1 DFF_1227_Q_reg ( .D(g22098), .SI(g2224), .SE(n8252), .CLK(n8439), .Q(
        test_so74), .QN(n8130) );
  SDFFX1 DFF_1228_Q_reg ( .D(g22115), .SI(test_si75), .SE(n8249), .CLK(n8436), 
        .Q(g2223), .QN(n7528) );
  SDFFX1 DFF_1229_Q_reg ( .D(g22099), .SI(g2223), .SE(n8249), .CLK(n8436), .Q(
        g2227), .QN(n7886) );
  SDFFX1 DFF_1230_Q_reg ( .D(g22116), .SI(g2227), .SE(n8250), .CLK(n8437), .Q(
        g2228), .QN(n7885) );
  SDFFX1 DFF_1231_Q_reg ( .D(g22138), .SI(g2228), .SE(n8250), .CLK(n8437), .Q(
        g2226), .QN(n7527) );
  SDFFX1 DFF_1232_Q_reg ( .D(g22117), .SI(g2226), .SE(n8250), .CLK(n8437), .Q(
        g2230), .QN(n7884) );
  SDFFX1 DFF_1233_Q_reg ( .D(g22139), .SI(g2230), .SE(n8250), .CLK(n8437), .Q(
        g2231), .QN(n7883) );
  SDFFX1 DFF_1234_Q_reg ( .D(g22153), .SI(g2231), .SE(n8250), .CLK(n8437), .Q(
        g2229), .QN(n7526) );
  SDFFX1 DFF_1235_Q_reg ( .D(g22140), .SI(g2229), .SE(n8250), .CLK(n8437), .Q(
        g2233), .QN(n7882) );
  SDFFX1 DFF_1236_Q_reg ( .D(g22154), .SI(g2233), .SE(n8250), .CLK(n8437), .Q(
        g2234), .QN(n7881) );
  SDFFX1 DFF_1237_Q_reg ( .D(g22171), .SI(g2234), .SE(n8250), .CLK(n8437), .Q(
        g2232), .QN(n7525) );
  SDFFX1 DFF_1238_Q_reg ( .D(g22155), .SI(g2232), .SE(n8250), .CLK(n8437), .Q(
        g2236), .QN(n7516) );
  SDFFX1 DFF_1239_Q_reg ( .D(g22172), .SI(g2236), .SE(n8250), .CLK(n8437), .Q(
        g2237), .QN(n7515) );
  SDFFX1 DFF_1240_Q_reg ( .D(g22184), .SI(g2237), .SE(n8251), .CLK(n8438), .Q(
        g2235), .QN(n7514) );
  SDFFX1 DFF_1241_Q_reg ( .D(g22173), .SI(g2235), .SE(n8251), .CLK(n8438), .Q(
        g2239), .QN(n7524) );
  SDFFX1 DFF_1242_Q_reg ( .D(g22185), .SI(g2239), .SE(n8251), .CLK(n8438), .Q(
        test_so75), .QN(n8129) );
  SDFFX1 DFF_1243_Q_reg ( .D(g22194), .SI(test_si76), .SE(n8249), .CLK(n8436), 
        .Q(g2238), .QN(n7523) );
  SDFFX1 DFF_1244_Q_reg ( .D(g25227), .SI(g2238), .SE(n8249), .CLK(n8436), .Q(
        g2245), .QN(n7590) );
  SDFFX1 DFF_1245_Q_reg ( .D(g25236), .SI(g2245), .SE(n8249), .CLK(n8436), .Q(
        g2246), .QN(n7589) );
  SDFFX1 DFF_1246_Q_reg ( .D(g25245), .SI(g2246), .SE(n8249), .CLK(n8436), .Q(
        g2244), .QN(n7588) );
  SDFFX1 DFF_1247_Q_reg ( .D(g25237), .SI(g2244), .SE(n8249), .CLK(n8436), .Q(
        g2248), .QN(n7587) );
  SDFFX1 DFF_1248_Q_reg ( .D(g25246), .SI(g2248), .SE(n8249), .CLK(n8436), .Q(
        g2249), .QN(n7586) );
  SDFFX1 DFF_1249_Q_reg ( .D(g25251), .SI(g2249), .SE(n8249), .CLK(n8436), .Q(
        g2247), .QN(n7585) );
  SDFFX1 DFF_1250_Q_reg ( .D(g25247), .SI(g2247), .SE(n8249), .CLK(n8436), .Q(
        g2251), .QN(n7584) );
  SDFFX1 DFF_1251_Q_reg ( .D(g25252), .SI(g2251), .SE(n8249), .CLK(n8436), .Q(
        g2252), .QN(n7583) );
  SDFFX1 DFF_1252_Q_reg ( .D(g25256), .SI(g2252), .SE(n8249), .CLK(n8436), .Q(
        g2250), .QN(n7582) );
  SDFFX1 DFF_1253_Q_reg ( .D(g25253), .SI(g2250), .SE(n8250), .CLK(n8437), .Q(
        g2254), .QN(n7581) );
  SDFFX1 DFF_1254_Q_reg ( .D(g25257), .SI(g2254), .SE(n8250), .CLK(n8437), .Q(
        g2255), .QN(n7580) );
  SDFFX1 DFF_1255_Q_reg ( .D(g25259), .SI(g2255), .SE(n8146), .CLK(n8333), .Q(
        g2253), .QN(n7579) );
  SDFFX1 DFF_1256_Q_reg ( .D(g30289), .SI(g2253), .SE(n8260), .CLK(n8447), .Q(
        g2261) );
  SDFFX1 DFF_1257_Q_reg ( .D(g30296), .SI(g2261), .SE(n8260), .CLK(n8447), .Q(
        test_so76) );
  SDFFX1 DFF_1258_Q_reg ( .D(g30300), .SI(test_si77), .SE(n8260), .CLK(n8447), 
        .Q(g2267) );
  SDFFX1 DFF_1259_Q_reg ( .D(g30660), .SI(g2267), .SE(n8260), .CLK(n8447), .Q(
        g2306) );
  SDFFX1 DFF_1260_Q_reg ( .D(g30666), .SI(g2306), .SE(n8261), .CLK(n8448), .Q(
        g2309) );
  SDFFX1 DFF_1261_Q_reg ( .D(g30672), .SI(g2309), .SE(n8261), .CLK(n8448), .Q(
        g2312) );
  SDFFX1 DFF_1262_Q_reg ( .D(g30690), .SI(g2312), .SE(n8261), .CLK(n8448), .Q(
        g2270) );
  SDFFX1 DFF_1263_Q_reg ( .D(g30693), .SI(g2270), .SE(n8261), .CLK(n8448), .Q(
        g2273) );
  SDFFX1 DFF_1264_Q_reg ( .D(g30695), .SI(g2273), .SE(n8252), .CLK(n8439), .Q(
        g2276) );
  SDFFX1 DFF_1265_Q_reg ( .D(g30667), .SI(g2276), .SE(n8252), .CLK(n8439), .Q(
        g2315) );
  SDFFX1 DFF_1266_Q_reg ( .D(g30673), .SI(g2315), .SE(n8252), .CLK(n8439), .Q(
        g2318) );
  SDFFX1 DFF_1267_Q_reg ( .D(g30679), .SI(g2318), .SE(n8252), .CLK(n8439), .Q(
        g2321) );
  SDFFX1 DFF_1268_Q_reg ( .D(g30301), .SI(g2321), .SE(n8252), .CLK(n8439), .Q(
        g2279) );
  SDFFX1 DFF_1269_Q_reg ( .D(g30303), .SI(g2279), .SE(n8252), .CLK(n8439), .Q(
        g2282) );
  SDFFX1 DFF_1270_Q_reg ( .D(g30304), .SI(g2282), .SE(n8252), .CLK(n8439), .Q(
        g2285) );
  SDFFX1 DFF_1271_Q_reg ( .D(g30274), .SI(g2285), .SE(n8252), .CLK(n8439), .Q(
        g2324) );
  SDFFX1 DFF_1272_Q_reg ( .D(g30282), .SI(g2324), .SE(n8252), .CLK(n8439), .Q(
        test_so77) );
  SDFFX1 DFF_1273_Q_reg ( .D(g30290), .SI(test_si78), .SE(n8253), .CLK(n8440), 
        .Q(g2330) );
  SDFFX1 DFF_1274_Q_reg ( .D(g30253), .SI(g2330), .SE(n8260), .CLK(n8447), .Q(
        g2288) );
  SDFFX1 DFF_1275_Q_reg ( .D(g30256), .SI(g2288), .SE(n8260), .CLK(n8447), .Q(
        g2291) );
  SDFFX1 DFF_1276_Q_reg ( .D(g30260), .SI(g2291), .SE(n8260), .CLK(n8447), .Q(
        g2294) );
  SDFFX1 DFF_1277_Q_reg ( .D(g30283), .SI(g2294), .SE(n8260), .CLK(n8447), .Q(
        g2333) );
  SDFFX1 DFF_1278_Q_reg ( .D(g30291), .SI(g2333), .SE(n8260), .CLK(n8447), .Q(
        g2336) );
  SDFFX1 DFF_1279_Q_reg ( .D(g30297), .SI(g2336), .SE(n8260), .CLK(n8447), .Q(
        g2339) );
  SDFFX1 DFF_1280_Q_reg ( .D(g30652), .SI(g2339), .SE(n8260), .CLK(n8447), .Q(
        g2297) );
  SDFFX1 DFF_1281_Q_reg ( .D(g30659), .SI(g2297), .SE(n8260), .CLK(n8447), .Q(
        g2300) );
  SDFFX1 DFF_1282_Q_reg ( .D(g30665), .SI(g2300), .SE(n8253), .CLK(n8440), .Q(
        g2303) );
  SDFFX1 DFF_1283_Q_reg ( .D(g30686), .SI(g2303), .SE(n8253), .CLK(n8440), .Q(
        g2342) );
  SDFFX1 DFF_1284_Q_reg ( .D(g30691), .SI(g2342), .SE(n8253), .CLK(n8440), .Q(
        g2345) );
  SDFFX1 DFF_1285_Q_reg ( .D(g30694), .SI(g2345), .SE(n8247), .CLK(n8434), .Q(
        g2348) );
  SDFFX1 DFF_1286_Q_reg ( .D(g25067), .SI(g2348), .SE(n8247), .CLK(n8434), .Q(
        g2160), .QN(n7702) );
  SDFFX1 DFF_1287_Q_reg ( .D(g25940), .SI(g2160), .SE(n8247), .CLK(n8434), .Q(
        test_so78) );
  SDFFX1 DFF_1288_Q_reg ( .D(g26532), .SI(test_si79), .SE(n8247), .CLK(n8434), 
        .Q(g2151), .QN(n7701) );
  SDFFX1 DFF_1289_Q_reg ( .D(g27131), .SI(g2151), .SE(n8247), .CLK(n8434), .Q(
        g2147), .QN(n8075) );
  SDFFX1 DFF_1290_Q_reg ( .D(g27621), .SI(g2147), .SE(n8247), .CLK(n8434), .Q(
        g2142), .QN(n7700) );
  SDFFX1 DFF_1291_Q_reg ( .D(g28148), .SI(g2142), .SE(n8247), .CLK(n8434), .Q(
        g2138), .QN(n8095) );
  SDFFX1 DFF_1292_Q_reg ( .D(g28637), .SI(g2138), .SE(n8247), .CLK(n8434), .Q(
        g2133), .QN(n7699) );
  SDFFX1 DFF_1293_Q_reg ( .D(g29112), .SI(g2133), .SE(n8247), .CLK(n8434), .Q(
        g2129), .QN(n8072) );
  SDFFX1 DFF_1294_Q_reg ( .D(g29357), .SI(g2129), .SE(n8248), .CLK(n8435), .Q(
        g2124), .QN(n7334) );
  SDFFX1 DFF_1295_Q_reg ( .D(g29582), .SI(g2124), .SE(n8248), .CLK(n8435), .Q(
        g2120), .QN(n7173) );
  SDFFX1 DFF_1296_Q_reg ( .D(n15), .SI(g2120), .SE(n8248), .CLK(n8435), .Q(
        g2256) );
  SDFFX1 DFF_1297_Q_reg ( .D(g2256), .SI(g2256), .SE(n8248), .CLK(n8435), .Q(
        g5637) );
  SDFFX1 DFF_1298_Q_reg ( .D(g5637), .SI(g5637), .SE(n8248), .CLK(n8435), .Q(
        g2257), .QN(n7718) );
  SDFFX1 DFF_1299_Q_reg ( .D(g2950), .SI(g2257), .SE(n8248), .CLK(n8435), .Q(
        g5555), .QN(n4516) );
  SDFFX1 DFF_1302_Q_reg ( .D(g5637), .SI(n4606), .SE(n8248), .CLK(n8435), .Q(
        test_so79), .QN(n8107) );
  SDFFX1 DFF_1303_Q_reg ( .D(g27276), .SI(test_si80), .SE(n8259), .CLK(n8446), 
        .Q(g2429), .QN(n7657) );
  SDFFX1 DFF_1304_Q_reg ( .D(g27291), .SI(g2429), .SE(n8259), .CLK(n8446), .Q(
        g2418), .QN(n7656) );
  SDFFX1 DFF_1305_Q_reg ( .D(g27307), .SI(g2418), .SE(n8259), .CLK(n8446), .Q(
        g2421), .QN(n7655) );
  SDFFX1 DFF_1306_Q_reg ( .D(g27292), .SI(g2421), .SE(n8259), .CLK(n8446), .Q(
        g2444), .QN(n7634) );
  SDFFX1 DFF_1307_Q_reg ( .D(g27308), .SI(g2444), .SE(n8259), .CLK(n8446), .Q(
        g2433), .QN(n7633) );
  SDFFX1 DFF_1308_Q_reg ( .D(g27322), .SI(g2433), .SE(n8259), .CLK(n8446), .Q(
        g2436), .QN(n7632) );
  SDFFX1 DFF_1309_Q_reg ( .D(g27309), .SI(g2436), .SE(n8259), .CLK(n8446), .Q(
        g2459), .QN(n7383) );
  SDFFX1 DFF_1310_Q_reg ( .D(g27323), .SI(g2459), .SE(n8259), .CLK(n8446), .Q(
        g2448), .QN(n7385) );
  SDFFX1 DFF_1311_Q_reg ( .D(g27334), .SI(g2448), .SE(n8259), .CLK(n8446), .Q(
        g2451), .QN(n7384) );
  SDFFX1 DFF_1312_Q_reg ( .D(g27324), .SI(g2451), .SE(n8259), .CLK(n8446), .Q(
        g2473), .QN(n7646) );
  SDFFX1 DFF_1313_Q_reg ( .D(g27335), .SI(g2473), .SE(n8259), .CLK(n8446), .Q(
        g2463), .QN(n7645) );
  SDFFX1 DFF_1314_Q_reg ( .D(g27342), .SI(g2463), .SE(n8253), .CLK(n8440), .Q(
        g2466), .QN(n7644) );
  SDFFX1 DFF_1315_Q_reg ( .D(g28763), .SI(g2466), .SE(n8253), .CLK(n8440), .Q(
        g2483) );
  SDFFX1 DFF_1316_Q_reg ( .D(g28773), .SI(g2483), .SE(n8258), .CLK(n8445), .Q(
        g2486) );
  SDFFX1 DFF_1317_Q_reg ( .D(g28782), .SI(g2486), .SE(n8258), .CLK(n8445), .Q(
        test_so80) );
  SDFFX1 DFF_1318_Q_reg ( .D(g29213), .SI(test_si81), .SE(n8253), .CLK(n8440), 
        .Q(g2492) );
  SDFFX1 DFF_1319_Q_reg ( .D(g29221), .SI(g2492), .SE(n8253), .CLK(n8440), .Q(
        g2495) );
  SDFFX1 DFF_1320_Q_reg ( .D(g29226), .SI(g2495), .SE(n8254), .CLK(n8441), .Q(
        g2498) );
  SDFFX1 DFF_1321_Q_reg ( .D(g28774), .SI(g2498), .SE(n8258), .CLK(n8445), .Q(
        g2502), .QN(n7678) );
  SDFFX1 DFF_1322_Q_reg ( .D(g28783), .SI(g2502), .SE(n8258), .CLK(n8445), .Q(
        g2503), .QN(n7668) );
  SDFFX1 DFF_1323_Q_reg ( .D(g28788), .SI(g2503), .SE(n8258), .CLK(n8445), .Q(
        g2501), .QN(n7677) );
  SDFFX1 DFF_1324_Q_reg ( .D(g26817), .SI(g2501), .SE(n8258), .CLK(n8445), .Q(
        g2504) );
  SDFFX1 DFF_1325_Q_reg ( .D(g26822), .SI(g2504), .SE(n8258), .CLK(n8445), .Q(
        g2507) );
  SDFFX1 DFF_1326_Q_reg ( .D(g26825), .SI(g2507), .SE(n8258), .CLK(n8445), .Q(
        g2510) );
  SDFFX1 DFF_1327_Q_reg ( .D(g26823), .SI(g2510), .SE(n8258), .CLK(n8445), .Q(
        g2513) );
  SDFFX1 DFF_1328_Q_reg ( .D(g26826), .SI(g2513), .SE(n8258), .CLK(n8445), .Q(
        g2516) );
  SDFFX1 DFF_1329_Q_reg ( .D(g26827), .SI(g2516), .SE(n8146), .CLK(n8333), .Q(
        g2519) );
  SDFFX1 DFF_1330_Q_reg ( .D(g27767), .SI(g2519), .SE(n8272), .CLK(n8459), .Q(
        g2523), .QN(n7676) );
  SDFFX1 DFF_1331_Q_reg ( .D(g27769), .SI(g2523), .SE(n8272), .CLK(n8459), .Q(
        g2524), .QN(n7667) );
  SDFFX1 DFF_1332_Q_reg ( .D(g27771), .SI(g2524), .SE(n8146), .CLK(n8333), .Q(
        test_so81), .QN(n8122) );
  SDFFX1 DFF_1333_Q_reg ( .D(g29618), .SI(test_si82), .SE(n8253), .CLK(n8440), 
        .Q(g2387), .QN(n7282) );
  SDFFX1 DFF_1334_Q_reg ( .D(g29621), .SI(g2387), .SE(n8253), .CLK(n8440), .Q(
        g2388), .QN(n7270) );
  SDFFX1 DFF_1335_Q_reg ( .D(g29623), .SI(g2388), .SE(n8253), .CLK(n8440), .Q(
        g2389), .QN(n7281) );
  SDFFX1 DFF_1336_Q_reg ( .D(g30707), .SI(g2389), .SE(n8253), .CLK(n8440), .Q(
        g2390), .QN(n7280) );
  SDFFX1 DFF_1337_Q_reg ( .D(g30709), .SI(g2390), .SE(n8247), .CLK(n8434), .Q(
        g2391), .QN(n7269) );
  SDFFX1 DFF_1338_Q_reg ( .D(g30566), .SI(g2391), .SE(n8248), .CLK(n8435), .Q(
        g2392), .QN(n7279) );
  SDFFX1 DFF_1339_Q_reg ( .D(g30505), .SI(g2392), .SE(n8247), .CLK(n8434), .Q(
        g2393), .QN(n7278) );
  SDFFX1 DFF_1340_Q_reg ( .D(g30341), .SI(g2393), .SE(n8248), .CLK(n8435), .Q(
        g2394), .QN(n7268) );
  SDFFX1 DFF_1341_Q_reg ( .D(g30356), .SI(g2394), .SE(n8248), .CLK(n8435), .Q(
        g2395), .QN(n7277) );
  SDFFX1 DFF_1342_Q_reg ( .D(g29182), .SI(g2395), .SE(n8261), .CLK(n8448), .Q(
        g2397), .QN(n7326) );
  SDFFX1 DFF_1343_Q_reg ( .D(g29185), .SI(g2397), .SE(n8261), .CLK(n8448), .Q(
        g2398), .QN(n7322) );
  SDFFX1 DFF_1344_Q_reg ( .D(g29187), .SI(g2398), .SE(n8261), .CLK(n8448), .Q(
        g2396), .QN(n7325) );
  SDFFX1 DFF_1345_Q_reg ( .D(g26672), .SI(g2396), .SE(n8261), .CLK(n8448), .Q(
        g2478), .QN(n7675) );
  SDFFX1 DFF_1346_Q_reg ( .D(g26676), .SI(g2478), .SE(n8261), .CLK(n8448), .Q(
        g2479), .QN(n7666) );
  SDFFX1 DFF_1347_Q_reg ( .D(g26025), .SI(g2479), .SE(n8261), .CLK(n8448), .Q(
        test_so82), .QN(n8128) );
  SDFFX1 DFF_1348_Q_reg ( .D(n4287), .SI(test_si83), .SE(n8153), .CLK(n8340), 
        .Q(g2525) );
  SDFFX1 DFF_1349_Q_reg ( .D(g2525), .SI(g2525), .SE(n8153), .CLK(n8340), .Q(
        n7946), .QN(DFF_1349_n1) );
  SDFFX1 DFF_1350_Q_reg ( .D(n4563), .SI(n7946), .SE(n8153), .CLK(n8340), .Q(
        g2527) );
  SDFFX1 DFF_1351_Q_reg ( .D(g2527), .SI(g2527), .SE(n8154), .CLK(n8341), .Q(
        n7945), .QN(DFF_1351_n1) );
  SDFFX1 DFF_1352_Q_reg ( .D(n4555), .SI(n7945), .SE(n8154), .CLK(n8341), .Q(
        g2529) );
  SDFFX1 DFF_1353_Q_reg ( .D(g2529), .SI(g2529), .SE(n8154), .CLK(n8341), .Q(
        n7944), .QN(DFF_1353_n1) );
  SDFFX1 DFF_1354_Q_reg ( .D(n4325), .SI(n7944), .SE(n8154), .CLK(n8341), .Q(
        g2355) );
  SDFFX1 DFF_1355_Q_reg ( .D(g2355), .SI(g2355), .SE(n8154), .CLK(n8341), .Q(
        n7943), .QN(DFF_1355_n1) );
  SDFFX1 DFF_1356_Q_reg ( .D(n4389), .SI(n7943), .SE(n8154), .CLK(n8341), .Q(
        g2357) );
  SDFFX1 DFF_1357_Q_reg ( .D(g2357), .SI(g2357), .SE(n8154), .CLK(n8341), .Q(
        n7942), .QN(DFF_1357_n1) );
  SDFFX1 DFF_1358_Q_reg ( .D(n4319), .SI(n7942), .SE(n8154), .CLK(n8341), .Q(
        g2359) );
  SDFFX1 DFF_1359_Q_reg ( .D(g2359), .SI(g2359), .SE(n8154), .CLK(n8341), .Q(
        n7941), .QN(DFF_1359_n1) );
  SDFFX1 DFF_1360_Q_reg ( .D(n4373), .SI(n7941), .SE(n8154), .CLK(n8341), .Q(
        g2361) );
  SDFFX1 DFF_1361_Q_reg ( .D(g2361), .SI(g2361), .SE(n8154), .CLK(n8341), .Q(
        n7940), .QN(DFF_1361_n1) );
  SDFFX1 DFF_1362_Q_reg ( .D(n4377), .SI(n7940), .SE(n8154), .CLK(n8341), .Q(
        test_so83) );
  SDFFX1 DFF_1363_Q_reg ( .D(test_so83), .SI(test_si84), .SE(n8155), .CLK(
        n8342), .Q(n7938), .QN(DFF_1363_n1) );
  SDFFX1 DFF_1364_Q_reg ( .D(g2878), .SI(n7938), .SE(n8170), .CLK(n8357), .Q(
        g2365) );
  SDFFX1 DFF_1365_Q_reg ( .D(g2365), .SI(g2365), .SE(n8170), .CLK(n8357), .Q(
        n7937), .QN(n4483) );
  SDFFX1 DFF_1366_Q_reg ( .D(n4285), .SI(n7937), .SE(n8259), .CLK(n8446), .Q(
        g2374), .QN(n4487) );
  SDFFX1 DFF_1367_Q_reg ( .D(g30055), .SI(g2374), .SE(n8264), .CLK(n8451), .Q(
        g2380) );
  SDFFX1 DFF_1378_Q_reg ( .D(n4275), .SI(g2380), .SE(n8261), .CLK(n8448), .Q(
        n7936), .QN(DFF_1378_n1) );
  SDFFX1 DFF_1379_Q_reg ( .D(g2429), .SI(n7936), .SE(n8261), .CLK(n8448), .Q(
        g2417) );
  SDFFX1 DFF_1380_Q_reg ( .D(g2417), .SI(g2417), .SE(n8262), .CLK(n8449), .Q(
        g2424) );
  SDFFX1 DFF_1381_Q_reg ( .D(g2418), .SI(g2424), .SE(n8262), .CLK(n8449), .Q(
        g2425) );
  SDFFX1 DFF_1382_Q_reg ( .D(g2425), .SI(g2425), .SE(n8262), .CLK(n8449), .Q(
        g2426) );
  SDFFX1 DFF_1383_Q_reg ( .D(g2421), .SI(g2426), .SE(n8262), .CLK(n8449), .Q(
        g2427) );
  SDFFX1 DFF_1384_Q_reg ( .D(g2427), .SI(g2427), .SE(n8262), .CLK(n8449), .Q(
        g2428) );
  SDFFX1 DFF_1385_Q_reg ( .D(g2444), .SI(g2428), .SE(n8262), .CLK(n8449), .Q(
        g2432) );
  SDFFX1 DFF_1386_Q_reg ( .D(g2432), .SI(g2432), .SE(n8262), .CLK(n8449), .Q(
        g2439) );
  SDFFX1 DFF_1387_Q_reg ( .D(g2433), .SI(g2439), .SE(n8262), .CLK(n8449), .Q(
        test_so84) );
  SDFFX1 DFF_1388_Q_reg ( .D(test_so84), .SI(test_si85), .SE(n8262), .CLK(
        n8449), .Q(g2441) );
  SDFFX1 DFF_1389_Q_reg ( .D(g2436), .SI(g2441), .SE(n8262), .CLK(n8449), .Q(
        g2442) );
  SDFFX1 DFF_1390_Q_reg ( .D(g2442), .SI(g2442), .SE(n8262), .CLK(n8449), .Q(
        g2443) );
  SDFFX1 DFF_1391_Q_reg ( .D(g2459), .SI(g2443), .SE(n8262), .CLK(n8449), .Q(
        g2447) );
  SDFFX1 DFF_1392_Q_reg ( .D(g2447), .SI(g2447), .SE(n8263), .CLK(n8450), .Q(
        g2454) );
  SDFFX1 DFF_1393_Q_reg ( .D(g2448), .SI(g2454), .SE(n8263), .CLK(n8450), .Q(
        g2455) );
  SDFFX1 DFF_1394_Q_reg ( .D(g2455), .SI(g2455), .SE(n8263), .CLK(n8450), .Q(
        g2456) );
  SDFFX1 DFF_1395_Q_reg ( .D(g2451), .SI(g2456), .SE(n8263), .CLK(n8450), .Q(
        g2457) );
  SDFFX1 DFF_1396_Q_reg ( .D(g2457), .SI(g2457), .SE(n8263), .CLK(n8450), .Q(
        g2458) );
  SDFFX1 DFF_1397_Q_reg ( .D(g2473), .SI(g2458), .SE(n8263), .CLK(n8450), .Q(
        g2462) );
  SDFFX1 DFF_1398_Q_reg ( .D(g2462), .SI(g2462), .SE(n8263), .CLK(n8450), .Q(
        g2469) );
  SDFFX1 DFF_1399_Q_reg ( .D(g2463), .SI(g2469), .SE(n8263), .CLK(n8450), .Q(
        g2470) );
  SDFFX1 DFF_1400_Q_reg ( .D(g2470), .SI(g2470), .SE(n8263), .CLK(n8450), .Q(
        g2471) );
  SDFFX1 DFF_1401_Q_reg ( .D(g2466), .SI(g2471), .SE(n8263), .CLK(n8450), .Q(
        g2472) );
  SDFFX1 DFF_1402_Q_reg ( .D(g2472), .SI(g2472), .SE(n8263), .CLK(n8450), .Q(
        test_so85) );
  SDFFX1 DFF_1403_Q_reg ( .D(n4598), .SI(test_si86), .SE(n8177), .CLK(n8364), 
        .Q(g5747) );
  SDFFX1 DFF_1404_Q_reg ( .D(g5747), .SI(g5747), .SE(n8177), .CLK(n8364), .Q(
        g5796) );
  SDFFX1 DFF_1405_Q_reg ( .D(g5796), .SI(g5796), .SE(n8177), .CLK(n8364), .Q(
        g2412) );
  SDFFX1 DFF_1406_Q_reg ( .D(n4598), .SI(g2412), .SE(n8177), .CLK(n8364), .Q(
        g7302), .QN(n4314) );
  SDFFX1 DFF_1407_Q_reg ( .D(g7302), .SI(g7302), .SE(n8177), .CLK(n8364), .Q(
        g7390), .QN(n4370) );
  SDFFX1 DFF_1408_Q_reg ( .D(g7390), .SI(g7390), .SE(n8177), .CLK(n8364), .Q(
        g2624), .QN(n4299) );
  SDFFX1 DFF_1409_Q_reg ( .D(n1431), .SI(g2624), .SE(n8178), .CLK(n8365), .Q(
        g2628), .QN(n7990) );
  SDFFX1 DFF_1410_Q_reg ( .D(g18780), .SI(g2628), .SE(n8178), .CLK(n8365), .Q(
        g2631), .QN(n4352) );
  SDFFX1 DFF_1411_Q_reg ( .D(g18820), .SI(g2631), .SE(n8178), .CLK(n8365), .Q(
        g2584), .QN(n4303) );
  SDFFX1 DFF_1412_Q_reg ( .D(n1427), .SI(g2584), .SE(n8256), .CLK(n8443), .Q(
        g2587) );
  SDFFX1 DFF_1413_Q_reg ( .D(g2587), .SI(g2587), .SE(n8256), .CLK(n8443), .Q(
        g2597) );
  SDFFX1 DFF_1414_Q_reg ( .D(g2597), .SI(g2597), .SE(n8256), .CLK(n8443), .Q(
        g2598) );
  SDFFX1 DFF_1415_Q_reg ( .D(g2530), .SI(g2598), .SE(n8256), .CLK(n8443), .Q(
        g2638) );
  SDFFX1 DFF_1416_Q_reg ( .D(g2638), .SI(g2638), .SE(n8256), .CLK(n8443), .Q(
        g2643) );
  SDFFX1 DFF_1417_Q_reg ( .D(g2533), .SI(g2643), .SE(n8256), .CLK(n8443), .Q(
        test_so86) );
  SDFFX1 DFF_1418_Q_reg ( .D(test_so86), .SI(test_si87), .SE(n8256), .CLK(
        n8443), .Q(g2645) );
  SDFFX1 DFF_1419_Q_reg ( .D(g2536), .SI(g2645), .SE(n8256), .CLK(n8443), .Q(
        g2646) );
  SDFFX1 DFF_1420_Q_reg ( .D(g2646), .SI(g2646), .SE(n8256), .CLK(n8443), .Q(
        g2647) );
  SDFFX1 DFF_1421_Q_reg ( .D(g2540), .SI(g2647), .SE(n8254), .CLK(n8441), .Q(
        g2648) );
  SDFFX1 DFF_1422_Q_reg ( .D(g2648), .SI(g2648), .SE(n8254), .CLK(n8441), .Q(
        g2639) );
  SDFFX1 DFF_1423_Q_reg ( .D(g2543), .SI(g2639), .SE(n8254), .CLK(n8441), .Q(
        g2640) );
  SDFFX1 DFF_1424_Q_reg ( .D(g2640), .SI(g2640), .SE(n8254), .CLK(n8441), .Q(
        g2641) );
  SDFFX1 DFF_1425_Q_reg ( .D(g2546), .SI(g2641), .SE(n8254), .CLK(n8441), .Q(
        g2642) );
  SDFFX1 DFF_1426_Q_reg ( .D(g2642), .SI(g2642), .SE(n8254), .CLK(n8441), .Q(
        g2564) );
  SDFFX1 DFF_1427_Q_reg ( .D(g2950), .SI(g2564), .SE(n8254), .CLK(n8441), .Q(
        g8087), .QN(n4456) );
  SDFFX1 DFF_1428_Q_reg ( .D(g8087), .SI(g8087), .SE(n8255), .CLK(n8442), .Q(
        g8167), .QN(n4455) );
  SDFFX1 DFF_1429_Q_reg ( .D(g8167), .SI(g8167), .SE(n8255), .CLK(n8442), .Q(
        g2560), .QN(n4463) );
  SDFFX1 DFF_1430_Q_reg ( .D(g23114), .SI(g2560), .SE(n8255), .CLK(n8442), .Q(
        g2561) );
  SDFFX1 DFF_1431_Q_reg ( .D(g23133), .SI(g2561), .SE(n8146), .CLK(n8333), .Q(
        g2562) );
  SDFFX1 DFF_1432_Q_reg ( .D(g21970), .SI(g2562), .SE(n8255), .CLK(n8442), .Q(
        test_so87) );
  SDFFX1 DFF_1433_Q_reg ( .D(g23407), .SI(test_si88), .SE(n8255), .CLK(n8442), 
        .Q(g2530) );
  SDFFX1 DFF_1434_Q_reg ( .D(g23418), .SI(g2530), .SE(n8255), .CLK(n8442), .Q(
        g2533) );
  SDFFX1 DFF_1435_Q_reg ( .D(g24209), .SI(g2533), .SE(n8255), .CLK(n8442), .Q(
        g2536) );
  SDFFX1 DFF_1436_Q_reg ( .D(g24214), .SI(g2536), .SE(n8257), .CLK(n8444), .Q(
        g2552) );
  SDFFX1 DFF_1437_Q_reg ( .D(g24226), .SI(g2552), .SE(n8257), .CLK(n8444), .Q(
        g2553) );
  SDFFX1 DFF_1438_Q_reg ( .D(g24238), .SI(g2553), .SE(n8257), .CLK(n8444), .Q(
        g2554) );
  SDFFX1 DFF_1439_Q_reg ( .D(g23132), .SI(g2554), .SE(n8254), .CLK(n8441), .Q(
        g2555) );
  SDFFX1 DFF_1440_Q_reg ( .D(g23047), .SI(g2555), .SE(n8254), .CLK(n8441), .Q(
        g2559) );
  SDFFX1 DFF_1441_Q_reg ( .D(g23076), .SI(g2559), .SE(n8254), .CLK(n8441), .Q(
        g2539) );
  SDFFX1 DFF_1442_Q_reg ( .D(g24225), .SI(g2539), .SE(n8254), .CLK(n8441), .Q(
        g2540) );
  SDFFX1 DFF_1443_Q_reg ( .D(g24237), .SI(g2540), .SE(n8255), .CLK(n8442), .Q(
        g2543) );
  SDFFX1 DFF_1444_Q_reg ( .D(g24250), .SI(g2543), .SE(n8255), .CLK(n8442), .Q(
        g2546) );
  SDFFX1 DFF_1445_Q_reg ( .D(n1406), .SI(g2546), .SE(n8255), .CLK(n8442), .Q(
        g2602) );
  SDFFX1 DFF_1446_Q_reg ( .D(g2602), .SI(g2602), .SE(n8255), .CLK(n8442), .Q(
        g2609) );
  SDFFX1 DFF_1447_Q_reg ( .D(g2609), .SI(g2609), .SE(n8255), .CLK(n8442), .Q(
        test_so88) );
  SDFFX1 DFF_1448_Q_reg ( .D(g13175), .SI(test_si89), .SE(n8257), .CLK(n8444), 
        .Q(g2617) );
  SDFFX1 DFF_1449_Q_reg ( .D(g2617), .SI(g2617), .SE(n8257), .CLK(n8444), .Q(
        n7930) );
  SDFFX1 DFF_1450_Q_reg ( .D(g30072), .SI(n7930), .SE(n8258), .CLK(n8445), .Q(
        n7929) );
  SDFFX1 DFF_1451_Q_reg ( .D(g13143), .SI(n7929), .SE(n8257), .CLK(n8444), .Q(
        g2623) );
  SDFFX1 DFF_1452_Q_reg ( .D(g2623), .SI(g2623), .SE(n8257), .CLK(n8444), .Q(
        g2574), .QN(n4543) );
  SDFFX1 DFF_1453_Q_reg ( .D(g13194), .SI(g2574), .SE(n8146), .CLK(n8333), .Q(
        g2632) );
  SDFFX1 DFF_1454_Q_reg ( .D(g2632), .SI(g2632), .SE(n8146), .CLK(n8333), .Q(
        g2633), .QN(n7761) );
  SDFFX1 DFF_1455_Q_reg ( .D(g27310), .SI(g2633), .SE(n8178), .CLK(n8365), .Q(
        g2650), .QN(n7338) );
  SDFFX1 DFF_1456_Q_reg ( .D(g27325), .SI(g2650), .SE(n8178), .CLK(n8365), .Q(
        g2651), .QN(n7340) );
  SDFFX1 DFF_1457_Q_reg ( .D(g27336), .SI(g2651), .SE(n8178), .CLK(n8365), .Q(
        g2649), .QN(n7339) );
  SDFFX1 DFF_1458_Q_reg ( .D(g27326), .SI(g2649), .SE(n8178), .CLK(n8365), .Q(
        g2653), .QN(n7350) );
  SDFFX1 DFF_1459_Q_reg ( .D(g27337), .SI(g2653), .SE(n8178), .CLK(n8365), .Q(
        g2654), .QN(n7352) );
  SDFFX1 DFF_1460_Q_reg ( .D(g27343), .SI(g2654), .SE(n8179), .CLK(n8366), .Q(
        g2652), .QN(n7351) );
  SDFFX1 DFF_1461_Q_reg ( .D(g27338), .SI(g2652), .SE(n8179), .CLK(n8366), .Q(
        g2656), .QN(n7177) );
  SDFFX1 DFF_1462_Q_reg ( .D(g27344), .SI(g2656), .SE(n8179), .CLK(n8366), .Q(
        test_so89), .QN(n8119) );
  SDFFX1 DFF_1463_Q_reg ( .D(g27347), .SI(test_si90), .SE(n8178), .CLK(n8365), 
        .Q(g2655), .QN(n7178) );
  SDFFX1 DFF_1464_Q_reg ( .D(g27345), .SI(g2655), .SE(n8178), .CLK(n8365), .Q(
        g2659), .QN(n7361) );
  SDFFX1 DFF_1465_Q_reg ( .D(g27348), .SI(g2659), .SE(n8178), .CLK(n8365), .Q(
        g2660), .QN(n7363) );
  SDFFX1 DFF_1466_Q_reg ( .D(g27354), .SI(g2660), .SE(n8178), .CLK(n8365), .Q(
        g2658), .QN(n7362) );
  SDFFX1 DFF_1467_Q_reg ( .D(g24527), .SI(g2658), .SE(n8256), .CLK(n8443), .Q(
        g2661) );
  SDFFX1 DFF_1468_Q_reg ( .D(g24537), .SI(g2661), .SE(n8256), .CLK(n8443), .Q(
        g2664) );
  SDFFX1 DFF_1469_Q_reg ( .D(g24547), .SI(g2664), .SE(n8256), .CLK(n8443), .Q(
        g2667) );
  SDFFX1 DFF_1470_Q_reg ( .D(g24538), .SI(g2667), .SE(n8257), .CLK(n8444), .Q(
        g2670) );
  SDFFX1 DFF_1471_Q_reg ( .D(g24548), .SI(g2670), .SE(n8257), .CLK(n8444), .Q(
        g2673) );
  SDFFX1 DFF_1472_Q_reg ( .D(g24557), .SI(g2673), .SE(n8257), .CLK(n8444), .Q(
        g2676) );
  SDFFX1 DFF_1473_Q_reg ( .D(g28364), .SI(g2676), .SE(n8257), .CLK(n8444), .Q(
        g2688) );
  SDFFX1 DFF_1474_Q_reg ( .D(g28368), .SI(g2688), .SE(n8257), .CLK(n8444), .Q(
        g2691) );
  SDFFX1 DFF_1475_Q_reg ( .D(g28371), .SI(g2691), .SE(n8170), .CLK(n8357), .Q(
        g2694) );
  SDFFX1 DFF_1476_Q_reg ( .D(g28358), .SI(g2694), .SE(n8263), .CLK(n8450), .Q(
        g2679) );
  SDFFX1 DFF_1477_Q_reg ( .D(g28363), .SI(g2679), .SE(n8264), .CLK(n8451), .Q(
        test_so90) );
  SDFFX1 DFF_1478_Q_reg ( .D(g28367), .SI(test_si91), .SE(n8264), .CLK(n8451), 
        .Q(g2685) );
  SDFFX1 DFF_1479_Q_reg ( .D(g26575), .SI(g2685), .SE(n8264), .CLK(n8451), .Q(
        g2565) );
  SDFFX1 DFF_1480_Q_reg ( .D(g26596), .SI(g2565), .SE(n8264), .CLK(n8451), .Q(
        g2568) );
  SDFFX1 DFF_1481_Q_reg ( .D(g26616), .SI(g2568), .SE(n8171), .CLK(n8358), .Q(
        g2571) );
  SDFFX1 DFF_1482_Q_reg ( .D(g2574), .SI(g2571), .SE(n8258), .CLK(n8445), .Q(
        g2580), .QN(n7501) );
  SDFFX1 DFF_1483_Q_reg ( .D(g22687), .SI(g2580), .SE(n8171), .CLK(n8358), .Q(
        n7926) );
  SDFFX1 DFF_1492_Q_reg ( .D(g30061), .SI(n7926), .SE(n8171), .CLK(n8358), .Q(
        g16437) );
  SDFFX1 DFF_1493_Q_reg ( .D(g16437), .SI(g16437), .SE(n8171), .CLK(n8358), 
        .Q(g2599), .QN(n8067) );
  SDFFX1 DFF_1494_Q_reg ( .D(DFF_1349_n1), .SI(g2599), .SE(n8171), .CLK(n8358), 
        .Q(n7925), .QN(DFF_1494_n1) );
  SDFFX1 DFF_1495_Q_reg ( .D(DFF_1351_n1), .SI(n7925), .SE(n8171), .CLK(n8358), 
        .Q(n7924), .QN(DFF_1495_n1) );
  SDFFX1 DFF_1496_Q_reg ( .D(DFF_1353_n1), .SI(n7924), .SE(n8171), .CLK(n8358), 
        .Q(n7923), .QN(DFF_1496_n1) );
  SDFFX1 DFF_1497_Q_reg ( .D(DFF_1355_n1), .SI(n7923), .SE(n8171), .CLK(n8358), 
        .Q(n7922), .QN(DFF_1497_n1) );
  SDFFX1 DFF_1498_Q_reg ( .D(DFF_1357_n1), .SI(n7922), .SE(n8171), .CLK(n8358), 
        .Q(n7921), .QN(DFF_1498_n1) );
  SDFFX1 DFF_1499_Q_reg ( .D(DFF_1359_n1), .SI(n7921), .SE(n8171), .CLK(n8358), 
        .Q(n7920), .QN(DFF_1499_n1) );
  SDFFX1 DFF_1500_Q_reg ( .D(DFF_1361_n1), .SI(n7920), .SE(n8171), .CLK(n8358), 
        .Q(test_so91), .QN(n7157) );
  SDFFX1 DFF_1501_Q_reg ( .D(DFF_1363_n1), .SI(test_si92), .SE(n8155), .CLK(
        n8342), .Q(g2611), .QN(n7156) );
  SDFFX1 DFF_1502_Q_reg ( .D(g24092), .SI(g2611), .SE(n8264), .CLK(n8451), .Q(
        g2612), .QN(n4490) );
  SDFFX1 DFF_1503_Q_reg ( .D(n4483), .SI(g2612), .SE(n8170), .CLK(n8357), .Q(
        n7918), .QN(n14379) );
  SDFFX1 DFF_1505_Q_reg ( .D(g7425), .SI(g7425), .SE(n8179), .CLK(n8366), .Q(
        g7487) );
  SDFFX1 DFF_1506_Q_reg ( .D(g7487), .SI(g7487), .SE(n8179), .CLK(n8366), .Q(
        g2703), .QN(n4292) );
  SDFFX1 DFF_1507_Q_reg ( .D(g16718), .SI(g2703), .SE(n8179), .CLK(n8366), .Q(
        g2704), .QN(n7757) );
  SDFFX1 DFF_1508_Q_reg ( .D(g20375), .SI(g2704), .SE(n8181), .CLK(n8368), .Q(
        g2733), .QN(n4426) );
  SDFFX1 DFF_1509_Q_reg ( .D(g20789), .SI(g2733), .SE(n8181), .CLK(n8368), .Q(
        g2714), .QN(n4398) );
  SDFFX1 DFF_1510_Q_reg ( .D(n1506), .SI(g2714), .SE(n8181), .CLK(n8368), .Q(
        g2707), .QN(n4472) );
  SDFFX1 DFF_1511_Q_reg ( .D(g23348), .SI(g2707), .SE(n8181), .CLK(n8368), .Q(
        g2727), .QN(n4419) );
  SDFFX1 DFF_1512_Q_reg ( .D(g24438), .SI(g2727), .SE(n8181), .CLK(n8368), .Q(
        g2720), .QN(n4408) );
  SDFFX1 DFF_1513_Q_reg ( .D(g25197), .SI(g2720), .SE(n8181), .CLK(n8368), .Q(
        g2734), .QN(n4397) );
  SDFFX1 DFF_1514_Q_reg ( .D(n1507), .SI(g2734), .SE(n8181), .CLK(n8368), .Q(
        g2746), .QN(n4407) );
  SDFFX1 DFF_1515_Q_reg ( .D(g26795), .SI(g2746), .SE(n8182), .CLK(n8369), .Q(
        test_so92), .QN(n8101) );
  SDFFX1 DFF_1516_Q_reg ( .D(g27243), .SI(test_si93), .SE(n8182), .CLK(n8369), 
        .Q(g2753), .QN(n4471) );
  SDFFX1 DFF_1517_Q_reg ( .D(g27724), .SI(g2753), .SE(n8182), .CLK(n8369), .Q(
        g2760), .QN(n4393) );
  SDFFX1 DFF_1518_Q_reg ( .D(g28328), .SI(g2760), .SE(n8182), .CLK(n8369), .Q(
        g2766), .QN(n4415) );
  SDFFX1 DFF_1519_Q_reg ( .D(g20918), .SI(g2766), .SE(n8182), .CLK(n8369), .Q(
        g2773), .QN(n7784) );
  SDFFX1 DFF_1520_Q_reg ( .D(g20939), .SI(g2773), .SE(n8182), .CLK(n8369), .Q(
        g2774), .QN(n7783) );
  SDFFX1 DFF_1521_Q_reg ( .D(g20962), .SI(g2774), .SE(n8182), .CLK(n8369), .Q(
        g2772), .QN(n7846) );
  SDFFX1 DFF_1522_Q_reg ( .D(g20940), .SI(g2772), .SE(n8184), .CLK(n8371), .Q(
        g2776), .QN(n7782) );
  SDFFX1 DFF_1523_Q_reg ( .D(g20963), .SI(g2776), .SE(n8184), .CLK(n8371), .Q(
        g2777), .QN(n7781) );
  SDFFX1 DFF_1524_Q_reg ( .D(g20981), .SI(g2777), .SE(n8184), .CLK(n8371), .Q(
        g2775), .QN(n7845) );
  SDFFX1 DFF_1525_Q_reg ( .D(g20964), .SI(g2775), .SE(n8184), .CLK(n8371), .Q(
        g2779), .QN(n7780) );
  SDFFX1 DFF_1526_Q_reg ( .D(g20982), .SI(g2779), .SE(n8184), .CLK(n8371), .Q(
        g2780), .QN(n7779) );
  SDFFX1 DFF_1527_Q_reg ( .D(g21004), .SI(g2780), .SE(n8184), .CLK(n8371), .Q(
        g2778), .QN(n7844) );
  SDFFX1 DFF_1528_Q_reg ( .D(g20983), .SI(g2778), .SE(n8184), .CLK(n8371), .Q(
        g2782), .QN(n7778) );
  SDFFX1 DFF_1529_Q_reg ( .D(g21005), .SI(g2782), .SE(n8184), .CLK(n8371), .Q(
        g2783), .QN(n7777) );
  SDFFX1 DFF_1530_Q_reg ( .D(g21025), .SI(g2783), .SE(n8184), .CLK(n8371), .Q(
        test_so93), .QN(n8131) );
  SDFFX1 DFF_1531_Q_reg ( .D(g21006), .SI(test_si94), .SE(n8181), .CLK(n8368), 
        .Q(g2785), .QN(n7776) );
  SDFFX1 DFF_1532_Q_reg ( .D(g21026), .SI(g2785), .SE(n8181), .CLK(n8368), .Q(
        g2786), .QN(n7775) );
  SDFFX1 DFF_1533_Q_reg ( .D(g21043), .SI(g2786), .SE(n8181), .CLK(n8368), .Q(
        g2784), .QN(n7843) );
  SDFFX1 DFF_1534_Q_reg ( .D(g21027), .SI(g2784), .SE(n8183), .CLK(n8370), .Q(
        g2788), .QN(n7774) );
  SDFFX1 DFF_1535_Q_reg ( .D(g21044), .SI(g2788), .SE(n8183), .CLK(n8370), .Q(
        g2789), .QN(n7773) );
  SDFFX1 DFF_1536_Q_reg ( .D(g21060), .SI(g2789), .SE(n8183), .CLK(n8370), .Q(
        g2787), .QN(n7842) );
  SDFFX1 DFF_1537_Q_reg ( .D(g21045), .SI(g2787), .SE(n8183), .CLK(n8370), .Q(
        g2791), .QN(n7772) );
  SDFFX1 DFF_1538_Q_reg ( .D(g21061), .SI(g2791), .SE(n8183), .CLK(n8370), .Q(
        g2792), .QN(n7771) );
  SDFFX1 DFF_1539_Q_reg ( .D(g21073), .SI(g2792), .SE(n8183), .CLK(n8370), .Q(
        g2790), .QN(n7841) );
  SDFFX1 DFF_1540_Q_reg ( .D(g21062), .SI(g2790), .SE(n8183), .CLK(n8370), .Q(
        g2794), .QN(n7770) );
  SDFFX1 DFF_1541_Q_reg ( .D(g21074), .SI(g2794), .SE(n8183), .CLK(n8370), .Q(
        g2795), .QN(n7769) );
  SDFFX1 DFF_1542_Q_reg ( .D(g21081), .SI(g2795), .SE(n8183), .CLK(n8370), .Q(
        g2793), .QN(n7840) );
  SDFFX1 DFF_1543_Q_reg ( .D(g21075), .SI(g2793), .SE(n8183), .CLK(n8370), .Q(
        g2797), .QN(n7768) );
  SDFFX1 DFF_1544_Q_reg ( .D(g21082), .SI(g2797), .SE(n8183), .CLK(n8370), .Q(
        g2798), .QN(n7767) );
  SDFFX1 DFF_1545_Q_reg ( .D(g21094), .SI(g2798), .SE(n8184), .CLK(n8371), .Q(
        test_so94), .QN(n8132) );
  SDFFX1 DFF_1546_Q_reg ( .D(g20919), .SI(test_si95), .SE(n8182), .CLK(n8369), 
        .Q(g2800), .QN(n7766) );
  SDFFX1 DFF_1547_Q_reg ( .D(g20941), .SI(g2800), .SE(n8182), .CLK(n8369), .Q(
        g2801), .QN(n7765) );
  SDFFX1 DFF_1548_Q_reg ( .D(g20965), .SI(g2801), .SE(n8182), .CLK(n8369), .Q(
        g2799), .QN(n7839) );
  SDFFX1 DFF_1549_Q_reg ( .D(g21007), .SI(g2799), .SE(n8182), .CLK(n8369), .Q(
        g2803), .QN(n8042) );
  SDFFX1 DFF_1550_Q_reg ( .D(g21028), .SI(g2803), .SE(n8182), .CLK(n8369), .Q(
        g2804), .QN(n7568) );
  SDFFX1 DFF_1551_Q_reg ( .D(g21046), .SI(g2804), .SE(n8183), .CLK(n8370), .Q(
        g2802) );
  SDFFX1 DFF_1552_Q_reg ( .D(g21029), .SI(g2802), .SE(n8264), .CLK(n8451), .Q(
        g2806), .QN(n7575) );
  SDFFX1 DFF_1553_Q_reg ( .D(g21047), .SI(g2806), .SE(n8264), .CLK(n8451), .Q(
        g2807), .QN(n7567) );
  SDFFX1 DFF_1554_Q_reg ( .D(g21063), .SI(g2807), .SE(n8264), .CLK(n8451), .Q(
        g2805), .QN(n7625) );
  SDFFX1 DFF_1555_Q_reg ( .D(g25272), .SI(g2805), .SE(n8264), .CLK(n8451), .Q(
        g2809), .QN(n7503) );
  SDFFX1 DFF_1556_Q_reg ( .D(g25280), .SI(g2809), .SE(n8264), .CLK(n8451), .Q(
        g2810), .QN(n7502) );
  SDFFX1 DFF_1557_Q_reg ( .D(g25288), .SI(g2810), .SE(n8171), .CLK(n8358), .Q(
        g2808), .QN(n7510) );
  SDFFX1 DFF_1558_Q_reg ( .D(g22269), .SI(g2808), .SE(n8172), .CLK(n8359), .Q(
        g2812), .QN(n7877) );
  SDFFX1 DFF_1559_Q_reg ( .D(g22284), .SI(g2812), .SE(n8181), .CLK(n8368), .Q(
        g2813), .QN(n7974) );
  SDFFX1 DFF_1560_Q_reg ( .D(g22299), .SI(g2813), .SE(n8181), .CLK(n8368), .Q(
        test_so95), .QN(n8116) );
  SDFFX1 DFF_1561_Q_reg ( .D(g20877), .SI(test_si96), .SE(n8172), .CLK(n8359), 
        .Q(n7913), .QN(DFF_1561_n1) );
  SDFFX1 DFF_1562_Q_reg ( .D(g20884), .SI(n7913), .SE(n8172), .CLK(n8359), .Q(
        n7912), .QN(DFF_1562_n1) );
  SDFFX1 DFF_1563_Q_reg ( .D(n4263_Tj_Payload), .SI(n7912), .SE(n8172), .CLK(
        n8359), .Q(n4598), .QN(n8049) );
  SDFFX1 DFF_1564_Q_reg ( .D(n4269), .SI(n4598), .SE(n8211), .CLK(n8398), .Q(
        g3043) );
  SDFFX1 DFF_1565_Q_reg ( .D(n4268), .SI(g3043), .SE(n8211), .CLK(n8398), .Q(
        g3044) );
  SDFFX1 DFF_1566_Q_reg ( .D(n4267), .SI(g3044), .SE(n8211), .CLK(n8398), .Q(
        g3045) );
  SDFFX1 DFF_1567_Q_reg ( .D(n4266), .SI(g3045), .SE(n8211), .CLK(n8398), .Q(
        g3046) );
  SDFFX1 DFF_1568_Q_reg ( .D(n4265), .SI(g3046), .SE(n8211), .CLK(n8398), .Q(
        g3047) );
  SDFFX1 DFF_1569_Q_reg ( .D(n4272), .SI(g3047), .SE(n8211), .CLK(n8398), .Q(
        g3048) );
  SDFFX1 DFF_1570_Q_reg ( .D(n4271), .SI(g3048), .SE(n8211), .CLK(n8398), .Q(
        g3049) );
  SDFFX1 DFF_1571_Q_reg ( .D(n4270), .SI(g3049), .SE(n8211), .CLK(n8398), .Q(
        g3050) );
  SDFFX1 DFF_1572_Q_reg ( .D(n4259), .SI(g3050), .SE(n8211), .CLK(n8398), .Q(
        g3051) );
  SDFFX1 DFF_1573_Q_reg ( .D(n4236), .SI(g3051), .SE(n8239), .CLK(n8426), .Q(
        g3052) );
  SDFFX1 DFF_1574_Q_reg ( .D(n4239), .SI(g3052), .SE(n8239), .CLK(n8426), .Q(
        g3053) );
  SDFFX1 DFF_1575_Q_reg ( .D(n4237), .SI(g3053), .SE(n8239), .CLK(n8426), .Q(
        test_so96) );
  SDFFX1 DFF_1576_Q_reg ( .D(n4234), .SI(test_si97), .SE(n8239), .CLK(n8426), 
        .Q(g3056) );
  SDFFX1 DFF_1577_Q_reg ( .D(n4233), .SI(g3056), .SE(n8239), .CLK(n8426), .Q(
        g3057) );
  SDFFX1 DFF_1578_Q_reg ( .D(n4238), .SI(g3057), .SE(n8239), .CLK(n8426), .Q(
        g3058) );
  SDFFX1 DFF_1579_Q_reg ( .D(n4235), .SI(g3058), .SE(n8239), .CLK(n8426), .Q(
        g3059) );
  SDFFX1 DFF_1580_Q_reg ( .D(n4240), .SI(g3059), .SE(n8239), .CLK(n8426), .Q(
        g3060) );
  SDFFX1 DFF_1581_Q_reg ( .D(n4232), .SI(g3060), .SE(n8239), .CLK(n8426), .Q(
        g3061) );
  SDFFX1 DFF_1582_Q_reg ( .D(n4245), .SI(g3061), .SE(n8264), .CLK(n8451), .Q(
        g3062) );
  SDFFX1 DFF_1583_Q_reg ( .D(n4248), .SI(g3062), .SE(n8265), .CLK(n8452), .Q(
        g3063) );
  SDFFX1 DFF_1584_Q_reg ( .D(n4246), .SI(g3063), .SE(n8265), .CLK(n8452), .Q(
        g3064) );
  SDFFX1 DFF_1585_Q_reg ( .D(n4243), .SI(g3064), .SE(n8265), .CLK(n8452), .Q(
        g3065) );
  SDFFX1 DFF_1586_Q_reg ( .D(n4242), .SI(g3065), .SE(n8265), .CLK(n8452), .Q(
        g3066) );
  SDFFX1 DFF_1587_Q_reg ( .D(n4247), .SI(g3066), .SE(n8265), .CLK(n8452), .Q(
        g3067) );
  SDFFX1 DFF_1588_Q_reg ( .D(n4244), .SI(g3067), .SE(n8265), .CLK(n8452), .Q(
        g3068) );
  SDFFX1 DFF_1589_Q_reg ( .D(n4249), .SI(g3068), .SE(n8265), .CLK(n8452), .Q(
        g3069) );
  SDFFX1 DFF_1590_Q_reg ( .D(n4241), .SI(g3069), .SE(n8265), .CLK(n8452), .Q(
        test_so97) );
  SDFFX1 DFF_1591_Q_reg ( .D(n4254), .SI(test_si98), .SE(n8267), .CLK(n8454), 
        .Q(g3071) );
  SDFFX1 DFF_1592_Q_reg ( .D(n4257), .SI(g3071), .SE(n8267), .CLK(n8454), .Q(
        g3072) );
  SDFFX1 DFF_1593_Q_reg ( .D(n4255), .SI(g3072), .SE(n8267), .CLK(n8454), .Q(
        g3073) );
  SDFFX1 DFF_1594_Q_reg ( .D(n4252), .SI(g3073), .SE(n8267), .CLK(n8454), .Q(
        g3074) );
  SDFFX1 DFF_1595_Q_reg ( .D(n4251), .SI(g3074), .SE(n8267), .CLK(n8454), .Q(
        g3075) );
  SDFFX1 DFF_1596_Q_reg ( .D(n4256), .SI(g3075), .SE(n8268), .CLK(n8455), .Q(
        g3076) );
  SDFFX1 DFF_1597_Q_reg ( .D(n4253), .SI(g3076), .SE(n8268), .CLK(n8455), .Q(
        g3077) );
  SDFFX1 DFF_1598_Q_reg ( .D(n4258), .SI(g3077), .SE(n8268), .CLK(n8455), .Q(
        g3078) );
  SDFFX1 DFF_1599_Q_reg ( .D(n4250), .SI(g3078), .SE(n8170), .CLK(n8357), .Q(
        g2997) );
  SDFFX1 DFF_1600_Q_reg ( .D(g25265), .SI(g2997), .SE(n8170), .CLK(n8357), .Q(
        g2993), .QN(n8050) );
  SDFFX1 DFF_1601_Q_reg ( .D(g26048), .SI(g2993), .SE(n8179), .CLK(n8366), .Q(
        n7909), .QN(n14387) );
  SDFFX1 DFF_1602_Q_reg ( .D(n1542), .SI(n7909), .SE(n8179), .CLK(n8366), .Q(
        g3006), .QN(n8053) );
  SDFFX1 DFF_1603_Q_reg ( .D(g24445), .SI(g3006), .SE(n8179), .CLK(n8366), .Q(
        g3002), .QN(n8052) );
  SDFFX1 DFF_1604_Q_reg ( .D(g25191), .SI(g3002), .SE(n8179), .CLK(n8366), .Q(
        g3013), .QN(n8073) );
  SDFFX1 DFF_1605_Q_reg ( .D(g26031), .SI(g3013), .SE(n8179), .CLK(n8366), .Q(
        test_so98) );
  SDFFX1 DFF_1606_Q_reg ( .D(g26786), .SI(test_si99), .SE(n8180), .CLK(n8367), 
        .Q(g3024), .QN(n8051) );
  SDFFX1 DFF_1607_Q_reg ( .D(n4262), .SI(g3024), .SE(n8265), .CLK(n8452), .Q(
        g3018), .QN(n4481) );
  SDFFX1 DFF_1608_Q_reg ( .D(n1544), .SI(g3018), .SE(n8265), .CLK(n8452), .Q(
        g3028), .QN(n4350) );
  SDFFX1 DFF_1609_Q_reg ( .D(g24446), .SI(g3028), .SE(n8267), .CLK(n8454), .Q(
        g3036), .QN(n4480) );
  SDFFX1 DFF_1610_Q_reg ( .D(g25202), .SI(g3036), .SE(n8265), .CLK(n8452), .Q(
        g3032), .QN(n7441) );
  SDFFX1 DFF_1611_Q_reg ( .D(g3234), .SI(g3032), .SE(n8265), .CLK(n8452), .Q(
        g5388) );
  SDFFX1 DFF_1612_Q_reg ( .D(g5388), .SI(g5388), .SE(n8266), .CLK(n8453), .Q(
        n7907), .QN(DFF_1612_n1) );
  SDFFX1 DFF_1613_Q_reg ( .D(g16496), .SI(n7907), .SE(n8266), .CLK(n8453), .Q(
        g2987), .QN(n4365) );
  SDFFX1 DFF_1614_Q_reg ( .D(g16824), .SI(g2987), .SE(n8266), .CLK(n8453), .Q(
        g8275) );
  SDFFX1 DFF_1615_Q_reg ( .D(g16844), .SI(g8275), .SE(n8266), .CLK(n8453), .Q(
        g8274), .QN(n8030) );
  SDFFX1 DFF_1616_Q_reg ( .D(g16853), .SI(g8274), .SE(n8266), .CLK(n8453), .Q(
        g8273), .QN(n14391) );
  SDFFX1 DFF_1617_Q_reg ( .D(g16860), .SI(g8273), .SE(n8266), .CLK(n8453), .Q(
        g8272), .QN(n14390) );
  SDFFX1 DFF_1618_Q_reg ( .D(g16803), .SI(g8272), .SE(n8266), .CLK(n8453), .Q(
        g8268), .QN(n14389) );
  SDFFX1 DFF_1619_Q_reg ( .D(g16835), .SI(g8268), .SE(n8266), .CLK(n8453), .Q(
        g8269), .QN(n8031) );
  SDFFX1 DFF_1620_Q_reg ( .D(g16851), .SI(g8269), .SE(n8266), .CLK(n8453), .Q(
        test_so99) );
  SDFFX1 DFF_1621_Q_reg ( .D(g16857), .SI(test_si100), .SE(n8266), .CLK(n8453), 
        .Q(g8271), .QN(n8029) );
  SDFFX1 DFF_1622_Q_reg ( .D(g16866), .SI(g8271), .SE(n8266), .CLK(n8453), .Q(
        g3083), .QN(n8034) );
  SDFFX1 DFF_1623_Q_reg ( .D(n4261), .SI(g3083), .SE(n8266), .CLK(n8453), .Q(
        g8267) );
  SDFFX1 DFF_1624_Q_reg ( .D(N995), .SI(g8267), .SE(n8267), .CLK(n8454), .Q(
        n4577), .QN(n7444) );
  SDFFX1 DFF_1625_Q_reg ( .D(g16845), .SI(n4577), .SE(n8267), .CLK(n8454), .Q(
        g8266), .QN(n14394) );
  SDFFX1 DFF_1626_Q_reg ( .D(g16854), .SI(g8266), .SE(n8267), .CLK(n8454), .Q(
        g8265), .QN(n14393) );
  SDFFX1 DFF_1627_Q_reg ( .D(g16861), .SI(g8265), .SE(n8267), .CLK(n8454), .Q(
        g8264), .QN(n7996) );
  SDFFX1 DFF_1628_Q_reg ( .D(g16880), .SI(g8264), .SE(n8267), .CLK(n8454), .Q(
        g8262) );
  SDFFX1 DFF_1629_Q_reg ( .D(g18755), .SI(g8262), .SE(n8267), .CLK(n8454), .Q(
        g8263), .QN(n7997) );
  SDFFX1 DFF_1630_Q_reg ( .D(g18804), .SI(g8263), .SE(n8268), .CLK(n8455), .Q(
        g8260), .QN(n7994) );
  SDFFX1 DFF_1631_Q_reg ( .D(g18837), .SI(g8260), .SE(n8268), .CLK(n8455), .Q(
        g8261), .QN(n14392) );
  SDFFX1 DFF_1632_Q_reg ( .D(g18868), .SI(g8261), .SE(n8268), .CLK(n8455), .Q(
        g8259), .QN(n7995) );
  SDFFX1 DFF_1633_Q_reg ( .D(g18907), .SI(g8259), .SE(n8268), .CLK(n8455), .Q(
        g2990), .QN(n8032) );
  SDFFX1 DFF_1634_Q_reg ( .D(N690), .SI(g2990), .SE(n8268), .CLK(n8455), .Q(
        n4578), .QN(n7443) );
  SDFFX1 DFF_1635_Q_reg ( .D(n4260), .SI(n4578), .SE(n8268), .CLK(n8455), .Q(
        test_so100) );
  SDFFX1 DFF_454_Q_reg ( .D(n4598), .SI(n8040), .SE(n8172), .CLK(n8359), .Q(
        g6677), .QN(n4309) );
  SDFFX1 DFF_804_Q_reg ( .D(n4598), .SI(test_si49), .SE(n8172), .CLK(n8359), 
        .Q(g6979), .QN(n4308) );
  SDFFX1 DFF_1154_Q_reg ( .D(n4598), .SI(n7960), .SE(n8172), .CLK(n8359), .Q(
        g7229), .QN(n4307) );
  SDFFX1 DFF_1504_Q_reg ( .D(n4598), .SI(n7918), .SE(n8179), .CLK(n8366), .Q(
        g7425), .QN(n4306) );
  SDFFX1 DFF_1300_Q_reg ( .D(g5555), .SI(g5555), .SE(n8248), .CLK(n8435), .Q(
        g7264), .QN(n4524) );
  SDFFX1 DFF_950_Q_reg ( .D(g5511), .SI(g5511), .SE(n8222), .CLK(n8409), .Q(
        g7014), .QN(n4525) );
  SDFFX1 DFF_951_Q_reg ( .D(g7014), .SI(g7014), .SE(n8222), .CLK(n8409), .Q(
        n4618), .QN(n4511) );
  SDFFX1 DFF_1301_Q_reg ( .D(g7264), .SI(g7264), .SE(n8248), .CLK(n8435), .Q(
        n4606), .QN(n4509) );
  SDFFX1 DFF_250_Q_reg ( .D(g5437), .SI(g5437), .SE(n8157), .CLK(n8344), .Q(
        g6447), .QN(n4499) );
  SDFFX1 DFF_249_Q_reg ( .D(g2950), .SI(g181), .SE(n8157), .CLK(n8344), .Q(
        g5437), .QN(n4520) );
  NOR2X0 Trojan1 ( .IN1(n155), .IN2(n3016), .QN(Tj_OUT1) );
  NOR2X0 Trojan2 ( .IN1(n3023), .IN2(n3000), .QN(Tj_OUT2) );
  NOR2X0 Trojan3 ( .IN1(n3008), .IN2(n3068), .QN(Tj_OUT3) );
  NOR2X0 Trojan4 ( .IN1(n3128), .IN2(n3036), .QN(Tj_OUT4) );
  AND4X1 Trojan1234_NOT ( .IN1(Tj_OUT1), .IN2(Tj_OUT2), .IN3(Tj_OUT3), .IN4(
        Tj_OUT4), .Q(Tj_OUT1234) );
  NOR2X0 Trojan5 ( .IN1(n162), .IN2(n184), .QN(Tj_OUT5) );
  NOR2X0 Trojan6 ( .IN1(n123), .IN2(n223), .QN(Tj_OUT6) );
  NOR2X0 Trojan7 ( .IN1(n2792), .IN2(n2632), .QN(Tj_OUT7) );
  NOR2X0 Trojan8 ( .IN1(n2351), .IN2(n2430), .QN(Tj_OUT8) );
  AND4X1 Trojan5678_NOT ( .IN1(Tj_OUT5), .IN2(Tj_OUT6), .IN3(Tj_OUT7), .IN4(
        Tj_OUT8), .Q(Tj_OUT5678) );
  AND2X1 Trojan_CLK_NOT ( .IN1(Tj_OUT1234), .IN2(Tj_OUT5678), .Q(Tj_Trigger)
         );
  OR2X1 Trojan_Payload ( .IN1(Tj_Trigger), .IN2(n4263), .Q(n4263_Tj_Payload)
         );
  NBUFFX2 U7976 ( .INP(n8316), .Z(n8143) );
  NBUFFX2 U7977 ( .INP(n8316), .Z(n8142) );
  NBUFFX2 U7978 ( .INP(n8275), .Z(n8266) );
  NBUFFX2 U7979 ( .INP(n8274), .Z(n8267) );
  NBUFFX2 U7980 ( .INP(n8275), .Z(n8265) );
  NBUFFX2 U7981 ( .INP(n8302), .Z(n8183) );
  NBUFFX2 U7982 ( .INP(n8303), .Z(n8182) );
  NBUFFX2 U7983 ( .INP(n8303), .Z(n8181) );
  NBUFFX2 U7984 ( .INP(n8306), .Z(n8171) );
  NBUFFX2 U7985 ( .INP(n8304), .Z(n8179) );
  NBUFFX2 U7986 ( .INP(n8278), .Z(n8257) );
  NBUFFX2 U7987 ( .INP(n8278), .Z(n8255) );
  NBUFFX2 U7988 ( .INP(n8278), .Z(n8256) );
  NBUFFX2 U7989 ( .INP(n8304), .Z(n8178) );
  NBUFFX2 U7990 ( .INP(n8276), .Z(n8263) );
  NBUFFX2 U7991 ( .INP(n8276), .Z(n8262) );
  NBUFFX2 U7992 ( .INP(n8275), .Z(n8264) );
  NBUFFX2 U7993 ( .INP(n8312), .Z(n8154) );
  NBUFFX2 U7994 ( .INP(n8279), .Z(n8254) );
  NBUFFX2 U7995 ( .INP(n8277), .Z(n8258) );
  NBUFFX2 U7996 ( .INP(n8277), .Z(n8259) );
  NBUFFX2 U7997 ( .INP(n8281), .Z(n8248) );
  NBUFFX2 U7998 ( .INP(n8279), .Z(n8253) );
  NBUFFX2 U7999 ( .INP(n8276), .Z(n8261) );
  NBUFFX2 U8000 ( .INP(n8277), .Z(n8260) );
  NBUFFX2 U8001 ( .INP(n8280), .Z(n8250) );
  NBUFFX2 U8002 ( .INP(n8280), .Z(n8249) );
  NBUFFX2 U8003 ( .INP(n8279), .Z(n8252) );
  NBUFFX2 U8004 ( .INP(n8281), .Z(n8247) );
  NBUFFX2 U8005 ( .INP(n8280), .Z(n8251) );
  NBUFFX2 U8006 ( .INP(n8281), .Z(n8246) );
  NBUFFX2 U8007 ( .INP(n8282), .Z(n8245) );
  NBUFFX2 U8008 ( .INP(n8282), .Z(n8244) );
  NBUFFX2 U8009 ( .INP(n8282), .Z(n8243) );
  NBUFFX2 U8010 ( .INP(n8283), .Z(n8242) );
  NBUFFX2 U8011 ( .INP(n8283), .Z(n8241) );
  NBUFFX2 U8012 ( .INP(n8283), .Z(n8240) );
  NBUFFX2 U8013 ( .INP(n8284), .Z(n8239) );
  NBUFFX2 U8014 ( .INP(n8284), .Z(n8238) );
  NBUFFX2 U8015 ( .INP(n8284), .Z(n8237) );
  NBUFFX2 U8016 ( .INP(n8285), .Z(n8236) );
  NBUFFX2 U8017 ( .INP(n8285), .Z(n8235) );
  NBUFFX2 U8018 ( .INP(n8285), .Z(n8234) );
  NBUFFX2 U8019 ( .INP(n8286), .Z(n8233) );
  NBUFFX2 U8020 ( .INP(n8286), .Z(n8232) );
  NBUFFX2 U8021 ( .INP(n8288), .Z(n8227) );
  NBUFFX2 U8022 ( .INP(n8287), .Z(n8229) );
  NBUFFX2 U8023 ( .INP(n8287), .Z(n8228) );
  NBUFFX2 U8024 ( .INP(n8286), .Z(n8231) );
  NBUFFX2 U8025 ( .INP(n8287), .Z(n8230) );
  NBUFFX2 U8026 ( .INP(n8290), .Z(n8221) );
  NBUFFX2 U8027 ( .INP(n8290), .Z(n8220) );
  NBUFFX2 U8028 ( .INP(n8288), .Z(n8226) );
  NBUFFX2 U8029 ( .INP(n8289), .Z(n8222) );
  NBUFFX2 U8030 ( .INP(n8288), .Z(n8225) );
  NBUFFX2 U8031 ( .INP(n8289), .Z(n8224) );
  NBUFFX2 U8032 ( .INP(n8289), .Z(n8223) );
  NBUFFX2 U8033 ( .INP(n8290), .Z(n8219) );
  NBUFFX2 U8034 ( .INP(n8291), .Z(n8218) );
  NBUFFX2 U8035 ( .INP(n8291), .Z(n8217) );
  NBUFFX2 U8036 ( .INP(n8291), .Z(n8216) );
  NBUFFX2 U8037 ( .INP(n8292), .Z(n8215) );
  NBUFFX2 U8038 ( .INP(n8292), .Z(n8214) );
  NBUFFX2 U8039 ( .INP(n8292), .Z(n8213) );
  NBUFFX2 U8040 ( .INP(n8293), .Z(n8212) );
  NBUFFX2 U8041 ( .INP(n8293), .Z(n8211) );
  NBUFFX2 U8042 ( .INP(n8293), .Z(n8210) );
  NBUFFX2 U8043 ( .INP(n8294), .Z(n8209) );
  NBUFFX2 U8044 ( .INP(n8294), .Z(n8208) );
  NBUFFX2 U8045 ( .INP(n8294), .Z(n8207) );
  NBUFFX2 U8046 ( .INP(n8295), .Z(n8206) );
  NBUFFX2 U8047 ( .INP(n8295), .Z(n8205) );
  NBUFFX2 U8048 ( .INP(n8295), .Z(n8204) );
  NBUFFX2 U8049 ( .INP(n8296), .Z(n8201) );
  NBUFFX2 U8050 ( .INP(n8297), .Z(n8200) );
  NBUFFX2 U8051 ( .INP(n8296), .Z(n8202) );
  NBUFFX2 U8052 ( .INP(n8297), .Z(n8198) );
  NBUFFX2 U8053 ( .INP(n8299), .Z(n8193) );
  NBUFFX2 U8054 ( .INP(n8297), .Z(n8199) );
  NBUFFX2 U8055 ( .INP(n8296), .Z(n8203) );
  NBUFFX2 U8056 ( .INP(n8299), .Z(n8194) );
  NBUFFX2 U8057 ( .INP(n8298), .Z(n8197) );
  NBUFFX2 U8058 ( .INP(n8298), .Z(n8196) );
  NBUFFX2 U8059 ( .INP(n8298), .Z(n8195) );
  NBUFFX2 U8060 ( .INP(n8299), .Z(n8192) );
  NBUFFX2 U8061 ( .INP(n8300), .Z(n8191) );
  NBUFFX2 U8062 ( .INP(n8300), .Z(n8190) );
  NBUFFX2 U8063 ( .INP(n8300), .Z(n8189) );
  NBUFFX2 U8064 ( .INP(n8301), .Z(n8188) );
  NBUFFX2 U8065 ( .INP(n8303), .Z(n8180) );
  NBUFFX2 U8066 ( .INP(n8306), .Z(n8172) );
  NBUFFX2 U8067 ( .INP(n8301), .Z(n8187) );
  NBUFFX2 U8068 ( .INP(n8301), .Z(n8186) );
  NBUFFX2 U8069 ( .INP(n8302), .Z(n8185) );
  NBUFFX2 U8070 ( .INP(n8302), .Z(n8184) );
  NBUFFX2 U8071 ( .INP(n8304), .Z(n8177) );
  NBUFFX2 U8072 ( .INP(n8305), .Z(n8176) );
  NBUFFX2 U8073 ( .INP(n8305), .Z(n8175) );
  NBUFFX2 U8074 ( .INP(n8305), .Z(n8174) );
  NBUFFX2 U8075 ( .INP(n8306), .Z(n8173) );
  NBUFFX2 U8076 ( .INP(n8307), .Z(n8168) );
  NBUFFX2 U8077 ( .INP(n8312), .Z(n8155) );
  NBUFFX2 U8078 ( .INP(n8307), .Z(n8169) );
  NBUFFX2 U8079 ( .INP(n8308), .Z(n8165) );
  NBUFFX2 U8080 ( .INP(n8308), .Z(n8167) );
  NBUFFX2 U8081 ( .INP(n8308), .Z(n8166) );
  NBUFFX2 U8082 ( .INP(n8311), .Z(n8157) );
  NBUFFX2 U8083 ( .INP(n8309), .Z(n8162) );
  NBUFFX2 U8084 ( .INP(n8309), .Z(n8164) );
  NBUFFX2 U8085 ( .INP(n8309), .Z(n8163) );
  NBUFFX2 U8086 ( .INP(n8311), .Z(n8158) );
  NBUFFX2 U8087 ( .INP(n8311), .Z(n8156) );
  NBUFFX2 U8088 ( .INP(n8310), .Z(n8159) );
  NBUFFX2 U8089 ( .INP(n8310), .Z(n8161) );
  NBUFFX2 U8090 ( .INP(n8310), .Z(n8160) );
  NBUFFX2 U8091 ( .INP(n8314), .Z(n8148) );
  NBUFFX2 U8092 ( .INP(n8314), .Z(n8147) );
  NBUFFX2 U8093 ( .INP(n8273), .Z(n8270) );
  NBUFFX2 U8094 ( .INP(n8315), .Z(n8146) );
  NBUFFX2 U8095 ( .INP(n8273), .Z(n8271) );
  NBUFFX2 U8096 ( .INP(n8274), .Z(n8269) );
  NBUFFX2 U8097 ( .INP(n8274), .Z(n8268) );
  NBUFFX2 U8098 ( .INP(n8307), .Z(n8170) );
  NBUFFX2 U8099 ( .INP(n8312), .Z(n8153) );
  NBUFFX2 U8100 ( .INP(n8313), .Z(n8152) );
  NBUFFX2 U8101 ( .INP(n8313), .Z(n8151) );
  NBUFFX2 U8102 ( .INP(n8313), .Z(n8150) );
  NBUFFX2 U8103 ( .INP(n8314), .Z(n8149) );
  NBUFFX2 U8104 ( .INP(n8315), .Z(n8145) );
  NBUFFX2 U8105 ( .INP(n8315), .Z(n8144) );
  NBUFFX2 U8106 ( .INP(n8503), .Z(n8330) );
  NBUFFX2 U8107 ( .INP(n8503), .Z(n8329) );
  NBUFFX2 U8108 ( .INP(n8462), .Z(n8453) );
  NBUFFX2 U8109 ( .INP(n8461), .Z(n8454) );
  NBUFFX2 U8110 ( .INP(n8462), .Z(n8452) );
  NBUFFX2 U8111 ( .INP(n8489), .Z(n8370) );
  NBUFFX2 U8112 ( .INP(n8490), .Z(n8369) );
  NBUFFX2 U8113 ( .INP(n8490), .Z(n8368) );
  NBUFFX2 U8114 ( .INP(n8493), .Z(n8358) );
  NBUFFX2 U8115 ( .INP(n8491), .Z(n8366) );
  NBUFFX2 U8116 ( .INP(n8465), .Z(n8444) );
  NBUFFX2 U8117 ( .INP(n8465), .Z(n8442) );
  NBUFFX2 U8118 ( .INP(n8465), .Z(n8443) );
  NBUFFX2 U8119 ( .INP(n8491), .Z(n8365) );
  NBUFFX2 U8120 ( .INP(n8463), .Z(n8450) );
  NBUFFX2 U8121 ( .INP(n8463), .Z(n8449) );
  NBUFFX2 U8122 ( .INP(n8462), .Z(n8451) );
  NBUFFX2 U8123 ( .INP(n8499), .Z(n8341) );
  NBUFFX2 U8124 ( .INP(n8466), .Z(n8441) );
  NBUFFX2 U8125 ( .INP(n8464), .Z(n8445) );
  NBUFFX2 U8126 ( .INP(n8464), .Z(n8446) );
  NBUFFX2 U8127 ( .INP(n8468), .Z(n8435) );
  NBUFFX2 U8128 ( .INP(n8466), .Z(n8440) );
  NBUFFX2 U8129 ( .INP(n8463), .Z(n8448) );
  NBUFFX2 U8130 ( .INP(n8464), .Z(n8447) );
  NBUFFX2 U8131 ( .INP(n8467), .Z(n8437) );
  NBUFFX2 U8132 ( .INP(n8467), .Z(n8436) );
  NBUFFX2 U8133 ( .INP(n8466), .Z(n8439) );
  NBUFFX2 U8134 ( .INP(n8468), .Z(n8434) );
  NBUFFX2 U8135 ( .INP(n8467), .Z(n8438) );
  NBUFFX2 U8136 ( .INP(n8468), .Z(n8433) );
  NBUFFX2 U8137 ( .INP(n8469), .Z(n8432) );
  NBUFFX2 U8138 ( .INP(n8469), .Z(n8431) );
  NBUFFX2 U8139 ( .INP(n8469), .Z(n8430) );
  NBUFFX2 U8140 ( .INP(n8470), .Z(n8429) );
  NBUFFX2 U8141 ( .INP(n8470), .Z(n8428) );
  NBUFFX2 U8142 ( .INP(n8470), .Z(n8427) );
  NBUFFX2 U8143 ( .INP(n8471), .Z(n8426) );
  NBUFFX2 U8144 ( .INP(n8471), .Z(n8425) );
  NBUFFX2 U8145 ( .INP(n8471), .Z(n8424) );
  NBUFFX2 U8146 ( .INP(n8472), .Z(n8423) );
  NBUFFX2 U8147 ( .INP(n8472), .Z(n8422) );
  NBUFFX2 U8148 ( .INP(n8472), .Z(n8421) );
  NBUFFX2 U8149 ( .INP(n8473), .Z(n8420) );
  NBUFFX2 U8150 ( .INP(n8473), .Z(n8419) );
  NBUFFX2 U8151 ( .INP(n8475), .Z(n8414) );
  NBUFFX2 U8152 ( .INP(n8474), .Z(n8416) );
  NBUFFX2 U8153 ( .INP(n8474), .Z(n8415) );
  NBUFFX2 U8154 ( .INP(n8473), .Z(n8418) );
  NBUFFX2 U8155 ( .INP(n8474), .Z(n8417) );
  NBUFFX2 U8156 ( .INP(n8477), .Z(n8408) );
  NBUFFX2 U8157 ( .INP(n8477), .Z(n8407) );
  NBUFFX2 U8158 ( .INP(n8475), .Z(n8413) );
  NBUFFX2 U8159 ( .INP(n8476), .Z(n8409) );
  NBUFFX2 U8160 ( .INP(n8475), .Z(n8412) );
  NBUFFX2 U8161 ( .INP(n8476), .Z(n8411) );
  NBUFFX2 U8162 ( .INP(n8476), .Z(n8410) );
  NBUFFX2 U8163 ( .INP(n8477), .Z(n8406) );
  NBUFFX2 U8164 ( .INP(n8478), .Z(n8405) );
  NBUFFX2 U8165 ( .INP(n8478), .Z(n8404) );
  NBUFFX2 U8166 ( .INP(n8478), .Z(n8403) );
  NBUFFX2 U8167 ( .INP(n8479), .Z(n8402) );
  NBUFFX2 U8168 ( .INP(n8479), .Z(n8401) );
  NBUFFX2 U8169 ( .INP(n8479), .Z(n8400) );
  NBUFFX2 U8170 ( .INP(n8480), .Z(n8399) );
  NBUFFX2 U8171 ( .INP(n8480), .Z(n8398) );
  NBUFFX2 U8172 ( .INP(n8480), .Z(n8397) );
  NBUFFX2 U8173 ( .INP(n8481), .Z(n8396) );
  NBUFFX2 U8174 ( .INP(n8481), .Z(n8395) );
  NBUFFX2 U8175 ( .INP(n8481), .Z(n8394) );
  NBUFFX2 U8176 ( .INP(n8482), .Z(n8393) );
  NBUFFX2 U8177 ( .INP(n8482), .Z(n8392) );
  NBUFFX2 U8178 ( .INP(n8482), .Z(n8391) );
  NBUFFX2 U8179 ( .INP(n8483), .Z(n8388) );
  NBUFFX2 U8180 ( .INP(n8484), .Z(n8387) );
  NBUFFX2 U8181 ( .INP(n8483), .Z(n8389) );
  NBUFFX2 U8182 ( .INP(n8484), .Z(n8385) );
  NBUFFX2 U8183 ( .INP(n8486), .Z(n8380) );
  NBUFFX2 U8184 ( .INP(n8484), .Z(n8386) );
  NBUFFX2 U8185 ( .INP(n8483), .Z(n8390) );
  NBUFFX2 U8186 ( .INP(n8486), .Z(n8381) );
  NBUFFX2 U8187 ( .INP(n8485), .Z(n8384) );
  NBUFFX2 U8188 ( .INP(n8485), .Z(n8383) );
  NBUFFX2 U8189 ( .INP(n8485), .Z(n8382) );
  NBUFFX2 U8190 ( .INP(n8486), .Z(n8379) );
  NBUFFX2 U8191 ( .INP(n8487), .Z(n8378) );
  NBUFFX2 U8192 ( .INP(n8487), .Z(n8377) );
  NBUFFX2 U8193 ( .INP(n8487), .Z(n8376) );
  NBUFFX2 U8194 ( .INP(n8488), .Z(n8375) );
  NBUFFX2 U8195 ( .INP(n8490), .Z(n8367) );
  NBUFFX2 U8196 ( .INP(n8493), .Z(n8359) );
  NBUFFX2 U8197 ( .INP(n8488), .Z(n8374) );
  NBUFFX2 U8198 ( .INP(n8488), .Z(n8373) );
  NBUFFX2 U8199 ( .INP(n8489), .Z(n8372) );
  NBUFFX2 U8200 ( .INP(n8489), .Z(n8371) );
  NBUFFX2 U8201 ( .INP(n8491), .Z(n8364) );
  NBUFFX2 U8202 ( .INP(n8492), .Z(n8363) );
  NBUFFX2 U8203 ( .INP(n8492), .Z(n8362) );
  NBUFFX2 U8204 ( .INP(n8492), .Z(n8361) );
  NBUFFX2 U8205 ( .INP(n8493), .Z(n8360) );
  NBUFFX2 U8206 ( .INP(n8494), .Z(n8355) );
  NBUFFX2 U8207 ( .INP(n8499), .Z(n8342) );
  NBUFFX2 U8208 ( .INP(n8494), .Z(n8356) );
  NBUFFX2 U8209 ( .INP(n8495), .Z(n8352) );
  NBUFFX2 U8210 ( .INP(n8495), .Z(n8354) );
  NBUFFX2 U8211 ( .INP(n8495), .Z(n8353) );
  NBUFFX2 U8212 ( .INP(n8498), .Z(n8344) );
  NBUFFX2 U8213 ( .INP(n8496), .Z(n8349) );
  NBUFFX2 U8214 ( .INP(n8496), .Z(n8351) );
  NBUFFX2 U8215 ( .INP(n8496), .Z(n8350) );
  NBUFFX2 U8216 ( .INP(n8498), .Z(n8345) );
  NBUFFX2 U8217 ( .INP(n8498), .Z(n8343) );
  NBUFFX2 U8218 ( .INP(n8497), .Z(n8346) );
  NBUFFX2 U8219 ( .INP(n8497), .Z(n8348) );
  NBUFFX2 U8220 ( .INP(n8497), .Z(n8347) );
  NBUFFX2 U8221 ( .INP(n8501), .Z(n8335) );
  NBUFFX2 U8222 ( .INP(n8501), .Z(n8334) );
  NBUFFX2 U8223 ( .INP(n8460), .Z(n8457) );
  NBUFFX2 U8224 ( .INP(n8502), .Z(n8333) );
  NBUFFX2 U8225 ( .INP(n8460), .Z(n8458) );
  NBUFFX2 U8226 ( .INP(n8461), .Z(n8456) );
  NBUFFX2 U8227 ( .INP(n8461), .Z(n8455) );
  NBUFFX2 U8228 ( .INP(n8494), .Z(n8357) );
  NBUFFX2 U8229 ( .INP(n8499), .Z(n8340) );
  NBUFFX2 U8230 ( .INP(n8500), .Z(n8339) );
  NBUFFX2 U8231 ( .INP(n8500), .Z(n8338) );
  NBUFFX2 U8232 ( .INP(n8500), .Z(n8337) );
  NBUFFX2 U8233 ( .INP(n8501), .Z(n8336) );
  NBUFFX2 U8234 ( .INP(n8502), .Z(n8332) );
  NBUFFX2 U8235 ( .INP(n8502), .Z(n8331) );
  NBUFFX2 U8236 ( .INP(n8273), .Z(n8272) );
  NBUFFX2 U8237 ( .INP(n8460), .Z(n8459) );
  NBUFFX2 U8238 ( .INP(n8512), .Z(n8462) );
  NBUFFX2 U8239 ( .INP(n8325), .Z(n8275) );
  NBUFFX2 U8240 ( .INP(n8512), .Z(n8463) );
  NBUFFX2 U8241 ( .INP(n8325), .Z(n8276) );
  NBUFFX2 U8242 ( .INP(n8512), .Z(n8460) );
  NBUFFX2 U8243 ( .INP(n8325), .Z(n8273) );
  NBUFFX2 U8244 ( .INP(n8512), .Z(n8461) );
  NBUFFX2 U8245 ( .INP(n8325), .Z(n8274) );
  NBUFFX2 U8246 ( .INP(n8511), .Z(n8465) );
  NBUFFX2 U8247 ( .INP(n8324), .Z(n8278) );
  NBUFFX2 U8248 ( .INP(n8511), .Z(n8464) );
  NBUFFX2 U8249 ( .INP(n8324), .Z(n8277) );
  NBUFFX2 U8250 ( .INP(n8511), .Z(n8466) );
  NBUFFX2 U8251 ( .INP(n8324), .Z(n8279) );
  NBUFFX2 U8252 ( .INP(n8511), .Z(n8467) );
  NBUFFX2 U8253 ( .INP(n8324), .Z(n8280) );
  NBUFFX2 U8254 ( .INP(n8511), .Z(n8468) );
  NBUFFX2 U8255 ( .INP(n8324), .Z(n8281) );
  NBUFFX2 U8256 ( .INP(n8510), .Z(n8469) );
  NBUFFX2 U8257 ( .INP(n8323), .Z(n8282) );
  NBUFFX2 U8258 ( .INP(n8510), .Z(n8470) );
  NBUFFX2 U8259 ( .INP(n8323), .Z(n8283) );
  NBUFFX2 U8260 ( .INP(n8510), .Z(n8471) );
  NBUFFX2 U8261 ( .INP(n8323), .Z(n8284) );
  NBUFFX2 U8262 ( .INP(n8510), .Z(n8472) );
  NBUFFX2 U8263 ( .INP(n8323), .Z(n8285) );
  NBUFFX2 U8264 ( .INP(n8510), .Z(n8473) );
  NBUFFX2 U8265 ( .INP(n8323), .Z(n8286) );
  NBUFFX2 U8266 ( .INP(n8509), .Z(n8474) );
  NBUFFX2 U8267 ( .INP(n8322), .Z(n8287) );
  NBUFFX2 U8268 ( .INP(n8509), .Z(n8475) );
  NBUFFX2 U8269 ( .INP(n8322), .Z(n8288) );
  NBUFFX2 U8270 ( .INP(n8509), .Z(n8476) );
  NBUFFX2 U8271 ( .INP(n8322), .Z(n8289) );
  NBUFFX2 U8272 ( .INP(n8509), .Z(n8477) );
  NBUFFX2 U8273 ( .INP(n8322), .Z(n8290) );
  NBUFFX2 U8274 ( .INP(n8509), .Z(n8478) );
  NBUFFX2 U8275 ( .INP(n8322), .Z(n8291) );
  NBUFFX2 U8276 ( .INP(n8508), .Z(n8479) );
  NBUFFX2 U8277 ( .INP(n8321), .Z(n8292) );
  NBUFFX2 U8278 ( .INP(n8508), .Z(n8480) );
  NBUFFX2 U8279 ( .INP(n8321), .Z(n8293) );
  NBUFFX2 U8280 ( .INP(n8508), .Z(n8481) );
  NBUFFX2 U8281 ( .INP(n8321), .Z(n8294) );
  NBUFFX2 U8282 ( .INP(n8508), .Z(n8482) );
  NBUFFX2 U8283 ( .INP(n8321), .Z(n8295) );
  NBUFFX2 U8284 ( .INP(n8507), .Z(n8484) );
  NBUFFX2 U8285 ( .INP(n8320), .Z(n8297) );
  NBUFFX2 U8286 ( .INP(n8508), .Z(n8483) );
  NBUFFX2 U8287 ( .INP(n8321), .Z(n8296) );
  NBUFFX2 U8288 ( .INP(n8507), .Z(n8485) );
  NBUFFX2 U8289 ( .INP(n8320), .Z(n8298) );
  NBUFFX2 U8290 ( .INP(n8507), .Z(n8486) );
  NBUFFX2 U8291 ( .INP(n8320), .Z(n8299) );
  NBUFFX2 U8292 ( .INP(n8507), .Z(n8487) );
  NBUFFX2 U8293 ( .INP(n8320), .Z(n8300) );
  NBUFFX2 U8294 ( .INP(n8506), .Z(n8490) );
  NBUFFX2 U8295 ( .INP(n8319), .Z(n8303) );
  NBUFFX2 U8296 ( .INP(n8507), .Z(n8488) );
  NBUFFX2 U8297 ( .INP(n8320), .Z(n8301) );
  NBUFFX2 U8298 ( .INP(n8506), .Z(n8489) );
  NBUFFX2 U8299 ( .INP(n8319), .Z(n8302) );
  NBUFFX2 U8300 ( .INP(n8506), .Z(n8491) );
  NBUFFX2 U8301 ( .INP(n8319), .Z(n8304) );
  NBUFFX2 U8302 ( .INP(n8506), .Z(n8492) );
  NBUFFX2 U8303 ( .INP(n8319), .Z(n8305) );
  NBUFFX2 U8304 ( .INP(n8506), .Z(n8493) );
  NBUFFX2 U8305 ( .INP(n8319), .Z(n8306) );
  NBUFFX2 U8306 ( .INP(n8505), .Z(n8495) );
  NBUFFX2 U8307 ( .INP(n8318), .Z(n8308) );
  NBUFFX2 U8308 ( .INP(n8505), .Z(n8496) );
  NBUFFX2 U8309 ( .INP(n8318), .Z(n8309) );
  NBUFFX2 U8310 ( .INP(n8505), .Z(n8498) );
  NBUFFX2 U8311 ( .INP(n8318), .Z(n8311) );
  NBUFFX2 U8312 ( .INP(n8505), .Z(n8497) );
  NBUFFX2 U8313 ( .INP(n8318), .Z(n8310) );
  NBUFFX2 U8314 ( .INP(n8505), .Z(n8494) );
  NBUFFX2 U8315 ( .INP(n8318), .Z(n8307) );
  NBUFFX2 U8316 ( .INP(n8504), .Z(n8499) );
  NBUFFX2 U8317 ( .INP(n8317), .Z(n8312) );
  NBUFFX2 U8318 ( .INP(n8504), .Z(n8500) );
  NBUFFX2 U8319 ( .INP(n8317), .Z(n8313) );
  NBUFFX2 U8320 ( .INP(n8504), .Z(n8501) );
  NBUFFX2 U8321 ( .INP(n8317), .Z(n8314) );
  NBUFFX2 U8322 ( .INP(n8504), .Z(n8502) );
  NBUFFX2 U8323 ( .INP(n8317), .Z(n8315) );
  NBUFFX2 U8324 ( .INP(n8504), .Z(n8503) );
  NBUFFX2 U8325 ( .INP(n8317), .Z(n8316) );
  NBUFFX2 U8326 ( .INP(n8328), .Z(n8317) );
  NBUFFX2 U8327 ( .INP(n8328), .Z(n8318) );
  NBUFFX2 U8328 ( .INP(n8328), .Z(n8319) );
  NBUFFX2 U8329 ( .INP(n8327), .Z(n8320) );
  NBUFFX2 U8330 ( .INP(n8327), .Z(n8321) );
  NBUFFX2 U8331 ( .INP(n8327), .Z(n8322) );
  NBUFFX2 U8332 ( .INP(n8326), .Z(n8323) );
  NBUFFX2 U8333 ( .INP(n8326), .Z(n8324) );
  NBUFFX2 U8334 ( .INP(n8326), .Z(n8325) );
  NBUFFX2 U8335 ( .INP(test_se), .Z(n8326) );
  NBUFFX2 U8336 ( .INP(test_se), .Z(n8327) );
  NBUFFX2 U8337 ( .INP(test_se), .Z(n8328) );
  NBUFFX2 U8338 ( .INP(n8515), .Z(n8504) );
  NBUFFX2 U8339 ( .INP(n8515), .Z(n8505) );
  NBUFFX2 U8340 ( .INP(n8515), .Z(n8506) );
  NBUFFX2 U8341 ( .INP(n8514), .Z(n8507) );
  NBUFFX2 U8342 ( .INP(n8514), .Z(n8508) );
  NBUFFX2 U8343 ( .INP(n8514), .Z(n8509) );
  NBUFFX2 U8344 ( .INP(n8513), .Z(n8510) );
  NBUFFX2 U8345 ( .INP(n8513), .Z(n8511) );
  NBUFFX2 U8346 ( .INP(n8513), .Z(n8512) );
  NBUFFX2 U8347 ( .INP(CK), .Z(n8513) );
  NBUFFX2 U8348 ( .INP(CK), .Z(n8514) );
  NBUFFX2 U8349 ( .INP(CK), .Z(n8515) );
  INVX0 U8350 ( .INP(n8516), .ZN(n971) );
  INVX0 U8351 ( .INP(n8517), .ZN(n913) );
  NAND3X0 U8352 ( .IN1(n8518), .IN2(n8519), .IN3(n8520), .QN(n8517) );
  NAND2X0 U8353 ( .IN1(n8521), .IN2(n4411), .QN(n8518) );
  NAND2X0 U8354 ( .IN1(g1346), .IN2(n8522), .QN(n8521) );
  NOR3X0 U8355 ( .IN1(n8523), .IN2(n8524), .IN3(n8525), .QN(n912) );
  NOR2X0 U8356 ( .IN1(n8526), .IN2(g1319), .QN(n8523) );
  NOR2X0 U8357 ( .IN1(n4402), .IN2(n8527), .QN(n8526) );
  NOR2X0 U8358 ( .IN1(n8524), .IN2(n8528), .QN(n883) );
  INVX0 U8359 ( .INP(n8529), .ZN(n8528) );
  NAND2X0 U8360 ( .IN1(n8530), .IN2(n7976), .QN(n8529) );
  INVX0 U8361 ( .INP(n8531), .ZN(n837) );
  NOR2X0 U8362 ( .IN1(n8532), .IN2(n8533), .QN(n8531) );
  NOR2X0 U8363 ( .IN1(g1236), .IN2(n7992), .QN(n8533) );
  INVX0 U8364 ( .INP(n8534), .ZN(n833) );
  INVX0 U8365 ( .INP(n8535), .ZN(n819) );
  INVX0 U8366 ( .INP(n8536), .ZN(n672) );
  INVX0 U8367 ( .INP(n8537), .ZN(n616) );
  NAND3X0 U8368 ( .IN1(n8538), .IN2(n8539), .IN3(n8540), .QN(n8537) );
  NAND2X0 U8369 ( .IN1(n8541), .IN2(n4413), .QN(n8538) );
  NAND2X0 U8370 ( .IN1(g660), .IN2(n8542), .QN(n8541) );
  INVX0 U8371 ( .INP(n8543), .ZN(n615) );
  NAND3X0 U8372 ( .IN1(n8544), .IN2(n8539), .IN3(n8545), .QN(n8543) );
  NAND2X0 U8373 ( .IN1(n8546), .IN2(n4478), .QN(n8544) );
  NAND2X0 U8374 ( .IN1(g640), .IN2(n8547), .QN(n8546) );
  NOR2X0 U8375 ( .IN1(n8548), .IN2(n8549), .QN(n586) );
  INVX0 U8376 ( .INP(n8550), .ZN(n8549) );
  NAND2X0 U8377 ( .IN1(n8551), .IN2(n7977), .QN(n8550) );
  INVX0 U8378 ( .INP(n8552), .ZN(n539) );
  NOR2X0 U8379 ( .IN1(n8553), .IN2(n8554), .QN(n8552) );
  NOR2X0 U8380 ( .IN1(g550), .IN2(n7993), .QN(n8554) );
  INVX0 U8381 ( .INP(n8555), .ZN(n534) );
  INVX0 U8382 ( .INP(n8556), .ZN(n533) );
  INVX0 U8383 ( .INP(n8557), .ZN(n532) );
  INVX0 U8384 ( .INP(n8558), .ZN(n518) );
  INVX0 U8385 ( .INP(n8559), .ZN(n494) );
  INVX0 U8386 ( .INP(n8560), .ZN(n472) );
  XNOR2X1 U8387 ( .IN1(n8033), .IN2(n8561), .Q(n4281) );
  XOR2X1 U8388 ( .IN1(n8562), .IN2(n8035), .Q(n4280) );
  NAND2X0 U8389 ( .IN1(g2879), .IN2(n8563), .QN(n4279) );
  NAND2X0 U8390 ( .IN1(DFF_18_n1), .IN2(g8021), .QN(n8563) );
  NOR2X0 U8391 ( .IN1(n8564), .IN2(n8565), .QN(n4278) );
  NOR2X0 U8392 ( .IN1(n8566), .IN2(n8567), .QN(n8565) );
  INVX0 U8393 ( .INP(n8568), .ZN(n8567) );
  NOR4X0 U8394 ( .IN1(n8569), .IN2(n8570), .IN3(n8571), .IN4(n8572), .QN(n8564) );
  NAND3X0 U8395 ( .IN1(n8573), .IN2(n8574), .IN3(n8575), .QN(n8572) );
  XOR2X1 U8396 ( .IN1(n7176), .IN2(n8576), .Q(n8575) );
  XOR2X1 U8397 ( .IN1(n8093), .IN2(n8577), .Q(n8574) );
  XOR2X1 U8398 ( .IN1(n8070), .IN2(n8578), .Q(n8573) );
  NAND3X0 U8399 ( .IN1(n8579), .IN2(n8580), .IN3(n8581), .QN(n8571) );
  XOR2X1 U8400 ( .IN1(n7711), .IN2(n8582), .Q(n8581) );
  XOR2X1 U8401 ( .IN1(g88), .IN2(n8583), .Q(n8580) );
  XOR2X1 U8402 ( .IN1(n7337), .IN2(n8584), .Q(n8579) );
  NAND3X0 U8403 ( .IN1(n8585), .IN2(n8586), .IN3(n8587), .QN(n8570) );
  XOR2X1 U8404 ( .IN1(n7712), .IN2(n8588), .Q(n8587) );
  XOR2X1 U8405 ( .IN1(n7713), .IN2(n8589), .Q(n8586) );
  XOR2X1 U8406 ( .IN1(n7714), .IN2(n8590), .Q(n8585) );
  NAND3X0 U8407 ( .IN1(n8591), .IN2(n8592), .IN3(n8593), .QN(n8569) );
  XOR2X1 U8408 ( .IN1(test_so15), .IN2(n8594), .Q(n8593) );
  NOR2X0 U8409 ( .IN1(n8595), .IN2(n8596), .QN(n4277) );
  NOR2X0 U8410 ( .IN1(n8597), .IN2(n8598), .QN(n8596) );
  NOR4X0 U8411 ( .IN1(n8599), .IN2(n8600), .IN3(n8601), .IN4(n8602), .QN(n8595) );
  NAND3X0 U8412 ( .IN1(n8603), .IN2(n8604), .IN3(n8605), .QN(n8602) );
  XOR2X1 U8413 ( .IN1(n8606), .IN2(n7709), .Q(n8605) );
  XOR2X1 U8414 ( .IN1(n8607), .IN2(n7336), .Q(n8604) );
  XOR2X1 U8415 ( .IN1(n8608), .IN2(n7175), .Q(n8603) );
  NAND3X0 U8416 ( .IN1(n8609), .IN2(n8610), .IN3(n8611), .QN(n8601) );
  XOR2X1 U8417 ( .IN1(n8612), .IN2(n8092), .Q(n8611) );
  XOR2X1 U8418 ( .IN1(n8613), .IN2(n7708), .Q(n8610) );
  XOR2X1 U8419 ( .IN1(n8614), .IN2(n7707), .Q(n8609) );
  NAND3X0 U8420 ( .IN1(n8615), .IN2(n8616), .IN3(n8617), .QN(n8600) );
  XOR2X1 U8421 ( .IN1(n8618), .IN2(n7710), .Q(n8617) );
  XOR2X1 U8422 ( .IN1(n8619), .IN2(n8085), .Q(n8616) );
  XOR2X1 U8423 ( .IN1(n8620), .IN2(n8091), .Q(n8615) );
  NAND3X0 U8424 ( .IN1(n8621), .IN2(n8591), .IN3(n8622), .QN(n8599) );
  XNOR2X1 U8425 ( .IN1(test_so36), .IN2(n8623), .Q(n8622) );
  NOR2X0 U8426 ( .IN1(n8624), .IN2(n8625), .QN(n4276) );
  NOR2X0 U8427 ( .IN1(n8626), .IN2(n8627), .QN(n8625) );
  INVX0 U8428 ( .INP(n8628), .ZN(n8627) );
  NOR2X0 U8429 ( .IN1(n8629), .IN2(n8630), .QN(n8624) );
  NAND4X0 U8430 ( .IN1(n8631), .IN2(n8632), .IN3(n8633), .IN4(n8634), .QN(
        n8630) );
  NOR3X0 U8431 ( .IN1(n8635), .IN2(n8636), .IN3(n8637), .QN(n8634) );
  XOR2X1 U8432 ( .IN1(n7703), .IN2(n8638), .Q(n8637) );
  XOR2X1 U8433 ( .IN1(n8071), .IN2(n8639), .Q(n8636) );
  XOR2X1 U8434 ( .IN1(n8069), .IN2(n8640), .Q(n8635) );
  XOR2X1 U8435 ( .IN1(g1453), .IN2(n8641), .Q(n8633) );
  XOR2X1 U8436 ( .IN1(n8094), .IN2(n8642), .Q(n8632) );
  XOR2X1 U8437 ( .IN1(n7174), .IN2(n8643), .Q(n8631) );
  NAND4X0 U8438 ( .IN1(n8644), .IN2(n8591), .IN3(n8645), .IN4(n8646), .QN(
        n8629) );
  NOR3X0 U8439 ( .IN1(n8647), .IN2(n8648), .IN3(n8649), .QN(n8646) );
  XNOR2X1 U8440 ( .IN1(n7705), .IN2(n8650), .Q(n8649) );
  XNOR2X1 U8441 ( .IN1(n7706), .IN2(n8651), .Q(n8648) );
  XOR2X1 U8442 ( .IN1(n7335), .IN2(n8652), .Q(n8647) );
  XOR2X1 U8443 ( .IN1(n7704), .IN2(n8653), .Q(n8645) );
  NOR2X0 U8444 ( .IN1(n8654), .IN2(n8655), .QN(n4275) );
  NOR2X0 U8445 ( .IN1(n8656), .IN2(n8657), .QN(n8655) );
  NOR4X0 U8446 ( .IN1(n8658), .IN2(n8659), .IN3(n8660), .IN4(n8661), .QN(n8654) );
  NAND3X0 U8447 ( .IN1(n8662), .IN2(n8663), .IN3(n8664), .QN(n8661) );
  XOR2X1 U8448 ( .IN1(n8665), .IN2(n8075), .Q(n8664) );
  XOR2X1 U8449 ( .IN1(n8666), .IN2(n8095), .Q(n8663) );
  XOR2X1 U8450 ( .IN1(n8667), .IN2(n7173), .Q(n8662) );
  NAND3X0 U8451 ( .IN1(n8668), .IN2(n8669), .IN3(n8670), .QN(n8660) );
  XOR2X1 U8452 ( .IN1(n8671), .IN2(n7699), .Q(n8670) );
  XOR2X1 U8453 ( .IN1(n8672), .IN2(n8072), .Q(n8669) );
  XOR2X1 U8454 ( .IN1(n8673), .IN2(n7702), .Q(n8668) );
  NAND3X0 U8455 ( .IN1(n8674), .IN2(n8675), .IN3(n8676), .QN(n8659) );
  XOR2X1 U8456 ( .IN1(n8677), .IN2(n7701), .Q(n8676) );
  XOR2X1 U8457 ( .IN1(n8678), .IN2(n7334), .Q(n8675) );
  XOR2X1 U8458 ( .IN1(n8679), .IN2(n7700), .Q(n8674) );
  NAND3X0 U8459 ( .IN1(n8680), .IN2(n8591), .IN3(n8681), .QN(n8658) );
  XOR2X1 U8460 ( .IN1(test_so78), .IN2(n8682), .Q(n8681) );
  NAND2X0 U8461 ( .IN1(n8683), .IN2(n8684), .QN(n4274) );
  INVX0 U8462 ( .INP(n8685), .ZN(n8684) );
  XNOR2X1 U8463 ( .IN1(n4330), .IN2(n4423), .Q(n8683) );
  NAND2X0 U8464 ( .IN1(n8686), .IN2(n8687), .QN(n4273) );
  NAND2X0 U8465 ( .IN1(n8688), .IN2(n8689), .QN(n8687) );
  NAND2X0 U8466 ( .IN1(n4482), .IN2(n8690), .QN(n8688) );
  NAND2X0 U8467 ( .IN1(n2426), .IN2(n8691), .QN(n4272) );
  NAND3X0 U8468 ( .IN1(n8692), .IN2(n8693), .IN3(n8694), .QN(n8691) );
  NAND2X0 U8469 ( .IN1(n8695), .IN2(n8696), .QN(n8693) );
  INVX0 U8470 ( .INP(n8697), .ZN(n8695) );
  NAND2X0 U8471 ( .IN1(n8698), .IN2(DFF_449_n1), .QN(n8692) );
  NAND2X0 U8472 ( .IN1(n8699), .IN2(n8700), .QN(n4271) );
  NAND2X0 U8473 ( .IN1(n2446), .IN2(n8701), .QN(n8700) );
  NAND3X0 U8474 ( .IN1(n8702), .IN2(n8703), .IN3(n8694), .QN(n8699) );
  NAND2X0 U8475 ( .IN1(n8704), .IN2(n8696), .QN(n8703) );
  INVX0 U8476 ( .INP(n8705), .ZN(n8704) );
  NAND2X0 U8477 ( .IN1(n7155), .IN2(n8698), .QN(n8702) );
  NAND2X0 U8478 ( .IN1(n8706), .IN2(n8707), .QN(n4270) );
  NAND2X0 U8479 ( .IN1(n2446), .IN2(n8708), .QN(n8707) );
  NAND3X0 U8480 ( .IN1(n8709), .IN2(n8710), .IN3(n8694), .QN(n8706) );
  NAND2X0 U8481 ( .IN1(n8711), .IN2(n8696), .QN(n8710) );
  NAND2X0 U8482 ( .IN1(n7154), .IN2(n8698), .QN(n8709) );
  NAND2X0 U8483 ( .IN1(n8712), .IN2(n8713), .QN(n4269) );
  NAND3X0 U8484 ( .IN1(n8714), .IN2(n8715), .IN3(n8694), .QN(n8713) );
  NAND2X0 U8485 ( .IN1(n8716), .IN2(n8696), .QN(n8715) );
  INVX0 U8486 ( .INP(n8717), .ZN(n8716) );
  NAND2X0 U8487 ( .IN1(n8698), .IN2(DFF_444_n1), .QN(n8714) );
  NAND3X0 U8488 ( .IN1(n2426), .IN2(n8718), .IN3(n2440), .QN(n4268) );
  NAND3X0 U8489 ( .IN1(n8719), .IN2(n8720), .IN3(n8694), .QN(n8718) );
  NAND2X0 U8490 ( .IN1(n8721), .IN2(n8696), .QN(n8720) );
  INVX0 U8491 ( .INP(n8722), .ZN(n8721) );
  NAND2X0 U8492 ( .IN1(n8698), .IN2(DFF_445_n1), .QN(n8719) );
  NAND3X0 U8493 ( .IN1(n2426), .IN2(n8723), .IN3(n2440), .QN(n4267) );
  NAND3X0 U8494 ( .IN1(n8724), .IN2(n8725), .IN3(n8694), .QN(n8723) );
  NAND2X0 U8495 ( .IN1(n8726), .IN2(n8696), .QN(n8725) );
  INVX0 U8496 ( .INP(n8727), .ZN(n8726) );
  NAND2X0 U8497 ( .IN1(n8698), .IN2(DFF_446_n1), .QN(n8724) );
  NAND2X0 U8498 ( .IN1(n8712), .IN2(n8728), .QN(n4266) );
  NAND3X0 U8499 ( .IN1(n8729), .IN2(n8730), .IN3(n8694), .QN(n8728) );
  NAND2X0 U8500 ( .IN1(n8731), .IN2(n8696), .QN(n8730) );
  NAND2X0 U8501 ( .IN1(n8698), .IN2(DFF_447_n1), .QN(n8729) );
  INVX0 U8502 ( .INP(n8732), .ZN(n8712) );
  NAND2X0 U8503 ( .IN1(n2426), .IN2(n8733), .QN(n8732) );
  NAND2X0 U8504 ( .IN1(n2446), .IN2(n2445), .QN(n8733) );
  NAND2X0 U8505 ( .IN1(n2426), .IN2(n8734), .QN(n4265) );
  NAND3X0 U8506 ( .IN1(n8735), .IN2(n8736), .IN3(n8694), .QN(n8734) );
  NAND2X0 U8507 ( .IN1(n8737), .IN2(n8696), .QN(n8736) );
  INVX0 U8508 ( .INP(n8738), .ZN(n8737) );
  NAND2X0 U8509 ( .IN1(n8698), .IN2(DFF_448_n1), .QN(n8735) );
  NAND2X0 U8510 ( .IN1(DFF_1562_n1), .IN2(n8739), .QN(n4263) );
  NAND2X0 U8511 ( .IN1(n8740), .IN2(n8741), .QN(n4262) );
  XOR2X1 U8512 ( .IN1(n4481), .IN2(n8742), .Q(n8740) );
  XNOR2X1 U8513 ( .IN1(n8743), .IN2(n8744), .Q(n4261) );
  XOR2X1 U8514 ( .IN1(n8744), .IN2(n8745), .Q(n4260) );
  INVX0 U8515 ( .INP(n8746), .ZN(n8745) );
  NOR2X0 U8516 ( .IN1(g3231), .IN2(n14386), .QN(n8744) );
  NAND3X0 U8517 ( .IN1(n8747), .IN2(n8748), .IN3(n8749), .QN(n4259) );
  NAND2X0 U8518 ( .IN1(test_so22), .IN2(n8750), .QN(n8749) );
  XOR2X1 U8519 ( .IN1(n8751), .IN2(n8752), .Q(n8750) );
  XNOR3X1 U8520 ( .IN1(n8738), .IN2(n8731), .IN3(n8753), .Q(n8752) );
  XNOR2X1 U8521 ( .IN1(n8722), .IN2(n8727), .Q(n8753) );
  NAND3X0 U8522 ( .IN1(n8754), .IN2(n8755), .IN3(n8756), .QN(n8727) );
  NAND2X0 U8523 ( .IN1(n8757), .IN2(n8758), .QN(n8755) );
  NAND2X0 U8524 ( .IN1(n8759), .IN2(n8760), .QN(n8754) );
  NAND3X0 U8525 ( .IN1(n8761), .IN2(n8762), .IN3(n8756), .QN(n8722) );
  NAND2X0 U8526 ( .IN1(n8763), .IN2(n8764), .QN(n8762) );
  NAND2X0 U8527 ( .IN1(n8765), .IN2(n8766), .QN(n8761) );
  INVX0 U8528 ( .INP(n8767), .ZN(n8731) );
  NAND3X0 U8529 ( .IN1(n8768), .IN2(n8769), .IN3(n8756), .QN(n8767) );
  NAND2X0 U8530 ( .IN1(n8770), .IN2(n8764), .QN(n8769) );
  NAND2X0 U8531 ( .IN1(n8765), .IN2(n8771), .QN(n8768) );
  NAND3X0 U8532 ( .IN1(n8772), .IN2(n8773), .IN3(n8774), .QN(n8738) );
  NAND2X0 U8533 ( .IN1(n8775), .IN2(n8758), .QN(n8773) );
  NAND2X0 U8534 ( .IN1(n8759), .IN2(n8776), .QN(n8772) );
  XNOR3X1 U8535 ( .IN1(n8717), .IN2(n8711), .IN3(n8777), .Q(n8751) );
  XNOR2X1 U8536 ( .IN1(n8697), .IN2(n8705), .Q(n8777) );
  NAND3X0 U8537 ( .IN1(n8778), .IN2(n8779), .IN3(n8774), .QN(n8705) );
  NAND2X0 U8538 ( .IN1(n8780), .IN2(n8758), .QN(n8779) );
  NAND2X0 U8539 ( .IN1(n8759), .IN2(n8781), .QN(n8778) );
  NAND3X0 U8540 ( .IN1(n8782), .IN2(n8783), .IN3(n8784), .QN(n8697) );
  NAND2X0 U8541 ( .IN1(n8785), .IN2(n8764), .QN(n8783) );
  NAND2X0 U8542 ( .IN1(n8765), .IN2(n8786), .QN(n8782) );
  INVX0 U8543 ( .INP(n8787), .ZN(n8711) );
  NAND3X0 U8544 ( .IN1(n8788), .IN2(n8789), .IN3(n8756), .QN(n8787) );
  NAND2X0 U8545 ( .IN1(n8790), .IN2(n8764), .QN(n8789) );
  NAND2X0 U8546 ( .IN1(n8765), .IN2(n8791), .QN(n8788) );
  NAND3X0 U8547 ( .IN1(n8792), .IN2(n8793), .IN3(n8756), .QN(n8717) );
  NAND2X0 U8548 ( .IN1(n8794), .IN2(n8758), .QN(n8793) );
  NAND2X0 U8549 ( .IN1(n8759), .IN2(n8795), .QN(n8792) );
  NAND4X0 U8550 ( .IN1(n8694), .IN2(n8698), .IN3(n8796), .IN4(n8797), .QN(
        n8748) );
  NAND2X0 U8551 ( .IN1(n14378), .IN2(n8798), .QN(n8797) );
  NAND2X0 U8552 ( .IN1(n4492), .IN2(g3229), .QN(n8796) );
  NOR2X0 U8553 ( .IN1(n8696), .IN2(n8560), .QN(n8698) );
  NAND2X0 U8554 ( .IN1(n8799), .IN2(g557), .QN(n8747) );
  XOR2X1 U8555 ( .IN1(n8701), .IN2(n8708), .Q(n8799) );
  NAND3X0 U8556 ( .IN1(n8800), .IN2(n8801), .IN3(n8784), .QN(n8708) );
  INVX0 U8557 ( .INP(n8802), .ZN(n8784) );
  NAND2X0 U8558 ( .IN1(n8756), .IN2(n8803), .QN(n8802) );
  NAND2X0 U8559 ( .IN1(n8804), .IN2(n8764), .QN(n8803) );
  NAND2X0 U8560 ( .IN1(n8805), .IN2(n8764), .QN(n8801) );
  NAND2X0 U8561 ( .IN1(n8765), .IN2(n8806), .QN(n8800) );
  NOR2X0 U8562 ( .IN1(n8764), .IN2(n8804), .QN(n8765) );
  NAND3X0 U8563 ( .IN1(n8807), .IN2(n8808), .IN3(n8774), .QN(n8701) );
  INVX0 U8564 ( .INP(n8809), .ZN(n8774) );
  NAND2X0 U8565 ( .IN1(n8756), .IN2(n2430), .QN(n8809) );
  NOR2X0 U8566 ( .IN1(n8560), .IN2(n4541), .QN(n8756) );
  NAND3X0 U8567 ( .IN1(n8810), .IN2(n7756), .IN3(n8811), .QN(n8560) );
  NOR2X0 U8568 ( .IN1(g563), .IN2(n8812), .QN(n8811) );
  NOR2X0 U8569 ( .IN1(n4298), .IN2(g499), .QN(n8812) );
  INVX0 U8570 ( .INP(g21851), .ZN(n8810) );
  NAND2X0 U8571 ( .IN1(n8813), .IN2(n8758), .QN(n8808) );
  NAND2X0 U8572 ( .IN1(n8759), .IN2(n8814), .QN(n8807) );
  NOR2X0 U8573 ( .IN1(n8758), .IN2(n8804), .QN(n8759) );
  NAND2X0 U8574 ( .IN1(n8815), .IN2(n8816), .QN(n4258) );
  NAND2X0 U8575 ( .IN1(n2361), .IN2(n8817), .QN(n8816) );
  NAND3X0 U8576 ( .IN1(n8818), .IN2(n8819), .IN3(n8820), .QN(n8815) );
  NAND2X0 U8577 ( .IN1(n8821), .IN2(n8822), .QN(n8819) );
  NAND2X0 U8578 ( .IN1(n7156), .IN2(n8823), .QN(n8818) );
  NAND3X0 U8579 ( .IN1(n8824), .IN2(n8825), .IN3(n2375), .QN(n4257) );
  NAND3X0 U8580 ( .IN1(n8826), .IN2(n8827), .IN3(n8820), .QN(n8824) );
  NAND2X0 U8581 ( .IN1(n8828), .IN2(n8822), .QN(n8827) );
  INVX0 U8582 ( .INP(n8829), .ZN(n8828) );
  NAND2X0 U8583 ( .IN1(n8823), .IN2(DFF_1495_n1), .QN(n8826) );
  NAND2X0 U8584 ( .IN1(n8825), .IN2(n8830), .QN(n4256) );
  NAND3X0 U8585 ( .IN1(n8831), .IN2(n8832), .IN3(n8820), .QN(n8830) );
  NAND2X0 U8586 ( .IN1(n8833), .IN2(n8822), .QN(n8832) );
  NAND2X0 U8587 ( .IN1(n8823), .IN2(DFF_1499_n1), .QN(n8831) );
  NAND3X0 U8588 ( .IN1(n8834), .IN2(n8825), .IN3(n2375), .QN(n4255) );
  NAND3X0 U8589 ( .IN1(n8835), .IN2(n8836), .IN3(n8820), .QN(n8834) );
  NAND2X0 U8590 ( .IN1(n8837), .IN2(n8822), .QN(n8836) );
  NAND2X0 U8591 ( .IN1(n8823), .IN2(DFF_1496_n1), .QN(n8835) );
  NAND2X0 U8592 ( .IN1(n8838), .IN2(n8839), .QN(n4254) );
  NAND3X0 U8593 ( .IN1(n8840), .IN2(n8841), .IN3(n8820), .QN(n8839) );
  NAND2X0 U8594 ( .IN1(n8842), .IN2(n8822), .QN(n8841) );
  NAND2X0 U8595 ( .IN1(n8823), .IN2(DFF_1494_n1), .QN(n8840) );
  NAND2X0 U8596 ( .IN1(n8843), .IN2(n8844), .QN(n4253) );
  NAND2X0 U8597 ( .IN1(n2361), .IN2(n8845), .QN(n8844) );
  NAND3X0 U8598 ( .IN1(n8846), .IN2(n8847), .IN3(n8820), .QN(n8843) );
  NAND2X0 U8599 ( .IN1(n8848), .IN2(n8822), .QN(n8847) );
  INVX0 U8600 ( .INP(n8849), .ZN(n8848) );
  NAND2X0 U8601 ( .IN1(n8823), .IN2(n7157), .QN(n8846) );
  NAND2X0 U8602 ( .IN1(n8838), .IN2(n8850), .QN(n4252) );
  NAND3X0 U8603 ( .IN1(n8851), .IN2(n8852), .IN3(n8820), .QN(n8850) );
  NAND2X0 U8604 ( .IN1(n8853), .IN2(n8822), .QN(n8852) );
  INVX0 U8605 ( .INP(n8854), .ZN(n8853) );
  NAND2X0 U8606 ( .IN1(n8823), .IN2(DFF_1497_n1), .QN(n8851) );
  INVX0 U8607 ( .INP(n8855), .ZN(n8838) );
  NAND2X0 U8608 ( .IN1(n8825), .IN2(n8856), .QN(n8855) );
  NAND2X0 U8609 ( .IN1(n2361), .IN2(n2374), .QN(n8856) );
  NAND2X0 U8610 ( .IN1(n8825), .IN2(n8857), .QN(n4251) );
  NAND3X0 U8611 ( .IN1(n8858), .IN2(n8859), .IN3(n8820), .QN(n8857) );
  NAND2X0 U8612 ( .IN1(n8860), .IN2(n8822), .QN(n8859) );
  INVX0 U8613 ( .INP(n8861), .ZN(n8860) );
  NAND2X0 U8614 ( .IN1(n8823), .IN2(DFF_1498_n1), .QN(n8858) );
  NAND2X0 U8615 ( .IN1(n2361), .IN2(n8862), .QN(n8825) );
  NAND3X0 U8616 ( .IN1(n8863), .IN2(n8864), .IN3(n8865), .QN(n4250) );
  NAND2X0 U8617 ( .IN1(n8866), .IN2(g2584), .QN(n8865) );
  XOR3X1 U8618 ( .IN1(n8867), .IN2(n8868), .IN3(n8869), .Q(n8866) );
  XOR3X1 U8619 ( .IN1(n8861), .IN2(n8854), .IN3(n8870), .Q(n8869) );
  XOR2X1 U8620 ( .IN1(n8849), .IN2(n8842), .Q(n8870) );
  INVX0 U8621 ( .INP(n8871), .ZN(n8842) );
  NAND3X0 U8622 ( .IN1(n8872), .IN2(n8873), .IN3(n8874), .QN(n8871) );
  NAND2X0 U8623 ( .IN1(n8875), .IN2(n8876), .QN(n8873) );
  NAND2X0 U8624 ( .IN1(n8877), .IN2(n8878), .QN(n8872) );
  NAND3X0 U8625 ( .IN1(n8879), .IN2(n8880), .IN3(n8881), .QN(n8849) );
  NAND2X0 U8626 ( .IN1(n8882), .IN2(n8876), .QN(n8880) );
  NAND2X0 U8627 ( .IN1(n8877), .IN2(n8883), .QN(n8879) );
  NAND3X0 U8628 ( .IN1(n8884), .IN2(n8885), .IN3(n8874), .QN(n8854) );
  NAND2X0 U8629 ( .IN1(n8886), .IN2(n8887), .QN(n8885) );
  NAND2X0 U8630 ( .IN1(n8888), .IN2(n8889), .QN(n8884) );
  NAND3X0 U8631 ( .IN1(n8890), .IN2(n8891), .IN3(n8881), .QN(n8861) );
  NAND2X0 U8632 ( .IN1(n8892), .IN2(n8876), .QN(n8891) );
  NAND2X0 U8633 ( .IN1(n8877), .IN2(n8893), .QN(n8890) );
  XOR2X1 U8634 ( .IN1(n8829), .IN2(n8821), .Q(n8868) );
  INVX0 U8635 ( .INP(n8894), .ZN(n8821) );
  NAND3X0 U8636 ( .IN1(n8895), .IN2(n8896), .IN3(n8874), .QN(n8894) );
  NAND2X0 U8637 ( .IN1(n8897), .IN2(n8887), .QN(n8896) );
  NAND2X0 U8638 ( .IN1(n8888), .IN2(n8898), .QN(n8895) );
  NAND3X0 U8639 ( .IN1(n8899), .IN2(n8900), .IN3(n8874), .QN(n8829) );
  NAND2X0 U8640 ( .IN1(n8901), .IN2(n8887), .QN(n8900) );
  NAND2X0 U8641 ( .IN1(n8888), .IN2(n8902), .QN(n8899) );
  XOR2X1 U8642 ( .IN1(n8833), .IN2(n8837), .Q(n8867) );
  INVX0 U8643 ( .INP(n8903), .ZN(n8837) );
  NAND3X0 U8644 ( .IN1(n8904), .IN2(n8905), .IN3(n8874), .QN(n8903) );
  NAND2X0 U8645 ( .IN1(n8906), .IN2(n8876), .QN(n8905) );
  NAND2X0 U8646 ( .IN1(n8877), .IN2(n8907), .QN(n8904) );
  NOR3X0 U8647 ( .IN1(n8908), .IN2(n8909), .IN3(n8910), .QN(n8833) );
  NOR2X0 U8648 ( .IN1(n8911), .IN2(n8912), .QN(n8909) );
  INVX0 U8649 ( .INP(n8913), .ZN(n8908) );
  NAND2X0 U8650 ( .IN1(n8888), .IN2(n8911), .QN(n8913) );
  NAND4X0 U8651 ( .IN1(n8820), .IN2(n8823), .IN3(n8914), .IN4(n8915), .QN(
        n8864) );
  NAND2X0 U8652 ( .IN1(n14379), .IN2(n8798), .QN(n8915) );
  NAND2X0 U8653 ( .IN1(n4490), .IN2(g3229), .QN(n8914) );
  NOR2X0 U8654 ( .IN1(n8862), .IN2(n8822), .QN(n8823) );
  NAND2X0 U8655 ( .IN1(n8916), .IN2(g2631), .QN(n8863) );
  XOR2X1 U8656 ( .IN1(n8817), .IN2(n8845), .Q(n8916) );
  NAND3X0 U8657 ( .IN1(n8917), .IN2(n8918), .IN3(n8881), .QN(n8845) );
  INVX0 U8658 ( .INP(n8919), .ZN(n8881) );
  NAND2X0 U8659 ( .IN1(n8874), .IN2(n2351), .QN(n8919) );
  NAND2X0 U8660 ( .IN1(n8920), .IN2(n8876), .QN(n8918) );
  NAND2X0 U8661 ( .IN1(n8877), .IN2(n8921), .QN(n8917) );
  NOR2X0 U8662 ( .IN1(n8876), .IN2(n8922), .QN(n8877) );
  NAND3X0 U8663 ( .IN1(n8923), .IN2(n8924), .IN3(n8925), .QN(n8817) );
  INVX0 U8664 ( .INP(n8910), .ZN(n8925) );
  NAND2X0 U8665 ( .IN1(n8874), .IN2(n8926), .QN(n8910) );
  NAND2X0 U8666 ( .IN1(n8922), .IN2(n8887), .QN(n8926) );
  NOR2X0 U8667 ( .IN1(n8862), .IN2(n4543), .QN(n8874) );
  NAND2X0 U8668 ( .IN1(n8927), .IN2(n7761), .QN(n8862) );
  NOR2X0 U8669 ( .IN1(g2637), .IN2(g30072), .QN(n8927) );
  NAND2X0 U8670 ( .IN1(n8928), .IN2(n8887), .QN(n8924) );
  NAND2X0 U8671 ( .IN1(n8888), .IN2(n8929), .QN(n8923) );
  NOR2X0 U8672 ( .IN1(n8887), .IN2(n8922), .QN(n8888) );
  NAND2X0 U8673 ( .IN1(n8930), .IN2(n8931), .QN(n4249) );
  NAND2X0 U8674 ( .IN1(n2289), .IN2(n8932), .QN(n8931) );
  NAND3X0 U8675 ( .IN1(n8933), .IN2(n8934), .IN3(n8935), .QN(n8930) );
  NAND2X0 U8676 ( .IN1(n8936), .IN2(n8937), .QN(n8934) );
  NAND2X0 U8677 ( .IN1(n7158), .IN2(n8938), .QN(n8933) );
  NAND3X0 U8678 ( .IN1(n2275), .IN2(n8939), .IN3(n2303), .QN(n4248) );
  NAND3X0 U8679 ( .IN1(n8940), .IN2(n8941), .IN3(n8935), .QN(n8939) );
  NAND2X0 U8680 ( .IN1(n8942), .IN2(n8937), .QN(n8941) );
  INVX0 U8681 ( .INP(n8943), .ZN(n8942) );
  NAND2X0 U8682 ( .IN1(n8938), .IN2(DFF_1145_n1), .QN(n8940) );
  NAND2X0 U8683 ( .IN1(n2275), .IN2(n8944), .QN(n4247) );
  NAND3X0 U8684 ( .IN1(n8945), .IN2(n8946), .IN3(n8935), .QN(n8944) );
  NAND2X0 U8685 ( .IN1(n8947), .IN2(n8937), .QN(n8946) );
  NAND2X0 U8686 ( .IN1(n8938), .IN2(DFF_1149_n1), .QN(n8945) );
  NAND3X0 U8687 ( .IN1(n2275), .IN2(n8948), .IN3(n2303), .QN(n4246) );
  NAND3X0 U8688 ( .IN1(n8949), .IN2(n8950), .IN3(n8935), .QN(n8948) );
  NAND2X0 U8689 ( .IN1(n8951), .IN2(n8937), .QN(n8950) );
  NAND2X0 U8690 ( .IN1(n8938), .IN2(DFF_1146_n1), .QN(n8949) );
  NAND2X0 U8691 ( .IN1(n8952), .IN2(n8953), .QN(n4245) );
  NAND3X0 U8692 ( .IN1(n8954), .IN2(n8955), .IN3(n8935), .QN(n8953) );
  NAND2X0 U8693 ( .IN1(n8956), .IN2(n8937), .QN(n8955) );
  NAND2X0 U8694 ( .IN1(n8938), .IN2(DFF_1144_n1), .QN(n8954) );
  NAND2X0 U8695 ( .IN1(n8957), .IN2(n8958), .QN(n4244) );
  NAND2X0 U8696 ( .IN1(n2289), .IN2(n8959), .QN(n8958) );
  NAND3X0 U8697 ( .IN1(n8960), .IN2(n8961), .IN3(n8935), .QN(n8957) );
  NAND2X0 U8698 ( .IN1(n8962), .IN2(n8937), .QN(n8961) );
  INVX0 U8699 ( .INP(n8963), .ZN(n8962) );
  NAND2X0 U8700 ( .IN1(n7159), .IN2(n8938), .QN(n8960) );
  NAND2X0 U8701 ( .IN1(n8952), .IN2(n8964), .QN(n4243) );
  NAND3X0 U8702 ( .IN1(n8965), .IN2(n8966), .IN3(n8935), .QN(n8964) );
  NAND2X0 U8703 ( .IN1(n8967), .IN2(n8937), .QN(n8966) );
  INVX0 U8704 ( .INP(n8968), .ZN(n8967) );
  NAND2X0 U8705 ( .IN1(n8938), .IN2(DFF_1147_n1), .QN(n8965) );
  INVX0 U8706 ( .INP(n8969), .ZN(n8952) );
  NAND2X0 U8707 ( .IN1(n2275), .IN2(n8970), .QN(n8969) );
  NAND2X0 U8708 ( .IN1(n2289), .IN2(n2302), .QN(n8970) );
  NAND2X0 U8709 ( .IN1(n2275), .IN2(n8971), .QN(n4242) );
  NAND3X0 U8710 ( .IN1(n8972), .IN2(n8973), .IN3(n8935), .QN(n8971) );
  NAND2X0 U8711 ( .IN1(n8974), .IN2(n8937), .QN(n8973) );
  INVX0 U8712 ( .INP(n8975), .ZN(n8974) );
  NAND2X0 U8713 ( .IN1(n8938), .IN2(DFF_1148_n1), .QN(n8972) );
  NAND3X0 U8714 ( .IN1(n8976), .IN2(n8977), .IN3(n8978), .QN(n4241) );
  NAND2X0 U8715 ( .IN1(n8979), .IN2(g1890), .QN(n8978) );
  XOR3X1 U8716 ( .IN1(n8980), .IN2(n8981), .IN3(n8982), .Q(n8979) );
  XOR3X1 U8717 ( .IN1(n8975), .IN2(n8968), .IN3(n8983), .Q(n8982) );
  XOR2X1 U8718 ( .IN1(n8963), .IN2(n8956), .Q(n8983) );
  INVX0 U8719 ( .INP(n8984), .ZN(n8956) );
  NAND3X0 U8720 ( .IN1(n8985), .IN2(n8986), .IN3(n8987), .QN(n8984) );
  NAND2X0 U8721 ( .IN1(n8988), .IN2(n8989), .QN(n8986) );
  NAND2X0 U8722 ( .IN1(n8990), .IN2(n8991), .QN(n8985) );
  NAND3X0 U8723 ( .IN1(n8992), .IN2(n8993), .IN3(n8994), .QN(n8963) );
  NAND2X0 U8724 ( .IN1(n8995), .IN2(n8989), .QN(n8993) );
  NAND2X0 U8725 ( .IN1(n8990), .IN2(n8996), .QN(n8992) );
  NAND3X0 U8726 ( .IN1(n8997), .IN2(n8998), .IN3(n8987), .QN(n8968) );
  INVX0 U8727 ( .INP(n8999), .ZN(n8998) );
  NOR2X0 U8728 ( .IN1(n9000), .IN2(n9001), .QN(n8999) );
  NAND2X0 U8729 ( .IN1(n9002), .IN2(n9000), .QN(n8997) );
  NAND3X0 U8730 ( .IN1(n9003), .IN2(n9004), .IN3(n8994), .QN(n8975) );
  NAND2X0 U8731 ( .IN1(n9005), .IN2(n8989), .QN(n9004) );
  NAND2X0 U8732 ( .IN1(n8990), .IN2(n9006), .QN(n9003) );
  XOR2X1 U8733 ( .IN1(n8943), .IN2(n8936), .Q(n8981) );
  INVX0 U8734 ( .INP(n9007), .ZN(n8936) );
  NAND3X0 U8735 ( .IN1(n9008), .IN2(n9009), .IN3(n8987), .QN(n9007) );
  NAND2X0 U8736 ( .IN1(n9010), .IN2(n9011), .QN(n9009) );
  NAND2X0 U8737 ( .IN1(n9002), .IN2(n9012), .QN(n9008) );
  NAND3X0 U8738 ( .IN1(n9013), .IN2(n9014), .IN3(n8987), .QN(n8943) );
  NAND2X0 U8739 ( .IN1(n9015), .IN2(n9011), .QN(n9014) );
  NAND2X0 U8740 ( .IN1(n9002), .IN2(n9016), .QN(n9013) );
  XOR2X1 U8741 ( .IN1(n8947), .IN2(n8951), .Q(n8980) );
  INVX0 U8742 ( .INP(n9017), .ZN(n8951) );
  NAND3X0 U8743 ( .IN1(n9018), .IN2(n9019), .IN3(n8987), .QN(n9017) );
  NAND2X0 U8744 ( .IN1(n9020), .IN2(n8989), .QN(n9019) );
  NAND2X0 U8745 ( .IN1(n8990), .IN2(n9021), .QN(n9018) );
  NOR3X0 U8746 ( .IN1(n9022), .IN2(n9023), .IN3(n9024), .QN(n8947) );
  NOR2X0 U8747 ( .IN1(n9025), .IN2(n9001), .QN(n9023) );
  INVX0 U8748 ( .INP(n9026), .ZN(n9022) );
  NAND2X0 U8749 ( .IN1(n9002), .IN2(n9025), .QN(n9026) );
  NAND4X0 U8750 ( .IN1(n8935), .IN2(n8938), .IN3(n9027), .IN4(n9028), .QN(
        n8977) );
  NAND2X0 U8751 ( .IN1(g3229), .IN2(n8111), .QN(n9028) );
  NAND2X0 U8752 ( .IN1(n14380), .IN2(n8798), .QN(n9027) );
  NOR2X0 U8753 ( .IN1(n8559), .IN2(n8937), .QN(n8938) );
  NAND2X0 U8754 ( .IN1(n9029), .IN2(g1937), .QN(n8976) );
  XOR2X1 U8755 ( .IN1(n8932), .IN2(n8959), .Q(n9029) );
  NAND3X0 U8756 ( .IN1(n9030), .IN2(n9031), .IN3(n8994), .QN(n8959) );
  INVX0 U8757 ( .INP(n9032), .ZN(n8994) );
  NAND2X0 U8758 ( .IN1(n8987), .IN2(n9033), .QN(n9032) );
  NAND2X0 U8759 ( .IN1(n9034), .IN2(n8989), .QN(n9033) );
  NAND2X0 U8760 ( .IN1(n9035), .IN2(n8989), .QN(n9031) );
  NAND2X0 U8761 ( .IN1(n8990), .IN2(n9036), .QN(n9030) );
  NOR2X0 U8762 ( .IN1(n8989), .IN2(n9034), .QN(n8990) );
  NAND3X0 U8763 ( .IN1(n9037), .IN2(n9038), .IN3(n9039), .QN(n8932) );
  INVX0 U8764 ( .INP(n9024), .ZN(n9039) );
  NAND2X0 U8765 ( .IN1(n8987), .IN2(n9040), .QN(n9024) );
  NAND2X0 U8766 ( .IN1(n9034), .IN2(n9011), .QN(n9040) );
  NOR2X0 U8767 ( .IN1(n8559), .IN2(n4545), .QN(n8987) );
  NAND2X0 U8768 ( .IN1(n9041), .IN2(n7762), .QN(n8559) );
  NOR2X0 U8769 ( .IN1(g1943), .IN2(n516), .QN(n9041) );
  NAND2X0 U8770 ( .IN1(n9042), .IN2(n9011), .QN(n9038) );
  NAND2X0 U8771 ( .IN1(n9002), .IN2(n9043), .QN(n9037) );
  NOR2X0 U8772 ( .IN1(n9011), .IN2(n9034), .QN(n9002) );
  INVX0 U8773 ( .INP(n9044), .ZN(n9034) );
  NAND2X0 U8774 ( .IN1(n9045), .IN2(n9046), .QN(n4240) );
  NAND2X0 U8775 ( .IN1(n2217), .IN2(n9047), .QN(n9046) );
  NAND3X0 U8776 ( .IN1(n9048), .IN2(n9049), .IN3(n9050), .QN(n9045) );
  NAND2X0 U8777 ( .IN1(n9051), .IN2(n9052), .QN(n9049) );
  NAND2X0 U8778 ( .IN1(n7160), .IN2(n9053), .QN(n9048) );
  NAND3X0 U8779 ( .IN1(n9054), .IN2(n9055), .IN3(n2231), .QN(n4239) );
  NAND3X0 U8780 ( .IN1(n9056), .IN2(n9057), .IN3(n9050), .QN(n9054) );
  NAND2X0 U8781 ( .IN1(n9058), .IN2(n9052), .QN(n9057) );
  INVX0 U8782 ( .INP(n9059), .ZN(n9058) );
  NAND2X0 U8783 ( .IN1(n9053), .IN2(DFF_795_n1), .QN(n9056) );
  NAND2X0 U8784 ( .IN1(n9055), .IN2(n9060), .QN(n4238) );
  NAND3X0 U8785 ( .IN1(n9061), .IN2(n9062), .IN3(n9050), .QN(n9060) );
  NAND2X0 U8786 ( .IN1(n9063), .IN2(n9052), .QN(n9062) );
  NAND2X0 U8787 ( .IN1(n9053), .IN2(DFF_799_n1), .QN(n9061) );
  NAND3X0 U8788 ( .IN1(n9064), .IN2(n9055), .IN3(n2231), .QN(n4237) );
  NAND3X0 U8789 ( .IN1(n9065), .IN2(n9066), .IN3(n9050), .QN(n9064) );
  NAND2X0 U8790 ( .IN1(n9067), .IN2(n9052), .QN(n9066) );
  NAND2X0 U8791 ( .IN1(n9053), .IN2(DFF_796_n1), .QN(n9065) );
  NAND2X0 U8792 ( .IN1(n9068), .IN2(n9069), .QN(n4236) );
  NAND3X0 U8793 ( .IN1(n9070), .IN2(n9071), .IN3(n9050), .QN(n9069) );
  NAND2X0 U8794 ( .IN1(n9072), .IN2(n9052), .QN(n9071) );
  NAND2X0 U8795 ( .IN1(n9053), .IN2(DFF_794_n1), .QN(n9070) );
  NAND2X0 U8796 ( .IN1(n9073), .IN2(n9074), .QN(n4235) );
  NAND2X0 U8797 ( .IN1(n2217), .IN2(n9075), .QN(n9074) );
  NAND3X0 U8798 ( .IN1(n9076), .IN2(n9077), .IN3(n9050), .QN(n9073) );
  NAND2X0 U8799 ( .IN1(n9078), .IN2(n9052), .QN(n9077) );
  INVX0 U8800 ( .INP(n9079), .ZN(n9078) );
  NAND2X0 U8801 ( .IN1(n7161), .IN2(n9053), .QN(n9076) );
  NAND2X0 U8802 ( .IN1(n9068), .IN2(n9080), .QN(n4234) );
  NAND3X0 U8803 ( .IN1(n9081), .IN2(n9082), .IN3(n9050), .QN(n9080) );
  NAND2X0 U8804 ( .IN1(n9083), .IN2(n9052), .QN(n9082) );
  INVX0 U8805 ( .INP(n9084), .ZN(n9083) );
  NAND2X0 U8806 ( .IN1(n9053), .IN2(DFF_797_n1), .QN(n9081) );
  INVX0 U8807 ( .INP(n9085), .ZN(n9068) );
  NAND2X0 U8808 ( .IN1(n9055), .IN2(n9086), .QN(n9085) );
  NAND2X0 U8809 ( .IN1(n2217), .IN2(n2230), .QN(n9086) );
  NAND2X0 U8810 ( .IN1(n9055), .IN2(n9087), .QN(n4233) );
  NAND3X0 U8811 ( .IN1(n9088), .IN2(n9089), .IN3(n9050), .QN(n9087) );
  NAND2X0 U8812 ( .IN1(n9090), .IN2(n9052), .QN(n9089) );
  INVX0 U8813 ( .INP(n9091), .ZN(n9090) );
  NAND2X0 U8814 ( .IN1(n9053), .IN2(DFF_798_n1), .QN(n9088) );
  NAND2X0 U8815 ( .IN1(n2217), .IN2(n9092), .QN(n9055) );
  NAND3X0 U8816 ( .IN1(n9093), .IN2(n9094), .IN3(n9095), .QN(n4232) );
  NAND2X0 U8817 ( .IN1(n9096), .IN2(g1196), .QN(n9095) );
  XOR3X1 U8818 ( .IN1(n9097), .IN2(n9098), .IN3(n9099), .Q(n9096) );
  XOR3X1 U8819 ( .IN1(n9091), .IN2(n9084), .IN3(n9100), .Q(n9099) );
  XOR2X1 U8820 ( .IN1(n9079), .IN2(n9072), .Q(n9100) );
  INVX0 U8821 ( .INP(n9101), .ZN(n9072) );
  NAND3X0 U8822 ( .IN1(n9102), .IN2(n9103), .IN3(n9104), .QN(n9101) );
  NAND2X0 U8823 ( .IN1(n9105), .IN2(n9106), .QN(n9103) );
  NAND2X0 U8824 ( .IN1(n9107), .IN2(n9108), .QN(n9102) );
  NAND3X0 U8825 ( .IN1(n9109), .IN2(n9110), .IN3(n9111), .QN(n9079) );
  NAND2X0 U8826 ( .IN1(n9112), .IN2(n9106), .QN(n9110) );
  NAND2X0 U8827 ( .IN1(n9107), .IN2(n9113), .QN(n9109) );
  NAND3X0 U8828 ( .IN1(n9114), .IN2(n9115), .IN3(n9104), .QN(n9084) );
  NAND2X0 U8829 ( .IN1(n9116), .IN2(n9117), .QN(n9115) );
  NAND2X0 U8830 ( .IN1(n9118), .IN2(n9119), .QN(n9114) );
  NAND3X0 U8831 ( .IN1(n9120), .IN2(n9121), .IN3(n9111), .QN(n9091) );
  NAND2X0 U8832 ( .IN1(n9122), .IN2(n9106), .QN(n9121) );
  NAND2X0 U8833 ( .IN1(n9107), .IN2(n9123), .QN(n9120) );
  XOR2X1 U8834 ( .IN1(n9059), .IN2(n9051), .Q(n9098) );
  INVX0 U8835 ( .INP(n9124), .ZN(n9051) );
  NAND3X0 U8836 ( .IN1(n9125), .IN2(n9126), .IN3(n9104), .QN(n9124) );
  INVX0 U8837 ( .INP(n9127), .ZN(n9126) );
  NOR2X0 U8838 ( .IN1(n9128), .IN2(n9129), .QN(n9127) );
  NAND2X0 U8839 ( .IN1(n9118), .IN2(n9128), .QN(n9125) );
  NAND3X0 U8840 ( .IN1(n9130), .IN2(n9131), .IN3(n9104), .QN(n9059) );
  NAND2X0 U8841 ( .IN1(n9132), .IN2(n9117), .QN(n9131) );
  NAND2X0 U8842 ( .IN1(n9118), .IN2(n9133), .QN(n9130) );
  XOR2X1 U8843 ( .IN1(n9063), .IN2(n9067), .Q(n9097) );
  INVX0 U8844 ( .INP(n9134), .ZN(n9067) );
  NAND3X0 U8845 ( .IN1(n9135), .IN2(n9136), .IN3(n9104), .QN(n9134) );
  NAND2X0 U8846 ( .IN1(n9137), .IN2(n9106), .QN(n9136) );
  NAND2X0 U8847 ( .IN1(n9107), .IN2(n9138), .QN(n9135) );
  NOR3X0 U8848 ( .IN1(n9139), .IN2(n9140), .IN3(n9141), .QN(n9063) );
  NOR2X0 U8849 ( .IN1(n9142), .IN2(n9129), .QN(n9140) );
  INVX0 U8850 ( .INP(n9143), .ZN(n9139) );
  NAND2X0 U8851 ( .IN1(n9118), .IN2(n9142), .QN(n9143) );
  NAND4X0 U8852 ( .IN1(n9050), .IN2(n9053), .IN3(n9144), .IN4(n9145), .QN(
        n9094) );
  NAND2X0 U8853 ( .IN1(n4489), .IN2(g3229), .QN(n9145) );
  NAND2X0 U8854 ( .IN1(n8798), .IN2(n14381), .QN(n9144) );
  NOR2X0 U8855 ( .IN1(n9092), .IN2(n9052), .QN(n9053) );
  NAND2X0 U8856 ( .IN1(n9146), .IN2(g1243), .QN(n9093) );
  XOR2X1 U8857 ( .IN1(n9047), .IN2(n9075), .Q(n9146) );
  NAND3X0 U8858 ( .IN1(n9147), .IN2(n9148), .IN3(n9111), .QN(n9075) );
  INVX0 U8859 ( .INP(n9149), .ZN(n9111) );
  NAND2X0 U8860 ( .IN1(n9104), .IN2(n9150), .QN(n9149) );
  NAND2X0 U8861 ( .IN1(n9151), .IN2(n9106), .QN(n9150) );
  NAND2X0 U8862 ( .IN1(n9152), .IN2(n9106), .QN(n9148) );
  NAND2X0 U8863 ( .IN1(n9107), .IN2(n9153), .QN(n9147) );
  NOR2X0 U8864 ( .IN1(n9106), .IN2(n9151), .QN(n9107) );
  NAND3X0 U8865 ( .IN1(n9154), .IN2(n9155), .IN3(n9156), .QN(n9047) );
  INVX0 U8866 ( .INP(n9141), .ZN(n9156) );
  NAND2X0 U8867 ( .IN1(n9104), .IN2(n9157), .QN(n9141) );
  NAND2X0 U8868 ( .IN1(n9151), .IN2(n9117), .QN(n9157) );
  NOR2X0 U8869 ( .IN1(n9092), .IN2(n4548), .QN(n9104) );
  NAND2X0 U8870 ( .IN1(n9158), .IN2(n7763), .QN(n9092) );
  NOR2X0 U8871 ( .IN1(g1249), .IN2(n517), .QN(n9158) );
  NAND2X0 U8872 ( .IN1(n9159), .IN2(n9117), .QN(n9155) );
  NAND2X0 U8873 ( .IN1(n9118), .IN2(n9160), .QN(n9154) );
  NOR2X0 U8874 ( .IN1(n9117), .IN2(n9151), .QN(n9118) );
  INVX0 U8875 ( .INP(n9161), .ZN(n9151) );
  INVX0 U8876 ( .INP(n9162), .ZN(n3938) );
  NAND2X0 U8877 ( .IN1(n3896), .IN2(g88), .QN(n4528) );
  NAND2X0 U8878 ( .IN1(n3890), .IN2(g1462), .QN(n4527) );
  NAND2X0 U8879 ( .IN1(n3887), .IN2(test_so78), .QN(n4526) );
  NAND2X0 U8880 ( .IN1(n3692), .IN2(test_so15), .QN(n4521) );
  NAND2X0 U8881 ( .IN1(n3686), .IN2(g1453), .QN(n4523) );
  NAND2X0 U8882 ( .IN1(n3683), .IN2(g2147), .QN(n4522) );
  INVX0 U8883 ( .INP(n9163), .ZN(n328) );
  NAND2X0 U8884 ( .IN1(n9164), .IN2(n9165), .QN(n3254) );
  NAND2X0 U8885 ( .IN1(n9166), .IN2(n9167), .QN(n9164) );
  INVX0 U8886 ( .INP(n9168), .ZN(n9166) );
  NAND4X0 U8887 ( .IN1(n9169), .IN2(n9170), .IN3(n9171), .IN4(g309), .QN(n3023) );
  INVX0 U8888 ( .INP(n9172), .ZN(n9171) );
  NAND4X0 U8889 ( .IN1(n9173), .IN2(n9174), .IN3(n9175), .IN4(g996), .QN(n3016) );
  INVX0 U8890 ( .INP(n9176), .ZN(n9175) );
  NAND4X0 U8891 ( .IN1(n9177), .IN2(n9178), .IN3(n9179), .IN4(g1690), .QN(
        n3008) );
  INVX0 U8892 ( .INP(n9180), .ZN(n9179) );
  NAND4X0 U8893 ( .IN1(test_so79), .IN2(n9181), .IN3(n9182), .IN4(n9183), .QN(
        n3000) );
  INVX0 U8894 ( .INP(n9184), .ZN(n9183) );
  INVX0 U8895 ( .INP(g24734), .ZN(n298) );
  INVX0 U8896 ( .INP(g25435), .ZN(n289) );
  XOR2X1 U8897 ( .IN1(n9185), .IN2(n9186), .Q(n2800) );
  NAND2X0 U8898 ( .IN1(n9187), .IN2(n9188), .QN(n9185) );
  NAND2X0 U8899 ( .IN1(n9186), .IN2(n9189), .QN(n9188) );
  NAND3X0 U8900 ( .IN1(n9190), .IN2(n9191), .IN3(n9192), .QN(n9189) );
  NAND2X0 U8901 ( .IN1(n9193), .IN2(n9194), .QN(n9191) );
  NAND3X0 U8902 ( .IN1(n9195), .IN2(g996), .IN3(n9196), .QN(n9190) );
  NAND3X0 U8903 ( .IN1(n9197), .IN2(n9192), .IN3(n9198), .QN(n9187) );
  XOR2X1 U8904 ( .IN1(n8584), .IN2(n9199), .Q(n2719) );
  XOR2X1 U8905 ( .IN1(n9200), .IN2(n9201), .Q(n2686) );
  XOR2X1 U8906 ( .IN1(n8678), .IN2(n9202), .Q(n2671) );
  INVX0 U8907 ( .INP(g26135), .ZN(n263) );
  XOR2X1 U8908 ( .IN1(n9194), .IN2(n9203), .Q(n2616) );
  NAND2X0 U8909 ( .IN1(n9204), .IN2(n9205), .QN(n9203) );
  NAND2X0 U8910 ( .IN1(n9206), .IN2(n9207), .QN(n9205) );
  NAND4X0 U8911 ( .IN1(n9208), .IN2(n9209), .IN3(n9210), .IN4(n9192), .QN(
        n9204) );
  NAND3X0 U8912 ( .IN1(n9186), .IN2(n9211), .IN3(n9197), .QN(n9210) );
  INVX0 U8913 ( .INP(n9212), .ZN(n9197) );
  NAND3X0 U8914 ( .IN1(n9213), .IN2(n9194), .IN3(n3102), .QN(n9212) );
  NAND2X0 U8915 ( .IN1(n9214), .IN2(n9194), .QN(n9209) );
  NAND2X0 U8916 ( .IN1(n9215), .IN2(n9196), .QN(n9208) );
  NAND2X0 U8917 ( .IN1(n9216), .IN2(n9217), .QN(n9215) );
  NAND2X0 U8918 ( .IN1(n9186), .IN2(n9218), .QN(n9217) );
  NAND3X0 U8919 ( .IN1(n9219), .IN2(n9211), .IN3(n9220), .QN(n9218) );
  INVX0 U8920 ( .INP(n9193), .ZN(n9220) );
  NAND2X0 U8921 ( .IN1(n9221), .IN2(n9222), .QN(n9193) );
  NAND2X0 U8922 ( .IN1(n9223), .IN2(n3102), .QN(n9222) );
  INVX0 U8923 ( .INP(n9213), .ZN(n9223) );
  NAND2X0 U8924 ( .IN1(n9224), .IN2(n9225), .QN(n9219) );
  NAND2X0 U8925 ( .IN1(n9226), .IN2(n9198), .QN(n9216) );
  NAND2X0 U8926 ( .IN1(n2632), .IN2(n9221), .QN(n9226) );
  NOR2X0 U8927 ( .IN1(n8696), .IN2(n8694), .QN(n2446) );
  NOR2X0 U8928 ( .IN1(g557), .IN2(n9227), .QN(n8694) );
  INVX0 U8929 ( .INP(n9228), .ZN(n9227) );
  NAND2X0 U8930 ( .IN1(n8054), .IN2(n8108), .QN(n9228) );
  NAND2X0 U8931 ( .IN1(n8108), .IN2(n9229), .QN(n8696) );
  NAND2X0 U8932 ( .IN1(n4360), .IN2(n8054), .QN(n9229) );
  NAND2X0 U8933 ( .IN1(g499), .IN2(n9230), .QN(n2445) );
  NAND4X0 U8934 ( .IN1(n9231), .IN2(n9232), .IN3(n9233), .IN4(n9234), .QN(
        n9230) );
  NAND2X0 U8935 ( .IN1(n7513), .IN2(g629), .QN(n9233) );
  NAND2X0 U8936 ( .IN1(n7509), .IN2(g6677), .QN(n9232) );
  NAND2X0 U8937 ( .IN1(n7508), .IN2(g6911), .QN(n9231) );
  NAND2X0 U8938 ( .IN1(n8804), .IN2(n8758), .QN(n2430) );
  INVX0 U8939 ( .INP(n9234), .ZN(n8804) );
  NAND4X0 U8940 ( .IN1(n9235), .IN2(n8781), .IN3(n9236), .IN4(n9237), .QN(
        n9234) );
  NOR4X0 U8941 ( .IN1(n9238), .IN2(n8760), .IN3(n8795), .IN4(n8766), .QN(n9237) );
  NAND3X0 U8942 ( .IN1(n8770), .IN2(n9239), .IN3(n8790), .QN(n9238) );
  NAND3X0 U8943 ( .IN1(n9240), .IN2(n9241), .IN3(n9242), .QN(n9239) );
  NAND2X0 U8944 ( .IN1(n7977), .IN2(g6911), .QN(n9242) );
  NAND2X0 U8945 ( .IN1(n7989), .IN2(g629), .QN(n9241) );
  NAND2X0 U8946 ( .IN1(n7880), .IN2(g6677), .QN(n9240) );
  NOR3X0 U8947 ( .IN1(n8775), .IN2(n8785), .IN3(n9243), .QN(n9236) );
  NOR2X0 U8948 ( .IN1(n8813), .IN2(n8805), .QN(n9235) );
  INVX0 U8949 ( .INP(n8814), .ZN(n8813) );
  NAND2X0 U8950 ( .IN1(g2574), .IN2(n9244), .QN(n2374) );
  NAND4X0 U8951 ( .IN1(n9245), .IN2(n9246), .IN3(n9247), .IN4(n9248), .QN(
        n9244) );
  NAND2X0 U8952 ( .IN1(n7510), .IN2(g2703), .QN(n9247) );
  NAND2X0 U8953 ( .IN1(n7503), .IN2(g7425), .QN(n9246) );
  NAND2X0 U8954 ( .IN1(n7502), .IN2(g7487), .QN(n9245) );
  NOR2X0 U8955 ( .IN1(n8822), .IN2(n8820), .QN(n2361) );
  NOR2X0 U8956 ( .IN1(g2631), .IN2(n9249), .QN(n8820) );
  INVX0 U8957 ( .INP(n9250), .ZN(n9249) );
  NAND2X0 U8958 ( .IN1(n8067), .IN2(n4303), .QN(n9250) );
  NAND2X0 U8959 ( .IN1(n4303), .IN2(n9251), .QN(n8822) );
  NAND2X0 U8960 ( .IN1(n4352), .IN2(n8067), .QN(n9251) );
  NAND2X0 U8961 ( .IN1(n8922), .IN2(n8876), .QN(n2351) );
  INVX0 U8962 ( .INP(n9248), .ZN(n8922) );
  NAND4X0 U8963 ( .IN1(n9252), .IN2(n8911), .IN3(n9253), .IN4(n9254), .QN(
        n9248) );
  NOR4X0 U8964 ( .IN1(n9255), .IN2(n8907), .IN3(n8878), .IN4(n8902), .QN(n9254) );
  NAND3X0 U8965 ( .IN1(n8886), .IN2(n9256), .IN3(n8897), .QN(n9255) );
  NAND3X0 U8966 ( .IN1(n9257), .IN2(n9258), .IN3(n9259), .QN(n9256) );
  NAND2X0 U8967 ( .IN1(n7974), .IN2(g7487), .QN(n9259) );
  NAND2X0 U8968 ( .IN1(g2703), .IN2(n8116), .QN(n9258) );
  NAND2X0 U8969 ( .IN1(n7877), .IN2(g7425), .QN(n9257) );
  NOR3X0 U8970 ( .IN1(n8892), .IN2(n8928), .IN3(n9260), .QN(n9253) );
  NOR2X0 U8971 ( .IN1(n8920), .IN2(n8882), .QN(n9252) );
  INVX0 U8972 ( .INP(n8921), .ZN(n8920) );
  NAND2X0 U8973 ( .IN1(g1880), .IN2(n9261), .QN(n2302) );
  NAND4X0 U8974 ( .IN1(n9262), .IN2(n9263), .IN3(n9264), .IN4(n9044), .QN(
        n9261) );
  NAND4X0 U8975 ( .IN1(n9265), .IN2(n9025), .IN3(n9266), .IN4(n9267), .QN(
        n9044) );
  NOR4X0 U8976 ( .IN1(n9268), .IN2(n9012), .IN3(n9000), .IN4(n9021), .QN(n9267) );
  NAND3X0 U8977 ( .IN1(n9015), .IN2(n9269), .IN3(n8988), .QN(n9268) );
  NAND3X0 U8978 ( .IN1(n9270), .IN2(n9271), .IN3(n9272), .QN(n9269) );
  NAND2X0 U8979 ( .IN1(n7975), .IN2(g7357), .QN(n9272) );
  NAND2X0 U8980 ( .IN1(n7981), .IN2(g2009), .QN(n9271) );
  NAND2X0 U8981 ( .IN1(n7878), .IN2(g7229), .QN(n9270) );
  INVX0 U8982 ( .INP(n9016), .ZN(n9015) );
  NOR3X0 U8983 ( .IN1(n9005), .IN2(n9042), .IN3(n9273), .QN(n9266) );
  NOR2X0 U8984 ( .IN1(n9035), .IN2(n8995), .QN(n9265) );
  INVX0 U8985 ( .INP(n9036), .ZN(n9035) );
  NAND2X0 U8986 ( .IN1(n7511), .IN2(g2009), .QN(n9264) );
  NAND2X0 U8987 ( .IN1(n7505), .IN2(g7229), .QN(n9263) );
  NAND2X0 U8988 ( .IN1(n7504), .IN2(g7357), .QN(n9262) );
  NOR2X0 U8989 ( .IN1(n8937), .IN2(n8935), .QN(n2289) );
  NOR2X0 U8990 ( .IN1(g1937), .IN2(n9274), .QN(n8935) );
  INVX0 U8991 ( .INP(n9275), .ZN(n9274) );
  NAND2X0 U8992 ( .IN1(n8064), .IN2(n4297), .QN(n9275) );
  NAND2X0 U8993 ( .IN1(n4297), .IN2(n9276), .QN(n8937) );
  NAND2X0 U8994 ( .IN1(n4311), .IN2(n8064), .QN(n9276) );
  NAND2X0 U8995 ( .IN1(g1186), .IN2(n9277), .QN(n2230) );
  NAND4X0 U8996 ( .IN1(n9278), .IN2(n9279), .IN3(n9280), .IN4(n9161), .QN(
        n9277) );
  NAND4X0 U8997 ( .IN1(n9281), .IN2(n9142), .IN3(n9282), .IN4(n9283), .QN(
        n9161) );
  NOR4X0 U8998 ( .IN1(n9284), .IN2(n9128), .IN3(n9119), .IN4(n9138), .QN(n9283) );
  NAND3X0 U8999 ( .IN1(n9132), .IN2(n9285), .IN3(n9105), .QN(n9284) );
  NAND3X0 U9000 ( .IN1(n9286), .IN2(n9287), .IN3(n9288), .QN(n9285) );
  NAND2X0 U9001 ( .IN1(n7976), .IN2(g7161), .QN(n9288) );
  NAND2X0 U9002 ( .IN1(n7982), .IN2(g1315), .QN(n9287) );
  NAND2X0 U9003 ( .IN1(n7879), .IN2(g6979), .QN(n9286) );
  INVX0 U9004 ( .INP(n9133), .ZN(n9132) );
  NOR3X0 U9005 ( .IN1(n9122), .IN2(n9159), .IN3(n9289), .QN(n9282) );
  NOR2X0 U9006 ( .IN1(n9152), .IN2(n9112), .QN(n9281) );
  NAND2X0 U9007 ( .IN1(n7512), .IN2(g1315), .QN(n9280) );
  NAND2X0 U9008 ( .IN1(n7507), .IN2(g6979), .QN(n9279) );
  NAND2X0 U9009 ( .IN1(n7506), .IN2(g7161), .QN(n9278) );
  INVX0 U9010 ( .INP(n9290), .ZN(n223) );
  NOR2X0 U9011 ( .IN1(n9052), .IN2(n9050), .QN(n2217) );
  NOR2X0 U9012 ( .IN1(g1243), .IN2(n9291), .QN(n9050) );
  INVX0 U9013 ( .INP(n9292), .ZN(n9291) );
  NAND2X0 U9014 ( .IN1(n8063), .IN2(n4304), .QN(n9292) );
  NAND2X0 U9015 ( .IN1(n4304), .IN2(n9293), .QN(n9052) );
  NAND2X0 U9016 ( .IN1(n4353), .IN2(n8063), .QN(n9293) );
  INVX0 U9017 ( .INP(n9294), .ZN(n184) );
  INVX0 U9018 ( .INP(n9295), .ZN(n162) );
  INVX0 U9019 ( .INP(n9296), .ZN(n1544) );
  NAND3X0 U9020 ( .IN1(n9297), .IN2(n1547), .IN3(n8741), .QN(n9296) );
  NAND2X0 U9021 ( .IN1(n9298), .IN2(n4350), .QN(n9297) );
  NAND2X0 U9022 ( .IN1(g3018), .IN2(n8742), .QN(n9298) );
  INVX0 U9023 ( .INP(n9299), .ZN(n1542) );
  NAND3X0 U9024 ( .IN1(n9300), .IN2(n4066), .IN3(n9301), .QN(n9299) );
  NAND2X0 U9025 ( .IN1(n9302), .IN2(n8053), .QN(n9301) );
  NAND2X0 U9026 ( .IN1(n7909), .IN2(n9303), .QN(n9302) );
  INVX0 U9027 ( .INP(n9304), .ZN(n1507) );
  NAND3X0 U9028 ( .IN1(n9305), .IN2(n9306), .IN3(n9307), .QN(n9304) );
  NAND2X0 U9029 ( .IN1(n9308), .IN2(n4407), .QN(n9305) );
  NAND2X0 U9030 ( .IN1(g2734), .IN2(n9309), .QN(n9308) );
  INVX0 U9031 ( .INP(n9310), .ZN(n1506) );
  NAND3X0 U9032 ( .IN1(n9311), .IN2(n9306), .IN3(n9312), .QN(n9310) );
  NAND2X0 U9033 ( .IN1(n9313), .IN2(n4472), .QN(n9311) );
  NAND2X0 U9034 ( .IN1(g2714), .IN2(n9314), .QN(n9313) );
  INVX0 U9035 ( .INP(n9315), .ZN(n1431) );
  NOR2X0 U9036 ( .IN1(n9316), .IN2(n9317), .QN(n9315) );
  NOR2X0 U9037 ( .IN1(g2624), .IN2(n7990), .QN(n9317) );
  INVX0 U9038 ( .INP(n9318), .ZN(n1427) );
  INVX0 U9039 ( .INP(n9319), .ZN(n1406) );
  INVX0 U9040 ( .INP(n9320), .ZN(n1269) );
  INVX0 U9041 ( .INP(n9321), .ZN(n123) );
  NOR3X0 U9042 ( .IN1(n9322), .IN2(n9323), .IN3(n9324), .QN(n1223) );
  NOR2X0 U9043 ( .IN1(n9325), .IN2(g2052), .QN(n9322) );
  NOR2X0 U9044 ( .IN1(n4399), .IN2(n9326), .QN(n9325) );
  INVX0 U9045 ( .INP(n9327), .ZN(n1222) );
  NAND3X0 U9046 ( .IN1(n9328), .IN2(n9329), .IN3(n9330), .QN(n9327) );
  NAND2X0 U9047 ( .IN1(n9331), .IN2(n4474), .QN(n9328) );
  NAND2X0 U9048 ( .IN1(g2020), .IN2(n9332), .QN(n9331) );
  NOR2X0 U9049 ( .IN1(n9323), .IN2(n9333), .QN(n1194) );
  INVX0 U9050 ( .INP(n9334), .ZN(n9333) );
  NAND2X0 U9051 ( .IN1(n9335), .IN2(n7975), .QN(n9334) );
  INVX0 U9052 ( .INP(n9336), .ZN(n1149) );
  NOR2X0 U9053 ( .IN1(n9337), .IN2(n9338), .QN(n9336) );
  NOR2X0 U9054 ( .IN1(g1930), .IN2(n7991), .QN(n9338) );
  INVX0 U9055 ( .INP(n9339), .ZN(n1145) );
  INVX0 U9056 ( .INP(n9340), .ZN(n1122) );
  INVX0 U9057 ( .INP(g27380), .ZN(n102) );
  NAND2X0 U9058 ( .IN1(n9341), .IN2(n9342), .QN(g30801) );
  INVX0 U9059 ( .INP(n9343), .ZN(n9342) );
  NOR2X0 U9060 ( .IN1(g3109), .IN2(n4334), .QN(n9343) );
  NAND2X0 U9061 ( .IN1(g30072), .IN2(g3109), .QN(n9341) );
  NAND2X0 U9062 ( .IN1(n9344), .IN2(n9345), .QN(g30798) );
  NAND2X0 U9063 ( .IN1(n4383), .IN2(g3107), .QN(n9345) );
  NAND2X0 U9064 ( .IN1(g30072), .IN2(g8030), .QN(n9344) );
  NAND2X0 U9065 ( .IN1(n9346), .IN2(n9347), .QN(g30796) );
  NAND2X0 U9066 ( .IN1(n4382), .IN2(g3106), .QN(n9347) );
  NAND2X0 U9067 ( .IN1(g30072), .IN2(g8106), .QN(n9346) );
  NAND2X0 U9068 ( .IN1(n9348), .IN2(n9349), .QN(g30709) );
  NAND2X0 U9069 ( .IN1(n9350), .IN2(g7264), .QN(n9349) );
  NAND2X0 U9070 ( .IN1(n4524), .IN2(g2391), .QN(n9348) );
  NAND2X0 U9071 ( .IN1(n9351), .IN2(n9352), .QN(g30708) );
  NAND2X0 U9072 ( .IN1(n9353), .IN2(n4618), .QN(n9352) );
  NAND2X0 U9073 ( .IN1(n4511), .IN2(g1698), .QN(n9351) );
  NAND2X0 U9074 ( .IN1(n9354), .IN2(n9355), .QN(g30707) );
  NAND2X0 U9075 ( .IN1(n9350), .IN2(g5555), .QN(n9355) );
  NAND2X0 U9076 ( .IN1(n4516), .IN2(g2390), .QN(n9354) );
  NAND2X0 U9077 ( .IN1(n9356), .IN2(n9357), .QN(g30706) );
  NAND2X0 U9078 ( .IN1(n9353), .IN2(g7014), .QN(n9357) );
  NAND2X0 U9079 ( .IN1(n4525), .IN2(g1697), .QN(n9356) );
  NAND2X0 U9080 ( .IN1(n9358), .IN2(n9359), .QN(g30705) );
  NAND2X0 U9081 ( .IN1(n4381), .IN2(g1004), .QN(n9359) );
  NAND2X0 U9082 ( .IN1(n2594), .IN2(g1088), .QN(n9358) );
  NAND2X0 U9083 ( .IN1(n9360), .IN2(n9361), .QN(g30704) );
  NAND2X0 U9084 ( .IN1(n9353), .IN2(g5511), .QN(n9361) );
  INVX0 U9085 ( .INP(n9362), .ZN(n9353) );
  NAND2X0 U9086 ( .IN1(n9363), .IN2(n9364), .QN(n9362) );
  XOR2X1 U9087 ( .IN1(n9365), .IN2(n9366), .Q(n9363) );
  NAND2X0 U9088 ( .IN1(n9367), .IN2(n9368), .QN(n9366) );
  NAND2X0 U9089 ( .IN1(n9369), .IN2(n9370), .QN(n9368) );
  NAND4X0 U9090 ( .IN1(n9371), .IN2(n9372), .IN3(n9373), .IN4(n9374), .QN(
        n9367) );
  NAND3X0 U9091 ( .IN1(n9375), .IN2(n9376), .IN3(n9377), .QN(n9373) );
  NAND2X0 U9092 ( .IN1(n9378), .IN2(n9365), .QN(n9372) );
  INVX0 U9093 ( .INP(n9379), .ZN(n9378) );
  NAND2X0 U9094 ( .IN1(n9380), .IN2(n9381), .QN(n9371) );
  NAND2X0 U9095 ( .IN1(n9382), .IN2(n9383), .QN(n9380) );
  NAND2X0 U9096 ( .IN1(n9375), .IN2(n9384), .QN(n9383) );
  NAND3X0 U9097 ( .IN1(n9385), .IN2(n9376), .IN3(n9386), .QN(n9384) );
  INVX0 U9098 ( .INP(n9387), .ZN(n9386) );
  NAND3X0 U9099 ( .IN1(n9388), .IN2(n9379), .IN3(n9389), .QN(n9385) );
  NAND2X0 U9100 ( .IN1(n9390), .IN2(n9391), .QN(n9382) );
  NAND2X0 U9101 ( .IN1(n9392), .IN2(n9393), .QN(n9390) );
  NAND2X0 U9102 ( .IN1(n9389), .IN2(n9388), .QN(n9392) );
  NAND2X0 U9103 ( .IN1(n4518), .IN2(g1696), .QN(n9360) );
  NAND2X0 U9104 ( .IN1(n9394), .IN2(n9395), .QN(g30703) );
  NAND2X0 U9105 ( .IN1(n4364), .IN2(g1003), .QN(n9395) );
  NAND2X0 U9106 ( .IN1(n2594), .IN2(g6712), .QN(n9394) );
  NAND2X0 U9107 ( .IN1(n9396), .IN2(n9397), .QN(g30702) );
  NAND2X0 U9108 ( .IN1(n9398), .IN2(n4640), .QN(n9397) );
  NAND2X0 U9109 ( .IN1(n4506), .IN2(g317), .QN(n9396) );
  NAND2X0 U9110 ( .IN1(n9399), .IN2(n9400), .QN(g30701) );
  NAND2X0 U9111 ( .IN1(n4363), .IN2(g1002), .QN(n9400) );
  NAND2X0 U9112 ( .IN1(n2594), .IN2(g5472), .QN(n9399) );
  NAND2X0 U9113 ( .IN1(n9401), .IN2(n9402), .QN(g30700) );
  NAND2X0 U9114 ( .IN1(n9398), .IN2(g6447), .QN(n9402) );
  NAND2X0 U9115 ( .IN1(test_so18), .IN2(n4499), .QN(n9401) );
  NAND2X0 U9116 ( .IN1(n9403), .IN2(n9404), .QN(g30699) );
  NAND2X0 U9117 ( .IN1(n9398), .IN2(g5437), .QN(n9404) );
  INVX0 U9118 ( .INP(n9405), .ZN(n9398) );
  NAND2X0 U9119 ( .IN1(n9406), .IN2(n9407), .QN(n9405) );
  XOR2X1 U9120 ( .IN1(n9408), .IN2(n9409), .Q(n9406) );
  NAND2X0 U9121 ( .IN1(n9410), .IN2(n9411), .QN(n9409) );
  NAND2X0 U9122 ( .IN1(n9412), .IN2(n9413), .QN(n9411) );
  NAND4X0 U9123 ( .IN1(n9414), .IN2(n9415), .IN3(n9416), .IN4(n9417), .QN(
        n9410) );
  NAND3X0 U9124 ( .IN1(n9418), .IN2(n9419), .IN3(n9420), .QN(n9416) );
  NAND2X0 U9125 ( .IN1(n9421), .IN2(n9408), .QN(n9415) );
  INVX0 U9126 ( .INP(n9422), .ZN(n9421) );
  NAND2X0 U9127 ( .IN1(n9423), .IN2(n9424), .QN(n9414) );
  NAND2X0 U9128 ( .IN1(n9425), .IN2(n9426), .QN(n9423) );
  NAND2X0 U9129 ( .IN1(n9418), .IN2(n9427), .QN(n9426) );
  NAND3X0 U9130 ( .IN1(n9428), .IN2(n9419), .IN3(n9429), .QN(n9427) );
  INVX0 U9131 ( .INP(n9430), .ZN(n9429) );
  NAND3X0 U9132 ( .IN1(n9431), .IN2(n9422), .IN3(n9432), .QN(n9428) );
  NAND2X0 U9133 ( .IN1(n9433), .IN2(n9434), .QN(n9425) );
  NAND2X0 U9134 ( .IN1(n9435), .IN2(n9436), .QN(n9433) );
  NAND2X0 U9135 ( .IN1(n9432), .IN2(n9431), .QN(n9435) );
  NAND2X0 U9136 ( .IN1(n4520), .IN2(g315), .QN(n9403) );
  NAND2X0 U9137 ( .IN1(n9437), .IN2(n9438), .QN(g30695) );
  NAND2X0 U9138 ( .IN1(n4367), .IN2(g2276), .QN(n9438) );
  NAND2X0 U9139 ( .IN1(n9439), .IN2(g2241), .QN(n9437) );
  NAND2X0 U9140 ( .IN1(n9440), .IN2(n9441), .QN(g30694) );
  NAND2X0 U9141 ( .IN1(n4367), .IN2(g2348), .QN(n9441) );
  NAND2X0 U9142 ( .IN1(n9442), .IN2(g2241), .QN(n9440) );
  NAND2X0 U9143 ( .IN1(n9443), .IN2(n9444), .QN(g30693) );
  NAND2X0 U9144 ( .IN1(g2273), .IN2(n8097), .QN(n9444) );
  NAND2X0 U9145 ( .IN1(test_so73), .IN2(n9439), .QN(n9443) );
  NAND2X0 U9146 ( .IN1(n9445), .IN2(n9446), .QN(g30692) );
  NAND2X0 U9147 ( .IN1(n4368), .IN2(g1582), .QN(n9446) );
  NAND2X0 U9148 ( .IN1(n9447), .IN2(g1547), .QN(n9445) );
  NAND2X0 U9149 ( .IN1(n9448), .IN2(n9449), .QN(g30691) );
  NAND2X0 U9150 ( .IN1(g2345), .IN2(n8097), .QN(n9449) );
  NAND2X0 U9151 ( .IN1(n9442), .IN2(test_so73), .QN(n9448) );
  NAND2X0 U9152 ( .IN1(n9450), .IN2(n9451), .QN(g30690) );
  NAND2X0 U9153 ( .IN1(n4324), .IN2(g2270), .QN(n9451) );
  NAND2X0 U9154 ( .IN1(n9439), .IN2(g6837), .QN(n9450) );
  NAND3X0 U9155 ( .IN1(n9452), .IN2(n9453), .IN3(n9454), .QN(n9439) );
  NAND2X0 U9156 ( .IN1(n9455), .IN2(n9456), .QN(n9453) );
  XOR2X1 U9157 ( .IN1(n9457), .IN2(n9458), .Q(n9455) );
  NAND2X0 U9158 ( .IN1(n9459), .IN2(g2175), .QN(n9452) );
  NAND2X0 U9159 ( .IN1(n9460), .IN2(n9461), .QN(g30689) );
  NAND2X0 U9160 ( .IN1(n4368), .IN2(g1654), .QN(n9461) );
  NAND2X0 U9161 ( .IN1(n9462), .IN2(g1547), .QN(n9460) );
  NAND2X0 U9162 ( .IN1(n9463), .IN2(n9464), .QN(g30688) );
  NAND2X0 U9163 ( .IN1(n4515), .IN2(g1579), .QN(n9464) );
  NAND2X0 U9164 ( .IN1(n9447), .IN2(g6782), .QN(n9463) );
  NAND2X0 U9165 ( .IN1(n9465), .IN2(n9466), .QN(g30687) );
  NAND2X0 U9166 ( .IN1(g888), .IN2(n8096), .QN(n9466) );
  NAND2X0 U9167 ( .IN1(test_so31), .IN2(n9467), .QN(n9465) );
  NAND2X0 U9168 ( .IN1(n9468), .IN2(n9469), .QN(g30686) );
  NAND2X0 U9169 ( .IN1(n4324), .IN2(g2342), .QN(n9469) );
  NAND2X0 U9170 ( .IN1(n9442), .IN2(g6837), .QN(n9468) );
  INVX0 U9171 ( .INP(n9470), .ZN(n9442) );
  NAND3X0 U9172 ( .IN1(n9471), .IN2(n9472), .IN3(n9473), .QN(n9470) );
  NAND2X0 U9173 ( .IN1(n9459), .IN2(n9474), .QN(n9473) );
  NAND2X0 U9174 ( .IN1(n9475), .IN2(n9456), .QN(n9471) );
  XOR2X1 U9175 ( .IN1(n8667), .IN2(n2669), .Q(n9475) );
  NAND2X0 U9176 ( .IN1(n9476), .IN2(n9477), .QN(g30684) );
  NAND2X0 U9177 ( .IN1(n4515), .IN2(g1651), .QN(n9477) );
  NAND2X0 U9178 ( .IN1(n9462), .IN2(g6782), .QN(n9476) );
  NAND2X0 U9179 ( .IN1(n9478), .IN2(n9479), .QN(g30683) );
  NAND2X0 U9180 ( .IN1(n4317), .IN2(g1576), .QN(n9479) );
  NAND2X0 U9181 ( .IN1(n9447), .IN2(g6573), .QN(n9478) );
  NAND3X0 U9182 ( .IN1(n9480), .IN2(n9481), .IN3(n9482), .QN(n9447) );
  NAND2X0 U9183 ( .IN1(n9483), .IN2(n9484), .QN(n9481) );
  XNOR2X1 U9184 ( .IN1(n9485), .IN2(n8650), .Q(n9483) );
  NAND2X0 U9185 ( .IN1(n9486), .IN2(g1481), .QN(n9480) );
  NAND2X0 U9186 ( .IN1(n9487), .IN2(n9488), .QN(g30682) );
  NAND2X0 U9187 ( .IN1(g960), .IN2(n8096), .QN(n9488) );
  NAND2X0 U9188 ( .IN1(n9489), .IN2(test_so31), .QN(n9487) );
  NAND2X0 U9189 ( .IN1(n9490), .IN2(n9491), .QN(g30681) );
  NAND2X0 U9190 ( .IN1(n4312), .IN2(g885), .QN(n9491) );
  NAND2X0 U9191 ( .IN1(n9467), .IN2(g6518), .QN(n9490) );
  NAND2X0 U9192 ( .IN1(n9492), .IN2(n9493), .QN(g30680) );
  NAND2X0 U9193 ( .IN1(n4369), .IN2(g201), .QN(n9493) );
  NAND2X0 U9194 ( .IN1(n9494), .IN2(g165), .QN(n9492) );
  NAND2X0 U9195 ( .IN1(n9495), .IN2(n9496), .QN(g30679) );
  NAND2X0 U9196 ( .IN1(n4367), .IN2(g2321), .QN(n9496) );
  NAND2X0 U9197 ( .IN1(n9497), .IN2(g2241), .QN(n9495) );
  NAND2X0 U9198 ( .IN1(n9498), .IN2(n9499), .QN(g30678) );
  NAND2X0 U9199 ( .IN1(n4317), .IN2(g1648), .QN(n9499) );
  NAND2X0 U9200 ( .IN1(n9462), .IN2(g6573), .QN(n9498) );
  INVX0 U9201 ( .INP(n9500), .ZN(n9462) );
  NAND3X0 U9202 ( .IN1(n9501), .IN2(n9502), .IN3(n9503), .QN(n9500) );
  NAND2X0 U9203 ( .IN1(n9486), .IN2(n9504), .QN(n9503) );
  NAND2X0 U9204 ( .IN1(n9505), .IN2(n9484), .QN(n9501) );
  XOR2X1 U9205 ( .IN1(n8643), .IN2(n2684), .Q(n9505) );
  NAND2X0 U9206 ( .IN1(n9506), .IN2(n9507), .QN(g30677) );
  NAND2X0 U9207 ( .IN1(n4312), .IN2(g957), .QN(n9507) );
  NAND2X0 U9208 ( .IN1(n9489), .IN2(g6518), .QN(n9506) );
  NAND2X0 U9209 ( .IN1(n9508), .IN2(n9509), .QN(g30676) );
  NAND2X0 U9210 ( .IN1(n4323), .IN2(g882), .QN(n9509) );
  NAND2X0 U9211 ( .IN1(n9467), .IN2(g6368), .QN(n9508) );
  NAND3X0 U9212 ( .IN1(n9510), .IN2(n9511), .IN3(n9512), .QN(n9467) );
  NAND2X0 U9213 ( .IN1(n9513), .IN2(g793), .QN(n9512) );
  NAND2X0 U9214 ( .IN1(n9514), .IN2(n9515), .QN(n9510) );
  XOR2X1 U9215 ( .IN1(n9516), .IN2(n9517), .Q(n9514) );
  NAND2X0 U9216 ( .IN1(n9518), .IN2(n9519), .QN(g30675) );
  NAND2X0 U9217 ( .IN1(n4369), .IN2(g273), .QN(n9519) );
  NAND2X0 U9218 ( .IN1(n9520), .IN2(g165), .QN(n9518) );
  NAND2X0 U9219 ( .IN1(n9521), .IN2(n9522), .QN(g30674) );
  NAND2X0 U9220 ( .IN1(n4512), .IN2(g198), .QN(n9522) );
  NAND2X0 U9221 ( .IN1(n9494), .IN2(g6313), .QN(n9521) );
  NAND2X0 U9222 ( .IN1(n9523), .IN2(n9524), .QN(g30673) );
  NAND2X0 U9223 ( .IN1(g2318), .IN2(n8097), .QN(n9524) );
  NAND2X0 U9224 ( .IN1(n9497), .IN2(test_so73), .QN(n9523) );
  NAND2X0 U9225 ( .IN1(n9525), .IN2(n9526), .QN(g30672) );
  NAND2X0 U9226 ( .IN1(n4367), .IN2(g2312), .QN(n9526) );
  NAND2X0 U9227 ( .IN1(n9527), .IN2(g2241), .QN(n9525) );
  NAND2X0 U9228 ( .IN1(n9528), .IN2(n9529), .QN(g30671) );
  NAND2X0 U9229 ( .IN1(n4368), .IN2(g1627), .QN(n9529) );
  NAND2X0 U9230 ( .IN1(n9530), .IN2(g1547), .QN(n9528) );
  NAND2X0 U9231 ( .IN1(n9531), .IN2(n9532), .QN(g30670) );
  NAND2X0 U9232 ( .IN1(n4323), .IN2(g954), .QN(n9532) );
  NAND2X0 U9233 ( .IN1(n9489), .IN2(g6368), .QN(n9531) );
  INVX0 U9234 ( .INP(n9533), .ZN(n9489) );
  NAND3X0 U9235 ( .IN1(n9534), .IN2(n9535), .IN3(n9536), .QN(n9533) );
  NAND2X0 U9236 ( .IN1(n9537), .IN2(n9513), .QN(n9536) );
  NAND2X0 U9237 ( .IN1(n9515), .IN2(n9538), .QN(n9534) );
  XOR2X1 U9238 ( .IN1(n9539), .IN2(n9540), .Q(n9538) );
  NOR2X0 U9239 ( .IN1(n9541), .IN2(n9542), .QN(n9540) );
  XOR2X1 U9240 ( .IN1(n9543), .IN2(n8607), .Q(n9541) );
  NAND2X0 U9241 ( .IN1(n9544), .IN2(n9545), .QN(g30669) );
  NAND2X0 U9242 ( .IN1(n4512), .IN2(g270), .QN(n9545) );
  NAND2X0 U9243 ( .IN1(n9520), .IN2(g6313), .QN(n9544) );
  NAND2X0 U9244 ( .IN1(n9546), .IN2(n9547), .QN(g30668) );
  NAND2X0 U9245 ( .IN1(n4318), .IN2(g195), .QN(n9547) );
  NAND2X0 U9246 ( .IN1(n9494), .IN2(g6231), .QN(n9546) );
  NAND3X0 U9247 ( .IN1(n9548), .IN2(n9549), .IN3(n9550), .QN(n9494) );
  NAND2X0 U9248 ( .IN1(n9551), .IN2(g105), .QN(n9550) );
  NAND2X0 U9249 ( .IN1(n9552), .IN2(n9553), .QN(n9548) );
  XNOR2X1 U9250 ( .IN1(n9554), .IN2(n8589), .Q(n9552) );
  NAND2X0 U9251 ( .IN1(n9555), .IN2(n9556), .QN(g30667) );
  NAND2X0 U9252 ( .IN1(n4324), .IN2(g2315), .QN(n9556) );
  NAND2X0 U9253 ( .IN1(n9497), .IN2(g6837), .QN(n9555) );
  INVX0 U9254 ( .INP(n9557), .ZN(n9497) );
  NAND3X0 U9255 ( .IN1(n9558), .IN2(n9472), .IN3(n9559), .QN(n9557) );
  NAND2X0 U9256 ( .IN1(n9459), .IN2(n4389), .QN(n9559) );
  NAND2X0 U9257 ( .IN1(n9456), .IN2(n9560), .QN(n9558) );
  XOR2X1 U9258 ( .IN1(n9561), .IN2(n9562), .Q(n9560) );
  NAND2X0 U9259 ( .IN1(n9563), .IN2(n9564), .QN(g30666) );
  NAND2X0 U9260 ( .IN1(g2309), .IN2(n8097), .QN(n9564) );
  NAND2X0 U9261 ( .IN1(n9527), .IN2(test_so73), .QN(n9563) );
  NAND2X0 U9262 ( .IN1(n9565), .IN2(n9566), .QN(g30665) );
  NAND2X0 U9263 ( .IN1(n4367), .IN2(g2303), .QN(n9566) );
  NAND2X0 U9264 ( .IN1(n9567), .IN2(g2241), .QN(n9565) );
  NAND2X0 U9265 ( .IN1(n9568), .IN2(n9569), .QN(g30664) );
  NAND2X0 U9266 ( .IN1(n4515), .IN2(g1624), .QN(n9569) );
  NAND2X0 U9267 ( .IN1(n9530), .IN2(g6782), .QN(n9568) );
  NAND2X0 U9268 ( .IN1(n9570), .IN2(n9571), .QN(g30663) );
  NAND2X0 U9269 ( .IN1(n4368), .IN2(g1618), .QN(n9571) );
  NAND2X0 U9270 ( .IN1(n9572), .IN2(g1547), .QN(n9570) );
  NAND2X0 U9271 ( .IN1(n9573), .IN2(n9574), .QN(g30662) );
  NAND2X0 U9272 ( .IN1(g933), .IN2(n8096), .QN(n9574) );
  NAND2X0 U9273 ( .IN1(n9575), .IN2(test_so31), .QN(n9573) );
  NAND2X0 U9274 ( .IN1(n9576), .IN2(n9577), .QN(g30661) );
  NAND2X0 U9275 ( .IN1(n4318), .IN2(g267), .QN(n9577) );
  NAND2X0 U9276 ( .IN1(n9520), .IN2(g6231), .QN(n9576) );
  INVX0 U9277 ( .INP(n9578), .ZN(n9520) );
  NAND3X0 U9278 ( .IN1(n9579), .IN2(n9580), .IN3(n9581), .QN(n9578) );
  NAND2X0 U9279 ( .IN1(n9582), .IN2(n9551), .QN(n9581) );
  NAND2X0 U9280 ( .IN1(n9583), .IN2(n9553), .QN(n9579) );
  XOR2X1 U9281 ( .IN1(n8576), .IN2(n2717), .Q(n9583) );
  NAND2X0 U9282 ( .IN1(n9584), .IN2(n9585), .QN(g30660) );
  NAND2X0 U9283 ( .IN1(n4324), .IN2(g2306), .QN(n9585) );
  NAND2X0 U9284 ( .IN1(n9527), .IN2(g6837), .QN(n9584) );
  INVX0 U9285 ( .INP(n9586), .ZN(n9527) );
  NAND3X0 U9286 ( .IN1(n9587), .IN2(n9472), .IN3(n9588), .QN(n9586) );
  NAND2X0 U9287 ( .IN1(n9459), .IN2(n4373), .QN(n9588) );
  NAND2X0 U9288 ( .IN1(n9589), .IN2(n4529), .QN(n9472) );
  NAND2X0 U9289 ( .IN1(n9456), .IN2(n9590), .QN(n9587) );
  XOR2X1 U9290 ( .IN1(n8682), .IN2(n9591), .Q(n9590) );
  INVX0 U9291 ( .INP(n9592), .ZN(n8682) );
  NAND2X0 U9292 ( .IN1(n9593), .IN2(n9594), .QN(g30659) );
  NAND2X0 U9293 ( .IN1(g2300), .IN2(n8097), .QN(n9594) );
  NAND2X0 U9294 ( .IN1(test_so73), .IN2(n9567), .QN(n9593) );
  NAND2X0 U9295 ( .IN1(n9595), .IN2(n9596), .QN(g30658) );
  NAND2X0 U9296 ( .IN1(n9530), .IN2(g6573), .QN(n9596) );
  INVX0 U9297 ( .INP(n9597), .ZN(n9530) );
  NAND3X0 U9298 ( .IN1(n9598), .IN2(n9502), .IN3(n9599), .QN(n9597) );
  NAND2X0 U9299 ( .IN1(n9486), .IN2(n4390), .QN(n9599) );
  NAND2X0 U9300 ( .IN1(n9484), .IN2(n9600), .QN(n9598) );
  XOR2X1 U9301 ( .IN1(n9601), .IN2(n8641), .Q(n9600) );
  NAND2X0 U9302 ( .IN1(test_so55), .IN2(n4317), .QN(n9595) );
  NAND2X0 U9303 ( .IN1(n9602), .IN2(n9603), .QN(g30657) );
  NAND2X0 U9304 ( .IN1(n4515), .IN2(g1615), .QN(n9603) );
  NAND2X0 U9305 ( .IN1(n9572), .IN2(g6782), .QN(n9602) );
  NAND2X0 U9306 ( .IN1(n9604), .IN2(n9605), .QN(g30656) );
  NAND2X0 U9307 ( .IN1(n4368), .IN2(g1609), .QN(n9605) );
  NAND2X0 U9308 ( .IN1(n9606), .IN2(g1547), .QN(n9604) );
  NAND2X0 U9309 ( .IN1(n9607), .IN2(n9608), .QN(g30655) );
  NAND2X0 U9310 ( .IN1(n4312), .IN2(g930), .QN(n9608) );
  NAND2X0 U9311 ( .IN1(n9575), .IN2(g6518), .QN(n9607) );
  NAND2X0 U9312 ( .IN1(n9609), .IN2(n9610), .QN(g30654) );
  NAND2X0 U9313 ( .IN1(test_so34), .IN2(n8096), .QN(n9610) );
  NAND2X0 U9314 ( .IN1(n9611), .IN2(test_so31), .QN(n9609) );
  NAND2X0 U9315 ( .IN1(n9612), .IN2(n9613), .QN(g30653) );
  NAND2X0 U9316 ( .IN1(n4369), .IN2(g246), .QN(n9613) );
  NAND2X0 U9317 ( .IN1(n9614), .IN2(g165), .QN(n9612) );
  NAND2X0 U9318 ( .IN1(n9615), .IN2(n9616), .QN(g30652) );
  NAND2X0 U9319 ( .IN1(n4324), .IN2(g2297), .QN(n9616) );
  NAND2X0 U9320 ( .IN1(n9567), .IN2(g6837), .QN(n9615) );
  NAND3X0 U9321 ( .IN1(n9617), .IN2(n9618), .IN3(n9454), .QN(n9567) );
  NAND2X0 U9322 ( .IN1(n9589), .IN2(n9619), .QN(n9454) );
  NAND2X0 U9323 ( .IN1(n9620), .IN2(n9456), .QN(n9618) );
  XNOR2X1 U9324 ( .IN1(n2670), .IN2(n8678), .Q(n9620) );
  NAND2X0 U9325 ( .IN1(n9621), .IN2(n9622), .QN(n2670) );
  XOR2X1 U9326 ( .IN1(n8672), .IN2(n9202), .Q(n9622) );
  NAND2X0 U9327 ( .IN1(n9459), .IN2(n9623), .QN(n9617) );
  NAND2X0 U9328 ( .IN1(n9624), .IN2(n9625), .QN(g30651) );
  NAND2X0 U9329 ( .IN1(n4317), .IN2(g1612), .QN(n9625) );
  NAND2X0 U9330 ( .IN1(n9572), .IN2(g6573), .QN(n9624) );
  INVX0 U9331 ( .INP(n9626), .ZN(n9572) );
  NAND3X0 U9332 ( .IN1(n9627), .IN2(n9502), .IN3(n9628), .QN(n9626) );
  NAND2X0 U9333 ( .IN1(n9486), .IN2(n4374), .QN(n9628) );
  NAND2X0 U9334 ( .IN1(n9629), .IN2(n4530), .QN(n9502) );
  NAND2X0 U9335 ( .IN1(n9484), .IN2(n9630), .QN(n9627) );
  XOR2X1 U9336 ( .IN1(n8640), .IN2(n9631), .Q(n9630) );
  NAND2X0 U9337 ( .IN1(n9632), .IN2(n9633), .QN(g30650) );
  NAND2X0 U9338 ( .IN1(test_so56), .IN2(n4515), .QN(n9633) );
  NAND2X0 U9339 ( .IN1(n9606), .IN2(g6782), .QN(n9632) );
  NAND2X0 U9340 ( .IN1(n9634), .IN2(n9635), .QN(g30649) );
  NAND2X0 U9341 ( .IN1(n4323), .IN2(g927), .QN(n9635) );
  NAND2X0 U9342 ( .IN1(n9575), .IN2(g6368), .QN(n9634) );
  INVX0 U9343 ( .INP(n9636), .ZN(n9575) );
  NAND3X0 U9344 ( .IN1(n9637), .IN2(n9535), .IN3(n9638), .QN(n9636) );
  NAND2X0 U9345 ( .IN1(n4391), .IN2(n9513), .QN(n9638) );
  NAND2X0 U9346 ( .IN1(n9515), .IN2(n9639), .QN(n9637) );
  XNOR2X1 U9347 ( .IN1(n8620), .IN2(n9640), .Q(n9639) );
  NAND2X0 U9348 ( .IN1(n9641), .IN2(n9642), .QN(g30648) );
  NAND2X0 U9349 ( .IN1(n4312), .IN2(g921), .QN(n9642) );
  NAND2X0 U9350 ( .IN1(n9611), .IN2(g6518), .QN(n9641) );
  NAND2X0 U9351 ( .IN1(n9643), .IN2(n9644), .QN(g30647) );
  NAND2X0 U9352 ( .IN1(g915), .IN2(n8096), .QN(n9644) );
  NAND2X0 U9353 ( .IN1(test_so31), .IN2(n9645), .QN(n9643) );
  NAND2X0 U9354 ( .IN1(n9646), .IN2(n9647), .QN(g30646) );
  NAND2X0 U9355 ( .IN1(n4512), .IN2(g243), .QN(n9647) );
  NAND2X0 U9356 ( .IN1(n9614), .IN2(g6313), .QN(n9646) );
  NAND2X0 U9357 ( .IN1(n9648), .IN2(n9649), .QN(g30645) );
  NAND2X0 U9358 ( .IN1(n4369), .IN2(g237), .QN(n9649) );
  NAND2X0 U9359 ( .IN1(n9650), .IN2(g165), .QN(n9648) );
  NAND2X0 U9360 ( .IN1(n9651), .IN2(n9652), .QN(g30644) );
  NAND2X0 U9361 ( .IN1(n4317), .IN2(g1603), .QN(n9652) );
  NAND2X0 U9362 ( .IN1(n9606), .IN2(g6573), .QN(n9651) );
  NAND3X0 U9363 ( .IN1(n9653), .IN2(n9654), .IN3(n9482), .QN(n9606) );
  NAND2X0 U9364 ( .IN1(n9629), .IN2(n9655), .QN(n9482) );
  NAND2X0 U9365 ( .IN1(n9656), .IN2(n9484), .QN(n9654) );
  XOR2X1 U9366 ( .IN1(n2685), .IN2(n8652), .Q(n9656) );
  NAND2X0 U9367 ( .IN1(n9657), .IN2(n9658), .QN(n2685) );
  XOR2X1 U9368 ( .IN1(n9659), .IN2(n9201), .Q(n9658) );
  NAND2X0 U9369 ( .IN1(n9486), .IN2(n9660), .QN(n9653) );
  NAND2X0 U9370 ( .IN1(n9661), .IN2(n9662), .QN(g30643) );
  NAND2X0 U9371 ( .IN1(n4323), .IN2(g918), .QN(n9662) );
  NAND2X0 U9372 ( .IN1(n9611), .IN2(g6368), .QN(n9661) );
  INVX0 U9373 ( .INP(n9663), .ZN(n9611) );
  NAND3X0 U9374 ( .IN1(n9664), .IN2(n9535), .IN3(n9665), .QN(n9663) );
  NAND2X0 U9375 ( .IN1(n4375), .IN2(n9513), .QN(n9665) );
  NAND3X0 U9376 ( .IN1(n9666), .IN2(n9543), .IN3(n9667), .QN(n9535) );
  NAND2X0 U9377 ( .IN1(n9515), .IN2(n9668), .QN(n9664) );
  XNOR2X1 U9378 ( .IN1(n8619), .IN2(n9669), .Q(n9668) );
  NAND2X0 U9379 ( .IN1(n9670), .IN2(n9671), .QN(g30642) );
  NAND2X0 U9380 ( .IN1(n4312), .IN2(g912), .QN(n9671) );
  NAND2X0 U9381 ( .IN1(n9645), .IN2(g6518), .QN(n9670) );
  NAND2X0 U9382 ( .IN1(n9672), .IN2(n9673), .QN(g30641) );
  NAND2X0 U9383 ( .IN1(n4318), .IN2(g240), .QN(n9673) );
  NAND2X0 U9384 ( .IN1(n9614), .IN2(g6231), .QN(n9672) );
  INVX0 U9385 ( .INP(n9674), .ZN(n9614) );
  NAND3X0 U9386 ( .IN1(n9675), .IN2(n9580), .IN3(n9676), .QN(n9674) );
  NAND2X0 U9387 ( .IN1(n4392), .IN2(n9551), .QN(n9676) );
  NAND2X0 U9388 ( .IN1(n9553), .IN2(n9677), .QN(n9675) );
  XOR2X1 U9389 ( .IN1(n8594), .IN2(n9678), .Q(n9677) );
  NAND2X0 U9390 ( .IN1(n9679), .IN2(n9680), .QN(g30640) );
  NAND2X0 U9391 ( .IN1(n4512), .IN2(g234), .QN(n9680) );
  NAND2X0 U9392 ( .IN1(n9650), .IN2(g6313), .QN(n9679) );
  NAND2X0 U9393 ( .IN1(n9681), .IN2(n9682), .QN(g30639) );
  NAND2X0 U9394 ( .IN1(n4369), .IN2(g228), .QN(n9682) );
  NAND2X0 U9395 ( .IN1(n9683), .IN2(g165), .QN(n9681) );
  NAND2X0 U9396 ( .IN1(n9684), .IN2(n9685), .QN(g30638) );
  NAND2X0 U9397 ( .IN1(n4323), .IN2(g909), .QN(n9685) );
  NAND2X0 U9398 ( .IN1(n9645), .IN2(g6368), .QN(n9684) );
  NAND3X0 U9399 ( .IN1(n9686), .IN2(n9511), .IN3(n9687), .QN(n9645) );
  NAND2X0 U9400 ( .IN1(n9513), .IN2(n9688), .QN(n9687) );
  NAND3X0 U9401 ( .IN1(n9666), .IN2(n9689), .IN3(n9667), .QN(n9511) );
  NAND2X0 U9402 ( .IN1(n9690), .IN2(n9515), .QN(n9686) );
  XNOR2X1 U9403 ( .IN1(n9542), .IN2(n8607), .Q(n9690) );
  NAND2X0 U9404 ( .IN1(n9691), .IN2(n9692), .QN(n9542) );
  XOR2X1 U9405 ( .IN1(n8623), .IN2(n9689), .Q(n9692) );
  NAND2X0 U9406 ( .IN1(n9693), .IN2(n9694), .QN(g30637) );
  NAND2X0 U9407 ( .IN1(n4318), .IN2(g231), .QN(n9694) );
  NAND2X0 U9408 ( .IN1(n9650), .IN2(g6231), .QN(n9693) );
  INVX0 U9409 ( .INP(n9695), .ZN(n9650) );
  NAND3X0 U9410 ( .IN1(n9696), .IN2(n9580), .IN3(n9697), .QN(n9695) );
  NAND2X0 U9411 ( .IN1(n4376), .IN2(n9551), .QN(n9697) );
  NAND3X0 U9412 ( .IN1(n9698), .IN2(n9699), .IN3(n9700), .QN(n9580) );
  NAND2X0 U9413 ( .IN1(n9553), .IN2(n9701), .QN(n9696) );
  XOR2X1 U9414 ( .IN1(n8583), .IN2(n9702), .Q(n9701) );
  NAND2X0 U9415 ( .IN1(n9703), .IN2(n9704), .QN(g30636) );
  NAND2X0 U9416 ( .IN1(n4512), .IN2(g225), .QN(n9704) );
  NAND2X0 U9417 ( .IN1(n9683), .IN2(g6313), .QN(n9703) );
  NAND2X0 U9418 ( .IN1(n9705), .IN2(n9706), .QN(g30635) );
  NAND2X0 U9419 ( .IN1(n4318), .IN2(g222), .QN(n9706) );
  NAND2X0 U9420 ( .IN1(n9683), .IN2(g6231), .QN(n9705) );
  NAND3X0 U9421 ( .IN1(n9707), .IN2(n9549), .IN3(n9708), .QN(n9683) );
  NAND2X0 U9422 ( .IN1(n9551), .IN2(n9709), .QN(n9708) );
  NAND3X0 U9423 ( .IN1(n9698), .IN2(n9199), .IN3(n9700), .QN(n9549) );
  NAND2X0 U9424 ( .IN1(n9710), .IN2(n9553), .QN(n9707) );
  XOR2X1 U9425 ( .IN1(n2718), .IN2(n9711), .Q(n9710) );
  NAND2X0 U9426 ( .IN1(n9712), .IN2(n9713), .QN(n2718) );
  XOR2X1 U9427 ( .IN1(n8578), .IN2(n9199), .Q(n9713) );
  NAND2X0 U9428 ( .IN1(n9714), .IN2(n9715), .QN(g30566) );
  NAND2X0 U9429 ( .IN1(n9350), .IN2(n4606), .QN(n9715) );
  INVX0 U9430 ( .INP(n9716), .ZN(n9350) );
  NAND2X0 U9431 ( .IN1(n9717), .IN2(n9718), .QN(n9716) );
  XOR2X1 U9432 ( .IN1(n9719), .IN2(n9720), .Q(n9717) );
  NAND2X0 U9433 ( .IN1(n9721), .IN2(n9722), .QN(n9720) );
  NAND2X0 U9434 ( .IN1(n9723), .IN2(n9724), .QN(n9722) );
  NAND4X0 U9435 ( .IN1(n9725), .IN2(n9726), .IN3(n9727), .IN4(n9728), .QN(
        n9721) );
  NAND3X0 U9436 ( .IN1(n9729), .IN2(n9730), .IN3(n9731), .QN(n9727) );
  NAND2X0 U9437 ( .IN1(n9732), .IN2(n9719), .QN(n9726) );
  INVX0 U9438 ( .INP(n9733), .ZN(n9732) );
  NAND2X0 U9439 ( .IN1(n9734), .IN2(n9735), .QN(n9725) );
  NAND2X0 U9440 ( .IN1(n9736), .IN2(n9737), .QN(n9734) );
  NAND2X0 U9441 ( .IN1(n9729), .IN2(n9738), .QN(n9737) );
  NAND3X0 U9442 ( .IN1(n9739), .IN2(n9730), .IN3(n9740), .QN(n9738) );
  INVX0 U9443 ( .INP(n9741), .ZN(n9740) );
  NAND2X0 U9444 ( .IN1(n9733), .IN2(n9742), .QN(n9739) );
  NAND2X0 U9445 ( .IN1(n9743), .IN2(n9744), .QN(n9736) );
  NAND2X0 U9446 ( .IN1(n2792), .IN2(n9745), .QN(n9743) );
  NAND2X0 U9447 ( .IN1(n4509), .IN2(g2392), .QN(n9714) );
  NAND2X0 U9448 ( .IN1(n9746), .IN2(n9747), .QN(g30505) );
  NAND2X0 U9449 ( .IN1(n9748), .IN2(g5555), .QN(n9747) );
  NAND2X0 U9450 ( .IN1(n4516), .IN2(g2393), .QN(n9746) );
  NAND2X0 U9451 ( .IN1(n9749), .IN2(n9750), .QN(g30503) );
  NAND2X0 U9452 ( .IN1(n9751), .IN2(g7014), .QN(n9750) );
  NAND2X0 U9453 ( .IN1(n4525), .IN2(g1700), .QN(n9749) );
  NAND2X0 U9454 ( .IN1(n9752), .IN2(n9753), .QN(g30500) );
  NAND2X0 U9455 ( .IN1(n2798), .IN2(g1088), .QN(n9753) );
  NAND2X0 U9456 ( .IN1(test_so39), .IN2(n4381), .QN(n9752) );
  NAND2X0 U9457 ( .IN1(n9754), .IN2(n9755), .QN(g30487) );
  NAND2X0 U9458 ( .IN1(n9751), .IN2(g5511), .QN(n9755) );
  NAND2X0 U9459 ( .IN1(n4518), .IN2(g1699), .QN(n9754) );
  NAND2X0 U9460 ( .IN1(n9756), .IN2(n9757), .QN(g30485) );
  NAND2X0 U9461 ( .IN1(n4364), .IN2(g1006), .QN(n9757) );
  NAND2X0 U9462 ( .IN1(n2798), .IN2(g6712), .QN(n9756) );
  NAND2X0 U9463 ( .IN1(n9758), .IN2(n9759), .QN(g30482) );
  NAND2X0 U9464 ( .IN1(n9760), .IN2(n4640), .QN(n9759) );
  NAND2X0 U9465 ( .IN1(n4506), .IN2(g320), .QN(n9758) );
  NAND2X0 U9466 ( .IN1(n9761), .IN2(n9762), .QN(g30470) );
  NAND2X0 U9467 ( .IN1(n4363), .IN2(g1005), .QN(n9762) );
  NAND2X0 U9468 ( .IN1(n2798), .IN2(g5472), .QN(n9761) );
  NAND2X0 U9469 ( .IN1(n9763), .IN2(n9764), .QN(g30468) );
  NAND2X0 U9470 ( .IN1(n9760), .IN2(g6447), .QN(n9764) );
  NAND2X0 U9471 ( .IN1(n4499), .IN2(g319), .QN(n9763) );
  NAND2X0 U9472 ( .IN1(n9765), .IN2(n9766), .QN(g30455) );
  NAND2X0 U9473 ( .IN1(n9760), .IN2(g5437), .QN(n9766) );
  INVX0 U9474 ( .INP(n9767), .ZN(n9760) );
  NAND2X0 U9475 ( .IN1(n9768), .IN2(n9407), .QN(n9767) );
  XOR2X1 U9476 ( .IN1(n9769), .IN2(n9418), .Q(n9768) );
  NAND2X0 U9477 ( .IN1(n9770), .IN2(n9771), .QN(n9769) );
  NAND2X0 U9478 ( .IN1(n9418), .IN2(n9772), .QN(n9771) );
  NAND3X0 U9479 ( .IN1(n9773), .IN2(n9774), .IN3(n9417), .QN(n9772) );
  NAND2X0 U9480 ( .IN1(n9430), .IN2(n9408), .QN(n9774) );
  NAND2X0 U9481 ( .IN1(n9436), .IN2(n9775), .QN(n9430) );
  NAND2X0 U9482 ( .IN1(n9776), .IN2(n3130), .QN(n9775) );
  INVX0 U9483 ( .INP(n9777), .ZN(n9776) );
  NAND3X0 U9484 ( .IN1(n9778), .IN2(g309), .IN3(n9424), .QN(n9773) );
  INVX0 U9485 ( .INP(n9779), .ZN(n9778) );
  NAND3X0 U9486 ( .IN1(n9420), .IN2(n9417), .IN3(n9434), .QN(n9770) );
  INVX0 U9487 ( .INP(n9780), .ZN(n9420) );
  NAND3X0 U9488 ( .IN1(n9777), .IN2(n9408), .IN3(n3130), .QN(n9780) );
  NAND2X0 U9489 ( .IN1(n4520), .IN2(g318), .QN(n9765) );
  NAND2X0 U9490 ( .IN1(n9781), .IN2(n9782), .QN(g30356) );
  NAND2X0 U9491 ( .IN1(n9748), .IN2(n4606), .QN(n9782) );
  NAND2X0 U9492 ( .IN1(n4509), .IN2(g2395), .QN(n9781) );
  NAND2X0 U9493 ( .IN1(n9783), .IN2(n9784), .QN(g30341) );
  NAND2X0 U9494 ( .IN1(n9748), .IN2(g7264), .QN(n9784) );
  INVX0 U9495 ( .INP(n9785), .ZN(n9748) );
  NAND2X0 U9496 ( .IN1(n9786), .IN2(n9718), .QN(n9785) );
  XOR2X1 U9497 ( .IN1(n9787), .IN2(n9729), .Q(n9786) );
  NAND2X0 U9498 ( .IN1(n9788), .IN2(n9789), .QN(n9787) );
  NAND2X0 U9499 ( .IN1(n9729), .IN2(n9790), .QN(n9789) );
  NAND3X0 U9500 ( .IN1(n9791), .IN2(n9792), .IN3(n9728), .QN(n9790) );
  NAND2X0 U9501 ( .IN1(n9741), .IN2(n9719), .QN(n9792) );
  NAND2X0 U9502 ( .IN1(n9745), .IN2(n9793), .QN(n9741) );
  NAND2X0 U9503 ( .IN1(n9794), .IN2(n3038), .QN(n9793) );
  INVX0 U9504 ( .INP(n9795), .ZN(n9794) );
  NAND3X0 U9505 ( .IN1(n9796), .IN2(test_so79), .IN3(n9735), .QN(n9791) );
  NAND3X0 U9506 ( .IN1(n9731), .IN2(n9728), .IN3(n9744), .QN(n9788) );
  INVX0 U9507 ( .INP(n9797), .ZN(n9731) );
  NAND3X0 U9508 ( .IN1(n9795), .IN2(n9719), .IN3(n3038), .QN(n9797) );
  NAND2X0 U9509 ( .IN1(n4524), .IN2(g2394), .QN(n9783) );
  NAND2X0 U9510 ( .IN1(n9798), .IN2(n9799), .QN(g30338) );
  NAND2X0 U9511 ( .IN1(n9751), .IN2(n4618), .QN(n9799) );
  INVX0 U9512 ( .INP(n9800), .ZN(n9751) );
  NAND2X0 U9513 ( .IN1(n9801), .IN2(n9364), .QN(n9800) );
  XOR2X1 U9514 ( .IN1(n9802), .IN2(n9375), .Q(n9801) );
  NAND2X0 U9515 ( .IN1(n9803), .IN2(n9804), .QN(n9802) );
  NAND2X0 U9516 ( .IN1(n9375), .IN2(n9805), .QN(n9804) );
  NAND3X0 U9517 ( .IN1(n9806), .IN2(n9807), .IN3(n9374), .QN(n9805) );
  NAND2X0 U9518 ( .IN1(n9387), .IN2(n9365), .QN(n9807) );
  NAND2X0 U9519 ( .IN1(n9393), .IN2(n9808), .QN(n9387) );
  NAND2X0 U9520 ( .IN1(n9809), .IN2(n3070), .QN(n9808) );
  INVX0 U9521 ( .INP(n9810), .ZN(n9809) );
  NAND3X0 U9522 ( .IN1(n9811), .IN2(g1690), .IN3(n9381), .QN(n9806) );
  INVX0 U9523 ( .INP(n9812), .ZN(n9811) );
  NAND3X0 U9524 ( .IN1(n9377), .IN2(n9374), .IN3(n9391), .QN(n9803) );
  INVX0 U9525 ( .INP(n9813), .ZN(n9377) );
  NAND3X0 U9526 ( .IN1(n9810), .IN2(n9365), .IN3(n3070), .QN(n9813) );
  NAND2X0 U9527 ( .IN1(n4511), .IN2(g1701), .QN(n9798) );
  NAND2X0 U9528 ( .IN1(n9814), .IN2(n9815), .QN(g30304) );
  NAND2X0 U9529 ( .IN1(n4367), .IN2(g2285), .QN(n9815) );
  NAND2X0 U9530 ( .IN1(n9816), .IN2(g2241), .QN(n9814) );
  NAND2X0 U9531 ( .IN1(n9817), .IN2(n9818), .QN(g30303) );
  NAND2X0 U9532 ( .IN1(g2282), .IN2(n8097), .QN(n9818) );
  NAND2X0 U9533 ( .IN1(test_so73), .IN2(n9816), .QN(n9817) );
  NAND2X0 U9534 ( .IN1(n9819), .IN2(n9820), .QN(g30302) );
  NAND2X0 U9535 ( .IN1(n4368), .IN2(g1591), .QN(n9820) );
  NAND2X0 U9536 ( .IN1(n9821), .IN2(g1547), .QN(n9819) );
  NAND2X0 U9537 ( .IN1(n9822), .IN2(n9823), .QN(g30301) );
  NAND2X0 U9538 ( .IN1(n4324), .IN2(g2279), .QN(n9823) );
  NAND2X0 U9539 ( .IN1(n9816), .IN2(g6837), .QN(n9822) );
  NAND2X0 U9540 ( .IN1(n9824), .IN2(n9825), .QN(n9816) );
  NAND2X0 U9541 ( .IN1(n9826), .IN2(n9456), .QN(n9825) );
  XOR2X1 U9542 ( .IN1(n9827), .IN2(n9828), .Q(n9826) );
  NAND2X0 U9543 ( .IN1(n9459), .IN2(g2185), .QN(n9824) );
  NAND2X0 U9544 ( .IN1(n9829), .IN2(n9830), .QN(g30300) );
  NAND2X0 U9545 ( .IN1(n4367), .IN2(g2267), .QN(n9830) );
  NAND2X0 U9546 ( .IN1(n9831), .IN2(g2241), .QN(n9829) );
  NAND2X0 U9547 ( .IN1(n9832), .IN2(n9833), .QN(g30299) );
  NAND2X0 U9548 ( .IN1(n4515), .IN2(g1588), .QN(n9833) );
  NAND2X0 U9549 ( .IN1(n9821), .IN2(g6782), .QN(n9832) );
  NAND2X0 U9550 ( .IN1(n9834), .IN2(n9835), .QN(g30298) );
  NAND2X0 U9551 ( .IN1(g897), .IN2(n8096), .QN(n9835) );
  NAND2X0 U9552 ( .IN1(test_so31), .IN2(n9836), .QN(n9834) );
  NAND2X0 U9553 ( .IN1(n9837), .IN2(n9838), .QN(g30297) );
  NAND2X0 U9554 ( .IN1(n4367), .IN2(g2339), .QN(n9838) );
  NAND2X0 U9555 ( .IN1(n9839), .IN2(g2241), .QN(n9837) );
  NAND2X0 U9556 ( .IN1(n9840), .IN2(n9841), .QN(g30296) );
  NAND2X0 U9557 ( .IN1(test_so76), .IN2(n8097), .QN(n9841) );
  NAND2X0 U9558 ( .IN1(test_so73), .IN2(n9831), .QN(n9840) );
  NAND2X0 U9559 ( .IN1(n9842), .IN2(n9843), .QN(g30295) );
  NAND2X0 U9560 ( .IN1(n4317), .IN2(g1585), .QN(n9843) );
  NAND2X0 U9561 ( .IN1(n9821), .IN2(g6573), .QN(n9842) );
  NAND2X0 U9562 ( .IN1(n9844), .IN2(n9845), .QN(n9821) );
  NAND2X0 U9563 ( .IN1(n9846), .IN2(n9484), .QN(n9845) );
  XNOR2X1 U9564 ( .IN1(n9847), .IN2(n8653), .Q(n9846) );
  NAND2X0 U9565 ( .IN1(n9486), .IN2(g1491), .QN(n9844) );
  NAND2X0 U9566 ( .IN1(n9848), .IN2(n9849), .QN(g30294) );
  NAND2X0 U9567 ( .IN1(n4368), .IN2(g1573), .QN(n9849) );
  NAND2X0 U9568 ( .IN1(n9850), .IN2(g1547), .QN(n9848) );
  NAND2X0 U9569 ( .IN1(n9851), .IN2(n9852), .QN(g30293) );
  NAND2X0 U9570 ( .IN1(n4312), .IN2(g894), .QN(n9852) );
  NAND2X0 U9571 ( .IN1(n9836), .IN2(g6518), .QN(n9851) );
  NAND2X0 U9572 ( .IN1(n9853), .IN2(n9854), .QN(g30292) );
  NAND2X0 U9573 ( .IN1(n4369), .IN2(g210), .QN(n9854) );
  NAND2X0 U9574 ( .IN1(n9855), .IN2(g165), .QN(n9853) );
  NAND2X0 U9575 ( .IN1(n9856), .IN2(n9857), .QN(g30291) );
  NAND2X0 U9576 ( .IN1(g2336), .IN2(n8097), .QN(n9857) );
  NAND2X0 U9577 ( .IN1(test_so73), .IN2(n9839), .QN(n9856) );
  NAND2X0 U9578 ( .IN1(n9858), .IN2(n9859), .QN(g30290) );
  NAND2X0 U9579 ( .IN1(n4367), .IN2(g2330), .QN(n9859) );
  NAND2X0 U9580 ( .IN1(n9860), .IN2(g2241), .QN(n9858) );
  NAND2X0 U9581 ( .IN1(n9861), .IN2(n9862), .QN(g30289) );
  NAND2X0 U9582 ( .IN1(n4324), .IN2(g2261), .QN(n9862) );
  NAND2X0 U9583 ( .IN1(n9831), .IN2(g6837), .QN(n9861) );
  NAND2X0 U9584 ( .IN1(n9863), .IN2(n9864), .QN(n9831) );
  NAND2X0 U9585 ( .IN1(n9456), .IN2(n9865), .QN(n9864) );
  XOR2X1 U9586 ( .IN1(n9866), .IN2(n9867), .Q(n9865) );
  NAND2X0 U9587 ( .IN1(n9459), .IN2(g2165), .QN(n9863) );
  NAND2X0 U9588 ( .IN1(n9868), .IN2(n9869), .QN(g30288) );
  NAND2X0 U9589 ( .IN1(n4368), .IN2(g1645), .QN(n9869) );
  NAND2X0 U9590 ( .IN1(n9870), .IN2(g1547), .QN(n9868) );
  NAND2X0 U9591 ( .IN1(n9871), .IN2(n9872), .QN(g30287) );
  NAND2X0 U9592 ( .IN1(n4515), .IN2(g1570), .QN(n9872) );
  NAND2X0 U9593 ( .IN1(n9850), .IN2(g6782), .QN(n9871) );
  NAND2X0 U9594 ( .IN1(n9873), .IN2(n9874), .QN(g30286) );
  NAND2X0 U9595 ( .IN1(n4323), .IN2(g891), .QN(n9874) );
  NAND2X0 U9596 ( .IN1(n9836), .IN2(g6368), .QN(n9873) );
  NAND2X0 U9597 ( .IN1(n9875), .IN2(n9876), .QN(n9836) );
  NAND2X0 U9598 ( .IN1(n9877), .IN2(n9515), .QN(n9876) );
  XOR2X1 U9599 ( .IN1(n9878), .IN2(n9879), .Q(n9877) );
  INVX0 U9600 ( .INP(n9880), .ZN(n9875) );
  NOR2X0 U9601 ( .IN1(n9667), .IN2(n4327), .QN(n9880) );
  NAND2X0 U9602 ( .IN1(n9881), .IN2(n9882), .QN(g30285) );
  NAND2X0 U9603 ( .IN1(g879), .IN2(n8096), .QN(n9882) );
  NAND2X0 U9604 ( .IN1(test_so31), .IN2(n9883), .QN(n9881) );
  NAND2X0 U9605 ( .IN1(n9884), .IN2(n9885), .QN(g30284) );
  NAND2X0 U9606 ( .IN1(n4512), .IN2(g207), .QN(n9885) );
  NAND2X0 U9607 ( .IN1(n9855), .IN2(g6313), .QN(n9884) );
  NAND2X0 U9608 ( .IN1(n9886), .IN2(n9887), .QN(g30283) );
  NAND2X0 U9609 ( .IN1(n4324), .IN2(g2333), .QN(n9887) );
  NAND2X0 U9610 ( .IN1(n9839), .IN2(g6837), .QN(n9886) );
  NAND2X0 U9611 ( .IN1(n9888), .IN2(n9889), .QN(n9839) );
  NAND3X0 U9612 ( .IN1(n9456), .IN2(n9890), .IN3(n9891), .QN(n9889) );
  XOR2X1 U9613 ( .IN1(n8672), .IN2(n9621), .Q(n9891) );
  NOR2X0 U9614 ( .IN1(n9892), .IN2(n9893), .QN(n9621) );
  XOR2X1 U9615 ( .IN1(n9894), .IN2(n9202), .Q(n9893) );
  NAND2X0 U9616 ( .IN1(n9459), .IN2(g2200), .QN(n9888) );
  NAND2X0 U9617 ( .IN1(n9895), .IN2(n9896), .QN(g30282) );
  NAND2X0 U9618 ( .IN1(test_so77), .IN2(n8097), .QN(n9896) );
  NAND2X0 U9619 ( .IN1(test_so73), .IN2(n9860), .QN(n9895) );
  NAND2X0 U9620 ( .IN1(n9897), .IN2(n9898), .QN(g30281) );
  NAND2X0 U9621 ( .IN1(n4515), .IN2(g1642), .QN(n9898) );
  NAND2X0 U9622 ( .IN1(n9870), .IN2(g6782), .QN(n9897) );
  NAND2X0 U9623 ( .IN1(n9899), .IN2(n9900), .QN(g30280) );
  NAND2X0 U9624 ( .IN1(n4368), .IN2(g1636), .QN(n9900) );
  NAND2X0 U9625 ( .IN1(n9901), .IN2(g1547), .QN(n9899) );
  NAND2X0 U9626 ( .IN1(n9902), .IN2(n9903), .QN(g30279) );
  NAND2X0 U9627 ( .IN1(n4317), .IN2(g1567), .QN(n9903) );
  NAND2X0 U9628 ( .IN1(n9850), .IN2(g6573), .QN(n9902) );
  NAND2X0 U9629 ( .IN1(n9904), .IN2(n9905), .QN(n9850) );
  NAND2X0 U9630 ( .IN1(n9484), .IN2(n9906), .QN(n9905) );
  XOR2X1 U9631 ( .IN1(n8651), .IN2(n9907), .Q(n9906) );
  NAND2X0 U9632 ( .IN1(n9486), .IN2(g1471), .QN(n9904) );
  NAND2X0 U9633 ( .IN1(n9908), .IN2(n9909), .QN(g30278) );
  NAND2X0 U9634 ( .IN1(g951), .IN2(n8096), .QN(n9909) );
  NAND2X0 U9635 ( .IN1(test_so31), .IN2(n9910), .QN(n9908) );
  NAND2X0 U9636 ( .IN1(n9911), .IN2(n9912), .QN(g30277) );
  NAND2X0 U9637 ( .IN1(n4312), .IN2(g876), .QN(n9912) );
  NAND2X0 U9638 ( .IN1(n9883), .IN2(g6518), .QN(n9911) );
  NAND2X0 U9639 ( .IN1(n9913), .IN2(n9914), .QN(g30276) );
  NAND2X0 U9640 ( .IN1(n4318), .IN2(g204), .QN(n9914) );
  NAND2X0 U9641 ( .IN1(n9855), .IN2(g6231), .QN(n9913) );
  NAND2X0 U9642 ( .IN1(n9915), .IN2(n9916), .QN(n9855) );
  NAND2X0 U9643 ( .IN1(n9917), .IN2(n9553), .QN(n9916) );
  XNOR2X1 U9644 ( .IN1(n9918), .IN2(n8588), .Q(n9917) );
  NAND2X0 U9645 ( .IN1(n9551), .IN2(g113), .QN(n9915) );
  NAND2X0 U9646 ( .IN1(n9919), .IN2(n9920), .QN(g30275) );
  NAND2X0 U9647 ( .IN1(n4369), .IN2(g192), .QN(n9920) );
  NAND2X0 U9648 ( .IN1(n9921), .IN2(g165), .QN(n9919) );
  NAND2X0 U9649 ( .IN1(n9922), .IN2(n9923), .QN(g30274) );
  NAND2X0 U9650 ( .IN1(n4324), .IN2(g2324), .QN(n9923) );
  NAND2X0 U9651 ( .IN1(n9860), .IN2(g6837), .QN(n9922) );
  NAND2X0 U9652 ( .IN1(n9924), .IN2(n9925), .QN(n9860) );
  NAND3X0 U9653 ( .IN1(n9456), .IN2(n9890), .IN3(n9926), .QN(n9925) );
  XOR2X1 U9654 ( .IN1(n8666), .IN2(n9927), .Q(n9926) );
  INVX0 U9655 ( .INP(n9589), .ZN(n9890) );
  NAND2X0 U9656 ( .IN1(n9459), .IN2(g2190), .QN(n9924) );
  NAND2X0 U9657 ( .IN1(n9928), .IN2(n9929), .QN(g30273) );
  NAND2X0 U9658 ( .IN1(n4317), .IN2(g1639), .QN(n9929) );
  NAND2X0 U9659 ( .IN1(n9870), .IN2(g6573), .QN(n9928) );
  NAND2X0 U9660 ( .IN1(n9930), .IN2(n9931), .QN(n9870) );
  NAND3X0 U9661 ( .IN1(n9484), .IN2(n9932), .IN3(n9933), .QN(n9931) );
  XOR2X1 U9662 ( .IN1(n9659), .IN2(n9657), .Q(n9933) );
  NOR2X0 U9663 ( .IN1(n9934), .IN2(n9935), .QN(n9657) );
  XOR2X1 U9664 ( .IN1(n8638), .IN2(n9201), .Q(n9935) );
  NAND2X0 U9665 ( .IN1(n9486), .IN2(g1506), .QN(n9930) );
  NAND2X0 U9666 ( .IN1(n9936), .IN2(n9937), .QN(g30272) );
  NAND2X0 U9667 ( .IN1(n4515), .IN2(g1633), .QN(n9937) );
  NAND2X0 U9668 ( .IN1(n9901), .IN2(g6782), .QN(n9936) );
  NAND2X0 U9669 ( .IN1(n9938), .IN2(n9939), .QN(g30271) );
  NAND2X0 U9670 ( .IN1(n4312), .IN2(g948), .QN(n9939) );
  NAND2X0 U9671 ( .IN1(n9910), .IN2(g6518), .QN(n9938) );
  NAND2X0 U9672 ( .IN1(n9940), .IN2(n9941), .QN(g30270) );
  NAND2X0 U9673 ( .IN1(g942), .IN2(n8096), .QN(n9941) );
  NAND2X0 U9674 ( .IN1(test_so31), .IN2(n9942), .QN(n9940) );
  NAND2X0 U9675 ( .IN1(n9943), .IN2(n9944), .QN(g30269) );
  NAND2X0 U9676 ( .IN1(n4323), .IN2(g873), .QN(n9944) );
  NAND2X0 U9677 ( .IN1(n9883), .IN2(g6368), .QN(n9943) );
  NAND2X0 U9678 ( .IN1(n9945), .IN2(n9946), .QN(n9883) );
  NAND2X0 U9679 ( .IN1(n9515), .IN2(n9947), .QN(n9946) );
  XNOR2X1 U9680 ( .IN1(n8618), .IN2(n9948), .Q(n9947) );
  NAND2X0 U9681 ( .IN1(n9513), .IN2(g785), .QN(n9945) );
  NAND2X0 U9682 ( .IN1(n9949), .IN2(n9950), .QN(g30268) );
  NAND2X0 U9683 ( .IN1(n4369), .IN2(g264), .QN(n9950) );
  NAND2X0 U9684 ( .IN1(n9951), .IN2(g165), .QN(n9949) );
  NAND2X0 U9685 ( .IN1(n9952), .IN2(n9953), .QN(g30267) );
  NAND2X0 U9686 ( .IN1(test_so13), .IN2(n4512), .QN(n9953) );
  NAND2X0 U9687 ( .IN1(n9921), .IN2(g6313), .QN(n9952) );
  NAND2X0 U9688 ( .IN1(n9954), .IN2(n9955), .QN(g30266) );
  NAND2X0 U9689 ( .IN1(n4317), .IN2(g1630), .QN(n9955) );
  NAND2X0 U9690 ( .IN1(n9901), .IN2(g6573), .QN(n9954) );
  NAND2X0 U9691 ( .IN1(n9956), .IN2(n9957), .QN(n9901) );
  NAND3X0 U9692 ( .IN1(n9484), .IN2(n9932), .IN3(n9958), .QN(n9957) );
  XOR2X1 U9693 ( .IN1(n8642), .IN2(n9959), .Q(n9958) );
  INVX0 U9694 ( .INP(n9629), .ZN(n9932) );
  NAND2X0 U9695 ( .IN1(n9486), .IN2(g1496), .QN(n9956) );
  NAND2X0 U9696 ( .IN1(n9960), .IN2(n9961), .QN(g30265) );
  NAND2X0 U9697 ( .IN1(test_so35), .IN2(n4323), .QN(n9961) );
  NAND2X0 U9698 ( .IN1(n9910), .IN2(g6368), .QN(n9960) );
  NAND2X0 U9699 ( .IN1(n9962), .IN2(n9963), .QN(n9910) );
  NAND2X0 U9700 ( .IN1(n9964), .IN2(n9515), .QN(n9963) );
  XOR2X1 U9701 ( .IN1(n8623), .IN2(n9691), .Q(n9964) );
  NOR2X0 U9702 ( .IN1(n9965), .IN2(n9966), .QN(n9691) );
  XOR2X1 U9703 ( .IN1(n9967), .IN2(n9689), .Q(n9966) );
  NAND2X0 U9704 ( .IN1(n9513), .IN2(g813), .QN(n9962) );
  NAND2X0 U9705 ( .IN1(n9968), .IN2(n9969), .QN(g30264) );
  NAND2X0 U9706 ( .IN1(n4312), .IN2(g939), .QN(n9969) );
  NAND2X0 U9707 ( .IN1(n9942), .IN2(g6518), .QN(n9968) );
  NAND2X0 U9708 ( .IN1(n9970), .IN2(n9971), .QN(g30263) );
  NAND2X0 U9709 ( .IN1(n4512), .IN2(g261), .QN(n9971) );
  NAND2X0 U9710 ( .IN1(n9951), .IN2(g6313), .QN(n9970) );
  NAND2X0 U9711 ( .IN1(n9972), .IN2(n9973), .QN(g30262) );
  NAND2X0 U9712 ( .IN1(n4369), .IN2(test_so14), .QN(n9973) );
  NAND2X0 U9713 ( .IN1(n9974), .IN2(g165), .QN(n9972) );
  NAND2X0 U9714 ( .IN1(n9975), .IN2(n9976), .QN(g30261) );
  NAND2X0 U9715 ( .IN1(n4318), .IN2(g186), .QN(n9976) );
  NAND2X0 U9716 ( .IN1(n9921), .IN2(g6231), .QN(n9975) );
  NAND2X0 U9717 ( .IN1(n9977), .IN2(n9978), .QN(n9921) );
  NAND2X0 U9718 ( .IN1(n9553), .IN2(n9979), .QN(n9978) );
  XOR2X1 U9719 ( .IN1(n4513), .IN2(n9980), .Q(n9979) );
  NAND2X0 U9720 ( .IN1(n9551), .IN2(g97), .QN(n9977) );
  NAND2X0 U9721 ( .IN1(n9981), .IN2(n9982), .QN(g30260) );
  NAND2X0 U9722 ( .IN1(n4367), .IN2(g2294), .QN(n9982) );
  NAND2X0 U9723 ( .IN1(n9983), .IN2(g2241), .QN(n9981) );
  NAND2X0 U9724 ( .IN1(n9984), .IN2(n9985), .QN(g30259) );
  NAND2X0 U9725 ( .IN1(n4323), .IN2(g936), .QN(n9985) );
  NAND2X0 U9726 ( .IN1(n9942), .IN2(g6368), .QN(n9984) );
  NAND2X0 U9727 ( .IN1(n9986), .IN2(n9987), .QN(n9942) );
  NAND2X0 U9728 ( .IN1(n9988), .IN2(n9515), .QN(n9987) );
  XOR2X1 U9729 ( .IN1(n8612), .IN2(n9989), .Q(n9988) );
  NAND2X0 U9730 ( .IN1(n9513), .IN2(g805), .QN(n9986) );
  NAND2X0 U9731 ( .IN1(n9990), .IN2(n9991), .QN(g30258) );
  NAND2X0 U9732 ( .IN1(n4318), .IN2(g258), .QN(n9991) );
  NAND2X0 U9733 ( .IN1(n9951), .IN2(g6231), .QN(n9990) );
  NAND2X0 U9734 ( .IN1(n9992), .IN2(n9993), .QN(n9951) );
  NAND2X0 U9735 ( .IN1(n9994), .IN2(n9553), .QN(n9993) );
  XOR2X1 U9736 ( .IN1(n8578), .IN2(n9712), .Q(n9994) );
  NOR2X0 U9737 ( .IN1(n9995), .IN2(n9996), .QN(n9712) );
  XOR2X1 U9738 ( .IN1(n8582), .IN2(n9699), .Q(n9996) );
  NAND2X0 U9739 ( .IN1(n9551), .IN2(g125), .QN(n9992) );
  NAND2X0 U9740 ( .IN1(n9997), .IN2(n9998), .QN(g30257) );
  NAND2X0 U9741 ( .IN1(n4512), .IN2(g252), .QN(n9998) );
  NAND2X0 U9742 ( .IN1(n9974), .IN2(g6313), .QN(n9997) );
  NAND2X0 U9743 ( .IN1(n9999), .IN2(n10000), .QN(g30256) );
  NAND2X0 U9744 ( .IN1(g2291), .IN2(n8097), .QN(n10000) );
  NAND2X0 U9745 ( .IN1(test_so73), .IN2(n9983), .QN(n9999) );
  NAND2X0 U9746 ( .IN1(n10001), .IN2(n10002), .QN(g30255) );
  NAND2X0 U9747 ( .IN1(n4368), .IN2(g1600), .QN(n10002) );
  NAND2X0 U9748 ( .IN1(n10003), .IN2(g1547), .QN(n10001) );
  NAND2X0 U9749 ( .IN1(n10004), .IN2(n10005), .QN(g30254) );
  NAND2X0 U9750 ( .IN1(n4318), .IN2(g249), .QN(n10005) );
  NAND2X0 U9751 ( .IN1(n9974), .IN2(g6231), .QN(n10004) );
  NAND2X0 U9752 ( .IN1(n10006), .IN2(n10007), .QN(n9974) );
  NAND2X0 U9753 ( .IN1(n10008), .IN2(n9553), .QN(n10007) );
  XOR2X1 U9754 ( .IN1(n8577), .IN2(n10009), .Q(n10008) );
  NAND2X0 U9755 ( .IN1(n9551), .IN2(g117), .QN(n10006) );
  NAND2X0 U9756 ( .IN1(n10010), .IN2(n10011), .QN(g30253) );
  NAND2X0 U9757 ( .IN1(n4324), .IN2(g2288), .QN(n10011) );
  NAND2X0 U9758 ( .IN1(n9983), .IN2(g6837), .QN(n10010) );
  NAND2X0 U9759 ( .IN1(n10012), .IN2(n10013), .QN(n9983) );
  NAND2X0 U9760 ( .IN1(n10014), .IN2(n9456), .QN(n10013) );
  XOR2X1 U9761 ( .IN1(n9892), .IN2(n9894), .Q(n10014) );
  NAND2X0 U9762 ( .IN1(n9927), .IN2(n10015), .QN(n9892) );
  XOR2X1 U9763 ( .IN1(n8666), .IN2(n9202), .Q(n10015) );
  NOR2X0 U9764 ( .IN1(n9827), .IN2(n10016), .QN(n9927) );
  XOR2X1 U9765 ( .IN1(n9828), .IN2(n9202), .Q(n10016) );
  INVX0 U9766 ( .INP(n8679), .ZN(n9828) );
  NAND2X0 U9767 ( .IN1(n9561), .IN2(n10017), .QN(n9827) );
  XOR2X1 U9768 ( .IN1(n8665), .IN2(n9202), .Q(n10017) );
  NOR2X0 U9769 ( .IN1(n9457), .IN2(n10018), .QN(n9561) );
  XOR2X1 U9770 ( .IN1(n9458), .IN2(n9202), .Q(n10018) );
  NAND2X0 U9771 ( .IN1(n9591), .IN2(n10019), .QN(n9457) );
  XOR2X1 U9772 ( .IN1(n9592), .IN2(n9202), .Q(n10019) );
  NOR2X0 U9773 ( .IN1(n10020), .IN2(n9867), .QN(n9591) );
  XOR2X1 U9774 ( .IN1(n9866), .IN2(n9202), .Q(n10020) );
  NAND2X0 U9775 ( .IN1(n9459), .IN2(g2195), .QN(n10012) );
  NOR2X0 U9776 ( .IN1(n9589), .IN2(n9456), .QN(n9459) );
  NOR2X0 U9777 ( .IN1(n10021), .IN2(n10022), .QN(n9456) );
  NOR2X0 U9778 ( .IN1(n10023), .IN2(n10024), .QN(n10022) );
  NOR2X0 U9779 ( .IN1(n9619), .IN2(n10025), .QN(n10024) );
  NOR2X0 U9780 ( .IN1(n10021), .IN2(n10023), .QN(n9589) );
  NAND2X0 U9781 ( .IN1(n10026), .IN2(n10027), .QN(n10023) );
  NAND2X0 U9782 ( .IN1(n10028), .IN2(n8656), .QN(n10027) );
  NAND4X0 U9783 ( .IN1(n9562), .IN2(n10029), .IN3(n10030), .IN4(n10031), .QN(
        n8656) );
  NOR3X0 U9784 ( .IN1(n8677), .IN2(n9592), .IN3(n8678), .QN(n10031) );
  INVX0 U9785 ( .INP(n10032), .ZN(n10030) );
  INVX0 U9786 ( .INP(n8667), .ZN(n10029) );
  INVX0 U9787 ( .INP(n8665), .ZN(n9562) );
  INVX0 U9788 ( .INP(n10025), .ZN(n10028) );
  NOR4X0 U9789 ( .IN1(n10032), .IN2(n9458), .IN3(n9619), .IN4(n10033), .QN(
        n10025) );
  NAND4X0 U9790 ( .IN1(n8665), .IN2(n8667), .IN3(n9592), .IN4(n8678), .QN(
        n10033) );
  INVX0 U9791 ( .INP(n4529), .ZN(n9619) );
  INVX0 U9792 ( .INP(n8677), .ZN(n9458) );
  NAND4X0 U9793 ( .IN1(n10034), .IN2(n9894), .IN3(n10035), .IN4(n9866), .QN(
        n10032) );
  INVX0 U9794 ( .INP(n8673), .ZN(n9866) );
  NOR2X0 U9795 ( .IN1(n8679), .IN2(n8672), .QN(n10035) );
  INVX0 U9796 ( .INP(n8671), .ZN(n9894) );
  INVX0 U9797 ( .INP(n8666), .ZN(n10034) );
  INVX0 U9798 ( .INP(n9867), .ZN(n10026) );
  NOR2X0 U9799 ( .IN1(n10036), .IN2(n4529), .QN(n9867) );
  INVX0 U9800 ( .INP(n9202), .ZN(n4529) );
  NAND3X0 U9801 ( .IN1(n10037), .IN2(n9718), .IN3(n10038), .QN(n10021) );
  NAND2X0 U9802 ( .IN1(n10039), .IN2(n9728), .QN(n10038) );
  NAND2X0 U9803 ( .IN1(n10040), .IN2(n9742), .QN(n10037) );
  INVX0 U9804 ( .INP(n2792), .ZN(n9742) );
  NAND2X0 U9805 ( .IN1(n10041), .IN2(n10042), .QN(n2792) );
  NAND3X0 U9806 ( .IN1(n10043), .IN2(n10044), .IN3(n10045), .QN(n10042) );
  NAND2X0 U9807 ( .IN1(n7322), .IN2(n10046), .QN(n10045) );
  NAND2X0 U9808 ( .IN1(n7325), .IN2(n10047), .QN(n10044) );
  NAND2X0 U9809 ( .IN1(n7326), .IN2(n10048), .QN(n10043) );
  NAND2X0 U9810 ( .IN1(n10049), .IN2(n10050), .QN(n10040) );
  NAND3X0 U9811 ( .IN1(n9735), .IN2(n9728), .IN3(n9796), .QN(n10050) );
  NAND2X0 U9812 ( .IN1(n10051), .IN2(n10052), .QN(g30252) );
  NAND2X0 U9813 ( .IN1(n4515), .IN2(g1597), .QN(n10052) );
  NAND2X0 U9814 ( .IN1(n10003), .IN2(g6782), .QN(n10051) );
  NAND2X0 U9815 ( .IN1(n10053), .IN2(n10054), .QN(g30251) );
  NAND2X0 U9816 ( .IN1(g906), .IN2(n8096), .QN(n10054) );
  NAND2X0 U9817 ( .IN1(test_so31), .IN2(n10055), .QN(n10053) );
  NAND2X0 U9818 ( .IN1(n10056), .IN2(n10057), .QN(g30250) );
  NAND2X0 U9819 ( .IN1(n4317), .IN2(g1594), .QN(n10057) );
  NAND2X0 U9820 ( .IN1(n10003), .IN2(g6573), .QN(n10056) );
  NAND2X0 U9821 ( .IN1(n10058), .IN2(n10059), .QN(n10003) );
  NAND2X0 U9822 ( .IN1(n10060), .IN2(n9484), .QN(n10059) );
  XOR2X1 U9823 ( .IN1(n9934), .IN2(n8638), .Q(n10060) );
  NAND2X0 U9824 ( .IN1(n9959), .IN2(n10061), .QN(n9934) );
  XOR2X1 U9825 ( .IN1(n8642), .IN2(n9201), .Q(n10061) );
  NOR2X0 U9826 ( .IN1(n9847), .IN2(n10062), .QN(n9959) );
  XNOR2X1 U9827 ( .IN1(n8653), .IN2(n9201), .Q(n10062) );
  NAND2X0 U9828 ( .IN1(n9601), .IN2(n10063), .QN(n9847) );
  XOR2X1 U9829 ( .IN1(n10064), .IN2(n9201), .Q(n10063) );
  NOR2X0 U9830 ( .IN1(n9485), .IN2(n10065), .QN(n9601) );
  XOR2X1 U9831 ( .IN1(n8650), .IN2(n4530), .Q(n10065) );
  NAND2X0 U9832 ( .IN1(n9631), .IN2(n10066), .QN(n9485) );
  XOR2X1 U9833 ( .IN1(n10067), .IN2(n9201), .Q(n10066) );
  NOR2X0 U9834 ( .IN1(n10068), .IN2(n10069), .QN(n9631) );
  XOR2X1 U9835 ( .IN1(n8651), .IN2(n4530), .Q(n10068) );
  NAND2X0 U9836 ( .IN1(n9486), .IN2(g1501), .QN(n10058) );
  NOR2X0 U9837 ( .IN1(n9629), .IN2(n9484), .QN(n9486) );
  NOR2X0 U9838 ( .IN1(n10070), .IN2(n10071), .QN(n9484) );
  NOR2X0 U9839 ( .IN1(n10072), .IN2(n10073), .QN(n10071) );
  NOR2X0 U9840 ( .IN1(n9655), .IN2(n10074), .QN(n10073) );
  INVX0 U9841 ( .INP(n10075), .ZN(n10074) );
  INVX0 U9842 ( .INP(n4530), .ZN(n9655) );
  NOR2X0 U9843 ( .IN1(n10070), .IN2(n10072), .QN(n9629) );
  NAND2X0 U9844 ( .IN1(n9907), .IN2(n10076), .QN(n10072) );
  NAND2X0 U9845 ( .IN1(n10075), .IN2(n8626), .QN(n10076) );
  NAND4X0 U9846 ( .IN1(n8641), .IN2(n10077), .IN3(n10078), .IN4(n10079), .QN(
        n8626) );
  NOR3X0 U9847 ( .IN1(n10067), .IN2(n8650), .IN3(n9200), .QN(n10079) );
  NAND4X0 U9848 ( .IN1(n10078), .IN2(n8650), .IN3(n4530), .IN4(n10080), .QN(
        n10075) );
  NOR4X0 U9849 ( .IN1(n8641), .IN2(n10077), .IN3(n8640), .IN4(n8652), .QN(
        n10080) );
  INVX0 U9850 ( .INP(n10064), .ZN(n8641) );
  INVX0 U9851 ( .INP(n10081), .ZN(n10078) );
  NAND4X0 U9852 ( .IN1(n10082), .IN2(n8638), .IN3(n10083), .IN4(n8639), .QN(
        n10081) );
  NOR2X0 U9853 ( .IN1(n8653), .IN2(n8651), .QN(n10083) );
  INVX0 U9854 ( .INP(n10084), .ZN(n8638) );
  INVX0 U9855 ( .INP(n10069), .ZN(n9907) );
  NOR2X0 U9856 ( .IN1(n8628), .IN2(n4530), .QN(n10069) );
  INVX0 U9857 ( .INP(n9201), .ZN(n4530) );
  NAND3X0 U9858 ( .IN1(n10085), .IN2(n9364), .IN3(n10086), .QN(n10070) );
  NAND2X0 U9859 ( .IN1(n10087), .IN2(n9374), .QN(n10086) );
  NAND2X0 U9860 ( .IN1(n10088), .IN2(n9388), .QN(n10085) );
  NAND3X0 U9861 ( .IN1(n10089), .IN2(n10090), .IN3(n10091), .QN(n9388) );
  NAND2X0 U9862 ( .IN1(n7323), .IN2(n10092), .QN(n10091) );
  NAND2X0 U9863 ( .IN1(n7327), .IN2(n10093), .QN(n10090) );
  NAND2X0 U9864 ( .IN1(n7328), .IN2(n10094), .QN(n10089) );
  NAND2X0 U9865 ( .IN1(n3068), .IN2(n10095), .QN(n10088) );
  NAND2X0 U9866 ( .IN1(n10096), .IN2(n9381), .QN(n10095) );
  NAND2X0 U9867 ( .IN1(n10097), .IN2(n10098), .QN(g30249) );
  NAND2X0 U9868 ( .IN1(n4312), .IN2(g903), .QN(n10098) );
  NAND2X0 U9869 ( .IN1(n10055), .IN2(g6518), .QN(n10097) );
  NAND2X0 U9870 ( .IN1(n10099), .IN2(n10100), .QN(g30248) );
  NAND2X0 U9871 ( .IN1(n4369), .IN2(g219), .QN(n10100) );
  NAND2X0 U9872 ( .IN1(n10101), .IN2(g165), .QN(n10099) );
  NAND2X0 U9873 ( .IN1(n10102), .IN2(n10103), .QN(g30247) );
  NAND2X0 U9874 ( .IN1(n4323), .IN2(g900), .QN(n10103) );
  NAND2X0 U9875 ( .IN1(n10055), .IN2(g6368), .QN(n10102) );
  NAND2X0 U9876 ( .IN1(n10104), .IN2(n10105), .QN(n10055) );
  NAND2X0 U9877 ( .IN1(n10106), .IN2(n9515), .QN(n10105) );
  INVX0 U9878 ( .INP(n10107), .ZN(n9515) );
  NAND2X0 U9879 ( .IN1(n9667), .IN2(n10108), .QN(n10107) );
  NAND2X0 U9880 ( .IN1(n9666), .IN2(n10109), .QN(n10108) );
  NAND2X0 U9881 ( .IN1(n9543), .IN2(n10110), .QN(n10109) );
  NOR2X0 U9882 ( .IN1(n9948), .IN2(n10111), .QN(n9666) );
  INVX0 U9883 ( .INP(n10112), .ZN(n10111) );
  NAND2X0 U9884 ( .IN1(n10110), .IN2(n8597), .QN(n10112) );
  NAND4X0 U9885 ( .IN1(n9517), .IN2(n9539), .IN3(n10113), .IN4(n10114), .QN(
        n8597) );
  NOR3X0 U9886 ( .IN1(n8607), .IN2(n8619), .IN3(n8620), .QN(n10114) );
  INVX0 U9887 ( .INP(n8608), .ZN(n9539) );
  NAND4X0 U9888 ( .IN1(n10113), .IN2(n8620), .IN3(n9543), .IN4(n10115), .QN(
        n10110) );
  INVX0 U9889 ( .INP(n10116), .ZN(n10115) );
  NAND4X0 U9890 ( .IN1(n8607), .IN2(n8606), .IN3(n8608), .IN4(n8619), .QN(
        n10116) );
  INVX0 U9891 ( .INP(n10117), .ZN(n10113) );
  NAND4X0 U9892 ( .IN1(n10118), .IN2(n9967), .IN3(n10119), .IN4(n9879), .QN(
        n10117) );
  NOR2X0 U9893 ( .IN1(n8623), .IN2(n8618), .QN(n10119) );
  INVX0 U9894 ( .INP(n8612), .ZN(n10118) );
  INVX0 U9895 ( .INP(n9513), .ZN(n9667) );
  XOR2X1 U9896 ( .IN1(n9965), .IN2(n9967), .Q(n10106) );
  INVX0 U9897 ( .INP(n8614), .ZN(n9967) );
  NAND2X0 U9898 ( .IN1(n9989), .IN2(n10120), .QN(n9965) );
  XOR2X1 U9899 ( .IN1(n8612), .IN2(n9689), .Q(n10120) );
  NOR2X0 U9900 ( .IN1(n9878), .IN2(n10121), .QN(n9989) );
  XOR2X1 U9901 ( .IN1(n9879), .IN2(n9689), .Q(n10121) );
  INVX0 U9902 ( .INP(n8613), .ZN(n9879) );
  NAND2X0 U9903 ( .IN1(n9640), .IN2(n10122), .QN(n9878) );
  XOR2X1 U9904 ( .IN1(n8620), .IN2(n9689), .Q(n10122) );
  NOR2X0 U9905 ( .IN1(n9516), .IN2(n10123), .QN(n9640) );
  XOR2X1 U9906 ( .IN1(n9517), .IN2(n9689), .Q(n10123) );
  INVX0 U9907 ( .INP(n8606), .ZN(n9517) );
  NAND2X0 U9908 ( .IN1(n9669), .IN2(n10124), .QN(n9516) );
  XOR2X1 U9909 ( .IN1(n8619), .IN2(n9689), .Q(n10124) );
  NOR2X0 U9910 ( .IN1(n10125), .IN2(n9948), .QN(n9669) );
  NOR2X0 U9911 ( .IN1(n10126), .IN2(n9543), .QN(n9948) );
  XNOR2X1 U9912 ( .IN1(n8618), .IN2(n9689), .Q(n10125) );
  NAND2X0 U9913 ( .IN1(n9513), .IN2(g809), .QN(n10104) );
  NAND3X0 U9914 ( .IN1(n10127), .IN2(n10128), .IN3(n10129), .QN(n9513) );
  NAND2X0 U9915 ( .IN1(n10130), .IN2(n9192), .QN(n10129) );
  NAND2X0 U9916 ( .IN1(n10131), .IN2(n9225), .QN(n10127) );
  INVX0 U9917 ( .INP(n2632), .ZN(n9225) );
  NAND2X0 U9918 ( .IN1(n10132), .IN2(n10133), .QN(n2632) );
  NAND3X0 U9919 ( .IN1(n10134), .IN2(n10135), .IN3(n10136), .QN(n10133) );
  NAND2X0 U9920 ( .IN1(n7329), .IN2(g1088), .QN(n10136) );
  NAND2X0 U9921 ( .IN1(n7330), .IN2(g5472), .QN(n10135) );
  NAND2X0 U9922 ( .IN1(n7324), .IN2(g6712), .QN(n10134) );
  NAND2X0 U9923 ( .IN1(n10137), .IN2(n10138), .QN(n10131) );
  NAND3X0 U9924 ( .IN1(n9196), .IN2(n9192), .IN3(n9195), .QN(n10138) );
  NAND2X0 U9925 ( .IN1(n10139), .IN2(n10140), .QN(g30246) );
  NAND2X0 U9926 ( .IN1(n4512), .IN2(g216), .QN(n10140) );
  NAND2X0 U9927 ( .IN1(n10101), .IN2(g6313), .QN(n10139) );
  NAND2X0 U9928 ( .IN1(n10141), .IN2(n10142), .QN(g30245) );
  NAND2X0 U9929 ( .IN1(n4318), .IN2(g213), .QN(n10142) );
  NAND2X0 U9930 ( .IN1(n10101), .IN2(g6231), .QN(n10141) );
  NAND2X0 U9931 ( .IN1(n10143), .IN2(n10144), .QN(n10101) );
  NAND2X0 U9932 ( .IN1(n10145), .IN2(n9553), .QN(n10144) );
  INVX0 U9933 ( .INP(n10146), .ZN(n9553) );
  NAND2X0 U9934 ( .IN1(n9700), .IN2(n10147), .QN(n10146) );
  NAND2X0 U9935 ( .IN1(n9698), .IN2(n10148), .QN(n10147) );
  NAND2X0 U9936 ( .IN1(n9699), .IN2(n10149), .QN(n10148) );
  NOR2X0 U9937 ( .IN1(n9980), .IN2(n10150), .QN(n9698) );
  INVX0 U9938 ( .INP(n10151), .ZN(n10150) );
  NAND2X0 U9939 ( .IN1(n10149), .IN2(n8566), .QN(n10151) );
  NAND4X0 U9940 ( .IN1(n10152), .IN2(n9711), .IN3(n10153), .IN4(n10154), .QN(
        n8566) );
  NOR3X0 U9941 ( .IN1(n10155), .IN2(n10156), .IN3(n8589), .QN(n10154) );
  NAND4X0 U9942 ( .IN1(n10153), .IN2(n8589), .IN3(n9699), .IN4(n10157), .QN(
        n10149) );
  NOR4X0 U9943 ( .IN1(n8594), .IN2(n10152), .IN3(n8583), .IN4(n9711), .QN(
        n10157) );
  NOR4X0 U9944 ( .IN1(n8582), .IN2(n8588), .IN3(n8577), .IN4(n10158), .QN(
        n10153) );
  NAND2X0 U9945 ( .IN1(n10159), .IN2(n4513), .QN(n10158) );
  INVX0 U9946 ( .INP(n9551), .ZN(n9700) );
  XNOR2X1 U9947 ( .IN1(n9995), .IN2(n8582), .Q(n10145) );
  NAND2X0 U9948 ( .IN1(n10009), .IN2(n10160), .QN(n9995) );
  XOR2X1 U9949 ( .IN1(n8577), .IN2(n9199), .Q(n10160) );
  NOR2X0 U9950 ( .IN1(n9918), .IN2(n10161), .QN(n10009) );
  XNOR2X1 U9951 ( .IN1(n8588), .IN2(n9199), .Q(n10161) );
  NAND2X0 U9952 ( .IN1(n9678), .IN2(n10162), .QN(n9918) );
  XOR2X1 U9953 ( .IN1(n10156), .IN2(n9199), .Q(n10162) );
  NOR2X0 U9954 ( .IN1(n9554), .IN2(n10163), .QN(n9678) );
  XNOR2X1 U9955 ( .IN1(n8589), .IN2(n9199), .Q(n10163) );
  NAND2X0 U9956 ( .IN1(n9702), .IN2(n10164), .QN(n9554) );
  XOR2X1 U9957 ( .IN1(n10155), .IN2(n9199), .Q(n10164) );
  NOR2X0 U9958 ( .IN1(n10165), .IN2(n9980), .QN(n9702) );
  NOR2X0 U9959 ( .IN1(n8568), .IN2(n9699), .QN(n9980) );
  INVX0 U9960 ( .INP(n9199), .ZN(n9699) );
  XOR2X1 U9961 ( .IN1(n4513), .IN2(n9199), .Q(n10165) );
  INVX0 U9962 ( .INP(n8590), .ZN(n4513) );
  NAND3X0 U9963 ( .IN1(n10166), .IN2(n10167), .IN3(n10168), .QN(n8590) );
  NAND2X0 U9964 ( .IN1(test_so13), .IN2(g6313), .QN(n10168) );
  NAND2X0 U9965 ( .IN1(g6231), .IN2(g186), .QN(n10167) );
  NAND2X0 U9966 ( .IN1(g165), .IN2(g192), .QN(n10166) );
  NAND2X0 U9967 ( .IN1(n9551), .IN2(g121), .QN(n10143) );
  NAND3X0 U9968 ( .IN1(n10169), .IN2(n9407), .IN3(n10170), .QN(n9551) );
  NAND2X0 U9969 ( .IN1(n10171), .IN2(n9417), .QN(n10170) );
  NAND2X0 U9970 ( .IN1(n10172), .IN2(n9431), .QN(n10169) );
  NAND3X0 U9971 ( .IN1(n10173), .IN2(n10174), .IN3(n10175), .QN(n9431) );
  NAND2X0 U9972 ( .IN1(n7333), .IN2(n10176), .QN(n10175) );
  NAND2X0 U9973 ( .IN1(n7332), .IN2(n10177), .QN(n10174) );
  NAND2X0 U9974 ( .IN1(n7331), .IN2(n10178), .QN(n10173) );
  NAND2X0 U9975 ( .IN1(n3128), .IN2(n10179), .QN(n10172) );
  NAND2X0 U9976 ( .IN1(n10180), .IN2(n9424), .QN(n10179) );
  NAND2X0 U9977 ( .IN1(n10181), .IN2(n10182), .QN(g30072) );
  NAND2X0 U9978 ( .IN1(g2574), .IN2(n7930), .QN(n10182) );
  NAND2X0 U9979 ( .IN1(n4543), .IN2(n10183), .QN(n10181) );
  NAND2X0 U9980 ( .IN1(n10184), .IN2(n10185), .QN(n10183) );
  NAND2X0 U9981 ( .IN1(n516), .IN2(n10186), .QN(n10185) );
  NAND2X0 U9982 ( .IN1(n10187), .IN2(n7929), .QN(n10184) );
  NAND2X0 U9983 ( .IN1(n10188), .IN2(n10189), .QN(g30061) );
  NAND2X0 U9984 ( .IN1(g2580), .IN2(n7926), .QN(n10189) );
  NAND2X0 U9985 ( .IN1(n7501), .IN2(n10190), .QN(n10188) );
  NAND2X0 U9986 ( .IN1(n10191), .IN2(n10192), .QN(n10190) );
  NAND2X0 U9987 ( .IN1(n4370), .IN2(g16437), .QN(n10192) );
  NAND2X0 U9988 ( .IN1(n531), .IN2(g7390), .QN(n10191) );
  INVX0 U9989 ( .INP(n10193), .ZN(n531) );
  NAND2X0 U9990 ( .IN1(n10194), .IN2(n10195), .QN(n10193) );
  NAND2X0 U9991 ( .IN1(g1886), .IN2(DFF_1133_n1), .QN(n10195) );
  NAND2X0 U9992 ( .IN1(n4493), .IN2(n10196), .QN(n10194) );
  NAND2X0 U9993 ( .IN1(n10197), .IN2(n10198), .QN(n10196) );
  NAND2X0 U9994 ( .IN1(n4315), .IN2(DFF_1142_n1), .QN(n10198) );
  NAND2X0 U9995 ( .IN1(n8557), .IN2(g7194), .QN(n10197) );
  NAND2X0 U9996 ( .IN1(n10199), .IN2(n10200), .QN(n8557) );
  NAND2X0 U9997 ( .IN1(g1192), .IN2(DFF_783_n1), .QN(n10200) );
  NAND2X0 U9998 ( .IN1(n4454), .IN2(n10201), .QN(n10199) );
  NAND2X0 U9999 ( .IN1(n10202), .IN2(n10203), .QN(n10201) );
  NAND2X0 U10000 ( .IN1(n4316), .IN2(DFF_792_n1), .QN(n10203) );
  NAND2X0 U10001 ( .IN1(n8556), .IN2(g6944), .QN(n10202) );
  NAND2X0 U10002 ( .IN1(n10204), .IN2(n10205), .QN(n8556) );
  NAND2X0 U10003 ( .IN1(n7418), .IN2(g506), .QN(n10205) );
  NAND3X0 U10004 ( .IN1(n8048), .IN2(n4372), .IN3(n4570), .QN(n10204) );
  NAND2X0 U10005 ( .IN1(n10206), .IN2(n10207), .QN(g30055) );
  NAND2X0 U10006 ( .IN1(n4487), .IN2(DFF_1378_n1), .QN(n10207) );
  NAND2X0 U10007 ( .IN1(n10208), .IN2(g2374), .QN(n10206) );
  NAND2X0 U10008 ( .IN1(n10209), .IN2(n10210), .QN(n10208) );
  NAND2X0 U10009 ( .IN1(n456), .IN2(g7264), .QN(n10210) );
  INVX0 U10010 ( .INP(n10211), .ZN(n456) );
  NAND2X0 U10011 ( .IN1(n10212), .IN2(n10213), .QN(n10211) );
  NAND2X0 U10012 ( .IN1(n4488), .IN2(n7978), .QN(n10213) );
  NAND3X0 U10013 ( .IN1(n10214), .IN2(n10215), .IN3(g1680), .QN(n10212) );
  NAND2X0 U10014 ( .IN1(g7014), .IN2(n457), .QN(n10215) );
  INVX0 U10015 ( .INP(n10216), .ZN(n457) );
  NAND2X0 U10016 ( .IN1(n10217), .IN2(n10218), .QN(n10216) );
  NAND2X0 U10017 ( .IN1(n4432), .IN2(n8017), .QN(n10218) );
  NAND2X0 U10018 ( .IN1(n10219), .IN2(g986), .QN(n10217) );
  NAND2X0 U10019 ( .IN1(n10220), .IN2(n10221), .QN(n10219) );
  NAND2X0 U10020 ( .IN1(n4364), .IN2(n7717), .QN(n10221) );
  INVX0 U10021 ( .INP(n10222), .ZN(n10220) );
  NOR2X0 U10022 ( .IN1(g21346), .IN2(n4364), .QN(n10222) );
  NAND2X0 U10023 ( .IN1(n4525), .IN2(g1686), .QN(n10214) );
  NAND2X0 U10024 ( .IN1(n4524), .IN2(g2380), .QN(n10209) );
  NAND2X0 U10025 ( .IN1(n10223), .IN2(n10224), .QN(g29941) );
  NAND2X0 U10026 ( .IN1(n4494), .IN2(g3105), .QN(n10224) );
  NAND2X0 U10027 ( .IN1(n516), .IN2(g3109), .QN(n10223) );
  NAND2X0 U10028 ( .IN1(n10225), .IN2(n10226), .QN(g29939) );
  NAND2X0 U10029 ( .IN1(n4383), .IN2(g3104), .QN(n10226) );
  NAND2X0 U10030 ( .IN1(n516), .IN2(g8030), .QN(n10225) );
  NAND2X0 U10031 ( .IN1(n10227), .IN2(n10228), .QN(g29936) );
  NAND2X0 U10032 ( .IN1(n4382), .IN2(g3103), .QN(n10228) );
  NAND2X0 U10033 ( .IN1(n516), .IN2(g8106), .QN(n10227) );
  INVX0 U10034 ( .INP(n10229), .ZN(n516) );
  NAND2X0 U10035 ( .IN1(n10230), .IN2(n10231), .QN(n10229) );
  NAND2X0 U10036 ( .IN1(g1880), .IN2(DFF_1099_n1), .QN(n10231) );
  NAND3X0 U10037 ( .IN1(n10232), .IN2(n10233), .IN3(n4545), .QN(n10230) );
  NAND2X0 U10038 ( .IN1(n517), .IN2(n10234), .QN(n10233) );
  NAND2X0 U10039 ( .IN1(n10235), .IN2(n7971), .QN(n10232) );
  NAND2X0 U10040 ( .IN1(n10236), .IN2(n10237), .QN(g29623) );
  NAND2X0 U10041 ( .IN1(n10238), .IN2(n4606), .QN(n10237) );
  NAND2X0 U10042 ( .IN1(n4509), .IN2(g2389), .QN(n10236) );
  NAND2X0 U10043 ( .IN1(n10239), .IN2(n10240), .QN(g29621) );
  NAND2X0 U10044 ( .IN1(n10238), .IN2(g7264), .QN(n10240) );
  NAND2X0 U10045 ( .IN1(n4524), .IN2(g2388), .QN(n10239) );
  NAND2X0 U10046 ( .IN1(n10241), .IN2(n10242), .QN(g29620) );
  NAND2X0 U10047 ( .IN1(n10243), .IN2(n4618), .QN(n10242) );
  NAND2X0 U10048 ( .IN1(n4511), .IN2(g1695), .QN(n10241) );
  NAND2X0 U10049 ( .IN1(n10244), .IN2(n10245), .QN(g29618) );
  NAND2X0 U10050 ( .IN1(n10238), .IN2(g5555), .QN(n10245) );
  INVX0 U10051 ( .INP(n10246), .ZN(n10238) );
  NAND2X0 U10052 ( .IN1(n9718), .IN2(n10247), .QN(n10246) );
  NAND2X0 U10053 ( .IN1(n10248), .IN2(n9202), .QN(n10247) );
  NAND3X0 U10054 ( .IN1(n9723), .IN2(n9719), .IN3(n9729), .QN(n9202) );
  NAND3X0 U10055 ( .IN1(n9728), .IN2(n10249), .IN3(n10049), .QN(n10248) );
  NAND2X0 U10056 ( .IN1(n10041), .IN2(n10250), .QN(n9718) );
  NAND2X0 U10057 ( .IN1(n4516), .IN2(g2387), .QN(n10244) );
  NAND2X0 U10058 ( .IN1(n10251), .IN2(n10252), .QN(g29617) );
  NAND2X0 U10059 ( .IN1(n10243), .IN2(g7014), .QN(n10252) );
  NAND2X0 U10060 ( .IN1(n4525), .IN2(g1694), .QN(n10251) );
  NAND2X0 U10061 ( .IN1(n10253), .IN2(n10254), .QN(g29616) );
  NAND2X0 U10062 ( .IN1(n4381), .IN2(g1001), .QN(n10254) );
  NAND2X0 U10063 ( .IN1(n10255), .IN2(g1088), .QN(n10253) );
  NAND2X0 U10064 ( .IN1(n10256), .IN2(n10257), .QN(g29613) );
  NAND2X0 U10065 ( .IN1(n10243), .IN2(g5511), .QN(n10257) );
  INVX0 U10066 ( .INP(n10258), .ZN(n10243) );
  NAND2X0 U10067 ( .IN1(n9364), .IN2(n10259), .QN(n10258) );
  NAND2X0 U10068 ( .IN1(n10260), .IN2(n9201), .QN(n10259) );
  NAND3X0 U10069 ( .IN1(n9369), .IN2(n9365), .IN3(n9375), .QN(n9201) );
  NAND3X0 U10070 ( .IN1(n9374), .IN2(n9812), .IN3(n10261), .QN(n10260) );
  NAND2X0 U10071 ( .IN1(n9389), .IN2(n10262), .QN(n9364) );
  NAND2X0 U10072 ( .IN1(n4518), .IN2(g1693), .QN(n10256) );
  NAND2X0 U10073 ( .IN1(n10263), .IN2(n10264), .QN(g29612) );
  NAND2X0 U10074 ( .IN1(n4364), .IN2(g1000), .QN(n10264) );
  NAND2X0 U10075 ( .IN1(n10255), .IN2(g6712), .QN(n10263) );
  NAND2X0 U10076 ( .IN1(n10265), .IN2(n10266), .QN(g29611) );
  NAND2X0 U10077 ( .IN1(n10267), .IN2(n4640), .QN(n10266) );
  NAND2X0 U10078 ( .IN1(n4506), .IN2(g314), .QN(n10265) );
  NAND2X0 U10079 ( .IN1(n10268), .IN2(n10269), .QN(g29609) );
  NAND2X0 U10080 ( .IN1(n4363), .IN2(g999), .QN(n10269) );
  NAND2X0 U10081 ( .IN1(n10255), .IN2(g5472), .QN(n10268) );
  NOR2X0 U10082 ( .IN1(n10270), .IN2(n163), .QN(n10255) );
  INVX0 U10083 ( .INP(n10128), .ZN(n163) );
  NAND2X0 U10084 ( .IN1(n10132), .IN2(n10271), .QN(n10128) );
  NOR2X0 U10085 ( .IN1(n9543), .IN2(n10272), .QN(n10270) );
  NOR3X0 U10086 ( .IN1(n9195), .IN2(n9206), .IN3(n10273), .QN(n10272) );
  INVX0 U10087 ( .INP(n9689), .ZN(n9543) );
  NAND3X0 U10088 ( .IN1(n9206), .IN2(n9194), .IN3(n9186), .QN(n9689) );
  NAND2X0 U10089 ( .IN1(n10274), .IN2(n10275), .QN(g29608) );
  NAND2X0 U10090 ( .IN1(n10267), .IN2(g6447), .QN(n10275) );
  NAND2X0 U10091 ( .IN1(n4499), .IN2(g313), .QN(n10274) );
  NAND2X0 U10092 ( .IN1(n10276), .IN2(n10277), .QN(g29606) );
  NAND2X0 U10093 ( .IN1(n10267), .IN2(g5437), .QN(n10277) );
  INVX0 U10094 ( .INP(n10278), .ZN(n10267) );
  NAND2X0 U10095 ( .IN1(n9407), .IN2(n10279), .QN(n10278) );
  NAND2X0 U10096 ( .IN1(n10280), .IN2(n9199), .QN(n10279) );
  NAND3X0 U10097 ( .IN1(n9412), .IN2(n9408), .IN3(n9418), .QN(n9199) );
  NAND3X0 U10098 ( .IN1(n9417), .IN2(n9779), .IN3(n10281), .QN(n10280) );
  NAND2X0 U10099 ( .IN1(n9432), .IN2(n10282), .QN(n9407) );
  NAND2X0 U10100 ( .IN1(n4520), .IN2(g312), .QN(n10276) );
  NOR2X0 U10101 ( .IN1(n10283), .IN2(n10284), .QN(g29582) );
  XNOR2X1 U10102 ( .IN1(n7173), .IN2(n2981), .Q(n10284) );
  NOR2X0 U10103 ( .IN1(n10285), .IN2(n10286), .QN(g29581) );
  XNOR2X1 U10104 ( .IN1(n7174), .IN2(n2984), .Q(n10286) );
  NOR2X0 U10105 ( .IN1(n10287), .IN2(n10288), .QN(g29580) );
  XNOR2X1 U10106 ( .IN1(n7175), .IN2(n2987), .Q(n10288) );
  NOR2X0 U10107 ( .IN1(n10289), .IN2(n10290), .QN(g29579) );
  XNOR2X1 U10108 ( .IN1(n7176), .IN2(n2990), .Q(n10290) );
  NOR2X0 U10109 ( .IN1(n10283), .IN2(n10291), .QN(g29357) );
  XNOR2X1 U10110 ( .IN1(n7334), .IN2(n2982), .Q(n10291) );
  NAND2X0 U10111 ( .IN1(n3159), .IN2(g2129), .QN(n2982) );
  NOR2X0 U10112 ( .IN1(n10285), .IN2(n10292), .QN(g29355) );
  XNOR2X1 U10113 ( .IN1(n7335), .IN2(n2985), .Q(n10292) );
  NAND2X0 U10114 ( .IN1(n3163), .IN2(g1435), .QN(n2985) );
  NOR2X0 U10115 ( .IN1(n10287), .IN2(n10293), .QN(g29354) );
  XNOR2X1 U10116 ( .IN1(n7336), .IN2(n2988), .Q(n10293) );
  NAND2X0 U10117 ( .IN1(n3167), .IN2(test_so36), .QN(n2988) );
  NOR2X0 U10118 ( .IN1(n10289), .IN2(n10294), .QN(g29353) );
  XNOR2X1 U10119 ( .IN1(n7337), .IN2(n2991), .Q(n10294) );
  NAND2X0 U10120 ( .IN1(n3171), .IN2(g61), .QN(n2991) );
  NAND2X0 U10121 ( .IN1(n10295), .IN2(n10296), .QN(g29226) );
  NAND2X0 U10122 ( .IN1(n10297), .IN2(n4606), .QN(n10296) );
  NAND2X0 U10123 ( .IN1(n4509), .IN2(g2498), .QN(n10295) );
  NAND2X0 U10124 ( .IN1(n10298), .IN2(n10299), .QN(g29221) );
  NAND2X0 U10125 ( .IN1(n10297), .IN2(g7264), .QN(n10299) );
  NAND2X0 U10126 ( .IN1(n4524), .IN2(g2495), .QN(n10298) );
  NAND2X0 U10127 ( .IN1(n10300), .IN2(n10301), .QN(g29218) );
  NAND2X0 U10128 ( .IN1(n10302), .IN2(n4618), .QN(n10301) );
  NAND2X0 U10129 ( .IN1(n4511), .IN2(g1804), .QN(n10300) );
  NAND2X0 U10130 ( .IN1(n10303), .IN2(n10304), .QN(g29213) );
  NAND2X0 U10131 ( .IN1(n10297), .IN2(g5555), .QN(n10304) );
  XOR2X1 U10132 ( .IN1(n10305), .IN2(n10306), .Q(n10297) );
  NAND3X0 U10133 ( .IN1(test_so79), .IN2(n10307), .IN3(n10308), .QN(n10305) );
  XOR2X1 U10134 ( .IN1(n10309), .IN2(n10306), .Q(n10308) );
  NAND2X0 U10135 ( .IN1(n10310), .IN2(n9184), .QN(n10307) );
  NAND2X0 U10136 ( .IN1(n10039), .IN2(n10306), .QN(n9184) );
  NAND2X0 U10137 ( .IN1(n10311), .IN2(n10312), .QN(n10310) );
  NAND2X0 U10138 ( .IN1(n4516), .IN2(g2492), .QN(n10303) );
  NAND2X0 U10139 ( .IN1(n10313), .IN2(n10314), .QN(g29212) );
  NAND2X0 U10140 ( .IN1(n10302), .IN2(g7014), .QN(n10314) );
  NAND2X0 U10141 ( .IN1(n4525), .IN2(g1801), .QN(n10313) );
  NAND2X0 U10142 ( .IN1(n10315), .IN2(n10316), .QN(g29209) );
  NAND2X0 U10143 ( .IN1(n4381), .IN2(g1110), .QN(n10316) );
  NAND2X0 U10144 ( .IN1(n10317), .IN2(g1088), .QN(n10315) );
  NAND2X0 U10145 ( .IN1(n10318), .IN2(n10319), .QN(g29205) );
  NAND2X0 U10146 ( .IN1(n10302), .IN2(g5511), .QN(n10319) );
  XOR2X1 U10147 ( .IN1(n10320), .IN2(n10321), .Q(n10302) );
  NAND3X0 U10148 ( .IN1(n10322), .IN2(g1690), .IN3(n10323), .QN(n10320) );
  XOR2X1 U10149 ( .IN1(n4284), .IN2(n9177), .Q(n10323) );
  NAND2X0 U10150 ( .IN1(n10324), .IN2(n9180), .QN(n10322) );
  NAND2X0 U10151 ( .IN1(n10087), .IN2(n10321), .QN(n9180) );
  NAND2X0 U10152 ( .IN1(n10325), .IN2(n10326), .QN(n10324) );
  NAND2X0 U10153 ( .IN1(n4518), .IN2(g1798), .QN(n10318) );
  NAND2X0 U10154 ( .IN1(n10327), .IN2(n10328), .QN(g29204) );
  NAND2X0 U10155 ( .IN1(n4364), .IN2(g1107), .QN(n10328) );
  NAND2X0 U10156 ( .IN1(n10317), .IN2(g6712), .QN(n10327) );
  NAND2X0 U10157 ( .IN1(n10329), .IN2(n10330), .QN(g29201) );
  NAND2X0 U10158 ( .IN1(n10331), .IN2(n4640), .QN(n10330) );
  NAND2X0 U10159 ( .IN1(n4506), .IN2(g423), .QN(n10329) );
  NAND2X0 U10160 ( .IN1(n10332), .IN2(n10333), .QN(g29198) );
  NAND2X0 U10161 ( .IN1(n4363), .IN2(g1104), .QN(n10333) );
  NAND2X0 U10162 ( .IN1(n10317), .IN2(g5472), .QN(n10332) );
  XOR2X1 U10163 ( .IN1(n10334), .IN2(n10335), .Q(n10317) );
  NAND3X0 U10164 ( .IN1(n10336), .IN2(g996), .IN3(n10337), .QN(n10334) );
  XOR2X1 U10165 ( .IN1(n10338), .IN2(n10335), .Q(n10337) );
  NAND2X0 U10166 ( .IN1(n10339), .IN2(n9176), .QN(n10336) );
  NAND2X0 U10167 ( .IN1(n10130), .IN2(n10335), .QN(n9176) );
  NAND2X0 U10168 ( .IN1(n10340), .IN2(n10341), .QN(n10339) );
  NAND2X0 U10169 ( .IN1(n10342), .IN2(n10343), .QN(g29197) );
  NAND2X0 U10170 ( .IN1(n10331), .IN2(g6447), .QN(n10343) );
  NAND2X0 U10171 ( .IN1(n4499), .IN2(g420), .QN(n10342) );
  NAND2X0 U10172 ( .IN1(n10344), .IN2(n10345), .QN(g29194) );
  NAND2X0 U10173 ( .IN1(n10331), .IN2(g5437), .QN(n10345) );
  XOR2X1 U10174 ( .IN1(n10346), .IN2(n10347), .Q(n10331) );
  NAND3X0 U10175 ( .IN1(n10348), .IN2(g309), .IN3(n10349), .QN(n10346) );
  XOR2X1 U10176 ( .IN1(n4282), .IN2(n9169), .Q(n10349) );
  NAND2X0 U10177 ( .IN1(n10350), .IN2(n9172), .QN(n10348) );
  NAND2X0 U10178 ( .IN1(n10171), .IN2(n10347), .QN(n9172) );
  NAND2X0 U10179 ( .IN1(n10351), .IN2(n10352), .QN(n10350) );
  NAND2X0 U10180 ( .IN1(n4520), .IN2(g417), .QN(n10344) );
  NAND2X0 U10181 ( .IN1(n10353), .IN2(n10354), .QN(g29187) );
  NAND2X0 U10182 ( .IN1(n10355), .IN2(g2396), .QN(n10354) );
  NAND2X0 U10183 ( .IN1(n10356), .IN2(n10047), .QN(n10355) );
  NAND2X0 U10184 ( .IN1(n10357), .IN2(n10047), .QN(n10353) );
  NAND2X0 U10185 ( .IN1(n10358), .IN2(n10359), .QN(g29185) );
  NAND2X0 U10186 ( .IN1(n10360), .IN2(g2398), .QN(n10359) );
  NAND2X0 U10187 ( .IN1(n10356), .IN2(n10046), .QN(n10360) );
  NAND2X0 U10188 ( .IN1(n10357), .IN2(n10046), .QN(n10358) );
  NAND2X0 U10189 ( .IN1(n10361), .IN2(n10362), .QN(g29184) );
  NAND2X0 U10190 ( .IN1(n10363), .IN2(g1702), .QN(n10362) );
  NAND2X0 U10191 ( .IN1(n10364), .IN2(n10093), .QN(n10363) );
  NAND2X0 U10192 ( .IN1(n10365), .IN2(n10093), .QN(n10361) );
  NAND2X0 U10193 ( .IN1(n10366), .IN2(n10367), .QN(g29182) );
  NAND2X0 U10194 ( .IN1(n10368), .IN2(g2397), .QN(n10367) );
  NAND2X0 U10195 ( .IN1(n10356), .IN2(n10048), .QN(n10368) );
  NAND2X0 U10196 ( .IN1(n10357), .IN2(n10048), .QN(n10366) );
  NOR2X0 U10197 ( .IN1(n10369), .IN2(n10356), .QN(n10357) );
  NOR2X0 U10198 ( .IN1(n10369), .IN2(n10370), .QN(n10356) );
  INVX0 U10199 ( .INP(n10371), .ZN(n10370) );
  NAND2X0 U10200 ( .IN1(n3036), .IN2(n10372), .QN(n10371) );
  NAND4X0 U10201 ( .IN1(n9796), .IN2(n10041), .IN3(n9729), .IN4(n9728), .QN(
        n10372) );
  INVX0 U10202 ( .INP(n10249), .ZN(n9796) );
  NAND2X0 U10203 ( .IN1(n9733), .IN2(n9730), .QN(n10249) );
  NAND2X0 U10204 ( .IN1(n3038), .IN2(n10373), .QN(n9730) );
  NAND3X0 U10205 ( .IN1(n10374), .IN2(n10375), .IN3(n10376), .QN(n10373) );
  NAND3X0 U10206 ( .IN1(n10377), .IN2(n10378), .IN3(n10379), .QN(n10376) );
  NAND2X0 U10207 ( .IN1(n10380), .IN2(n10381), .QN(n10377) );
  NAND3X0 U10208 ( .IN1(n10382), .IN2(n10383), .IN3(n10384), .QN(n10375) );
  NAND2X0 U10209 ( .IN1(n10385), .IN2(n10386), .QN(n10383) );
  NAND2X0 U10210 ( .IN1(n10387), .IN2(n10380), .QN(n10382) );
  NAND3X0 U10211 ( .IN1(n10388), .IN2(n10389), .IN3(n10390), .QN(n10374) );
  NAND2X0 U10212 ( .IN1(n10386), .IN2(n10380), .QN(n10389) );
  INVX0 U10213 ( .INP(n10391), .ZN(n10380) );
  INVX0 U10214 ( .INP(n10379), .ZN(n10386) );
  NAND2X0 U10215 ( .IN1(n10385), .IN2(n10381), .QN(n10388) );
  INVX0 U10216 ( .INP(n10384), .ZN(n10381) );
  NAND2X0 U10217 ( .IN1(n3038), .IN2(n10392), .QN(n9733) );
  NAND3X0 U10218 ( .IN1(n10393), .IN2(n10394), .IN3(n10395), .QN(n10392) );
  NAND3X0 U10219 ( .IN1(n10396), .IN2(n10397), .IN3(n10398), .QN(n10395) );
  NAND2X0 U10220 ( .IN1(n10399), .IN2(n10400), .QN(n10397) );
  NAND2X0 U10221 ( .IN1(n10401), .IN2(n10402), .QN(n10396) );
  NAND3X0 U10222 ( .IN1(n10403), .IN2(n10404), .IN3(n10405), .QN(n10394) );
  NAND2X0 U10223 ( .IN1(n10401), .IN2(n10400), .QN(n10404) );
  NAND2X0 U10224 ( .IN1(n10406), .IN2(n10402), .QN(n10403) );
  NAND3X0 U10225 ( .IN1(n10407), .IN2(n10408), .IN3(n10409), .QN(n10393) );
  INVX0 U10226 ( .INP(n10401), .ZN(n10409) );
  NAND2X0 U10227 ( .IN1(n10399), .IN2(n10402), .QN(n10408) );
  INVX0 U10228 ( .INP(n10410), .ZN(n10402) );
  NAND2X0 U10229 ( .IN1(n10400), .IN2(n10406), .QN(n10407) );
  INVX0 U10230 ( .INP(n10398), .ZN(n10406) );
  INVX0 U10231 ( .INP(n10411), .ZN(n10400) );
  NAND2X0 U10232 ( .IN1(n10412), .IN2(n10041), .QN(n3036) );
  INVX0 U10233 ( .INP(n10413), .ZN(n10041) );
  INVX0 U10234 ( .INP(n10414), .ZN(n10369) );
  NAND2X0 U10235 ( .IN1(n10415), .IN2(n10416), .QN(n10414) );
  NAND3X0 U10236 ( .IN1(n3038), .IN2(n9795), .IN3(n10049), .QN(n10416) );
  NAND4X0 U10237 ( .IN1(n10401), .IN2(n10399), .IN3(n10417), .IN4(n10418), 
        .QN(n9795) );
  NOR4X0 U10238 ( .IN1(n10378), .IN2(n10379), .IN3(n10391), .IN4(n10384), .QN(
        n10418) );
  XNOR2X1 U10239 ( .IN1(n8666), .IN2(n4555), .Q(n10384) );
  NAND3X0 U10240 ( .IN1(n10419), .IN2(n10420), .IN3(n10421), .QN(n8666) );
  NAND2X0 U10241 ( .IN1(test_so77), .IN2(test_so73), .QN(n10421) );
  NAND2X0 U10242 ( .IN1(g6837), .IN2(g2324), .QN(n10420) );
  NAND2X0 U10243 ( .IN1(g2241), .IN2(g2330), .QN(n10419) );
  XNOR2X1 U10244 ( .IN1(n8665), .IN2(n4389), .Q(n10391) );
  NAND3X0 U10245 ( .IN1(n10422), .IN2(n10423), .IN3(n10424), .QN(n8665) );
  NAND2X0 U10246 ( .IN1(test_so73), .IN2(g2318), .QN(n10424) );
  NAND2X0 U10247 ( .IN1(g6837), .IN2(g2315), .QN(n10423) );
  NAND2X0 U10248 ( .IN1(g2241), .IN2(g2321), .QN(n10422) );
  XNOR2X1 U10249 ( .IN1(n9592), .IN2(n4373), .Q(n10379) );
  NAND3X0 U10250 ( .IN1(n10425), .IN2(n10426), .IN3(n10427), .QN(n9592) );
  NAND2X0 U10251 ( .IN1(test_so73), .IN2(g2309), .QN(n10427) );
  NAND2X0 U10252 ( .IN1(g6837), .IN2(g2306), .QN(n10426) );
  NAND2X0 U10253 ( .IN1(g2241), .IN2(g2312), .QN(n10425) );
  NAND2X0 U10254 ( .IN1(n10387), .IN2(n10385), .QN(n10378) );
  XOR2X1 U10255 ( .IN1(n8672), .IN2(n4287), .Q(n10385) );
  NAND3X0 U10256 ( .IN1(n10428), .IN2(n10429), .IN3(n10430), .QN(n8672) );
  NAND2X0 U10257 ( .IN1(test_so73), .IN2(g2336), .QN(n10430) );
  NAND2X0 U10258 ( .IN1(g6837), .IN2(g2333), .QN(n10429) );
  NAND2X0 U10259 ( .IN1(g2241), .IN2(g2339), .QN(n10428) );
  INVX0 U10260 ( .INP(n10390), .ZN(n10387) );
  XNOR2X1 U10261 ( .IN1(n8667), .IN2(n9474), .Q(n10390) );
  NAND3X0 U10262 ( .IN1(n10431), .IN2(n10432), .IN3(n10433), .QN(n8667) );
  NAND2X0 U10263 ( .IN1(test_so73), .IN2(g2345), .QN(n10433) );
  NAND2X0 U10264 ( .IN1(g6837), .IN2(g2342), .QN(n10432) );
  NAND2X0 U10265 ( .IN1(g2241), .IN2(g2348), .QN(n10431) );
  NOR3X0 U10266 ( .IN1(n10411), .IN2(n10410), .IN3(n10398), .QN(n10417) );
  XNOR2X1 U10267 ( .IN1(n8673), .IN2(n4377), .Q(n10398) );
  NAND3X0 U10268 ( .IN1(n10434), .IN2(n10435), .IN3(n10436), .QN(n8673) );
  NAND2X0 U10269 ( .IN1(test_so76), .IN2(test_so73), .QN(n10436) );
  NAND2X0 U10270 ( .IN1(g6837), .IN2(g2261), .QN(n10435) );
  NAND2X0 U10271 ( .IN1(g2241), .IN2(g2267), .QN(n10434) );
  XNOR2X1 U10272 ( .IN1(n8671), .IN2(n4563), .Q(n10410) );
  NAND3X0 U10273 ( .IN1(n10437), .IN2(n10438), .IN3(n10439), .QN(n8671) );
  NAND2X0 U10274 ( .IN1(test_so73), .IN2(g2291), .QN(n10439) );
  NAND2X0 U10275 ( .IN1(g6837), .IN2(g2288), .QN(n10438) );
  NAND2X0 U10276 ( .IN1(g2241), .IN2(g2294), .QN(n10437) );
  XNOR2X1 U10277 ( .IN1(n8677), .IN2(n4319), .Q(n10411) );
  NAND3X0 U10278 ( .IN1(n10440), .IN2(n10441), .IN3(n10442), .QN(n8677) );
  NAND2X0 U10279 ( .IN1(test_so73), .IN2(g2273), .QN(n10442) );
  NAND2X0 U10280 ( .IN1(g6837), .IN2(g2270), .QN(n10441) );
  NAND2X0 U10281 ( .IN1(g2241), .IN2(g2276), .QN(n10440) );
  INVX0 U10282 ( .INP(n10405), .ZN(n10399) );
  XNOR2X1 U10283 ( .IN1(n8679), .IN2(n4325), .Q(n10405) );
  NAND3X0 U10284 ( .IN1(n10443), .IN2(n10444), .IN3(n10445), .QN(n8679) );
  NAND2X0 U10285 ( .IN1(test_so73), .IN2(g2282), .QN(n10445) );
  NAND2X0 U10286 ( .IN1(g6837), .IN2(g2279), .QN(n10444) );
  NAND2X0 U10287 ( .IN1(g2241), .IN2(g2285), .QN(n10443) );
  XOR2X1 U10288 ( .IN1(n8678), .IN2(n10446), .Q(n10401) );
  NAND3X0 U10289 ( .IN1(n10447), .IN2(n10448), .IN3(n10449), .QN(n8678) );
  NAND2X0 U10290 ( .IN1(test_so73), .IN2(g2300), .QN(n10449) );
  NAND2X0 U10291 ( .IN1(g6837), .IN2(g2297), .QN(n10448) );
  NAND2X0 U10292 ( .IN1(g2241), .IN2(g2303), .QN(n10447) );
  NAND2X0 U10293 ( .IN1(test_so79), .IN2(n10412), .QN(n10415) );
  NAND2X0 U10294 ( .IN1(n10450), .IN2(n10451), .QN(g29181) );
  NAND2X0 U10295 ( .IN1(n10452), .IN2(g1704), .QN(n10451) );
  NAND2X0 U10296 ( .IN1(n10364), .IN2(n10092), .QN(n10452) );
  NAND2X0 U10297 ( .IN1(n10365), .IN2(n10092), .QN(n10450) );
  NAND2X0 U10298 ( .IN1(n10453), .IN2(n10454), .QN(g29179) );
  NAND2X0 U10299 ( .IN1(n10455), .IN2(g1008), .QN(n10454) );
  NAND2X0 U10300 ( .IN1(n10456), .IN2(g1088), .QN(n10455) );
  NAND2X0 U10301 ( .IN1(n10457), .IN2(g1088), .QN(n10453) );
  NAND2X0 U10302 ( .IN1(n10458), .IN2(n10459), .QN(g29178) );
  NAND2X0 U10303 ( .IN1(n10460), .IN2(g1703), .QN(n10459) );
  NAND2X0 U10304 ( .IN1(n10364), .IN2(n10094), .QN(n10460) );
  NAND2X0 U10305 ( .IN1(n10365), .IN2(n10094), .QN(n10458) );
  NOR2X0 U10306 ( .IN1(n10461), .IN2(n10364), .QN(n10365) );
  NOR2X0 U10307 ( .IN1(n10461), .IN2(n10462), .QN(n10364) );
  INVX0 U10308 ( .INP(n10463), .ZN(n10462) );
  NAND2X0 U10309 ( .IN1(n3068), .IN2(n10464), .QN(n10463) );
  NAND2X0 U10310 ( .IN1(n10096), .IN2(n9375), .QN(n10464) );
  NOR3X0 U10311 ( .IN1(n10465), .IN2(n9369), .IN3(n9812), .QN(n10096) );
  NAND2X0 U10312 ( .IN1(n9379), .IN2(n9376), .QN(n9812) );
  NAND2X0 U10313 ( .IN1(n3070), .IN2(n10466), .QN(n9376) );
  NAND3X0 U10314 ( .IN1(n10467), .IN2(n10468), .IN3(n10469), .QN(n10466) );
  NAND3X0 U10315 ( .IN1(n10470), .IN2(n10471), .IN3(n10472), .QN(n10469) );
  NAND2X0 U10316 ( .IN1(n10473), .IN2(n10474), .QN(n10471) );
  NAND3X0 U10317 ( .IN1(n10475), .IN2(n10476), .IN3(n10477), .QN(n10468) );
  NAND2X0 U10318 ( .IN1(n10474), .IN2(n10478), .QN(n10476) );
  NAND2X0 U10319 ( .IN1(n10473), .IN2(n10479), .QN(n10475) );
  INVX0 U10320 ( .INP(n10480), .ZN(n10473) );
  NAND3X0 U10321 ( .IN1(n10481), .IN2(n10482), .IN3(n10480), .QN(n10467) );
  NAND2X0 U10322 ( .IN1(n10478), .IN2(n10479), .QN(n10482) );
  INVX0 U10323 ( .INP(n10472), .ZN(n10478) );
  NAND2X0 U10324 ( .IN1(n10474), .IN2(n10483), .QN(n10481) );
  INVX0 U10325 ( .INP(n10484), .ZN(n10474) );
  NAND2X0 U10326 ( .IN1(n3070), .IN2(n10485), .QN(n9379) );
  NAND3X0 U10327 ( .IN1(n10486), .IN2(n10487), .IN3(n10488), .QN(n10485) );
  NAND3X0 U10328 ( .IN1(n10489), .IN2(n10490), .IN3(n10491), .QN(n10488) );
  NAND2X0 U10329 ( .IN1(n10492), .IN2(n10493), .QN(n10490) );
  NAND2X0 U10330 ( .IN1(n10494), .IN2(n10495), .QN(n10489) );
  NAND3X0 U10331 ( .IN1(n10496), .IN2(n10497), .IN3(n10498), .QN(n10487) );
  NAND2X0 U10332 ( .IN1(n10494), .IN2(n10493), .QN(n10497) );
  NAND2X0 U10333 ( .IN1(n10499), .IN2(n10495), .QN(n10496) );
  NAND3X0 U10334 ( .IN1(n10500), .IN2(n10501), .IN3(n10502), .QN(n10486) );
  NAND2X0 U10335 ( .IN1(n10492), .IN2(n10495), .QN(n10501) );
  NAND2X0 U10336 ( .IN1(n10493), .IN2(n10499), .QN(n10500) );
  NAND2X0 U10337 ( .IN1(n10503), .IN2(n9389), .QN(n3068) );
  INVX0 U10338 ( .INP(n10465), .ZN(n9389) );
  INVX0 U10339 ( .INP(n10504), .ZN(n10461) );
  NAND2X0 U10340 ( .IN1(n10505), .IN2(n10506), .QN(n10504) );
  NAND2X0 U10341 ( .IN1(n10503), .IN2(g1690), .QN(n10506) );
  NAND3X0 U10342 ( .IN1(n3070), .IN2(n9810), .IN3(n10261), .QN(n10505) );
  NAND4X0 U10343 ( .IN1(n10494), .IN2(n10492), .IN3(n10507), .IN4(n10508), 
        .QN(n9810) );
  NOR4X0 U10344 ( .IN1(n10472), .IN2(n10470), .IN3(n10484), .IN4(n10480), .QN(
        n10508) );
  XNOR2X1 U10345 ( .IN1(n10509), .IN2(n10077), .Q(n10480) );
  INVX0 U10346 ( .INP(n8643), .ZN(n10077) );
  NAND3X0 U10347 ( .IN1(n10510), .IN2(n10511), .IN3(n10512), .QN(n8643) );
  NAND2X0 U10348 ( .IN1(g6782), .IN2(g1651), .QN(n10512) );
  NAND2X0 U10349 ( .IN1(g6573), .IN2(g1648), .QN(n10511) );
  NAND2X0 U10350 ( .IN1(g1547), .IN2(g1654), .QN(n10510) );
  XNOR2X1 U10351 ( .IN1(g1506), .IN2(n8639), .Q(n10484) );
  INVX0 U10352 ( .INP(n9659), .ZN(n8639) );
  NAND3X0 U10353 ( .IN1(n10513), .IN2(n10514), .IN3(n10515), .QN(n9659) );
  NAND2X0 U10354 ( .IN1(g6782), .IN2(g1642), .QN(n10515) );
  NAND2X0 U10355 ( .IN1(g6573), .IN2(g1639), .QN(n10514) );
  NAND2X0 U10356 ( .IN1(g1547), .IN2(g1645), .QN(n10513) );
  NAND2X0 U10357 ( .IN1(n10483), .IN2(n10479), .QN(n10470) );
  XOR2X1 U10358 ( .IN1(n4390), .IN2(n10064), .Q(n10479) );
  NAND3X0 U10359 ( .IN1(n10516), .IN2(n10517), .IN3(n10518), .QN(n10064) );
  NAND2X0 U10360 ( .IN1(g6782), .IN2(g1624), .QN(n10518) );
  NAND2X0 U10361 ( .IN1(test_so55), .IN2(g6573), .QN(n10517) );
  NAND2X0 U10362 ( .IN1(g1547), .IN2(g1627), .QN(n10516) );
  INVX0 U10363 ( .INP(n10477), .ZN(n10483) );
  XNOR2X1 U10364 ( .IN1(g1496), .IN2(n10082), .Q(n10477) );
  INVX0 U10365 ( .INP(n8642), .ZN(n10082) );
  NAND3X0 U10366 ( .IN1(n10519), .IN2(n10520), .IN3(n10521), .QN(n8642) );
  NAND2X0 U10367 ( .IN1(g6782), .IN2(g1633), .QN(n10521) );
  NAND2X0 U10368 ( .IN1(g6573), .IN2(g1630), .QN(n10520) );
  NAND2X0 U10369 ( .IN1(g1547), .IN2(g1636), .QN(n10519) );
  XOR2X1 U10370 ( .IN1(n4374), .IN2(n8640), .Q(n10472) );
  INVX0 U10371 ( .INP(n10067), .ZN(n8640) );
  NAND3X0 U10372 ( .IN1(n10522), .IN2(n10523), .IN3(n10524), .QN(n10067) );
  NAND2X0 U10373 ( .IN1(g6782), .IN2(g1615), .QN(n10524) );
  NAND2X0 U10374 ( .IN1(g6573), .IN2(g1612), .QN(n10523) );
  NAND2X0 U10375 ( .IN1(g1547), .IN2(g1618), .QN(n10522) );
  INVX0 U10376 ( .INP(n10525), .ZN(n10507) );
  NAND3X0 U10377 ( .IN1(n10493), .IN2(n10495), .IN3(n10499), .QN(n10525) );
  INVX0 U10378 ( .INP(n10491), .ZN(n10499) );
  XOR2X1 U10379 ( .IN1(g1471), .IN2(n8651), .Q(n10491) );
  NAND3X0 U10380 ( .IN1(n10526), .IN2(n10527), .IN3(n10528), .QN(n8651) );
  NAND2X0 U10381 ( .IN1(g6782), .IN2(g1570), .QN(n10528) );
  NAND2X0 U10382 ( .IN1(g6573), .IN2(g1567), .QN(n10527) );
  NAND2X0 U10383 ( .IN1(g1547), .IN2(g1573), .QN(n10526) );
  XOR2X1 U10384 ( .IN1(n4565), .IN2(n10084), .Q(n10495) );
  NAND3X0 U10385 ( .IN1(n10529), .IN2(n10530), .IN3(n10531), .QN(n10084) );
  NAND2X0 U10386 ( .IN1(g6782), .IN2(g1597), .QN(n10531) );
  NAND2X0 U10387 ( .IN1(g6573), .IN2(g1594), .QN(n10530) );
  NAND2X0 U10388 ( .IN1(g1547), .IN2(g1600), .QN(n10529) );
  XNOR2X1 U10389 ( .IN1(g1481), .IN2(n8650), .Q(n10493) );
  NAND3X0 U10390 ( .IN1(n10532), .IN2(n10533), .IN3(n10534), .QN(n8650) );
  NAND2X0 U10391 ( .IN1(g6782), .IN2(g1579), .QN(n10534) );
  NAND2X0 U10392 ( .IN1(g6573), .IN2(g1576), .QN(n10533) );
  NAND2X0 U10393 ( .IN1(g1547), .IN2(g1582), .QN(n10532) );
  INVX0 U10394 ( .INP(n10498), .ZN(n10492) );
  XOR2X1 U10395 ( .IN1(g1491), .IN2(n8653), .Q(n10498) );
  NAND3X0 U10396 ( .IN1(n10535), .IN2(n10536), .IN3(n10537), .QN(n8653) );
  NAND2X0 U10397 ( .IN1(g6782), .IN2(g1588), .QN(n10537) );
  NAND2X0 U10398 ( .IN1(g6573), .IN2(g1585), .QN(n10536) );
  NAND2X0 U10399 ( .IN1(g1547), .IN2(g1591), .QN(n10535) );
  INVX0 U10400 ( .INP(n10502), .ZN(n10494) );
  XNOR2X1 U10401 ( .IN1(n9660), .IN2(n8652), .Q(n10502) );
  INVX0 U10402 ( .INP(n9200), .ZN(n8652) );
  NAND3X0 U10403 ( .IN1(n10538), .IN2(n10539), .IN3(n10540), .QN(n9200) );
  NAND2X0 U10404 ( .IN1(test_so56), .IN2(g6782), .QN(n10540) );
  NAND2X0 U10405 ( .IN1(g6573), .IN2(g1603), .QN(n10539) );
  NAND2X0 U10406 ( .IN1(g1547), .IN2(g1609), .QN(n10538) );
  NAND2X0 U10407 ( .IN1(n10541), .IN2(n10542), .QN(g29173) );
  NAND2X0 U10408 ( .IN1(n10543), .IN2(g1010), .QN(n10542) );
  NAND2X0 U10409 ( .IN1(n10456), .IN2(g6712), .QN(n10543) );
  NAND2X0 U10410 ( .IN1(n10457), .IN2(g6712), .QN(n10541) );
  NAND2X0 U10411 ( .IN1(n10544), .IN2(n10545), .QN(g29172) );
  NAND2X0 U10412 ( .IN1(n10546), .IN2(g321), .QN(n10545) );
  NAND2X0 U10413 ( .IN1(n10547), .IN2(n10178), .QN(n10546) );
  NAND2X0 U10414 ( .IN1(n10548), .IN2(n10178), .QN(n10544) );
  NAND2X0 U10415 ( .IN1(n10549), .IN2(n10550), .QN(g29170) );
  NAND2X0 U10416 ( .IN1(n10551), .IN2(g1009), .QN(n10550) );
  NAND2X0 U10417 ( .IN1(n10456), .IN2(g5472), .QN(n10551) );
  INVX0 U10418 ( .INP(n155), .ZN(n10456) );
  NAND2X0 U10419 ( .IN1(n10457), .IN2(g5472), .QN(n10549) );
  INVX0 U10420 ( .INP(n10552), .ZN(n10457) );
  NAND2X0 U10421 ( .IN1(n10553), .IN2(n155), .QN(n10552) );
  NAND3X0 U10422 ( .IN1(n10553), .IN2(n10554), .IN3(n10132), .QN(n155) );
  INVX0 U10423 ( .INP(n10555), .ZN(n10132) );
  NAND2X0 U10424 ( .IN1(n10137), .IN2(n10556), .QN(n10554) );
  NAND3X0 U10425 ( .IN1(n9186), .IN2(n9192), .IN3(n9195), .QN(n10556) );
  NOR2X0 U10426 ( .IN1(n10557), .IN2(n9214), .QN(n9195) );
  INVX0 U10427 ( .INP(n9224), .ZN(n9214) );
  NAND2X0 U10428 ( .IN1(n3102), .IN2(n10558), .QN(n9224) );
  NAND3X0 U10429 ( .IN1(n10559), .IN2(n10560), .IN3(n10561), .QN(n10558) );
  NAND3X0 U10430 ( .IN1(n10562), .IN2(n10563), .IN3(n10564), .QN(n10561) );
  NAND2X0 U10431 ( .IN1(n10565), .IN2(n10566), .QN(n10563) );
  NAND2X0 U10432 ( .IN1(n10567), .IN2(n10568), .QN(n10562) );
  NAND3X0 U10433 ( .IN1(n10569), .IN2(n10570), .IN3(n10571), .QN(n10560) );
  NAND2X0 U10434 ( .IN1(n10572), .IN2(n10565), .QN(n10570) );
  NAND2X0 U10435 ( .IN1(n10568), .IN2(n10566), .QN(n10569) );
  NAND3X0 U10436 ( .IN1(n10573), .IN2(n10574), .IN3(n10575), .QN(n10559) );
  NAND2X0 U10437 ( .IN1(n10572), .IN2(n10568), .QN(n10574) );
  INVX0 U10438 ( .INP(n10576), .ZN(n10568) );
  NAND2X0 U10439 ( .IN1(n10565), .IN2(n10567), .QN(n10573) );
  INVX0 U10440 ( .INP(n10571), .ZN(n10567) );
  INVX0 U10441 ( .INP(n10577), .ZN(n10565) );
  INVX0 U10442 ( .INP(n9211), .ZN(n10557) );
  NAND2X0 U10443 ( .IN1(n3102), .IN2(n10578), .QN(n9211) );
  NAND3X0 U10444 ( .IN1(n10579), .IN2(n10580), .IN3(n10581), .QN(n10578) );
  NAND3X0 U10445 ( .IN1(n10582), .IN2(n10583), .IN3(n10584), .QN(n10581) );
  NAND2X0 U10446 ( .IN1(n10585), .IN2(n10586), .QN(n10583) );
  NAND2X0 U10447 ( .IN1(n10587), .IN2(n10588), .QN(n10582) );
  NAND3X0 U10448 ( .IN1(n10589), .IN2(n10590), .IN3(n10591), .QN(n10580) );
  NAND2X0 U10449 ( .IN1(n10585), .IN2(n10588), .QN(n10590) );
  NAND2X0 U10450 ( .IN1(n10592), .IN2(n10587), .QN(n10589) );
  NAND3X0 U10451 ( .IN1(n10593), .IN2(n10594), .IN3(n10595), .QN(n10579) );
  NAND2X0 U10452 ( .IN1(n10587), .IN2(n10586), .QN(n10593) );
  NAND2X0 U10453 ( .IN1(n10596), .IN2(n10597), .QN(n10553) );
  NAND2X0 U10454 ( .IN1(n10273), .IN2(g996), .QN(n10597) );
  NAND3X0 U10455 ( .IN1(n3102), .IN2(n9213), .IN3(n10137), .QN(n10596) );
  NAND4X0 U10456 ( .IN1(n10588), .IN2(n10586), .IN3(n10598), .IN4(n10599), 
        .QN(n9213) );
  NOR4X0 U10457 ( .IN1(n10594), .IN2(n10564), .IN3(n10600), .IN4(n10577), .QN(
        n10599) );
  XNOR2X1 U10458 ( .IN1(n8614), .IN2(n4567), .Q(n10577) );
  NAND3X0 U10459 ( .IN1(n10601), .IN2(n10602), .IN3(n10603), .QN(n8614) );
  NAND2X0 U10460 ( .IN1(test_so31), .IN2(g906), .QN(n10603) );
  NAND2X0 U10461 ( .IN1(g6518), .IN2(g903), .QN(n10602) );
  NAND2X0 U10462 ( .IN1(g6368), .IN2(g900), .QN(n10601) );
  INVX0 U10463 ( .INP(n10587), .ZN(n10600) );
  XOR2X1 U10464 ( .IN1(n8623), .IN2(n4289), .Q(n10587) );
  NAND3X0 U10465 ( .IN1(n10604), .IN2(n10605), .IN3(n10606), .QN(n8623) );
  NAND2X0 U10466 ( .IN1(test_so31), .IN2(g951), .QN(n10606) );
  NAND2X0 U10467 ( .IN1(g6518), .IN2(g948), .QN(n10605) );
  NAND2X0 U10468 ( .IN1(test_so35), .IN2(g6368), .QN(n10604) );
  INVX0 U10469 ( .INP(n10572), .ZN(n10564) );
  XOR2X1 U10470 ( .IN1(n8618), .IN2(n4379), .Q(n10572) );
  NAND3X0 U10471 ( .IN1(n10607), .IN2(n10608), .IN3(n10609), .QN(n8618) );
  NAND2X0 U10472 ( .IN1(test_so31), .IN2(g879), .QN(n10609) );
  NAND2X0 U10473 ( .IN1(g6518), .IN2(g876), .QN(n10608) );
  NAND2X0 U10474 ( .IN1(g6368), .IN2(g873), .QN(n10607) );
  NAND2X0 U10475 ( .IN1(n10592), .IN2(n10585), .QN(n10594) );
  XOR2X1 U10476 ( .IN1(n8620), .IN2(n4391), .Q(n10585) );
  NAND3X0 U10477 ( .IN1(n10610), .IN2(n10611), .IN3(n10612), .QN(n8620) );
  NAND2X0 U10478 ( .IN1(test_so31), .IN2(g933), .QN(n10612) );
  NAND2X0 U10479 ( .IN1(g6518), .IN2(g930), .QN(n10611) );
  NAND2X0 U10480 ( .IN1(g6368), .IN2(g927), .QN(n10610) );
  INVX0 U10481 ( .INP(n10584), .ZN(n10592) );
  XNOR2X1 U10482 ( .IN1(n8619), .IN2(n4375), .Q(n10584) );
  NAND3X0 U10483 ( .IN1(n10613), .IN2(n10614), .IN3(n10615), .QN(n8619) );
  NAND2X0 U10484 ( .IN1(test_so34), .IN2(test_so31), .QN(n10615) );
  NAND2X0 U10485 ( .IN1(g6518), .IN2(g921), .QN(n10614) );
  NAND2X0 U10486 ( .IN1(g6368), .IN2(g918), .QN(n10613) );
  NOR3X0 U10487 ( .IN1(n10571), .IN2(n10575), .IN3(n10576), .QN(n10598) );
  XNOR2X1 U10488 ( .IN1(n8606), .IN2(n4321), .Q(n10576) );
  NAND3X0 U10489 ( .IN1(n10616), .IN2(n10617), .IN3(n10618), .QN(n8606) );
  NAND2X0 U10490 ( .IN1(test_so31), .IN2(g888), .QN(n10618) );
  NAND2X0 U10491 ( .IN1(g6518), .IN2(g885), .QN(n10617) );
  NAND2X0 U10492 ( .IN1(g6368), .IN2(g882), .QN(n10616) );
  INVX0 U10493 ( .INP(n10566), .ZN(n10575) );
  XOR2X1 U10494 ( .IN1(n8607), .IN2(n10619), .Q(n10566) );
  NAND3X0 U10495 ( .IN1(n10620), .IN2(n10621), .IN3(n10622), .QN(n8607) );
  NAND2X0 U10496 ( .IN1(test_so31), .IN2(g915), .QN(n10622) );
  NAND2X0 U10497 ( .IN1(g6518), .IN2(g912), .QN(n10621) );
  NAND2X0 U10498 ( .IN1(g6368), .IN2(g909), .QN(n10620) );
  XNOR2X1 U10499 ( .IN1(n8613), .IN2(n4327), .Q(n10571) );
  NAND3X0 U10500 ( .IN1(n10623), .IN2(n10624), .IN3(n10625), .QN(n8613) );
  NAND2X0 U10501 ( .IN1(test_so31), .IN2(g897), .QN(n10625) );
  NAND2X0 U10502 ( .IN1(g6518), .IN2(g894), .QN(n10624) );
  NAND2X0 U10503 ( .IN1(g6368), .IN2(g891), .QN(n10623) );
  INVX0 U10504 ( .INP(n10591), .ZN(n10586) );
  XNOR2X1 U10505 ( .IN1(n8612), .IN2(n4559), .Q(n10591) );
  NAND3X0 U10506 ( .IN1(n10626), .IN2(n10627), .IN3(n10628), .QN(n8612) );
  NAND2X0 U10507 ( .IN1(test_so31), .IN2(g942), .QN(n10628) );
  NAND2X0 U10508 ( .IN1(g6518), .IN2(g939), .QN(n10627) );
  NAND2X0 U10509 ( .IN1(g6368), .IN2(g936), .QN(n10626) );
  INVX0 U10510 ( .INP(n10595), .ZN(n10588) );
  XNOR2X1 U10511 ( .IN1(n8608), .IN2(n9537), .Q(n10595) );
  NAND3X0 U10512 ( .IN1(n10629), .IN2(n10630), .IN3(n10631), .QN(n8608) );
  NAND2X0 U10513 ( .IN1(test_so31), .IN2(g960), .QN(n10631) );
  NAND2X0 U10514 ( .IN1(g6518), .IN2(g957), .QN(n10630) );
  NAND2X0 U10515 ( .IN1(g6368), .IN2(g954), .QN(n10629) );
  NAND2X0 U10516 ( .IN1(n10632), .IN2(n10633), .QN(g29169) );
  NAND2X0 U10517 ( .IN1(n10634), .IN2(g323), .QN(n10633) );
  NAND2X0 U10518 ( .IN1(n10547), .IN2(n10177), .QN(n10634) );
  NAND2X0 U10519 ( .IN1(n10548), .IN2(n10177), .QN(n10632) );
  NAND2X0 U10520 ( .IN1(n10635), .IN2(n10636), .QN(g29167) );
  NAND2X0 U10521 ( .IN1(n10637), .IN2(g322), .QN(n10636) );
  NAND2X0 U10522 ( .IN1(n10547), .IN2(n10176), .QN(n10637) );
  NAND2X0 U10523 ( .IN1(n10548), .IN2(n10176), .QN(n10635) );
  NOR2X0 U10524 ( .IN1(n10638), .IN2(n10547), .QN(n10548) );
  NOR2X0 U10525 ( .IN1(n10638), .IN2(n10639), .QN(n10547) );
  INVX0 U10526 ( .INP(n10640), .ZN(n10639) );
  NAND2X0 U10527 ( .IN1(n3128), .IN2(n10641), .QN(n10640) );
  NAND2X0 U10528 ( .IN1(n10180), .IN2(n9418), .QN(n10641) );
  NOR3X0 U10529 ( .IN1(n10642), .IN2(n9412), .IN3(n9779), .QN(n10180) );
  NAND2X0 U10530 ( .IN1(n9422), .IN2(n9419), .QN(n9779) );
  NAND2X0 U10531 ( .IN1(n3130), .IN2(n10643), .QN(n9419) );
  NAND3X0 U10532 ( .IN1(n10644), .IN2(n10645), .IN3(n10646), .QN(n10643) );
  NAND3X0 U10533 ( .IN1(n10647), .IN2(n10648), .IN3(n10649), .QN(n10646) );
  NAND2X0 U10534 ( .IN1(n10650), .IN2(n10651), .QN(n10648) );
  NAND2X0 U10535 ( .IN1(n10652), .IN2(n10653), .QN(n10647) );
  NAND3X0 U10536 ( .IN1(n10654), .IN2(n10655), .IN3(n10656), .QN(n10645) );
  INVX0 U10537 ( .INP(n10653), .ZN(n10656) );
  NAND2X0 U10538 ( .IN1(n10651), .IN2(n10657), .QN(n10655) );
  NAND2X0 U10539 ( .IN1(n10650), .IN2(n10652), .QN(n10654) );
  NAND3X0 U10540 ( .IN1(n10658), .IN2(n10659), .IN3(n10660), .QN(n10644) );
  NAND2X0 U10541 ( .IN1(n10657), .IN2(n10652), .QN(n10659) );
  NAND2X0 U10542 ( .IN1(n10651), .IN2(n10653), .QN(n10658) );
  NAND2X0 U10543 ( .IN1(n3130), .IN2(n10661), .QN(n9422) );
  NAND3X0 U10544 ( .IN1(n10662), .IN2(n10663), .IN3(n10664), .QN(n10661) );
  NAND3X0 U10545 ( .IN1(n10665), .IN2(n10666), .IN3(n10667), .QN(n10664) );
  NAND2X0 U10546 ( .IN1(n10668), .IN2(n10669), .QN(n10666) );
  NAND2X0 U10547 ( .IN1(n10670), .IN2(n10671), .QN(n10665) );
  NAND3X0 U10548 ( .IN1(n10672), .IN2(n10673), .IN3(n10674), .QN(n10663) );
  NAND2X0 U10549 ( .IN1(n10670), .IN2(n10669), .QN(n10673) );
  INVX0 U10550 ( .INP(n10675), .ZN(n10670) );
  NAND3X0 U10551 ( .IN1(n10676), .IN2(n10677), .IN3(n10675), .QN(n10662) );
  NAND2X0 U10552 ( .IN1(n10668), .IN2(n10671), .QN(n10677) );
  INVX0 U10553 ( .INP(n10674), .ZN(n10668) );
  NAND2X0 U10554 ( .IN1(n10669), .IN2(n10678), .QN(n10676) );
  INVX0 U10555 ( .INP(n10679), .ZN(n10669) );
  NAND2X0 U10556 ( .IN1(n10680), .IN2(n9432), .QN(n3128) );
  INVX0 U10557 ( .INP(n10642), .ZN(n9432) );
  INVX0 U10558 ( .INP(n10681), .ZN(n10638) );
  NAND2X0 U10559 ( .IN1(n10682), .IN2(n10683), .QN(n10681) );
  NAND2X0 U10560 ( .IN1(n10680), .IN2(g309), .QN(n10683) );
  NAND3X0 U10561 ( .IN1(n3130), .IN2(n9777), .IN3(n10281), .QN(n10682) );
  NAND4X0 U10562 ( .IN1(n10650), .IN2(n10651), .IN3(n10684), .IN4(n10685), 
        .QN(n9777) );
  NOR4X0 U10563 ( .IN1(n10679), .IN2(n10672), .IN3(n10674), .IN4(n10675), .QN(
        n10685) );
  XNOR2X1 U10564 ( .IN1(n9709), .IN2(n9711), .Q(n10675) );
  INVX0 U10565 ( .INP(n8584), .ZN(n9711) );
  NAND3X0 U10566 ( .IN1(n10686), .IN2(n10687), .IN3(n10688), .QN(n8584) );
  NAND2X0 U10567 ( .IN1(g6313), .IN2(g225), .QN(n10688) );
  NAND2X0 U10568 ( .IN1(g6231), .IN2(g222), .QN(n10687) );
  NAND2X0 U10569 ( .IN1(g165), .IN2(g228), .QN(n10686) );
  XOR2X1 U10570 ( .IN1(g113), .IN2(n8588), .Q(n10674) );
  NAND3X0 U10571 ( .IN1(n10689), .IN2(n10690), .IN3(n10691), .QN(n8588) );
  NAND2X0 U10572 ( .IN1(g6313), .IN2(g207), .QN(n10691) );
  NAND2X0 U10573 ( .IN1(g6231), .IN2(g204), .QN(n10690) );
  NAND2X0 U10574 ( .IN1(g165), .IN2(g210), .QN(n10689) );
  NAND2X0 U10575 ( .IN1(n10678), .IN2(n10671), .QN(n10672) );
  XOR2X1 U10576 ( .IN1(n4569), .IN2(n8582), .Q(n10671) );
  NAND3X0 U10577 ( .IN1(n10692), .IN2(n10693), .IN3(n10694), .QN(n8582) );
  NAND2X0 U10578 ( .IN1(g6313), .IN2(g216), .QN(n10694) );
  NAND2X0 U10579 ( .IN1(g6231), .IN2(g213), .QN(n10693) );
  NAND2X0 U10580 ( .IN1(g165), .IN2(g219), .QN(n10692) );
  INVX0 U10581 ( .INP(n10667), .ZN(n10678) );
  XOR2X1 U10582 ( .IN1(n4513), .IN2(n4380), .Q(n10667) );
  XOR2X1 U10583 ( .IN1(g105), .IN2(n8589), .Q(n10679) );
  NAND3X0 U10584 ( .IN1(n10695), .IN2(n10696), .IN3(n10697), .QN(n8589) );
  NAND2X0 U10585 ( .IN1(g6313), .IN2(g198), .QN(n10697) );
  NAND2X0 U10586 ( .IN1(g6231), .IN2(g195), .QN(n10696) );
  NAND2X0 U10587 ( .IN1(g165), .IN2(g201), .QN(n10695) );
  INVX0 U10588 ( .INP(n10698), .ZN(n10684) );
  NAND3X0 U10589 ( .IN1(n10657), .IN2(n10652), .IN3(n10653), .QN(n10698) );
  XNOR2X1 U10590 ( .IN1(n4561), .IN2(n10699), .Q(n10653) );
  INVX0 U10591 ( .INP(n8577), .ZN(n10699) );
  NAND3X0 U10592 ( .IN1(n10700), .IN2(n10701), .IN3(n10702), .QN(n8577) );
  NAND2X0 U10593 ( .IN1(g6313), .IN2(g252), .QN(n10702) );
  NAND2X0 U10594 ( .IN1(g6231), .IN2(g249), .QN(n10701) );
  NAND2X0 U10595 ( .IN1(test_so14), .IN2(g165), .QN(n10700) );
  XNOR2X1 U10596 ( .IN1(n4392), .IN2(n8594), .Q(n10652) );
  INVX0 U10597 ( .INP(n10156), .ZN(n8594) );
  NAND3X0 U10598 ( .IN1(n10703), .IN2(n10704), .IN3(n10705), .QN(n10156) );
  NAND2X0 U10599 ( .IN1(g6313), .IN2(g243), .QN(n10705) );
  NAND2X0 U10600 ( .IN1(g6231), .IN2(g240), .QN(n10704) );
  NAND2X0 U10601 ( .IN1(g165), .IN2(g246), .QN(n10703) );
  INVX0 U10602 ( .INP(n10649), .ZN(n10657) );
  XOR2X1 U10603 ( .IN1(n4376), .IN2(n8583), .Q(n10649) );
  INVX0 U10604 ( .INP(n10155), .ZN(n8583) );
  NAND3X0 U10605 ( .IN1(n10706), .IN2(n10707), .IN3(n10708), .QN(n10155) );
  NAND2X0 U10606 ( .IN1(g6313), .IN2(g234), .QN(n10708) );
  NAND2X0 U10607 ( .IN1(g6231), .IN2(g231), .QN(n10707) );
  NAND2X0 U10608 ( .IN1(g165), .IN2(g237), .QN(n10706) );
  XOR2X1 U10609 ( .IN1(g125), .IN2(n10159), .Q(n10651) );
  INVX0 U10610 ( .INP(n8578), .ZN(n10159) );
  NAND3X0 U10611 ( .IN1(n10709), .IN2(n10710), .IN3(n10711), .QN(n8578) );
  NAND2X0 U10612 ( .IN1(g6313), .IN2(g261), .QN(n10711) );
  NAND2X0 U10613 ( .IN1(g6231), .IN2(g258), .QN(n10710) );
  NAND2X0 U10614 ( .IN1(g165), .IN2(g264), .QN(n10709) );
  INVX0 U10615 ( .INP(n10660), .ZN(n10650) );
  XNOR2X1 U10616 ( .IN1(n10712), .IN2(n10152), .Q(n10660) );
  INVX0 U10617 ( .INP(n8576), .ZN(n10152) );
  NAND3X0 U10618 ( .IN1(n10713), .IN2(n10714), .IN3(n10715), .QN(n8576) );
  NAND2X0 U10619 ( .IN1(g6313), .IN2(g270), .QN(n10715) );
  NAND2X0 U10620 ( .IN1(g6231), .IN2(g267), .QN(n10714) );
  NAND2X0 U10621 ( .IN1(g165), .IN2(g273), .QN(n10713) );
  NOR2X0 U10622 ( .IN1(n10283), .IN2(n10716), .QN(g29112) );
  XOR2X1 U10623 ( .IN1(n8072), .IN2(n3159), .Q(n10716) );
  NOR2X0 U10624 ( .IN1(n10285), .IN2(n10717), .QN(g29111) );
  XOR2X1 U10625 ( .IN1(n8071), .IN2(n3163), .Q(n10717) );
  NOR2X0 U10626 ( .IN1(n10287), .IN2(n10718), .QN(g29110) );
  XNOR2X1 U10627 ( .IN1(n3167), .IN2(test_so36), .Q(n10718) );
  NOR2X0 U10628 ( .IN1(n10289), .IN2(n10719), .QN(g29109) );
  XOR2X1 U10629 ( .IN1(n8070), .IN2(n3171), .Q(n10719) );
  NAND2X0 U10630 ( .IN1(n10720), .IN2(n10721), .QN(g28788) );
  NAND2X0 U10631 ( .IN1(n10722), .IN2(g2501), .QN(n10721) );
  NAND2X0 U10632 ( .IN1(n10723), .IN2(n10047), .QN(n10722) );
  NAND2X0 U10633 ( .IN1(n10724), .IN2(n10047), .QN(n10720) );
  NAND2X0 U10634 ( .IN1(n10725), .IN2(n10726), .QN(g28783) );
  NAND2X0 U10635 ( .IN1(n10727), .IN2(g2503), .QN(n10726) );
  NAND2X0 U10636 ( .IN1(n10723), .IN2(n10046), .QN(n10727) );
  NAND2X0 U10637 ( .IN1(n10724), .IN2(n10046), .QN(n10725) );
  NAND2X0 U10638 ( .IN1(n10728), .IN2(n10729), .QN(g28782) );
  NAND2X0 U10639 ( .IN1(n4606), .IN2(n10730), .QN(n10729) );
  NAND2X0 U10640 ( .IN1(n4509), .IN2(test_so80), .QN(n10728) );
  NAND2X0 U10641 ( .IN1(n10731), .IN2(n10732), .QN(g28778) );
  NAND2X0 U10642 ( .IN1(n10733), .IN2(g1807), .QN(n10732) );
  NAND2X0 U10643 ( .IN1(n10734), .IN2(n10093), .QN(n10733) );
  NAND2X0 U10644 ( .IN1(n10735), .IN2(n10093), .QN(n10731) );
  NAND2X0 U10645 ( .IN1(n10736), .IN2(n10737), .QN(g28774) );
  NAND2X0 U10646 ( .IN1(n10738), .IN2(g2502), .QN(n10737) );
  NAND2X0 U10647 ( .IN1(n10723), .IN2(n10048), .QN(n10738) );
  INVX0 U10648 ( .INP(n10739), .ZN(n10723) );
  NAND3X0 U10649 ( .IN1(test_so79), .IN2(n10740), .IN3(n10741), .QN(n10739) );
  NAND2X0 U10650 ( .IN1(n10724), .IN2(n10048), .QN(n10736) );
  INVX0 U10651 ( .INP(n10742), .ZN(n10724) );
  NAND2X0 U10652 ( .IN1(n10743), .IN2(n10744), .QN(g28773) );
  NAND2X0 U10653 ( .IN1(g7264), .IN2(n10730), .QN(n10744) );
  NAND2X0 U10654 ( .IN1(n4524), .IN2(g2486), .QN(n10743) );
  NAND2X0 U10655 ( .IN1(n10745), .IN2(n10746), .QN(g28772) );
  NAND2X0 U10656 ( .IN1(n10747), .IN2(g1809), .QN(n10746) );
  NAND2X0 U10657 ( .IN1(n10734), .IN2(n10092), .QN(n10747) );
  NAND2X0 U10658 ( .IN1(n10735), .IN2(n10092), .QN(n10745) );
  NAND2X0 U10659 ( .IN1(n10748), .IN2(n10749), .QN(g28771) );
  NAND2X0 U10660 ( .IN1(n4618), .IN2(n10750), .QN(n10749) );
  NAND2X0 U10661 ( .IN1(n4511), .IN2(g1795), .QN(n10748) );
  NAND2X0 U10662 ( .IN1(n10751), .IN2(n10752), .QN(g28767) );
  NAND2X0 U10663 ( .IN1(n10753), .IN2(g1113), .QN(n10752) );
  NAND2X0 U10664 ( .IN1(n10754), .IN2(g1088), .QN(n10753) );
  NAND2X0 U10665 ( .IN1(n10755), .IN2(g1088), .QN(n10751) );
  NAND2X0 U10666 ( .IN1(n10756), .IN2(n10757), .QN(g28763) );
  NAND2X0 U10667 ( .IN1(g5555), .IN2(n10730), .QN(n10757) );
  NAND2X0 U10668 ( .IN1(n10742), .IN2(n10758), .QN(n10730) );
  NAND2X0 U10669 ( .IN1(n10759), .IN2(n10312), .QN(n10758) );
  NAND2X0 U10670 ( .IN1(test_so79), .IN2(n10760), .QN(n10759) );
  NAND2X0 U10671 ( .IN1(n10741), .IN2(n10740), .QN(n10760) );
  INVX0 U10672 ( .INP(n10311), .ZN(n10741) );
  NAND3X0 U10673 ( .IN1(n10761), .IN2(n10762), .IN3(n10763), .QN(n10311) );
  NAND2X0 U10674 ( .IN1(n7668), .IN2(n10046), .QN(n10763) );
  NAND2X0 U10675 ( .IN1(n7677), .IN2(n10047), .QN(n10762) );
  NAND2X0 U10676 ( .IN1(n7678), .IN2(n10048), .QN(n10761) );
  NAND3X0 U10677 ( .IN1(n9182), .IN2(n10740), .IN3(test_so79), .QN(n10742) );
  NAND2X0 U10678 ( .IN1(n10764), .IN2(n10765), .QN(n10740) );
  NAND2X0 U10679 ( .IN1(n10309), .IN2(n4285), .QN(n10765) );
  NAND3X0 U10680 ( .IN1(n9181), .IN2(n9745), .IN3(n10306), .QN(n10764) );
  INVX0 U10681 ( .INP(n10039), .ZN(n9745) );
  NOR2X0 U10682 ( .IN1(n9320), .IN2(n7718), .QN(n10039) );
  NAND3X0 U10683 ( .IN1(n10766), .IN2(n10767), .IN3(n10768), .QN(n9320) );
  NAND2X0 U10684 ( .IN1(n7589), .IN2(test_so73), .QN(n10768) );
  NAND2X0 U10685 ( .IN1(n7590), .IN2(g6837), .QN(n10767) );
  NAND2X0 U10686 ( .IN1(n7588), .IN2(g2241), .QN(n10766) );
  INVX0 U10687 ( .INP(n10309), .ZN(n9181) );
  NAND3X0 U10688 ( .IN1(n10769), .IN2(n9623), .IN3(n10770), .QN(n10309) );
  INVX0 U10689 ( .INP(n10312), .ZN(n9182) );
  NAND3X0 U10690 ( .IN1(n10771), .IN2(n10772), .IN3(n10773), .QN(n10312) );
  NAND2X0 U10691 ( .IN1(g5555), .IN2(g2483), .QN(n10773) );
  NAND2X0 U10692 ( .IN1(test_so80), .IN2(n4606), .QN(n10772) );
  NAND2X0 U10693 ( .IN1(g7264), .IN2(g2486), .QN(n10771) );
  NAND2X0 U10694 ( .IN1(n4516), .IN2(g2483), .QN(n10756) );
  NAND2X0 U10695 ( .IN1(n10774), .IN2(n10775), .QN(g28761) );
  NAND2X0 U10696 ( .IN1(n10776), .IN2(g1808), .QN(n10775) );
  NAND2X0 U10697 ( .IN1(n10734), .IN2(n10094), .QN(n10776) );
  INVX0 U10698 ( .INP(n10777), .ZN(n10734) );
  NAND3X0 U10699 ( .IN1(n10778), .IN2(g1690), .IN3(n10779), .QN(n10777) );
  NAND2X0 U10700 ( .IN1(n10735), .IN2(n10094), .QN(n10774) );
  INVX0 U10701 ( .INP(n10780), .ZN(n10735) );
  NAND2X0 U10702 ( .IN1(n10781), .IN2(n10782), .QN(g28760) );
  NAND2X0 U10703 ( .IN1(g7014), .IN2(n10750), .QN(n10782) );
  NAND2X0 U10704 ( .IN1(n4525), .IN2(g1792), .QN(n10781) );
  NAND2X0 U10705 ( .IN1(n10783), .IN2(n10784), .QN(g28759) );
  NAND2X0 U10706 ( .IN1(n10785), .IN2(g1115), .QN(n10784) );
  NAND2X0 U10707 ( .IN1(n10754), .IN2(g6712), .QN(n10785) );
  NAND2X0 U10708 ( .IN1(n10755), .IN2(g6712), .QN(n10783) );
  NAND2X0 U10709 ( .IN1(n10786), .IN2(n10787), .QN(g28758) );
  NAND2X0 U10710 ( .IN1(n4381), .IN2(g1101), .QN(n10787) );
  NAND2X0 U10711 ( .IN1(n10788), .IN2(g1088), .QN(n10786) );
  NAND2X0 U10712 ( .IN1(n10789), .IN2(n10790), .QN(g28754) );
  NAND2X0 U10713 ( .IN1(n10791), .IN2(g426), .QN(n10790) );
  NAND2X0 U10714 ( .IN1(n10792), .IN2(n10178), .QN(n10791) );
  NAND2X0 U10715 ( .IN1(n10793), .IN2(n10178), .QN(n10789) );
  NAND2X0 U10716 ( .IN1(n10794), .IN2(n10795), .QN(g28749) );
  NAND2X0 U10717 ( .IN1(g5511), .IN2(n10750), .QN(n10795) );
  NAND2X0 U10718 ( .IN1(n10780), .IN2(n10796), .QN(n10750) );
  NAND2X0 U10719 ( .IN1(n10797), .IN2(n10326), .QN(n10796) );
  NAND2X0 U10720 ( .IN1(g1690), .IN2(n10798), .QN(n10797) );
  NAND2X0 U10721 ( .IN1(n10779), .IN2(n10778), .QN(n10798) );
  INVX0 U10722 ( .INP(n10325), .ZN(n10779) );
  NAND3X0 U10723 ( .IN1(n10799), .IN2(n10800), .IN3(n10801), .QN(n10325) );
  NAND2X0 U10724 ( .IN1(n7671), .IN2(n10092), .QN(n10801) );
  NAND2X0 U10725 ( .IN1(n7682), .IN2(n10093), .QN(n10800) );
  NAND2X0 U10726 ( .IN1(n7683), .IN2(n10094), .QN(n10799) );
  NAND3X0 U10727 ( .IN1(n10778), .IN2(g1690), .IN3(n9178), .QN(n10780) );
  INVX0 U10728 ( .INP(n10326), .ZN(n9178) );
  NAND3X0 U10729 ( .IN1(n10802), .IN2(n10803), .IN3(n10804), .QN(n10326) );
  NAND2X0 U10730 ( .IN1(g5511), .IN2(g1789), .QN(n10804) );
  NAND2X0 U10731 ( .IN1(n4618), .IN2(g1795), .QN(n10803) );
  NAND2X0 U10732 ( .IN1(g7014), .IN2(g1792), .QN(n10802) );
  NAND2X0 U10733 ( .IN1(n10805), .IN2(n10806), .QN(n10778) );
  NAND2X0 U10734 ( .IN1(n10807), .IN2(n4284), .QN(n10806) );
  NAND3X0 U10735 ( .IN1(n9177), .IN2(n9393), .IN3(n10321), .QN(n10805) );
  INVX0 U10736 ( .INP(n10087), .ZN(n9393) );
  NOR2X0 U10737 ( .IN1(n8516), .IN2(n7719), .QN(n10087) );
  NAND3X0 U10738 ( .IN1(n10808), .IN2(n10809), .IN3(n10810), .QN(n8516) );
  NAND2X0 U10739 ( .IN1(n7600), .IN2(g6782), .QN(n10810) );
  NAND2X0 U10740 ( .IN1(n7601), .IN2(g6573), .QN(n10809) );
  NAND2X0 U10741 ( .IN1(n7599), .IN2(g1547), .QN(n10808) );
  INVX0 U10742 ( .INP(n10807), .ZN(n9177) );
  NAND3X0 U10743 ( .IN1(n10509), .IN2(n9660), .IN3(n10811), .QN(n10807) );
  NAND2X0 U10744 ( .IN1(n4518), .IN2(g1789), .QN(n10794) );
  NAND2X0 U10745 ( .IN1(n10812), .IN2(n10813), .QN(g28747) );
  NAND2X0 U10746 ( .IN1(n10814), .IN2(g1114), .QN(n10813) );
  NAND2X0 U10747 ( .IN1(n10754), .IN2(g5472), .QN(n10814) );
  INVX0 U10748 ( .INP(n10815), .ZN(n10754) );
  NAND3X0 U10749 ( .IN1(n10816), .IN2(g996), .IN3(n10817), .QN(n10815) );
  NAND2X0 U10750 ( .IN1(n10755), .IN2(g5472), .QN(n10812) );
  INVX0 U10751 ( .INP(n10818), .ZN(n10755) );
  NAND2X0 U10752 ( .IN1(n10819), .IN2(n10820), .QN(g28746) );
  NAND2X0 U10753 ( .IN1(n4364), .IN2(g1098), .QN(n10820) );
  NAND2X0 U10754 ( .IN1(n10788), .IN2(g6712), .QN(n10819) );
  NAND2X0 U10755 ( .IN1(n10821), .IN2(n10822), .QN(g28745) );
  NAND2X0 U10756 ( .IN1(n10823), .IN2(g428), .QN(n10822) );
  NAND2X0 U10757 ( .IN1(n10792), .IN2(n10177), .QN(n10823) );
  NAND2X0 U10758 ( .IN1(n10793), .IN2(n10177), .QN(n10821) );
  NAND2X0 U10759 ( .IN1(n10824), .IN2(n10825), .QN(g28744) );
  NAND2X0 U10760 ( .IN1(n4640), .IN2(n10826), .QN(n10825) );
  NAND2X0 U10761 ( .IN1(n4506), .IN2(g414), .QN(n10824) );
  NAND2X0 U10762 ( .IN1(n10827), .IN2(n10828), .QN(g28738) );
  NAND2X0 U10763 ( .IN1(n4363), .IN2(g1095), .QN(n10828) );
  NAND2X0 U10764 ( .IN1(n10788), .IN2(g5472), .QN(n10827) );
  NAND2X0 U10765 ( .IN1(n10818), .IN2(n10829), .QN(n10788) );
  NAND2X0 U10766 ( .IN1(n10830), .IN2(n10341), .QN(n10829) );
  NAND2X0 U10767 ( .IN1(g996), .IN2(n10831), .QN(n10830) );
  NAND2X0 U10768 ( .IN1(n10817), .IN2(n10816), .QN(n10831) );
  INVX0 U10769 ( .INP(n10340), .ZN(n10817) );
  NAND3X0 U10770 ( .IN1(n10832), .IN2(n10833), .IN3(n10834), .QN(n10340) );
  NAND2X0 U10771 ( .IN1(n7688), .IN2(g1088), .QN(n10834) );
  NAND2X0 U10772 ( .IN1(n7689), .IN2(g5472), .QN(n10833) );
  NAND2X0 U10773 ( .IN1(n7674), .IN2(g6712), .QN(n10832) );
  NAND3X0 U10774 ( .IN1(n10816), .IN2(g996), .IN3(n9174), .QN(n10818) );
  INVX0 U10775 ( .INP(n10341), .ZN(n9174) );
  NAND3X0 U10776 ( .IN1(n10835), .IN2(n10836), .IN3(n10837), .QN(n10341) );
  NAND2X0 U10777 ( .IN1(g1088), .IN2(g1101), .QN(n10837) );
  NAND2X0 U10778 ( .IN1(g5472), .IN2(g1095), .QN(n10836) );
  NAND2X0 U10779 ( .IN1(g6712), .IN2(g1098), .QN(n10835) );
  NAND2X0 U10780 ( .IN1(n10838), .IN2(n10839), .QN(n10816) );
  NAND2X0 U10781 ( .IN1(n10338), .IN2(n4283), .QN(n10839) );
  NAND3X0 U10782 ( .IN1(n9173), .IN2(n9221), .IN3(n10335), .QN(n10838) );
  INVX0 U10783 ( .INP(n10130), .ZN(n9221) );
  NOR2X0 U10784 ( .IN1(n8536), .IN2(n7720), .QN(n10130) );
  NAND3X0 U10785 ( .IN1(n10840), .IN2(n10841), .IN3(n10842), .QN(n8536) );
  NAND2X0 U10786 ( .IN1(test_so31), .IN2(n7611), .QN(n10842) );
  NAND2X0 U10787 ( .IN1(g6518), .IN2(n8117), .QN(n10841) );
  NAND2X0 U10788 ( .IN1(n7612), .IN2(g6368), .QN(n10840) );
  INVX0 U10789 ( .INP(n10338), .ZN(n9173) );
  NAND3X0 U10790 ( .IN1(n10843), .IN2(n9688), .IN3(n10844), .QN(n10338) );
  NAND2X0 U10791 ( .IN1(n10845), .IN2(n10846), .QN(g28736) );
  NAND2X0 U10792 ( .IN1(test_so17), .IN2(n10847), .QN(n10846) );
  NAND2X0 U10793 ( .IN1(n10792), .IN2(n10176), .QN(n10847) );
  INVX0 U10794 ( .INP(n10848), .ZN(n10792) );
  NAND3X0 U10795 ( .IN1(n10849), .IN2(g309), .IN3(n10850), .QN(n10848) );
  NAND2X0 U10796 ( .IN1(n10793), .IN2(n10176), .QN(n10845) );
  INVX0 U10797 ( .INP(n10851), .ZN(n10793) );
  NAND2X0 U10798 ( .IN1(n10852), .IN2(n10853), .QN(g28735) );
  NAND2X0 U10799 ( .IN1(g6447), .IN2(n10826), .QN(n10853) );
  NAND2X0 U10800 ( .IN1(n4499), .IN2(g411), .QN(n10852) );
  NAND2X0 U10801 ( .IN1(n10854), .IN2(n10855), .QN(g28732) );
  NAND2X0 U10802 ( .IN1(g5437), .IN2(n10826), .QN(n10855) );
  NAND2X0 U10803 ( .IN1(n10851), .IN2(n10856), .QN(n10826) );
  NAND2X0 U10804 ( .IN1(n10857), .IN2(n10352), .QN(n10856) );
  NAND2X0 U10805 ( .IN1(g309), .IN2(n10858), .QN(n10857) );
  NAND2X0 U10806 ( .IN1(n10850), .IN2(n10849), .QN(n10858) );
  INVX0 U10807 ( .INP(n10351), .ZN(n10850) );
  NAND3X0 U10808 ( .IN1(n10859), .IN2(n10860), .IN3(n10861), .QN(n10351) );
  NAND2X0 U10809 ( .IN1(n10176), .IN2(n8118), .QN(n10861) );
  NAND2X0 U10810 ( .IN1(n7697), .IN2(n10177), .QN(n10860) );
  NAND2X0 U10811 ( .IN1(n7696), .IN2(n10178), .QN(n10859) );
  NAND3X0 U10812 ( .IN1(n10849), .IN2(g309), .IN3(n9170), .QN(n10851) );
  INVX0 U10813 ( .INP(n10352), .ZN(n9170) );
  NAND3X0 U10814 ( .IN1(n10862), .IN2(n10863), .IN3(n10864), .QN(n10352) );
  NAND2X0 U10815 ( .IN1(g5437), .IN2(g408), .QN(n10864) );
  NAND2X0 U10816 ( .IN1(n4640), .IN2(g414), .QN(n10863) );
  NAND2X0 U10817 ( .IN1(g6447), .IN2(g411), .QN(n10862) );
  NAND2X0 U10818 ( .IN1(n10865), .IN2(n10866), .QN(n10849) );
  NAND2X0 U10819 ( .IN1(n10867), .IN2(n4282), .QN(n10866) );
  NAND3X0 U10820 ( .IN1(n9169), .IN2(n9436), .IN3(n10347), .QN(n10865) );
  INVX0 U10821 ( .INP(n10171), .ZN(n9436) );
  NOR2X0 U10822 ( .IN1(n9163), .IN2(n7721), .QN(n10171) );
  NAND3X0 U10823 ( .IN1(n10868), .IN2(n10869), .IN3(n10870), .QN(n9163) );
  NAND2X0 U10824 ( .IN1(n7623), .IN2(g6313), .QN(n10870) );
  NAND2X0 U10825 ( .IN1(n7624), .IN2(g6231), .QN(n10869) );
  NAND2X0 U10826 ( .IN1(n7622), .IN2(g165), .QN(n10868) );
  INVX0 U10827 ( .INP(n10867), .ZN(n9169) );
  NAND3X0 U10828 ( .IN1(n10712), .IN2(n9709), .IN3(n10871), .QN(n10867) );
  NAND2X0 U10829 ( .IN1(n4520), .IN2(g408), .QN(n10854) );
  NOR2X0 U10830 ( .IN1(n8548), .IN2(n10872), .QN(g28668) );
  XNOR2X1 U10831 ( .IN1(n4418), .IN2(n10873), .Q(n10872) );
  NAND2X0 U10832 ( .IN1(n10874), .IN2(g686), .QN(n10873) );
  NOR2X0 U10833 ( .IN1(n10283), .IN2(n10875), .QN(g28637) );
  XNOR2X1 U10834 ( .IN1(n7699), .IN2(n3160), .Q(n10875) );
  NAND2X0 U10835 ( .IN1(n3424), .IN2(g2138), .QN(n3160) );
  NOR2X0 U10836 ( .IN1(n10285), .IN2(n10876), .QN(g28636) );
  XNOR2X1 U10837 ( .IN1(n7703), .IN2(n3164), .Q(n10876) );
  NAND2X0 U10838 ( .IN1(n3427), .IN2(g1444), .QN(n3164) );
  NOR2X0 U10839 ( .IN1(n10287), .IN2(n10877), .QN(g28635) );
  XNOR2X1 U10840 ( .IN1(n7707), .IN2(n3168), .Q(n10877) );
  NAND2X0 U10841 ( .IN1(n3430), .IN2(g758), .QN(n3168) );
  NOR2X0 U10842 ( .IN1(n10289), .IN2(n10878), .QN(g28634) );
  XNOR2X1 U10843 ( .IN1(n7711), .IN2(n3172), .Q(n10878) );
  NAND2X0 U10844 ( .IN1(n3433), .IN2(g70), .QN(n3172) );
  NAND2X0 U10845 ( .IN1(n10879), .IN2(n10880), .QN(g28425) );
  NAND2X0 U10846 ( .IN1(n4494), .IN2(g3102), .QN(n10880) );
  NAND2X0 U10847 ( .IN1(n517), .IN2(g3109), .QN(n10879) );
  NAND2X0 U10848 ( .IN1(n10881), .IN2(n10882), .QN(g28421) );
  NAND2X0 U10849 ( .IN1(n4383), .IN2(test_so7), .QN(n10882) );
  NAND2X0 U10850 ( .IN1(n517), .IN2(g8030), .QN(n10881) );
  NAND2X0 U10851 ( .IN1(n10883), .IN2(n10884), .QN(g28420) );
  INVX0 U10852 ( .INP(n10885), .ZN(n10884) );
  NOR2X0 U10853 ( .IN1(g8106), .IN2(n4342), .QN(n10885) );
  NAND2X0 U10854 ( .IN1(n517), .IN2(g8106), .QN(n10883) );
  INVX0 U10855 ( .INP(n10886), .ZN(n517) );
  NAND2X0 U10856 ( .IN1(n10887), .IN2(n10888), .QN(n10886) );
  NAND2X0 U10857 ( .IN1(n7153), .IN2(g1186), .QN(n10888) );
  NAND3X0 U10858 ( .IN1(n10889), .IN2(n10890), .IN3(n4548), .QN(n10887) );
  NAND2X0 U10859 ( .IN1(g6750), .IN2(g21851), .QN(n10890) );
  NAND2X0 U10860 ( .IN1(n4371), .IN2(n4361), .QN(n10889) );
  NAND2X0 U10861 ( .IN1(n10891), .IN2(n10892), .QN(g28371) );
  NAND2X0 U10862 ( .IN1(n4299), .IN2(g2694), .QN(n10892) );
  NAND2X0 U10863 ( .IN1(n10893), .IN2(g2624), .QN(n10891) );
  NAND2X0 U10864 ( .IN1(n10894), .IN2(n10895), .QN(g28368) );
  NAND2X0 U10865 ( .IN1(n4370), .IN2(g2691), .QN(n10895) );
  NAND2X0 U10866 ( .IN1(n10893), .IN2(g7390), .QN(n10894) );
  NAND2X0 U10867 ( .IN1(n10896), .IN2(n10897), .QN(g28367) );
  NAND2X0 U10868 ( .IN1(n4299), .IN2(g2685), .QN(n10897) );
  NAND2X0 U10869 ( .IN1(n10898), .IN2(g2624), .QN(n10896) );
  NAND2X0 U10870 ( .IN1(n10899), .IN2(n10900), .QN(g28366) );
  NAND2X0 U10871 ( .IN1(n4366), .IN2(g2000), .QN(n10900) );
  NAND2X0 U10872 ( .IN1(n10901), .IN2(g1930), .QN(n10899) );
  NAND2X0 U10873 ( .IN1(n10902), .IN2(n10903), .QN(g28364) );
  NAND2X0 U10874 ( .IN1(n4314), .IN2(g2688), .QN(n10903) );
  NAND2X0 U10875 ( .IN1(n10893), .IN2(n10186), .QN(n10902) );
  NAND2X0 U10876 ( .IN1(n10904), .IN2(n10905), .QN(n10893) );
  NAND2X0 U10877 ( .IN1(n3252), .IN2(n10906), .QN(n10905) );
  NAND2X0 U10878 ( .IN1(n8887), .IN2(n10907), .QN(n10904) );
  NAND2X0 U10879 ( .IN1(n10908), .IN2(n10909), .QN(g28363) );
  NAND2X0 U10880 ( .IN1(n10898), .IN2(g7390), .QN(n10909) );
  NAND2X0 U10881 ( .IN1(n4370), .IN2(test_so90), .QN(n10908) );
  NAND2X0 U10882 ( .IN1(n10910), .IN2(n10911), .QN(g28362) );
  NAND2X0 U10883 ( .IN1(n4315), .IN2(g1997), .QN(n10911) );
  NAND2X0 U10884 ( .IN1(n10901), .IN2(g7194), .QN(n10910) );
  NAND2X0 U10885 ( .IN1(n10912), .IN2(n10913), .QN(g28361) );
  NAND2X0 U10886 ( .IN1(n4366), .IN2(g1991), .QN(n10913) );
  NAND2X0 U10887 ( .IN1(n10914), .IN2(g1930), .QN(n10912) );
  NAND2X0 U10888 ( .IN1(n10915), .IN2(n10916), .QN(g28360) );
  NAND2X0 U10889 ( .IN1(n4300), .IN2(g1306), .QN(n10916) );
  NAND2X0 U10890 ( .IN1(n10917), .IN2(g1236), .QN(n10915) );
  NAND2X0 U10891 ( .IN1(n10918), .IN2(n10919), .QN(g28358) );
  NAND2X0 U10892 ( .IN1(g7302), .IN2(n10898), .QN(n10919) );
  NAND2X0 U10893 ( .IN1(n10920), .IN2(n10921), .QN(n10898) );
  NAND2X0 U10894 ( .IN1(n8876), .IN2(n10907), .QN(n10921) );
  NAND4X0 U10895 ( .IN1(n10922), .IN2(n9165), .IN3(n9167), .IN4(n10906), .QN(
        n10920) );
  INVX0 U10896 ( .INP(n10923), .ZN(n9167) );
  NAND3X0 U10897 ( .IN1(n10924), .IN2(n10925), .IN3(n10926), .QN(n10923) );
  NAND3X0 U10898 ( .IN1(n10927), .IN2(n10928), .IN3(n10929), .QN(n10926) );
  NAND2X0 U10899 ( .IN1(n10930), .IN2(n10931), .QN(n10929) );
  NAND2X0 U10900 ( .IN1(n10932), .IN2(n10933), .QN(n10931) );
  NAND2X0 U10901 ( .IN1(n10934), .IN2(n10935), .QN(n10928) );
  NAND2X0 U10902 ( .IN1(n10936), .IN2(n10937), .QN(n10927) );
  NAND2X0 U10903 ( .IN1(n10938), .IN2(n10939), .QN(n10936) );
  NAND2X0 U10904 ( .IN1(n10940), .IN2(n10933), .QN(n10925) );
  NAND2X0 U10905 ( .IN1(n10941), .IN2(n10942), .QN(n10940) );
  NAND2X0 U10906 ( .IN1(n10943), .IN2(n10944), .QN(n10942) );
  NAND2X0 U10907 ( .IN1(n10945), .IN2(n10946), .QN(n10943) );
  NAND2X0 U10908 ( .IN1(n10947), .IN2(n10948), .QN(n10946) );
  NAND2X0 U10909 ( .IN1(n10949), .IN2(n10950), .QN(n10941) );
  NAND2X0 U10910 ( .IN1(n10951), .IN2(n10952), .QN(n10924) );
  NAND2X0 U10911 ( .IN1(n10953), .IN2(n10954), .QN(n10952) );
  NAND2X0 U10912 ( .IN1(n10955), .IN2(n10956), .QN(n10954) );
  NAND2X0 U10913 ( .IN1(n10957), .IN2(n10958), .QN(n10956) );
  NAND3X0 U10914 ( .IN1(n10930), .IN2(n10959), .IN3(n10947), .QN(n10958) );
  INVX0 U10915 ( .INP(n10949), .ZN(n10957) );
  NAND2X0 U10916 ( .IN1(n10960), .IN2(n10961), .QN(n10949) );
  NAND2X0 U10917 ( .IN1(n10938), .IN2(n10937), .QN(n10961) );
  NAND2X0 U10918 ( .IN1(n10962), .IN2(n10934), .QN(n10960) );
  NAND2X0 U10919 ( .IN1(n10963), .IN2(n10964), .QN(n10953) );
  NAND2X0 U10920 ( .IN1(n10939), .IN2(n10965), .QN(n10963) );
  NAND2X0 U10921 ( .IN1(n10935), .IN2(n10937), .QN(n10965) );
  NAND2X0 U10922 ( .IN1(n9168), .IN2(n10966), .QN(n9165) );
  NAND2X0 U10923 ( .IN1(n1396), .IN2(n10967), .QN(n10922) );
  INVX0 U10924 ( .INP(n10966), .ZN(n10967) );
  INVX0 U10925 ( .INP(n10968), .ZN(n1396) );
  NAND3X0 U10926 ( .IN1(n10969), .IN2(n10970), .IN3(n10971), .QN(n10968) );
  NAND2X0 U10927 ( .IN1(n10972), .IN2(n10937), .QN(n10971) );
  NAND2X0 U10928 ( .IN1(n10973), .IN2(n10974), .QN(n10972) );
  NAND3X0 U10929 ( .IN1(n10955), .IN2(n10930), .IN3(n10975), .QN(n10974) );
  INVX0 U10930 ( .INP(n10935), .ZN(n10975) );
  NAND2X0 U10931 ( .IN1(n10951), .IN2(n10976), .QN(n10973) );
  NAND3X0 U10932 ( .IN1(n10977), .IN2(n10978), .IN3(n10979), .QN(n10976) );
  NAND2X0 U10933 ( .IN1(n10947), .IN2(n10944), .QN(n10979) );
  NAND3X0 U10934 ( .IN1(n10959), .IN2(n10950), .IN3(n10935), .QN(n10978) );
  NAND2X0 U10935 ( .IN1(n10980), .IN2(n10962), .QN(n10977) );
  NAND3X0 U10936 ( .IN1(n10981), .IN2(n10944), .IN3(n10938), .QN(n10970) );
  NAND2X0 U10937 ( .IN1(n10982), .IN2(n10983), .QN(n10981) );
  NAND2X0 U10938 ( .IN1(n10934), .IN2(n10939), .QN(n10983) );
  NAND2X0 U10939 ( .IN1(n10951), .IN2(n10930), .QN(n10982) );
  INVX0 U10940 ( .INP(n10933), .ZN(n10951) );
  NAND2X0 U10941 ( .IN1(n10984), .IN2(n10933), .QN(n10969) );
  NAND3X0 U10942 ( .IN1(n10985), .IN2(n10986), .IN3(n10987), .QN(n10933) );
  NAND2X0 U10943 ( .IN1(g5796), .IN2(g2426), .QN(n10987) );
  NAND2X0 U10944 ( .IN1(g5747), .IN2(g2424), .QN(n10986) );
  NAND2X0 U10945 ( .IN1(g2412), .IN2(g2428), .QN(n10985) );
  NAND2X0 U10946 ( .IN1(n10988), .IN2(n10989), .QN(n10984) );
  NAND2X0 U10947 ( .IN1(n10962), .IN2(n10964), .QN(n10989) );
  NOR2X0 U10948 ( .IN1(n10947), .IN2(n10938), .QN(n10962) );
  NAND2X0 U10949 ( .IN1(n10934), .IN2(n10990), .QN(n10988) );
  NAND3X0 U10950 ( .IN1(n10948), .IN2(n10991), .IN3(n10992), .QN(n10990) );
  NAND2X0 U10951 ( .IN1(n10980), .IN2(n10947), .QN(n10992) );
  INVX0 U10952 ( .INP(n10939), .ZN(n10947) );
  NAND3X0 U10953 ( .IN1(n10993), .IN2(n10994), .IN3(n10995), .QN(n10939) );
  NAND2X0 U10954 ( .IN1(g5796), .IN2(g2456), .QN(n10995) );
  NAND2X0 U10955 ( .IN1(g5747), .IN2(g2454), .QN(n10994) );
  NAND2X0 U10956 ( .IN1(g2412), .IN2(g2458), .QN(n10993) );
  NAND2X0 U10957 ( .IN1(n10996), .IN2(n10955), .QN(n10991) );
  INVX0 U10958 ( .INP(n10945), .ZN(n10996) );
  NAND3X0 U10959 ( .IN1(n10935), .IN2(n10959), .IN3(n10930), .QN(n10945) );
  NAND3X0 U10960 ( .IN1(n10997), .IN2(n10998), .IN3(n10999), .QN(n10935) );
  NAND2X0 U10961 ( .IN1(g5796), .IN2(g2471), .QN(n10999) );
  NAND2X0 U10962 ( .IN1(g5747), .IN2(g2469), .QN(n10998) );
  NAND2X0 U10963 ( .IN1(test_so85), .IN2(g2412), .QN(n10997) );
  NAND2X0 U10964 ( .IN1(n10938), .IN2(n10950), .QN(n10948) );
  INVX0 U10965 ( .INP(n10959), .ZN(n10938) );
  NAND3X0 U10966 ( .IN1(n11000), .IN2(n11001), .IN3(n11002), .QN(n10959) );
  NAND2X0 U10967 ( .IN1(g5796), .IN2(g2441), .QN(n11002) );
  NAND2X0 U10968 ( .IN1(g5747), .IN2(g2439), .QN(n11001) );
  NAND2X0 U10969 ( .IN1(g2412), .IN2(g2443), .QN(n11000) );
  NAND2X0 U10970 ( .IN1(n4314), .IN2(g2679), .QN(n10918) );
  NAND2X0 U10971 ( .IN1(n11003), .IN2(n11004), .QN(g28357) );
  NAND2X0 U10972 ( .IN1(n4296), .IN2(g1994), .QN(n11004) );
  NAND2X0 U10973 ( .IN1(n10901), .IN2(n10234), .QN(n11003) );
  NAND2X0 U10974 ( .IN1(n11005), .IN2(n11006), .QN(n10901) );
  NAND2X0 U10975 ( .IN1(n9011), .IN2(n10907), .QN(n11006) );
  NAND4X0 U10976 ( .IN1(n11007), .IN2(n11008), .IN3(n11009), .IN4(n10906), 
        .QN(n11005) );
  NAND2X0 U10977 ( .IN1(n11010), .IN2(n11011), .QN(n11007) );
  INVX0 U10978 ( .INP(n11012), .ZN(n11010) );
  NAND2X0 U10979 ( .IN1(n11013), .IN2(n11014), .QN(g28356) );
  NAND2X0 U10980 ( .IN1(n4315), .IN2(g1988), .QN(n11014) );
  NAND2X0 U10981 ( .IN1(n10914), .IN2(g7194), .QN(n11013) );
  NAND2X0 U10982 ( .IN1(n11015), .IN2(n11016), .QN(g28355) );
  NAND2X0 U10983 ( .IN1(n4316), .IN2(g1303), .QN(n11016) );
  NAND2X0 U10984 ( .IN1(n10917), .IN2(g6944), .QN(n11015) );
  NAND2X0 U10985 ( .IN1(n11017), .IN2(n11018), .QN(g28354) );
  NAND2X0 U10986 ( .IN1(n4300), .IN2(g1297), .QN(n11018) );
  NAND2X0 U10987 ( .IN1(n11019), .IN2(g1236), .QN(n11017) );
  NAND2X0 U10988 ( .IN1(n11020), .IN2(n11021), .QN(g28353) );
  NAND2X0 U10989 ( .IN1(n11022), .IN2(g550), .QN(n11021) );
  NAND2X0 U10990 ( .IN1(test_so26), .IN2(n4313), .QN(n11020) );
  NAND2X0 U10991 ( .IN1(n11023), .IN2(n11024), .QN(g28352) );
  NAND2X0 U10992 ( .IN1(g7052), .IN2(n10914), .QN(n11024) );
  NAND2X0 U10993 ( .IN1(n11025), .IN2(n11026), .QN(n10914) );
  NAND2X0 U10994 ( .IN1(n8989), .IN2(n10907), .QN(n11026) );
  NAND4X0 U10995 ( .IN1(n11008), .IN2(n11027), .IN3(n11011), .IN4(n10906), 
        .QN(n11025) );
  INVX0 U10996 ( .INP(n11028), .ZN(n11011) );
  NAND4X0 U10997 ( .IN1(n11029), .IN2(n11030), .IN3(n11031), .IN4(n11032), 
        .QN(n11028) );
  NAND2X0 U10998 ( .IN1(n11033), .IN2(n11034), .QN(n11032) );
  NAND2X0 U10999 ( .IN1(n11035), .IN2(n11036), .QN(n11034) );
  NAND2X0 U11000 ( .IN1(n11037), .IN2(n11038), .QN(n11036) );
  INVX0 U11001 ( .INP(n11039), .ZN(n11038) );
  NAND2X0 U11002 ( .IN1(n11040), .IN2(n11041), .QN(n11035) );
  NAND3X0 U11003 ( .IN1(n11042), .IN2(n11043), .IN3(n11044), .QN(n11031) );
  NAND2X0 U11004 ( .IN1(n11039), .IN2(n11045), .QN(n11043) );
  NAND2X0 U11005 ( .IN1(n11041), .IN2(n11046), .QN(n11045) );
  NAND2X0 U11006 ( .IN1(n11047), .IN2(n11048), .QN(n11041) );
  NAND2X0 U11007 ( .IN1(n11049), .IN2(n11050), .QN(n11048) );
  NOR2X0 U11008 ( .IN1(n11051), .IN2(n11052), .QN(n11039) );
  NOR2X0 U11009 ( .IN1(n11053), .IN2(n11050), .QN(n11052) );
  NOR2X0 U11010 ( .IN1(n11047), .IN2(n11054), .QN(n11051) );
  NAND2X0 U11011 ( .IN1(n11054), .IN2(n11055), .QN(n11030) );
  NAND2X0 U11012 ( .IN1(n11056), .IN2(n11057), .QN(n11055) );
  NAND3X0 U11013 ( .IN1(n11058), .IN2(n11059), .IN3(n11060), .QN(n11057) );
  NAND2X0 U11014 ( .IN1(n11061), .IN2(n11062), .QN(n11056) );
  NAND2X0 U11015 ( .IN1(n11046), .IN2(n11063), .QN(n11061) );
  NAND2X0 U11016 ( .IN1(n11064), .IN2(n11044), .QN(n11063) );
  NAND3X0 U11017 ( .IN1(n11065), .IN2(n11053), .IN3(n11050), .QN(n11029) );
  NAND2X0 U11018 ( .IN1(n11066), .IN2(n11067), .QN(n11065) );
  NAND2X0 U11019 ( .IN1(n11047), .IN2(n11068), .QN(n11067) );
  NAND2X0 U11020 ( .IN1(n11046), .IN2(n11069), .QN(n11068) );
  NAND2X0 U11021 ( .IN1(n11060), .IN2(n11059), .QN(n11066) );
  NAND2X0 U11022 ( .IN1(n11070), .IN2(n11009), .QN(n11027) );
  INVX0 U11023 ( .INP(n11071), .ZN(n11009) );
  NAND3X0 U11024 ( .IN1(n11072), .IN2(n11073), .IN3(n11074), .QN(n11071) );
  NAND2X0 U11025 ( .IN1(n11075), .IN2(n11044), .QN(n11074) );
  NAND2X0 U11026 ( .IN1(n11076), .IN2(n11077), .QN(n11075) );
  NAND2X0 U11027 ( .IN1(n11040), .IN2(n11058), .QN(n11077) );
  INVX0 U11028 ( .INP(n11064), .ZN(n11040) );
  NAND2X0 U11029 ( .IN1(n11054), .IN2(n11078), .QN(n11076) );
  NAND3X0 U11030 ( .IN1(n11079), .IN2(n11080), .IN3(n11081), .QN(n11078) );
  NAND2X0 U11031 ( .IN1(n11060), .IN2(n11053), .QN(n11081) );
  NAND2X0 U11032 ( .IN1(n11082), .IN2(n11083), .QN(n11080) );
  NAND2X0 U11033 ( .IN1(n11084), .IN2(n11037), .QN(n11079) );
  NAND3X0 U11034 ( .IN1(n11085), .IN2(n11053), .IN3(n11042), .QN(n11073) );
  NAND2X0 U11035 ( .IN1(n11086), .IN2(n11087), .QN(n11085) );
  NAND2X0 U11036 ( .IN1(n11033), .IN2(n11046), .QN(n11087) );
  NAND2X0 U11037 ( .IN1(n11054), .IN2(n11047), .QN(n11086) );
  INVX0 U11038 ( .INP(n11050), .ZN(n11054) );
  NAND2X0 U11039 ( .IN1(n11088), .IN2(n11050), .QN(n11072) );
  NAND3X0 U11040 ( .IN1(n11089), .IN2(n11090), .IN3(n11091), .QN(n11050) );
  NAND2X0 U11041 ( .IN1(test_so63), .IN2(g1730), .QN(n11091) );
  NAND2X0 U11042 ( .IN1(g1718), .IN2(g1734), .QN(n11090) );
  NAND2X0 U11043 ( .IN1(g5738), .IN2(g1732), .QN(n11089) );
  NAND2X0 U11044 ( .IN1(n11092), .IN2(n11093), .QN(n11088) );
  NAND2X0 U11045 ( .IN1(n11037), .IN2(n11062), .QN(n11093) );
  NOR2X0 U11046 ( .IN1(n11060), .IN2(n11042), .QN(n11037) );
  NAND2X0 U11047 ( .IN1(n11033), .IN2(n11094), .QN(n11092) );
  NAND3X0 U11048 ( .IN1(n11095), .IN2(n11096), .IN3(n11097), .QN(n11094) );
  NAND2X0 U11049 ( .IN1(n11084), .IN2(n11060), .QN(n11097) );
  INVX0 U11050 ( .INP(n11046), .ZN(n11060) );
  NAND3X0 U11051 ( .IN1(n11098), .IN2(n11099), .IN3(n11100), .QN(n11046) );
  NAND2X0 U11052 ( .IN1(test_so63), .IN2(g1760), .QN(n11100) );
  NAND2X0 U11053 ( .IN1(g1718), .IN2(g1764), .QN(n11099) );
  NAND2X0 U11054 ( .IN1(g5738), .IN2(g1762), .QN(n11098) );
  NAND2X0 U11055 ( .IN1(n11058), .IN2(n11082), .QN(n11096) );
  INVX0 U11056 ( .INP(n11069), .ZN(n11082) );
  NAND2X0 U11057 ( .IN1(n11064), .IN2(n11059), .QN(n11069) );
  NAND3X0 U11058 ( .IN1(n11101), .IN2(n11102), .IN3(n11103), .QN(n11064) );
  NAND2X0 U11059 ( .IN1(test_so63), .IN2(g1775), .QN(n11103) );
  NAND2X0 U11060 ( .IN1(g1718), .IN2(g1705), .QN(n11102) );
  NAND2X0 U11061 ( .IN1(g5738), .IN2(g1777), .QN(n11101) );
  NAND2X0 U11062 ( .IN1(n11042), .IN2(n11083), .QN(n11095) );
  INVX0 U11063 ( .INP(n11059), .ZN(n11042) );
  NAND3X0 U11064 ( .IN1(n11104), .IN2(n11105), .IN3(n11106), .QN(n11059) );
  NAND2X0 U11065 ( .IN1(test_so63), .IN2(g1745), .QN(n11106) );
  NAND2X0 U11066 ( .IN1(g1718), .IN2(g1749), .QN(n11105) );
  NAND2X0 U11067 ( .IN1(g5738), .IN2(g1747), .QN(n11104) );
  INVX0 U11068 ( .INP(n11107), .ZN(n11070) );
  NAND2X0 U11069 ( .IN1(n11012), .IN2(n11107), .QN(n11008) );
  NAND2X0 U11070 ( .IN1(n4296), .IN2(g1985), .QN(n11023) );
  NAND2X0 U11071 ( .IN1(n11108), .IN2(n11109), .QN(g28351) );
  NAND2X0 U11072 ( .IN1(n4371), .IN2(g1300), .QN(n11109) );
  NAND2X0 U11073 ( .IN1(n10917), .IN2(n11110), .QN(n11108) );
  NAND2X0 U11074 ( .IN1(n11111), .IN2(n11112), .QN(n10917) );
  NAND2X0 U11075 ( .IN1(n9117), .IN2(n10907), .QN(n11112) );
  NAND4X0 U11076 ( .IN1(n11113), .IN2(n11114), .IN3(n11115), .IN4(n10906), 
        .QN(n11111) );
  NAND2X0 U11077 ( .IN1(n11116), .IN2(n11117), .QN(n11113) );
  INVX0 U11078 ( .INP(n11118), .ZN(n11116) );
  NAND2X0 U11079 ( .IN1(n11119), .IN2(n11120), .QN(g28350) );
  NAND2X0 U11080 ( .IN1(n4316), .IN2(g1294), .QN(n11120) );
  NAND2X0 U11081 ( .IN1(n11019), .IN2(g6944), .QN(n11119) );
  NAND2X0 U11082 ( .IN1(n11121), .IN2(n11122), .QN(g28349) );
  NAND2X0 U11083 ( .IN1(n4372), .IN2(g617), .QN(n11122) );
  NAND2X0 U11084 ( .IN1(n11022), .IN2(g6642), .QN(n11121) );
  NAND2X0 U11085 ( .IN1(n11123), .IN2(n11124), .QN(g28348) );
  NAND2X0 U11086 ( .IN1(n4313), .IN2(g611), .QN(n11124) );
  NAND2X0 U11087 ( .IN1(n11125), .IN2(g550), .QN(n11123) );
  NAND2X0 U11088 ( .IN1(n11126), .IN2(n11127), .QN(g28346) );
  NAND2X0 U11089 ( .IN1(g6750), .IN2(n11019), .QN(n11127) );
  NAND2X0 U11090 ( .IN1(n11128), .IN2(n11129), .QN(n11019) );
  NAND2X0 U11091 ( .IN1(n9106), .IN2(n10907), .QN(n11129) );
  NAND4X0 U11092 ( .IN1(n11114), .IN2(n11130), .IN3(n11117), .IN4(n10906), 
        .QN(n11128) );
  INVX0 U11093 ( .INP(n11131), .ZN(n11117) );
  NAND4X0 U11094 ( .IN1(n11132), .IN2(n11133), .IN3(n11134), .IN4(n11135), 
        .QN(n11131) );
  NAND2X0 U11095 ( .IN1(n11136), .IN2(n11137), .QN(n11135) );
  NAND2X0 U11096 ( .IN1(n11138), .IN2(n11139), .QN(n11137) );
  NAND2X0 U11097 ( .IN1(n11140), .IN2(n11141), .QN(n11139) );
  INVX0 U11098 ( .INP(n11142), .ZN(n11141) );
  NAND2X0 U11099 ( .IN1(n11143), .IN2(n11144), .QN(n11138) );
  NAND3X0 U11100 ( .IN1(n11145), .IN2(n11146), .IN3(n11147), .QN(n11134) );
  NAND2X0 U11101 ( .IN1(n11142), .IN2(n11148), .QN(n11146) );
  NAND2X0 U11102 ( .IN1(n11144), .IN2(n11149), .QN(n11148) );
  NAND2X0 U11103 ( .IN1(n11150), .IN2(n11151), .QN(n11144) );
  NAND2X0 U11104 ( .IN1(n11152), .IN2(n11153), .QN(n11151) );
  NOR2X0 U11105 ( .IN1(n11154), .IN2(n11155), .QN(n11142) );
  NOR2X0 U11106 ( .IN1(n11156), .IN2(n11153), .QN(n11155) );
  NOR2X0 U11107 ( .IN1(n11150), .IN2(n11157), .QN(n11154) );
  NAND2X0 U11108 ( .IN1(n11157), .IN2(n11158), .QN(n11133) );
  NAND2X0 U11109 ( .IN1(n11159), .IN2(n11160), .QN(n11158) );
  NAND3X0 U11110 ( .IN1(n11161), .IN2(n11162), .IN3(n11163), .QN(n11160) );
  NAND2X0 U11111 ( .IN1(n11164), .IN2(n11165), .QN(n11159) );
  NAND2X0 U11112 ( .IN1(n11149), .IN2(n11166), .QN(n11164) );
  NAND2X0 U11113 ( .IN1(n11167), .IN2(n11147), .QN(n11166) );
  NAND3X0 U11114 ( .IN1(n11168), .IN2(n11156), .IN3(n11153), .QN(n11132) );
  NAND2X0 U11115 ( .IN1(n11169), .IN2(n11170), .QN(n11168) );
  NAND2X0 U11116 ( .IN1(n11150), .IN2(n11171), .QN(n11170) );
  NAND2X0 U11117 ( .IN1(n11149), .IN2(n11172), .QN(n11171) );
  NAND2X0 U11118 ( .IN1(n11163), .IN2(n11162), .QN(n11169) );
  NAND2X0 U11119 ( .IN1(n11173), .IN2(n11115), .QN(n11130) );
  INVX0 U11120 ( .INP(n11174), .ZN(n11115) );
  NAND3X0 U11121 ( .IN1(n11175), .IN2(n11176), .IN3(n11177), .QN(n11174) );
  NAND2X0 U11122 ( .IN1(n11178), .IN2(n11147), .QN(n11177) );
  NAND2X0 U11123 ( .IN1(n11179), .IN2(n11180), .QN(n11178) );
  NAND2X0 U11124 ( .IN1(n11143), .IN2(n11161), .QN(n11180) );
  INVX0 U11125 ( .INP(n11167), .ZN(n11143) );
  NAND2X0 U11126 ( .IN1(n11157), .IN2(n11181), .QN(n11179) );
  NAND3X0 U11127 ( .IN1(n11182), .IN2(n11183), .IN3(n11184), .QN(n11181) );
  NAND2X0 U11128 ( .IN1(n11163), .IN2(n11156), .QN(n11184) );
  NAND2X0 U11129 ( .IN1(n11185), .IN2(n11186), .QN(n11183) );
  NAND2X0 U11130 ( .IN1(n11187), .IN2(n11140), .QN(n11182) );
  NAND3X0 U11131 ( .IN1(n11188), .IN2(n11156), .IN3(n11145), .QN(n11176) );
  NAND2X0 U11132 ( .IN1(n11189), .IN2(n11190), .QN(n11188) );
  NAND2X0 U11133 ( .IN1(n11136), .IN2(n11149), .QN(n11190) );
  NAND2X0 U11134 ( .IN1(n11157), .IN2(n11150), .QN(n11189) );
  INVX0 U11135 ( .INP(n11153), .ZN(n11157) );
  NAND2X0 U11136 ( .IN1(n11191), .IN2(n11153), .QN(n11175) );
  NAND3X0 U11137 ( .IN1(n11192), .IN2(n11193), .IN3(n11194), .QN(n11153) );
  NAND2X0 U11138 ( .IN1(g5686), .IN2(g1038), .QN(n11194) );
  NAND2X0 U11139 ( .IN1(g5657), .IN2(g1036), .QN(n11193) );
  NAND2X0 U11140 ( .IN1(g1024), .IN2(g1040), .QN(n11192) );
  NAND2X0 U11141 ( .IN1(n11195), .IN2(n11196), .QN(n11191) );
  NAND2X0 U11142 ( .IN1(n11140), .IN2(n11165), .QN(n11196) );
  NOR2X0 U11143 ( .IN1(n11163), .IN2(n11145), .QN(n11140) );
  NAND2X0 U11144 ( .IN1(n11136), .IN2(n11197), .QN(n11195) );
  NAND3X0 U11145 ( .IN1(n11198), .IN2(n11199), .IN3(n11200), .QN(n11197) );
  NAND2X0 U11146 ( .IN1(n11187), .IN2(n11163), .QN(n11200) );
  INVX0 U11147 ( .INP(n11149), .ZN(n11163) );
  NAND3X0 U11148 ( .IN1(n11201), .IN2(n11202), .IN3(n11203), .QN(n11149) );
  NAND2X0 U11149 ( .IN1(g5686), .IN2(g1068), .QN(n11203) );
  NAND2X0 U11150 ( .IN1(g5657), .IN2(g1066), .QN(n11202) );
  NAND2X0 U11151 ( .IN1(g1024), .IN2(g1070), .QN(n11201) );
  NAND2X0 U11152 ( .IN1(n11161), .IN2(n11185), .QN(n11199) );
  INVX0 U11153 ( .INP(n11172), .ZN(n11185) );
  NAND2X0 U11154 ( .IN1(n11167), .IN2(n11162), .QN(n11172) );
  NAND3X0 U11155 ( .IN1(n11204), .IN2(n11205), .IN3(n11206), .QN(n11167) );
  NAND2X0 U11156 ( .IN1(g5686), .IN2(g1083), .QN(n11206) );
  NAND2X0 U11157 ( .IN1(g5657), .IN2(g1081), .QN(n11205) );
  NAND2X0 U11158 ( .IN1(g1024), .IN2(g1011), .QN(n11204) );
  NAND2X0 U11159 ( .IN1(n11145), .IN2(n11186), .QN(n11198) );
  INVX0 U11160 ( .INP(n11162), .ZN(n11145) );
  NAND3X0 U11161 ( .IN1(n11207), .IN2(n11208), .IN3(n11209), .QN(n11162) );
  NAND2X0 U11162 ( .IN1(g5686), .IN2(g1053), .QN(n11209) );
  NAND2X0 U11163 ( .IN1(g5657), .IN2(g1051), .QN(n11208) );
  NAND2X0 U11164 ( .IN1(g1024), .IN2(g1055), .QN(n11207) );
  INVX0 U11165 ( .INP(n11210), .ZN(n11173) );
  NAND2X0 U11166 ( .IN1(n11118), .IN2(n11210), .QN(n11114) );
  NAND2X0 U11167 ( .IN1(n4371), .IN2(g1291), .QN(n11126) );
  NAND2X0 U11168 ( .IN1(n11211), .IN2(n11212), .QN(g28345) );
  NAND2X0 U11169 ( .IN1(n4298), .IN2(g614), .QN(n11212) );
  NAND2X0 U11170 ( .IN1(n11022), .IN2(n11213), .QN(n11211) );
  NAND2X0 U11171 ( .IN1(n11214), .IN2(n11215), .QN(n11022) );
  NAND2X0 U11172 ( .IN1(n8764), .IN2(n10907), .QN(n11215) );
  NAND4X0 U11173 ( .IN1(n11216), .IN2(n11217), .IN3(n11218), .IN4(n10906), 
        .QN(n11214) );
  NAND2X0 U11174 ( .IN1(n11219), .IN2(n11220), .QN(n11216) );
  INVX0 U11175 ( .INP(n11221), .ZN(n11219) );
  NAND2X0 U11176 ( .IN1(n11222), .IN2(n11223), .QN(g28344) );
  NAND2X0 U11177 ( .IN1(n4372), .IN2(g608), .QN(n11223) );
  NAND2X0 U11178 ( .IN1(n11125), .IN2(g6642), .QN(n11222) );
  NAND2X0 U11179 ( .IN1(n11224), .IN2(n11225), .QN(g28342) );
  NAND2X0 U11180 ( .IN1(g6485), .IN2(n11125), .QN(n11225) );
  NAND2X0 U11181 ( .IN1(n11226), .IN2(n11227), .QN(n11125) );
  NAND2X0 U11182 ( .IN1(n8758), .IN2(n10907), .QN(n11227) );
  NAND4X0 U11183 ( .IN1(n11217), .IN2(n11228), .IN3(n11220), .IN4(n10906), 
        .QN(n11226) );
  INVX0 U11184 ( .INP(n11229), .ZN(n11220) );
  NAND4X0 U11185 ( .IN1(n11230), .IN2(n11231), .IN3(n11232), .IN4(n11233), 
        .QN(n11229) );
  NAND2X0 U11186 ( .IN1(n11234), .IN2(n11235), .QN(n11233) );
  NAND2X0 U11187 ( .IN1(n11236), .IN2(n11237), .QN(n11235) );
  NAND2X0 U11188 ( .IN1(n11238), .IN2(n11239), .QN(n11237) );
  INVX0 U11189 ( .INP(n11240), .ZN(n11239) );
  NAND2X0 U11190 ( .IN1(n11241), .IN2(n11242), .QN(n11236) );
  NAND3X0 U11191 ( .IN1(n11243), .IN2(n11244), .IN3(n11245), .QN(n11232) );
  NAND2X0 U11192 ( .IN1(n11240), .IN2(n11246), .QN(n11244) );
  NAND2X0 U11193 ( .IN1(n11242), .IN2(n11247), .QN(n11246) );
  NAND2X0 U11194 ( .IN1(n11248), .IN2(n11249), .QN(n11242) );
  NAND2X0 U11195 ( .IN1(n11250), .IN2(n11251), .QN(n11249) );
  NOR2X0 U11196 ( .IN1(n11252), .IN2(n11253), .QN(n11240) );
  NOR2X0 U11197 ( .IN1(n11254), .IN2(n11251), .QN(n11253) );
  NOR2X0 U11198 ( .IN1(n11248), .IN2(n11255), .QN(n11252) );
  NAND2X0 U11199 ( .IN1(n11255), .IN2(n11256), .QN(n11231) );
  NAND2X0 U11200 ( .IN1(n11257), .IN2(n11258), .QN(n11256) );
  NAND3X0 U11201 ( .IN1(n11259), .IN2(n11260), .IN3(n11261), .QN(n11258) );
  NAND2X0 U11202 ( .IN1(n11262), .IN2(n11263), .QN(n11257) );
  NAND2X0 U11203 ( .IN1(n11247), .IN2(n11264), .QN(n11262) );
  NAND2X0 U11204 ( .IN1(n11265), .IN2(n11245), .QN(n11264) );
  NAND3X0 U11205 ( .IN1(n11266), .IN2(n11254), .IN3(n11251), .QN(n11230) );
  NAND2X0 U11206 ( .IN1(n11267), .IN2(n11268), .QN(n11266) );
  NAND2X0 U11207 ( .IN1(n11248), .IN2(n11269), .QN(n11268) );
  NAND2X0 U11208 ( .IN1(n11247), .IN2(n11270), .QN(n11269) );
  NAND2X0 U11209 ( .IN1(n11261), .IN2(n11260), .QN(n11267) );
  NAND2X0 U11210 ( .IN1(n11271), .IN2(n11218), .QN(n11228) );
  INVX0 U11211 ( .INP(n11272), .ZN(n11218) );
  NAND3X0 U11212 ( .IN1(n11273), .IN2(n11274), .IN3(n11275), .QN(n11272) );
  NAND2X0 U11213 ( .IN1(n11276), .IN2(n11245), .QN(n11275) );
  NAND2X0 U11214 ( .IN1(n11277), .IN2(n11278), .QN(n11276) );
  NAND2X0 U11215 ( .IN1(n11241), .IN2(n11259), .QN(n11278) );
  INVX0 U11216 ( .INP(n11265), .ZN(n11241) );
  NAND2X0 U11217 ( .IN1(n11255), .IN2(n11279), .QN(n11277) );
  NAND3X0 U11218 ( .IN1(n11280), .IN2(n11281), .IN3(n11282), .QN(n11279) );
  NAND2X0 U11219 ( .IN1(n11261), .IN2(n11254), .QN(n11282) );
  NAND2X0 U11220 ( .IN1(n11283), .IN2(n11284), .QN(n11281) );
  NAND2X0 U11221 ( .IN1(n11285), .IN2(n11238), .QN(n11280) );
  NAND3X0 U11222 ( .IN1(n11286), .IN2(n11254), .IN3(n11243), .QN(n11274) );
  NAND2X0 U11223 ( .IN1(n11287), .IN2(n11288), .QN(n11286) );
  NAND2X0 U11224 ( .IN1(n11234), .IN2(n11247), .QN(n11288) );
  NAND2X0 U11225 ( .IN1(n11255), .IN2(n11248), .QN(n11287) );
  INVX0 U11226 ( .INP(n11251), .ZN(n11255) );
  NAND2X0 U11227 ( .IN1(n11289), .IN2(n11251), .QN(n11273) );
  NAND3X0 U11228 ( .IN1(n11290), .IN2(n11291), .IN3(n11292), .QN(n11251) );
  NAND2X0 U11229 ( .IN1(g5648), .IN2(g351), .QN(n11292) );
  NAND2X0 U11230 ( .IN1(g5629), .IN2(g349), .QN(n11291) );
  NAND2X0 U11231 ( .IN1(g337), .IN2(g353), .QN(n11290) );
  NAND2X0 U11232 ( .IN1(n11293), .IN2(n11294), .QN(n11289) );
  NAND2X0 U11233 ( .IN1(n11238), .IN2(n11263), .QN(n11294) );
  NOR2X0 U11234 ( .IN1(n11261), .IN2(n11243), .QN(n11238) );
  NAND2X0 U11235 ( .IN1(n11234), .IN2(n11295), .QN(n11293) );
  NAND3X0 U11236 ( .IN1(n11296), .IN2(n11297), .IN3(n11298), .QN(n11295) );
  NAND2X0 U11237 ( .IN1(n11285), .IN2(n11261), .QN(n11298) );
  INVX0 U11238 ( .INP(n11247), .ZN(n11261) );
  NAND3X0 U11239 ( .IN1(n11299), .IN2(n11300), .IN3(n11301), .QN(n11247) );
  NAND2X0 U11240 ( .IN1(g5648), .IN2(g381), .QN(n11301) );
  NAND2X0 U11241 ( .IN1(g5629), .IN2(g379), .QN(n11300) );
  NAND2X0 U11242 ( .IN1(g337), .IN2(g383), .QN(n11299) );
  NAND2X0 U11243 ( .IN1(n11259), .IN2(n11283), .QN(n11297) );
  INVX0 U11244 ( .INP(n11270), .ZN(n11283) );
  NAND2X0 U11245 ( .IN1(n11265), .IN2(n11260), .QN(n11270) );
  NAND3X0 U11246 ( .IN1(n11302), .IN2(n11303), .IN3(n11304), .QN(n11265) );
  NAND2X0 U11247 ( .IN1(g5648), .IN2(g396), .QN(n11304) );
  NAND2X0 U11248 ( .IN1(g5629), .IN2(g394), .QN(n11303) );
  NAND2X0 U11249 ( .IN1(g337), .IN2(g324), .QN(n11302) );
  NAND2X0 U11250 ( .IN1(n11243), .IN2(n11284), .QN(n11296) );
  INVX0 U11251 ( .INP(n11260), .ZN(n11243) );
  NAND3X0 U11252 ( .IN1(n11305), .IN2(n11306), .IN3(n11307), .QN(n11260) );
  NAND2X0 U11253 ( .IN1(g5648), .IN2(g366), .QN(n11307) );
  NAND2X0 U11254 ( .IN1(g5629), .IN2(g364), .QN(n11306) );
  NAND2X0 U11255 ( .IN1(g337), .IN2(g368), .QN(n11305) );
  INVX0 U11256 ( .INP(n11308), .ZN(n11271) );
  NAND2X0 U11257 ( .IN1(n11221), .IN2(n11308), .QN(n11217) );
  NAND2X0 U11258 ( .IN1(n4298), .IN2(g605), .QN(n11224) );
  NOR2X0 U11259 ( .IN1(n11309), .IN2(n11310), .QN(g28328) );
  XNOR2X1 U11260 ( .IN1(n4415), .IN2(n11311), .Q(n11310) );
  NAND2X0 U11261 ( .IN1(n11312), .IN2(g2760), .QN(n11311) );
  NOR2X0 U11262 ( .IN1(n9323), .IN2(n11313), .QN(g28325) );
  XNOR2X1 U11263 ( .IN1(n4416), .IN2(n11314), .Q(n11313) );
  NAND2X0 U11264 ( .IN1(test_so70), .IN2(n11315), .QN(n11314) );
  NOR2X0 U11265 ( .IN1(n8524), .IN2(n11316), .QN(g28321) );
  XNOR2X1 U11266 ( .IN1(n4417), .IN2(n11317), .Q(n11316) );
  NAND2X0 U11267 ( .IN1(n11318), .IN2(g1372), .QN(n11317) );
  NOR2X0 U11268 ( .IN1(n8548), .IN2(n11319), .QN(g28199) );
  XOR2X1 U11269 ( .IN1(n4396), .IN2(n10874), .Q(n11319) );
  NOR2X0 U11270 ( .IN1(n10283), .IN2(n11320), .QN(g28148) );
  XOR2X1 U11271 ( .IN1(n8095), .IN2(n3424), .Q(n11320) );
  NOR2X0 U11272 ( .IN1(n10285), .IN2(n11321), .QN(g28147) );
  XOR2X1 U11273 ( .IN1(n8094), .IN2(n3427), .Q(n11321) );
  NOR2X0 U11274 ( .IN1(n10287), .IN2(n11322), .QN(g28146) );
  XOR2X1 U11275 ( .IN1(n8092), .IN2(n3430), .Q(n11322) );
  NOR2X0 U11276 ( .IN1(n10289), .IN2(n11323), .QN(g28145) );
  XOR2X1 U11277 ( .IN1(n8093), .IN2(n3433), .Q(n11323) );
  NAND2X0 U11278 ( .IN1(n11324), .IN2(n11325), .QN(g27771) );
  NAND2X0 U11279 ( .IN1(test_so81), .IN2(n11326), .QN(n11325) );
  NAND2X0 U11280 ( .IN1(n11327), .IN2(n10047), .QN(n11326) );
  NAND2X0 U11281 ( .IN1(n11328), .IN2(n10047), .QN(n11324) );
  NAND2X0 U11282 ( .IN1(n11329), .IN2(n11330), .QN(g27769) );
  NAND2X0 U11283 ( .IN1(n11331), .IN2(g2524), .QN(n11330) );
  NAND2X0 U11284 ( .IN1(n11327), .IN2(n10046), .QN(n11331) );
  NAND2X0 U11285 ( .IN1(n11328), .IN2(n10046), .QN(n11329) );
  NAND2X0 U11286 ( .IN1(n11332), .IN2(n11333), .QN(g27768) );
  NAND2X0 U11287 ( .IN1(n11334), .IN2(g1828), .QN(n11333) );
  NAND2X0 U11288 ( .IN1(n11335), .IN2(n10093), .QN(n11334) );
  NAND2X0 U11289 ( .IN1(n11336), .IN2(n10093), .QN(n11332) );
  NAND2X0 U11290 ( .IN1(n11337), .IN2(n11338), .QN(g27767) );
  NAND2X0 U11291 ( .IN1(n11339), .IN2(g2523), .QN(n11338) );
  NAND2X0 U11292 ( .IN1(n11327), .IN2(n10048), .QN(n11339) );
  NOR2X0 U11293 ( .IN1(n11340), .IN2(n11341), .QN(n11327) );
  NAND2X0 U11294 ( .IN1(n11328), .IN2(n10048), .QN(n11337) );
  INVX0 U11295 ( .INP(n11342), .ZN(n11328) );
  NAND4X0 U11296 ( .IN1(test_so79), .IN2(n11343), .IN3(n11344), .IN4(n11345), 
        .QN(n11342) );
  NAND2X0 U11297 ( .IN1(n11346), .IN2(n11347), .QN(n11345) );
  NAND2X0 U11298 ( .IN1(n11348), .IN2(n11349), .QN(n11344) );
  NAND2X0 U11299 ( .IN1(n11350), .IN2(n11351), .QN(n11343) );
  NAND2X0 U11300 ( .IN1(n11352), .IN2(n11353), .QN(g27766) );
  NAND2X0 U11301 ( .IN1(n11354), .IN2(g1830), .QN(n11353) );
  NAND2X0 U11302 ( .IN1(n11335), .IN2(n10092), .QN(n11354) );
  NAND2X0 U11303 ( .IN1(n11336), .IN2(n10092), .QN(n11352) );
  NAND2X0 U11304 ( .IN1(n11355), .IN2(n11356), .QN(g27765) );
  NAND2X0 U11305 ( .IN1(n11357), .IN2(g1134), .QN(n11356) );
  NAND2X0 U11306 ( .IN1(n11358), .IN2(g1088), .QN(n11357) );
  NAND2X0 U11307 ( .IN1(n11359), .IN2(g1088), .QN(n11355) );
  NAND2X0 U11308 ( .IN1(n11360), .IN2(n11361), .QN(g27764) );
  NAND2X0 U11309 ( .IN1(n11362), .IN2(g1829), .QN(n11361) );
  NAND2X0 U11310 ( .IN1(n11335), .IN2(n10094), .QN(n11362) );
  NOR2X0 U11311 ( .IN1(n11363), .IN2(n11364), .QN(n11335) );
  NAND2X0 U11312 ( .IN1(n11336), .IN2(n10094), .QN(n11360) );
  INVX0 U11313 ( .INP(n11365), .ZN(n11336) );
  NAND4X0 U11314 ( .IN1(n11366), .IN2(g1690), .IN3(n11367), .IN4(n11368), .QN(
        n11365) );
  NAND2X0 U11315 ( .IN1(n11369), .IN2(n11370), .QN(n11368) );
  NAND2X0 U11316 ( .IN1(n11371), .IN2(n11372), .QN(n11367) );
  NAND2X0 U11317 ( .IN1(n11373), .IN2(n11374), .QN(n11366) );
  NAND2X0 U11318 ( .IN1(n11375), .IN2(n11376), .QN(g27763) );
  NAND2X0 U11319 ( .IN1(n11377), .IN2(g1136), .QN(n11376) );
  NAND2X0 U11320 ( .IN1(n11358), .IN2(g6712), .QN(n11377) );
  NAND2X0 U11321 ( .IN1(n11359), .IN2(g6712), .QN(n11375) );
  NAND2X0 U11322 ( .IN1(n11378), .IN2(n11379), .QN(g27762) );
  NAND2X0 U11323 ( .IN1(n11380), .IN2(g447), .QN(n11379) );
  NAND2X0 U11324 ( .IN1(n11381), .IN2(n10178), .QN(n11380) );
  NAND2X0 U11325 ( .IN1(n11382), .IN2(n10178), .QN(n11378) );
  NAND2X0 U11326 ( .IN1(n11383), .IN2(n11384), .QN(g27761) );
  NAND2X0 U11327 ( .IN1(n11385), .IN2(g1135), .QN(n11384) );
  NAND2X0 U11328 ( .IN1(n11358), .IN2(g5472), .QN(n11385) );
  NOR2X0 U11329 ( .IN1(n11386), .IN2(n11387), .QN(n11358) );
  NAND2X0 U11330 ( .IN1(n11359), .IN2(g5472), .QN(n11383) );
  INVX0 U11331 ( .INP(n11388), .ZN(n11359) );
  NAND4X0 U11332 ( .IN1(n11389), .IN2(g996), .IN3(n11390), .IN4(n11391), .QN(
        n11388) );
  NAND2X0 U11333 ( .IN1(n11392), .IN2(n11393), .QN(n11391) );
  NAND2X0 U11334 ( .IN1(n11394), .IN2(n11395), .QN(n11390) );
  NAND2X0 U11335 ( .IN1(n11396), .IN2(n11397), .QN(n11389) );
  NAND2X0 U11336 ( .IN1(n11398), .IN2(n11399), .QN(g27760) );
  NAND2X0 U11337 ( .IN1(n11400), .IN2(g449), .QN(n11399) );
  NAND2X0 U11338 ( .IN1(n11381), .IN2(n10177), .QN(n11400) );
  NAND2X0 U11339 ( .IN1(n11382), .IN2(n10177), .QN(n11398) );
  NAND2X0 U11340 ( .IN1(n11401), .IN2(n11402), .QN(g27759) );
  NAND2X0 U11341 ( .IN1(n11403), .IN2(g448), .QN(n11402) );
  NAND2X0 U11342 ( .IN1(n11381), .IN2(n10176), .QN(n11403) );
  NOR2X0 U11343 ( .IN1(n11404), .IN2(n11405), .QN(n11381) );
  NAND2X0 U11344 ( .IN1(n11382), .IN2(n10176), .QN(n11401) );
  INVX0 U11345 ( .INP(n11406), .ZN(n11382) );
  NAND4X0 U11346 ( .IN1(n11407), .IN2(g309), .IN3(n11408), .IN4(n11409), .QN(
        n11406) );
  NAND2X0 U11347 ( .IN1(n11410), .IN2(n11411), .QN(n11409) );
  NAND2X0 U11348 ( .IN1(n11412), .IN2(n11413), .QN(n11408) );
  NAND2X0 U11349 ( .IN1(n11414), .IN2(n11415), .QN(n11407) );
  NOR2X0 U11350 ( .IN1(n11309), .IN2(n11416), .QN(g27724) );
  XOR2X1 U11351 ( .IN1(n4393), .IN2(n11312), .Q(n11416) );
  NOR2X0 U11352 ( .IN1(n9323), .IN2(n11417), .QN(g27722) );
  XOR2X1 U11353 ( .IN1(n8106), .IN2(n11315), .Q(n11417) );
  NOR2X0 U11354 ( .IN1(n8524), .IN2(n11418), .QN(g27718) );
  XOR2X1 U11355 ( .IN1(n4395), .IN2(n11318), .Q(n11418) );
  NOR3X0 U11356 ( .IN1(n11419), .IN2(n9323), .IN3(n11315), .QN(g27682) );
  NOR3X0 U11357 ( .IN1(n4468), .IN2(n4473), .IN3(n11420), .QN(n11315) );
  NOR2X0 U11358 ( .IN1(n11421), .IN2(g2059), .QN(n11419) );
  NOR2X0 U11359 ( .IN1(n4468), .IN2(n11420), .QN(n11421) );
  INVX0 U11360 ( .INP(n9324), .ZN(n11420) );
  NOR3X0 U11361 ( .IN1(n11422), .IN2(n8524), .IN3(n11318), .QN(g27678) );
  NOR3X0 U11362 ( .IN1(n4469), .IN2(n4475), .IN3(n8520), .QN(n11318) );
  NOR2X0 U11363 ( .IN1(n11423), .IN2(g1365), .QN(n11422) );
  NOR2X0 U11364 ( .IN1(n4469), .IN2(n8520), .QN(n11423) );
  NOR3X0 U11365 ( .IN1(n11424), .IN2(n8548), .IN3(n10874), .QN(g27672) );
  NOR3X0 U11366 ( .IN1(n8540), .IN2(n4477), .IN3(n8105), .QN(n10874) );
  NOR2X0 U11367 ( .IN1(n11425), .IN2(g679), .QN(n11424) );
  NOR2X0 U11368 ( .IN1(n8540), .IN2(n8105), .QN(n11425) );
  NOR2X0 U11369 ( .IN1(n10283), .IN2(n11426), .QN(g27621) );
  XOR2X1 U11370 ( .IN1(n11427), .IN2(n7700), .Q(n11426) );
  NOR2X0 U11371 ( .IN1(n10285), .IN2(n11428), .QN(g27612) );
  XOR2X1 U11372 ( .IN1(n11429), .IN2(n7704), .Q(n11428) );
  NOR2X0 U11373 ( .IN1(n10287), .IN2(n11430), .QN(g27603) );
  XNOR2X1 U11374 ( .IN1(n7708), .IN2(n3431), .Q(n11430) );
  NAND2X0 U11375 ( .IN1(n3689), .IN2(g767), .QN(n3431) );
  NOR2X0 U11376 ( .IN1(n10289), .IN2(n11431), .QN(g27594) );
  XOR2X1 U11377 ( .IN1(n11432), .IN2(n7712), .Q(n11431) );
  NAND4X0 U11378 ( .IN1(n11433), .IN2(n11434), .IN3(n3700), .IN4(n11435), .QN(
        g27380) );
  NOR4X0 U11379 ( .IN1(n11436), .IN2(n11437), .IN3(n11438), .IN4(n11439), .QN(
        n11435) );
  NOR2X0 U11380 ( .IN1(n4424), .IN2(n11440), .QN(n11439) );
  NOR2X0 U11381 ( .IN1(n11441), .IN2(n11442), .QN(n11438) );
  NOR2X0 U11382 ( .IN1(n11443), .IN2(n3705), .QN(n11441) );
  NOR3X0 U11383 ( .IN1(g185), .IN2(n4405), .IN3(n11444), .QN(n11443) );
  NOR4X0 U11384 ( .IN1(n11445), .IN2(n11446), .IN3(n11444), .IN4(n11447), .QN(
        n11437) );
  NOR2X0 U11385 ( .IN1(n14384), .IN2(n11448), .QN(n11446) );
  NOR2X0 U11386 ( .IN1(n14382), .IN2(n11449), .QN(n11445) );
  INVX0 U11387 ( .INP(n11450), .ZN(n11434) );
  NOR2X0 U11388 ( .IN1(n11451), .IN2(n14385), .QN(n11450) );
  NAND2X0 U11389 ( .IN1(n7442), .IN2(n11452), .QN(n11433) );
  NAND2X0 U11390 ( .IN1(n11453), .IN2(n11454), .QN(g27354) );
  INVX0 U11391 ( .INP(n11455), .ZN(n11454) );
  NOR2X0 U11392 ( .IN1(n11456), .IN2(n7362), .QN(n11455) );
  NAND2X0 U11393 ( .IN1(n11456), .IN2(n11457), .QN(n11453) );
  NAND2X0 U11394 ( .IN1(n11458), .IN2(n11459), .QN(g27348) );
  NAND2X0 U11395 ( .IN1(n11460), .IN2(g2660), .QN(n11459) );
  NAND2X0 U11396 ( .IN1(n11461), .IN2(n11457), .QN(n11458) );
  NAND2X0 U11397 ( .IN1(n11462), .IN2(n11463), .QN(g27347) );
  INVX0 U11398 ( .INP(n11464), .ZN(n11463) );
  NOR2X0 U11399 ( .IN1(n11456), .IN2(n7178), .QN(n11464) );
  NAND2X0 U11400 ( .IN1(n11456), .IN2(n11465), .QN(n11462) );
  NAND2X0 U11401 ( .IN1(n11466), .IN2(n11467), .QN(g27346) );
  INVX0 U11402 ( .INP(n11468), .ZN(n11467) );
  NOR2X0 U11403 ( .IN1(n11469), .IN2(n7364), .QN(n11468) );
  NAND2X0 U11404 ( .IN1(n11469), .IN2(n11470), .QN(n11466) );
  NAND2X0 U11405 ( .IN1(n11471), .IN2(n11472), .QN(g27345) );
  INVX0 U11406 ( .INP(n11473), .ZN(n11472) );
  NOR2X0 U11407 ( .IN1(n11474), .IN2(n7361), .QN(n11473) );
  NAND2X0 U11408 ( .IN1(n11474), .IN2(n11457), .QN(n11471) );
  NAND3X0 U11409 ( .IN1(n10955), .IN2(n10930), .IN3(n11475), .QN(n11457) );
  INVX0 U11410 ( .INP(n10944), .ZN(n10955) );
  NAND2X0 U11411 ( .IN1(n11476), .IN2(n11477), .QN(g27344) );
  NAND2X0 U11412 ( .IN1(test_so89), .IN2(n11460), .QN(n11477) );
  NAND2X0 U11413 ( .IN1(n11461), .IN2(n11465), .QN(n11476) );
  NAND2X0 U11414 ( .IN1(n11478), .IN2(n11479), .QN(g27343) );
  INVX0 U11415 ( .INP(n11480), .ZN(n11479) );
  NOR2X0 U11416 ( .IN1(n11456), .IN2(n7351), .QN(n11480) );
  NAND2X0 U11417 ( .IN1(n11456), .IN2(n11481), .QN(n11478) );
  NAND2X0 U11418 ( .IN1(n11482), .IN2(n11483), .QN(g27342) );
  INVX0 U11419 ( .INP(n11484), .ZN(n11483) );
  NOR2X0 U11420 ( .IN1(n11485), .IN2(n7644), .QN(n11484) );
  NAND2X0 U11421 ( .IN1(n11485), .IN2(n11486), .QN(n11482) );
  NAND2X0 U11422 ( .IN1(n11487), .IN2(n11488), .QN(g27341) );
  INVX0 U11423 ( .INP(n11489), .ZN(n11488) );
  NOR2X0 U11424 ( .IN1(n11490), .IN2(n7365), .QN(n11489) );
  NAND2X0 U11425 ( .IN1(n11490), .IN2(n11470), .QN(n11487) );
  NAND2X0 U11426 ( .IN1(n11491), .IN2(n11492), .QN(g27340) );
  INVX0 U11427 ( .INP(n11493), .ZN(n11492) );
  NOR2X0 U11428 ( .IN1(n11469), .IN2(n7180), .QN(n11493) );
  NAND2X0 U11429 ( .IN1(n11469), .IN2(n11494), .QN(n11491) );
  NAND2X0 U11430 ( .IN1(n11495), .IN2(n11496), .QN(g27339) );
  NAND2X0 U11431 ( .IN1(n11497), .IN2(g1270), .QN(n11496) );
  NAND2X0 U11432 ( .IN1(n11498), .IN2(n11499), .QN(n11495) );
  NAND2X0 U11433 ( .IN1(n11500), .IN2(n11501), .QN(g27338) );
  INVX0 U11434 ( .INP(n11502), .ZN(n11501) );
  NOR2X0 U11435 ( .IN1(n11474), .IN2(n7177), .QN(n11502) );
  NAND2X0 U11436 ( .IN1(n11474), .IN2(n11465), .QN(n11500) );
  INVX0 U11437 ( .INP(n11503), .ZN(n11465) );
  NAND2X0 U11438 ( .IN1(n11504), .IN2(n11505), .QN(n11503) );
  NAND2X0 U11439 ( .IN1(n11506), .IN2(n10980), .QN(n11505) );
  NAND2X0 U11440 ( .IN1(n11475), .IN2(n10944), .QN(n11504) );
  INVX0 U11441 ( .INP(n11506), .ZN(n11475) );
  NAND2X0 U11442 ( .IN1(n11507), .IN2(n11508), .QN(g27337) );
  NAND2X0 U11443 ( .IN1(n11460), .IN2(g2654), .QN(n11508) );
  NAND2X0 U11444 ( .IN1(n11461), .IN2(n11481), .QN(n11507) );
  NAND2X0 U11445 ( .IN1(n11509), .IN2(n11510), .QN(g27336) );
  INVX0 U11446 ( .INP(n11511), .ZN(n11510) );
  NOR2X0 U11447 ( .IN1(n11456), .IN2(n7339), .QN(n11511) );
  NAND2X0 U11448 ( .IN1(n11456), .IN2(n11512), .QN(n11509) );
  NOR2X0 U11449 ( .IN1(n11513), .IN2(n4299), .QN(n11456) );
  NAND2X0 U11450 ( .IN1(n11514), .IN2(n11515), .QN(g27335) );
  INVX0 U11451 ( .INP(n11516), .ZN(n11515) );
  NOR2X0 U11452 ( .IN1(n11517), .IN2(n7645), .QN(n11516) );
  NAND2X0 U11453 ( .IN1(n11517), .IN2(n11486), .QN(n11514) );
  NAND2X0 U11454 ( .IN1(n11518), .IN2(n11519), .QN(g27334) );
  INVX0 U11455 ( .INP(n11520), .ZN(n11519) );
  NOR2X0 U11456 ( .IN1(n11485), .IN2(n7384), .QN(n11520) );
  NAND2X0 U11457 ( .IN1(n11485), .IN2(n11521), .QN(n11518) );
  NAND2X0 U11458 ( .IN1(n11522), .IN2(n11523), .QN(g27333) );
  NAND2X0 U11459 ( .IN1(n11524), .IN2(n11470), .QN(n11523) );
  NAND2X0 U11460 ( .IN1(n11525), .IN2(n11058), .QN(n11470) );
  NOR2X0 U11461 ( .IN1(n11053), .IN2(n11083), .QN(n11058) );
  INVX0 U11462 ( .INP(n11526), .ZN(n11522) );
  NOR2X0 U11463 ( .IN1(n8109), .IN2(n11524), .QN(n11526) );
  NAND2X0 U11464 ( .IN1(n11527), .IN2(n11528), .QN(g27332) );
  INVX0 U11465 ( .INP(n11529), .ZN(n11528) );
  NOR2X0 U11466 ( .IN1(n11490), .IN2(n7181), .QN(n11529) );
  NAND2X0 U11467 ( .IN1(n11490), .IN2(n11494), .QN(n11527) );
  NAND2X0 U11468 ( .IN1(n11530), .IN2(n11531), .QN(g27331) );
  INVX0 U11469 ( .INP(n11532), .ZN(n11531) );
  NOR2X0 U11470 ( .IN1(n11469), .IN2(n7354), .QN(n11532) );
  NAND2X0 U11471 ( .IN1(n11469), .IN2(n11533), .QN(n11530) );
  NAND2X0 U11472 ( .IN1(n11534), .IN2(n11535), .QN(g27330) );
  INVX0 U11473 ( .INP(n11536), .ZN(n11535) );
  NOR2X0 U11474 ( .IN1(n11537), .IN2(n7647), .QN(n11536) );
  NAND2X0 U11475 ( .IN1(n11537), .IN2(n11538), .QN(n11534) );
  NAND2X0 U11476 ( .IN1(n11539), .IN2(n11540), .QN(g27329) );
  NAND2X0 U11477 ( .IN1(n11541), .IN2(n11499), .QN(n11540) );
  INVX0 U11478 ( .INP(n11542), .ZN(n11539) );
  NOR2X0 U11479 ( .IN1(n11541), .IN2(n7368), .QN(n11542) );
  NAND2X0 U11480 ( .IN1(n11543), .IN2(n11544), .QN(g27328) );
  NAND2X0 U11481 ( .IN1(test_so46), .IN2(n11497), .QN(n11544) );
  NAND2X0 U11482 ( .IN1(n11498), .IN2(n11545), .QN(n11543) );
  NAND2X0 U11483 ( .IN1(n11546), .IN2(n11547), .QN(g27327) );
  INVX0 U11484 ( .INP(n11548), .ZN(n11547) );
  NOR2X0 U11485 ( .IN1(n11549), .IN2(n7370), .QN(n11548) );
  NAND2X0 U11486 ( .IN1(n11549), .IN2(n11550), .QN(n11546) );
  NAND2X0 U11487 ( .IN1(n11551), .IN2(n11552), .QN(g27326) );
  INVX0 U11488 ( .INP(n11553), .ZN(n11552) );
  NOR2X0 U11489 ( .IN1(n11474), .IN2(n7350), .QN(n11553) );
  NAND2X0 U11490 ( .IN1(n11474), .IN2(n11481), .QN(n11551) );
  INVX0 U11491 ( .INP(n11554), .ZN(n11481) );
  NAND2X0 U11492 ( .IN1(n11555), .IN2(n11556), .QN(n11554) );
  NAND2X0 U11493 ( .IN1(n11506), .IN2(n10950), .QN(n11555) );
  XNOR2X1 U11494 ( .IN1(n8798), .IN2(n10934), .Q(n11506) );
  NAND2X0 U11495 ( .IN1(n11557), .IN2(n11558), .QN(g27325) );
  NAND2X0 U11496 ( .IN1(n11460), .IN2(g2651), .QN(n11558) );
  INVX0 U11497 ( .INP(n11461), .ZN(n11460) );
  NAND2X0 U11498 ( .IN1(n11461), .IN2(n11512), .QN(n11557) );
  NOR2X0 U11499 ( .IN1(n11513), .IN2(n4370), .QN(n11461) );
  NAND2X0 U11500 ( .IN1(n11559), .IN2(n11560), .QN(g27324) );
  INVX0 U11501 ( .INP(n11561), .ZN(n11560) );
  NOR2X0 U11502 ( .IN1(n11562), .IN2(n7646), .QN(n11561) );
  NAND2X0 U11503 ( .IN1(n11562), .IN2(n11486), .QN(n11559) );
  NAND3X0 U11504 ( .IN1(n11563), .IN2(n11564), .IN3(n11565), .QN(n11486) );
  NAND2X0 U11505 ( .IN1(n11566), .IN2(n11567), .QN(g27323) );
  INVX0 U11506 ( .INP(n11568), .ZN(n11567) );
  NOR2X0 U11507 ( .IN1(n11517), .IN2(n7385), .QN(n11568) );
  NAND2X0 U11508 ( .IN1(n11517), .IN2(n11521), .QN(n11566) );
  NAND2X0 U11509 ( .IN1(n11569), .IN2(n11570), .QN(g27322) );
  INVX0 U11510 ( .INP(n11571), .ZN(n11570) );
  NOR2X0 U11511 ( .IN1(n11485), .IN2(n7632), .QN(n11571) );
  NAND2X0 U11512 ( .IN1(n11572), .IN2(n11485), .QN(n11569) );
  NAND2X0 U11513 ( .IN1(n11573), .IN2(n11574), .QN(g27321) );
  INVX0 U11514 ( .INP(n11575), .ZN(n11574) );
  NOR2X0 U11515 ( .IN1(n11524), .IN2(n7179), .QN(n11575) );
  NAND2X0 U11516 ( .IN1(n11524), .IN2(n11494), .QN(n11573) );
  INVX0 U11517 ( .INP(n11576), .ZN(n11494) );
  NAND2X0 U11518 ( .IN1(n11577), .IN2(n11578), .QN(n11576) );
  NAND2X0 U11519 ( .IN1(n11579), .IN2(n11084), .QN(n11578) );
  NAND2X0 U11520 ( .IN1(n11525), .IN2(n11053), .QN(n11577) );
  INVX0 U11521 ( .INP(n11579), .ZN(n11525) );
  NAND2X0 U11522 ( .IN1(n11580), .IN2(n11581), .QN(g27320) );
  INVX0 U11523 ( .INP(n11582), .ZN(n11581) );
  NOR2X0 U11524 ( .IN1(n11490), .IN2(n7355), .QN(n11582) );
  NAND2X0 U11525 ( .IN1(n11490), .IN2(n11533), .QN(n11580) );
  NAND2X0 U11526 ( .IN1(n11583), .IN2(n11584), .QN(g27319) );
  INVX0 U11527 ( .INP(n11585), .ZN(n11584) );
  NOR2X0 U11528 ( .IN1(n11469), .IN2(n7342), .QN(n11585) );
  NAND2X0 U11529 ( .IN1(n11469), .IN2(n11586), .QN(n11583) );
  NOR2X0 U11530 ( .IN1(n11587), .IN2(n4366), .QN(n11469) );
  NAND2X0 U11531 ( .IN1(n11588), .IN2(n11589), .QN(g27318) );
  NAND2X0 U11532 ( .IN1(n11590), .IN2(n11538), .QN(n11589) );
  NAND2X0 U11533 ( .IN1(test_so58), .IN2(n11591), .QN(n11588) );
  NAND2X0 U11534 ( .IN1(n11592), .IN2(n11593), .QN(g27317) );
  INVX0 U11535 ( .INP(n11594), .ZN(n11593) );
  NOR2X0 U11536 ( .IN1(n11537), .IN2(n7387), .QN(n11594) );
  NAND2X0 U11537 ( .IN1(n11537), .IN2(n11595), .QN(n11592) );
  NAND2X0 U11538 ( .IN1(n11596), .IN2(n11597), .QN(g27316) );
  NAND2X0 U11539 ( .IN1(n11598), .IN2(n11499), .QN(n11597) );
  NAND2X0 U11540 ( .IN1(n11599), .IN2(n11161), .QN(n11499) );
  NOR2X0 U11541 ( .IN1(n11156), .IN2(n11186), .QN(n11161) );
  NAND2X0 U11542 ( .IN1(n11600), .IN2(g1271), .QN(n11596) );
  NAND2X0 U11543 ( .IN1(n11601), .IN2(n11602), .QN(g27315) );
  INVX0 U11544 ( .INP(n11603), .ZN(n11602) );
  NOR2X0 U11545 ( .IN1(n11541), .IN2(n7183), .QN(n11603) );
  NAND2X0 U11546 ( .IN1(n11541), .IN2(n11545), .QN(n11601) );
  NAND2X0 U11547 ( .IN1(n11604), .IN2(n11605), .QN(g27314) );
  NAND2X0 U11548 ( .IN1(n11497), .IN2(g1264), .QN(n11605) );
  NAND2X0 U11549 ( .IN1(n11498), .IN2(n11606), .QN(n11604) );
  NAND2X0 U11550 ( .IN1(n11607), .IN2(n11608), .QN(g27313) );
  INVX0 U11551 ( .INP(n11609), .ZN(n11608) );
  NOR2X0 U11552 ( .IN1(n11610), .IN2(n7649), .QN(n11609) );
  NAND2X0 U11553 ( .IN1(n11610), .IN2(n11611), .QN(n11607) );
  NAND2X0 U11554 ( .IN1(n11612), .IN2(n11613), .QN(g27312) );
  NAND2X0 U11555 ( .IN1(n11614), .IN2(n11550), .QN(n11613) );
  NAND2X0 U11556 ( .IN1(n11615), .IN2(g586), .QN(n11612) );
  NAND2X0 U11557 ( .IN1(n11616), .IN2(n11617), .QN(g27311) );
  INVX0 U11558 ( .INP(n11618), .ZN(n11617) );
  NOR2X0 U11559 ( .IN1(n11549), .IN2(n7185), .QN(n11618) );
  NAND2X0 U11560 ( .IN1(n11549), .IN2(n11619), .QN(n11616) );
  NAND2X0 U11561 ( .IN1(n11620), .IN2(n11621), .QN(g27310) );
  INVX0 U11562 ( .INP(n11622), .ZN(n11621) );
  NOR2X0 U11563 ( .IN1(n11474), .IN2(n7338), .QN(n11622) );
  NAND2X0 U11564 ( .IN1(n11474), .IN2(n11512), .QN(n11620) );
  NOR2X0 U11565 ( .IN1(n11623), .IN2(n11624), .QN(n11512) );
  NOR2X0 U11566 ( .IN1(n11625), .IN2(g3229), .QN(n11624) );
  INVX0 U11567 ( .INP(n11626), .ZN(n11625) );
  NAND2X0 U11568 ( .IN1(n11556), .IN2(n11627), .QN(n11626) );
  NAND2X0 U11569 ( .IN1(n10932), .IN2(n10937), .QN(n11627) );
  INVX0 U11570 ( .INP(n10964), .ZN(n10932) );
  NAND2X0 U11571 ( .IN1(n10930), .IN2(n10944), .QN(n11556) );
  INVX0 U11572 ( .INP(n10950), .ZN(n10930) );
  NOR2X0 U11573 ( .IN1(n8798), .IN2(n11628), .QN(n11623) );
  NOR2X0 U11574 ( .IN1(n10964), .IN2(n11629), .QN(n11628) );
  NOR2X0 U11575 ( .IN1(n10934), .IN2(n11630), .QN(n11629) );
  NOR2X0 U11576 ( .IN1(n10950), .IN2(n10980), .QN(n11630) );
  NOR2X0 U11577 ( .IN1(n10944), .IN2(n10964), .QN(n10980) );
  NAND3X0 U11578 ( .IN1(n11631), .IN2(n11632), .IN3(n11633), .QN(n10944) );
  NAND2X0 U11579 ( .IN1(n7352), .IN2(g7390), .QN(n11633) );
  NAND2X0 U11580 ( .IN1(n7351), .IN2(g2624), .QN(n11632) );
  NAND2X0 U11581 ( .IN1(n7350), .IN2(n10186), .QN(n11631) );
  NAND3X0 U11582 ( .IN1(n11634), .IN2(n11635), .IN3(n11636), .QN(n10950) );
  NAND2X0 U11583 ( .IN1(g7390), .IN2(n8119), .QN(n11636) );
  NAND2X0 U11584 ( .IN1(n7178), .IN2(g2624), .QN(n11635) );
  NAND2X0 U11585 ( .IN1(n7177), .IN2(n10186), .QN(n11634) );
  INVX0 U11586 ( .INP(n10937), .ZN(n10934) );
  NAND3X0 U11587 ( .IN1(n11637), .IN2(n11638), .IN3(n11639), .QN(n10937) );
  NAND2X0 U11588 ( .IN1(n7340), .IN2(g7390), .QN(n11639) );
  NAND2X0 U11589 ( .IN1(n7339), .IN2(g2624), .QN(n11638) );
  NAND2X0 U11590 ( .IN1(n7338), .IN2(n10186), .QN(n11637) );
  NAND3X0 U11591 ( .IN1(n11640), .IN2(n11641), .IN3(n11642), .QN(n10964) );
  NAND2X0 U11592 ( .IN1(n7363), .IN2(g7390), .QN(n11642) );
  NAND2X0 U11593 ( .IN1(n7362), .IN2(g2624), .QN(n11641) );
  NAND2X0 U11594 ( .IN1(n7361), .IN2(n10186), .QN(n11640) );
  NOR2X0 U11595 ( .IN1(n10187), .IN2(n11513), .QN(n11474) );
  INVX0 U11596 ( .INP(g22687), .ZN(n11513) );
  INVX0 U11597 ( .INP(g7302), .ZN(n10187) );
  NAND2X0 U11598 ( .IN1(n11643), .IN2(n11644), .QN(g27309) );
  INVX0 U11599 ( .INP(n11645), .ZN(n11644) );
  NOR2X0 U11600 ( .IN1(n11562), .IN2(n7383), .QN(n11645) );
  NAND2X0 U11601 ( .IN1(n11562), .IN2(n11521), .QN(n11643) );
  INVX0 U11602 ( .INP(n11646), .ZN(n11521) );
  NAND2X0 U11603 ( .IN1(n11647), .IN2(n11648), .QN(n11646) );
  NAND2X0 U11604 ( .IN1(n11563), .IN2(n11649), .QN(n11648) );
  NAND3X0 U11605 ( .IN1(n11650), .IN2(n11651), .IN3(n11564), .QN(n11647) );
  NAND2X0 U11606 ( .IN1(n11652), .IN2(n11653), .QN(g27308) );
  INVX0 U11607 ( .INP(n11654), .ZN(n11653) );
  NOR2X0 U11608 ( .IN1(n11517), .IN2(n7633), .QN(n11654) );
  NAND2X0 U11609 ( .IN1(n11572), .IN2(n11517), .QN(n11652) );
  NAND2X0 U11610 ( .IN1(n11655), .IN2(n11656), .QN(g27307) );
  INVX0 U11611 ( .INP(n11657), .ZN(n11656) );
  NOR2X0 U11612 ( .IN1(n11485), .IN2(n7655), .QN(n11657) );
  NAND2X0 U11613 ( .IN1(n11658), .IN2(n11485), .QN(n11655) );
  NOR2X0 U11614 ( .IN1(n11659), .IN2(n4509), .QN(n11485) );
  NAND2X0 U11615 ( .IN1(n11660), .IN2(n11661), .QN(g27306) );
  INVX0 U11616 ( .INP(n11662), .ZN(n11661) );
  NOR2X0 U11617 ( .IN1(n11524), .IN2(n7353), .QN(n11662) );
  NAND2X0 U11618 ( .IN1(n11524), .IN2(n11533), .QN(n11660) );
  INVX0 U11619 ( .INP(n11663), .ZN(n11533) );
  NAND2X0 U11620 ( .IN1(n11664), .IN2(n11665), .QN(n11663) );
  NAND2X0 U11621 ( .IN1(n11579), .IN2(n11083), .QN(n11664) );
  XNOR2X1 U11622 ( .IN1(n8798), .IN2(n11033), .Q(n11579) );
  NAND2X0 U11623 ( .IN1(n11666), .IN2(n11667), .QN(g27305) );
  INVX0 U11624 ( .INP(n11668), .ZN(n11667) );
  NOR2X0 U11625 ( .IN1(n11490), .IN2(n7343), .QN(n11668) );
  NAND2X0 U11626 ( .IN1(n11490), .IN2(n11586), .QN(n11666) );
  NOR2X0 U11627 ( .IN1(n11587), .IN2(n4315), .QN(n11490) );
  NAND2X0 U11628 ( .IN1(n11669), .IN2(n11670), .QN(g27304) );
  NAND2X0 U11629 ( .IN1(n11671), .IN2(n11538), .QN(n11670) );
  NAND3X0 U11630 ( .IN1(n11672), .IN2(n11673), .IN3(n11674), .QN(n11538) );
  INVX0 U11631 ( .INP(n11675), .ZN(n11669) );
  NOR2X0 U11632 ( .IN1(n11671), .IN2(n7648), .QN(n11675) );
  NAND2X0 U11633 ( .IN1(n11676), .IN2(n11677), .QN(g27303) );
  NAND2X0 U11634 ( .IN1(n11591), .IN2(g1754), .QN(n11677) );
  NAND2X0 U11635 ( .IN1(n11590), .IN2(n11595), .QN(n11676) );
  NAND2X0 U11636 ( .IN1(n11678), .IN2(n11679), .QN(g27302) );
  INVX0 U11637 ( .INP(n11680), .ZN(n11679) );
  NOR2X0 U11638 ( .IN1(n11537), .IN2(n7635), .QN(n11680) );
  NAND2X0 U11639 ( .IN1(n11681), .IN2(n11537), .QN(n11678) );
  NAND2X0 U11640 ( .IN1(n11682), .IN2(n11683), .QN(g27301) );
  NAND2X0 U11641 ( .IN1(n11600), .IN2(g1268), .QN(n11683) );
  NAND2X0 U11642 ( .IN1(n11598), .IN2(n11545), .QN(n11682) );
  INVX0 U11643 ( .INP(n11684), .ZN(n11545) );
  NAND2X0 U11644 ( .IN1(n11685), .IN2(n11686), .QN(n11684) );
  NAND2X0 U11645 ( .IN1(n11687), .IN2(n11187), .QN(n11686) );
  NAND2X0 U11646 ( .IN1(n11599), .IN2(n11156), .QN(n11685) );
  INVX0 U11647 ( .INP(n11687), .ZN(n11599) );
  NAND2X0 U11648 ( .IN1(n11688), .IN2(n11689), .QN(g27300) );
  INVX0 U11649 ( .INP(n11690), .ZN(n11689) );
  NOR2X0 U11650 ( .IN1(n11541), .IN2(n7358), .QN(n11690) );
  NAND2X0 U11651 ( .IN1(n11541), .IN2(n11606), .QN(n11688) );
  NAND2X0 U11652 ( .IN1(n11691), .IN2(n11692), .QN(g27299) );
  NAND2X0 U11653 ( .IN1(n11497), .IN2(g1261), .QN(n11692) );
  NAND2X0 U11654 ( .IN1(n11498), .IN2(n11693), .QN(n11691) );
  INVX0 U11655 ( .INP(n11497), .ZN(n11498) );
  NAND2X0 U11656 ( .IN1(g1236), .IN2(g22615), .QN(n11497) );
  NAND2X0 U11657 ( .IN1(n11694), .IN2(n11695), .QN(g27298) );
  INVX0 U11658 ( .INP(n11696), .ZN(n11695) );
  NOR2X0 U11659 ( .IN1(n11697), .IN2(n7650), .QN(n11696) );
  NAND2X0 U11660 ( .IN1(n11697), .IN2(n11611), .QN(n11694) );
  NAND2X0 U11661 ( .IN1(n11698), .IN2(n11699), .QN(g27297) );
  INVX0 U11662 ( .INP(n11700), .ZN(n11699) );
  NOR2X0 U11663 ( .IN1(n11610), .IN2(n7390), .QN(n11700) );
  NAND2X0 U11664 ( .IN1(n11610), .IN2(n11701), .QN(n11698) );
  NAND2X0 U11665 ( .IN1(n11702), .IN2(n11703), .QN(g27296) );
  NAND2X0 U11666 ( .IN1(n11704), .IN2(n11550), .QN(n11703) );
  NAND2X0 U11667 ( .IN1(n11705), .IN2(n11259), .QN(n11550) );
  NOR2X0 U11668 ( .IN1(n11254), .IN2(n11284), .QN(n11259) );
  NAND2X0 U11669 ( .IN1(n11706), .IN2(g585), .QN(n11702) );
  NAND2X0 U11670 ( .IN1(n11707), .IN2(n11708), .QN(g27295) );
  NAND2X0 U11671 ( .IN1(n11615), .IN2(g583), .QN(n11708) );
  NAND2X0 U11672 ( .IN1(n11614), .IN2(n11619), .QN(n11707) );
  NAND2X0 U11673 ( .IN1(n11709), .IN2(n11710), .QN(g27294) );
  INVX0 U11674 ( .INP(n11711), .ZN(n11710) );
  NOR2X0 U11675 ( .IN1(n11549), .IN2(n7360), .QN(n11711) );
  NAND2X0 U11676 ( .IN1(n11549), .IN2(n11712), .QN(n11709) );
  NAND2X0 U11677 ( .IN1(n11713), .IN2(n11714), .QN(g27293) );
  NAND2X0 U11678 ( .IN1(n11715), .IN2(g391), .QN(n11714) );
  NAND2X0 U11679 ( .IN1(n11716), .IN2(n11717), .QN(n11713) );
  NAND2X0 U11680 ( .IN1(n11718), .IN2(n11719), .QN(g27292) );
  INVX0 U11681 ( .INP(n11720), .ZN(n11719) );
  NOR2X0 U11682 ( .IN1(n11562), .IN2(n7634), .QN(n11720) );
  NAND2X0 U11683 ( .IN1(n11572), .IN2(n11562), .QN(n11718) );
  NAND2X0 U11684 ( .IN1(n11721), .IN2(n11722), .QN(n11572) );
  NAND2X0 U11685 ( .IN1(n11565), .IN2(n11564), .QN(n11722) );
  INVX0 U11686 ( .INP(n11649), .ZN(n11564) );
  NAND2X0 U11687 ( .IN1(n11563), .IN2(n11723), .QN(n11721) );
  INVX0 U11688 ( .INP(n11651), .ZN(n11563) );
  XOR2X1 U11689 ( .IN1(n8798), .IN2(n11724), .Q(n11651) );
  NAND2X0 U11690 ( .IN1(n11725), .IN2(n11726), .QN(g27291) );
  INVX0 U11691 ( .INP(n11727), .ZN(n11726) );
  NOR2X0 U11692 ( .IN1(n11517), .IN2(n7656), .QN(n11727) );
  NAND2X0 U11693 ( .IN1(n11658), .IN2(n11517), .QN(n11725) );
  NOR2X0 U11694 ( .IN1(n11659), .IN2(n11728), .QN(n11517) );
  INVX0 U11695 ( .INP(g7264), .ZN(n11728) );
  NAND2X0 U11696 ( .IN1(n11729), .IN2(n11730), .QN(g27290) );
  INVX0 U11697 ( .INP(n11731), .ZN(n11730) );
  NOR2X0 U11698 ( .IN1(n11524), .IN2(n7341), .QN(n11731) );
  NAND2X0 U11699 ( .IN1(n11524), .IN2(n11586), .QN(n11729) );
  NOR2X0 U11700 ( .IN1(n11732), .IN2(n11733), .QN(n11586) );
  NOR2X0 U11701 ( .IN1(n11734), .IN2(g3229), .QN(n11733) );
  INVX0 U11702 ( .INP(n11735), .ZN(n11734) );
  NAND2X0 U11703 ( .IN1(n11665), .IN2(n11736), .QN(n11735) );
  NAND2X0 U11704 ( .IN1(n11049), .IN2(n11044), .QN(n11736) );
  INVX0 U11705 ( .INP(n11062), .ZN(n11049) );
  NAND2X0 U11706 ( .IN1(n11047), .IN2(n11053), .QN(n11665) );
  INVX0 U11707 ( .INP(n11083), .ZN(n11047) );
  NOR2X0 U11708 ( .IN1(n8798), .IN2(n11737), .QN(n11732) );
  NOR2X0 U11709 ( .IN1(n11062), .IN2(n11738), .QN(n11737) );
  NOR2X0 U11710 ( .IN1(n11033), .IN2(n11739), .QN(n11738) );
  NOR2X0 U11711 ( .IN1(n11083), .IN2(n11084), .QN(n11739) );
  NOR2X0 U11712 ( .IN1(n11062), .IN2(n11053), .QN(n11084) );
  NAND3X0 U11713 ( .IN1(n11740), .IN2(n11741), .IN3(n11742), .QN(n11053) );
  NAND2X0 U11714 ( .IN1(n7354), .IN2(g1930), .QN(n11742) );
  NAND2X0 U11715 ( .IN1(n7353), .IN2(n10234), .QN(n11741) );
  NAND2X0 U11716 ( .IN1(n7355), .IN2(g7194), .QN(n11740) );
  NAND3X0 U11717 ( .IN1(n11743), .IN2(n11744), .IN3(n11745), .QN(n11083) );
  NAND2X0 U11718 ( .IN1(n7180), .IN2(g1930), .QN(n11745) );
  NAND2X0 U11719 ( .IN1(n7179), .IN2(n10234), .QN(n11744) );
  NAND2X0 U11720 ( .IN1(n7181), .IN2(g7194), .QN(n11743) );
  INVX0 U11721 ( .INP(n11044), .ZN(n11033) );
  NAND3X0 U11722 ( .IN1(n11746), .IN2(n11747), .IN3(n11748), .QN(n11044) );
  NAND2X0 U11723 ( .IN1(n7342), .IN2(g1930), .QN(n11748) );
  NAND2X0 U11724 ( .IN1(n7341), .IN2(n10234), .QN(n11747) );
  NAND2X0 U11725 ( .IN1(n7343), .IN2(g7194), .QN(n11746) );
  NAND3X0 U11726 ( .IN1(n11749), .IN2(n11750), .IN3(n11751), .QN(n11062) );
  NAND2X0 U11727 ( .IN1(n7364), .IN2(g1930), .QN(n11751) );
  NAND2X0 U11728 ( .IN1(n10234), .IN2(n8109), .QN(n11750) );
  NAND2X0 U11729 ( .IN1(n7365), .IN2(g7194), .QN(n11749) );
  NOR2X0 U11730 ( .IN1(n10235), .IN2(n11587), .QN(n11524) );
  INVX0 U11731 ( .INP(g22651), .ZN(n11587) );
  INVX0 U11732 ( .INP(g7052), .ZN(n10235) );
  NAND2X0 U11733 ( .IN1(n11752), .IN2(n11753), .QN(g27289) );
  INVX0 U11734 ( .INP(n11754), .ZN(n11753) );
  NOR2X0 U11735 ( .IN1(n11671), .IN2(n7386), .QN(n11754) );
  NAND2X0 U11736 ( .IN1(n11671), .IN2(n11595), .QN(n11752) );
  INVX0 U11737 ( .INP(n11755), .ZN(n11595) );
  NAND2X0 U11738 ( .IN1(n11756), .IN2(n11757), .QN(n11755) );
  NAND2X0 U11739 ( .IN1(n11672), .IN2(n11758), .QN(n11757) );
  NAND3X0 U11740 ( .IN1(n11759), .IN2(n11760), .IN3(n11673), .QN(n11756) );
  NAND2X0 U11741 ( .IN1(n11761), .IN2(n11762), .QN(g27288) );
  NAND2X0 U11742 ( .IN1(n11591), .IN2(g1739), .QN(n11762) );
  NAND2X0 U11743 ( .IN1(n11681), .IN2(n11590), .QN(n11761) );
  NAND2X0 U11744 ( .IN1(n11763), .IN2(n11764), .QN(g27287) );
  INVX0 U11745 ( .INP(n11765), .ZN(n11764) );
  NOR2X0 U11746 ( .IN1(n11537), .IN2(n7658), .QN(n11765) );
  NAND2X0 U11747 ( .IN1(n11766), .IN2(n11537), .QN(n11763) );
  INVX0 U11748 ( .INP(n11767), .ZN(n11537) );
  NAND2X0 U11749 ( .IN1(n11768), .IN2(n10093), .QN(n11767) );
  NAND2X0 U11750 ( .IN1(n11769), .IN2(n11770), .QN(g27286) );
  NAND2X0 U11751 ( .IN1(n11600), .IN2(g1265), .QN(n11770) );
  NAND2X0 U11752 ( .IN1(n11598), .IN2(n11606), .QN(n11769) );
  INVX0 U11753 ( .INP(n11771), .ZN(n11606) );
  NAND2X0 U11754 ( .IN1(n11772), .IN2(n11773), .QN(n11771) );
  NAND2X0 U11755 ( .IN1(n11687), .IN2(n11186), .QN(n11772) );
  XNOR2X1 U11756 ( .IN1(n8798), .IN2(n11136), .Q(n11687) );
  NAND2X0 U11757 ( .IN1(n11774), .IN2(n11775), .QN(g27285) );
  INVX0 U11758 ( .INP(n11776), .ZN(n11775) );
  NOR2X0 U11759 ( .IN1(n11541), .IN2(n7346), .QN(n11776) );
  NAND2X0 U11760 ( .IN1(n11541), .IN2(n11693), .QN(n11774) );
  NOR2X0 U11761 ( .IN1(n4316), .IN2(n11777), .QN(n11541) );
  INVX0 U11762 ( .INP(g22615), .ZN(n11777) );
  NAND2X0 U11763 ( .IN1(n11778), .IN2(n11779), .QN(g27284) );
  NAND2X0 U11764 ( .IN1(n11780), .IN2(g1085), .QN(n11779) );
  NAND2X0 U11765 ( .IN1(n11781), .IN2(n11611), .QN(n11778) );
  NAND3X0 U11766 ( .IN1(n11782), .IN2(n11783), .IN3(n11784), .QN(n11611) );
  NAND2X0 U11767 ( .IN1(n11785), .IN2(n11786), .QN(g27283) );
  INVX0 U11768 ( .INP(n11787), .ZN(n11786) );
  NOR2X0 U11769 ( .IN1(n11697), .IN2(n7389), .QN(n11787) );
  NAND2X0 U11770 ( .IN1(n11697), .IN2(n11701), .QN(n11785) );
  NAND2X0 U11771 ( .IN1(n11788), .IN2(n11789), .QN(g27282) );
  INVX0 U11772 ( .INP(n11790), .ZN(n11789) );
  NOR2X0 U11773 ( .IN1(n11610), .IN2(n7638), .QN(n11790) );
  NAND2X0 U11774 ( .IN1(n11791), .IN2(n11610), .QN(n11788) );
  NAND2X0 U11775 ( .IN1(n11792), .IN2(n11793), .QN(g27281) );
  NAND2X0 U11776 ( .IN1(n11706), .IN2(g582), .QN(n11793) );
  NAND2X0 U11777 ( .IN1(n11704), .IN2(n11619), .QN(n11792) );
  INVX0 U11778 ( .INP(n11794), .ZN(n11619) );
  NAND2X0 U11779 ( .IN1(n11795), .IN2(n11796), .QN(n11794) );
  NAND2X0 U11780 ( .IN1(n11797), .IN2(n11285), .QN(n11796) );
  NAND2X0 U11781 ( .IN1(n11705), .IN2(n11254), .QN(n11795) );
  INVX0 U11782 ( .INP(n11797), .ZN(n11705) );
  NAND2X0 U11783 ( .IN1(n11798), .IN2(n11799), .QN(g27280) );
  NAND2X0 U11784 ( .IN1(test_so25), .IN2(n11615), .QN(n11799) );
  NAND2X0 U11785 ( .IN1(n11614), .IN2(n11712), .QN(n11798) );
  NAND2X0 U11786 ( .IN1(n11800), .IN2(n11801), .QN(g27279) );
  INVX0 U11787 ( .INP(n11802), .ZN(n11801) );
  NOR2X0 U11788 ( .IN1(n11549), .IN2(n7348), .QN(n11802) );
  NAND2X0 U11789 ( .IN1(n11549), .IN2(n11803), .QN(n11800) );
  NOR2X0 U11790 ( .IN1(n4313), .IN2(n11804), .QN(n11549) );
  NAND2X0 U11791 ( .IN1(n11805), .IN2(n11806), .QN(g27278) );
  NAND2X0 U11792 ( .IN1(n11807), .IN2(g388), .QN(n11806) );
  NAND2X0 U11793 ( .IN1(n11808), .IN2(n11717), .QN(n11805) );
  NAND2X0 U11794 ( .IN1(n11809), .IN2(n11810), .QN(g27277) );
  NAND2X0 U11795 ( .IN1(n11715), .IN2(g376), .QN(n11810) );
  NAND2X0 U11796 ( .IN1(n11716), .IN2(n11811), .QN(n11809) );
  NAND2X0 U11797 ( .IN1(n11812), .IN2(n11813), .QN(g27276) );
  INVX0 U11798 ( .INP(n11814), .ZN(n11813) );
  NOR2X0 U11799 ( .IN1(n11562), .IN2(n7657), .QN(n11814) );
  NAND2X0 U11800 ( .IN1(n11658), .IN2(n11562), .QN(n11812) );
  NOR2X0 U11801 ( .IN1(n11659), .IN2(n11815), .QN(n11562) );
  INVX0 U11802 ( .INP(g5555), .ZN(n11815) );
  NAND2X0 U11803 ( .IN1(n8680), .IN2(n11816), .QN(n11659) );
  NAND2X0 U11804 ( .IN1(n11817), .IN2(n8657), .QN(n11816) );
  INVX0 U11805 ( .INP(n10036), .ZN(n8657) );
  INVX0 U11806 ( .INP(n11818), .ZN(n11658) );
  NAND3X0 U11807 ( .IN1(n11819), .IN2(n11820), .IN3(n11821), .QN(n11818) );
  NAND2X0 U11808 ( .IN1(g3229), .IN2(n11822), .QN(n11821) );
  INVX0 U11809 ( .INP(n11823), .ZN(n11820) );
  NOR2X0 U11810 ( .IN1(n11824), .IN2(g3229), .QN(n11823) );
  NAND3X0 U11811 ( .IN1(n11650), .IN2(n11724), .IN3(n11824), .QN(n11819) );
  NAND2X0 U11812 ( .IN1(n11565), .IN2(n11649), .QN(n11824) );
  NAND3X0 U11813 ( .IN1(n11825), .IN2(n11826), .IN3(n11827), .QN(n11649) );
  NAND2X0 U11814 ( .IN1(n7633), .IN2(n10046), .QN(n11827) );
  NAND2X0 U11815 ( .IN1(n7632), .IN2(n10047), .QN(n11826) );
  NAND2X0 U11816 ( .IN1(n7634), .IN2(n10048), .QN(n11825) );
  INVX0 U11817 ( .INP(n11723), .ZN(n11565) );
  NAND3X0 U11818 ( .IN1(n11828), .IN2(n11829), .IN3(n11830), .QN(n11723) );
  NAND2X0 U11819 ( .IN1(n7385), .IN2(n10046), .QN(n11830) );
  NAND2X0 U11820 ( .IN1(n7384), .IN2(n10047), .QN(n11829) );
  NAND2X0 U11821 ( .IN1(n7383), .IN2(n10048), .QN(n11828) );
  NAND3X0 U11822 ( .IN1(n11831), .IN2(n11832), .IN3(n11833), .QN(n11724) );
  NAND2X0 U11823 ( .IN1(n7656), .IN2(n10046), .QN(n11833) );
  NAND2X0 U11824 ( .IN1(n7655), .IN2(n10047), .QN(n11832) );
  NAND2X0 U11825 ( .IN1(n7657), .IN2(n10048), .QN(n11831) );
  INVX0 U11826 ( .INP(n11822), .ZN(n11650) );
  NAND3X0 U11827 ( .IN1(n11834), .IN2(n11835), .IN3(n11836), .QN(n11822) );
  NAND2X0 U11828 ( .IN1(n7645), .IN2(n10046), .QN(n11836) );
  NAND2X0 U11829 ( .IN1(n7644), .IN2(n10047), .QN(n11835) );
  NAND2X0 U11830 ( .IN1(n7646), .IN2(n10048), .QN(n11834) );
  NAND2X0 U11831 ( .IN1(n11837), .IN2(n11838), .QN(g27275) );
  INVX0 U11832 ( .INP(n11839), .ZN(n11838) );
  NOR2X0 U11833 ( .IN1(n11671), .IN2(n7637), .QN(n11839) );
  NAND2X0 U11834 ( .IN1(n11681), .IN2(n11671), .QN(n11837) );
  NAND2X0 U11835 ( .IN1(n11840), .IN2(n11841), .QN(n11681) );
  NAND2X0 U11836 ( .IN1(n11674), .IN2(n11673), .QN(n11841) );
  INVX0 U11837 ( .INP(n11758), .ZN(n11673) );
  NAND2X0 U11838 ( .IN1(n11672), .IN2(n11842), .QN(n11840) );
  INVX0 U11839 ( .INP(n11760), .ZN(n11672) );
  XOR2X1 U11840 ( .IN1(n8798), .IN2(n11843), .Q(n11760) );
  NAND2X0 U11841 ( .IN1(n11844), .IN2(n11845), .QN(g27274) );
  NAND2X0 U11842 ( .IN1(n11591), .IN2(g1724), .QN(n11845) );
  NAND2X0 U11843 ( .IN1(n11766), .IN2(n11590), .QN(n11844) );
  INVX0 U11844 ( .INP(n11591), .ZN(n11590) );
  NAND2X0 U11845 ( .IN1(n11768), .IN2(g7014), .QN(n11591) );
  NAND2X0 U11846 ( .IN1(n11846), .IN2(n11847), .QN(g27273) );
  NAND2X0 U11847 ( .IN1(n11600), .IN2(g1262), .QN(n11847) );
  NAND2X0 U11848 ( .IN1(n11598), .IN2(n11693), .QN(n11846) );
  NOR2X0 U11849 ( .IN1(n11848), .IN2(n11849), .QN(n11693) );
  NOR2X0 U11850 ( .IN1(n11850), .IN2(g3229), .QN(n11849) );
  INVX0 U11851 ( .INP(n11851), .ZN(n11850) );
  NAND2X0 U11852 ( .IN1(n11773), .IN2(n11852), .QN(n11851) );
  NAND2X0 U11853 ( .IN1(n11152), .IN2(n11147), .QN(n11852) );
  INVX0 U11854 ( .INP(n11165), .ZN(n11152) );
  NAND2X0 U11855 ( .IN1(n11150), .IN2(n11156), .QN(n11773) );
  INVX0 U11856 ( .INP(n11186), .ZN(n11150) );
  NOR2X0 U11857 ( .IN1(n8798), .IN2(n11853), .QN(n11848) );
  NOR2X0 U11858 ( .IN1(n11165), .IN2(n11854), .QN(n11853) );
  NOR2X0 U11859 ( .IN1(n11136), .IN2(n11855), .QN(n11854) );
  NOR2X0 U11860 ( .IN1(n11186), .IN2(n11187), .QN(n11855) );
  NOR2X0 U11861 ( .IN1(n11165), .IN2(n11156), .QN(n11187) );
  NAND3X0 U11862 ( .IN1(n11856), .IN2(n11857), .IN3(n11858), .QN(n11156) );
  NAND2X0 U11863 ( .IN1(n7356), .IN2(n11110), .QN(n11858) );
  NAND2X0 U11864 ( .IN1(n7357), .IN2(g1236), .QN(n11857) );
  NAND2X0 U11865 ( .IN1(n7358), .IN2(g6944), .QN(n11856) );
  NAND3X0 U11866 ( .IN1(n11859), .IN2(n11860), .IN3(n11861), .QN(n11186) );
  NAND2X0 U11867 ( .IN1(n7182), .IN2(n11110), .QN(n11861) );
  NAND2X0 U11868 ( .IN1(g1236), .IN2(n8120), .QN(n11860) );
  NAND2X0 U11869 ( .IN1(n7183), .IN2(g6944), .QN(n11859) );
  INVX0 U11870 ( .INP(n11147), .ZN(n11136) );
  NAND3X0 U11871 ( .IN1(n11862), .IN2(n11863), .IN3(n11864), .QN(n11147) );
  NAND2X0 U11872 ( .IN1(n7344), .IN2(n11110), .QN(n11864) );
  NAND2X0 U11873 ( .IN1(n7345), .IN2(g1236), .QN(n11863) );
  NAND2X0 U11874 ( .IN1(n7346), .IN2(g6944), .QN(n11862) );
  NAND3X0 U11875 ( .IN1(n11865), .IN2(n11866), .IN3(n11867), .QN(n11165) );
  NAND2X0 U11876 ( .IN1(n7366), .IN2(n11110), .QN(n11867) );
  NAND2X0 U11877 ( .IN1(n7367), .IN2(g1236), .QN(n11866) );
  NAND2X0 U11878 ( .IN1(n7368), .IN2(g6944), .QN(n11865) );
  INVX0 U11879 ( .INP(n11600), .ZN(n11598) );
  NAND2X0 U11880 ( .IN1(g6750), .IN2(g22615), .QN(n11600) );
  NAND2X0 U11881 ( .IN1(n11868), .IN2(n11869), .QN(g27272) );
  NAND2X0 U11882 ( .IN1(test_so37), .IN2(n11780), .QN(n11869) );
  NAND2X0 U11883 ( .IN1(n11781), .IN2(n11701), .QN(n11868) );
  INVX0 U11884 ( .INP(n11870), .ZN(n11701) );
  NAND2X0 U11885 ( .IN1(n11871), .IN2(n11872), .QN(n11870) );
  NAND2X0 U11886 ( .IN1(n11782), .IN2(n11873), .QN(n11872) );
  NAND3X0 U11887 ( .IN1(n11874), .IN2(n11875), .IN3(n11783), .QN(n11871) );
  NAND2X0 U11888 ( .IN1(n11876), .IN2(n11877), .QN(g27271) );
  INVX0 U11889 ( .INP(n11878), .ZN(n11877) );
  NOR2X0 U11890 ( .IN1(n11697), .IN2(n7639), .QN(n11878) );
  NAND2X0 U11891 ( .IN1(n11791), .IN2(n11697), .QN(n11876) );
  NAND2X0 U11892 ( .IN1(n11879), .IN2(n11880), .QN(g27270) );
  INVX0 U11893 ( .INP(n11881), .ZN(n11880) );
  NOR2X0 U11894 ( .IN1(n11610), .IN2(n7661), .QN(n11881) );
  NAND2X0 U11895 ( .IN1(n11882), .IN2(n11610), .QN(n11879) );
  NOR2X0 U11896 ( .IN1(n11883), .IN2(n4381), .QN(n11610) );
  NAND2X0 U11897 ( .IN1(n11884), .IN2(n11885), .QN(g27269) );
  NAND2X0 U11898 ( .IN1(n11706), .IN2(g579), .QN(n11885) );
  NAND2X0 U11899 ( .IN1(n11704), .IN2(n11712), .QN(n11884) );
  INVX0 U11900 ( .INP(n11886), .ZN(n11712) );
  NAND2X0 U11901 ( .IN1(n11887), .IN2(n11888), .QN(n11886) );
  NAND2X0 U11902 ( .IN1(n11797), .IN2(n11284), .QN(n11887) );
  XNOR2X1 U11903 ( .IN1(n8798), .IN2(n11234), .Q(n11797) );
  NAND2X0 U11904 ( .IN1(n11889), .IN2(n11890), .QN(g27268) );
  NAND2X0 U11905 ( .IN1(n11615), .IN2(g577), .QN(n11890) );
  INVX0 U11906 ( .INP(n11614), .ZN(n11615) );
  NAND2X0 U11907 ( .IN1(n11614), .IN2(n11803), .QN(n11889) );
  NOR2X0 U11908 ( .IN1(n4372), .IN2(n11804), .QN(n11614) );
  INVX0 U11909 ( .INP(g22578), .ZN(n11804) );
  NAND2X0 U11910 ( .IN1(n11891), .IN2(n11892), .QN(g27267) );
  NAND2X0 U11911 ( .IN1(n11893), .IN2(g398), .QN(n11892) );
  NAND2X0 U11912 ( .IN1(n11894), .IN2(n11717), .QN(n11891) );
  NAND3X0 U11913 ( .IN1(n11895), .IN2(n11896), .IN3(n11897), .QN(n11717) );
  NAND2X0 U11914 ( .IN1(n11898), .IN2(n11899), .QN(g27266) );
  NAND2X0 U11915 ( .IN1(n11807), .IN2(g373), .QN(n11899) );
  NAND2X0 U11916 ( .IN1(n11808), .IN2(n11811), .QN(n11898) );
  NAND2X0 U11917 ( .IN1(n11900), .IN2(n11901), .QN(g27265) );
  NAND2X0 U11918 ( .IN1(n11715), .IN2(g361), .QN(n11901) );
  NAND2X0 U11919 ( .IN1(n11902), .IN2(n11716), .QN(n11900) );
  NAND2X0 U11920 ( .IN1(n11903), .IN2(n11904), .QN(g27264) );
  INVX0 U11921 ( .INP(n11905), .ZN(n11904) );
  NOR2X0 U11922 ( .IN1(n11671), .IN2(n7660), .QN(n11905) );
  NAND2X0 U11923 ( .IN1(n11766), .IN2(n11671), .QN(n11903) );
  INVX0 U11924 ( .INP(n11906), .ZN(n11671) );
  NAND2X0 U11925 ( .IN1(n11768), .IN2(g5511), .QN(n11906) );
  NOR2X0 U11926 ( .IN1(n11907), .IN2(n11908), .QN(n11768) );
  NOR2X0 U11927 ( .IN1(n8591), .IN2(n8628), .QN(n11908) );
  INVX0 U11928 ( .INP(n11909), .ZN(n11766) );
  NAND3X0 U11929 ( .IN1(n11910), .IN2(n11911), .IN3(n11912), .QN(n11909) );
  NAND2X0 U11930 ( .IN1(g3229), .IN2(n11913), .QN(n11912) );
  INVX0 U11931 ( .INP(n11914), .ZN(n11911) );
  NOR2X0 U11932 ( .IN1(n11915), .IN2(g3229), .QN(n11914) );
  NAND3X0 U11933 ( .IN1(n11759), .IN2(n11843), .IN3(n11915), .QN(n11910) );
  NAND2X0 U11934 ( .IN1(n11674), .IN2(n11758), .QN(n11915) );
  NAND3X0 U11935 ( .IN1(n11916), .IN2(n11917), .IN3(n11918), .QN(n11758) );
  NAND2X0 U11936 ( .IN1(n7636), .IN2(n10092), .QN(n11918) );
  NAND2X0 U11937 ( .IN1(n7635), .IN2(n10093), .QN(n11917) );
  NAND2X0 U11938 ( .IN1(n7637), .IN2(n10094), .QN(n11916) );
  INVX0 U11939 ( .INP(n11842), .ZN(n11674) );
  NAND3X0 U11940 ( .IN1(n11919), .IN2(n11920), .IN3(n11921), .QN(n11842) );
  NAND2X0 U11941 ( .IN1(n7388), .IN2(n10092), .QN(n11921) );
  NAND2X0 U11942 ( .IN1(n7387), .IN2(n10093), .QN(n11920) );
  NAND2X0 U11943 ( .IN1(n7386), .IN2(n10094), .QN(n11919) );
  NAND3X0 U11944 ( .IN1(n11922), .IN2(n11923), .IN3(n11924), .QN(n11843) );
  NAND2X0 U11945 ( .IN1(n7659), .IN2(n10092), .QN(n11924) );
  NAND2X0 U11946 ( .IN1(n7658), .IN2(n10093), .QN(n11923) );
  NAND2X0 U11947 ( .IN1(n7660), .IN2(n10094), .QN(n11922) );
  INVX0 U11948 ( .INP(n11913), .ZN(n11759) );
  NAND3X0 U11949 ( .IN1(n11925), .IN2(n11926), .IN3(n11927), .QN(n11913) );
  NAND2X0 U11950 ( .IN1(n10092), .IN2(n8113), .QN(n11927) );
  NAND2X0 U11951 ( .IN1(n7647), .IN2(n10093), .QN(n11926) );
  NAND2X0 U11952 ( .IN1(n7648), .IN2(n10094), .QN(n11925) );
  NAND2X0 U11953 ( .IN1(n11928), .IN2(n11929), .QN(g27263) );
  NAND2X0 U11954 ( .IN1(n11780), .IN2(g1056), .QN(n11929) );
  NAND2X0 U11955 ( .IN1(n11791), .IN2(n11781), .QN(n11928) );
  NAND2X0 U11956 ( .IN1(n11930), .IN2(n11931), .QN(n11791) );
  NAND2X0 U11957 ( .IN1(n11784), .IN2(n11783), .QN(n11931) );
  INVX0 U11958 ( .INP(n11873), .ZN(n11783) );
  NAND2X0 U11959 ( .IN1(n11782), .IN2(n11932), .QN(n11930) );
  INVX0 U11960 ( .INP(n11875), .ZN(n11782) );
  XOR2X1 U11961 ( .IN1(n8798), .IN2(n11933), .Q(n11875) );
  NAND2X0 U11962 ( .IN1(n11934), .IN2(n11935), .QN(g27262) );
  INVX0 U11963 ( .INP(n11936), .ZN(n11935) );
  NOR2X0 U11964 ( .IN1(n11697), .IN2(n7662), .QN(n11936) );
  NAND2X0 U11965 ( .IN1(n11882), .IN2(n11697), .QN(n11934) );
  NOR2X0 U11966 ( .IN1(n11883), .IN2(n4364), .QN(n11697) );
  NAND2X0 U11967 ( .IN1(n11937), .IN2(n11938), .QN(g27261) );
  NAND2X0 U11968 ( .IN1(n11706), .IN2(g576), .QN(n11938) );
  NAND2X0 U11969 ( .IN1(n11704), .IN2(n11803), .QN(n11937) );
  NOR2X0 U11970 ( .IN1(n11939), .IN2(n11940), .QN(n11803) );
  NOR2X0 U11971 ( .IN1(n11941), .IN2(g3229), .QN(n11940) );
  INVX0 U11972 ( .INP(n11942), .ZN(n11941) );
  NAND2X0 U11973 ( .IN1(n11888), .IN2(n11943), .QN(n11942) );
  NAND2X0 U11974 ( .IN1(n11250), .IN2(n11245), .QN(n11943) );
  INVX0 U11975 ( .INP(n11263), .ZN(n11250) );
  NAND2X0 U11976 ( .IN1(n11248), .IN2(n11254), .QN(n11888) );
  INVX0 U11977 ( .INP(n11284), .ZN(n11248) );
  NOR2X0 U11978 ( .IN1(n8798), .IN2(n11944), .QN(n11939) );
  NOR2X0 U11979 ( .IN1(n11263), .IN2(n11945), .QN(n11944) );
  NOR2X0 U11980 ( .IN1(n11234), .IN2(n11946), .QN(n11945) );
  NOR2X0 U11981 ( .IN1(n11284), .IN2(n11285), .QN(n11946) );
  NOR2X0 U11982 ( .IN1(n11263), .IN2(n11254), .QN(n11285) );
  NAND3X0 U11983 ( .IN1(n11947), .IN2(n11948), .IN3(n11949), .QN(n11254) );
  NAND2X0 U11984 ( .IN1(g6642), .IN2(n8121), .QN(n11949) );
  NAND2X0 U11985 ( .IN1(n7359), .IN2(n11213), .QN(n11948) );
  NAND2X0 U11986 ( .IN1(n7360), .IN2(g550), .QN(n11947) );
  NAND3X0 U11987 ( .IN1(n11950), .IN2(n11951), .IN3(n11952), .QN(n11284) );
  NAND2X0 U11988 ( .IN1(n7186), .IN2(g6642), .QN(n11952) );
  NAND2X0 U11989 ( .IN1(n7184), .IN2(n11213), .QN(n11951) );
  NAND2X0 U11990 ( .IN1(n7185), .IN2(g550), .QN(n11950) );
  INVX0 U11991 ( .INP(n11245), .ZN(n11234) );
  NAND3X0 U11992 ( .IN1(n11953), .IN2(n11954), .IN3(n11955), .QN(n11245) );
  NAND2X0 U11993 ( .IN1(n7349), .IN2(g6642), .QN(n11955) );
  NAND2X0 U11994 ( .IN1(n7347), .IN2(n11213), .QN(n11954) );
  NAND2X0 U11995 ( .IN1(n7348), .IN2(g550), .QN(n11953) );
  NAND3X0 U11996 ( .IN1(n11956), .IN2(n11957), .IN3(n11958), .QN(n11263) );
  NAND2X0 U11997 ( .IN1(n7371), .IN2(g6642), .QN(n11958) );
  NAND2X0 U11998 ( .IN1(n7369), .IN2(n11213), .QN(n11957) );
  NAND2X0 U11999 ( .IN1(n7370), .IN2(g550), .QN(n11956) );
  INVX0 U12000 ( .INP(n11706), .ZN(n11704) );
  NAND2X0 U12001 ( .IN1(g6485), .IN2(g22578), .QN(n11706) );
  NAND2X0 U12002 ( .IN1(n11959), .IN2(n11960), .QN(g27260) );
  NAND2X0 U12003 ( .IN1(n11893), .IN2(g384), .QN(n11960) );
  NAND2X0 U12004 ( .IN1(n11894), .IN2(n11811), .QN(n11959) );
  INVX0 U12005 ( .INP(n11961), .ZN(n11811) );
  NAND2X0 U12006 ( .IN1(n11962), .IN2(n11963), .QN(n11961) );
  NAND2X0 U12007 ( .IN1(n11895), .IN2(n11964), .QN(n11963) );
  NAND3X0 U12008 ( .IN1(n11965), .IN2(n11966), .IN3(n11896), .QN(n11962) );
  NAND2X0 U12009 ( .IN1(n11967), .IN2(n11968), .QN(g27259) );
  NAND2X0 U12010 ( .IN1(n11807), .IN2(g358), .QN(n11968) );
  NAND2X0 U12011 ( .IN1(n11902), .IN2(n11808), .QN(n11967) );
  NAND2X0 U12012 ( .IN1(n11969), .IN2(n11970), .QN(g27258) );
  NAND2X0 U12013 ( .IN1(test_so16), .IN2(n11715), .QN(n11970) );
  NAND2X0 U12014 ( .IN1(n11971), .IN2(n11716), .QN(n11969) );
  INVX0 U12015 ( .INP(n11715), .ZN(n11716) );
  NAND2X0 U12016 ( .IN1(n11972), .IN2(n10178), .QN(n11715) );
  NAND2X0 U12017 ( .IN1(n11973), .IN2(n11974), .QN(g27257) );
  NAND2X0 U12018 ( .IN1(n11780), .IN2(g1041), .QN(n11974) );
  INVX0 U12019 ( .INP(n11781), .ZN(n11780) );
  NAND2X0 U12020 ( .IN1(n11882), .IN2(n11781), .QN(n11973) );
  NOR2X0 U12021 ( .IN1(n11883), .IN2(n4363), .QN(n11781) );
  NAND2X0 U12022 ( .IN1(n8621), .IN2(n11975), .QN(n11883) );
  NAND2X0 U12023 ( .IN1(n11817), .IN2(n8598), .QN(n11975) );
  INVX0 U12024 ( .INP(n10126), .ZN(n8598) );
  INVX0 U12025 ( .INP(n11976), .ZN(n11882) );
  NAND3X0 U12026 ( .IN1(n11977), .IN2(n11978), .IN3(n11979), .QN(n11976) );
  NAND2X0 U12027 ( .IN1(g3229), .IN2(n11980), .QN(n11979) );
  INVX0 U12028 ( .INP(n11981), .ZN(n11978) );
  NOR2X0 U12029 ( .IN1(n11982), .IN2(g3229), .QN(n11981) );
  NAND3X0 U12030 ( .IN1(n11874), .IN2(n11933), .IN3(n11982), .QN(n11977) );
  NAND2X0 U12031 ( .IN1(n11784), .IN2(n11873), .QN(n11982) );
  NAND3X0 U12032 ( .IN1(n11983), .IN2(n11984), .IN3(n11985), .QN(n11873) );
  NAND2X0 U12033 ( .IN1(n7638), .IN2(g1088), .QN(n11985) );
  NAND2X0 U12034 ( .IN1(n7640), .IN2(g5472), .QN(n11984) );
  NAND2X0 U12035 ( .IN1(n7639), .IN2(g6712), .QN(n11983) );
  INVX0 U12036 ( .INP(n11932), .ZN(n11784) );
  NAND3X0 U12037 ( .IN1(n11986), .IN2(n11987), .IN3(n11988), .QN(n11932) );
  NAND2X0 U12038 ( .IN1(n7390), .IN2(g1088), .QN(n11988) );
  NAND2X0 U12039 ( .IN1(g5472), .IN2(n8114), .QN(n11987) );
  NAND2X0 U12040 ( .IN1(n7389), .IN2(g6712), .QN(n11986) );
  NAND3X0 U12041 ( .IN1(n11989), .IN2(n11990), .IN3(n11991), .QN(n11933) );
  NAND2X0 U12042 ( .IN1(n7661), .IN2(g1088), .QN(n11991) );
  NAND2X0 U12043 ( .IN1(n7663), .IN2(g5472), .QN(n11990) );
  NAND2X0 U12044 ( .IN1(n7662), .IN2(g6712), .QN(n11989) );
  INVX0 U12045 ( .INP(n11980), .ZN(n11874) );
  NAND3X0 U12046 ( .IN1(n11992), .IN2(n11993), .IN3(n11994), .QN(n11980) );
  NAND2X0 U12047 ( .IN1(n7649), .IN2(g1088), .QN(n11994) );
  NAND2X0 U12048 ( .IN1(n7651), .IN2(g5472), .QN(n11993) );
  NAND2X0 U12049 ( .IN1(n7650), .IN2(g6712), .QN(n11992) );
  NAND2X0 U12050 ( .IN1(n11995), .IN2(n11996), .QN(g27256) );
  NAND2X0 U12051 ( .IN1(n11893), .IN2(g369), .QN(n11996) );
  NAND2X0 U12052 ( .IN1(n11902), .IN2(n11894), .QN(n11995) );
  NAND2X0 U12053 ( .IN1(n11997), .IN2(n11998), .QN(n11902) );
  NAND2X0 U12054 ( .IN1(n11897), .IN2(n11896), .QN(n11998) );
  INVX0 U12055 ( .INP(n11964), .ZN(n11896) );
  NAND2X0 U12056 ( .IN1(n11895), .IN2(n11999), .QN(n11997) );
  INVX0 U12057 ( .INP(n11966), .ZN(n11895) );
  XOR2X1 U12058 ( .IN1(n8798), .IN2(n12000), .Q(n11966) );
  NAND2X0 U12059 ( .IN1(n12001), .IN2(n12002), .QN(g27255) );
  NAND2X0 U12060 ( .IN1(n11807), .IN2(g343), .QN(n12002) );
  NAND2X0 U12061 ( .IN1(n11971), .IN2(n11808), .QN(n12001) );
  INVX0 U12062 ( .INP(n11807), .ZN(n11808) );
  NAND2X0 U12063 ( .IN1(n11972), .IN2(g6447), .QN(n11807) );
  NAND2X0 U12064 ( .IN1(n12003), .IN2(n12004), .QN(g27253) );
  NAND2X0 U12065 ( .IN1(n11893), .IN2(g354), .QN(n12004) );
  NAND2X0 U12066 ( .IN1(n11971), .IN2(n11894), .QN(n12003) );
  INVX0 U12067 ( .INP(n11893), .ZN(n11894) );
  NAND2X0 U12068 ( .IN1(n11972), .IN2(g5437), .QN(n11893) );
  NOR2X0 U12069 ( .IN1(n12005), .IN2(n12006), .QN(n11972) );
  NOR2X0 U12070 ( .IN1(n8591), .IN2(n8568), .QN(n12006) );
  INVX0 U12071 ( .INP(n12007), .ZN(n11971) );
  NAND3X0 U12072 ( .IN1(n12008), .IN2(n12009), .IN3(n12010), .QN(n12007) );
  NAND2X0 U12073 ( .IN1(g3229), .IN2(n12011), .QN(n12010) );
  INVX0 U12074 ( .INP(n12012), .ZN(n12009) );
  NOR2X0 U12075 ( .IN1(n12013), .IN2(g3229), .QN(n12012) );
  NAND3X0 U12076 ( .IN1(n11965), .IN2(n12000), .IN3(n12013), .QN(n12008) );
  NAND2X0 U12077 ( .IN1(n11897), .IN2(n11964), .QN(n12013) );
  NAND3X0 U12078 ( .IN1(n12014), .IN2(n12015), .IN3(n12016), .QN(n11964) );
  NAND2X0 U12079 ( .IN1(n7643), .IN2(n10176), .QN(n12016) );
  NAND2X0 U12080 ( .IN1(n7642), .IN2(n10177), .QN(n12015) );
  NAND2X0 U12081 ( .IN1(n7641), .IN2(n10178), .QN(n12014) );
  INVX0 U12082 ( .INP(n11999), .ZN(n11897) );
  NAND3X0 U12083 ( .IN1(n12017), .IN2(n12018), .IN3(n12019), .QN(n11999) );
  NAND2X0 U12084 ( .IN1(n7391), .IN2(n10176), .QN(n12019) );
  NAND2X0 U12085 ( .IN1(n7393), .IN2(n10177), .QN(n12018) );
  NAND2X0 U12086 ( .IN1(n7392), .IN2(n10178), .QN(n12017) );
  NAND3X0 U12087 ( .IN1(n12020), .IN2(n12021), .IN3(n12022), .QN(n12000) );
  NAND2X0 U12088 ( .IN1(n7665), .IN2(n10176), .QN(n12022) );
  NAND2X0 U12089 ( .IN1(n7664), .IN2(n10177), .QN(n12021) );
  NAND2X0 U12090 ( .IN1(n10178), .IN2(n8115), .QN(n12020) );
  INVX0 U12091 ( .INP(n12011), .ZN(n11965) );
  NAND3X0 U12092 ( .IN1(n12023), .IN2(n12024), .IN3(n12025), .QN(n12011) );
  NAND2X0 U12093 ( .IN1(n7654), .IN2(n10176), .QN(n12025) );
  NAND2X0 U12094 ( .IN1(n7653), .IN2(n10177), .QN(n12024) );
  NAND2X0 U12095 ( .IN1(n7652), .IN2(n10178), .QN(n12023) );
  NOR3X0 U12096 ( .IN1(n12026), .IN2(n11309), .IN3(n11312), .QN(g27243) );
  NOR3X0 U12097 ( .IN1(n9307), .IN2(n4471), .IN3(n8101), .QN(n11312) );
  NOR2X0 U12098 ( .IN1(n12027), .IN2(g2753), .QN(n12026) );
  NOR2X0 U12099 ( .IN1(n9307), .IN2(n8101), .QN(n12027) );
  NOR3X0 U12100 ( .IN1(n11427), .IN2(n10283), .IN3(n12028), .QN(g27131) );
  NOR2X0 U12101 ( .IN1(n3683), .IN2(g2147), .QN(n12028) );
  INVX0 U12102 ( .INP(n4522), .ZN(n11427) );
  NOR3X0 U12103 ( .IN1(n11429), .IN2(n10285), .IN3(n12029), .QN(g27129) );
  NOR2X0 U12104 ( .IN1(n3686), .IN2(g1453), .QN(n12029) );
  INVX0 U12105 ( .INP(n4523), .ZN(n11429) );
  NOR2X0 U12106 ( .IN1(n10287), .IN2(n12030), .QN(g27123) );
  XOR2X1 U12107 ( .IN1(n8091), .IN2(n3689), .Q(n12030) );
  NOR3X0 U12108 ( .IN1(n11432), .IN2(n10289), .IN3(n12031), .QN(g27120) );
  NOR2X0 U12109 ( .IN1(n3692), .IN2(test_so15), .QN(n12031) );
  INVX0 U12110 ( .INP(n4521), .ZN(n11432) );
  NAND2X0 U12111 ( .IN1(n12032), .IN2(n12033), .QN(g26827) );
  NAND2X0 U12112 ( .IN1(n12034), .IN2(n4606), .QN(n12033) );
  NAND2X0 U12113 ( .IN1(n4509), .IN2(g2519), .QN(n12032) );
  NAND2X0 U12114 ( .IN1(n12035), .IN2(n12036), .QN(g26826) );
  NAND2X0 U12115 ( .IN1(n12034), .IN2(g7264), .QN(n12036) );
  NAND2X0 U12116 ( .IN1(n4524), .IN2(g2516), .QN(n12035) );
  NAND2X0 U12117 ( .IN1(n12037), .IN2(n12038), .QN(g26825) );
  NAND2X0 U12118 ( .IN1(n4606), .IN2(n12039), .QN(n12038) );
  NAND2X0 U12119 ( .IN1(n4509), .IN2(g2510), .QN(n12037) );
  NAND2X0 U12120 ( .IN1(n12040), .IN2(n12041), .QN(g26824) );
  NAND2X0 U12121 ( .IN1(n12042), .IN2(n4618), .QN(n12041) );
  NAND2X0 U12122 ( .IN1(test_so59), .IN2(n4511), .QN(n12040) );
  NAND2X0 U12123 ( .IN1(n12043), .IN2(n12044), .QN(g26823) );
  NAND2X0 U12124 ( .IN1(n12034), .IN2(g5555), .QN(n12044) );
  XOR2X1 U12125 ( .IN1(n12045), .IN2(n11350), .Q(n12034) );
  NAND2X0 U12126 ( .IN1(n12046), .IN2(n11340), .QN(n12045) );
  NAND3X0 U12127 ( .IN1(n12047), .IN2(n12048), .IN3(n12049), .QN(n11340) );
  NAND2X0 U12128 ( .IN1(n7667), .IN2(n10046), .QN(n12049) );
  NAND2X0 U12129 ( .IN1(n10047), .IN2(n8122), .QN(n12048) );
  NAND2X0 U12130 ( .IN1(n7676), .IN2(n10048), .QN(n12047) );
  INVX0 U12131 ( .INP(n11341), .ZN(n12046) );
  NAND3X0 U12132 ( .IN1(n12050), .IN2(n12051), .IN3(test_so79), .QN(n11341) );
  NAND2X0 U12133 ( .IN1(n12052), .IN2(n11351), .QN(n12051) );
  NAND2X0 U12134 ( .IN1(n11350), .IN2(n11346), .QN(n12052) );
  INVX0 U12135 ( .INP(n11347), .ZN(n11350) );
  NAND2X0 U12136 ( .IN1(n11348), .IN2(n12053), .QN(n12050) );
  NAND2X0 U12137 ( .IN1(n11349), .IN2(n11347), .QN(n12053) );
  INVX0 U12138 ( .INP(n11351), .ZN(n11348) );
  NAND2X0 U12139 ( .IN1(n4516), .IN2(g2513), .QN(n12043) );
  NAND2X0 U12140 ( .IN1(n12054), .IN2(n12055), .QN(g26822) );
  NAND2X0 U12141 ( .IN1(g7264), .IN2(n12039), .QN(n12055) );
  NAND2X0 U12142 ( .IN1(n4524), .IN2(g2507), .QN(n12054) );
  NAND2X0 U12143 ( .IN1(n12056), .IN2(n12057), .QN(g26821) );
  NAND2X0 U12144 ( .IN1(n12042), .IN2(g7014), .QN(n12057) );
  NAND2X0 U12145 ( .IN1(n4525), .IN2(g1822), .QN(n12056) );
  NAND2X0 U12146 ( .IN1(n12058), .IN2(n12059), .QN(g26820) );
  NAND2X0 U12147 ( .IN1(n4618), .IN2(n12060), .QN(n12059) );
  NAND2X0 U12148 ( .IN1(n4511), .IN2(g1816), .QN(n12058) );
  NAND2X0 U12149 ( .IN1(n12061), .IN2(n12062), .QN(g26818) );
  NAND2X0 U12150 ( .IN1(n4381), .IN2(g1131), .QN(n12062) );
  NAND2X0 U12151 ( .IN1(n12063), .IN2(g1088), .QN(n12061) );
  NAND2X0 U12152 ( .IN1(n12064), .IN2(n12065), .QN(g26817) );
  NAND2X0 U12153 ( .IN1(g5555), .IN2(n12039), .QN(n12065) );
  NAND2X0 U12154 ( .IN1(n12066), .IN2(n12067), .QN(n12039) );
  NAND2X0 U12155 ( .IN1(n11351), .IN2(n8107), .QN(n12067) );
  NAND3X0 U12156 ( .IN1(n12068), .IN2(n12069), .IN3(n12070), .QN(n11351) );
  NAND2X0 U12157 ( .IN1(g5555), .IN2(g2504), .QN(n12070) );
  NAND2X0 U12158 ( .IN1(n4606), .IN2(g2510), .QN(n12069) );
  NAND2X0 U12159 ( .IN1(g7264), .IN2(g2507), .QN(n12068) );
  NAND2X0 U12160 ( .IN1(n11346), .IN2(test_so79), .QN(n12066) );
  INVX0 U12161 ( .INP(n11349), .ZN(n11346) );
  NAND2X0 U12162 ( .IN1(n10770), .IN2(n12071), .QN(n11349) );
  NAND3X0 U12163 ( .IN1(n12072), .IN2(n12073), .IN3(n12074), .QN(n12071) );
  NAND2X0 U12164 ( .IN1(n7580), .IN2(test_so73), .QN(n12074) );
  NAND2X0 U12165 ( .IN1(n7581), .IN2(g6837), .QN(n12073) );
  NAND2X0 U12166 ( .IN1(n7579), .IN2(g2241), .QN(n12072) );
  INVX0 U12167 ( .INP(n12075), .ZN(n10770) );
  NAND2X0 U12168 ( .IN1(n4516), .IN2(g2504), .QN(n12064) );
  NAND2X0 U12169 ( .IN1(n12076), .IN2(n12077), .QN(g26816) );
  NAND2X0 U12170 ( .IN1(n12042), .IN2(g5511), .QN(n12077) );
  XOR2X1 U12171 ( .IN1(n11370), .IN2(n12078), .Q(n12042) );
  NOR2X0 U12172 ( .IN1(n12079), .IN2(n11364), .QN(n12078) );
  NAND3X0 U12173 ( .IN1(n12080), .IN2(n12081), .IN3(g1690), .QN(n11364) );
  NAND2X0 U12174 ( .IN1(n12082), .IN2(n11374), .QN(n12081) );
  NAND2X0 U12175 ( .IN1(n11373), .IN2(n11369), .QN(n12082) );
  INVX0 U12176 ( .INP(n11370), .ZN(n11373) );
  NAND2X0 U12177 ( .IN1(n11371), .IN2(n12083), .QN(n12080) );
  NAND2X0 U12178 ( .IN1(n11372), .IN2(n11370), .QN(n12083) );
  INVX0 U12179 ( .INP(n11374), .ZN(n11371) );
  INVX0 U12180 ( .INP(n11363), .ZN(n12079) );
  NAND3X0 U12181 ( .IN1(n12084), .IN2(n12085), .IN3(n12086), .QN(n11363) );
  NAND2X0 U12182 ( .IN1(n7670), .IN2(n10092), .QN(n12086) );
  NAND2X0 U12183 ( .IN1(n7680), .IN2(n10093), .QN(n12085) );
  NAND2X0 U12184 ( .IN1(n7681), .IN2(n10094), .QN(n12084) );
  NAND2X0 U12185 ( .IN1(n4518), .IN2(g1819), .QN(n12076) );
  NAND2X0 U12186 ( .IN1(n12087), .IN2(n12088), .QN(g26815) );
  NAND2X0 U12187 ( .IN1(g7014), .IN2(n12060), .QN(n12088) );
  NAND2X0 U12188 ( .IN1(n4525), .IN2(g1813), .QN(n12087) );
  NAND2X0 U12189 ( .IN1(n12089), .IN2(n12090), .QN(g26814) );
  NAND2X0 U12190 ( .IN1(n4364), .IN2(g1128), .QN(n12090) );
  NAND2X0 U12191 ( .IN1(n12063), .IN2(g6712), .QN(n12089) );
  NAND2X0 U12192 ( .IN1(n12091), .IN2(n12092), .QN(g26813) );
  NAND2X0 U12193 ( .IN1(n4381), .IN2(g1122), .QN(n12092) );
  NAND2X0 U12194 ( .IN1(n12093), .IN2(g1088), .QN(n12091) );
  NAND2X0 U12195 ( .IN1(n12094), .IN2(n12095), .QN(g26812) );
  NAND2X0 U12196 ( .IN1(n12096), .IN2(n4640), .QN(n12095) );
  NAND2X0 U12197 ( .IN1(n4506), .IN2(g444), .QN(n12094) );
  NAND2X0 U12198 ( .IN1(n12097), .IN2(n12098), .QN(g26811) );
  NAND2X0 U12199 ( .IN1(g5511), .IN2(n12060), .QN(n12098) );
  NAND2X0 U12200 ( .IN1(n12099), .IN2(n12100), .QN(n12060) );
  NAND2X0 U12201 ( .IN1(n4386), .IN2(n11374), .QN(n12100) );
  NAND3X0 U12202 ( .IN1(n12101), .IN2(n12102), .IN3(n12103), .QN(n11374) );
  NAND2X0 U12203 ( .IN1(g5511), .IN2(g1810), .QN(n12103) );
  NAND2X0 U12204 ( .IN1(n4618), .IN2(g1816), .QN(n12102) );
  NAND2X0 U12205 ( .IN1(g7014), .IN2(g1813), .QN(n12101) );
  NAND2X0 U12206 ( .IN1(n11369), .IN2(g1690), .QN(n12099) );
  INVX0 U12207 ( .INP(n11372), .ZN(n11369) );
  NAND2X0 U12208 ( .IN1(n10811), .IN2(n12104), .QN(n11372) );
  NAND3X0 U12209 ( .IN1(n12105), .IN2(n12106), .IN3(n12107), .QN(n12104) );
  NAND2X0 U12210 ( .IN1(n7592), .IN2(g6782), .QN(n12107) );
  NAND2X0 U12211 ( .IN1(n7593), .IN2(g6573), .QN(n12106) );
  NAND2X0 U12212 ( .IN1(n7591), .IN2(g1547), .QN(n12105) );
  INVX0 U12213 ( .INP(n12108), .ZN(n10811) );
  NAND2X0 U12214 ( .IN1(n4518), .IN2(g1810), .QN(n12097) );
  NAND2X0 U12215 ( .IN1(n12109), .IN2(n12110), .QN(g26810) );
  NAND2X0 U12216 ( .IN1(n4363), .IN2(g1125), .QN(n12110) );
  NAND2X0 U12217 ( .IN1(n12063), .IN2(g5472), .QN(n12109) );
  XOR2X1 U12218 ( .IN1(n12111), .IN2(n11396), .Q(n12063) );
  NAND2X0 U12219 ( .IN1(n12112), .IN2(n11386), .QN(n12111) );
  NAND3X0 U12220 ( .IN1(n12113), .IN2(n12114), .IN3(n12115), .QN(n11386) );
  NAND2X0 U12221 ( .IN1(n7686), .IN2(g1088), .QN(n12115) );
  NAND2X0 U12222 ( .IN1(n7687), .IN2(g5472), .QN(n12114) );
  NAND2X0 U12223 ( .IN1(n7673), .IN2(g6712), .QN(n12113) );
  INVX0 U12224 ( .INP(n11387), .ZN(n12112) );
  NAND3X0 U12225 ( .IN1(n12116), .IN2(n12117), .IN3(g996), .QN(n11387) );
  NAND2X0 U12226 ( .IN1(n12118), .IN2(n11397), .QN(n12117) );
  NAND2X0 U12227 ( .IN1(n11396), .IN2(n11392), .QN(n12118) );
  INVX0 U12228 ( .INP(n11393), .ZN(n11396) );
  NAND2X0 U12229 ( .IN1(n11394), .IN2(n12119), .QN(n12116) );
  NAND2X0 U12230 ( .IN1(n11395), .IN2(n11393), .QN(n12119) );
  INVX0 U12231 ( .INP(n11397), .ZN(n11394) );
  NAND2X0 U12232 ( .IN1(n12120), .IN2(n12121), .QN(g26809) );
  NAND2X0 U12233 ( .IN1(n12093), .IN2(g6712), .QN(n12121) );
  NAND2X0 U12234 ( .IN1(n4364), .IN2(test_so38), .QN(n12120) );
  NAND2X0 U12235 ( .IN1(n12122), .IN2(n12123), .QN(g26808) );
  NAND2X0 U12236 ( .IN1(n12096), .IN2(g6447), .QN(n12123) );
  NAND2X0 U12237 ( .IN1(n4499), .IN2(g441), .QN(n12122) );
  NAND2X0 U12238 ( .IN1(n12124), .IN2(n12125), .QN(g26807) );
  NAND2X0 U12239 ( .IN1(n4640), .IN2(n12126), .QN(n12125) );
  NAND2X0 U12240 ( .IN1(n4506), .IN2(g435), .QN(n12124) );
  NAND2X0 U12241 ( .IN1(n12127), .IN2(n12128), .QN(g26806) );
  NAND2X0 U12242 ( .IN1(n4363), .IN2(g1116), .QN(n12128) );
  NAND2X0 U12243 ( .IN1(n12093), .IN2(g5472), .QN(n12127) );
  NAND2X0 U12244 ( .IN1(n12129), .IN2(n12130), .QN(n12093) );
  NAND2X0 U12245 ( .IN1(n4387), .IN2(n11397), .QN(n12130) );
  NAND3X0 U12246 ( .IN1(n12131), .IN2(n12132), .IN3(n12133), .QN(n11397) );
  NAND2X0 U12247 ( .IN1(g1088), .IN2(g1122), .QN(n12133) );
  NAND2X0 U12248 ( .IN1(g5472), .IN2(g1116), .QN(n12132) );
  NAND2X0 U12249 ( .IN1(test_so38), .IN2(g6712), .QN(n12131) );
  NAND2X0 U12250 ( .IN1(n11392), .IN2(g996), .QN(n12129) );
  INVX0 U12251 ( .INP(n11395), .ZN(n11392) );
  NAND2X0 U12252 ( .IN1(n10844), .IN2(n12134), .QN(n11395) );
  NAND3X0 U12253 ( .IN1(n12135), .IN2(n12136), .IN3(n12137), .QN(n12134) );
  NAND2X0 U12254 ( .IN1(n7602), .IN2(test_so31), .QN(n12137) );
  NAND2X0 U12255 ( .IN1(n7603), .IN2(g6518), .QN(n12136) );
  NAND2X0 U12256 ( .IN1(n7604), .IN2(g6368), .QN(n12135) );
  INVX0 U12257 ( .INP(n12138), .ZN(n10844) );
  NAND2X0 U12258 ( .IN1(n12139), .IN2(n12140), .QN(g26805) );
  NAND2X0 U12259 ( .IN1(n12096), .IN2(g5437), .QN(n12140) );
  XOR2X1 U12260 ( .IN1(n11411), .IN2(n12141), .Q(n12096) );
  NOR2X0 U12261 ( .IN1(n12142), .IN2(n11405), .QN(n12141) );
  NAND3X0 U12262 ( .IN1(n12143), .IN2(n12144), .IN3(g309), .QN(n11405) );
  NAND2X0 U12263 ( .IN1(n12145), .IN2(n11415), .QN(n12144) );
  NAND2X0 U12264 ( .IN1(n11414), .IN2(n11410), .QN(n12145) );
  INVX0 U12265 ( .INP(n11411), .ZN(n11414) );
  NAND2X0 U12266 ( .IN1(n11412), .IN2(n12146), .QN(n12143) );
  NAND2X0 U12267 ( .IN1(n11413), .IN2(n11411), .QN(n12146) );
  INVX0 U12268 ( .INP(n11415), .ZN(n11412) );
  INVX0 U12269 ( .INP(n11404), .ZN(n12142) );
  NAND3X0 U12270 ( .IN1(n12147), .IN2(n12148), .IN3(n12149), .QN(n11404) );
  NAND2X0 U12271 ( .IN1(n7695), .IN2(n10176), .QN(n12149) );
  NAND2X0 U12272 ( .IN1(n7694), .IN2(n10177), .QN(n12148) );
  NAND2X0 U12273 ( .IN1(n7693), .IN2(n10178), .QN(n12147) );
  NAND2X0 U12274 ( .IN1(n4520), .IN2(g438), .QN(n12139) );
  NAND2X0 U12275 ( .IN1(n12150), .IN2(n12151), .QN(g26804) );
  NAND2X0 U12276 ( .IN1(g6447), .IN2(n12126), .QN(n12151) );
  NAND2X0 U12277 ( .IN1(n4499), .IN2(g432), .QN(n12150) );
  NAND2X0 U12278 ( .IN1(n12152), .IN2(n12153), .QN(g26803) );
  NAND2X0 U12279 ( .IN1(g5437), .IN2(n12126), .QN(n12153) );
  NAND2X0 U12280 ( .IN1(n12154), .IN2(n12155), .QN(n12126) );
  NAND2X0 U12281 ( .IN1(n4388), .IN2(n11415), .QN(n12155) );
  NAND3X0 U12282 ( .IN1(n12156), .IN2(n12157), .IN3(n12158), .QN(n11415) );
  NAND2X0 U12283 ( .IN1(g5437), .IN2(g429), .QN(n12158) );
  NAND2X0 U12284 ( .IN1(n4640), .IN2(g435), .QN(n12157) );
  NAND2X0 U12285 ( .IN1(g6447), .IN2(g432), .QN(n12156) );
  NAND2X0 U12286 ( .IN1(n11410), .IN2(g309), .QN(n12154) );
  INVX0 U12287 ( .INP(n11413), .ZN(n11410) );
  NAND2X0 U12288 ( .IN1(n10871), .IN2(n12159), .QN(n11413) );
  NAND3X0 U12289 ( .IN1(n12160), .IN2(n12161), .IN3(n12162), .QN(n12159) );
  NAND2X0 U12290 ( .IN1(n7614), .IN2(g6313), .QN(n12162) );
  NAND2X0 U12291 ( .IN1(n7615), .IN2(g6231), .QN(n12161) );
  NAND2X0 U12292 ( .IN1(n7613), .IN2(g165), .QN(n12160) );
  INVX0 U12293 ( .INP(n12163), .ZN(n10871) );
  NAND2X0 U12294 ( .IN1(n4520), .IN2(g429), .QN(n12152) );
  NOR2X0 U12295 ( .IN1(n8685), .IN2(n12164), .QN(g26798) );
  XNOR2X1 U12296 ( .IN1(n4355), .IN2(n12165), .Q(n12164) );
  NAND2X0 U12297 ( .IN1(n12166), .IN2(g2900), .QN(n12165) );
  NOR2X0 U12298 ( .IN1(n11309), .IN2(n12167), .QN(g26795) );
  XOR2X1 U12299 ( .IN1(n9307), .IN2(test_so92), .Q(n12167) );
  NAND3X0 U12300 ( .IN1(g2734), .IN2(g2746), .IN3(n9309), .QN(n9307) );
  NOR2X0 U12301 ( .IN1(n9323), .IN2(n12168), .QN(g26789) );
  XOR2X1 U12302 ( .IN1(n4468), .IN2(n9324), .Q(n12168) );
  NOR3X0 U12303 ( .IN1(n4399), .IN2(n4409), .IN3(n9326), .QN(n9324) );
  INVX0 U12304 ( .INP(n12169), .ZN(n9326) );
  NOR2X0 U12305 ( .IN1(n12170), .IN2(n12171), .QN(g26786) );
  XOR2X1 U12306 ( .IN1(g3024), .IN2(n3741), .Q(n12170) );
  NOR2X0 U12307 ( .IN1(n8524), .IN2(n12172), .QN(g26781) );
  XNOR2X1 U12308 ( .IN1(n4469), .IN2(n8520), .Q(n12172) );
  NAND3X0 U12309 ( .IN1(g1346), .IN2(g1358), .IN3(n8522), .QN(n8520) );
  NOR2X0 U12310 ( .IN1(n8548), .IN2(n12173), .QN(g26776) );
  XOR2X1 U12311 ( .IN1(n8540), .IN2(test_so28), .Q(n12173) );
  NAND3X0 U12312 ( .IN1(g660), .IN2(g672), .IN3(n8542), .QN(n8540) );
  NAND2X0 U12313 ( .IN1(n12174), .IN2(n12175), .QN(g26676) );
  NAND2X0 U12314 ( .IN1(n12176), .IN2(g2479), .QN(n12175) );
  NAND2X0 U12315 ( .IN1(n9290), .IN2(n10046), .QN(n12176) );
  NAND2X0 U12316 ( .IN1(n12177), .IN2(n10046), .QN(n12174) );
  NAND2X0 U12317 ( .IN1(n12178), .IN2(n12179), .QN(g26675) );
  NAND2X0 U12318 ( .IN1(n12180), .IN2(g1783), .QN(n12179) );
  NAND2X0 U12319 ( .IN1(n9321), .IN2(n10093), .QN(n12180) );
  NAND2X0 U12320 ( .IN1(n12181), .IN2(n10093), .QN(n12178) );
  NAND2X0 U12321 ( .IN1(n12182), .IN2(n12183), .QN(g26672) );
  NAND2X0 U12322 ( .IN1(n12184), .IN2(g2478), .QN(n12183) );
  NAND2X0 U12323 ( .IN1(n9290), .IN2(n10048), .QN(n12184) );
  NAND2X0 U12324 ( .IN1(n12177), .IN2(n10048), .QN(n12182) );
  NAND2X0 U12325 ( .IN1(n12185), .IN2(n12186), .QN(g26670) );
  NAND2X0 U12326 ( .IN1(n12187), .IN2(g1785), .QN(n12186) );
  NAND2X0 U12327 ( .IN1(n9321), .IN2(n10092), .QN(n12187) );
  NAND2X0 U12328 ( .IN1(n12181), .IN2(n10092), .QN(n12185) );
  NAND2X0 U12329 ( .IN1(n12188), .IN2(n12189), .QN(g26669) );
  NAND2X0 U12330 ( .IN1(n12190), .IN2(g1089), .QN(n12189) );
  NAND2X0 U12331 ( .IN1(n9295), .IN2(g1088), .QN(n12190) );
  NAND2X0 U12332 ( .IN1(n12191), .IN2(g1088), .QN(n12188) );
  NAND2X0 U12333 ( .IN1(n12192), .IN2(n12193), .QN(g26667) );
  NAND2X0 U12334 ( .IN1(test_so60), .IN2(n12194), .QN(n12193) );
  NAND2X0 U12335 ( .IN1(n9321), .IN2(n10094), .QN(n12194) );
  NAND2X0 U12336 ( .IN1(n12181), .IN2(n10094), .QN(n12192) );
  NOR2X0 U12337 ( .IN1(n9321), .IN2(n4386), .QN(n12181) );
  NOR3X0 U12338 ( .IN1(n10465), .IN2(n4386), .IN3(n10262), .QN(n9321) );
  NAND3X0 U12339 ( .IN1(n12195), .IN2(n12196), .IN3(n12197), .QN(n10262) );
  NAND2X0 U12340 ( .IN1(n7669), .IN2(n10092), .QN(n12197) );
  NAND2X0 U12341 ( .IN1(n7679), .IN2(n10093), .QN(n12196) );
  NAND2X0 U12342 ( .IN1(n10094), .IN2(n8123), .QN(n12195) );
  NAND4X0 U12343 ( .IN1(n12198), .IN2(n12199), .IN3(n12200), .IN4(n12201), 
        .QN(n10465) );
  NOR4X0 U12344 ( .IN1(n12202), .IN2(n12203), .IN3(n12204), .IN4(n12205), .QN(
        n12201) );
  XNOR2X1 U12345 ( .IN1(n4374), .IN2(n12206), .Q(n12205) );
  NAND3X0 U12346 ( .IN1(n12207), .IN2(n12208), .IN3(n12209), .QN(n12206) );
  NAND2X0 U12347 ( .IN1(n7908), .IN2(g6782), .QN(n12209) );
  NAND2X0 U12348 ( .IN1(g6573), .IN2(n8110), .QN(n12208) );
  NAND2X0 U12349 ( .IN1(n7542), .IN2(g1547), .QN(n12207) );
  XOR2X1 U12350 ( .IN1(g1481), .IN2(n12210), .Q(n12204) );
  NAND3X0 U12351 ( .IN1(n12211), .IN2(n12212), .IN3(n12213), .QN(n12210) );
  NAND2X0 U12352 ( .IN1(n7905), .IN2(g6782), .QN(n12213) );
  NAND2X0 U12353 ( .IN1(n7906), .IN2(g6573), .QN(n12212) );
  NAND2X0 U12354 ( .IN1(n7541), .IN2(g1547), .QN(n12211) );
  XOR2X1 U12355 ( .IN1(n9660), .IN2(n12214), .Q(n12203) );
  NAND3X0 U12356 ( .IN1(n12215), .IN2(n12216), .IN3(n12217), .QN(n12214) );
  NAND2X0 U12357 ( .IN1(n7518), .IN2(g6782), .QN(n12217) );
  NAND2X0 U12358 ( .IN1(n7519), .IN2(g6573), .QN(n12216) );
  NAND2X0 U12359 ( .IN1(n7517), .IN2(g1547), .QN(n12215) );
  NAND3X0 U12360 ( .IN1(n12218), .IN2(n3070), .IN3(n12219), .QN(n12202) );
  XOR2X1 U12361 ( .IN1(n12220), .IN2(n4378), .Q(n12219) );
  NAND3X0 U12362 ( .IN1(n12221), .IN2(n12222), .IN3(n12223), .QN(n12220) );
  NAND2X0 U12363 ( .IN1(n7910), .IN2(g6782), .QN(n12223) );
  NAND2X0 U12364 ( .IN1(n7911), .IN2(g6573), .QN(n12222) );
  NAND2X0 U12365 ( .IN1(n7543), .IN2(g1547), .QN(n12221) );
  XOR2X1 U12366 ( .IN1(n12224), .IN2(n9504), .Q(n12218) );
  NAND3X0 U12367 ( .IN1(n12225), .IN2(n12226), .IN3(n12227), .QN(n12224) );
  NAND2X0 U12368 ( .IN1(n7534), .IN2(g6782), .QN(n12227) );
  NAND2X0 U12369 ( .IN1(n7535), .IN2(g6573), .QN(n12226) );
  NAND2X0 U12370 ( .IN1(n7533), .IN2(g1547), .QN(n12225) );
  NOR3X0 U12371 ( .IN1(n12228), .IN2(n12229), .IN3(n12230), .QN(n12200) );
  XOR2X1 U12372 ( .IN1(g1501), .IN2(n12231), .Q(n12230) );
  NAND3X0 U12373 ( .IN1(n12232), .IN2(n12233), .IN3(n12234), .QN(n12231) );
  NAND2X0 U12374 ( .IN1(g6782), .IN2(n8124), .QN(n12234) );
  NAND2X0 U12375 ( .IN1(n7898), .IN2(g6573), .QN(n12233) );
  NAND2X0 U12376 ( .IN1(n7537), .IN2(g1547), .QN(n12232) );
  XOR2X1 U12377 ( .IN1(g1496), .IN2(n12235), .Q(n12229) );
  NAND3X0 U12378 ( .IN1(n12236), .IN2(n12237), .IN3(n12238), .QN(n12235) );
  NAND2X0 U12379 ( .IN1(n7899), .IN2(g6782), .QN(n12238) );
  NAND2X0 U12380 ( .IN1(n7900), .IN2(g6573), .QN(n12237) );
  NAND2X0 U12381 ( .IN1(n7538), .IN2(g1547), .QN(n12236) );
  XNOR2X1 U12382 ( .IN1(n4390), .IN2(n12239), .Q(n12228) );
  NAND3X0 U12383 ( .IN1(n12240), .IN2(n12241), .IN3(n12242), .QN(n12239) );
  NAND2X0 U12384 ( .IN1(n7903), .IN2(g6782), .QN(n12242) );
  NAND2X0 U12385 ( .IN1(n7904), .IN2(g6573), .QN(n12241) );
  NAND2X0 U12386 ( .IN1(n7540), .IN2(g1547), .QN(n12240) );
  XOR2X1 U12387 ( .IN1(n12243), .IN2(n4288), .Q(n12199) );
  NAND3X0 U12388 ( .IN1(n12244), .IN2(n12245), .IN3(n12246), .QN(n12243) );
  NAND2X0 U12389 ( .IN1(n7896), .IN2(g6782), .QN(n12246) );
  NAND2X0 U12390 ( .IN1(n7897), .IN2(g6573), .QN(n12245) );
  NAND2X0 U12391 ( .IN1(n7536), .IN2(g1547), .QN(n12244) );
  XOR2X1 U12392 ( .IN1(n12247), .IN2(n4326), .Q(n12198) );
  NAND3X0 U12393 ( .IN1(n12248), .IN2(n12249), .IN3(n12250), .QN(n12247) );
  NAND2X0 U12394 ( .IN1(n7901), .IN2(g6782), .QN(n12250) );
  NAND2X0 U12395 ( .IN1(n7902), .IN2(g6573), .QN(n12249) );
  NAND2X0 U12396 ( .IN1(n7539), .IN2(g1547), .QN(n12248) );
  NAND2X0 U12397 ( .IN1(n12251), .IN2(n12252), .QN(g26665) );
  NAND2X0 U12398 ( .IN1(n12253), .IN2(g1091), .QN(n12252) );
  NAND2X0 U12399 ( .IN1(n9295), .IN2(g6712), .QN(n12253) );
  NAND2X0 U12400 ( .IN1(n12191), .IN2(g6712), .QN(n12251) );
  NAND2X0 U12401 ( .IN1(n12254), .IN2(n12255), .QN(g26664) );
  NAND2X0 U12402 ( .IN1(n12256), .IN2(g402), .QN(n12255) );
  NAND2X0 U12403 ( .IN1(n9294), .IN2(n10178), .QN(n12256) );
  NAND2X0 U12404 ( .IN1(n12257), .IN2(n10178), .QN(n12254) );
  NAND2X0 U12405 ( .IN1(n12258), .IN2(n12259), .QN(g26661) );
  NAND2X0 U12406 ( .IN1(n12260), .IN2(g1090), .QN(n12259) );
  NAND2X0 U12407 ( .IN1(n9295), .IN2(g5472), .QN(n12260) );
  NAND2X0 U12408 ( .IN1(n12191), .IN2(g5472), .QN(n12258) );
  NOR2X0 U12409 ( .IN1(n9295), .IN2(n4387), .QN(n12191) );
  NOR3X0 U12410 ( .IN1(n10555), .IN2(n4387), .IN3(n10271), .QN(n9295) );
  NAND3X0 U12411 ( .IN1(n12261), .IN2(n12262), .IN3(n12263), .QN(n10271) );
  NAND2X0 U12412 ( .IN1(n7684), .IN2(g1088), .QN(n12263) );
  NAND2X0 U12413 ( .IN1(n7685), .IN2(g5472), .QN(n12262) );
  NAND2X0 U12414 ( .IN1(n7672), .IN2(g6712), .QN(n12261) );
  NAND4X0 U12415 ( .IN1(n12264), .IN2(n12265), .IN3(n12266), .IN4(n12267), 
        .QN(n10555) );
  NOR4X0 U12416 ( .IN1(n12268), .IN2(n12269), .IN3(n12270), .IN4(n12271), .QN(
        n12267) );
  XNOR2X1 U12417 ( .IN1(n4375), .IN2(n12272), .Q(n12271) );
  NAND3X0 U12418 ( .IN1(n12273), .IN2(n12274), .IN3(n12275), .QN(n12272) );
  NAND2X0 U12419 ( .IN1(n7556), .IN2(test_so31), .QN(n12275) );
  NAND2X0 U12420 ( .IN1(n7935), .IN2(g6518), .QN(n12274) );
  NAND2X0 U12421 ( .IN1(n7939), .IN2(g6368), .QN(n12273) );
  XOR2X1 U12422 ( .IN1(g785), .IN2(n12276), .Q(n12270) );
  NAND3X0 U12423 ( .IN1(n12277), .IN2(n12278), .IN3(n12279), .QN(n12276) );
  NAND2X0 U12424 ( .IN1(n7557), .IN2(test_so31), .QN(n12279) );
  NAND2X0 U12425 ( .IN1(n7947), .IN2(g6518), .QN(n12278) );
  NAND2X0 U12426 ( .IN1(n7948), .IN2(g6368), .QN(n12277) );
  XOR2X1 U12427 ( .IN1(n10843), .IN2(n12280), .Q(n12269) );
  NAND3X0 U12428 ( .IN1(n12281), .IN2(n12282), .IN3(n12283), .QN(n12280) );
  NAND2X0 U12429 ( .IN1(n7544), .IN2(test_so31), .QN(n12283) );
  NAND2X0 U12430 ( .IN1(n7545), .IN2(g6518), .QN(n12282) );
  NAND2X0 U12431 ( .IN1(n7546), .IN2(g6368), .QN(n12281) );
  NAND3X0 U12432 ( .IN1(n12284), .IN2(n3102), .IN3(n12285), .QN(n12268) );
  XOR2X1 U12433 ( .IN1(n12286), .IN2(n4321), .Q(n12285) );
  NAND3X0 U12434 ( .IN1(n12287), .IN2(n12288), .IN3(n12289), .QN(n12286) );
  NAND2X0 U12435 ( .IN1(n7555), .IN2(test_so31), .QN(n12289) );
  NAND2X0 U12436 ( .IN1(n7933), .IN2(g6518), .QN(n12288) );
  NAND2X0 U12437 ( .IN1(n7934), .IN2(g6368), .QN(n12287) );
  XOR2X1 U12438 ( .IN1(n12290), .IN2(n10619), .Q(n12284) );
  NAND3X0 U12439 ( .IN1(n12291), .IN2(n12292), .IN3(n12293), .QN(n12290) );
  NAND2X0 U12440 ( .IN1(n7547), .IN2(test_so31), .QN(n12293) );
  NAND2X0 U12441 ( .IN1(n7548), .IN2(g6518), .QN(n12292) );
  NAND2X0 U12442 ( .IN1(n7549), .IN2(g6368), .QN(n12291) );
  NOR3X0 U12443 ( .IN1(n12294), .IN2(n12295), .IN3(n12296), .QN(n12266) );
  XOR2X1 U12444 ( .IN1(g809), .IN2(n12297), .Q(n12296) );
  NAND3X0 U12445 ( .IN1(n12298), .IN2(n12299), .IN3(n12300), .QN(n12297) );
  NAND2X0 U12446 ( .IN1(n7551), .IN2(test_so31), .QN(n12300) );
  NAND2X0 U12447 ( .IN1(n7916), .IN2(g6518), .QN(n12299) );
  NAND2X0 U12448 ( .IN1(n7917), .IN2(g6368), .QN(n12298) );
  XOR2X1 U12449 ( .IN1(g805), .IN2(n12301), .Q(n12295) );
  NAND3X0 U12450 ( .IN1(n12302), .IN2(n12303), .IN3(n12304), .QN(n12301) );
  NAND2X0 U12451 ( .IN1(n7552), .IN2(test_so31), .QN(n12304) );
  NAND2X0 U12452 ( .IN1(n7919), .IN2(g6518), .QN(n12303) );
  NAND2X0 U12453 ( .IN1(g6368), .IN2(n8125), .QN(n12302) );
  XNOR2X1 U12454 ( .IN1(n4391), .IN2(n12305), .Q(n12294) );
  NAND3X0 U12455 ( .IN1(n12306), .IN2(n12307), .IN3(n12308), .QN(n12305) );
  NAND2X0 U12456 ( .IN1(n7554), .IN2(test_so31), .QN(n12308) );
  NAND2X0 U12457 ( .IN1(n7931), .IN2(g6518), .QN(n12307) );
  NAND2X0 U12458 ( .IN1(n7932), .IN2(g6368), .QN(n12306) );
  XOR2X1 U12459 ( .IN1(n12309), .IN2(n4289), .Q(n12265) );
  NAND3X0 U12460 ( .IN1(n12310), .IN2(n12311), .IN3(n12312), .QN(n12309) );
  NAND2X0 U12461 ( .IN1(n7550), .IN2(test_so31), .QN(n12312) );
  NAND2X0 U12462 ( .IN1(n7914), .IN2(g6518), .QN(n12311) );
  NAND2X0 U12463 ( .IN1(n7915), .IN2(g6368), .QN(n12310) );
  XOR2X1 U12464 ( .IN1(n12313), .IN2(n4327), .Q(n12264) );
  NAND3X0 U12465 ( .IN1(n12314), .IN2(n12315), .IN3(n12316), .QN(n12313) );
  NAND2X0 U12466 ( .IN1(n7553), .IN2(test_so31), .QN(n12316) );
  NAND2X0 U12467 ( .IN1(n7927), .IN2(g6518), .QN(n12315) );
  NAND2X0 U12468 ( .IN1(n7928), .IN2(g6368), .QN(n12314) );
  NAND2X0 U12469 ( .IN1(n12317), .IN2(n12318), .QN(g26659) );
  NAND2X0 U12470 ( .IN1(n12319), .IN2(g404), .QN(n12318) );
  NAND2X0 U12471 ( .IN1(n9294), .IN2(n10177), .QN(n12319) );
  NAND2X0 U12472 ( .IN1(n12257), .IN2(n10177), .QN(n12317) );
  NAND2X0 U12473 ( .IN1(n12320), .IN2(n12321), .QN(g26655) );
  NAND2X0 U12474 ( .IN1(n12322), .IN2(g403), .QN(n12321) );
  NAND2X0 U12475 ( .IN1(n9294), .IN2(n10176), .QN(n12322) );
  NAND2X0 U12476 ( .IN1(n12257), .IN2(n10176), .QN(n12320) );
  NOR2X0 U12477 ( .IN1(n9294), .IN2(n4388), .QN(n12257) );
  NOR3X0 U12478 ( .IN1(n10642), .IN2(n4388), .IN3(n10282), .QN(n9294) );
  NAND3X0 U12479 ( .IN1(n12323), .IN2(n12324), .IN3(n12325), .QN(n10282) );
  NAND2X0 U12480 ( .IN1(n7692), .IN2(n10176), .QN(n12325) );
  NAND2X0 U12481 ( .IN1(n7691), .IN2(n10177), .QN(n12324) );
  NAND2X0 U12482 ( .IN1(n7690), .IN2(n10178), .QN(n12323) );
  NAND4X0 U12483 ( .IN1(n12326), .IN2(n12327), .IN3(n12328), .IN4(n12329), 
        .QN(n10642) );
  NOR4X0 U12484 ( .IN1(n12330), .IN2(n12331), .IN3(n12332), .IN4(n12333), .QN(
        n12329) );
  XNOR2X1 U12485 ( .IN1(n4376), .IN2(n12334), .Q(n12333) );
  NAND3X0 U12486 ( .IN1(n12335), .IN2(n12336), .IN3(n12337), .QN(n12334) );
  NAND2X0 U12487 ( .IN1(n7969), .IN2(g6313), .QN(n12337) );
  NAND2X0 U12488 ( .IN1(n7970), .IN2(g6231), .QN(n12336) );
  NAND2X0 U12489 ( .IN1(n7565), .IN2(g165), .QN(n12335) );
  XOR2X1 U12490 ( .IN1(g97), .IN2(n12338), .Q(n12332) );
  NAND3X0 U12491 ( .IN1(n12339), .IN2(n12340), .IN3(n12341), .QN(n12338) );
  NAND2X0 U12492 ( .IN1(n7972), .IN2(g6313), .QN(n12341) );
  NAND2X0 U12493 ( .IN1(n7973), .IN2(g6231), .QN(n12340) );
  NAND2X0 U12494 ( .IN1(n7566), .IN2(g165), .QN(n12339) );
  XOR2X1 U12495 ( .IN1(n10712), .IN2(n12342), .Q(n12331) );
  NAND3X0 U12496 ( .IN1(n12343), .IN2(n12344), .IN3(n12345), .QN(n12342) );
  NAND2X0 U12497 ( .IN1(n7559), .IN2(g6313), .QN(n12345) );
  NAND2X0 U12498 ( .IN1(g6231), .IN2(n8126), .QN(n12344) );
  NAND2X0 U12499 ( .IN1(n7558), .IN2(g165), .QN(n12343) );
  NAND3X0 U12500 ( .IN1(n12346), .IN2(n3130), .IN3(n12347), .QN(n12330) );
  XOR2X1 U12501 ( .IN1(n12348), .IN2(n4322), .Q(n12347) );
  NAND3X0 U12502 ( .IN1(n12349), .IN2(n12350), .IN3(n12351), .QN(n12348) );
  NAND2X0 U12503 ( .IN1(n7959), .IN2(g6313), .QN(n12351) );
  NAND2X0 U12504 ( .IN1(n7961), .IN2(g6231), .QN(n12350) );
  NAND2X0 U12505 ( .IN1(n7564), .IN2(g165), .QN(n12349) );
  XOR2X1 U12506 ( .IN1(n12352), .IN2(n12353), .Q(n12346) );
  NAND3X0 U12507 ( .IN1(n12354), .IN2(n12355), .IN3(n12356), .QN(n12352) );
  NAND2X0 U12508 ( .IN1(n7521), .IN2(g6313), .QN(n12356) );
  NAND2X0 U12509 ( .IN1(n7522), .IN2(g6231), .QN(n12355) );
  NAND2X0 U12510 ( .IN1(n7520), .IN2(g165), .QN(n12354) );
  NOR3X0 U12511 ( .IN1(n12357), .IN2(n12358), .IN3(n12359), .QN(n12328) );
  XNOR2X1 U12512 ( .IN1(n4569), .IN2(n12360), .Q(n12359) );
  NAND3X0 U12513 ( .IN1(n12361), .IN2(n12362), .IN3(n12363), .QN(n12360) );
  NAND2X0 U12514 ( .IN1(n7951), .IN2(g6313), .QN(n12363) );
  NAND2X0 U12515 ( .IN1(n7952), .IN2(g6231), .QN(n12362) );
  NAND2X0 U12516 ( .IN1(n7561), .IN2(g165), .QN(n12361) );
  XNOR2X1 U12517 ( .IN1(n4561), .IN2(n12364), .Q(n12358) );
  NAND3X0 U12518 ( .IN1(n12365), .IN2(n12366), .IN3(n12367), .QN(n12364) );
  NAND2X0 U12519 ( .IN1(n7953), .IN2(g6313), .QN(n12367) );
  NAND2X0 U12520 ( .IN1(n7954), .IN2(g6231), .QN(n12366) );
  NAND2X0 U12521 ( .IN1(n7562), .IN2(g165), .QN(n12365) );
  XNOR2X1 U12522 ( .IN1(n4392), .IN2(n12368), .Q(n12357) );
  NAND3X0 U12523 ( .IN1(n12369), .IN2(n12370), .IN3(n12371), .QN(n12368) );
  NAND2X0 U12524 ( .IN1(n7957), .IN2(g6313), .QN(n12371) );
  NAND2X0 U12525 ( .IN1(n7958), .IN2(g6231), .QN(n12370) );
  NAND2X0 U12526 ( .IN1(g165), .IN2(n8127), .QN(n12369) );
  XOR2X1 U12527 ( .IN1(n12372), .IN2(n4290), .Q(n12327) );
  NAND3X0 U12528 ( .IN1(n12373), .IN2(n12374), .IN3(n12375), .QN(n12372) );
  NAND2X0 U12529 ( .IN1(n7949), .IN2(g6313), .QN(n12375) );
  NAND2X0 U12530 ( .IN1(n7950), .IN2(g6231), .QN(n12374) );
  NAND2X0 U12531 ( .IN1(n7560), .IN2(g165), .QN(n12373) );
  XOR2X1 U12532 ( .IN1(n12376), .IN2(n4328), .Q(n12326) );
  NAND3X0 U12533 ( .IN1(n12377), .IN2(n12378), .IN3(n12379), .QN(n12376) );
  NAND2X0 U12534 ( .IN1(n7955), .IN2(g6313), .QN(n12379) );
  NAND2X0 U12535 ( .IN1(n7956), .IN2(g6231), .QN(n12378) );
  NAND2X0 U12536 ( .IN1(n7563), .IN2(g165), .QN(n12377) );
  NAND2X0 U12537 ( .IN1(n12380), .IN2(n12381), .QN(g26616) );
  NAND2X0 U12538 ( .IN1(n4299), .IN2(g2571), .QN(n12381) );
  NAND2X0 U12539 ( .IN1(n12382), .IN2(g2624), .QN(n12380) );
  NAND2X0 U12540 ( .IN1(n12383), .IN2(n12384), .QN(g26596) );
  NAND2X0 U12541 ( .IN1(n4370), .IN2(g2568), .QN(n12384) );
  NAND2X0 U12542 ( .IN1(n12382), .IN2(g7390), .QN(n12383) );
  NAND2X0 U12543 ( .IN1(n12385), .IN2(n12386), .QN(g26592) );
  NAND2X0 U12544 ( .IN1(n4366), .IN2(g1877), .QN(n12386) );
  NAND2X0 U12545 ( .IN1(n12387), .IN2(g1930), .QN(n12385) );
  NAND2X0 U12546 ( .IN1(n12388), .IN2(n12389), .QN(g26575) );
  NAND2X0 U12547 ( .IN1(n4314), .IN2(g2565), .QN(n12389) );
  NAND2X0 U12548 ( .IN1(n12382), .IN2(n10186), .QN(n12388) );
  NOR3X0 U12549 ( .IN1(n8887), .IN2(n4303), .IN3(n12390), .QN(n12382) );
  NAND2X0 U12550 ( .IN1(n12391), .IN2(n12392), .QN(g26573) );
  NAND2X0 U12551 ( .IN1(n4315), .IN2(g1874), .QN(n12392) );
  NAND2X0 U12552 ( .IN1(n12387), .IN2(g7194), .QN(n12391) );
  NAND2X0 U12553 ( .IN1(n12393), .IN2(n12394), .QN(g26569) );
  NAND2X0 U12554 ( .IN1(n4300), .IN2(g1183), .QN(n12394) );
  NAND2X0 U12555 ( .IN1(n12395), .IN2(g1236), .QN(n12393) );
  NAND2X0 U12556 ( .IN1(n12396), .IN2(n12397), .QN(g26559) );
  NAND2X0 U12557 ( .IN1(n12387), .IN2(n10234), .QN(n12397) );
  NOR3X0 U12558 ( .IN1(n9011), .IN2(n4297), .IN3(n12398), .QN(n12387) );
  NAND2X0 U12559 ( .IN1(test_so68), .IN2(n4296), .QN(n12396) );
  NAND2X0 U12560 ( .IN1(n12399), .IN2(n12400), .QN(g26557) );
  NAND2X0 U12561 ( .IN1(n4316), .IN2(g1180), .QN(n12400) );
  NAND2X0 U12562 ( .IN1(n12395), .IN2(g6944), .QN(n12399) );
  NAND2X0 U12563 ( .IN1(n12401), .IN2(n12402), .QN(g26553) );
  NAND2X0 U12564 ( .IN1(n4313), .IN2(g496), .QN(n12402) );
  NAND2X0 U12565 ( .IN1(n12403), .IN2(g550), .QN(n12401) );
  NAND2X0 U12566 ( .IN1(n12404), .IN2(n12405), .QN(g26547) );
  NAND2X0 U12567 ( .IN1(n12395), .IN2(n11110), .QN(n12405) );
  NOR3X0 U12568 ( .IN1(n9117), .IN2(n4304), .IN3(n12406), .QN(n12395) );
  NAND2X0 U12569 ( .IN1(test_so47), .IN2(n4371), .QN(n12404) );
  NAND2X0 U12570 ( .IN1(n12407), .IN2(n12408), .QN(g26545) );
  NAND2X0 U12571 ( .IN1(n4372), .IN2(g493), .QN(n12408) );
  NAND2X0 U12572 ( .IN1(n12403), .IN2(g6642), .QN(n12407) );
  NAND2X0 U12573 ( .IN1(n12409), .IN2(n12410), .QN(g26541) );
  NAND2X0 U12574 ( .IN1(n4298), .IN2(g490), .QN(n12410) );
  NAND2X0 U12575 ( .IN1(n12403), .IN2(n11213), .QN(n12409) );
  NOR3X0 U12576 ( .IN1(n8108), .IN2(n8764), .IN3(n12411), .QN(n12403) );
  NOR2X0 U12577 ( .IN1(n10283), .IN2(n12412), .QN(g26532) );
  XOR2X1 U12578 ( .IN1(n12413), .IN2(n7701), .Q(n12412) );
  NOR2X0 U12579 ( .IN1(n10285), .IN2(n12414), .QN(g26531) );
  XOR2X1 U12580 ( .IN1(n12415), .IN2(n7705), .Q(n12414) );
  NOR2X0 U12581 ( .IN1(n10287), .IN2(n12416), .QN(g26530) );
  XNOR2X1 U12582 ( .IN1(n7709), .IN2(n3690), .Q(n12416) );
  NAND2X0 U12583 ( .IN1(n3893), .IN2(g776), .QN(n3690) );
  NOR2X0 U12584 ( .IN1(n10289), .IN2(n12417), .QN(g26529) );
  XOR2X1 U12585 ( .IN1(n12418), .IN2(n7713), .Q(n12417) );
  NAND4X0 U12586 ( .IN1(n3700), .IN2(n12419), .IN3(n12420), .IN4(n12421), .QN(
        g26149) );
  NOR4X0 U12587 ( .IN1(n12422), .IN2(n12423), .IN3(n12424), .IN4(n12425), .QN(
        n12421) );
  NOR2X0 U12588 ( .IN1(n4441), .IN2(n12426), .QN(n12425) );
  NOR2X0 U12589 ( .IN1(n4338), .IN2(n12427), .QN(n12424) );
  NOR2X0 U12590 ( .IN1(n11451), .IN2(DFF_156_n1), .QN(n12423) );
  NAND3X0 U12591 ( .IN1(n12428), .IN2(n12429), .IN3(n12430), .QN(n12422) );
  NAND2X0 U12592 ( .IN1(n3936), .IN2(n12431), .QN(n12430) );
  NAND4X0 U12593 ( .IN1(n12432), .IN2(n12433), .IN3(n12434), .IN4(n12435), 
        .QN(n12431) );
  NAND2X0 U12594 ( .IN1(n12436), .IN2(g3088), .QN(n12435) );
  NAND2X0 U12595 ( .IN1(n12437), .IN2(g3164), .QN(n12434) );
  NAND2X0 U12596 ( .IN1(n12438), .IN2(g3158), .QN(n12433) );
  NAND2X0 U12597 ( .IN1(n12439), .IN2(g3182), .QN(n12432) );
  NAND2X0 U12598 ( .IN1(n12440), .IN2(g3167), .QN(n12429) );
  NAND2X0 U12599 ( .IN1(n3939), .IN2(n12441), .QN(n12428) );
  NAND3X0 U12600 ( .IN1(n12442), .IN2(n12443), .IN3(n12444), .QN(n12441) );
  NAND2X0 U12601 ( .IN1(n3940), .IN2(g3185), .QN(n12444) );
  NAND2X0 U12602 ( .IN1(test_so8), .IN2(n12445), .QN(n12443) );
  NAND2X0 U12603 ( .IN1(n12446), .IN2(g3155), .QN(n12442) );
  NOR3X0 U12604 ( .IN1(n12447), .IN2(n12448), .IN3(n12449), .QN(n12420) );
  NOR2X0 U12605 ( .IN1(n4444), .IN2(n12450), .QN(n12449) );
  NOR2X0 U12606 ( .IN1(n4450), .IN2(n12451), .QN(n12448) );
  NOR2X0 U12607 ( .IN1(n12452), .IN2(DFF_149_n1), .QN(n12447) );
  NAND2X0 U12608 ( .IN1(n11452), .IN2(n8086), .QN(n12419) );
  NAND4X0 U12609 ( .IN1(n12453), .IN2(n3700), .IN3(n12454), .IN4(n12455), .QN(
        g26135) );
  NOR4X0 U12610 ( .IN1(n12456), .IN2(n12457), .IN3(n12458), .IN4(n12459), .QN(
        n12455) );
  NOR2X0 U12611 ( .IN1(n4447), .IN2(n12427), .QN(n12459) );
  NOR2X0 U12612 ( .IN1(n12460), .IN2(n12461), .QN(n12458) );
  INVX0 U12613 ( .INP(n3936), .ZN(n12461) );
  NOR4X0 U12614 ( .IN1(n12462), .IN2(n12463), .IN3(n12464), .IN4(n12465), .QN(
        n12460) );
  NOR2X0 U12615 ( .IN1(n4438), .IN2(n11442), .QN(n12465) );
  INVX0 U12616 ( .INP(n12466), .ZN(n12464) );
  NAND2X0 U12617 ( .IN1(g3098), .IN2(n12438), .QN(n12466) );
  NOR2X0 U12618 ( .IN1(n4342), .IN2(n12467), .QN(n12463) );
  INVX0 U12619 ( .INP(n12437), .ZN(n12467) );
  NOR2X0 U12620 ( .IN1(n4334), .IN2(n12468), .QN(n12462) );
  INVX0 U12621 ( .INP(n12436), .ZN(n12468) );
  NOR2X0 U12622 ( .IN1(n4343), .IN2(n12426), .QN(n12457) );
  NAND4X0 U12623 ( .IN1(n12469), .IN2(n12470), .IN3(n12471), .IN4(n12472), 
        .QN(n12456) );
  NAND2X0 U12624 ( .IN1(test_so10), .IN2(n12473), .QN(n12472) );
  NAND2X0 U12625 ( .IN1(test_so7), .IN2(n12440), .QN(n12471) );
  NAND2X0 U12626 ( .IN1(n11436), .IN2(n12474), .QN(n12470) );
  INVX0 U12627 ( .INP(n12475), .ZN(n11436) );
  NAND2X0 U12628 ( .IN1(n3939), .IN2(n12476), .QN(n12469) );
  NAND3X0 U12629 ( .IN1(n12477), .IN2(n12478), .IN3(n12479), .QN(n12476) );
  NAND2X0 U12630 ( .IN1(n3940), .IN2(g3107), .QN(n12479) );
  NAND2X0 U12631 ( .IN1(n12445), .IN2(g3105), .QN(n12478) );
  NAND2X0 U12632 ( .IN1(n12446), .IN2(g3097), .QN(n12477) );
  NOR3X0 U12633 ( .IN1(n12480), .IN2(n12481), .IN3(n12482), .QN(n12454) );
  NOR2X0 U12634 ( .IN1(n4452), .IN2(n12451), .QN(n12482) );
  NOR2X0 U12635 ( .IN1(n11451), .IN2(DFF_155_n1), .QN(n12481) );
  NOR2X0 U12636 ( .IN1(n4443), .IN2(n12450), .QN(n12480) );
  NOR2X0 U12637 ( .IN1(n12483), .IN2(n12484), .QN(n12453) );
  NOR2X0 U12638 ( .IN1(n12485), .IN2(g3128), .QN(n12484) );
  NOR2X0 U12639 ( .IN1(n14384), .IN2(n12452), .QN(n12483) );
  NAND4X0 U12640 ( .IN1(n12486), .IN2(n3700), .IN3(n12487), .IN4(n12488), .QN(
        g26104) );
  NOR4X0 U12641 ( .IN1(n12489), .IN2(n12490), .IN3(n12491), .IN4(n12492), .QN(
        n12488) );
  NOR2X0 U12642 ( .IN1(n4448), .IN2(n12427), .QN(n12492) );
  NAND3X0 U12643 ( .IN1(n12493), .IN2(n4406), .IN3(n3933), .QN(n12427) );
  NOR2X0 U12644 ( .IN1(n11449), .IN2(n12475), .QN(n12491) );
  NAND2X0 U12645 ( .IN1(n12446), .IN2(n3705), .QN(n12475) );
  INVX0 U12646 ( .INP(n12494), .ZN(n11449) );
  NOR2X0 U12647 ( .IN1(n4344), .IN2(n12426), .QN(n12490) );
  NAND2X0 U12648 ( .IN1(n12495), .IN2(n4329), .QN(n12426) );
  NAND4X0 U12649 ( .IN1(n12496), .IN2(n12497), .IN3(n12498), .IN4(n12499), 
        .QN(n12489) );
  NAND2X0 U12650 ( .IN1(n12473), .IN2(g3142), .QN(n12499) );
  INVX0 U12651 ( .INP(n11440), .ZN(n12473) );
  NAND3X0 U12652 ( .IN1(n3940), .IN2(g3204), .IN3(n4073), .QN(n11440) );
  NAND2X0 U12653 ( .IN1(n12440), .IN2(g3086), .QN(n12498) );
  NOR2X0 U12654 ( .IN1(n11444), .IN2(n12500), .QN(n12440) );
  NAND2X0 U12655 ( .IN1(n3939), .IN2(n12501), .QN(n12497) );
  NAND3X0 U12656 ( .IN1(n12502), .IN2(n12503), .IN3(n12504), .QN(n12501) );
  NAND2X0 U12657 ( .IN1(n3940), .IN2(g3095), .QN(n12504) );
  NAND2X0 U12658 ( .IN1(n12445), .IN2(g3093), .QN(n12503) );
  NAND2X0 U12659 ( .IN1(test_so6), .IN2(n12446), .QN(n12502) );
  NAND2X0 U12660 ( .IN1(n3936), .IN2(n12505), .QN(n12496) );
  NAND4X0 U12661 ( .IN1(n12506), .IN2(n12507), .IN3(n12508), .IN4(n12509), 
        .QN(n12505) );
  NAND2X0 U12662 ( .IN1(n12436), .IN2(g3096), .QN(n12509) );
  NOR2X0 U12663 ( .IN1(n4329), .IN2(n4406), .QN(n12436) );
  NAND2X0 U12664 ( .IN1(n12437), .IN2(g3085), .QN(n12508) );
  NOR2X0 U12665 ( .IN1(g3201), .IN2(n4329), .QN(n12437) );
  NAND2X0 U12666 ( .IN1(n12438), .IN2(g3211), .QN(n12507) );
  NAND2X0 U12667 ( .IN1(n12439), .IN2(g3094), .QN(n12506) );
  NOR3X0 U12668 ( .IN1(n12510), .IN2(n12511), .IN3(n12512), .QN(n12487) );
  NOR2X0 U12669 ( .IN1(n4451), .IN2(n12451), .QN(n12512) );
  NAND2X0 U12670 ( .IN1(n12495), .IN2(g3207), .QN(n12451) );
  NOR3X0 U12671 ( .IN1(g3201), .IN2(n4405), .IN3(n11444), .QN(n12495) );
  INVX0 U12672 ( .INP(n12493), .ZN(n11444) );
  NOR2X0 U12673 ( .IN1(n9162), .IN2(n8036), .QN(n12493) );
  NAND2X0 U12674 ( .IN1(n285), .IN2(g3197), .QN(n9162) );
  INVX0 U12675 ( .INP(n12513), .ZN(n285) );
  NAND3X0 U12676 ( .IN1(DFF_132_n1), .IN2(DFF_131_n1), .IN3(DFF_134_n1), .QN(
        n12513) );
  NOR2X0 U12677 ( .IN1(n14386), .IN2(n11451), .QN(n12511) );
  NAND3X0 U12678 ( .IN1(n4073), .IN2(g3204), .IN3(n12445), .QN(n11451) );
  INVX0 U12679 ( .INP(n11447), .ZN(n12445) );
  NAND2X0 U12680 ( .IN1(n12439), .IN2(n4405), .QN(n11447) );
  INVX0 U12681 ( .INP(n11442), .ZN(n12439) );
  NAND2X0 U12682 ( .IN1(n4329), .IN2(g3201), .QN(n11442) );
  NOR2X0 U12683 ( .IN1(n4445), .IN2(n12450), .QN(n12510) );
  NAND3X0 U12684 ( .IN1(n3939), .IN2(n4406), .IN3(n3933), .QN(n12450) );
  INVX0 U12685 ( .INP(n12514), .ZN(n3933) );
  NAND2X0 U12686 ( .IN1(n4405), .IN2(g3207), .QN(n12514) );
  NOR2X0 U12687 ( .IN1(n12515), .IN2(n12516), .QN(n12486) );
  NOR2X0 U12688 ( .IN1(n12485), .IN2(DFF_140_n1), .QN(n12516) );
  NOR2X0 U12689 ( .IN1(n14382), .IN2(n12452), .QN(n12515) );
  NAND2X0 U12690 ( .IN1(n8739), .IN2(n12517), .QN(g26048) );
  NAND2X0 U12691 ( .IN1(n12518), .IN2(n9300), .QN(n12517) );
  XOR2X1 U12692 ( .IN1(n7909), .IN2(n9303), .Q(n12518) );
  NOR2X0 U12693 ( .IN1(n8685), .IN2(n12519), .QN(g26037) );
  XOR2X1 U12694 ( .IN1(n4291), .IN2(n12166), .Q(n12519) );
  NOR2X0 U12695 ( .IN1(n12520), .IN2(n12171), .QN(g26031) );
  XOR2X1 U12696 ( .IN1(test_so98), .IN2(n3742), .Q(n12520) );
  NAND2X0 U12697 ( .IN1(n4065), .IN2(g3013), .QN(n3742) );
  NAND2X0 U12698 ( .IN1(n12521), .IN2(n12522), .QN(g26025) );
  NAND2X0 U12699 ( .IN1(test_so82), .IN2(n12523), .QN(n12522) );
  NAND2X0 U12700 ( .IN1(n9290), .IN2(n10047), .QN(n12523) );
  NAND2X0 U12701 ( .IN1(n12177), .IN2(n10047), .QN(n12521) );
  NOR2X0 U12702 ( .IN1(n8107), .IN2(n9290), .QN(n12177) );
  NOR3X0 U12703 ( .IN1(n8107), .IN2(n10413), .IN3(n10250), .QN(n9290) );
  NAND3X0 U12704 ( .IN1(n12524), .IN2(n12525), .IN3(n12526), .QN(n10250) );
  NAND2X0 U12705 ( .IN1(n7666), .IN2(n10046), .QN(n12526) );
  NAND2X0 U12706 ( .IN1(n10047), .IN2(n8128), .QN(n12525) );
  NAND2X0 U12707 ( .IN1(n7675), .IN2(n10048), .QN(n12524) );
  NAND4X0 U12708 ( .IN1(n12527), .IN2(n12528), .IN3(n12529), .IN4(n12530), 
        .QN(n10413) );
  NOR4X0 U12709 ( .IN1(n12531), .IN2(n12532), .IN3(n12533), .IN4(n12534), .QN(
        n12530) );
  XOR2X1 U12710 ( .IN1(g2170), .IN2(n12535), .Q(n12534) );
  NAND3X0 U12711 ( .IN1(n12536), .IN2(n12537), .IN3(n12538), .QN(n12535) );
  NAND2X0 U12712 ( .IN1(n7892), .IN2(test_so73), .QN(n12538) );
  NAND2X0 U12713 ( .IN1(n7893), .IN2(g6837), .QN(n12537) );
  NAND2X0 U12714 ( .IN1(n7531), .IN2(g2241), .QN(n12536) );
  XOR2X1 U12715 ( .IN1(g2165), .IN2(n12539), .Q(n12533) );
  NAND3X0 U12716 ( .IN1(n12540), .IN2(n12541), .IN3(n12542), .QN(n12539) );
  NAND2X0 U12717 ( .IN1(n7894), .IN2(test_so73), .QN(n12542) );
  NAND2X0 U12718 ( .IN1(n7895), .IN2(g6837), .QN(n12541) );
  NAND2X0 U12719 ( .IN1(n7532), .IN2(g2241), .QN(n12540) );
  XOR2X1 U12720 ( .IN1(n10769), .IN2(n12543), .Q(n12532) );
  NAND3X0 U12721 ( .IN1(n12544), .IN2(n12545), .IN3(n12546), .QN(n12543) );
  NAND2X0 U12722 ( .IN1(test_so73), .IN2(n8129), .QN(n12546) );
  NAND2X0 U12723 ( .IN1(n7524), .IN2(g6837), .QN(n12545) );
  NAND2X0 U12724 ( .IN1(n7523), .IN2(g2241), .QN(n12544) );
  NAND3X0 U12725 ( .IN1(n12547), .IN2(n3038), .IN3(n12548), .QN(n12531) );
  XOR2X1 U12726 ( .IN1(n12549), .IN2(n4319), .Q(n12548) );
  NAND3X0 U12727 ( .IN1(n12550), .IN2(n12551), .IN3(n12552), .QN(n12549) );
  NAND2X0 U12728 ( .IN1(n7890), .IN2(test_so73), .QN(n12552) );
  NAND2X0 U12729 ( .IN1(n7891), .IN2(g6837), .QN(n12551) );
  NAND2X0 U12730 ( .IN1(n7530), .IN2(g2241), .QN(n12550) );
  XOR2X1 U12731 ( .IN1(n12553), .IN2(n10446), .Q(n12547) );
  NAND3X0 U12732 ( .IN1(n12554), .IN2(n12555), .IN3(n12556), .QN(n12553) );
  NAND2X0 U12733 ( .IN1(n7515), .IN2(test_so73), .QN(n12556) );
  NAND2X0 U12734 ( .IN1(n7516), .IN2(g6837), .QN(n12555) );
  NAND2X0 U12735 ( .IN1(n7514), .IN2(g2241), .QN(n12554) );
  NOR3X0 U12736 ( .IN1(n12557), .IN2(n12558), .IN3(n12559), .QN(n12529) );
  XOR2X1 U12737 ( .IN1(g2195), .IN2(n12560), .Q(n12559) );
  NAND3X0 U12738 ( .IN1(n12561), .IN2(n12562), .IN3(n12563), .QN(n12560) );
  NAND2X0 U12739 ( .IN1(n7883), .IN2(test_so73), .QN(n12563) );
  NAND2X0 U12740 ( .IN1(n7884), .IN2(g6837), .QN(n12562) );
  NAND2X0 U12741 ( .IN1(n7526), .IN2(g2241), .QN(n12561) );
  XOR2X1 U12742 ( .IN1(g2190), .IN2(n12564), .Q(n12558) );
  NAND3X0 U12743 ( .IN1(n12565), .IN2(n12566), .IN3(n12567), .QN(n12564) );
  NAND2X0 U12744 ( .IN1(n7885), .IN2(test_so73), .QN(n12567) );
  NAND2X0 U12745 ( .IN1(n7886), .IN2(g6837), .QN(n12566) );
  NAND2X0 U12746 ( .IN1(n7527), .IN2(g2241), .QN(n12565) );
  XOR2X1 U12747 ( .IN1(g2180), .IN2(n12568), .Q(n12557) );
  NAND3X0 U12748 ( .IN1(n12569), .IN2(n12570), .IN3(n12571), .QN(n12568) );
  NAND2X0 U12749 ( .IN1(n7888), .IN2(test_so73), .QN(n12571) );
  NAND2X0 U12750 ( .IN1(n7889), .IN2(g6837), .QN(n12570) );
  NAND2X0 U12751 ( .IN1(n7529), .IN2(g2241), .QN(n12569) );
  XOR2X1 U12752 ( .IN1(n12572), .IN2(n4287), .Q(n12528) );
  NAND3X0 U12753 ( .IN1(n12573), .IN2(n12574), .IN3(n12575), .QN(n12572) );
  NAND2X0 U12754 ( .IN1(n7881), .IN2(test_so73), .QN(n12575) );
  NAND2X0 U12755 ( .IN1(n7882), .IN2(g6837), .QN(n12574) );
  NAND2X0 U12756 ( .IN1(n7525), .IN2(g2241), .QN(n12573) );
  XOR2X1 U12757 ( .IN1(n12576), .IN2(n4325), .Q(n12527) );
  NAND3X0 U12758 ( .IN1(n12577), .IN2(n12578), .IN3(n12579), .QN(n12576) );
  NAND2X0 U12759 ( .IN1(test_so73), .IN2(n8130), .QN(n12579) );
  NAND2X0 U12760 ( .IN1(n7887), .IN2(g6837), .QN(n12578) );
  NAND2X0 U12761 ( .IN1(n7528), .IN2(g2241), .QN(n12577) );
  NOR3X0 U12762 ( .IN1(n12413), .IN2(n10283), .IN3(n12580), .QN(g25940) );
  NOR2X0 U12763 ( .IN1(n3887), .IN2(test_so78), .QN(n12580) );
  INVX0 U12764 ( .INP(n4526), .ZN(n12413) );
  NOR3X0 U12765 ( .IN1(n12415), .IN2(n10285), .IN3(n12581), .QN(g25938) );
  NOR2X0 U12766 ( .IN1(n3890), .IN2(g1462), .QN(n12581) );
  INVX0 U12767 ( .INP(n4527), .ZN(n12415) );
  NOR2X0 U12768 ( .IN1(n10287), .IN2(n12582), .QN(g25935) );
  XOR2X1 U12769 ( .IN1(n8085), .IN2(n3893), .Q(n12582) );
  NOR3X0 U12770 ( .IN1(n12418), .IN2(n10289), .IN3(n12583), .QN(g25932) );
  NOR2X0 U12771 ( .IN1(n3896), .IN2(g88), .QN(n12583) );
  INVX0 U12772 ( .INP(n4528), .ZN(n12418) );
  NAND2X0 U12773 ( .IN1(n12584), .IN2(n12585), .QN(g25489) );
  NAND2X0 U12774 ( .IN1(n12586), .IN2(n8112), .QN(n12585) );
  NAND2X0 U12775 ( .IN1(n12587), .IN2(n12588), .QN(n12586) );
  NAND2X0 U12776 ( .IN1(n4424), .IN2(n12589), .QN(n12588) );
  NAND2X0 U12777 ( .IN1(n11448), .IN2(g3142), .QN(n12589) );
  INVX0 U12778 ( .INP(n12474), .ZN(n11448) );
  NAND2X0 U12779 ( .IN1(n7444), .IN2(n7443), .QN(n12474) );
  NAND2X0 U12780 ( .IN1(n4301), .IN2(n12494), .QN(n12587) );
  NAND2X0 U12781 ( .IN1(DFF_15_n1), .IN2(DFF_16_n1), .QN(n12494) );
  NAND4X0 U12782 ( .IN1(g3151), .IN2(g3097), .IN3(g3142), .IN4(test_so10), 
        .QN(n12584) );
  NAND2X0 U12783 ( .IN1(n12590), .IN2(n12591), .QN(g25452) );
  NAND2X0 U12784 ( .IN1(n4494), .IN2(g3099), .QN(n12591) );
  NAND2X0 U12785 ( .IN1(g21851), .IN2(g3109), .QN(n12590) );
  NAND2X0 U12786 ( .IN1(n12592), .IN2(n12593), .QN(g25451) );
  NAND2X0 U12787 ( .IN1(n4383), .IN2(g3098), .QN(n12593) );
  NAND2X0 U12788 ( .IN1(g21851), .IN2(g8030), .QN(n12592) );
  NAND2X0 U12789 ( .IN1(n12594), .IN2(n12595), .QN(g25450) );
  NAND2X0 U12790 ( .IN1(n4382), .IN2(g3097), .QN(n12595) );
  NAND2X0 U12791 ( .IN1(g21851), .IN2(g8106), .QN(n12594) );
  NAND3X0 U12792 ( .IN1(n12596), .IN2(n12597), .IN3(n3700), .QN(g25442) );
  NAND2X0 U12793 ( .IN1(n12598), .IN2(g3111), .QN(n12597) );
  NAND2X0 U12794 ( .IN1(n11452), .IN2(g3124), .QN(n12596) );
  NAND3X0 U12795 ( .IN1(n12599), .IN2(n12600), .IN3(n3700), .QN(g25435) );
  NAND2X0 U12796 ( .IN1(n12598), .IN2(g3110), .QN(n12600) );
  NAND2X0 U12797 ( .IN1(n11452), .IN2(DFF_144_n1), .QN(n12599) );
  NAND3X0 U12798 ( .IN1(n12601), .IN2(n12602), .IN3(n3700), .QN(g25420) );
  NAND2X0 U12799 ( .IN1(n12598), .IN2(g3112), .QN(n12602) );
  INVX0 U12800 ( .INP(n12452), .ZN(n12598) );
  NAND3X0 U12801 ( .IN1(n12446), .IN2(g3204), .IN3(n4073), .QN(n12452) );
  INVX0 U12802 ( .INP(n12500), .ZN(n12446) );
  NAND2X0 U12803 ( .IN1(n12438), .IN2(n4405), .QN(n12500) );
  NOR2X0 U12804 ( .IN1(g3201), .IN2(g3207), .QN(n12438) );
  NAND2X0 U12805 ( .IN1(test_so9), .IN2(n11452), .QN(n12601) );
  NAND2X0 U12806 ( .IN1(n12603), .IN2(n12604), .QN(g25288) );
  NAND2X0 U12807 ( .IN1(n12605), .IN2(g2808), .QN(n12604) );
  NAND2X0 U12808 ( .IN1(n12606), .IN2(n12607), .QN(n12603) );
  NAND2X0 U12809 ( .IN1(n12608), .IN2(n12609), .QN(g25280) );
  NAND2X0 U12810 ( .IN1(n12610), .IN2(g2810), .QN(n12609) );
  NAND2X0 U12811 ( .IN1(n12611), .IN2(n12606), .QN(n12608) );
  NAND2X0 U12812 ( .IN1(n12612), .IN2(n12613), .QN(g25279) );
  NAND2X0 U12813 ( .IN1(n12614), .IN2(g2114), .QN(n12613) );
  NAND2X0 U12814 ( .IN1(n12615), .IN2(n12616), .QN(n12612) );
  NAND2X0 U12815 ( .IN1(n12617), .IN2(n12618), .QN(g25272) );
  NAND2X0 U12816 ( .IN1(n12619), .IN2(g2809), .QN(n12618) );
  NAND2X0 U12817 ( .IN1(n12620), .IN2(n12606), .QN(n12617) );
  INVX0 U12818 ( .INP(n12621), .ZN(n12606) );
  NAND4X0 U12819 ( .IN1(n9260), .IN2(n12622), .IN3(n12623), .IN4(n12624), .QN(
        n12621) );
  NAND2X0 U12820 ( .IN1(n8042), .IN2(g7425), .QN(n12624) );
  NOR2X0 U12821 ( .IN1(n12625), .IN2(n12626), .QN(n12623) );
  NOR2X0 U12822 ( .IN1(n4292), .IN2(g2802), .QN(n12626) );
  NOR4X0 U12823 ( .IN1(n12627), .IN2(n12628), .IN3(n12629), .IN4(n12630), .QN(
        n12625) );
  XNOR2X1 U12824 ( .IN1(n4419), .IN2(n8911), .Q(n12630) );
  NAND3X0 U12825 ( .IN1(n12631), .IN2(n12632), .IN3(n12633), .QN(n8911) );
  NAND2X0 U12826 ( .IN1(n7779), .IN2(g7487), .QN(n12633) );
  NAND2X0 U12827 ( .IN1(n7844), .IN2(g2703), .QN(n12632) );
  NAND2X0 U12828 ( .IN1(n7780), .IN2(g7425), .QN(n12631) );
  XOR2X1 U12829 ( .IN1(n4471), .IN2(n8875), .Q(n12629) );
  INVX0 U12830 ( .INP(n8878), .ZN(n8875) );
  NAND3X0 U12831 ( .IN1(n12634), .IN2(n12635), .IN3(n12636), .QN(n8878) );
  NAND2X0 U12832 ( .IN1(n7769), .IN2(g7487), .QN(n12636) );
  NAND2X0 U12833 ( .IN1(n7840), .IN2(g2703), .QN(n12635) );
  NAND2X0 U12834 ( .IN1(n7770), .IN2(g7425), .QN(n12634) );
  NAND3X0 U12835 ( .IN1(n12637), .IN2(n12638), .IN3(n12639), .QN(n12628) );
  XOR2X1 U12836 ( .IN1(g2734), .IN2(n8886), .Q(n12639) );
  INVX0 U12837 ( .INP(n8889), .ZN(n8886) );
  NAND3X0 U12838 ( .IN1(n12640), .IN2(n12641), .IN3(n12642), .QN(n8889) );
  NAND2X0 U12839 ( .IN1(n7775), .IN2(g7487), .QN(n12642) );
  NAND2X0 U12840 ( .IN1(n7843), .IN2(g2703), .QN(n12641) );
  NAND2X0 U12841 ( .IN1(n7776), .IN2(g7425), .QN(n12640) );
  XOR2X1 U12842 ( .IN1(g2714), .IN2(n8897), .Q(n12638) );
  INVX0 U12843 ( .INP(n8898), .ZN(n8897) );
  NAND3X0 U12844 ( .IN1(n12643), .IN2(n12644), .IN3(n12645), .QN(n8898) );
  NAND2X0 U12845 ( .IN1(n7783), .IN2(g7487), .QN(n12645) );
  NAND2X0 U12846 ( .IN1(n7846), .IN2(g2703), .QN(n12644) );
  NAND2X0 U12847 ( .IN1(n7784), .IN2(g7425), .QN(n12643) );
  XOR2X1 U12848 ( .IN1(g2720), .IN2(n8892), .Q(n12637) );
  INVX0 U12849 ( .INP(n8893), .ZN(n8892) );
  NAND3X0 U12850 ( .IN1(n12646), .IN2(n12647), .IN3(n12648), .QN(n8893) );
  NAND2X0 U12851 ( .IN1(n7777), .IN2(g7487), .QN(n12648) );
  NAND2X0 U12852 ( .IN1(g2703), .IN2(n8131), .QN(n12647) );
  NAND2X0 U12853 ( .IN1(n7778), .IN2(g7425), .QN(n12646) );
  NAND4X0 U12854 ( .IN1(n12649), .IN2(n12650), .IN3(n12651), .IN4(n12652), 
        .QN(n12627) );
  XOR2X1 U12855 ( .IN1(g2707), .IN2(n8882), .Q(n12652) );
  INVX0 U12856 ( .INP(n8883), .ZN(n8882) );
  NAND3X0 U12857 ( .IN1(n12653), .IN2(n12654), .IN3(n12655), .QN(n8883) );
  NAND2X0 U12858 ( .IN1(n7781), .IN2(g7487), .QN(n12655) );
  NAND2X0 U12859 ( .IN1(n7845), .IN2(g2703), .QN(n12654) );
  NAND2X0 U12860 ( .IN1(n7782), .IN2(g7425), .QN(n12653) );
  NOR2X0 U12861 ( .IN1(n12656), .IN2(n12657), .QN(n12651) );
  XOR2X1 U12862 ( .IN1(n4393), .IN2(n8928), .Q(n12657) );
  INVX0 U12863 ( .INP(n8929), .ZN(n8928) );
  NAND3X0 U12864 ( .IN1(n12658), .IN2(n12659), .IN3(n12660), .QN(n8929) );
  NAND2X0 U12865 ( .IN1(n7767), .IN2(g7487), .QN(n12660) );
  NAND2X0 U12866 ( .IN1(g2703), .IN2(n8132), .QN(n12659) );
  NAND2X0 U12867 ( .IN1(n7768), .IN2(g7425), .QN(n12658) );
  XOR2X1 U12868 ( .IN1(n8101), .IN2(n8901), .Q(n12656) );
  INVX0 U12869 ( .INP(n8902), .ZN(n8901) );
  NAND3X0 U12870 ( .IN1(n12661), .IN2(n12662), .IN3(n12663), .QN(n8902) );
  NAND2X0 U12871 ( .IN1(n7771), .IN2(g7487), .QN(n12663) );
  NAND2X0 U12872 ( .IN1(n7841), .IN2(g2703), .QN(n12662) );
  NAND2X0 U12873 ( .IN1(n7772), .IN2(g7425), .QN(n12661) );
  XOR2X1 U12874 ( .IN1(n4415), .IN2(n8921), .Q(n12650) );
  NAND3X0 U12875 ( .IN1(n12664), .IN2(n12665), .IN3(n12666), .QN(n8921) );
  NAND2X0 U12876 ( .IN1(n7765), .IN2(g7487), .QN(n12666) );
  NAND2X0 U12877 ( .IN1(n7839), .IN2(g2703), .QN(n12665) );
  NAND2X0 U12878 ( .IN1(n7766), .IN2(g7425), .QN(n12664) );
  XOR2X1 U12879 ( .IN1(g2746), .IN2(n8906), .Q(n12649) );
  INVX0 U12880 ( .INP(n8907), .ZN(n8906) );
  NAND3X0 U12881 ( .IN1(n12667), .IN2(n12668), .IN3(n12669), .QN(n8907) );
  NAND2X0 U12882 ( .IN1(n7773), .IN2(g7487), .QN(n12669) );
  NAND2X0 U12883 ( .IN1(n7842), .IN2(g2703), .QN(n12668) );
  NAND2X0 U12884 ( .IN1(n7774), .IN2(g7425), .QN(n12667) );
  NAND2X0 U12885 ( .IN1(n7568), .IN2(g7487), .QN(n12622) );
  INVX0 U12886 ( .INP(n12670), .ZN(n9260) );
  NAND3X0 U12887 ( .IN1(n12671), .IN2(n12672), .IN3(n12673), .QN(n12670) );
  NAND2X0 U12888 ( .IN1(n7567), .IN2(g7487), .QN(n12673) );
  NAND2X0 U12889 ( .IN1(n7625), .IN2(g2703), .QN(n12672) );
  NAND2X0 U12890 ( .IN1(n7575), .IN2(g7425), .QN(n12671) );
  NAND2X0 U12891 ( .IN1(n12674), .IN2(n12675), .QN(g25271) );
  NAND2X0 U12892 ( .IN1(n9335), .IN2(g2116), .QN(n12675) );
  NAND2X0 U12893 ( .IN1(n12676), .IN2(n12615), .QN(n12674) );
  NAND2X0 U12894 ( .IN1(n12677), .IN2(n12678), .QN(g25270) );
  INVX0 U12895 ( .INP(n12679), .ZN(n12678) );
  NOR2X0 U12896 ( .IN1(n12680), .IN2(n7512), .QN(n12679) );
  NAND2X0 U12897 ( .IN1(n12681), .IN2(n12680), .QN(n12677) );
  NAND2X0 U12898 ( .IN1(n12682), .IN2(n12683), .QN(g25268) );
  NAND2X0 U12899 ( .IN1(n12684), .IN2(g2115), .QN(n12683) );
  NAND2X0 U12900 ( .IN1(n12685), .IN2(n12615), .QN(n12682) );
  INVX0 U12901 ( .INP(n12686), .ZN(n12615) );
  NAND4X0 U12902 ( .IN1(n9273), .IN2(n12687), .IN3(n12688), .IN4(n12689), .QN(
        n12686) );
  NAND2X0 U12903 ( .IN1(n8041), .IN2(g7229), .QN(n12689) );
  NOR2X0 U12904 ( .IN1(n12690), .IN2(n12691), .QN(n12688) );
  NOR2X0 U12905 ( .IN1(n4293), .IN2(g2108), .QN(n12691) );
  NOR4X0 U12906 ( .IN1(n12692), .IN2(n12693), .IN3(n12694), .IN4(n12695), .QN(
        n12690) );
  XNOR2X1 U12907 ( .IN1(n4420), .IN2(n9025), .Q(n12695) );
  NAND3X0 U12908 ( .IN1(n12696), .IN2(n12697), .IN3(n12698), .QN(n9025) );
  NAND2X0 U12909 ( .IN1(n7797), .IN2(g7357), .QN(n12698) );
  NAND2X0 U12910 ( .IN1(n7854), .IN2(g2009), .QN(n12697) );
  NAND2X0 U12911 ( .IN1(n7798), .IN2(g7229), .QN(n12696) );
  XNOR2X1 U12912 ( .IN1(n4399), .IN2(n9000), .Q(n12694) );
  NAND3X0 U12913 ( .IN1(n12699), .IN2(n12700), .IN3(n12701), .QN(n9000) );
  NAND2X0 U12914 ( .IN1(g7357), .IN2(n8133), .QN(n12701) );
  NAND2X0 U12915 ( .IN1(n7852), .IN2(g2009), .QN(n12700) );
  NAND2X0 U12916 ( .IN1(n7794), .IN2(g7229), .QN(n12699) );
  NAND3X0 U12917 ( .IN1(n12702), .IN2(n12703), .IN3(n12704), .QN(n12693) );
  XOR2X1 U12918 ( .IN1(n4468), .IN2(n9016), .Q(n12704) );
  NAND3X0 U12919 ( .IN1(n12705), .IN2(n12706), .IN3(n12707), .QN(n9016) );
  NAND2X0 U12920 ( .IN1(n7790), .IN2(g7357), .QN(n12707) );
  NAND2X0 U12921 ( .IN1(n7850), .IN2(g2009), .QN(n12706) );
  NAND2X0 U12922 ( .IN1(n7791), .IN2(g7229), .QN(n12705) );
  XOR2X1 U12923 ( .IN1(g2059), .IN2(n8988), .Q(n12703) );
  INVX0 U12924 ( .INP(n8991), .ZN(n8988) );
  NAND3X0 U12925 ( .IN1(n12708), .IN2(n12709), .IN3(n12710), .QN(n8991) );
  NAND2X0 U12926 ( .IN1(n7788), .IN2(g7357), .QN(n12710) );
  NAND2X0 U12927 ( .IN1(n7849), .IN2(g2009), .QN(n12709) );
  NAND2X0 U12928 ( .IN1(n7789), .IN2(g7229), .QN(n12708) );
  XOR2X1 U12929 ( .IN1(g2020), .IN2(n9010), .Q(n12702) );
  INVX0 U12930 ( .INP(n9012), .ZN(n9010) );
  NAND3X0 U12931 ( .IN1(n12711), .IN2(n12712), .IN3(n12713), .QN(n9012) );
  NAND2X0 U12932 ( .IN1(n7801), .IN2(g7357), .QN(n12713) );
  NAND2X0 U12933 ( .IN1(n7856), .IN2(g2009), .QN(n12712) );
  NAND2X0 U12934 ( .IN1(n7802), .IN2(g7229), .QN(n12711) );
  NAND4X0 U12935 ( .IN1(n12714), .IN2(n12715), .IN3(n12716), .IN4(n12717), 
        .QN(n12692) );
  XOR2X1 U12936 ( .IN1(g2013), .IN2(n8995), .Q(n12717) );
  INVX0 U12937 ( .INP(n8996), .ZN(n8995) );
  NAND3X0 U12938 ( .IN1(n12718), .IN2(n12719), .IN3(n12720), .QN(n8996) );
  NAND2X0 U12939 ( .IN1(n7799), .IN2(g7357), .QN(n12720) );
  NAND2X0 U12940 ( .IN1(n7855), .IN2(g2009), .QN(n12719) );
  NAND2X0 U12941 ( .IN1(n7800), .IN2(g7229), .QN(n12718) );
  NOR2X0 U12942 ( .IN1(n12721), .IN2(n12722), .QN(n12716) );
  XOR2X1 U12943 ( .IN1(n4409), .IN2(n9020), .Q(n12722) );
  INVX0 U12944 ( .INP(n9021), .ZN(n9020) );
  NAND3X0 U12945 ( .IN1(n12723), .IN2(n12724), .IN3(n12725), .QN(n9021) );
  NAND2X0 U12946 ( .IN1(n7792), .IN2(g7357), .QN(n12725) );
  NAND2X0 U12947 ( .IN1(n7851), .IN2(g2009), .QN(n12724) );
  NAND2X0 U12948 ( .IN1(n7793), .IN2(g7229), .QN(n12723) );
  XOR2X1 U12949 ( .IN1(n8106), .IN2(n9042), .Q(n12721) );
  INVX0 U12950 ( .INP(n9043), .ZN(n9042) );
  NAND3X0 U12951 ( .IN1(n12726), .IN2(n12727), .IN3(n12728), .QN(n9043) );
  NAND2X0 U12952 ( .IN1(n7786), .IN2(g7357), .QN(n12728) );
  NAND2X0 U12953 ( .IN1(n7848), .IN2(g2009), .QN(n12727) );
  NAND2X0 U12954 ( .IN1(n7787), .IN2(g7229), .QN(n12726) );
  XOR2X1 U12955 ( .IN1(n4416), .IN2(n9036), .Q(n12715) );
  NAND3X0 U12956 ( .IN1(n12729), .IN2(n12730), .IN3(n12731), .QN(n9036) );
  NAND2X0 U12957 ( .IN1(g7357), .IN2(n8134), .QN(n12731) );
  NAND2X0 U12958 ( .IN1(n7847), .IN2(g2009), .QN(n12730) );
  NAND2X0 U12959 ( .IN1(n7785), .IN2(g7229), .QN(n12729) );
  XOR2X1 U12960 ( .IN1(g2026), .IN2(n9005), .Q(n12714) );
  INVX0 U12961 ( .INP(n9006), .ZN(n9005) );
  NAND3X0 U12962 ( .IN1(n12732), .IN2(n12733), .IN3(n12734), .QN(n9006) );
  NAND2X0 U12963 ( .IN1(n7795), .IN2(g7357), .QN(n12734) );
  NAND2X0 U12964 ( .IN1(n7853), .IN2(g2009), .QN(n12733) );
  NAND2X0 U12965 ( .IN1(n7796), .IN2(g7229), .QN(n12732) );
  NAND2X0 U12966 ( .IN1(n7570), .IN2(g7357), .QN(n12687) );
  INVX0 U12967 ( .INP(n12735), .ZN(n9273) );
  NAND3X0 U12968 ( .IN1(n12736), .IN2(n12737), .IN3(n12738), .QN(n12735) );
  NAND2X0 U12969 ( .IN1(n7569), .IN2(g7357), .QN(n12738) );
  NAND2X0 U12970 ( .IN1(n7627), .IN2(g2009), .QN(n12737) );
  NAND2X0 U12971 ( .IN1(n7576), .IN2(g7229), .QN(n12736) );
  NAND2X0 U12972 ( .IN1(n12739), .IN2(n12740), .QN(g25267) );
  NAND2X0 U12973 ( .IN1(n8530), .IN2(g1422), .QN(n12740) );
  NAND2X0 U12974 ( .IN1(n12741), .IN2(n12681), .QN(n12739) );
  NAND2X0 U12975 ( .IN1(n12742), .IN2(n12743), .QN(g25266) );
  NAND2X0 U12976 ( .IN1(n12744), .IN2(g734), .QN(n12743) );
  NAND2X0 U12977 ( .IN1(n12745), .IN2(n12746), .QN(n12742) );
  NAND2X0 U12978 ( .IN1(n12747), .IN2(n12748), .QN(g25265) );
  NAND2X0 U12979 ( .IN1(n12171), .IN2(n8739), .QN(n12748) );
  NAND2X0 U12980 ( .IN1(n12749), .IN2(n9300), .QN(n12747) );
  XOR2X1 U12981 ( .IN1(n8050), .IN2(n8049), .Q(n12749) );
  NAND2X0 U12982 ( .IN1(n12750), .IN2(n12751), .QN(g25263) );
  NAND2X0 U12983 ( .IN1(n12752), .IN2(g1421), .QN(n12751) );
  NAND2X0 U12984 ( .IN1(n12753), .IN2(n12681), .QN(n12750) );
  INVX0 U12985 ( .INP(n12754), .ZN(n12681) );
  NAND4X0 U12986 ( .IN1(n9289), .IN2(n12755), .IN3(n12756), .IN4(n12757), .QN(
        n12754) );
  NAND2X0 U12987 ( .IN1(n8039), .IN2(g6979), .QN(n12757) );
  NOR2X0 U12988 ( .IN1(n12758), .IN2(n12759), .QN(n12756) );
  NOR2X0 U12989 ( .IN1(test_so51), .IN2(n4294), .QN(n12759) );
  NOR4X0 U12990 ( .IN1(n12760), .IN2(n12761), .IN3(n12762), .IN4(n12763), .QN(
        n12758) );
  XOR2X1 U12991 ( .IN1(n4412), .IN2(n9122), .Q(n12763) );
  INVX0 U12992 ( .INP(n9123), .ZN(n9122) );
  NAND3X0 U12993 ( .IN1(n12764), .IN2(n12765), .IN3(n12766), .QN(n9123) );
  NAND2X0 U12994 ( .IN1(n7814), .IN2(g7161), .QN(n12766) );
  NAND2X0 U12995 ( .IN1(n7863), .IN2(g1315), .QN(n12765) );
  NAND2X0 U12996 ( .IN1(n7815), .IN2(g6979), .QN(n12764) );
  XOR2X1 U12997 ( .IN1(n4417), .IN2(n9152), .Q(n12762) );
  INVX0 U12998 ( .INP(n9153), .ZN(n9152) );
  NAND3X0 U12999 ( .IN1(n12767), .IN2(n12768), .IN3(n12769), .QN(n9153) );
  NAND2X0 U13000 ( .IN1(n7803), .IN2(g7161), .QN(n12769) );
  NAND2X0 U13001 ( .IN1(n7857), .IN2(g1315), .QN(n12768) );
  NAND2X0 U13002 ( .IN1(n7804), .IN2(g6979), .QN(n12767) );
  NAND3X0 U13003 ( .IN1(n12770), .IN2(n12771), .IN3(n12772), .QN(n12761) );
  XOR2X1 U13004 ( .IN1(g1358), .IN2(n9137), .Q(n12772) );
  INVX0 U13005 ( .INP(n9138), .ZN(n9137) );
  NAND3X0 U13006 ( .IN1(n12773), .IN2(n12774), .IN3(n12775), .QN(n9138) );
  NAND2X0 U13007 ( .IN1(g7161), .IN2(n8135), .QN(n12775) );
  NAND2X0 U13008 ( .IN1(n7861), .IN2(g1315), .QN(n12774) );
  NAND2X0 U13009 ( .IN1(n7811), .IN2(g6979), .QN(n12773) );
  XOR2X1 U13010 ( .IN1(g1372), .IN2(n9159), .Q(n12771) );
  INVX0 U13011 ( .INP(n9160), .ZN(n9159) );
  NAND3X0 U13012 ( .IN1(n12776), .IN2(n12777), .IN3(n12778), .QN(n9160) );
  NAND2X0 U13013 ( .IN1(n7805), .IN2(g7161), .QN(n12778) );
  NAND2X0 U13014 ( .IN1(n7858), .IN2(g1315), .QN(n12777) );
  NAND2X0 U13015 ( .IN1(n7806), .IN2(g6979), .QN(n12776) );
  XOR2X1 U13016 ( .IN1(g1319), .IN2(n9112), .Q(n12770) );
  INVX0 U13017 ( .INP(n9113), .ZN(n9112) );
  NAND3X0 U13018 ( .IN1(n12779), .IN2(n12780), .IN3(n12781), .QN(n9113) );
  NAND2X0 U13019 ( .IN1(n7818), .IN2(g7161), .QN(n12781) );
  NAND2X0 U13020 ( .IN1(n7865), .IN2(g1315), .QN(n12780) );
  NAND2X0 U13021 ( .IN1(n7819), .IN2(g6979), .QN(n12779) );
  NAND4X0 U13022 ( .IN1(n12782), .IN2(n12783), .IN3(n12784), .IN4(n12785), 
        .QN(n12760) );
  XOR2X1 U13023 ( .IN1(n4469), .IN2(n9133), .Q(n12785) );
  NAND3X0 U13024 ( .IN1(n12786), .IN2(n12787), .IN3(n12788), .QN(n9133) );
  NAND2X0 U13025 ( .IN1(n7809), .IN2(g7161), .QN(n12788) );
  NAND2X0 U13026 ( .IN1(n7860), .IN2(g1315), .QN(n12787) );
  NAND2X0 U13027 ( .IN1(n7810), .IN2(g6979), .QN(n12786) );
  NOR2X0 U13028 ( .IN1(n12789), .IN2(n12790), .QN(n12784) );
  XNOR2X1 U13029 ( .IN1(n4402), .IN2(n9128), .Q(n12790) );
  NAND3X0 U13030 ( .IN1(n12791), .IN2(n12792), .IN3(n12793), .QN(n9128) );
  NAND2X0 U13031 ( .IN1(n7820), .IN2(g7161), .QN(n12793) );
  NAND2X0 U13032 ( .IN1(n7866), .IN2(g1315), .QN(n12792) );
  NAND2X0 U13033 ( .IN1(g6979), .IN2(n8136), .QN(n12791) );
  XOR2X1 U13034 ( .IN1(n4475), .IN2(n9105), .Q(n12789) );
  INVX0 U13035 ( .INP(n9108), .ZN(n9105) );
  NAND3X0 U13036 ( .IN1(n12794), .IN2(n12795), .IN3(n12796), .QN(n9108) );
  NAND2X0 U13037 ( .IN1(n7807), .IN2(g7161), .QN(n12796) );
  NAND2X0 U13038 ( .IN1(n7859), .IN2(g1315), .QN(n12795) );
  NAND2X0 U13039 ( .IN1(n7808), .IN2(g6979), .QN(n12794) );
  XOR2X1 U13040 ( .IN1(g1346), .IN2(n9116), .Q(n12783) );
  INVX0 U13041 ( .INP(n9119), .ZN(n9116) );
  NAND3X0 U13042 ( .IN1(n12797), .IN2(n12798), .IN3(n12799), .QN(n9119) );
  NAND2X0 U13043 ( .IN1(n7812), .IN2(g7161), .QN(n12799) );
  NAND2X0 U13044 ( .IN1(n7862), .IN2(g1315), .QN(n12798) );
  NAND2X0 U13045 ( .IN1(n7813), .IN2(g6979), .QN(n12797) );
  XOR2X1 U13046 ( .IN1(n4421), .IN2(n9142), .Q(n12782) );
  NAND3X0 U13047 ( .IN1(n12800), .IN2(n12801), .IN3(n12802), .QN(n9142) );
  NAND2X0 U13048 ( .IN1(n7816), .IN2(g7161), .QN(n12802) );
  NAND2X0 U13049 ( .IN1(n7864), .IN2(g1315), .QN(n12801) );
  NAND2X0 U13050 ( .IN1(n7817), .IN2(g6979), .QN(n12800) );
  NAND2X0 U13051 ( .IN1(n7572), .IN2(g7161), .QN(n12755) );
  INVX0 U13052 ( .INP(n12803), .ZN(n9289) );
  NAND3X0 U13053 ( .IN1(n12804), .IN2(n12805), .IN3(n12806), .QN(n12803) );
  NAND2X0 U13054 ( .IN1(n7571), .IN2(g7161), .QN(n12806) );
  NAND2X0 U13055 ( .IN1(n7629), .IN2(g1315), .QN(n12805) );
  NAND2X0 U13056 ( .IN1(n7577), .IN2(g6979), .QN(n12804) );
  NAND2X0 U13057 ( .IN1(n12807), .IN2(n12808), .QN(g25262) );
  NAND2X0 U13058 ( .IN1(n8551), .IN2(g736), .QN(n12808) );
  NAND2X0 U13059 ( .IN1(n12809), .IN2(n12745), .QN(n12807) );
  NAND2X0 U13060 ( .IN1(n12810), .IN2(n12811), .QN(g25260) );
  NAND2X0 U13061 ( .IN1(n12812), .IN2(g735), .QN(n12811) );
  NAND2X0 U13062 ( .IN1(n12813), .IN2(n12745), .QN(n12810) );
  INVX0 U13063 ( .INP(n12814), .ZN(n12745) );
  NAND4X0 U13064 ( .IN1(n9243), .IN2(n12815), .IN3(n12816), .IN4(n12817), .QN(
        n12814) );
  NAND2X0 U13065 ( .IN1(n8038), .IN2(g6677), .QN(n12817) );
  NOR2X0 U13066 ( .IN1(n12818), .IN2(n12819), .QN(n12816) );
  NOR2X0 U13067 ( .IN1(n4295), .IN2(g728), .QN(n12819) );
  NOR4X0 U13068 ( .IN1(n12820), .IN2(n12821), .IN3(n12822), .IN4(n12823), .QN(
        n12818) );
  XOR2X1 U13069 ( .IN1(n4422), .IN2(n8785), .Q(n12823) );
  INVX0 U13070 ( .INP(n8786), .ZN(n8785) );
  NAND3X0 U13071 ( .IN1(n12824), .IN2(n12825), .IN3(n12826), .QN(n8786) );
  NAND2X0 U13072 ( .IN1(n7833), .IN2(g6911), .QN(n12826) );
  NAND2X0 U13073 ( .IN1(n7874), .IN2(g629), .QN(n12825) );
  NAND2X0 U13074 ( .IN1(n7834), .IN2(g6677), .QN(n12824) );
  XOR2X1 U13075 ( .IN1(n4477), .IN2(n8794), .Q(n12822) );
  INVX0 U13076 ( .INP(n8795), .ZN(n8794) );
  NAND3X0 U13077 ( .IN1(n12827), .IN2(n12828), .IN3(n12829), .QN(n8795) );
  NAND2X0 U13078 ( .IN1(n7824), .IN2(g6911), .QN(n12829) );
  NAND2X0 U13079 ( .IN1(n7869), .IN2(g629), .QN(n12828) );
  NAND2X0 U13080 ( .IN1(n7825), .IN2(g6677), .QN(n12827) );
  NAND3X0 U13081 ( .IN1(n12830), .IN2(n12831), .IN3(n12832), .QN(n12821) );
  XOR2X1 U13082 ( .IN1(g660), .IN2(n8770), .Q(n12832) );
  INVX0 U13083 ( .INP(n8771), .ZN(n8770) );
  NAND3X0 U13084 ( .IN1(n12833), .IN2(n12834), .IN3(n12835), .QN(n8771) );
  NAND2X0 U13085 ( .IN1(n7830), .IN2(g6911), .QN(n12835) );
  NAND2X0 U13086 ( .IN1(n7872), .IN2(g629), .QN(n12834) );
  NAND2X0 U13087 ( .IN1(g6677), .IN2(n8137), .QN(n12833) );
  XOR2X1 U13088 ( .IN1(g640), .IN2(n8790), .Q(n12831) );
  INVX0 U13089 ( .INP(n8791), .ZN(n8790) );
  NAND3X0 U13090 ( .IN1(n12836), .IN2(n12837), .IN3(n12838), .QN(n8791) );
  NAND2X0 U13091 ( .IN1(n7837), .IN2(g6911), .QN(n12838) );
  NAND2X0 U13092 ( .IN1(n7876), .IN2(g629), .QN(n12837) );
  NAND2X0 U13093 ( .IN1(n7838), .IN2(g6677), .QN(n12836) );
  XOR2X1 U13094 ( .IN1(g646), .IN2(n8775), .Q(n12830) );
  INVX0 U13095 ( .INP(n8776), .ZN(n8775) );
  NAND3X0 U13096 ( .IN1(n12839), .IN2(n12840), .IN3(n12841), .QN(n8776) );
  NAND2X0 U13097 ( .IN1(n7831), .IN2(g6911), .QN(n12841) );
  NAND2X0 U13098 ( .IN1(n7873), .IN2(g629), .QN(n12840) );
  NAND2X0 U13099 ( .IN1(n7832), .IN2(g6677), .QN(n12839) );
  NAND4X0 U13100 ( .IN1(n12842), .IN2(n12843), .IN3(n12844), .IN4(n12845), 
        .QN(n12820) );
  XOR2X1 U13101 ( .IN1(g633), .IN2(n8780), .Q(n12845) );
  INVX0 U13102 ( .INP(n8781), .ZN(n8780) );
  NAND3X0 U13103 ( .IN1(n12846), .IN2(n12847), .IN3(n12848), .QN(n8781) );
  NAND2X0 U13104 ( .IN1(n7835), .IN2(g6911), .QN(n12848) );
  NAND2X0 U13105 ( .IN1(n7875), .IN2(g629), .QN(n12847) );
  NAND2X0 U13106 ( .IN1(n7836), .IN2(g6677), .QN(n12846) );
  NOR2X0 U13107 ( .IN1(n12849), .IN2(n12850), .QN(n12844) );
  XOR2X1 U13108 ( .IN1(n4396), .IN2(n8805), .Q(n12850) );
  INVX0 U13109 ( .INP(n8806), .ZN(n8805) );
  NAND3X0 U13110 ( .IN1(n12851), .IN2(n12852), .IN3(n12853), .QN(n8806) );
  NAND2X0 U13111 ( .IN1(n7822), .IN2(g6911), .QN(n12853) );
  NAND2X0 U13112 ( .IN1(n7868), .IN2(g629), .QN(n12852) );
  NAND2X0 U13113 ( .IN1(n7823), .IN2(g6677), .QN(n12851) );
  XOR2X1 U13114 ( .IN1(n8105), .IN2(n8763), .Q(n12849) );
  INVX0 U13115 ( .INP(n8766), .ZN(n8763) );
  NAND3X0 U13116 ( .IN1(n12854), .IN2(n12855), .IN3(n12856), .QN(n8766) );
  NAND2X0 U13117 ( .IN1(n7826), .IN2(g6911), .QN(n12856) );
  NAND2X0 U13118 ( .IN1(n7870), .IN2(g629), .QN(n12855) );
  NAND2X0 U13119 ( .IN1(n7827), .IN2(g6677), .QN(n12854) );
  XOR2X1 U13120 ( .IN1(n4418), .IN2(n8814), .Q(n12843) );
  NAND3X0 U13121 ( .IN1(n12857), .IN2(n12858), .IN3(n12859), .QN(n8814) );
  NAND2X0 U13122 ( .IN1(g6911), .IN2(n8138), .QN(n12859) );
  NAND2X0 U13123 ( .IN1(n7867), .IN2(g629), .QN(n12858) );
  NAND2X0 U13124 ( .IN1(n7821), .IN2(g6677), .QN(n12857) );
  XOR2X1 U13125 ( .IN1(g672), .IN2(n8757), .Q(n12842) );
  INVX0 U13126 ( .INP(n8760), .ZN(n8757) );
  NAND3X0 U13127 ( .IN1(n12860), .IN2(n12861), .IN3(n12862), .QN(n8760) );
  NAND2X0 U13128 ( .IN1(n7828), .IN2(g6911), .QN(n12862) );
  NAND2X0 U13129 ( .IN1(n7871), .IN2(g629), .QN(n12861) );
  NAND2X0 U13130 ( .IN1(n7829), .IN2(g6677), .QN(n12860) );
  NAND2X0 U13131 ( .IN1(n7574), .IN2(g6911), .QN(n12815) );
  INVX0 U13132 ( .INP(n12863), .ZN(n9243) );
  NAND3X0 U13133 ( .IN1(n12864), .IN2(n12865), .IN3(n12866), .QN(n12863) );
  NAND2X0 U13134 ( .IN1(n7573), .IN2(g6911), .QN(n12866) );
  NAND2X0 U13135 ( .IN1(n7630), .IN2(g629), .QN(n12865) );
  NAND2X0 U13136 ( .IN1(n7578), .IN2(g6677), .QN(n12864) );
  NAND2X0 U13137 ( .IN1(n12867), .IN2(n12868), .QN(g25259) );
  INVX0 U13138 ( .INP(n12869), .ZN(n12868) );
  NOR2X0 U13139 ( .IN1(n12870), .IN2(n7579), .QN(n12869) );
  NAND2X0 U13140 ( .IN1(n12870), .IN2(n12075), .QN(n12867) );
  NAND2X0 U13141 ( .IN1(n12871), .IN2(n12872), .QN(g25257) );
  INVX0 U13142 ( .INP(n12873), .ZN(n12872) );
  NOR2X0 U13143 ( .IN1(n12874), .IN2(n7580), .QN(n12873) );
  NAND2X0 U13144 ( .IN1(n12874), .IN2(n12075), .QN(n12871) );
  NAND2X0 U13145 ( .IN1(n12875), .IN2(n12876), .QN(g25256) );
  NAND2X0 U13146 ( .IN1(n12870), .IN2(n4377), .QN(n12876) );
  INVX0 U13147 ( .INP(n12877), .ZN(n12875) );
  NOR2X0 U13148 ( .IN1(n12870), .IN2(n7582), .QN(n12877) );
  NAND2X0 U13149 ( .IN1(n12878), .IN2(n12879), .QN(g25255) );
  NAND2X0 U13150 ( .IN1(n12880), .IN2(n12108), .QN(n12879) );
  NAND2X0 U13151 ( .IN1(n12881), .IN2(g1559), .QN(n12878) );
  NAND2X0 U13152 ( .IN1(n12882), .IN2(n12883), .QN(g25253) );
  INVX0 U13153 ( .INP(n12884), .ZN(n12883) );
  NOR2X0 U13154 ( .IN1(n12885), .IN2(n7581), .QN(n12884) );
  NAND2X0 U13155 ( .IN1(n12885), .IN2(n12075), .QN(n12882) );
  NAND4X0 U13156 ( .IN1(g2200), .IN2(g2175), .IN3(n12886), .IN4(n12887), .QN(
        n12075) );
  NOR4X0 U13157 ( .IN1(n4563), .IN2(n4555), .IN3(n4389), .IN4(n4377), .QN(
        n12887) );
  NOR2X0 U13158 ( .IN1(n4373), .IN2(n4325), .QN(n12886) );
  NAND2X0 U13159 ( .IN1(n12888), .IN2(n12889), .QN(g25252) );
  NAND2X0 U13160 ( .IN1(n12874), .IN2(n4377), .QN(n12889) );
  INVX0 U13161 ( .INP(n12890), .ZN(n12888) );
  NOR2X0 U13162 ( .IN1(n12874), .IN2(n7583), .QN(n12890) );
  NAND2X0 U13163 ( .IN1(n12891), .IN2(n12892), .QN(g25251) );
  NAND2X0 U13164 ( .IN1(n12870), .IN2(n4373), .QN(n12892) );
  INVX0 U13165 ( .INP(n12893), .ZN(n12891) );
  NOR2X0 U13166 ( .IN1(n12870), .IN2(n7585), .QN(n12893) );
  NAND2X0 U13167 ( .IN1(n12894), .IN2(n12895), .QN(g25250) );
  INVX0 U13168 ( .INP(n12896), .ZN(n12895) );
  NOR2X0 U13169 ( .IN1(n12897), .IN2(n7592), .QN(n12896) );
  NAND2X0 U13170 ( .IN1(n12897), .IN2(n12108), .QN(n12894) );
  NAND2X0 U13171 ( .IN1(n12898), .IN2(n12899), .QN(g25249) );
  NAND2X0 U13172 ( .IN1(n12880), .IN2(n4378), .QN(n12899) );
  NAND2X0 U13173 ( .IN1(n12881), .IN2(g1556), .QN(n12898) );
  NAND2X0 U13174 ( .IN1(n12900), .IN2(n12901), .QN(g25248) );
  INVX0 U13175 ( .INP(n12902), .ZN(n12901) );
  NOR2X0 U13176 ( .IN1(n12903), .IN2(n7602), .QN(n12902) );
  NAND2X0 U13177 ( .IN1(n12903), .IN2(n12138), .QN(n12900) );
  NAND2X0 U13178 ( .IN1(n12904), .IN2(n12905), .QN(g25247) );
  NAND2X0 U13179 ( .IN1(n12885), .IN2(n4377), .QN(n12905) );
  INVX0 U13180 ( .INP(n12906), .ZN(n12904) );
  NOR2X0 U13181 ( .IN1(n12885), .IN2(n7584), .QN(n12906) );
  NAND2X0 U13182 ( .IN1(n12907), .IN2(n12908), .QN(g25246) );
  NAND2X0 U13183 ( .IN1(n12874), .IN2(n4373), .QN(n12908) );
  INVX0 U13184 ( .INP(n12909), .ZN(n12907) );
  NOR2X0 U13185 ( .IN1(n12874), .IN2(n7586), .QN(n12909) );
  NAND2X0 U13186 ( .IN1(n12910), .IN2(n12911), .QN(g25245) );
  NAND2X0 U13187 ( .IN1(n12912), .IN2(n12870), .QN(n12911) );
  INVX0 U13188 ( .INP(n12913), .ZN(n12910) );
  NOR2X0 U13189 ( .IN1(n12870), .IN2(n7588), .QN(n12913) );
  NOR2X0 U13190 ( .IN1(n12914), .IN2(n4367), .QN(n12870) );
  NAND2X0 U13191 ( .IN1(n12915), .IN2(n12916), .QN(g25244) );
  INVX0 U13192 ( .INP(n12917), .ZN(n12916) );
  NOR2X0 U13193 ( .IN1(n12918), .IN2(n7593), .QN(n12917) );
  NAND2X0 U13194 ( .IN1(n12918), .IN2(n12108), .QN(n12915) );
  NAND4X0 U13195 ( .IN1(g1506), .IN2(g1481), .IN3(n12919), .IN4(n12920), .QN(
        n12108) );
  NOR4X0 U13196 ( .IN1(n4565), .IN2(n4557), .IN3(n4390), .IN4(n4378), .QN(
        n12920) );
  NOR2X0 U13197 ( .IN1(n4374), .IN2(n4326), .QN(n12919) );
  NAND2X0 U13198 ( .IN1(n12921), .IN2(n12922), .QN(g25243) );
  NAND2X0 U13199 ( .IN1(n12897), .IN2(n4378), .QN(n12922) );
  INVX0 U13200 ( .INP(n12923), .ZN(n12921) );
  NOR2X0 U13201 ( .IN1(n12897), .IN2(n7595), .QN(n12923) );
  NAND2X0 U13202 ( .IN1(n12924), .IN2(n12925), .QN(g25242) );
  NAND2X0 U13203 ( .IN1(test_so54), .IN2(n12881), .QN(n12925) );
  NAND2X0 U13204 ( .IN1(n12880), .IN2(n4374), .QN(n12924) );
  NAND2X0 U13205 ( .IN1(n12926), .IN2(n12927), .QN(g25241) );
  NAND2X0 U13206 ( .IN1(n12928), .IN2(n12138), .QN(n12927) );
  NAND2X0 U13207 ( .IN1(n12929), .IN2(g867), .QN(n12926) );
  NAND2X0 U13208 ( .IN1(n12930), .IN2(n12931), .QN(g25240) );
  NAND2X0 U13209 ( .IN1(n4379), .IN2(n12903), .QN(n12931) );
  INVX0 U13210 ( .INP(n12932), .ZN(n12930) );
  NOR2X0 U13211 ( .IN1(n12903), .IN2(n7605), .QN(n12932) );
  NAND2X0 U13212 ( .IN1(n12933), .IN2(n12934), .QN(g25239) );
  INVX0 U13213 ( .INP(n12935), .ZN(n12934) );
  NOR2X0 U13214 ( .IN1(n12936), .IN2(n7613), .QN(n12935) );
  NAND2X0 U13215 ( .IN1(n12936), .IN2(n12163), .QN(n12933) );
  NAND2X0 U13216 ( .IN1(n12937), .IN2(n12938), .QN(g25237) );
  NAND2X0 U13217 ( .IN1(n12885), .IN2(n4373), .QN(n12938) );
  INVX0 U13218 ( .INP(n12939), .ZN(n12937) );
  NOR2X0 U13219 ( .IN1(n12885), .IN2(n7587), .QN(n12939) );
  NAND2X0 U13220 ( .IN1(n12940), .IN2(n12941), .QN(g25236) );
  NAND2X0 U13221 ( .IN1(n12912), .IN2(n12874), .QN(n12941) );
  INVX0 U13222 ( .INP(n12942), .ZN(n12940) );
  NOR2X0 U13223 ( .IN1(n12874), .IN2(n7589), .QN(n12942) );
  NOR2X0 U13224 ( .IN1(n12914), .IN2(n8097), .QN(n12874) );
  NAND2X0 U13225 ( .IN1(n12943), .IN2(n12944), .QN(g25235) );
  NAND2X0 U13226 ( .IN1(n12918), .IN2(n4378), .QN(n12944) );
  INVX0 U13227 ( .INP(n12945), .ZN(n12943) );
  NOR2X0 U13228 ( .IN1(n12918), .IN2(n7596), .QN(n12945) );
  NAND2X0 U13229 ( .IN1(n12946), .IN2(n12947), .QN(g25234) );
  NAND2X0 U13230 ( .IN1(n12897), .IN2(n4374), .QN(n12947) );
  INVX0 U13231 ( .INP(n12948), .ZN(n12946) );
  NOR2X0 U13232 ( .IN1(n12897), .IN2(n7597), .QN(n12948) );
  NAND2X0 U13233 ( .IN1(n12949), .IN2(n12950), .QN(g25233) );
  NAND2X0 U13234 ( .IN1(n12951), .IN2(n12880), .QN(n12950) );
  INVX0 U13235 ( .INP(n12881), .ZN(n12880) );
  NAND2X0 U13236 ( .IN1(n12881), .IN2(g1550), .QN(n12949) );
  NAND2X0 U13237 ( .IN1(n15), .IN2(g1547), .QN(n12881) );
  NAND2X0 U13238 ( .IN1(n12952), .IN2(n12953), .QN(g25232) );
  INVX0 U13239 ( .INP(n12954), .ZN(n12953) );
  NOR2X0 U13240 ( .IN1(n12955), .IN2(n7604), .QN(n12954) );
  NAND2X0 U13241 ( .IN1(n12955), .IN2(n12138), .QN(n12952) );
  NAND4X0 U13242 ( .IN1(g813), .IN2(g793), .IN3(n12956), .IN4(n12957), .QN(
        n12138) );
  NOR4X0 U13243 ( .IN1(n4567), .IN2(n4559), .IN3(n4391), .IN4(n4379), .QN(
        n12957) );
  NOR2X0 U13244 ( .IN1(n4375), .IN2(n4327), .QN(n12956) );
  NAND2X0 U13245 ( .IN1(n12958), .IN2(n12959), .QN(g25231) );
  NAND2X0 U13246 ( .IN1(n4379), .IN2(n12928), .QN(n12959) );
  NAND2X0 U13247 ( .IN1(n12929), .IN2(g864), .QN(n12958) );
  NAND2X0 U13248 ( .IN1(n12960), .IN2(n12961), .QN(g25230) );
  NAND2X0 U13249 ( .IN1(n12903), .IN2(n4375), .QN(n12961) );
  INVX0 U13250 ( .INP(n12962), .ZN(n12960) );
  NOR2X0 U13251 ( .IN1(n12903), .IN2(n7608), .QN(n12962) );
  NAND2X0 U13252 ( .IN1(n12963), .IN2(n12964), .QN(g25229) );
  INVX0 U13253 ( .INP(n12965), .ZN(n12964) );
  NOR2X0 U13254 ( .IN1(n12966), .IN2(n7614), .QN(n12965) );
  NAND2X0 U13255 ( .IN1(n12966), .IN2(n12163), .QN(n12963) );
  NAND2X0 U13256 ( .IN1(n12967), .IN2(n12968), .QN(g25228) );
  NAND2X0 U13257 ( .IN1(n4380), .IN2(n12936), .QN(n12968) );
  INVX0 U13258 ( .INP(n12969), .ZN(n12967) );
  NOR2X0 U13259 ( .IN1(n12936), .IN2(n7616), .QN(n12969) );
  NAND2X0 U13260 ( .IN1(n12970), .IN2(n12971), .QN(g25227) );
  INVX0 U13261 ( .INP(n12972), .ZN(n12971) );
  NOR2X0 U13262 ( .IN1(n12885), .IN2(n7590), .QN(n12972) );
  NAND2X0 U13263 ( .IN1(n12912), .IN2(n12885), .QN(n12970) );
  NOR2X0 U13264 ( .IN1(n12914), .IN2(n4324), .QN(n12885) );
  NOR4X0 U13265 ( .IN1(g2195), .IN2(g2190), .IN3(n4287), .IN4(n4325), .QN(
        n12912) );
  NAND2X0 U13266 ( .IN1(n12973), .IN2(n12974), .QN(g25225) );
  NAND2X0 U13267 ( .IN1(n12918), .IN2(n4374), .QN(n12974) );
  INVX0 U13268 ( .INP(n12975), .ZN(n12973) );
  NOR2X0 U13269 ( .IN1(n12918), .IN2(n7598), .QN(n12975) );
  NAND2X0 U13270 ( .IN1(n12976), .IN2(n12977), .QN(g25224) );
  NAND2X0 U13271 ( .IN1(n12951), .IN2(n12897), .QN(n12977) );
  INVX0 U13272 ( .INP(n12978), .ZN(n12976) );
  NOR2X0 U13273 ( .IN1(n12897), .IN2(n7600), .QN(n12978) );
  NOR2X0 U13274 ( .IN1(n12914), .IN2(n4515), .QN(n12897) );
  NAND2X0 U13275 ( .IN1(n12979), .IN2(n12980), .QN(g25223) );
  NAND2X0 U13276 ( .IN1(n12955), .IN2(n4379), .QN(n12980) );
  INVX0 U13277 ( .INP(n12981), .ZN(n12979) );
  NOR2X0 U13278 ( .IN1(n12955), .IN2(n7607), .QN(n12981) );
  NAND2X0 U13279 ( .IN1(n12982), .IN2(n12983), .QN(g25222) );
  NAND2X0 U13280 ( .IN1(n12928), .IN2(n4375), .QN(n12983) );
  NAND2X0 U13281 ( .IN1(n12929), .IN2(g861), .QN(n12982) );
  NAND2X0 U13282 ( .IN1(n12984), .IN2(n12985), .QN(g25221) );
  NAND2X0 U13283 ( .IN1(n12986), .IN2(n12903), .QN(n12985) );
  INVX0 U13284 ( .INP(n12987), .ZN(n12984) );
  NOR2X0 U13285 ( .IN1(n12903), .IN2(n7611), .QN(n12987) );
  NOR2X0 U13286 ( .IN1(n12914), .IN2(n8096), .QN(n12903) );
  NAND2X0 U13287 ( .IN1(n12988), .IN2(n12989), .QN(g25220) );
  INVX0 U13288 ( .INP(n12990), .ZN(n12989) );
  NOR2X0 U13289 ( .IN1(n12991), .IN2(n7615), .QN(n12990) );
  NAND2X0 U13290 ( .IN1(n12991), .IN2(n12163), .QN(n12988) );
  NAND4X0 U13291 ( .IN1(g125), .IN2(g105), .IN3(n12992), .IN4(n12993), .QN(
        n12163) );
  NOR4X0 U13292 ( .IN1(n4569), .IN2(n4561), .IN3(n4392), .IN4(n4380), .QN(
        n12993) );
  NOR2X0 U13293 ( .IN1(n4376), .IN2(n4328), .QN(n12992) );
  NAND2X0 U13294 ( .IN1(n12994), .IN2(n12995), .QN(g25219) );
  NAND2X0 U13295 ( .IN1(n4380), .IN2(n12966), .QN(n12995) );
  INVX0 U13296 ( .INP(n12996), .ZN(n12994) );
  NOR2X0 U13297 ( .IN1(n12966), .IN2(n7617), .QN(n12996) );
  NAND2X0 U13298 ( .IN1(n12997), .IN2(n12998), .QN(g25218) );
  NAND2X0 U13299 ( .IN1(n12936), .IN2(n4376), .QN(n12998) );
  INVX0 U13300 ( .INP(n12999), .ZN(n12997) );
  NOR2X0 U13301 ( .IN1(n12936), .IN2(n7619), .QN(n12999) );
  NAND2X0 U13302 ( .IN1(n13000), .IN2(n13001), .QN(g25217) );
  INVX0 U13303 ( .INP(n13002), .ZN(n13001) );
  NOR2X0 U13304 ( .IN1(n12918), .IN2(n7601), .QN(n13002) );
  NAND2X0 U13305 ( .IN1(n12951), .IN2(n12918), .QN(n13000) );
  NOR2X0 U13306 ( .IN1(n12914), .IN2(n4317), .QN(n12918) );
  NOR4X0 U13307 ( .IN1(g1501), .IN2(g1496), .IN3(n4288), .IN4(n4326), .QN(
        n12951) );
  NAND2X0 U13308 ( .IN1(n13003), .IN2(n13004), .QN(g25215) );
  NAND2X0 U13309 ( .IN1(n12955), .IN2(n4375), .QN(n13004) );
  INVX0 U13310 ( .INP(n13005), .ZN(n13003) );
  NOR2X0 U13311 ( .IN1(n12955), .IN2(n7610), .QN(n13005) );
  NAND2X0 U13312 ( .IN1(n13006), .IN2(n13007), .QN(g25214) );
  NAND2X0 U13313 ( .IN1(test_so33), .IN2(n12929), .QN(n13007) );
  NAND2X0 U13314 ( .IN1(n12986), .IN2(n12928), .QN(n13006) );
  INVX0 U13315 ( .INP(n12929), .ZN(n12928) );
  NAND2X0 U13316 ( .IN1(n15), .IN2(g6518), .QN(n12929) );
  INVX0 U13317 ( .INP(n12914), .ZN(n15) );
  NAND2X0 U13318 ( .IN1(n13008), .IN2(n13009), .QN(g25213) );
  NAND2X0 U13319 ( .IN1(n12991), .IN2(n4380), .QN(n13009) );
  INVX0 U13320 ( .INP(n13010), .ZN(n13008) );
  NOR2X0 U13321 ( .IN1(n12991), .IN2(n7618), .QN(n13010) );
  NAND2X0 U13322 ( .IN1(n13011), .IN2(n13012), .QN(g25212) );
  NAND2X0 U13323 ( .IN1(n12966), .IN2(n4376), .QN(n13012) );
  INVX0 U13324 ( .INP(n13013), .ZN(n13011) );
  NOR2X0 U13325 ( .IN1(n12966), .IN2(n7620), .QN(n13013) );
  NAND2X0 U13326 ( .IN1(n13014), .IN2(n13015), .QN(g25211) );
  NAND2X0 U13327 ( .IN1(n13016), .IN2(n12936), .QN(n13015) );
  INVX0 U13328 ( .INP(n13017), .ZN(n13014) );
  NOR2X0 U13329 ( .IN1(n12936), .IN2(n7622), .QN(n13017) );
  NOR2X0 U13330 ( .IN1(n12914), .IN2(n4369), .QN(n12936) );
  NAND2X0 U13331 ( .IN1(n13018), .IN2(n13019), .QN(g25209) );
  INVX0 U13332 ( .INP(n13020), .ZN(n13019) );
  NOR2X0 U13333 ( .IN1(n12955), .IN2(n7612), .QN(n13020) );
  NAND2X0 U13334 ( .IN1(n12986), .IN2(n12955), .QN(n13018) );
  NOR2X0 U13335 ( .IN1(n12914), .IN2(n4323), .QN(n12955) );
  NOR4X0 U13336 ( .IN1(g805), .IN2(g809), .IN3(n4289), .IN4(n4327), .QN(n12986) );
  NAND2X0 U13337 ( .IN1(n13021), .IN2(n13022), .QN(g25207) );
  NAND2X0 U13338 ( .IN1(n12991), .IN2(n4376), .QN(n13022) );
  INVX0 U13339 ( .INP(n13023), .ZN(n13021) );
  NOR2X0 U13340 ( .IN1(n12991), .IN2(n7621), .QN(n13023) );
  NAND2X0 U13341 ( .IN1(n13024), .IN2(n13025), .QN(g25206) );
  NAND2X0 U13342 ( .IN1(n13016), .IN2(n12966), .QN(n13025) );
  INVX0 U13343 ( .INP(n13026), .ZN(n13024) );
  NOR2X0 U13344 ( .IN1(n12966), .IN2(n7623), .QN(n13026) );
  NOR2X0 U13345 ( .IN1(n12914), .IN2(n4512), .QN(n12966) );
  NAND2X0 U13346 ( .IN1(n13027), .IN2(n13028), .QN(g25204) );
  INVX0 U13347 ( .INP(n13029), .ZN(n13028) );
  NOR2X0 U13348 ( .IN1(n12991), .IN2(n7624), .QN(n13029) );
  NAND2X0 U13349 ( .IN1(n13016), .IN2(n12991), .QN(n13027) );
  NOR2X0 U13350 ( .IN1(n12914), .IN2(n4318), .QN(n12991) );
  NAND4X0 U13351 ( .IN1(n7715), .IN2(n11817), .IN3(n8037), .IN4(n13030), .QN(
        n12914) );
  NOR4X0 U13352 ( .IN1(n4349), .IN2(n4330), .IN3(g2912), .IN4(g2917), .QN(
        n13030) );
  NOR4X0 U13353 ( .IN1(g121), .IN2(g117), .IN3(n4290), .IN4(n4328), .QN(n13016) );
  NOR2X0 U13354 ( .IN1(n13031), .IN2(n13032), .QN(g25202) );
  XOR2X1 U13355 ( .IN1(n7441), .IN2(n13033), .Q(n13032) );
  NOR3X0 U13356 ( .IN1(n8685), .IN2(n4057), .IN3(n12166), .QN(g25201) );
  NOR2X0 U13357 ( .IN1(n4058), .IN2(n4305), .QN(n12166) );
  NAND2X0 U13358 ( .IN1(n13034), .IN2(g2892), .QN(n4058) );
  NOR2X0 U13359 ( .IN1(n13035), .IN2(n13036), .QN(g25199) );
  XOR2X1 U13360 ( .IN1(n7715), .IN2(n13037), .Q(n13036) );
  NOR2X0 U13361 ( .IN1(n11309), .IN2(n13038), .QN(g25197) );
  XOR2X1 U13362 ( .IN1(n4397), .IN2(n9309), .Q(n13038) );
  NOR2X0 U13363 ( .IN1(n9323), .IN2(n13039), .QN(g25194) );
  XOR2X1 U13364 ( .IN1(n4399), .IN2(n12169), .Q(n13039) );
  NOR2X0 U13365 ( .IN1(n12171), .IN2(n13040), .QN(g25191) );
  XOR2X1 U13366 ( .IN1(n8073), .IN2(n4065), .Q(n13040) );
  NOR2X0 U13367 ( .IN1(n8524), .IN2(n13041), .QN(g25189) );
  XOR2X1 U13368 ( .IN1(n4401), .IN2(n8522), .Q(n13041) );
  NOR2X0 U13369 ( .IN1(n8548), .IN2(n13042), .QN(g25185) );
  XOR2X1 U13370 ( .IN1(n4403), .IN2(n8542), .Q(n13042) );
  NOR2X0 U13371 ( .IN1(n10283), .IN2(n13043), .QN(g25067) );
  XNOR2X1 U13372 ( .IN1(n7702), .IN2(n3888), .Q(n13043) );
  NAND2X0 U13373 ( .IN1(g2241), .IN2(n8591), .QN(n3888) );
  INVX0 U13374 ( .INP(n13044), .ZN(n10283) );
  NAND2X0 U13375 ( .IN1(n13045), .IN2(n11817), .QN(n13044) );
  NOR2X0 U13376 ( .IN1(n10285), .IN2(n13046), .QN(g25056) );
  XNOR2X1 U13377 ( .IN1(n7706), .IN2(n3891), .Q(n13046) );
  NAND2X0 U13378 ( .IN1(g1547), .IN2(n8591), .QN(n3891) );
  INVX0 U13379 ( .INP(n13047), .ZN(n10285) );
  NAND2X0 U13380 ( .IN1(n13048), .IN2(n11817), .QN(n13047) );
  NOR2X0 U13381 ( .IN1(n10287), .IN2(n13049), .QN(g25042) );
  XNOR2X1 U13382 ( .IN1(n7710), .IN2(n3894), .Q(n13049) );
  NAND2X0 U13383 ( .IN1(test_so31), .IN2(n8591), .QN(n3894) );
  INVX0 U13384 ( .INP(n13050), .ZN(n10287) );
  NAND2X0 U13385 ( .IN1(n13051), .IN2(n11817), .QN(n13050) );
  INVX0 U13386 ( .INP(n8591), .ZN(n11817) );
  NOR2X0 U13387 ( .IN1(n10289), .IN2(n13052), .QN(g25027) );
  XNOR2X1 U13388 ( .IN1(n7714), .IN2(n3897), .Q(n13052) );
  NAND2X0 U13389 ( .IN1(g165), .IN2(n8591), .QN(n3897) );
  NOR2X0 U13390 ( .IN1(n13053), .IN2(n8591), .QN(n10289) );
  NAND4X0 U13391 ( .IN1(n7764), .IN2(n4431), .IN3(n13054), .IN4(n4355), .QN(
        n8591) );
  INVX0 U13392 ( .INP(n13055), .ZN(n13054) );
  NAND2X0 U13393 ( .IN1(n4291), .IN2(n4305), .QN(n13055) );
  NAND2X0 U13394 ( .IN1(n3700), .IN2(n13056), .QN(g24734) );
  NAND2X0 U13395 ( .IN1(n11452), .IN2(DFF_146_n1), .QN(n13056) );
  INVX0 U13396 ( .INP(n12485), .ZN(n11452) );
  NAND2X0 U13397 ( .IN1(n3940), .IN2(n3705), .QN(n12485) );
  NAND2X0 U13398 ( .IN1(n13057), .IN2(n13058), .QN(g24557) );
  NAND2X0 U13399 ( .IN1(n9316), .IN2(n9168), .QN(n13058) );
  NAND2X0 U13400 ( .IN1(n4299), .IN2(g2676), .QN(n13057) );
  NAND2X0 U13401 ( .IN1(n13059), .IN2(n13060), .QN(g24548) );
  NAND2X0 U13402 ( .IN1(n4370), .IN2(g2673), .QN(n13060) );
  NAND3X0 U13403 ( .IN1(n9168), .IN2(n10907), .IN3(g7390), .QN(n13059) );
  NAND2X0 U13404 ( .IN1(n13061), .IN2(n13062), .QN(g24547) );
  NAND2X0 U13405 ( .IN1(n9316), .IN2(n10966), .QN(n13062) );
  NOR2X0 U13406 ( .IN1(n10906), .IN2(n4299), .QN(n9316) );
  NAND2X0 U13407 ( .IN1(n4299), .IN2(g2667), .QN(n13061) );
  NAND2X0 U13408 ( .IN1(n13063), .IN2(n13064), .QN(g24545) );
  NAND2X0 U13409 ( .IN1(n9337), .IN2(n11012), .QN(n13064) );
  NAND2X0 U13410 ( .IN1(n4366), .IN2(g1982), .QN(n13063) );
  NAND2X0 U13411 ( .IN1(n13065), .IN2(n13066), .QN(g24538) );
  NAND3X0 U13412 ( .IN1(n9168), .IN2(n10907), .IN3(g7302), .QN(n13066) );
  NAND4X0 U13413 ( .IN1(n13067), .IN2(n13068), .IN3(n13069), .IN4(n13070), 
        .QN(n9168) );
  NAND3X0 U13414 ( .IN1(n9319), .IN2(g185), .IN3(test_so88), .QN(n13070) );
  NAND3X0 U13415 ( .IN1(n13071), .IN2(n13072), .IN3(n13073), .QN(n9319) );
  NAND2X0 U13416 ( .IN1(g7390), .IN2(g2641), .QN(n13073) );
  NAND2X0 U13417 ( .IN1(g2624), .IN2(g2564), .QN(n13072) );
  NAND2X0 U13418 ( .IN1(n10186), .IN2(g2639), .QN(n13071) );
  NAND2X0 U13419 ( .IN1(g2624), .IN2(g2676), .QN(n13069) );
  NAND2X0 U13420 ( .IN1(n10186), .IN2(g2670), .QN(n13068) );
  NAND2X0 U13421 ( .IN1(g7390), .IN2(g2673), .QN(n13067) );
  NAND2X0 U13422 ( .IN1(n4314), .IN2(g2670), .QN(n13065) );
  NAND2X0 U13423 ( .IN1(n13074), .IN2(n13075), .QN(g24537) );
  NAND2X0 U13424 ( .IN1(n4370), .IN2(g2664), .QN(n13075) );
  NAND3X0 U13425 ( .IN1(n10966), .IN2(n10907), .IN3(g7390), .QN(n13074) );
  NAND2X0 U13426 ( .IN1(n13076), .IN2(n13077), .QN(g24535) );
  NAND2X0 U13427 ( .IN1(n4315), .IN2(g1979), .QN(n13077) );
  NAND3X0 U13428 ( .IN1(n11012), .IN2(n10907), .IN3(g7194), .QN(n13076) );
  NAND2X0 U13429 ( .IN1(n13078), .IN2(n13079), .QN(g24534) );
  NAND2X0 U13430 ( .IN1(n9337), .IN2(n11107), .QN(n13079) );
  NOR2X0 U13431 ( .IN1(n10906), .IN2(n4366), .QN(n9337) );
  NAND2X0 U13432 ( .IN1(n4366), .IN2(g1973), .QN(n13078) );
  NAND2X0 U13433 ( .IN1(n13080), .IN2(n13081), .QN(g24532) );
  NAND2X0 U13434 ( .IN1(n8532), .IN2(n11118), .QN(n13081) );
  NAND2X0 U13435 ( .IN1(n4300), .IN2(g1288), .QN(n13080) );
  NAND2X0 U13436 ( .IN1(n13082), .IN2(n13083), .QN(g24527) );
  NAND2X0 U13437 ( .IN1(n4314), .IN2(g2661), .QN(n13083) );
  NAND3X0 U13438 ( .IN1(n10966), .IN2(n10907), .IN3(n10186), .QN(n13082) );
  NAND4X0 U13439 ( .IN1(n13084), .IN2(n13085), .IN3(n13086), .IN4(n13087), 
        .QN(n10966) );
  NAND3X0 U13440 ( .IN1(g185), .IN2(g2598), .IN3(n9318), .QN(n13087) );
  NAND3X0 U13441 ( .IN1(n13088), .IN2(n13089), .IN3(n13090), .QN(n9318) );
  NAND2X0 U13442 ( .IN1(g7390), .IN2(g2645), .QN(n13090) );
  NAND2X0 U13443 ( .IN1(g7302), .IN2(g2643), .QN(n13089) );
  NAND2X0 U13444 ( .IN1(g2624), .IN2(g2647), .QN(n13088) );
  NAND2X0 U13445 ( .IN1(g7302), .IN2(g2661), .QN(n13086) );
  NAND2X0 U13446 ( .IN1(g2624), .IN2(g2667), .QN(n13085) );
  NAND2X0 U13447 ( .IN1(g7390), .IN2(g2664), .QN(n13084) );
  NAND2X0 U13448 ( .IN1(n13091), .IN2(n13092), .QN(g24525) );
  NAND3X0 U13449 ( .IN1(n11012), .IN2(n10907), .IN3(g7052), .QN(n13092) );
  NAND4X0 U13450 ( .IN1(n13093), .IN2(n13094), .IN3(n13095), .IN4(n13096), 
        .QN(n11012) );
  NAND3X0 U13451 ( .IN1(g185), .IN2(g1922), .IN3(n9340), .QN(n13096) );
  NAND3X0 U13452 ( .IN1(n13097), .IN2(n13098), .IN3(n13099), .QN(n9340) );
  NAND2X0 U13453 ( .IN1(g1930), .IN2(g1870), .QN(n13099) );
  NAND2X0 U13454 ( .IN1(n10234), .IN2(g1945), .QN(n13098) );
  NAND2X0 U13455 ( .IN1(g7194), .IN2(g1947), .QN(n13097) );
  NAND2X0 U13456 ( .IN1(n10234), .IN2(g1976), .QN(n13095) );
  NAND2X0 U13457 ( .IN1(g7194), .IN2(g1979), .QN(n13094) );
  NAND2X0 U13458 ( .IN1(g1930), .IN2(g1982), .QN(n13093) );
  NAND2X0 U13459 ( .IN1(n4296), .IN2(g1976), .QN(n13091) );
  NAND2X0 U13460 ( .IN1(n13100), .IN2(n13101), .QN(g24524) );
  NAND2X0 U13461 ( .IN1(n4315), .IN2(g1970), .QN(n13101) );
  NAND3X0 U13462 ( .IN1(n11107), .IN2(n10907), .IN3(g7194), .QN(n13100) );
  NAND2X0 U13463 ( .IN1(n13102), .IN2(n13103), .QN(g24522) );
  NAND2X0 U13464 ( .IN1(n4316), .IN2(g1285), .QN(n13103) );
  NAND3X0 U13465 ( .IN1(n11118), .IN2(n10907), .IN3(g6944), .QN(n13102) );
  NAND2X0 U13466 ( .IN1(n13104), .IN2(n13105), .QN(g24521) );
  NAND2X0 U13467 ( .IN1(n8532), .IN2(n11210), .QN(n13105) );
  NOR2X0 U13468 ( .IN1(n10906), .IN2(n4300), .QN(n8532) );
  NAND2X0 U13469 ( .IN1(n4300), .IN2(g1279), .QN(n13104) );
  NAND2X0 U13470 ( .IN1(n13106), .IN2(n13107), .QN(g24519) );
  NAND2X0 U13471 ( .IN1(n8553), .IN2(n11221), .QN(n13107) );
  NAND2X0 U13472 ( .IN1(n4313), .IN2(g602), .QN(n13106) );
  NAND2X0 U13473 ( .IN1(n13108), .IN2(n13109), .QN(g24513) );
  NAND2X0 U13474 ( .IN1(n4296), .IN2(g1967), .QN(n13109) );
  NAND3X0 U13475 ( .IN1(n11107), .IN2(n10907), .IN3(n10234), .QN(n13108) );
  NAND4X0 U13476 ( .IN1(n13110), .IN2(n13111), .IN3(n13112), .IN4(n13113), 
        .QN(n11107) );
  NAND3X0 U13477 ( .IN1(g185), .IN2(g1904), .IN3(n9339), .QN(n13113) );
  NAND3X0 U13478 ( .IN1(n13114), .IN2(n13115), .IN3(n13116), .QN(n9339) );
  NAND2X0 U13479 ( .IN1(g1930), .IN2(g1953), .QN(n13116) );
  NAND2X0 U13480 ( .IN1(g7052), .IN2(g1949), .QN(n13115) );
  NAND2X0 U13481 ( .IN1(g7194), .IN2(g1951), .QN(n13114) );
  NAND2X0 U13482 ( .IN1(g7052), .IN2(g1967), .QN(n13112) );
  NAND2X0 U13483 ( .IN1(g7194), .IN2(g1970), .QN(n13111) );
  NAND2X0 U13484 ( .IN1(g1930), .IN2(g1973), .QN(n13110) );
  NAND2X0 U13485 ( .IN1(n13117), .IN2(n13118), .QN(g24511) );
  NAND3X0 U13486 ( .IN1(n11118), .IN2(n10907), .IN3(g6750), .QN(n13118) );
  NAND4X0 U13487 ( .IN1(n13119), .IN2(n13120), .IN3(n13121), .IN4(n13122), 
        .QN(n11118) );
  NAND3X0 U13488 ( .IN1(n8534), .IN2(g185), .IN3(test_so45), .QN(n13122) );
  NAND3X0 U13489 ( .IN1(n13123), .IN2(n13124), .IN3(n13125), .QN(n8534) );
  NAND2X0 U13490 ( .IN1(g6944), .IN2(g1253), .QN(n13125) );
  NAND2X0 U13491 ( .IN1(g6750), .IN2(g1251), .QN(n13124) );
  NAND2X0 U13492 ( .IN1(g1236), .IN2(g1176), .QN(n13123) );
  NAND2X0 U13493 ( .IN1(g1236), .IN2(g1288), .QN(n13121) );
  NAND2X0 U13494 ( .IN1(g6944), .IN2(g1285), .QN(n13120) );
  NAND2X0 U13495 ( .IN1(n11110), .IN2(g1282), .QN(n13119) );
  NAND2X0 U13496 ( .IN1(n4371), .IN2(g1282), .QN(n13117) );
  NAND2X0 U13497 ( .IN1(n13126), .IN2(n13127), .QN(g24510) );
  NAND2X0 U13498 ( .IN1(n4316), .IN2(g1276), .QN(n13127) );
  NAND3X0 U13499 ( .IN1(n11210), .IN2(n10907), .IN3(g6944), .QN(n13126) );
  NAND2X0 U13500 ( .IN1(n13128), .IN2(n13129), .QN(g24508) );
  NAND2X0 U13501 ( .IN1(n4372), .IN2(g599), .QN(n13129) );
  NAND3X0 U13502 ( .IN1(n11221), .IN2(n10907), .IN3(g6642), .QN(n13128) );
  NAND2X0 U13503 ( .IN1(n13130), .IN2(n13131), .QN(g24507) );
  NAND2X0 U13504 ( .IN1(n8553), .IN2(n11308), .QN(n13131) );
  NOR2X0 U13505 ( .IN1(n10906), .IN2(n4313), .QN(n8553) );
  NAND2X0 U13506 ( .IN1(n4313), .IN2(g593), .QN(n13130) );
  NAND2X0 U13507 ( .IN1(n13132), .IN2(n13133), .QN(g24501) );
  NAND2X0 U13508 ( .IN1(n4371), .IN2(g1273), .QN(n13133) );
  NAND3X0 U13509 ( .IN1(n11210), .IN2(n10907), .IN3(n11110), .QN(n13132) );
  NAND4X0 U13510 ( .IN1(n13134), .IN2(n13135), .IN3(n13136), .IN4(n13137), 
        .QN(n11210) );
  NAND3X0 U13511 ( .IN1(g185), .IN2(g1210), .IN3(n8535), .QN(n13137) );
  NAND3X0 U13512 ( .IN1(n13138), .IN2(n13139), .IN3(n13140), .QN(n8535) );
  NAND2X0 U13513 ( .IN1(n11110), .IN2(g1255), .QN(n13140) );
  NAND2X0 U13514 ( .IN1(g1236), .IN2(g1259), .QN(n13139) );
  NAND2X0 U13515 ( .IN1(g6944), .IN2(g1257), .QN(n13138) );
  NAND2X0 U13516 ( .IN1(g6750), .IN2(g1273), .QN(n13136) );
  NAND2X0 U13517 ( .IN1(g1236), .IN2(g1279), .QN(n13135) );
  NAND2X0 U13518 ( .IN1(g6944), .IN2(g1276), .QN(n13134) );
  NAND2X0 U13519 ( .IN1(n13141), .IN2(n13142), .QN(g24499) );
  NAND3X0 U13520 ( .IN1(n11221), .IN2(n10907), .IN3(g6485), .QN(n13142) );
  NAND4X0 U13521 ( .IN1(n13143), .IN2(n13144), .IN3(n13145), .IN4(n13146), 
        .QN(n11221) );
  NAND3X0 U13522 ( .IN1(g185), .IN2(g542), .IN3(n8558), .QN(n13146) );
  NAND3X0 U13523 ( .IN1(n13147), .IN2(n13148), .IN3(n13149), .QN(n8558) );
  NAND2X0 U13524 ( .IN1(g6642), .IN2(g567), .QN(n13149) );
  NAND2X0 U13525 ( .IN1(n11213), .IN2(g565), .QN(n13148) );
  NAND2X0 U13526 ( .IN1(g550), .IN2(g489), .QN(n13147) );
  NAND2X0 U13527 ( .IN1(g6485), .IN2(g596), .QN(n13145) );
  NAND2X0 U13528 ( .IN1(g550), .IN2(g602), .QN(n13144) );
  NAND2X0 U13529 ( .IN1(g6642), .IN2(g599), .QN(n13143) );
  NAND2X0 U13530 ( .IN1(n4298), .IN2(g596), .QN(n13141) );
  NAND2X0 U13531 ( .IN1(n13150), .IN2(n13151), .QN(g24498) );
  NAND2X0 U13532 ( .IN1(n4372), .IN2(g590), .QN(n13151) );
  NAND3X0 U13533 ( .IN1(n11308), .IN2(n10907), .IN3(g6642), .QN(n13150) );
  NAND2X0 U13534 ( .IN1(n13152), .IN2(n13153), .QN(g24491) );
  NAND2X0 U13535 ( .IN1(n4298), .IN2(g587), .QN(n13153) );
  NAND3X0 U13536 ( .IN1(n11308), .IN2(n10907), .IN3(n11213), .QN(n13152) );
  INVX0 U13537 ( .INP(n10906), .ZN(n10907) );
  NOR4X0 U13538 ( .IN1(n4350), .IN2(n4481), .IN3(n13154), .IN4(n13155), .QN(
        n10906) );
  NAND2X0 U13539 ( .IN1(n4480), .IN2(n7441), .QN(n13155) );
  NAND4X0 U13540 ( .IN1(n13156), .IN2(n13157), .IN3(n13158), .IN4(n13159), 
        .QN(n11308) );
  NAND3X0 U13541 ( .IN1(g185), .IN2(g524), .IN3(n8555), .QN(n13159) );
  NAND3X0 U13542 ( .IN1(n13160), .IN2(n13161), .IN3(n13162), .QN(n8555) );
  NAND2X0 U13543 ( .IN1(g6642), .IN2(g571), .QN(n13162) );
  NAND2X0 U13544 ( .IN1(g6485), .IN2(g569), .QN(n13161) );
  NAND2X0 U13545 ( .IN1(g550), .IN2(g573), .QN(n13160) );
  NAND2X0 U13546 ( .IN1(n11213), .IN2(g587), .QN(n13158) );
  NAND2X0 U13547 ( .IN1(g550), .IN2(g593), .QN(n13157) );
  NAND2X0 U13548 ( .IN1(g6642), .IN2(g590), .QN(n13156) );
  NOR3X0 U13549 ( .IN1(n13163), .IN2(n13037), .IN3(n13035), .QN(g24476) );
  NOR3X0 U13550 ( .IN1(n4349), .IN2(n4479), .IN3(n8689), .QN(n13037) );
  NOR2X0 U13551 ( .IN1(n13164), .IN2(g2924), .QN(n13163) );
  NOR2X0 U13552 ( .IN1(n4479), .IN2(n8689), .QN(n13164) );
  NOR2X0 U13553 ( .IN1(n8685), .IN2(n13165), .QN(g24473) );
  XOR2X1 U13554 ( .IN1(n7764), .IN2(n13034), .Q(n13165) );
  NOR3X0 U13555 ( .IN1(n13033), .IN2(n4101), .IN3(n13031), .QN(g24446) );
  INVX0 U13556 ( .INP(n8741), .ZN(n13031) );
  NAND2X0 U13557 ( .IN1(n12171), .IN2(n13166), .QN(n8741) );
  NAND2X0 U13558 ( .IN1(n13167), .IN2(n8739), .QN(n13166) );
  INVX0 U13559 ( .INP(g3234), .ZN(n8739) );
  NAND4X0 U13560 ( .IN1(n4350), .IN2(n4480), .IN3(g3018), .IN4(g3032), .QN(
        n13167) );
  NOR2X0 U13561 ( .IN1(n1547), .IN2(n4480), .QN(n13033) );
  NAND3X0 U13562 ( .IN1(g3028), .IN2(g3018), .IN3(n8742), .QN(n1547) );
  NOR2X0 U13563 ( .IN1(n12171), .IN2(n13168), .QN(g24445) );
  XNOR2X1 U13564 ( .IN1(n8052), .IN2(n4066), .Q(n13168) );
  NAND3X0 U13565 ( .IN1(g3006), .IN2(n7909), .IN3(n9303), .QN(n4066) );
  NOR2X0 U13566 ( .IN1(n8050), .IN2(n8049), .QN(n9303) );
  INVX0 U13567 ( .INP(n9300), .ZN(n12171) );
  NOR2X0 U13568 ( .IN1(g3234), .IN2(n8742), .QN(n9300) );
  NOR2X0 U13569 ( .IN1(n13154), .IN2(n8049), .QN(n8742) );
  NAND4X0 U13570 ( .IN1(n8050), .IN2(g3024), .IN3(n8053), .IN4(n13169), .QN(
        n13154) );
  NOR4X0 U13571 ( .IN1(test_so98), .IN2(n14387), .IN3(n8073), .IN4(n8052), 
        .QN(n13169) );
  NOR3X0 U13572 ( .IN1(n13170), .IN2(n11309), .IN3(n9309), .QN(g24438) );
  NOR3X0 U13573 ( .IN1(n4408), .IN2(n4419), .IN3(n9312), .QN(n9309) );
  NOR2X0 U13574 ( .IN1(n13171), .IN2(g2720), .QN(n13170) );
  NOR2X0 U13575 ( .IN1(n4419), .IN2(n9312), .QN(n13171) );
  NOR3X0 U13576 ( .IN1(n13172), .IN2(n9323), .IN3(n12169), .QN(g24434) );
  NOR3X0 U13577 ( .IN1(n4410), .IN2(n4420), .IN3(n9330), .QN(n12169) );
  NOR2X0 U13578 ( .IN1(n13173), .IN2(g2026), .QN(n13172) );
  NOR2X0 U13579 ( .IN1(n4420), .IN2(n9330), .QN(n13173) );
  NOR3X0 U13580 ( .IN1(n13174), .IN2(n8524), .IN3(n8522), .QN(g24430) );
  NOR3X0 U13581 ( .IN1(n4412), .IN2(n4421), .IN3(n13175), .QN(n8522) );
  NOR2X0 U13582 ( .IN1(n13176), .IN2(g1332), .QN(n13174) );
  NOR2X0 U13583 ( .IN1(n4421), .IN2(n13175), .QN(n13176) );
  INVX0 U13584 ( .INP(n8525), .ZN(n13175) );
  NOR3X0 U13585 ( .IN1(n13177), .IN2(n8548), .IN3(n8542), .QN(g24426) );
  NOR3X0 U13586 ( .IN1(n4414), .IN2(n4422), .IN3(n8545), .QN(n8542) );
  NOR2X0 U13587 ( .IN1(n13178), .IN2(g646), .QN(n13177) );
  NOR2X0 U13588 ( .IN1(n4422), .IN2(n8545), .QN(n13178) );
  NAND2X0 U13589 ( .IN1(n13179), .IN2(n13180), .QN(g24250) );
  NAND2X0 U13590 ( .IN1(n4463), .IN2(g2546), .QN(n13180) );
  NAND2X0 U13591 ( .IN1(n10036), .IN2(g2560), .QN(n13179) );
  NAND2X0 U13592 ( .IN1(n13181), .IN2(n13182), .QN(g24243) );
  NAND2X0 U13593 ( .IN1(n4464), .IN2(g1852), .QN(n13182) );
  NAND2X0 U13594 ( .IN1(n8628), .IN2(g1866), .QN(n13181) );
  NAND2X0 U13595 ( .IN1(n13183), .IN2(n13184), .QN(g24238) );
  NAND2X0 U13596 ( .IN1(n4463), .IN2(g2554), .QN(n13184) );
  NAND2X0 U13597 ( .IN1(n10412), .IN2(g2560), .QN(n13183) );
  NAND2X0 U13598 ( .IN1(n13185), .IN2(n13186), .QN(g24237) );
  NAND2X0 U13599 ( .IN1(n4455), .IN2(g2543), .QN(n13186) );
  NAND2X0 U13600 ( .IN1(n10036), .IN2(g8167), .QN(n13185) );
  NAND2X0 U13601 ( .IN1(n13187), .IN2(n13188), .QN(g24235) );
  NAND2X0 U13602 ( .IN1(n4465), .IN2(g1158), .QN(n13188) );
  NAND2X0 U13603 ( .IN1(n10126), .IN2(g1172), .QN(n13187) );
  NAND2X0 U13604 ( .IN1(n13189), .IN2(n13190), .QN(g24231) );
  NAND2X0 U13605 ( .IN1(n4464), .IN2(g1860), .QN(n13190) );
  NAND2X0 U13606 ( .IN1(n10503), .IN2(g1866), .QN(n13189) );
  NAND2X0 U13607 ( .IN1(n13191), .IN2(n13192), .QN(g24230) );
  NAND2X0 U13608 ( .IN1(n4457), .IN2(g1849), .QN(n13192) );
  NAND2X0 U13609 ( .IN1(n8628), .IN2(g8082), .QN(n13191) );
  NAND2X0 U13610 ( .IN1(n13193), .IN2(n13194), .QN(g24228) );
  NAND2X0 U13611 ( .IN1(n4466), .IN2(g471), .QN(n13194) );
  NAND2X0 U13612 ( .IN1(n8568), .IN2(g485), .QN(n13193) );
  NAND2X0 U13613 ( .IN1(n13195), .IN2(n13196), .QN(g24226) );
  NAND2X0 U13614 ( .IN1(n4455), .IN2(g2553), .QN(n13196) );
  NAND2X0 U13615 ( .IN1(n10412), .IN2(g8167), .QN(n13195) );
  NAND2X0 U13616 ( .IN1(n13197), .IN2(n13198), .QN(g24225) );
  NAND2X0 U13617 ( .IN1(n4456), .IN2(g2540), .QN(n13198) );
  NAND2X0 U13618 ( .IN1(n10036), .IN2(g8087), .QN(n13197) );
  NOR2X0 U13619 ( .IN1(n9724), .IN2(n9728), .QN(n10036) );
  NAND2X0 U13620 ( .IN1(n9729), .IN2(n9735), .QN(n9724) );
  INVX0 U13621 ( .INP(n9744), .ZN(n9729) );
  NAND2X0 U13622 ( .IN1(n13199), .IN2(n13200), .QN(g24223) );
  NAND2X0 U13623 ( .IN1(n4465), .IN2(g1166), .QN(n13200) );
  NAND2X0 U13624 ( .IN1(n10273), .IN2(g1172), .QN(n13199) );
  NAND2X0 U13625 ( .IN1(n13201), .IN2(n13202), .QN(g24222) );
  NAND2X0 U13626 ( .IN1(n4459), .IN2(g1155), .QN(n13202) );
  NAND2X0 U13627 ( .IN1(n10126), .IN2(g8007), .QN(n13201) );
  NAND2X0 U13628 ( .IN1(n13203), .IN2(n13204), .QN(g24219) );
  NAND2X0 U13629 ( .IN1(n4457), .IN2(g1859), .QN(n13204) );
  NAND2X0 U13630 ( .IN1(n10503), .IN2(g8082), .QN(n13203) );
  NAND2X0 U13631 ( .IN1(n13205), .IN2(n13206), .QN(g24218) );
  NAND2X0 U13632 ( .IN1(n4458), .IN2(g1846), .QN(n13206) );
  NAND2X0 U13633 ( .IN1(n8628), .IN2(g8012), .QN(n13205) );
  NOR2X0 U13634 ( .IN1(n9370), .IN2(n9374), .QN(n8628) );
  NAND2X0 U13635 ( .IN1(n9375), .IN2(n9381), .QN(n9370) );
  INVX0 U13636 ( .INP(n9391), .ZN(n9375) );
  NAND2X0 U13637 ( .IN1(n13207), .IN2(n13208), .QN(g24216) );
  NAND2X0 U13638 ( .IN1(n4466), .IN2(g479), .QN(n13208) );
  NAND2X0 U13639 ( .IN1(n10680), .IN2(g485), .QN(n13207) );
  NAND2X0 U13640 ( .IN1(n13209), .IN2(n13210), .QN(g24215) );
  NAND2X0 U13641 ( .IN1(n8568), .IN2(g7956), .QN(n13210) );
  NAND2X0 U13642 ( .IN1(test_so24), .IN2(n4461), .QN(n13209) );
  NAND2X0 U13643 ( .IN1(n13211), .IN2(n13212), .QN(g24214) );
  NAND2X0 U13644 ( .IN1(n4456), .IN2(g2552), .QN(n13212) );
  NAND2X0 U13645 ( .IN1(n10412), .IN2(g8087), .QN(n13211) );
  INVX0 U13646 ( .INP(n10049), .ZN(n10412) );
  NAND3X0 U13647 ( .IN1(n9728), .IN2(n9744), .IN3(n9735), .QN(n10049) );
  INVX0 U13648 ( .INP(n9719), .ZN(n9735) );
  NAND2X0 U13649 ( .IN1(n13213), .IN2(n13214), .QN(g24213) );
  NAND2X0 U13650 ( .IN1(n4459), .IN2(g1165), .QN(n13214) );
  NAND2X0 U13651 ( .IN1(n10273), .IN2(g8007), .QN(n13213) );
  NAND2X0 U13652 ( .IN1(n13215), .IN2(n13216), .QN(g24212) );
  NAND2X0 U13653 ( .IN1(n4460), .IN2(g1152), .QN(n13216) );
  NAND2X0 U13654 ( .IN1(n10126), .IN2(g7961), .QN(n13215) );
  NOR2X0 U13655 ( .IN1(n9207), .IN2(n9192), .QN(n10126) );
  NAND2X0 U13656 ( .IN1(n9186), .IN2(n9196), .QN(n9207) );
  INVX0 U13657 ( .INP(n9198), .ZN(n9186) );
  NAND2X0 U13658 ( .IN1(n13217), .IN2(n13218), .QN(g24209) );
  NAND2X0 U13659 ( .IN1(n4463), .IN2(g2536), .QN(n13218) );
  NAND2X0 U13660 ( .IN1(n13219), .IN2(g2560), .QN(n13217) );
  NAND2X0 U13661 ( .IN1(n13220), .IN2(n13221), .QN(g24208) );
  NAND2X0 U13662 ( .IN1(n4458), .IN2(g1858), .QN(n13221) );
  NAND2X0 U13663 ( .IN1(n10503), .IN2(g8012), .QN(n13220) );
  INVX0 U13664 ( .INP(n10261), .ZN(n10503) );
  NAND3X0 U13665 ( .IN1(n9374), .IN2(n9391), .IN3(n9381), .QN(n10261) );
  INVX0 U13666 ( .INP(n9365), .ZN(n9381) );
  NAND2X0 U13667 ( .IN1(n13222), .IN2(n13223), .QN(g24207) );
  NAND2X0 U13668 ( .IN1(n4461), .IN2(g478), .QN(n13223) );
  NAND2X0 U13669 ( .IN1(n10680), .IN2(g7956), .QN(n13222) );
  NAND2X0 U13670 ( .IN1(n13224), .IN2(n13225), .QN(g24206) );
  NAND2X0 U13671 ( .IN1(g465), .IN2(n8100), .QN(n13225) );
  NAND2X0 U13672 ( .IN1(test_so23), .IN2(n8568), .QN(n13224) );
  NOR2X0 U13673 ( .IN1(n9413), .IN2(n9417), .QN(n8568) );
  NAND2X0 U13674 ( .IN1(n9418), .IN2(n9424), .QN(n9413) );
  INVX0 U13675 ( .INP(n9434), .ZN(n9418) );
  NAND2X0 U13676 ( .IN1(n13226), .IN2(n13227), .QN(g24182) );
  NAND2X0 U13677 ( .IN1(n4464), .IN2(g1842), .QN(n13227) );
  NAND2X0 U13678 ( .IN1(n11907), .IN2(g1866), .QN(n13226) );
  NAND2X0 U13679 ( .IN1(n13228), .IN2(n13229), .QN(g24181) );
  NAND2X0 U13680 ( .IN1(n4460), .IN2(g1164), .QN(n13229) );
  NAND2X0 U13681 ( .IN1(n10273), .IN2(g7961), .QN(n13228) );
  INVX0 U13682 ( .INP(n10137), .ZN(n10273) );
  NAND3X0 U13683 ( .IN1(n9192), .IN2(n9198), .IN3(n9196), .QN(n10137) );
  INVX0 U13684 ( .INP(n9194), .ZN(n9196) );
  NAND2X0 U13685 ( .IN1(n13230), .IN2(n13231), .QN(g24179) );
  NAND2X0 U13686 ( .IN1(n4465), .IN2(g1148), .QN(n13231) );
  NAND2X0 U13687 ( .IN1(n13232), .IN2(g1172), .QN(n13230) );
  NAND2X0 U13688 ( .IN1(n13233), .IN2(n13234), .QN(g24178) );
  NAND2X0 U13689 ( .IN1(g477), .IN2(n8100), .QN(n13234) );
  NAND2X0 U13690 ( .IN1(test_so23), .IN2(n10680), .QN(n13233) );
  INVX0 U13691 ( .INP(n10281), .ZN(n10680) );
  NAND3X0 U13692 ( .IN1(n9417), .IN2(n9434), .IN3(n9424), .QN(n10281) );
  INVX0 U13693 ( .INP(n9408), .ZN(n9424) );
  NAND2X0 U13694 ( .IN1(n13235), .IN2(n13236), .QN(g24174) );
  NAND2X0 U13695 ( .IN1(n4466), .IN2(g461), .QN(n13236) );
  NAND2X0 U13696 ( .IN1(n12005), .IN2(g485), .QN(n13235) );
  NAND2X0 U13697 ( .IN1(n13237), .IN2(n13238), .QN(g24092) );
  NAND2X0 U13698 ( .IN1(g3229), .IN2(n4483), .QN(n13238) );
  NAND2X0 U13699 ( .IN1(n8798), .IN2(g2380), .QN(n13237) );
  NAND2X0 U13700 ( .IN1(n13239), .IN2(n13240), .QN(g24083) );
  NAND2X0 U13701 ( .IN1(g3229), .IN2(n4484), .QN(n13240) );
  NAND2X0 U13702 ( .IN1(n8798), .IN2(g1686), .QN(n13239) );
  NAND2X0 U13703 ( .IN1(n13241), .IN2(n13242), .QN(g24072) );
  NAND2X0 U13704 ( .IN1(g3229), .IN2(n4486), .QN(n13242) );
  NAND2X0 U13705 ( .IN1(n8798), .IN2(g992), .QN(n13241) );
  NAND2X0 U13706 ( .IN1(n13243), .IN2(n13244), .QN(g24059) );
  NAND2X0 U13707 ( .IN1(g3229), .IN2(n4485), .QN(n13244) );
  NAND2X0 U13708 ( .IN1(n8798), .IN2(g305), .QN(n13243) );
  INVX0 U13709 ( .INP(g3229), .ZN(n8798) );
  NAND2X0 U13710 ( .IN1(n13245), .IN2(n13246), .QN(g23418) );
  NAND2X0 U13711 ( .IN1(n4455), .IN2(g2533), .QN(n13246) );
  NAND2X0 U13712 ( .IN1(n13219), .IN2(g8167), .QN(n13245) );
  NAND2X0 U13713 ( .IN1(n13247), .IN2(n13248), .QN(g23413) );
  NAND2X0 U13714 ( .IN1(n11907), .IN2(g8082), .QN(n13248) );
  NAND2X0 U13715 ( .IN1(test_so65), .IN2(n4457), .QN(n13247) );
  NAND2X0 U13716 ( .IN1(n13249), .IN2(n13250), .QN(g23407) );
  NAND2X0 U13717 ( .IN1(n4456), .IN2(g2530), .QN(n13250) );
  NAND2X0 U13718 ( .IN1(n13219), .IN2(g8087), .QN(n13249) );
  INVX0 U13719 ( .INP(n8680), .ZN(n13219) );
  NAND3X0 U13720 ( .IN1(n9719), .IN2(n9744), .IN3(n9723), .QN(n8680) );
  INVX0 U13721 ( .INP(n9728), .ZN(n9723) );
  NAND3X0 U13722 ( .IN1(n13251), .IN2(n13252), .IN3(n13253), .QN(n9728) );
  NAND2X0 U13723 ( .IN1(n7270), .IN2(n10046), .QN(n13253) );
  NAND2X0 U13724 ( .IN1(n7281), .IN2(n10047), .QN(n13252) );
  NAND2X0 U13725 ( .IN1(n7282), .IN2(n10048), .QN(n13251) );
  NAND3X0 U13726 ( .IN1(n13254), .IN2(n13255), .IN3(n13256), .QN(n9744) );
  NAND2X0 U13727 ( .IN1(n7268), .IN2(n10046), .QN(n13256) );
  NAND2X0 U13728 ( .IN1(n7277), .IN2(n10047), .QN(n13255) );
  NAND2X0 U13729 ( .IN1(n7278), .IN2(n10048), .QN(n13254) );
  NAND3X0 U13730 ( .IN1(n13257), .IN2(n13258), .IN3(n13259), .QN(n9719) );
  NAND2X0 U13731 ( .IN1(n7269), .IN2(n10046), .QN(n13259) );
  INVX0 U13732 ( .INP(n4524), .ZN(n10046) );
  NAND2X0 U13733 ( .IN1(n7279), .IN2(n10047), .QN(n13258) );
  INVX0 U13734 ( .INP(n4509), .ZN(n10047) );
  NAND2X0 U13735 ( .IN1(n7280), .IN2(n10048), .QN(n13257) );
  INVX0 U13736 ( .INP(n4516), .ZN(n10048) );
  NAND2X0 U13737 ( .IN1(n13260), .IN2(n13261), .QN(g23406) );
  NAND2X0 U13738 ( .IN1(n4459), .IN2(g1145), .QN(n13261) );
  NAND2X0 U13739 ( .IN1(n13232), .IN2(g8007), .QN(n13260) );
  NAND2X0 U13740 ( .IN1(n13262), .IN2(n13263), .QN(g23400) );
  NAND2X0 U13741 ( .IN1(n4458), .IN2(g1836), .QN(n13263) );
  NAND2X0 U13742 ( .IN1(n11907), .IN2(g8012), .QN(n13262) );
  INVX0 U13743 ( .INP(n8644), .ZN(n11907) );
  NAND3X0 U13744 ( .IN1(n9365), .IN2(n9391), .IN3(n9369), .QN(n8644) );
  INVX0 U13745 ( .INP(n9374), .ZN(n9369) );
  NAND3X0 U13746 ( .IN1(n13264), .IN2(n13265), .IN3(n13266), .QN(n9374) );
  NAND2X0 U13747 ( .IN1(n7273), .IN2(n10092), .QN(n13266) );
  NAND2X0 U13748 ( .IN1(n7287), .IN2(n10093), .QN(n13265) );
  NAND2X0 U13749 ( .IN1(n7288), .IN2(n10094), .QN(n13264) );
  NAND3X0 U13750 ( .IN1(n13267), .IN2(n13268), .IN3(n13269), .QN(n9391) );
  NAND2X0 U13751 ( .IN1(n7271), .IN2(n10092), .QN(n13269) );
  NAND2X0 U13752 ( .IN1(n7283), .IN2(n10093), .QN(n13268) );
  NAND2X0 U13753 ( .IN1(n7284), .IN2(n10094), .QN(n13267) );
  NAND3X0 U13754 ( .IN1(n13270), .IN2(n13271), .IN3(n13272), .QN(n9365) );
  NAND2X0 U13755 ( .IN1(n7272), .IN2(n10092), .QN(n13272) );
  INVX0 U13756 ( .INP(n4525), .ZN(n10092) );
  NAND2X0 U13757 ( .IN1(n7285), .IN2(n10093), .QN(n13271) );
  INVX0 U13758 ( .INP(n4511), .ZN(n10093) );
  NAND2X0 U13759 ( .IN1(n7286), .IN2(n10094), .QN(n13270) );
  INVX0 U13760 ( .INP(n4518), .ZN(n10094) );
  NAND2X0 U13761 ( .IN1(n13273), .IN2(n13274), .QN(g23399) );
  NAND2X0 U13762 ( .IN1(n4461), .IN2(g458), .QN(n13274) );
  NAND2X0 U13763 ( .IN1(n12005), .IN2(g7956), .QN(n13273) );
  NAND2X0 U13764 ( .IN1(n13275), .IN2(n13276), .QN(g23392) );
  NAND2X0 U13765 ( .IN1(n4460), .IN2(g1142), .QN(n13276) );
  NAND2X0 U13766 ( .IN1(n13232), .IN2(g7961), .QN(n13275) );
  INVX0 U13767 ( .INP(n8621), .ZN(n13232) );
  NAND3X0 U13768 ( .IN1(n9194), .IN2(n9198), .IN3(n9206), .QN(n8621) );
  INVX0 U13769 ( .INP(n9192), .ZN(n9206) );
  NAND3X0 U13770 ( .IN1(n13277), .IN2(n13278), .IN3(n13279), .QN(n9192) );
  NAND2X0 U13771 ( .IN1(n7292), .IN2(g1088), .QN(n13279) );
  NAND2X0 U13772 ( .IN1(n7293), .IN2(g5472), .QN(n13278) );
  NAND2X0 U13773 ( .IN1(n7276), .IN2(g6712), .QN(n13277) );
  NAND3X0 U13774 ( .IN1(n13280), .IN2(n13281), .IN3(n13282), .QN(n9198) );
  NAND2X0 U13775 ( .IN1(g1088), .IN2(n8139), .QN(n13282) );
  NAND2X0 U13776 ( .IN1(n7289), .IN2(g5472), .QN(n13281) );
  NAND2X0 U13777 ( .IN1(n7274), .IN2(g6712), .QN(n13280) );
  NAND3X0 U13778 ( .IN1(n13283), .IN2(n13284), .IN3(n13285), .QN(n9194) );
  NAND2X0 U13779 ( .IN1(n7290), .IN2(g1088), .QN(n13285) );
  NAND2X0 U13780 ( .IN1(n7291), .IN2(g5472), .QN(n13284) );
  NAND2X0 U13781 ( .IN1(n7275), .IN2(g6712), .QN(n13283) );
  NAND2X0 U13782 ( .IN1(n13286), .IN2(n13287), .QN(g23385) );
  NAND2X0 U13783 ( .IN1(g455), .IN2(n8100), .QN(n13287) );
  NAND2X0 U13784 ( .IN1(n12005), .IN2(test_so23), .QN(n13286) );
  INVX0 U13785 ( .INP(n8592), .ZN(n12005) );
  NAND3X0 U13786 ( .IN1(n9408), .IN2(n9434), .IN3(n9412), .QN(n8592) );
  INVX0 U13787 ( .INP(n9417), .ZN(n9412) );
  NAND3X0 U13788 ( .IN1(n13288), .IN2(n13289), .IN3(n13290), .QN(n9417) );
  NAND2X0 U13789 ( .IN1(n7301), .IN2(n10176), .QN(n13290) );
  NAND2X0 U13790 ( .IN1(n7300), .IN2(n10177), .QN(n13289) );
  NAND2X0 U13791 ( .IN1(n7299), .IN2(n10178), .QN(n13288) );
  NAND3X0 U13792 ( .IN1(n13291), .IN2(n13292), .IN3(n13293), .QN(n9434) );
  NAND2X0 U13793 ( .IN1(n7296), .IN2(n10176), .QN(n13293) );
  NAND2X0 U13794 ( .IN1(n7295), .IN2(n10177), .QN(n13292) );
  NAND2X0 U13795 ( .IN1(n7294), .IN2(n10178), .QN(n13291) );
  NAND3X0 U13796 ( .IN1(n13294), .IN2(n13295), .IN3(n13296), .QN(n9408) );
  NAND2X0 U13797 ( .IN1(n7298), .IN2(n10176), .QN(n13296) );
  INVX0 U13798 ( .INP(n4520), .ZN(n10176) );
  NAND2X0 U13799 ( .IN1(n10177), .IN2(n8140), .QN(n13295) );
  INVX0 U13800 ( .INP(n4499), .ZN(n10177) );
  NAND2X0 U13801 ( .IN1(n7297), .IN2(n10178), .QN(n13294) );
  INVX0 U13802 ( .INP(n4506), .ZN(n10178) );
  NOR3X0 U13803 ( .IN1(n8685), .IN2(n4122), .IN3(n13034), .QN(g23358) );
  NOR2X0 U13804 ( .IN1(n10), .IN2(n4431), .QN(n13034) );
  NAND2X0 U13805 ( .IN1(n13297), .IN2(g2888), .QN(n10) );
  NOR2X0 U13806 ( .IN1(n13035), .IN2(n13298), .QN(g23357) );
  XOR2X1 U13807 ( .IN1(g2917), .IN2(n8689), .Q(n13298) );
  NAND2X0 U13808 ( .IN1(n13299), .IN2(g2912), .QN(n8689) );
  INVX0 U13809 ( .INP(n8690), .ZN(n13299) );
  INVX0 U13810 ( .INP(n8686), .ZN(n13035) );
  NAND2X0 U13811 ( .IN1(n8685), .IN2(n13300), .QN(n8686) );
  NAND2X0 U13812 ( .IN1(n14383), .IN2(n13301), .QN(n13300) );
  NAND4X0 U13813 ( .IN1(n4479), .IN2(n4349), .IN3(g2912), .IN4(g2920), .QN(
        n13301) );
  NOR2X0 U13814 ( .IN1(n11309), .IN2(n13302), .QN(g23348) );
  XNOR2X1 U13815 ( .IN1(n4419), .IN2(n9312), .Q(n13302) );
  NAND3X0 U13816 ( .IN1(g2714), .IN2(g2707), .IN3(n9314), .QN(n9312) );
  NOR2X0 U13817 ( .IN1(n9323), .IN2(n13303), .QN(g23339) );
  XNOR2X1 U13818 ( .IN1(n4420), .IN2(n9330), .Q(n13303) );
  NAND3X0 U13819 ( .IN1(g2020), .IN2(g2013), .IN3(n9332), .QN(n9330) );
  NOR2X0 U13820 ( .IN1(n8524), .IN2(n13304), .QN(g23329) );
  XOR2X1 U13821 ( .IN1(n4421), .IN2(n8525), .Q(n13304) );
  NOR3X0 U13822 ( .IN1(n4402), .IN2(n4476), .IN3(n8527), .QN(n8525) );
  NOR2X0 U13823 ( .IN1(n8548), .IN2(n13305), .QN(g23324) );
  XNOR2X1 U13824 ( .IN1(n4422), .IN2(n8545), .Q(n13305) );
  NAND3X0 U13825 ( .IN1(g640), .IN2(g633), .IN3(n8547), .QN(n8545) );
  NAND2X0 U13826 ( .IN1(n13306), .IN2(n13307), .QN(g23137) );
  NAND2X0 U13827 ( .IN1(n4464), .IN2(g1869), .QN(n13307) );
  NAND2X0 U13828 ( .IN1(n11370), .IN2(g1866), .QN(n13306) );
  NAND2X0 U13829 ( .IN1(n13308), .IN2(n13309), .QN(g23133) );
  NAND2X0 U13830 ( .IN1(n4455), .IN2(g2562), .QN(n13309) );
  NAND2X0 U13831 ( .IN1(n11347), .IN2(g8167), .QN(n13308) );
  NAND2X0 U13832 ( .IN1(n13310), .IN2(n13311), .QN(g23132) );
  NAND2X0 U13833 ( .IN1(n4456), .IN2(g2555), .QN(n13311) );
  NAND2X0 U13834 ( .IN1(n10306), .IN2(g8087), .QN(n13310) );
  NAND2X0 U13835 ( .IN1(n13312), .IN2(n13313), .QN(g23126) );
  NAND2X0 U13836 ( .IN1(n4465), .IN2(g1175), .QN(n13313) );
  NAND2X0 U13837 ( .IN1(n11393), .IN2(g1172), .QN(n13312) );
  NAND2X0 U13838 ( .IN1(n13314), .IN2(n13315), .QN(g23124) );
  NAND2X0 U13839 ( .IN1(n4457), .IN2(g1868), .QN(n13315) );
  NAND2X0 U13840 ( .IN1(n11370), .IN2(g8082), .QN(n13314) );
  NAND2X0 U13841 ( .IN1(n13316), .IN2(n13317), .QN(g23123) );
  NAND2X0 U13842 ( .IN1(n4458), .IN2(g1861), .QN(n13317) );
  NAND2X0 U13843 ( .IN1(n10321), .IN2(g8012), .QN(n13316) );
  NAND2X0 U13844 ( .IN1(n13318), .IN2(n13319), .QN(g23117) );
  NAND2X0 U13845 ( .IN1(n4466), .IN2(g488), .QN(n13319) );
  NAND2X0 U13846 ( .IN1(n11411), .IN2(g485), .QN(n13318) );
  NAND2X0 U13847 ( .IN1(n13320), .IN2(n13321), .QN(g23114) );
  NAND2X0 U13848 ( .IN1(n4456), .IN2(g2561), .QN(n13321) );
  NAND2X0 U13849 ( .IN1(n11347), .IN2(g8087), .QN(n13320) );
  NAND2X0 U13850 ( .IN1(n13322), .IN2(n13323), .QN(g23111) );
  NAND2X0 U13851 ( .IN1(test_so44), .IN2(n4459), .QN(n13323) );
  NAND2X0 U13852 ( .IN1(n11393), .IN2(g8007), .QN(n13322) );
  NAND2X0 U13853 ( .IN1(n13324), .IN2(n13325), .QN(g23110) );
  NAND2X0 U13854 ( .IN1(n4460), .IN2(g1167), .QN(n13325) );
  NAND2X0 U13855 ( .IN1(n10335), .IN2(g7961), .QN(n13324) );
  NAND2X0 U13856 ( .IN1(n13326), .IN2(n13327), .QN(g23097) );
  NAND2X0 U13857 ( .IN1(n4458), .IN2(g1867), .QN(n13327) );
  NAND2X0 U13858 ( .IN1(n11370), .IN2(g8012), .QN(n13326) );
  NAND3X0 U13859 ( .IN1(n13328), .IN2(n13329), .IN3(n13330), .QN(n11370) );
  NAND2X0 U13860 ( .IN1(g5511), .IN2(g1819), .QN(n13330) );
  NAND2X0 U13861 ( .IN1(test_so59), .IN2(n4618), .QN(n13329) );
  NAND2X0 U13862 ( .IN1(g7014), .IN2(g1822), .QN(n13328) );
  NAND2X0 U13863 ( .IN1(n13331), .IN2(n13332), .QN(g23093) );
  NAND2X0 U13864 ( .IN1(n4461), .IN2(g487), .QN(n13332) );
  NAND2X0 U13865 ( .IN1(n11411), .IN2(g7956), .QN(n13331) );
  NAND2X0 U13866 ( .IN1(n13333), .IN2(n13334), .QN(g23092) );
  NAND2X0 U13867 ( .IN1(g480), .IN2(n8100), .QN(n13334) );
  NAND2X0 U13868 ( .IN1(test_so23), .IN2(n10347), .QN(n13333) );
  NAND2X0 U13869 ( .IN1(n13335), .IN2(n13336), .QN(g23081) );
  NAND2X0 U13870 ( .IN1(n4460), .IN2(g1173), .QN(n13336) );
  NAND2X0 U13871 ( .IN1(n11393), .IN2(g7961), .QN(n13335) );
  NAND3X0 U13872 ( .IN1(n13337), .IN2(n13338), .IN3(n13339), .QN(n11393) );
  NAND2X0 U13873 ( .IN1(g1088), .IN2(g1131), .QN(n13339) );
  NAND2X0 U13874 ( .IN1(g5472), .IN2(g1125), .QN(n13338) );
  NAND2X0 U13875 ( .IN1(g6712), .IN2(g1128), .QN(n13337) );
  NAND2X0 U13876 ( .IN1(n13340), .IN2(n13341), .QN(g23076) );
  NAND2X0 U13877 ( .IN1(n4463), .IN2(g2539), .QN(n13341) );
  NAND2X0 U13878 ( .IN1(n10306), .IN2(g2560), .QN(n13340) );
  NAND2X0 U13879 ( .IN1(n13342), .IN2(n13343), .QN(g23067) );
  NAND2X0 U13880 ( .IN1(g486), .IN2(n8100), .QN(n13343) );
  NAND2X0 U13881 ( .IN1(test_so23), .IN2(n11411), .QN(n13342) );
  NAND3X0 U13882 ( .IN1(n13344), .IN2(n13345), .IN3(n13346), .QN(n11411) );
  NAND2X0 U13883 ( .IN1(g5437), .IN2(g438), .QN(n13346) );
  NAND2X0 U13884 ( .IN1(n4640), .IN2(g444), .QN(n13345) );
  NAND2X0 U13885 ( .IN1(g6447), .IN2(g441), .QN(n13344) );
  NAND2X0 U13886 ( .IN1(n13347), .IN2(n13348), .QN(g23058) );
  NAND2X0 U13887 ( .IN1(n4464), .IN2(g1845), .QN(n13348) );
  NAND2X0 U13888 ( .IN1(n10321), .IN2(g1866), .QN(n13347) );
  NAND2X0 U13889 ( .IN1(n13349), .IN2(n13350), .QN(g23047) );
  NAND2X0 U13890 ( .IN1(n4455), .IN2(g2559), .QN(n13350) );
  NAND2X0 U13891 ( .IN1(n10306), .IN2(g8167), .QN(n13349) );
  INVX0 U13892 ( .INP(n4285), .ZN(n10306) );
  NAND3X0 U13893 ( .IN1(n13351), .IN2(n13352), .IN3(n13353), .QN(n4285) );
  NAND2X0 U13894 ( .IN1(g5555), .IN2(g2492), .QN(n13353) );
  NAND2X0 U13895 ( .IN1(n4606), .IN2(g2498), .QN(n13352) );
  NAND2X0 U13896 ( .IN1(g7264), .IN2(g2495), .QN(n13351) );
  NAND2X0 U13897 ( .IN1(n13354), .IN2(n13355), .QN(g23039) );
  NAND2X0 U13898 ( .IN1(n4465), .IN2(g1151), .QN(n13355) );
  NAND2X0 U13899 ( .IN1(n10335), .IN2(g1172), .QN(n13354) );
  NAND2X0 U13900 ( .IN1(n13356), .IN2(n13357), .QN(g23030) );
  NAND2X0 U13901 ( .IN1(n4457), .IN2(g1865), .QN(n13357) );
  NAND2X0 U13902 ( .IN1(n10321), .IN2(g8082), .QN(n13356) );
  INVX0 U13903 ( .INP(n4284), .ZN(n10321) );
  NAND3X0 U13904 ( .IN1(n13358), .IN2(n13359), .IN3(n13360), .QN(n4284) );
  NAND2X0 U13905 ( .IN1(g5511), .IN2(g1798), .QN(n13360) );
  NAND2X0 U13906 ( .IN1(n4618), .IN2(g1804), .QN(n13359) );
  NAND2X0 U13907 ( .IN1(g7014), .IN2(g1801), .QN(n13358) );
  NAND2X0 U13908 ( .IN1(n13361), .IN2(n13362), .QN(g23022) );
  NAND2X0 U13909 ( .IN1(n4466), .IN2(g464), .QN(n13362) );
  NAND2X0 U13910 ( .IN1(n10347), .IN2(g485), .QN(n13361) );
  NAND2X0 U13911 ( .IN1(n13363), .IN2(n13364), .QN(g23014) );
  NAND2X0 U13912 ( .IN1(n4459), .IN2(g1171), .QN(n13364) );
  NAND2X0 U13913 ( .IN1(n10335), .IN2(g8007), .QN(n13363) );
  INVX0 U13914 ( .INP(n4283), .ZN(n10335) );
  NAND3X0 U13915 ( .IN1(n13365), .IN2(n13366), .IN3(n13367), .QN(n4283) );
  NAND2X0 U13916 ( .IN1(g1088), .IN2(g1110), .QN(n13367) );
  NAND2X0 U13917 ( .IN1(g5472), .IN2(g1104), .QN(n13366) );
  NAND2X0 U13918 ( .IN1(g6712), .IN2(g1107), .QN(n13365) );
  NAND2X0 U13919 ( .IN1(n13368), .IN2(n13369), .QN(g23000) );
  NAND2X0 U13920 ( .IN1(n4461), .IN2(g484), .QN(n13369) );
  NAND2X0 U13921 ( .IN1(n10347), .IN2(g7956), .QN(n13368) );
  INVX0 U13922 ( .INP(n4282), .ZN(n10347) );
  NAND3X0 U13923 ( .IN1(n13370), .IN2(n13371), .IN3(n13372), .QN(n4282) );
  NAND2X0 U13924 ( .IN1(g5437), .IN2(g417), .QN(n13372) );
  NAND2X0 U13925 ( .IN1(n4640), .IN2(g423), .QN(n13371) );
  NAND2X0 U13926 ( .IN1(g6447), .IN2(g420), .QN(n13370) );
  NAND2X0 U13927 ( .IN1(n13373), .IN2(n13374), .QN(g22687) );
  NAND3X0 U13928 ( .IN1(n8887), .IN2(g2584), .IN3(n13375), .QN(n13374) );
  INVX0 U13929 ( .INP(n12390), .ZN(n13375) );
  NAND2X0 U13930 ( .IN1(n13376), .IN2(n13377), .QN(n13373) );
  NAND2X0 U13931 ( .IN1(n8876), .IN2(n12390), .QN(n13376) );
  NAND3X0 U13932 ( .IN1(n13378), .IN2(n13379), .IN3(n13380), .QN(n12390) );
  NAND2X0 U13933 ( .IN1(g7390), .IN2(g2568), .QN(n13380) );
  NAND2X0 U13934 ( .IN1(g2624), .IN2(g2571), .QN(n13379) );
  NAND2X0 U13935 ( .IN1(n10186), .IN2(g2565), .QN(n13378) );
  NAND2X0 U13936 ( .IN1(n13381), .IN2(n13382), .QN(g22651) );
  NAND3X0 U13937 ( .IN1(n9011), .IN2(g1890), .IN3(n13383), .QN(n13382) );
  INVX0 U13938 ( .INP(n12398), .ZN(n13383) );
  NAND2X0 U13939 ( .IN1(n13384), .IN2(n13377), .QN(n13381) );
  NAND2X0 U13940 ( .IN1(n8989), .IN2(n12398), .QN(n13384) );
  NAND3X0 U13941 ( .IN1(n13385), .IN2(n13386), .IN3(n13387), .QN(n12398) );
  NAND2X0 U13942 ( .IN1(g1930), .IN2(g1877), .QN(n13387) );
  NAND2X0 U13943 ( .IN1(test_so68), .IN2(n10234), .QN(n13386) );
  NAND2X0 U13944 ( .IN1(g7194), .IN2(g1874), .QN(n13385) );
  NAND2X0 U13945 ( .IN1(n13388), .IN2(n13389), .QN(g22615) );
  NAND3X0 U13946 ( .IN1(n9117), .IN2(g1196), .IN3(n13390), .QN(n13389) );
  INVX0 U13947 ( .INP(n12406), .ZN(n13390) );
  NAND2X0 U13948 ( .IN1(n13391), .IN2(n13377), .QN(n13388) );
  NAND2X0 U13949 ( .IN1(n9106), .IN2(n12406), .QN(n13391) );
  NAND3X0 U13950 ( .IN1(n13392), .IN2(n13393), .IN3(n13394), .QN(n12406) );
  NAND2X0 U13951 ( .IN1(test_so47), .IN2(n11110), .QN(n13394) );
  NAND2X0 U13952 ( .IN1(g1236), .IN2(g1183), .QN(n13393) );
  NAND2X0 U13953 ( .IN1(g6944), .IN2(g1180), .QN(n13392) );
  NAND2X0 U13954 ( .IN1(n13395), .IN2(n13396), .QN(g22578) );
  NAND3X0 U13955 ( .IN1(test_so22), .IN2(n8764), .IN3(n13397), .QN(n13396) );
  INVX0 U13956 ( .INP(n12411), .ZN(n13397) );
  NAND2X0 U13957 ( .IN1(n13398), .IN2(n13377), .QN(n13395) );
  NAND2X0 U13958 ( .IN1(n8758), .IN2(n12411), .QN(n13398) );
  NAND3X0 U13959 ( .IN1(n13399), .IN2(n13400), .IN3(n13401), .QN(n12411) );
  NAND2X0 U13960 ( .IN1(g6642), .IN2(g493), .QN(n13401) );
  NAND2X0 U13961 ( .IN1(g6485), .IN2(g490), .QN(n13400) );
  NAND2X0 U13962 ( .IN1(g550), .IN2(g496), .QN(n13399) );
  NOR2X0 U13963 ( .IN1(n13402), .IN2(n13403), .QN(g22299) );
  NOR2X0 U13964 ( .IN1(n12607), .IN2(test_so95), .QN(n13403) );
  NOR2X0 U13965 ( .IN1(n11309), .IN2(n13404), .QN(g22284) );
  INVX0 U13966 ( .INP(n13405), .ZN(n13404) );
  NAND2X0 U13967 ( .IN1(n12610), .IN2(n7974), .QN(n13405) );
  NOR2X0 U13968 ( .IN1(n13406), .IN2(n13407), .QN(g22280) );
  NOR2X0 U13969 ( .IN1(n12616), .IN2(g2117), .QN(n13407) );
  NOR2X0 U13970 ( .IN1(n13408), .IN2(n13409), .QN(g22269) );
  INVX0 U13971 ( .INP(n13410), .ZN(n13409) );
  NAND2X0 U13972 ( .IN1(n12619), .IN2(n7877), .QN(n13410) );
  NOR2X0 U13973 ( .IN1(n13411), .IN2(n13412), .QN(g22263) );
  NOR2X0 U13974 ( .IN1(n12680), .IN2(g1423), .QN(n13412) );
  NOR2X0 U13975 ( .IN1(n13413), .IN2(n13414), .QN(g22249) );
  INVX0 U13976 ( .INP(n13415), .ZN(n13414) );
  NAND2X0 U13977 ( .IN1(n12684), .IN2(n7878), .QN(n13415) );
  NOR2X0 U13978 ( .IN1(n13416), .IN2(n13417), .QN(g22242) );
  NOR2X0 U13979 ( .IN1(n12746), .IN2(g737), .QN(n13417) );
  NOR2X0 U13980 ( .IN1(n13418), .IN2(n13419), .QN(g22234) );
  INVX0 U13981 ( .INP(n13420), .ZN(n13419) );
  NAND2X0 U13982 ( .IN1(n12752), .IN2(n7879), .QN(n13420) );
  NOR2X0 U13983 ( .IN1(n13421), .IN2(n13422), .QN(g22218) );
  INVX0 U13984 ( .INP(n13423), .ZN(n13422) );
  NAND2X0 U13985 ( .IN1(n12812), .IN2(n7880), .QN(n13423) );
  NAND2X0 U13986 ( .IN1(n13424), .IN2(n13425), .QN(g22200) );
  NAND2X0 U13987 ( .IN1(n13045), .IN2(n4373), .QN(n13425) );
  INVX0 U13988 ( .INP(n13426), .ZN(n13424) );
  NOR2X0 U13989 ( .IN1(n13045), .IN2(n7531), .QN(n13426) );
  NAND2X0 U13990 ( .IN1(n13427), .IN2(n13428), .QN(g22194) );
  INVX0 U13991 ( .INP(n13429), .ZN(n13428) );
  NOR2X0 U13992 ( .IN1(n13045), .IN2(n7523), .QN(n13429) );
  NAND2X0 U13993 ( .IN1(n13045), .IN2(n9474), .QN(n13427) );
  NAND2X0 U13994 ( .IN1(n13430), .IN2(n13431), .QN(g22193) );
  NAND2X0 U13995 ( .IN1(n13432), .IN2(n4373), .QN(n13431) );
  NAND2X0 U13996 ( .IN1(n13433), .IN2(g2210), .QN(n13430) );
  NAND2X0 U13997 ( .IN1(n13434), .IN2(n13435), .QN(g22192) );
  NAND2X0 U13998 ( .IN1(n13045), .IN2(n4377), .QN(n13435) );
  INVX0 U13999 ( .INP(n13436), .ZN(n13434) );
  NOR2X0 U14000 ( .IN1(n13045), .IN2(n7532), .QN(n13436) );
  NAND2X0 U14001 ( .IN1(n13437), .IN2(n13438), .QN(g22191) );
  NAND2X0 U14002 ( .IN1(n13048), .IN2(n4374), .QN(n13438) );
  INVX0 U14003 ( .INP(n13439), .ZN(n13437) );
  NOR2X0 U14004 ( .IN1(n13048), .IN2(n7542), .QN(n13439) );
  NAND2X0 U14005 ( .IN1(n13440), .IN2(n13441), .QN(g22185) );
  NAND2X0 U14006 ( .IN1(test_so75), .IN2(n13433), .QN(n13441) );
  NAND2X0 U14007 ( .IN1(n13432), .IN2(n9474), .QN(n13440) );
  NAND2X0 U14008 ( .IN1(n13442), .IN2(n13443), .QN(g22184) );
  INVX0 U14009 ( .INP(n13444), .ZN(n13443) );
  NOR2X0 U14010 ( .IN1(n13045), .IN2(n7514), .QN(n13444) );
  NAND2X0 U14011 ( .IN1(n10446), .IN2(n13045), .QN(n13442) );
  NAND2X0 U14012 ( .IN1(n13445), .IN2(n13446), .QN(g22183) );
  NAND2X0 U14013 ( .IN1(n13447), .IN2(n4373), .QN(n13446) );
  INVX0 U14014 ( .INP(n13448), .ZN(n13445) );
  NOR2X0 U14015 ( .IN1(n13447), .IN2(n7893), .QN(n13448) );
  NAND2X0 U14016 ( .IN1(n13449), .IN2(n13450), .QN(g22182) );
  NAND2X0 U14017 ( .IN1(n13432), .IN2(n4377), .QN(n13450) );
  NAND2X0 U14018 ( .IN1(n13433), .IN2(g2207), .QN(n13449) );
  NAND2X0 U14019 ( .IN1(n13451), .IN2(n13452), .QN(g22180) );
  INVX0 U14020 ( .INP(n13453), .ZN(n13452) );
  NOR2X0 U14021 ( .IN1(n13048), .IN2(n7533), .QN(n13453) );
  NAND2X0 U14022 ( .IN1(n13048), .IN2(n9504), .QN(n13451) );
  NAND2X0 U14023 ( .IN1(n13454), .IN2(n13455), .QN(g22179) );
  NAND2X0 U14024 ( .IN1(n13456), .IN2(n4374), .QN(n13455) );
  NAND2X0 U14025 ( .IN1(n13457), .IN2(g1516), .QN(n13454) );
  NAND2X0 U14026 ( .IN1(n13458), .IN2(n13459), .QN(g22178) );
  NAND2X0 U14027 ( .IN1(n13048), .IN2(n4378), .QN(n13459) );
  INVX0 U14028 ( .INP(n13460), .ZN(n13458) );
  NOR2X0 U14029 ( .IN1(n13048), .IN2(n7543), .QN(n13460) );
  NAND2X0 U14030 ( .IN1(n13461), .IN2(n13462), .QN(g22177) );
  NAND2X0 U14031 ( .IN1(n13051), .IN2(n4375), .QN(n13462) );
  INVX0 U14032 ( .INP(n13463), .ZN(n13461) );
  NOR2X0 U14033 ( .IN1(n13051), .IN2(n7556), .QN(n13463) );
  NAND2X0 U14034 ( .IN1(n13464), .IN2(n13465), .QN(g22173) );
  INVX0 U14035 ( .INP(n13466), .ZN(n13465) );
  NOR2X0 U14036 ( .IN1(n13447), .IN2(n7524), .QN(n13466) );
  NAND2X0 U14037 ( .IN1(n13447), .IN2(n9474), .QN(n13464) );
  INVX0 U14038 ( .INP(n10769), .ZN(n9474) );
  NAND3X0 U14039 ( .IN1(n13467), .IN2(n13468), .IN3(n13469), .QN(n10769) );
  NAND2X0 U14040 ( .IN1(n7586), .IN2(test_so73), .QN(n13469) );
  NAND2X0 U14041 ( .IN1(n7587), .IN2(g6837), .QN(n13468) );
  NAND2X0 U14042 ( .IN1(n7585), .IN2(g2241), .QN(n13467) );
  NAND2X0 U14043 ( .IN1(n13470), .IN2(n13471), .QN(g22172) );
  NAND2X0 U14044 ( .IN1(n13433), .IN2(g2237), .QN(n13471) );
  NAND2X0 U14045 ( .IN1(n10446), .IN2(n13432), .QN(n13470) );
  NAND2X0 U14046 ( .IN1(n13472), .IN2(n13473), .QN(g22171) );
  NAND2X0 U14047 ( .IN1(n13045), .IN2(n4287), .QN(n13473) );
  INVX0 U14048 ( .INP(n13474), .ZN(n13472) );
  NOR2X0 U14049 ( .IN1(n13045), .IN2(n7525), .QN(n13474) );
  NAND2X0 U14050 ( .IN1(n13475), .IN2(n13476), .QN(g22170) );
  NAND2X0 U14051 ( .IN1(n13447), .IN2(n4377), .QN(n13476) );
  INVX0 U14052 ( .INP(n13477), .ZN(n13475) );
  NOR2X0 U14053 ( .IN1(n13447), .IN2(n7895), .QN(n13477) );
  NAND2X0 U14054 ( .IN1(n13478), .IN2(n13479), .QN(g22169) );
  NAND2X0 U14055 ( .IN1(n13457), .IN2(g1546), .QN(n13479) );
  NAND2X0 U14056 ( .IN1(n13456), .IN2(n9504), .QN(n13478) );
  NAND2X0 U14057 ( .IN1(n13480), .IN2(n13481), .QN(g22168) );
  INVX0 U14058 ( .INP(n13482), .ZN(n13481) );
  NOR2X0 U14059 ( .IN1(n13048), .IN2(n7517), .QN(n13482) );
  NAND2X0 U14060 ( .IN1(n13483), .IN2(n13048), .QN(n13480) );
  NAND2X0 U14061 ( .IN1(n13484), .IN2(n13485), .QN(g22167) );
  INVX0 U14062 ( .INP(n13486), .ZN(n13485) );
  NOR2X0 U14063 ( .IN1(n8110), .IN2(n13487), .QN(n13486) );
  NAND2X0 U14064 ( .IN1(n13487), .IN2(n4374), .QN(n13484) );
  NAND2X0 U14065 ( .IN1(n13488), .IN2(n13489), .QN(g22166) );
  NAND2X0 U14066 ( .IN1(n13456), .IN2(n4378), .QN(n13489) );
  NAND2X0 U14067 ( .IN1(n13457), .IN2(g1513), .QN(n13488) );
  NAND2X0 U14068 ( .IN1(n13490), .IN2(n13491), .QN(g22164) );
  INVX0 U14069 ( .INP(n13492), .ZN(n13491) );
  NOR2X0 U14070 ( .IN1(n13051), .IN2(n7544), .QN(n13492) );
  NAND2X0 U14071 ( .IN1(n13051), .IN2(n9537), .QN(n13490) );
  NAND2X0 U14072 ( .IN1(n13493), .IN2(n13494), .QN(g22163) );
  NAND2X0 U14073 ( .IN1(n13495), .IN2(n4375), .QN(n13494) );
  INVX0 U14074 ( .INP(n13496), .ZN(n13493) );
  NOR2X0 U14075 ( .IN1(n13495), .IN2(n7935), .QN(n13496) );
  NAND2X0 U14076 ( .IN1(n13497), .IN2(n13498), .QN(g22162) );
  NAND2X0 U14077 ( .IN1(n4379), .IN2(n13051), .QN(n13498) );
  INVX0 U14078 ( .INP(n13499), .ZN(n13497) );
  NOR2X0 U14079 ( .IN1(n13051), .IN2(n7557), .QN(n13499) );
  NAND2X0 U14080 ( .IN1(n13500), .IN2(n13501), .QN(g22161) );
  NAND2X0 U14081 ( .IN1(n13502), .IN2(n4376), .QN(n13501) );
  NAND2X0 U14082 ( .IN1(n13053), .IN2(g132), .QN(n13500) );
  NAND2X0 U14083 ( .IN1(n13503), .IN2(n13504), .QN(g22155) );
  INVX0 U14084 ( .INP(n13505), .ZN(n13504) );
  NOR2X0 U14085 ( .IN1(n13447), .IN2(n7516), .QN(n13505) );
  NAND2X0 U14086 ( .IN1(n13447), .IN2(n10446), .QN(n13503) );
  INVX0 U14087 ( .INP(n9623), .ZN(n10446) );
  NAND3X0 U14088 ( .IN1(n13506), .IN2(n13507), .IN3(n13508), .QN(n9623) );
  NAND2X0 U14089 ( .IN1(n7583), .IN2(test_so73), .QN(n13508) );
  NAND2X0 U14090 ( .IN1(n7584), .IN2(g6837), .QN(n13507) );
  NAND2X0 U14091 ( .IN1(n7582), .IN2(g2241), .QN(n13506) );
  NAND2X0 U14092 ( .IN1(n13509), .IN2(n13510), .QN(g22154) );
  NAND2X0 U14093 ( .IN1(n13432), .IN2(n4287), .QN(n13510) );
  NAND2X0 U14094 ( .IN1(n13433), .IN2(g2234), .QN(n13509) );
  NAND2X0 U14095 ( .IN1(n13511), .IN2(n13512), .QN(g22153) );
  NAND2X0 U14096 ( .IN1(n13045), .IN2(n4563), .QN(n13512) );
  INVX0 U14097 ( .INP(n13513), .ZN(n13511) );
  NOR2X0 U14098 ( .IN1(n13045), .IN2(n7526), .QN(n13513) );
  NAND2X0 U14099 ( .IN1(n13514), .IN2(n13515), .QN(g22152) );
  INVX0 U14100 ( .INP(n13516), .ZN(n13515) );
  NOR2X0 U14101 ( .IN1(n13487), .IN2(n7535), .QN(n13516) );
  NAND2X0 U14102 ( .IN1(n13487), .IN2(n9504), .QN(n13514) );
  INVX0 U14103 ( .INP(n10509), .ZN(n9504) );
  NAND3X0 U14104 ( .IN1(n13517), .IN2(n13518), .IN3(n13519), .QN(n10509) );
  NAND2X0 U14105 ( .IN1(n7597), .IN2(g6782), .QN(n13519) );
  NAND2X0 U14106 ( .IN1(n7598), .IN2(g6573), .QN(n13518) );
  NAND2X0 U14107 ( .IN1(g1547), .IN2(n8141), .QN(n13517) );
  NAND2X0 U14108 ( .IN1(n13520), .IN2(n13521), .QN(g22151) );
  NAND2X0 U14109 ( .IN1(n13457), .IN2(g1543), .QN(n13521) );
  NAND2X0 U14110 ( .IN1(n13483), .IN2(n13456), .QN(n13520) );
  NAND2X0 U14111 ( .IN1(n13522), .IN2(n13523), .QN(g22150) );
  NAND2X0 U14112 ( .IN1(n13048), .IN2(n4288), .QN(n13523) );
  INVX0 U14113 ( .INP(n13524), .ZN(n13522) );
  NOR2X0 U14114 ( .IN1(n13048), .IN2(n7536), .QN(n13524) );
  NAND2X0 U14115 ( .IN1(n13525), .IN2(n13526), .QN(g22149) );
  NAND2X0 U14116 ( .IN1(n13487), .IN2(n4378), .QN(n13526) );
  INVX0 U14117 ( .INP(n13527), .ZN(n13525) );
  NOR2X0 U14118 ( .IN1(n13487), .IN2(n7911), .QN(n13527) );
  NAND2X0 U14119 ( .IN1(n13528), .IN2(n13529), .QN(g22148) );
  INVX0 U14120 ( .INP(n13530), .ZN(n13529) );
  NOR2X0 U14121 ( .IN1(n13495), .IN2(n7545), .QN(n13530) );
  NAND2X0 U14122 ( .IN1(n13495), .IN2(n9537), .QN(n13528) );
  NAND2X0 U14123 ( .IN1(n13531), .IN2(n13532), .QN(g22147) );
  INVX0 U14124 ( .INP(n13533), .ZN(n13532) );
  NOR2X0 U14125 ( .IN1(n13051), .IN2(n7547), .QN(n13533) );
  NAND2X0 U14126 ( .IN1(n10619), .IN2(n13051), .QN(n13531) );
  NAND2X0 U14127 ( .IN1(n13534), .IN2(n13535), .QN(g22146) );
  NAND2X0 U14128 ( .IN1(n13536), .IN2(n4375), .QN(n13535) );
  NAND2X0 U14129 ( .IN1(n13537), .IN2(g821), .QN(n13534) );
  NAND2X0 U14130 ( .IN1(n13538), .IN2(n13539), .QN(g22145) );
  NAND2X0 U14131 ( .IN1(n13495), .IN2(n4379), .QN(n13539) );
  INVX0 U14132 ( .INP(n13540), .ZN(n13538) );
  NOR2X0 U14133 ( .IN1(n13495), .IN2(n7947), .QN(n13540) );
  NAND2X0 U14134 ( .IN1(n13541), .IN2(n13542), .QN(g22143) );
  NAND2X0 U14135 ( .IN1(n13053), .IN2(g162), .QN(n13542) );
  NAND2X0 U14136 ( .IN1(n13502), .IN2(n9582), .QN(n13541) );
  NAND2X0 U14137 ( .IN1(n13543), .IN2(n13544), .QN(g22142) );
  NAND2X0 U14138 ( .IN1(n13545), .IN2(n4376), .QN(n13544) );
  INVX0 U14139 ( .INP(n13546), .ZN(n13543) );
  NOR2X0 U14140 ( .IN1(n13545), .IN2(n7969), .QN(n13546) );
  NAND2X0 U14141 ( .IN1(n13547), .IN2(n13548), .QN(g22141) );
  NAND2X0 U14142 ( .IN1(n4380), .IN2(n13502), .QN(n13548) );
  NAND2X0 U14143 ( .IN1(n13053), .IN2(g129), .QN(n13547) );
  NAND2X0 U14144 ( .IN1(n13549), .IN2(n13550), .QN(g22140) );
  NAND2X0 U14145 ( .IN1(n13447), .IN2(n4287), .QN(n13550) );
  INVX0 U14146 ( .INP(n13551), .ZN(n13549) );
  NOR2X0 U14147 ( .IN1(n13447), .IN2(n7882), .QN(n13551) );
  NAND2X0 U14148 ( .IN1(n13552), .IN2(n13553), .QN(g22139) );
  NAND2X0 U14149 ( .IN1(n13432), .IN2(n4563), .QN(n13553) );
  NAND2X0 U14150 ( .IN1(n13433), .IN2(g2231), .QN(n13552) );
  NAND2X0 U14151 ( .IN1(n13554), .IN2(n13555), .QN(g22138) );
  NAND2X0 U14152 ( .IN1(n13045), .IN2(n4555), .QN(n13555) );
  INVX0 U14153 ( .INP(n13556), .ZN(n13554) );
  NOR2X0 U14154 ( .IN1(n13045), .IN2(n7527), .QN(n13556) );
  NAND2X0 U14155 ( .IN1(n13557), .IN2(n13558), .QN(g22132) );
  INVX0 U14156 ( .INP(n13559), .ZN(n13558) );
  NOR2X0 U14157 ( .IN1(n13487), .IN2(n7519), .QN(n13559) );
  NAND2X0 U14158 ( .IN1(n13487), .IN2(n13483), .QN(n13557) );
  INVX0 U14159 ( .INP(n9660), .ZN(n13483) );
  NAND3X0 U14160 ( .IN1(n13560), .IN2(n13561), .IN3(n13562), .QN(n9660) );
  NAND2X0 U14161 ( .IN1(n7595), .IN2(g6782), .QN(n13562) );
  NAND2X0 U14162 ( .IN1(n7596), .IN2(g6573), .QN(n13561) );
  NAND2X0 U14163 ( .IN1(n7594), .IN2(g1547), .QN(n13560) );
  NAND2X0 U14164 ( .IN1(n13563), .IN2(n13564), .QN(g22131) );
  NAND2X0 U14165 ( .IN1(n13456), .IN2(n4288), .QN(n13564) );
  NAND2X0 U14166 ( .IN1(n13457), .IN2(g1540), .QN(n13563) );
  NAND2X0 U14167 ( .IN1(n13565), .IN2(n13566), .QN(g22130) );
  NAND2X0 U14168 ( .IN1(n13048), .IN2(n4565), .QN(n13566) );
  INVX0 U14169 ( .INP(n13567), .ZN(n13565) );
  NOR2X0 U14170 ( .IN1(n13048), .IN2(n7537), .QN(n13567) );
  NAND2X0 U14171 ( .IN1(n13568), .IN2(n13569), .QN(g22129) );
  NAND2X0 U14172 ( .IN1(n13537), .IN2(g851), .QN(n13569) );
  NAND2X0 U14173 ( .IN1(n13536), .IN2(n9537), .QN(n13568) );
  INVX0 U14174 ( .INP(n10843), .ZN(n9537) );
  NAND3X0 U14175 ( .IN1(n13570), .IN2(n13571), .IN3(n13572), .QN(n10843) );
  NAND2X0 U14176 ( .IN1(n7608), .IN2(test_so31), .QN(n13572) );
  NAND2X0 U14177 ( .IN1(n7609), .IN2(g6518), .QN(n13571) );
  NAND2X0 U14178 ( .IN1(n7610), .IN2(g6368), .QN(n13570) );
  NAND2X0 U14179 ( .IN1(n13573), .IN2(n13574), .QN(g22128) );
  INVX0 U14180 ( .INP(n13575), .ZN(n13574) );
  NOR2X0 U14181 ( .IN1(n13495), .IN2(n7548), .QN(n13575) );
  NAND2X0 U14182 ( .IN1(n10619), .IN2(n13495), .QN(n13573) );
  NAND2X0 U14183 ( .IN1(n13576), .IN2(n13577), .QN(g22127) );
  NAND2X0 U14184 ( .IN1(n4289), .IN2(n13051), .QN(n13577) );
  INVX0 U14185 ( .INP(n13578), .ZN(n13576) );
  NOR2X0 U14186 ( .IN1(n13051), .IN2(n7550), .QN(n13578) );
  NAND2X0 U14187 ( .IN1(n13579), .IN2(n13580), .QN(g22126) );
  NAND2X0 U14188 ( .IN1(n13536), .IN2(n4379), .QN(n13580) );
  NAND2X0 U14189 ( .IN1(n13537), .IN2(g818), .QN(n13579) );
  NAND2X0 U14190 ( .IN1(n13581), .IN2(n13582), .QN(g22125) );
  INVX0 U14191 ( .INP(n13583), .ZN(n13582) );
  NOR2X0 U14192 ( .IN1(n13545), .IN2(n7559), .QN(n13583) );
  NAND2X0 U14193 ( .IN1(n13545), .IN2(n9582), .QN(n13581) );
  NAND2X0 U14194 ( .IN1(n13584), .IN2(n13585), .QN(g22124) );
  NAND2X0 U14195 ( .IN1(n13053), .IN2(g159), .QN(n13585) );
  NAND2X0 U14196 ( .IN1(n12353), .IN2(n13502), .QN(n13584) );
  NAND2X0 U14197 ( .IN1(n13586), .IN2(n13587), .QN(g22123) );
  NAND2X0 U14198 ( .IN1(n13588), .IN2(n4376), .QN(n13587) );
  NAND2X0 U14199 ( .IN1(n13589), .IN2(g133), .QN(n13586) );
  NAND2X0 U14200 ( .IN1(n13590), .IN2(n13591), .QN(g22122) );
  NAND2X0 U14201 ( .IN1(n13545), .IN2(n4380), .QN(n13591) );
  INVX0 U14202 ( .INP(n13592), .ZN(n13590) );
  NOR2X0 U14203 ( .IN1(n13545), .IN2(n7972), .QN(n13592) );
  NAND2X0 U14204 ( .IN1(n13593), .IN2(n13594), .QN(g22117) );
  NAND2X0 U14205 ( .IN1(n13447), .IN2(n4563), .QN(n13594) );
  INVX0 U14206 ( .INP(n13595), .ZN(n13593) );
  NOR2X0 U14207 ( .IN1(n13447), .IN2(n7884), .QN(n13595) );
  NAND2X0 U14208 ( .IN1(n13596), .IN2(n13597), .QN(g22116) );
  NAND2X0 U14209 ( .IN1(n13432), .IN2(n4555), .QN(n13597) );
  NAND2X0 U14210 ( .IN1(n13433), .IN2(g2228), .QN(n13596) );
  NAND2X0 U14211 ( .IN1(n13598), .IN2(n13599), .QN(g22115) );
  NAND2X0 U14212 ( .IN1(n13045), .IN2(n4325), .QN(n13599) );
  INVX0 U14213 ( .INP(n13600), .ZN(n13598) );
  NOR2X0 U14214 ( .IN1(n13045), .IN2(n7528), .QN(n13600) );
  NAND2X0 U14215 ( .IN1(n13601), .IN2(n13602), .QN(g22114) );
  NAND2X0 U14216 ( .IN1(n13487), .IN2(n4288), .QN(n13602) );
  INVX0 U14217 ( .INP(n13603), .ZN(n13601) );
  NOR2X0 U14218 ( .IN1(n13487), .IN2(n7897), .QN(n13603) );
  NAND2X0 U14219 ( .IN1(n13604), .IN2(n13605), .QN(g22113) );
  NAND2X0 U14220 ( .IN1(test_so53), .IN2(n13457), .QN(n13605) );
  NAND2X0 U14221 ( .IN1(n13456), .IN2(n4565), .QN(n13604) );
  NAND2X0 U14222 ( .IN1(n13606), .IN2(n13607), .QN(g22112) );
  NAND2X0 U14223 ( .IN1(n13048), .IN2(n4557), .QN(n13607) );
  INVX0 U14224 ( .INP(n13608), .ZN(n13606) );
  NOR2X0 U14225 ( .IN1(n13048), .IN2(n7538), .QN(n13608) );
  NAND2X0 U14226 ( .IN1(n13609), .IN2(n13610), .QN(g22106) );
  NAND2X0 U14227 ( .IN1(n13537), .IN2(g848), .QN(n13610) );
  NAND2X0 U14228 ( .IN1(n13536), .IN2(n10619), .QN(n13609) );
  INVX0 U14229 ( .INP(n9688), .ZN(n10619) );
  NAND3X0 U14230 ( .IN1(n13611), .IN2(n13612), .IN3(n13613), .QN(n9688) );
  NAND2X0 U14231 ( .IN1(n7605), .IN2(test_so31), .QN(n13613) );
  NAND2X0 U14232 ( .IN1(n7606), .IN2(g6518), .QN(n13612) );
  NAND2X0 U14233 ( .IN1(n7607), .IN2(g6368), .QN(n13611) );
  NAND2X0 U14234 ( .IN1(n13614), .IN2(n13615), .QN(g22105) );
  NAND2X0 U14235 ( .IN1(n4289), .IN2(n13495), .QN(n13615) );
  INVX0 U14236 ( .INP(n13616), .ZN(n13614) );
  NOR2X0 U14237 ( .IN1(n13495), .IN2(n7914), .QN(n13616) );
  NAND2X0 U14238 ( .IN1(n13617), .IN2(n13618), .QN(g22104) );
  NAND2X0 U14239 ( .IN1(n13051), .IN2(n4567), .QN(n13618) );
  INVX0 U14240 ( .INP(n13619), .ZN(n13617) );
  NOR2X0 U14241 ( .IN1(n13051), .IN2(n7551), .QN(n13619) );
  NAND2X0 U14242 ( .IN1(n13620), .IN2(n13621), .QN(g22103) );
  NAND2X0 U14243 ( .IN1(test_so12), .IN2(n13589), .QN(n13621) );
  NAND2X0 U14244 ( .IN1(n13588), .IN2(n9582), .QN(n13620) );
  INVX0 U14245 ( .INP(n10712), .ZN(n9582) );
  NAND3X0 U14246 ( .IN1(n13622), .IN2(n13623), .IN3(n13624), .QN(n10712) );
  NAND2X0 U14247 ( .IN1(n7620), .IN2(g6313), .QN(n13624) );
  NAND2X0 U14248 ( .IN1(n7621), .IN2(g6231), .QN(n13623) );
  NAND2X0 U14249 ( .IN1(n7619), .IN2(g165), .QN(n13622) );
  NAND2X0 U14250 ( .IN1(n13625), .IN2(n13626), .QN(g22102) );
  INVX0 U14251 ( .INP(n13627), .ZN(n13626) );
  NOR2X0 U14252 ( .IN1(n13545), .IN2(n7521), .QN(n13627) );
  NAND2X0 U14253 ( .IN1(n12353), .IN2(n13545), .QN(n13625) );
  NAND2X0 U14254 ( .IN1(n13628), .IN2(n13629), .QN(g22101) );
  NAND2X0 U14255 ( .IN1(n4290), .IN2(n13502), .QN(n13629) );
  NAND2X0 U14256 ( .IN1(n13053), .IN2(g156), .QN(n13628) );
  NAND2X0 U14257 ( .IN1(n13630), .IN2(n13631), .QN(g22100) );
  NAND2X0 U14258 ( .IN1(n13588), .IN2(n4380), .QN(n13631) );
  NAND2X0 U14259 ( .IN1(n13589), .IN2(g130), .QN(n13630) );
  NAND2X0 U14260 ( .IN1(n13632), .IN2(n13633), .QN(g22099) );
  NAND2X0 U14261 ( .IN1(n13447), .IN2(n4555), .QN(n13633) );
  INVX0 U14262 ( .INP(n13634), .ZN(n13632) );
  NOR2X0 U14263 ( .IN1(n13447), .IN2(n7886), .QN(n13634) );
  NAND2X0 U14264 ( .IN1(n13635), .IN2(n13636), .QN(g22098) );
  NAND2X0 U14265 ( .IN1(test_so74), .IN2(n13433), .QN(n13636) );
  NAND2X0 U14266 ( .IN1(n13432), .IN2(n4325), .QN(n13635) );
  NAND2X0 U14267 ( .IN1(n13637), .IN2(n13638), .QN(g22097) );
  NAND2X0 U14268 ( .IN1(n13045), .IN2(n4389), .QN(n13638) );
  INVX0 U14269 ( .INP(n13639), .ZN(n13637) );
  NOR2X0 U14270 ( .IN1(n13045), .IN2(n7529), .QN(n13639) );
  NAND2X0 U14271 ( .IN1(n13640), .IN2(n13641), .QN(g22092) );
  NAND2X0 U14272 ( .IN1(n13487), .IN2(n4565), .QN(n13641) );
  INVX0 U14273 ( .INP(n13642), .ZN(n13640) );
  NOR2X0 U14274 ( .IN1(n13487), .IN2(n7898), .QN(n13642) );
  NAND2X0 U14275 ( .IN1(n13643), .IN2(n13644), .QN(g22091) );
  NAND2X0 U14276 ( .IN1(n13456), .IN2(n4557), .QN(n13644) );
  NAND2X0 U14277 ( .IN1(n13457), .IN2(g1534), .QN(n13643) );
  NAND2X0 U14278 ( .IN1(n13645), .IN2(n13646), .QN(g22090) );
  NAND2X0 U14279 ( .IN1(n13048), .IN2(n4326), .QN(n13646) );
  INVX0 U14280 ( .INP(n13647), .ZN(n13645) );
  NOR2X0 U14281 ( .IN1(n13048), .IN2(n7539), .QN(n13647) );
  NAND2X0 U14282 ( .IN1(n13648), .IN2(n13649), .QN(g22089) );
  NAND2X0 U14283 ( .IN1(n4289), .IN2(n13536), .QN(n13649) );
  NAND2X0 U14284 ( .IN1(n13537), .IN2(g845), .QN(n13648) );
  NAND2X0 U14285 ( .IN1(n13650), .IN2(n13651), .QN(g22088) );
  NAND2X0 U14286 ( .IN1(n13495), .IN2(n4567), .QN(n13651) );
  INVX0 U14287 ( .INP(n13652), .ZN(n13650) );
  NOR2X0 U14288 ( .IN1(n13495), .IN2(n7916), .QN(n13652) );
  NAND2X0 U14289 ( .IN1(n13653), .IN2(n13654), .QN(g22087) );
  NAND2X0 U14290 ( .IN1(n13051), .IN2(n4559), .QN(n13654) );
  INVX0 U14291 ( .INP(n13655), .ZN(n13653) );
  NOR2X0 U14292 ( .IN1(n13051), .IN2(n7552), .QN(n13655) );
  NAND2X0 U14293 ( .IN1(n13656), .IN2(n13657), .QN(g22081) );
  NAND2X0 U14294 ( .IN1(n13589), .IN2(g160), .QN(n13657) );
  NAND2X0 U14295 ( .IN1(n13588), .IN2(n12353), .QN(n13656) );
  INVX0 U14296 ( .INP(n9709), .ZN(n12353) );
  NAND3X0 U14297 ( .IN1(n13658), .IN2(n13659), .IN3(n13660), .QN(n9709) );
  NAND2X0 U14298 ( .IN1(n7617), .IN2(g6313), .QN(n13660) );
  NAND2X0 U14299 ( .IN1(n7618), .IN2(g6231), .QN(n13659) );
  NAND2X0 U14300 ( .IN1(n7616), .IN2(g165), .QN(n13658) );
  NAND2X0 U14301 ( .IN1(n13661), .IN2(n13662), .QN(g22080) );
  NAND2X0 U14302 ( .IN1(n4290), .IN2(n13545), .QN(n13662) );
  INVX0 U14303 ( .INP(n13663), .ZN(n13661) );
  NOR2X0 U14304 ( .IN1(n13545), .IN2(n7949), .QN(n13663) );
  NAND2X0 U14305 ( .IN1(n13664), .IN2(n13665), .QN(g22079) );
  NAND2X0 U14306 ( .IN1(n13502), .IN2(n4569), .QN(n13665) );
  NAND2X0 U14307 ( .IN1(n13053), .IN2(g153), .QN(n13664) );
  NAND2X0 U14308 ( .IN1(n13666), .IN2(n13667), .QN(g22078) );
  NAND2X0 U14309 ( .IN1(n13447), .IN2(n4325), .QN(n13667) );
  INVX0 U14310 ( .INP(n13668), .ZN(n13666) );
  NOR2X0 U14311 ( .IN1(n13447), .IN2(n7887), .QN(n13668) );
  NAND2X0 U14312 ( .IN1(n13669), .IN2(n13670), .QN(g22077) );
  NAND2X0 U14313 ( .IN1(n13432), .IN2(n4389), .QN(n13670) );
  NAND2X0 U14314 ( .IN1(n13433), .IN2(g2222), .QN(n13669) );
  NAND2X0 U14315 ( .IN1(n13671), .IN2(n13672), .QN(g22076) );
  NAND2X0 U14316 ( .IN1(n13045), .IN2(n4319), .QN(n13672) );
  INVX0 U14317 ( .INP(n13673), .ZN(n13671) );
  NOR2X0 U14318 ( .IN1(n13045), .IN2(n7530), .QN(n13673) );
  NOR2X0 U14319 ( .IN1(n4367), .IN2(n7718), .QN(n13045) );
  NAND2X0 U14320 ( .IN1(n13674), .IN2(n13675), .QN(g22075) );
  NAND2X0 U14321 ( .IN1(n13487), .IN2(n4557), .QN(n13675) );
  INVX0 U14322 ( .INP(n13676), .ZN(n13674) );
  NOR2X0 U14323 ( .IN1(n13487), .IN2(n7900), .QN(n13676) );
  NAND2X0 U14324 ( .IN1(n13677), .IN2(n13678), .QN(g22074) );
  NAND2X0 U14325 ( .IN1(n13456), .IN2(n4326), .QN(n13678) );
  NAND2X0 U14326 ( .IN1(n13457), .IN2(g1531), .QN(n13677) );
  NAND2X0 U14327 ( .IN1(n13679), .IN2(n13680), .QN(g22073) );
  NAND2X0 U14328 ( .IN1(n13048), .IN2(n4390), .QN(n13680) );
  INVX0 U14329 ( .INP(n13681), .ZN(n13679) );
  NOR2X0 U14330 ( .IN1(n13048), .IN2(n7540), .QN(n13681) );
  NAND2X0 U14331 ( .IN1(n13682), .IN2(n13683), .QN(g22068) );
  NAND2X0 U14332 ( .IN1(n13536), .IN2(n4567), .QN(n13683) );
  NAND2X0 U14333 ( .IN1(n13537), .IN2(g842), .QN(n13682) );
  NAND2X0 U14334 ( .IN1(n13684), .IN2(n13685), .QN(g22067) );
  NAND2X0 U14335 ( .IN1(n13495), .IN2(n4559), .QN(n13685) );
  INVX0 U14336 ( .INP(n13686), .ZN(n13684) );
  NOR2X0 U14337 ( .IN1(n13495), .IN2(n7919), .QN(n13686) );
  NAND2X0 U14338 ( .IN1(n13687), .IN2(n13688), .QN(g22066) );
  NAND2X0 U14339 ( .IN1(n4327), .IN2(n13051), .QN(n13688) );
  INVX0 U14340 ( .INP(n13689), .ZN(n13687) );
  NOR2X0 U14341 ( .IN1(n13051), .IN2(n7553), .QN(n13689) );
  NAND2X0 U14342 ( .IN1(n13690), .IN2(n13691), .QN(g22065) );
  NAND2X0 U14343 ( .IN1(n4290), .IN2(n13588), .QN(n13691) );
  NAND2X0 U14344 ( .IN1(n13589), .IN2(g157), .QN(n13690) );
  NAND2X0 U14345 ( .IN1(n13692), .IN2(n13693), .QN(g22064) );
  NAND2X0 U14346 ( .IN1(n13545), .IN2(n4569), .QN(n13693) );
  INVX0 U14347 ( .INP(n13694), .ZN(n13692) );
  NOR2X0 U14348 ( .IN1(n13545), .IN2(n7951), .QN(n13694) );
  NAND2X0 U14349 ( .IN1(n13695), .IN2(n13696), .QN(g22063) );
  NAND2X0 U14350 ( .IN1(n13502), .IN2(n4561), .QN(n13696) );
  NAND2X0 U14351 ( .IN1(n13053), .IN2(g150), .QN(n13695) );
  NAND2X0 U14352 ( .IN1(n13697), .IN2(n13698), .QN(g22061) );
  NAND2X0 U14353 ( .IN1(n13447), .IN2(n4389), .QN(n13698) );
  INVX0 U14354 ( .INP(n13699), .ZN(n13697) );
  NOR2X0 U14355 ( .IN1(n13447), .IN2(n7889), .QN(n13699) );
  NAND2X0 U14356 ( .IN1(n13700), .IN2(n13701), .QN(g22060) );
  NAND2X0 U14357 ( .IN1(n13432), .IN2(n4319), .QN(n13701) );
  NAND2X0 U14358 ( .IN1(n13433), .IN2(g2219), .QN(n13700) );
  INVX0 U14359 ( .INP(n13432), .ZN(n13433) );
  NOR2X0 U14360 ( .IN1(n8097), .IN2(n7718), .QN(n13432) );
  NAND2X0 U14361 ( .IN1(n13702), .IN2(n13703), .QN(g22059) );
  NAND2X0 U14362 ( .IN1(n13487), .IN2(n4326), .QN(n13703) );
  INVX0 U14363 ( .INP(n13704), .ZN(n13702) );
  NOR2X0 U14364 ( .IN1(n13487), .IN2(n7902), .QN(n13704) );
  NAND2X0 U14365 ( .IN1(n13705), .IN2(n13706), .QN(g22058) );
  NAND2X0 U14366 ( .IN1(n13456), .IN2(n4390), .QN(n13706) );
  NAND2X0 U14367 ( .IN1(n13457), .IN2(g1528), .QN(n13705) );
  NAND2X0 U14368 ( .IN1(n13707), .IN2(n13708), .QN(g22057) );
  NAND2X0 U14369 ( .IN1(n13048), .IN2(n4320), .QN(n13708) );
  INVX0 U14370 ( .INP(n13709), .ZN(n13707) );
  NOR2X0 U14371 ( .IN1(n13048), .IN2(n7541), .QN(n13709) );
  NOR2X0 U14372 ( .IN1(n4368), .IN2(n7719), .QN(n13048) );
  NAND2X0 U14373 ( .IN1(n13710), .IN2(n13711), .QN(g22056) );
  NAND2X0 U14374 ( .IN1(test_so32), .IN2(n13537), .QN(n13711) );
  NAND2X0 U14375 ( .IN1(n13536), .IN2(n4559), .QN(n13710) );
  NAND2X0 U14376 ( .IN1(n13712), .IN2(n13713), .QN(g22055) );
  NAND2X0 U14377 ( .IN1(n4327), .IN2(n13495), .QN(n13713) );
  INVX0 U14378 ( .INP(n13714), .ZN(n13712) );
  NOR2X0 U14379 ( .IN1(n13495), .IN2(n7927), .QN(n13714) );
  NAND2X0 U14380 ( .IN1(n13715), .IN2(n13716), .QN(g22054) );
  NAND2X0 U14381 ( .IN1(n13051), .IN2(n4391), .QN(n13716) );
  INVX0 U14382 ( .INP(n13717), .ZN(n13715) );
  NOR2X0 U14383 ( .IN1(n13051), .IN2(n7554), .QN(n13717) );
  NAND2X0 U14384 ( .IN1(n13718), .IN2(n13719), .QN(g22049) );
  NAND2X0 U14385 ( .IN1(n13588), .IN2(n4569), .QN(n13719) );
  NAND2X0 U14386 ( .IN1(n13589), .IN2(g154), .QN(n13718) );
  NAND2X0 U14387 ( .IN1(n13720), .IN2(n13721), .QN(g22048) );
  NAND2X0 U14388 ( .IN1(n13545), .IN2(n4561), .QN(n13721) );
  INVX0 U14389 ( .INP(n13722), .ZN(n13720) );
  NOR2X0 U14390 ( .IN1(n13545), .IN2(n7953), .QN(n13722) );
  NAND2X0 U14391 ( .IN1(n13723), .IN2(n13724), .QN(g22047) );
  NAND2X0 U14392 ( .IN1(n4328), .IN2(n13502), .QN(n13724) );
  NAND2X0 U14393 ( .IN1(n13053), .IN2(g147), .QN(n13723) );
  NAND2X0 U14394 ( .IN1(n13725), .IN2(n13726), .QN(g22045) );
  NAND2X0 U14395 ( .IN1(n13447), .IN2(n4319), .QN(n13726) );
  INVX0 U14396 ( .INP(n13727), .ZN(n13725) );
  NOR2X0 U14397 ( .IN1(n13447), .IN2(n7891), .QN(n13727) );
  NOR2X0 U14398 ( .IN1(n4324), .IN2(n7718), .QN(n13447) );
  NAND2X0 U14399 ( .IN1(n13728), .IN2(n13729), .QN(g22044) );
  NAND2X0 U14400 ( .IN1(n13487), .IN2(n4390), .QN(n13729) );
  INVX0 U14401 ( .INP(n13730), .ZN(n13728) );
  NOR2X0 U14402 ( .IN1(n13487), .IN2(n7904), .QN(n13730) );
  NAND2X0 U14403 ( .IN1(n13731), .IN2(n13732), .QN(g22043) );
  NAND2X0 U14404 ( .IN1(n13456), .IN2(n4320), .QN(n13732) );
  NAND2X0 U14405 ( .IN1(n13457), .IN2(g1525), .QN(n13731) );
  INVX0 U14406 ( .INP(n13456), .ZN(n13457) );
  NOR2X0 U14407 ( .IN1(n4515), .IN2(n7719), .QN(n13456) );
  NAND2X0 U14408 ( .IN1(n13733), .IN2(n13734), .QN(g22042) );
  NAND2X0 U14409 ( .IN1(n4327), .IN2(n13536), .QN(n13734) );
  NAND2X0 U14410 ( .IN1(n13537), .IN2(g836), .QN(n13733) );
  NAND2X0 U14411 ( .IN1(n13735), .IN2(n13736), .QN(g22041) );
  NAND2X0 U14412 ( .IN1(n13495), .IN2(n4391), .QN(n13736) );
  INVX0 U14413 ( .INP(n13737), .ZN(n13735) );
  NOR2X0 U14414 ( .IN1(n13495), .IN2(n7931), .QN(n13737) );
  NAND2X0 U14415 ( .IN1(n13738), .IN2(n13739), .QN(g22040) );
  NAND2X0 U14416 ( .IN1(n4321), .IN2(n13051), .QN(n13739) );
  INVX0 U14417 ( .INP(n13740), .ZN(n13738) );
  NOR2X0 U14418 ( .IN1(n13051), .IN2(n7555), .QN(n13740) );
  NOR2X0 U14419 ( .IN1(n8096), .IN2(n7720), .QN(n13051) );
  NAND2X0 U14420 ( .IN1(n13741), .IN2(n13742), .QN(g22039) );
  NAND2X0 U14421 ( .IN1(n13588), .IN2(n4561), .QN(n13742) );
  NAND2X0 U14422 ( .IN1(n13589), .IN2(g151), .QN(n13741) );
  NAND2X0 U14423 ( .IN1(n13743), .IN2(n13744), .QN(g22038) );
  NAND2X0 U14424 ( .IN1(n4328), .IN2(n13545), .QN(n13744) );
  INVX0 U14425 ( .INP(n13745), .ZN(n13743) );
  NOR2X0 U14426 ( .IN1(n13545), .IN2(n7955), .QN(n13745) );
  NAND2X0 U14427 ( .IN1(n13746), .IN2(n13747), .QN(g22037) );
  NAND2X0 U14428 ( .IN1(test_so11), .IN2(n13053), .QN(n13747) );
  NAND2X0 U14429 ( .IN1(n13502), .IN2(n4392), .QN(n13746) );
  NAND2X0 U14430 ( .IN1(n13748), .IN2(n13749), .QN(g22035) );
  NAND2X0 U14431 ( .IN1(n13487), .IN2(n4320), .QN(n13749) );
  INVX0 U14432 ( .INP(n13750), .ZN(n13748) );
  NOR2X0 U14433 ( .IN1(n13487), .IN2(n7906), .QN(n13750) );
  NOR2X0 U14434 ( .IN1(n4317), .IN2(n7719), .QN(n13487) );
  NAND2X0 U14435 ( .IN1(n13751), .IN2(n13752), .QN(g22034) );
  NAND2X0 U14436 ( .IN1(n13536), .IN2(n4391), .QN(n13752) );
  NAND2X0 U14437 ( .IN1(n13537), .IN2(g833), .QN(n13751) );
  NAND2X0 U14438 ( .IN1(n13753), .IN2(n13754), .QN(g22033) );
  NAND2X0 U14439 ( .IN1(n4321), .IN2(n13495), .QN(n13754) );
  INVX0 U14440 ( .INP(n13755), .ZN(n13753) );
  NOR2X0 U14441 ( .IN1(n13495), .IN2(n7933), .QN(n13755) );
  NOR2X0 U14442 ( .IN1(n4312), .IN2(n7720), .QN(n13495) );
  NAND2X0 U14443 ( .IN1(n13756), .IN2(n13757), .QN(g22032) );
  NAND2X0 U14444 ( .IN1(n4328), .IN2(n13588), .QN(n13757) );
  NAND2X0 U14445 ( .IN1(n13589), .IN2(g148), .QN(n13756) );
  NAND2X0 U14446 ( .IN1(n13758), .IN2(n13759), .QN(g22031) );
  NAND2X0 U14447 ( .IN1(n13545), .IN2(n4392), .QN(n13759) );
  INVX0 U14448 ( .INP(n13760), .ZN(n13758) );
  NOR2X0 U14449 ( .IN1(n13545), .IN2(n7957), .QN(n13760) );
  NAND2X0 U14450 ( .IN1(n13761), .IN2(n13762), .QN(g22030) );
  NAND2X0 U14451 ( .IN1(n4322), .IN2(n13502), .QN(n13762) );
  NAND2X0 U14452 ( .IN1(n13053), .IN2(g141), .QN(n13761) );
  INVX0 U14453 ( .INP(n13502), .ZN(n13053) );
  NOR2X0 U14454 ( .IN1(n4369), .IN2(n7721), .QN(n13502) );
  NAND2X0 U14455 ( .IN1(n13763), .IN2(n13764), .QN(g22029) );
  NAND2X0 U14456 ( .IN1(n4321), .IN2(n13536), .QN(n13764) );
  NAND2X0 U14457 ( .IN1(n13537), .IN2(g830), .QN(n13763) );
  INVX0 U14458 ( .INP(n13536), .ZN(n13537) );
  NOR2X0 U14459 ( .IN1(n4323), .IN2(n7720), .QN(n13536) );
  NAND2X0 U14460 ( .IN1(n13765), .IN2(n13766), .QN(g22028) );
  NAND2X0 U14461 ( .IN1(n13588), .IN2(n4392), .QN(n13766) );
  NAND2X0 U14462 ( .IN1(n13589), .IN2(g145), .QN(n13765) );
  NAND2X0 U14463 ( .IN1(n13767), .IN2(n13768), .QN(g22027) );
  NAND2X0 U14464 ( .IN1(n4322), .IN2(n13545), .QN(n13768) );
  INVX0 U14465 ( .INP(n13769), .ZN(n13767) );
  NOR2X0 U14466 ( .IN1(n13545), .IN2(n7959), .QN(n13769) );
  NOR2X0 U14467 ( .IN1(n4512), .IN2(n7721), .QN(n13545) );
  NOR2X0 U14468 ( .IN1(n8685), .IN2(n13770), .QN(g22026) );
  XOR2X1 U14469 ( .IN1(n8037), .IN2(n13297), .Q(n13770) );
  NOR2X0 U14470 ( .IN1(n4423), .IN2(n4330), .QN(n13297) );
  NAND2X0 U14471 ( .IN1(n14383), .IN2(n8690), .QN(n8685) );
  NAND4X0 U14472 ( .IN1(n4182), .IN2(n4431), .IN3(n4330), .IN4(n13771), .QN(
        n8690) );
  NOR4X0 U14473 ( .IN1(n8037), .IN2(n4423), .IN3(n4355), .IN4(g2900), .QN(
        n13771) );
  NAND2X0 U14474 ( .IN1(n13772), .IN2(n13773), .QN(g22025) );
  NAND2X0 U14475 ( .IN1(n4322), .IN2(n13588), .QN(n13773) );
  NAND2X0 U14476 ( .IN1(n13589), .IN2(g142), .QN(n13772) );
  INVX0 U14477 ( .INP(n13588), .ZN(n13589) );
  NOR2X0 U14478 ( .IN1(n4318), .IN2(n7721), .QN(n13588) );
  NAND2X0 U14479 ( .IN1(n13774), .IN2(n13775), .QN(g21970) );
  NAND2X0 U14480 ( .IN1(test_so87), .IN2(n4463), .QN(n13775) );
  NAND2X0 U14481 ( .IN1(n11347), .IN2(g2560), .QN(n13774) );
  NAND3X0 U14482 ( .IN1(n13776), .IN2(n13777), .IN3(n13778), .QN(n11347) );
  NAND2X0 U14483 ( .IN1(g5555), .IN2(g2513), .QN(n13778) );
  NAND2X0 U14484 ( .IN1(n4606), .IN2(g2519), .QN(n13777) );
  NAND2X0 U14485 ( .IN1(g7264), .IN2(g2516), .QN(n13776) );
  NAND2X0 U14486 ( .IN1(n13779), .IN2(n13780), .QN(g21882) );
  NAND2X0 U14487 ( .IN1(n4351), .IN2(g2878), .QN(n13780) );
  NAND2X0 U14488 ( .IN1(n13781), .IN2(g2879), .QN(n13779) );
  NAND2X0 U14489 ( .IN1(n13782), .IN2(n13783), .QN(g21880) );
  NAND2X0 U14490 ( .IN1(n4351), .IN2(g2877), .QN(n13783) );
  NAND2X0 U14491 ( .IN1(n13784), .IN2(g2879), .QN(n13782) );
  NAND2X0 U14492 ( .IN1(n13785), .IN2(n13786), .QN(g21878) );
  NAND2X0 U14493 ( .IN1(test_so4), .IN2(g2879), .QN(n13786) );
  NAND2X0 U14494 ( .IN1(n13781), .IN2(n4351), .QN(n13785) );
  XNOR2X1 U14495 ( .IN1(n8561), .IN2(n13787), .Q(n13781) );
  XOR3X1 U14496 ( .IN1(n13788), .IN2(n13789), .IN3(n13790), .Q(n8561) );
  XOR3X1 U14497 ( .IN1(n8023), .IN2(n8022), .IN3(n13791), .Q(n13790) );
  XOR2X1 U14498 ( .IN1(g2981), .IN2(test_so2), .Q(n13791) );
  XOR2X1 U14499 ( .IN1(n8014), .IN2(n8013), .Q(n13789) );
  XOR2X1 U14500 ( .IN1(n8016), .IN2(n8015), .Q(n13788) );
  NAND2X0 U14501 ( .IN1(n13792), .IN2(n13793), .QN(g21851) );
  NAND2X0 U14502 ( .IN1(g499), .IN2(g544), .QN(n13793) );
  NAND3X0 U14503 ( .IN1(n4298), .IN2(g548), .IN3(n4541), .QN(n13792) );
  NAND2X0 U14504 ( .IN1(n13794), .IN2(n13795), .QN(g21346) );
  NAND2X0 U14505 ( .IN1(n14388), .IN2(DFF_328_n1), .QN(n13795) );
  INVX0 U14506 ( .INP(n13796), .ZN(n13794) );
  NOR3X0 U14507 ( .IN1(g6447), .IN2(n7445), .IN3(n14388), .QN(n13796) );
  NAND2X0 U14508 ( .IN1(n13797), .IN2(n13798), .QN(g21094) );
  NAND2X0 U14509 ( .IN1(test_so94), .IN2(n12605), .QN(n13798) );
  NAND2X0 U14510 ( .IN1(n4393), .IN2(n12607), .QN(n13797) );
  NAND2X0 U14511 ( .IN1(n13799), .IN2(n13800), .QN(g21082) );
  NAND2X0 U14512 ( .IN1(n4393), .IN2(n12611), .QN(n13800) );
  NAND2X0 U14513 ( .IN1(n12610), .IN2(g2798), .QN(n13799) );
  NAND2X0 U14514 ( .IN1(n13801), .IN2(n13802), .QN(g21081) );
  NAND2X0 U14515 ( .IN1(n12607), .IN2(n4471), .QN(n13802) );
  NAND2X0 U14516 ( .IN1(n12605), .IN2(g2793), .QN(n13801) );
  NAND2X0 U14517 ( .IN1(n13803), .IN2(n13804), .QN(g21080) );
  NAND2X0 U14518 ( .IN1(n12616), .IN2(n8106), .QN(n13804) );
  NAND2X0 U14519 ( .IN1(n12614), .IN2(g2102), .QN(n13803) );
  NAND2X0 U14520 ( .IN1(n13805), .IN2(n13806), .QN(g21075) );
  NAND2X0 U14521 ( .IN1(n4393), .IN2(n12620), .QN(n13806) );
  NAND2X0 U14522 ( .IN1(n12619), .IN2(g2797), .QN(n13805) );
  NAND2X0 U14523 ( .IN1(n13807), .IN2(n13808), .QN(g21074) );
  NAND2X0 U14524 ( .IN1(n12611), .IN2(n4471), .QN(n13808) );
  NAND2X0 U14525 ( .IN1(n12610), .IN2(g2795), .QN(n13807) );
  NAND2X0 U14526 ( .IN1(n13809), .IN2(n13810), .QN(g21073) );
  NAND2X0 U14527 ( .IN1(n12607), .IN2(n8101), .QN(n13810) );
  NAND2X0 U14528 ( .IN1(n12605), .IN2(g2790), .QN(n13809) );
  NAND2X0 U14529 ( .IN1(n13811), .IN2(n13812), .QN(g21072) );
  NAND2X0 U14530 ( .IN1(n12676), .IN2(n8106), .QN(n13812) );
  NAND2X0 U14531 ( .IN1(n9335), .IN2(g2104), .QN(n13811) );
  NAND2X0 U14532 ( .IN1(n13813), .IN2(n13814), .QN(g21071) );
  NAND2X0 U14533 ( .IN1(n12616), .IN2(n4473), .QN(n13814) );
  NAND2X0 U14534 ( .IN1(n12614), .IN2(g2099), .QN(n13813) );
  NAND2X0 U14535 ( .IN1(n13815), .IN2(n13816), .QN(g21070) );
  NAND2X0 U14536 ( .IN1(n4395), .IN2(n12680), .QN(n13816) );
  INVX0 U14537 ( .INP(n13817), .ZN(n13815) );
  NOR2X0 U14538 ( .IN1(n12680), .IN2(n7858), .QN(n13817) );
  NAND2X0 U14539 ( .IN1(n13818), .IN2(n13819), .QN(g21063) );
  NAND2X0 U14540 ( .IN1(n13820), .IN2(g2805), .QN(n13819) );
  NAND2X0 U14541 ( .IN1(n13402), .IN2(n13821), .QN(n13818) );
  NAND2X0 U14542 ( .IN1(n13822), .IN2(n13823), .QN(g21062) );
  NAND2X0 U14543 ( .IN1(n12620), .IN2(n4471), .QN(n13823) );
  NAND2X0 U14544 ( .IN1(n12619), .IN2(g2794), .QN(n13822) );
  NAND2X0 U14545 ( .IN1(n13824), .IN2(n13825), .QN(g21061) );
  NAND2X0 U14546 ( .IN1(n12611), .IN2(n8101), .QN(n13825) );
  NAND2X0 U14547 ( .IN1(n12610), .IN2(g2792), .QN(n13824) );
  NAND2X0 U14548 ( .IN1(n13826), .IN2(n13827), .QN(g21060) );
  NAND2X0 U14549 ( .IN1(n12607), .IN2(n4407), .QN(n13827) );
  NAND2X0 U14550 ( .IN1(n12605), .IN2(g2787), .QN(n13826) );
  NAND2X0 U14551 ( .IN1(n13828), .IN2(n13829), .QN(g21056) );
  NAND2X0 U14552 ( .IN1(n12685), .IN2(n8106), .QN(n13829) );
  NAND2X0 U14553 ( .IN1(n12684), .IN2(g2103), .QN(n13828) );
  NAND2X0 U14554 ( .IN1(n13830), .IN2(n13831), .QN(g21055) );
  NAND2X0 U14555 ( .IN1(n12676), .IN2(n4473), .QN(n13831) );
  NAND2X0 U14556 ( .IN1(n9335), .IN2(g2101), .QN(n13830) );
  NAND2X0 U14557 ( .IN1(n13832), .IN2(n13833), .QN(g21054) );
  NAND2X0 U14558 ( .IN1(n4468), .IN2(n12616), .QN(n13833) );
  NAND2X0 U14559 ( .IN1(n12614), .IN2(g2096), .QN(n13832) );
  NAND2X0 U14560 ( .IN1(n13834), .IN2(n13835), .QN(g21053) );
  NAND2X0 U14561 ( .IN1(n4395), .IN2(n12741), .QN(n13835) );
  NAND2X0 U14562 ( .IN1(n8530), .IN2(g1410), .QN(n13834) );
  NAND2X0 U14563 ( .IN1(n13836), .IN2(n13837), .QN(g21052) );
  NAND2X0 U14564 ( .IN1(n12680), .IN2(n4475), .QN(n13837) );
  INVX0 U14565 ( .INP(n13838), .ZN(n13836) );
  NOR2X0 U14566 ( .IN1(n12680), .IN2(n7859), .QN(n13838) );
  NAND2X0 U14567 ( .IN1(n13839), .IN2(n13840), .QN(g21051) );
  NAND2X0 U14568 ( .IN1(n4396), .IN2(n12746), .QN(n13840) );
  NAND2X0 U14569 ( .IN1(n12744), .IN2(g722), .QN(n13839) );
  NAND2X0 U14570 ( .IN1(n13841), .IN2(n13842), .QN(g21047) );
  NAND2X0 U14571 ( .IN1(n9306), .IN2(g2807), .QN(n13842) );
  NAND2X0 U14572 ( .IN1(n11309), .IN2(n13821), .QN(n13841) );
  NAND2X0 U14573 ( .IN1(n13843), .IN2(n13844), .QN(g21046) );
  NAND2X0 U14574 ( .IN1(n13820), .IN2(g2802), .QN(n13844) );
  NAND2X0 U14575 ( .IN1(n13402), .IN2(n8912), .QN(n13843) );
  INVX0 U14576 ( .INP(n13820), .ZN(n13402) );
  NAND2X0 U14577 ( .IN1(g2703), .IN2(g2704), .QN(n13820) );
  NAND2X0 U14578 ( .IN1(n13845), .IN2(n13846), .QN(g21045) );
  NAND2X0 U14579 ( .IN1(n12620), .IN2(n8101), .QN(n13846) );
  NAND2X0 U14580 ( .IN1(n12619), .IN2(g2791), .QN(n13845) );
  NAND2X0 U14581 ( .IN1(n13847), .IN2(n13848), .QN(g21044) );
  NAND2X0 U14582 ( .IN1(n12611), .IN2(n4407), .QN(n13848) );
  NAND2X0 U14583 ( .IN1(n12610), .IN2(g2789), .QN(n13847) );
  NAND2X0 U14584 ( .IN1(n13849), .IN2(n13850), .QN(g21043) );
  NAND2X0 U14585 ( .IN1(n4397), .IN2(n12607), .QN(n13850) );
  NAND2X0 U14586 ( .IN1(n12605), .IN2(g2784), .QN(n13849) );
  NAND2X0 U14587 ( .IN1(n13851), .IN2(n13852), .QN(g21042) );
  NAND2X0 U14588 ( .IN1(n13853), .IN2(g2111), .QN(n13852) );
  NAND2X0 U14589 ( .IN1(n13406), .IN2(n13854), .QN(n13851) );
  NAND2X0 U14590 ( .IN1(n13855), .IN2(n13856), .QN(g21041) );
  NAND2X0 U14591 ( .IN1(n12685), .IN2(n4473), .QN(n13856) );
  NAND2X0 U14592 ( .IN1(n12684), .IN2(g2100), .QN(n13855) );
  NAND2X0 U14593 ( .IN1(n13857), .IN2(n13858), .QN(g21040) );
  NAND2X0 U14594 ( .IN1(n4468), .IN2(n12676), .QN(n13858) );
  NAND2X0 U14595 ( .IN1(n9335), .IN2(g2098), .QN(n13857) );
  NAND2X0 U14596 ( .IN1(n13859), .IN2(n13860), .QN(g21039) );
  NAND2X0 U14597 ( .IN1(n12616), .IN2(n4409), .QN(n13860) );
  NAND2X0 U14598 ( .IN1(n12614), .IN2(g2093), .QN(n13859) );
  NAND2X0 U14599 ( .IN1(n13861), .IN2(n13862), .QN(g21035) );
  NAND2X0 U14600 ( .IN1(n4395), .IN2(n12753), .QN(n13862) );
  NAND2X0 U14601 ( .IN1(n12752), .IN2(g1409), .QN(n13861) );
  NAND2X0 U14602 ( .IN1(n13863), .IN2(n13864), .QN(g21034) );
  NAND2X0 U14603 ( .IN1(n12741), .IN2(n4475), .QN(n13864) );
  NAND2X0 U14604 ( .IN1(n8530), .IN2(g1407), .QN(n13863) );
  NAND2X0 U14605 ( .IN1(n13865), .IN2(n13866), .QN(g21033) );
  NAND2X0 U14606 ( .IN1(n4469), .IN2(n12680), .QN(n13866) );
  INVX0 U14607 ( .INP(n13867), .ZN(n13865) );
  NOR2X0 U14608 ( .IN1(n12680), .IN2(n7860), .QN(n13867) );
  NAND2X0 U14609 ( .IN1(n13868), .IN2(n13869), .QN(g21032) );
  NAND2X0 U14610 ( .IN1(n4396), .IN2(n12809), .QN(n13869) );
  NAND2X0 U14611 ( .IN1(n8551), .IN2(g724), .QN(n13868) );
  NAND2X0 U14612 ( .IN1(n13870), .IN2(n13871), .QN(g21031) );
  NAND2X0 U14613 ( .IN1(n12746), .IN2(n4477), .QN(n13871) );
  NAND2X0 U14614 ( .IN1(n12744), .IN2(g719), .QN(n13870) );
  NAND2X0 U14615 ( .IN1(n13872), .IN2(n13873), .QN(g21029) );
  INVX0 U14616 ( .INP(n13874), .ZN(n13873) );
  NOR2X0 U14617 ( .IN1(n13408), .IN2(n7575), .QN(n13874) );
  NAND2X0 U14618 ( .IN1(n13408), .IN2(n13821), .QN(n13872) );
  INVX0 U14619 ( .INP(n8876), .ZN(n13821) );
  NAND3X0 U14620 ( .IN1(n13875), .IN2(n13876), .IN3(n13877), .QN(n8876) );
  NAND2X0 U14621 ( .IN1(test_so90), .IN2(g7390), .QN(n13877) );
  NAND2X0 U14622 ( .IN1(g7302), .IN2(g2679), .QN(n13876) );
  NAND2X0 U14623 ( .IN1(g2624), .IN2(g2685), .QN(n13875) );
  NAND2X0 U14624 ( .IN1(n13878), .IN2(n13879), .QN(g21028) );
  NAND2X0 U14625 ( .IN1(n9306), .IN2(g2804), .QN(n13879) );
  NAND2X0 U14626 ( .IN1(n11309), .IN2(n8912), .QN(n13878) );
  NAND2X0 U14627 ( .IN1(n13880), .IN2(n13881), .QN(g21027) );
  NAND2X0 U14628 ( .IN1(n12620), .IN2(n4407), .QN(n13881) );
  NAND2X0 U14629 ( .IN1(n12619), .IN2(g2788), .QN(n13880) );
  NAND2X0 U14630 ( .IN1(n13882), .IN2(n13883), .QN(g21026) );
  NAND2X0 U14631 ( .IN1(n4397), .IN2(n12611), .QN(n13883) );
  NAND2X0 U14632 ( .IN1(n12610), .IN2(g2786), .QN(n13882) );
  NAND2X0 U14633 ( .IN1(n13884), .IN2(n13885), .QN(g21025) );
  NAND2X0 U14634 ( .IN1(test_so93), .IN2(n12605), .QN(n13885) );
  NAND2X0 U14635 ( .IN1(n12607), .IN2(n4408), .QN(n13884) );
  NAND2X0 U14636 ( .IN1(n13886), .IN2(n13887), .QN(g21023) );
  NAND2X0 U14637 ( .IN1(n9329), .IN2(g2113), .QN(n13887) );
  NAND2X0 U14638 ( .IN1(n9323), .IN2(n13854), .QN(n13886) );
  NAND2X0 U14639 ( .IN1(n13888), .IN2(n13889), .QN(g21022) );
  NAND2X0 U14640 ( .IN1(n13853), .IN2(g2108), .QN(n13889) );
  INVX0 U14641 ( .INP(n13406), .ZN(n13853) );
  NAND2X0 U14642 ( .IN1(n13406), .IN2(n9001), .QN(n13888) );
  NOR2X0 U14643 ( .IN1(n4293), .IN2(n7758), .QN(n13406) );
  NAND2X0 U14644 ( .IN1(n13890), .IN2(n13891), .QN(g21021) );
  NAND2X0 U14645 ( .IN1(n4468), .IN2(n12685), .QN(n13891) );
  NAND2X0 U14646 ( .IN1(n12684), .IN2(g2097), .QN(n13890) );
  NAND2X0 U14647 ( .IN1(n13892), .IN2(n13893), .QN(g21020) );
  NAND2X0 U14648 ( .IN1(n12676), .IN2(n4409), .QN(n13893) );
  NAND2X0 U14649 ( .IN1(n9335), .IN2(g2095), .QN(n13892) );
  NAND2X0 U14650 ( .IN1(n13894), .IN2(n13895), .QN(g21019) );
  NAND2X0 U14651 ( .IN1(n4399), .IN2(n12616), .QN(n13895) );
  NAND2X0 U14652 ( .IN1(n12614), .IN2(g2090), .QN(n13894) );
  NAND2X0 U14653 ( .IN1(n13896), .IN2(n13897), .QN(g21018) );
  NAND2X0 U14654 ( .IN1(n13898), .IN2(g1417), .QN(n13897) );
  NAND2X0 U14655 ( .IN1(n13411), .IN2(n13899), .QN(n13896) );
  NAND2X0 U14656 ( .IN1(n13900), .IN2(n13901), .QN(g21017) );
  NAND2X0 U14657 ( .IN1(n12753), .IN2(n4475), .QN(n13901) );
  NAND2X0 U14658 ( .IN1(n12752), .IN2(g1406), .QN(n13900) );
  NAND2X0 U14659 ( .IN1(n13902), .IN2(n13903), .QN(g21016) );
  NAND2X0 U14660 ( .IN1(n4469), .IN2(n12741), .QN(n13903) );
  NAND2X0 U14661 ( .IN1(n8530), .IN2(g1404), .QN(n13902) );
  NAND2X0 U14662 ( .IN1(n13904), .IN2(n13905), .QN(g21015) );
  NAND2X0 U14663 ( .IN1(n12680), .IN2(n4411), .QN(n13905) );
  INVX0 U14664 ( .INP(n13906), .ZN(n13904) );
  NOR2X0 U14665 ( .IN1(n12680), .IN2(n7861), .QN(n13906) );
  NAND2X0 U14666 ( .IN1(n13907), .IN2(n13908), .QN(g21011) );
  NAND2X0 U14667 ( .IN1(n4396), .IN2(n12813), .QN(n13908) );
  NAND2X0 U14668 ( .IN1(n12812), .IN2(g723), .QN(n13907) );
  NAND2X0 U14669 ( .IN1(n13909), .IN2(n13910), .QN(g21010) );
  NAND2X0 U14670 ( .IN1(n12809), .IN2(n4477), .QN(n13910) );
  NAND2X0 U14671 ( .IN1(n8551), .IN2(g721), .QN(n13909) );
  NAND2X0 U14672 ( .IN1(n13911), .IN2(n13912), .QN(g21009) );
  NAND2X0 U14673 ( .IN1(n12746), .IN2(n8105), .QN(n13912) );
  NAND2X0 U14674 ( .IN1(n12744), .IN2(g716), .QN(n13911) );
  NAND2X0 U14675 ( .IN1(n13913), .IN2(n13914), .QN(g21007) );
  INVX0 U14676 ( .INP(n13915), .ZN(n13914) );
  NOR2X0 U14677 ( .IN1(n13408), .IN2(n8042), .QN(n13915) );
  NAND2X0 U14678 ( .IN1(n13408), .IN2(n8912), .QN(n13913) );
  INVX0 U14679 ( .INP(n8887), .ZN(n8912) );
  NAND3X0 U14680 ( .IN1(n13916), .IN2(n13917), .IN3(n13918), .QN(n8887) );
  NAND2X0 U14681 ( .IN1(g7390), .IN2(g2691), .QN(n13918) );
  NAND2X0 U14682 ( .IN1(g2624), .IN2(g2694), .QN(n13917) );
  NAND2X0 U14683 ( .IN1(n10186), .IN2(g2688), .QN(n13916) );
  INVX0 U14684 ( .INP(n4314), .ZN(n10186) );
  NOR2X0 U14685 ( .IN1(n4306), .IN2(n7757), .QN(n13408) );
  NAND2X0 U14686 ( .IN1(n13919), .IN2(n13920), .QN(g21006) );
  NAND2X0 U14687 ( .IN1(n4397), .IN2(n12620), .QN(n13920) );
  NAND2X0 U14688 ( .IN1(n12619), .IN2(g2785), .QN(n13919) );
  NAND2X0 U14689 ( .IN1(n13921), .IN2(n13922), .QN(g21005) );
  NAND2X0 U14690 ( .IN1(n12611), .IN2(n4408), .QN(n13922) );
  NAND2X0 U14691 ( .IN1(n12610), .IN2(g2783), .QN(n13921) );
  NAND2X0 U14692 ( .IN1(n13923), .IN2(n13924), .QN(g21004) );
  NAND2X0 U14693 ( .IN1(n4419), .IN2(n12607), .QN(n13924) );
  NAND2X0 U14694 ( .IN1(n12605), .IN2(g2778), .QN(n13923) );
  NAND2X0 U14695 ( .IN1(n13925), .IN2(n13926), .QN(g21003) );
  INVX0 U14696 ( .INP(n13927), .ZN(n13926) );
  NOR2X0 U14697 ( .IN1(n13413), .IN2(n7576), .QN(n13927) );
  NAND2X0 U14698 ( .IN1(n13413), .IN2(n13854), .QN(n13925) );
  INVX0 U14699 ( .INP(n8989), .ZN(n13854) );
  NAND3X0 U14700 ( .IN1(n13928), .IN2(n13929), .IN3(n13930), .QN(n8989) );
  NAND2X0 U14701 ( .IN1(g1930), .IN2(g1991), .QN(n13930) );
  NAND2X0 U14702 ( .IN1(g7052), .IN2(g1985), .QN(n13929) );
  NAND2X0 U14703 ( .IN1(g7194), .IN2(g1988), .QN(n13928) );
  NAND2X0 U14704 ( .IN1(n13931), .IN2(n13932), .QN(g21002) );
  NAND2X0 U14705 ( .IN1(n9329), .IN2(g2110), .QN(n13932) );
  INVX0 U14706 ( .INP(n9323), .ZN(n9329) );
  NAND2X0 U14707 ( .IN1(n9323), .IN2(n9001), .QN(n13931) );
  NAND2X0 U14708 ( .IN1(n13933), .IN2(n13934), .QN(g21001) );
  NAND2X0 U14709 ( .IN1(n12685), .IN2(n4409), .QN(n13934) );
  NAND2X0 U14710 ( .IN1(n12684), .IN2(g2094), .QN(n13933) );
  NAND2X0 U14711 ( .IN1(n13935), .IN2(n13936), .QN(g21000) );
  NAND2X0 U14712 ( .IN1(test_so71), .IN2(n9335), .QN(n13936) );
  NAND2X0 U14713 ( .IN1(n4399), .IN2(n12676), .QN(n13935) );
  NAND2X0 U14714 ( .IN1(n13937), .IN2(n13938), .QN(g20999) );
  NAND2X0 U14715 ( .IN1(n12616), .IN2(n4410), .QN(n13938) );
  NAND2X0 U14716 ( .IN1(n12614), .IN2(g2087), .QN(n13937) );
  NAND2X0 U14717 ( .IN1(n13939), .IN2(n13940), .QN(g20997) );
  NAND2X0 U14718 ( .IN1(n8519), .IN2(g1419), .QN(n13940) );
  NAND2X0 U14719 ( .IN1(n8524), .IN2(n13899), .QN(n13939) );
  NAND2X0 U14720 ( .IN1(n13941), .IN2(n13942), .QN(g20996) );
  NAND2X0 U14721 ( .IN1(test_so51), .IN2(n13898), .QN(n13942) );
  INVX0 U14722 ( .INP(n13411), .ZN(n13898) );
  NAND2X0 U14723 ( .IN1(n13411), .IN2(n9129), .QN(n13941) );
  NOR2X0 U14724 ( .IN1(n4294), .IN2(n7759), .QN(n13411) );
  NAND2X0 U14725 ( .IN1(n13943), .IN2(n13944), .QN(g20995) );
  NAND2X0 U14726 ( .IN1(n4469), .IN2(n12753), .QN(n13944) );
  NAND2X0 U14727 ( .IN1(n12752), .IN2(g1403), .QN(n13943) );
  NAND2X0 U14728 ( .IN1(n13945), .IN2(n13946), .QN(g20994) );
  NAND2X0 U14729 ( .IN1(test_so50), .IN2(n8530), .QN(n13946) );
  NAND2X0 U14730 ( .IN1(n12741), .IN2(n4411), .QN(n13945) );
  NAND2X0 U14731 ( .IN1(n13947), .IN2(n13948), .QN(g20993) );
  NAND2X0 U14732 ( .IN1(n4401), .IN2(n12680), .QN(n13948) );
  INVX0 U14733 ( .INP(n13949), .ZN(n13947) );
  NOR2X0 U14734 ( .IN1(n12680), .IN2(n7862), .QN(n13949) );
  NAND2X0 U14735 ( .IN1(n13950), .IN2(n13951), .QN(g20992) );
  NAND2X0 U14736 ( .IN1(n13952), .IN2(g731), .QN(n13951) );
  NAND2X0 U14737 ( .IN1(n13416), .IN2(n13953), .QN(n13950) );
  NAND2X0 U14738 ( .IN1(n13954), .IN2(n13955), .QN(g20991) );
  NAND2X0 U14739 ( .IN1(n12813), .IN2(n4477), .QN(n13955) );
  NAND2X0 U14740 ( .IN1(n12812), .IN2(g720), .QN(n13954) );
  NAND2X0 U14741 ( .IN1(n13956), .IN2(n13957), .QN(g20990) );
  NAND2X0 U14742 ( .IN1(n12809), .IN2(n8105), .QN(n13957) );
  NAND2X0 U14743 ( .IN1(n8551), .IN2(g718), .QN(n13956) );
  NAND2X0 U14744 ( .IN1(n13958), .IN2(n13959), .QN(g20989) );
  NAND2X0 U14745 ( .IN1(n12746), .IN2(n4413), .QN(n13959) );
  NAND2X0 U14746 ( .IN1(n12744), .IN2(g713), .QN(n13958) );
  NAND2X0 U14747 ( .IN1(n13960), .IN2(n13961), .QN(g20983) );
  NAND2X0 U14748 ( .IN1(n12620), .IN2(n4408), .QN(n13961) );
  NAND2X0 U14749 ( .IN1(n12619), .IN2(g2782), .QN(n13960) );
  NAND2X0 U14750 ( .IN1(n13962), .IN2(n13963), .QN(g20982) );
  NAND2X0 U14751 ( .IN1(n4419), .IN2(n12611), .QN(n13963) );
  NAND2X0 U14752 ( .IN1(n12610), .IN2(g2780), .QN(n13962) );
  NAND2X0 U14753 ( .IN1(n13964), .IN2(n13965), .QN(g20981) );
  NAND2X0 U14754 ( .IN1(n12607), .IN2(n4472), .QN(n13965) );
  NAND2X0 U14755 ( .IN1(n12605), .IN2(g2775), .QN(n13964) );
  NAND2X0 U14756 ( .IN1(n13966), .IN2(n13967), .QN(g20980) );
  INVX0 U14757 ( .INP(n13968), .ZN(n13967) );
  NOR2X0 U14758 ( .IN1(n13413), .IN2(n8041), .QN(n13968) );
  NAND2X0 U14759 ( .IN1(n13413), .IN2(n9001), .QN(n13966) );
  INVX0 U14760 ( .INP(n9011), .ZN(n9001) );
  NAND3X0 U14761 ( .IN1(n13969), .IN2(n13970), .IN3(n13971), .QN(n9011) );
  NAND2X0 U14762 ( .IN1(g1930), .IN2(g2000), .QN(n13971) );
  NAND2X0 U14763 ( .IN1(n10234), .IN2(g1994), .QN(n13970) );
  INVX0 U14764 ( .INP(n4296), .ZN(n10234) );
  NAND2X0 U14765 ( .IN1(g7194), .IN2(g1997), .QN(n13969) );
  NOR2X0 U14766 ( .IN1(n4307), .IN2(n7758), .QN(n13413) );
  NAND2X0 U14767 ( .IN1(n13972), .IN2(n13973), .QN(g20979) );
  NAND2X0 U14768 ( .IN1(n4399), .IN2(n12685), .QN(n13973) );
  NAND2X0 U14769 ( .IN1(n12684), .IN2(g2091), .QN(n13972) );
  NAND2X0 U14770 ( .IN1(n13974), .IN2(n13975), .QN(g20978) );
  NAND2X0 U14771 ( .IN1(n12676), .IN2(n4410), .QN(n13975) );
  NAND2X0 U14772 ( .IN1(n9335), .IN2(g2089), .QN(n13974) );
  NAND2X0 U14773 ( .IN1(n13976), .IN2(n13977), .QN(g20977) );
  NAND2X0 U14774 ( .IN1(n4420), .IN2(n12616), .QN(n13977) );
  NAND2X0 U14775 ( .IN1(n12614), .IN2(g2084), .QN(n13976) );
  NAND2X0 U14776 ( .IN1(n13978), .IN2(n13979), .QN(g20976) );
  INVX0 U14777 ( .INP(n13980), .ZN(n13979) );
  NOR2X0 U14778 ( .IN1(n13418), .IN2(n7577), .QN(n13980) );
  NAND2X0 U14779 ( .IN1(n13418), .IN2(n13899), .QN(n13978) );
  INVX0 U14780 ( .INP(n9106), .ZN(n13899) );
  NAND3X0 U14781 ( .IN1(n13981), .IN2(n13982), .IN3(n13983), .QN(n9106) );
  NAND2X0 U14782 ( .IN1(g6944), .IN2(g1294), .QN(n13983) );
  NAND2X0 U14783 ( .IN1(g6750), .IN2(g1291), .QN(n13982) );
  NAND2X0 U14784 ( .IN1(g1236), .IN2(g1297), .QN(n13981) );
  NAND2X0 U14785 ( .IN1(n13984), .IN2(n13985), .QN(g20975) );
  NAND2X0 U14786 ( .IN1(n8519), .IN2(g1416), .QN(n13985) );
  INVX0 U14787 ( .INP(n8524), .ZN(n8519) );
  NAND2X0 U14788 ( .IN1(n8524), .IN2(n9129), .QN(n13984) );
  NAND2X0 U14789 ( .IN1(n13986), .IN2(n13987), .QN(g20974) );
  NAND2X0 U14790 ( .IN1(n12753), .IN2(n4411), .QN(n13987) );
  NAND2X0 U14791 ( .IN1(n12752), .IN2(g1400), .QN(n13986) );
  NAND2X0 U14792 ( .IN1(n13988), .IN2(n13989), .QN(g20973) );
  NAND2X0 U14793 ( .IN1(n4401), .IN2(n12741), .QN(n13989) );
  NAND2X0 U14794 ( .IN1(n8530), .IN2(g1398), .QN(n13988) );
  NAND2X0 U14795 ( .IN1(n13990), .IN2(n13991), .QN(g20972) );
  NAND2X0 U14796 ( .IN1(n12680), .IN2(n4412), .QN(n13991) );
  INVX0 U14797 ( .INP(n13992), .ZN(n13990) );
  NOR2X0 U14798 ( .IN1(n12680), .IN2(n7863), .QN(n13992) );
  NAND2X0 U14799 ( .IN1(n13993), .IN2(n13994), .QN(g20970) );
  NAND2X0 U14800 ( .IN1(n8539), .IN2(g733), .QN(n13994) );
  NAND2X0 U14801 ( .IN1(n8548), .IN2(n13953), .QN(n13993) );
  NAND2X0 U14802 ( .IN1(n13995), .IN2(n13996), .QN(g20969) );
  NAND2X0 U14803 ( .IN1(n13952), .IN2(g728), .QN(n13996) );
  INVX0 U14804 ( .INP(n13416), .ZN(n13952) );
  NAND2X0 U14805 ( .IN1(n13416), .IN2(n13997), .QN(n13995) );
  NOR2X0 U14806 ( .IN1(n4295), .IN2(n7760), .QN(n13416) );
  NAND2X0 U14807 ( .IN1(n13998), .IN2(n13999), .QN(g20968) );
  NAND2X0 U14808 ( .IN1(n12813), .IN2(n8105), .QN(n13999) );
  NAND2X0 U14809 ( .IN1(n12812), .IN2(g717), .QN(n13998) );
  NAND2X0 U14810 ( .IN1(n14000), .IN2(n14001), .QN(g20967) );
  NAND2X0 U14811 ( .IN1(n12809), .IN2(n4413), .QN(n14001) );
  NAND2X0 U14812 ( .IN1(n8551), .IN2(g715), .QN(n14000) );
  NAND2X0 U14813 ( .IN1(n14002), .IN2(n14003), .QN(g20966) );
  NAND2X0 U14814 ( .IN1(n4403), .IN2(n12746), .QN(n14003) );
  NAND2X0 U14815 ( .IN1(n12744), .IN2(g710), .QN(n14002) );
  NAND2X0 U14816 ( .IN1(n14004), .IN2(n14005), .QN(g20965) );
  NAND2X0 U14817 ( .IN1(n4415), .IN2(n12607), .QN(n14005) );
  NAND2X0 U14818 ( .IN1(n12605), .IN2(g2799), .QN(n14004) );
  NAND2X0 U14819 ( .IN1(n14006), .IN2(n14007), .QN(g20964) );
  NAND2X0 U14820 ( .IN1(n4419), .IN2(n12620), .QN(n14007) );
  NAND2X0 U14821 ( .IN1(n12619), .IN2(g2779), .QN(n14006) );
  NAND2X0 U14822 ( .IN1(n14008), .IN2(n14009), .QN(g20963) );
  NAND2X0 U14823 ( .IN1(n12611), .IN2(n4472), .QN(n14009) );
  NAND2X0 U14824 ( .IN1(n12610), .IN2(g2777), .QN(n14008) );
  NAND2X0 U14825 ( .IN1(n14010), .IN2(n14011), .QN(g20962) );
  NAND2X0 U14826 ( .IN1(n4398), .IN2(n12607), .QN(n14011) );
  INVX0 U14827 ( .INP(n12605), .ZN(n12607) );
  NAND2X0 U14828 ( .IN1(n12605), .IN2(g2772), .QN(n14010) );
  NAND2X0 U14829 ( .IN1(n14012), .IN2(n9314), .QN(n12605) );
  NAND2X0 U14830 ( .IN1(n14013), .IN2(n14014), .QN(g20955) );
  NAND2X0 U14831 ( .IN1(n12685), .IN2(n4410), .QN(n14014) );
  NAND2X0 U14832 ( .IN1(n12684), .IN2(g2088), .QN(n14013) );
  NAND2X0 U14833 ( .IN1(n14015), .IN2(n14016), .QN(g20954) );
  NAND2X0 U14834 ( .IN1(n4420), .IN2(n12676), .QN(n14016) );
  NAND2X0 U14835 ( .IN1(n9335), .IN2(g2086), .QN(n14015) );
  NAND2X0 U14836 ( .IN1(n14017), .IN2(n14018), .QN(g20953) );
  NAND2X0 U14837 ( .IN1(n12616), .IN2(n4474), .QN(n14018) );
  NAND2X0 U14838 ( .IN1(n12614), .IN2(g2081), .QN(n14017) );
  NAND2X0 U14839 ( .IN1(n14019), .IN2(n14020), .QN(g20952) );
  INVX0 U14840 ( .INP(n14021), .ZN(n14020) );
  NOR2X0 U14841 ( .IN1(n13418), .IN2(n8039), .QN(n14021) );
  NAND2X0 U14842 ( .IN1(n13418), .IN2(n9129), .QN(n14019) );
  INVX0 U14843 ( .INP(n9117), .ZN(n9129) );
  NAND3X0 U14844 ( .IN1(n14022), .IN2(n14023), .IN3(n14024), .QN(n9117) );
  NAND2X0 U14845 ( .IN1(n11110), .IN2(g1300), .QN(n14024) );
  INVX0 U14846 ( .INP(n4371), .ZN(n11110) );
  NAND2X0 U14847 ( .IN1(g1236), .IN2(g1306), .QN(n14023) );
  NAND2X0 U14848 ( .IN1(g6944), .IN2(g1303), .QN(n14022) );
  NOR2X0 U14849 ( .IN1(n4308), .IN2(n7759), .QN(n13418) );
  NAND2X0 U14850 ( .IN1(n14025), .IN2(n14026), .QN(g20951) );
  NAND2X0 U14851 ( .IN1(n4401), .IN2(n12753), .QN(n14026) );
  NAND2X0 U14852 ( .IN1(n12752), .IN2(g1397), .QN(n14025) );
  NAND2X0 U14853 ( .IN1(n14027), .IN2(n14028), .QN(g20950) );
  NAND2X0 U14854 ( .IN1(n12741), .IN2(n4412), .QN(n14028) );
  NAND2X0 U14855 ( .IN1(n8530), .IN2(g1395), .QN(n14027) );
  NAND2X0 U14856 ( .IN1(n14029), .IN2(n14030), .QN(g20949) );
  NAND2X0 U14857 ( .IN1(n4421), .IN2(n12680), .QN(n14030) );
  INVX0 U14858 ( .INP(n14031), .ZN(n14029) );
  NOR2X0 U14859 ( .IN1(n12680), .IN2(n7864), .QN(n14031) );
  NAND2X0 U14860 ( .IN1(n14032), .IN2(n14033), .QN(g20948) );
  INVX0 U14861 ( .INP(n14034), .ZN(n14033) );
  NOR2X0 U14862 ( .IN1(n13421), .IN2(n7578), .QN(n14034) );
  NAND2X0 U14863 ( .IN1(n13421), .IN2(n13953), .QN(n14032) );
  INVX0 U14864 ( .INP(n8758), .ZN(n13953) );
  NAND3X0 U14865 ( .IN1(n14035), .IN2(n14036), .IN3(n14037), .QN(n8758) );
  NAND2X0 U14866 ( .IN1(g6642), .IN2(g608), .QN(n14037) );
  NAND2X0 U14867 ( .IN1(n11213), .IN2(g605), .QN(n14036) );
  INVX0 U14868 ( .INP(n4298), .ZN(n11213) );
  NAND2X0 U14869 ( .IN1(g550), .IN2(g611), .QN(n14035) );
  NAND2X0 U14870 ( .IN1(n14038), .IN2(n14039), .QN(g20947) );
  NAND2X0 U14871 ( .IN1(n8539), .IN2(g730), .QN(n14039) );
  INVX0 U14872 ( .INP(n8548), .ZN(n8539) );
  NAND2X0 U14873 ( .IN1(n8548), .IN2(n13997), .QN(n14038) );
  NAND2X0 U14874 ( .IN1(n14040), .IN2(n14041), .QN(g20946) );
  NAND2X0 U14875 ( .IN1(n12813), .IN2(n4413), .QN(n14041) );
  NAND2X0 U14876 ( .IN1(n12812), .IN2(g714), .QN(n14040) );
  NAND2X0 U14877 ( .IN1(n14042), .IN2(n14043), .QN(g20945) );
  NAND2X0 U14878 ( .IN1(n4403), .IN2(n12809), .QN(n14043) );
  NAND2X0 U14879 ( .IN1(n8551), .IN2(g712), .QN(n14042) );
  NAND2X0 U14880 ( .IN1(n14044), .IN2(n14045), .QN(g20944) );
  NAND2X0 U14881 ( .IN1(n12746), .IN2(n4414), .QN(n14045) );
  NAND2X0 U14882 ( .IN1(n12744), .IN2(g707), .QN(n14044) );
  NAND2X0 U14883 ( .IN1(n14046), .IN2(n14047), .QN(g20941) );
  NAND2X0 U14884 ( .IN1(n4415), .IN2(n12611), .QN(n14047) );
  NAND2X0 U14885 ( .IN1(n12610), .IN2(g2801), .QN(n14046) );
  NAND2X0 U14886 ( .IN1(n14048), .IN2(n14049), .QN(g20940) );
  NAND2X0 U14887 ( .IN1(n12620), .IN2(n4472), .QN(n14049) );
  NAND2X0 U14888 ( .IN1(n12619), .IN2(g2776), .QN(n14048) );
  NAND2X0 U14889 ( .IN1(n14050), .IN2(n14051), .QN(g20939) );
  NAND2X0 U14890 ( .IN1(n4398), .IN2(n12611), .QN(n14051) );
  INVX0 U14891 ( .INP(n12610), .ZN(n12611) );
  NAND2X0 U14892 ( .IN1(n12610), .IN2(g2774), .QN(n14050) );
  NAND3X0 U14893 ( .IN1(n4426), .IN2(g7487), .IN3(n14012), .QN(n12610) );
  NAND2X0 U14894 ( .IN1(n14052), .IN2(n14053), .QN(g20937) );
  NAND2X0 U14895 ( .IN1(n4416), .IN2(n12616), .QN(n14053) );
  NAND2X0 U14896 ( .IN1(n12614), .IN2(g2105), .QN(n14052) );
  NAND2X0 U14897 ( .IN1(n14054), .IN2(n14055), .QN(g20936) );
  NAND2X0 U14898 ( .IN1(n4420), .IN2(n12685), .QN(n14055) );
  NAND2X0 U14899 ( .IN1(n12684), .IN2(g2085), .QN(n14054) );
  NAND2X0 U14900 ( .IN1(n14056), .IN2(n14057), .QN(g20935) );
  NAND2X0 U14901 ( .IN1(n12676), .IN2(n4474), .QN(n14057) );
  NAND2X0 U14902 ( .IN1(n9335), .IN2(g2083), .QN(n14056) );
  NAND2X0 U14903 ( .IN1(n14058), .IN2(n14059), .QN(g20934) );
  NAND2X0 U14904 ( .IN1(n4400), .IN2(n12616), .QN(n14059) );
  INVX0 U14905 ( .INP(n12614), .ZN(n12616) );
  NAND2X0 U14906 ( .IN1(n12614), .IN2(g2078), .QN(n14058) );
  NAND2X0 U14907 ( .IN1(n14060), .IN2(n9332), .QN(n12614) );
  NAND2X0 U14908 ( .IN1(n14061), .IN2(n14062), .QN(g20927) );
  NAND2X0 U14909 ( .IN1(n12753), .IN2(n4412), .QN(n14062) );
  NAND2X0 U14910 ( .IN1(n12752), .IN2(g1394), .QN(n14061) );
  NAND2X0 U14911 ( .IN1(n14063), .IN2(n14064), .QN(g20926) );
  NAND2X0 U14912 ( .IN1(n4421), .IN2(n12741), .QN(n14064) );
  NAND2X0 U14913 ( .IN1(n8530), .IN2(g1392), .QN(n14063) );
  NAND2X0 U14914 ( .IN1(n14065), .IN2(n14066), .QN(g20925) );
  NAND2X0 U14915 ( .IN1(n12680), .IN2(n4476), .QN(n14066) );
  INVX0 U14916 ( .INP(n14067), .ZN(n14065) );
  NOR2X0 U14917 ( .IN1(n12680), .IN2(n7865), .QN(n14067) );
  NAND2X0 U14918 ( .IN1(n14068), .IN2(n14069), .QN(g20924) );
  INVX0 U14919 ( .INP(n14070), .ZN(n14069) );
  NOR2X0 U14920 ( .IN1(n13421), .IN2(n8038), .QN(n14070) );
  NAND2X0 U14921 ( .IN1(n13421), .IN2(n13997), .QN(n14068) );
  INVX0 U14922 ( .INP(n8764), .ZN(n13997) );
  NAND3X0 U14923 ( .IN1(n14071), .IN2(n14072), .IN3(n14073), .QN(n8764) );
  NAND2X0 U14924 ( .IN1(g6642), .IN2(g617), .QN(n14073) );
  NAND2X0 U14925 ( .IN1(g6485), .IN2(g614), .QN(n14072) );
  NAND2X0 U14926 ( .IN1(test_so26), .IN2(g550), .QN(n14071) );
  NOR2X0 U14927 ( .IN1(n4309), .IN2(n7760), .QN(n13421) );
  NAND2X0 U14928 ( .IN1(n14074), .IN2(n14075), .QN(g20923) );
  NAND2X0 U14929 ( .IN1(test_so29), .IN2(n12812), .QN(n14075) );
  NAND2X0 U14930 ( .IN1(n4403), .IN2(n12813), .QN(n14074) );
  NAND2X0 U14931 ( .IN1(n14076), .IN2(n14077), .QN(g20922) );
  NAND2X0 U14932 ( .IN1(n12809), .IN2(n4414), .QN(n14077) );
  NAND2X0 U14933 ( .IN1(n8551), .IN2(g709), .QN(n14076) );
  NAND2X0 U14934 ( .IN1(n14078), .IN2(n14079), .QN(g20921) );
  NAND2X0 U14935 ( .IN1(n4422), .IN2(n12746), .QN(n14079) );
  NAND2X0 U14936 ( .IN1(n12744), .IN2(g704), .QN(n14078) );
  NAND2X0 U14937 ( .IN1(n14080), .IN2(n14081), .QN(g20919) );
  NAND2X0 U14938 ( .IN1(n4415), .IN2(n12620), .QN(n14081) );
  NAND2X0 U14939 ( .IN1(n12619), .IN2(g2800), .QN(n14080) );
  NAND2X0 U14940 ( .IN1(n14082), .IN2(n14083), .QN(g20918) );
  NAND2X0 U14941 ( .IN1(n4398), .IN2(n12620), .QN(n14083) );
  INVX0 U14942 ( .INP(n12619), .ZN(n12620) );
  NAND2X0 U14943 ( .IN1(n12619), .IN2(g2773), .QN(n14082) );
  NAND3X0 U14944 ( .IN1(n4426), .IN2(g7425), .IN3(n14012), .QN(n12619) );
  NOR2X0 U14945 ( .IN1(n4490), .IN2(n8067), .QN(n14012) );
  NAND2X0 U14946 ( .IN1(n14084), .IN2(n14085), .QN(g20917) );
  NAND2X0 U14947 ( .IN1(test_so72), .IN2(n9335), .QN(n14085) );
  NAND2X0 U14948 ( .IN1(n4416), .IN2(n12676), .QN(n14084) );
  NAND2X0 U14949 ( .IN1(n14086), .IN2(n14087), .QN(g20916) );
  NAND2X0 U14950 ( .IN1(n12685), .IN2(n4474), .QN(n14087) );
  NAND2X0 U14951 ( .IN1(n12684), .IN2(g2082), .QN(n14086) );
  NAND2X0 U14952 ( .IN1(n14088), .IN2(n14089), .QN(g20915) );
  NAND2X0 U14953 ( .IN1(n4400), .IN2(n12676), .QN(n14089) );
  INVX0 U14954 ( .INP(n9335), .ZN(n12676) );
  NAND2X0 U14955 ( .IN1(n9335), .IN2(g2080), .QN(n14088) );
  NAND3X0 U14956 ( .IN1(n4427), .IN2(g7357), .IN3(n14060), .QN(n9335) );
  NAND2X0 U14957 ( .IN1(n14090), .IN2(n14091), .QN(g20913) );
  NAND2X0 U14958 ( .IN1(n4417), .IN2(n12680), .QN(n14091) );
  INVX0 U14959 ( .INP(n14092), .ZN(n14090) );
  NOR2X0 U14960 ( .IN1(n12680), .IN2(n7857), .QN(n14092) );
  NAND2X0 U14961 ( .IN1(n14093), .IN2(n14094), .QN(g20912) );
  NAND2X0 U14962 ( .IN1(n4421), .IN2(n12753), .QN(n14094) );
  NAND2X0 U14963 ( .IN1(n12752), .IN2(g1391), .QN(n14093) );
  NAND2X0 U14964 ( .IN1(n14095), .IN2(n14096), .QN(g20911) );
  NAND2X0 U14965 ( .IN1(n12741), .IN2(n4476), .QN(n14096) );
  NAND2X0 U14966 ( .IN1(n8530), .IN2(g1389), .QN(n14095) );
  NAND2X0 U14967 ( .IN1(n14097), .IN2(n14098), .QN(g20910) );
  NAND2X0 U14968 ( .IN1(n4402), .IN2(n12680), .QN(n14098) );
  INVX0 U14969 ( .INP(n14099), .ZN(n14097) );
  NOR2X0 U14970 ( .IN1(n12680), .IN2(n7866), .QN(n14099) );
  NOR2X0 U14971 ( .IN1(n14100), .IN2(n8527), .QN(n12680) );
  INVX0 U14972 ( .INP(n14101), .ZN(n14100) );
  NAND2X0 U14973 ( .IN1(n14102), .IN2(n14103), .QN(g20903) );
  NAND2X0 U14974 ( .IN1(n12813), .IN2(n4414), .QN(n14103) );
  NAND2X0 U14975 ( .IN1(n12812), .IN2(g708), .QN(n14102) );
  NAND2X0 U14976 ( .IN1(n14104), .IN2(n14105), .QN(g20902) );
  NAND2X0 U14977 ( .IN1(n4422), .IN2(n12809), .QN(n14105) );
  NAND2X0 U14978 ( .IN1(n8551), .IN2(g706), .QN(n14104) );
  NAND2X0 U14979 ( .IN1(n14106), .IN2(n14107), .QN(g20901) );
  NAND2X0 U14980 ( .IN1(n12746), .IN2(n4478), .QN(n14107) );
  NAND2X0 U14981 ( .IN1(n12744), .IN2(g701), .QN(n14106) );
  NAND2X0 U14982 ( .IN1(n14108), .IN2(n14109), .QN(g20900) );
  NAND2X0 U14983 ( .IN1(n4416), .IN2(n12685), .QN(n14109) );
  NAND2X0 U14984 ( .IN1(n12684), .IN2(g2106), .QN(n14108) );
  NAND2X0 U14985 ( .IN1(n14110), .IN2(n14111), .QN(g20899) );
  NAND2X0 U14986 ( .IN1(n4400), .IN2(n12685), .QN(n14111) );
  INVX0 U14987 ( .INP(n12684), .ZN(n12685) );
  NAND2X0 U14988 ( .IN1(n12684), .IN2(g2079), .QN(n14110) );
  NAND3X0 U14989 ( .IN1(n4427), .IN2(g7229), .IN3(n14060), .QN(n12684) );
  NOR2X0 U14990 ( .IN1(n8111), .IN2(n8064), .QN(n14060) );
  NAND2X0 U14991 ( .IN1(n14112), .IN2(n14113), .QN(g20898) );
  NAND2X0 U14992 ( .IN1(n4417), .IN2(n12741), .QN(n14113) );
  NAND2X0 U14993 ( .IN1(n8530), .IN2(g1413), .QN(n14112) );
  NAND2X0 U14994 ( .IN1(n14114), .IN2(n14115), .QN(g20897) );
  NAND2X0 U14995 ( .IN1(n12753), .IN2(n4476), .QN(n14115) );
  NAND2X0 U14996 ( .IN1(n12752), .IN2(g1388), .QN(n14114) );
  NAND2X0 U14997 ( .IN1(n14116), .IN2(n14117), .QN(g20896) );
  NAND2X0 U14998 ( .IN1(n4402), .IN2(n12741), .QN(n14117) );
  INVX0 U14999 ( .INP(n8530), .ZN(n12741) );
  NAND2X0 U15000 ( .IN1(n8530), .IN2(g1386), .QN(n14116) );
  NAND3X0 U15001 ( .IN1(n4428), .IN2(g7161), .IN3(n14101), .QN(n8530) );
  NAND2X0 U15002 ( .IN1(n14118), .IN2(n14119), .QN(g20894) );
  NAND2X0 U15003 ( .IN1(n4418), .IN2(n12746), .QN(n14119) );
  NAND2X0 U15004 ( .IN1(n12744), .IN2(g725), .QN(n14118) );
  NAND2X0 U15005 ( .IN1(n14120), .IN2(n14121), .QN(g20893) );
  NAND2X0 U15006 ( .IN1(n4422), .IN2(n12813), .QN(n14121) );
  NAND2X0 U15007 ( .IN1(n12812), .IN2(g705), .QN(n14120) );
  NAND2X0 U15008 ( .IN1(n14122), .IN2(n14123), .QN(g20892) );
  NAND2X0 U15009 ( .IN1(n12809), .IN2(n4478), .QN(n14123) );
  NAND2X0 U15010 ( .IN1(n8551), .IN2(g703), .QN(n14122) );
  NAND2X0 U15011 ( .IN1(n14124), .IN2(n14125), .QN(g20891) );
  NAND2X0 U15012 ( .IN1(n4404), .IN2(n12746), .QN(n14125) );
  INVX0 U15013 ( .INP(n12744), .ZN(n12746) );
  NAND2X0 U15014 ( .IN1(n12744), .IN2(g698), .QN(n14124) );
  NAND2X0 U15015 ( .IN1(n14126), .IN2(n8547), .QN(n12744) );
  NOR2X0 U15016 ( .IN1(g3234), .IN2(DFF_1561_n1), .QN(g20884) );
  NAND2X0 U15017 ( .IN1(n14127), .IN2(n14128), .QN(g20883) );
  NAND2X0 U15018 ( .IN1(n4417), .IN2(n12753), .QN(n14128) );
  NAND2X0 U15019 ( .IN1(n12752), .IN2(g1412), .QN(n14127) );
  NAND2X0 U15020 ( .IN1(n14129), .IN2(n14130), .QN(g20882) );
  NAND2X0 U15021 ( .IN1(test_so49), .IN2(n12752), .QN(n14130) );
  NAND2X0 U15022 ( .IN1(n4402), .IN2(n12753), .QN(n14129) );
  INVX0 U15023 ( .INP(n12752), .ZN(n12753) );
  NAND3X0 U15024 ( .IN1(n4428), .IN2(g6979), .IN3(n14101), .QN(n12752) );
  NOR2X0 U15025 ( .IN1(n4489), .IN2(n8063), .QN(n14101) );
  NAND2X0 U15026 ( .IN1(n14131), .IN2(n14132), .QN(g20881) );
  NAND2X0 U15027 ( .IN1(test_so30), .IN2(n8551), .QN(n14132) );
  NAND2X0 U15028 ( .IN1(n4418), .IN2(n12809), .QN(n14131) );
  NAND2X0 U15029 ( .IN1(n14133), .IN2(n14134), .QN(g20880) );
  NAND2X0 U15030 ( .IN1(n12813), .IN2(n4478), .QN(n14134) );
  NAND2X0 U15031 ( .IN1(n12812), .IN2(g702), .QN(n14133) );
  NAND2X0 U15032 ( .IN1(n14135), .IN2(n14136), .QN(g20879) );
  NAND2X0 U15033 ( .IN1(n4404), .IN2(n12809), .QN(n14136) );
  INVX0 U15034 ( .INP(n8551), .ZN(n12809) );
  NAND2X0 U15035 ( .IN1(n8551), .IN2(g700), .QN(n14135) );
  NAND3X0 U15036 ( .IN1(n4429), .IN2(g6911), .IN3(n14126), .QN(n8551) );
  NAND2X0 U15037 ( .IN1(n14137), .IN2(n14138), .QN(g20876) );
  NAND2X0 U15038 ( .IN1(n4418), .IN2(n12813), .QN(n14138) );
  NAND2X0 U15039 ( .IN1(n12812), .IN2(g726), .QN(n14137) );
  NAND2X0 U15040 ( .IN1(n14139), .IN2(n14140), .QN(g20875) );
  NAND2X0 U15041 ( .IN1(n4404), .IN2(n12813), .QN(n14140) );
  INVX0 U15042 ( .INP(n12812), .ZN(n12813) );
  NAND2X0 U15043 ( .IN1(n12812), .IN2(g699), .QN(n14139) );
  NAND3X0 U15044 ( .IN1(n4429), .IN2(g6677), .IN3(n14126), .QN(n12812) );
  NOR2X0 U15045 ( .IN1(n4492), .IN2(n8054), .QN(n14126) );
  NAND2X0 U15046 ( .IN1(n14141), .IN2(n14142), .QN(g20874) );
  NAND2X0 U15047 ( .IN1(g2879), .IN2(g8096), .QN(n14142) );
  NAND2X0 U15048 ( .IN1(n4351), .IN2(n13784), .QN(n14141) );
  XOR2X1 U15049 ( .IN1(n8562), .IN2(n13787), .Q(n13784) );
  NOR2X0 U15050 ( .IN1(g3231), .IN2(n14385), .QN(n13787) );
  XOR3X1 U15051 ( .IN1(n14143), .IN2(n14144), .IN3(n14145), .Q(n8562) );
  XOR3X1 U15052 ( .IN1(n8010), .IN2(n8002), .IN3(n14146), .Q(n14145) );
  XOR2X1 U15053 ( .IN1(g2944), .IN2(n8012), .Q(n14146) );
  XOR2X1 U15054 ( .IN1(n7999), .IN2(n7998), .Q(n14144) );
  XOR2X1 U15055 ( .IN1(n8001), .IN2(n8000), .Q(n14143) );
  NOR2X0 U15056 ( .IN1(n11309), .IN2(n14147), .QN(g20789) );
  XOR2X1 U15057 ( .IN1(n4398), .IN2(n9314), .Q(n14147) );
  NOR2X0 U15058 ( .IN1(g2733), .IN2(n4292), .QN(n9314) );
  INVX0 U15059 ( .INP(n9306), .ZN(n11309) );
  NAND2X0 U15060 ( .IN1(g7487), .IN2(g2704), .QN(n9306) );
  NOR2X0 U15061 ( .IN1(n9323), .IN2(n14148), .QN(g20752) );
  XOR2X1 U15062 ( .IN1(n4400), .IN2(n9332), .Q(n14148) );
  NOR2X0 U15063 ( .IN1(g2039), .IN2(n4293), .QN(n9332) );
  NOR2X0 U15064 ( .IN1(n4357), .IN2(n7758), .QN(n9323) );
  NOR2X0 U15065 ( .IN1(n8524), .IN2(n14149), .QN(g20717) );
  XNOR2X1 U15066 ( .IN1(n4402), .IN2(n8527), .Q(n14149) );
  NAND2X0 U15067 ( .IN1(n4428), .IN2(g1315), .QN(n8527) );
  NOR2X0 U15068 ( .IN1(n4358), .IN2(n7759), .QN(n8524) );
  NOR2X0 U15069 ( .IN1(n8548), .IN2(n14150), .QN(g20682) );
  XOR2X1 U15070 ( .IN1(n4404), .IN2(n8547), .Q(n14150) );
  NOR2X0 U15071 ( .IN1(g659), .IN2(n4295), .QN(n8547) );
  NOR2X0 U15072 ( .IN1(n4359), .IN2(n7760), .QN(n8548) );
  NAND2X0 U15073 ( .IN1(n14151), .IN2(n14152), .QN(g20417) );
  NAND2X0 U15074 ( .IN1(n4351), .IN2(g2963), .QN(n14152) );
  NAND2X0 U15075 ( .IN1(g2879), .IN2(g7334), .QN(n14151) );
  NAND2X0 U15076 ( .IN1(n14153), .IN2(n14154), .QN(g20376) );
  NAND2X0 U15077 ( .IN1(test_so2), .IN2(n4351), .QN(n14154) );
  NAND2X0 U15078 ( .IN1(g2879), .IN2(g6895), .QN(n14153) );
  NAND2X0 U15079 ( .IN1(n14155), .IN2(n14156), .QN(g20375) );
  NAND2X0 U15080 ( .IN1(n4292), .IN2(g2733), .QN(n14156) );
  NAND2X0 U15081 ( .IN1(n14157), .IN2(g2703), .QN(n14155) );
  NAND2X0 U15082 ( .IN1(n14158), .IN2(n14159), .QN(g20353) );
  NAND2X0 U15083 ( .IN1(n4293), .IN2(g2039), .QN(n14159) );
  NAND2X0 U15084 ( .IN1(n14157), .IN2(g2009), .QN(n14158) );
  NAND2X0 U15085 ( .IN1(n14160), .IN2(n14161), .QN(g20343) );
  NAND2X0 U15086 ( .IN1(n4351), .IN2(g2969), .QN(n14161) );
  NAND2X0 U15087 ( .IN1(g2879), .IN2(g6442), .QN(n14160) );
  NAND2X0 U15088 ( .IN1(n14162), .IN2(n14163), .QN(g20333) );
  NAND2X0 U15089 ( .IN1(n4294), .IN2(g1345), .QN(n14163) );
  NAND2X0 U15090 ( .IN1(n14157), .IN2(g1315), .QN(n14162) );
  NAND2X0 U15091 ( .IN1(n14164), .IN2(n14165), .QN(g20314) );
  NAND2X0 U15092 ( .IN1(n4295), .IN2(g659), .QN(n14165) );
  NAND2X0 U15093 ( .IN1(n14157), .IN2(g629), .QN(n14164) );
  INVX0 U15094 ( .INP(n13377), .ZN(n14157) );
  NAND4X0 U15095 ( .IN1(n8073), .IN2(n8052), .IN3(n14166), .IN4(n8051), .QN(
        n13377) );
  NOR2X0 U15096 ( .IN1(test_so98), .IN2(g3006), .QN(n14166) );
  NAND2X0 U15097 ( .IN1(n14167), .IN2(n14168), .QN(g20310) );
  NAND2X0 U15098 ( .IN1(n4351), .IN2(g2972), .QN(n14168) );
  NAND2X0 U15099 ( .IN1(g2879), .IN2(g6225), .QN(n14167) );
  NAND2X0 U15100 ( .IN1(n14169), .IN2(n14170), .QN(g19184) );
  NAND2X0 U15101 ( .IN1(n4351), .IN2(g2975), .QN(n14170) );
  NAND2X0 U15102 ( .IN1(g2879), .IN2(g4590), .QN(n14169) );
  NAND2X0 U15103 ( .IN1(n14171), .IN2(n14172), .QN(g19178) );
  NAND2X0 U15104 ( .IN1(n4351), .IN2(g2935), .QN(n14172) );
  NAND2X0 U15105 ( .IN1(test_so5), .IN2(g2879), .QN(n14171) );
  NAND2X0 U15106 ( .IN1(n14173), .IN2(n14174), .QN(g19173) );
  NAND2X0 U15107 ( .IN1(n4351), .IN2(g2978), .QN(n14174) );
  NAND2X0 U15108 ( .IN1(g2879), .IN2(g4323), .QN(n14173) );
  NAND2X0 U15109 ( .IN1(n14175), .IN2(n14176), .QN(g19172) );
  NAND2X0 U15110 ( .IN1(n4351), .IN2(g2953), .QN(n14176) );
  NAND2X0 U15111 ( .IN1(g2879), .IN2(g4321), .QN(n14175) );
  NAND2X0 U15112 ( .IN1(n14177), .IN2(n14178), .QN(g19167) );
  NAND2X0 U15113 ( .IN1(n4351), .IN2(g2938), .QN(n14178) );
  NAND2X0 U15114 ( .IN1(g2879), .IN2(g4200), .QN(n14177) );
  NAND2X0 U15115 ( .IN1(n14179), .IN2(n14180), .QN(g19163) );
  NAND2X0 U15116 ( .IN1(n4351), .IN2(g2981), .QN(n14180) );
  NAND2X0 U15117 ( .IN1(g2879), .IN2(g4090), .QN(n14179) );
  NAND2X0 U15118 ( .IN1(n14181), .IN2(n14182), .QN(g19162) );
  NAND2X0 U15119 ( .IN1(n4351), .IN2(g2956), .QN(n14182) );
  NAND2X0 U15120 ( .IN1(g2879), .IN2(g4088), .QN(n14181) );
  NAND2X0 U15121 ( .IN1(n14183), .IN2(n14184), .QN(g19157) );
  NAND2X0 U15122 ( .IN1(n4351), .IN2(g2941), .QN(n14184) );
  NAND2X0 U15123 ( .IN1(g2879), .IN2(g3993), .QN(n14183) );
  NAND2X0 U15124 ( .IN1(n14185), .IN2(n14186), .QN(g19154) );
  NAND2X0 U15125 ( .IN1(n4351), .IN2(g2874), .QN(n14186) );
  NAND2X0 U15126 ( .IN1(test_so3), .IN2(g2879), .QN(n14185) );
  NAND2X0 U15127 ( .IN1(n14187), .IN2(n14188), .QN(g19153) );
  NAND2X0 U15128 ( .IN1(n4351), .IN2(g2959), .QN(n14188) );
  NAND2X0 U15129 ( .IN1(g2879), .IN2(g8249), .QN(n14187) );
  NAND2X0 U15130 ( .IN1(n14189), .IN2(n14190), .QN(g19149) );
  NAND2X0 U15131 ( .IN1(n4351), .IN2(g2944), .QN(n14190) );
  NAND2X0 U15132 ( .IN1(g2879), .IN2(g8175), .QN(n14189) );
  NAND2X0 U15133 ( .IN1(n14191), .IN2(n14192), .QN(g19144) );
  NAND2X0 U15134 ( .IN1(n4351), .IN2(g2947), .QN(n14192) );
  NAND2X0 U15135 ( .IN1(g2879), .IN2(g8023), .QN(n14191) );
  NAND2X0 U15136 ( .IN1(n14193), .IN2(n14194), .QN(g18975) );
  NAND2X0 U15137 ( .IN1(n4351), .IN2(g2195), .QN(n14194) );
  NAND2X0 U15138 ( .IN1(g2879), .IN2(g2981), .QN(n14193) );
  NAND2X0 U15139 ( .IN1(n14195), .IN2(n14196), .QN(g18968) );
  NAND2X0 U15140 ( .IN1(n4351), .IN2(g2190), .QN(n14196) );
  NAND2X0 U15141 ( .IN1(g2879), .IN2(g2978), .QN(n14195) );
  NAND2X0 U15142 ( .IN1(n14197), .IN2(n14198), .QN(g18957) );
  NAND2X0 U15143 ( .IN1(n4351), .IN2(g2165), .QN(n14198) );
  NAND2X0 U15144 ( .IN1(g2879), .IN2(g2963), .QN(n14197) );
  NAND2X0 U15145 ( .IN1(n14199), .IN2(n14200), .QN(g18942) );
  NAND2X0 U15146 ( .IN1(g2879), .IN2(g2975), .QN(n14200) );
  NAND2X0 U15147 ( .IN1(n4351), .IN2(g2185), .QN(n14199) );
  NAND2X0 U15148 ( .IN1(n14201), .IN2(n14202), .QN(g18907) );
  NAND2X0 U15149 ( .IN1(n4365), .IN2(g3061), .QN(n14202) );
  NAND2X0 U15150 ( .IN1(g2987), .IN2(g2997), .QN(n14201) );
  NAND2X0 U15151 ( .IN1(n14203), .IN2(n14204), .QN(g18906) );
  NAND2X0 U15152 ( .IN1(n4351), .IN2(g2180), .QN(n14204) );
  NAND2X0 U15153 ( .IN1(g2879), .IN2(g2972), .QN(n14203) );
  NAND2X0 U15154 ( .IN1(n14205), .IN2(n14206), .QN(g18885) );
  NAND2X0 U15155 ( .IN1(g2879), .IN2(g2874), .QN(n14206) );
  NAND2X0 U15156 ( .IN1(n4351), .IN2(g2200), .QN(n14205) );
  NAND2X0 U15157 ( .IN1(n14207), .IN2(n14208), .QN(g18883) );
  NAND2X0 U15158 ( .IN1(n4351), .IN2(g1471), .QN(n14208) );
  NAND2X0 U15159 ( .IN1(g2879), .IN2(g2935), .QN(n14207) );
  NAND2X0 U15160 ( .IN1(n14209), .IN2(n14210), .QN(g18868) );
  NAND2X0 U15161 ( .IN1(n4365), .IN2(g3060), .QN(n14210) );
  NAND2X0 U15162 ( .IN1(g2987), .IN2(g3078), .QN(n14209) );
  NAND2X0 U15163 ( .IN1(n14211), .IN2(n14212), .QN(g18867) );
  NAND2X0 U15164 ( .IN1(g2879), .IN2(g2969), .QN(n14212) );
  NAND2X0 U15165 ( .IN1(n4351), .IN2(g2175), .QN(n14211) );
  NAND2X0 U15166 ( .IN1(n14213), .IN2(n14214), .QN(g18866) );
  NAND2X0 U15167 ( .IN1(n4351), .IN2(g1476), .QN(n14214) );
  NAND2X0 U15168 ( .IN1(g2879), .IN2(g2938), .QN(n14213) );
  NAND2X0 U15169 ( .IN1(n14215), .IN2(n14216), .QN(g18852) );
  NAND2X0 U15170 ( .IN1(g2879), .IN2(g2941), .QN(n14216) );
  NAND2X0 U15171 ( .IN1(n4351), .IN2(g1481), .QN(n14215) );
  NAND2X0 U15172 ( .IN1(n14217), .IN2(n14218), .QN(g18837) );
  NAND2X0 U15173 ( .IN1(n4365), .IN2(g3059), .QN(n14218) );
  NAND2X0 U15174 ( .IN1(g2987), .IN2(g3077), .QN(n14217) );
  NAND2X0 U15175 ( .IN1(n14219), .IN2(n14220), .QN(g18836) );
  NAND2X0 U15176 ( .IN1(n4351), .IN2(g2170), .QN(n14220) );
  NAND2X0 U15177 ( .IN1(test_so2), .IN2(g2879), .QN(n14219) );
  NAND2X0 U15178 ( .IN1(n14221), .IN2(n14222), .QN(g18835) );
  NAND2X0 U15179 ( .IN1(n4351), .IN2(g1486), .QN(n14222) );
  NAND2X0 U15180 ( .IN1(g2879), .IN2(g2944), .QN(n14221) );
  NAND2X0 U15181 ( .IN1(n14223), .IN2(n14224), .QN(g18821) );
  NAND2X0 U15182 ( .IN1(g2879), .IN2(g2947), .QN(n14224) );
  NAND2X0 U15183 ( .IN1(n4351), .IN2(g1491), .QN(n14223) );
  NAND2X0 U15184 ( .IN1(n14225), .IN2(n14226), .QN(g18820) );
  NAND2X0 U15185 ( .IN1(n4299), .IN2(g2584), .QN(n14226) );
  NAND2X0 U15186 ( .IN1(g2624), .IN2(g2631), .QN(n14225) );
  NAND2X0 U15187 ( .IN1(n14227), .IN2(n14228), .QN(g18804) );
  NAND2X0 U15188 ( .IN1(n4365), .IN2(g3058), .QN(n14228) );
  NAND2X0 U15189 ( .IN1(g2987), .IN2(g3076), .QN(n14227) );
  NAND2X0 U15190 ( .IN1(n14229), .IN2(n14230), .QN(g18803) );
  NAND2X0 U15191 ( .IN1(n4351), .IN2(g1496), .QN(n14230) );
  NAND2X0 U15192 ( .IN1(g2879), .IN2(g2953), .QN(n14229) );
  NAND2X0 U15193 ( .IN1(n14231), .IN2(n14232), .QN(g18794) );
  NAND2X0 U15194 ( .IN1(g1937), .IN2(g1930), .QN(n14232) );
  NAND2X0 U15195 ( .IN1(n4366), .IN2(g1890), .QN(n14231) );
  NAND2X0 U15196 ( .IN1(n14233), .IN2(n14234), .QN(g18782) );
  NAND2X0 U15197 ( .IN1(g3109), .IN2(g559), .QN(n14234) );
  NAND2X0 U15198 ( .IN1(n4494), .IN2(g3084), .QN(n14233) );
  NAND2X0 U15199 ( .IN1(n14235), .IN2(n14236), .QN(g18781) );
  NAND2X0 U15200 ( .IN1(n4351), .IN2(g1501), .QN(n14236) );
  NAND2X0 U15201 ( .IN1(g2879), .IN2(g2956), .QN(n14235) );
  NAND2X0 U15202 ( .IN1(n14237), .IN2(n14238), .QN(g18780) );
  NAND2X0 U15203 ( .IN1(n4299), .IN2(g2631), .QN(n14238) );
  NAND2X0 U15204 ( .IN1(n7990), .IN2(g2624), .QN(n14237) );
  NAND2X0 U15205 ( .IN1(n14239), .IN2(n14240), .QN(g18763) );
  NAND2X0 U15206 ( .IN1(n4300), .IN2(g1196), .QN(n14240) );
  NAND2X0 U15207 ( .IN1(g1236), .IN2(g1243), .QN(n14239) );
  NAND2X0 U15208 ( .IN1(n14241), .IN2(n14242), .QN(g18755) );
  NAND2X0 U15209 ( .IN1(n4365), .IN2(g3057), .QN(n14242) );
  NAND2X0 U15210 ( .IN1(g2987), .IN2(g3075), .QN(n14241) );
  NAND2X0 U15211 ( .IN1(n14243), .IN2(n14244), .QN(g18754) );
  NAND2X0 U15212 ( .IN1(g2879), .IN2(g2959), .QN(n14244) );
  NAND2X0 U15213 ( .IN1(n4351), .IN2(g1506), .QN(n14243) );
  NAND2X0 U15214 ( .IN1(n14245), .IN2(n14246), .QN(g18743) );
  NAND2X0 U15215 ( .IN1(n7991), .IN2(g1930), .QN(n14246) );
  NAND2X0 U15216 ( .IN1(n4366), .IN2(g1937), .QN(n14245) );
  NAND2X0 U15217 ( .IN1(n14247), .IN2(n14248), .QN(g18726) );
  NAND2X0 U15218 ( .IN1(test_so22), .IN2(n4313), .QN(n14248) );
  NAND2X0 U15219 ( .IN1(g550), .IN2(g557), .QN(n14247) );
  NAND2X0 U15220 ( .IN1(n14249), .IN2(n14250), .QN(g18719) );
  NAND2X0 U15221 ( .IN1(n4383), .IN2(g3211), .QN(n14250) );
  NAND2X0 U15222 ( .IN1(g8030), .IN2(g559), .QN(n14249) );
  NAND2X0 U15223 ( .IN1(n14251), .IN2(n14252), .QN(g18707) );
  NAND2X0 U15224 ( .IN1(n4300), .IN2(g1243), .QN(n14252) );
  NAND2X0 U15225 ( .IN1(n7992), .IN2(g1236), .QN(n14251) );
  NAND2X0 U15226 ( .IN1(n14253), .IN2(n14254), .QN(g18678) );
  NAND2X0 U15227 ( .IN1(n4313), .IN2(g557), .QN(n14254) );
  NAND2X0 U15228 ( .IN1(n7993), .IN2(g550), .QN(n14253) );
  NAND2X0 U15229 ( .IN1(n14255), .IN2(n14256), .QN(g18669) );
  NAND2X0 U15230 ( .IN1(n4382), .IN2(test_so6), .QN(n14256) );
  NAND2X0 U15231 ( .IN1(g8106), .IN2(g559), .QN(n14255) );
  NAND2X0 U15232 ( .IN1(n14257), .IN2(n14258), .QN(g17429) );
  NAND2X0 U15233 ( .IN1(g3109), .IN2(g2574), .QN(n14258) );
  NAND2X0 U15234 ( .IN1(n4494), .IN2(g3088), .QN(n14257) );
  NAND2X0 U15235 ( .IN1(n14259), .IN2(n14260), .QN(g17383) );
  NAND2X0 U15236 ( .IN1(n4494), .IN2(test_so8), .QN(n14260) );
  NAND2X0 U15237 ( .IN1(g3109), .IN2(g1880), .QN(n14259) );
  NAND2X0 U15238 ( .IN1(n14261), .IN2(n14262), .QN(g17341) );
  NAND2X0 U15239 ( .IN1(n4383), .IN2(g3185), .QN(n14262) );
  NAND2X0 U15240 ( .IN1(g8030), .IN2(g2574), .QN(n14261) );
  NAND2X0 U15241 ( .IN1(n14263), .IN2(n14264), .QN(g17340) );
  NAND2X0 U15242 ( .IN1(g3109), .IN2(g1186), .QN(n14264) );
  NAND2X0 U15243 ( .IN1(n4494), .IN2(g3170), .QN(n14263) );
  NAND2X0 U15244 ( .IN1(n14265), .IN2(n14266), .QN(g17303) );
  NAND2X0 U15245 ( .IN1(n4383), .IN2(g3176), .QN(n14266) );
  NAND2X0 U15246 ( .IN1(g8030), .IN2(g1880), .QN(n14265) );
  NAND2X0 U15247 ( .IN1(n14267), .IN2(n14268), .QN(g17302) );
  NAND2X0 U15248 ( .IN1(g3109), .IN2(g499), .QN(n14268) );
  NAND2X0 U15249 ( .IN1(n4494), .IN2(g3161), .QN(n14267) );
  NAND2X0 U15250 ( .IN1(n14269), .IN2(n14270), .QN(g17271) );
  NAND2X0 U15251 ( .IN1(n4382), .IN2(g3182), .QN(n14270) );
  NAND2X0 U15252 ( .IN1(g8106), .IN2(g2574), .QN(n14269) );
  NAND2X0 U15253 ( .IN1(n14271), .IN2(n14272), .QN(g17270) );
  NAND2X0 U15254 ( .IN1(g8030), .IN2(g1186), .QN(n14272) );
  NAND2X0 U15255 ( .IN1(n4383), .IN2(g3167), .QN(n14271) );
  NAND2X0 U15256 ( .IN1(n14273), .IN2(n14274), .QN(g17269) );
  NAND2X0 U15257 ( .IN1(g3109), .IN2(g2633), .QN(n14274) );
  NAND2X0 U15258 ( .IN1(n4494), .IN2(g3096), .QN(n14273) );
  NAND2X0 U15259 ( .IN1(n14275), .IN2(n14276), .QN(g17248) );
  NAND2X0 U15260 ( .IN1(g8106), .IN2(g1880), .QN(n14276) );
  NAND2X0 U15261 ( .IN1(n4382), .IN2(g3173), .QN(n14275) );
  NAND2X0 U15262 ( .IN1(n14277), .IN2(n14278), .QN(g17247) );
  NAND2X0 U15263 ( .IN1(n4383), .IN2(g3158), .QN(n14278) );
  NAND2X0 U15264 ( .IN1(g8030), .IN2(g499), .QN(n14277) );
  NAND2X0 U15265 ( .IN1(n14279), .IN2(n14280), .QN(g17246) );
  NAND2X0 U15266 ( .IN1(g3109), .IN2(g1939), .QN(n14280) );
  NAND2X0 U15267 ( .IN1(n4494), .IN2(g3093), .QN(n14279) );
  NAND2X0 U15268 ( .IN1(n14281), .IN2(n14282), .QN(g17236) );
  NAND2X0 U15269 ( .IN1(g8106), .IN2(g1186), .QN(n14282) );
  NAND2X0 U15270 ( .IN1(n4382), .IN2(g3164), .QN(n14281) );
  NAND2X0 U15271 ( .IN1(n14283), .IN2(n14284), .QN(g17235) );
  NAND2X0 U15272 ( .IN1(n4383), .IN2(g3095), .QN(n14284) );
  NAND2X0 U15273 ( .IN1(g8030), .IN2(g2633), .QN(n14283) );
  NAND2X0 U15274 ( .IN1(n14285), .IN2(n14286), .QN(g17234) );
  NAND2X0 U15275 ( .IN1(g3109), .IN2(g1245), .QN(n14286) );
  NAND2X0 U15276 ( .IN1(n4494), .IN2(g3087), .QN(n14285) );
  NAND2X0 U15277 ( .IN1(n14287), .IN2(n14288), .QN(g17229) );
  NAND2X0 U15278 ( .IN1(n4382), .IN2(g3155), .QN(n14288) );
  NAND2X0 U15279 ( .IN1(g8106), .IN2(g499), .QN(n14287) );
  NAND2X0 U15280 ( .IN1(n14289), .IN2(n14290), .QN(g17228) );
  NAND2X0 U15281 ( .IN1(n4383), .IN2(g3092), .QN(n14290) );
  NAND2X0 U15282 ( .IN1(g8030), .IN2(g1939), .QN(n14289) );
  NAND2X0 U15283 ( .IN1(n14291), .IN2(n14292), .QN(g17226) );
  NAND2X0 U15284 ( .IN1(n4382), .IN2(g3094), .QN(n14292) );
  NAND2X0 U15285 ( .IN1(g8106), .IN2(g2633), .QN(n14291) );
  NAND2X0 U15286 ( .IN1(n14293), .IN2(n14294), .QN(g17225) );
  NAND2X0 U15287 ( .IN1(g8030), .IN2(g1245), .QN(n14294) );
  NAND2X0 U15288 ( .IN1(n4383), .IN2(g3086), .QN(n14293) );
  NAND2X0 U15289 ( .IN1(n14295), .IN2(n14296), .QN(g17224) );
  NAND2X0 U15290 ( .IN1(n4382), .IN2(g3091), .QN(n14296) );
  NAND2X0 U15291 ( .IN1(g8106), .IN2(g1939), .QN(n14295) );
  NAND2X0 U15292 ( .IN1(n14297), .IN2(n14298), .QN(g17222) );
  NAND2X0 U15293 ( .IN1(g8106), .IN2(g1245), .QN(n14298) );
  NAND2X0 U15294 ( .IN1(n4382), .IN2(g3085), .QN(n14297) );
  NAND2X0 U15295 ( .IN1(n14299), .IN2(n14300), .QN(g16880) );
  NAND2X0 U15296 ( .IN1(n4365), .IN2(g3056), .QN(n14300) );
  NAND2X0 U15297 ( .IN1(g2987), .IN2(g3074), .QN(n14299) );
  NAND2X0 U15298 ( .IN1(n14301), .IN2(n14302), .QN(g16866) );
  NAND2X0 U15299 ( .IN1(n4365), .IN2(g3051), .QN(n14302) );
  NAND2X0 U15300 ( .IN1(test_so97), .IN2(g2987), .QN(n14301) );
  NAND2X0 U15301 ( .IN1(n14303), .IN2(n14304), .QN(g16861) );
  NAND2X0 U15302 ( .IN1(test_so96), .IN2(n4365), .QN(n14304) );
  NAND2X0 U15303 ( .IN1(g2987), .IN2(g3073), .QN(n14303) );
  NAND2X0 U15304 ( .IN1(n14305), .IN2(n14306), .QN(g16860) );
  NAND2X0 U15305 ( .IN1(n4365), .IN2(g3046), .QN(n14306) );
  NAND2X0 U15306 ( .IN1(g2987), .IN2(g3065), .QN(n14305) );
  NAND2X0 U15307 ( .IN1(n14307), .IN2(n14308), .QN(g16857) );
  NAND2X0 U15308 ( .IN1(n4365), .IN2(g3050), .QN(n14308) );
  NAND2X0 U15309 ( .IN1(g2987), .IN2(g3069), .QN(n14307) );
  NAND2X0 U15310 ( .IN1(n14309), .IN2(n14310), .QN(g16854) );
  NAND2X0 U15311 ( .IN1(n4365), .IN2(g3053), .QN(n14310) );
  NAND2X0 U15312 ( .IN1(g2987), .IN2(g3072), .QN(n14309) );
  NAND2X0 U15313 ( .IN1(n14311), .IN2(n14312), .QN(g16853) );
  NAND2X0 U15314 ( .IN1(n4365), .IN2(g3045), .QN(n14312) );
  NAND2X0 U15315 ( .IN1(g2987), .IN2(g3064), .QN(n14311) );
  NAND2X0 U15316 ( .IN1(n14313), .IN2(n14314), .QN(g16851) );
  NAND2X0 U15317 ( .IN1(n4365), .IN2(g3049), .QN(n14314) );
  NAND2X0 U15318 ( .IN1(g2987), .IN2(g3068), .QN(n14313) );
  NAND2X0 U15319 ( .IN1(n14315), .IN2(n14316), .QN(g16845) );
  NAND2X0 U15320 ( .IN1(n4365), .IN2(g3052), .QN(n14316) );
  NAND2X0 U15321 ( .IN1(g2987), .IN2(g3071), .QN(n14315) );
  NAND2X0 U15322 ( .IN1(n14317), .IN2(n14318), .QN(g16844) );
  NAND2X0 U15323 ( .IN1(n4365), .IN2(g3044), .QN(n14318) );
  NAND2X0 U15324 ( .IN1(g2987), .IN2(g3063), .QN(n14317) );
  NAND2X0 U15325 ( .IN1(n14319), .IN2(n14320), .QN(g16835) );
  NAND2X0 U15326 ( .IN1(n4365), .IN2(g3048), .QN(n14320) );
  NAND2X0 U15327 ( .IN1(g2987), .IN2(g3067), .QN(n14319) );
  NAND2X0 U15328 ( .IN1(n14321), .IN2(n14322), .QN(g16824) );
  NAND2X0 U15329 ( .IN1(n4365), .IN2(g3043), .QN(n14322) );
  NAND2X0 U15330 ( .IN1(g2987), .IN2(g3062), .QN(n14321) );
  NOR2X0 U15331 ( .IN1(g51), .IN2(DFF_1_n1), .QN(g16823) );
  NAND2X0 U15332 ( .IN1(n14323), .IN2(n14324), .QN(g16803) );
  NAND2X0 U15333 ( .IN1(n4365), .IN2(g3047), .QN(n14324) );
  NAND2X0 U15334 ( .IN1(g2987), .IN2(g3066), .QN(n14323) );
  NOR2X0 U15335 ( .IN1(n4423), .IN2(g51), .QN(g16802) );
  NAND2X0 U15336 ( .IN1(n14325), .IN2(n14326), .QN(g16718) );
  NAND2X0 U15337 ( .IN1(n4292), .IN2(g2704), .QN(n14326) );
  NAND2X0 U15338 ( .IN1(g2703), .IN2(g2584), .QN(n14325) );
  NAND2X0 U15339 ( .IN1(n14327), .IN2(n14328), .QN(g16692) );
  NAND2X0 U15340 ( .IN1(n4293), .IN2(g2010), .QN(n14328) );
  NAND2X0 U15341 ( .IN1(g2009), .IN2(g1890), .QN(n14327) );
  NAND2X0 U15342 ( .IN1(n14329), .IN2(n14330), .QN(g16671) );
  NAND2X0 U15343 ( .IN1(n4294), .IN2(g1316), .QN(n14330) );
  NAND2X0 U15344 ( .IN1(g1315), .IN2(g1196), .QN(n14329) );
  NAND2X0 U15345 ( .IN1(n14331), .IN2(n14332), .QN(g16654) );
  NAND2X0 U15346 ( .IN1(n4295), .IN2(g630), .QN(n14332) );
  NAND2X0 U15347 ( .IN1(test_so22), .IN2(g629), .QN(n14331) );
  NAND2X0 U15348 ( .IN1(n14333), .IN2(g2987), .QN(g16496) );
  NAND2X0 U15349 ( .IN1(DFF_1612_n1), .IN2(g5388), .QN(n14333) );
  NOR3X0 U15350 ( .IN1(n14334), .IN2(n14335), .IN3(n14336), .QN(g13194) );
  NOR2X0 U15351 ( .IN1(n4314), .IN2(test_so87), .QN(n14336) );
  NOR2X0 U15352 ( .IN1(n4370), .IN2(g2561), .QN(n14335) );
  NOR2X0 U15353 ( .IN1(n4299), .IN2(g2562), .QN(n14334) );
  NOR3X0 U15354 ( .IN1(n14337), .IN2(n14338), .IN3(n14339), .QN(g13182) );
  NOR2X0 U15355 ( .IN1(n4366), .IN2(g1868), .QN(n14339) );
  NOR2X0 U15356 ( .IN1(n4296), .IN2(g1869), .QN(n14338) );
  NOR2X0 U15357 ( .IN1(n4315), .IN2(g1867), .QN(n14337) );
  NOR3X0 U15358 ( .IN1(n14340), .IN2(n14341), .IN3(n14342), .QN(g13175) );
  NOR2X0 U15359 ( .IN1(n4299), .IN2(g2553), .QN(n14342) );
  NOR2X0 U15360 ( .IN1(n4314), .IN2(g2554), .QN(n14341) );
  NOR2X0 U15361 ( .IN1(n4370), .IN2(g2552), .QN(n14340) );
  NOR3X0 U15362 ( .IN1(n14343), .IN2(n14344), .IN3(n14345), .QN(g13171) );
  NOR2X0 U15363 ( .IN1(n4300), .IN2(test_so44), .QN(n14345) );
  NOR2X0 U15364 ( .IN1(n4316), .IN2(g1173), .QN(n14344) );
  NOR2X0 U15365 ( .IN1(n4371), .IN2(g1175), .QN(n14343) );
  NOR3X0 U15366 ( .IN1(n14346), .IN2(n14347), .IN3(n14348), .QN(g13164) );
  NOR2X0 U15367 ( .IN1(n4366), .IN2(g1859), .QN(n14348) );
  NOR2X0 U15368 ( .IN1(n4296), .IN2(g1860), .QN(n14347) );
  NOR2X0 U15369 ( .IN1(n4315), .IN2(g1858), .QN(n14346) );
  NOR3X0 U15370 ( .IN1(n14349), .IN2(n14350), .IN3(n14351), .QN(g13160) );
  NOR2X0 U15371 ( .IN1(n4313), .IN2(g487), .QN(n14351) );
  NOR2X0 U15372 ( .IN1(n4298), .IN2(g488), .QN(n14350) );
  NOR2X0 U15373 ( .IN1(n4372), .IN2(g486), .QN(n14349) );
  NOR3X0 U15374 ( .IN1(n14352), .IN2(n14353), .IN3(n14354), .QN(g13155) );
  NOR2X0 U15375 ( .IN1(n4300), .IN2(g1165), .QN(n14354) );
  NOR2X0 U15376 ( .IN1(n4371), .IN2(g1166), .QN(n14353) );
  NOR2X0 U15377 ( .IN1(n4316), .IN2(g1164), .QN(n14352) );
  NOR3X0 U15378 ( .IN1(n14355), .IN2(n14356), .IN3(n14357), .QN(g13149) );
  NOR2X0 U15379 ( .IN1(n4313), .IN2(g478), .QN(n14357) );
  NOR2X0 U15380 ( .IN1(n4298), .IN2(g479), .QN(n14356) );
  NOR2X0 U15381 ( .IN1(n4372), .IN2(g477), .QN(n14355) );
  NOR3X0 U15382 ( .IN1(n14358), .IN2(n14359), .IN3(n14360), .QN(g13143) );
  NOR2X0 U15383 ( .IN1(n4299), .IN2(g2559), .QN(n14360) );
  NOR2X0 U15384 ( .IN1(n4314), .IN2(g2539), .QN(n14359) );
  NOR2X0 U15385 ( .IN1(n4370), .IN2(g2555), .QN(n14358) );
  NOR3X0 U15386 ( .IN1(n14361), .IN2(n14362), .IN3(n14363), .QN(g13135) );
  NOR2X0 U15387 ( .IN1(n4366), .IN2(g1865), .QN(n14363) );
  NOR2X0 U15388 ( .IN1(n4296), .IN2(g1845), .QN(n14362) );
  NOR2X0 U15389 ( .IN1(n4315), .IN2(g1861), .QN(n14361) );
  NOR3X0 U15390 ( .IN1(n14364), .IN2(n14365), .IN3(n14366), .QN(g13124) );
  NOR2X0 U15391 ( .IN1(n4300), .IN2(g1171), .QN(n14366) );
  NOR2X0 U15392 ( .IN1(n4371), .IN2(g1151), .QN(n14365) );
  NOR2X0 U15393 ( .IN1(n4316), .IN2(g1167), .QN(n14364) );
  NOR3X0 U15394 ( .IN1(n14367), .IN2(n14368), .IN3(n14369), .QN(g13111) );
  NOR2X0 U15395 ( .IN1(n4313), .IN2(g484), .QN(n14369) );
  NOR2X0 U15396 ( .IN1(n4298), .IN2(g464), .QN(n14368) );
  NOR2X0 U15397 ( .IN1(n4372), .IN2(g480), .QN(n14367) );
  XOR2X1 U15398 ( .IN1(n8034), .IN2(n8743), .Q(N995) );
  XNOR3X1 U15399 ( .IN1(n14370), .IN2(n14371), .IN3(n14372), .Q(n8743) );
  XOR3X1 U15400 ( .IN1(n14389), .IN2(n14390), .IN3(n14373), .Q(n14372) );
  XOR2X1 U15401 ( .IN1(g8275), .IN2(test_so99), .Q(n14373) );
  XOR2X1 U15402 ( .IN1(n8030), .IN2(n8029), .Q(n14371) );
  XOR2X1 U15403 ( .IN1(n14391), .IN2(n8031), .Q(n14370) );
  XOR2X1 U15404 ( .IN1(n8746), .IN2(n8032), .Q(N690) );
  XOR3X1 U15405 ( .IN1(n14374), .IN2(n14375), .IN3(n14376), .Q(n8746) );
  XOR3X1 U15406 ( .IN1(n14393), .IN2(n14394), .IN3(n14377), .Q(n14376) );
  XOR2X1 U15407 ( .IN1(g8262), .IN2(n14392), .Q(n14377) );
  XOR2X1 U15408 ( .IN1(n7995), .IN2(n7994), .Q(n14375) );
  XOR2X1 U15409 ( .IN1(n7997), .IN2(n7996), .Q(n14374) );
  NOR2X0 U3772_U2 ( .IN1(n2230), .IN2(n2217), .QN(U3772_n1) );
  INVX0 U3772_U1 ( .INP(U3772_n1), .ZN(n2231) );
  NOR2X0 U3776_U2 ( .IN1(n2374), .IN2(n2361), .QN(U3776_n1) );
  INVX0 U3776_U1 ( .INP(U3776_n1), .ZN(n2375) );
  NOR2X0 U3777_U2 ( .IN1(g51), .IN2(DFF_2_n1), .QN(U3777_n1) );
  INVX0 U3777_U1 ( .INP(U3777_n1), .ZN(n4264) );
  NOR2X0 U3778_U2 ( .IN1(n2445), .IN2(n2446), .QN(U3778_n1) );
  INVX0 U3778_U1 ( .INP(U3778_n1), .ZN(n2440) );
  NOR2X0 U3779_U2 ( .IN1(n472), .IN2(n2446), .QN(U3779_n1) );
  INVX0 U3779_U1 ( .INP(U3779_n1), .ZN(n2426) );
  NOR2X0 U3780_U2 ( .IN1(n2670), .IN2(n2671), .QN(U3780_n1) );
  INVX0 U3780_U1 ( .INP(U3780_n1), .ZN(n2669) );
  NOR2X0 U3781_U2 ( .IN1(n2685), .IN2(n2686), .QN(U3781_n1) );
  INVX0 U3781_U1 ( .INP(U3781_n1), .ZN(n2684) );
  NOR2X0 U3782_U2 ( .IN1(n2718), .IN2(n2719), .QN(U3782_n1) );
  INVX0 U3782_U1 ( .INP(U3782_n1), .ZN(n2717) );
  NOR2X0 U3783_U2 ( .IN1(n2982), .IN2(g2124), .QN(U3783_n1) );
  INVX0 U3783_U1 ( .INP(U3783_n1), .ZN(n2981) );
  NOR2X0 U3784_U2 ( .IN1(n2985), .IN2(g1430), .QN(U3784_n1) );
  INVX0 U3784_U1 ( .INP(U3784_n1), .ZN(n2984) );
  NOR2X0 U3785_U2 ( .IN1(n2988), .IN2(g744), .QN(U3785_n1) );
  INVX0 U3785_U1 ( .INP(U3785_n1), .ZN(n2987) );
  NOR2X0 U3786_U2 ( .IN1(n2991), .IN2(g56), .QN(U3786_n1) );
  INVX0 U3786_U1 ( .INP(U3786_n1), .ZN(n2990) );
  NOR2X0 U3787_U2 ( .IN1(n3742), .IN2(test_so98), .QN(U3787_n1) );
  INVX0 U3787_U1 ( .INP(U3787_n1), .ZN(n3741) );
  NOR2X0 U3901_U2 ( .IN1(n2302), .IN2(n2289), .QN(U3901_n1) );
  INVX0 U3901_U1 ( .INP(U3901_n1), .ZN(n2303) );
  NOR2X0 U3902_U2 ( .IN1(n494), .IN2(n2289), .QN(U3902_n1) );
  INVX0 U3902_U1 ( .INP(U3902_n1), .ZN(n2275) );
  INVX0 U4467_U2 ( .INP(n1396), .ZN(U4467_n1) );
  NOR2X0 U4467_U1 ( .IN1(n3254), .IN2(U4467_n1), .QN(n3252) );
  INVX0 U4904_U2 ( .INP(n2800), .ZN(U4904_n1) );
  NOR2X0 U4904_U1 ( .IN1(n163), .IN2(U4904_n1), .QN(n2798) );
  INVX0 U4930_U2 ( .INP(n2616), .ZN(U4930_n1) );
  NOR2X0 U4930_U1 ( .IN1(n163), .IN2(U4930_n1), .QN(n2594) );
  INVX0 U5128_U2 ( .INP(n3933), .ZN(U5128_n1) );
  NOR2X0 U5128_U1 ( .IN1(n4406), .IN2(U5128_n1), .QN(n3940) );
  INVX0 U5141_U2 ( .INP(n3939), .ZN(U5141_n1) );
  NOR2X0 U5141_U1 ( .IN1(n4405), .IN2(U5141_n1), .QN(n3936) );
  INVX0 U5749_U2 ( .INP(g2133), .ZN(U5749_n1) );
  NOR2X0 U5749_U1 ( .IN1(n3160), .IN2(U5749_n1), .QN(n3159) );
  INVX0 U5750_U2 ( .INP(g1439), .ZN(U5750_n1) );
  NOR2X0 U5750_U1 ( .IN1(n3164), .IN2(U5750_n1), .QN(n3163) );
  INVX0 U5751_U2 ( .INP(g753), .ZN(U5751_n1) );
  NOR2X0 U5751_U1 ( .IN1(n3168), .IN2(U5751_n1), .QN(n3167) );
  INVX0 U5752_U2 ( .INP(g65), .ZN(U5752_n1) );
  NOR2X0 U5752_U1 ( .IN1(n3172), .IN2(U5752_n1), .QN(n3171) );
  INVX0 U5753_U2 ( .INP(g2142), .ZN(U5753_n1) );
  NOR2X0 U5753_U1 ( .IN1(n4522), .IN2(U5753_n1), .QN(n3424) );
  INVX0 U5754_U2 ( .INP(g2151), .ZN(U5754_n1) );
  NOR2X0 U5754_U1 ( .IN1(n4526), .IN2(U5754_n1), .QN(n3683) );
  INVX0 U5755_U2 ( .INP(g2160), .ZN(U5755_n1) );
  NOR2X0 U5755_U1 ( .IN1(n3888), .IN2(U5755_n1), .QN(n3887) );
  INVX0 U5756_U2 ( .INP(g1448), .ZN(U5756_n1) );
  NOR2X0 U5756_U1 ( .IN1(n4523), .IN2(U5756_n1), .QN(n3427) );
  INVX0 U5757_U2 ( .INP(g1457), .ZN(U5757_n1) );
  NOR2X0 U5757_U1 ( .IN1(n4527), .IN2(U5757_n1), .QN(n3686) );
  INVX0 U5758_U2 ( .INP(g1466), .ZN(U5758_n1) );
  NOR2X0 U5758_U1 ( .IN1(n3891), .IN2(U5758_n1), .QN(n3890) );
  INVX0 U5759_U2 ( .INP(g762), .ZN(U5759_n1) );
  NOR2X0 U5759_U1 ( .IN1(n3431), .IN2(U5759_n1), .QN(n3430) );
  INVX0 U5760_U2 ( .INP(g771), .ZN(U5760_n1) );
  NOR2X0 U5760_U1 ( .IN1(n3690), .IN2(U5760_n1), .QN(n3689) );
  INVX0 U5761_U2 ( .INP(g780), .ZN(U5761_n1) );
  NOR2X0 U5761_U1 ( .IN1(n3894), .IN2(U5761_n1), .QN(n3893) );
  INVX0 U5762_U2 ( .INP(g74), .ZN(U5762_n1) );
  NOR2X0 U5762_U1 ( .IN1(n4521), .IN2(U5762_n1), .QN(n3433) );
  INVX0 U5763_U2 ( .INP(g83), .ZN(U5763_n1) );
  NOR2X0 U5763_U1 ( .IN1(n4528), .IN2(U5763_n1), .QN(n3692) );
  INVX0 U5764_U2 ( .INP(g92), .ZN(U5764_n1) );
  NOR2X0 U5764_U1 ( .IN1(n3897), .IN2(U5764_n1), .QN(n3896) );
  INVX0 U5882_U2 ( .INP(n1547), .ZN(U5882_n1) );
  NOR2X0 U5882_U1 ( .IN1(g3036), .IN2(U5882_n1), .QN(n4101) );
  INVX0 U5939_U2 ( .INP(g2257), .ZN(U5939_n1) );
  NOR2X0 U5939_U1 ( .IN1(n1269), .IN2(U5939_n1), .QN(n3038) );
  INVX0 U5940_U2 ( .INP(g1563), .ZN(U5940_n1) );
  NOR2X0 U5940_U1 ( .IN1(n971), .IN2(U5940_n1), .QN(n3070) );
  INVX0 U5941_U2 ( .INP(g869), .ZN(U5941_n1) );
  NOR2X0 U5941_U1 ( .IN1(n672), .IN2(U5941_n1), .QN(n3102) );
  INVX0 U5942_U2 ( .INP(g181), .ZN(U5942_n1) );
  NOR2X0 U5942_U1 ( .IN1(n328), .IN2(U5942_n1), .QN(n3130) );
  INVX0 U6140_U2 ( .INP(g3002), .ZN(U6140_n1) );
  NOR2X0 U6140_U1 ( .IN1(n4066), .IN2(U6140_n1), .QN(n4065) );
  INVX0 U6460_U2 ( .INP(g3233), .ZN(U6460_n1) );
  NOR2X0 U6460_U1 ( .IN1(g3230), .IN2(U6460_n1), .QN(n3700) );
  INVX0 U6470_U2 ( .INP(g2892), .ZN(U6470_n1) );
  NOR2X0 U6470_U1 ( .IN1(n4305), .IN2(U6470_n1), .QN(n4182) );
  INVX0 U6562_U2 ( .INP(n3938), .ZN(U6562_n1) );
  NOR2X0 U6562_U1 ( .IN1(g3204), .IN2(U6562_n1), .QN(n3939) );
  INVX0 U6563_U2 ( .INP(n4073), .ZN(U6563_n1) );
  NOR2X0 U6563_U1 ( .IN1(g3204), .IN2(U6563_n1), .QN(n3705) );
  INVX0 U6718_U2 ( .INP(n285), .ZN(U6718_n1) );
  NOR2X0 U6718_U1 ( .IN1(g3197), .IN2(U6718_n1), .QN(n4073) );
  INVX0 U7116_U2 ( .INP(n4058), .ZN(U7116_n1) );
  NOR2X0 U7116_U1 ( .IN1(g2903), .IN2(U7116_n1), .QN(n4057) );
  INVX0 U7118_U2 ( .INP(n10), .ZN(U7118_n1) );
  NOR2X0 U7118_U1 ( .IN1(g2896), .IN2(U7118_n1), .QN(n4122) );
  INVX0 U7293_U2 ( .INP(n4598), .ZN(U7293_n1) );
  NOR2X0 U7293_U1 ( .IN1(g3234), .IN2(U7293_n1), .QN(g20877) );
endmodule

