module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n595_, new_n614_, new_n445_, new_n699_, new_n236_, new_n479_, new_n608_, new_n847_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n368_, new_n738_, new_n439_, new_n827_, new_n283_, new_n390_, new_n743_, new_n779_, new_n241_, new_n641_, new_n339_, new_n365_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n246_, new_n682_, new_n812_, new_n679_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n419_, new_n728_, new_n624_, new_n534_, new_n819_, new_n637_, new_n451_, new_n489_, new_n424_, new_n804_, new_n853_, new_n602_, new_n695_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n642_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n500_, new_n786_, new_n799_, new_n317_, new_n344_, new_n287_, new_n504_, new_n742_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n774_, new_n716_, new_n701_, new_n792_, new_n257_, new_n481_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n766_, new_n272_, new_n282_, new_n634_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n849_, new_n855_, new_n606_, new_n589_, new_n350_, new_n655_, new_n759_, new_n630_, new_n385_, new_n829_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n764_, new_n683_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n530_, new_n318_, new_n622_, new_n629_, new_n702_, new_n833_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n763_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n674_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n423_, new_n498_, new_n492_, new_n496_, new_n650_, new_n708_, new_n750_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n506_, new_n680_, new_n256_, new_n778_, new_n452_, new_n381_, new_n656_, new_n820_, new_n771_, new_n388_, new_n508_, new_n714_, new_n483_, new_n394_, new_n299_, new_n657_, new_n652_, new_n314_, new_n582_, new_n363_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n398_, new_n301_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n541_, new_n458_, new_n854_, new_n447_, new_n267_, new_n473_, new_n790_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n621_, new_n846_, new_n349_, new_n488_, new_n524_, new_n705_, new_n848_, new_n277_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n438_, new_n696_, new_n632_, new_n671_, new_n528_, new_n572_, new_n850_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n805_, new_n559_, new_n762_, new_n838_, new_n233_, new_n469_, new_n391_, new_n437_, new_n295_, new_n359_, new_n794_, new_n628_, new_n409_, new_n745_, new_n457_, new_n553_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n448_, new_n276_, new_n688_, new_n384_, new_n410_, new_n851_, new_n543_, new_n775_, new_n371_, new_n509_, new_n454_, new_n296_, new_n661_, new_n308_, new_n633_, new_n797_, new_n232_, new_n784_, new_n724_, new_n860_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n809_, new_n654_, new_n713_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n749_, new_n310_, new_n275_, new_n352_, new_n575_, new_n839_, new_n485_, new_n525_, new_n562_, new_n578_, new_n810_, new_n808_, new_n493_, new_n547_, new_n264_, new_n665_, new_n800_, new_n379_, new_n719_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n824_, new_n520_, new_n253_, new_n717_, new_n403_, new_n237_, new_n825_, new_n858_, new_n557_, new_n260_, new_n251_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n748_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n513_, new_n592_, new_n726_, new_n558_, new_n231_, new_n219_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n428_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n755_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n856_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n499_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n468_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n737_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n337_, new_n623_, new_n446_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n519_, new_n563_, new_n662_, new_n440_, new_n733_, new_n531_, new_n593_, new_n252_, new_n585_, new_n751_, new_n312_, new_n535_, new_n372_, new_n725_, new_n814_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n408_, new_n470_, new_n769_, new_n651_, new_n433_, new_n435_, new_n776_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n815_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n712_, new_n550_, new_n269_, new_n512_, new_n788_, new_n841_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n818_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n754_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n803_, new_n727_, new_n375_, new_n294_, new_n760_, new_n627_, new_n704_, new_n567_, new_n576_, new_n831_, new_n791_, new_n357_, new_n320_, new_n780_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n490_, new_n560_, new_n358_, new_n348_, new_n610_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n226_, new_n802_, new_n697_, new_n709_, new_n373_, new_n540_, new_n434_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n551_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n521_, new_n793_, new_n406_, new_n828_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n573_, new_n765_, new_n405_;

not g000 ( new_n215_, N75 );
nand g001 ( new_n216_, N29, N42 );
nor g002 ( N388, new_n216_, new_n215_ );
not g003 ( new_n218_, N80 );
nand g004 ( new_n219_, N29, N36 );
nor g005 ( N389, new_n219_, new_n218_ );
not g006 ( new_n221_, N42 );
nor g007 ( new_n222_, new_n219_, new_n221_ );
xor g008 ( N390, new_n222_, keyIn_0_6 );
nand g009 ( new_n224_, N85, N86 );
not g010 ( N391, new_n224_ );
not g011 ( new_n226_, N17 );
nand g012 ( new_n227_, N1, N8 );
not g013 ( new_n228_, new_n227_ );
nand g014 ( new_n229_, new_n228_, N13 );
nor g015 ( N418, new_n229_, new_n226_ );
xor g016 ( new_n231_, new_n222_, keyIn_0_0 );
nand g017 ( new_n232_, N1, N26 );
nand g018 ( new_n233_, N13, N17 );
nor g019 ( new_n234_, new_n232_, new_n233_ );
nand g020 ( N419, new_n231_, new_n234_ );
nand g021 ( new_n236_, N59, N75 );
not g022 ( new_n237_, new_n236_ );
nand g023 ( N420, new_n237_, N80 );
nand g024 ( new_n239_, N36, N59 );
nor g025 ( new_n240_, new_n239_, new_n218_ );
xnor g026 ( new_n241_, new_n240_, keyIn_0_8 );
xnor g027 ( N421, new_n241_, keyIn_0_19 );
nor g028 ( new_n243_, new_n239_, new_n221_ );
xnor g029 ( N422, new_n243_, keyIn_0_9 );
not g030 ( new_n245_, N90 );
nor g031 ( new_n246_, N87, N88 );
nor g032 ( new_n247_, new_n246_, new_n245_ );
xor g033 ( N423, new_n247_, keyIn_0_20 );
not g034 ( new_n249_, new_n231_ );
nand g035 ( N446, new_n249_, new_n234_ );
not g036 ( new_n251_, keyIn_0_1 );
not g037 ( new_n252_, new_n232_ );
nand g038 ( new_n253_, new_n252_, N51 );
nand g039 ( new_n254_, new_n253_, new_n251_ );
not g040 ( new_n255_, N51 );
nor g041 ( new_n256_, new_n232_, new_n255_ );
nand g042 ( new_n257_, new_n256_, keyIn_0_1 );
nand g043 ( N447, new_n254_, new_n257_ );
not g044 ( new_n259_, N55 );
nor g045 ( new_n260_, new_n229_, new_n259_ );
xnor g046 ( new_n261_, new_n260_, keyIn_0_3 );
nand g047 ( new_n262_, N29, N68 );
xor g048 ( new_n263_, new_n262_, keyIn_0_4 );
nand g049 ( new_n264_, new_n261_, new_n263_ );
xor g050 ( N448, new_n264_, keyIn_0_27 );
not g051 ( new_n266_, N74 );
nand g052 ( new_n267_, N59, N68 );
nor g053 ( new_n268_, new_n267_, new_n266_ );
xnor g054 ( new_n269_, new_n268_, keyIn_0_5 );
nand g055 ( new_n270_, new_n261_, new_n269_ );
xnor g056 ( N449, new_n270_, keyIn_0_28 );
not g057 ( new_n272_, N89 );
nor g058 ( new_n273_, new_n246_, new_n272_ );
xor g059 ( N450, new_n273_, keyIn_0_29 );
not g060 ( new_n275_, N130 );
nand g061 ( new_n276_, N101, N106 );
xnor g062 ( new_n277_, new_n276_, keyIn_0_10 );
nor g063 ( new_n278_, N101, N106 );
xor g064 ( new_n279_, new_n278_, keyIn_0_11 );
nor g065 ( new_n280_, new_n279_, new_n277_ );
xnor g066 ( new_n281_, new_n280_, keyIn_0_22 );
xnor g067 ( new_n282_, N91, N96 );
xnor g068 ( new_n283_, new_n282_, keyIn_0_21 );
nor g069 ( new_n284_, new_n281_, new_n283_ );
not g070 ( new_n285_, new_n284_ );
nor g071 ( new_n286_, new_n285_, keyIn_0_30 );
nand g072 ( new_n287_, new_n285_, keyIn_0_30 );
nand g073 ( new_n288_, new_n281_, new_n283_ );
nand g074 ( new_n289_, new_n287_, new_n288_ );
nor g075 ( new_n290_, new_n289_, new_n286_ );
not g076 ( new_n291_, new_n290_ );
nor g077 ( new_n292_, new_n291_, new_n275_ );
not g078 ( new_n293_, new_n292_ );
nand g079 ( new_n294_, new_n293_, keyIn_0_44 );
not g080 ( new_n295_, new_n294_ );
nor g081 ( new_n296_, new_n290_, N130 );
nor g082 ( new_n297_, new_n296_, keyIn_0_45 );
nor g083 ( new_n298_, new_n295_, new_n297_ );
nor g084 ( new_n299_, new_n293_, keyIn_0_44 );
nand g085 ( new_n300_, new_n296_, keyIn_0_45 );
not g086 ( new_n301_, new_n300_ );
nor g087 ( new_n302_, new_n299_, new_n301_ );
nand g088 ( new_n303_, new_n298_, new_n302_ );
nor g089 ( new_n304_, new_n303_, keyIn_0_57 );
nand g090 ( new_n305_, new_n303_, keyIn_0_57 );
not g091 ( new_n306_, N135 );
not g092 ( new_n307_, keyIn_0_12 );
nor g093 ( new_n308_, N121, N126 );
nand g094 ( new_n309_, new_n308_, new_n307_ );
nor g095 ( new_n310_, new_n308_, new_n307_ );
not g096 ( new_n311_, keyIn_0_31 );
nand g097 ( new_n312_, N121, N126 );
nand g098 ( new_n313_, new_n312_, new_n311_ );
nor g099 ( new_n314_, new_n310_, new_n313_ );
nand g100 ( new_n315_, new_n314_, new_n309_ );
xor g101 ( new_n316_, N111, N116 );
xnor g102 ( new_n317_, new_n316_, keyIn_0_23 );
xnor g103 ( new_n318_, new_n317_, new_n315_ );
not g104 ( new_n319_, new_n318_ );
nand g105 ( new_n320_, new_n319_, new_n306_ );
xor g106 ( new_n321_, new_n320_, keyIn_0_46 );
nand g107 ( new_n322_, new_n318_, N135 );
nand g108 ( new_n323_, new_n321_, new_n322_ );
xnor g109 ( new_n324_, new_n323_, keyIn_0_53 );
nand g110 ( new_n325_, new_n305_, new_n324_ );
nor g111 ( new_n326_, new_n325_, new_n304_ );
xnor g112 ( new_n327_, new_n326_, keyIn_0_63 );
not g113 ( new_n328_, new_n303_ );
nor g114 ( new_n329_, new_n328_, new_n324_ );
nor g115 ( N767, new_n327_, new_n329_ );
not g116 ( new_n331_, keyIn_0_64 );
not g117 ( new_n332_, keyIn_0_62 );
not g118 ( new_n333_, N207 );
xnor g119 ( new_n334_, N183, N189 );
xnor g120 ( new_n335_, new_n334_, keyIn_0_25 );
xnor g121 ( new_n336_, N195, N201 );
xnor g122 ( new_n337_, new_n336_, keyIn_0_26 );
xnor g123 ( new_n338_, new_n335_, new_n337_ );
not g124 ( new_n339_, new_n338_ );
nor g125 ( new_n340_, new_n339_, new_n333_ );
not g126 ( new_n341_, new_n340_ );
nor g127 ( new_n342_, new_n341_, keyIn_0_51 );
nand g128 ( new_n343_, new_n341_, keyIn_0_51 );
not g129 ( new_n344_, new_n343_ );
nor g130 ( new_n345_, new_n338_, N207 );
nor g131 ( new_n346_, new_n344_, new_n345_ );
not g132 ( new_n347_, new_n346_ );
nor g133 ( new_n348_, new_n347_, new_n342_ );
nand g134 ( new_n349_, new_n348_, new_n332_ );
nor g135 ( new_n350_, new_n348_, new_n332_ );
xor g136 ( new_n351_, N171, N177 );
nand g137 ( new_n352_, N159, N165 );
xnor g138 ( new_n353_, new_n351_, new_n352_ );
nor g139 ( new_n354_, N159, N165 );
nor g140 ( new_n355_, new_n354_, keyIn_0_15 );
xnor g141 ( new_n356_, new_n353_, new_n355_ );
xnor g142 ( new_n357_, new_n356_, new_n275_ );
xnor g143 ( new_n358_, new_n357_, keyIn_0_61 );
nor g144 ( new_n359_, new_n350_, new_n358_ );
nand g145 ( new_n360_, new_n359_, new_n349_ );
nor g146 ( new_n361_, new_n360_, new_n331_ );
nand g147 ( new_n362_, new_n360_, new_n331_ );
not g148 ( new_n363_, new_n348_ );
nand g149 ( new_n364_, new_n363_, new_n357_ );
nand g150 ( new_n365_, new_n362_, new_n364_ );
nor g151 ( N768, new_n365_, new_n361_ );
not g152 ( new_n367_, N261 );
not g153 ( new_n368_, N201 );
not g154 ( new_n369_, keyIn_0_56 );
not g155 ( new_n370_, keyIn_0_50 );
not g156 ( new_n371_, keyIn_0_36 );
nand g157 ( new_n372_, N17, N51 );
not g158 ( new_n373_, new_n372_ );
nand g159 ( new_n374_, new_n228_, new_n373_ );
nand g160 ( new_n375_, new_n374_, keyIn_0_2 );
not g161 ( new_n376_, keyIn_0_2 );
nor g162 ( new_n377_, new_n227_, new_n372_ );
nand g163 ( new_n378_, new_n377_, new_n376_ );
nand g164 ( new_n379_, new_n375_, new_n378_ );
not g165 ( new_n380_, keyIn_0_7 );
nand g166 ( new_n381_, N42, N59 );
not g167 ( new_n382_, new_n381_ );
nand g168 ( new_n383_, new_n382_, N75 );
nand g169 ( new_n384_, new_n383_, new_n380_ );
nor g170 ( new_n385_, new_n381_, new_n215_ );
nand g171 ( new_n386_, new_n385_, keyIn_0_7 );
nand g172 ( new_n387_, new_n384_, new_n386_ );
nand g173 ( new_n388_, new_n379_, new_n387_ );
nand g174 ( new_n389_, N17, N42 );
not g175 ( new_n390_, new_n389_ );
nand g176 ( new_n391_, new_n226_, new_n221_ );
nand g177 ( new_n392_, N59, N156 );
not g178 ( new_n393_, new_n392_ );
nand g179 ( new_n394_, new_n391_, new_n393_ );
nor g180 ( new_n395_, new_n394_, new_n390_ );
nand g181 ( new_n396_, N447, new_n395_ );
nand g182 ( new_n397_, new_n388_, new_n396_ );
xnor g183 ( new_n398_, new_n397_, new_n371_ );
nand g184 ( new_n399_, new_n398_, N126 );
nand g185 ( new_n400_, new_n399_, new_n370_ );
not g186 ( new_n401_, N126 );
xnor g187 ( new_n402_, new_n397_, keyIn_0_36 );
nor g188 ( new_n403_, new_n402_, new_n401_ );
nand g189 ( new_n404_, new_n403_, keyIn_0_50 );
nand g190 ( new_n405_, new_n404_, new_n400_ );
xnor g191 ( new_n406_, new_n256_, new_n251_ );
xnor g192 ( new_n407_, new_n392_, keyIn_0_14 );
nand g193 ( new_n408_, new_n407_, N17 );
nor g194 ( new_n409_, new_n406_, new_n408_ );
nand g195 ( new_n410_, new_n409_, keyIn_0_35 );
not g196 ( new_n411_, keyIn_0_35 );
not g197 ( new_n412_, keyIn_0_14 );
xnor g198 ( new_n413_, new_n392_, new_n412_ );
nor g199 ( new_n414_, new_n413_, new_n226_ );
nand g200 ( new_n415_, new_n414_, N447 );
nand g201 ( new_n416_, new_n415_, new_n411_ );
nand g202 ( new_n417_, new_n410_, new_n416_ );
nand g203 ( new_n418_, new_n417_, N1 );
nand g204 ( new_n419_, new_n418_, N153 );
nand g205 ( new_n420_, new_n405_, new_n419_ );
nor g206 ( new_n421_, new_n420_, new_n369_ );
nand g207 ( new_n422_, new_n420_, new_n369_ );
nand g208 ( new_n423_, N29, N75 );
nor g209 ( new_n424_, new_n423_, new_n218_ );
not g210 ( new_n425_, new_n424_ );
nor g211 ( new_n426_, new_n406_, new_n425_ );
xor g212 ( new_n427_, keyIn_0_24, N268 );
nor g213 ( new_n428_, new_n427_, new_n259_ );
nand g214 ( new_n429_, new_n426_, new_n428_ );
nand g215 ( new_n430_, new_n422_, new_n429_ );
nor g216 ( new_n431_, new_n430_, new_n421_ );
nand g217 ( new_n432_, new_n431_, new_n368_ );
not g218 ( new_n433_, new_n421_ );
not g219 ( new_n434_, new_n430_ );
nand g220 ( new_n435_, new_n434_, new_n433_ );
nand g221 ( new_n436_, new_n435_, N201 );
nand g222 ( new_n437_, new_n436_, new_n432_ );
xor g223 ( new_n438_, new_n437_, keyIn_0_82 );
nor g224 ( new_n439_, new_n438_, new_n367_ );
nand g225 ( new_n440_, new_n439_, keyIn_0_93 );
not g226 ( new_n441_, keyIn_0_93 );
not g227 ( new_n442_, new_n439_ );
nand g228 ( new_n443_, new_n442_, new_n441_ );
not g229 ( new_n444_, new_n443_ );
nand g230 ( new_n445_, new_n438_, new_n367_ );
nand g231 ( new_n446_, new_n445_, N219 );
nor g232 ( new_n447_, new_n444_, new_n446_ );
nand g233 ( new_n448_, new_n447_, new_n440_ );
not g234 ( new_n449_, new_n438_ );
nand g235 ( new_n450_, new_n449_, N228 );
not g236 ( new_n451_, N237 );
nor g237 ( new_n452_, new_n436_, new_n451_ );
nand g238 ( new_n453_, new_n435_, N246 );
nand g239 ( new_n454_, N42, N72 );
not g240 ( new_n455_, new_n454_ );
nand g241 ( new_n456_, new_n455_, N73 );
nor g242 ( new_n457_, new_n456_, new_n267_ );
nand g243 ( new_n458_, new_n261_, new_n457_ );
xnor g244 ( new_n459_, new_n458_, keyIn_0_33 );
not g245 ( new_n460_, new_n459_ );
nand g246 ( new_n461_, new_n460_, N201 );
not g247 ( new_n462_, keyIn_0_18 );
nand g248 ( new_n463_, N255, N267 );
nor g249 ( new_n464_, new_n463_, new_n462_ );
nand g250 ( new_n465_, new_n463_, new_n462_ );
nand g251 ( new_n466_, N121, N210 );
nand g252 ( new_n467_, new_n465_, new_n466_ );
nor g253 ( new_n468_, new_n467_, new_n464_ );
nand g254 ( new_n469_, new_n461_, new_n468_ );
not g255 ( new_n470_, new_n469_ );
nand g256 ( new_n471_, new_n453_, new_n470_ );
nor g257 ( new_n472_, new_n452_, new_n471_ );
nand g258 ( new_n473_, new_n450_, new_n472_ );
not g259 ( new_n474_, new_n473_ );
nand g260 ( N850, new_n448_, new_n474_ );
not g261 ( new_n476_, N189 );
nand g262 ( new_n477_, new_n418_, N146 );
xnor g263 ( new_n478_, new_n477_, keyIn_0_48 );
nand g264 ( new_n479_, new_n398_, N116 );
nand g265 ( new_n480_, new_n479_, new_n429_ );
not g266 ( new_n481_, new_n480_ );
nand g267 ( new_n482_, new_n478_, new_n481_ );
xnor g268 ( new_n483_, new_n482_, keyIn_0_60 );
nand g269 ( new_n484_, new_n483_, new_n476_ );
nand g270 ( new_n485_, new_n484_, keyIn_0_70 );
not g271 ( new_n486_, keyIn_0_70 );
not g272 ( new_n487_, keyIn_0_60 );
nand g273 ( new_n488_, new_n482_, new_n487_ );
not g274 ( new_n489_, keyIn_0_48 );
xnor g275 ( new_n490_, new_n477_, new_n489_ );
nor g276 ( new_n491_, new_n490_, new_n480_ );
nand g277 ( new_n492_, new_n491_, keyIn_0_60 );
nand g278 ( new_n493_, new_n492_, new_n488_ );
nor g279 ( new_n494_, new_n493_, N189 );
nand g280 ( new_n495_, new_n494_, new_n486_ );
nand g281 ( new_n496_, new_n485_, new_n495_ );
not g282 ( new_n497_, keyIn_0_72 );
nand g283 ( new_n498_, new_n418_, N149 );
xor g284 ( new_n499_, new_n498_, keyIn_0_49 );
xnor g285 ( new_n500_, new_n429_, keyIn_0_43 );
not g286 ( new_n501_, N121 );
nor g287 ( new_n502_, new_n402_, new_n501_ );
nor g288 ( new_n503_, new_n502_, new_n500_ );
nand g289 ( new_n504_, new_n499_, new_n503_ );
nor g290 ( new_n505_, new_n504_, N195 );
xnor g291 ( new_n506_, new_n505_, new_n497_ );
not g292 ( new_n507_, new_n506_ );
nand g293 ( new_n508_, new_n432_, N261 );
not g294 ( new_n509_, new_n508_ );
nand g295 ( new_n510_, new_n509_, new_n507_ );
nand g296 ( new_n511_, new_n504_, N195 );
xnor g297 ( new_n512_, new_n511_, keyIn_0_71 );
xor g298 ( new_n513_, new_n512_, keyIn_0_80 );
nand g299 ( new_n514_, new_n513_, new_n510_ );
nand g300 ( new_n515_, new_n514_, new_n496_ );
not g301 ( new_n516_, keyIn_0_95 );
nor g302 ( new_n517_, new_n436_, new_n506_ );
nand g303 ( new_n518_, new_n517_, new_n496_ );
nor g304 ( new_n519_, new_n518_, new_n516_ );
nand g305 ( new_n520_, new_n518_, new_n516_ );
nor g306 ( new_n521_, new_n483_, new_n476_ );
xnor g307 ( new_n522_, new_n521_, keyIn_0_90 );
nand g308 ( new_n523_, new_n520_, new_n522_ );
nor g309 ( new_n524_, new_n523_, new_n519_ );
nand g310 ( new_n525_, new_n524_, new_n515_ );
not g311 ( new_n526_, N183 );
nand g312 ( new_n527_, new_n418_, N143 );
not g313 ( new_n528_, new_n527_ );
nand g314 ( new_n529_, new_n398_, N111 );
xor g315 ( new_n530_, new_n429_, keyIn_0_42 );
nand g316 ( new_n531_, new_n529_, new_n530_ );
nor g317 ( new_n532_, new_n531_, new_n528_ );
nor g318 ( new_n533_, new_n532_, new_n526_ );
not g319 ( new_n534_, new_n533_ );
nand g320 ( new_n535_, new_n532_, new_n526_ );
nand g321 ( new_n536_, new_n534_, new_n535_ );
xor g322 ( new_n537_, new_n536_, keyIn_0_79 );
xor g323 ( new_n538_, new_n525_, new_n537_ );
nor g324 ( new_n539_, new_n538_, keyIn_0_103 );
nand g325 ( new_n540_, new_n538_, keyIn_0_103 );
nand g326 ( new_n541_, new_n540_, N219 );
nor g327 ( new_n542_, new_n541_, new_n539_ );
xor g328 ( new_n543_, new_n542_, keyIn_0_106 );
not g329 ( new_n544_, keyIn_0_89 );
not g330 ( new_n545_, N228 );
nor g331 ( new_n546_, new_n537_, new_n545_ );
nand g332 ( new_n547_, new_n546_, new_n544_ );
not g333 ( new_n548_, new_n546_ );
nand g334 ( new_n549_, new_n548_, keyIn_0_89 );
xor g335 ( new_n550_, new_n533_, keyIn_0_78 );
nand g336 ( new_n551_, new_n550_, N237 );
nand g337 ( new_n552_, new_n549_, new_n551_ );
not g338 ( new_n553_, new_n552_ );
nand g339 ( new_n554_, new_n553_, new_n547_ );
nor g340 ( new_n555_, new_n554_, keyIn_0_98 );
nand g341 ( new_n556_, new_n554_, keyIn_0_98 );
not g342 ( new_n557_, N246 );
nor g343 ( new_n558_, new_n532_, new_n557_ );
nand g344 ( new_n559_, new_n460_, N183 );
nand g345 ( new_n560_, N106, N210 );
nand g346 ( new_n561_, new_n559_, new_n560_ );
nor g347 ( new_n562_, new_n558_, new_n561_ );
nand g348 ( new_n563_, new_n556_, new_n562_ );
nor g349 ( new_n564_, new_n563_, new_n555_ );
nand g350 ( new_n565_, new_n543_, new_n564_ );
xor g351 ( N863, new_n565_, keyIn_0_120 );
not g352 ( new_n567_, keyIn_0_111 );
xor g353 ( new_n568_, new_n510_, keyIn_0_83 );
xor g354 ( new_n569_, new_n513_, keyIn_0_91 );
xor g355 ( new_n570_, new_n517_, keyIn_0_94 );
nand g356 ( new_n571_, new_n569_, new_n570_ );
nor g357 ( new_n572_, new_n571_, new_n568_ );
xnor g358 ( new_n573_, new_n572_, keyIn_0_99 );
not g359 ( new_n574_, new_n521_ );
nand g360 ( new_n575_, new_n496_, new_n574_ );
nor g361 ( new_n576_, new_n573_, new_n575_ );
nand g362 ( new_n577_, new_n573_, new_n575_ );
nand g363 ( new_n578_, new_n577_, N219 );
nor g364 ( new_n579_, new_n578_, new_n576_ );
nand g365 ( new_n580_, N111, N210 );
not g366 ( new_n581_, new_n580_ );
nor g367 ( new_n582_, new_n579_, new_n581_ );
nand g368 ( new_n583_, new_n582_, new_n567_ );
nor g369 ( new_n584_, new_n582_, new_n567_ );
not g370 ( new_n585_, new_n575_ );
nand g371 ( new_n586_, new_n585_, N228 );
nor g372 ( new_n587_, new_n574_, new_n451_ );
nand g373 ( new_n588_, new_n493_, N246 );
nand g374 ( new_n589_, new_n460_, N189 );
nand g375 ( new_n590_, N255, N259 );
nand g376 ( new_n591_, new_n589_, new_n590_ );
not g377 ( new_n592_, new_n591_ );
nand g378 ( new_n593_, new_n588_, new_n592_ );
nor g379 ( new_n594_, new_n587_, new_n593_ );
nand g380 ( new_n595_, new_n586_, new_n594_ );
nor g381 ( new_n596_, new_n584_, new_n595_ );
nand g382 ( N864, new_n596_, new_n583_ );
not g383 ( new_n598_, N219 );
nand g384 ( new_n599_, new_n507_, new_n512_ );
nand g385 ( new_n600_, new_n508_, new_n436_ );
xnor g386 ( new_n601_, new_n600_, new_n599_ );
xnor g387 ( new_n602_, new_n601_, keyIn_0_104 );
nor g388 ( new_n603_, new_n602_, new_n598_ );
nor g389 ( new_n604_, new_n513_, new_n451_ );
nor g390 ( new_n605_, new_n599_, new_n545_ );
xor g391 ( new_n606_, new_n605_, keyIn_0_92 );
nor g392 ( new_n607_, new_n606_, new_n604_ );
xnor g393 ( new_n608_, new_n607_, keyIn_0_100 );
nand g394 ( new_n609_, new_n504_, N246 );
nand g395 ( new_n610_, N255, N260 );
nand g396 ( new_n611_, new_n609_, new_n610_ );
xor g397 ( new_n612_, new_n611_, keyIn_0_81 );
nand g398 ( new_n613_, new_n460_, N195 );
nand g399 ( new_n614_, N116, N210 );
xnor g400 ( new_n615_, new_n614_, keyIn_0_17 );
nand g401 ( new_n616_, new_n613_, new_n615_ );
nor g402 ( new_n617_, new_n612_, new_n616_ );
nand g403 ( new_n618_, new_n608_, new_n617_ );
nor g404 ( new_n619_, new_n618_, new_n603_ );
xnor g405 ( N865, new_n619_, keyIn_0_117 );
not g406 ( new_n621_, keyIn_0_102 );
nand g407 ( new_n622_, new_n525_, new_n535_ );
xnor g408 ( new_n623_, new_n622_, keyIn_0_101 );
nor g409 ( new_n624_, new_n623_, new_n550_ );
nand g410 ( new_n625_, new_n624_, new_n621_ );
not g411 ( new_n626_, new_n550_ );
not g412 ( new_n627_, keyIn_0_101 );
xnor g413 ( new_n628_, new_n622_, new_n627_ );
nand g414 ( new_n629_, new_n628_, new_n626_ );
nand g415 ( new_n630_, new_n629_, keyIn_0_102 );
nand g416 ( new_n631_, new_n625_, new_n630_ );
not g417 ( new_n632_, N177 );
nor g418 ( new_n633_, new_n413_, new_n259_ );
nand g419 ( new_n634_, new_n633_, N447 );
xnor g420 ( new_n635_, new_n634_, keyIn_0_34 );
not g421 ( new_n636_, new_n635_ );
nand g422 ( new_n637_, new_n636_, N153 );
nor g423 ( new_n638_, new_n226_, N268 );
nand g424 ( new_n639_, new_n426_, new_n638_ );
nand g425 ( new_n640_, new_n637_, new_n639_ );
nor g426 ( new_n641_, new_n640_, keyIn_0_47 );
nand g427 ( new_n642_, new_n640_, keyIn_0_47 );
not g428 ( new_n643_, N106 );
nor g429 ( new_n644_, new_n402_, new_n643_ );
nand g430 ( new_n645_, N138, N152 );
xnor g431 ( new_n646_, new_n645_, keyIn_0_13 );
nor g432 ( new_n647_, new_n644_, new_n646_ );
nand g433 ( new_n648_, new_n642_, new_n647_ );
nor g434 ( new_n649_, new_n648_, new_n641_ );
xor g435 ( new_n650_, new_n649_, keyIn_0_59 );
not g436 ( new_n651_, new_n650_ );
nand g437 ( new_n652_, new_n651_, new_n632_ );
xnor g438 ( new_n653_, new_n652_, keyIn_0_69 );
not g439 ( new_n654_, new_n653_ );
nand g440 ( new_n655_, new_n631_, new_n654_ );
nand g441 ( new_n656_, new_n398_, N101 );
nand g442 ( new_n657_, N17, N138 );
nand g443 ( new_n658_, new_n656_, new_n657_ );
xor g444 ( new_n659_, new_n658_, keyIn_0_55 );
nand g445 ( new_n660_, new_n636_, N149 );
nor g446 ( new_n661_, new_n660_, keyIn_0_41 );
nand g447 ( new_n662_, new_n660_, keyIn_0_41 );
nand g448 ( new_n663_, new_n662_, new_n639_ );
nor g449 ( new_n664_, new_n663_, new_n661_ );
nand g450 ( new_n665_, new_n659_, new_n664_ );
nor g451 ( new_n666_, new_n665_, N171 );
xnor g452 ( new_n667_, new_n666_, keyIn_0_68 );
nor g453 ( new_n668_, new_n655_, new_n667_ );
not g454 ( new_n669_, N165 );
nand g455 ( new_n670_, new_n636_, N146 );
nor g456 ( new_n671_, new_n670_, keyIn_0_39 );
xor g457 ( new_n672_, new_n639_, keyIn_0_40 );
nand g458 ( new_n673_, N51, N138 );
not g459 ( new_n674_, new_n673_ );
nor g460 ( new_n675_, new_n672_, new_n674_ );
not g461 ( new_n676_, new_n675_ );
nor g462 ( new_n677_, new_n676_, new_n671_ );
not g463 ( new_n678_, new_n677_ );
nand g464 ( new_n679_, new_n398_, N96 );
nand g465 ( new_n680_, new_n670_, keyIn_0_39 );
nand g466 ( new_n681_, new_n680_, new_n679_ );
nor g467 ( new_n682_, new_n678_, new_n681_ );
nand g468 ( new_n683_, new_n682_, new_n669_ );
xnor g469 ( new_n684_, new_n683_, keyIn_0_66 );
not g470 ( new_n685_, new_n684_ );
nand g471 ( new_n686_, new_n668_, new_n685_ );
not g472 ( new_n687_, new_n667_ );
nor g473 ( new_n688_, new_n651_, new_n632_ );
nand g474 ( new_n689_, new_n687_, new_n688_ );
nand g475 ( new_n690_, new_n665_, N171 );
xnor g476 ( new_n691_, new_n690_, keyIn_0_67 );
nand g477 ( new_n692_, new_n689_, new_n691_ );
nand g478 ( new_n693_, new_n692_, new_n685_ );
nor g479 ( new_n694_, new_n682_, new_n669_ );
not g480 ( new_n695_, new_n694_ );
nand g481 ( new_n696_, new_n693_, new_n695_ );
not g482 ( new_n697_, new_n696_ );
nand g483 ( new_n698_, new_n686_, new_n697_ );
not g484 ( new_n699_, N159 );
nand g485 ( new_n700_, new_n398_, N91 );
nand g486 ( new_n701_, N8, N138 );
nand g487 ( new_n702_, new_n700_, new_n701_ );
xor g488 ( new_n703_, new_n702_, keyIn_0_54 );
not g489 ( new_n704_, keyIn_0_37 );
nand g490 ( new_n705_, new_n636_, N143 );
nor g491 ( new_n706_, new_n705_, new_n704_ );
nand g492 ( new_n707_, new_n705_, new_n704_ );
xnor g493 ( new_n708_, new_n639_, keyIn_0_38 );
nand g494 ( new_n709_, new_n707_, new_n708_ );
nor g495 ( new_n710_, new_n709_, new_n706_ );
nand g496 ( new_n711_, new_n703_, new_n710_ );
xor g497 ( new_n712_, new_n711_, keyIn_0_58 );
not g498 ( new_n713_, new_n712_ );
nand g499 ( new_n714_, new_n713_, new_n699_ );
xnor g500 ( new_n715_, new_n714_, keyIn_0_65 );
nand g501 ( new_n716_, new_n698_, new_n715_ );
xnor g502 ( new_n717_, new_n716_, keyIn_0_114 );
nand g503 ( new_n718_, new_n712_, N159 );
xnor g504 ( new_n719_, new_n718_, keyIn_0_73 );
nand g505 ( new_n720_, new_n717_, new_n719_ );
xnor g506 ( N866, new_n720_, keyIn_0_118 );
nor g507 ( new_n722_, new_n653_, new_n688_ );
nor g508 ( new_n723_, new_n631_, new_n722_ );
nand g509 ( new_n724_, new_n723_, keyIn_0_105 );
nor g510 ( new_n725_, new_n723_, keyIn_0_105 );
not g511 ( new_n726_, new_n631_ );
not g512 ( new_n727_, new_n722_ );
nor g513 ( new_n728_, new_n726_, new_n727_ );
nor g514 ( new_n729_, new_n725_, new_n728_ );
nand g515 ( new_n730_, new_n729_, new_n724_ );
xnor g516 ( new_n731_, new_n730_, keyIn_0_110 );
nand g517 ( new_n732_, new_n731_, N219 );
nor g518 ( new_n733_, new_n727_, new_n545_ );
nand g519 ( new_n734_, new_n688_, N237 );
nor g520 ( new_n735_, new_n651_, new_n557_ );
nand g521 ( new_n736_, new_n460_, N177 );
xnor g522 ( new_n737_, new_n736_, keyIn_0_52 );
nand g523 ( new_n738_, N101, N210 );
nand g524 ( new_n739_, new_n737_, new_n738_ );
nor g525 ( new_n740_, new_n735_, new_n739_ );
nand g526 ( new_n741_, new_n740_, new_n734_ );
nor g527 ( new_n742_, new_n733_, new_n741_ );
nand g528 ( new_n743_, new_n732_, new_n742_ );
xnor g529 ( N874, new_n743_, keyIn_0_123 );
not g530 ( new_n745_, keyIn_0_124 );
not g531 ( new_n746_, keyIn_0_115 );
not g532 ( new_n747_, keyIn_0_112 );
nand g533 ( new_n748_, new_n715_, new_n718_ );
xnor g534 ( new_n749_, new_n748_, keyIn_0_74 );
nor g535 ( new_n750_, new_n698_, new_n749_ );
nand g536 ( new_n751_, new_n750_, new_n747_ );
not g537 ( new_n752_, new_n751_ );
not g538 ( new_n753_, new_n698_ );
not g539 ( new_n754_, new_n749_ );
nand g540 ( new_n755_, new_n753_, new_n754_ );
nand g541 ( new_n756_, new_n755_, keyIn_0_112 );
nand g542 ( new_n757_, new_n698_, new_n749_ );
nand g543 ( new_n758_, new_n756_, new_n757_ );
nor g544 ( new_n759_, new_n758_, new_n752_ );
nand g545 ( new_n760_, new_n759_, new_n746_ );
nor g546 ( new_n761_, new_n750_, new_n747_ );
not g547 ( new_n762_, new_n757_ );
nor g548 ( new_n763_, new_n761_, new_n762_ );
nand g549 ( new_n764_, new_n763_, new_n751_ );
nand g550 ( new_n765_, new_n764_, keyIn_0_115 );
nand g551 ( new_n766_, new_n760_, new_n765_ );
nand g552 ( new_n767_, new_n766_, N219 );
nand g553 ( new_n768_, new_n427_, N210 );
xor g554 ( new_n769_, new_n768_, keyIn_0_32 );
nand g555 ( new_n770_, new_n767_, new_n769_ );
xnor g556 ( new_n771_, new_n770_, keyIn_0_121 );
nor g557 ( new_n772_, new_n754_, new_n545_ );
nor g558 ( new_n773_, new_n719_, new_n451_ );
not g559 ( new_n774_, new_n773_ );
nor g560 ( new_n775_, new_n774_, keyIn_0_84 );
nand g561 ( new_n776_, new_n774_, keyIn_0_84 );
nor g562 ( new_n777_, new_n713_, new_n557_ );
nor g563 ( new_n778_, new_n459_, new_n699_ );
nor g564 ( new_n779_, new_n777_, new_n778_ );
nand g565 ( new_n780_, new_n776_, new_n779_ );
nor g566 ( new_n781_, new_n780_, new_n775_ );
not g567 ( new_n782_, new_n781_ );
nor g568 ( new_n783_, new_n772_, new_n782_ );
nand g569 ( new_n784_, new_n771_, new_n783_ );
xnor g570 ( new_n785_, new_n784_, new_n745_ );
nand g571 ( new_n786_, new_n785_, keyIn_0_125 );
not g572 ( new_n787_, keyIn_0_125 );
nand g573 ( new_n788_, new_n784_, keyIn_0_124 );
not g574 ( new_n789_, keyIn_0_121 );
xnor g575 ( new_n790_, new_n770_, new_n789_ );
not g576 ( new_n791_, new_n783_ );
nor g577 ( new_n792_, new_n790_, new_n791_ );
nand g578 ( new_n793_, new_n792_, new_n745_ );
nand g579 ( new_n794_, new_n793_, new_n788_ );
nand g580 ( new_n795_, new_n794_, new_n787_ );
nand g581 ( N878, new_n786_, new_n795_ );
not g582 ( new_n797_, keyIn_0_119 );
not g583 ( new_n798_, keyIn_0_107 );
nand g584 ( new_n799_, new_n668_, new_n798_ );
nor g585 ( new_n800_, new_n668_, new_n798_ );
xnor g586 ( new_n801_, new_n689_, keyIn_0_96 );
xor g587 ( new_n802_, new_n691_, keyIn_0_86 );
nand g588 ( new_n803_, new_n801_, new_n802_ );
nor g589 ( new_n804_, new_n800_, new_n803_ );
nand g590 ( new_n805_, new_n804_, new_n799_ );
xnor g591 ( new_n806_, new_n805_, keyIn_0_108 );
nor g592 ( new_n807_, new_n684_, new_n694_ );
nor g593 ( new_n808_, new_n806_, new_n807_ );
nand g594 ( new_n809_, new_n806_, new_n807_ );
nand g595 ( new_n810_, new_n809_, N219 );
nor g596 ( new_n811_, new_n810_, new_n808_ );
nand g597 ( new_n812_, new_n811_, new_n797_ );
nor g598 ( new_n813_, new_n811_, new_n797_ );
not g599 ( new_n814_, keyIn_0_85 );
not g600 ( new_n815_, new_n807_ );
nor g601 ( new_n816_, new_n815_, new_n545_ );
nand g602 ( new_n817_, new_n816_, new_n814_ );
nor g603 ( new_n818_, new_n816_, new_n814_ );
nor g604 ( new_n819_, new_n682_, new_n557_ );
nor g605 ( new_n820_, new_n459_, new_n669_ );
nor g606 ( new_n821_, new_n819_, new_n820_ );
xor g607 ( new_n822_, new_n821_, keyIn_0_75 );
nor g608 ( new_n823_, new_n695_, new_n451_ );
nand g609 ( new_n824_, N91, N210 );
xnor g610 ( new_n825_, new_n824_, keyIn_0_16 );
nor g611 ( new_n826_, new_n823_, new_n825_ );
nand g612 ( new_n827_, new_n822_, new_n826_ );
nor g613 ( new_n828_, new_n818_, new_n827_ );
nand g614 ( new_n829_, new_n828_, new_n817_ );
nor g615 ( new_n830_, new_n813_, new_n829_ );
nand g616 ( new_n831_, new_n830_, new_n812_ );
xor g617 ( N879, new_n831_, keyIn_0_126 );
not g618 ( new_n833_, keyIn_0_122 );
xor g619 ( new_n834_, new_n688_, keyIn_0_88 );
nand g620 ( new_n835_, new_n655_, new_n834_ );
xnor g621 ( new_n836_, new_n835_, keyIn_0_109 );
nand g622 ( new_n837_, new_n687_, new_n691_ );
xnor g623 ( new_n838_, new_n837_, keyIn_0_76 );
nor g624 ( new_n839_, new_n836_, new_n838_ );
xnor g625 ( new_n840_, new_n839_, keyIn_0_113 );
nand g626 ( new_n841_, new_n836_, new_n838_ );
nand g627 ( new_n842_, new_n840_, new_n841_ );
xnor g628 ( new_n843_, new_n842_, keyIn_0_116 );
nand g629 ( new_n844_, new_n843_, N219 );
nand g630 ( new_n845_, N96, N210 );
nand g631 ( new_n846_, new_n844_, new_n845_ );
nor g632 ( new_n847_, new_n846_, new_n833_ );
nand g633 ( new_n848_, new_n846_, new_n833_ );
nand g634 ( new_n849_, new_n838_, N228 );
xor g635 ( new_n850_, new_n849_, keyIn_0_87 );
nor g636 ( new_n851_, new_n691_, new_n451_ );
nor g637 ( new_n852_, new_n850_, new_n851_ );
xor g638 ( new_n853_, new_n852_, keyIn_0_97 );
nand g639 ( new_n854_, new_n665_, N246 );
nand g640 ( new_n855_, new_n460_, N171 );
nand g641 ( new_n856_, new_n854_, new_n855_ );
xor g642 ( new_n857_, new_n856_, keyIn_0_77 );
nor g643 ( new_n858_, new_n853_, new_n857_ );
nand g644 ( new_n859_, new_n848_, new_n858_ );
nor g645 ( new_n860_, new_n859_, new_n847_ );
xnor g646 ( N880, new_n860_, keyIn_0_127 );
endmodule