module add_mul_sub_8_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, operation_0_, 
        operation_1_, Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, 
        Result_5_, Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, 
        Result_11_, Result_12_, Result_13_, Result_14_, Result_15_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_,
         b_4_, b_5_, b_6_, b_7_, operation_0_, operation_1_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_;
  wire   n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186;

  OR3_X1 U587 ( .A1(n571), .A2(n572), .A3(n573), .ZN(Result_9_) );
  AND2_X1 U588 ( .A1(n574), .A2(n575), .ZN(n573) );
  XNOR2_X1 U589 ( .A(n576), .B(n577), .ZN(n575) );
  XOR2_X1 U590 ( .A(n578), .B(n579), .Z(n577) );
  AND2_X1 U591 ( .A1(n580), .A2(n581), .ZN(n572) );
  OR3_X1 U592 ( .A1(n582), .A2(n583), .A3(n584), .ZN(n581) );
  AND2_X1 U593 ( .A1(n585), .A2(n586), .ZN(n584) );
  INV_X1 U594 ( .A(n587), .ZN(n586) );
  AND2_X1 U595 ( .A1(n588), .A2(n589), .ZN(n583) );
  INV_X1 U596 ( .A(n590), .ZN(n589) );
  AND2_X1 U597 ( .A1(n591), .A2(n592), .ZN(n582) );
  AND2_X1 U598 ( .A1(n593), .A2(n594), .ZN(n571) );
  INV_X1 U599 ( .A(n580), .ZN(n594) );
  AND2_X1 U600 ( .A1(n595), .A2(n596), .ZN(n580) );
  OR2_X1 U601 ( .A1(a_1_), .A2(b_1_), .ZN(n595) );
  OR3_X1 U602 ( .A1(n597), .A2(n598), .A3(n599), .ZN(n593) );
  AND2_X1 U603 ( .A1(n585), .A2(n587), .ZN(n599) );
  AND2_X1 U604 ( .A1(n588), .A2(n590), .ZN(n598) );
  AND2_X1 U605 ( .A1(n600), .A2(n591), .ZN(n597) );
  INV_X1 U606 ( .A(n592), .ZN(n600) );
  OR3_X1 U607 ( .A1(n601), .A2(n602), .A3(n603), .ZN(Result_8_) );
  AND2_X1 U608 ( .A1(n574), .A2(n604), .ZN(n603) );
  XNOR2_X1 U609 ( .A(n605), .B(n606), .ZN(n604) );
  XOR2_X1 U610 ( .A(n607), .B(n608), .Z(n606) );
  AND2_X1 U611 ( .A1(n609), .A2(n610), .ZN(n602) );
  INV_X1 U612 ( .A(n611), .ZN(n610) );
  OR3_X1 U613 ( .A1(n612), .A2(n613), .A3(n614), .ZN(n609) );
  AND2_X1 U614 ( .A1(n615), .A2(n585), .ZN(n614) );
  INV_X1 U615 ( .A(n616), .ZN(n615) );
  AND2_X1 U616 ( .A1(n617), .A2(n588), .ZN(n613) );
  INV_X1 U617 ( .A(n618), .ZN(n617) );
  AND2_X1 U618 ( .A1(n591), .A2(n619), .ZN(n612) );
  AND2_X1 U619 ( .A1(n611), .A2(n620), .ZN(n601) );
  OR3_X1 U620 ( .A1(n621), .A2(n622), .A3(n623), .ZN(n620) );
  AND2_X1 U621 ( .A1(n585), .A2(n616), .ZN(n623) );
  AND2_X1 U622 ( .A1(n588), .A2(n618), .ZN(n622) );
  AND2_X1 U623 ( .A1(n624), .A2(n591), .ZN(n621) );
  INV_X1 U624 ( .A(n619), .ZN(n624) );
  OR2_X1 U625 ( .A1(n625), .A2(n626), .ZN(n619) );
  AND2_X1 U626 ( .A1(n627), .A2(n628), .ZN(n626) );
  AND2_X1 U627 ( .A1(n592), .A2(n596), .ZN(n625) );
  OR2_X1 U628 ( .A1(n629), .A2(n630), .ZN(n592) );
  AND2_X1 U629 ( .A1(n631), .A2(n632), .ZN(n629) );
  AND2_X1 U630 ( .A1(n633), .A2(n634), .ZN(n611) );
  OR2_X1 U631 ( .A1(n635), .A2(n636), .ZN(Result_7_) );
  AND2_X1 U632 ( .A1(n574), .A2(n637), .ZN(n635) );
  XOR2_X1 U633 ( .A(n638), .B(n639), .Z(n637) );
  OR2_X1 U634 ( .A1(n640), .A2(n636), .ZN(Result_6_) );
  AND3_X1 U635 ( .A1(n641), .A2(n642), .A3(n574), .ZN(n640) );
  OR2_X1 U636 ( .A1(n643), .A2(n644), .ZN(n641) );
  XOR2_X1 U637 ( .A(n645), .B(n646), .Z(n644) );
  INV_X1 U638 ( .A(n647), .ZN(n643) );
  OR2_X1 U639 ( .A1(n638), .A2(n639), .ZN(n647) );
  OR2_X1 U640 ( .A1(n648), .A2(n636), .ZN(Result_5_) );
  AND2_X1 U641 ( .A1(n574), .A2(n649), .ZN(n648) );
  XOR2_X1 U642 ( .A(n650), .B(n651), .Z(n649) );
  OR2_X1 U643 ( .A1(n652), .A2(n636), .ZN(Result_4_) );
  AND2_X1 U644 ( .A1(n574), .A2(n653), .ZN(n652) );
  XNOR2_X1 U645 ( .A(n654), .B(n655), .ZN(n653) );
  OR2_X1 U646 ( .A1(n656), .A2(n636), .ZN(Result_3_) );
  AND2_X1 U647 ( .A1(n574), .A2(n657), .ZN(n656) );
  XOR2_X1 U648 ( .A(n658), .B(n659), .Z(n657) );
  AND2_X1 U649 ( .A1(n660), .A2(n661), .ZN(n659) );
  OR2_X1 U650 ( .A1(n662), .A2(n663), .ZN(n661) );
  AND2_X1 U651 ( .A1(n664), .A2(n665), .ZN(n663) );
  INV_X1 U652 ( .A(n666), .ZN(n660) );
  OR2_X1 U653 ( .A1(n667), .A2(n636), .ZN(Result_2_) );
  AND2_X1 U654 ( .A1(n668), .A2(n574), .ZN(n667) );
  XOR2_X1 U655 ( .A(n669), .B(n670), .Z(n668) );
  OR2_X1 U656 ( .A1(n671), .A2(n636), .ZN(Result_1_) );
  AND2_X1 U657 ( .A1(n574), .A2(n672), .ZN(n671) );
  XOR2_X1 U658 ( .A(n673), .B(n674), .Z(n672) );
  AND2_X1 U659 ( .A1(n675), .A2(n676), .ZN(n674) );
  OR2_X1 U660 ( .A1(n677), .A2(n678), .ZN(n676) );
  AND2_X1 U661 ( .A1(n679), .A2(n680), .ZN(n677) );
  INV_X1 U662 ( .A(n681), .ZN(n675) );
  OR2_X1 U663 ( .A1(n682), .A2(n683), .ZN(Result_15_) );
  AND2_X1 U664 ( .A1(n574), .A2(n684), .ZN(n683) );
  AND2_X1 U665 ( .A1(n685), .A2(n686), .ZN(n682) );
  OR3_X1 U666 ( .A1(n585), .A2(n588), .A3(n591), .ZN(n686) );
  OR2_X1 U667 ( .A1(n687), .A2(n688), .ZN(n685) );
  OR3_X1 U668 ( .A1(n689), .A2(n690), .A3(n691), .ZN(Result_14_) );
  AND2_X1 U669 ( .A1(n574), .A2(n692), .ZN(n691) );
  OR4_X1 U670 ( .A1(n693), .A2(n694), .A3(n695), .A4(n696), .ZN(n692) );
  AND2_X1 U671 ( .A1(n687), .A2(b_6_), .ZN(n696) );
  AND2_X1 U672 ( .A1(n697), .A2(a_7_), .ZN(n695) );
  AND2_X1 U673 ( .A1(n688), .A2(a_6_), .ZN(n694) );
  AND2_X1 U674 ( .A1(n698), .A2(b_7_), .ZN(n693) );
  AND2_X1 U675 ( .A1(n699), .A2(n700), .ZN(n690) );
  OR3_X1 U676 ( .A1(n701), .A2(n702), .A3(n703), .ZN(n700) );
  AND2_X1 U677 ( .A1(n585), .A2(n688), .ZN(n703) );
  AND2_X1 U678 ( .A1(n588), .A2(n687), .ZN(n702) );
  AND2_X1 U679 ( .A1(n591), .A2(n684), .ZN(n701) );
  INV_X1 U680 ( .A(n704), .ZN(n699) );
  AND2_X1 U681 ( .A1(n705), .A2(n704), .ZN(n689) );
  OR2_X1 U682 ( .A1(n697), .A2(n698), .ZN(n704) );
  OR3_X1 U683 ( .A1(n706), .A2(n707), .A3(n708), .ZN(n705) );
  AND2_X1 U684 ( .A1(n585), .A2(n709), .ZN(n708) );
  INV_X1 U685 ( .A(n688), .ZN(n709) );
  AND2_X1 U686 ( .A1(n588), .A2(n710), .ZN(n707) );
  AND2_X1 U687 ( .A1(n591), .A2(n711), .ZN(n706) );
  OR3_X1 U688 ( .A1(n712), .A2(n713), .A3(n714), .ZN(Result_13_) );
  AND2_X1 U689 ( .A1(n574), .A2(n715), .ZN(n714) );
  XNOR2_X1 U690 ( .A(n716), .B(n717), .ZN(n715) );
  XOR2_X1 U691 ( .A(n718), .B(n719), .Z(n717) );
  AND2_X1 U692 ( .A1(n720), .A2(n721), .ZN(n713) );
  OR3_X1 U693 ( .A1(n722), .A2(n723), .A3(n724), .ZN(n721) );
  AND2_X1 U694 ( .A1(n585), .A2(n725), .ZN(n724) );
  AND2_X1 U695 ( .A1(n588), .A2(n726), .ZN(n723) );
  AND2_X1 U696 ( .A1(n591), .A2(n727), .ZN(n722) );
  INV_X1 U697 ( .A(n728), .ZN(n720) );
  AND2_X1 U698 ( .A1(n728), .A2(n729), .ZN(n712) );
  OR3_X1 U699 ( .A1(n730), .A2(n731), .A3(n732), .ZN(n729) );
  AND2_X1 U700 ( .A1(n585), .A2(n733), .ZN(n732) );
  INV_X1 U701 ( .A(n725), .ZN(n733) );
  AND2_X1 U702 ( .A1(n588), .A2(n734), .ZN(n731) );
  AND2_X1 U703 ( .A1(n591), .A2(n735), .ZN(n730) );
  XNOR2_X1 U704 ( .A(b_5_), .B(n736), .ZN(n728) );
  OR3_X1 U705 ( .A1(n737), .A2(n738), .A3(n739), .ZN(Result_12_) );
  AND2_X1 U706 ( .A1(n574), .A2(n740), .ZN(n739) );
  XNOR2_X1 U707 ( .A(n741), .B(n742), .ZN(n740) );
  XOR2_X1 U708 ( .A(n743), .B(n744), .Z(n742) );
  AND2_X1 U709 ( .A1(n745), .A2(n746), .ZN(n738) );
  OR3_X1 U710 ( .A1(n747), .A2(n748), .A3(n749), .ZN(n746) );
  AND2_X1 U711 ( .A1(n585), .A2(n750), .ZN(n749) );
  AND2_X1 U712 ( .A1(n588), .A2(n751), .ZN(n748) );
  AND2_X1 U713 ( .A1(n752), .A2(n591), .ZN(n747) );
  INV_X1 U714 ( .A(n753), .ZN(n752) );
  INV_X1 U715 ( .A(n754), .ZN(n745) );
  AND2_X1 U716 ( .A1(n754), .A2(n755), .ZN(n737) );
  OR3_X1 U717 ( .A1(n756), .A2(n757), .A3(n758), .ZN(n755) );
  AND2_X1 U718 ( .A1(n585), .A2(n759), .ZN(n758) );
  INV_X1 U719 ( .A(n750), .ZN(n759) );
  AND2_X1 U720 ( .A1(n588), .A2(n760), .ZN(n757) );
  INV_X1 U721 ( .A(n751), .ZN(n760) );
  AND2_X1 U722 ( .A1(n591), .A2(n753), .ZN(n756) );
  XNOR2_X1 U723 ( .A(b_4_), .B(n761), .ZN(n754) );
  OR3_X1 U724 ( .A1(n762), .A2(n763), .A3(n764), .ZN(Result_11_) );
  AND2_X1 U725 ( .A1(n574), .A2(n765), .ZN(n764) );
  XNOR2_X1 U726 ( .A(n766), .B(n767), .ZN(n765) );
  XOR2_X1 U727 ( .A(n768), .B(n769), .Z(n767) );
  AND2_X1 U728 ( .A1(n770), .A2(n771), .ZN(n763) );
  OR3_X1 U729 ( .A1(n772), .A2(n773), .A3(n774), .ZN(n771) );
  AND2_X1 U730 ( .A1(n585), .A2(n775), .ZN(n774) );
  INV_X1 U731 ( .A(n776), .ZN(n775) );
  AND2_X1 U732 ( .A1(n588), .A2(n777), .ZN(n773) );
  INV_X1 U733 ( .A(n778), .ZN(n777) );
  AND2_X1 U734 ( .A1(n591), .A2(n779), .ZN(n772) );
  INV_X1 U735 ( .A(n780), .ZN(n770) );
  AND2_X1 U736 ( .A1(n781), .A2(n780), .ZN(n762) );
  OR2_X1 U737 ( .A1(n782), .A2(n783), .ZN(n780) );
  OR3_X1 U738 ( .A1(n784), .A2(n785), .A3(n786), .ZN(n781) );
  AND2_X1 U739 ( .A1(n585), .A2(n776), .ZN(n786) );
  AND2_X1 U740 ( .A1(n588), .A2(n778), .ZN(n785) );
  AND2_X1 U741 ( .A1(n787), .A2(n591), .ZN(n784) );
  INV_X1 U742 ( .A(n779), .ZN(n787) );
  OR3_X1 U743 ( .A1(n788), .A2(n789), .A3(n790), .ZN(Result_10_) );
  AND2_X1 U744 ( .A1(n574), .A2(n791), .ZN(n790) );
  XNOR2_X1 U745 ( .A(n792), .B(n793), .ZN(n791) );
  XOR2_X1 U746 ( .A(n794), .B(n795), .Z(n793) );
  AND2_X1 U747 ( .A1(n796), .A2(n797), .ZN(n789) );
  OR3_X1 U748 ( .A1(n798), .A2(n799), .A3(n800), .ZN(n797) );
  AND2_X1 U749 ( .A1(n585), .A2(n801), .ZN(n800) );
  INV_X1 U750 ( .A(n802), .ZN(n801) );
  AND2_X1 U751 ( .A1(n588), .A2(n803), .ZN(n799) );
  INV_X1 U752 ( .A(n804), .ZN(n803) );
  AND2_X1 U753 ( .A1(n591), .A2(n631), .ZN(n798) );
  INV_X1 U754 ( .A(n805), .ZN(n796) );
  AND2_X1 U755 ( .A1(n806), .A2(n805), .ZN(n788) );
  OR2_X1 U756 ( .A1(n630), .A2(n807), .ZN(n805) );
  AND2_X1 U757 ( .A1(n808), .A2(n809), .ZN(n630) );
  OR3_X1 U758 ( .A1(n810), .A2(n811), .A3(n812), .ZN(n806) );
  AND2_X1 U759 ( .A1(n585), .A2(n802), .ZN(n812) );
  AND2_X1 U760 ( .A1(n588), .A2(n804), .ZN(n811) );
  AND2_X1 U761 ( .A1(n813), .A2(n591), .ZN(n810) );
  AND2_X1 U762 ( .A1(n814), .A2(n815), .ZN(n591) );
  INV_X1 U763 ( .A(n631), .ZN(n813) );
  OR2_X1 U764 ( .A1(n816), .A2(n782), .ZN(n631) );
  AND2_X1 U765 ( .A1(n817), .A2(n818), .ZN(n782) );
  AND2_X1 U766 ( .A1(n779), .A2(n819), .ZN(n816) );
  OR2_X1 U767 ( .A1(n820), .A2(n821), .ZN(n779) );
  AND2_X1 U768 ( .A1(n761), .A2(n822), .ZN(n821) );
  AND2_X1 U769 ( .A1(n753), .A2(n823), .ZN(n820) );
  OR2_X1 U770 ( .A1(n824), .A2(n825), .ZN(n753) );
  AND2_X1 U771 ( .A1(n736), .A2(n826), .ZN(n825) );
  AND2_X1 U772 ( .A1(n735), .A2(n827), .ZN(n824) );
  INV_X1 U773 ( .A(n727), .ZN(n735) );
  OR2_X1 U774 ( .A1(n828), .A2(n829), .ZN(n727) );
  AND2_X1 U775 ( .A1(n684), .A2(n830), .ZN(n828) );
  OR2_X1 U776 ( .A1(a_6_), .A2(b_6_), .ZN(n830) );
  OR2_X1 U777 ( .A1(n831), .A2(n636), .ZN(Result_0_) );
  OR2_X1 U778 ( .A1(n832), .A2(n833), .ZN(n636) );
  AND2_X1 U779 ( .A1(n585), .A2(n834), .ZN(n833) );
  OR2_X1 U780 ( .A1(n835), .A2(n836), .ZN(n834) );
  AND2_X1 U781 ( .A1(n616), .A2(n633), .ZN(n835) );
  INV_X1 U782 ( .A(n837), .ZN(n633) );
  OR2_X1 U783 ( .A1(n838), .A2(n839), .ZN(n616) );
  AND2_X1 U784 ( .A1(n587), .A2(n627), .ZN(n839) );
  AND2_X1 U785 ( .A1(b_1_), .A2(n840), .ZN(n838) );
  OR2_X1 U786 ( .A1(n627), .A2(n587), .ZN(n840) );
  OR2_X1 U787 ( .A1(n841), .A2(n842), .ZN(n587) );
  AND2_X1 U788 ( .A1(n802), .A2(n808), .ZN(n842) );
  AND2_X1 U789 ( .A1(b_2_), .A2(n843), .ZN(n841) );
  OR2_X1 U790 ( .A1(n808), .A2(n802), .ZN(n843) );
  OR2_X1 U791 ( .A1(n844), .A2(n845), .ZN(n802) );
  AND2_X1 U792 ( .A1(n776), .A2(n817), .ZN(n845) );
  AND2_X1 U793 ( .A1(b_3_), .A2(n846), .ZN(n844) );
  OR2_X1 U794 ( .A1(n817), .A2(n776), .ZN(n846) );
  OR2_X1 U795 ( .A1(n847), .A2(n848), .ZN(n776) );
  AND2_X1 U796 ( .A1(n750), .A2(n761), .ZN(n848) );
  AND2_X1 U797 ( .A1(b_4_), .A2(n849), .ZN(n847) );
  OR2_X1 U798 ( .A1(n761), .A2(n750), .ZN(n849) );
  OR2_X1 U799 ( .A1(n850), .A2(n851), .ZN(n750) );
  AND2_X1 U800 ( .A1(n725), .A2(n736), .ZN(n851) );
  AND2_X1 U801 ( .A1(b_5_), .A2(n852), .ZN(n850) );
  OR2_X1 U802 ( .A1(n736), .A2(n725), .ZN(n852) );
  OR2_X1 U803 ( .A1(n853), .A2(n697), .ZN(n725) );
  AND2_X1 U804 ( .A1(n688), .A2(n854), .ZN(n853) );
  AND2_X1 U805 ( .A1(n855), .A2(b_7_), .ZN(n688) );
  AND2_X1 U806 ( .A1(n815), .A2(operation_1_), .ZN(n585) );
  INV_X1 U807 ( .A(operation_0_), .ZN(n815) );
  AND3_X1 U808 ( .A1(n856), .A2(n634), .A3(n588), .ZN(n832) );
  AND2_X1 U809 ( .A1(n814), .A2(operation_0_), .ZN(n588) );
  INV_X1 U810 ( .A(operation_1_), .ZN(n814) );
  INV_X1 U811 ( .A(n836), .ZN(n634) );
  AND2_X1 U812 ( .A1(n857), .A2(b_0_), .ZN(n836) );
  OR2_X1 U813 ( .A1(n837), .A2(n618), .ZN(n856) );
  OR2_X1 U814 ( .A1(n858), .A2(n859), .ZN(n618) );
  AND2_X1 U815 ( .A1(a_1_), .A2(n590), .ZN(n859) );
  AND2_X1 U816 ( .A1(n860), .A2(n628), .ZN(n858) );
  OR2_X1 U817 ( .A1(a_1_), .A2(n590), .ZN(n860) );
  OR2_X1 U818 ( .A1(n861), .A2(n862), .ZN(n590) );
  AND2_X1 U819 ( .A1(a_2_), .A2(n804), .ZN(n862) );
  AND2_X1 U820 ( .A1(n863), .A2(n809), .ZN(n861) );
  OR2_X1 U821 ( .A1(a_2_), .A2(n804), .ZN(n863) );
  OR2_X1 U822 ( .A1(n864), .A2(n865), .ZN(n804) );
  AND2_X1 U823 ( .A1(a_3_), .A2(n778), .ZN(n865) );
  AND2_X1 U824 ( .A1(n866), .A2(n818), .ZN(n864) );
  OR2_X1 U825 ( .A1(a_3_), .A2(n778), .ZN(n866) );
  OR2_X1 U826 ( .A1(n867), .A2(n868), .ZN(n778) );
  AND2_X1 U827 ( .A1(a_4_), .A2(n751), .ZN(n868) );
  AND2_X1 U828 ( .A1(n869), .A2(n822), .ZN(n867) );
  OR2_X1 U829 ( .A1(a_4_), .A2(n751), .ZN(n869) );
  OR2_X1 U830 ( .A1(n870), .A2(n871), .ZN(n751) );
  AND2_X1 U831 ( .A1(a_5_), .A2(n726), .ZN(n871) );
  AND2_X1 U832 ( .A1(n872), .A2(n826), .ZN(n870) );
  OR2_X1 U833 ( .A1(a_5_), .A2(n726), .ZN(n872) );
  INV_X1 U834 ( .A(n734), .ZN(n726) );
  AND2_X1 U835 ( .A1(n854), .A2(n873), .ZN(n734) );
  OR2_X1 U836 ( .A1(n710), .A2(n697), .ZN(n873) );
  AND2_X1 U837 ( .A1(n874), .A2(b_6_), .ZN(n697) );
  INV_X1 U838 ( .A(n687), .ZN(n710) );
  AND2_X1 U839 ( .A1(n875), .A2(a_7_), .ZN(n687) );
  INV_X1 U840 ( .A(n698), .ZN(n854) );
  AND2_X1 U841 ( .A1(n876), .A2(a_6_), .ZN(n698) );
  AND2_X1 U842 ( .A1(n877), .A2(a_0_), .ZN(n837) );
  AND2_X1 U843 ( .A1(n574), .A2(n878), .ZN(n831) );
  OR3_X1 U844 ( .A1(n681), .A2(n879), .A3(n880), .ZN(n878) );
  AND2_X1 U845 ( .A1(n881), .A2(a_0_), .ZN(n880) );
  INV_X1 U846 ( .A(n882), .ZN(n881) );
  AND2_X1 U847 ( .A1(n673), .A2(n678), .ZN(n879) );
  AND2_X1 U848 ( .A1(n669), .A2(n670), .ZN(n673) );
  XNOR2_X1 U849 ( .A(n680), .B(n883), .ZN(n670) );
  OR2_X1 U850 ( .A1(n884), .A2(n885), .ZN(n669) );
  OR2_X1 U851 ( .A1(n886), .A2(n666), .ZN(n884) );
  AND3_X1 U852 ( .A1(n665), .A2(n664), .A3(n662), .ZN(n666) );
  INV_X1 U853 ( .A(n887), .ZN(n664) );
  AND2_X1 U854 ( .A1(n658), .A2(n662), .ZN(n886) );
  INV_X1 U855 ( .A(n888), .ZN(n662) );
  OR2_X1 U856 ( .A1(n889), .A2(n885), .ZN(n888) );
  INV_X1 U857 ( .A(n890), .ZN(n885) );
  OR2_X1 U858 ( .A1(n891), .A2(n892), .ZN(n890) );
  AND2_X1 U859 ( .A1(n891), .A2(n892), .ZN(n889) );
  OR2_X1 U860 ( .A1(n893), .A2(n894), .ZN(n892) );
  AND2_X1 U861 ( .A1(n895), .A2(n896), .ZN(n894) );
  AND2_X1 U862 ( .A1(n897), .A2(n898), .ZN(n893) );
  OR2_X1 U863 ( .A1(n896), .A2(n895), .ZN(n898) );
  XOR2_X1 U864 ( .A(n899), .B(n900), .Z(n891) );
  XOR2_X1 U865 ( .A(n901), .B(n902), .Z(n900) );
  AND2_X1 U866 ( .A1(n903), .A2(n655), .ZN(n658) );
  XNOR2_X1 U867 ( .A(n665), .B(n887), .ZN(n655) );
  OR2_X1 U868 ( .A1(n904), .A2(n905), .ZN(n887) );
  AND2_X1 U869 ( .A1(n906), .A2(n907), .ZN(n905) );
  AND2_X1 U870 ( .A1(n908), .A2(n909), .ZN(n904) );
  OR2_X1 U871 ( .A1(n907), .A2(n906), .ZN(n909) );
  XOR2_X1 U872 ( .A(n910), .B(n897), .Z(n665) );
  XOR2_X1 U873 ( .A(n911), .B(n912), .Z(n897) );
  XOR2_X1 U874 ( .A(n913), .B(n914), .Z(n912) );
  XNOR2_X1 U875 ( .A(n896), .B(n895), .ZN(n910) );
  OR2_X1 U876 ( .A1(n915), .A2(n916), .ZN(n895) );
  AND2_X1 U877 ( .A1(n917), .A2(n918), .ZN(n916) );
  AND2_X1 U878 ( .A1(n919), .A2(n920), .ZN(n915) );
  OR2_X1 U879 ( .A1(n918), .A2(n917), .ZN(n920) );
  OR2_X1 U880 ( .A1(n818), .A2(n857), .ZN(n896) );
  INV_X1 U881 ( .A(n654), .ZN(n903) );
  AND2_X1 U882 ( .A1(n921), .A2(n922), .ZN(n654) );
  OR2_X1 U883 ( .A1(n650), .A2(n651), .ZN(n922) );
  OR2_X1 U884 ( .A1(n923), .A2(n924), .ZN(n651) );
  INV_X1 U885 ( .A(n921), .ZN(n924) );
  AND2_X1 U886 ( .A1(n925), .A2(n926), .ZN(n923) );
  AND2_X1 U887 ( .A1(n642), .A2(n927), .ZN(n650) );
  OR4_X1 U888 ( .A1(n639), .A2(n638), .A3(n928), .A4(n929), .ZN(n642) );
  AND2_X1 U889 ( .A1(n645), .A2(n646), .ZN(n929) );
  INV_X1 U890 ( .A(n927), .ZN(n928) );
  OR2_X1 U891 ( .A1(n645), .A2(n646), .ZN(n927) );
  OR2_X1 U892 ( .A1(n930), .A2(n931), .ZN(n646) );
  AND2_X1 U893 ( .A1(n932), .A2(n933), .ZN(n931) );
  AND2_X1 U894 ( .A1(n934), .A2(n935), .ZN(n930) );
  OR2_X1 U895 ( .A1(n933), .A2(n932), .ZN(n935) );
  XOR2_X1 U896 ( .A(n936), .B(n937), .Z(n645) );
  XOR2_X1 U897 ( .A(n938), .B(n939), .Z(n937) );
  OR2_X1 U898 ( .A1(n940), .A2(n941), .ZN(n638) );
  AND2_X1 U899 ( .A1(n608), .A2(n607), .ZN(n941) );
  AND2_X1 U900 ( .A1(n605), .A2(n942), .ZN(n940) );
  OR2_X1 U901 ( .A1(n607), .A2(n608), .ZN(n942) );
  OR2_X1 U902 ( .A1(n875), .A2(n857), .ZN(n608) );
  OR2_X1 U903 ( .A1(n943), .A2(n944), .ZN(n607) );
  AND2_X1 U904 ( .A1(n579), .A2(n578), .ZN(n944) );
  AND2_X1 U905 ( .A1(n576), .A2(n945), .ZN(n943) );
  OR2_X1 U906 ( .A1(n578), .A2(n579), .ZN(n945) );
  OR2_X1 U907 ( .A1(n875), .A2(n627), .ZN(n579) );
  OR2_X1 U908 ( .A1(n946), .A2(n947), .ZN(n578) );
  AND2_X1 U909 ( .A1(n795), .A2(n794), .ZN(n947) );
  AND2_X1 U910 ( .A1(n792), .A2(n948), .ZN(n946) );
  OR2_X1 U911 ( .A1(n795), .A2(n794), .ZN(n948) );
  OR2_X1 U912 ( .A1(n949), .A2(n950), .ZN(n794) );
  AND2_X1 U913 ( .A1(n769), .A2(n768), .ZN(n950) );
  AND2_X1 U914 ( .A1(n766), .A2(n951), .ZN(n949) );
  OR2_X1 U915 ( .A1(n769), .A2(n768), .ZN(n951) );
  OR2_X1 U916 ( .A1(n952), .A2(n953), .ZN(n768) );
  AND2_X1 U917 ( .A1(n744), .A2(n743), .ZN(n953) );
  AND2_X1 U918 ( .A1(n741), .A2(n954), .ZN(n952) );
  OR2_X1 U919 ( .A1(n744), .A2(n743), .ZN(n954) );
  OR2_X1 U920 ( .A1(n955), .A2(n956), .ZN(n743) );
  AND2_X1 U921 ( .A1(n719), .A2(n718), .ZN(n956) );
  AND2_X1 U922 ( .A1(n716), .A2(n957), .ZN(n955) );
  OR2_X1 U923 ( .A1(n719), .A2(n718), .ZN(n957) );
  OR2_X1 U924 ( .A1(n736), .A2(n875), .ZN(n718) );
  OR2_X1 U925 ( .A1(n711), .A2(n958), .ZN(n719) );
  INV_X1 U926 ( .A(n829), .ZN(n958) );
  INV_X1 U927 ( .A(n684), .ZN(n711) );
  AND2_X1 U928 ( .A1(a_7_), .A2(b_7_), .ZN(n684) );
  XOR2_X1 U929 ( .A(n959), .B(n829), .Z(n716) );
  AND2_X1 U930 ( .A1(a_6_), .A2(b_6_), .ZN(n829) );
  OR2_X1 U931 ( .A1(n761), .A2(n875), .ZN(n744) );
  XNOR2_X1 U932 ( .A(n960), .B(n961), .ZN(n741) );
  XNOR2_X1 U933 ( .A(n962), .B(n963), .ZN(n960) );
  OR2_X1 U934 ( .A1(n817), .A2(n875), .ZN(n769) );
  XOR2_X1 U935 ( .A(n964), .B(n965), .Z(n766) );
  XOR2_X1 U936 ( .A(n966), .B(n967), .Z(n965) );
  OR2_X1 U937 ( .A1(n808), .A2(n875), .ZN(n795) );
  INV_X1 U938 ( .A(b_7_), .ZN(n875) );
  XOR2_X1 U939 ( .A(n968), .B(n969), .Z(n792) );
  XOR2_X1 U940 ( .A(n970), .B(n971), .Z(n969) );
  XOR2_X1 U941 ( .A(n972), .B(n973), .Z(n576) );
  XOR2_X1 U942 ( .A(n974), .B(n975), .Z(n973) );
  XOR2_X1 U943 ( .A(n976), .B(n977), .Z(n605) );
  XOR2_X1 U944 ( .A(n978), .B(n979), .Z(n977) );
  XOR2_X1 U945 ( .A(n934), .B(n980), .Z(n639) );
  XOR2_X1 U946 ( .A(n933), .B(n932), .Z(n980) );
  OR2_X1 U947 ( .A1(n876), .A2(n857), .ZN(n932) );
  OR2_X1 U948 ( .A1(n981), .A2(n982), .ZN(n933) );
  AND2_X1 U949 ( .A1(n979), .A2(n978), .ZN(n982) );
  AND2_X1 U950 ( .A1(n976), .A2(n983), .ZN(n981) );
  OR2_X1 U951 ( .A1(n978), .A2(n979), .ZN(n983) );
  OR2_X1 U952 ( .A1(n876), .A2(n627), .ZN(n979) );
  OR2_X1 U953 ( .A1(n984), .A2(n985), .ZN(n978) );
  AND2_X1 U954 ( .A1(n975), .A2(n974), .ZN(n985) );
  AND2_X1 U955 ( .A1(n972), .A2(n986), .ZN(n984) );
  OR2_X1 U956 ( .A1(n974), .A2(n975), .ZN(n986) );
  OR2_X1 U957 ( .A1(n876), .A2(n808), .ZN(n975) );
  OR2_X1 U958 ( .A1(n987), .A2(n988), .ZN(n974) );
  AND2_X1 U959 ( .A1(n971), .A2(n970), .ZN(n988) );
  AND2_X1 U960 ( .A1(n968), .A2(n989), .ZN(n987) );
  OR2_X1 U961 ( .A1(n971), .A2(n970), .ZN(n989) );
  OR2_X1 U962 ( .A1(n990), .A2(n991), .ZN(n970) );
  AND2_X1 U963 ( .A1(n967), .A2(n966), .ZN(n991) );
  AND2_X1 U964 ( .A1(n964), .A2(n992), .ZN(n990) );
  OR2_X1 U965 ( .A1(n967), .A2(n966), .ZN(n992) );
  OR2_X1 U966 ( .A1(n993), .A2(n994), .ZN(n966) );
  AND2_X1 U967 ( .A1(n962), .A2(n963), .ZN(n994) );
  AND2_X1 U968 ( .A1(n961), .A2(n995), .ZN(n993) );
  OR2_X1 U969 ( .A1(n962), .A2(n963), .ZN(n995) );
  OR3_X1 U970 ( .A1(n855), .A2(n996), .A3(n876), .ZN(n963) );
  OR2_X1 U971 ( .A1(n736), .A2(n876), .ZN(n962) );
  XNOR2_X1 U972 ( .A(n996), .B(n997), .ZN(n961) );
  OR2_X1 U973 ( .A1(n874), .A2(n826), .ZN(n996) );
  OR2_X1 U974 ( .A1(n761), .A2(n876), .ZN(n967) );
  XOR2_X1 U975 ( .A(n998), .B(n999), .Z(n964) );
  XOR2_X1 U976 ( .A(n827), .B(n1000), .Z(n999) );
  OR2_X1 U977 ( .A1(n817), .A2(n876), .ZN(n971) );
  INV_X1 U978 ( .A(b_6_), .ZN(n876) );
  XOR2_X1 U979 ( .A(n1001), .B(n1002), .Z(n968) );
  XOR2_X1 U980 ( .A(n1003), .B(n1004), .Z(n1002) );
  XOR2_X1 U981 ( .A(n1005), .B(n1006), .Z(n972) );
  XOR2_X1 U982 ( .A(n1007), .B(n1008), .Z(n1006) );
  XOR2_X1 U983 ( .A(n1009), .B(n1010), .Z(n976) );
  XOR2_X1 U984 ( .A(n1011), .B(n1012), .Z(n1010) );
  XOR2_X1 U985 ( .A(n1013), .B(n1014), .Z(n934) );
  XOR2_X1 U986 ( .A(n1015), .B(n1016), .Z(n1014) );
  OR2_X1 U987 ( .A1(n925), .A2(n926), .ZN(n921) );
  OR2_X1 U988 ( .A1(n1017), .A2(n1018), .ZN(n926) );
  AND2_X1 U989 ( .A1(n936), .A2(n939), .ZN(n1018) );
  AND2_X1 U990 ( .A1(n1019), .A2(n938), .ZN(n1017) );
  OR2_X1 U991 ( .A1(n1020), .A2(n1021), .ZN(n938) );
  AND2_X1 U992 ( .A1(n1016), .A2(n1015), .ZN(n1021) );
  AND2_X1 U993 ( .A1(n1013), .A2(n1022), .ZN(n1020) );
  OR2_X1 U994 ( .A1(n1015), .A2(n1016), .ZN(n1022) );
  OR2_X1 U995 ( .A1(n826), .A2(n627), .ZN(n1016) );
  OR2_X1 U996 ( .A1(n1023), .A2(n1024), .ZN(n1015) );
  AND2_X1 U997 ( .A1(n1012), .A2(n1011), .ZN(n1024) );
  AND2_X1 U998 ( .A1(n1009), .A2(n1025), .ZN(n1023) );
  OR2_X1 U999 ( .A1(n1011), .A2(n1012), .ZN(n1025) );
  OR2_X1 U1000 ( .A1(n826), .A2(n808), .ZN(n1012) );
  OR2_X1 U1001 ( .A1(n1026), .A2(n1027), .ZN(n1011) );
  AND2_X1 U1002 ( .A1(n1008), .A2(n1007), .ZN(n1027) );
  AND2_X1 U1003 ( .A1(n1005), .A2(n1028), .ZN(n1026) );
  OR2_X1 U1004 ( .A1(n1007), .A2(n1008), .ZN(n1028) );
  OR2_X1 U1005 ( .A1(n826), .A2(n817), .ZN(n1008) );
  OR2_X1 U1006 ( .A1(n1029), .A2(n1030), .ZN(n1007) );
  AND2_X1 U1007 ( .A1(n1004), .A2(n1003), .ZN(n1030) );
  AND2_X1 U1008 ( .A1(n1001), .A2(n1031), .ZN(n1029) );
  OR2_X1 U1009 ( .A1(n1004), .A2(n1003), .ZN(n1031) );
  OR2_X1 U1010 ( .A1(n1032), .A2(n1033), .ZN(n1003) );
  AND2_X1 U1011 ( .A1(n1000), .A2(n827), .ZN(n1033) );
  AND2_X1 U1012 ( .A1(n998), .A2(n1034), .ZN(n1032) );
  OR2_X1 U1013 ( .A1(n1000), .A2(n827), .ZN(n1034) );
  OR2_X1 U1014 ( .A1(n736), .A2(n826), .ZN(n827) );
  OR2_X1 U1015 ( .A1(n959), .A2(n1035), .ZN(n1000) );
  OR2_X1 U1016 ( .A1(n855), .A2(n826), .ZN(n959) );
  XNOR2_X1 U1017 ( .A(n1036), .B(n1035), .ZN(n998) );
  OR2_X1 U1018 ( .A1(n874), .A2(n822), .ZN(n1035) );
  OR2_X1 U1019 ( .A1(n818), .A2(n855), .ZN(n1036) );
  OR2_X1 U1020 ( .A1(n761), .A2(n826), .ZN(n1004) );
  XNOR2_X1 U1021 ( .A(n1037), .B(n1038), .ZN(n1001) );
  XNOR2_X1 U1022 ( .A(n1039), .B(n1040), .ZN(n1037) );
  XNOR2_X1 U1023 ( .A(n1041), .B(n1042), .ZN(n1005) );
  XNOR2_X1 U1024 ( .A(n823), .B(n1043), .ZN(n1041) );
  XOR2_X1 U1025 ( .A(n1044), .B(n1045), .Z(n1009) );
  XOR2_X1 U1026 ( .A(n1046), .B(n1047), .Z(n1045) );
  XOR2_X1 U1027 ( .A(n1048), .B(n1049), .Z(n1013) );
  XOR2_X1 U1028 ( .A(n1050), .B(n1051), .Z(n1049) );
  OR2_X1 U1029 ( .A1(n939), .A2(n936), .ZN(n1019) );
  XOR2_X1 U1030 ( .A(n1052), .B(n1053), .Z(n936) );
  XOR2_X1 U1031 ( .A(n1054), .B(n1055), .Z(n1053) );
  OR2_X1 U1032 ( .A1(n826), .A2(n857), .ZN(n939) );
  INV_X1 U1033 ( .A(b_5_), .ZN(n826) );
  XOR2_X1 U1034 ( .A(n908), .B(n1056), .Z(n925) );
  XOR2_X1 U1035 ( .A(n907), .B(n906), .Z(n1056) );
  OR2_X1 U1036 ( .A1(n822), .A2(n857), .ZN(n906) );
  OR2_X1 U1037 ( .A1(n1057), .A2(n1058), .ZN(n907) );
  AND2_X1 U1038 ( .A1(n1052), .A2(n1055), .ZN(n1058) );
  AND2_X1 U1039 ( .A1(n1059), .A2(n1054), .ZN(n1057) );
  OR2_X1 U1040 ( .A1(n1060), .A2(n1061), .ZN(n1054) );
  AND2_X1 U1041 ( .A1(n1051), .A2(n1050), .ZN(n1061) );
  AND2_X1 U1042 ( .A1(n1048), .A2(n1062), .ZN(n1060) );
  OR2_X1 U1043 ( .A1(n1050), .A2(n1051), .ZN(n1062) );
  OR2_X1 U1044 ( .A1(n822), .A2(n808), .ZN(n1051) );
  OR2_X1 U1045 ( .A1(n1063), .A2(n1064), .ZN(n1050) );
  AND2_X1 U1046 ( .A1(n1047), .A2(n1046), .ZN(n1064) );
  AND2_X1 U1047 ( .A1(n1044), .A2(n1065), .ZN(n1063) );
  OR2_X1 U1048 ( .A1(n1046), .A2(n1047), .ZN(n1065) );
  OR2_X1 U1049 ( .A1(n822), .A2(n817), .ZN(n1047) );
  OR2_X1 U1050 ( .A1(n1066), .A2(n1067), .ZN(n1046) );
  AND2_X1 U1051 ( .A1(n1043), .A2(n823), .ZN(n1067) );
  AND2_X1 U1052 ( .A1(n1042), .A2(n1068), .ZN(n1066) );
  OR2_X1 U1053 ( .A1(n823), .A2(n1043), .ZN(n1068) );
  OR2_X1 U1054 ( .A1(n1069), .A2(n1070), .ZN(n1043) );
  AND2_X1 U1055 ( .A1(n1038), .A2(n1040), .ZN(n1070) );
  AND2_X1 U1056 ( .A1(n1071), .A2(n1039), .ZN(n1069) );
  OR2_X1 U1057 ( .A1(n1072), .A2(n1073), .ZN(n1039) );
  AND2_X1 U1058 ( .A1(n1074), .A2(n1075), .ZN(n1072) );
  OR2_X1 U1059 ( .A1(n1038), .A2(n1040), .ZN(n1071) );
  OR2_X1 U1060 ( .A1(n1075), .A2(n997), .ZN(n1040) );
  OR2_X1 U1061 ( .A1(n855), .A2(n822), .ZN(n997) );
  OR2_X1 U1062 ( .A1(n736), .A2(n822), .ZN(n1038) );
  OR2_X1 U1063 ( .A1(n761), .A2(n822), .ZN(n823) );
  XOR2_X1 U1064 ( .A(n1076), .B(n1073), .Z(n1042) );
  INV_X1 U1065 ( .A(n1077), .ZN(n1073) );
  XNOR2_X1 U1066 ( .A(n1078), .B(n1079), .ZN(n1076) );
  XNOR2_X1 U1067 ( .A(n1080), .B(n1081), .ZN(n1044) );
  XNOR2_X1 U1068 ( .A(n1082), .B(n1083), .ZN(n1080) );
  XNOR2_X1 U1069 ( .A(n1084), .B(n1085), .ZN(n1048) );
  XNOR2_X1 U1070 ( .A(n819), .B(n1086), .ZN(n1084) );
  OR2_X1 U1071 ( .A1(n1055), .A2(n1052), .ZN(n1059) );
  XNOR2_X1 U1072 ( .A(n1087), .B(n1088), .ZN(n1052) );
  XNOR2_X1 U1073 ( .A(n1089), .B(n1090), .ZN(n1087) );
  OR2_X1 U1074 ( .A1(n822), .A2(n627), .ZN(n1055) );
  INV_X1 U1075 ( .A(b_4_), .ZN(n822) );
  XNOR2_X1 U1076 ( .A(n1091), .B(n919), .ZN(n908) );
  XNOR2_X1 U1077 ( .A(n1092), .B(n1093), .ZN(n919) );
  XNOR2_X1 U1078 ( .A(n632), .B(n1094), .ZN(n1092) );
  XNOR2_X1 U1079 ( .A(n918), .B(n917), .ZN(n1091) );
  OR2_X1 U1080 ( .A1(n1095), .A2(n1096), .ZN(n917) );
  AND2_X1 U1081 ( .A1(n1090), .A2(n1089), .ZN(n1096) );
  AND2_X1 U1082 ( .A1(n1088), .A2(n1097), .ZN(n1095) );
  OR2_X1 U1083 ( .A1(n1089), .A2(n1090), .ZN(n1097) );
  OR2_X1 U1084 ( .A1(n1098), .A2(n1099), .ZN(n1090) );
  AND2_X1 U1085 ( .A1(n1086), .A2(n819), .ZN(n1099) );
  AND2_X1 U1086 ( .A1(n1085), .A2(n1100), .ZN(n1098) );
  OR2_X1 U1087 ( .A1(n819), .A2(n1086), .ZN(n1100) );
  OR2_X1 U1088 ( .A1(n1101), .A2(n1102), .ZN(n1086) );
  AND2_X1 U1089 ( .A1(n1083), .A2(n1082), .ZN(n1102) );
  AND2_X1 U1090 ( .A1(n1081), .A2(n1103), .ZN(n1101) );
  OR2_X1 U1091 ( .A1(n1082), .A2(n1083), .ZN(n1103) );
  OR2_X1 U1092 ( .A1(n1104), .A2(n1105), .ZN(n1083) );
  AND2_X1 U1093 ( .A1(n1077), .A2(n1079), .ZN(n1105) );
  AND2_X1 U1094 ( .A1(n1106), .A2(n1078), .ZN(n1104) );
  OR2_X1 U1095 ( .A1(n1107), .A2(n1108), .ZN(n1078) );
  INV_X1 U1096 ( .A(n1109), .ZN(n1108) );
  AND2_X1 U1097 ( .A1(n1110), .A2(n1111), .ZN(n1107) );
  OR2_X1 U1098 ( .A1(n1079), .A2(n1077), .ZN(n1106) );
  OR2_X1 U1099 ( .A1(n1074), .A2(n1075), .ZN(n1077) );
  OR2_X1 U1100 ( .A1(n874), .A2(n818), .ZN(n1075) );
  OR2_X1 U1101 ( .A1(n855), .A2(n809), .ZN(n1074) );
  OR2_X1 U1102 ( .A1(n818), .A2(n736), .ZN(n1079) );
  OR2_X1 U1103 ( .A1(n818), .A2(n761), .ZN(n1082) );
  XNOR2_X1 U1104 ( .A(n1112), .B(n1113), .ZN(n1081) );
  XNOR2_X1 U1105 ( .A(n1114), .B(n1109), .ZN(n1112) );
  INV_X1 U1106 ( .A(n783), .ZN(n819) );
  AND2_X1 U1107 ( .A1(b_3_), .A2(a_3_), .ZN(n783) );
  XNOR2_X1 U1108 ( .A(n1115), .B(n1116), .ZN(n1085) );
  XNOR2_X1 U1109 ( .A(n1117), .B(n1118), .ZN(n1115) );
  OR2_X1 U1110 ( .A1(n818), .A2(n808), .ZN(n1089) );
  XNOR2_X1 U1111 ( .A(n1119), .B(n1120), .ZN(n1088) );
  XNOR2_X1 U1112 ( .A(n1121), .B(n1122), .ZN(n1119) );
  OR2_X1 U1113 ( .A1(n818), .A2(n627), .ZN(n918) );
  INV_X1 U1114 ( .A(b_3_), .ZN(n818) );
  AND3_X1 U1115 ( .A1(n680), .A2(n678), .A3(n679), .ZN(n681) );
  INV_X1 U1116 ( .A(n883), .ZN(n679) );
  OR2_X1 U1117 ( .A1(n1123), .A2(n1124), .ZN(n883) );
  AND2_X1 U1118 ( .A1(n902), .A2(n901), .ZN(n1124) );
  AND2_X1 U1119 ( .A1(n899), .A2(n1125), .ZN(n1123) );
  OR2_X1 U1120 ( .A1(n901), .A2(n902), .ZN(n1125) );
  OR2_X1 U1121 ( .A1(n809), .A2(n857), .ZN(n902) );
  OR2_X1 U1122 ( .A1(n1126), .A2(n1127), .ZN(n901) );
  AND2_X1 U1123 ( .A1(n914), .A2(n913), .ZN(n1127) );
  AND2_X1 U1124 ( .A1(n911), .A2(n1128), .ZN(n1126) );
  OR2_X1 U1125 ( .A1(n913), .A2(n914), .ZN(n1128) );
  OR2_X1 U1126 ( .A1(n809), .A2(n627), .ZN(n914) );
  OR2_X1 U1127 ( .A1(n1129), .A2(n1130), .ZN(n913) );
  AND2_X1 U1128 ( .A1(n1094), .A2(n632), .ZN(n1130) );
  AND2_X1 U1129 ( .A1(n1093), .A2(n1131), .ZN(n1129) );
  OR2_X1 U1130 ( .A1(n632), .A2(n1094), .ZN(n1131) );
  OR2_X1 U1131 ( .A1(n1132), .A2(n1133), .ZN(n1094) );
  AND2_X1 U1132 ( .A1(n1121), .A2(n1122), .ZN(n1133) );
  AND2_X1 U1133 ( .A1(n1120), .A2(n1134), .ZN(n1132) );
  OR2_X1 U1134 ( .A1(n1122), .A2(n1121), .ZN(n1134) );
  OR2_X1 U1135 ( .A1(n1135), .A2(n1136), .ZN(n1121) );
  AND2_X1 U1136 ( .A1(n1118), .A2(n1117), .ZN(n1136) );
  AND2_X1 U1137 ( .A1(n1116), .A2(n1137), .ZN(n1135) );
  OR2_X1 U1138 ( .A1(n1117), .A2(n1118), .ZN(n1137) );
  OR2_X1 U1139 ( .A1(n809), .A2(n761), .ZN(n1118) );
  OR2_X1 U1140 ( .A1(n1138), .A2(n1139), .ZN(n1117) );
  AND2_X1 U1141 ( .A1(n1113), .A2(n1109), .ZN(n1139) );
  AND2_X1 U1142 ( .A1(n1140), .A2(n1114), .ZN(n1138) );
  OR2_X1 U1143 ( .A1(n1141), .A2(n1142), .ZN(n1114) );
  INV_X1 U1144 ( .A(n1143), .ZN(n1142) );
  AND2_X1 U1145 ( .A1(n1144), .A2(n1145), .ZN(n1141) );
  OR2_X1 U1146 ( .A1(n855), .A2(n877), .ZN(n1144) );
  OR2_X1 U1147 ( .A1(n1109), .A2(n1113), .ZN(n1140) );
  OR2_X1 U1148 ( .A1(n809), .A2(n736), .ZN(n1113) );
  OR2_X1 U1149 ( .A1(n1110), .A2(n1111), .ZN(n1109) );
  OR2_X1 U1150 ( .A1(n874), .A2(n809), .ZN(n1111) );
  OR2_X1 U1151 ( .A1(n855), .A2(n628), .ZN(n1110) );
  XNOR2_X1 U1152 ( .A(n1146), .B(n1143), .ZN(n1116) );
  OR2_X1 U1153 ( .A1(n1147), .A2(n1148), .ZN(n1146) );
  INV_X1 U1154 ( .A(n1149), .ZN(n1148) );
  AND2_X1 U1155 ( .A1(n1150), .A2(n1151), .ZN(n1147) );
  OR2_X1 U1156 ( .A1(n874), .A2(n877), .ZN(n1150) );
  OR2_X1 U1157 ( .A1(n809), .A2(n817), .ZN(n1122) );
  INV_X1 U1158 ( .A(b_2_), .ZN(n809) );
  XOR2_X1 U1159 ( .A(n1152), .B(n1153), .Z(n1120) );
  XOR2_X1 U1160 ( .A(n1154), .B(n1155), .Z(n1152) );
  INV_X1 U1161 ( .A(n807), .ZN(n632) );
  AND2_X1 U1162 ( .A1(b_2_), .A2(a_2_), .ZN(n807) );
  XOR2_X1 U1163 ( .A(n1156), .B(n1157), .Z(n1093) );
  XOR2_X1 U1164 ( .A(n1158), .B(n1159), .Z(n1157) );
  XOR2_X1 U1165 ( .A(n1160), .B(n1161), .Z(n911) );
  XOR2_X1 U1166 ( .A(n1162), .B(n1163), .Z(n1161) );
  XNOR2_X1 U1167 ( .A(n1164), .B(n1165), .ZN(n899) );
  XNOR2_X1 U1168 ( .A(n596), .B(n1166), .ZN(n1164) );
  XOR2_X1 U1169 ( .A(n1167), .B(n882), .Z(n678) );
  OR2_X1 U1170 ( .A1(n1168), .A2(n1169), .ZN(n882) );
  AND2_X1 U1171 ( .A1(n1170), .A2(n1171), .ZN(n1169) );
  AND2_X1 U1172 ( .A1(n1172), .A2(n1173), .ZN(n1168) );
  OR2_X1 U1173 ( .A1(n1171), .A2(n1170), .ZN(n1172) );
  OR2_X1 U1174 ( .A1(n877), .A2(n857), .ZN(n1167) );
  XNOR2_X1 U1175 ( .A(n1170), .B(n1174), .ZN(n680) );
  XOR2_X1 U1176 ( .A(n1171), .B(n1173), .Z(n1174) );
  OR2_X1 U1177 ( .A1(n628), .A2(n857), .ZN(n1173) );
  INV_X1 U1178 ( .A(a_0_), .ZN(n857) );
  OR2_X1 U1179 ( .A1(n1175), .A2(n1176), .ZN(n1171) );
  AND2_X1 U1180 ( .A1(n1165), .A2(n1166), .ZN(n1176) );
  AND2_X1 U1181 ( .A1(n1177), .A2(n596), .ZN(n1175) );
  OR2_X1 U1182 ( .A1(n628), .A2(n627), .ZN(n596) );
  OR2_X1 U1183 ( .A1(n1166), .A2(n1165), .ZN(n1177) );
  OR2_X1 U1184 ( .A1(n808), .A2(n877), .ZN(n1165) );
  OR2_X1 U1185 ( .A1(n1178), .A2(n1179), .ZN(n1166) );
  AND2_X1 U1186 ( .A1(n1160), .A2(n1162), .ZN(n1179) );
  AND2_X1 U1187 ( .A1(n1180), .A2(n1163), .ZN(n1178) );
  OR2_X1 U1188 ( .A1(n817), .A2(n877), .ZN(n1163) );
  OR2_X1 U1189 ( .A1(n1162), .A2(n1160), .ZN(n1180) );
  OR2_X1 U1190 ( .A1(n628), .A2(n808), .ZN(n1160) );
  INV_X1 U1191 ( .A(a_2_), .ZN(n808) );
  OR2_X1 U1192 ( .A1(n1181), .A2(n1182), .ZN(n1162) );
  AND2_X1 U1193 ( .A1(n1156), .A2(n1158), .ZN(n1182) );
  AND2_X1 U1194 ( .A1(n1183), .A2(n1159), .ZN(n1181) );
  OR2_X1 U1195 ( .A1(n628), .A2(n817), .ZN(n1159) );
  INV_X1 U1196 ( .A(a_3_), .ZN(n817) );
  OR2_X1 U1197 ( .A1(n1158), .A2(n1156), .ZN(n1183) );
  OR2_X1 U1198 ( .A1(n761), .A2(n877), .ZN(n1156) );
  OR2_X1 U1199 ( .A1(n1184), .A2(n1185), .ZN(n1158) );
  AND2_X1 U1200 ( .A1(n1153), .A2(n1155), .ZN(n1185) );
  AND2_X1 U1201 ( .A1(n1154), .A2(n1186), .ZN(n1184) );
  OR2_X1 U1202 ( .A1(n1155), .A2(n1153), .ZN(n1186) );
  OR2_X1 U1203 ( .A1(n736), .A2(n877), .ZN(n1153) );
  OR2_X1 U1204 ( .A1(n628), .A2(n761), .ZN(n1155) );
  INV_X1 U1205 ( .A(a_4_), .ZN(n761) );
  AND2_X1 U1206 ( .A1(n1149), .A2(n1143), .ZN(n1154) );
  OR3_X1 U1207 ( .A1(n855), .A2(n877), .A3(n1145), .ZN(n1143) );
  OR2_X1 U1208 ( .A1(n874), .A2(n628), .ZN(n1145) );
  INV_X1 U1209 ( .A(a_7_), .ZN(n855) );
  OR3_X1 U1210 ( .A1(n874), .A2(n877), .A3(n1151), .ZN(n1149) );
  OR2_X1 U1211 ( .A1(n628), .A2(n736), .ZN(n1151) );
  INV_X1 U1212 ( .A(a_5_), .ZN(n736) );
  INV_X1 U1213 ( .A(b_1_), .ZN(n628) );
  INV_X1 U1214 ( .A(a_6_), .ZN(n874) );
  OR2_X1 U1215 ( .A1(n627), .A2(n877), .ZN(n1170) );
  INV_X1 U1216 ( .A(b_0_), .ZN(n877) );
  INV_X1 U1217 ( .A(a_1_), .ZN(n627) );
  AND2_X1 U1218 ( .A1(operation_0_), .A2(operation_1_), .ZN(n574) );
endmodule

