module s15850 ( CK, g100, g101, g102, g103, g10377, g10379, g104, g10455, 
        g10457, g10459, g10461, g10463, g10465, g10628, g10801, g109, g11163, 
        g11206, g11489, g1170, g1173, g1176, g1179, g1182, g1185, g1188, g1191, 
        g1194, g1197, g1200, g1203, g1696, g1700, g1712, g18, g1957, g1960, 
        g1961, g23, g2355, g2601, g2602, g2603, g2604, g2605, g2606, g2607, 
        g2608, g2609, g2610, g2611, g2612, g2648, g27, g28, g29, g2986, g30, 
        g3007, g3069, g31, g3327, g41, g4171, g4172, g4173, g4174, g4175, 
        g4176, g4177, g4178, g4179, g4180, g4181, g4191, g4192, g4193, g4194, 
        g4195, g4196, g4197, g4198, g4199, g42, g4200, g4201, g4202, g4203, 
        g4204, g4205, g4206, g4207, g4208, g4209, g4210, g4211, g4212, g4213, 
        g4214, g4215, g4216, g43, g44, g45, g46, g47, g48, g4887, g4888, g5101, 
        g5105, g5658, g5659, g5816, g6253, g6254, g6255, g6256, g6257, g6258, 
        g6259, g6260, g6261, g6262, g6263, g6264, g6265, g6266, g6267, g6268, 
        g6269, g6270, g6271, g6272, g6273, g6274, g6275, g6276, g6277, g6278, 
        g6279, g6280, g6281, g6282, g6283, g6284, g6285, g6842, g6920, g6926, 
        g6932, g6942, g6949, g6955, g741, g742, g743, g744, g750, g7744, g8061, 
        g8062, g82, g8271, g83, g8313, g8316, g8318, g8323, g8328, g8331, 
        g8335, g8340, g8347, g8349, g8352, g84, g85, g8561, g8562, g8563, 
        g8564, g8565, g8566, g86, g87, g872, g873, g877, g88, g881, g886, g889, 
        g89, g892, g895, g8976, g8977, g8978, g8979, g898, g8980, g8981, g8982, 
        g8983, g8984, g8985, g8986, g90, g901, g904, g907, g91, g910, g913, 
        g916, g919, g92, g922, g925, g93, g94, g9451, g95, g96, g99, g9961, 
        test_se, test_si1, test_so1, test_si2, test_so2, test_si3, test_so3, 
        test_si4, test_so4, test_si5, test_so5, test_si6, test_so6, test_si7, 
        test_so7, test_si8, test_so8, test_si9, test_so9, test_si10, test_so10
 );
  input CK, g100, g101, g102, g103, g104, g109, g1170, g1173, g1176, g1179,
         g1182, g1185, g1188, g1191, g1194, g1197, g1200, g1203, g1696, g1700,
         g1712, g18, g1960, g1961, g23, g27, g28, g29, g30, g31, g41, g42, g43,
         g44, g45, g46, g47, g48, g741, g742, g743, g744, g750, g82, g83, g84,
         g85, g86, g87, g872, g873, g877, g88, g881, g886, g889, g89, g892,
         g895, g898, g90, g901, g904, g907, g91, g910, g913, g916, g919, g92,
         g922, g925, g93, g94, g95, g96, g99, test_se, test_si1, test_si2,
         test_si3, test_si4, test_si5, test_si6, test_si7, test_si8, test_si9,
         test_si10;
  output g10377, g10379, g10455, g10457, g10459, g10461, g10463, g10465,
         g10628, g10801, g11163, g11206, g11489, g1957, g2355, g2601, g2602,
         g2603, g2604, g2605, g2606, g2607, g2608, g2609, g2610, g2611, g2612,
         g2648, g2986, g3007, g3069, g3327, g4171, g4172, g4173, g4174, g4175,
         g4176, g4177, g4178, g4179, g4180, g4181, g4191, g4192, g4193, g4194,
         g4195, g4196, g4197, g4198, g4199, g4200, g4201, g4202, g4203, g4204,
         g4205, g4206, g4207, g4208, g4209, g4210, g4211, g4212, g4213, g4214,
         g4215, g4216, g4887, g4888, g5101, g5105, g5658, g5659, g5816, g6253,
         g6254, g6255, g6256, g6257, g6258, g6259, g6260, g6261, g6262, g6263,
         g6264, g6265, g6266, g6267, g6268, g6269, g6270, g6271, g6272, g6273,
         g6274, g6275, g6276, g6277, g6278, g6279, g6280, g6281, g6282, g6283,
         g6284, g6285, g6842, g6920, g6926, g6932, g6942, g6949, g6955, g7744,
         g8061, g8062, g8271, g8313, g8316, g8318, g8323, g8328, g8331, g8335,
         g8340, g8347, g8349, g8352, g8561, g8562, g8563, g8564, g8565, g8566,
         g8976, g8977, g8978, g8979, g8980, g8981, g8982, g8983, g8984, g8985,
         g8986, g9451, g9961, test_so1, test_so2, test_so3, test_so4, test_so5,
         test_so6, test_so7, test_so8, test_so9, test_so10;
  wire   g100, g101, g102, g103, g104, g1170, g1173, g1176, g1179, g1182,
         g1185, g1188, g1191, g1194, g1197, g1203, g18, g1960, g1961, g27, g28,
         g29, g30, g31, g41, g42, g43, g44, g45, g46, g47, g48, g5816, g82,
         g83, g84, g85, g8561, g8562, g8563, g8564, g8565, g8566, g86, g87,
         g872, g873, g88, g886, g889, g89, g892, g895, g898, g90, g901, g904,
         g907, g91, g910, g913, g916, g919, g92, g922, g925, g93, g94, g9451,
         g95, g96, g99, test_so10, g10722, g10664, g1289, g8943, g1882, n1663,
         g255, g312, g11257, g452, g7032, g123, g6830, g207, g8920, g713,
         g4340, g1153, n1686, g4239, g1744, g6538, g1558, g8887, g695, g11372,
         g461, n1594, g8260, g940, g11391, g976, g8432, g709, n1719, g6088,
         g1092, g6478, g1574, g6795, g1864, g11320, g369, g6500, g1580, g5392,
         g1736, g10663, n1637, g10782, n3065, g6216, g1424, g1737, g10858,
         g1672, g5914, g1077, g7590, g1231, g6656, g4, g6728, g5126, g1104,
         n1658, g7290, g1304, g6841, g243, g8041, g1499, g8766, g1444, n3064,
         g8019, g6545, g1543, g256, g315, g6533, g1534, g8820, g622, n1713,
         g8941, g1927, g10859, g1660, g6922, g278, g8772, g1436, g8433, g718,
         g6526, g10793, g554, g11333, g496, n1689, g11392, g981, n1720, g794,
         g829, g6093, g1095, g8889, g704, g7302, g1265, g6525, g1786, g8429,
         g682, g7292, g1296, g6621, g7134, n3062, g260, g327, g6333, g1389,
         g6826, g1371, g1955, g1956, g10860, g1675, g11483, g354, g6392, g113,
         g7626, g639, n1692, g10866, g1684, g8193, g1639, g6983, g1791, n1702,
         g6839, g248, g4076, g1707, g4293, g1759, g11482, g351, g6507, g1604,
         g6096, g1098, g8250, g932, g8282, g1896, g8435, g736, g6924, g1019,
         g6819, n3061, g746, g745, g6244, g1419, n1602, g6627, g32, n1865,
         g6071, g1086, g8046, g1486, g10707, g1730, g6198, g1504, g8051, g1470,
         g8024, g822, g10862, g1678, g8050, g174, g7133, g1766, g7930, g1801,
         g6832, g186, g11308, g959, g6918, g8769, g1407, g6909, g1868, g4940,
         g5404, g1718, n1611, g11265, g396, g6930, g1015, g10726, n1650, g4891,
         n3059, n1874, g6224, g1415, g7586, g1227, g10770, g1721, n3058, n3057,
         g6934, g284, g11256, g426, g6824, g219, g1360, n3056, g6126, g806,
         g8767, g1428, g6546, g1564, g4238, g1741, g6823, g225, g6928, g281,
         g11602, g1308, g9721, g611, n1609, g4890, n3055, n1586, g1217, g6524,
         g1589, g8045, g1466, g6469, g1571, g6471, g1861, g6821, n3054, g11514,
         g1448, g1133, n1706, g11610, g1333, g7843, g153, g11310, g962, g5536,
         g11331, g486, n1621, g11380, g471, n1606, g6838, g1397, g8288, g1950,
         g755, g756, n3053, g10855, g1101, g549, g10898, g105, g10865, g1669,
         g6822, g6528, g1531, g6180, g1458, n1703, g10718, g572, g6912, g1011,
         g10719, n3051, g6234, g1411, g6099, g1074, g11259, g444, g8039, g1474,
         g6059, g1080, g5396, g1713, n1610, g262, g333, g6906, g269, g11266,
         g401, g11294, g1857, n1682, g5421, g9, g8649, g664, g11312, g965,
         g6840, g1400, g254, g309, g7202, g814, g6834, g231, g10795, g557,
         g875, g869, g6831, g1383, g8060, g158, g4893, g627, g7244, g1023,
         g6026, g259, n3050, g11608, g1327, g7660, g654, g6911, g293, g11640,
         g1346, g8777, g1633, g4274, g1753, g1508, n1707, g7297, g1240, g11326,
         g538, g11269, g416, g11325, g542, g10864, g1681, g11290, g374, g10798,
         g563, g8284, g1914, g11328, g530, g10800, g575, g8944, g1936, n1694,
         g7183, g4465, g1356, g1317, g11484, g357, g11263, g386, g6501, g1601,
         g6757, g166, g11334, g501, n1690, g6042, g8384, g1840, g6653, g257,
         g318, g5763, g5849, n3048, g6929, g302, g11488, g342, g7299, g1250,
         g4330, g1163, g1958, n3047, g7257, g1032, g8775, g1432, g5770, g1453,
         n1628, g11486, g363, g261, g330, g4338, g1157, g4500, n3046, g10721,
         n3045, g8147, g928, g6038, g11337, g516, n1620, g6045, g7191, g826,
         g861, g8774, g1627, g7293, g1292, g6907, g290, g4903, n3044, n1873,
         g6123, g6506, g1583, g11376, g466, n1646, g6542, g1561, g6551, g1546,
         g6901, g287, g10797, g560, g8505, g617, n1645, n1631, g11647, g336,
         g11340, g456, n1641, g253, g305, n1681, g11625, g345, g636, g8, g6502,
         N599, g6049, g8945, g1945, n1697, g4231, g1738, g8040, g1478, n3042,
         g6155, g1690, n1653, g8043, g1482, g5173, g1110, n1677, g6916, g296,
         g10861, g1663, g8431, g700, g4309, g1762, g11485, g360, g6334, g192,
         g10767, g1657, g8923, g722, n1693, g7189, g10799, g566, g6747, n3041,
         g6080, g1089, g3381, g5910, g1071, g11393, g986, n1722, g11349, g971,
         g6439, g143, g9266, g1814, n1608, g1212, g8940, g1918, g7705, g9269,
         g1822, n1643, g6820, g237, g8042, g1462, g6759, g178, g11487, g366,
         g802, g837, g9124, g599, n1644, g11293, g1854, g11298, g944, g8287,
         g1941, g8047, g170, g6205, g1520, n1710, g8885, g686, n1676, g11305,
         g953, g5556, n3040, g2478, g1765, g10711, g1733, g7303, g5194, g1610,
         g7541, g1796, n1626, g11607, g1324, g6541, g1540, g6827, n3038,
         g11332, g491, n1691, g4902, n3037, g6828, g213, g6516, g1781, n1659,
         g8938, g1900, n1675, g7298, g1245, n3036, n3035, g8048, g148, g798,
         g833, g8285, g1923, n1718, g8254, g936, g11604, g1314, g849, g11636,
         g1336, g6910, g272, g8173, g1806, g8245, n1716, g8281, g1887, g10724,
         n3034, g11314, g968, g4905, n3033, g1137, n1597, g8937, g1891, n1657,
         g7300, g1255, g6002, n1588, g874, g9110, g591, n1607, g8926, g731,
         n1696, g8631, g7632, g1218, g9150, g605, n1593, g6531, g6786, g182,
         g11303, g950, g4477, g1129, n1705, g857, g11258, g448, g9272, g1828,
         n1605, g10773, g1727, g6470, g1592, g5083, g1703, g8286, g1932, g8773,
         g1624, g6054, g11260, g440, g11338, g476, n1599, g5918, g119, n1613,
         g8922, g668, n1662, g8049, g139, g4342, g1149, n1685, g10720, n3031,
         g6755, n3030, g6897, g263, g7709, g818, g4255, g1747, g5543, n1622,
         g6915, g275, g6513, g1524, g6480, g1577, g6733, g810, g11264, g391,
         g8973, g658, n1615, g6833, g1386, g5996, n1587, g4473, g1125, n1708,
         g5755, g201, n1619, g7295, g1280, n1862, g6068, g1083, g7137, g650,
         n1709, g8779, g1636, g853, g11270, g421, g5529, g11306, g956, g11291,
         g378, g4283, g1756, g841, g6894, g1027, g6902, g1003, g8765, g1403,
         g1145, n1617, g5148, g1107, n1614, g7581, g1223, g11267, g406, g10936,
         g1811, n1699, g10784, n3029, g10765, g1654, g6332, g197, n1678, g6479,
         g1595, g6537, g1537, g8434, g727, g6908, g6243, n1717, g11324, g481,
         n1680, n1647, g11609, g1330, g845, g8244, g8194, g1512, n3027,
         DFF_436_n1, g8052, g1490, g4325, g1166, g11481, g348, n3026, g7301,
         g1260, g6035, g8059, g131, n3025, g6015, g258, g11330, g521, n1698,
         g11605, g1318, g8921, g1872, n1616, g8883, g677, n1656, n3024, g6523,
         g1549, g11300, g947, g9555, g1834, n1655, g6481, g1598, g4471, g1121,
         n1618, g11606, g1321, g11335, g506, n1600, g10791, g546, g8939, g1909,
         g6529, g1552, g10776, g1687, g6514, g1586, g324, g1141, n1660, g11639,
         g1341, g4089, g1710, g10785, n3023, g6179, n3022, g8053, g135, g11329,
         g525, n1695, g6515, g1607, g321, g7204, g11443, g1275, g11603, g8770,
         g1615, g11292, g382, g6331, n3020, g6900, g266, g7294, g1284, n1864,
         g6829, n3019, g8428, g673, n3018, g8054, g162, g11268, g411, g11262,
         g431, n1876, g8283, g1905, g6193, g1515, n1627, g8776, g1630, g7143,
         g6898, g991, n1871, g7291, g1300, g11478, g339, g6000, g4264, g1750,
         g8768, g1440, g10863, g1666, g6522, g1528, g11641, g1351, n1721,
         g10780, n3017, g8044, g127, n1704, g11579, g1618, g7296, g1235, g6923,
         g299, g11261, g435, n1878, g6638, g6534, g1555, g6895, g995, g8771,
         g1621, g4506, n3016, g7441, g643, n1612, g8055, g1494, g6468, g1567,
         g8430, g691, g11327, g534, g6508, g1776, n1715, g10717, g569, g4334,
         g1160, n1585, g6679, g1, g11336, g511, n1679, g10771, g1724, g5445,
         g12, g8559, g1878, g7219, g5390, n1654, n1512, n1486, n1485, n1545,
         n1530, n1420, n1855, n1239, n1566, n1567, n1479, n1858, n1480, n1478,
         n1137, n1195, n1404, n1262, n1227, n1450, n916, n822, n958, n918,
         n1159, n812, n1056, n1258, n817, n837, n804, n1016, n1380, n926,
         n1385, n1391, n1564, n1231, n1226, n1232, n1260, n1107, n1154, n1093,
         n1214, n931, n962, n902, n1147, n1193, n1153, n1125, n1099, n857,
         n806, n808, n1097, n1123, n1151, n1090, n1161, n967, n921, n1055,
         n1150, n1096, n1098, n1213, n1152, n836, n838, Tg1_OUT1, Tg1_OUT2,
         Tg1_OUT3, Tg1_OUT4, Tg1_OUT5, Tg1_OUT6, Tg1_OUT7, Tg1_OUT8, Tg2_OUT1,
         Tg2_OUT2, Tg2_OUT3, Tg2_OUT4, Tg2_OUT5, Tg2_OUT6, Tg2_OUT7, Tg2_OUT8,
         test_se_NOT, Trigger_select, n1, n6, n9, n13, n25, n29, n30, n32, n45,
         n72, n74, n103, n104, n145, n160, n178, n187, n225, n250, n252, n269,
         n316, n352, n369, n371, n407, n444, n499, n503, n519, n521, n524,
         n525, n529, n530, n534, n535, n2605, n2606, n2628, n2629, n2649,
         n2650, n2651, n2657, n2696, n2714, n2721, n2739, n2740, n2741, n2742,
         n2745, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2792, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2855, n2856, n2857, n2858, n2859, n2860, n2862,
         n2864, n2865, n2866, n2869, n2870, n2871, n2872, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2885, n2886, n2887, n2888, n2889, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3021, n3028, n3032, n3039, n3043, n3049,
         n3052, n3060, n3063, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         U1586_n1, U1754_n1, U1798_n1, U1839_n1, U1843_n1, U1877_n1, U1908_n1,
         U1909_n1, U1987_n1, U2031_n1, U2035_n1, U2418_n1, U2468_n1, U2478_n1,
         U2488_n1, U2533_n1, U2534_n1, U2639_n1, U2641_n1, U2654_n1, U2658_n1,
         U2683_n1, U2699_n1, U2846_n1, U2847_n1, U2848_n1, U2859_n1, U2860_n1,
         U2861_n1, U2867_n1, U2879_n1, U2881_n1, U2882_n1, U2883_n1, U2884_n1,
         U2885_n1, U2886_n1, U2887_n1, U2888_n1, U2889_n1, U2890_n1, U2891_n1,
         U2892_n1, U2893_n1, U2894_n1, U2895_n1, U2896_n1, U2897_n1, U2898_n1,
         U2899_n1, U2900_n1, U2901_n1, U2902_n1, U3090_n1, U3092_n1, U3094_n1,
         U3096_n1, U3098_n1, U3124_n1, U3171_n1;
  assign g11489 = 1'b0;
  assign g6280 = g100;
  assign g6281 = g101;
  assign g6282 = g102;
  assign g6283 = g103;
  assign g6284 = g104;
  assign g4205 = g1170;
  assign g4209 = g1173;
  assign g4210 = g1176;
  assign g4211 = g1179;
  assign g4212 = g1182;
  assign g4213 = g1185;
  assign g4214 = g1188;
  assign g4215 = g1191;
  assign g4216 = g1194;
  assign g4206 = g1197;
  assign g4208 = g1203;
  assign g2355 = g18;
  assign g4888 = g1960;
  assign g4887 = g1961;
  assign g7744 = g27;
  assign g6285 = g28;
  assign g6253 = g29;
  assign g6254 = g30;
  assign g6255 = g31;
  assign g6256 = g41;
  assign g6257 = g42;
  assign g6258 = g43;
  assign g6259 = g44;
  assign g6260 = g45;
  assign g6261 = g46;
  assign g6262 = g47;
  assign g6263 = g48;
  assign g8271 = g5816;
  assign g6264 = g82;
  assign g6265 = g83;
  assign g6266 = g84;
  assign g6267 = g85;
  assign g6920 = g8561;
  assign g6926 = g8562;
  assign g6932 = g8563;
  assign g6942 = g8564;
  assign g6949 = g8565;
  assign g6955 = g8566;
  assign g6268 = g86;
  assign g6269 = g87;
  assign g5101 = g872;
  assign g8061 = g872;
  assign g5105 = g873;
  assign g8062 = g873;
  assign g6270 = g88;
  assign g4191 = g886;
  assign g4192 = g889;
  assign g6271 = g89;
  assign g4193 = g892;
  assign g4194 = g895;
  assign g4195 = g898;
  assign g6272 = g90;
  assign g4197 = g901;
  assign g4198 = g904;
  assign g4199 = g907;
  assign g6273 = g91;
  assign g4200 = g910;
  assign g4201 = g913;
  assign g4202 = g916;
  assign g4203 = g919;
  assign g6274 = g92;
  assign g4204 = g922;
  assign g4196 = g925;
  assign g6275 = g93;
  assign g6276 = g94;
  assign g9961 = g9451;
  assign g6277 = g95;
  assign g6278 = g96;
  assign g6279 = g99;
  assign g8984 = test_so10;

  SDFFX1 DFF_0_Q_reg ( .D(n1), .SI(test_si1), .SE(n2994), .CLK(n3075), .Q(
        g1289), .QN(n2844) );
  SDFFX1 DFF_1_Q_reg ( .D(g8943), .SI(g1289), .SE(n2972), .CLK(n3085), .Q(
        g1882), .QN(n1663) );
  SDFFX1 DFF_2_Q_reg ( .D(g255), .SI(g1882), .SE(n2935), .CLK(n3104), .Q(g312), 
        .QN(n2797) );
  SDFFX1 DFF_3_Q_reg ( .D(g11257), .SI(g312), .SE(n2985), .CLK(n3079), .Q(g452) );
  SDFFX1 DFF_4_Q_reg ( .D(g7032), .SI(g452), .SE(n2974), .CLK(n3084), .Q(g123)
         );
  SDFFX1 DFF_5_Q_reg ( .D(g6830), .SI(g123), .SE(n2974), .CLK(n3084), .Q(g207), 
        .QN(n2878) );
  SDFFX1 DFF_6_Q_reg ( .D(g8920), .SI(g207), .SE(n2988), .CLK(n3078), .Q(g713)
         );
  SDFFX1 DFF_7_Q_reg ( .D(g4340), .SI(g713), .SE(n2987), .CLK(n3078), .Q(g1153), .QN(n1686) );
  SDFFX1 DFF_9_Q_reg ( .D(g4239), .SI(g1153), .SE(n2910), .CLK(n3117), .Q(
        g1744) );
  SDFFX1 DFF_10_Q_reg ( .D(g6538), .SI(g1744), .SE(n2910), .CLK(n3117), .Q(
        g1558) );
  SDFFX1 DFF_11_Q_reg ( .D(g8887), .SI(g1558), .SE(n2988), .CLK(n3078), .Q(
        g695), .QN(n2850) );
  SDFFX1 DFF_12_Q_reg ( .D(g11372), .SI(g695), .SE(n2926), .CLK(n3108), .Q(
        g461), .QN(n1594) );
  SDFFX1 DFF_13_Q_reg ( .D(g8260), .SI(g461), .SE(n2926), .CLK(n3108), .Q(g940) );
  SDFFX1 DFF_14_Q_reg ( .D(g11391), .SI(g940), .SE(n2926), .CLK(n3109), .Q(
        g976), .QN(n2892) );
  SDFFX1 DFF_15_Q_reg ( .D(g8432), .SI(g976), .SE(n2926), .CLK(n3109), .Q(g709), .QN(n1719) );
  SDFFX1 DFF_16_Q_reg ( .D(g6088), .SI(g709), .SE(n2959), .CLK(n3092), .Q(
        g1092) );
  SDFFX1 DFF_17_Q_reg ( .D(g6478), .SI(g1092), .SE(n2916), .CLK(n3113), .Q(
        g1574) );
  SDFFX1 DFF_18_Q_reg ( .D(g6795), .SI(g1574), .SE(n2916), .CLK(n3114), .Q(
        g1864) );
  SDFFX1 DFF_19_Q_reg ( .D(g11320), .SI(g1864), .SE(n2916), .CLK(n3114), .Q(
        g369), .QN(n2894) );
  SDFFX1 DFF_20_Q_reg ( .D(g6500), .SI(g369), .SE(n2958), .CLK(n3092), .Q(
        g1580) );
  SDFFX1 DFF_21_Q_reg ( .D(g5392), .SI(g1580), .SE(n2958), .CLK(n3093), .Q(
        g1736) );
  SDFFX1 DFF_22_Q_reg ( .D(g10663), .SI(g1736), .SE(n2958), .CLK(n3093), .Q(
        n1637) );
  SDFFX1 DFF_23_Q_reg ( .D(g10782), .SI(n1637), .SE(n2958), .CLK(n3093), .Q(
        n3065) );
  SDFFX1 DFF_24_Q_reg ( .D(g6216), .SI(n3065), .SE(n2929), .CLK(n3107), .Q(
        g1424) );
  SDFFX1 DFF_25_Q_reg ( .D(g1736), .SI(g1424), .SE(n2929), .CLK(n3107), .Q(
        g1737), .QN(n2849) );
  SDFFX1 DFF_26_Q_reg ( .D(g10858), .SI(g1737), .SE(n2993), .CLK(n3075), .Q(
        g1672) );
  SDFFX1 DFF_27_Q_reg ( .D(g5914), .SI(g1672), .SE(n2993), .CLK(n3075), .Q(
        g1077) );
  SDFFX1 DFF_28_Q_reg ( .D(g7590), .SI(g1077), .SE(n2944), .CLK(n3100), .Q(
        g1231), .QN(n2881) );
  SDFFX1 DFF_29_Q_reg ( .D(g6656), .SI(g1231), .SE(n2976), .CLK(n3084), .Q(g4)
         );
  SDFFX1 DFF_30_Q_reg ( .D(g6728), .SI(g4), .SE(n2976), .CLK(n3084), .Q(g4177)
         );
  SDFFX1 DFF_31_Q_reg ( .D(g5126), .SI(g4177), .SE(n2976), .CLK(n3084), .Q(
        g1104), .QN(n1658) );
  SDFFX1 DFF_32_Q_reg ( .D(g7290), .SI(g1104), .SE(n2979), .CLK(n3082), .Q(
        g1304), .QN(n2756) );
  SDFFX1 DFF_33_Q_reg ( .D(g6841), .SI(g1304), .SE(n2962), .CLK(n3091), .Q(
        g243) );
  SDFFX1 DFF_34_Q_reg ( .D(g8041), .SI(g243), .SE(n2969), .CLK(n3087), .Q(
        g1499), .QN(n2792) );
  SDFFX1 DFF_36_Q_reg ( .D(g8766), .SI(g1499), .SE(n2948), .CLK(n3098), .Q(
        g1444), .QN(n2832) );
  SDFFX1 DFF_37_Q_reg ( .D(n13), .SI(g1444), .SE(n2947), .CLK(n3098), .Q(n3064) );
  SDFFX1 DFF_38_Q_reg ( .D(g8019), .SI(n3064), .SE(n2945), .CLK(n3099), .Q(
        g4180), .QN(n2883) );
  SDFFX1 DFF_39_Q_reg ( .D(g6545), .SI(g4180), .SE(n2940), .CLK(n3102), .Q(
        g1543) );
  SDFFX1 DFF_41_Q_reg ( .D(g256), .SI(g1543), .SE(n2940), .CLK(n3102), .Q(g315), .QN(n2816) );
  SDFFX1 DFF_42_Q_reg ( .D(g6533), .SI(g315), .SE(n2939), .CLK(n3102), .Q(
        g1534) );
  SDFFX1 DFF_43_Q_reg ( .D(g8820), .SI(g1534), .SE(n2939), .CLK(n3102), .Q(
        g622), .QN(n1713) );
  SDFFX1 DFF_44_Q_reg ( .D(g8941), .SI(g622), .SE(n2972), .CLK(n3085), .Q(
        g1927) );
  SDFFX1 DFF_45_Q_reg ( .D(g10859), .SI(g1927), .SE(n2919), .CLK(n3112), .Q(
        g1660) );
  SDFFX1 DFF_46_Q_reg ( .D(g6922), .SI(g1660), .SE(n2970), .CLK(n3087), .Q(
        g278) );
  SDFFX1 DFF_47_Q_reg ( .D(g8772), .SI(g278), .SE(n2970), .CLK(n3087), .Q(
        g1436), .QN(n2829) );
  SDFFX1 DFF_48_Q_reg ( .D(g8433), .SI(g1436), .SE(n2926), .CLK(n3109), .Q(
        g718), .QN(n2696) );
  SDFFX1 DFF_49_Q_reg ( .D(g6526), .SI(g718), .SE(n2925), .CLK(n3109), .Q(
        g8985) );
  SDFFX1 DFF_50_Q_reg ( .D(g10793), .SI(g8985), .SE(n2919), .CLK(n3112), .Q(
        g554) );
  SDFFX1 DFF_51_Q_reg ( .D(g11333), .SI(g554), .SE(n2919), .CLK(n3112), .Q(
        g496), .QN(n1689) );
  SDFFX1 DFF_52_Q_reg ( .D(g11392), .SI(g496), .SE(n2984), .CLK(n3080), .Q(
        g981), .QN(n1720) );
  SDFFX1 DFF_53_Q_reg ( .D(n2896), .SI(g981), .SE(n2984), .CLK(n3079), .Q(
        g3007) );
  SDFFX1 DFF_54_Q_reg ( .D(g1713), .SI(g3007), .SE(n2964), .CLK(n3089), .Q(
        test_so1) );
  SDFFX1 DFF_55_Q_reg ( .D(g794), .SI(test_si2), .SE(n2982), .CLK(n3080), .Q(
        g829) );
  SDFFX1 DFF_56_Q_reg ( .D(g6093), .SI(g829), .SE(n2918), .CLK(n3112), .Q(
        g1095) );
  SDFFX1 DFF_57_Q_reg ( .D(g8889), .SI(g1095), .SE(n2911), .CLK(n3116), .Q(
        g704), .QN(n2796) );
  SDFFX1 DFF_58_Q_reg ( .D(g7302), .SI(g704), .SE(n2979), .CLK(n3082), .Q(
        g1265), .QN(n2752) );
  SDFFX1 DFF_59_Q_reg ( .D(g6525), .SI(g1265), .SE(n2943), .CLK(n3100), .Q(
        g1786), .QN(n2853) );
  SDFFX1 DFF_60_Q_reg ( .D(g8429), .SI(g1786), .SE(n2954), .CLK(n3094), .Q(
        g682), .QN(n2864) );
  SDFFX1 DFF_61_Q_reg ( .D(g7292), .SI(g682), .SE(n2978), .CLK(n3082), .Q(
        g1296), .QN(n2754) );
  SDFFX1 DFF_62_Q_reg ( .D(g104), .SI(g1296), .SE(n2978), .CLK(n3082), .Q(
        g2602) );
  SDFFX1 DFF_63_Q_reg ( .D(g6621), .SI(g2602), .SE(n2950), .CLK(n3097), .Q(
        g8977) );
  SDFFX1 DFF_64_Q_reg ( .D(g7134), .SI(g8977), .SE(n2938), .CLK(n3102), .Q(
        n3062), .QN(n5133) );
  SDFFX1 DFF_65_Q_reg ( .D(g260), .SI(n3062), .SE(n2938), .CLK(n3102), .Q(g327), .QN(n2782) );
  SDFFX1 DFF_66_Q_reg ( .D(g6333), .SI(g327), .SE(n2938), .CLK(n3102), .Q(
        g1389) );
  SDFFX1 DFF_67_Q_reg ( .D(g6826), .SI(g1389), .SE(n2938), .CLK(n3103), .Q(
        g1371) );
  SDFFX1 DFF_68_Q_reg ( .D(g1955), .SI(g1371), .SE(n2936), .CLK(n3104), .Q(
        g1956) );
  SDFFX1 DFF_69_Q_reg ( .D(g10860), .SI(g1956), .SE(n2919), .CLK(n3112), .Q(
        g1675) );
  SDFFX1 DFF_70_Q_reg ( .D(g11483), .SI(g1675), .SE(n2957), .CLK(n3093), .Q(
        g354) );
  SDFFX1 DFF_71_Q_reg ( .D(g6392), .SI(g354), .SE(n2957), .CLK(n3093), .Q(g113) );
  SDFFX1 DFF_72_Q_reg ( .D(g7626), .SI(g113), .SE(n2956), .CLK(n3093), .Q(g639), .QN(n1692) );
  SDFFX1 DFF_73_Q_reg ( .D(g10866), .SI(g639), .SE(n2932), .CLK(n3105), .Q(
        g1684) );
  SDFFX1 DFF_74_Q_reg ( .D(g8193), .SI(g1684), .SE(n2932), .CLK(n3106), .Q(
        g1639) );
  SDFFX1 DFF_75_Q_reg ( .D(g6983), .SI(g1639), .SE(n2932), .CLK(n3106), .Q(
        g1791), .QN(n1702) );
  SDFFX1 DFF_76_Q_reg ( .D(g6839), .SI(g1791), .SE(n2927), .CLK(n3108), .Q(
        g248) );
  SDFFX1 DFF_77_Q_reg ( .D(g4076), .SI(g248), .SE(n2927), .CLK(n3108), .Q(
        g1707), .QN(n2848) );
  SDFFX1 DFF_78_Q_reg ( .D(g4293), .SI(g1707), .SE(n2920), .CLK(n3111), .Q(
        g1759) );
  SDFFX1 DFF_79_Q_reg ( .D(g11482), .SI(g1759), .SE(n2952), .CLK(n3096), .Q(
        g351) );
  SDFFX1 DFF_80_Q_reg ( .D(g1956), .SI(g351), .SE(n2951), .CLK(n3096), .Q(
        g1957) );
  SDFFX1 DFF_81_Q_reg ( .D(g6507), .SI(g1957), .SE(n2951), .CLK(n3096), .Q(
        g1604) );
  SDFFX1 DFF_82_Q_reg ( .D(g6096), .SI(g1604), .SE(n2951), .CLK(n3096), .Q(
        g1098) );
  SDFFX1 DFF_83_Q_reg ( .D(g8250), .SI(g1098), .SE(n2923), .CLK(n3110), .Q(
        g932) );
  SDFFX1 DFF_85_Q_reg ( .D(g8282), .SI(g932), .SE(n2917), .CLK(n3113), .Q(
        g1896) );
  SDFFX1 DFF_86_Q_reg ( .D(g8435), .SI(g1896), .SE(n2955), .CLK(n3094), .Q(
        g736), .QN(n2808) );
  SDFFX1 DFF_87_Q_reg ( .D(g6924), .SI(g736), .SE(n2951), .CLK(n3096), .Q(
        g1019), .QN(n2742) );
  SDFFX1 DFF_88_Q_reg ( .D(g6819), .SI(g1019), .SE(n2951), .CLK(n3096), .Q(
        n3061), .QN(n5137) );
  SDFFX1 DFF_89_Q_reg ( .D(g746), .SI(n3061), .SE(n2950), .CLK(n3096), .Q(g745), .QN(n2649) );
  SDFFX1 DFF_90_Q_reg ( .D(g6244), .SI(g745), .SE(n2950), .CLK(n3096), .Q(
        g1419), .QN(n1602) );
  SDFFX1 DFF_91_Q_reg ( .D(g6627), .SI(g1419), .SE(n2950), .CLK(n3097), .Q(
        g8979) );
  SDFFX1 DFF_92_Q_reg ( .D(n2895), .SI(g8979), .SE(n2949), .CLK(n3097), .Q(g32) );
  SDFFX1 DFF_93_Q_reg ( .D(g3007), .SI(g32), .SE(n2949), .CLK(n3097), .Q(n1865), .QN(n5139) );
  SDFFX1 DFF_94_Q_reg ( .D(g6071), .SI(n1865), .SE(n2911), .CLK(n3116), .Q(
        g1086) );
  SDFFX1 DFF_95_Q_reg ( .D(g8046), .SI(g1086), .SE(n2975), .CLK(n3084), .Q(
        g1486), .QN(n2765) );
  SDFFX1 DFF_96_Q_reg ( .D(g10707), .SI(g1486), .SE(n2941), .CLK(n3101), .Q(
        g1730) );
  SDFFX1 DFF_97_Q_reg ( .D(g6198), .SI(g1730), .SE(n2941), .CLK(n3101), .Q(
        g1504) );
  SDFFX1 DFF_98_Q_reg ( .D(g8051), .SI(g1504), .SE(n2963), .CLK(n3090), .Q(
        g1470), .QN(n2803) );
  SDFFX1 DFF_99_Q_reg ( .D(g8024), .SI(g1470), .SE(n2963), .CLK(n3090), .Q(
        g822), .QN(n2855) );
  SDFFX1 DFF_100_Q_reg ( .D(g29), .SI(g822), .SE(n2962), .CLK(n3090), .Q(g2609) );
  SDFFX1 DFF_101_Q_reg ( .D(g10862), .SI(g2609), .SE(n2921), .CLK(n3111), .Q(
        g1678) );
  SDFFX1 DFF_102_Q_reg ( .D(g8050), .SI(g1678), .SE(n2915), .CLK(n3114), .Q(
        g174), .QN(n2842) );
  SDFFX1 DFF_103_Q_reg ( .D(g7133), .SI(g174), .SE(n2964), .CLK(n3089), .Q(
        g1766), .QN(n2860) );
  SDFFX1 DFF_104_Q_reg ( .D(g7930), .SI(g1766), .SE(n2931), .CLK(n3106), .Q(
        g1801), .QN(n2840) );
  SDFFX1 DFF_105_Q_reg ( .D(g6832), .SI(g1801), .SE(n2931), .CLK(n3106), .Q(
        g186) );
  SDFFX1 DFF_106_Q_reg ( .D(g11308), .SI(g186), .SE(n2910), .CLK(n3116), .Q(
        g959) );
  SDFFX1 DFF_108_Q_reg ( .D(g6918), .SI(g959), .SE(n2910), .CLK(n3117), .Q(
        test_so2) );
  SDFFX1 DFF_109_Q_reg ( .D(g8769), .SI(test_si3), .SE(n2930), .CLK(n3107), 
        .Q(g1407) );
  SDFFX1 DFF_111_Q_reg ( .D(g6909), .SI(g1407), .SE(n2946), .CLK(n3098), .Q(
        g1868) );
  SDFFX1 DFF_112_Q_reg ( .D(g4940), .SI(g1868), .SE(n2946), .CLK(n3098), .Q(
        g4173), .QN(n2871) );
  SDFFX1 DFF_113_Q_reg ( .D(g5404), .SI(g4173), .SE(n2941), .CLK(n3101), .Q(
        g1718), .QN(n1611) );
  SDFFX1 DFF_114_Q_reg ( .D(g11265), .SI(g1718), .SE(n2986), .CLK(n3078), .Q(
        g396), .QN(n2779) );
  SDFFX1 DFF_115_Q_reg ( .D(g6930), .SI(g396), .SE(n2913), .CLK(n3115), .Q(
        g1015), .QN(n2741) );
  SDFFX1 DFF_116_Q_reg ( .D(g10726), .SI(g1015), .SE(n2913), .CLK(n3115), .Q(
        n1650) );
  SDFFX1 DFF_117_Q_reg ( .D(g4891), .SI(n1650), .SE(n2989), .CLK(n3077), .Q(
        n3059), .QN(n1874) );
  SDFFX1 DFF_118_Q_reg ( .D(g6224), .SI(n3059), .SE(n2916), .CLK(n3113), .Q(
        g1415), .QN(n2657) );
  SDFFX1 DFF_119_Q_reg ( .D(g7586), .SI(g1415), .SE(n2993), .CLK(n3075), .Q(
        g1227), .QN(n2650) );
  SDFFX1 DFF_120_Q_reg ( .D(g10770), .SI(g1227), .SE(n2993), .CLK(n3075), .Q(
        g1721) );
  SDFFX1 DFF_121_Q_reg ( .D(g2986), .SI(g1721), .SE(n2925), .CLK(n3109), .Q(
        n3058) );
  SDFFX1 DFF_122_Q_reg ( .D(n2902), .SI(n3058), .SE(n2917), .CLK(n3113), .Q(
        n3057) );
  SDFFX1 DFF_123_Q_reg ( .D(g6934), .SI(n3057), .SE(n2909), .CLK(n3117), .Q(
        g284) );
  SDFFX1 DFF_124_Q_reg ( .D(g11256), .SI(g284), .SE(n2987), .CLK(n3078), .Q(
        g426), .QN(n2815) );
  SDFFX1 DFF_125_Q_reg ( .D(g6824), .SI(g426), .SE(n2938), .CLK(n3103), .Q(
        g219), .QN(n2880) );
  SDFFX1 DFF_126_Q_reg ( .D(g1360), .SI(g219), .SE(n2937), .CLK(n3103), .Q(
        n3056), .QN(n2907) );
  SDFFX1 DFF_127_Q_reg ( .D(g6126), .SI(n3056), .SE(n2937), .CLK(n3103), .Q(
        g806), .QN(n2859) );
  SDFFX1 DFF_128_Q_reg ( .D(g8767), .SI(g806), .SE(n2937), .CLK(n3103), .Q(
        g1428), .QN(n2831) );
  SDFFX1 DFF_129_Q_reg ( .D(g102), .SI(g1428), .SE(n2937), .CLK(n3103), .Q(
        g2605) );
  SDFFX1 DFF_130_Q_reg ( .D(g6546), .SI(g2605), .SE(n2909), .CLK(n3117), .Q(
        g1564) );
  SDFFX1 DFF_131_Q_reg ( .D(g4238), .SI(g1564), .SE(n2909), .CLK(n3117), .Q(
        g1741) );
  SDFFX1 DFF_132_Q_reg ( .D(g6823), .SI(g1741), .SE(n2991), .CLK(n3076), .Q(
        g225), .QN(n2877) );
  SDFFX1 DFF_133_Q_reg ( .D(g6928), .SI(g225), .SE(n2915), .CLK(n3114), .Q(
        g281) );
  SDFFX1 DFF_134_Q_reg ( .D(g11602), .SI(g281), .SE(n2914), .CLK(n3114), .Q(
        g1308) );
  SDFFX1 DFF_135_Q_reg ( .D(g9721), .SI(g1308), .SE(n2955), .CLK(n3094), .Q(
        g611), .QN(n1609) );
  SDFFX1 DFF_136_Q_reg ( .D(g4890), .SI(g611), .SE(n2989), .CLK(n3077), .Q(
        n3055) );
  SDFFX1 DFF_137_Q_reg ( .D(n1586), .SI(n3055), .SE(n2989), .CLK(n3077), .Q(
        g1217) );
  SDFFX1 DFF_138_Q_reg ( .D(g6524), .SI(g1217), .SE(n2937), .CLK(n3103), .Q(
        g1589) );
  SDFFX1 DFF_139_Q_reg ( .D(g8045), .SI(g1589), .SE(n2947), .CLK(n3098), .Q(
        g1466), .QN(n2769) );
  SDFFX1 DFF_140_Q_reg ( .D(g6469), .SI(g1466), .SE(n2947), .CLK(n3098), .Q(
        g1571) );
  SDFFX1 DFF_141_Q_reg ( .D(g6471), .SI(g1571), .SE(n2947), .CLK(n3098), .Q(
        g1861), .QN(n2839) );
  SDFFX1 DFF_142_Q_reg ( .D(g6821), .SI(g1861), .SE(n2947), .CLK(n3098), .Q(
        n3054), .QN(n5136) );
  SDFFX1 DFF_143_Q_reg ( .D(g11514), .SI(n3054), .SE(n2957), .CLK(n3093), .Q(
        g1448), .QN(n2771) );
  SDFFX1 DFF_145_Q_reg ( .D(n187), .SI(g1448), .SE(n2957), .CLK(n3093), .Q(
        g1133), .QN(n1706) );
  SDFFX1 DFF_146_Q_reg ( .D(g11610), .SI(g1133), .SE(n2993), .CLK(n3075), .Q(
        g1333) );
  SDFFX1 DFF_147_Q_reg ( .D(g7843), .SI(g1333), .SE(n2974), .CLK(n3085), .Q(
        g153), .QN(n2789) );
  SDFFX1 DFF_148_Q_reg ( .D(g11310), .SI(g153), .SE(n2952), .CLK(n3095), .Q(
        g962) );
  SDFFX1 DFF_149_Q_reg ( .D(g5536), .SI(g962), .SE(n2952), .CLK(n3095), .Q(
        g4175) );
  SDFFX1 DFF_150_Q_reg ( .D(g28), .SI(g4175), .SE(n2952), .CLK(n3095), .Q(
        g2603) );
  SDFFX1 DFF_151_Q_reg ( .D(g11331), .SI(g2603), .SE(n2952), .CLK(n3096), .Q(
        g486), .QN(n1621) );
  SDFFX1 DFF_152_Q_reg ( .D(g11380), .SI(g486), .SE(n2928), .CLK(n3108), .Q(
        g471), .QN(n1606) );
  SDFFX1 DFF_153_Q_reg ( .D(g6838), .SI(g471), .SE(n2927), .CLK(n3108), .Q(
        g1397) );
  SDFFX1 DFF_154_Q_reg ( .D(g103), .SI(g1397), .SE(n2927), .CLK(n3108), .Q(
        g2606) );
  SDFFX1 DFF_155_Q_reg ( .D(g8288), .SI(g2606), .SE(n2973), .CLK(n3085), .Q(
        g1950), .QN(n2810) );
  SDFFX1 DFF_156_Q_reg ( .D(g755), .SI(g1950), .SE(n2968), .CLK(n3088), .Q(
        g756) );
  SDFFX1 DFF_157_Q_reg ( .D(n160), .SI(g756), .SE(n2989), .CLK(n3077), .Q(
        n3053) );
  SDFFX1 DFF_159_Q_reg ( .D(g10855), .SI(g1101), .SE(n2941), .CLK(n3101), .Q(
        g549) );
  SDFFX1 DFF_161_Q_reg ( .D(g10898), .SI(g549), .SE(n2991), .CLK(n3076), .Q(
        g105), .QN(n2893) );
  SDFFX1 DFF_162_Q_reg ( .D(g10865), .SI(g105), .SE(n2991), .CLK(n3076), .Q(
        g1669) );
  SDFFX1 DFF_163_Q_reg ( .D(g6822), .SI(g1669), .SE(n2991), .CLK(n3076), .Q(
        test_so3) );
  SDFFX1 DFF_164_Q_reg ( .D(g6528), .SI(test_si4), .SE(n2940), .CLK(n3102), 
        .Q(g1531) );
  SDFFX1 DFF_165_Q_reg ( .D(g6180), .SI(g1531), .SE(n2969), .CLK(n3087), .Q(
        g1458), .QN(n1703) );
  SDFFX1 DFF_166_Q_reg ( .D(g10718), .SI(g1458), .SE(n2941), .CLK(n3101), .Q(
        g572) );
  SDFFX1 DFF_167_Q_reg ( .D(g6912), .SI(g572), .SE(n2959), .CLK(n3092), .Q(
        g1011), .QN(n2776) );
  SDFFX1 DFF_168_Q_reg ( .D(g10719), .SI(g1011), .SE(n2958), .CLK(n3092), .Q(
        n3051) );
  SDFFX1 DFF_169_Q_reg ( .D(g6234), .SI(n3051), .SE(n2958), .CLK(n3092), .Q(
        g1411) );
  SDFFX1 DFF_170_Q_reg ( .D(g6099), .SI(g1411), .SE(n2914), .CLK(n3115), .Q(
        g1074) );
  SDFFX1 DFF_171_Q_reg ( .D(g11259), .SI(g1074), .SE(n2985), .CLK(n3079), .Q(
        g444) );
  SDFFX1 DFF_172_Q_reg ( .D(g8039), .SI(g444), .SE(n2991), .CLK(n3076), .Q(
        g1474), .QN(n2802) );
  SDFFX1 DFF_173_Q_reg ( .D(g6059), .SI(g1474), .SE(n2965), .CLK(n3089), .Q(
        g1080) );
  SDFFX1 DFF_174_Q_reg ( .D(g5396), .SI(g1080), .SE(n2965), .CLK(n3089), .Q(
        g1713), .QN(n1610) );
  SDFFX1 DFF_175_Q_reg ( .D(g262), .SI(g1713), .SE(n2933), .CLK(n3105), .Q(
        g333), .QN(n2799) );
  SDFFX1 DFF_176_Q_reg ( .D(g6906), .SI(g333), .SE(n2924), .CLK(n3110), .Q(
        g269) );
  SDFFX1 DFF_177_Q_reg ( .D(g11266), .SI(g269), .SE(n2986), .CLK(n3078), .Q(
        g401), .QN(n2783) );
  SDFFX1 DFF_178_Q_reg ( .D(g11294), .SI(g401), .SE(n2968), .CLK(n3087), .Q(
        g1857), .QN(n1682) );
  SDFFX1 DFF_179_Q_reg ( .D(g5421), .SI(g1857), .SE(n2968), .CLK(n3087), .Q(g9) );
  SDFFX1 DFF_180_Q_reg ( .D(g8649), .SI(g9), .SE(n2954), .CLK(n3094), .Q(g664), 
        .QN(n2856) );
  SDFFX1 DFF_181_Q_reg ( .D(g11312), .SI(g664), .SE(n2962), .CLK(n3090), .Q(
        g965) );
  SDFFX1 DFF_182_Q_reg ( .D(g6840), .SI(g965), .SE(n2962), .CLK(n3091), .Q(
        g1400) );
  SDFFX1 DFF_183_Q_reg ( .D(g254), .SI(g1400), .SE(n2953), .CLK(n3095), .Q(
        g309), .QN(n2606) );
  SDFFX1 DFF_184_Q_reg ( .D(g7202), .SI(g309), .SE(n2953), .CLK(n3095), .Q(
        g814), .QN(n2858) );
  SDFFX1 DFF_185_Q_reg ( .D(g6834), .SI(g814), .SE(n2946), .CLK(n3098), .Q(
        g231), .QN(n2879) );
  SDFFX1 DFF_186_Q_reg ( .D(g10795), .SI(g231), .SE(n2929), .CLK(n3107), .Q(
        g557) );
  SDFFX1 DFF_187_Q_reg ( .D(g103), .SI(g557), .SE(n2929), .CLK(n3107), .Q(
        g2612) );
  SDFFX1 DFF_188_Q_reg ( .D(g875), .SI(g2612), .SE(n2928), .CLK(n3107), .Q(
        g869) );
  SDFFX1 DFF_189_Q_reg ( .D(g6831), .SI(g869), .SE(n2928), .CLK(n3107), .Q(
        g1383) );
  SDFFX1 DFF_190_Q_reg ( .D(g8060), .SI(g1383), .SE(n2922), .CLK(n3111), .Q(
        g158), .QN(n2768) );
  SDFFX1 DFF_191_Q_reg ( .D(g4893), .SI(g158), .SE(n2990), .CLK(n3077), .Q(
        g627) );
  SDFFX1 DFF_192_Q_reg ( .D(g7244), .SI(g627), .SE(n2918), .CLK(n3113), .Q(
        g1023), .QN(n2721) );
  SDFFX1 DFF_193_Q_reg ( .D(g6026), .SI(g1023), .SE(n2915), .CLK(n3114), .Q(
        g259) );
  SDFFX1 DFF_194_Q_reg ( .D(g3069), .SI(g259), .SE(n2915), .CLK(n3114), .Q(
        n3050) );
  SDFFX1 DFF_195_Q_reg ( .D(g11608), .SI(n3050), .SE(n2915), .CLK(n3114), .Q(
        g1327) );
  SDFFX1 DFF_196_Q_reg ( .D(g7660), .SI(g1327), .SE(n2955), .CLK(n3094), .Q(
        g654), .QN(n2836) );
  SDFFX1 DFF_197_Q_reg ( .D(g6911), .SI(g654), .SE(n2912), .CLK(n3116), .Q(
        g293) );
  SDFFX1 DFF_198_Q_reg ( .D(g11640), .SI(g293), .SE(n2963), .CLK(n3090), .Q(
        g1346), .QN(n2820) );
  SDFFX1 DFF_199_Q_reg ( .D(g8777), .SI(g1346), .SE(n2963), .CLK(n3090), .Q(
        g1633) );
  SDFFX1 DFF_200_Q_reg ( .D(g4274), .SI(g1633), .SE(n2932), .CLK(n3106), .Q(
        g1753) );
  SDFFX1 DFF_201_Q_reg ( .D(n2898), .SI(g1753), .SE(n2931), .CLK(n3106), .Q(
        g1508), .QN(n1707) );
  SDFFX1 DFF_202_Q_reg ( .D(g7297), .SI(g1508), .SE(n2980), .CLK(n3081), .Q(
        g1240), .QN(n2813) );
  SDFFX1 DFF_203_Q_reg ( .D(g11326), .SI(g1240), .SE(n2923), .CLK(n3110), .Q(
        g538), .QN(n2806) );
  SDFFX1 DFF_204_Q_reg ( .D(g11269), .SI(g538), .SE(n2986), .CLK(n3079), .Q(
        g416), .QN(n2757) );
  SDFFX1 DFF_205_Q_reg ( .D(g11325), .SI(g416), .SE(n2924), .CLK(n3110), .Q(
        g542), .QN(n2807) );
  SDFFX1 DFF_206_Q_reg ( .D(g10864), .SI(g542), .SE(n2923), .CLK(n3110), .Q(
        g1681) );
  SDFFX1 DFF_207_Q_reg ( .D(g11290), .SI(g1681), .SE(n2916), .CLK(n3114), .Q(
        g374), .QN(n2740) );
  SDFFX1 DFF_208_Q_reg ( .D(g10798), .SI(g374), .SE(n2915), .CLK(n3114), .Q(
        g563) );
  SDFFX1 DFF_209_Q_reg ( .D(g8284), .SI(g563), .SE(n2914), .CLK(n3114), .Q(
        g1914), .QN(n2745) );
  SDFFX1 DFF_210_Q_reg ( .D(g11328), .SI(g1914), .SE(n2954), .CLK(n3095), .Q(
        g530), .QN(n2804) );
  SDFFX1 DFF_211_Q_reg ( .D(g10800), .SI(g530), .SE(n2953), .CLK(n3095), .Q(
        g575) );
  SDFFX1 DFF_212_Q_reg ( .D(g8944), .SI(g575), .SE(n2971), .CLK(n3086), .Q(
        g1936), .QN(n1694) );
  SDFFX1 DFF_213_Q_reg ( .D(g7183), .SI(g1936), .SE(n2949), .CLK(n3097), .Q(
        g8978) );
  SDFFX1 DFF_214_Q_reg ( .D(g4465), .SI(g8978), .SE(n2948), .CLK(n3097), .Q(
        test_so4), .QN(n2906) );
  SDFFX1 DFF_215_Q_reg ( .D(g1356), .SI(test_si5), .SE(n2983), .CLK(n3080), 
        .Q(g1317), .QN(n2889) );
  SDFFX1 DFF_216_Q_reg ( .D(g11484), .SI(g1317), .SE(n2949), .CLK(n3097), .Q(
        g357) );
  SDFFX1 DFF_217_Q_reg ( .D(g11263), .SI(g357), .SE(n2987), .CLK(n3078), .Q(
        g386), .QN(n2781) );
  SDFFX1 DFF_218_Q_reg ( .D(g6501), .SI(g386), .SE(n2934), .CLK(n3104), .Q(
        g1601) );
  SDFFX1 DFF_220_Q_reg ( .D(g6757), .SI(g1601), .SE(n2934), .CLK(n3105), .Q(
        g166), .QN(n2766) );
  SDFFX1 DFF_221_Q_reg ( .D(g11334), .SI(g166), .SE(n2934), .CLK(n3105), .Q(
        g501), .QN(n1690) );
  SDFFX1 DFF_222_Q_reg ( .D(g6042), .SI(g501), .SE(n2934), .CLK(n3105), .Q(
        g262) );
  SDFFX1 DFF_223_Q_reg ( .D(g8384), .SI(g262), .SE(n2918), .CLK(n3113), .Q(
        g1840), .QN(n2809) );
  SDFFX1 DFF_224_Q_reg ( .D(g6653), .SI(g1840), .SE(n2918), .CLK(n3113), .Q(
        g8983) );
  SDFFX1 DFF_225_Q_reg ( .D(g257), .SI(g8983), .SE(n2917), .CLK(n3113), .Q(
        g318), .QN(n2780) );
  SDFFX1 DFF_226_Q_reg ( .D(g5763), .SI(g318), .SE(n2983), .CLK(n3080), .Q(
        g1356) );
  SDFFX1 DFF_227_Q_reg ( .D(g5849), .SI(g1356), .SE(n2982), .CLK(n3080), .Q(
        g794), .QN(n2866) );
  SDFFX1 DFF_228_Q_reg ( .D(g10722), .SI(g794), .SE(n2982), .CLK(n3080), .Q(
        n3048) );
  SDFFX1 DFF_229_Q_reg ( .D(g6929), .SI(n3048), .SE(n2924), .CLK(n3110), .Q(
        g302) );
  SDFFX1 DFF_230_Q_reg ( .D(g11488), .SI(g302), .SE(n2914), .CLK(n3115), .Q(
        g342) );
  SDFFX1 DFF_231_Q_reg ( .D(g7299), .SI(g342), .SE(n2980), .CLK(n3082), .Q(
        g1250), .QN(n2777) );
  SDFFX1 DFF_232_Q_reg ( .D(g4330), .SI(g1250), .SE(n2979), .CLK(n3082), .Q(
        g1163), .QN(n2786) );
  SDFFX1 DFF_233_Q_reg ( .D(g1958), .SI(g1163), .SE(n2960), .CLK(n3092), .Q(
        n3047), .QN(g5816) );
  SDFFX1 DFF_234_Q_reg ( .D(g7257), .SI(n3047), .SE(n2993), .CLK(n3075), .Q(
        g1032), .QN(n2888) );
  SDFFX1 DFF_235_Q_reg ( .D(g8775), .SI(g1032), .SE(n2988), .CLK(n3077), .Q(
        g1432), .QN(n2772) );
  SDFFX1 DFF_237_Q_reg ( .D(g5770), .SI(g1432), .SE(n2969), .CLK(n3087), .Q(
        g1453), .QN(n1628) );
  SDFFX1 DFF_238_Q_reg ( .D(g11486), .SI(g1453), .SE(n2933), .CLK(n3105), .Q(
        g363) );
  SDFFX1 DFF_239_Q_reg ( .D(g261), .SI(g363), .SE(n2933), .CLK(n3105), .Q(g330), .QN(n2605) );
  SDFFX1 DFF_240_Q_reg ( .D(g4338), .SI(g330), .SE(n2933), .CLK(n3105), .Q(
        g1157), .QN(n2784) );
  SDFFX1 DFF_241_Q_reg ( .D(g4500), .SI(g1157), .SE(n2932), .CLK(n3105), .Q(
        n3046), .QN(n5141) );
  SDFFX1 DFF_242_Q_reg ( .D(g10721), .SI(n3046), .SE(n2932), .CLK(n3105), .Q(
        n3045) );
  SDFFX1 DFF_243_Q_reg ( .D(g8147), .SI(n3045), .SE(n2925), .CLK(n3109), .Q(
        g928) );
  SDFFX1 DFF_244_Q_reg ( .D(g6038), .SI(g928), .SE(n2925), .CLK(n3109), .Q(
        g261) );
  SDFFX1 DFF_245_Q_reg ( .D(g11337), .SI(g261), .SE(n2925), .CLK(n3109), .Q(
        g516), .QN(n1620) );
  SDFFX1 DFF_246_Q_reg ( .D(g6045), .SI(g516), .SE(n2953), .CLK(n3095), .Q(
        g254) );
  SDFFX1 DFF_247_Q_reg ( .D(g7191), .SI(g254), .SE(n2946), .CLK(n3099), .Q(
        g4178), .QN(n2869) );
  SDFFX1 DFF_248_Q_reg ( .D(g826), .SI(g4178), .SE(n2911), .CLK(n3116), .Q(
        g861) );
  SDFFX1 DFF_249_Q_reg ( .D(g8774), .SI(g861), .SE(n2910), .CLK(n3116), .Q(
        g1627) );
  SDFFX1 DFF_250_Q_reg ( .D(g7293), .SI(g1627), .SE(n2978), .CLK(n3083), .Q(
        g1292), .QN(n2753) );
  SDFFX1 DFF_251_Q_reg ( .D(g6907), .SI(g1292), .SE(n2978), .CLK(n3083), .Q(
        g290) );
  SDFFX1 DFF_252_Q_reg ( .D(g4903), .SI(g290), .SE(n2978), .CLK(n3083), .Q(
        n3044), .QN(n1873) );
  SDFFX1 DFF_253_Q_reg ( .D(g6123), .SI(n3044), .SE(n2946), .CLK(n3099), .Q(
        g4176), .QN(n2870) );
  SDFFX1 DFF_254_Q_reg ( .D(g6506), .SI(g4176), .SE(n2929), .CLK(n3107), .Q(
        g1583) );
  SDFFX1 DFF_255_Q_reg ( .D(g11376), .SI(g1583), .SE(n2923), .CLK(n3110), .Q(
        g466), .QN(n1646) );
  SDFFX1 DFF_256_Q_reg ( .D(g6542), .SI(g466), .SE(n2969), .CLK(n3087), .Q(
        g1561) );
  SDFFX1 DFF_258_Q_reg ( .D(g6551), .SI(g1561), .SE(n2971), .CLK(n3086), .Q(
        g1546) );
  SDFFX1 DFF_259_Q_reg ( .D(g6901), .SI(g1546), .SE(n2970), .CLK(n3086), .Q(
        g287) );
  SDFFX1 DFF_260_Q_reg ( .D(g10797), .SI(g287), .SE(n2970), .CLK(n3086), .Q(
        g560) );
  SDFFX1 DFF_261_Q_reg ( .D(g8505), .SI(g560), .SE(n2955), .CLK(n3094), .Q(
        g617), .QN(n1645) );
  SDFFX1 DFF_262_Q_reg ( .D(n2900), .SI(g617), .SE(n2955), .CLK(n3094), .Q(
        n1631) );
  SDFFX1 DFF_263_Q_reg ( .D(g11647), .SI(n1631), .SE(n2966), .CLK(n3088), .Q(
        g336) );
  SDFFX1 DFF_264_Q_reg ( .D(g11340), .SI(g336), .SE(n2927), .CLK(n3108), .Q(
        g456), .QN(n1641) );
  SDFFX1 DFF_265_Q_reg ( .D(g253), .SI(g456), .SE(n2926), .CLK(n3108), .Q(g305), .QN(n1681) );
  SDFFX1 DFF_266_Q_reg ( .D(g11625), .SI(g305), .SE(n2909), .CLK(n3117), .Q(
        g345) );
  SDFFX1 DFF_267_Q_reg ( .D(g636), .SI(g345), .SE(n2987), .CLK(n3078), .Q(g8)
         );
  SDFFX1 DFF_268_Q_reg ( .D(g6502), .SI(g8), .SE(n2964), .CLK(n3089), .Q(
        test_so5), .QN(n2904) );
  SDFFX1 DFF_269_Q_reg ( .D(N599), .SI(test_si6), .SE(n2945), .CLK(n3099), .Q(
        g2648) );
  SDFFX1 DFF_270_Q_reg ( .D(g6049), .SI(g2648), .SE(n2935), .CLK(n3104), .Q(
        g255) );
  SDFFX1 DFF_271_Q_reg ( .D(g8945), .SI(g255), .SE(n2971), .CLK(n3086), .Q(
        g1945), .QN(n1697) );
  SDFFX1 DFF_272_Q_reg ( .D(g4231), .SI(g1945), .SE(n2971), .CLK(n3086), .Q(
        g1738) );
  SDFFX1 DFF_273_Q_reg ( .D(g8040), .SI(g1738), .SE(n2971), .CLK(n3086), .Q(
        g1478), .QN(n2835) );
  SDFFX1 DFF_275_Q_reg ( .D(n521), .SI(g1478), .SE(n2971), .CLK(n3086), .Q(
        n3042) );
  SDFFX1 DFF_276_Q_reg ( .D(g6155), .SI(n3042), .SE(n2927), .CLK(n3108), .Q(
        g1690), .QN(n1653) );
  SDFFX1 DFF_277_Q_reg ( .D(g8043), .SI(g1690), .SE(n2976), .CLK(n3083), .Q(
        g1482), .QN(n2770) );
  SDFFX1 DFF_278_Q_reg ( .D(g5173), .SI(g1482), .SE(n2936), .CLK(n3103), .Q(
        g1110), .QN(n1677) );
  SDFFX1 DFF_279_Q_reg ( .D(g6916), .SI(g1110), .SE(n2912), .CLK(n3116), .Q(
        g296) );
  SDFFX1 DFF_280_Q_reg ( .D(g10861), .SI(g296), .SE(n2988), .CLK(n3077), .Q(
        g1663) );
  SDFFX1 DFF_281_Q_reg ( .D(g8431), .SI(g1663), .SE(n2988), .CLK(n3078), .Q(
        g700) );
  SDFFX1 DFF_282_Q_reg ( .D(g4309), .SI(g700), .SE(n2959), .CLK(n3092), .Q(
        g1762) );
  SDFFX1 DFF_283_Q_reg ( .D(g11485), .SI(g1762), .SE(n2959), .CLK(n3092), .Q(
        g360) );
  SDFFX1 DFF_284_Q_reg ( .D(g6334), .SI(g360), .SE(n2936), .CLK(n3104), .Q(
        g192) );
  SDFFX1 DFF_285_Q_reg ( .D(g10767), .SI(g192), .SE(n2990), .CLK(n3076), .Q(
        g1657) );
  SDFFX1 DFF_286_Q_reg ( .D(g8923), .SI(g1657), .SE(n2990), .CLK(n3077), .Q(
        g722), .QN(n1693) );
  SDFFX1 DFF_287_Q_reg ( .D(g7189), .SI(g722), .SE(n2948), .CLK(n3097), .Q(
        g8980) );
  SDFFX1 DFF_288_Q_reg ( .D(g10799), .SI(g8980), .SE(n2975), .CLK(n3084), .Q(
        g566) );
  SDFFX1 DFF_289_Q_reg ( .D(g6747), .SI(g566), .SE(n2992), .CLK(n3076), .Q(
        n3041) );
  SDFFX1 DFF_290_Q_reg ( .D(g6080), .SI(n3041), .SE(n2992), .CLK(n3076), .Q(
        g1089) );
  SDFFX1 DFF_291_Q_reg ( .D(g3381), .SI(g1089), .SE(n2925), .CLK(n3109), .Q(
        g2986), .QN(n2628) );
  SDFFX1 DFF_292_Q_reg ( .D(g5910), .SI(g2986), .SE(n2918), .CLK(n3112), .Q(
        g1071) );
  SDFFX1 DFF_293_Q_reg ( .D(g11393), .SI(g1071), .SE(n2984), .CLK(n3079), .Q(
        g986), .QN(n1722) );
  SDFFX1 DFF_294_Q_reg ( .D(g11349), .SI(g986), .SE(n2984), .CLK(n3080), .Q(
        g971), .QN(n2891) );
  SDFFX1 DFF_295_Q_reg ( .D(g83), .SI(g971), .SE(n2984), .CLK(n3080), .Q(g1955) );
  SDFFX1 DFF_296_Q_reg ( .D(g6439), .SI(g1955), .SE(n2930), .CLK(n3107), .Q(
        g143), .QN(n2790) );
  SDFFX1 DFF_297_Q_reg ( .D(g9266), .SI(g143), .SE(n2945), .CLK(n3099), .Q(
        g1814), .QN(n1608) );
  SDFFX1 DFF_299_Q_reg ( .D(g1217), .SI(g1814), .SE(n2944), .CLK(n3099), .Q(
        g1212), .QN(n2882) );
  SDFFX1 DFF_300_Q_reg ( .D(g8940), .SI(g1212), .SE(n2972), .CLK(n3086), .Q(
        g1918), .QN(n2795) );
  SDFFX1 DFF_301_Q_reg ( .D(g7705), .SI(g1918), .SE(n2945), .CLK(n3099), .Q(
        g4179) );
  SDFFX1 DFF_302_Q_reg ( .D(g9269), .SI(g4179), .SE(n2945), .CLK(n3099), .Q(
        g1822), .QN(n1643) );
  SDFFX1 DFF_303_Q_reg ( .D(g6820), .SI(g1822), .SE(n2951), .CLK(n3096), .Q(
        g237) );
  SDFFX1 DFF_304_Q_reg ( .D(g756), .SI(g237), .SE(n2950), .CLK(n3096), .Q(g746), .QN(n2838) );
  SDFFX1 DFF_306_Q_reg ( .D(g8042), .SI(g746), .SE(n2935), .CLK(n3104), .Q(
        g1462), .QN(n2834) );
  SDFFX1 DFF_307_Q_reg ( .D(g6759), .SI(g1462), .SE(n2930), .CLK(n3106), .Q(
        g178) );
  SDFFX1 DFF_308_Q_reg ( .D(g11487), .SI(g178), .SE(n2923), .CLK(n3110), .Q(
        g366) );
  SDFFX1 DFF_309_Q_reg ( .D(g802), .SI(g366), .SE(n2922), .CLK(n3110), .Q(g837) );
  SDFFX1 DFF_310_Q_reg ( .D(g9124), .SI(g837), .SE(n2939), .CLK(n3102), .Q(
        g599), .QN(n1644) );
  SDFFX1 DFF_311_Q_reg ( .D(g11293), .SI(g599), .SE(n2973), .CLK(n3085), .Q(
        g1854) );
  SDFFX1 DFF_312_Q_reg ( .D(g11298), .SI(g1854), .SE(n2973), .CLK(n3085), .Q(
        g944) );
  SDFFX1 DFF_313_Q_reg ( .D(g8287), .SI(g944), .SE(n2973), .CLK(n3085), .Q(
        g1941), .QN(n2747) );
  SDFFX1 DFF_314_Q_reg ( .D(g8047), .SI(g1941), .SE(n2974), .CLK(n3084), .Q(
        g170), .QN(n2843) );
  SDFFX1 DFF_315_Q_reg ( .D(g6205), .SI(g170), .SE(n2917), .CLK(n3113), .Q(
        g1520), .QN(n1710) );
  SDFFX1 DFF_316_Q_reg ( .D(g8885), .SI(g1520), .SE(n2960), .CLK(n3091), .Q(
        g686), .QN(n1676) );
  SDFFX1 DFF_317_Q_reg ( .D(g11305), .SI(g686), .SE(n2960), .CLK(n3092), .Q(
        g953) );
  SDFFX1 DFF_318_Q_reg ( .D(g5556), .SI(g953), .SE(n2960), .CLK(n3092), .Q(
        g1958) );
  SDFFX1 DFF_319_Q_reg ( .D(g10664), .SI(g1958), .SE(n2959), .CLK(n3092), .Q(
        n3040) );
  SDFFX1 DFF_320_Q_reg ( .D(g2478), .SI(n3040), .SE(n2959), .CLK(n3092), .Q(
        g1765), .QN(n2886) );
  SDFFX1 DFF_321_Q_reg ( .D(g10711), .SI(g1765), .SE(n2940), .CLK(n3101), .Q(
        g1733) );
  SDFFX1 DFF_322_Q_reg ( .D(g7303), .SI(g1733), .SE(n2979), .CLK(n3082), .Q(
        test_so6), .QN(n2905) );
  SDFFX1 DFF_323_Q_reg ( .D(g5194), .SI(test_si7), .SE(n2943), .CLK(n3100), 
        .Q(g1610), .QN(n2885) );
  SDFFX1 DFF_324_Q_reg ( .D(g7541), .SI(g1610), .SE(n2920), .CLK(n3111), .Q(
        g1796), .QN(n1626) );
  SDFFX1 DFF_325_Q_reg ( .D(g11607), .SI(g1796), .SE(n2920), .CLK(n3112), .Q(
        g1324) );
  SDFFX1 DFF_326_Q_reg ( .D(g6541), .SI(g1324), .SE(n2975), .CLK(n3084), .Q(
        g1540) );
  SDFFX1 DFF_327_Q_reg ( .D(g6827), .SI(g1540), .SE(n2938), .CLK(n3103), .Q(
        n3038) );
  SDFFX1 DFF_328_Q_reg ( .D(n2901), .SI(n3038), .SE(n2983), .CLK(n3080), .Q(
        g3069), .QN(n2629) );
  SDFFX1 DFF_329_Q_reg ( .D(g11332), .SI(g3069), .SE(n2952), .CLK(n3096), .Q(
        g491), .QN(n1691) );
  SDFFX1 DFF_330_Q_reg ( .D(g4902), .SI(g491), .SE(n2977), .CLK(n3083), .Q(
        n3037) );
  SDFFX1 DFF_331_Q_reg ( .D(g6828), .SI(n3037), .SE(n2977), .CLK(n3083), .Q(
        g213) );
  SDFFX1 DFF_332_Q_reg ( .D(g6516), .SI(g213), .SE(n2942), .CLK(n3100), .Q(
        g1781), .QN(n1659) );
  SDFFX1 DFF_333_Q_reg ( .D(g8938), .SI(g1781), .SE(n2911), .CLK(n3116), .Q(
        g1900), .QN(n1675) );
  SDFFX1 DFF_334_Q_reg ( .D(g7298), .SI(g1900), .SE(n2980), .CLK(n3082), .Q(
        g1245), .QN(n2774) );
  SDFFX1 DFF_335_Q_reg ( .D(n6), .SI(g1245), .SE(n2980), .CLK(n3082), .Q(n3036), .QN(n5140) );
  SDFFX1 DFF_336_Q_reg ( .D(n178), .SI(n3036), .SE(n2989), .CLK(n3077), .Q(
        n3035) );
  SDFFX1 DFF_337_Q_reg ( .D(g8048), .SI(n3035), .SE(n2930), .CLK(n3106), .Q(
        g148) );
  SDFFX1 DFF_338_Q_reg ( .D(g798), .SI(g148), .SE(n2930), .CLK(n3107), .Q(g833) );
  SDFFX1 DFF_339_Q_reg ( .D(g8285), .SI(g833), .SE(n2972), .CLK(n3086), .Q(
        g1923), .QN(n1718) );
  SDFFX1 DFF_340_Q_reg ( .D(g8254), .SI(g1923), .SE(n2923), .CLK(n3110), .Q(
        g936) );
  SDFFX1 DFF_342_Q_reg ( .D(g11604), .SI(g936), .SE(n2964), .CLK(n3090), .Q(
        g1314) );
  SDFFX1 DFF_343_Q_reg ( .D(g814), .SI(g1314), .SE(n2963), .CLK(n3090), .Q(
        g849) );
  SDFFX1 DFF_344_Q_reg ( .D(g11636), .SI(g849), .SE(n2963), .CLK(n3090), .Q(
        g1336), .QN(n2821) );
  SDFFX1 DFF_345_Q_reg ( .D(g6910), .SI(g1336), .SE(n2974), .CLK(n3085), .Q(
        g272) );
  SDFFX1 DFF_346_Q_reg ( .D(g8173), .SI(g272), .SE(n2974), .CLK(n3085), .Q(
        g1806), .QN(n2841) );
  SDFFX1 DFF_347_Q_reg ( .D(g8245), .SI(g1806), .SE(n2911), .CLK(n3116), .Q(
        g826), .QN(n1716) );
  SDFFX1 DFF_349_Q_reg ( .D(g8281), .SI(g826), .SE(n2973), .CLK(n3085), .Q(
        g1887) );
  SDFFX1 DFF_350_Q_reg ( .D(g10724), .SI(g1887), .SE(n2968), .CLK(n3087), .Q(
        n3034) );
  SDFFX1 DFF_351_Q_reg ( .D(g11314), .SI(n3034), .SE(n2910), .CLK(n3116), .Q(
        g968) );
  SDFFX1 DFF_352_Q_reg ( .D(g4905), .SI(g968), .SE(n2977), .CLK(n3083), .Q(
        n3033), .QN(n5135) );
  SDFFX1 DFF_353_Q_reg ( .D(n352), .SI(n3033), .SE(n2977), .CLK(n3083), .Q(
        g1137), .QN(n1597) );
  SDFFX1 DFF_354_Q_reg ( .D(g8937), .SI(g1137), .SE(n2972), .CLK(n3085), .Q(
        g1891), .QN(n1657) );
  SDFFX1 DFF_355_Q_reg ( .D(g7300), .SI(g1891), .SE(n2979), .CLK(n3082), .Q(
        g1255), .QN(n2749) );
  SDFFX1 DFF_356_Q_reg ( .D(g6002), .SI(g1255), .SE(n2928), .CLK(n3107), .Q(
        g257) );
  SDFFX1 DFF_357_Q_reg ( .D(n1588), .SI(g257), .SE(n2928), .CLK(n3108), .Q(
        g874) );
  SDFFX1 DFF_358_Q_reg ( .D(g9110), .SI(g874), .SE(n2990), .CLK(n3077), .Q(
        g591), .QN(n1607) );
  SDFFX1 DFF_359_Q_reg ( .D(g8926), .SI(g591), .SE(n2987), .CLK(n3078), .Q(
        g731), .QN(n1696) );
  SDFFX1 DFF_360_Q_reg ( .D(g8631), .SI(g731), .SE(n2987), .CLK(n3078), .Q(
        g636) );
  SDFFX1 DFF_361_Q_reg ( .D(g7632), .SI(g636), .SE(n2994), .CLK(n3075), .Q(
        g1218), .QN(n2887) );
  SDFFX1 DFF_362_Q_reg ( .D(g9150), .SI(g1218), .SE(n2939), .CLK(n3102), .Q(
        g605), .QN(n1593) );
  SDFFX1 DFF_363_Q_reg ( .D(g6531), .SI(g605), .SE(n2939), .CLK(n3102), .Q(
        g8986) );
  SDFFX1 DFF_364_Q_reg ( .D(g6786), .SI(g8986), .SE(n2930), .CLK(n3106), .Q(
        g182), .QN(n2788) );
  SDFFX1 DFF_365_Q_reg ( .D(g11303), .SI(g182), .SE(n2922), .CLK(n3110), .Q(
        g950) );
  SDFFX1 DFF_366_Q_reg ( .D(g4477), .SI(g950), .SE(n2922), .CLK(n3110), .Q(
        g1129), .QN(n1705) );
  SDFFX1 DFF_367_Q_reg ( .D(g822), .SI(g1129), .SE(n2962), .CLK(n3090), .Q(
        g857) );
  SDFFX1 DFF_368_Q_reg ( .D(g11258), .SI(g857), .SE(n2985), .CLK(n3079), .Q(
        g448) );
  SDFFX1 DFF_369_Q_reg ( .D(g9272), .SI(g448), .SE(n2944), .CLK(n3100), .Q(
        g1828), .QN(n1605) );
  SDFFX1 DFF_370_Q_reg ( .D(g10773), .SI(g1828), .SE(n2944), .CLK(n3100), .Q(
        g1727) );
  SDFFX1 DFF_371_Q_reg ( .D(g6470), .SI(g1727), .SE(n2943), .CLK(n3100), .Q(
        g1592) );
  SDFFX1 DFF_372_Q_reg ( .D(g5083), .SI(g1592), .SE(n2943), .CLK(n3100), .Q(
        g1703), .QN(n2852) );
  SDFFX1 DFF_373_Q_reg ( .D(g8286), .SI(g1703), .SE(n2909), .CLK(n3117), .Q(
        g1932), .QN(n2748) );
  SDFFX1 DFF_374_Q_reg ( .D(g8773), .SI(g1932), .SE(n2976), .CLK(n3083), .Q(
        g1624) );
  SDFFX1 DFF_376_Q_reg ( .D(g6054), .SI(g1624), .SE(n2966), .CLK(n3088), .Q(
        test_so7) );
  SDFFX1 DFF_377_Q_reg ( .D(g101), .SI(test_si8), .SE(n2994), .CLK(n3075), .Q(
        g2601) );
  SDFFX1 DFF_378_Q_reg ( .D(g11260), .SI(g2601), .SE(n2985), .CLK(n3079), .Q(
        g440) );
  SDFFX1 DFF_379_Q_reg ( .D(g11338), .SI(g440), .SE(n2924), .CLK(n3109), .Q(
        g476), .QN(n1599) );
  SDFFX1 DFF_380_Q_reg ( .D(g5918), .SI(g476), .SE(n2924), .CLK(n3109), .Q(
        g119), .QN(n1613) );
  SDFFX1 DFF_381_Q_reg ( .D(g8922), .SI(g119), .SE(n2913), .CLK(n3115), .Q(
        g668), .QN(n1662) );
  SDFFX1 DFF_382_Q_reg ( .D(g8049), .SI(g668), .SE(n2913), .CLK(n3115), .Q(
        g139), .QN(n2763) );
  SDFFX1 DFF_383_Q_reg ( .D(g4342), .SI(g139), .SE(n2913), .CLK(n3115), .Q(
        g1149), .QN(n1685) );
  SDFFX1 DFF_384_Q_reg ( .D(g10720), .SI(g1149), .SE(n2912), .CLK(n3115), .Q(
        n3031) );
  SDFFX1 DFF_385_Q_reg ( .D(g6755), .SI(n3031), .SE(n2977), .CLK(n3083), .Q(
        n3030) );
  SDFFX1 DFF_386_Q_reg ( .D(g6897), .SI(n3030), .SE(n2924), .CLK(n3109), .Q(
        g263) );
  SDFFX1 DFF_387_Q_reg ( .D(g7709), .SI(g263), .SE(n2953), .CLK(n3095), .Q(
        g818), .QN(n2846) );
  SDFFX1 DFF_388_Q_reg ( .D(g4255), .SI(g818), .SE(n2914), .CLK(n3115), .Q(
        g1747) );
  SDFFX1 DFF_389_Q_reg ( .D(g5543), .SI(g1747), .SE(n2982), .CLK(n3081), .Q(
        g802), .QN(n1622) );
  SDFFX1 DFF_390_Q_reg ( .D(g6915), .SI(g802), .SE(n2922), .CLK(n3111), .Q(
        g275) );
  SDFFX1 DFF_391_Q_reg ( .D(g6513), .SI(g275), .SE(n2922), .CLK(n3111), .Q(
        g1524) );
  SDFFX1 DFF_392_Q_reg ( .D(g6480), .SI(g1524), .SE(n2921), .CLK(n3111), .Q(
        g1577) );
  SDFFX1 DFF_393_Q_reg ( .D(g6733), .SI(g1577), .SE(n2982), .CLK(n3081), .Q(
        g810), .QN(n2847) );
  SDFFX1 DFF_394_Q_reg ( .D(g11264), .SI(g810), .SE(n2986), .CLK(n3078), .Q(
        g391), .QN(n2817) );
  SDFFX1 DFF_395_Q_reg ( .D(g8973), .SI(g391), .SE(n2956), .CLK(n3093), .Q(
        g658), .QN(n1615) );
  SDFFX1 DFF_396_Q_reg ( .D(g6833), .SI(g658), .SE(n2956), .CLK(n3093), .Q(
        g1386) );
  SDFFX1 DFF_397_Q_reg ( .D(g5996), .SI(g1386), .SE(n2931), .CLK(n3106), .Q(
        g253) );
  SDFFX1 DFF_398_Q_reg ( .D(n1587), .SI(g253), .SE(n2931), .CLK(n3106), .Q(
        g875) );
  SDFFX1 DFF_399_Q_reg ( .D(g4473), .SI(g875), .SE(n2931), .CLK(n3106), .Q(
        g1125), .QN(n1708) );
  SDFFX1 DFF_400_Q_reg ( .D(g5755), .SI(g1125), .SE(n2956), .CLK(n3094), .Q(
        g201), .QN(n1619) );
  SDFFX1 DFF_401_Q_reg ( .D(g7295), .SI(g201), .SE(n2956), .CLK(n3094), .Q(
        g1280), .QN(n1862) );
  SDFFX1 DFF_402_Q_reg ( .D(g6068), .SI(g1280), .SE(n2956), .CLK(n3094), .Q(
        g1083) );
  SDFFX1 DFF_403_Q_reg ( .D(g7137), .SI(g1083), .SE(n2955), .CLK(n3094), .Q(
        g650), .QN(n1709) );
  SDFFX1 DFF_404_Q_reg ( .D(g8779), .SI(g650), .SE(n2947), .CLK(n3098), .Q(
        g1636) );
  SDFFX1 DFF_405_Q_reg ( .D(g818), .SI(g1636), .SE(n2953), .CLK(n3095), .Q(
        g853) );
  SDFFX1 DFF_406_Q_reg ( .D(g11270), .SI(g853), .SE(n2985), .CLK(n3079), .Q(
        g421), .QN(n2798) );
  SDFFX1 DFF_407_Q_reg ( .D(g5529), .SI(g421), .SE(n2946), .CLK(n3099), .Q(
        g4174), .QN(n2872) );
  SDFFX1 DFF_408_Q_reg ( .D(g11306), .SI(g4174), .SE(n2981), .CLK(n3081), .Q(
        g956) );
  SDFFX1 DFF_409_Q_reg ( .D(g11291), .SI(g956), .SE(n2981), .CLK(n3081), .Q(
        g378), .QN(n2739) );
  SDFFX1 DFF_410_Q_reg ( .D(g4283), .SI(g378), .SE(n2920), .CLK(n3112), .Q(
        g1756) );
  SDFFX1 DFF_411_Q_reg ( .D(g29), .SI(g1756), .SE(n2920), .CLK(n3112), .Q(
        g2604) );
  SDFFX1 DFF_412_Q_reg ( .D(g806), .SI(g2604), .SE(n2919), .CLK(n3112), .Q(
        g841) );
  SDFFX1 DFF_413_Q_reg ( .D(g6894), .SI(g841), .SE(n2966), .CLK(n3088), .Q(
        g1027), .QN(n2845) );
  SDFFX1 DFF_414_Q_reg ( .D(g6902), .SI(g1027), .SE(n2966), .CLK(n3089), .Q(
        g1003), .QN(n2814) );
  SDFFX1 DFF_415_Q_reg ( .D(g8765), .SI(g1003), .SE(n2966), .CLK(n3089), .Q(
        g1403), .QN(n2773) );
  SDFFX1 DFF_416_Q_reg ( .D(n407), .SI(g1403), .SE(n2966), .CLK(n3089), .Q(
        g1145), .QN(n1617) );
  SDFFX1 DFF_417_Q_reg ( .D(g5148), .SI(g1145), .SE(n2937), .CLK(n3103), .Q(
        g1107), .QN(n1614) );
  SDFFX1 DFF_418_Q_reg ( .D(g7581), .SI(g1107), .SE(n2936), .CLK(n3103), .Q(
        g1223), .QN(n2651) );
  SDFFX1 DFF_419_Q_reg ( .D(g11267), .SI(g1223), .SE(n2986), .CLK(n3079), .Q(
        g406), .QN(n2751) );
  SDFFX1 DFF_420_Q_reg ( .D(g10936), .SI(g406), .SE(n2943), .CLK(n3100), .Q(
        g1811), .QN(n1699) );
  SDFFX1 DFF_421_Q_reg ( .D(g10784), .SI(g1811), .SE(n2942), .CLK(n3100), .Q(
        n3029) );
  SDFFX1 DFF_423_Q_reg ( .D(g10765), .SI(n3029), .SE(n2992), .CLK(n3075), .Q(
        g1654) );
  SDFFX1 DFF_424_Q_reg ( .D(g6332), .SI(g1654), .SE(n2992), .CLK(n3075), .Q(
        g197), .QN(n1678) );
  SDFFX1 DFF_425_Q_reg ( .D(g6479), .SI(g197), .SE(n2988), .CLK(n3077), .Q(
        g1595) );
  SDFFX1 DFF_426_Q_reg ( .D(g6537), .SI(g1595), .SE(n2921), .CLK(n3111), .Q(
        g1537) );
  SDFFX1 DFF_427_Q_reg ( .D(g8434), .SI(g1537), .SE(n2921), .CLK(n3111), .Q(
        g727) );
  SDFFX1 DFF_428_Q_reg ( .D(g6908), .SI(g727), .SE(n2992), .CLK(n3076), .Q(
        test_so8) );
  SDFFX1 DFF_429_Q_reg ( .D(g6243), .SI(test_si9), .SE(n2948), .CLK(n3098), 
        .Q(g798), .QN(n1717) );
  SDFFX1 DFF_430_Q_reg ( .D(g11324), .SI(g798), .SE(n2965), .CLK(n3089), .Q(
        g481), .QN(n1680) );
  SDFFX1 DFF_431_Q_reg ( .D(n316), .SI(g481), .SE(n2950), .CLK(n3097), .Q(
        g4172), .QN(n1647) );
  SDFFX1 DFF_432_Q_reg ( .D(g11609), .SI(g4172), .SE(n2920), .CLK(n3111), .Q(
        g1330) );
  SDFFX1 DFF_433_Q_reg ( .D(g810), .SI(g1330), .SE(n2982), .CLK(n3081), .Q(
        g845) );
  SDFFX1 DFF_434_Q_reg ( .D(g8244), .SI(g845), .SE(n2945), .CLK(n3099), .Q(
        g4181), .QN(n2865) );
  SDFFX1 DFF_435_Q_reg ( .D(g8194), .SI(g4181), .SE(n2936), .CLK(n3103), .Q(
        g1512) );
  SDFFX1 DFF_436_Q_reg ( .D(g113), .SI(g1512), .SE(n2936), .CLK(n3104), .Q(
        n3027), .QN(DFF_436_n1) );
  SDFFX1 DFF_437_Q_reg ( .D(g8052), .SI(n3027), .SE(n2921), .CLK(n3111), .Q(
        g1490), .QN(n2833) );
  SDFFX1 DFF_438_Q_reg ( .D(g4325), .SI(g1490), .SE(n2921), .CLK(n3111), .Q(
        g1166), .QN(n2787) );
  SDFFX1 DFF_440_Q_reg ( .D(g11481), .SI(g1166), .SE(n2965), .CLK(n3089), .Q(
        g348) );
  SDFFX1 DFF_441_Q_reg ( .D(g874), .SI(g348), .SE(n2928), .CLK(n3108), .Q(
        n3026), .QN(n2908) );
  SDFFX1 DFF_442_Q_reg ( .D(g7301), .SI(n3026), .SE(n2979), .CLK(n3082), .Q(
        g1260), .QN(n2750) );
  SDFFX1 DFF_443_Q_reg ( .D(g6035), .SI(g1260), .SE(n2975), .CLK(n3084), .Q(
        g260) );
  SDFFX1 DFF_444_Q_reg ( .D(g8059), .SI(g260), .SE(n2962), .CLK(n3091), .Q(
        g131), .QN(n2762) );
  SDFFX1 DFF_445_Q_reg ( .D(g1854), .SI(g131), .SE(n2961), .CLK(n3091), .Q(
        n3025) );
  SDFFX1 DFF_446_Q_reg ( .D(g6015), .SI(n3025), .SE(n2961), .CLK(n3091), .Q(
        g258) );
  SDFFX1 DFF_447_Q_reg ( .D(g11330), .SI(g258), .SE(n2961), .CLK(n3091), .Q(
        g521), .QN(n1698) );
  SDFFX1 DFF_448_Q_reg ( .D(g11605), .SI(g521), .SE(n2961), .CLK(n3091), .Q(
        g1318) );
  SDFFX1 DFF_449_Q_reg ( .D(g8921), .SI(g1318), .SE(n2961), .CLK(n3091), .Q(
        g1872), .QN(n1616) );
  SDFFX1 DFF_450_Q_reg ( .D(g8883), .SI(g1872), .SE(n2961), .CLK(n3091), .Q(
        g677), .QN(n1656) );
  SDFFX1 DFF_451_Q_reg ( .D(g28), .SI(g677), .SE(n2960), .CLK(n3091), .Q(g2608) );
  SDFFX1 DFF_452_Q_reg ( .D(n30), .SI(g2608), .SE(n2960), .CLK(n3091), .Q(
        n3024) );
  SDFFX1 DFF_453_Q_reg ( .D(g6523), .SI(n3024), .SE(n2990), .CLK(n3076), .Q(
        g1549) );
  SDFFX1 DFF_454_Q_reg ( .D(g11300), .SI(g1549), .SE(n2990), .CLK(n3076), .Q(
        g947) );
  SDFFX1 DFF_455_Q_reg ( .D(g9555), .SI(g947), .SE(n2972), .CLK(n3086), .Q(
        g1834), .QN(n1655) );
  SDFFX1 DFF_456_Q_reg ( .D(g6481), .SI(g1834), .SE(n2970), .CLK(n3087), .Q(
        g1598) );
  SDFFX1 DFF_457_Q_reg ( .D(g4471), .SI(g1598), .SE(n2969), .CLK(n3087), .Q(
        g1121), .QN(n1618) );
  SDFFX1 DFF_458_Q_reg ( .D(g11606), .SI(g1121), .SE(n2943), .CLK(n3100), .Q(
        g1321) );
  SDFFX1 DFF_459_Q_reg ( .D(g11335), .SI(g1321), .SE(n2933), .CLK(n3105), .Q(
        g506), .QN(n1600) );
  SDFFX1 DFF_460_Q_reg ( .D(g10791), .SI(g506), .SE(n2933), .CLK(n3105), .Q(
        g546) );
  SDFFX1 DFF_461_Q_reg ( .D(g8939), .SI(g546), .SE(n2968), .CLK(n3088), .Q(
        g1909), .QN(n2851) );
  SDFFX1 DFF_462_Q_reg ( .D(g83), .SI(g1909), .SE(n2968), .CLK(n3088), .Q(g755) );
  SDFFX1 DFF_463_Q_reg ( .D(g6529), .SI(g755), .SE(n2967), .CLK(n3088), .Q(
        g1552) );
  SDFFX1 DFF_464_Q_reg ( .D(g101), .SI(g1552), .SE(n2967), .CLK(n3088), .Q(
        g2610) );
  SDFFX1 DFF_465_Q_reg ( .D(g10776), .SI(g2610), .SE(n2967), .CLK(n3088), .Q(
        g1687) );
  SDFFX1 DFF_466_Q_reg ( .D(g6514), .SI(g1687), .SE(n2967), .CLK(n3088), .Q(
        g1586) );
  SDFFX1 DFF_467_Q_reg ( .D(g259), .SI(g1586), .SE(n2967), .CLK(n3088), .Q(
        g324), .QN(n2778) );
  SDFFX1 DFF_468_Q_reg ( .D(n444), .SI(g324), .SE(n2967), .CLK(n3088), .Q(
        g1141), .QN(n1660) );
  SDFFX1 DFF_470_Q_reg ( .D(g11639), .SI(g1141), .SE(n2944), .CLK(n3099), .Q(
        g1341), .QN(n2819) );
  SDFFX1 DFF_471_Q_reg ( .D(g4089), .SI(g1341), .SE(n2944), .CLK(n3099), .Q(
        g1710) );
  SDFFX1 DFF_472_Q_reg ( .D(g10785), .SI(g1710), .SE(n2942), .CLK(n3100), .Q(
        n3023) );
  SDFFX1 DFF_473_Q_reg ( .D(g6179), .SI(n3023), .SE(n2992), .CLK(n3075), .Q(
        n3022), .QN(n5134) );
  SDFFX1 DFF_474_Q_reg ( .D(g8053), .SI(n3022), .SE(n2912), .CLK(n3115), .Q(
        g135), .QN(n2764) );
  SDFFX1 DFF_475_Q_reg ( .D(g11329), .SI(g135), .SE(n2912), .CLK(n3115), .Q(
        g525), .QN(n1695) );
  SDFFX1 DFF_476_Q_reg ( .D(g104), .SI(g525), .SE(n2912), .CLK(n3116), .Q(
        g2607) );
  SDFFX1 DFF_477_Q_reg ( .D(g6515), .SI(g2607), .SE(n2957), .CLK(n3093), .Q(
        g1607) );
  SDFFX1 DFF_478_Q_reg ( .D(g258), .SI(g1607), .SE(n2957), .CLK(n3093), .Q(
        g321), .QN(n2818) );
  SDFFX1 DFF_479_Q_reg ( .D(g7204), .SI(g321), .SE(n2948), .CLK(n3097), .Q(
        g8982) );
  SDFFX1 DFF_480_Q_reg ( .D(g11443), .SI(g8982), .SE(n2980), .CLK(n3081), .Q(
        g1275), .QN(n2811) );
  SDFFX1 DFF_481_Q_reg ( .D(g11603), .SI(g1275), .SE(n2964), .CLK(n3090), .Q(
        test_so9) );
  SDFFX1 DFF_482_Q_reg ( .D(g8770), .SI(test_si10), .SE(n2929), .CLK(n3107), 
        .Q(g1615) );
  SDFFX1 DFF_483_Q_reg ( .D(g11292), .SI(g1615), .SE(n2981), .CLK(n3081), .Q(
        g382) );
  SDFFX1 DFF_484_Q_reg ( .D(g6331), .SI(g382), .SE(n2981), .CLK(n3081), .Q(
        n3020) );
  SDFFX1 DFF_485_Q_reg ( .D(g6900), .SI(n3020), .SE(n2981), .CLK(n3081), .Q(
        g266) );
  SDFFX1 DFF_486_Q_reg ( .D(g7294), .SI(g266), .SE(n2981), .CLK(n3081), .Q(
        g1284), .QN(n1864) );
  SDFFX1 DFF_487_Q_reg ( .D(g6829), .SI(g1284), .SE(n2976), .CLK(n3083), .Q(
        n3019) );
  SDFFX1 DFF_488_Q_reg ( .D(g8428), .SI(n3019), .SE(n2954), .CLK(n3094), .Q(
        g673), .QN(n2714) );
  SDFFX1 DFF_489_Q_reg ( .D(n269), .SI(g673), .SE(n2977), .CLK(n3083), .Q(
        n3018) );
  SDFFX1 DFF_490_Q_reg ( .D(g8054), .SI(n3018), .SE(n2970), .CLK(n3086), .Q(
        g162), .QN(n2767) );
  SDFFX1 DFF_491_Q_reg ( .D(g11268), .SI(g162), .SE(n2986), .CLK(n3079), .Q(
        g411), .QN(n2800) );
  SDFFX1 DFF_492_Q_reg ( .D(g11262), .SI(g411), .SE(n2984), .CLK(n3079), .Q(
        g431), .QN(n1876) );
  SDFFX1 DFF_493_Q_reg ( .D(g8283), .SI(g431), .SE(n2917), .CLK(n3113), .Q(
        g1905), .QN(n2862) );
  SDFFX1 DFF_494_Q_reg ( .D(g6193), .SI(g1905), .SE(n2917), .CLK(n3113), .Q(
        g1515), .QN(n1627) );
  SDFFX1 DFF_495_Q_reg ( .D(g8776), .SI(g1515), .SE(n2991), .CLK(n3076), .Q(
        g1630) );
  SDFFX1 DFF_496_Q_reg ( .D(g7143), .SI(g1630), .SE(n2949), .CLK(n3097), .Q(
        g8976) );
  SDFFX1 DFF_497_Q_reg ( .D(g6898), .SI(g8976), .SE(n2913), .CLK(n3115), .Q(
        g991), .QN(n1871) );
  SDFFX1 DFF_498_Q_reg ( .D(g7291), .SI(g991), .SE(n2978), .CLK(n3082), .Q(
        g1300), .QN(n2755) );
  SDFFX1 DFF_499_Q_reg ( .D(g11478), .SI(g1300), .SE(n2935), .CLK(n3104), .Q(
        g339) );
  SDFFX1 DFF_500_Q_reg ( .D(g6000), .SI(g339), .SE(n2935), .CLK(n3104), .Q(
        g256) );
  SDFFX1 DFF_501_Q_reg ( .D(g4264), .SI(g256), .SE(n2935), .CLK(n3104), .Q(
        g1750) );
  SDFFX1 DFF_502_Q_reg ( .D(g102), .SI(g1750), .SE(n2934), .CLK(n3104), .Q(
        g2611) );
  SDFFX1 DFF_503_Q_reg ( .D(g8768), .SI(g2611), .SE(n2934), .CLK(n3104), .Q(
        g1440), .QN(n2830) );
  SDFFX1 DFF_504_Q_reg ( .D(g10863), .SI(g1440), .SE(n2983), .CLK(n3080), .Q(
        g1666) );
  SDFFX1 DFF_505_Q_reg ( .D(g6522), .SI(g1666), .SE(n2983), .CLK(n3080), .Q(
        g1528) );
  SDFFX1 DFF_506_Q_reg ( .D(g11641), .SI(g1528), .SE(n2983), .CLK(n3080), .Q(
        g1351), .QN(n1721) );
  SDFFX1 DFF_507_Q_reg ( .D(g10780), .SI(g1351), .SE(n2942), .CLK(n3101), .Q(
        n3017) );
  SDFFX1 DFF_508_Q_reg ( .D(g8044), .SI(n3017), .SE(n2911), .CLK(n3116), .Q(
        g127), .QN(n1704) );
  SDFFX1 DFF_509_Q_reg ( .D(g11579), .SI(g127), .SE(n2969), .CLK(n3087), .Q(
        g1618) );
  SDFFX1 DFF_510_Q_reg ( .D(g7296), .SI(g1618), .SE(n2980), .CLK(n3081), .Q(
        g1235), .QN(n2775) );
  SDFFX1 DFF_511_Q_reg ( .D(g6923), .SI(g1235), .SE(n2918), .CLK(n3112), .Q(
        g299) );
  SDFFX1 DFF_512_Q_reg ( .D(g11261), .SI(g299), .SE(n2985), .CLK(n3079), .Q(
        g435), .QN(n1878) );
  SDFFX1 DFF_513_Q_reg ( .D(g6638), .SI(g435), .SE(n2949), .CLK(n3097), .Q(
        g8981) );
  SDFFX1 DFF_514_Q_reg ( .D(g6534), .SI(g8981), .SE(n2914), .CLK(n3114), .Q(
        g1555) );
  SDFFX1 DFF_515_Q_reg ( .D(g6895), .SI(g1555), .SE(n2909), .CLK(n3117), .Q(
        g995), .QN(n2812) );
  SDFFX1 DFF_516_Q_reg ( .D(g8771), .SI(g995), .SE(n2975), .CLK(n3084), .Q(
        g1621) );
  SDFFX1 DFF_517_Q_reg ( .D(g4506), .SI(g1621), .SE(n2975), .CLK(n3084), .Q(
        n3016), .QN(n5138) );
  SDFFX1 DFF_518_Q_reg ( .D(g7441), .SI(n3016), .SE(n2939), .CLK(n3102), .Q(
        g643), .QN(n1612) );
  SDFFX1 DFF_519_Q_reg ( .D(g8055), .SI(g643), .SE(n2919), .CLK(n3112), .Q(
        g1494), .QN(n2801) );
  SDFFX1 DFF_520_Q_reg ( .D(g6468), .SI(g1494), .SE(n2916), .CLK(n3113), .Q(
        g1567) );
  SDFFX1 DFF_521_Q_reg ( .D(g8430), .SI(g1567), .SE(n2954), .CLK(n3095), .Q(
        g691) );
  SDFFX1 DFF_522_Q_reg ( .D(g11327), .SI(g691), .SE(n2954), .CLK(n3095), .Q(
        g534), .QN(n2805) );
  SDFFX1 DFF_523_Q_reg ( .D(g6508), .SI(g534), .SE(n2964), .CLK(n3090), .Q(
        g1776), .QN(n1715) );
  SDFFX1 DFF_524_Q_reg ( .D(g10717), .SI(g1776), .SE(n2942), .CLK(n3101), .Q(
        g569) );
  SDFFX1 DFF_525_Q_reg ( .D(g4334), .SI(g569), .SE(n2942), .CLK(n3101), .Q(
        g1160), .QN(n2785) );
  SDFFX1 DFF_526_Q_reg ( .D(n1585), .SI(g1160), .SE(n2941), .CLK(n3101), .Q(
        g1360) );
  SDFFX1 DFF_528_Q_reg ( .D(g6679), .SI(g1360), .SE(n2965), .CLK(n3089), .Q(g1) );
  SDFFX1 DFF_529_Q_reg ( .D(g11336), .SI(g1), .SE(n2965), .CLK(n3089), .Q(g511), .QN(n1679) );
  SDFFX1 DFF_530_Q_reg ( .D(g10771), .SI(g511), .SE(n2940), .CLK(n3101), .Q(
        g1724) );
  SDFFX1 DFF_531_Q_reg ( .D(g5445), .SI(g1724), .SE(n2940), .CLK(n3101), .Q(
        g12) );
  SDFFX1 DFF_532_Q_reg ( .D(g8559), .SI(g12), .SE(n2973), .CLK(n3085), .Q(
        g1878), .QN(n2857) );
  SDFFX1 DFF_533_Q_reg ( .D(g7219), .SI(g1878), .SE(n2948), .CLK(n3098), .Q(
        test_so10) );
  SDFFX1 DFF_158_Q_reg ( .D(g5390), .SI(n3053), .SE(n2989), .CLK(n3077), .Q(
        g1101), .QN(n1654) );
  AND2X2 Tg1_Trojan1 ( .IN1(g6179), .IN2(n30), .Q(Tg1_OUT1) );
  AND2X2 Tg1_Trojan2 ( .IN1(n29), .IN2(n145), .Q(Tg1_OUT2) );
  AND2X2 Tg1_Trojan3 ( .IN1(n1226), .IN2(n1858), .Q(Tg1_OUT3) );
  AND2X2 Tg1_Trojan4 ( .IN1(g5556), .IN2(n32), .Q(Tg1_OUT4) );
  AND4X1 Tg1_Trojan1234 ( .IN1(Tg1_OUT1), .IN2(Tg1_OUT2), .IN3(Tg1_OUT3), 
        .IN4(Tg1_OUT4) );
  NOR2X0 Tg1_Trojan5 ( .IN1(n1391), .IN2(n931), .QN(Tg1_OUT5) );
  NOR2X0 Tg1_Trojan6 ( .IN1(n857), .IN2(n902), .QN(Tg1_OUT6) );
  NOR2X0 Tg1_Trojan7 ( .IN1(n1239), .IN2(n1239), .QN(Tg1_OUT7) );
  NOR2X0 Tg1_Trojan8 ( .IN1(n1055), .IN2(n1016), .QN(Tg1_OUT8) );
  AND4X1 Tg1_Trojan5678 ( .IN1(Tg1_OUT5), .IN2(Tg1_OUT6), .IN3(Tg1_OUT7), 
        .IN4(Tg1_OUT8) );
  AND2X2 Tg2_Trojan1 ( .IN1(n45), .IN2(n25), .Q(Tg2_OUT1) );
  AND2X2 Tg2_Trojan2 ( .IN1(n25), .IN2(n25), .Q(Tg2_OUT2) );
  AND2X2 Tg2_Trojan3 ( .IN1(n25), .IN2(n25), .Q(Tg2_OUT3) );
  AND2X2 Tg2_Trojan4 ( .IN1(n25), .IN2(n25), .Q(Tg2_OUT4) );
  AND4X1 Tg2_Trojan1234 ( .IN1(Tg2_OUT1), .IN2(Tg2_OUT2), .IN3(Tg2_OUT3), 
        .IN4(Tg2_OUT4) );
  AND2X2 Tg2_Trojan5 ( .IN1(n1161), .IN2(n1154), .Q(Tg2_OUT5) );
  AND2X2 Tg2_Trojan6 ( .IN1(n103), .IN2(n72), .Q(Tg2_OUT6) );
  AND2X2 Tg2_Trojan7 ( .IN1(n74), .IN2(n1107), .Q(Tg2_OUT7) );
  AND2X2 Tg2_Trojan8 ( .IN1(n250), .IN2(n2899), .Q(Tg2_OUT8) );
  AND4X1 Tg2_Trojan5678 ( .IN1(Tg2_OUT5), .IN2(Tg2_OUT6), .IN3(Tg2_OUT7), 
        .IN4(Tg2_OUT8) );
  INVX0 TrojanINVtest_se ( .INP(n2994), .ZN(test_se_NOT) );
  AND2X2 Trojan_Trigger ( .IN1(1'b1), .IN2(test_se_NOT), .Q(Trigger_select) );
  MUX21X2 Trojan_Paylaod ( .IN1(g1200), .IN2(n371), .S(Trigger_select), .Q(
        g4207) );
  NBUFFX2 U2957 ( .INP(n3126), .Z(n3076) );
  NBUFFX2 U2958 ( .INP(n3126), .Z(n3077) );
  NBUFFX2 U2959 ( .INP(n3126), .Z(n3075) );
  NBUFFX2 U2960 ( .INP(n3124), .Z(n3083) );
  NBUFFX2 U2961 ( .INP(n3124), .Z(n3086) );
  NBUFFX2 U2962 ( .INP(n3125), .Z(n3081) );
  NBUFFX2 U2963 ( .INP(n3123), .Z(n3088) );
  NBUFFX2 U2964 ( .INP(n3122), .Z(n3095) );
  NBUFFX2 U2965 ( .INP(n3118), .Z(n3115) );
  NBUFFX2 U2966 ( .INP(n3123), .Z(n3090) );
  NBUFFX2 U2967 ( .INP(n3121), .Z(n3101) );
  NBUFFX2 U2968 ( .INP(n3119), .Z(n3110) );
  NBUFFX2 U2969 ( .INP(n3122), .Z(n3096) );
  NBUFFX2 U2970 ( .INP(n3119), .Z(n3111) );
  NBUFFX2 U2971 ( .INP(n3120), .Z(n3106) );
  NBUFFX2 U2972 ( .INP(n3120), .Z(n3105) );
  NBUFFX2 U2973 ( .INP(n3120), .Z(n3103) );
  NBUFFX2 U2974 ( .INP(n3122), .Z(n3097) );
  NBUFFX2 U2975 ( .INP(n3122), .Z(n3094) );
  NBUFFX2 U2976 ( .INP(n3118), .Z(n3116) );
  NBUFFX2 U2977 ( .INP(n3123), .Z(n3089) );
  NBUFFX2 U2978 ( .INP(n3125), .Z(n3080) );
  NBUFFX2 U2979 ( .INP(n3119), .Z(n3112) );
  NBUFFX2 U2980 ( .INP(n3121), .Z(n3102) );
  NBUFFX2 U2981 ( .INP(n3121), .Z(n3099) );
  NBUFFX2 U2982 ( .INP(n3121), .Z(n3098) );
  NBUFFX2 U2983 ( .INP(n3124), .Z(n3087) );
  NBUFFX2 U2984 ( .INP(n3123), .Z(n3091) );
  NBUFFX2 U2985 ( .INP(n3125), .Z(n3082) );
  NBUFFX2 U2986 ( .INP(n3121), .Z(n3100) );
  NBUFFX2 U2987 ( .INP(n3120), .Z(n3107) );
  NBUFFX2 U2988 ( .INP(n3122), .Z(n3093) );
  NBUFFX2 U2989 ( .INP(n3118), .Z(n3114) );
  NBUFFX2 U2990 ( .INP(n3118), .Z(n3113) );
  NBUFFX2 U2991 ( .INP(n3123), .Z(n3092) );
  NBUFFX2 U2992 ( .INP(n3119), .Z(n3109) );
  NBUFFX2 U2993 ( .INP(n3119), .Z(n3108) );
  NBUFFX2 U2994 ( .INP(n3125), .Z(n3078) );
  NBUFFX2 U2995 ( .INP(n3124), .Z(n3084) );
  NBUFFX2 U2996 ( .INP(n3125), .Z(n3079) );
  NBUFFX2 U2997 ( .INP(n3120), .Z(n3104) );
  NBUFFX2 U2998 ( .INP(n3124), .Z(n3085) );
  NBUFFX2 U2999 ( .INP(n3118), .Z(n3117) );
  NBUFFX2 U3000 ( .INP(n3060), .Z(n2909) );
  NBUFFX2 U3001 ( .INP(n3060), .Z(n2910) );
  NBUFFX2 U3002 ( .INP(n3052), .Z(n2911) );
  NBUFFX2 U3003 ( .INP(n3052), .Z(n2912) );
  NBUFFX2 U3004 ( .INP(n3052), .Z(n2913) );
  NBUFFX2 U3005 ( .INP(n3049), .Z(n2914) );
  NBUFFX2 U3006 ( .INP(n3049), .Z(n2915) );
  NBUFFX2 U3007 ( .INP(n3049), .Z(n2916) );
  NBUFFX2 U3008 ( .INP(n3043), .Z(n2917) );
  NBUFFX2 U3009 ( .INP(n3043), .Z(n2918) );
  NBUFFX2 U3010 ( .INP(n3043), .Z(n2919) );
  NBUFFX2 U3011 ( .INP(n3039), .Z(n2920) );
  NBUFFX2 U3012 ( .INP(n3039), .Z(n2921) );
  NBUFFX2 U3013 ( .INP(n3039), .Z(n2922) );
  NBUFFX2 U3014 ( .INP(n3032), .Z(n2923) );
  NBUFFX2 U3015 ( .INP(n3032), .Z(n2924) );
  NBUFFX2 U3016 ( .INP(n3032), .Z(n2925) );
  NBUFFX2 U3017 ( .INP(n3028), .Z(n2926) );
  NBUFFX2 U3018 ( .INP(n3028), .Z(n2927) );
  NBUFFX2 U3019 ( .INP(n3028), .Z(n2928) );
  NBUFFX2 U3020 ( .INP(n3021), .Z(n2929) );
  NBUFFX2 U3021 ( .INP(n3021), .Z(n2930) );
  NBUFFX2 U3022 ( .INP(n3021), .Z(n2931) );
  NBUFFX2 U3023 ( .INP(n3015), .Z(n2932) );
  NBUFFX2 U3024 ( .INP(n3015), .Z(n2933) );
  NBUFFX2 U3025 ( .INP(n3015), .Z(n2934) );
  NBUFFX2 U3026 ( .INP(n3014), .Z(n2935) );
  NBUFFX2 U3027 ( .INP(n3014), .Z(n2936) );
  NBUFFX2 U3028 ( .INP(n3014), .Z(n2937) );
  NBUFFX2 U3029 ( .INP(n3013), .Z(n2938) );
  NBUFFX2 U3030 ( .INP(n3013), .Z(n2939) );
  NBUFFX2 U3031 ( .INP(n3013), .Z(n2940) );
  NBUFFX2 U3032 ( .INP(n3012), .Z(n2941) );
  NBUFFX2 U3033 ( .INP(n3012), .Z(n2942) );
  NBUFFX2 U3034 ( .INP(n3012), .Z(n2943) );
  NBUFFX2 U3035 ( .INP(n3011), .Z(n2944) );
  NBUFFX2 U3036 ( .INP(n3011), .Z(n2945) );
  NBUFFX2 U3037 ( .INP(n3011), .Z(n2946) );
  NBUFFX2 U3038 ( .INP(n3010), .Z(n2947) );
  NBUFFX2 U3039 ( .INP(n3010), .Z(n2948) );
  NBUFFX2 U3040 ( .INP(n3010), .Z(n2949) );
  NBUFFX2 U3041 ( .INP(n3009), .Z(n2950) );
  NBUFFX2 U3042 ( .INP(n3009), .Z(n2951) );
  NBUFFX2 U3043 ( .INP(n3009), .Z(n2952) );
  NBUFFX2 U3044 ( .INP(n3008), .Z(n2953) );
  NBUFFX2 U3045 ( .INP(n3008), .Z(n2954) );
  NBUFFX2 U3046 ( .INP(n3008), .Z(n2955) );
  NBUFFX2 U3047 ( .INP(n3007), .Z(n2956) );
  NBUFFX2 U3048 ( .INP(n3007), .Z(n2957) );
  NBUFFX2 U3049 ( .INP(n3007), .Z(n2958) );
  NBUFFX2 U3050 ( .INP(n3006), .Z(n2959) );
  NBUFFX2 U3051 ( .INP(n3006), .Z(n2960) );
  NBUFFX2 U3052 ( .INP(n3006), .Z(n2961) );
  NBUFFX2 U3053 ( .INP(n3005), .Z(n2962) );
  NBUFFX2 U3054 ( .INP(n3005), .Z(n2963) );
  NBUFFX2 U3055 ( .INP(n3005), .Z(n2964) );
  NBUFFX2 U3056 ( .INP(n3004), .Z(n2965) );
  NBUFFX2 U3057 ( .INP(n3004), .Z(n2966) );
  NBUFFX2 U3058 ( .INP(n3004), .Z(n2967) );
  NBUFFX2 U3059 ( .INP(n3003), .Z(n2968) );
  NBUFFX2 U3060 ( .INP(n3003), .Z(n2969) );
  NBUFFX2 U3061 ( .INP(n3003), .Z(n2970) );
  NBUFFX2 U3062 ( .INP(n3002), .Z(n2971) );
  NBUFFX2 U3063 ( .INP(n3002), .Z(n2972) );
  NBUFFX2 U3064 ( .INP(n3002), .Z(n2973) );
  NBUFFX2 U3065 ( .INP(n3001), .Z(n2974) );
  NBUFFX2 U3066 ( .INP(n3001), .Z(n2975) );
  NBUFFX2 U3067 ( .INP(n3001), .Z(n2976) );
  NBUFFX2 U3068 ( .INP(n3000), .Z(n2977) );
  NBUFFX2 U3069 ( .INP(n3000), .Z(n2978) );
  NBUFFX2 U3070 ( .INP(n3000), .Z(n2979) );
  NBUFFX2 U3071 ( .INP(n2999), .Z(n2980) );
  NBUFFX2 U3072 ( .INP(n2999), .Z(n2981) );
  NBUFFX2 U3073 ( .INP(n2999), .Z(n2982) );
  NBUFFX2 U3074 ( .INP(n2998), .Z(n2983) );
  NBUFFX2 U3075 ( .INP(n2998), .Z(n2984) );
  NBUFFX2 U3076 ( .INP(n2998), .Z(n2985) );
  NBUFFX2 U3077 ( .INP(n2997), .Z(n2986) );
  NBUFFX2 U3078 ( .INP(n2997), .Z(n2987) );
  NBUFFX2 U3079 ( .INP(n2997), .Z(n2988) );
  NBUFFX2 U3080 ( .INP(n2996), .Z(n2989) );
  NBUFFX2 U3081 ( .INP(n2996), .Z(n2990) );
  NBUFFX2 U3082 ( .INP(n2996), .Z(n2991) );
  NBUFFX2 U3083 ( .INP(n2995), .Z(n2992) );
  NBUFFX2 U3084 ( .INP(n2995), .Z(n2993) );
  NBUFFX2 U3085 ( .INP(n2995), .Z(n2994) );
  NBUFFX2 U3086 ( .INP(n3074), .Z(n2995) );
  NBUFFX2 U3087 ( .INP(n3074), .Z(n2996) );
  NBUFFX2 U3088 ( .INP(n3073), .Z(n2997) );
  NBUFFX2 U3089 ( .INP(n3073), .Z(n2998) );
  NBUFFX2 U3091 ( .INP(n3073), .Z(n2999) );
  NBUFFX2 U3093 ( .INP(n3072), .Z(n3000) );
  NBUFFX2 U3095 ( .INP(n3072), .Z(n3001) );
  NBUFFX2 U3097 ( .INP(n3072), .Z(n3002) );
  NBUFFX2 U3099 ( .INP(n3071), .Z(n3003) );
  NBUFFX2 U3100 ( .INP(n3071), .Z(n3004) );
  NBUFFX2 U3101 ( .INP(n3071), .Z(n3005) );
  NBUFFX2 U3102 ( .INP(n3070), .Z(n3006) );
  NBUFFX2 U3103 ( .INP(n3070), .Z(n3007) );
  NBUFFX2 U3104 ( .INP(n3070), .Z(n3008) );
  NBUFFX2 U3105 ( .INP(n3069), .Z(n3009) );
  NBUFFX2 U3106 ( .INP(n3069), .Z(n3010) );
  NBUFFX2 U3107 ( .INP(n3069), .Z(n3011) );
  NBUFFX2 U3108 ( .INP(n3068), .Z(n3012) );
  NBUFFX2 U3109 ( .INP(n3068), .Z(n3013) );
  NBUFFX2 U3110 ( .INP(n3068), .Z(n3014) );
  NBUFFX2 U3111 ( .INP(n3067), .Z(n3015) );
  NBUFFX2 U3112 ( .INP(n3067), .Z(n3021) );
  NBUFFX2 U3113 ( .INP(n3067), .Z(n3028) );
  NBUFFX2 U3114 ( .INP(n3066), .Z(n3032) );
  NBUFFX2 U3115 ( .INP(n3066), .Z(n3039) );
  NBUFFX2 U3116 ( .INP(n3066), .Z(n3043) );
  NBUFFX2 U3117 ( .INP(n3063), .Z(n3049) );
  NBUFFX2 U3118 ( .INP(n3063), .Z(n3052) );
  NBUFFX2 U3119 ( .INP(n3063), .Z(n3060) );
  NBUFFX2 U3120 ( .INP(test_se), .Z(n3063) );
  NBUFFX2 U3121 ( .INP(n3070), .Z(n3066) );
  NBUFFX2 U3122 ( .INP(n3006), .Z(n3067) );
  NBUFFX2 U3123 ( .INP(n3007), .Z(n3068) );
  NBUFFX2 U3125 ( .INP(n3008), .Z(n3069) );
  NBUFFX2 U3126 ( .INP(test_se), .Z(n3070) );
  NBUFFX2 U3127 ( .INP(test_se), .Z(n3071) );
  NBUFFX2 U3128 ( .INP(n3060), .Z(n3072) );
  NBUFFX2 U3129 ( .INP(test_se), .Z(n3073) );
  NBUFFX2 U3130 ( .INP(n3063), .Z(n3074) );
  NBUFFX2 U3131 ( .INP(n3129), .Z(n3118) );
  NBUFFX2 U3132 ( .INP(n3129), .Z(n3119) );
  NBUFFX2 U3133 ( .INP(n3129), .Z(n3120) );
  NBUFFX2 U3134 ( .INP(n3128), .Z(n3121) );
  NBUFFX2 U3135 ( .INP(n3128), .Z(n3122) );
  NBUFFX2 U3136 ( .INP(n3128), .Z(n3123) );
  NBUFFX2 U3137 ( .INP(n3127), .Z(n3124) );
  NBUFFX2 U3138 ( .INP(n3127), .Z(n3125) );
  NBUFFX2 U3139 ( .INP(n3127), .Z(n3126) );
  NBUFFX2 U3140 ( .INP(CK), .Z(n3127) );
  NBUFFX2 U3141 ( .INP(CK), .Z(n3128) );
  NBUFFX2 U3142 ( .INP(CK), .Z(n3129) );
  OR2X1 U3144 ( .IN1(n3130), .IN2(n3131), .Q(n962) );
  AND2X1 U3145 ( .IN1(n3132), .IN2(n1696), .Q(n3131) );
  AND2X1 U3146 ( .IN1(n3133), .IN2(g731), .Q(n3130) );
  OR2X1 U3147 ( .IN1(n3134), .IN2(n3135), .Q(n9) );
  AND2X1 U3148 ( .IN1(n3136), .IN2(n1697), .Q(n3135) );
  INVX0 U3149 ( .INP(n3137), .ZN(n3136) );
  INVX0 U3150 ( .INP(n3138), .ZN(n3134) );
  OR2X1 U3151 ( .IN1(n857), .IN2(n1697), .Q(n3138) );
  AND2X1 U3152 ( .IN1(n804), .IN2(n3139), .Q(n838) );
  INVX0 U3153 ( .INP(n3140), .ZN(n534) );
  INVX0 U3154 ( .INP(n3141), .ZN(n524) );
  INVX0 U3155 ( .INP(n3142), .ZN(n499) );
  INVX0 U3156 ( .INP(n3143), .ZN(n444) );
  OR2X1 U3157 ( .IN1(n519), .IN2(n1660), .Q(n3143) );
  AND2X1 U3158 ( .IN1(g109), .IN2(g1145), .Q(n407) );
  AND2X1 U3159 ( .IN1(g109), .IN2(g1137), .Q(n352) );
  INVX0 U3160 ( .INP(n3144), .ZN(n316) );
  OR2X1 U3161 ( .IN1(n3145), .IN2(n2838), .Q(n3144) );
  AND2X1 U3162 ( .IN1(n3146), .IN2(n3147), .Q(n3145) );
  OR2X1 U3163 ( .IN1(g750), .IN2(n1647), .Q(n3146) );
  INVX0 U3164 ( .INP(n3148), .ZN(n2896) );
  OR2X1 U3165 ( .IN1(n3149), .IN2(n1722), .Q(n3148) );
  INVX0 U3166 ( .INP(n3150), .ZN(n269) );
  AND2X1 U3167 ( .IN1(g109), .IN2(g1133), .Q(n187) );
  OR2X1 U3168 ( .IN1(n2900), .IN2(g627), .Q(n178) );
  INVX0 U3169 ( .INP(n3151), .ZN(n160) );
  OR2X1 U3170 ( .IN1(n3152), .IN2(n3153), .Q(n1588) );
  OR2X1 U3172 ( .IN1(g42), .IN2(n3154), .Q(n3153) );
  OR2X1 U3173 ( .IN1(n3154), .IN2(n3155), .Q(n1587) );
  OR2X1 U3174 ( .IN1(n3156), .IN2(n3155), .Q(n1586) );
  OR2X1 U3175 ( .IN1(n3152), .IN2(n3157), .Q(n1585) );
  OR2X1 U3176 ( .IN1(g42), .IN2(n3156), .Q(n3157) );
  OR2X1 U3177 ( .IN1(n2871), .IN2(n2872), .Q(n1214) );
  OR2X1 U3178 ( .IN1(n2870), .IN2(n3158), .Q(n1153) );
  INVX0 U3179 ( .INP(n1193), .ZN(n3158) );
  OR2X1 U3180 ( .IN1(n2859), .IN2(n3159), .Q(n1151) );
  OR2X1 U3181 ( .IN1(n2869), .IN2(n3160), .Q(n1099) );
  INVX0 U3182 ( .INP(n1125), .ZN(n3160) );
  OR2X1 U3183 ( .IN1(n2858), .IN2(n3161), .Q(n1097) );
  INVX0 U3184 ( .INP(n1123), .ZN(n3161) );
  INVX0 U3185 ( .INP(n3162), .ZN(n104) );
  INVX0 U3186 ( .INP(n3163), .ZN(n1) );
  AND2X1 U3187 ( .IN1(n2844), .IN2(n2882), .Q(n3163) );
  AND2X1 U3188 ( .IN1(g18), .IN2(n3164), .Q(g9721) );
  XNOR2X1 U3189 ( .IN1(g611), .IN2(n3165), .Q(n3164) );
  AND2X1 U3190 ( .IN1(n3166), .IN2(n3167), .Q(n3165) );
  OR2X1 U3191 ( .IN1(n3168), .IN2(n3169), .Q(n3166) );
  AND2X1 U3192 ( .IN1(n1645), .IN2(n3170), .Q(n3168) );
  OR2X1 U3193 ( .IN1(n804), .IN2(n3171), .Q(n3170) );
  AND2X1 U3194 ( .IN1(n3172), .IN2(g18), .Q(g9555) );
  AND2X1 U3195 ( .IN1(n3173), .IN2(n3174), .Q(n3172) );
  OR2X1 U3196 ( .IN1(n806), .IN2(g1834), .Q(n3174) );
  OR2X1 U3197 ( .IN1(n1655), .IN2(n3175), .Q(n3173) );
  INVX0 U3198 ( .INP(n3176), .ZN(n3175) );
  AND2X1 U3199 ( .IN1(n808), .IN2(n926), .Q(n3176) );
  OR2X1 U3200 ( .IN1(n3177), .IN2(g1840), .Q(n808) );
  AND2X1 U3201 ( .IN1(n252), .IN2(n3178), .Q(n3177) );
  INVX0 U3202 ( .INP(n3179), .ZN(n252) );
  OR2X1 U3203 ( .IN1(n3180), .IN2(n3181), .Q(g9451) );
  OR2X1 U3204 ( .IN1(g31), .IN2(g30), .Q(n3181) );
  AND2X1 U3205 ( .IN1(n3182), .IN2(g18), .Q(g9272) );
  AND2X1 U3206 ( .IN1(n3183), .IN2(n3184), .Q(n3182) );
  OR2X1 U3207 ( .IN1(n1605), .IN2(n3185), .Q(n3184) );
  OR2X1 U3208 ( .IN1(g1828), .IN2(n3186), .Q(n3183) );
  INVX0 U3209 ( .INP(n3187), .ZN(n3186) );
  AND2X1 U3210 ( .IN1(n3188), .IN2(n3185), .Q(n3187) );
  OR2X1 U3211 ( .IN1(n3189), .IN2(n3178), .Q(n3185) );
  AND2X1 U3212 ( .IN1(n3190), .IN2(n3191), .Q(n3189) );
  OR2X1 U3213 ( .IN1(n1643), .IN2(n817), .Q(n3191) );
  INVX0 U3214 ( .INP(n3192), .ZN(n3190) );
  AND2X1 U3215 ( .IN1(n3193), .IN2(g18), .Q(g9269) );
  XNOR2X1 U3216 ( .IN1(n1643), .IN2(n3194), .Q(n3193) );
  AND2X1 U3217 ( .IN1(n812), .IN2(n3195), .Q(n3194) );
  OR2X1 U3218 ( .IN1(n3196), .IN2(n3197), .Q(n3195) );
  OR2X1 U3219 ( .IN1(n3198), .IN2(n3199), .Q(n3197) );
  AND2X1 U3220 ( .IN1(n1643), .IN2(n3200), .Q(n3196) );
  AND2X1 U3221 ( .IN1(n3201), .IN2(g18), .Q(g9266) );
  XNOR2X1 U3222 ( .IN1(n3202), .IN2(g1814), .Q(n3201) );
  OR2X1 U3223 ( .IN1(n3203), .IN2(n3178), .Q(n3202) );
  AND2X1 U3224 ( .IN1(n3204), .IN2(n3205), .Q(n3203) );
  OR2X1 U3225 ( .IN1(n817), .IN2(g1822), .Q(n3205) );
  INVX0 U3226 ( .INP(n3200), .ZN(n817) );
  AND2X1 U3227 ( .IN1(n3206), .IN2(n3179), .Q(n3204) );
  AND2X1 U3228 ( .IN1(n3207), .IN2(g18), .Q(g9150) );
  AND2X1 U3229 ( .IN1(n3208), .IN2(n3209), .Q(n3207) );
  INVX0 U3230 ( .INP(n3210), .ZN(n3209) );
  AND2X1 U3231 ( .IN1(g605), .IN2(n3211), .Q(n3210) );
  OR2X1 U3232 ( .IN1(g605), .IN2(n3212), .Q(n3208) );
  OR2X1 U3233 ( .IN1(n3213), .IN2(n3211), .Q(n3212) );
  OR2X1 U3234 ( .IN1(n3214), .IN2(n3215), .Q(n3211) );
  AND2X1 U3235 ( .IN1(n804), .IN2(n3216), .Q(n3214) );
  OR2X1 U3236 ( .IN1(n3217), .IN2(n3218), .Q(n3216) );
  OR2X1 U3237 ( .IN1(n3219), .IN2(n3220), .Q(n3218) );
  AND2X1 U3238 ( .IN1(n3221), .IN2(g599), .Q(n3217) );
  AND2X1 U3239 ( .IN1(g18), .IN2(n3222), .Q(g9124) );
  XNOR2X1 U3240 ( .IN1(n836), .IN2(g599), .Q(n3222) );
  AND2X1 U3241 ( .IN1(g18), .IN2(n3223), .Q(g9110) );
  XNOR2X1 U3242 ( .IN1(g591), .IN2(n3224), .Q(n3223) );
  AND2X1 U3243 ( .IN1(n837), .IN2(n3225), .Q(n3224) );
  OR2X1 U3244 ( .IN1(n3226), .IN2(n3227), .Q(n3225) );
  AND2X1 U3245 ( .IN1(n3228), .IN2(n3171), .Q(n3226) );
  OR2X1 U3246 ( .IN1(n3229), .IN2(n3230), .Q(n837) );
  OR2X1 U3247 ( .IN1(g599), .IN2(n3227), .Q(n3230) );
  OR2X1 U3248 ( .IN1(n3231), .IN2(n3232), .Q(g8973) );
  AND2X1 U3249 ( .IN1(n3233), .IN2(n3234), .Q(n3231) );
  XOR2X1 U3250 ( .IN1(n3235), .IN2(n1615), .Q(n3233) );
  OR2X1 U3251 ( .IN1(n3236), .IN2(n3237), .Q(n3235) );
  AND2X1 U3252 ( .IN1(n2856), .IN2(n3238), .Q(n3236) );
  OR2X1 U3253 ( .IN1(n3239), .IN2(n3240), .Q(g8945) );
  AND2X1 U3254 ( .IN1(n3241), .IN2(n3242), .Q(n3239) );
  XOR2X1 U3255 ( .IN1(n1697), .IN2(n3243), .Q(n3241) );
  AND2X1 U3256 ( .IN1(n3244), .IN2(n3245), .Q(n3243) );
  OR2X1 U3257 ( .IN1(n2810), .IN2(n3246), .Q(n3245) );
  OR2X1 U3258 ( .IN1(n3247), .IN2(n3248), .Q(n3244) );
  OR2X1 U3259 ( .IN1(n3249), .IN2(n3250), .Q(n3248) );
  AND2X1 U3260 ( .IN1(n3137), .IN2(n857), .Q(n3250) );
  OR2X1 U3261 ( .IN1(n1694), .IN2(n3251), .Q(n857) );
  OR2X1 U3262 ( .IN1(n3252), .IN2(n3253), .Q(n3137) );
  OR2X1 U3263 ( .IN1(g1927), .IN2(n3254), .Q(n3253) );
  OR2X1 U3264 ( .IN1(g1918), .IN2(g1909), .Q(n3254) );
  OR2X1 U3265 ( .IN1(g1936), .IN2(n3255), .Q(n3252) );
  OR2X1 U3266 ( .IN1(n3256), .IN2(g1900), .Q(n3255) );
  OR2X1 U3267 ( .IN1(n3257), .IN2(n3240), .Q(g8944) );
  AND2X1 U3268 ( .IN1(n3258), .IN2(n3242), .Q(n3257) );
  XNOR2X1 U3269 ( .IN1(n3259), .IN2(g1936), .Q(n3258) );
  OR2X1 U3270 ( .IN1(n3260), .IN2(n3249), .Q(n3259) );
  AND2X1 U3271 ( .IN1(n3261), .IN2(n3262), .Q(n3260) );
  OR2X1 U3272 ( .IN1(g1927), .IN2(n3263), .Q(n3262) );
  AND2X1 U3273 ( .IN1(n3264), .IN2(n3265), .Q(n3261) );
  OR2X1 U3274 ( .IN1(n3251), .IN2(n3247), .Q(n3265) );
  OR2X1 U3275 ( .IN1(n3266), .IN2(n3267), .Q(n3251) );
  INVX0 U3276 ( .INP(n3268), .ZN(n3267) );
  AND2X1 U3277 ( .IN1(n3269), .IN2(n921), .Q(n3268) );
  OR2X1 U3278 ( .IN1(n1675), .IN2(n3270), .Q(n3266) );
  OR2X1 U3279 ( .IN1(n2851), .IN2(n2795), .Q(n3270) );
  OR2X1 U3280 ( .IN1(n2747), .IN2(n3246), .Q(n3264) );
  OR2X1 U3281 ( .IN1(n3271), .IN2(n3240), .Q(g8943) );
  AND2X1 U3282 ( .IN1(n3272), .IN2(n3242), .Q(n3271) );
  XNOR2X1 U3283 ( .IN1(n1663), .IN2(n3273), .Q(n3272) );
  AND2X1 U3284 ( .IN1(n3274), .IN2(n3275), .Q(n3273) );
  AND2X1 U3285 ( .IN1(n3276), .IN2(n3277), .Q(n3274) );
  OR2X1 U3286 ( .IN1(n3246), .IN2(g1887), .Q(n3277) );
  OR2X1 U3287 ( .IN1(n3247), .IN2(n3278), .Q(n3276) );
  XNOR2X1 U3288 ( .IN1(n3279), .IN2(n1616), .Q(n3278) );
  OR2X1 U3289 ( .IN1(n3280), .IN2(n3240), .Q(g8941) );
  AND2X1 U3290 ( .IN1(n3281), .IN2(n3242), .Q(n3280) );
  XNOR2X1 U3291 ( .IN1(n3282), .IN2(g1927), .Q(n3281) );
  OR2X1 U3292 ( .IN1(n3283), .IN2(n3249), .Q(n3282) );
  AND2X1 U3293 ( .IN1(n3284), .IN2(n3285), .Q(n3283) );
  OR2X1 U3294 ( .IN1(n2795), .IN2(n3286), .Q(n3285) );
  AND2X1 U3295 ( .IN1(n3287), .IN2(n3263), .Q(n3284) );
  OR2X1 U3296 ( .IN1(g1918), .IN2(n3288), .Q(n3263) );
  OR2X1 U3297 ( .IN1(n3246), .IN2(n2748), .Q(n3287) );
  OR2X1 U3298 ( .IN1(n3289), .IN2(n3240), .Q(g8940) );
  AND2X1 U3299 ( .IN1(n3290), .IN2(n3242), .Q(n3289) );
  XNOR2X1 U3300 ( .IN1(n3291), .IN2(g1918), .Q(n3290) );
  OR2X1 U3301 ( .IN1(n3292), .IN2(n3249), .Q(n3291) );
  AND2X1 U3302 ( .IN1(n3293), .IN2(n3294), .Q(n3292) );
  OR2X1 U3303 ( .IN1(n3246), .IN2(n1718), .Q(n3294) );
  AND2X1 U3304 ( .IN1(n3286), .IN2(n3288), .Q(n3293) );
  OR2X1 U3305 ( .IN1(n3295), .IN2(n3296), .Q(n3288) );
  OR2X1 U3306 ( .IN1(g1900), .IN2(g1909), .Q(n3296) );
  OR2X1 U3307 ( .IN1(n3297), .IN2(n3298), .Q(n3286) );
  OR2X1 U3308 ( .IN1(n2851), .IN2(n1675), .Q(n3298) );
  OR2X1 U3309 ( .IN1(n3299), .IN2(n3240), .Q(g8939) );
  AND2X1 U3310 ( .IN1(n3300), .IN2(n3242), .Q(n3299) );
  XNOR2X1 U3311 ( .IN1(n3301), .IN2(g1909), .Q(n3300) );
  OR2X1 U3312 ( .IN1(n3302), .IN2(n3249), .Q(n3301) );
  AND2X1 U3313 ( .IN1(n3303), .IN2(n3304), .Q(n3302) );
  OR2X1 U3314 ( .IN1(n3246), .IN2(n2745), .Q(n3304) );
  AND2X1 U3315 ( .IN1(n3305), .IN2(n3306), .Q(n3303) );
  OR2X1 U3316 ( .IN1(n1675), .IN2(n3297), .Q(n3306) );
  OR2X1 U3317 ( .IN1(g1900), .IN2(n3295), .Q(n3305) );
  OR2X1 U3318 ( .IN1(n3307), .IN2(n3240), .Q(g8938) );
  AND2X1 U3319 ( .IN1(n3308), .IN2(n3242), .Q(n3307) );
  XNOR2X1 U3320 ( .IN1(n3309), .IN2(g1900), .Q(n3308) );
  OR2X1 U3321 ( .IN1(n3310), .IN2(n3249), .Q(n3309) );
  AND2X1 U3322 ( .IN1(n3311), .IN2(n3312), .Q(n3310) );
  OR2X1 U3323 ( .IN1(n3246), .IN2(n2862), .Q(n3312) );
  AND2X1 U3324 ( .IN1(n3297), .IN2(n3295), .Q(n3311) );
  OR2X1 U3325 ( .IN1(n3256), .IN2(n3247), .Q(n3295) );
  INVX0 U3326 ( .INP(n3313), .ZN(n3256) );
  AND2X1 U3327 ( .IN1(n3314), .IN2(n3315), .Q(n3313) );
  AND2X1 U3328 ( .IN1(n1657), .IN2(n1663), .Q(n3315) );
  OR2X1 U3329 ( .IN1(n3247), .IN2(n3316), .Q(n3297) );
  OR2X1 U3330 ( .IN1(n1657), .IN2(n3317), .Q(n3316) );
  OR2X1 U3331 ( .IN1(n3318), .IN2(n3240), .Q(g8937) );
  AND2X1 U3332 ( .IN1(n3319), .IN2(n3242), .Q(n3318) );
  XNOR2X1 U3333 ( .IN1(n1657), .IN2(n3320), .Q(n3319) );
  OR2X1 U3334 ( .IN1(n3321), .IN2(n3322), .Q(n3320) );
  AND2X1 U3335 ( .IN1(n3323), .IN2(n3246), .Q(n3322) );
  AND2X1 U3336 ( .IN1(n3324), .IN2(n3275), .Q(n3323) );
  INVX0 U3337 ( .INP(n3249), .ZN(n3275) );
  OR2X1 U3338 ( .IN1(n3325), .IN2(n3269), .Q(n3324) );
  INVX0 U3339 ( .INP(n3317), .ZN(n3269) );
  OR2X1 U3340 ( .IN1(n3279), .IN2(n3326), .Q(n3317) );
  OR2X1 U3341 ( .IN1(n1663), .IN2(n1616), .Q(n3326) );
  AND2X1 U3342 ( .IN1(n3314), .IN2(n1663), .Q(n3325) );
  AND2X1 U3343 ( .IN1(n1616), .IN2(n3279), .Q(n3314) );
  INVX0 U3344 ( .INP(n3327), .ZN(n3279) );
  OR2X1 U3345 ( .IN1(n3328), .IN2(n3192), .Q(n3327) );
  OR2X1 U3346 ( .IN1(n3329), .IN2(n3198), .Q(n3192) );
  AND2X1 U3347 ( .IN1(n1605), .IN2(n3330), .Q(n3329) );
  AND2X1 U3348 ( .IN1(n1643), .IN2(g1814), .Q(n3328) );
  AND2X1 U3349 ( .IN1(n3247), .IN2(g1896), .Q(n3321) );
  OR2X1 U3350 ( .IN1(n3331), .IN2(n3232), .Q(g8926) );
  AND2X1 U3351 ( .IN1(n3234), .IN2(n3332), .Q(n3331) );
  XOR2X1 U3352 ( .IN1(g731), .IN2(n32), .Q(n3332) );
  OR2X1 U3353 ( .IN1(n3333), .IN2(n3334), .Q(n32) );
  AND2X1 U3354 ( .IN1(n3335), .IN2(n3336), .Q(n3334) );
  OR2X1 U3355 ( .IN1(n3133), .IN2(n3132), .Q(n3336) );
  INVX0 U3356 ( .INP(n3337), .ZN(n3132) );
  OR2X1 U3357 ( .IN1(n3338), .IN2(n3339), .Q(n3337) );
  OR2X1 U3358 ( .IN1(g713), .IN2(n3340), .Q(n3339) );
  OR2X1 U3359 ( .IN1(g704), .IN2(g695), .Q(n3340) );
  OR2X1 U3360 ( .IN1(n3341), .IN2(n3342), .Q(n3338) );
  INVX0 U3361 ( .INP(n3343), .ZN(n3342) );
  AND2X1 U3362 ( .IN1(n1676), .IN2(n1693), .Q(n3343) );
  INVX0 U3363 ( .INP(n902), .ZN(n3133) );
  OR2X1 U3364 ( .IN1(n1693), .IN2(n3344), .Q(n902) );
  AND2X1 U3365 ( .IN1(g736), .IN2(n3238), .Q(n3333) );
  OR2X1 U3366 ( .IN1(n3345), .IN2(n3232), .Q(g8923) );
  AND2X1 U3367 ( .IN1(n3346), .IN2(n3234), .Q(n3345) );
  XNOR2X1 U3368 ( .IN1(n1693), .IN2(n3347), .Q(n3346) );
  AND2X1 U3369 ( .IN1(n3348), .IN2(n3349), .Q(n3347) );
  OR2X1 U3370 ( .IN1(n3350), .IN2(n3351), .Q(n3349) );
  OR2X1 U3371 ( .IN1(n3352), .IN2(n3353), .Q(n3351) );
  INVX0 U3372 ( .INP(n3354), .ZN(n3353) );
  OR2X1 U3373 ( .IN1(n3238), .IN2(n3344), .Q(n3354) );
  OR2X1 U3374 ( .IN1(n3355), .IN2(n3356), .Q(n3344) );
  OR2X1 U3375 ( .IN1(n3357), .IN2(n3358), .Q(n3356) );
  INVX0 U3376 ( .INP(n967), .ZN(n3358) );
  OR2X1 U3377 ( .IN1(n1676), .IN2(n3359), .Q(n3355) );
  OR2X1 U3378 ( .IN1(n2850), .IN2(n2796), .Q(n3359) );
  AND2X1 U3379 ( .IN1(n3238), .IN2(g727), .Q(n3352) );
  INVX0 U3380 ( .INP(n3360), .ZN(n3350) );
  OR2X1 U3381 ( .IN1(n3361), .IN2(g713), .Q(n3360) );
  OR2X1 U3382 ( .IN1(n3362), .IN2(n3232), .Q(g8922) );
  AND2X1 U3383 ( .IN1(n3363), .IN2(n3234), .Q(n3362) );
  XOR2X1 U3384 ( .IN1(n3364), .IN2(n1662), .Q(n3363) );
  OR2X1 U3385 ( .IN1(n3237), .IN2(n3365), .Q(n3364) );
  OR2X1 U3386 ( .IN1(n3366), .IN2(n3367), .Q(n3365) );
  AND2X1 U3387 ( .IN1(n3368), .IN2(n3369), .Q(n3367) );
  XNOR2X1 U3388 ( .IN1(n1615), .IN2(n3370), .Q(n3368) );
  AND2X1 U3389 ( .IN1(n2714), .IN2(n3238), .Q(n3366) );
  OR2X1 U3390 ( .IN1(n3371), .IN2(n3240), .Q(g8921) );
  AND2X1 U3391 ( .IN1(n3372), .IN2(n3373), .Q(n3240) );
  AND2X1 U3392 ( .IN1(n3188), .IN2(n916), .Q(n3373) );
  INVX0 U3393 ( .INP(n3374), .ZN(n3372) );
  OR2X1 U3394 ( .IN1(n3198), .IN2(n3242), .Q(n3374) );
  AND2X1 U3395 ( .IN1(n3375), .IN2(n3242), .Q(n3371) );
  AND2X1 U3396 ( .IN1(n3178), .IN2(n3188), .Q(n3242) );
  INVX0 U3397 ( .INP(n812), .ZN(n3178) );
  XOR2X1 U3398 ( .IN1(n3376), .IN2(n1616), .Q(n3375) );
  OR2X1 U3399 ( .IN1(n3377), .IN2(n3249), .Q(n3376) );
  AND2X1 U3400 ( .IN1(n918), .IN2(n3246), .Q(n3249) );
  INVX0 U3401 ( .INP(n3247), .ZN(n3246) );
  OR2X1 U3402 ( .IN1(n503), .IN2(n3378), .Q(n918) );
  AND2X1 U3403 ( .IN1(n3379), .IN2(n3179), .Q(n3378) );
  OR2X1 U3404 ( .IN1(g1840), .IN2(n3380), .Q(n3179) );
  OR2X1 U3405 ( .IN1(n1655), .IN2(n1608), .Q(n3380) );
  OR2X1 U3406 ( .IN1(n3381), .IN2(n1682), .Q(n3379) );
  AND2X1 U3407 ( .IN1(n1643), .IN2(n1605), .Q(n3381) );
  AND2X1 U3408 ( .IN1(n2857), .IN2(n3247), .Q(n3377) );
  OR2X1 U3409 ( .IN1(n3382), .IN2(n250), .Q(n3247) );
  AND2X1 U3410 ( .IN1(n926), .IN2(g1840), .Q(n3382) );
  OR2X1 U3411 ( .IN1(n3383), .IN2(n3232), .Q(g8920) );
  AND2X1 U3412 ( .IN1(n3384), .IN2(n3234), .Q(n3383) );
  XNOR2X1 U3413 ( .IN1(n931), .IN2(g713), .Q(n3384) );
  OR2X1 U3414 ( .IN1(n3385), .IN2(n3237), .Q(n931) );
  AND2X1 U3415 ( .IN1(n3386), .IN2(n3387), .Q(n3385) );
  OR2X1 U3416 ( .IN1(n2796), .IN2(n3388), .Q(n3387) );
  AND2X1 U3417 ( .IN1(n3389), .IN2(n3361), .Q(n3386) );
  OR2X1 U3418 ( .IN1(g704), .IN2(n3390), .Q(n3361) );
  OR2X1 U3419 ( .IN1(n3369), .IN2(n2696), .Q(n3389) );
  OR2X1 U3420 ( .IN1(n3391), .IN2(n3232), .Q(g8889) );
  AND2X1 U3421 ( .IN1(n3392), .IN2(n3234), .Q(n3391) );
  XNOR2X1 U3422 ( .IN1(n45), .IN2(n2796), .Q(n3392) );
  AND2X1 U3423 ( .IN1(n3393), .IN2(n3348), .Q(n45) );
  INVX0 U3424 ( .INP(n3394), .ZN(n3393) );
  AND2X1 U3425 ( .IN1(n3395), .IN2(n3396), .Q(n3394) );
  OR2X1 U3426 ( .IN1(n3369), .IN2(n1719), .Q(n3396) );
  AND2X1 U3427 ( .IN1(n3388), .IN2(n3390), .Q(n3395) );
  OR2X1 U3428 ( .IN1(n3397), .IN2(n3398), .Q(n3390) );
  OR2X1 U3429 ( .IN1(g686), .IN2(g695), .Q(n3398) );
  OR2X1 U3430 ( .IN1(n3399), .IN2(n3400), .Q(n3388) );
  OR2X1 U3431 ( .IN1(n2850), .IN2(n1676), .Q(n3400) );
  OR2X1 U3432 ( .IN1(n3401), .IN2(n3232), .Q(g8887) );
  AND2X1 U3433 ( .IN1(n3402), .IN2(n3234), .Q(n3401) );
  XNOR2X1 U3434 ( .IN1(n2850), .IN2(n3403), .Q(n3402) );
  AND2X1 U3435 ( .IN1(n3404), .IN2(n3348), .Q(n3403) );
  OR2X1 U3436 ( .IN1(n3405), .IN2(n3406), .Q(n3404) );
  OR2X1 U3437 ( .IN1(n3407), .IN2(n3408), .Q(n3406) );
  AND2X1 U3438 ( .IN1(n3409), .IN2(n1676), .Q(n3408) );
  AND2X1 U3439 ( .IN1(n3410), .IN2(g686), .Q(n3407) );
  AND2X1 U3440 ( .IN1(n3238), .IN2(g700), .Q(n3405) );
  OR2X1 U3441 ( .IN1(n3411), .IN2(n3232), .Q(g8885) );
  AND2X1 U3442 ( .IN1(n3412), .IN2(n3234), .Q(n3411) );
  XNOR2X1 U3443 ( .IN1(n1676), .IN2(n3413), .Q(n3412) );
  AND2X1 U3444 ( .IN1(n3414), .IN2(n3348), .Q(n3413) );
  OR2X1 U3445 ( .IN1(n3415), .IN2(n3416), .Q(n3414) );
  OR2X1 U3446 ( .IN1(n3409), .IN2(n3410), .Q(n3416) );
  INVX0 U3447 ( .INP(n3399), .ZN(n3410) );
  OR2X1 U3448 ( .IN1(n3238), .IN2(n3417), .Q(n3399) );
  OR2X1 U3449 ( .IN1(n1656), .IN2(n3357), .Q(n3417) );
  INVX0 U3450 ( .INP(n3397), .ZN(n3409) );
  OR2X1 U3451 ( .IN1(n3238), .IN2(n3341), .Q(n3397) );
  OR2X1 U3452 ( .IN1(n3418), .IN2(g677), .Q(n3341) );
  AND2X1 U3453 ( .IN1(n3238), .IN2(g691), .Q(n3415) );
  INVX0 U3454 ( .INP(n3369), .ZN(n3238) );
  OR2X1 U3455 ( .IN1(n3419), .IN2(n3232), .Q(g8883) );
  INVX0 U3456 ( .INP(n3420), .ZN(n3232) );
  OR2X1 U3457 ( .IN1(n3421), .IN2(n3422), .Q(n3420) );
  OR2X1 U3458 ( .IN1(n3213), .IN2(n3139), .Q(n3422) );
  OR2X1 U3459 ( .IN1(n3234), .IN2(n3423), .Q(n3421) );
  INVX0 U3460 ( .INP(n3171), .ZN(n3423) );
  AND2X1 U3461 ( .IN1(n3234), .IN2(n3424), .Q(n3419) );
  XNOR2X1 U3462 ( .IN1(g677), .IN2(n3425), .Q(n3424) );
  AND2X1 U3463 ( .IN1(n3426), .IN2(n3427), .Q(n3425) );
  OR2X1 U3464 ( .IN1(n3428), .IN2(n3429), .Q(n3427) );
  INVX0 U3465 ( .INP(n3335), .ZN(n3429) );
  AND2X1 U3466 ( .IN1(n3348), .IN2(n3369), .Q(n3335) );
  INVX0 U3467 ( .INP(n3237), .ZN(n3348) );
  AND2X1 U3468 ( .IN1(n958), .IN2(n3369), .Q(n3237) );
  OR2X1 U3469 ( .IN1(n3430), .IN2(n3169), .Q(n958) );
  AND2X1 U3470 ( .IN1(n3431), .IN2(n3171), .Q(n3430) );
  OR2X1 U3471 ( .IN1(n3432), .IN2(n1692), .Q(n3431) );
  AND2X1 U3472 ( .IN1(n1644), .IN2(n1593), .Q(n3432) );
  AND2X1 U3473 ( .IN1(n3357), .IN2(n3418), .Q(n3428) );
  INVX0 U3474 ( .INP(n3433), .ZN(n3418) );
  AND2X1 U3475 ( .IN1(n1662), .IN2(n3434), .Q(n3433) );
  AND2X1 U3476 ( .IN1(n3435), .IN2(n1615), .Q(n3434) );
  OR2X1 U3477 ( .IN1(n3435), .IN2(n3436), .Q(n3357) );
  OR2X1 U3478 ( .IN1(n1662), .IN2(n1615), .Q(n3436) );
  INVX0 U3479 ( .INP(n3370), .ZN(n3435) );
  OR2X1 U3480 ( .IN1(n3437), .IN2(n3220), .Q(n3370) );
  AND2X1 U3481 ( .IN1(n3438), .IN2(n1593), .Q(n3220) );
  AND2X1 U3482 ( .IN1(n1644), .IN2(n3439), .Q(n3437) );
  OR2X1 U3483 ( .IN1(n2864), .IN2(n3369), .Q(n3426) );
  AND2X1 U3484 ( .IN1(n3440), .IN2(n3441), .Q(n3369) );
  OR2X1 U3485 ( .IN1(n3442), .IN2(n3215), .Q(g8820) );
  INVX0 U3486 ( .INP(n3167), .ZN(n3215) );
  OR2X1 U3487 ( .IN1(g622), .IN2(n3443), .Q(n3167) );
  OR2X1 U3488 ( .IN1(n3227), .IN2(n3171), .Q(n3443) );
  AND2X1 U3489 ( .IN1(n3444), .IN2(g622), .Q(n3442) );
  OR2X1 U3490 ( .IN1(n3445), .IN2(n3234), .Q(n3444) );
  AND2X1 U3491 ( .IN1(n3227), .IN2(n3446), .Q(n3234) );
  INVX0 U3492 ( .INP(n804), .ZN(n3227) );
  AND2X1 U3493 ( .IN1(n3446), .IN2(n3171), .Q(n3445) );
  OR2X1 U3494 ( .IN1(g617), .IN2(n3447), .Q(n3171) );
  OR2X1 U3495 ( .IN1(n1609), .IN2(n1607), .Q(n3447) );
  OR2X1 U3496 ( .IN1(n3448), .IN2(n3449), .Q(g8779) );
  AND2X1 U3497 ( .IN1(n3450), .IN2(n3451), .Q(n3449) );
  AND2X1 U3498 ( .IN1(n371), .IN2(g1636), .Q(n3448) );
  OR2X1 U3499 ( .IN1(n3452), .IN2(n3453), .Q(g8777) );
  AND2X1 U3500 ( .IN1(n3454), .IN2(n3451), .Q(n3453) );
  AND2X1 U3501 ( .IN1(n371), .IN2(g1633), .Q(n3452) );
  OR2X1 U3502 ( .IN1(n3455), .IN2(n3456), .Q(g8776) );
  AND2X1 U3503 ( .IN1(n3457), .IN2(n3451), .Q(n3456) );
  AND2X1 U3504 ( .IN1(n371), .IN2(g1630), .Q(n3455) );
  AND2X1 U3505 ( .IN1(n3458), .IN2(g109), .Q(g8775) );
  XNOR2X1 U3506 ( .IN1(n2829), .IN2(n3459), .Q(n3458) );
  OR2X1 U3507 ( .IN1(n3460), .IN2(n3461), .Q(g8774) );
  AND2X1 U3508 ( .IN1(n3459), .IN2(n3451), .Q(n3461) );
  OR2X1 U3509 ( .IN1(n3462), .IN2(n3463), .Q(n3459) );
  OR2X1 U3510 ( .IN1(n3464), .IN2(n3465), .Q(n3463) );
  AND2X1 U3511 ( .IN1(n3466), .IN2(n1706), .Q(n3465) );
  AND2X1 U3512 ( .IN1(n3467), .IN2(n3468), .Q(n3466) );
  AND2X1 U3513 ( .IN1(n1654), .IN2(g1107), .Q(n3467) );
  AND2X1 U3514 ( .IN1(n3469), .IN2(g1133), .Q(n3464) );
  AND2X1 U3515 ( .IN1(n3470), .IN2(n3471), .Q(n3469) );
  OR2X1 U3516 ( .IN1(n3472), .IN2(n3473), .Q(n3470) );
  OR2X1 U3517 ( .IN1(n1614), .IN2(g1101), .Q(n3473) );
  AND2X1 U3518 ( .IN1(n371), .IN2(g1627), .Q(n3460) );
  OR2X1 U3519 ( .IN1(n3474), .IN2(n3475), .Q(g8773) );
  AND2X1 U3520 ( .IN1(n3476), .IN2(n3451), .Q(n3475) );
  AND2X1 U3521 ( .IN1(n371), .IN2(g1624), .Q(n3474) );
  AND2X1 U3522 ( .IN1(n3477), .IN2(g109), .Q(g8772) );
  XNOR2X1 U3523 ( .IN1(n2830), .IN2(n3457), .Q(n3477) );
  OR2X1 U3524 ( .IN1(n3478), .IN2(n3479), .Q(n3457) );
  OR2X1 U3525 ( .IN1(n3480), .IN2(n3481), .Q(n3479) );
  AND2X1 U3526 ( .IN1(n3482), .IN2(n1597), .Q(n3481) );
  AND2X1 U3527 ( .IN1(n3483), .IN2(n3468), .Q(n3482) );
  AND2X1 U3528 ( .IN1(g1107), .IN2(g1101), .Q(n3483) );
  AND2X1 U3529 ( .IN1(n3484), .IN2(g1137), .Q(n3480) );
  AND2X1 U3530 ( .IN1(n3485), .IN2(n3471), .Q(n3484) );
  OR2X1 U3531 ( .IN1(n3472), .IN2(n3486), .Q(n3485) );
  OR2X1 U3532 ( .IN1(n1654), .IN2(n1614), .Q(n3486) );
  OR2X1 U3533 ( .IN1(n3487), .IN2(n3488), .Q(g8771) );
  AND2X1 U3534 ( .IN1(n3489), .IN2(n3451), .Q(n3488) );
  AND2X1 U3535 ( .IN1(n371), .IN2(g1621), .Q(n3487) );
  OR2X1 U3536 ( .IN1(n3490), .IN2(n3491), .Q(g8770) );
  AND2X1 U3537 ( .IN1(n3492), .IN2(n3451), .Q(n3491) );
  AND2X1 U3538 ( .IN1(n371), .IN2(g1615), .Q(n3490) );
  AND2X1 U3539 ( .IN1(n3493), .IN2(g109), .Q(g8769) );
  XNOR2X1 U3540 ( .IN1(n2831), .IN2(n3492), .Q(n3493) );
  OR2X1 U3541 ( .IN1(n3494), .IN2(n3495), .Q(n3492) );
  OR2X1 U3542 ( .IN1(n3496), .IN2(n3497), .Q(n3495) );
  AND2X1 U3543 ( .IN1(n3498), .IN2(n1618), .Q(n3497) );
  AND2X1 U3544 ( .IN1(n3468), .IN2(n3499), .Q(n3498) );
  AND2X1 U3545 ( .IN1(n3471), .IN2(n3500), .Q(n3468) );
  AND2X1 U3546 ( .IN1(n3501), .IN2(g1121), .Q(n3496) );
  AND2X1 U3547 ( .IN1(n3502), .IN2(n3471), .Q(n3501) );
  OR2X1 U3548 ( .IN1(n3503), .IN2(n3472), .Q(n3502) );
  INVX0 U3549 ( .INP(n3500), .ZN(n3472) );
  AND2X1 U3550 ( .IN1(n3504), .IN2(g109), .Q(g8768) );
  XNOR2X1 U3551 ( .IN1(n2832), .IN2(n3454), .Q(n3504) );
  OR2X1 U3552 ( .IN1(n3505), .IN2(n3506), .Q(n3454) );
  AND2X1 U3553 ( .IN1(n3507), .IN2(n3471), .Q(n3505) );
  XNOR2X1 U3554 ( .IN1(n1660), .IN2(n3508), .Q(n3507) );
  AND2X1 U3555 ( .IN1(n3509), .IN2(n1658), .Q(n3508) );
  AND2X1 U3556 ( .IN1(n3510), .IN2(g109), .Q(g8767) );
  XNOR2X1 U3557 ( .IN1(n2773), .IN2(n3489), .Q(n3510) );
  OR2X1 U3558 ( .IN1(n3511), .IN2(n3512), .Q(n3489) );
  AND2X1 U3559 ( .IN1(n3513), .IN2(n3471), .Q(n3511) );
  XOR2X1 U3560 ( .IN1(n3514), .IN2(n1708), .Q(n3513) );
  OR2X1 U3561 ( .IN1(g1101), .IN2(n3515), .Q(n3514) );
  AND2X1 U3562 ( .IN1(n3516), .IN2(g109), .Q(g8766) );
  XNOR2X1 U3563 ( .IN1(n2771), .IN2(n3450), .Q(n3516) );
  OR2X1 U3564 ( .IN1(n3517), .IN2(n3518), .Q(n3450) );
  AND2X1 U3565 ( .IN1(n3519), .IN2(n3471), .Q(n3517) );
  XNOR2X1 U3566 ( .IN1(n3520), .IN2(g1145), .Q(n3519) );
  OR2X1 U3567 ( .IN1(n1677), .IN2(n3521), .Q(n3520) );
  AND2X1 U3568 ( .IN1(n3522), .IN2(g109), .Q(g8765) );
  XNOR2X1 U3569 ( .IN1(n2772), .IN2(n3476), .Q(n3522) );
  OR2X1 U3570 ( .IN1(n3523), .IN2(n3524), .Q(n3476) );
  AND2X1 U3571 ( .IN1(n3525), .IN2(n3471), .Q(n3523) );
  XOR2X1 U3572 ( .IN1(n3526), .IN2(n1705), .Q(n3525) );
  OR2X1 U3573 ( .IN1(n1654), .IN2(n3515), .Q(n3526) );
  OR2X1 U3574 ( .IN1(g1110), .IN2(n3527), .Q(n3515) );
  OR2X1 U3575 ( .IN1(n1614), .IN2(g1104), .Q(n3527) );
  OR2X1 U3576 ( .IN1(n3528), .IN2(n3529), .Q(g8649) );
  INVX0 U3577 ( .INP(n3530), .ZN(n3529) );
  AND2X1 U3578 ( .IN1(n3446), .IN2(n3531), .Q(n3530) );
  AND2X1 U3579 ( .IN1(n1016), .IN2(g664), .Q(n3528) );
  OR2X1 U3580 ( .IN1(n3532), .IN2(n3533), .Q(g8631) );
  AND2X1 U3581 ( .IN1(n3534), .IN2(n3446), .Q(n3533) );
  OR2X1 U3582 ( .IN1(n3535), .IN2(n3536), .Q(n3534) );
  AND2X1 U3583 ( .IN1(n3537), .IN2(g636), .Q(n3536) );
  OR2X1 U3584 ( .IN1(n3538), .IN2(n3539), .Q(n3537) );
  OR2X1 U3585 ( .IN1(n3540), .IN2(n3151), .Q(n3539) );
  OR2X1 U3586 ( .IN1(n2900), .IN2(n1874), .Q(n3151) );
  AND2X1 U3587 ( .IN1(n3541), .IN2(n3542), .Q(n3540) );
  AND2X1 U3588 ( .IN1(n3543), .IN2(n3229), .Q(n3542) );
  AND2X1 U3589 ( .IN1(n1609), .IN2(n1644), .Q(n3541) );
  XOR2X1 U3590 ( .IN1(n3544), .IN2(n3545), .Q(n3538) );
  AND2X1 U3591 ( .IN1(g255), .IN2(g622), .Q(n3545) );
  OR2X1 U3592 ( .IN1(n3546), .IN2(n3547), .Q(n3544) );
  AND2X1 U3593 ( .IN1(n3548), .IN2(n1692), .Q(n3547) );
  AND2X1 U3594 ( .IN1(n1609), .IN2(n3229), .Q(n3548) );
  INVX0 U3595 ( .INP(n3221), .ZN(n3229) );
  AND2X1 U3596 ( .IN1(n3228), .IN2(g639), .Q(n3546) );
  INVX0 U3597 ( .INP(n3438), .ZN(n3228) );
  AND2X1 U3598 ( .IN1(n3219), .IN2(n1713), .Q(n3535) );
  AND2X1 U3599 ( .IN1(n3213), .IN2(n3549), .Q(n3532) );
  OR2X1 U3600 ( .IN1(n3550), .IN2(n3551), .Q(n3549) );
  OR2X1 U3601 ( .IN1(n1716), .IN2(n3552), .Q(n3551) );
  AND2X1 U3602 ( .IN1(n3553), .IN2(n3554), .Q(n3552) );
  OR2X1 U3603 ( .IN1(n2847), .IN2(n2858), .Q(n3554) );
  OR2X1 U3604 ( .IN1(n2846), .IN2(n2855), .Q(n3553) );
  AND2X1 U3605 ( .IN1(n3555), .IN2(n3556), .Q(n3550) );
  OR2X1 U3606 ( .IN1(n1622), .IN2(n2859), .Q(n3555) );
  OR2X1 U3607 ( .IN1(n3557), .IN2(n3558), .Q(g8566) );
  AND2X1 U3608 ( .IN1(g1690), .IN2(g1687), .Q(n3558) );
  AND2X1 U3609 ( .IN1(n1653), .IN2(g1669), .Q(n3557) );
  OR2X1 U3610 ( .IN1(n3559), .IN2(n3560), .Q(g8565) );
  AND2X1 U3611 ( .IN1(g1690), .IN2(g1684), .Q(n3560) );
  AND2X1 U3612 ( .IN1(n1653), .IN2(g1666), .Q(n3559) );
  OR2X1 U3613 ( .IN1(n3561), .IN2(n3562), .Q(g8564) );
  AND2X1 U3614 ( .IN1(g1690), .IN2(g1681), .Q(n3562) );
  AND2X1 U3615 ( .IN1(n1653), .IN2(g1663), .Q(n3561) );
  OR2X1 U3616 ( .IN1(n3563), .IN2(n3564), .Q(g8563) );
  AND2X1 U3617 ( .IN1(g1690), .IN2(g1678), .Q(n3564) );
  AND2X1 U3618 ( .IN1(n1653), .IN2(g1660), .Q(n3563) );
  OR2X1 U3619 ( .IN1(n3565), .IN2(n3566), .Q(g8562) );
  AND2X1 U3620 ( .IN1(g1690), .IN2(g1675), .Q(n3566) );
  AND2X1 U3621 ( .IN1(n1653), .IN2(g1657), .Q(n3565) );
  OR2X1 U3622 ( .IN1(n3567), .IN2(n3568), .Q(g8561) );
  AND2X1 U3623 ( .IN1(g1690), .IN2(g1672), .Q(n3568) );
  AND2X1 U3624 ( .IN1(n1653), .IN2(g1654), .Q(n3567) );
  OR2X1 U3625 ( .IN1(n3569), .IN2(n3570), .Q(g8559) );
  OR2X1 U3626 ( .IN1(n3571), .IN2(n3572), .Q(n3570) );
  AND2X1 U3627 ( .IN1(n3573), .IN2(g1878), .Q(n3572) );
  AND2X1 U3628 ( .IN1(g18), .IN2(n3574), .Q(g8505) );
  XNOR2X1 U3629 ( .IN1(g617), .IN2(n3575), .Q(n3574) );
  AND2X1 U3630 ( .IN1(n3440), .IN2(n3531), .Q(n3575) );
  OR2X1 U3631 ( .IN1(n2808), .IN2(n1016), .Q(n3531) );
  OR2X1 U3632 ( .IN1(n3576), .IN2(n3577), .Q(n3440) );
  OR2X1 U3633 ( .IN1(n3543), .IN2(g611), .Q(n3577) );
  OR2X1 U3634 ( .IN1(g617), .IN2(n3578), .Q(n3543) );
  OR2X1 U3635 ( .IN1(n1607), .IN2(g605), .Q(n3578) );
  OR2X1 U3636 ( .IN1(g599), .IN2(n3169), .Q(n3576) );
  OR2X1 U3637 ( .IN1(n3579), .IN2(n3580), .Q(g8435) );
  AND2X1 U3638 ( .IN1(n3581), .IN2(g727), .Q(n3580) );
  AND2X1 U3639 ( .IN1(n3582), .IN2(g736), .Q(n3579) );
  OR2X1 U3640 ( .IN1(n3583), .IN2(n3584), .Q(g8434) );
  AND2X1 U3641 ( .IN1(n3581), .IN2(g718), .Q(n3584) );
  AND2X1 U3642 ( .IN1(n3582), .IN2(g727), .Q(n3583) );
  OR2X1 U3643 ( .IN1(n3585), .IN2(n3586), .Q(g8433) );
  AND2X1 U3644 ( .IN1(n3581), .IN2(g709), .Q(n3586) );
  AND2X1 U3645 ( .IN1(n3582), .IN2(g718), .Q(n3585) );
  OR2X1 U3646 ( .IN1(n3587), .IN2(n3588), .Q(g8432) );
  AND2X1 U3647 ( .IN1(n3581), .IN2(g700), .Q(n3588) );
  AND2X1 U3648 ( .IN1(n3582), .IN2(g709), .Q(n3587) );
  OR2X1 U3649 ( .IN1(n3589), .IN2(n3590), .Q(g8431) );
  AND2X1 U3650 ( .IN1(n3581), .IN2(g691), .Q(n3590) );
  AND2X1 U3651 ( .IN1(n3582), .IN2(g700), .Q(n3589) );
  OR2X1 U3652 ( .IN1(n3591), .IN2(n3592), .Q(g8430) );
  AND2X1 U3653 ( .IN1(n3581), .IN2(g682), .Q(n3592) );
  AND2X1 U3654 ( .IN1(n3582), .IN2(g691), .Q(n3591) );
  OR2X1 U3655 ( .IN1(n3593), .IN2(n3594), .Q(g8429) );
  AND2X1 U3656 ( .IN1(n3581), .IN2(g673), .Q(n3594) );
  AND2X1 U3657 ( .IN1(n3582), .IN2(g682), .Q(n3593) );
  OR2X1 U3658 ( .IN1(n3595), .IN2(n3596), .Q(g8428) );
  AND2X1 U3659 ( .IN1(n3581), .IN2(g664), .Q(n3596) );
  INVX0 U3660 ( .INP(n1016), .ZN(n3581) );
  AND2X1 U3661 ( .IN1(n3582), .IN2(g673), .Q(n3595) );
  AND2X1 U3662 ( .IN1(n3446), .IN2(n1016), .Q(n3582) );
  OR2X1 U3663 ( .IN1(g611), .IN2(n3441), .Q(n1016) );
  OR2X1 U3664 ( .IN1(n1645), .IN2(n3169), .Q(n3441) );
  AND2X1 U3665 ( .IN1(g18), .IN2(n3597), .Q(g8384) );
  XNOR2X1 U3666 ( .IN1(n2809), .IN2(n3598), .Q(n3597) );
  OR2X1 U3667 ( .IN1(n3571), .IN2(n250), .Q(n3598) );
  INVX0 U3668 ( .INP(n3599), .ZN(n250) );
  OR2X1 U3669 ( .IN1(n3600), .IN2(n3601), .Q(n3599) );
  OR2X1 U3670 ( .IN1(n503), .IN2(g1822), .Q(n3601) );
  AND2X1 U3671 ( .IN1(n3602), .IN2(g1950), .Q(n3571) );
  OR2X1 U3672 ( .IN1(g82), .IN2(g8986), .Q(g8352) );
  OR2X1 U3673 ( .IN1(g82), .IN2(g8985), .Q(g8349) );
  OR2X1 U3674 ( .IN1(g82), .IN2(g8976), .Q(g8347) );
  OR2X1 U3675 ( .IN1(g82), .IN2(test_so10), .Q(g8340) );
  OR2X1 U3676 ( .IN1(g82), .IN2(g8983), .Q(g8335) );
  OR2X1 U3677 ( .IN1(g82), .IN2(g8982), .Q(g8331) );
  OR2X1 U3678 ( .IN1(g82), .IN2(g8981), .Q(g8328) );
  OR2X1 U3679 ( .IN1(g82), .IN2(g8980), .Q(g8323) );
  OR2X1 U3680 ( .IN1(g82), .IN2(g8979), .Q(g8318) );
  OR2X1 U3681 ( .IN1(g82), .IN2(g8978), .Q(g8316) );
  OR2X1 U3682 ( .IN1(g82), .IN2(g8977), .Q(g8313) );
  OR2X1 U3683 ( .IN1(n3603), .IN2(n3604), .Q(g8288) );
  AND2X1 U3684 ( .IN1(n3602), .IN2(g1941), .Q(n3604) );
  AND2X1 U3685 ( .IN1(n3605), .IN2(g1950), .Q(n3603) );
  OR2X1 U3686 ( .IN1(n3606), .IN2(n3607), .Q(g8287) );
  AND2X1 U3687 ( .IN1(n3602), .IN2(g1932), .Q(n3607) );
  AND2X1 U3688 ( .IN1(n3605), .IN2(g1941), .Q(n3606) );
  OR2X1 U3689 ( .IN1(n3608), .IN2(n3609), .Q(g8286) );
  AND2X1 U3690 ( .IN1(n3602), .IN2(g1923), .Q(n3609) );
  AND2X1 U3691 ( .IN1(n3605), .IN2(g1932), .Q(n3608) );
  OR2X1 U3692 ( .IN1(n3610), .IN2(n3611), .Q(g8285) );
  AND2X1 U3693 ( .IN1(n3602), .IN2(g1914), .Q(n3611) );
  AND2X1 U3694 ( .IN1(n3605), .IN2(g1923), .Q(n3610) );
  OR2X1 U3695 ( .IN1(n3612), .IN2(n3613), .Q(g8284) );
  AND2X1 U3696 ( .IN1(n3602), .IN2(g1905), .Q(n3613) );
  AND2X1 U3697 ( .IN1(n3605), .IN2(g1914), .Q(n3612) );
  OR2X1 U3698 ( .IN1(n3614), .IN2(n3615), .Q(g8283) );
  AND2X1 U3699 ( .IN1(n3602), .IN2(g1896), .Q(n3615) );
  AND2X1 U3700 ( .IN1(n3605), .IN2(g1905), .Q(n3614) );
  OR2X1 U3701 ( .IN1(n3616), .IN2(n3617), .Q(g8282) );
  AND2X1 U3702 ( .IN1(n3602), .IN2(g1887), .Q(n3617) );
  AND2X1 U3703 ( .IN1(n3605), .IN2(g1896), .Q(n3616) );
  OR2X1 U3704 ( .IN1(n3618), .IN2(n3619), .Q(g8281) );
  AND2X1 U3705 ( .IN1(n3602), .IN2(g1878), .Q(n3619) );
  INVX0 U3706 ( .INP(n3573), .ZN(n3602) );
  AND2X1 U3707 ( .IN1(n3605), .IN2(g1887), .Q(n3618) );
  AND2X1 U3708 ( .IN1(n3188), .IN2(n3573), .Q(n3605) );
  OR2X1 U3709 ( .IN1(g1834), .IN2(n3620), .Q(n3573) );
  OR2X1 U3710 ( .IN1(n2809), .IN2(n503), .Q(n3620) );
  AND2X1 U3711 ( .IN1(n3621), .IN2(g940), .Q(g8260) );
  AND2X1 U3712 ( .IN1(n3621), .IN2(g936), .Q(g8254) );
  AND2X1 U3713 ( .IN1(n3621), .IN2(g932), .Q(g8250) );
  AND2X1 U3714 ( .IN1(n3622), .IN2(n3623), .Q(g8245) );
  XOR2X1 U3715 ( .IN1(n3624), .IN2(n1716), .Q(n3622) );
  OR2X1 U3716 ( .IN1(n2855), .IN2(n3625), .Q(n3624) );
  INVX0 U3717 ( .INP(n1090), .ZN(n3625) );
  AND2X1 U3718 ( .IN1(n3626), .IN2(n3627), .Q(g8244) );
  AND2X1 U3719 ( .IN1(n3628), .IN2(n3629), .Q(n3626) );
  INVX0 U3720 ( .INP(n3630), .ZN(n3628) );
  AND2X1 U3721 ( .IN1(n3631), .IN2(n2865), .Q(n3630) );
  OR2X1 U3722 ( .IN1(n3632), .IN2(n2883), .Q(n3631) );
  OR2X1 U3723 ( .IN1(n3633), .IN2(n3634), .Q(g8194) );
  AND2X1 U3724 ( .IN1(n3635), .IN2(n3451), .Q(n3634) );
  XNOR2X1 U3725 ( .IN1(n5138), .IN2(n3636), .Q(n3635) );
  AND2X1 U3726 ( .IN1(n3509), .IN2(g1104), .Q(n3636) );
  AND2X1 U3727 ( .IN1(g1110), .IN2(n3637), .Q(n3509) );
  AND2X1 U3728 ( .IN1(n371), .IN2(g1512), .Q(n3633) );
  OR2X1 U3729 ( .IN1(n3638), .IN2(n3639), .Q(g8193) );
  AND2X1 U3730 ( .IN1(n3640), .IN2(n3451), .Q(n3639) );
  XNOR2X1 U3731 ( .IN1(n2906), .IN2(n3641), .Q(n3640) );
  AND2X1 U3732 ( .IN1(n3500), .IN2(n3637), .Q(n3641) );
  AND2X1 U3733 ( .IN1(n1614), .IN2(n1654), .Q(n3637) );
  AND2X1 U3734 ( .IN1(g1104), .IN2(n1677), .Q(n3500) );
  AND2X1 U3735 ( .IN1(n371), .IN2(g1639), .Q(n3638) );
  AND2X1 U3736 ( .IN1(n1610), .IN2(n3642), .Q(g8173) );
  OR2X1 U3737 ( .IN1(n3643), .IN2(n3644), .Q(n3642) );
  AND2X1 U3738 ( .IN1(n3645), .IN2(g1806), .Q(n3644) );
  OR2X1 U3739 ( .IN1(n369), .IN2(n1055), .Q(n3645) );
  AND2X1 U3740 ( .IN1(n3646), .IN2(n1056), .Q(n3643) );
  AND2X1 U3741 ( .IN1(n1055), .IN2(g1801), .Q(n3646) );
  OR2X1 U3742 ( .IN1(n3162), .IN2(n3647), .Q(n1055) );
  OR2X1 U3743 ( .IN1(n2841), .IN2(n2840), .Q(n3647) );
  OR2X1 U3744 ( .IN1(n1626), .IN2(n3648), .Q(n3162) );
  AND2X1 U3745 ( .IN1(n3621), .IN2(g928), .Q(g8147) );
  AND2X1 U3746 ( .IN1(g109), .IN2(n3649), .Q(n3621) );
  INVX0 U3747 ( .INP(n3650), .ZN(n3649) );
  AND2X1 U3748 ( .IN1(n3651), .IN2(n3652), .Q(n3650) );
  AND2X1 U3749 ( .IN1(n3653), .IN2(DFF_436_n1), .Q(n3651) );
  AND2X1 U3750 ( .IN1(n3654), .IN2(g109), .Q(g8060) );
  XNOR2X1 U3751 ( .IN1(n2767), .IN2(g6002), .Q(n3654) );
  AND2X1 U3752 ( .IN1(n3655), .IN2(g109), .Q(g8059) );
  XNOR2X1 U3753 ( .IN1(n2764), .IN2(g6042), .Q(n3655) );
  AND2X1 U3754 ( .IN1(n3656), .IN2(g109), .Q(g8055) );
  XOR2X1 U3755 ( .IN1(g1490), .IN2(n3657), .Q(n3656) );
  AND2X1 U3756 ( .IN1(n3658), .IN2(g109), .Q(g8054) );
  XNOR2X1 U3757 ( .IN1(n2842), .IN2(g6015), .Q(n3658) );
  AND2X1 U3758 ( .IN1(n3659), .IN2(g109), .Q(g8053) );
  XNOR2X1 U3759 ( .IN1(n2763), .IN2(g6045), .Q(n3659) );
  AND2X1 U3760 ( .IN1(n3660), .IN2(g109), .Q(g8052) );
  XNOR2X1 U3761 ( .IN1(n2765), .IN2(n3661), .Q(n3660) );
  AND2X1 U3762 ( .IN1(n3662), .IN2(g109), .Q(g8051) );
  XNOR2X1 U3763 ( .IN1(n2769), .IN2(n3663), .Q(n3662) );
  AND2X1 U3764 ( .IN1(n3664), .IN2(g109), .Q(g8050) );
  XNOR2X1 U3765 ( .IN1(n2843), .IN2(g6026), .Q(n3664) );
  AND2X1 U3766 ( .IN1(n3665), .IN2(g109), .Q(g8049) );
  XNOR2X1 U3767 ( .IN1(n2766), .IN2(g6049), .Q(n3665) );
  AND2X1 U3768 ( .IN1(n3666), .IN2(g109), .Q(g8048) );
  XNOR2X1 U3769 ( .IN1(n2789), .IN2(g5996), .Q(n3666) );
  AND2X1 U3770 ( .IN1(n3667), .IN2(g109), .Q(g8047) );
  XNOR2X1 U3771 ( .IN1(n1704), .IN2(g6035), .Q(n3667) );
  AND2X1 U3772 ( .IN1(n3668), .IN2(g109), .Q(g8046) );
  XNOR2X1 U3773 ( .IN1(n2770), .IN2(n3669), .Q(n3668) );
  AND2X1 U3774 ( .IN1(n3670), .IN2(g109), .Q(g8045) );
  XNOR2X1 U3775 ( .IN1(n2834), .IN2(n3671), .Q(n3670) );
  AND2X1 U3776 ( .IN1(n3672), .IN2(g109), .Q(g8044) );
  XNOR2X1 U3777 ( .IN1(n2762), .IN2(g6038), .Q(n3672) );
  AND2X1 U3778 ( .IN1(n3673), .IN2(g109), .Q(g8043) );
  XNOR2X1 U3779 ( .IN1(n2835), .IN2(n3674), .Q(n3673) );
  AND2X1 U3780 ( .IN1(n3675), .IN2(g109), .Q(g8042) );
  XNOR2X1 U3781 ( .IN1(n1703), .IN2(n3676), .Q(n3675) );
  AND2X1 U3782 ( .IN1(n3677), .IN2(g109), .Q(g8041) );
  XNOR2X1 U3783 ( .IN1(n2801), .IN2(n3678), .Q(n3677) );
  AND2X1 U3784 ( .IN1(n3679), .IN2(g109), .Q(g8040) );
  XNOR2X1 U3785 ( .IN1(n2802), .IN2(n3680), .Q(n3679) );
  AND2X1 U3786 ( .IN1(n3681), .IN2(g109), .Q(g8039) );
  XNOR2X1 U3787 ( .IN1(n2803), .IN2(n3682), .Q(n3681) );
  AND2X1 U3788 ( .IN1(n3683), .IN2(n3623), .Q(g8024) );
  XNOR2X1 U3789 ( .IN1(n1090), .IN2(n2855), .Q(n3683) );
  AND2X1 U3790 ( .IN1(n3684), .IN2(n3627), .Q(g8019) );
  XNOR2X1 U3791 ( .IN1(n2883), .IN2(n1093), .Q(n3684) );
  AND2X1 U3792 ( .IN1(n3685), .IN2(n1610), .Q(g7930) );
  XNOR2X1 U3793 ( .IN1(n1056), .IN2(n2840), .Q(n3685) );
  AND2X1 U3794 ( .IN1(n3686), .IN2(g109), .Q(g7843) );
  XNOR2X1 U3795 ( .IN1(n2768), .IN2(g6000), .Q(n3686) );
  AND2X1 U3796 ( .IN1(n3687), .IN2(n3623), .Q(g7709) );
  INVX0 U3797 ( .INP(n3688), .ZN(n3687) );
  OR2X1 U3798 ( .IN1(n1090), .IN2(n1096), .Q(n3688) );
  INVX0 U3799 ( .INP(n3689), .ZN(g7705) );
  OR2X1 U3800 ( .IN1(n3690), .IN2(n3691), .Q(n3689) );
  OR2X1 U3801 ( .IN1(n1093), .IN2(n1098), .Q(n3690) );
  OR2X1 U3802 ( .IN1(n3692), .IN2(n3693), .Q(g7660) );
  OR2X1 U3803 ( .IN1(n3694), .IN2(n3213), .Q(n3693) );
  INVX0 U3804 ( .INP(n3695), .ZN(n3692) );
  OR2X1 U3805 ( .IN1(n3696), .IN2(n2836), .Q(n3695) );
  AND2X1 U3806 ( .IN1(n3697), .IN2(n3698), .Q(g7632) );
  AND2X1 U3807 ( .IN1(n3699), .IN2(n3700), .Q(n3697) );
  INVX0 U3808 ( .INP(n3701), .ZN(n3699) );
  AND2X1 U3809 ( .IN1(n3702), .IN2(n2887), .Q(n3701) );
  OR2X1 U3810 ( .IN1(n3213), .IN2(n3703), .Q(g7626) );
  OR2X1 U3811 ( .IN1(n3704), .IN2(n3705), .Q(n3703) );
  AND2X1 U3812 ( .IN1(n3706), .IN2(n1692), .Q(n3705) );
  AND2X1 U3813 ( .IN1(n3694), .IN2(n3707), .Q(n3706) );
  OR2X1 U3814 ( .IN1(n3139), .IN2(n3708), .Q(n3707) );
  OR2X1 U3815 ( .IN1(n3221), .IN2(n3438), .Q(n3708) );
  AND2X1 U3816 ( .IN1(g599), .IN2(n1607), .Q(n3438) );
  AND2X1 U3817 ( .IN1(g591), .IN2(g605), .Q(n3221) );
  OR2X1 U3818 ( .IN1(n3709), .IN2(n3219), .Q(n3139) );
  AND2X1 U3819 ( .IN1(n1644), .IN2(n3710), .Q(n3219) );
  AND2X1 U3820 ( .IN1(g605), .IN2(n1607), .Q(n3710) );
  AND2X1 U3821 ( .IN1(n1593), .IN2(g599), .Q(n3709) );
  AND2X1 U3822 ( .IN1(n3169), .IN2(g639), .Q(n3704) );
  AND2X1 U3823 ( .IN1(n3698), .IN2(n3711), .Q(g7590) );
  INVX0 U3824 ( .INP(n3712), .ZN(n3711) );
  AND2X1 U3825 ( .IN1(n3713), .IN2(n2881), .Q(n3712) );
  AND2X1 U3826 ( .IN1(n3698), .IN2(n3714), .Q(g7586) );
  OR2X1 U3827 ( .IN1(n3715), .IN2(n1107), .Q(n3714) );
  INVX0 U3828 ( .INP(n3716), .ZN(n1107) );
  OR2X1 U3829 ( .IN1(n3700), .IN2(n3717), .Q(n3716) );
  OR2X1 U3830 ( .IN1(n2651), .IN2(n3718), .Q(n3717) );
  INVX0 U3831 ( .INP(n3719), .ZN(n3718) );
  AND2X1 U3832 ( .IN1(n3713), .IN2(g1227), .Q(n3715) );
  OR2X1 U3833 ( .IN1(n3702), .IN2(n3720), .Q(n3713) );
  OR2X1 U3834 ( .IN1(n3721), .IN2(n3719), .Q(n3720) );
  AND2X1 U3835 ( .IN1(n3722), .IN2(n3698), .Q(g7581) );
  XOR2X1 U3836 ( .IN1(n3700), .IN2(n2651), .Q(n3722) );
  OR2X1 U3837 ( .IN1(n3702), .IN2(n3723), .Q(n3700) );
  OR2X1 U3838 ( .IN1(n2887), .IN2(n3721), .Q(n3723) );
  AND2X1 U3839 ( .IN1(n3724), .IN2(n1610), .Q(g7541) );
  AND2X1 U3840 ( .IN1(n3725), .IN2(n3726), .Q(n3724) );
  OR2X1 U3841 ( .IN1(n1626), .IN2(n3727), .Q(n3726) );
  INVX0 U3842 ( .INP(n1056), .ZN(n3727) );
  OR2X1 U3843 ( .IN1(n103), .IN2(g1796), .Q(n3725) );
  INVX0 U3844 ( .INP(n3728), .ZN(n103) );
  OR2X1 U3845 ( .IN1(n3729), .IN2(n3730), .Q(g7441) );
  OR2X1 U3846 ( .IN1(n3731), .IN2(n3213), .Q(n3730) );
  INVX0 U3847 ( .INP(n3732), .ZN(n3729) );
  OR2X1 U3848 ( .IN1(g627), .IN2(n1612), .Q(n3732) );
  OR2X1 U3849 ( .IN1(n3733), .IN2(n3734), .Q(g7303) );
  AND2X1 U3850 ( .IN1(n3735), .IN2(g1265), .Q(n3734) );
  AND2X1 U3851 ( .IN1(n3736), .IN2(test_so6), .Q(n3733) );
  OR2X1 U3852 ( .IN1(n3737), .IN2(n3738), .Q(g7302) );
  AND2X1 U3853 ( .IN1(n3735), .IN2(g1260), .Q(n3738) );
  AND2X1 U3854 ( .IN1(n3736), .IN2(g1265), .Q(n3737) );
  OR2X1 U3855 ( .IN1(n3739), .IN2(n3740), .Q(g7301) );
  AND2X1 U3856 ( .IN1(n3735), .IN2(g1255), .Q(n3740) );
  AND2X1 U3857 ( .IN1(n3736), .IN2(g1260), .Q(n3739) );
  OR2X1 U3858 ( .IN1(n3741), .IN2(n3742), .Q(g7300) );
  AND2X1 U3859 ( .IN1(n3735), .IN2(g1250), .Q(n3742) );
  AND2X1 U3860 ( .IN1(n3736), .IN2(g1255), .Q(n3741) );
  OR2X1 U3861 ( .IN1(n3743), .IN2(n3744), .Q(g7299) );
  AND2X1 U3862 ( .IN1(n3735), .IN2(g1245), .Q(n3744) );
  AND2X1 U3863 ( .IN1(n3736), .IN2(g1250), .Q(n3743) );
  OR2X1 U3864 ( .IN1(n3745), .IN2(n3746), .Q(g7298) );
  AND2X1 U3865 ( .IN1(n3735), .IN2(g1240), .Q(n3746) );
  AND2X1 U3866 ( .IN1(n3736), .IN2(g1245), .Q(n3745) );
  OR2X1 U3867 ( .IN1(n3747), .IN2(n3748), .Q(g7297) );
  AND2X1 U3868 ( .IN1(n3735), .IN2(g1235), .Q(n3748) );
  AND2X1 U3869 ( .IN1(n3736), .IN2(g1240), .Q(n3747) );
  OR2X1 U3870 ( .IN1(n3749), .IN2(n3750), .Q(g7296) );
  AND2X1 U3871 ( .IN1(n3735), .IN2(g1275), .Q(n3750) );
  AND2X1 U3872 ( .IN1(n3736), .IN2(g1235), .Q(n3749) );
  OR2X1 U3873 ( .IN1(n3751), .IN2(n3752), .Q(g7295) );
  AND2X1 U3874 ( .IN1(n3735), .IN2(g1284), .Q(n3752) );
  AND2X1 U3875 ( .IN1(n3736), .IN2(g1280), .Q(n3751) );
  OR2X1 U3876 ( .IN1(n3753), .IN2(n3754), .Q(g7294) );
  AND2X1 U3877 ( .IN1(n3735), .IN2(g1292), .Q(n3754) );
  AND2X1 U3878 ( .IN1(n3736), .IN2(g1284), .Q(n3753) );
  OR2X1 U3879 ( .IN1(n3755), .IN2(n3756), .Q(g7293) );
  AND2X1 U3880 ( .IN1(n3735), .IN2(g1296), .Q(n3756) );
  AND2X1 U3881 ( .IN1(n3736), .IN2(g1292), .Q(n3755) );
  OR2X1 U3882 ( .IN1(n3757), .IN2(n3758), .Q(g7292) );
  AND2X1 U3883 ( .IN1(n3735), .IN2(g1300), .Q(n3758) );
  AND2X1 U3884 ( .IN1(n3736), .IN2(g1296), .Q(n3757) );
  OR2X1 U3885 ( .IN1(n3759), .IN2(n3760), .Q(g7291) );
  AND2X1 U3886 ( .IN1(n3735), .IN2(g1304), .Q(n3760) );
  AND2X1 U3887 ( .IN1(n3736), .IN2(g1300), .Q(n3759) );
  OR2X1 U3888 ( .IN1(n3761), .IN2(n3762), .Q(g7290) );
  AND2X1 U3889 ( .IN1(n3735), .IN2(test_so6), .Q(n3762) );
  AND2X1 U3890 ( .IN1(n3736), .IN2(g1304), .Q(n3761) );
  OR2X1 U3891 ( .IN1(n3763), .IN2(n3764), .Q(g7257) );
  INVX0 U3892 ( .INP(n3765), .ZN(n3764) );
  OR2X1 U3893 ( .IN1(n3451), .IN2(n2888), .Q(n3765) );
  AND2X1 U3894 ( .IN1(n3451), .IN2(g1077), .Q(n3763) );
  OR2X1 U3895 ( .IN1(n3766), .IN2(n3767), .Q(g7244) );
  AND2X1 U3896 ( .IN1(n371), .IN2(g1023), .Q(n3767) );
  AND2X1 U3897 ( .IN1(n3451), .IN2(g1071), .Q(n3766) );
  OR2X1 U3898 ( .IN1(n3768), .IN2(test_so10), .Q(g7219) );
  OR2X1 U3899 ( .IN1(n3768), .IN2(g8982), .Q(g7204) );
  AND2X1 U3900 ( .IN1(n3769), .IN2(n3623), .Q(g7202) );
  XNOR2X1 U3901 ( .IN1(n1123), .IN2(n2858), .Q(n3769) );
  AND2X1 U3902 ( .IN1(n3770), .IN2(n3627), .Q(g7191) );
  XNOR2X1 U3903 ( .IN1(n1125), .IN2(n2869), .Q(n3770) );
  OR2X1 U3904 ( .IN1(n3768), .IN2(g8980), .Q(g7189) );
  OR2X1 U3905 ( .IN1(n3768), .IN2(g8978), .Q(g7183) );
  OR2X1 U3906 ( .IN1(n3768), .IN2(g8976), .Q(g7143) );
  AND2X1 U3907 ( .IN1(n3771), .IN2(n3772), .Q(g7137) );
  OR2X1 U3908 ( .IN1(n3773), .IN2(n3696), .Q(n3772) );
  INVX0 U3909 ( .INP(n3774), .ZN(n3773) );
  OR2X1 U3910 ( .IN1(n3775), .IN2(n1709), .Q(n3774) );
  AND2X1 U3911 ( .IN1(n3771), .IN2(n3776), .Q(g7134) );
  OR2X1 U3912 ( .IN1(n3777), .IN2(n3775), .Q(n3776) );
  INVX0 U3913 ( .INP(n3778), .ZN(n3777) );
  OR2X1 U3914 ( .IN1(n3731), .IN2(n5133), .Q(n3778) );
  AND2X1 U3915 ( .IN1(n3446), .IN2(n3169), .Q(n3771) );
  INVX0 U3916 ( .INP(n3694), .ZN(n3169) );
  AND2X1 U3917 ( .IN1(n3696), .IN2(n2836), .Q(n3694) );
  AND2X1 U3918 ( .IN1(n3775), .IN2(n1709), .Q(n3696) );
  AND2X1 U3919 ( .IN1(n3731), .IN2(n5133), .Q(n3775) );
  AND2X1 U3920 ( .IN1(g627), .IN2(n1612), .Q(n3731) );
  OR2X1 U3921 ( .IN1(n3779), .IN2(g1713), .Q(g7133) );
  AND2X1 U3922 ( .IN1(n3780), .IN2(n3781), .Q(n3779) );
  INVX0 U3923 ( .INP(n3782), .ZN(n3781) );
  OR2X1 U3924 ( .IN1(n2903), .IN2(g1766), .Q(n3780) );
  OR2X1 U3925 ( .IN1(n3783), .IN2(n145), .Q(g7032) );
  INVX0 U3926 ( .INP(n3784), .ZN(n145) );
  OR2X1 U3927 ( .IN1(n3785), .IN2(n3786), .Q(n3784) );
  OR2X1 U3928 ( .IN1(n3787), .IN2(n3788), .Q(n3786) );
  OR2X1 U3929 ( .IN1(n3789), .IN2(n3790), .Q(n3788) );
  OR2X1 U3930 ( .IN1(g143), .IN2(g148), .Q(n3790) );
  OR2X1 U3931 ( .IN1(g158), .IN2(g153), .Q(n3789) );
  OR2X1 U3932 ( .IN1(n3791), .IN2(n3792), .Q(n3787) );
  OR2X1 U3933 ( .IN1(g135), .IN2(g162), .Q(n3792) );
  OR2X1 U3934 ( .IN1(g131), .IN2(g139), .Q(n3791) );
  OR2X1 U3935 ( .IN1(n3793), .IN2(n3794), .Q(n3785) );
  OR2X1 U3936 ( .IN1(n3795), .IN2(n3796), .Q(n3794) );
  OR2X1 U3937 ( .IN1(g119), .IN2(g127), .Q(n3796) );
  OR2X1 U3938 ( .IN1(n3797), .IN2(n3798), .Q(n3795) );
  INVX0 U3939 ( .INP(g6786), .ZN(n3797) );
  OR2X1 U3940 ( .IN1(n3799), .IN2(n3800), .Q(n3793) );
  OR2X1 U3941 ( .IN1(n2788), .IN2(n2766), .Q(n3800) );
  OR2X1 U3942 ( .IN1(n2843), .IN2(n2842), .Q(n3799) );
  AND2X1 U3943 ( .IN1(g109), .IN2(g123), .Q(n3783) );
  AND2X1 U3944 ( .IN1(n1610), .IN2(n3801), .Q(g6983) );
  OR2X1 U3945 ( .IN1(n3802), .IN2(n3803), .Q(n3801) );
  AND2X1 U3946 ( .IN1(n3728), .IN2(g1791), .Q(n3803) );
  OR2X1 U3947 ( .IN1(n369), .IN2(n3648), .Q(n3728) );
  AND2X1 U3948 ( .IN1(n3804), .IN2(n2899), .Q(n3802) );
  AND2X1 U3949 ( .IN1(n3648), .IN2(g1786), .Q(n3804) );
  OR2X1 U3950 ( .IN1(n3805), .IN2(n3806), .Q(n3648) );
  OR2X1 U3951 ( .IN1(n1659), .IN2(n3807), .Q(n3806) );
  OR2X1 U3952 ( .IN1(n3808), .IN2(n3809), .Q(g6934) );
  AND2X1 U3953 ( .IN1(n3810), .IN2(g170), .Q(n3809) );
  AND2X1 U3954 ( .IN1(n3811), .IN2(g284), .Q(n3808) );
  OR2X1 U3955 ( .IN1(n3812), .IN2(n3813), .Q(g6930) );
  AND2X1 U3956 ( .IN1(n371), .IN2(g1015), .Q(n3813) );
  AND2X1 U3957 ( .IN1(n3451), .IN2(g1074), .Q(n3812) );
  OR2X1 U3958 ( .IN1(n3814), .IN2(n3815), .Q(g6929) );
  AND2X1 U3959 ( .IN1(n3810), .IN2(g143), .Q(n3815) );
  AND2X1 U3960 ( .IN1(n3811), .IN2(g302), .Q(n3814) );
  OR2X1 U3961 ( .IN1(n3816), .IN2(n3817), .Q(g6928) );
  AND2X1 U3962 ( .IN1(n3810), .IN2(g174), .Q(n3817) );
  AND2X1 U3963 ( .IN1(n3811), .IN2(g281), .Q(n3816) );
  OR2X1 U3964 ( .IN1(n3818), .IN2(n3819), .Q(g6924) );
  AND2X1 U3965 ( .IN1(n371), .IN2(g1019), .Q(n3819) );
  AND2X1 U3966 ( .IN1(n3451), .IN2(g1098), .Q(n3818) );
  OR2X1 U3967 ( .IN1(n3820), .IN2(n3821), .Q(g6923) );
  AND2X1 U3968 ( .IN1(n3810), .IN2(g166), .Q(n3821) );
  AND2X1 U3969 ( .IN1(n3811), .IN2(g299), .Q(n3820) );
  OR2X1 U3970 ( .IN1(n3822), .IN2(n3823), .Q(g6922) );
  AND2X1 U3971 ( .IN1(n3810), .IN2(g162), .Q(n3823) );
  AND2X1 U3972 ( .IN1(n3811), .IN2(g278), .Q(n3822) );
  OR2X1 U3973 ( .IN1(n3824), .IN2(n3825), .Q(g6918) );
  AND2X1 U3974 ( .IN1(test_so2), .IN2(n371), .Q(n3825) );
  AND2X1 U3975 ( .IN1(n3451), .IN2(g1095), .Q(n3824) );
  OR2X1 U3976 ( .IN1(n3826), .IN2(n3827), .Q(g6916) );
  AND2X1 U3977 ( .IN1(n3810), .IN2(g139), .Q(n3827) );
  AND2X1 U3978 ( .IN1(n3811), .IN2(g296), .Q(n3826) );
  OR2X1 U3979 ( .IN1(n3828), .IN2(n3829), .Q(g6915) );
  AND2X1 U3980 ( .IN1(n3810), .IN2(g158), .Q(n3829) );
  AND2X1 U3981 ( .IN1(n3811), .IN2(g275), .Q(n3828) );
  OR2X1 U3982 ( .IN1(n3830), .IN2(n3831), .Q(g6912) );
  AND2X1 U3983 ( .IN1(n371), .IN2(g1011), .Q(n3831) );
  AND2X1 U3984 ( .IN1(n3451), .IN2(g1092), .Q(n3830) );
  OR2X1 U3985 ( .IN1(n3832), .IN2(n3833), .Q(g6911) );
  AND2X1 U3986 ( .IN1(n3810), .IN2(g135), .Q(n3833) );
  AND2X1 U3987 ( .IN1(n3811), .IN2(g293), .Q(n3832) );
  OR2X1 U3988 ( .IN1(n3834), .IN2(n3835), .Q(g6910) );
  AND2X1 U3989 ( .IN1(n3810), .IN2(g153), .Q(n3835) );
  AND2X1 U3990 ( .IN1(n3811), .IN2(g272), .Q(n3834) );
  OR2X1 U3991 ( .IN1(n3836), .IN2(n3837), .Q(g6909) );
  INVX0 U3992 ( .INP(n3838), .ZN(n3837) );
  AND2X1 U3993 ( .IN1(n3839), .IN2(g1868), .Q(n3836) );
  OR2X1 U3994 ( .IN1(n3840), .IN2(n3841), .Q(g6908) );
  AND2X1 U3995 ( .IN1(test_so8), .IN2(n371), .Q(n3841) );
  AND2X1 U3996 ( .IN1(n3451), .IN2(g1089), .Q(n3840) );
  OR2X1 U3997 ( .IN1(n3842), .IN2(n3843), .Q(g6907) );
  AND2X1 U3998 ( .IN1(n3810), .IN2(g131), .Q(n3843) );
  AND2X1 U3999 ( .IN1(n3811), .IN2(g290), .Q(n3842) );
  OR2X1 U4000 ( .IN1(n3844), .IN2(n3845), .Q(g6906) );
  AND2X1 U4001 ( .IN1(n3810), .IN2(g148), .Q(n3845) );
  AND2X1 U4002 ( .IN1(n3811), .IN2(g269), .Q(n3844) );
  OR2X1 U4003 ( .IN1(n3846), .IN2(n3847), .Q(g6902) );
  AND2X1 U4004 ( .IN1(n371), .IN2(g1003), .Q(n3847) );
  AND2X1 U4005 ( .IN1(n3451), .IN2(g1086), .Q(n3846) );
  OR2X1 U4006 ( .IN1(n3848), .IN2(n3849), .Q(g6901) );
  AND2X1 U4007 ( .IN1(n3810), .IN2(g127), .Q(n3849) );
  AND2X1 U4008 ( .IN1(n3811), .IN2(g287), .Q(n3848) );
  OR2X1 U4009 ( .IN1(n3850), .IN2(n3851), .Q(g6900) );
  AND2X1 U4010 ( .IN1(n3810), .IN2(g178), .Q(n3851) );
  AND2X1 U4011 ( .IN1(n3811), .IN2(g266), .Q(n3850) );
  OR2X1 U4012 ( .IN1(n3852), .IN2(n3853), .Q(g6898) );
  INVX0 U4013 ( .INP(n3854), .ZN(n3853) );
  OR2X1 U4014 ( .IN1(n3451), .IN2(n1871), .Q(n3854) );
  AND2X1 U4015 ( .IN1(n3451), .IN2(g1083), .Q(n3852) );
  OR2X1 U4016 ( .IN1(n3855), .IN2(n3856), .Q(g6897) );
  INVX0 U4017 ( .INP(n3857), .ZN(n3856) );
  OR2X1 U4018 ( .IN1(n3811), .IN2(n2788), .Q(n3857) );
  AND2X1 U4019 ( .IN1(n3811), .IN2(g263), .Q(n3855) );
  INVX0 U4020 ( .INP(n3810), .ZN(n3811) );
  OR2X1 U4021 ( .IN1(n519), .IN2(n3858), .Q(n3810) );
  AND2X1 U4022 ( .IN1(n1613), .IN2(n1137), .Q(n3858) );
  INVX0 U4023 ( .INP(n3798), .ZN(n1137) );
  OR2X1 U4024 ( .IN1(n5134), .IN2(n3471), .Q(n3798) );
  OR2X1 U4025 ( .IN1(n3859), .IN2(n3860), .Q(g6895) );
  AND2X1 U4026 ( .IN1(n371), .IN2(g995), .Q(n3860) );
  AND2X1 U4027 ( .IN1(n3451), .IN2(g1080), .Q(n3859) );
  OR2X1 U4028 ( .IN1(n3861), .IN2(n3862), .Q(g6894) );
  AND2X1 U4029 ( .IN1(n371), .IN2(g1027), .Q(n3862) );
  AND2X1 U4030 ( .IN1(test_so7), .IN2(n3451), .Q(n3861) );
  AND2X1 U4031 ( .IN1(n3863), .IN2(n3864), .Q(g6842) );
  AND2X1 U4032 ( .IN1(g109), .IN2(g1400), .Q(g6841) );
  AND2X1 U4033 ( .IN1(g109), .IN2(g248), .Q(g6840) );
  AND2X1 U4034 ( .IN1(g109), .IN2(g1397), .Q(g6839) );
  INVX0 U4035 ( .INP(n3865), .ZN(g6834) );
  OR2X1 U4036 ( .IN1(n519), .IN2(n5136), .Q(n3865) );
  AND2X1 U4037 ( .IN1(g109), .IN2(n3019), .Q(g6830) );
  AND2X1 U4038 ( .IN1(g109), .IN2(n3038), .Q(g6828) );
  INVX0 U4039 ( .INP(n3866), .ZN(g6820) );
  OR2X1 U4040 ( .IN1(n519), .IN2(n5137), .Q(n3866) );
  AND2X1 U4041 ( .IN1(n3838), .IN2(n3867), .Q(g6795) );
  OR2X1 U4042 ( .IN1(n3868), .IN2(n1147), .Q(n3867) );
  INVX0 U4043 ( .INP(n3839), .ZN(n1147) );
  OR2X1 U4044 ( .IN1(g1861), .IN2(n3869), .Q(n3839) );
  OR2X1 U4045 ( .IN1(n5135), .IN2(g1864), .Q(n3869) );
  AND2X1 U4046 ( .IN1(n3870), .IN2(g1864), .Q(n3868) );
  OR2X1 U4047 ( .IN1(n5135), .IN2(g1861), .Q(n3870) );
  OR2X1 U4048 ( .IN1(n2902), .IN2(n3033), .Q(g6755) );
  AND2X1 U4049 ( .IN1(n3871), .IN2(n5134), .Q(g6747) );
  AND2X1 U4050 ( .IN1(n3872), .IN2(g109), .Q(n3871) );
  OR2X1 U4051 ( .IN1(n3041), .IN2(n3024), .Q(n3872) );
  AND2X1 U4052 ( .IN1(n3873), .IN2(n3623), .Q(g6733) );
  INVX0 U4053 ( .INP(n3874), .ZN(n3873) );
  OR2X1 U4054 ( .IN1(n1123), .IN2(n1150), .Q(n3874) );
  INVX0 U4055 ( .INP(n3875), .ZN(g6728) );
  OR2X1 U4056 ( .IN1(n3876), .IN2(n3691), .Q(n3875) );
  OR2X1 U4057 ( .IN1(n1125), .IN2(n1152), .Q(n3876) );
  OR2X1 U4058 ( .IN1(n3877), .IN2(n3878), .Q(g6679) );
  AND2X1 U4059 ( .IN1(g109), .IN2(g1), .Q(n3878) );
  AND2X1 U4060 ( .IN1(n1154), .IN2(n74), .Q(n3877) );
  INVX0 U4061 ( .INP(n3879), .ZN(n74) );
  OR2X1 U4062 ( .IN1(n3880), .IN2(n3881), .Q(n3879) );
  OR2X1 U4063 ( .IN1(n3882), .IN2(n3883), .Q(n3881) );
  OR2X1 U4064 ( .IN1(g1411), .IN2(g1403), .Q(n3883) );
  OR2X1 U4065 ( .IN1(g1415), .IN2(g1407), .Q(n3882) );
  OR2X1 U4066 ( .IN1(n3884), .IN2(n3885), .Q(n3880) );
  OR2X1 U4067 ( .IN1(n2830), .IN2(n2829), .Q(n3885) );
  OR2X1 U4068 ( .IN1(n2832), .IN2(n2831), .Q(n3884) );
  AND2X1 U4069 ( .IN1(n3886), .IN2(n3887), .Q(n1154) );
  AND2X1 U4070 ( .IN1(g6234), .IN2(n3888), .Q(n3887) );
  AND2X1 U4071 ( .IN1(g1419), .IN2(n1159), .Q(n3888) );
  INVX0 U4072 ( .INP(n3889), .ZN(n3886) );
  OR2X1 U4073 ( .IN1(n3890), .IN2(n3891), .Q(n3889) );
  OR2X1 U4074 ( .IN1(n1710), .IN2(n1627), .Q(n3891) );
  OR2X1 U4075 ( .IN1(n2772), .IN2(n2771), .Q(n3890) );
  OR2X1 U4076 ( .IN1(n3892), .IN2(n3893), .Q(g6656) );
  AND2X1 U4077 ( .IN1(g109), .IN2(g4), .Q(n3893) );
  AND2X1 U4078 ( .IN1(n1161), .IN2(n72), .Q(n3892) );
  INVX0 U4079 ( .INP(n3894), .ZN(n72) );
  OR2X1 U4080 ( .IN1(n3895), .IN2(n3896), .Q(n3894) );
  OR2X1 U4081 ( .IN1(n3897), .IN2(n3898), .Q(n3896) );
  OR2X1 U4082 ( .IN1(g1482), .IN2(g1499), .Q(n3898) );
  OR2X1 U4083 ( .IN1(g1486), .IN2(g1466), .Q(n3897) );
  OR2X1 U4084 ( .IN1(n3899), .IN2(n3900), .Q(n3895) );
  OR2X1 U4085 ( .IN1(n2833), .IN2(g1458), .Q(n3900) );
  OR2X1 U4086 ( .IN1(n2835), .IN2(n2834), .Q(n3899) );
  AND2X1 U4087 ( .IN1(n3901), .IN2(n3902), .Q(n1161) );
  AND2X1 U4088 ( .IN1(n1159), .IN2(n3903), .Q(n3902) );
  AND2X1 U4089 ( .IN1(g1453), .IN2(n2898), .Q(n3903) );
  AND2X1 U4090 ( .IN1(g1504), .IN2(g109), .Q(n2898) );
  INVX0 U4091 ( .INP(n3904), .ZN(n3901) );
  OR2X1 U4092 ( .IN1(n3905), .IN2(n3906), .Q(n3904) );
  OR2X1 U4093 ( .IN1(n2801), .IN2(n1707), .Q(n3906) );
  OR2X1 U4094 ( .IN1(n2803), .IN2(n2802), .Q(n3905) );
  AND2X1 U4095 ( .IN1(n3147), .IN2(g8983), .Q(g6653) );
  AND2X1 U4096 ( .IN1(n3147), .IN2(g8981), .Q(g6638) );
  AND2X1 U4097 ( .IN1(n3147), .IN2(g8979), .Q(g6627) );
  AND2X1 U4098 ( .IN1(n3147), .IN2(g8977), .Q(g6621) );
  OR2X1 U4099 ( .IN1(n3907), .IN2(n3908), .Q(g6551) );
  AND2X1 U4100 ( .IN1(n3909), .IN2(g1478), .Q(n3908) );
  AND2X1 U4101 ( .IN1(n3910), .IN2(g1546), .Q(n3907) );
  OR2X1 U4102 ( .IN1(n3911), .IN2(n3912), .Q(g6546) );
  AND2X1 U4103 ( .IN1(n3909), .IN2(g1453), .Q(n3912) );
  AND2X1 U4104 ( .IN1(n3910), .IN2(g1564), .Q(n3911) );
  OR2X1 U4105 ( .IN1(n3913), .IN2(n3914), .Q(g6545) );
  AND2X1 U4106 ( .IN1(n3909), .IN2(g1482), .Q(n3914) );
  AND2X1 U4107 ( .IN1(n3910), .IN2(g1543), .Q(n3913) );
  OR2X1 U4108 ( .IN1(n3915), .IN2(n3916), .Q(g6542) );
  AND2X1 U4109 ( .IN1(n3909), .IN2(g1458), .Q(n3916) );
  AND2X1 U4110 ( .IN1(n3910), .IN2(g1561), .Q(n3915) );
  OR2X1 U4111 ( .IN1(n3917), .IN2(n3918), .Q(g6541) );
  AND2X1 U4112 ( .IN1(n3909), .IN2(g1486), .Q(n3918) );
  AND2X1 U4113 ( .IN1(n3910), .IN2(g1540), .Q(n3917) );
  OR2X1 U4114 ( .IN1(n3919), .IN2(n3920), .Q(g6538) );
  AND2X1 U4115 ( .IN1(n3909), .IN2(g1462), .Q(n3920) );
  AND2X1 U4116 ( .IN1(n3910), .IN2(g1558), .Q(n3919) );
  OR2X1 U4117 ( .IN1(n3921), .IN2(n3922), .Q(g6537) );
  AND2X1 U4118 ( .IN1(n3909), .IN2(g1490), .Q(n3922) );
  AND2X1 U4119 ( .IN1(n3910), .IN2(g1537), .Q(n3921) );
  OR2X1 U4120 ( .IN1(n3923), .IN2(n3924), .Q(g6534) );
  AND2X1 U4121 ( .IN1(n3909), .IN2(g1466), .Q(n3924) );
  AND2X1 U4122 ( .IN1(n3910), .IN2(g1555), .Q(n3923) );
  OR2X1 U4123 ( .IN1(n3925), .IN2(n3926), .Q(g6533) );
  AND2X1 U4124 ( .IN1(n3909), .IN2(g1494), .Q(n3926) );
  AND2X1 U4125 ( .IN1(n3910), .IN2(g1534), .Q(n3925) );
  AND2X1 U4126 ( .IN1(n3147), .IN2(g8986), .Q(g6531) );
  OR2X1 U4127 ( .IN1(n3927), .IN2(n3928), .Q(g6529) );
  AND2X1 U4128 ( .IN1(n3909), .IN2(g1470), .Q(n3928) );
  AND2X1 U4129 ( .IN1(n3910), .IN2(g1552), .Q(n3927) );
  OR2X1 U4130 ( .IN1(n3929), .IN2(n3930), .Q(g6528) );
  AND2X1 U4131 ( .IN1(n3909), .IN2(g1499), .Q(n3930) );
  AND2X1 U4132 ( .IN1(n3910), .IN2(g1531), .Q(n3929) );
  AND2X1 U4133 ( .IN1(n3147), .IN2(g8985), .Q(g6526) );
  AND2X1 U4134 ( .IN1(n3931), .IN2(n1610), .Q(g6525) );
  XNOR2X1 U4135 ( .IN1(n2899), .IN2(n2853), .Q(n3931) );
  OR2X1 U4136 ( .IN1(n3932), .IN2(n3933), .Q(g6524) );
  AND2X1 U4137 ( .IN1(n3909), .IN2(g1428), .Q(n3933) );
  AND2X1 U4138 ( .IN1(n3910), .IN2(g1589), .Q(n3932) );
  OR2X1 U4139 ( .IN1(n3934), .IN2(n3935), .Q(g6523) );
  AND2X1 U4140 ( .IN1(n3909), .IN2(g1474), .Q(n3935) );
  AND2X1 U4141 ( .IN1(n3910), .IN2(g1549), .Q(n3934) );
  OR2X1 U4142 ( .IN1(n3936), .IN2(n3937), .Q(g6522) );
  AND2X1 U4143 ( .IN1(n3909), .IN2(g1504), .Q(n3937) );
  AND2X1 U4144 ( .IN1(n3910), .IN2(g1528), .Q(n3936) );
  AND2X1 U4145 ( .IN1(n3938), .IN2(n1610), .Q(g6516) );
  INVX0 U4146 ( .INP(n3939), .ZN(n3938) );
  OR2X1 U4147 ( .IN1(n3940), .IN2(n2899), .Q(n3939) );
  INVX0 U4148 ( .INP(n3941), .ZN(n2899) );
  OR2X1 U4149 ( .IN1(n1659), .IN2(n3942), .Q(n3941) );
  AND2X1 U4150 ( .IN1(n3942), .IN2(n1659), .Q(n3940) );
  OR2X1 U4151 ( .IN1(n3943), .IN2(n3944), .Q(g6515) );
  AND2X1 U4152 ( .IN1(n3909), .IN2(g1448), .Q(n3944) );
  AND2X1 U4153 ( .IN1(n3910), .IN2(g1607), .Q(n3943) );
  OR2X1 U4154 ( .IN1(n3945), .IN2(n3946), .Q(g6514) );
  AND2X1 U4155 ( .IN1(n3909), .IN2(g1407), .Q(n3946) );
  AND2X1 U4156 ( .IN1(n3910), .IN2(g1586), .Q(n3945) );
  OR2X1 U4157 ( .IN1(n3947), .IN2(n3948), .Q(g6513) );
  AND2X1 U4158 ( .IN1(n3909), .IN2(g1508), .Q(n3948) );
  AND2X1 U4159 ( .IN1(n3910), .IN2(g1524), .Q(n3947) );
  AND2X1 U4160 ( .IN1(n1610), .IN2(n3949), .Q(g6508) );
  OR2X1 U4161 ( .IN1(n3950), .IN2(n3951), .Q(n3949) );
  AND2X1 U4162 ( .IN1(n3942), .IN2(g1776), .Q(n3951) );
  OR2X1 U4163 ( .IN1(n369), .IN2(n3807), .Q(n3942) );
  AND2X1 U4164 ( .IN1(n3952), .IN2(n3782), .Q(n3950) );
  AND2X1 U4165 ( .IN1(test_so5), .IN2(n3807), .Q(n3952) );
  OR2X1 U4166 ( .IN1(n3953), .IN2(n3954), .Q(g6507) );
  AND2X1 U4167 ( .IN1(n3909), .IN2(g1444), .Q(n3954) );
  AND2X1 U4168 ( .IN1(n3910), .IN2(g1604), .Q(n3953) );
  OR2X1 U4169 ( .IN1(n3955), .IN2(n3956), .Q(g6506) );
  AND2X1 U4170 ( .IN1(n3909), .IN2(g1424), .Q(n3956) );
  AND2X1 U4171 ( .IN1(n3910), .IN2(g1583), .Q(n3955) );
  AND2X1 U4172 ( .IN1(n1610), .IN2(n3957), .Q(g6502) );
  XNOR2X1 U4173 ( .IN1(n2904), .IN2(n3782), .Q(n3957) );
  AND2X1 U4174 ( .IN1(g1766), .IN2(n2903), .Q(n3782) );
  OR2X1 U4175 ( .IN1(n3958), .IN2(n3959), .Q(g6501) );
  AND2X1 U4176 ( .IN1(n3909), .IN2(g1440), .Q(n3959) );
  AND2X1 U4177 ( .IN1(n3910), .IN2(g1601), .Q(n3958) );
  OR2X1 U4178 ( .IN1(n3960), .IN2(n3961), .Q(g6500) );
  AND2X1 U4179 ( .IN1(n3909), .IN2(g1411), .Q(n3961) );
  AND2X1 U4180 ( .IN1(n3910), .IN2(g1580), .Q(n3960) );
  OR2X1 U4181 ( .IN1(n3962), .IN2(n3963), .Q(g6481) );
  AND2X1 U4182 ( .IN1(n3909), .IN2(g1436), .Q(n3963) );
  AND2X1 U4183 ( .IN1(n3910), .IN2(g1598), .Q(n3962) );
  OR2X1 U4184 ( .IN1(n3964), .IN2(n3965), .Q(g6480) );
  AND2X1 U4185 ( .IN1(n3909), .IN2(g1419), .Q(n3965) );
  AND2X1 U4186 ( .IN1(n3910), .IN2(g1577), .Q(n3964) );
  OR2X1 U4187 ( .IN1(n3966), .IN2(n3967), .Q(g6479) );
  AND2X1 U4188 ( .IN1(n3909), .IN2(g1432), .Q(n3967) );
  AND2X1 U4189 ( .IN1(n3910), .IN2(g1595), .Q(n3966) );
  OR2X1 U4190 ( .IN1(n3968), .IN2(n3969), .Q(g6478) );
  AND2X1 U4191 ( .IN1(n3909), .IN2(g1515), .Q(n3969) );
  AND2X1 U4192 ( .IN1(n3910), .IN2(g1574), .Q(n3968) );
  AND2X1 U4193 ( .IN1(n3838), .IN2(n3970), .Q(g6471) );
  XNOR2X1 U4194 ( .IN1(n3033), .IN2(n2839), .Q(n3970) );
  OR2X1 U4195 ( .IN1(n3971), .IN2(n3972), .Q(g6470) );
  AND2X1 U4196 ( .IN1(n3909), .IN2(g1403), .Q(n3972) );
  AND2X1 U4197 ( .IN1(n3910), .IN2(g1592), .Q(n3971) );
  OR2X1 U4198 ( .IN1(n3973), .IN2(n3974), .Q(g6469) );
  AND2X1 U4199 ( .IN1(n3909), .IN2(g1520), .Q(n3974) );
  AND2X1 U4200 ( .IN1(n3910), .IN2(g1571), .Q(n3973) );
  OR2X1 U4201 ( .IN1(n3975), .IN2(n3976), .Q(g6468) );
  AND2X1 U4202 ( .IN1(n3909), .IN2(g1415), .Q(n3976) );
  AND2X1 U4203 ( .IN1(n3910), .IN2(g1567), .Q(n3975) );
  INVX0 U4204 ( .INP(n3909), .ZN(n3910) );
  OR2X1 U4205 ( .IN1(n1159), .IN2(n519), .Q(n3909) );
  AND2X1 U4206 ( .IN1(n3977), .IN2(g109), .Q(g6439) );
  XOR2X1 U4207 ( .IN1(n3978), .IN2(n3979), .Q(n3977) );
  XNOR2X1 U4208 ( .IN1(g153), .IN2(n2788), .Q(n3979) );
  XNOR2X1 U4209 ( .IN1(g148), .IN2(n2790), .Q(n3978) );
  AND2X1 U4210 ( .IN1(n3980), .IN2(n3652), .Q(g6392) );
  OR2X1 U4211 ( .IN1(n519), .IN2(n3653), .Q(n3980) );
  INVX0 U4212 ( .INP(g881), .ZN(n3653) );
  AND2X1 U4213 ( .IN1(g109), .IN2(g1389), .Q(g6334) );
  AND2X1 U4214 ( .IN1(g109), .IN2(n3020), .Q(g6332) );
  OR2X1 U4215 ( .IN1(n3981), .IN2(n3982), .Q(g6243) );
  XOR2X1 U4216 ( .IN1(n2866), .IN2(n1717), .Q(n3982) );
  AND2X1 U4217 ( .IN1(g109), .IN2(g1520), .Q(g6224) );
  AND2X1 U4218 ( .IN1(g109), .IN2(g1515), .Q(g6205) );
  AND2X1 U4219 ( .IN1(g109), .IN2(g1453), .Q(g6180) );
  AND2X1 U4220 ( .IN1(n30), .IN2(n3041), .Q(g6179) );
  AND2X1 U4221 ( .IN1(n3983), .IN2(g6331), .Q(n30) );
  OR2X1 U4222 ( .IN1(n3984), .IN2(n3985), .Q(g6155) );
  AND2X1 U4223 ( .IN1(n3986), .IN2(n1653), .Q(n3985) );
  AND2X1 U4224 ( .IN1(g1700), .IN2(g1707), .Q(n3986) );
  AND2X1 U4225 ( .IN1(g4076), .IN2(g1690), .Q(n3984) );
  AND2X1 U4226 ( .IN1(n3987), .IN2(n3623), .Q(g6126) );
  INVX0 U4227 ( .INP(n3981), .ZN(n3623) );
  XOR2X1 U4228 ( .IN1(n3159), .IN2(n2859), .Q(n3987) );
  AND2X1 U4229 ( .IN1(n3988), .IN2(n3627), .Q(g6123) );
  XNOR2X1 U4230 ( .IN1(n1193), .IN2(n2870), .Q(n3988) );
  OR2X1 U4231 ( .IN1(n3989), .IN2(n3990), .Q(g6099) );
  AND2X1 U4232 ( .IN1(n3991), .IN2(g1074), .Q(n3990) );
  AND2X1 U4233 ( .IN1(n3992), .IN2(g342), .Q(n3989) );
  OR2X1 U4234 ( .IN1(n3993), .IN2(n3994), .Q(g6096) );
  AND2X1 U4235 ( .IN1(n3991), .IN2(g1098), .Q(n3994) );
  AND2X1 U4236 ( .IN1(n3992), .IN2(g366), .Q(n3993) );
  OR2X1 U4237 ( .IN1(n3995), .IN2(n3996), .Q(g6093) );
  AND2X1 U4238 ( .IN1(n3991), .IN2(g1095), .Q(n3996) );
  AND2X1 U4239 ( .IN1(n3992), .IN2(g363), .Q(n3995) );
  OR2X1 U4240 ( .IN1(n3997), .IN2(n3998), .Q(g6088) );
  AND2X1 U4241 ( .IN1(n3991), .IN2(g1092), .Q(n3998) );
  AND2X1 U4242 ( .IN1(n3992), .IN2(g360), .Q(n3997) );
  OR2X1 U4243 ( .IN1(n3999), .IN2(n4000), .Q(g6080) );
  AND2X1 U4244 ( .IN1(n3991), .IN2(g1089), .Q(n4000) );
  AND2X1 U4245 ( .IN1(n3992), .IN2(g357), .Q(n3999) );
  OR2X1 U4246 ( .IN1(n4001), .IN2(n4002), .Q(g6071) );
  AND2X1 U4247 ( .IN1(n3991), .IN2(g1086), .Q(n4002) );
  AND2X1 U4248 ( .IN1(n3992), .IN2(g354), .Q(n4001) );
  OR2X1 U4249 ( .IN1(n4003), .IN2(n4004), .Q(g6068) );
  AND2X1 U4250 ( .IN1(n3991), .IN2(g1083), .Q(n4004) );
  AND2X1 U4251 ( .IN1(n3992), .IN2(g351), .Q(n4003) );
  OR2X1 U4252 ( .IN1(n4005), .IN2(n4006), .Q(g6059) );
  AND2X1 U4253 ( .IN1(n3991), .IN2(g1080), .Q(n4006) );
  AND2X1 U4254 ( .IN1(n3992), .IN2(g348), .Q(n4005) );
  OR2X1 U4255 ( .IN1(n4007), .IN2(n4008), .Q(g6054) );
  AND2X1 U4256 ( .IN1(test_so7), .IN2(n3991), .Q(n4008) );
  AND2X1 U4257 ( .IN1(n3992), .IN2(g336), .Q(n4007) );
  OR2X1 U4258 ( .IN1(n4009), .IN2(n4010), .Q(g6049) );
  AND2X1 U4259 ( .IN1(n3471), .IN2(g549), .Q(n4010) );
  OR2X1 U4260 ( .IN1(n4011), .IN2(n4012), .Q(g6045) );
  AND2X1 U4261 ( .IN1(n3471), .IN2(g575), .Q(n4012) );
  OR2X1 U4262 ( .IN1(n4013), .IN2(n4014), .Q(g6042) );
  AND2X1 U4263 ( .IN1(n3471), .IN2(g572), .Q(n4014) );
  OR2X1 U4264 ( .IN1(n4015), .IN2(n3518), .Q(g6038) );
  AND2X1 U4265 ( .IN1(n3471), .IN2(g569), .Q(n4015) );
  OR2X1 U4266 ( .IN1(n4016), .IN2(n3506), .Q(g6035) );
  AND2X1 U4267 ( .IN1(n3471), .IN2(g566), .Q(n4016) );
  OR2X1 U4268 ( .IN1(n4017), .IN2(n3478), .Q(g6026) );
  AND2X1 U4269 ( .IN1(n3471), .IN2(g563), .Q(n4017) );
  OR2X1 U4270 ( .IN1(n4018), .IN2(n3462), .Q(g6015) );
  AND2X1 U4271 ( .IN1(n3471), .IN2(g560), .Q(n4018) );
  OR2X1 U4272 ( .IN1(n4019), .IN2(n3524), .Q(g6002) );
  AND2X1 U4273 ( .IN1(n3471), .IN2(g557), .Q(n4019) );
  OR2X1 U4274 ( .IN1(n4020), .IN2(n3512), .Q(g6000) );
  AND2X1 U4275 ( .IN1(n3471), .IN2(g554), .Q(n4020) );
  OR2X1 U4276 ( .IN1(n4021), .IN2(n3494), .Q(g5996) );
  AND2X1 U4277 ( .IN1(n3471), .IN2(g546), .Q(n4021) );
  OR2X1 U4278 ( .IN1(n4022), .IN2(n1195), .Q(g5918) );
  AND2X1 U4279 ( .IN1(g109), .IN2(g119), .Q(n4022) );
  OR2X1 U4280 ( .IN1(n4023), .IN2(n4024), .Q(g5914) );
  AND2X1 U4281 ( .IN1(n3991), .IN2(g1077), .Q(n4024) );
  AND2X1 U4282 ( .IN1(n3992), .IN2(g345), .Q(n4023) );
  OR2X1 U4283 ( .IN1(n4025), .IN2(n4026), .Q(g5910) );
  AND2X1 U4284 ( .IN1(n3991), .IN2(g1071), .Q(n4026) );
  AND2X1 U4285 ( .IN1(n3992), .IN2(g339), .Q(n4025) );
  AND2X1 U4286 ( .IN1(n4027), .IN2(g109), .Q(g5770) );
  XOR2X1 U4287 ( .IN1(n4028), .IN2(n4029), .Q(n4027) );
  XNOR2X1 U4288 ( .IN1(g1508), .IN2(n1628), .Q(n4029) );
  XNOR2X1 U4289 ( .IN1(g1494), .IN2(n2792), .Q(n4028) );
  AND2X1 U4290 ( .IN1(n4030), .IN2(n4031), .Q(g5763) );
  OR2X1 U4291 ( .IN1(n5140), .IN2(n519), .Q(n4030) );
  OR2X1 U4292 ( .IN1(n4032), .IN2(n4033), .Q(g5755) );
  AND2X1 U4293 ( .IN1(n4034), .IN2(n1678), .Q(n4033) );
  AND2X1 U4294 ( .IN1(n4035), .IN2(n4036), .Q(n4034) );
  OR2X1 U4295 ( .IN1(n4037), .IN2(n4038), .Q(n4036) );
  AND2X1 U4296 ( .IN1(n1619), .IN2(g109), .Q(n4037) );
  OR2X1 U4297 ( .IN1(g6331), .IN2(n4039), .Q(n4035) );
  AND2X1 U4298 ( .IN1(g201), .IN2(g109), .Q(g6331) );
  AND2X1 U4299 ( .IN1(g6333), .IN2(n4040), .Q(n4032) );
  XNOR2X1 U4300 ( .IN1(n1619), .IN2(n4038), .Q(n4040) );
  INVX0 U4301 ( .INP(n4039), .ZN(n4038) );
  XOR2X1 U4302 ( .IN1(n4041), .IN2(g1389), .Q(n4039) );
  OR2X1 U4303 ( .IN1(n29), .IN2(g1386), .Q(n4041) );
  AND2X1 U4304 ( .IN1(n3983), .IN2(n1619), .Q(n29) );
  INVX0 U4305 ( .INP(n4042), .ZN(n3983) );
  OR2X1 U4306 ( .IN1(n4043), .IN2(n4044), .Q(n4042) );
  OR2X1 U4307 ( .IN1(n4045), .IN2(n4046), .Q(n4044) );
  OR2X1 U4308 ( .IN1(n4047), .IN2(n4048), .Q(n4046) );
  OR2X1 U4309 ( .IN1(g1383), .IN2(n3020), .Q(n4048) );
  OR2X1 U4310 ( .IN1(n3019), .IN2(n4049), .Q(n4047) );
  OR2X1 U4311 ( .IN1(g1371), .IN2(n3038), .Q(n4049) );
  INVX0 U4312 ( .INP(n4050), .ZN(n4045) );
  AND2X1 U4313 ( .IN1(n4051), .IN2(n4052), .Q(n4050) );
  AND2X1 U4314 ( .IN1(n5136), .IN2(n4053), .Q(n4052) );
  AND2X1 U4315 ( .IN1(n2880), .IN2(n5137), .Q(n4053) );
  AND2X1 U4316 ( .IN1(n2879), .IN2(n4054), .Q(n4051) );
  AND2X1 U4317 ( .IN1(n2877), .IN2(n2878), .Q(n4054) );
  OR2X1 U4318 ( .IN1(n4055), .IN2(n4056), .Q(n4043) );
  OR2X1 U4319 ( .IN1(n4057), .IN2(n4058), .Q(n4056) );
  OR2X1 U4320 ( .IN1(g186), .IN2(n4059), .Q(n4058) );
  OR2X1 U4321 ( .IN1(g213), .IN2(g237), .Q(n4059) );
  OR2X1 U4322 ( .IN1(g1386), .IN2(n4060), .Q(n4057) );
  OR2X1 U4323 ( .IN1(g192), .IN2(g243), .Q(n4060) );
  OR2X1 U4324 ( .IN1(n4061), .IN2(n4062), .Q(n4055) );
  OR2X1 U4325 ( .IN1(g1397), .IN2(n4063), .Q(n4062) );
  OR2X1 U4326 ( .IN1(g1400), .IN2(g197), .Q(n4063) );
  OR2X1 U4327 ( .IN1(g1389), .IN2(n4064), .Q(n4061) );
  OR2X1 U4328 ( .IN1(test_so3), .IN2(g248), .Q(n4064) );
  AND2X1 U4329 ( .IN1(g197), .IN2(g109), .Q(g6333) );
  AND2X1 U4330 ( .IN1(n4065), .IN2(g744), .Q(g5659) );
  AND2X1 U4331 ( .IN1(g743), .IN2(g109), .Q(n4065) );
  AND2X1 U4332 ( .IN1(n4066), .IN2(g742), .Q(g5658) );
  AND2X1 U4333 ( .IN1(g741), .IN2(g109), .Q(n4066) );
  AND2X1 U4334 ( .IN1(n4067), .IN2(n4068), .Q(g5556) );
  AND2X1 U4335 ( .IN1(n4069), .IN2(n4070), .Q(n4068) );
  AND2X1 U4336 ( .IN1(g1806), .IN2(g1707), .Q(n4070) );
  AND2X1 U4337 ( .IN1(g1690), .IN2(g1801), .Q(n4069) );
  INVX0 U4338 ( .INP(n4071), .ZN(n4067) );
  OR2X1 U4339 ( .IN1(n4072), .IN2(n4073), .Q(n4071) );
  OR2X1 U4340 ( .IN1(n3807), .IN2(n1626), .Q(n4073) );
  OR2X1 U4341 ( .IN1(n2904), .IN2(n4074), .Q(n3807) );
  OR2X1 U4342 ( .IN1(n2860), .IN2(n1715), .Q(n4074) );
  OR2X1 U4343 ( .IN1(g1781), .IN2(n3805), .Q(n4072) );
  AND2X1 U4344 ( .IN1(n4075), .IN2(n3159), .Q(g5543) );
  OR2X1 U4345 ( .IN1(n1622), .IN2(n3556), .Q(n3159) );
  OR2X1 U4346 ( .IN1(n1717), .IN2(n2866), .Q(n3556) );
  INVX0 U4347 ( .INP(n4076), .ZN(n4075) );
  AND2X1 U4348 ( .IN1(n4077), .IN2(n4078), .Q(n4076) );
  OR2X1 U4349 ( .IN1(g5849), .IN2(n1717), .Q(n4078) );
  OR2X1 U4350 ( .IN1(n2866), .IN2(n3981), .Q(g5849) );
  OR2X1 U4351 ( .IN1(n3981), .IN2(n1622), .Q(n4077) );
  OR2X1 U4352 ( .IN1(n519), .IN2(n4079), .Q(n3981) );
  OR2X1 U4353 ( .IN1(n2838), .IN2(n2649), .Q(n4079) );
  INVX0 U4354 ( .INP(n4080), .ZN(g5536) );
  OR2X1 U4355 ( .IN1(n4081), .IN2(n3691), .Q(n4080) );
  OR2X1 U4356 ( .IN1(n1193), .IN2(n1213), .Q(n4081) );
  OR2X1 U4357 ( .IN1(n4082), .IN2(n4083), .Q(g5529) );
  INVX0 U4358 ( .INP(n4084), .ZN(n4083) );
  OR2X1 U4359 ( .IN1(n4085), .IN2(g4174), .Q(n4084) );
  OR2X1 U4360 ( .IN1(n3691), .IN2(n2871), .Q(n4085) );
  AND2X1 U4361 ( .IN1(g4940), .IN2(g4174), .Q(n4082) );
  OR2X1 U4362 ( .IN1(n4086), .IN2(n1195), .Q(g5445) );
  AND2X1 U4363 ( .IN1(g109), .IN2(g12), .Q(n4086) );
  OR2X1 U4364 ( .IN1(n4087), .IN2(n1195), .Q(g5421) );
  AND2X1 U4365 ( .IN1(g109), .IN2(g9), .Q(n4087) );
  OR2X1 U4366 ( .IN1(n4088), .IN2(n4089), .Q(g5404) );
  AND2X1 U4367 ( .IN1(n371), .IN2(g1718), .Q(n4089) );
  AND2X1 U4368 ( .IN1(n3451), .IN2(g1713), .Q(n4088) );
  OR2X1 U4369 ( .IN1(n4090), .IN2(n4091), .Q(g5396) );
  AND2X1 U4370 ( .IN1(n371), .IN2(g1713), .Q(n4091) );
  AND2X1 U4371 ( .IN1(n3451), .IN2(g1710), .Q(n4090) );
  AND2X1 U4372 ( .IN1(n4092), .IN2(g1101), .Q(g5390) );
  AND2X1 U4373 ( .IN1(n4092), .IN2(g1110), .Q(g5173) );
  AND2X1 U4374 ( .IN1(n4092), .IN2(g1107), .Q(g5148) );
  AND2X1 U4375 ( .IN1(n4092), .IN2(g1104), .Q(g5126) );
  AND2X1 U4376 ( .IN1(g109), .IN2(n2907), .Q(n4092) );
  AND2X1 U4377 ( .IN1(n4093), .IN2(n4094), .Q(g5083) );
  AND2X1 U4378 ( .IN1(n371), .IN2(n3863), .Q(n4093) );
  INVX0 U4379 ( .INP(g4089), .ZN(n3863) );
  AND2X1 U4380 ( .IN1(n3627), .IN2(n2871), .Q(g4940) );
  INVX0 U4381 ( .INP(n3691), .ZN(n3627) );
  OR2X1 U4382 ( .IN1(test_so1), .IN2(n519), .Q(n3691) );
  AND2X1 U4383 ( .IN1(n4095), .IN2(n3018), .Q(g4905) );
  AND2X1 U4384 ( .IN1(n4095), .IN2(n3037), .Q(g4903) );
  AND2X1 U4385 ( .IN1(n4095), .IN2(n3030), .Q(g4902) );
  INVX0 U4386 ( .INP(n2902), .ZN(n4095) );
  AND2X1 U4387 ( .IN1(n4096), .IN2(n3053), .Q(g4893) );
  AND2X1 U4388 ( .IN1(n4096), .IN2(n3055), .Q(g4891) );
  AND2X1 U4389 ( .IN1(n4096), .IN2(n3035), .Q(g4890) );
  INVX0 U4390 ( .INP(n2900), .ZN(n4096) );
  OR2X1 U4391 ( .IN1(n4097), .IN2(n3213), .Q(n2900) );
  INVX0 U4392 ( .INP(n3446), .ZN(n3213) );
  OR2X1 U4393 ( .IN1(n3439), .IN2(n4098), .Q(n3446) );
  OR2X1 U4394 ( .IN1(g599), .IN2(g611), .Q(n4098) );
  OR2X1 U4395 ( .IN1(g605), .IN2(g591), .Q(n3439) );
  AND2X1 U4396 ( .IN1(n1607), .IN2(g611), .Q(n4097) );
  AND2X1 U4397 ( .IN1(g109), .IN2(n3016), .Q(g4506) );
  AND2X1 U4398 ( .IN1(n371), .IN2(n3046), .Q(g4500) );
  INVX0 U4399 ( .INP(n4099), .ZN(g4477) );
  OR2X1 U4400 ( .IN1(n519), .IN2(n1705), .Q(n4099) );
  INVX0 U4401 ( .INP(n4100), .ZN(g4473) );
  OR2X1 U4402 ( .IN1(n519), .IN2(n1708), .Q(n4100) );
  AND2X1 U4403 ( .IN1(g109), .IN2(g1121), .Q(g4471) );
  AND2X1 U4404 ( .IN1(test_so4), .IN2(g109), .Q(g4465) );
  AND2X1 U4405 ( .IN1(g109), .IN2(g1149), .Q(g4342) );
  AND2X1 U4406 ( .IN1(g109), .IN2(g1153), .Q(g4340) );
  OR2X1 U4407 ( .IN1(n4101), .IN2(n4102), .Q(g4309) );
  AND2X1 U4408 ( .IN1(n4103), .IN2(g1762), .Q(n4102) );
  AND2X1 U4409 ( .IN1(n4104), .IN2(g1806), .Q(n4101) );
  OR2X1 U4410 ( .IN1(n4105), .IN2(n4106), .Q(g4293) );
  AND2X1 U4411 ( .IN1(n4103), .IN2(g1759), .Q(n4106) );
  AND2X1 U4412 ( .IN1(n4104), .IN2(g1801), .Q(n4105) );
  OR2X1 U4413 ( .IN1(n4107), .IN2(n4108), .Q(g4283) );
  AND2X1 U4414 ( .IN1(n4103), .IN2(g1756), .Q(n4108) );
  AND2X1 U4415 ( .IN1(n4104), .IN2(g1796), .Q(n4107) );
  OR2X1 U4416 ( .IN1(n4109), .IN2(n4110), .Q(g4274) );
  AND2X1 U4417 ( .IN1(n4103), .IN2(g1753), .Q(n4110) );
  AND2X1 U4418 ( .IN1(n4104), .IN2(g1791), .Q(n4109) );
  OR2X1 U4419 ( .IN1(n4111), .IN2(n4112), .Q(g4264) );
  AND2X1 U4420 ( .IN1(n4103), .IN2(g1750), .Q(n4112) );
  AND2X1 U4421 ( .IN1(n4104), .IN2(g1786), .Q(n4111) );
  OR2X1 U4422 ( .IN1(n4113), .IN2(n4114), .Q(g4255) );
  AND2X1 U4423 ( .IN1(n4103), .IN2(g1747), .Q(n4114) );
  AND2X1 U4424 ( .IN1(n4104), .IN2(g1781), .Q(n4113) );
  OR2X1 U4425 ( .IN1(n4115), .IN2(n4116), .Q(g4239) );
  AND2X1 U4426 ( .IN1(n4103), .IN2(g1744), .Q(n4116) );
  AND2X1 U4427 ( .IN1(n4104), .IN2(g1776), .Q(n4115) );
  OR2X1 U4428 ( .IN1(n4117), .IN2(n4118), .Q(g4238) );
  AND2X1 U4429 ( .IN1(n4103), .IN2(g1741), .Q(n4118) );
  AND2X1 U4430 ( .IN1(n4104), .IN2(test_so5), .Q(n4117) );
  OR2X1 U4431 ( .IN1(n4119), .IN2(n4120), .Q(g4231) );
  AND2X1 U4432 ( .IN1(n4103), .IN2(g1738), .Q(n4120) );
  AND2X1 U4433 ( .IN1(n4104), .IN2(g1766), .Q(n4119) );
  OR2X1 U4434 ( .IN1(n521), .IN2(n3042), .Q(g4089) );
  INVX0 U4435 ( .INP(g1700), .ZN(n521) );
  AND2X1 U4436 ( .IN1(g1700), .IN2(n2848), .Q(g4076) );
  AND2X1 U4437 ( .IN1(n4121), .IN2(n4122), .Q(g3381) );
  AND2X1 U4438 ( .IN1(g936), .IN2(g940), .Q(n4122) );
  AND2X1 U4439 ( .IN1(g932), .IN2(g928), .Q(n4121) );
  INVX0 U4440 ( .INP(g23), .ZN(g3327) );
  AND2X1 U4441 ( .IN1(n2885), .IN2(n2849), .Q(g2478) );
  OR2X1 U4442 ( .IN1(n4123), .IN2(n4124), .Q(g11647) );
  AND2X1 U4443 ( .IN1(n3768), .IN2(n4125), .Q(n4124) );
  OR2X1 U4444 ( .IN1(n4126), .IN2(n4127), .Q(n4125) );
  AND2X1 U4445 ( .IN1(n4128), .IN2(n4129), .Q(n4127) );
  AND2X1 U4446 ( .IN1(n4130), .IN2(n4131), .Q(n4126) );
  INVX0 U4447 ( .INP(n4128), .ZN(n4131) );
  AND2X1 U4448 ( .IN1(n3147), .IN2(g336), .Q(n4123) );
  AND2X1 U4449 ( .IN1(n4132), .IN2(n4133), .Q(g11641) );
  INVX0 U4450 ( .INP(n4134), .ZN(n4132) );
  AND2X1 U4451 ( .IN1(n4135), .IN2(n4136), .Q(n4134) );
  OR2X1 U4452 ( .IN1(n1226), .IN2(n1721), .Q(n4136) );
  AND2X1 U4453 ( .IN1(n6), .IN2(n2901), .Q(n1226) );
  OR2X1 U4454 ( .IN1(n4137), .IN2(n2901), .Q(n4135) );
  AND2X1 U4455 ( .IN1(g1351), .IN2(n225), .Q(n2901) );
  INVX0 U4456 ( .INP(n4138), .ZN(n225) );
  AND2X1 U4457 ( .IN1(n4139), .IN2(n4133), .Q(g11640) );
  OR2X1 U4458 ( .IN1(n4140), .IN2(n4141), .Q(n4139) );
  AND2X1 U4459 ( .IN1(n1232), .IN2(n1231), .Q(n4141) );
  AND2X1 U4460 ( .IN1(n4137), .IN2(g1346), .Q(n4140) );
  OR2X1 U4461 ( .IN1(n1227), .IN2(n4138), .Q(n4137) );
  OR2X1 U4462 ( .IN1(n2819), .IN2(n4142), .Q(n4138) );
  OR2X1 U4463 ( .IN1(n2821), .IN2(n2820), .Q(n4142) );
  AND2X1 U4464 ( .IN1(n4143), .IN2(n4133), .Q(g11639) );
  XOR2X1 U4465 ( .IN1(n1231), .IN2(g1341), .Q(n4143) );
  AND2X1 U4466 ( .IN1(n4144), .IN2(n4133), .Q(g11636) );
  OR2X1 U4467 ( .IN1(n4145), .IN2(n3698), .Q(n4133) );
  AND2X1 U4468 ( .IN1(g109), .IN2(n2882), .Q(n3698) );
  AND2X1 U4469 ( .IN1(n4146), .IN2(g109), .Q(n4145) );
  OR2X1 U4470 ( .IN1(n4147), .IN2(n3036), .Q(n4146) );
  XNOR2X1 U4471 ( .IN1(n6), .IN2(n2821), .Q(n4144) );
  INVX0 U4472 ( .INP(n1227), .ZN(n6) );
  OR2X1 U4473 ( .IN1(n4148), .IN2(n4149), .Q(g11625) );
  AND2X1 U4474 ( .IN1(n3768), .IN2(n4150), .Q(n4149) );
  XOR2X1 U4475 ( .IN1(n4130), .IN2(n4129), .Q(n4150) );
  AND2X1 U4476 ( .IN1(n4151), .IN2(n4152), .Q(n4129) );
  OR2X1 U4477 ( .IN1(n4153), .IN2(n25), .Q(n4152) );
  XOR2X1 U4478 ( .IN1(n4154), .IN2(n4155), .Q(n4153) );
  OR2X1 U4479 ( .IN1(g461), .IN2(n4156), .Q(n4155) );
  OR2X1 U4480 ( .IN1(n1239), .IN2(n1681), .Q(n4151) );
  XOR2X1 U4481 ( .IN1(n4157), .IN2(n4158), .Q(n4130) );
  XOR2X1 U4482 ( .IN1(n4159), .IN2(n4160), .Q(n4158) );
  XOR2X1 U4483 ( .IN1(n4161), .IN2(n4162), .Q(n4160) );
  XOR2X1 U4484 ( .IN1(n4163), .IN2(n4164), .Q(n4162) );
  XOR2X1 U4485 ( .IN1(n4165), .IN2(n4166), .Q(n4161) );
  XOR2X1 U4486 ( .IN1(n4167), .IN2(n4168), .Q(n4159) );
  XOR2X1 U4487 ( .IN1(n4169), .IN2(n4170), .Q(n4168) );
  XOR2X1 U4488 ( .IN1(n4171), .IN2(n4172), .Q(n4167) );
  AND2X1 U4489 ( .IN1(n3147), .IN2(g345), .Q(n4148) );
  OR2X1 U4490 ( .IN1(n4173), .IN2(n4174), .Q(g11610) );
  AND2X1 U4491 ( .IN1(n4175), .IN2(g1333), .Q(n4174) );
  AND2X1 U4492 ( .IN1(n4176), .IN2(g1806), .Q(n4173) );
  OR2X1 U4493 ( .IN1(n4177), .IN2(n4178), .Q(g11609) );
  AND2X1 U4494 ( .IN1(n4175), .IN2(g1330), .Q(n4178) );
  AND2X1 U4495 ( .IN1(n4176), .IN2(g1801), .Q(n4177) );
  OR2X1 U4496 ( .IN1(n4179), .IN2(n4180), .Q(g11608) );
  AND2X1 U4497 ( .IN1(n4175), .IN2(g1327), .Q(n4180) );
  AND2X1 U4498 ( .IN1(n4176), .IN2(g1796), .Q(n4179) );
  OR2X1 U4499 ( .IN1(n4181), .IN2(n4182), .Q(g11607) );
  AND2X1 U4500 ( .IN1(n4175), .IN2(g1324), .Q(n4182) );
  AND2X1 U4501 ( .IN1(n4176), .IN2(g1791), .Q(n4181) );
  OR2X1 U4502 ( .IN1(n4183), .IN2(n4184), .Q(g11606) );
  AND2X1 U4503 ( .IN1(n4175), .IN2(g1321), .Q(n4184) );
  AND2X1 U4504 ( .IN1(n4176), .IN2(g1786), .Q(n4183) );
  OR2X1 U4505 ( .IN1(n4185), .IN2(n4186), .Q(g11605) );
  AND2X1 U4506 ( .IN1(n4175), .IN2(g1318), .Q(n4186) );
  AND2X1 U4507 ( .IN1(n4176), .IN2(g1781), .Q(n4185) );
  OR2X1 U4508 ( .IN1(n4187), .IN2(n4188), .Q(g11604) );
  AND2X1 U4509 ( .IN1(n4175), .IN2(g1314), .Q(n4188) );
  AND2X1 U4510 ( .IN1(n4176), .IN2(g1776), .Q(n4187) );
  OR2X1 U4511 ( .IN1(n4189), .IN2(n4190), .Q(g11603) );
  AND2X1 U4512 ( .IN1(n4176), .IN2(test_so5), .Q(n4190) );
  AND2X1 U4513 ( .IN1(test_so9), .IN2(n4175), .Q(n4189) );
  OR2X1 U4514 ( .IN1(n4191), .IN2(n4192), .Q(g11602) );
  AND2X1 U4515 ( .IN1(n4175), .IN2(g1308), .Q(n4192) );
  AND2X1 U4516 ( .IN1(n4176), .IN2(g1766), .Q(n4191) );
  INVX0 U4517 ( .INP(n4175), .ZN(n4176) );
  OR2X1 U4518 ( .IN1(n2889), .IN2(n1227), .Q(n4175) );
  OR2X1 U4519 ( .IN1(n3702), .IN2(n4193), .Q(n1227) );
  OR2X1 U4520 ( .IN1(n4194), .IN2(n4195), .Q(n4193) );
  AND2X1 U4521 ( .IN1(n4196), .IN2(n4197), .Q(n4194) );
  AND2X1 U4522 ( .IN1(n4198), .IN2(n4199), .Q(n4197) );
  AND2X1 U4523 ( .IN1(n4200), .IN2(n4201), .Q(n4199) );
  XNOR2X1 U4524 ( .IN1(test_so2), .IN2(g1255), .Q(n4201) );
  AND2X1 U4525 ( .IN1(n4202), .IN2(n4203), .Q(n4200) );
  XNOR2X1 U4526 ( .IN1(n2905), .IN2(n2721), .Q(n4203) );
  XNOR2X1 U4527 ( .IN1(n4204), .IN2(n4205), .Q(n4202) );
  AND2X1 U4528 ( .IN1(n4206), .IN2(n4207), .Q(n4198) );
  XNOR2X1 U4529 ( .IN1(test_so8), .IN2(g1245), .Q(n4207) );
  XNOR2X1 U4530 ( .IN1(n2776), .IN2(n2777), .Q(n4206) );
  AND2X1 U4531 ( .IN1(n4208), .IN2(n4209), .Q(n4196) );
  AND2X1 U4532 ( .IN1(n4210), .IN2(n4211), .Q(n4209) );
  XNOR2X1 U4533 ( .IN1(n2742), .IN2(n2750), .Q(n4211) );
  AND2X1 U4534 ( .IN1(n4212), .IN2(n4213), .Q(n4210) );
  XNOR2X1 U4535 ( .IN1(n1871), .IN2(n2775), .Q(n4213) );
  XNOR2X1 U4536 ( .IN1(n2812), .IN2(n2811), .Q(n4212) );
  AND2X1 U4537 ( .IN1(n4214), .IN2(n4215), .Q(n4208) );
  XNOR2X1 U4538 ( .IN1(n2814), .IN2(n2813), .Q(n4215) );
  XNOR2X1 U4539 ( .IN1(n2741), .IN2(n2752), .Q(n4214) );
  OR2X1 U4540 ( .IN1(n4216), .IN2(n4217), .Q(g11579) );
  AND2X1 U4541 ( .IN1(n4218), .IN2(n3451), .Q(n4217) );
  XNOR2X1 U4542 ( .IN1(n2885), .IN2(n4219), .Q(n4218) );
  OR2X1 U4543 ( .IN1(n4220), .IN2(n4221), .Q(n4219) );
  AND2X1 U4544 ( .IN1(n1260), .IN2(n4222), .Q(n4221) );
  AND2X1 U4545 ( .IN1(n4223), .IN2(n4224), .Q(n4220) );
  OR2X1 U4546 ( .IN1(n1258), .IN2(n4225), .Q(n4224) );
  INVX0 U4547 ( .INP(n1262), .ZN(n4225) );
  OR2X1 U4548 ( .IN1(n4226), .IN2(n4227), .Q(n1262) );
  AND2X1 U4549 ( .IN1(n4227), .IN2(n4226), .Q(n1258) );
  INVX0 U4550 ( .INP(n4228), .ZN(n4226) );
  OR2X1 U4551 ( .IN1(n4229), .IN2(n4230), .Q(n4228) );
  AND2X1 U4552 ( .IN1(n1685), .IN2(n4231), .Q(n4230) );
  OR2X1 U4553 ( .IN1(n4232), .IN2(g1153), .Q(n4231) );
  AND2X1 U4554 ( .IN1(n4233), .IN2(n4234), .Q(n4232) );
  AND2X1 U4555 ( .IN1(n4235), .IN2(n4236), .Q(n4234) );
  AND2X1 U4556 ( .IN1(n4237), .IN2(n4238), .Q(n4236) );
  AND2X1 U4557 ( .IN1(n1597), .IN2(n2906), .Q(n4238) );
  AND2X1 U4558 ( .IN1(n1618), .IN2(n1617), .Q(n4237) );
  AND2X1 U4559 ( .IN1(n4239), .IN2(n1706), .Q(n4235) );
  AND2X1 U4560 ( .IN1(n1705), .IN2(n1660), .Q(n4239) );
  AND2X1 U4561 ( .IN1(n4240), .IN2(n4241), .Q(n4233) );
  AND2X1 U4562 ( .IN1(n4242), .IN2(n2785), .Q(n4241) );
  AND2X1 U4563 ( .IN1(n2784), .IN2(n1708), .Q(n4242) );
  AND2X1 U4564 ( .IN1(n4243), .IN2(n5138), .Q(n4240) );
  AND2X1 U4565 ( .IN1(n2787), .IN2(n2786), .Q(n4243) );
  AND2X1 U4566 ( .IN1(n1686), .IN2(g1149), .Q(n4229) );
  OR2X1 U4567 ( .IN1(n3521), .IN2(g1110), .Q(n4227) );
  OR2X1 U4568 ( .IN1(n3503), .IN2(g1104), .Q(n3521) );
  INVX0 U4569 ( .INP(n3499), .ZN(n3503) );
  AND2X1 U4570 ( .IN1(g1101), .IN2(n1614), .Q(n3499) );
  AND2X1 U4571 ( .IN1(n371), .IN2(g1618), .Q(n4216) );
  OR2X1 U4572 ( .IN1(n4244), .IN2(n4245), .Q(g11514) );
  AND2X1 U4573 ( .IN1(g6193), .IN2(n4246), .Q(n4245) );
  INVX0 U4574 ( .INP(n4247), .ZN(n4246) );
  AND2X1 U4575 ( .IN1(g1419), .IN2(g109), .Q(g6193) );
  AND2X1 U4576 ( .IN1(n4248), .IN2(n4247), .Q(n4244) );
  XNOR2X1 U4577 ( .IN1(n4249), .IN2(n4250), .Q(n4247) );
  XNOR2X1 U4578 ( .IN1(g1448), .IN2(n2657), .Q(n4250) );
  XNOR2X1 U4579 ( .IN1(n4222), .IN2(n1627), .Q(n4249) );
  INVX0 U4580 ( .INP(n4223), .ZN(n4222) );
  OR2X1 U4581 ( .IN1(n4251), .IN2(n4252), .Q(n4223) );
  AND2X1 U4582 ( .IN1(n4253), .IN2(n3471), .Q(n4252) );
  OR2X1 U4583 ( .IN1(n4254), .IN2(n4255), .Q(n4253) );
  AND2X1 U4584 ( .IN1(n4256), .IN2(n4257), .Q(n4255) );
  OR2X1 U4585 ( .IN1(g10726), .IN2(n4258), .Q(n4256) );
  AND2X1 U4586 ( .IN1(n4259), .IN2(n1699), .Q(n4254) );
  INVX0 U4587 ( .INP(n4257), .ZN(n4259) );
  OR2X1 U4588 ( .IN1(n4260), .IN2(n4261), .Q(n4257) );
  OR2X1 U4589 ( .IN1(n3029), .IN2(n3023), .Q(n4261) );
  OR2X1 U4590 ( .IN1(n3017), .IN2(n3065), .Q(n4260) );
  AND2X1 U4591 ( .IN1(g18), .IN2(g201), .Q(n4251) );
  AND2X1 U4592 ( .IN1(n1602), .IN2(g109), .Q(n4248) );
  OR2X1 U4593 ( .IN1(n4262), .IN2(n4263), .Q(g11488) );
  AND2X1 U4594 ( .IN1(n3768), .IN2(n4164), .Q(n4263) );
  OR2X1 U4595 ( .IN1(n4264), .IN2(n4265), .Q(n4164) );
  AND2X1 U4596 ( .IN1(n4266), .IN2(n1239), .Q(n4265) );
  XNOR2X1 U4597 ( .IN1(n4267), .IN2(g516), .Q(n4266) );
  OR2X1 U4598 ( .IN1(n1641), .IN2(n4268), .Q(n4267) );
  AND2X1 U4599 ( .IN1(n25), .IN2(g309), .Q(n4264) );
  AND2X1 U4600 ( .IN1(n3147), .IN2(g342), .Q(n4262) );
  OR2X1 U4601 ( .IN1(n4269), .IN2(n4270), .Q(g11487) );
  AND2X1 U4602 ( .IN1(n3768), .IN2(n4163), .Q(n4270) );
  OR2X1 U4603 ( .IN1(n4271), .IN2(n4272), .Q(n4163) );
  AND2X1 U4604 ( .IN1(n4273), .IN2(n1239), .Q(n4272) );
  XNOR2X1 U4605 ( .IN1(n4274), .IN2(g511), .Q(n4273) );
  OR2X1 U4606 ( .IN1(g456), .IN2(n4268), .Q(n4274) );
  OR2X1 U4607 ( .IN1(g461), .IN2(n4275), .Q(n4268) );
  OR2X1 U4608 ( .IN1(n1606), .IN2(g466), .Q(n4275) );
  AND2X1 U4609 ( .IN1(n25), .IN2(g333), .Q(n4271) );
  AND2X1 U4610 ( .IN1(n3147), .IN2(g366), .Q(n4269) );
  OR2X1 U4611 ( .IN1(n4276), .IN2(n4277), .Q(g11486) );
  AND2X1 U4612 ( .IN1(n3768), .IN2(n4166), .Q(n4277) );
  OR2X1 U4613 ( .IN1(n4278), .IN2(n4279), .Q(n4166) );
  AND2X1 U4614 ( .IN1(n4280), .IN2(n1239), .Q(n4279) );
  XNOR2X1 U4615 ( .IN1(n4281), .IN2(g506), .Q(n4280) );
  OR2X1 U4616 ( .IN1(g471), .IN2(n4282), .Q(n4281) );
  AND2X1 U4617 ( .IN1(n25), .IN2(g330), .Q(n4278) );
  AND2X1 U4618 ( .IN1(n3147), .IN2(g363), .Q(n4276) );
  OR2X1 U4619 ( .IN1(n4283), .IN2(n4284), .Q(g11485) );
  AND2X1 U4620 ( .IN1(n3768), .IN2(n4172), .Q(n4284) );
  OR2X1 U4621 ( .IN1(n4285), .IN2(n4286), .Q(n4172) );
  AND2X1 U4622 ( .IN1(n4287), .IN2(n1239), .Q(n4286) );
  XNOR2X1 U4623 ( .IN1(n1690), .IN2(n4288), .Q(n4287) );
  AND2X1 U4624 ( .IN1(n4289), .IN2(g461), .Q(n4288) );
  AND2X1 U4625 ( .IN1(n25), .IN2(g327), .Q(n4285) );
  AND2X1 U4626 ( .IN1(n3147), .IN2(g360), .Q(n4283) );
  OR2X1 U4627 ( .IN1(n4290), .IN2(n4291), .Q(g11484) );
  AND2X1 U4628 ( .IN1(n3768), .IN2(n4171), .Q(n4291) );
  OR2X1 U4629 ( .IN1(n4292), .IN2(n4293), .Q(n4171) );
  AND2X1 U4630 ( .IN1(n4294), .IN2(n1239), .Q(n4293) );
  XNOR2X1 U4631 ( .IN1(n4295), .IN2(g496), .Q(n4294) );
  OR2X1 U4632 ( .IN1(n4296), .IN2(n4297), .Q(n4295) );
  OR2X1 U4633 ( .IN1(g471), .IN2(g461), .Q(n4297) );
  AND2X1 U4634 ( .IN1(n25), .IN2(g324), .Q(n4292) );
  AND2X1 U4635 ( .IN1(n3147), .IN2(g357), .Q(n4290) );
  OR2X1 U4636 ( .IN1(n4298), .IN2(n4299), .Q(g11483) );
  AND2X1 U4637 ( .IN1(n3768), .IN2(n4170), .Q(n4299) );
  OR2X1 U4638 ( .IN1(n4300), .IN2(n4301), .Q(n4170) );
  AND2X1 U4639 ( .IN1(n4302), .IN2(n1239), .Q(n4301) );
  XNOR2X1 U4640 ( .IN1(n1691), .IN2(n4303), .Q(n4302) );
  AND2X1 U4641 ( .IN1(n4289), .IN2(n1594), .Q(n4303) );
  AND2X1 U4642 ( .IN1(n1641), .IN2(n4304), .Q(n4289) );
  AND2X1 U4643 ( .IN1(g466), .IN2(n1606), .Q(n4304) );
  AND2X1 U4644 ( .IN1(n25), .IN2(g321), .Q(n4300) );
  AND2X1 U4645 ( .IN1(n3147), .IN2(g354), .Q(n4298) );
  OR2X1 U4646 ( .IN1(n4305), .IN2(n4306), .Q(g11482) );
  AND2X1 U4647 ( .IN1(n3768), .IN2(n4157), .Q(n4306) );
  OR2X1 U4648 ( .IN1(n4307), .IN2(n4308), .Q(n4157) );
  AND2X1 U4649 ( .IN1(n4309), .IN2(n1239), .Q(n4308) );
  XNOR2X1 U4650 ( .IN1(n4310), .IN2(g486), .Q(n4309) );
  OR2X1 U4651 ( .IN1(n1594), .IN2(n4156), .Q(n4310) );
  OR2X1 U4652 ( .IN1(g466), .IN2(n4311), .Q(n4156) );
  OR2X1 U4653 ( .IN1(n1641), .IN2(g471), .Q(n4311) );
  AND2X1 U4654 ( .IN1(n25), .IN2(g318), .Q(n4307) );
  AND2X1 U4655 ( .IN1(n3147), .IN2(g351), .Q(n4305) );
  OR2X1 U4656 ( .IN1(n4312), .IN2(n4313), .Q(g11481) );
  AND2X1 U4657 ( .IN1(n3768), .IN2(n4169), .Q(n4313) );
  OR2X1 U4658 ( .IN1(n4314), .IN2(n4315), .Q(n4169) );
  AND2X1 U4659 ( .IN1(n4316), .IN2(n1239), .Q(n4315) );
  XNOR2X1 U4660 ( .IN1(n4317), .IN2(g481), .Q(n4316) );
  OR2X1 U4661 ( .IN1(g471), .IN2(n4318), .Q(n4317) );
  AND2X1 U4662 ( .IN1(n25), .IN2(g315), .Q(n4314) );
  AND2X1 U4663 ( .IN1(n3147), .IN2(g348), .Q(n4312) );
  OR2X1 U4664 ( .IN1(n4319), .IN2(n4320), .Q(g11478) );
  AND2X1 U4665 ( .IN1(n3768), .IN2(n4165), .Q(n4320) );
  OR2X1 U4666 ( .IN1(n4321), .IN2(n4322), .Q(n4165) );
  AND2X1 U4667 ( .IN1(n4323), .IN2(n1239), .Q(n4322) );
  XNOR2X1 U4668 ( .IN1(n4324), .IN2(g476), .Q(n4323) );
  OR2X1 U4669 ( .IN1(n1606), .IN2(n4318), .Q(n4324) );
  OR2X1 U4670 ( .IN1(g456), .IN2(n4325), .Q(n4318) );
  OR2X1 U4671 ( .IN1(n1594), .IN2(g466), .Q(n4325) );
  AND2X1 U4672 ( .IN1(n25), .IN2(g312), .Q(n4321) );
  AND2X1 U4673 ( .IN1(n3147), .IN2(g339), .Q(n4319) );
  INVX0 U4674 ( .INP(n3768), .ZN(n3147) );
  AND2X1 U4675 ( .IN1(g750), .IN2(n1647), .Q(n3768) );
  OR2X1 U4676 ( .IN1(n4326), .IN2(n4327), .Q(g11443) );
  AND2X1 U4677 ( .IN1(n3736), .IN2(g1275), .Q(n4327) );
  AND2X1 U4678 ( .IN1(g109), .IN2(n3702), .Q(n3736) );
  AND2X1 U4679 ( .IN1(n3735), .IN2(n4204), .Q(n4326) );
  OR2X1 U4680 ( .IN1(n4328), .IN2(n4329), .Q(n4204) );
  AND2X1 U4681 ( .IN1(n4330), .IN2(n3721), .Q(n4329) );
  INVX0 U4682 ( .INP(n4195), .ZN(n3721) );
  OR2X1 U4683 ( .IN1(n4331), .IN2(n4332), .Q(n4330) );
  AND2X1 U4684 ( .IN1(n1862), .IN2(n4333), .Q(n4332) );
  OR2X1 U4685 ( .IN1(n4334), .IN2(g1284), .Q(n4333) );
  AND2X1 U4686 ( .IN1(n4335), .IN2(n4336), .Q(n4334) );
  AND2X1 U4687 ( .IN1(n4337), .IN2(n4338), .Q(n4336) );
  AND2X1 U4688 ( .IN1(n4339), .IN2(n4340), .Q(n4338) );
  AND2X1 U4689 ( .IN1(n2749), .IN2(n2905), .Q(n4340) );
  AND2X1 U4690 ( .IN1(n2752), .IN2(n2750), .Q(n4339) );
  AND2X1 U4691 ( .IN1(n4341), .IN2(n2755), .Q(n4337) );
  AND2X1 U4692 ( .IN1(n2754), .IN2(n2753), .Q(n4341) );
  AND2X1 U4693 ( .IN1(n4342), .IN2(n4343), .Q(n4335) );
  AND2X1 U4694 ( .IN1(n4344), .IN2(n2775), .Q(n4343) );
  AND2X1 U4695 ( .IN1(n2774), .IN2(n2756), .Q(n4344) );
  AND2X1 U4696 ( .IN1(n4345), .IN2(n2813), .Q(n4342) );
  AND2X1 U4697 ( .IN1(n2811), .IN2(n2777), .Q(n4345) );
  AND2X1 U4698 ( .IN1(n1864), .IN2(g1280), .Q(n4331) );
  AND2X1 U4699 ( .IN1(n4205), .IN2(n4195), .Q(n4328) );
  OR2X1 U4700 ( .IN1(n2881), .IN2(n3719), .Q(n4195) );
  OR2X1 U4701 ( .IN1(n2650), .IN2(n4346), .Q(n3719) );
  OR2X1 U4702 ( .IN1(n2887), .IN2(n2651), .Q(n4346) );
  XNOR2X1 U4703 ( .IN1(n4347), .IN2(g1027), .Q(n4205) );
  OR2X1 U4704 ( .IN1(n4128), .IN2(n2888), .Q(n4347) );
  INVX0 U4705 ( .INP(n3702), .ZN(n3735) );
  OR2X1 U4706 ( .IN1(g1713), .IN2(n4348), .Q(n3702) );
  OR2X1 U4707 ( .IN1(n2844), .IN2(n371), .Q(n4348) );
  AND2X1 U4708 ( .IN1(n4349), .IN2(n4350), .Q(g11393) );
  XNOR2X1 U4709 ( .IN1(n4351), .IN2(g986), .Q(n4349) );
  AND2X1 U4710 ( .IN1(n4352), .IN2(n4350), .Q(g11392) );
  OR2X1 U4711 ( .IN1(n4353), .IN2(n4354), .Q(n4352) );
  AND2X1 U4712 ( .IN1(n4351), .IN2(g981), .Q(n4354) );
  OR2X1 U4713 ( .IN1(n3149), .IN2(n4355), .Q(n4351) );
  AND2X1 U4714 ( .IN1(n4356), .IN2(n4357), .Q(n4353) );
  AND2X1 U4715 ( .IN1(n3149), .IN2(g976), .Q(n4356) );
  OR2X1 U4716 ( .IN1(n1720), .IN2(n4358), .Q(n3149) );
  OR2X1 U4717 ( .IN1(n2892), .IN2(n2891), .Q(n4358) );
  AND2X1 U4718 ( .IN1(n4359), .IN2(n4350), .Q(g11391) );
  XNOR2X1 U4719 ( .IN1(n4357), .IN2(n2892), .Q(n4359) );
  AND2X1 U4720 ( .IN1(n4360), .IN2(n4361), .Q(g11380) );
  OR2X1 U4721 ( .IN1(n4362), .IN2(g471), .Q(n4361) );
  AND2X1 U4722 ( .IN1(n4363), .IN2(n4364), .Q(n4362) );
  AND2X1 U4723 ( .IN1(n4360), .IN2(n4365), .Q(g11376) );
  OR2X1 U4724 ( .IN1(n4366), .IN2(n4367), .Q(n4365) );
  AND2X1 U4725 ( .IN1(n4368), .IN2(g466), .Q(n4367) );
  OR2X1 U4726 ( .IN1(n4282), .IN2(n4369), .Q(n4368) );
  AND2X1 U4727 ( .IN1(n4370), .IN2(n4371), .Q(n4366) );
  AND2X1 U4728 ( .IN1(g461), .IN2(g456), .Q(n4371) );
  AND2X1 U4729 ( .IN1(n4363), .IN2(n4282), .Q(n4370) );
  AND2X1 U4730 ( .IN1(n4372), .IN2(n4360), .Q(g11372) );
  XNOR2X1 U4731 ( .IN1(n4373), .IN2(g461), .Q(n4372) );
  OR2X1 U4732 ( .IN1(n1641), .IN2(n4369), .Q(n4373) );
  AND2X1 U4733 ( .IN1(n4374), .IN2(n4375), .Q(g11349) );
  OR2X1 U4734 ( .IN1(n13), .IN2(g971), .Q(n4375) );
  AND2X1 U4735 ( .IN1(n4376), .IN2(n4350), .Q(n4374) );
  OR2X1 U4736 ( .IN1(n4377), .IN2(n2897), .Q(n4350) );
  AND2X1 U4737 ( .IN1(g109), .IN2(n4378), .Q(n2897) );
  OR2X1 U4738 ( .IN1(n3064), .IN2(n4379), .Q(n4378) );
  AND2X1 U4739 ( .IN1(g3007), .IN2(n5139), .Q(n4379) );
  INVX0 U4740 ( .INP(n4357), .ZN(n4376) );
  AND2X1 U4741 ( .IN1(g971), .IN2(n13), .Q(n4357) );
  INVX0 U4742 ( .INP(n4355), .ZN(n13) );
  OR2X1 U4743 ( .IN1(n4380), .IN2(n4381), .Q(n4355) );
  OR2X1 U4744 ( .IN1(n25), .IN2(n4382), .Q(n4381) );
  AND2X1 U4745 ( .IN1(n4383), .IN2(n4384), .Q(n4382) );
  AND2X1 U4746 ( .IN1(n4385), .IN2(n4386), .Q(n4384) );
  AND2X1 U4747 ( .IN1(n4387), .IN2(n4388), .Q(n4386) );
  XNOR2X1 U4748 ( .IN1(n2797), .IN2(n2798), .Q(n4388) );
  AND2X1 U4749 ( .IN1(n4389), .IN2(n4390), .Q(n4387) );
  XNOR2X1 U4750 ( .IN1(n2799), .IN2(n2800), .Q(n4390) );
  XNOR2X1 U4751 ( .IN1(n2782), .IN2(n2783), .Q(n4389) );
  AND2X1 U4752 ( .IN1(n4391), .IN2(n4392), .Q(n4385) );
  XNOR2X1 U4753 ( .IN1(n2606), .IN2(n2757), .Q(n4392) );
  XOR2X1 U4754 ( .IN1(n1681), .IN2(n4393), .Q(n4391) );
  AND2X1 U4755 ( .IN1(n4394), .IN2(n4395), .Q(n4383) );
  AND2X1 U4756 ( .IN1(n4396), .IN2(n4397), .Q(n4395) );
  XNOR2X1 U4757 ( .IN1(n2778), .IN2(n2779), .Q(n4397) );
  AND2X1 U4758 ( .IN1(n4398), .IN2(n4399), .Q(n4396) );
  XNOR2X1 U4759 ( .IN1(n2816), .IN2(n2815), .Q(n4399) );
  XNOR2X1 U4760 ( .IN1(n2605), .IN2(n2751), .Q(n4398) );
  AND2X1 U4761 ( .IN1(n4400), .IN2(n4401), .Q(n4394) );
  XNOR2X1 U4762 ( .IN1(n2818), .IN2(n2817), .Q(n4401) );
  XNOR2X1 U4763 ( .IN1(n2780), .IN2(n2781), .Q(n4400) );
  AND2X1 U4764 ( .IN1(n4402), .IN2(n4360), .Q(g11340) );
  AND2X1 U4765 ( .IN1(g109), .IN2(n2908), .Q(n4360) );
  XNOR2X1 U4766 ( .IN1(n4363), .IN2(n1641), .Q(n4402) );
  INVX0 U4767 ( .INP(n4369), .ZN(n4363) );
  OR2X1 U4768 ( .IN1(n25), .IN2(n4403), .Q(n4369) );
  AND2X1 U4769 ( .IN1(n4364), .IN2(g471), .Q(n4403) );
  INVX0 U4770 ( .INP(n4282), .ZN(n4364) );
  OR2X1 U4771 ( .IN1(n1594), .IN2(n4296), .Q(n4282) );
  OR2X1 U4772 ( .IN1(n1646), .IN2(n1641), .Q(n4296) );
  OR2X1 U4773 ( .IN1(n4404), .IN2(n4405), .Q(g11338) );
  AND2X1 U4774 ( .IN1(n1239), .IN2(g516), .Q(n4405) );
  AND2X1 U4775 ( .IN1(n25), .IN2(g476), .Q(n4404) );
  OR2X1 U4776 ( .IN1(n4406), .IN2(n4407), .Q(g11337) );
  AND2X1 U4777 ( .IN1(n1239), .IN2(g511), .Q(n4407) );
  AND2X1 U4778 ( .IN1(n25), .IN2(g516), .Q(n4406) );
  OR2X1 U4779 ( .IN1(n4408), .IN2(n4409), .Q(g11336) );
  AND2X1 U4780 ( .IN1(n1239), .IN2(g506), .Q(n4409) );
  AND2X1 U4781 ( .IN1(n25), .IN2(g511), .Q(n4408) );
  OR2X1 U4782 ( .IN1(n4410), .IN2(n4411), .Q(g11335) );
  AND2X1 U4783 ( .IN1(n1239), .IN2(g501), .Q(n4411) );
  AND2X1 U4784 ( .IN1(n25), .IN2(g506), .Q(n4410) );
  OR2X1 U4785 ( .IN1(n4412), .IN2(n4413), .Q(g11334) );
  AND2X1 U4786 ( .IN1(n1239), .IN2(g496), .Q(n4413) );
  AND2X1 U4787 ( .IN1(n25), .IN2(g501), .Q(n4412) );
  OR2X1 U4788 ( .IN1(n4414), .IN2(n4415), .Q(g11333) );
  AND2X1 U4789 ( .IN1(n1239), .IN2(g491), .Q(n4415) );
  AND2X1 U4790 ( .IN1(n25), .IN2(g496), .Q(n4414) );
  OR2X1 U4791 ( .IN1(n4416), .IN2(n4417), .Q(g11332) );
  AND2X1 U4792 ( .IN1(n1239), .IN2(g486), .Q(n4417) );
  AND2X1 U4793 ( .IN1(n25), .IN2(g491), .Q(n4416) );
  OR2X1 U4794 ( .IN1(n4418), .IN2(n4419), .Q(g11331) );
  AND2X1 U4795 ( .IN1(n1239), .IN2(g481), .Q(n4419) );
  AND2X1 U4796 ( .IN1(n25), .IN2(g486), .Q(n4418) );
  OR2X1 U4797 ( .IN1(n4420), .IN2(n4421), .Q(g11330) );
  AND2X1 U4798 ( .IN1(n1239), .IN2(g525), .Q(n4421) );
  AND2X1 U4799 ( .IN1(n25), .IN2(g521), .Q(n4420) );
  OR2X1 U4800 ( .IN1(n4422), .IN2(n4423), .Q(g11329) );
  AND2X1 U4801 ( .IN1(n1239), .IN2(g530), .Q(n4423) );
  AND2X1 U4802 ( .IN1(n25), .IN2(g525), .Q(n4422) );
  OR2X1 U4803 ( .IN1(n4424), .IN2(n4425), .Q(g11328) );
  AND2X1 U4804 ( .IN1(n1239), .IN2(g534), .Q(n4425) );
  AND2X1 U4805 ( .IN1(n25), .IN2(g530), .Q(n4424) );
  OR2X1 U4806 ( .IN1(n4426), .IN2(n4427), .Q(g11327) );
  AND2X1 U4807 ( .IN1(n1239), .IN2(g538), .Q(n4427) );
  AND2X1 U4808 ( .IN1(n25), .IN2(g534), .Q(n4426) );
  OR2X1 U4809 ( .IN1(n4428), .IN2(n4429), .Q(g11326) );
  AND2X1 U4810 ( .IN1(n1239), .IN2(g542), .Q(n4429) );
  AND2X1 U4811 ( .IN1(n25), .IN2(g538), .Q(n4428) );
  OR2X1 U4812 ( .IN1(n4430), .IN2(n4431), .Q(g11325) );
  AND2X1 U4813 ( .IN1(n1239), .IN2(g476), .Q(n4431) );
  AND2X1 U4814 ( .IN1(n25), .IN2(g542), .Q(n4430) );
  OR2X1 U4815 ( .IN1(n4432), .IN2(n4433), .Q(g11324) );
  AND2X1 U4816 ( .IN1(n4154), .IN2(n1239), .Q(n4433) );
  OR2X1 U4817 ( .IN1(n4434), .IN2(n4435), .Q(n4154) );
  AND2X1 U4818 ( .IN1(n1698), .IN2(n4436), .Q(n4435) );
  OR2X1 U4819 ( .IN1(n4437), .IN2(g525), .Q(n4436) );
  AND2X1 U4820 ( .IN1(n4438), .IN2(n4439), .Q(n4437) );
  AND2X1 U4821 ( .IN1(n4440), .IN2(n4441), .Q(n4439) );
  AND2X1 U4822 ( .IN1(n4442), .IN2(n4443), .Q(n4441) );
  AND2X1 U4823 ( .IN1(n1600), .IN2(n1599), .Q(n4443) );
  AND2X1 U4824 ( .IN1(n1621), .IN2(n1620), .Q(n4442) );
  AND2X1 U4825 ( .IN1(n4444), .IN2(n1689), .Q(n4440) );
  AND2X1 U4826 ( .IN1(n1680), .IN2(n1679), .Q(n4444) );
  AND2X1 U4827 ( .IN1(n4445), .IN2(n4446), .Q(n4438) );
  AND2X1 U4828 ( .IN1(n4447), .IN2(n2804), .Q(n4446) );
  AND2X1 U4829 ( .IN1(n1691), .IN2(n1690), .Q(n4447) );
  AND2X1 U4830 ( .IN1(n4448), .IN2(n2807), .Q(n4445) );
  AND2X1 U4831 ( .IN1(n2806), .IN2(n2805), .Q(n4448) );
  AND2X1 U4832 ( .IN1(n1695), .IN2(g521), .Q(n4434) );
  AND2X1 U4833 ( .IN1(n25), .IN2(g481), .Q(n4432) );
  AND2X1 U4834 ( .IN1(n4449), .IN2(n4377), .Q(g11320) );
  AND2X1 U4835 ( .IN1(n4450), .IN2(n4451), .Q(n4449) );
  OR2X1 U4836 ( .IN1(n4452), .IN2(g369), .Q(n4450) );
  AND2X1 U4837 ( .IN1(n1239), .IN2(n4380), .Q(n4452) );
  OR2X1 U4838 ( .IN1(n4453), .IN2(n4454), .Q(g11314) );
  AND2X1 U4839 ( .IN1(n4455), .IN2(g968), .Q(n4454) );
  AND2X1 U4840 ( .IN1(n1855), .IN2(g861), .Q(n4453) );
  OR2X1 U4841 ( .IN1(n4456), .IN2(n4457), .Q(g11312) );
  AND2X1 U4842 ( .IN1(g965), .IN2(n4455), .Q(n4457) );
  AND2X1 U4843 ( .IN1(n1855), .IN2(g857), .Q(n4456) );
  OR2X1 U4844 ( .IN1(n4458), .IN2(n4459), .Q(g11310) );
  AND2X1 U4845 ( .IN1(g962), .IN2(n4455), .Q(n4459) );
  AND2X1 U4846 ( .IN1(n1855), .IN2(g853), .Q(n4458) );
  OR2X1 U4847 ( .IN1(n4460), .IN2(n4461), .Q(g11308) );
  AND2X1 U4848 ( .IN1(n4455), .IN2(g959), .Q(n4461) );
  AND2X1 U4849 ( .IN1(n1855), .IN2(g849), .Q(n4460) );
  OR2X1 U4850 ( .IN1(n4462), .IN2(n4463), .Q(g11306) );
  AND2X1 U4851 ( .IN1(n4455), .IN2(g956), .Q(n4463) );
  AND2X1 U4852 ( .IN1(n1855), .IN2(g845), .Q(n4462) );
  OR2X1 U4853 ( .IN1(n4464), .IN2(n4465), .Q(g11305) );
  AND2X1 U4854 ( .IN1(n4455), .IN2(g953), .Q(n4465) );
  AND2X1 U4855 ( .IN1(n1855), .IN2(g841), .Q(n4464) );
  OR2X1 U4856 ( .IN1(n4466), .IN2(n4467), .Q(g11303) );
  AND2X1 U4857 ( .IN1(n4455), .IN2(g950), .Q(n4467) );
  AND2X1 U4858 ( .IN1(n1855), .IN2(g837), .Q(n4466) );
  OR2X1 U4859 ( .IN1(n4468), .IN2(n4469), .Q(g11300) );
  AND2X1 U4860 ( .IN1(n4455), .IN2(g947), .Q(n4469) );
  AND2X1 U4861 ( .IN1(n1855), .IN2(g833), .Q(n4468) );
  OR2X1 U4862 ( .IN1(n4470), .IN2(n4471), .Q(g11298) );
  AND2X1 U4863 ( .IN1(n1855), .IN2(g829), .Q(n4471) );
  AND2X1 U4864 ( .IN1(n4455), .IN2(g944), .Q(n4470) );
  INVX0 U4865 ( .INP(n1855), .ZN(n4455) );
  OR2X1 U4866 ( .IN1(n4472), .IN2(n4473), .Q(g11294) );
  OR2X1 U4867 ( .IN1(n4474), .IN2(n4475), .Q(n4473) );
  AND2X1 U4868 ( .IN1(n4476), .IN2(n1682), .Q(n4475) );
  AND2X1 U4869 ( .IN1(n926), .IN2(n4477), .Q(n4476) );
  OR2X1 U4870 ( .IN1(n4478), .IN2(n4479), .Q(n4477) );
  OR2X1 U4871 ( .IN1(n3199), .IN2(n3200), .Q(n4479) );
  AND2X1 U4872 ( .IN1(g1828), .IN2(g1814), .Q(n3200) );
  OR2X1 U4873 ( .IN1(n3198), .IN2(n3330), .Q(n4478) );
  AND2X1 U4874 ( .IN1(n3838), .IN2(g1857), .Q(n4474) );
  AND2X1 U4875 ( .IN1(n503), .IN2(n3188), .Q(n3838) );
  INVX0 U4876 ( .INP(n926), .ZN(n503) );
  AND2X1 U4877 ( .IN1(n4480), .IN2(n3569), .Q(n4472) );
  AND2X1 U4878 ( .IN1(n4481), .IN2(n4482), .Q(n4480) );
  OR2X1 U4879 ( .IN1(n1653), .IN2(n4483), .Q(n4482) );
  OR2X1 U4880 ( .IN1(n4484), .IN2(n4485), .Q(n4483) );
  AND2X1 U4881 ( .IN1(n4486), .IN2(n4487), .Q(n4485) );
  OR2X1 U4882 ( .IN1(n4488), .IN2(n4489), .Q(n4486) );
  INVX0 U4883 ( .INP(n4490), .ZN(n4484) );
  OR2X1 U4884 ( .IN1(n4491), .IN2(n4492), .Q(n4490) );
  AND2X1 U4885 ( .IN1(g10721), .IN2(g10722), .Q(n4491) );
  OR2X1 U4886 ( .IN1(g1690), .IN2(n4493), .Q(n4481) );
  OR2X1 U4887 ( .IN1(n4494), .IN2(n4495), .Q(n4493) );
  AND2X1 U4888 ( .IN1(n4496), .IN2(n3805), .Q(n4495) );
  OR2X1 U4889 ( .IN1(n1702), .IN2(n2853), .Q(n3805) );
  OR2X1 U4890 ( .IN1(n1626), .IN2(n2840), .Q(n4496) );
  AND2X1 U4891 ( .IN1(n4497), .IN2(n4498), .Q(n4494) );
  OR2X1 U4892 ( .IN1(n1659), .IN2(n1715), .Q(n4498) );
  OR2X1 U4893 ( .IN1(n2860), .IN2(n2904), .Q(n4497) );
  OR2X1 U4894 ( .IN1(n4499), .IN2(n4500), .Q(g11293) );
  AND2X1 U4895 ( .IN1(n4501), .IN2(n3569), .Q(n4500) );
  OR2X1 U4896 ( .IN1(n4502), .IN2(n4503), .Q(n4501) );
  AND2X1 U4897 ( .IN1(n1653), .IN2(n2841), .Q(n4503) );
  AND2X1 U4898 ( .IN1(n4504), .IN2(g1690), .Q(n4502) );
  AND2X1 U4899 ( .IN1(n4505), .IN2(n3188), .Q(n4499) );
  OR2X1 U4900 ( .IN1(n4506), .IN2(n3198), .Q(n4505) );
  AND2X1 U4901 ( .IN1(n1608), .IN2(n4507), .Q(n3198) );
  AND2X1 U4902 ( .IN1(g1828), .IN2(n1643), .Q(n4507) );
  AND2X1 U4903 ( .IN1(n4508), .IN2(g1854), .Q(n4506) );
  OR2X1 U4904 ( .IN1(n4509), .IN2(n4510), .Q(n4508) );
  OR2X1 U4905 ( .IN1(n4511), .IN2(n3150), .Q(n4510) );
  OR2X1 U4906 ( .IN1(n2902), .IN2(n1873), .Q(n3150) );
  OR2X1 U4907 ( .IN1(n4512), .IN2(n3569), .Q(n2902) );
  INVX0 U4908 ( .INP(n3188), .ZN(n3569) );
  OR2X1 U4909 ( .IN1(n4513), .IN2(n4514), .Q(n3188) );
  OR2X1 U4910 ( .IN1(g1814), .IN2(g1834), .Q(n4514) );
  OR2X1 U4911 ( .IN1(g1828), .IN2(g1822), .Q(n4513) );
  AND2X1 U4912 ( .IN1(n1608), .IN2(g1834), .Q(n4512) );
  AND2X1 U4913 ( .IN1(n4515), .IN2(n4516), .Q(n4511) );
  AND2X1 U4914 ( .IN1(n822), .IN2(n3206), .Q(n4516) );
  INVX0 U4915 ( .INP(n3199), .ZN(n822) );
  AND2X1 U4916 ( .IN1(g1822), .IN2(n1605), .Q(n3199) );
  AND2X1 U4917 ( .IN1(n1380), .IN2(n3600), .Q(n4515) );
  OR2X1 U4918 ( .IN1(n4517), .IN2(n4518), .Q(n3600) );
  OR2X1 U4919 ( .IN1(g1828), .IN2(g1834), .Q(n4518) );
  OR2X1 U4920 ( .IN1(n1608), .IN2(g1840), .Q(n4517) );
  OR2X1 U4921 ( .IN1(n4519), .IN2(n4520), .Q(n4509) );
  AND2X1 U4922 ( .IN1(n1682), .IN2(n4521), .Q(n4520) );
  XNOR2X1 U4923 ( .IN1(n1380), .IN2(n4522), .Q(n4521) );
  AND2X1 U4924 ( .IN1(n4523), .IN2(g1857), .Q(n4519) );
  XNOR2X1 U4925 ( .IN1(n3206), .IN2(n4522), .Q(n4523) );
  INVX0 U4926 ( .INP(n3330), .ZN(n3206) );
  AND2X1 U4927 ( .IN1(g1822), .IN2(n1608), .Q(n3330) );
  AND2X1 U4928 ( .IN1(n4377), .IN2(n4524), .Q(g11292) );
  OR2X1 U4929 ( .IN1(n4525), .IN2(g382), .Q(n4524) );
  AND2X1 U4930 ( .IN1(n4377), .IN2(n4526), .Q(g11291) );
  INVX0 U4931 ( .INP(n4527), .ZN(n4526) );
  AND2X1 U4932 ( .IN1(n4528), .IN2(n4529), .Q(n4527) );
  OR2X1 U4933 ( .IN1(n4525), .IN2(n2739), .Q(n4529) );
  AND2X1 U4934 ( .IN1(n1239), .IN2(n4530), .Q(n4525) );
  AND2X1 U4935 ( .IN1(n4380), .IN2(n4531), .Q(n4530) );
  OR2X1 U4936 ( .IN1(n4532), .IN2(n4451), .Q(n4528) );
  OR2X1 U4937 ( .IN1(n4531), .IN2(n2740), .Q(n4532) );
  INVX0 U4938 ( .INP(n1385), .ZN(n4531) );
  OR2X1 U4939 ( .IN1(n2739), .IN2(n4533), .Q(n1385) );
  OR2X1 U4940 ( .IN1(n2894), .IN2(n2740), .Q(n4533) );
  AND2X1 U4941 ( .IN1(n4534), .IN2(n4377), .Q(g11290) );
  INVX0 U4942 ( .INP(n4535), .ZN(n4377) );
  OR2X1 U4943 ( .IN1(n519), .IN2(g869), .Q(n4535) );
  XOR2X1 U4944 ( .IN1(n4451), .IN2(n2740), .Q(n4534) );
  OR2X1 U4945 ( .IN1(n25), .IN2(n4536), .Q(n4451) );
  OR2X1 U4946 ( .IN1(n2894), .IN2(n1420), .Q(n4536) );
  OR2X1 U4947 ( .IN1(n4537), .IN2(n4538), .Q(g11270) );
  AND2X1 U4948 ( .IN1(n1239), .IN2(g416), .Q(n4538) );
  AND2X1 U4949 ( .IN1(n25), .IN2(g421), .Q(n4537) );
  OR2X1 U4950 ( .IN1(n4539), .IN2(n4540), .Q(g11269) );
  AND2X1 U4951 ( .IN1(n1239), .IN2(g411), .Q(n4540) );
  AND2X1 U4952 ( .IN1(n25), .IN2(g416), .Q(n4539) );
  OR2X1 U4953 ( .IN1(n4541), .IN2(n4542), .Q(g11268) );
  AND2X1 U4954 ( .IN1(n1239), .IN2(g406), .Q(n4542) );
  AND2X1 U4955 ( .IN1(n25), .IN2(g411), .Q(n4541) );
  OR2X1 U4956 ( .IN1(n4543), .IN2(n4544), .Q(g11267) );
  AND2X1 U4957 ( .IN1(n1239), .IN2(g401), .Q(n4544) );
  AND2X1 U4958 ( .IN1(n25), .IN2(g406), .Q(n4543) );
  OR2X1 U4959 ( .IN1(n4545), .IN2(n4546), .Q(g11266) );
  AND2X1 U4960 ( .IN1(n1239), .IN2(g396), .Q(n4546) );
  AND2X1 U4961 ( .IN1(n25), .IN2(g401), .Q(n4545) );
  OR2X1 U4962 ( .IN1(n4547), .IN2(n4548), .Q(g11265) );
  AND2X1 U4963 ( .IN1(n1239), .IN2(g391), .Q(n4548) );
  AND2X1 U4964 ( .IN1(n25), .IN2(g396), .Q(n4547) );
  OR2X1 U4965 ( .IN1(n4549), .IN2(n4550), .Q(g11264) );
  AND2X1 U4966 ( .IN1(n1239), .IN2(g386), .Q(n4550) );
  AND2X1 U4967 ( .IN1(n25), .IN2(g391), .Q(n4549) );
  OR2X1 U4968 ( .IN1(n4551), .IN2(n4552), .Q(g11263) );
  AND2X1 U4969 ( .IN1(n1239), .IN2(g426), .Q(n4552) );
  AND2X1 U4970 ( .IN1(n25), .IN2(g386), .Q(n4551) );
  OR2X1 U4971 ( .IN1(n4553), .IN2(n4554), .Q(g11262) );
  AND2X1 U4972 ( .IN1(n1239), .IN2(g435), .Q(n4554) );
  AND2X1 U4973 ( .IN1(n25), .IN2(g431), .Q(n4553) );
  OR2X1 U4974 ( .IN1(n4555), .IN2(n4556), .Q(g11261) );
  AND2X1 U4975 ( .IN1(n1239), .IN2(g440), .Q(n4556) );
  AND2X1 U4976 ( .IN1(n25), .IN2(g435), .Q(n4555) );
  OR2X1 U4977 ( .IN1(n4557), .IN2(n4558), .Q(g11260) );
  AND2X1 U4978 ( .IN1(n1239), .IN2(g444), .Q(n4558) );
  AND2X1 U4979 ( .IN1(n25), .IN2(g440), .Q(n4557) );
  OR2X1 U4980 ( .IN1(n4559), .IN2(n4560), .Q(g11259) );
  AND2X1 U4981 ( .IN1(n1239), .IN2(g448), .Q(n4560) );
  AND2X1 U4982 ( .IN1(n25), .IN2(g444), .Q(n4559) );
  OR2X1 U4983 ( .IN1(n4561), .IN2(n4562), .Q(g11258) );
  AND2X1 U4984 ( .IN1(n1239), .IN2(g452), .Q(n4562) );
  AND2X1 U4985 ( .IN1(n25), .IN2(g448), .Q(n4561) );
  OR2X1 U4986 ( .IN1(n4563), .IN2(n4564), .Q(g11257) );
  AND2X1 U4987 ( .IN1(n1239), .IN2(g421), .Q(n4564) );
  AND2X1 U4988 ( .IN1(n25), .IN2(g452), .Q(n4563) );
  OR2X1 U4989 ( .IN1(n4565), .IN2(n4566), .Q(g11256) );
  AND2X1 U4990 ( .IN1(n4393), .IN2(n1239), .Q(n4566) );
  INVX0 U4991 ( .INP(n4567), .ZN(n4393) );
  OR2X1 U4992 ( .IN1(n4568), .IN2(n4569), .Q(n4567) );
  AND2X1 U4993 ( .IN1(n4570), .IN2(n1420), .Q(n4569) );
  OR2X1 U4994 ( .IN1(n4571), .IN2(n4572), .Q(n4570) );
  AND2X1 U4995 ( .IN1(n4573), .IN2(n1878), .Q(n4572) );
  AND2X1 U4996 ( .IN1(n1876), .IN2(n4574), .Q(n4573) );
  OR2X1 U4997 ( .IN1(n4575), .IN2(n4576), .Q(n4574) );
  OR2X1 U4998 ( .IN1(n4577), .IN2(n4578), .Q(n4576) );
  OR2X1 U4999 ( .IN1(g391), .IN2(n4579), .Q(n4578) );
  OR2X1 U5000 ( .IN1(g386), .IN2(g426), .Q(n4579) );
  OR2X1 U5001 ( .IN1(g396), .IN2(n4580), .Q(n4577) );
  OR2X1 U5002 ( .IN1(g448), .IN2(g452), .Q(n4580) );
  OR2X1 U5003 ( .IN1(n4581), .IN2(n4582), .Q(n4575) );
  OR2X1 U5004 ( .IN1(g444), .IN2(n4583), .Q(n4582) );
  OR2X1 U5005 ( .IN1(g406), .IN2(g440), .Q(n4583) );
  OR2X1 U5006 ( .IN1(n4584), .IN2(n4585), .Q(n4581) );
  OR2X1 U5007 ( .IN1(g421), .IN2(g416), .Q(n4585) );
  OR2X1 U5008 ( .IN1(g411), .IN2(g401), .Q(n4584) );
  AND2X1 U5009 ( .IN1(g431), .IN2(g435), .Q(n4571) );
  AND2X1 U5010 ( .IN1(n1681), .IN2(n4380), .Q(n4568) );
  INVX0 U5011 ( .INP(n1420), .ZN(n4380) );
  AND2X1 U5012 ( .IN1(n25), .IN2(g426), .Q(n4565) );
  INVX0 U5013 ( .INP(n1239), .ZN(n25) );
  OR2X1 U5014 ( .IN1(n4586), .IN2(n4587), .Q(n1239) );
  OR2X1 U5015 ( .IN1(n4588), .IN2(n4589), .Q(n4587) );
  OR2X1 U5016 ( .IN1(g849), .IN2(g845), .Q(n4589) );
  OR2X1 U5017 ( .IN1(g853), .IN2(n4590), .Q(n4588) );
  OR2X1 U5018 ( .IN1(g841), .IN2(g857), .Q(n4590) );
  OR2X1 U5019 ( .IN1(n4591), .IN2(n4592), .Q(n4586) );
  OR2X1 U5020 ( .IN1(g837), .IN2(g861), .Q(n4592) );
  OR2X1 U5021 ( .IN1(g833), .IN2(n4593), .Q(n4591) );
  OR2X1 U5022 ( .IN1(n4594), .IN2(g829), .Q(n4593) );
  AND2X1 U5023 ( .IN1(n4595), .IN2(n4596), .Q(n4594) );
  OR2X1 U5024 ( .IN1(n519), .IN2(n4597), .Q(n4596) );
  AND2X1 U5025 ( .IN1(n4598), .IN2(n4599), .Q(n4597) );
  AND2X1 U5026 ( .IN1(n4600), .IN2(n4601), .Q(n4595) );
  AND2X1 U5027 ( .IN1(g10628), .IN2(n4602), .Q(g11206) );
  XOR2X1 U5028 ( .IN1(n4602), .IN2(n2895), .Q(g11163) );
  INVX0 U5029 ( .INP(n4603), .ZN(n4602) );
  OR2X1 U5030 ( .IN1(n4604), .IN2(n4605), .Q(n4603) );
  OR2X1 U5031 ( .IN1(n4606), .IN2(n4607), .Q(n4605) );
  AND2X1 U5032 ( .IN1(n4147), .IN2(g10724), .Q(n4607) );
  INVX0 U5033 ( .INP(n4031), .ZN(n4147) );
  OR2X1 U5034 ( .IN1(n3050), .IN2(n4608), .Q(n4031) );
  OR2X1 U5035 ( .IN1(n2629), .IN2(n519), .Q(n4608) );
  AND2X1 U5036 ( .IN1(n4609), .IN2(g109), .Q(n4606) );
  OR2X1 U5037 ( .IN1(n4610), .IN2(n4611), .Q(n4609) );
  OR2X1 U5038 ( .IN1(n4612), .IN2(n4613), .Q(n4611) );
  AND2X1 U5039 ( .IN1(g10664), .IN2(g2648), .Q(n4613) );
  AND2X1 U5040 ( .IN1(n4614), .IN2(n3036), .Q(n4612) );
  AND2X1 U5041 ( .IN1(n2893), .IN2(g10726), .Q(n4610) );
  AND2X1 U5042 ( .IN1(g5392), .IN2(g10663), .Q(n4604) );
  AND2X1 U5043 ( .IN1(g109), .IN2(n4104), .Q(g5392) );
  INVX0 U5044 ( .INP(n4103), .ZN(n4104) );
  OR2X1 U5045 ( .IN1(n2885), .IN2(n2886), .Q(n4103) );
  OR2X1 U5046 ( .IN1(n4615), .IN2(n4616), .Q(g10936) );
  AND2X1 U5047 ( .IN1(n1391), .IN2(n2903), .Q(n4616) );
  OR2X1 U5048 ( .IN1(n4617), .IN2(n4618), .Q(n1391) );
  OR2X1 U5049 ( .IN1(n4619), .IN2(n4601), .Q(n4618) );
  INVX0 U5050 ( .INP(n4614), .ZN(n4601) );
  OR2X1 U5051 ( .IN1(g10721), .IN2(n4258), .Q(n4617) );
  INVX0 U5052 ( .INP(n4620), .ZN(n4258) );
  INVX0 U5053 ( .INP(n4621), .ZN(n4615) );
  OR2X1 U5054 ( .IN1(n2903), .IN2(n1699), .Q(n4621) );
  OR2X1 U5055 ( .IN1(n4622), .IN2(n4623), .Q(g10898) );
  AND2X1 U5056 ( .IN1(n4624), .IN2(n3451), .Q(n4623) );
  OR2X1 U5057 ( .IN1(n4128), .IN2(n4625), .Q(n4624) );
  XOR2X1 U5058 ( .IN1(n4626), .IN2(n4627), .Q(n4625) );
  XNOR2X1 U5059 ( .IN1(test_so8), .IN2(g1019), .Q(n4627) );
  XOR2X1 U5060 ( .IN1(n4628), .IN2(n4629), .Q(n4626) );
  XOR2X1 U5061 ( .IN1(n4630), .IN2(n4631), .Q(n4629) );
  XNOR2X1 U5062 ( .IN1(g1023), .IN2(n1871), .Q(n4631) );
  XNOR2X1 U5063 ( .IN1(g1011), .IN2(n2741), .Q(n4630) );
  XOR2X1 U5064 ( .IN1(n4632), .IN2(n4633), .Q(n4628) );
  XNOR2X1 U5065 ( .IN1(g1003), .IN2(n2812), .Q(n4633) );
  XOR2X1 U5066 ( .IN1(test_so2), .IN2(n2845), .Q(n4632) );
  AND2X1 U5067 ( .IN1(n4634), .IN2(n4620), .Q(n4128) );
  OR2X1 U5068 ( .IN1(n3155), .IN2(n4635), .Q(n4620) );
  OR2X1 U5069 ( .IN1(g46), .IN2(n4636), .Q(n4635) );
  OR2X1 U5070 ( .IN1(n4637), .IN2(n3152), .Q(n3155) );
  OR2X1 U5071 ( .IN1(n4638), .IN2(n4639), .Q(n3152) );
  OR2X1 U5072 ( .IN1(g44), .IN2(g43), .Q(n4639) );
  OR2X1 U5073 ( .IN1(g48), .IN2(g45), .Q(n4638) );
  INVX0 U5074 ( .INP(n4640), .ZN(n4622) );
  OR2X1 U5075 ( .IN1(n3451), .IN2(n2893), .Q(n4640) );
  OR2X1 U5076 ( .IN1(n4641), .IN2(n4642), .Q(g10866) );
  AND2X1 U5077 ( .IN1(n371), .IN2(g1684), .Q(n4641) );
  OR2X1 U5078 ( .IN1(n4643), .IN2(n4644), .Q(g10865) );
  AND2X1 U5079 ( .IN1(n4645), .IN2(n3992), .Q(n4644) );
  AND2X1 U5080 ( .IN1(n1404), .IN2(n4646), .Q(n4645) );
  OR2X1 U5081 ( .IN1(n519), .IN2(g10722), .Q(n4646) );
  AND2X1 U5082 ( .IN1(n3991), .IN2(g1669), .Q(n4643) );
  OR2X1 U5083 ( .IN1(n4647), .IN2(n4648), .Q(g10864) );
  AND2X1 U5084 ( .IN1(n371), .IN2(g1681), .Q(n4647) );
  OR2X1 U5085 ( .IN1(n4649), .IN2(n4650), .Q(g10863) );
  AND2X1 U5086 ( .IN1(n4651), .IN2(n3992), .Q(n4650) );
  AND2X1 U5087 ( .IN1(n4652), .IN2(n4653), .Q(n4651) );
  OR2X1 U5088 ( .IN1(n4654), .IN2(g1718), .Q(n4652) );
  AND2X1 U5089 ( .IN1(n3991), .IN2(g1666), .Q(n4649) );
  OR2X1 U5090 ( .IN1(n4655), .IN2(n4656), .Q(g10862) );
  AND2X1 U5091 ( .IN1(n371), .IN2(g1678), .Q(n4655) );
  OR2X1 U5092 ( .IN1(n4657), .IN2(n4658), .Q(g10861) );
  AND2X1 U5093 ( .IN1(n4659), .IN2(n3992), .Q(n4658) );
  AND2X1 U5094 ( .IN1(n3991), .IN2(g1663), .Q(n4657) );
  OR2X1 U5095 ( .IN1(n4660), .IN2(n4661), .Q(g10860) );
  AND2X1 U5096 ( .IN1(n371), .IN2(g1675), .Q(n4660) );
  OR2X1 U5097 ( .IN1(n4662), .IN2(n4663), .Q(g10859) );
  AND2X1 U5098 ( .IN1(n4664), .IN2(n3992), .Q(n4663) );
  AND2X1 U5099 ( .IN1(n3991), .IN2(g1660), .Q(n4662) );
  OR2X1 U5100 ( .IN1(n4665), .IN2(n4666), .Q(g10858) );
  AND2X1 U5101 ( .IN1(n371), .IN2(g1672), .Q(n4665) );
  OR2X1 U5102 ( .IN1(n4667), .IN2(n4668), .Q(g10855) );
  AND2X1 U5103 ( .IN1(n4659), .IN2(n3451), .Q(n4668) );
  OR2X1 U5104 ( .IN1(n4669), .IN2(n4670), .Q(n4659) );
  AND2X1 U5105 ( .IN1(n3676), .IN2(n4671), .Q(n4670) );
  OR2X1 U5106 ( .IN1(n4009), .IN2(n4672), .Q(n3676) );
  AND2X1 U5107 ( .IN1(n3471), .IN2(g1512), .Q(n4672) );
  AND2X1 U5108 ( .IN1(g18), .IN2(g192), .Q(n4009) );
  AND2X1 U5109 ( .IN1(n4673), .IN2(n4653), .Q(n4669) );
  OR2X1 U5110 ( .IN1(n4674), .IN2(g1718), .Q(n4673) );
  AND2X1 U5111 ( .IN1(n371), .IN2(g549), .Q(n4667) );
  OR2X1 U5112 ( .IN1(n2895), .IN2(n3141), .Q(g10801) );
  XOR2X1 U5113 ( .IN1(n4675), .IN2(n4676), .Q(n2895) );
  XOR2X1 U5114 ( .IN1(n4677), .IN2(n4678), .Q(n4676) );
  OR2X1 U5115 ( .IN1(n4679), .IN2(g32), .Q(n4678) );
  INVX0 U5116 ( .INP(n4680), .ZN(n4679) );
  OR2X1 U5117 ( .IN1(n4598), .IN2(n4681), .Q(n4677) );
  OR2X1 U5118 ( .IN1(n4682), .IN2(n4683), .Q(n4681) );
  INVX0 U5119 ( .INP(n4684), .ZN(n4683) );
  OR2X1 U5120 ( .IN1(n4487), .IN2(g10726), .Q(n4684) );
  OR2X1 U5121 ( .IN1(n4634), .IN2(n4685), .Q(n4487) );
  AND2X1 U5122 ( .IN1(n4686), .IN2(g10726), .Q(n4682) );
  XNOR2X1 U5123 ( .IN1(g10663), .IN2(n4685), .Q(n4686) );
  AND2X1 U5124 ( .IN1(n4634), .IN2(n4687), .Q(n4598) );
  AND2X1 U5125 ( .IN1(n4489), .IN2(n4685), .Q(n4687) );
  INVX0 U5126 ( .INP(g10664), .ZN(n4685) );
  INVX0 U5127 ( .INP(g10726), .ZN(n4489) );
  INVX0 U5128 ( .INP(g10663), .ZN(n4634) );
  XNOR2X1 U5129 ( .IN1(n4688), .IN2(n1858), .Q(n4675) );
  XNOR2X1 U5130 ( .IN1(g10721), .IN2(g10722), .Q(n1858) );
  OR2X1 U5131 ( .IN1(n4599), .IN2(n4689), .Q(n4688) );
  OR2X1 U5132 ( .IN1(n4690), .IN2(n4691), .Q(n4689) );
  AND2X1 U5133 ( .IN1(n4492), .IN2(n4488), .Q(n4691) );
  AND2X1 U5134 ( .IN1(g10719), .IN2(g10720), .Q(n4492) );
  AND2X1 U5135 ( .IN1(n4692), .IN2(g10724), .Q(n4690) );
  XNOR2X1 U5136 ( .IN1(g10720), .IN2(n4504), .Q(n4692) );
  INVX0 U5137 ( .INP(g10719), .ZN(n4504) );
  INVX0 U5138 ( .INP(n4619), .ZN(n4599) );
  OR2X1 U5139 ( .IN1(g10719), .IN2(n4693), .Q(n4619) );
  OR2X1 U5140 ( .IN1(g10724), .IN2(g10720), .Q(n4693) );
  OR2X1 U5141 ( .IN1(n4694), .IN2(n4695), .Q(g10800) );
  AND2X1 U5142 ( .IN1(n4664), .IN2(n3451), .Q(n4695) );
  OR2X1 U5143 ( .IN1(n4696), .IN2(n4697), .Q(n4664) );
  AND2X1 U5144 ( .IN1(n3671), .IN2(n4671), .Q(n4697) );
  OR2X1 U5145 ( .IN1(n4011), .IN2(n4698), .Q(n3671) );
  AND2X1 U5146 ( .IN1(n3471), .IN2(g1636), .Q(n4698) );
  AND2X1 U5147 ( .IN1(g18), .IN2(g248), .Q(n4011) );
  AND2X1 U5148 ( .IN1(n4699), .IN2(n4653), .Q(n4696) );
  OR2X1 U5149 ( .IN1(g10719), .IN2(n4700), .Q(n4699) );
  AND2X1 U5150 ( .IN1(n371), .IN2(g575), .Q(n4694) );
  OR2X1 U5151 ( .IN1(n4701), .IN2(n4702), .Q(g10799) );
  AND2X1 U5152 ( .IN1(n371), .IN2(g566), .Q(n4701) );
  OR2X1 U5153 ( .IN1(n4703), .IN2(n4642), .Q(g10798) );
  AND2X1 U5154 ( .IN1(n4704), .IN2(n3451), .Q(n4642) );
  OR2X1 U5155 ( .IN1(n4705), .IN2(n4706), .Q(n4704) );
  AND2X1 U5156 ( .IN1(n1404), .IN2(n4707), .Q(n4706) );
  AND2X1 U5157 ( .IN1(n4671), .IN2(n3674), .Q(n4705) );
  OR2X1 U5158 ( .IN1(n4708), .IN2(n3478), .Q(n3674) );
  AND2X1 U5159 ( .IN1(g225), .IN2(g18), .Q(n3478) );
  AND2X1 U5160 ( .IN1(n3471), .IN2(g1624), .Q(n4708) );
  AND2X1 U5161 ( .IN1(n371), .IN2(g563), .Q(n4703) );
  OR2X1 U5162 ( .IN1(n4709), .IN2(n4648), .Q(g10797) );
  AND2X1 U5163 ( .IN1(n4710), .IN2(n3451), .Q(n4648) );
  OR2X1 U5164 ( .IN1(n4711), .IN2(n4712), .Q(n4710) );
  AND2X1 U5165 ( .IN1(n1404), .IN2(n4614), .Q(n4712) );
  AND2X1 U5166 ( .IN1(n4671), .IN2(n3669), .Q(n4711) );
  OR2X1 U5167 ( .IN1(n4713), .IN2(n3462), .Q(n3669) );
  AND2X1 U5168 ( .IN1(g219), .IN2(g18), .Q(n3462) );
  AND2X1 U5169 ( .IN1(n3471), .IN2(g1621), .Q(n4713) );
  AND2X1 U5170 ( .IN1(n371), .IN2(g560), .Q(n4709) );
  OR2X1 U5171 ( .IN1(n4714), .IN2(n4656), .Q(g10795) );
  AND2X1 U5172 ( .IN1(n4715), .IN2(n3451), .Q(n4656) );
  OR2X1 U5173 ( .IN1(n4716), .IN2(n4717), .Q(n4715) );
  AND2X1 U5174 ( .IN1(n1404), .IN2(n4654), .Q(n4717) );
  AND2X1 U5175 ( .IN1(n4671), .IN2(n3661), .Q(n4716) );
  OR2X1 U5176 ( .IN1(n4718), .IN2(n3524), .Q(n3661) );
  AND2X1 U5177 ( .IN1(g213), .IN2(g18), .Q(n3524) );
  AND2X1 U5178 ( .IN1(n3471), .IN2(g1615), .Q(n4718) );
  AND2X1 U5179 ( .IN1(n371), .IN2(g557), .Q(n4714) );
  OR2X1 U5180 ( .IN1(n4719), .IN2(n4661), .Q(g10793) );
  AND2X1 U5181 ( .IN1(n3451), .IN2(n4720), .Q(n4661) );
  AND2X1 U5182 ( .IN1(n4721), .IN2(n4722), .Q(n4720) );
  OR2X1 U5183 ( .IN1(n3657), .IN2(n4653), .Q(n4722) );
  OR2X1 U5184 ( .IN1(n4723), .IN2(n3512), .Q(n3657) );
  AND2X1 U5185 ( .IN1(g207), .IN2(g18), .Q(n3512) );
  AND2X1 U5186 ( .IN1(n3471), .IN2(g1639), .Q(n4723) );
  OR2X1 U5187 ( .IN1(n4724), .IN2(n4671), .Q(n4721) );
  OR2X1 U5188 ( .IN1(n4700), .IN2(g10720), .Q(n4724) );
  OR2X1 U5189 ( .IN1(n519), .IN2(g1718), .Q(n4700) );
  AND2X1 U5190 ( .IN1(n371), .IN2(g554), .Q(n4719) );
  OR2X1 U5191 ( .IN1(n4725), .IN2(n4666), .Q(g10791) );
  AND2X1 U5192 ( .IN1(n3451), .IN2(n4726), .Q(n4666) );
  OR2X1 U5193 ( .IN1(n4727), .IN2(n4728), .Q(n4726) );
  AND2X1 U5194 ( .IN1(n1404), .IN2(n4729), .Q(n4728) );
  AND2X1 U5195 ( .IN1(n3678), .IN2(n4671), .Q(n4727) );
  OR2X1 U5196 ( .IN1(n4730), .IN2(n3494), .Q(n3678) );
  AND2X1 U5197 ( .IN1(g186), .IN2(g18), .Q(n3494) );
  AND2X1 U5198 ( .IN1(n3471), .IN2(g1618), .Q(n4730) );
  AND2X1 U5199 ( .IN1(n371), .IN2(g546), .Q(n4725) );
  AND2X1 U5200 ( .IN1(n369), .IN2(n3023), .Q(g10785) );
  AND2X1 U5201 ( .IN1(n369), .IN2(n3029), .Q(g10784) );
  AND2X1 U5202 ( .IN1(n369), .IN2(n3065), .Q(g10782) );
  AND2X1 U5203 ( .IN1(n369), .IN2(n3017), .Q(g10780) );
  INVX0 U5204 ( .INP(n2903), .ZN(n369) );
  AND2X1 U5205 ( .IN1(n2852), .IN2(g1696), .Q(n2903) );
  OR2X1 U5206 ( .IN1(n4731), .IN2(n4702), .Q(g10776) );
  AND2X1 U5207 ( .IN1(n3451), .IN2(n4732), .Q(n4702) );
  OR2X1 U5208 ( .IN1(n4733), .IN2(n4734), .Q(n4732) );
  AND2X1 U5209 ( .IN1(g10726), .IN2(n1404), .Q(n4734) );
  OR2X1 U5210 ( .IN1(n4735), .IN2(n1450), .Q(n4733) );
  AND2X1 U5211 ( .IN1(n3680), .IN2(n4671), .Q(n4735) );
  OR2X1 U5212 ( .IN1(n4736), .IN2(n3506), .Q(n3680) );
  AND2X1 U5213 ( .IN1(g231), .IN2(g18), .Q(n3506) );
  AND2X1 U5214 ( .IN1(n3471), .IN2(g1627), .Q(n4736) );
  AND2X1 U5215 ( .IN1(n371), .IN2(g1687), .Q(n4731) );
  OR2X1 U5216 ( .IN1(n4737), .IN2(n4738), .Q(g10773) );
  AND2X1 U5217 ( .IN1(n4094), .IN2(g1727), .Q(n4738) );
  AND2X1 U5218 ( .IN1(n4739), .IN2(n4654), .Q(n4737) );
  OR2X1 U5219 ( .IN1(n4740), .IN2(n4741), .Q(g10771) );
  AND2X1 U5220 ( .IN1(n4674), .IN2(n4739), .Q(n4741) );
  AND2X1 U5221 ( .IN1(g109), .IN2(g10720), .Q(n4674) );
  AND2X1 U5222 ( .IN1(n4094), .IN2(g1724), .Q(n4740) );
  OR2X1 U5223 ( .IN1(n4742), .IN2(n4743), .Q(g10770) );
  AND2X1 U5224 ( .IN1(n4729), .IN2(n4739), .Q(n4743) );
  AND2X1 U5225 ( .IN1(g109), .IN2(g10719), .Q(n4729) );
  AND2X1 U5226 ( .IN1(n4094), .IN2(g1721), .Q(n4742) );
  OR2X1 U5227 ( .IN1(n4744), .IN2(n4745), .Q(g10767) );
  AND2X1 U5228 ( .IN1(n4746), .IN2(n3992), .Q(n4745) );
  AND2X1 U5229 ( .IN1(n3991), .IN2(g1657), .Q(n4744) );
  OR2X1 U5230 ( .IN1(n4747), .IN2(n4748), .Q(g10765) );
  AND2X1 U5231 ( .IN1(n3992), .IN2(n4749), .Q(n4748) );
  INVX0 U5232 ( .INP(n3991), .ZN(n3992) );
  AND2X1 U5233 ( .IN1(n3991), .IN2(g1654), .Q(n4747) );
  OR2X1 U5234 ( .IN1(g1696), .IN2(n2852), .Q(n3991) );
  OR2X1 U5235 ( .IN1(n4750), .IN2(n4751), .Q(g10718) );
  AND2X1 U5236 ( .IN1(n4746), .IN2(n3451), .Q(n4751) );
  OR2X1 U5237 ( .IN1(n4752), .IN2(n4753), .Q(n4746) );
  AND2X1 U5238 ( .IN1(n3663), .IN2(n4671), .Q(n4753) );
  OR2X1 U5239 ( .IN1(n4013), .IN2(n4754), .Q(n3663) );
  AND2X1 U5240 ( .IN1(n3471), .IN2(g1633), .Q(n4754) );
  AND2X1 U5241 ( .IN1(g18), .IN2(g243), .Q(n4013) );
  AND2X1 U5242 ( .IN1(n4755), .IN2(n4653), .Q(n4752) );
  OR2X1 U5243 ( .IN1(n4756), .IN2(g1718), .Q(n4755) );
  AND2X1 U5244 ( .IN1(g10664), .IN2(g109), .Q(n4756) );
  AND2X1 U5245 ( .IN1(n371), .IN2(g572), .Q(n4750) );
  OR2X1 U5246 ( .IN1(n4757), .IN2(n4758), .Q(g10717) );
  AND2X1 U5247 ( .IN1(n4749), .IN2(n3451), .Q(n4758) );
  OR2X1 U5248 ( .IN1(n4759), .IN2(n4760), .Q(n4749) );
  OR2X1 U5249 ( .IN1(n1450), .IN2(n4761), .Q(n4760) );
  AND2X1 U5250 ( .IN1(n4671), .IN2(n3682), .Q(n4761) );
  OR2X1 U5251 ( .IN1(n4762), .IN2(n3518), .Q(n3682) );
  AND2X1 U5252 ( .IN1(g237), .IN2(g18), .Q(n3518) );
  AND2X1 U5253 ( .IN1(n3471), .IN2(g1630), .Q(n4762) );
  INVX0 U5254 ( .INP(g18), .ZN(n3471) );
  AND2X1 U5255 ( .IN1(n1404), .IN2(g10663), .Q(n4759) );
  AND2X1 U5256 ( .IN1(n4653), .IN2(n1611), .Q(n1404) );
  INVX0 U5257 ( .INP(n4671), .ZN(n4653) );
  AND2X1 U5258 ( .IN1(n1611), .IN2(n5141), .Q(n4671) );
  AND2X1 U5259 ( .IN1(n371), .IN2(g569), .Q(n4757) );
  INVX0 U5260 ( .INP(n3451), .ZN(n371) );
  AND2X1 U5261 ( .IN1(n3864), .IN2(n2852), .Q(n3451) );
  OR2X1 U5262 ( .IN1(n4763), .IN2(n4764), .Q(g10711) );
  AND2X1 U5263 ( .IN1(n4739), .IN2(n4707), .Q(n4764) );
  INVX0 U5264 ( .INP(n4522), .ZN(n4707) );
  AND2X1 U5265 ( .IN1(g109), .IN2(n4488), .Q(n4522) );
  INVX0 U5266 ( .INP(g10724), .ZN(n4488) );
  AND2X1 U5267 ( .IN1(n4094), .IN2(g1733), .Q(n4763) );
  OR2X1 U5268 ( .IN1(n4765), .IN2(n4766), .Q(g10707) );
  AND2X1 U5269 ( .IN1(n4094), .IN2(g1730), .Q(n4766) );
  AND2X1 U5270 ( .IN1(n4739), .IN2(n4614), .Q(n4765) );
  INVX0 U5271 ( .INP(n4094), .ZN(n4739) );
  OR2X1 U5272 ( .IN1(n2852), .IN2(n3864), .Q(n4094) );
  INVX0 U5273 ( .INP(g1696), .ZN(n3864) );
  OR2X1 U5274 ( .IN1(n4767), .IN2(n4768), .Q(g10664) );
  OR2X1 U5275 ( .IN1(n4769), .IN2(n4770), .Q(n4768) );
  OR2X1 U5276 ( .IN1(n4771), .IN2(n4772), .Q(n4770) );
  OR2X1 U5277 ( .IN1(n4773), .IN2(n4774), .Q(n4772) );
  AND2X1 U5278 ( .IN1(g1191), .IN2(n4775), .Q(n4774) );
  AND2X1 U5279 ( .IN1(n4776), .IN2(n4777), .Q(n4773) );
  INVX0 U5280 ( .INP(n4775), .ZN(n4777) );
  AND2X1 U5281 ( .IN1(n4778), .IN2(n4779), .Q(n4776) );
  INVX0 U5282 ( .INP(n4780), .ZN(n4779) );
  OR2X1 U5283 ( .IN1(n4781), .IN2(n4782), .Q(n4780) );
  OR2X1 U5284 ( .IN1(n1480), .IN2(n1479), .Q(n4781) );
  AND2X1 U5285 ( .IN1(n4783), .IN2(n1478), .Q(n4778) );
  AND2X1 U5286 ( .IN1(n4784), .IN2(n4785), .Q(n4783) );
  INVX0 U5287 ( .INP(n4786), .ZN(n4785) );
  OR2X1 U5288 ( .IN1(n4787), .IN2(n4788), .Q(n4784) );
  AND2X1 U5289 ( .IN1(n4789), .IN2(n4790), .Q(n4787) );
  AND2X1 U5290 ( .IN1(test_so9), .IN2(n4782), .Q(n4771) );
  OR2X1 U5291 ( .IN1(n4791), .IN2(n4792), .Q(n4769) );
  AND2X1 U5292 ( .IN1(n4786), .IN2(g1741), .Q(n4792) );
  AND2X1 U5293 ( .IN1(n1486), .IN2(g1546), .Q(n4791) );
  OR2X1 U5294 ( .IN1(n4793), .IN2(n4794), .Q(n4767) );
  OR2X1 U5295 ( .IN1(n4795), .IN2(n4796), .Q(n4794) );
  AND2X1 U5296 ( .IN1(n1485), .IN2(g1589), .Q(n4796) );
  AND2X1 U5297 ( .IN1(n4680), .IN2(n3040), .Q(n4795) );
  OR2X1 U5298 ( .IN1(n4797), .IN2(n4798), .Q(n4793) );
  OR2X1 U5299 ( .IN1(n4799), .IN2(n4800), .Q(n4798) );
  AND2X1 U5300 ( .IN1(g919), .IN2(n4801), .Q(n4800) );
  AND2X1 U5301 ( .IN1(n4802), .IN2(g284), .Q(n4799) );
  AND2X1 U5302 ( .IN1(n4803), .IN2(g947), .Q(n4797) );
  AND2X1 U5303 ( .IN1(n4804), .IN2(n4805), .Q(g10628) );
  OR2X1 U5304 ( .IN1(n4600), .IN2(n3652), .Q(n4805) );
  OR2X1 U5305 ( .IN1(n3058), .IN2(n4806), .Q(n3652) );
  OR2X1 U5306 ( .IN1(n2628), .IN2(n519), .Q(n4806) );
  INVX0 U5307 ( .INP(n4654), .ZN(n4600) );
  AND2X1 U5308 ( .IN1(g109), .IN2(g10721), .Q(n4654) );
  OR2X1 U5309 ( .IN1(n4807), .IN2(n519), .Q(n4804) );
  INVX0 U5310 ( .INP(g109), .ZN(n519) );
  INVX0 U5311 ( .INP(n4808), .ZN(n4807) );
  OR2X1 U5312 ( .IN1(n4809), .IN2(n4810), .Q(n4808) );
  OR2X1 U5313 ( .IN1(n4811), .IN2(n4812), .Q(n4810) );
  AND2X1 U5314 ( .IN1(g881), .IN2(g10720), .Q(n4812) );
  AND2X1 U5315 ( .IN1(g877), .IN2(g10719), .Q(n4811) );
  OR2X1 U5316 ( .IN1(n4813), .IN2(n4814), .Q(n4809) );
  AND2X1 U5317 ( .IN1(n3064), .IN2(n4614), .Q(n4814) );
  AND2X1 U5318 ( .IN1(g109), .IN2(g10722), .Q(n4614) );
  OR2X1 U5319 ( .IN1(n4815), .IN2(n4816), .Q(g10722) );
  OR2X1 U5320 ( .IN1(n4817), .IN2(n4818), .Q(n4816) );
  OR2X1 U5321 ( .IN1(n4819), .IN2(n4820), .Q(n4818) );
  OR2X1 U5322 ( .IN1(n4821), .IN2(n4822), .Q(n4820) );
  AND2X1 U5323 ( .IN1(n1486), .IN2(g1534), .Q(n4822) );
  AND2X1 U5324 ( .IN1(n1485), .IN2(g1577), .Q(n4821) );
  OR2X1 U5325 ( .IN1(n4823), .IN2(n4824), .Q(n4819) );
  OR2X1 U5326 ( .IN1(n4825), .IN2(n4826), .Q(n4824) );
  AND2X1 U5327 ( .IN1(g1203), .IN2(n1512), .Q(n4826) );
  AND2X1 U5328 ( .IN1(n1480), .IN2(g1601), .Q(n4825) );
  AND2X1 U5329 ( .IN1(n1479), .IN2(g1558), .Q(n4823) );
  OR2X1 U5330 ( .IN1(n4827), .IN2(n4828), .Q(n4817) );
  OR2X1 U5331 ( .IN1(n4829), .IN2(n4830), .Q(n4828) );
  AND2X1 U5332 ( .IN1(n4680), .IN2(n3048), .Q(n4830) );
  AND2X1 U5333 ( .IN1(n4831), .IN2(g1753), .Q(n4829) );
  OR2X1 U5334 ( .IN1(n4832), .IN2(n4833), .Q(n4827) );
  OR2X1 U5335 ( .IN1(n4834), .IN2(n4835), .Q(n4833) );
  AND2X1 U5336 ( .IN1(g1179), .IN2(n4775), .Q(n4835) );
  AND2X1 U5337 ( .IN1(n4836), .IN2(g1324), .Q(n4834) );
  AND2X1 U5338 ( .IN1(n4786), .IN2(g1730), .Q(n4832) );
  OR2X1 U5339 ( .IN1(n4837), .IN2(n4838), .Q(n4815) );
  OR2X1 U5340 ( .IN1(n4839), .IN2(n4840), .Q(n4838) );
  OR2X1 U5341 ( .IN1(n4841), .IN2(n4842), .Q(n4840) );
  AND2X1 U5342 ( .IN1(n4782), .IN2(g1351), .Q(n4842) );
  AND2X1 U5343 ( .IN1(n4803), .IN2(g986), .Q(n4841) );
  OR2X1 U5344 ( .IN1(n4843), .IN2(n4844), .Q(n4839) );
  OR2X1 U5345 ( .IN1(n4845), .IN2(n4846), .Q(n4844) );
  AND2X1 U5346 ( .IN1(n4847), .IN2(g296), .Q(n4846) );
  AND2X1 U5347 ( .IN1(n4802), .IN2(g272), .Q(n4845) );
  AND2X1 U5348 ( .IN1(g907), .IN2(n4801), .Q(n4843) );
  OR2X1 U5349 ( .IN1(n4848), .IN2(n4849), .Q(n4837) );
  OR2X1 U5350 ( .IN1(n4850), .IN2(n4851), .Q(n4849) );
  OR2X1 U5351 ( .IN1(n4852), .IN2(n4853), .Q(n4851) );
  AND2X1 U5352 ( .IN1(n4854), .IN2(g8), .Q(n4853) );
  AND2X1 U5353 ( .IN1(g895), .IN2(n4855), .Q(n4852) );
  AND2X1 U5354 ( .IN1(n4856), .IN2(n1631), .Q(n4850) );
  OR2X1 U5355 ( .IN1(n4857), .IN2(n4858), .Q(n4848) );
  OR2X1 U5356 ( .IN1(n4859), .IN2(n4860), .Q(n4858) );
  AND2X1 U5357 ( .IN1(n4861), .IN2(g940), .Q(n4860) );
  AND2X1 U5358 ( .IN1(n3140), .IN2(g959), .Q(n4857) );
  AND2X1 U5359 ( .IN1(n4862), .IN2(n5139), .Q(n4813) );
  AND2X1 U5360 ( .IN1(g10724), .IN2(g3007), .Q(n4862) );
  OR2X1 U5361 ( .IN1(g10726), .IN2(n3141), .Q(g10465) );
  OR2X1 U5362 ( .IN1(n4863), .IN2(n4864), .Q(g10726) );
  OR2X1 U5363 ( .IN1(n4865), .IN2(n4866), .Q(n4864) );
  OR2X1 U5364 ( .IN1(n4867), .IN2(n4868), .Q(n4866) );
  OR2X1 U5365 ( .IN1(n4869), .IN2(n4870), .Q(n4868) );
  AND2X1 U5366 ( .IN1(n1485), .IN2(g1583), .Q(n4870) );
  AND2X1 U5367 ( .IN1(n1479), .IN2(g1564), .Q(n4869) );
  AND2X1 U5368 ( .IN1(n1486), .IN2(g1540), .Q(n4867) );
  OR2X1 U5369 ( .IN1(n4871), .IN2(n4872), .Q(n4865) );
  OR2X1 U5370 ( .IN1(n4873), .IN2(n4874), .Q(n4872) );
  AND2X1 U5371 ( .IN1(n4680), .IN2(n1650), .Q(n4874) );
  AND2X1 U5372 ( .IN1(n4831), .IN2(g1759), .Q(n4873) );
  AND2X1 U5373 ( .IN1(n1480), .IN2(g1607), .Q(n4871) );
  OR2X1 U5374 ( .IN1(n4875), .IN2(n4876), .Q(n4863) );
  OR2X1 U5375 ( .IN1(n4877), .IN2(n4878), .Q(n4876) );
  OR2X1 U5376 ( .IN1(n4879), .IN2(n4880), .Q(n4878) );
  AND2X1 U5377 ( .IN1(n4836), .IN2(g1330), .Q(n4880) );
  AND2X1 U5378 ( .IN1(g1185), .IN2(n4775), .Q(n4877) );
  OR2X1 U5379 ( .IN1(n4881), .IN2(n4882), .Q(n4875) );
  OR2X1 U5380 ( .IN1(n4883), .IN2(n4884), .Q(n4882) );
  AND2X1 U5381 ( .IN1(g913), .IN2(n4801), .Q(n4884) );
  AND2X1 U5382 ( .IN1(n4847), .IN2(g302), .Q(n4883) );
  OR2X1 U5383 ( .IN1(n4885), .IN2(n4886), .Q(n4881) );
  AND2X1 U5384 ( .IN1(n4802), .IN2(g278), .Q(n4886) );
  AND2X1 U5385 ( .IN1(n3140), .IN2(g965), .Q(n4885) );
  OR2X1 U5386 ( .IN1(g10724), .IN2(n3141), .Q(g10463) );
  OR2X1 U5387 ( .IN1(n4887), .IN2(n4888), .Q(g10724) );
  OR2X1 U5388 ( .IN1(n4889), .IN2(n4890), .Q(n4888) );
  OR2X1 U5389 ( .IN1(n4891), .IN2(n4892), .Q(n4890) );
  OR2X1 U5390 ( .IN1(n4893), .IN2(n4894), .Q(n4892) );
  AND2X1 U5391 ( .IN1(n1486), .IN2(g1537), .Q(n4894) );
  AND2X1 U5392 ( .IN1(n1485), .IN2(g1580), .Q(n4893) );
  OR2X1 U5393 ( .IN1(n4895), .IN2(n4896), .Q(n4891) );
  INVX0 U5394 ( .INP(n4897), .ZN(n4896) );
  AND2X1 U5395 ( .IN1(n4854), .IN2(n3025), .Q(n4895) );
  OR2X1 U5396 ( .IN1(n4898), .IN2(n4899), .Q(n4889) );
  OR2X1 U5397 ( .IN1(n4900), .IN2(n4901), .Q(n4899) );
  AND2X1 U5398 ( .IN1(n1479), .IN2(g1561), .Q(n4901) );
  AND2X1 U5399 ( .IN1(n1480), .IN2(g1604), .Q(n4900) );
  OR2X1 U5400 ( .IN1(n4902), .IN2(n4903), .Q(n4898) );
  AND2X1 U5401 ( .IN1(n4680), .IN2(n3034), .Q(n4903) );
  AND2X1 U5402 ( .IN1(n4831), .IN2(g1756), .Q(n4902) );
  OR2X1 U5403 ( .IN1(n4904), .IN2(n4905), .Q(n4887) );
  OR2X1 U5404 ( .IN1(n4906), .IN2(n4907), .Q(n4905) );
  OR2X1 U5405 ( .IN1(n4908), .IN2(n4909), .Q(n4907) );
  AND2X1 U5406 ( .IN1(n4786), .IN2(g1733), .Q(n4909) );
  AND2X1 U5407 ( .IN1(g1182), .IN2(n4775), .Q(n4908) );
  OR2X1 U5408 ( .IN1(n4910), .IN2(n4911), .Q(n4906) );
  AND2X1 U5409 ( .IN1(n4836), .IN2(g1327), .Q(n4911) );
  AND2X1 U5410 ( .IN1(g910), .IN2(n4801), .Q(n4910) );
  OR2X1 U5411 ( .IN1(n4912), .IN2(n4913), .Q(n4904) );
  OR2X1 U5412 ( .IN1(n4914), .IN2(n4915), .Q(n4913) );
  AND2X1 U5413 ( .IN1(n4847), .IN2(g299), .Q(n4915) );
  AND2X1 U5414 ( .IN1(n4802), .IN2(g275), .Q(n4914) );
  OR2X1 U5415 ( .IN1(n4916), .IN2(n4917), .Q(n4912) );
  AND2X1 U5416 ( .IN1(n4856), .IN2(n3057), .Q(n4917) );
  AND2X1 U5417 ( .IN1(n3140), .IN2(g962), .Q(n4916) );
  OR2X1 U5418 ( .IN1(g10721), .IN2(n3141), .Q(g10459) );
  OR2X1 U5419 ( .IN1(n4918), .IN2(n4919), .Q(g10721) );
  OR2X1 U5420 ( .IN1(n4920), .IN2(n4921), .Q(n4919) );
  OR2X1 U5421 ( .IN1(n4922), .IN2(n4923), .Q(n4921) );
  OR2X1 U5422 ( .IN1(n4924), .IN2(n4925), .Q(n4923) );
  AND2X1 U5423 ( .IN1(n1486), .IN2(g1531), .Q(n4925) );
  AND2X1 U5424 ( .IN1(n1485), .IN2(g1574), .Q(n4924) );
  OR2X1 U5425 ( .IN1(n4926), .IN2(n4927), .Q(n4922) );
  OR2X1 U5426 ( .IN1(n4928), .IN2(n4929), .Q(n4927) );
  AND2X1 U5427 ( .IN1(g1200), .IN2(n1512), .Q(n4929) );
  AND2X1 U5428 ( .IN1(n1480), .IN2(g1598), .Q(n4928) );
  AND2X1 U5429 ( .IN1(n1479), .IN2(g1555), .Q(n4926) );
  OR2X1 U5430 ( .IN1(n4930), .IN2(n4931), .Q(n4920) );
  OR2X1 U5431 ( .IN1(n4932), .IN2(n4933), .Q(n4931) );
  AND2X1 U5432 ( .IN1(n4680), .IN2(n3045), .Q(n4933) );
  AND2X1 U5433 ( .IN1(n4831), .IN2(g1750), .Q(n4932) );
  OR2X1 U5434 ( .IN1(n4934), .IN2(n4935), .Q(n4930) );
  OR2X1 U5435 ( .IN1(n4936), .IN2(n4937), .Q(n4935) );
  AND2X1 U5436 ( .IN1(g1176), .IN2(n4775), .Q(n4937) );
  AND2X1 U5437 ( .IN1(n4836), .IN2(g1321), .Q(n4936) );
  AND2X1 U5438 ( .IN1(n4786), .IN2(g1727), .Q(n4934) );
  OR2X1 U5439 ( .IN1(n4938), .IN2(n4939), .Q(n4918) );
  OR2X1 U5440 ( .IN1(n4940), .IN2(n4941), .Q(n4939) );
  OR2X1 U5441 ( .IN1(n4942), .IN2(n4943), .Q(n4941) );
  AND2X1 U5442 ( .IN1(n4782), .IN2(g1346), .Q(n4943) );
  AND2X1 U5443 ( .IN1(n4803), .IN2(g981), .Q(n4942) );
  OR2X1 U5444 ( .IN1(n4944), .IN2(n4945), .Q(n4940) );
  OR2X1 U5445 ( .IN1(n4946), .IN2(n4947), .Q(n4945) );
  AND2X1 U5446 ( .IN1(n4847), .IN2(g293), .Q(n4947) );
  AND2X1 U5447 ( .IN1(n4802), .IN2(g269), .Q(n4946) );
  AND2X1 U5448 ( .IN1(g904), .IN2(n4801), .Q(n4944) );
  OR2X1 U5449 ( .IN1(n4948), .IN2(n4949), .Q(n4938) );
  OR2X1 U5450 ( .IN1(n4950), .IN2(n4951), .Q(n4949) );
  OR2X1 U5451 ( .IN1(n4952), .IN2(n4953), .Q(n4951) );
  AND2X1 U5452 ( .IN1(n4854), .IN2(g1), .Q(n4953) );
  AND2X1 U5453 ( .IN1(g892), .IN2(n4855), .Q(n4952) );
  AND2X1 U5454 ( .IN1(n4856), .IN2(g9), .Q(n4950) );
  OR2X1 U5455 ( .IN1(n4954), .IN2(n4955), .Q(n4948) );
  OR2X1 U5456 ( .IN1(n4859), .IN2(n4956), .Q(n4955) );
  AND2X1 U5457 ( .IN1(n4861), .IN2(g936), .Q(n4956) );
  AND2X1 U5458 ( .IN1(n3140), .IN2(g956), .Q(n4954) );
  OR2X1 U5459 ( .IN1(g10720), .IN2(n3141), .Q(g10457) );
  OR2X1 U5460 ( .IN1(n4957), .IN2(n4958), .Q(g10720) );
  OR2X1 U5461 ( .IN1(n4959), .IN2(n4960), .Q(n4958) );
  OR2X1 U5462 ( .IN1(n4961), .IN2(n4962), .Q(n4960) );
  OR2X1 U5463 ( .IN1(n4963), .IN2(n4964), .Q(n4962) );
  AND2X1 U5464 ( .IN1(n1486), .IN2(g1528), .Q(n4964) );
  AND2X1 U5465 ( .IN1(n1485), .IN2(g1571), .Q(n4963) );
  OR2X1 U5466 ( .IN1(n4965), .IN2(n4966), .Q(n4961) );
  OR2X1 U5467 ( .IN1(n4967), .IN2(n4968), .Q(n4966) );
  AND2X1 U5468 ( .IN1(n1530), .IN2(g925), .Q(n4968) );
  AND2X1 U5469 ( .IN1(n1512), .IN2(g1197), .Q(n4967) );
  AND2X1 U5470 ( .IN1(n1479), .IN2(g1552), .Q(n4965) );
  OR2X1 U5471 ( .IN1(n4969), .IN2(n4970), .Q(n4959) );
  OR2X1 U5472 ( .IN1(n4971), .IN2(n4972), .Q(n4970) );
  OR2X1 U5473 ( .IN1(n4973), .IN2(n4974), .Q(n4972) );
  AND2X1 U5474 ( .IN1(n4680), .IN2(n3031), .Q(n4974) );
  AND2X1 U5475 ( .IN1(n4831), .IN2(g1747), .Q(n4973) );
  AND2X1 U5476 ( .IN1(n1480), .IN2(g1595), .Q(n4971) );
  OR2X1 U5477 ( .IN1(n4975), .IN2(n4976), .Q(n4969) );
  OR2X1 U5478 ( .IN1(n4977), .IN2(n4978), .Q(n4976) );
  AND2X1 U5479 ( .IN1(g1173), .IN2(n4775), .Q(n4978) );
  AND2X1 U5480 ( .IN1(n4836), .IN2(g1318), .Q(n4977) );
  AND2X1 U5481 ( .IN1(n4786), .IN2(g1724), .Q(n4975) );
  OR2X1 U5482 ( .IN1(n4979), .IN2(n4980), .Q(n4957) );
  OR2X1 U5483 ( .IN1(n4981), .IN2(n4982), .Q(n4980) );
  OR2X1 U5484 ( .IN1(n4983), .IN2(n4984), .Q(n4982) );
  AND2X1 U5485 ( .IN1(n4782), .IN2(g1341), .Q(n4984) );
  AND2X1 U5486 ( .IN1(n4803), .IN2(g976), .Q(n4983) );
  OR2X1 U5487 ( .IN1(n4985), .IN2(n4986), .Q(n4981) );
  OR2X1 U5488 ( .IN1(n4987), .IN2(n4988), .Q(n4986) );
  AND2X1 U5489 ( .IN1(n4847), .IN2(g290), .Q(n4988) );
  AND2X1 U5490 ( .IN1(n4802), .IN2(g266), .Q(n4987) );
  AND2X1 U5491 ( .IN1(g901), .IN2(n4801), .Q(n4985) );
  OR2X1 U5492 ( .IN1(n4989), .IN2(n4990), .Q(n4979) );
  OR2X1 U5493 ( .IN1(n4991), .IN2(n4992), .Q(n4990) );
  OR2X1 U5494 ( .IN1(n4993), .IN2(n4994), .Q(n4992) );
  AND2X1 U5495 ( .IN1(n4854), .IN2(g4), .Q(n4994) );
  AND2X1 U5496 ( .IN1(g889), .IN2(n4855), .Q(n4993) );
  AND2X1 U5497 ( .IN1(n4856), .IN2(g12), .Q(n4991) );
  OR2X1 U5498 ( .IN1(n4995), .IN2(n4996), .Q(n4989) );
  OR2X1 U5499 ( .IN1(n4859), .IN2(n4997), .Q(n4996) );
  AND2X1 U5500 ( .IN1(n4861), .IN2(g932), .Q(n4997) );
  AND2X1 U5501 ( .IN1(n3140), .IN2(g953), .Q(n4995) );
  OR2X1 U5502 ( .IN1(g10719), .IN2(n3141), .Q(g10455) );
  OR2X1 U5503 ( .IN1(n4998), .IN2(n4999), .Q(g10719) );
  OR2X1 U5504 ( .IN1(n5000), .IN2(n5001), .Q(n4999) );
  OR2X1 U5505 ( .IN1(n5002), .IN2(n5003), .Q(n5001) );
  OR2X1 U5506 ( .IN1(n5004), .IN2(n5005), .Q(n5003) );
  AND2X1 U5507 ( .IN1(n1486), .IN2(g1524), .Q(n5005) );
  AND2X1 U5508 ( .IN1(n1485), .IN2(g1567), .Q(n5004) );
  OR2X1 U5509 ( .IN1(n5006), .IN2(n5007), .Q(n5002) );
  OR2X1 U5510 ( .IN1(n5008), .IN2(n5009), .Q(n5007) );
  AND2X1 U5511 ( .IN1(g922), .IN2(n1530), .Q(n5009) );
  AND2X1 U5512 ( .IN1(g1194), .IN2(n1512), .Q(n5008) );
  AND2X1 U5513 ( .IN1(n1479), .IN2(g1549), .Q(n5006) );
  OR2X1 U5514 ( .IN1(n5010), .IN2(n5011), .Q(n5000) );
  OR2X1 U5515 ( .IN1(n5012), .IN2(n5013), .Q(n5011) );
  OR2X1 U5516 ( .IN1(n5014), .IN2(n5015), .Q(n5013) );
  AND2X1 U5517 ( .IN1(n4680), .IN2(n3051), .Q(n5015) );
  AND2X1 U5518 ( .IN1(n4831), .IN2(g1744), .Q(n5014) );
  AND2X1 U5519 ( .IN1(n1480), .IN2(g1592), .Q(n5012) );
  OR2X1 U5520 ( .IN1(n5016), .IN2(n5017), .Q(n5010) );
  OR2X1 U5521 ( .IN1(n5018), .IN2(n5019), .Q(n5017) );
  AND2X1 U5522 ( .IN1(g1170), .IN2(n4775), .Q(n5019) );
  AND2X1 U5523 ( .IN1(n4836), .IN2(g1314), .Q(n5018) );
  AND2X1 U5524 ( .IN1(n4786), .IN2(g1721), .Q(n5016) );
  OR2X1 U5525 ( .IN1(n5020), .IN2(n5021), .Q(n4998) );
  OR2X1 U5526 ( .IN1(n5022), .IN2(n5023), .Q(n5021) );
  OR2X1 U5527 ( .IN1(n5024), .IN2(n5025), .Q(n5023) );
  OR2X1 U5528 ( .IN1(n5026), .IN2(n5027), .Q(n5025) );
  AND2X1 U5529 ( .IN1(n4803), .IN2(g971), .Q(n5027) );
  AND2X1 U5530 ( .IN1(g898), .IN2(n4801), .Q(n5026) );
  INVX0 U5531 ( .INP(n5028), .ZN(n5024) );
  OR2X1 U5532 ( .IN1(n5029), .IN2(n2821), .Q(n5028) );
  OR2X1 U5533 ( .IN1(n5030), .IN2(n5031), .Q(n5022) );
  OR2X1 U5534 ( .IN1(n5032), .IN2(n5033), .Q(n5031) );
  AND2X1 U5535 ( .IN1(n4802), .IN2(g263), .Q(n5033) );
  AND2X1 U5536 ( .IN1(n4856), .IN2(g119), .Q(n5032) );
  AND2X1 U5537 ( .IN1(n4847), .IN2(g287), .Q(n5030) );
  INVX0 U5538 ( .INP(n5034), .ZN(n4847) );
  OR2X1 U5539 ( .IN1(n5035), .IN2(n5036), .Q(n5020) );
  OR2X1 U5540 ( .IN1(n5037), .IN2(n5038), .Q(n5036) );
  OR2X1 U5541 ( .IN1(n5039), .IN2(n5040), .Q(n5038) );
  AND2X1 U5542 ( .IN1(g886), .IN2(n4855), .Q(n5040) );
  AND2X1 U5543 ( .IN1(n3140), .IN2(g950), .Q(n5039) );
  AND2X1 U5544 ( .IN1(n4854), .IN2(g123), .Q(n5037) );
  OR2X1 U5545 ( .IN1(n5041), .IN2(n5042), .Q(n5035) );
  OR2X1 U5546 ( .IN1(n525), .IN2(n4859), .Q(n5042) );
  INVX0 U5547 ( .INP(n5043), .ZN(n4859) );
  OR2X1 U5548 ( .IN1(n5044), .IN2(n4897), .Q(n5043) );
  OR2X1 U5549 ( .IN1(n5045), .IN2(n4854), .Q(n4897) );
  AND2X1 U5550 ( .IN1(g42), .IN2(n5046), .Q(n4854) );
  OR2X1 U5551 ( .IN1(n5047), .IN2(n5048), .Q(n5045) );
  OR2X1 U5552 ( .IN1(n5049), .IN2(n3142), .Q(n5048) );
  OR2X1 U5553 ( .IN1(n5050), .IN2(n5051), .Q(n3142) );
  OR2X1 U5554 ( .IN1(n5052), .IN2(n5053), .Q(n5051) );
  OR2X1 U5555 ( .IN1(n5054), .IN2(n4680), .Q(n5053) );
  OR2X1 U5556 ( .IN1(n3140), .IN2(n4861), .Q(n5052) );
  AND2X1 U5557 ( .IN1(n535), .IN2(n5055), .Q(n3140) );
  OR2X1 U5558 ( .IN1(n5056), .IN2(n5057), .Q(n5050) );
  OR2X1 U5559 ( .IN1(n4801), .IN2(n4855), .Q(n5057) );
  INVX0 U5560 ( .INP(n5058), .ZN(n4855) );
  OR2X1 U5561 ( .IN1(n5059), .IN2(n5060), .Q(n5058) );
  OR2X1 U5562 ( .IN1(n5061), .IN2(n5062), .Q(n5060) );
  OR2X1 U5563 ( .IN1(n5063), .IN2(n4637), .Q(n5059) );
  OR2X1 U5564 ( .IN1(n1530), .IN2(n4803), .Q(n5056) );
  OR2X1 U5565 ( .IN1(n525), .IN2(n4856), .Q(n5047) );
  AND2X1 U5566 ( .IN1(n4637), .IN2(n5046), .Q(n4856) );
  INVX0 U5567 ( .INP(n5064), .ZN(n5046) );
  OR2X1 U5568 ( .IN1(n5065), .IN2(n5066), .Q(n5064) );
  OR2X1 U5569 ( .IN1(n5063), .IN2(n4788), .Q(n5066) );
  INVX0 U5570 ( .INP(g43), .ZN(n5063) );
  OR2X1 U5571 ( .IN1(g45), .IN2(g44), .Q(n5065) );
  OR2X1 U5572 ( .IN1(n1512), .IN2(n4782), .Q(n5044) );
  AND2X1 U5573 ( .IN1(n4861), .IN2(g928), .Q(n5041) );
  INVX0 U5574 ( .INP(n5067), .ZN(n4861) );
  OR2X1 U5575 ( .IN1(n5068), .IN2(n5069), .Q(n5067) );
  OR2X1 U5576 ( .IN1(n5061), .IN2(n5070), .Q(n5069) );
  OR2X1 U5577 ( .IN1(n4637), .IN2(n5071), .Q(n5068) );
  OR2X1 U5578 ( .IN1(g43), .IN2(n5072), .Q(n5071) );
  OR2X1 U5579 ( .IN1(g10663), .IN2(n3141), .Q(g10377) );
  OR2X1 U5580 ( .IN1(g30), .IN2(n4680), .Q(n3141) );
  OR2X1 U5581 ( .IN1(n5073), .IN2(n5074), .Q(g10663) );
  OR2X1 U5582 ( .IN1(n5075), .IN2(n5076), .Q(n5074) );
  OR2X1 U5583 ( .IN1(n5077), .IN2(n5078), .Q(n5076) );
  OR2X1 U5584 ( .IN1(n5079), .IN2(n5080), .Q(n5078) );
  AND2X1 U5585 ( .IN1(n1486), .IN2(g1543), .Q(n5080) );
  AND2X1 U5586 ( .IN1(n1485), .IN2(g1586), .Q(n5079) );
  OR2X1 U5587 ( .IN1(n5081), .IN2(n5082), .Q(n5077) );
  AND2X1 U5588 ( .IN1(n4879), .IN2(n5029), .Q(n5082) );
  INVX0 U5589 ( .INP(n4782), .ZN(n5029) );
  AND2X1 U5590 ( .IN1(n1478), .IN2(n5083), .Q(n4879) );
  INVX0 U5591 ( .INP(n5049), .ZN(n5083) );
  OR2X1 U5592 ( .IN1(n5084), .IN2(n5085), .Q(n5049) );
  OR2X1 U5593 ( .IN1(n4786), .IN2(n5086), .Q(n5085) );
  OR2X1 U5594 ( .IN1(n4836), .IN2(n4831), .Q(n5086) );
  OR2X1 U5595 ( .IN1(n4775), .IN2(n5087), .Q(n5084) );
  OR2X1 U5596 ( .IN1(n1567), .IN2(n1566), .Q(n5087) );
  OR2X1 U5597 ( .IN1(n5088), .IN2(n1479), .Q(n1566) );
  AND2X1 U5598 ( .IN1(n5089), .IN2(n530), .Q(n5088) );
  OR2X1 U5599 ( .IN1(n5090), .IN2(n1480), .Q(n1567) );
  AND2X1 U5600 ( .IN1(n530), .IN2(n5055), .Q(n1480) );
  AND2X1 U5601 ( .IN1(n5091), .IN2(n530), .Q(n5090) );
  INVX0 U5602 ( .INP(n4788), .ZN(n530) );
  AND2X1 U5603 ( .IN1(n4782), .IN2(g1308), .Q(n5081) );
  AND2X1 U5604 ( .IN1(n5091), .IN2(n529), .Q(n4782) );
  OR2X1 U5605 ( .IN1(n5092), .IN2(n5093), .Q(n5075) );
  OR2X1 U5606 ( .IN1(n5094), .IN2(n5095), .Q(n5093) );
  AND2X1 U5607 ( .IN1(n4831), .IN2(g1762), .Q(n5095) );
  AND2X1 U5608 ( .IN1(n4637), .IN2(n5096), .Q(n4831) );
  AND2X1 U5609 ( .IN1(n4786), .IN2(g1738), .Q(n5094) );
  AND2X1 U5610 ( .IN1(g42), .IN2(n5096), .Q(n4786) );
  AND2X1 U5611 ( .IN1(n529), .IN2(n5097), .Q(n5096) );
  AND2X1 U5612 ( .IN1(n5098), .IN2(g45), .Q(n5097) );
  AND2X1 U5613 ( .IN1(n4680), .IN2(n1637), .Q(n5092) );
  OR2X1 U5614 ( .IN1(n5099), .IN2(n5100), .Q(n5073) );
  OR2X1 U5615 ( .IN1(n5101), .IN2(n5102), .Q(n5100) );
  OR2X1 U5616 ( .IN1(n5103), .IN2(n5104), .Q(n5102) );
  AND2X1 U5617 ( .IN1(n4836), .IN2(g1333), .Q(n5104) );
  AND2X1 U5618 ( .IN1(n529), .IN2(n5055), .Q(n4836) );
  INVX0 U5619 ( .INP(n5105), .ZN(n5055) );
  OR2X1 U5620 ( .IN1(n5062), .IN2(n5106), .Q(n5105) );
  OR2X1 U5621 ( .IN1(g43), .IN2(g42), .Q(n5106) );
  AND2X1 U5622 ( .IN1(n4803), .IN2(g944), .Q(n5103) );
  AND2X1 U5623 ( .IN1(n535), .IN2(n5091), .Q(n4803) );
  INVX0 U5624 ( .INP(n4790), .ZN(n5091) );
  OR2X1 U5625 ( .IN1(n5062), .IN2(n5107), .Q(n4790) );
  OR2X1 U5626 ( .IN1(g43), .IN2(n4637), .Q(n5107) );
  OR2X1 U5627 ( .IN1(g44), .IN2(n5070), .Q(n5062) );
  INVX0 U5628 ( .INP(g45), .ZN(n5070) );
  AND2X1 U5629 ( .IN1(g1188), .IN2(n4775), .Q(n5101) );
  AND2X1 U5630 ( .IN1(n5089), .IN2(n529), .Q(n4775) );
  INVX0 U5631 ( .INP(n5108), .ZN(n529) );
  OR2X1 U5632 ( .IN1(n5109), .IN2(n3156), .Q(n5108) );
  OR2X1 U5633 ( .IN1(n5110), .IN2(n5111), .Q(n3156) );
  OR2X1 U5634 ( .IN1(g46), .IN2(n3180), .Q(n5111) );
  OR2X1 U5635 ( .IN1(n5112), .IN2(n5113), .Q(n5099) );
  OR2X1 U5636 ( .IN1(n5114), .IN2(n5115), .Q(n5113) );
  AND2X1 U5637 ( .IN1(g916), .IN2(n4801), .Q(n5115) );
  AND2X1 U5638 ( .IN1(n535), .IN2(n5089), .Q(n4801) );
  INVX0 U5639 ( .INP(n4789), .ZN(n5089) );
  OR2X1 U5640 ( .IN1(n4637), .IN2(n5116), .Q(n4789) );
  OR2X1 U5641 ( .IN1(g45), .IN2(n5117), .Q(n5116) );
  INVX0 U5642 ( .INP(g42), .ZN(n4637) );
  INVX0 U5643 ( .INP(n5061), .ZN(n535) );
  OR2X1 U5644 ( .IN1(n5109), .IN2(n3154), .Q(n5061) );
  OR2X1 U5645 ( .IN1(n5118), .IN2(n4636), .Q(n3154) );
  AND2X1 U5646 ( .IN1(n4802), .IN2(g281), .Q(n5114) );
  AND2X1 U5647 ( .IN1(n5034), .IN2(n5054), .Q(n4802) );
  INVX0 U5648 ( .INP(n5119), .ZN(n5054) );
  OR2X1 U5649 ( .IN1(g42), .IN2(n5119), .Q(n5034) );
  OR2X1 U5650 ( .IN1(n5120), .IN2(n5121), .Q(n5119) );
  OR2X1 U5651 ( .IN1(n5072), .IN2(n4788), .Q(n5121) );
  OR2X1 U5652 ( .IN1(n4636), .IN2(n5122), .Q(n4788) );
  OR2X1 U5653 ( .IN1(g46), .IN2(n5109), .Q(n5122) );
  OR2X1 U5654 ( .IN1(n3180), .IN2(g47), .Q(n4636) );
  INVX0 U5655 ( .INP(g44), .ZN(n5072) );
  OR2X1 U5656 ( .IN1(g45), .IN2(g43), .Q(n5120) );
  OR2X1 U5657 ( .IN1(n1564), .IN2(n525), .Q(n5112) );
  INVX0 U5658 ( .INP(n5123), .ZN(n525) );
  OR2X1 U5659 ( .IN1(n5124), .IN2(n5125), .Q(n5123) );
  OR2X1 U5660 ( .IN1(n5118), .IN2(n5110), .Q(n5125) );
  INVX0 U5661 ( .INP(g47), .ZN(n5110) );
  INVX0 U5662 ( .INP(g46), .ZN(n5118) );
  OR2X1 U5663 ( .IN1(n5109), .IN2(n5126), .Q(n5124) );
  OR2X1 U5664 ( .IN1(n1545), .IN2(n3180), .Q(n5126) );
  AND2X1 U5665 ( .IN1(n5127), .IN2(n5128), .Q(n3180) );
  OR2X1 U5666 ( .IN1(n4680), .IN2(n5109), .Q(n5128) );
  OR2X1 U5667 ( .IN1(g31), .IN2(n5129), .Q(n4680) );
  OR2X1 U5668 ( .IN1(n5130), .IN2(g30), .Q(n5127) );
  OR2X1 U5669 ( .IN1(g41), .IN2(g48), .Q(n5130) );
  OR2X1 U5670 ( .IN1(n5117), .IN2(n5131), .Q(n1545) );
  OR2X1 U5671 ( .IN1(g45), .IN2(g42), .Q(n5131) );
  INVX0 U5672 ( .INP(n5098), .ZN(n5117) );
  AND2X1 U5673 ( .IN1(g43), .IN2(g44), .Q(n5098) );
  OR2X1 U5674 ( .IN1(g41), .IN2(n5129), .Q(n5109) );
  INVX0 U5675 ( .INP(g48), .ZN(n5129) );
  XNOR2X1 U5676 ( .IN1(test_so1), .IN2(n3629), .Q(N599) );
  OR2X1 U5677 ( .IN1(n3632), .IN2(n5132), .Q(n3629) );
  OR2X1 U5678 ( .IN1(n2883), .IN2(n2865), .Q(n5132) );
  INVX0 U5679 ( .INP(n1093), .ZN(n3632) );
  OR2X1 U1550_U1 ( .IN1(g10722), .IN2(n524), .Q(g10461) );
  OR2X1 U1551_U1 ( .IN1(g10664), .IN2(n524), .Q(g10379) );
  INVX0 U1586_U2 ( .INP(n2897), .ZN(U1586_n1) );
  AND2X1 U1586_U1 ( .IN1(n13), .IN2(U1586_n1), .Q(n1855) );
  INVX0 U1754_U2 ( .INP(n1545), .ZN(U1754_n1) );
  AND2X1 U1754_U1 ( .IN1(n530), .IN2(U1754_n1), .Q(n1479) );
  INVX0 U1798_U2 ( .INP(n1480), .ZN(U1798_n1) );
  AND2X1 U1798_U1 ( .IN1(n1567), .IN2(U1798_n1), .Q(n1485) );
  INVX0 U1839_U2 ( .INP(n1479), .ZN(U1839_n1) );
  AND2X1 U1839_U1 ( .IN1(n1566), .IN2(U1839_n1), .Q(n1486) );
  INVX0 U1843_U2 ( .INP(n525), .ZN(U1843_n1) );
  AND2X1 U1843_U1 ( .IN1(n499), .IN2(U1843_n1), .Q(n1478) );
  INVX0 U1877_U2 ( .INP(n519), .ZN(U1877_n1) );
  AND2X1 U1877_U1 ( .IN1(n1137), .IN2(U1877_n1), .Q(n1195) );
  INVX0 U1908_U2 ( .INP(n1545), .ZN(U1908_n1) );
  AND2X1 U1908_U1 ( .IN1(n529), .IN2(U1908_n1), .Q(n1512) );
  INVX0 U1909_U2 ( .INP(n1545), .ZN(U1909_n1) );
  AND2X1 U1909_U1 ( .IN1(n535), .IN2(U1909_n1), .Q(n1530) );
  INVX0 U1987_U2 ( .INP(n252), .ZN(U1987_n1) );
  AND2X1 U1987_U1 ( .IN1(n822), .IN2(U1987_n1), .Q(n916) );
  INVX0 U2031_U2 ( .INP(n369), .ZN(U2031_n1) );
  AND2X1 U2031_U1 ( .IN1(n104), .IN2(U2031_n1), .Q(n1056) );
  INVX0 U2035_U2 ( .INP(g109), .ZN(U2035_n1) );
  AND2X1 U2035_U1 ( .IN1(n1404), .IN2(U2035_n1), .Q(n1450) );
  INVX0 U2418_U2 ( .INP(n534), .ZN(U2418_n1) );
  AND2X1 U2418_U1 ( .IN1(g968), .IN2(U2418_n1), .Q(n1564) );
  INVX0 U2468_U2 ( .INP(n1227), .ZN(U2468_n1) );
  AND2X1 U2468_U1 ( .IN1(g1336), .IN2(U2468_n1), .Q(n1231) );
  INVX0 U2478_U2 ( .INP(n225), .ZN(U2478_n1) );
  AND2X1 U2478_U1 ( .IN1(g1341), .IN2(U2478_n1), .Q(n1232) );
  INVX0 U2488_U2 ( .INP(n1258), .ZN(U2488_n1) );
  AND2X1 U2488_U1 ( .IN1(n1262), .IN2(U2488_n1), .Q(n1260) );
  INVX0 U2533_U2 ( .INP(n519), .ZN(U2533_n1) );
  AND2X1 U2533_U1 ( .IN1(g178), .IN2(U2533_n1), .Q(g6786) );
  INVX0 U2534_U2 ( .INP(n519), .ZN(U2534_n1) );
  AND2X1 U2534_U1 ( .IN1(g1424), .IN2(U2534_n1), .Q(g6234) );
  INVX0 U2639_U2 ( .INP(n958), .ZN(U2639_n1) );
  AND2X1 U2639_U1 ( .IN1(n962), .IN2(U2639_n1), .Q(n804) );
  INVX0 U2641_U2 ( .INP(g1868), .ZN(U2641_n1) );
  AND2X1 U2641_U1 ( .IN1(n1147), .IN2(U2641_n1), .Q(n926) );
  INVX0 U2654_U2 ( .INP(g750), .ZN(U2654_n1) );
  AND2X1 U2654_U1 ( .IN1(g746), .IN2(U2654_n1), .Q(g4171) );
  INVX0 U2658_U2 ( .INP(n918), .ZN(U2658_n1) );
  AND2X1 U2658_U1 ( .IN1(n9), .IN2(U2658_n1), .Q(n812) );
  INVX0 U2683_U2 ( .INP(n1385), .ZN(U2683_n1) );
  AND2X1 U2683_U1 ( .IN1(g382), .IN2(U2683_n1), .Q(n1420) );
  INVX0 U2699_U2 ( .INP(n503), .ZN(U2699_n1) );
  AND2X1 U2699_U1 ( .IN1(n808), .IN2(U2699_n1), .Q(n806) );
  INVX0 U2846_U2 ( .INP(n1214), .ZN(U2846_n1) );
  AND2X1 U2846_U1 ( .IN1(g4175), .IN2(U2846_n1), .Q(n1193) );
  INVX0 U2847_U2 ( .INP(n1153), .ZN(U2847_n1) );
  AND2X1 U2847_U1 ( .IN1(g4177), .IN2(U2847_n1), .Q(n1125) );
  INVX0 U2848_U2 ( .INP(n1099), .ZN(U2848_n1) );
  AND2X1 U2848_U1 ( .IN1(g4179), .IN2(U2848_n1), .Q(n1093) );
  INVX0 U2859_U2 ( .INP(g12), .ZN(U2859_n1) );
  AND2X1 U2859_U1 ( .IN1(n1137), .IN2(U2859_n1), .Q(n1159) );
  INVX0 U2860_U2 ( .INP(n1151), .ZN(U2860_n1) );
  AND2X1 U2860_U1 ( .IN1(g810), .IN2(U2860_n1), .Q(n1123) );
  INVX0 U2861_U2 ( .INP(n1097), .ZN(U2861_n1) );
  AND2X1 U2861_U1 ( .IN1(g818), .IN2(U2861_n1), .Q(n1090) );
  INVX0 U2867_U2 ( .INP(g1834), .ZN(U2867_n1) );
  AND2X1 U2867_U1 ( .IN1(n817), .IN2(U2867_n1), .Q(n1380) );
  INVX0 U2879_U2 ( .INP(n1656), .ZN(U2879_n1) );
  AND2X1 U2879_U1 ( .IN1(g713), .IN2(U2879_n1), .Q(n967) );
  INVX0 U2881_U2 ( .INP(n1657), .ZN(U2881_n1) );
  AND2X1 U2881_U1 ( .IN1(g1927), .IN2(U2881_n1), .Q(n921) );
  INVX0 U2882_U2 ( .INP(n519), .ZN(U2882_n1) );
  AND2X1 U2882_U1 ( .IN1(g1160), .IN2(U2882_n1), .Q(g4334) );
  INVX0 U2883_U2 ( .INP(n519), .ZN(U2883_n1) );
  AND2X1 U2883_U1 ( .IN1(g1166), .IN2(U2883_n1), .Q(g4325) );
  INVX0 U2884_U2 ( .INP(n519), .ZN(U2884_n1) );
  AND2X1 U2884_U1 ( .IN1(g148), .IN2(U2884_n1), .Q(g6759) );
  INVX0 U2885_U2 ( .INP(n519), .ZN(U2885_n1) );
  AND2X1 U2885_U1 ( .IN1(g1157), .IN2(U2885_n1), .Q(g4338) );
  INVX0 U2886_U2 ( .INP(n519), .ZN(U2886_n1) );
  AND2X1 U2886_U1 ( .IN1(g1163), .IN2(U2886_n1), .Q(g4330) );
  INVX0 U2887_U2 ( .INP(n519), .ZN(U2887_n1) );
  AND2X1 U2887_U1 ( .IN1(g237), .IN2(U2887_n1), .Q(g6821) );
  INVX0 U2888_U2 ( .INP(n519), .ZN(U2888_n1) );
  AND2X1 U2888_U1 ( .IN1(g1499), .IN2(U2888_n1), .Q(g6198) );
  INVX0 U2889_U2 ( .INP(n519), .ZN(U2889_n1) );
  AND2X1 U2889_U1 ( .IN1(g1411), .IN2(U2889_n1), .Q(g6244) );
  INVX0 U2890_U2 ( .INP(n519), .ZN(U2890_n1) );
  AND2X1 U2890_U1 ( .IN1(g225), .IN2(U2890_n1), .Q(g6826) );
  INVX0 U2891_U2 ( .INP(n519), .ZN(U2891_n1) );
  AND2X1 U2891_U1 ( .IN1(g1407), .IN2(U2891_n1), .Q(g6216) );
  INVX0 U2892_U2 ( .INP(n519), .ZN(U2892_n1) );
  AND2X1 U2892_U1 ( .IN1(g213), .IN2(U2892_n1), .Q(g6829) );
  INVX0 U2893_U2 ( .INP(n519), .ZN(U2893_n1) );
  AND2X1 U2893_U1 ( .IN1(g186), .IN2(U2893_n1), .Q(g6833) );
  INVX0 U2894_U2 ( .INP(n519), .ZN(U2894_n1) );
  AND2X1 U2894_U1 ( .IN1(g219), .IN2(U2894_n1), .Q(g6827) );
  INVX0 U2895_U2 ( .INP(n519), .ZN(U2895_n1) );
  AND2X1 U2895_U1 ( .IN1(g143), .IN2(U2895_n1), .Q(g6757) );
  INVX0 U2896_U2 ( .INP(n519), .ZN(U2896_n1) );
  AND2X1 U2896_U1 ( .IN1(g207), .IN2(U2896_n1), .Q(g6831) );
  INVX0 U2897_U2 ( .INP(n519), .ZN(U2897_n1) );
  AND2X1 U2897_U1 ( .IN1(g231), .IN2(U2897_n1), .Q(g6822) );
  INVX0 U2898_U2 ( .INP(n519), .ZN(U2898_n1) );
  AND2X1 U2898_U1 ( .IN1(g192), .IN2(U2898_n1), .Q(g6838) );
  INVX0 U2899_U2 ( .INP(n519), .ZN(U2899_n1) );
  AND2X1 U2899_U1 ( .IN1(test_so3), .IN2(U2899_n1), .Q(g6823) );
  INVX0 U2900_U2 ( .INP(n519), .ZN(U2900_n1) );
  AND2X1 U2900_U1 ( .IN1(g1371), .IN2(U2900_n1), .Q(g6824) );
  INVX0 U2901_U2 ( .INP(n519), .ZN(U2901_n1) );
  AND2X1 U2901_U1 ( .IN1(g1383), .IN2(U2901_n1), .Q(g6832) );
  INVX0 U2902_U2 ( .INP(n519), .ZN(U2902_n1) );
  AND2X1 U2902_U1 ( .IN1(g243), .IN2(U2902_n1), .Q(g6819) );
  INVX0 U3090_U2 ( .INP(g810), .ZN(U3090_n1) );
  AND2X1 U3090_U1 ( .IN1(n1151), .IN2(U3090_n1), .Q(n1150) );
  INVX0 U3092_U2 ( .INP(g818), .ZN(U3092_n1) );
  AND2X1 U3092_U1 ( .IN1(n1097), .IN2(U3092_n1), .Q(n1096) );
  INVX0 U3094_U2 ( .INP(g4179), .ZN(U3094_n1) );
  AND2X1 U3094_U1 ( .IN1(n1099), .IN2(U3094_n1), .Q(n1098) );
  INVX0 U3096_U2 ( .INP(g4175), .ZN(U3096_n1) );
  AND2X1 U3096_U1 ( .IN1(n1214), .IN2(U3096_n1), .Q(n1213) );
  INVX0 U3098_U2 ( .INP(g4177), .ZN(U3098_n1) );
  AND2X1 U3098_U1 ( .IN1(n1153), .IN2(U3098_n1), .Q(n1152) );
  INVX0 U3124_U2 ( .INP(n838), .ZN(U3124_n1) );
  AND2X1 U3124_U1 ( .IN1(n837), .IN2(U3124_n1), .Q(n836) );
  INVX0 U3171_U2 ( .INP(n2903), .ZN(U3171_n1) );
  AND2X1 U3171_U1 ( .IN1(g1610), .IN2(U3171_n1), .Q(g5194) );
endmodule

