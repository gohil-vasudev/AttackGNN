module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n318_, new_n155_, new_n384_, new_n163_, new_n410_, new_n445_, new_n236_, new_n238_, new_n148_, new_n321_, new_n440_, new_n443_, new_n324_, new_n122_, new_n250_, new_n288_, new_n371_, new_n252_, new_n421_, new_n202_, new_n262_, new_n296_, new_n160_, new_n308_, new_n271_, new_n274_, new_n372_, new_n242_, new_n368_, new_n232_, new_n218_, new_n258_, new_n307_, new_n190_, new_n439_, new_n176_, new_n305_, new_n420_, new_n156_, new_n223_, new_n283_, new_n306_, new_n291_, new_n366_, new_n261_, new_n390_, new_n241_, new_n309_, new_n408_, new_n186_, new_n339_, new_n213_, new_n134_, new_n197_, new_n205_, new_n323_, new_n365_, new_n386_, new_n259_, new_n362_, new_n389_, new_n401_, new_n433_, new_n435_, new_n206_, new_n429_, new_n227_, new_n355_, new_n353_, new_n222_, new_n416_, new_n432_, new_n265_, new_n246_, new_n170_, new_n370_, new_n400_, new_n256_, new_n328_, new_n266_, new_n367_, new_n278_, new_n304_, new_n381_, new_n173_, new_n220_, new_n388_, new_n268_, new_n217_, new_n269_, new_n374_, new_n376_, new_n194_, new_n380_, new_n214_, new_n394_, new_n299_, new_n138_, new_n424_, new_n142_, new_n310_, new_n275_, new_n188_, new_n139_, new_n240_, new_n413_, new_n314_, new_n352_, new_n442_, new_n363_, new_n412_, new_n165_, new_n123_, new_n127_, new_n211_, new_n342_, new_n441_, new_n327_, new_n216_, new_n177_, new_n431_, new_n196_, new_n280_, new_n264_, new_n426_, new_n319_, new_n235_, new_n379_, new_n273_, new_n398_, new_n224_, new_n301_, new_n169_, new_n270_, new_n338_, new_n395_, new_n383_, new_n317_, new_n210_, new_n343_, new_n143_, new_n344_, new_n447_, new_n207_, new_n267_, new_n145_, new_n287_, new_n253_, new_n140_, new_n336_, new_n247_, new_n377_, new_n403_, new_n237_, new_n330_, new_n375_, new_n234_, new_n427_, new_n294_, new_n187_, new_n260_, new_n311_, new_n393_, new_n418_, new_n251_, new_n189_, new_n300_, new_n292_, new_n195_, new_n263_, new_n411_, new_n215_, new_n331_, new_n334_, new_n152_, new_n341_, new_n378_, new_n157_, new_n182_, new_n407_, new_n153_, new_n357_, new_n320_, new_n349_, new_n244_, new_n172_, new_n133_, new_n277_, new_n257_, new_n245_, new_n402_, new_n212_, new_n151_, new_n286_, new_n404_, new_n335_, new_n347_, new_n364_, new_n449_, new_n193_, new_n219_, new_n231_, new_n313_, new_n239_, new_n382_, new_n272_, new_n282_, new_n396_, new_n198_, new_n201_, new_n428_, new_n438_, new_n128_, new_n192_, new_n199_, new_n146_, new_n358_, new_n208_, new_n348_, new_n360_, new_n414_, new_n159_, new_n322_, new_n228_, new_n315_, new_n302_, new_n191_, new_n326_, new_n289_, new_n179_, new_n225_, new_n164_, new_n425_, new_n230_, new_n175_, new_n226_, new_n281_, new_n397_, new_n430_, new_n436_, new_n185_, new_n387_, new_n399_, new_n373_, new_n171_, new_n248_, new_n350_, new_n121_, new_n415_, new_n221_, new_n243_, new_n385_, new_n200_, new_n345_, new_n434_, new_n298_, new_n422_, new_n184_, new_n154_, new_n255_, new_n329_, new_n249_, new_n233_, new_n284_, new_n293_, new_n178_, new_n168_, new_n174_, new_n297_, new_n279_, new_n361_, new_n150_, new_n295_, new_n359_, new_n354_, new_n392_, new_n444_, new_n166_, new_n137_, new_n162_, new_n183_, new_n409_, new_n303_, new_n161_, new_n340_, new_n285_, new_n406_, new_n423_, new_n356_, new_n333_, new_n229_, new_n209_, new_n337_, new_n351_, new_n290_, new_n203_, new_n316_, new_n204_, new_n446_, new_n325_, new_n181_, new_n369_, new_n417_, new_n180_, new_n448_, new_n276_;

and g000 ( N388, N29, N42, N75 );
and g001 ( N389, N29, N36, N80 );
not g002 ( new_n121_, N29 );
not g003 ( new_n122_, N36 );
not g004 ( new_n123_, N42 );
nor g005 ( N390, new_n121_, new_n122_, new_n123_ );
and g006 ( N391, N85, N86 );
and g007 ( N418, N1, N8, N13, N17 );
not g008 ( new_n127_, N390 );
and g009 ( new_n128_, N1, N13, N17, N26 );
nand g010 ( N419, new_n127_, new_n128_ );
nand g011 ( N420, N59, N75, N80 );
nand g012 ( N421, N36, N59, N80 );
nand g013 ( N422, N36, N42, N59 );
not g014 ( new_n133_, N90 );
nor g015 ( new_n134_, N87, N88 );
nor g016 ( N423, new_n134_, new_n133_ );
nand g017 ( N446, N390, new_n128_ );
not g018 ( new_n137_, keyIn_0_0 );
nand g019 ( new_n138_, new_n137_, N1, N26, N51 );
nand g020 ( new_n139_, N1, N26, N51 );
nand g021 ( new_n140_, new_n139_, keyIn_0_0 );
nand g022 ( N447, new_n140_, new_n138_ );
not g023 ( new_n142_, N68 );
nand g024 ( new_n143_, N1, N8, N13, N55 );
nor g025 ( N448, new_n143_, new_n121_, new_n142_ );
not g026 ( new_n145_, N74 );
nand g027 ( new_n146_, N59, N68 );
nor g028 ( N449, new_n143_, new_n145_, new_n146_ );
not g029 ( new_n148_, N89 );
nor g030 ( N450, new_n134_, new_n148_ );
xor g031 ( new_n150_, N111, N116 );
xnor g032 ( new_n151_, N121, N126 );
xnor g033 ( new_n152_, new_n150_, new_n151_ );
xnor g034 ( new_n153_, new_n152_, N135 );
xnor g035 ( new_n154_, N91, N96 );
xnor g036 ( new_n155_, N101, N106 );
xnor g037 ( new_n156_, new_n154_, new_n155_ );
xnor g038 ( new_n157_, new_n156_, N130 );
xnor g039 ( N767, new_n153_, new_n157_ );
xor g040 ( new_n159_, N183, N189 );
xnor g041 ( new_n160_, N195, N201 );
xnor g042 ( new_n161_, new_n159_, new_n160_ );
xnor g043 ( new_n162_, new_n161_, N207 );
xnor g044 ( new_n163_, N159, N165 );
xnor g045 ( new_n164_, N171, N177 );
xnor g046 ( new_n165_, new_n163_, new_n164_ );
xnor g047 ( new_n166_, new_n165_, N130 );
xnor g048 ( N768, new_n162_, new_n166_ );
not g049 ( new_n168_, keyIn_0_21 );
not g050 ( new_n169_, keyIn_0_17 );
not g051 ( new_n170_, keyIn_0_15 );
not g052 ( new_n171_, keyIn_0_10 );
not g053 ( new_n172_, keyIn_0_6 );
nand g054 ( new_n173_, N447, new_n172_ );
nand g055 ( new_n174_, new_n140_, keyIn_0_6, new_n138_ );
nand g056 ( new_n175_, new_n173_, new_n174_ );
nand g057 ( new_n176_, new_n175_, new_n171_ );
nand g058 ( new_n177_, new_n173_, keyIn_0_10, new_n174_ );
nand g059 ( new_n178_, new_n176_, new_n177_ );
not g060 ( new_n179_, N17 );
nand g061 ( new_n180_, new_n179_, new_n123_ );
nand g062 ( new_n181_, new_n180_, keyIn_0_4 );
or g063 ( new_n182_, keyIn_0_4, N17, N42 );
nand g064 ( new_n183_, new_n181_, new_n182_ );
nand g065 ( new_n184_, N17, N42 );
xnor g066 ( new_n185_, new_n184_, keyIn_0_5 );
nand g067 ( new_n186_, new_n183_, new_n185_, keyIn_0_9 );
nand g068 ( new_n187_, N59, N156 );
not g069 ( new_n188_, new_n187_ );
not g070 ( new_n189_, keyIn_0_9 );
nand g071 ( new_n190_, new_n183_, new_n185_ );
nand g072 ( new_n191_, new_n190_, new_n189_ );
and g073 ( new_n192_, new_n191_, new_n186_, new_n188_ );
nand g074 ( new_n193_, new_n192_, new_n170_, new_n178_ );
nand g075 ( new_n194_, new_n192_, new_n178_ );
nand g076 ( new_n195_, new_n194_, keyIn_0_15 );
nand g077 ( new_n196_, new_n195_, new_n193_ );
not g078 ( new_n197_, keyIn_0_11 );
nand g079 ( new_n198_, N42, N59, N75 );
xnor g080 ( new_n199_, new_n198_, keyIn_0_2 );
xnor g081 ( new_n200_, new_n199_, keyIn_0_8 );
and g082 ( new_n201_, N1, N8, N17, N51 );
xnor g083 ( new_n202_, new_n201_, keyIn_0_1 );
xnor g084 ( new_n203_, new_n202_, keyIn_0_7 );
nand g085 ( new_n204_, new_n203_, new_n200_ );
nand g086 ( new_n205_, new_n204_, new_n197_ );
nand g087 ( new_n206_, new_n203_, keyIn_0_11, new_n200_ );
nand g088 ( new_n207_, new_n205_, new_n206_ );
nand g089 ( new_n208_, new_n196_, new_n207_ );
nand g090 ( new_n209_, new_n208_, new_n169_ );
nand g091 ( new_n210_, new_n196_, new_n207_, keyIn_0_17 );
nand g092 ( new_n211_, new_n209_, new_n210_ );
nand g093 ( new_n212_, new_n211_, N126 );
xnor g094 ( new_n213_, new_n187_, keyIn_0_3 );
and g095 ( new_n214_, new_n178_, new_n213_ );
nand g096 ( new_n215_, new_n214_, N17 );
or g097 ( new_n216_, new_n215_, keyIn_0_16 );
nand g098 ( new_n217_, new_n215_, keyIn_0_16 );
nand g099 ( new_n218_, new_n216_, N1, new_n217_ );
nand g100 ( new_n219_, new_n218_, N153 );
nand g101 ( new_n220_, new_n212_, new_n168_, new_n219_ );
nand g102 ( new_n221_, new_n212_, new_n219_ );
nand g103 ( new_n222_, new_n221_, keyIn_0_21 );
not g104 ( new_n223_, N268 );
and g105 ( new_n224_, N29, new_n178_, N75, N80 );
nand g106 ( new_n225_, new_n224_, N55 );
or g107 ( new_n226_, new_n225_, keyIn_0_14 );
nand g108 ( new_n227_, new_n225_, keyIn_0_14 );
nand g109 ( new_n228_, new_n226_, new_n223_, new_n227_ );
xnor g110 ( new_n229_, new_n228_, keyIn_0_19 );
nand g111 ( new_n230_, new_n222_, new_n220_, new_n229_ );
nand g112 ( new_n231_, new_n230_, keyIn_0_23 );
not g113 ( new_n232_, keyIn_0_23 );
nand g114 ( new_n233_, new_n222_, new_n232_, new_n220_, new_n229_ );
and g115 ( new_n234_, new_n231_, N201, new_n233_ );
not g116 ( new_n235_, new_n234_ );
not g117 ( new_n236_, N201 );
nand g118 ( new_n237_, new_n231_, new_n233_ );
nand g119 ( new_n238_, new_n237_, new_n236_ );
nand g120 ( new_n239_, new_n235_, N261, new_n238_ );
and g121 ( new_n240_, new_n235_, new_n238_ );
or g122 ( new_n241_, new_n240_, N261 );
nand g123 ( new_n242_, new_n241_, N219, new_n239_ );
nand g124 ( new_n243_, new_n240_, N228 );
nand g125 ( new_n244_, new_n234_, N237 );
nand g126 ( new_n245_, new_n231_, N246, new_n233_ );
nand g127 ( new_n246_, N42, N72, N73 );
or g128 ( new_n247_, new_n143_, new_n246_, new_n146_ );
nor g129 ( new_n248_, new_n247_, new_n236_ );
and g130 ( new_n249_, N121, N210 );
and g131 ( new_n250_, N255, N267 );
nor g132 ( new_n251_, new_n248_, new_n249_, new_n250_ );
and g133 ( new_n252_, new_n244_, new_n245_, new_n251_ );
nand g134 ( new_n253_, new_n242_, new_n243_, new_n252_ );
xor g135 ( N850, new_n253_, keyIn_0_27 );
not g136 ( new_n255_, keyIn_0_25 );
not g137 ( new_n256_, N195 );
not g138 ( new_n257_, keyIn_0_22 );
not g139 ( new_n258_, keyIn_0_20 );
nand g140 ( new_n259_, new_n211_, N121 );
nand g141 ( new_n260_, new_n218_, N149 );
nand g142 ( new_n261_, new_n259_, new_n258_, new_n260_ );
nand g143 ( new_n262_, new_n259_, new_n260_ );
nand g144 ( new_n263_, new_n262_, keyIn_0_20 );
not g145 ( new_n264_, keyIn_0_18 );
xnor g146 ( new_n265_, new_n228_, new_n264_ );
nand g147 ( new_n266_, new_n263_, new_n261_, new_n265_ );
nand g148 ( new_n267_, new_n266_, new_n257_ );
nand g149 ( new_n268_, new_n263_, keyIn_0_22, new_n261_, new_n265_ );
nand g150 ( new_n269_, new_n267_, new_n268_ );
nand g151 ( new_n270_, new_n269_, new_n256_ );
nand g152 ( new_n271_, new_n211_, N116 );
nand g153 ( new_n272_, new_n218_, N146 );
nand g154 ( new_n273_, new_n271_, new_n228_, new_n272_ );
or g155 ( new_n274_, new_n273_, N189 );
nand g156 ( new_n275_, new_n270_, new_n234_, new_n255_, new_n274_ );
nand g157 ( new_n276_, new_n270_, new_n234_, new_n274_ );
nand g158 ( new_n277_, new_n276_, keyIn_0_25 );
nand g159 ( new_n278_, new_n277_, new_n275_ );
nand g160 ( new_n279_, new_n238_, new_n270_, N261, new_n274_ );
nand g161 ( new_n280_, new_n279_, keyIn_0_24 );
nor g162 ( new_n281_, new_n279_, keyIn_0_24 );
not g163 ( new_n282_, new_n269_ );
nand g164 ( new_n283_, new_n282_, N195, new_n274_ );
nand g165 ( new_n284_, new_n273_, N189 );
nand g166 ( new_n285_, new_n283_, new_n284_ );
nor g167 ( new_n286_, new_n281_, new_n285_ );
nand g168 ( new_n287_, new_n286_, keyIn_0_26, new_n278_, new_n280_ );
not g169 ( new_n288_, keyIn_0_26 );
not g170 ( new_n289_, keyIn_0_24 );
and g171 ( new_n290_, new_n238_, N261 );
nand g172 ( new_n291_, new_n290_, new_n289_, new_n270_, new_n274_ );
not g173 ( new_n292_, new_n285_ );
nand g174 ( new_n293_, new_n278_, new_n291_, new_n280_, new_n292_ );
nand g175 ( new_n294_, new_n293_, new_n288_ );
nand g176 ( new_n295_, new_n211_, N111 );
nand g177 ( new_n296_, new_n218_, N143 );
nand g178 ( new_n297_, new_n295_, new_n228_, new_n296_ );
nand g179 ( new_n298_, new_n297_, N183 );
or g180 ( new_n299_, new_n297_, N183 );
nand g181 ( new_n300_, new_n299_, new_n298_ );
nand g182 ( new_n301_, new_n294_, new_n287_, new_n300_ );
nand g183 ( new_n302_, new_n294_, new_n287_ );
nand g184 ( new_n303_, new_n302_, new_n298_, new_n299_ );
nand g185 ( new_n304_, new_n303_, N219, new_n301_ );
nand g186 ( new_n305_, new_n299_, N228, new_n298_ );
nand g187 ( new_n306_, new_n297_, N183, N237 );
nand g188 ( new_n307_, new_n297_, N246 );
not g189 ( new_n308_, N183 );
or g190 ( new_n309_, new_n247_, new_n308_ );
nand g191 ( new_n310_, N106, N210 );
and g192 ( new_n311_, new_n306_, new_n307_, new_n309_, new_n310_ );
nand g193 ( N863, new_n304_, new_n305_, new_n311_ );
nand g194 ( new_n313_, new_n282_, N195 );
or g195 ( new_n314_, new_n290_, new_n234_ );
nand g196 ( new_n315_, new_n314_, new_n270_ );
nand g197 ( new_n316_, new_n315_, new_n313_ );
nand g198 ( new_n317_, new_n274_, new_n284_ );
not g199 ( new_n318_, new_n317_ );
nand g200 ( new_n319_, new_n316_, new_n318_ );
nand g201 ( new_n320_, new_n315_, new_n313_, new_n317_ );
nand g202 ( new_n321_, new_n319_, N219, new_n320_ );
nand g203 ( new_n322_, new_n318_, N228 );
nand g204 ( new_n323_, new_n273_, N189, N237 );
nand g205 ( new_n324_, new_n273_, N246 );
not g206 ( new_n325_, N189 );
nor g207 ( new_n326_, new_n247_, new_n325_ );
and g208 ( new_n327_, N111, N210 );
and g209 ( new_n328_, N255, N259 );
nor g210 ( new_n329_, new_n326_, new_n327_, new_n328_ );
and g211 ( new_n330_, new_n323_, new_n324_, new_n329_ );
nand g212 ( new_n331_, new_n321_, new_n322_, new_n330_ );
xnor g213 ( N864, new_n331_, keyIn_0_30 );
and g214 ( new_n333_, new_n313_, new_n270_ );
or g215 ( new_n334_, new_n314_, new_n333_ );
nand g216 ( new_n335_, new_n314_, new_n333_ );
nand g217 ( new_n336_, new_n334_, N219, new_n335_ );
nand g218 ( new_n337_, new_n333_, N228 );
nand g219 ( new_n338_, new_n282_, N195, N237 );
nand g220 ( new_n339_, new_n282_, N246 );
nor g221 ( new_n340_, new_n247_, new_n256_ );
and g222 ( new_n341_, N116, N210 );
and g223 ( new_n342_, N255, N260 );
nor g224 ( new_n343_, new_n340_, new_n341_, new_n342_ );
and g225 ( new_n344_, new_n338_, new_n339_, new_n343_ );
nand g226 ( new_n345_, new_n336_, new_n337_, new_n344_ );
xor g227 ( N865, new_n345_, keyIn_0_31 );
not g228 ( new_n347_, keyIn_0_29 );
not g229 ( new_n348_, keyIn_0_28 );
nand g230 ( new_n349_, new_n302_, new_n299_ );
nand g231 ( new_n350_, new_n349_, new_n298_ );
nand g232 ( new_n351_, new_n211_, N96 );
nand g233 ( new_n352_, new_n214_, N55 );
xnor g234 ( new_n353_, new_n352_, keyIn_0_12 );
nand g235 ( new_n354_, new_n353_, N146 );
and g236 ( new_n355_, new_n224_, N17 );
nand g237 ( new_n356_, new_n355_, keyIn_0_13 );
or g238 ( new_n357_, new_n355_, keyIn_0_13 );
nand g239 ( new_n358_, new_n357_, new_n223_, new_n356_ );
nand g240 ( new_n359_, N51, N138 );
nand g241 ( new_n360_, new_n351_, new_n354_, new_n358_, new_n359_ );
or g242 ( new_n361_, new_n360_, N165 );
nand g243 ( new_n362_, new_n211_, N101 );
nand g244 ( new_n363_, new_n353_, N149 );
nand g245 ( new_n364_, N17, N138 );
nand g246 ( new_n365_, new_n362_, new_n358_, new_n363_, new_n364_ );
or g247 ( new_n366_, new_n365_, N171 );
nand g248 ( new_n367_, new_n211_, N106 );
nand g249 ( new_n368_, new_n353_, N153 );
nand g250 ( new_n369_, N138, N152 );
nand g251 ( new_n370_, new_n367_, new_n358_, new_n368_, new_n369_ );
or g252 ( new_n371_, new_n370_, N177 );
and g253 ( new_n372_, new_n361_, new_n366_, new_n371_ );
nand g254 ( new_n373_, new_n350_, new_n372_ );
nand g255 ( new_n374_, new_n373_, new_n348_ );
nand g256 ( new_n375_, new_n350_, keyIn_0_28, new_n372_ );
nand g257 ( new_n376_, new_n374_, new_n375_ );
nand g258 ( new_n377_, new_n361_, new_n366_, N177, new_n370_ );
nand g259 ( new_n378_, new_n361_, N171, new_n365_ );
nand g260 ( new_n379_, new_n360_, N165 );
and g261 ( new_n380_, new_n377_, new_n378_, new_n379_ );
nand g262 ( new_n381_, new_n376_, new_n347_, new_n380_ );
nand g263 ( new_n382_, new_n376_, new_n380_ );
nand g264 ( new_n383_, new_n382_, keyIn_0_29 );
nand g265 ( new_n384_, new_n211_, N91 );
nand g266 ( new_n385_, new_n353_, N143 );
nand g267 ( new_n386_, N8, N138 );
nand g268 ( new_n387_, new_n384_, new_n358_, new_n385_, new_n386_ );
or g269 ( new_n388_, new_n387_, N159 );
nand g270 ( new_n389_, new_n383_, new_n381_, new_n388_ );
nand g271 ( new_n390_, new_n387_, N159 );
nand g272 ( N866, new_n389_, new_n390_ );
nand g273 ( new_n392_, new_n370_, N177 );
nand g274 ( new_n393_, new_n371_, new_n392_ );
not g275 ( new_n394_, new_n393_ );
nand g276 ( new_n395_, new_n350_, new_n394_ );
nand g277 ( new_n396_, new_n349_, new_n298_, new_n393_ );
nand g278 ( new_n397_, new_n395_, N219, new_n396_ );
nand g279 ( new_n398_, new_n394_, N228 );
nand g280 ( new_n399_, new_n370_, N177, N237 );
nand g281 ( new_n400_, new_n370_, N246 );
not g282 ( new_n401_, N177 );
or g283 ( new_n402_, new_n247_, new_n401_ );
nand g284 ( new_n403_, N101, N210 );
and g285 ( new_n404_, new_n399_, new_n400_, new_n402_, new_n403_ );
nand g286 ( N874, new_n397_, new_n398_, new_n404_ );
nand g287 ( new_n406_, new_n383_, new_n381_ );
nand g288 ( new_n407_, new_n388_, new_n390_ );
nand g289 ( new_n408_, new_n406_, new_n407_ );
nand g290 ( new_n409_, new_n383_, new_n381_, new_n388_, new_n390_ );
nand g291 ( new_n410_, new_n408_, N219, new_n409_ );
and g292 ( new_n411_, new_n388_, N228, new_n390_ );
nand g293 ( new_n412_, new_n387_, N159, N237 );
nand g294 ( new_n413_, new_n387_, N246 );
not g295 ( new_n414_, N159 );
or g296 ( new_n415_, new_n247_, new_n414_ );
nand g297 ( new_n416_, N210, N268 );
nand g298 ( new_n417_, new_n412_, new_n413_, new_n415_, new_n416_ );
nor g299 ( new_n418_, new_n411_, new_n417_ );
nand g300 ( N878, new_n410_, new_n418_ );
nand g301 ( new_n420_, new_n365_, N171 );
nand g302 ( new_n421_, new_n350_, new_n371_ );
nand g303 ( new_n422_, new_n421_, new_n392_ );
nand g304 ( new_n423_, new_n422_, new_n366_ );
nand g305 ( new_n424_, new_n423_, new_n420_ );
nand g306 ( new_n425_, new_n361_, new_n379_ );
not g307 ( new_n426_, new_n425_ );
nand g308 ( new_n427_, new_n424_, new_n426_ );
nand g309 ( new_n428_, new_n423_, new_n420_, new_n425_ );
nand g310 ( new_n429_, new_n427_, N219, new_n428_ );
nand g311 ( new_n430_, new_n426_, N228 );
nand g312 ( new_n431_, new_n360_, N165, N237 );
nand g313 ( new_n432_, new_n360_, N246 );
not g314 ( new_n433_, N165 );
or g315 ( new_n434_, new_n247_, new_n433_ );
nand g316 ( new_n435_, N91, N210 );
and g317 ( new_n436_, new_n431_, new_n432_, new_n434_, new_n435_ );
nand g318 ( N879, new_n429_, new_n430_, new_n436_ );
nand g319 ( new_n438_, new_n366_, new_n420_ );
not g320 ( new_n439_, new_n438_ );
nand g321 ( new_n440_, new_n422_, new_n439_ );
nand g322 ( new_n441_, new_n421_, new_n392_, new_n438_ );
nand g323 ( new_n442_, new_n440_, N219, new_n441_ );
nand g324 ( new_n443_, new_n439_, N228 );
nand g325 ( new_n444_, new_n365_, N171, N237 );
nand g326 ( new_n445_, new_n365_, N246 );
not g327 ( new_n446_, N171 );
or g328 ( new_n447_, new_n247_, new_n446_ );
nand g329 ( new_n448_, N96, N210 );
and g330 ( new_n449_, new_n444_, new_n445_, new_n447_, new_n448_ );
nand g331 ( N880, new_n442_, new_n443_, new_n449_ );
endmodule