module add_mul_mix_32_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, 
        a_18_, a_19_, a_20_, a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, 
        a_28_, a_29_, a_30_, a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, 
        b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, 
        b_17_, b_18_, b_19_, b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, 
        b_27_, b_28_, b_29_, b_30_, b_31_, c_0_, c_1_, c_2_, c_3_, c_4_, c_5_, 
        c_6_, c_7_, c_8_, c_9_, c_10_, c_11_, c_12_, c_13_, c_14_, c_15_, 
        c_16_, c_17_, c_18_, c_19_, c_20_, c_21_, c_22_, c_23_, c_24_, c_25_, 
        c_26_, c_27_, c_28_, c_29_, c_30_, c_31_, d_0_, d_1_, d_2_, d_3_, d_4_, 
        d_5_, d_6_, d_7_, d_8_, d_9_, d_10_, d_11_, d_12_, d_13_, d_14_, d_15_, 
        d_16_, d_17_, d_18_, d_19_, d_20_, d_21_, d_22_, d_23_, d_24_, d_25_, 
        d_26_, d_27_, d_28_, d_29_, d_30_, d_31_, Result_0_, Result_1_, 
        Result_2_, Result_3_, Result_4_, Result_5_, Result_6_, Result_7_, 
        Result_8_, Result_9_, Result_10_, Result_11_, Result_12_, Result_13_, 
        Result_14_, Result_15_, Result_16_, Result_17_, Result_18_, Result_19_, 
        Result_20_, Result_21_, Result_22_, Result_23_, Result_24_, Result_25_, 
        Result_26_, Result_27_, Result_28_, Result_29_, Result_30_, Result_31_, 
        Result_32_, Result_33_, Result_34_, Result_35_, Result_36_, Result_37_, 
        Result_38_, Result_39_, Result_40_, Result_41_, Result_42_, Result_43_, 
        Result_44_, Result_45_, Result_46_, Result_47_, Result_48_, Result_49_, 
        Result_50_, Result_51_, Result_52_, Result_53_, Result_54_, Result_55_, 
        Result_56_, Result_57_, Result_58_, Result_59_, Result_60_, Result_61_, 
        Result_62_, Result_63_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, a_19_, a_20_,
         a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, a_29_, a_30_,
         a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_,
         b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, b_18_, b_19_,
         b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, b_28_, b_29_,
         b_30_, b_31_, c_0_, c_1_, c_2_, c_3_, c_4_, c_5_, c_6_, c_7_, c_8_,
         c_9_, c_10_, c_11_, c_12_, c_13_, c_14_, c_15_, c_16_, c_17_, c_18_,
         c_19_, c_20_, c_21_, c_22_, c_23_, c_24_, c_25_, c_26_, c_27_, c_28_,
         c_29_, c_30_, c_31_, d_0_, d_1_, d_2_, d_3_, d_4_, d_5_, d_6_, d_7_,
         d_8_, d_9_, d_10_, d_11_, d_12_, d_13_, d_14_, d_15_, d_16_, d_17_,
         d_18_, d_19_, d_20_, d_21_, d_22_, d_23_, d_24_, d_25_, d_26_, d_27_,
         d_28_, d_29_, d_30_, d_31_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_,
         Result_32_, Result_33_, Result_34_, Result_35_, Result_36_,
         Result_37_, Result_38_, Result_39_, Result_40_, Result_41_,
         Result_42_, Result_43_, Result_44_, Result_45_, Result_46_,
         Result_47_, Result_48_, Result_49_, Result_50_, Result_51_,
         Result_52_, Result_53_, Result_54_, Result_55_, Result_56_,
         Result_57_, Result_58_, Result_59_, Result_60_, Result_61_,
         Result_62_, Result_63_;
  wire   n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231;

  INV_X1 U7669 ( .A(n8518), .ZN(n7605) );
  INV_X1 U7670 ( .A(n7605), .ZN(n7606) );
  INV_X1 U7671 ( .A(n8023), .ZN(n7607) );
  INV_X1 U7672 ( .A(n7607), .ZN(n7608) );
  INV_X1 U7673 ( .A(n8056), .ZN(n7609) );
  INV_X1 U7674 ( .A(n7609), .ZN(n7610) );
  INV_X1 U7675 ( .A(n8105), .ZN(n7611) );
  INV_X1 U7676 ( .A(n7611), .ZN(n7612) );
  INV_X1 U7677 ( .A(n8152), .ZN(n7613) );
  INV_X1 U7678 ( .A(n7613), .ZN(n7614) );
  INV_X1 U7679 ( .A(n8644), .ZN(n7615) );
  INV_X1 U7680 ( .A(n7615), .ZN(n7616) );
  INV_X1 U7681 ( .A(n8639), .ZN(n7617) );
  INV_X1 U7682 ( .A(n7617), .ZN(n7618) );
  INV_X1 U7683 ( .A(n8634), .ZN(n7619) );
  INV_X1 U7684 ( .A(n7619), .ZN(n7620) );
  INV_X1 U7685 ( .A(n8629), .ZN(n7621) );
  INV_X1 U7686 ( .A(n7621), .ZN(n7622) );
  INV_X1 U7687 ( .A(n8624), .ZN(n7623) );
  INV_X1 U7688 ( .A(n7623), .ZN(n7624) );
  INV_X1 U7689 ( .A(n8619), .ZN(n7625) );
  INV_X1 U7690 ( .A(n7625), .ZN(n7626) );
  INV_X1 U7691 ( .A(n8614), .ZN(n7627) );
  INV_X1 U7692 ( .A(n7627), .ZN(n7628) );
  INV_X1 U7693 ( .A(n8609), .ZN(n7629) );
  INV_X1 U7694 ( .A(n7629), .ZN(n7630) );
  INV_X1 U7695 ( .A(n8604), .ZN(n7631) );
  INV_X1 U7696 ( .A(n7631), .ZN(n7632) );
  INV_X1 U7697 ( .A(n8599), .ZN(n7633) );
  INV_X1 U7698 ( .A(n7633), .ZN(n7634) );
  INV_X1 U7699 ( .A(n8594), .ZN(n7635) );
  INV_X1 U7700 ( .A(n7635), .ZN(n7636) );
  INV_X1 U7701 ( .A(n8589), .ZN(n7637) );
  INV_X1 U7702 ( .A(n7637), .ZN(n7638) );
  INV_X1 U7703 ( .A(n8584), .ZN(n7639) );
  INV_X1 U7704 ( .A(n7639), .ZN(n7640) );
  INV_X1 U7705 ( .A(n8579), .ZN(n7641) );
  INV_X1 U7706 ( .A(n7641), .ZN(n7642) );
  INV_X1 U7707 ( .A(n8574), .ZN(n7643) );
  INV_X1 U7708 ( .A(n7643), .ZN(n7644) );
  INV_X1 U7709 ( .A(n8569), .ZN(n7645) );
  INV_X1 U7710 ( .A(n7645), .ZN(n7646) );
  INV_X1 U7711 ( .A(n8564), .ZN(n7647) );
  INV_X1 U7712 ( .A(n7647), .ZN(n7648) );
  INV_X1 U7713 ( .A(n8559), .ZN(n7649) );
  INV_X1 U7714 ( .A(n7649), .ZN(n7650) );
  INV_X1 U7715 ( .A(n8554), .ZN(n7651) );
  INV_X1 U7716 ( .A(n7651), .ZN(n7652) );
  INV_X1 U7717 ( .A(n8549), .ZN(n7653) );
  INV_X1 U7718 ( .A(n7653), .ZN(n7654) );
  INV_X1 U7719 ( .A(n8544), .ZN(n7655) );
  INV_X1 U7720 ( .A(n7655), .ZN(n7656) );
  INV_X1 U7721 ( .A(n8539), .ZN(n7657) );
  INV_X1 U7722 ( .A(n7657), .ZN(n7658) );
  INV_X1 U7723 ( .A(n8534), .ZN(n7659) );
  INV_X1 U7724 ( .A(n7659), .ZN(n7660) );
  INV_X1 U7725 ( .A(n8529), .ZN(n7661) );
  INV_X1 U7726 ( .A(n7661), .ZN(n7662) );
  INV_X1 U7727 ( .A(n7960), .ZN(n7663) );
  INV_X1 U7728 ( .A(n7663), .ZN(n7664) );
  INV_X1 U7729 ( .A(n7694), .ZN(n7665) );
  INV_X1 U7730 ( .A(n14653), .ZN(n7666) );
  INV_X1 U7731 ( .A(n8523), .ZN(n7667) );
  XOR2_X1 U7732 ( .A(n7668), .B(n7669), .Z(Result_9_) );
  AND2_X1 U7733 ( .A1(n7670), .A2(n7671), .ZN(n7669) );
  OR2_X1 U7734 ( .A1(n7672), .A2(n7673), .ZN(n7671) );
  AND2_X1 U7735 ( .A1(n7674), .A2(n7675), .ZN(n7673) );
  INV_X1 U7736 ( .A(n7676), .ZN(n7670) );
  XOR2_X1 U7737 ( .A(n7677), .B(n7678), .Z(Result_8_) );
  XOR2_X1 U7738 ( .A(n7679), .B(n7680), .Z(Result_7_) );
  AND2_X1 U7739 ( .A1(n7681), .A2(n7682), .ZN(n7680) );
  OR2_X1 U7740 ( .A1(n7683), .A2(n7684), .ZN(n7682) );
  AND2_X1 U7741 ( .A1(n7685), .A2(n7686), .ZN(n7684) );
  INV_X1 U7742 ( .A(n7687), .ZN(n7681) );
  XOR2_X1 U7743 ( .A(n7688), .B(n7689), .Z(Result_6_) );
  AND2_X1 U7744 ( .A1(n7690), .A2(n7691), .ZN(Result_63_) );
  OR2_X1 U7745 ( .A1(n7692), .A2(n7693), .ZN(Result_62_) );
  AND2_X1 U7746 ( .A1(n7694), .A2(n7695), .ZN(n7693) );
  OR2_X1 U7747 ( .A1(n7696), .A2(n7697), .ZN(n7695) );
  AND2_X1 U7748 ( .A1(n7691), .A2(n7698), .ZN(n7696) );
  AND2_X1 U7749 ( .A1(n7690), .A2(n7699), .ZN(n7692) );
  OR2_X1 U7750 ( .A1(n7700), .A2(n7701), .ZN(n7699) );
  AND2_X1 U7751 ( .A1(n7665), .A2(n7703), .ZN(n7700) );
  XOR2_X1 U7752 ( .A(n7704), .B(n7705), .Z(Result_61_) );
  XNOR2_X1 U7753 ( .A(n7706), .B(n7707), .ZN(n7705) );
  XNOR2_X1 U7754 ( .A(n7708), .B(n7709), .ZN(Result_60_) );
  XOR2_X1 U7755 ( .A(n7710), .B(n7711), .Z(n7709) );
  XOR2_X1 U7756 ( .A(n7712), .B(n7713), .Z(Result_5_) );
  AND2_X1 U7757 ( .A1(n7714), .A2(n7715), .ZN(n7713) );
  OR2_X1 U7758 ( .A1(n7716), .A2(n7717), .ZN(n7715) );
  AND2_X1 U7759 ( .A1(n7718), .A2(n7719), .ZN(n7717) );
  INV_X1 U7760 ( .A(n7720), .ZN(n7714) );
  XNOR2_X1 U7761 ( .A(n7721), .B(n7722), .ZN(Result_59_) );
  XOR2_X1 U7762 ( .A(n7723), .B(n7724), .Z(n7722) );
  XNOR2_X1 U7763 ( .A(n7725), .B(n7726), .ZN(Result_58_) );
  XOR2_X1 U7764 ( .A(n7727), .B(n7728), .Z(n7726) );
  XNOR2_X1 U7765 ( .A(n7729), .B(n7730), .ZN(Result_57_) );
  XOR2_X1 U7766 ( .A(n7731), .B(n7732), .Z(n7730) );
  XNOR2_X1 U7767 ( .A(n7733), .B(n7734), .ZN(Result_56_) );
  XOR2_X1 U7768 ( .A(n7735), .B(n7736), .Z(n7734) );
  XNOR2_X1 U7769 ( .A(n7737), .B(n7738), .ZN(Result_55_) );
  XOR2_X1 U7770 ( .A(n7739), .B(n7740), .Z(n7738) );
  XNOR2_X1 U7771 ( .A(n7741), .B(n7742), .ZN(Result_54_) );
  XOR2_X1 U7772 ( .A(n7743), .B(n7744), .Z(n7742) );
  XNOR2_X1 U7773 ( .A(n7745), .B(n7746), .ZN(Result_53_) );
  XOR2_X1 U7774 ( .A(n7747), .B(n7748), .Z(n7746) );
  XNOR2_X1 U7775 ( .A(n7749), .B(n7750), .ZN(Result_52_) );
  XOR2_X1 U7776 ( .A(n7751), .B(n7752), .Z(n7750) );
  XNOR2_X1 U7777 ( .A(n7753), .B(n7754), .ZN(Result_51_) );
  XOR2_X1 U7778 ( .A(n7755), .B(n7756), .Z(n7754) );
  XNOR2_X1 U7779 ( .A(n7757), .B(n7758), .ZN(Result_50_) );
  XOR2_X1 U7780 ( .A(n7759), .B(n7760), .Z(n7758) );
  XOR2_X1 U7781 ( .A(n7761), .B(n7762), .Z(Result_4_) );
  XNOR2_X1 U7782 ( .A(n7763), .B(n7764), .ZN(Result_49_) );
  XOR2_X1 U7783 ( .A(n7765), .B(n7766), .Z(n7764) );
  XNOR2_X1 U7784 ( .A(n7767), .B(n7768), .ZN(Result_48_) );
  XOR2_X1 U7785 ( .A(n7769), .B(n7770), .Z(n7768) );
  XNOR2_X1 U7786 ( .A(n7771), .B(n7772), .ZN(Result_47_) );
  XOR2_X1 U7787 ( .A(n7773), .B(n7774), .Z(n7772) );
  XNOR2_X1 U7788 ( .A(n7775), .B(n7776), .ZN(Result_46_) );
  XOR2_X1 U7789 ( .A(n7777), .B(n7778), .Z(n7776) );
  XNOR2_X1 U7790 ( .A(n7779), .B(n7780), .ZN(Result_45_) );
  XOR2_X1 U7791 ( .A(n7781), .B(n7782), .Z(n7780) );
  XNOR2_X1 U7792 ( .A(n7783), .B(n7784), .ZN(Result_44_) );
  XOR2_X1 U7793 ( .A(n7785), .B(n7786), .Z(n7784) );
  XNOR2_X1 U7794 ( .A(n7787), .B(n7788), .ZN(Result_43_) );
  XOR2_X1 U7795 ( .A(n7789), .B(n7790), .Z(n7788) );
  XNOR2_X1 U7796 ( .A(n7791), .B(n7792), .ZN(Result_42_) );
  XOR2_X1 U7797 ( .A(n7793), .B(n7794), .Z(n7792) );
  XNOR2_X1 U7798 ( .A(n7795), .B(n7796), .ZN(Result_41_) );
  XOR2_X1 U7799 ( .A(n7797), .B(n7798), .Z(n7796) );
  XNOR2_X1 U7800 ( .A(n7799), .B(n7800), .ZN(Result_40_) );
  XOR2_X1 U7801 ( .A(n7801), .B(n7802), .Z(n7800) );
  XOR2_X1 U7802 ( .A(n7803), .B(n7804), .Z(Result_3_) );
  AND2_X1 U7803 ( .A1(n7805), .A2(n7806), .ZN(n7804) );
  OR2_X1 U7804 ( .A1(n7807), .A2(n7808), .ZN(n7806) );
  AND2_X1 U7805 ( .A1(n7809), .A2(n7810), .ZN(n7808) );
  INV_X1 U7806 ( .A(n7811), .ZN(n7805) );
  XNOR2_X1 U7807 ( .A(n7812), .B(n7813), .ZN(Result_39_) );
  XOR2_X1 U7808 ( .A(n7814), .B(n7815), .Z(n7813) );
  XNOR2_X1 U7809 ( .A(n7816), .B(n7817), .ZN(Result_38_) );
  XOR2_X1 U7810 ( .A(n7818), .B(n7819), .Z(n7817) );
  XNOR2_X1 U7811 ( .A(n7820), .B(n7821), .ZN(Result_37_) );
  XOR2_X1 U7812 ( .A(n7822), .B(n7823), .Z(n7821) );
  XNOR2_X1 U7813 ( .A(n7824), .B(n7825), .ZN(Result_36_) );
  XOR2_X1 U7814 ( .A(n7826), .B(n7827), .Z(n7825) );
  XNOR2_X1 U7815 ( .A(n7828), .B(n7829), .ZN(Result_35_) );
  XOR2_X1 U7816 ( .A(n7830), .B(n7831), .Z(n7829) );
  XNOR2_X1 U7817 ( .A(n7832), .B(n7833), .ZN(Result_34_) );
  XOR2_X1 U7818 ( .A(n7834), .B(n7835), .Z(n7833) );
  XNOR2_X1 U7819 ( .A(n7836), .B(n7837), .ZN(Result_33_) );
  XOR2_X1 U7820 ( .A(n7838), .B(n7839), .Z(n7837) );
  XNOR2_X1 U7821 ( .A(n7840), .B(n7841), .ZN(Result_32_) );
  XOR2_X1 U7822 ( .A(n7842), .B(n7843), .Z(n7841) );
  XNOR2_X1 U7823 ( .A(n7844), .B(n7845), .ZN(Result_31_) );
  AND2_X1 U7824 ( .A1(n7846), .A2(n7847), .ZN(Result_30_) );
  OR2_X1 U7825 ( .A1(n7848), .A2(n7849), .ZN(n7846) );
  AND2_X1 U7826 ( .A1(n7850), .A2(n7845), .ZN(n7848) );
  XOR2_X1 U7827 ( .A(n7851), .B(n7852), .Z(Result_2_) );
  XNOR2_X1 U7828 ( .A(n7853), .B(n7854), .ZN(Result_29_) );
  OR2_X1 U7829 ( .A1(n7855), .A2(n7856), .ZN(n7854) );
  INV_X1 U7830 ( .A(n7857), .ZN(n7856) );
  XOR2_X1 U7831 ( .A(n7858), .B(n7859), .Z(Result_28_) );
  OR2_X1 U7832 ( .A1(n7860), .A2(n7861), .ZN(n7858) );
  INV_X1 U7833 ( .A(n7862), .ZN(n7861) );
  XOR2_X1 U7834 ( .A(n7863), .B(n7864), .Z(Result_27_) );
  OR2_X1 U7835 ( .A1(n7865), .A2(n7866), .ZN(n7863) );
  INV_X1 U7836 ( .A(n7867), .ZN(n7866) );
  XOR2_X1 U7837 ( .A(n7868), .B(n7869), .Z(Result_26_) );
  OR2_X1 U7838 ( .A1(n7870), .A2(n7871), .ZN(n7868) );
  INV_X1 U7839 ( .A(n7872), .ZN(n7870) );
  XOR2_X1 U7840 ( .A(n7873), .B(n7874), .Z(Result_25_) );
  OR2_X1 U7841 ( .A1(n7875), .A2(n7876), .ZN(n7873) );
  INV_X1 U7842 ( .A(n7877), .ZN(n7876) );
  XOR2_X1 U7843 ( .A(n7878), .B(n7879), .Z(Result_24_) );
  OR2_X1 U7844 ( .A1(n7880), .A2(n7881), .ZN(n7878) );
  INV_X1 U7845 ( .A(n7882), .ZN(n7881) );
  XOR2_X1 U7846 ( .A(n7883), .B(n7884), .Z(Result_23_) );
  OR2_X1 U7847 ( .A1(n7885), .A2(n7886), .ZN(n7883) );
  INV_X1 U7848 ( .A(n7887), .ZN(n7886) );
  XOR2_X1 U7849 ( .A(n7888), .B(n7889), .Z(Result_22_) );
  OR2_X1 U7850 ( .A1(n7890), .A2(n7891), .ZN(n7888) );
  INV_X1 U7851 ( .A(n7892), .ZN(n7891) );
  XOR2_X1 U7852 ( .A(n7893), .B(n7894), .Z(Result_21_) );
  OR2_X1 U7853 ( .A1(n7895), .A2(n7896), .ZN(n7893) );
  XOR2_X1 U7854 ( .A(n7897), .B(n7898), .Z(Result_20_) );
  OR2_X1 U7855 ( .A1(n7899), .A2(n7900), .ZN(n7897) );
  INV_X1 U7856 ( .A(n7901), .ZN(n7900) );
  XOR2_X1 U7857 ( .A(n7902), .B(n7903), .Z(Result_1_) );
  AND2_X1 U7858 ( .A1(n7904), .A2(n7905), .ZN(n7903) );
  OR2_X1 U7859 ( .A1(n7906), .A2(n7907), .ZN(n7905) );
  AND2_X1 U7860 ( .A1(n7908), .A2(n7909), .ZN(n7906) );
  INV_X1 U7861 ( .A(n7910), .ZN(n7904) );
  XOR2_X1 U7862 ( .A(n7911), .B(n7912), .Z(Result_19_) );
  OR2_X1 U7863 ( .A1(n7913), .A2(n7914), .ZN(n7911) );
  INV_X1 U7864 ( .A(n7915), .ZN(n7914) );
  XOR2_X1 U7865 ( .A(n7916), .B(n7917), .Z(Result_18_) );
  OR2_X1 U7866 ( .A1(n7918), .A2(n7919), .ZN(n7916) );
  INV_X1 U7867 ( .A(n7920), .ZN(n7919) );
  XNOR2_X1 U7868 ( .A(n7921), .B(n7922), .ZN(Result_17_) );
  AND2_X1 U7869 ( .A1(n7923), .A2(n7924), .ZN(n7922) );
  INV_X1 U7870 ( .A(n7925), .ZN(n7924) );
  XNOR2_X1 U7871 ( .A(n7926), .B(n7927), .ZN(Result_16_) );
  AND2_X1 U7872 ( .A1(n7928), .A2(n7929), .ZN(n7927) );
  INV_X1 U7873 ( .A(n7930), .ZN(n7929) );
  XNOR2_X1 U7874 ( .A(n7931), .B(n7932), .ZN(Result_15_) );
  AND2_X1 U7875 ( .A1(n7933), .A2(n7934), .ZN(n7932) );
  INV_X1 U7876 ( .A(n7935), .ZN(n7934) );
  XOR2_X1 U7877 ( .A(n7936), .B(n7937), .Z(Result_14_) );
  XNOR2_X1 U7878 ( .A(n7938), .B(n7939), .ZN(n7936) );
  XOR2_X1 U7879 ( .A(n7940), .B(n7941), .Z(Result_13_) );
  XNOR2_X1 U7880 ( .A(n7942), .B(n7943), .ZN(n7940) );
  XNOR2_X1 U7881 ( .A(n7944), .B(n7945), .ZN(Result_12_) );
  XOR2_X1 U7882 ( .A(n7946), .B(n7947), .Z(n7944) );
  XNOR2_X1 U7883 ( .A(n7948), .B(n7949), .ZN(Result_11_) );
  XOR2_X1 U7884 ( .A(n7950), .B(n7951), .Z(n7948) );
  XOR2_X1 U7885 ( .A(n7952), .B(n7953), .Z(Result_10_) );
  OR2_X1 U7886 ( .A1(n7954), .A2(n7955), .ZN(n7952) );
  OR3_X1 U7887 ( .A1(n7910), .A2(n7956), .A3(n7957), .ZN(Result_0_) );
  INV_X1 U7888 ( .A(n7958), .ZN(n7957) );
  OR2_X1 U7889 ( .A1(n7959), .A2(n7664), .ZN(n7958) );
  AND2_X1 U7890 ( .A1(n7902), .A2(n7907), .ZN(n7956) );
  AND2_X1 U7891 ( .A1(n7851), .A2(n7852), .ZN(n7902) );
  XNOR2_X1 U7892 ( .A(n7909), .B(n7961), .ZN(n7852) );
  OR2_X1 U7893 ( .A1(n7962), .A2(n7963), .ZN(n7851) );
  OR2_X1 U7894 ( .A1(n7964), .A2(n7811), .ZN(n7962) );
  AND3_X1 U7895 ( .A1(n7810), .A2(n7809), .A3(n7807), .ZN(n7811) );
  INV_X1 U7896 ( .A(n7965), .ZN(n7809) );
  AND2_X1 U7897 ( .A1(n7803), .A2(n7807), .ZN(n7964) );
  INV_X1 U7898 ( .A(n7966), .ZN(n7807) );
  OR2_X1 U7899 ( .A1(n7967), .A2(n7963), .ZN(n7966) );
  INV_X1 U7900 ( .A(n7968), .ZN(n7963) );
  OR2_X1 U7901 ( .A1(n7969), .A2(n7970), .ZN(n7968) );
  AND2_X1 U7902 ( .A1(n7969), .A2(n7970), .ZN(n7967) );
  OR2_X1 U7903 ( .A1(n7971), .A2(n7972), .ZN(n7970) );
  AND2_X1 U7904 ( .A1(n7973), .A2(n7974), .ZN(n7972) );
  AND2_X1 U7905 ( .A1(n7975), .A2(n7976), .ZN(n7971) );
  OR2_X1 U7906 ( .A1(n7974), .A2(n7973), .ZN(n7976) );
  XOR2_X1 U7907 ( .A(n7977), .B(n7978), .Z(n7969) );
  XOR2_X1 U7908 ( .A(n7979), .B(n7980), .Z(n7978) );
  AND2_X1 U7909 ( .A1(n7761), .A2(n7762), .ZN(n7803) );
  XNOR2_X1 U7910 ( .A(n7810), .B(n7965), .ZN(n7762) );
  OR2_X1 U7911 ( .A1(n7981), .A2(n7982), .ZN(n7965) );
  AND2_X1 U7912 ( .A1(n7983), .A2(n7984), .ZN(n7982) );
  AND2_X1 U7913 ( .A1(n7985), .A2(n7986), .ZN(n7981) );
  OR2_X1 U7914 ( .A1(n7984), .A2(n7983), .ZN(n7986) );
  XNOR2_X1 U7915 ( .A(n7975), .B(n7987), .ZN(n7810) );
  XOR2_X1 U7916 ( .A(n7974), .B(n7973), .Z(n7987) );
  OR2_X1 U7917 ( .A1(n7988), .A2(n7664), .ZN(n7973) );
  OR2_X1 U7918 ( .A1(n7989), .A2(n7990), .ZN(n7974) );
  AND2_X1 U7919 ( .A1(n7991), .A2(n7992), .ZN(n7990) );
  AND2_X1 U7920 ( .A1(n7993), .A2(n7994), .ZN(n7989) );
  OR2_X1 U7921 ( .A1(n7992), .A2(n7991), .ZN(n7994) );
  XOR2_X1 U7922 ( .A(n7995), .B(n7996), .Z(n7975) );
  XOR2_X1 U7923 ( .A(n7997), .B(n7998), .Z(n7996) );
  OR2_X1 U7924 ( .A1(n7999), .A2(n8000), .ZN(n7761) );
  OR2_X1 U7925 ( .A1(n8001), .A2(n7720), .ZN(n7999) );
  AND3_X1 U7926 ( .A1(n7719), .A2(n7718), .A3(n7716), .ZN(n7720) );
  INV_X1 U7927 ( .A(n8002), .ZN(n7718) );
  AND2_X1 U7928 ( .A1(n7712), .A2(n7716), .ZN(n8001) );
  INV_X1 U7929 ( .A(n8003), .ZN(n7716) );
  OR2_X1 U7930 ( .A1(n8004), .A2(n8000), .ZN(n8003) );
  INV_X1 U7931 ( .A(n8005), .ZN(n8000) );
  OR2_X1 U7932 ( .A1(n8006), .A2(n8007), .ZN(n8005) );
  AND2_X1 U7933 ( .A1(n8006), .A2(n8007), .ZN(n8004) );
  OR2_X1 U7934 ( .A1(n8008), .A2(n8009), .ZN(n8007) );
  AND2_X1 U7935 ( .A1(n8010), .A2(n8011), .ZN(n8009) );
  AND2_X1 U7936 ( .A1(n8012), .A2(n8013), .ZN(n8008) );
  OR2_X1 U7937 ( .A1(n8011), .A2(n8010), .ZN(n8013) );
  XOR2_X1 U7938 ( .A(n7985), .B(n8014), .Z(n8006) );
  XOR2_X1 U7939 ( .A(n7984), .B(n7983), .Z(n8014) );
  OR2_X1 U7940 ( .A1(n8015), .A2(n7664), .ZN(n7983) );
  OR2_X1 U7941 ( .A1(n8016), .A2(n8017), .ZN(n7984) );
  AND2_X1 U7942 ( .A1(n8018), .A2(n8019), .ZN(n8017) );
  AND2_X1 U7943 ( .A1(n8020), .A2(n8021), .ZN(n8016) );
  OR2_X1 U7944 ( .A1(n8019), .A2(n8018), .ZN(n8021) );
  XOR2_X1 U7945 ( .A(n7993), .B(n8022), .Z(n7985) );
  XOR2_X1 U7946 ( .A(n7992), .B(n7991), .Z(n8022) );
  OR2_X1 U7947 ( .A1(n7988), .A2(n7608), .ZN(n7991) );
  OR2_X1 U7948 ( .A1(n8024), .A2(n8025), .ZN(n7992) );
  AND2_X1 U7949 ( .A1(n8026), .A2(n8027), .ZN(n8025) );
  AND2_X1 U7950 ( .A1(n8028), .A2(n8029), .ZN(n8024) );
  OR2_X1 U7951 ( .A1(n8027), .A2(n8026), .ZN(n8029) );
  XOR2_X1 U7952 ( .A(n8030), .B(n8031), .Z(n7993) );
  XOR2_X1 U7953 ( .A(n8032), .B(n8033), .Z(n8031) );
  AND2_X1 U7954 ( .A1(n7688), .A2(n7689), .ZN(n7712) );
  XNOR2_X1 U7955 ( .A(n7719), .B(n8002), .ZN(n7689) );
  OR2_X1 U7956 ( .A1(n8034), .A2(n8035), .ZN(n8002) );
  AND2_X1 U7957 ( .A1(n8036), .A2(n8037), .ZN(n8035) );
  AND2_X1 U7958 ( .A1(n8038), .A2(n8039), .ZN(n8034) );
  OR2_X1 U7959 ( .A1(n8037), .A2(n8036), .ZN(n8039) );
  XNOR2_X1 U7960 ( .A(n8012), .B(n8040), .ZN(n7719) );
  XOR2_X1 U7961 ( .A(n8011), .B(n8010), .Z(n8040) );
  OR2_X1 U7962 ( .A1(n8041), .A2(n7664), .ZN(n8010) );
  OR2_X1 U7963 ( .A1(n8042), .A2(n8043), .ZN(n8011) );
  AND2_X1 U7964 ( .A1(n8044), .A2(n8045), .ZN(n8043) );
  AND2_X1 U7965 ( .A1(n8046), .A2(n8047), .ZN(n8042) );
  OR2_X1 U7966 ( .A1(n8045), .A2(n8044), .ZN(n8047) );
  XOR2_X1 U7967 ( .A(n8020), .B(n8048), .Z(n8012) );
  XOR2_X1 U7968 ( .A(n8019), .B(n8018), .Z(n8048) );
  OR2_X1 U7969 ( .A1(n8015), .A2(n7608), .ZN(n8018) );
  OR2_X1 U7970 ( .A1(n8049), .A2(n8050), .ZN(n8019) );
  AND2_X1 U7971 ( .A1(n8051), .A2(n8052), .ZN(n8050) );
  AND2_X1 U7972 ( .A1(n8053), .A2(n8054), .ZN(n8049) );
  OR2_X1 U7973 ( .A1(n8052), .A2(n8051), .ZN(n8054) );
  XOR2_X1 U7974 ( .A(n8028), .B(n8055), .Z(n8020) );
  XOR2_X1 U7975 ( .A(n8027), .B(n8026), .Z(n8055) );
  OR2_X1 U7976 ( .A1(n7988), .A2(n7610), .ZN(n8026) );
  OR2_X1 U7977 ( .A1(n8057), .A2(n8058), .ZN(n8027) );
  AND2_X1 U7978 ( .A1(n8059), .A2(n8060), .ZN(n8058) );
  AND2_X1 U7979 ( .A1(n8061), .A2(n8062), .ZN(n8057) );
  OR2_X1 U7980 ( .A1(n8060), .A2(n8059), .ZN(n8062) );
  XOR2_X1 U7981 ( .A(n8063), .B(n8064), .Z(n8028) );
  XOR2_X1 U7982 ( .A(n8065), .B(n8066), .Z(n8064) );
  OR2_X1 U7983 ( .A1(n8067), .A2(n8068), .ZN(n7688) );
  OR2_X1 U7984 ( .A1(n8069), .A2(n7687), .ZN(n8067) );
  AND3_X1 U7985 ( .A1(n7686), .A2(n7685), .A3(n7683), .ZN(n7687) );
  INV_X1 U7986 ( .A(n8070), .ZN(n7685) );
  AND2_X1 U7987 ( .A1(n7679), .A2(n7683), .ZN(n8069) );
  INV_X1 U7988 ( .A(n8071), .ZN(n7683) );
  OR2_X1 U7989 ( .A1(n8072), .A2(n8068), .ZN(n8071) );
  INV_X1 U7990 ( .A(n8073), .ZN(n8068) );
  OR2_X1 U7991 ( .A1(n8074), .A2(n8075), .ZN(n8073) );
  AND2_X1 U7992 ( .A1(n8074), .A2(n8075), .ZN(n8072) );
  OR2_X1 U7993 ( .A1(n8076), .A2(n8077), .ZN(n8075) );
  AND2_X1 U7994 ( .A1(n8078), .A2(n8079), .ZN(n8077) );
  AND2_X1 U7995 ( .A1(n8080), .A2(n8081), .ZN(n8076) );
  OR2_X1 U7996 ( .A1(n8079), .A2(n8078), .ZN(n8081) );
  XOR2_X1 U7997 ( .A(n8038), .B(n8082), .Z(n8074) );
  XOR2_X1 U7998 ( .A(n8037), .B(n8036), .Z(n8082) );
  OR2_X1 U7999 ( .A1(n8083), .A2(n7664), .ZN(n8036) );
  OR2_X1 U8000 ( .A1(n8084), .A2(n8085), .ZN(n8037) );
  AND2_X1 U8001 ( .A1(n8086), .A2(n8087), .ZN(n8085) );
  AND2_X1 U8002 ( .A1(n8088), .A2(n8089), .ZN(n8084) );
  OR2_X1 U8003 ( .A1(n8087), .A2(n8086), .ZN(n8089) );
  XOR2_X1 U8004 ( .A(n8046), .B(n8090), .Z(n8038) );
  XOR2_X1 U8005 ( .A(n8045), .B(n8044), .Z(n8090) );
  OR2_X1 U8006 ( .A1(n8041), .A2(n7608), .ZN(n8044) );
  OR2_X1 U8007 ( .A1(n8091), .A2(n8092), .ZN(n8045) );
  AND2_X1 U8008 ( .A1(n8093), .A2(n8094), .ZN(n8092) );
  AND2_X1 U8009 ( .A1(n8095), .A2(n8096), .ZN(n8091) );
  OR2_X1 U8010 ( .A1(n8094), .A2(n8093), .ZN(n8096) );
  XOR2_X1 U8011 ( .A(n8053), .B(n8097), .Z(n8046) );
  XOR2_X1 U8012 ( .A(n8052), .B(n8051), .Z(n8097) );
  OR2_X1 U8013 ( .A1(n8015), .A2(n7610), .ZN(n8051) );
  OR2_X1 U8014 ( .A1(n8098), .A2(n8099), .ZN(n8052) );
  AND2_X1 U8015 ( .A1(n8100), .A2(n8101), .ZN(n8099) );
  AND2_X1 U8016 ( .A1(n8102), .A2(n8103), .ZN(n8098) );
  OR2_X1 U8017 ( .A1(n8101), .A2(n8100), .ZN(n8103) );
  XOR2_X1 U8018 ( .A(n8061), .B(n8104), .Z(n8053) );
  XOR2_X1 U8019 ( .A(n8060), .B(n8059), .Z(n8104) );
  OR2_X1 U8020 ( .A1(n7988), .A2(n7612), .ZN(n8059) );
  OR2_X1 U8021 ( .A1(n8106), .A2(n8107), .ZN(n8060) );
  AND2_X1 U8022 ( .A1(n8108), .A2(n8109), .ZN(n8107) );
  AND2_X1 U8023 ( .A1(n8110), .A2(n8111), .ZN(n8106) );
  OR2_X1 U8024 ( .A1(n8109), .A2(n8108), .ZN(n8111) );
  XOR2_X1 U8025 ( .A(n8112), .B(n8113), .Z(n8061) );
  XOR2_X1 U8026 ( .A(n8114), .B(n8115), .Z(n8113) );
  AND2_X1 U8027 ( .A1(n7677), .A2(n7678), .ZN(n7679) );
  XNOR2_X1 U8028 ( .A(n7686), .B(n8070), .ZN(n7678) );
  OR2_X1 U8029 ( .A1(n8116), .A2(n8117), .ZN(n8070) );
  AND2_X1 U8030 ( .A1(n8118), .A2(n8119), .ZN(n8117) );
  AND2_X1 U8031 ( .A1(n8120), .A2(n8121), .ZN(n8116) );
  OR2_X1 U8032 ( .A1(n8119), .A2(n8118), .ZN(n8121) );
  XNOR2_X1 U8033 ( .A(n8080), .B(n8122), .ZN(n7686) );
  XOR2_X1 U8034 ( .A(n8079), .B(n8078), .Z(n8122) );
  OR2_X1 U8035 ( .A1(n8123), .A2(n7664), .ZN(n8078) );
  OR2_X1 U8036 ( .A1(n8124), .A2(n8125), .ZN(n8079) );
  AND2_X1 U8037 ( .A1(n8126), .A2(n8127), .ZN(n8125) );
  AND2_X1 U8038 ( .A1(n8128), .A2(n8129), .ZN(n8124) );
  OR2_X1 U8039 ( .A1(n8127), .A2(n8126), .ZN(n8129) );
  XOR2_X1 U8040 ( .A(n8088), .B(n8130), .Z(n8080) );
  XOR2_X1 U8041 ( .A(n8087), .B(n8086), .Z(n8130) );
  OR2_X1 U8042 ( .A1(n8083), .A2(n7608), .ZN(n8086) );
  OR2_X1 U8043 ( .A1(n8131), .A2(n8132), .ZN(n8087) );
  AND2_X1 U8044 ( .A1(n8133), .A2(n8134), .ZN(n8132) );
  AND2_X1 U8045 ( .A1(n8135), .A2(n8136), .ZN(n8131) );
  OR2_X1 U8046 ( .A1(n8134), .A2(n8133), .ZN(n8136) );
  XOR2_X1 U8047 ( .A(n8095), .B(n8137), .Z(n8088) );
  XOR2_X1 U8048 ( .A(n8094), .B(n8093), .Z(n8137) );
  OR2_X1 U8049 ( .A1(n8041), .A2(n7610), .ZN(n8093) );
  OR2_X1 U8050 ( .A1(n8138), .A2(n8139), .ZN(n8094) );
  AND2_X1 U8051 ( .A1(n8140), .A2(n8141), .ZN(n8139) );
  AND2_X1 U8052 ( .A1(n8142), .A2(n8143), .ZN(n8138) );
  OR2_X1 U8053 ( .A1(n8141), .A2(n8140), .ZN(n8143) );
  XOR2_X1 U8054 ( .A(n8102), .B(n8144), .Z(n8095) );
  XOR2_X1 U8055 ( .A(n8101), .B(n8100), .Z(n8144) );
  OR2_X1 U8056 ( .A1(n8015), .A2(n7612), .ZN(n8100) );
  OR2_X1 U8057 ( .A1(n8145), .A2(n8146), .ZN(n8101) );
  AND2_X1 U8058 ( .A1(n8147), .A2(n8148), .ZN(n8146) );
  AND2_X1 U8059 ( .A1(n8149), .A2(n8150), .ZN(n8145) );
  OR2_X1 U8060 ( .A1(n8148), .A2(n8147), .ZN(n8150) );
  XOR2_X1 U8061 ( .A(n8110), .B(n8151), .Z(n8102) );
  XOR2_X1 U8062 ( .A(n8109), .B(n8108), .Z(n8151) );
  OR2_X1 U8063 ( .A1(n7988), .A2(n7614), .ZN(n8108) );
  OR2_X1 U8064 ( .A1(n8153), .A2(n8154), .ZN(n8109) );
  AND2_X1 U8065 ( .A1(n8155), .A2(n8156), .ZN(n8154) );
  AND2_X1 U8066 ( .A1(n8157), .A2(n8158), .ZN(n8153) );
  OR2_X1 U8067 ( .A1(n8156), .A2(n8155), .ZN(n8158) );
  XOR2_X1 U8068 ( .A(n8159), .B(n8160), .Z(n8110) );
  XOR2_X1 U8069 ( .A(n8161), .B(n8162), .Z(n8160) );
  OR2_X1 U8070 ( .A1(n8163), .A2(n8164), .ZN(n7677) );
  OR2_X1 U8071 ( .A1(n8165), .A2(n7676), .ZN(n8163) );
  AND3_X1 U8072 ( .A1(n7675), .A2(n7674), .A3(n7672), .ZN(n7676) );
  INV_X1 U8073 ( .A(n8166), .ZN(n7674) );
  AND2_X1 U8074 ( .A1(n7672), .A2(n7668), .ZN(n8165) );
  OR2_X1 U8075 ( .A1(n8167), .A2(n8168), .ZN(n7668) );
  AND2_X1 U8076 ( .A1(n7954), .A2(n7953), .ZN(n8168) );
  INV_X1 U8077 ( .A(n8169), .ZN(n7954) );
  AND2_X1 U8078 ( .A1(n7953), .A2(n7955), .ZN(n8167) );
  OR2_X1 U8079 ( .A1(n8170), .A2(n8171), .ZN(n7955) );
  AND2_X1 U8080 ( .A1(n8172), .A2(n7951), .ZN(n8171) );
  INV_X1 U8081 ( .A(n7949), .ZN(n8172) );
  AND2_X1 U8082 ( .A1(n7951), .A2(n7950), .ZN(n8170) );
  OR2_X1 U8083 ( .A1(n8173), .A2(n8174), .ZN(n7950) );
  AND2_X1 U8084 ( .A1(n8175), .A2(n7947), .ZN(n8174) );
  AND2_X1 U8085 ( .A1(n7947), .A2(n7946), .ZN(n8173) );
  OR2_X1 U8086 ( .A1(n8176), .A2(n8177), .ZN(n7946) );
  AND2_X1 U8087 ( .A1(n7941), .A2(n8178), .ZN(n8177) );
  INV_X1 U8088 ( .A(n8179), .ZN(n7941) );
  AND2_X1 U8089 ( .A1(n8178), .A2(n7942), .ZN(n8176) );
  OR2_X1 U8090 ( .A1(n8180), .A2(n8181), .ZN(n7942) );
  AND2_X1 U8091 ( .A1(n7937), .A2(n7939), .ZN(n8181) );
  AND2_X1 U8092 ( .A1(n7939), .A2(n8182), .ZN(n8180) );
  INV_X1 U8093 ( .A(n7938), .ZN(n8182) );
  AND2_X1 U8094 ( .A1(n7933), .A2(n8183), .ZN(n7938) );
  OR2_X1 U8095 ( .A1(n7931), .A2(n7935), .ZN(n8183) );
  AND2_X1 U8096 ( .A1(n8184), .A2(n8185), .ZN(n7935) );
  AND2_X1 U8097 ( .A1(n8186), .A2(n7928), .ZN(n7931) );
  OR3_X1 U8098 ( .A1(n8187), .A2(n8188), .A3(n8189), .ZN(n7928) );
  OR2_X1 U8099 ( .A1(n7926), .A2(n7930), .ZN(n8186) );
  AND2_X1 U8100 ( .A1(n8190), .A2(n8188), .ZN(n7930) );
  XNOR2_X1 U8101 ( .A(n8191), .B(n8192), .ZN(n8188) );
  OR2_X1 U8102 ( .A1(n8189), .A2(n8187), .ZN(n8190) );
  AND2_X1 U8103 ( .A1(n8193), .A2(n7923), .ZN(n7926) );
  OR3_X1 U8104 ( .A1(n8194), .A2(n8195), .A3(n8196), .ZN(n7923) );
  OR2_X1 U8105 ( .A1(n7921), .A2(n7925), .ZN(n8193) );
  AND2_X1 U8106 ( .A1(n8197), .A2(n8195), .ZN(n7925) );
  XNOR2_X1 U8107 ( .A(n8187), .B(n8189), .ZN(n8195) );
  OR2_X1 U8108 ( .A1(n8198), .A2(n8199), .ZN(n8189) );
  AND2_X1 U8109 ( .A1(n8200), .A2(n8201), .ZN(n8199) );
  AND2_X1 U8110 ( .A1(n8202), .A2(n8203), .ZN(n8198) );
  OR2_X1 U8111 ( .A1(n8200), .A2(n8201), .ZN(n8203) );
  XNOR2_X1 U8112 ( .A(n8204), .B(n8205), .ZN(n8187) );
  XNOR2_X1 U8113 ( .A(n8206), .B(n8207), .ZN(n8204) );
  OR2_X1 U8114 ( .A1(n8196), .A2(n8194), .ZN(n8197) );
  AND2_X1 U8115 ( .A1(n8208), .A2(n7920), .ZN(n7921) );
  OR3_X1 U8116 ( .A1(n8209), .A2(n8210), .A3(n8211), .ZN(n7920) );
  OR2_X1 U8117 ( .A1(n7917), .A2(n7918), .ZN(n8208) );
  AND2_X1 U8118 ( .A1(n8212), .A2(n8210), .ZN(n7918) );
  XNOR2_X1 U8119 ( .A(n8194), .B(n8196), .ZN(n8210) );
  OR2_X1 U8120 ( .A1(n8213), .A2(n8214), .ZN(n8196) );
  AND2_X1 U8121 ( .A1(n8215), .A2(n8216), .ZN(n8214) );
  AND2_X1 U8122 ( .A1(n8217), .A2(n8218), .ZN(n8213) );
  OR2_X1 U8123 ( .A1(n8215), .A2(n8216), .ZN(n8218) );
  XOR2_X1 U8124 ( .A(n8202), .B(n8219), .Z(n8194) );
  XOR2_X1 U8125 ( .A(n8201), .B(n8200), .Z(n8219) );
  OR2_X1 U8126 ( .A1(n8220), .A2(n7664), .ZN(n8200) );
  OR2_X1 U8127 ( .A1(n8221), .A2(n8222), .ZN(n8201) );
  AND2_X1 U8128 ( .A1(n8223), .A2(n8224), .ZN(n8222) );
  AND2_X1 U8129 ( .A1(n8225), .A2(n8226), .ZN(n8221) );
  OR2_X1 U8130 ( .A1(n8223), .A2(n8224), .ZN(n8226) );
  XNOR2_X1 U8131 ( .A(n8227), .B(n8228), .ZN(n8202) );
  XNOR2_X1 U8132 ( .A(n8229), .B(n8230), .ZN(n8227) );
  OR2_X1 U8133 ( .A1(n8211), .A2(n8209), .ZN(n8212) );
  AND2_X1 U8134 ( .A1(n8231), .A2(n7915), .ZN(n7917) );
  OR3_X1 U8135 ( .A1(n8232), .A2(n8233), .A3(n8234), .ZN(n7915) );
  OR2_X1 U8136 ( .A1(n7912), .A2(n7913), .ZN(n8231) );
  AND2_X1 U8137 ( .A1(n8235), .A2(n8233), .ZN(n7913) );
  XNOR2_X1 U8138 ( .A(n8209), .B(n8211), .ZN(n8233) );
  OR2_X1 U8139 ( .A1(n8236), .A2(n8237), .ZN(n8211) );
  AND2_X1 U8140 ( .A1(n8238), .A2(n8239), .ZN(n8237) );
  AND2_X1 U8141 ( .A1(n8240), .A2(n8241), .ZN(n8236) );
  OR2_X1 U8142 ( .A1(n8238), .A2(n8239), .ZN(n8241) );
  XOR2_X1 U8143 ( .A(n8217), .B(n8242), .Z(n8209) );
  XOR2_X1 U8144 ( .A(n8216), .B(n8215), .Z(n8242) );
  OR2_X1 U8145 ( .A1(n8243), .A2(n7664), .ZN(n8215) );
  OR2_X1 U8146 ( .A1(n8244), .A2(n8245), .ZN(n8216) );
  AND2_X1 U8147 ( .A1(n8246), .A2(n8247), .ZN(n8245) );
  AND2_X1 U8148 ( .A1(n8248), .A2(n8249), .ZN(n8244) );
  OR2_X1 U8149 ( .A1(n8246), .A2(n8247), .ZN(n8249) );
  XOR2_X1 U8150 ( .A(n8225), .B(n8250), .Z(n8217) );
  XOR2_X1 U8151 ( .A(n8224), .B(n8223), .Z(n8250) );
  OR2_X1 U8152 ( .A1(n7608), .A2(n8220), .ZN(n8223) );
  OR2_X1 U8153 ( .A1(n8251), .A2(n8252), .ZN(n8224) );
  AND2_X1 U8154 ( .A1(n8253), .A2(n8254), .ZN(n8252) );
  AND2_X1 U8155 ( .A1(n8255), .A2(n8256), .ZN(n8251) );
  OR2_X1 U8156 ( .A1(n8253), .A2(n8254), .ZN(n8256) );
  XOR2_X1 U8157 ( .A(n8257), .B(n8258), .Z(n8225) );
  XOR2_X1 U8158 ( .A(n8259), .B(n8260), .Z(n8258) );
  OR2_X1 U8159 ( .A1(n8234), .A2(n8232), .ZN(n8235) );
  AND2_X1 U8160 ( .A1(n8261), .A2(n7901), .ZN(n7912) );
  OR3_X1 U8161 ( .A1(n8262), .A2(n8263), .A3(n8264), .ZN(n7901) );
  OR2_X1 U8162 ( .A1(n7898), .A2(n7899), .ZN(n8261) );
  AND2_X1 U8163 ( .A1(n8265), .A2(n8263), .ZN(n7899) );
  XNOR2_X1 U8164 ( .A(n8232), .B(n8234), .ZN(n8263) );
  OR2_X1 U8165 ( .A1(n8266), .A2(n8267), .ZN(n8234) );
  AND2_X1 U8166 ( .A1(n8268), .A2(n8269), .ZN(n8267) );
  AND2_X1 U8167 ( .A1(n8270), .A2(n8271), .ZN(n8266) );
  OR2_X1 U8168 ( .A1(n8268), .A2(n8269), .ZN(n8271) );
  XOR2_X1 U8169 ( .A(n8240), .B(n8272), .Z(n8232) );
  XOR2_X1 U8170 ( .A(n8239), .B(n8238), .Z(n8272) );
  OR2_X1 U8171 ( .A1(n8273), .A2(n7664), .ZN(n8238) );
  OR2_X1 U8172 ( .A1(n8274), .A2(n8275), .ZN(n8239) );
  AND2_X1 U8173 ( .A1(n8276), .A2(n8277), .ZN(n8275) );
  AND2_X1 U8174 ( .A1(n8278), .A2(n8279), .ZN(n8274) );
  OR2_X1 U8175 ( .A1(n8276), .A2(n8277), .ZN(n8279) );
  XOR2_X1 U8176 ( .A(n8248), .B(n8280), .Z(n8240) );
  XOR2_X1 U8177 ( .A(n8247), .B(n8246), .Z(n8280) );
  OR2_X1 U8178 ( .A1(n7608), .A2(n8243), .ZN(n8246) );
  OR2_X1 U8179 ( .A1(n8281), .A2(n8282), .ZN(n8247) );
  AND2_X1 U8180 ( .A1(n8283), .A2(n8284), .ZN(n8282) );
  AND2_X1 U8181 ( .A1(n8285), .A2(n8286), .ZN(n8281) );
  OR2_X1 U8182 ( .A1(n8283), .A2(n8284), .ZN(n8286) );
  XOR2_X1 U8183 ( .A(n8255), .B(n8287), .Z(n8248) );
  XOR2_X1 U8184 ( .A(n8254), .B(n8253), .Z(n8287) );
  OR2_X1 U8185 ( .A1(n7610), .A2(n8220), .ZN(n8253) );
  OR2_X1 U8186 ( .A1(n8288), .A2(n8289), .ZN(n8254) );
  AND2_X1 U8187 ( .A1(n8290), .A2(n8291), .ZN(n8289) );
  AND2_X1 U8188 ( .A1(n8292), .A2(n8293), .ZN(n8288) );
  OR2_X1 U8189 ( .A1(n8290), .A2(n8291), .ZN(n8293) );
  XOR2_X1 U8190 ( .A(n8294), .B(n8295), .Z(n8255) );
  XOR2_X1 U8191 ( .A(n8296), .B(n8297), .Z(n8295) );
  OR2_X1 U8192 ( .A1(n8264), .A2(n8262), .ZN(n8265) );
  AND2_X1 U8193 ( .A1(n8298), .A2(n8299), .ZN(n7898) );
  INV_X1 U8194 ( .A(n7896), .ZN(n8299) );
  AND3_X1 U8195 ( .A1(n8300), .A2(n8301), .A3(n8302), .ZN(n7896) );
  OR2_X1 U8196 ( .A1(n7895), .A2(n7894), .ZN(n8298) );
  AND2_X1 U8197 ( .A1(n8303), .A2(n7892), .ZN(n7894) );
  OR3_X1 U8198 ( .A1(n8304), .A2(n8305), .A3(n8306), .ZN(n7892) );
  OR2_X1 U8199 ( .A1(n7889), .A2(n7890), .ZN(n8303) );
  AND2_X1 U8200 ( .A1(n8307), .A2(n8305), .ZN(n7890) );
  XNOR2_X1 U8201 ( .A(n8300), .B(n8302), .ZN(n8305) );
  OR2_X1 U8202 ( .A1(n8306), .A2(n8304), .ZN(n8307) );
  AND2_X1 U8203 ( .A1(n8308), .A2(n7887), .ZN(n7889) );
  OR3_X1 U8204 ( .A1(n8309), .A2(n8310), .A3(n8311), .ZN(n7887) );
  OR2_X1 U8205 ( .A1(n7884), .A2(n7885), .ZN(n8308) );
  AND2_X1 U8206 ( .A1(n8312), .A2(n8310), .ZN(n7885) );
  XNOR2_X1 U8207 ( .A(n8304), .B(n8306), .ZN(n8310) );
  OR2_X1 U8208 ( .A1(n8313), .A2(n8314), .ZN(n8306) );
  AND2_X1 U8209 ( .A1(n8315), .A2(n8316), .ZN(n8314) );
  AND2_X1 U8210 ( .A1(n8317), .A2(n8318), .ZN(n8313) );
  OR2_X1 U8211 ( .A1(n8315), .A2(n8316), .ZN(n8318) );
  XOR2_X1 U8212 ( .A(n8319), .B(n8320), .Z(n8304) );
  XOR2_X1 U8213 ( .A(n8321), .B(n8322), .Z(n8320) );
  OR2_X1 U8214 ( .A1(n8311), .A2(n8309), .ZN(n8312) );
  AND2_X1 U8215 ( .A1(n8323), .A2(n7882), .ZN(n7884) );
  OR3_X1 U8216 ( .A1(n8324), .A2(n8325), .A3(n8326), .ZN(n7882) );
  OR2_X1 U8217 ( .A1(n7879), .A2(n7880), .ZN(n8323) );
  AND2_X1 U8218 ( .A1(n8327), .A2(n8325), .ZN(n7880) );
  XNOR2_X1 U8219 ( .A(n8309), .B(n8311), .ZN(n8325) );
  OR2_X1 U8220 ( .A1(n8328), .A2(n8329), .ZN(n8311) );
  AND2_X1 U8221 ( .A1(n8330), .A2(n8331), .ZN(n8329) );
  AND2_X1 U8222 ( .A1(n8332), .A2(n8333), .ZN(n8328) );
  OR2_X1 U8223 ( .A1(n8330), .A2(n8331), .ZN(n8333) );
  XOR2_X1 U8224 ( .A(n8317), .B(n8334), .Z(n8309) );
  XOR2_X1 U8225 ( .A(n8316), .B(n8315), .Z(n8334) );
  OR2_X1 U8226 ( .A1(n8335), .A2(n7664), .ZN(n8315) );
  OR2_X1 U8227 ( .A1(n8336), .A2(n8337), .ZN(n8316) );
  AND2_X1 U8228 ( .A1(n8338), .A2(n8339), .ZN(n8337) );
  AND2_X1 U8229 ( .A1(n8340), .A2(n8341), .ZN(n8336) );
  OR2_X1 U8230 ( .A1(n8338), .A2(n8339), .ZN(n8341) );
  XOR2_X1 U8231 ( .A(n8342), .B(n8343), .Z(n8317) );
  XOR2_X1 U8232 ( .A(n8344), .B(n8345), .Z(n8343) );
  OR2_X1 U8233 ( .A1(n8326), .A2(n8324), .ZN(n8327) );
  AND2_X1 U8234 ( .A1(n8346), .A2(n7877), .ZN(n7879) );
  OR3_X1 U8235 ( .A1(n8347), .A2(n8348), .A3(n8349), .ZN(n7877) );
  OR2_X1 U8236 ( .A1(n7874), .A2(n7875), .ZN(n8346) );
  AND2_X1 U8237 ( .A1(n8350), .A2(n8348), .ZN(n7875) );
  XNOR2_X1 U8238 ( .A(n8324), .B(n8326), .ZN(n8348) );
  OR2_X1 U8239 ( .A1(n8351), .A2(n8352), .ZN(n8326) );
  AND2_X1 U8240 ( .A1(n8353), .A2(n8354), .ZN(n8352) );
  AND2_X1 U8241 ( .A1(n8355), .A2(n8356), .ZN(n8351) );
  OR2_X1 U8242 ( .A1(n8353), .A2(n8354), .ZN(n8356) );
  XOR2_X1 U8243 ( .A(n8332), .B(n8357), .Z(n8324) );
  XOR2_X1 U8244 ( .A(n8331), .B(n8330), .Z(n8357) );
  OR2_X1 U8245 ( .A1(n8358), .A2(n7664), .ZN(n8330) );
  OR2_X1 U8246 ( .A1(n8359), .A2(n8360), .ZN(n8331) );
  AND2_X1 U8247 ( .A1(n8361), .A2(n8362), .ZN(n8360) );
  AND2_X1 U8248 ( .A1(n8363), .A2(n8364), .ZN(n8359) );
  OR2_X1 U8249 ( .A1(n8361), .A2(n8362), .ZN(n8364) );
  XOR2_X1 U8250 ( .A(n8340), .B(n8365), .Z(n8332) );
  XOR2_X1 U8251 ( .A(n8339), .B(n8338), .Z(n8365) );
  OR2_X1 U8252 ( .A1(n7608), .A2(n8335), .ZN(n8338) );
  OR2_X1 U8253 ( .A1(n8366), .A2(n8367), .ZN(n8339) );
  AND2_X1 U8254 ( .A1(n8368), .A2(n8369), .ZN(n8367) );
  AND2_X1 U8255 ( .A1(n8370), .A2(n8371), .ZN(n8366) );
  OR2_X1 U8256 ( .A1(n8368), .A2(n8369), .ZN(n8371) );
  XOR2_X1 U8257 ( .A(n8372), .B(n8373), .Z(n8340) );
  XOR2_X1 U8258 ( .A(n8374), .B(n8375), .Z(n8373) );
  OR2_X1 U8259 ( .A1(n8349), .A2(n8347), .ZN(n8350) );
  AND2_X1 U8260 ( .A1(n8376), .A2(n7872), .ZN(n7874) );
  OR2_X1 U8261 ( .A1(n8377), .A2(n8378), .ZN(n7872) );
  OR2_X1 U8262 ( .A1(n7871), .A2(n7869), .ZN(n8376) );
  AND2_X1 U8263 ( .A1(n8379), .A2(n7867), .ZN(n7869) );
  OR2_X1 U8264 ( .A1(n8380), .A2(n8381), .ZN(n7867) );
  OR2_X1 U8265 ( .A1(n7864), .A2(n7865), .ZN(n8379) );
  AND2_X1 U8266 ( .A1(n8381), .A2(n8380), .ZN(n7865) );
  OR2_X1 U8267 ( .A1(n8382), .A2(n8383), .ZN(n8380) );
  INV_X1 U8268 ( .A(n8378), .ZN(n8383) );
  AND2_X1 U8269 ( .A1(n8384), .A2(n8385), .ZN(n8382) );
  OR2_X1 U8270 ( .A1(n8386), .A2(n8387), .ZN(n8381) );
  AND2_X1 U8271 ( .A1(n8388), .A2(n7862), .ZN(n7864) );
  OR2_X1 U8272 ( .A1(n8389), .A2(n8390), .ZN(n7862) );
  OR2_X1 U8273 ( .A1(n7859), .A2(n7860), .ZN(n8388) );
  AND2_X1 U8274 ( .A1(n8390), .A2(n8389), .ZN(n7860) );
  XNOR2_X1 U8275 ( .A(n8386), .B(n8387), .ZN(n8389) );
  OR2_X1 U8276 ( .A1(n8391), .A2(n8392), .ZN(n8387) );
  AND2_X1 U8277 ( .A1(n8393), .A2(n8394), .ZN(n8392) );
  AND2_X1 U8278 ( .A1(n8395), .A2(n8396), .ZN(n8391) );
  OR2_X1 U8279 ( .A1(n8393), .A2(n8394), .ZN(n8396) );
  XOR2_X1 U8280 ( .A(n8397), .B(n8398), .Z(n8386) );
  XOR2_X1 U8281 ( .A(n8399), .B(n8400), .Z(n8398) );
  AND2_X1 U8282 ( .A1(n8401), .A2(n7857), .ZN(n7859) );
  OR2_X1 U8283 ( .A1(n8402), .A2(n8403), .ZN(n7857) );
  OR2_X1 U8284 ( .A1(n7847), .A2(n7855), .ZN(n8401) );
  AND2_X1 U8285 ( .A1(n8403), .A2(n8402), .ZN(n7855) );
  OR2_X1 U8286 ( .A1(n8404), .A2(n8405), .ZN(n8402) );
  OR2_X1 U8287 ( .A1(n8406), .A2(n8407), .ZN(n8403) );
  INV_X1 U8288 ( .A(n8390), .ZN(n8407) );
  OR2_X1 U8289 ( .A1(n8408), .A2(n8409), .ZN(n8390) );
  AND2_X1 U8290 ( .A1(n8408), .A2(n8409), .ZN(n8406) );
  OR2_X1 U8291 ( .A1(n8410), .A2(n8411), .ZN(n8409) );
  AND2_X1 U8292 ( .A1(n8412), .A2(n8413), .ZN(n8411) );
  AND2_X1 U8293 ( .A1(n8414), .A2(n8415), .ZN(n8410) );
  OR2_X1 U8294 ( .A1(n8412), .A2(n8413), .ZN(n8415) );
  XOR2_X1 U8295 ( .A(n8395), .B(n8416), .Z(n8408) );
  XOR2_X1 U8296 ( .A(n8394), .B(n8393), .Z(n8416) );
  OR2_X1 U8297 ( .A1(n8417), .A2(n7664), .ZN(n8393) );
  OR2_X1 U8298 ( .A1(n8418), .A2(n8419), .ZN(n8394) );
  AND2_X1 U8299 ( .A1(n8420), .A2(n8421), .ZN(n8419) );
  AND2_X1 U8300 ( .A1(n8422), .A2(n8423), .ZN(n8418) );
  OR2_X1 U8301 ( .A1(n8420), .A2(n8421), .ZN(n8423) );
  XOR2_X1 U8302 ( .A(n8424), .B(n8425), .Z(n8395) );
  XOR2_X1 U8303 ( .A(n8426), .B(n8427), .Z(n8425) );
  INV_X1 U8304 ( .A(n7853), .ZN(n7847) );
  AND3_X1 U8305 ( .A1(n7845), .A2(n7849), .A3(n7850), .ZN(n7853) );
  INV_X1 U8306 ( .A(n7844), .ZN(n7850) );
  OR2_X1 U8307 ( .A1(n8428), .A2(n8429), .ZN(n7844) );
  AND2_X1 U8308 ( .A1(n7843), .A2(n7842), .ZN(n8429) );
  AND2_X1 U8309 ( .A1(n7840), .A2(n8430), .ZN(n8428) );
  OR2_X1 U8310 ( .A1(n7843), .A2(n7842), .ZN(n8430) );
  OR2_X1 U8311 ( .A1(n8431), .A2(n8432), .ZN(n7842) );
  AND2_X1 U8312 ( .A1(n7839), .A2(n7838), .ZN(n8432) );
  AND2_X1 U8313 ( .A1(n7836), .A2(n8433), .ZN(n8431) );
  OR2_X1 U8314 ( .A1(n7839), .A2(n7838), .ZN(n8433) );
  OR2_X1 U8315 ( .A1(n8434), .A2(n8435), .ZN(n7838) );
  AND2_X1 U8316 ( .A1(n7835), .A2(n7834), .ZN(n8435) );
  AND2_X1 U8317 ( .A1(n7832), .A2(n8436), .ZN(n8434) );
  OR2_X1 U8318 ( .A1(n7835), .A2(n7834), .ZN(n8436) );
  OR2_X1 U8319 ( .A1(n8437), .A2(n8438), .ZN(n7834) );
  AND2_X1 U8320 ( .A1(n7831), .A2(n7830), .ZN(n8438) );
  AND2_X1 U8321 ( .A1(n7828), .A2(n8439), .ZN(n8437) );
  OR2_X1 U8322 ( .A1(n7831), .A2(n7830), .ZN(n8439) );
  OR2_X1 U8323 ( .A1(n8440), .A2(n8441), .ZN(n7830) );
  AND2_X1 U8324 ( .A1(n7827), .A2(n7826), .ZN(n8441) );
  AND2_X1 U8325 ( .A1(n7824), .A2(n8442), .ZN(n8440) );
  OR2_X1 U8326 ( .A1(n7827), .A2(n7826), .ZN(n8442) );
  OR2_X1 U8327 ( .A1(n8443), .A2(n8444), .ZN(n7826) );
  AND2_X1 U8328 ( .A1(n7823), .A2(n7822), .ZN(n8444) );
  AND2_X1 U8329 ( .A1(n7820), .A2(n8445), .ZN(n8443) );
  OR2_X1 U8330 ( .A1(n7823), .A2(n7822), .ZN(n8445) );
  OR2_X1 U8331 ( .A1(n8446), .A2(n8447), .ZN(n7822) );
  AND2_X1 U8332 ( .A1(n7819), .A2(n7818), .ZN(n8447) );
  AND2_X1 U8333 ( .A1(n7816), .A2(n8448), .ZN(n8446) );
  OR2_X1 U8334 ( .A1(n7819), .A2(n7818), .ZN(n8448) );
  OR2_X1 U8335 ( .A1(n8449), .A2(n8450), .ZN(n7818) );
  AND2_X1 U8336 ( .A1(n7815), .A2(n7814), .ZN(n8450) );
  AND2_X1 U8337 ( .A1(n7812), .A2(n8451), .ZN(n8449) );
  OR2_X1 U8338 ( .A1(n7815), .A2(n7814), .ZN(n8451) );
  OR2_X1 U8339 ( .A1(n8452), .A2(n8453), .ZN(n7814) );
  AND2_X1 U8340 ( .A1(n7802), .A2(n7801), .ZN(n8453) );
  AND2_X1 U8341 ( .A1(n7799), .A2(n8454), .ZN(n8452) );
  OR2_X1 U8342 ( .A1(n7802), .A2(n7801), .ZN(n8454) );
  OR2_X1 U8343 ( .A1(n8455), .A2(n8456), .ZN(n7801) );
  AND2_X1 U8344 ( .A1(n7798), .A2(n7797), .ZN(n8456) );
  AND2_X1 U8345 ( .A1(n7795), .A2(n8457), .ZN(n8455) );
  OR2_X1 U8346 ( .A1(n7798), .A2(n7797), .ZN(n8457) );
  OR2_X1 U8347 ( .A1(n8458), .A2(n8459), .ZN(n7797) );
  AND2_X1 U8348 ( .A1(n7794), .A2(n7793), .ZN(n8459) );
  AND2_X1 U8349 ( .A1(n7791), .A2(n8460), .ZN(n8458) );
  OR2_X1 U8350 ( .A1(n7794), .A2(n7793), .ZN(n8460) );
  OR2_X1 U8351 ( .A1(n8461), .A2(n8462), .ZN(n7793) );
  AND2_X1 U8352 ( .A1(n7790), .A2(n7789), .ZN(n8462) );
  AND2_X1 U8353 ( .A1(n7787), .A2(n8463), .ZN(n8461) );
  OR2_X1 U8354 ( .A1(n7790), .A2(n7789), .ZN(n8463) );
  OR2_X1 U8355 ( .A1(n8464), .A2(n8465), .ZN(n7789) );
  AND2_X1 U8356 ( .A1(n7786), .A2(n7785), .ZN(n8465) );
  AND2_X1 U8357 ( .A1(n7783), .A2(n8466), .ZN(n8464) );
  OR2_X1 U8358 ( .A1(n7786), .A2(n7785), .ZN(n8466) );
  OR2_X1 U8359 ( .A1(n8467), .A2(n8468), .ZN(n7785) );
  AND2_X1 U8360 ( .A1(n7782), .A2(n7781), .ZN(n8468) );
  AND2_X1 U8361 ( .A1(n7779), .A2(n8469), .ZN(n8467) );
  OR2_X1 U8362 ( .A1(n7782), .A2(n7781), .ZN(n8469) );
  OR2_X1 U8363 ( .A1(n8470), .A2(n8471), .ZN(n7781) );
  AND2_X1 U8364 ( .A1(n7778), .A2(n7777), .ZN(n8471) );
  AND2_X1 U8365 ( .A1(n7775), .A2(n8472), .ZN(n8470) );
  OR2_X1 U8366 ( .A1(n7778), .A2(n7777), .ZN(n8472) );
  OR2_X1 U8367 ( .A1(n8473), .A2(n8474), .ZN(n7777) );
  AND2_X1 U8368 ( .A1(n7774), .A2(n7773), .ZN(n8474) );
  AND2_X1 U8369 ( .A1(n7771), .A2(n8475), .ZN(n8473) );
  OR2_X1 U8370 ( .A1(n7774), .A2(n7773), .ZN(n8475) );
  OR2_X1 U8371 ( .A1(n8476), .A2(n8477), .ZN(n7773) );
  AND2_X1 U8372 ( .A1(n7770), .A2(n7769), .ZN(n8477) );
  AND2_X1 U8373 ( .A1(n7767), .A2(n8478), .ZN(n8476) );
  OR2_X1 U8374 ( .A1(n7770), .A2(n7769), .ZN(n8478) );
  OR2_X1 U8375 ( .A1(n8479), .A2(n8480), .ZN(n7769) );
  AND2_X1 U8376 ( .A1(n7766), .A2(n7765), .ZN(n8480) );
  AND2_X1 U8377 ( .A1(n7763), .A2(n8481), .ZN(n8479) );
  OR2_X1 U8378 ( .A1(n7766), .A2(n7765), .ZN(n8481) );
  OR2_X1 U8379 ( .A1(n8482), .A2(n8483), .ZN(n7765) );
  AND2_X1 U8380 ( .A1(n7760), .A2(n7759), .ZN(n8483) );
  AND2_X1 U8381 ( .A1(n7757), .A2(n8484), .ZN(n8482) );
  OR2_X1 U8382 ( .A1(n7760), .A2(n7759), .ZN(n8484) );
  OR2_X1 U8383 ( .A1(n8485), .A2(n8486), .ZN(n7759) );
  AND2_X1 U8384 ( .A1(n7756), .A2(n7755), .ZN(n8486) );
  AND2_X1 U8385 ( .A1(n7753), .A2(n8487), .ZN(n8485) );
  OR2_X1 U8386 ( .A1(n7756), .A2(n7755), .ZN(n8487) );
  OR2_X1 U8387 ( .A1(n8488), .A2(n8489), .ZN(n7755) );
  AND2_X1 U8388 ( .A1(n7752), .A2(n7751), .ZN(n8489) );
  AND2_X1 U8389 ( .A1(n7749), .A2(n8490), .ZN(n8488) );
  OR2_X1 U8390 ( .A1(n7752), .A2(n7751), .ZN(n8490) );
  OR2_X1 U8391 ( .A1(n8491), .A2(n8492), .ZN(n7751) );
  AND2_X1 U8392 ( .A1(n7748), .A2(n7747), .ZN(n8492) );
  AND2_X1 U8393 ( .A1(n7745), .A2(n8493), .ZN(n8491) );
  OR2_X1 U8394 ( .A1(n7748), .A2(n7747), .ZN(n8493) );
  OR2_X1 U8395 ( .A1(n8494), .A2(n8495), .ZN(n7747) );
  AND2_X1 U8396 ( .A1(n7744), .A2(n7743), .ZN(n8495) );
  AND2_X1 U8397 ( .A1(n7741), .A2(n8496), .ZN(n8494) );
  OR2_X1 U8398 ( .A1(n7744), .A2(n7743), .ZN(n8496) );
  OR2_X1 U8399 ( .A1(n8497), .A2(n8498), .ZN(n7743) );
  AND2_X1 U8400 ( .A1(n7740), .A2(n7739), .ZN(n8498) );
  AND2_X1 U8401 ( .A1(n7737), .A2(n8499), .ZN(n8497) );
  OR2_X1 U8402 ( .A1(n7740), .A2(n7739), .ZN(n8499) );
  OR2_X1 U8403 ( .A1(n8500), .A2(n8501), .ZN(n7739) );
  AND2_X1 U8404 ( .A1(n7736), .A2(n7735), .ZN(n8501) );
  AND2_X1 U8405 ( .A1(n7733), .A2(n8502), .ZN(n8500) );
  OR2_X1 U8406 ( .A1(n7736), .A2(n7735), .ZN(n8502) );
  OR2_X1 U8407 ( .A1(n8503), .A2(n8504), .ZN(n7735) );
  AND2_X1 U8408 ( .A1(n7732), .A2(n7731), .ZN(n8504) );
  AND2_X1 U8409 ( .A1(n7729), .A2(n8505), .ZN(n8503) );
  OR2_X1 U8410 ( .A1(n7732), .A2(n7731), .ZN(n8505) );
  OR2_X1 U8411 ( .A1(n8506), .A2(n8507), .ZN(n7731) );
  AND2_X1 U8412 ( .A1(n7728), .A2(n7727), .ZN(n8507) );
  AND2_X1 U8413 ( .A1(n7725), .A2(n8508), .ZN(n8506) );
  OR2_X1 U8414 ( .A1(n7728), .A2(n7727), .ZN(n8508) );
  OR2_X1 U8415 ( .A1(n8509), .A2(n8510), .ZN(n7727) );
  AND2_X1 U8416 ( .A1(n7724), .A2(n7723), .ZN(n8510) );
  AND2_X1 U8417 ( .A1(n7721), .A2(n8511), .ZN(n8509) );
  OR2_X1 U8418 ( .A1(n7724), .A2(n7723), .ZN(n8511) );
  OR2_X1 U8419 ( .A1(n8512), .A2(n8513), .ZN(n7723) );
  AND2_X1 U8420 ( .A1(n7711), .A2(n7710), .ZN(n8513) );
  AND2_X1 U8421 ( .A1(n7708), .A2(n8514), .ZN(n8512) );
  OR2_X1 U8422 ( .A1(n7711), .A2(n7710), .ZN(n8514) );
  OR2_X1 U8423 ( .A1(n8515), .A2(n8516), .ZN(n7710) );
  AND2_X1 U8424 ( .A1(n7704), .A2(n7707), .ZN(n8516) );
  AND2_X1 U8425 ( .A1(n7706), .A2(n8517), .ZN(n8515) );
  OR2_X1 U8426 ( .A1(n7704), .A2(n7707), .ZN(n8517) );
  OR2_X1 U8427 ( .A1(n8518), .A2(n7698), .ZN(n7707) );
  OR3_X1 U8428 ( .A1(n7702), .A2(n8519), .A3(n7698), .ZN(n7704) );
  INV_X1 U8429 ( .A(n8520), .ZN(n7706) );
  OR2_X1 U8430 ( .A1(n8521), .A2(n8522), .ZN(n8520) );
  AND2_X1 U8431 ( .A1(n8523), .A2(n8524), .ZN(n8522) );
  OR2_X1 U8432 ( .A1(n8525), .A2(n7697), .ZN(n8524) );
  AND2_X1 U8433 ( .A1(n7665), .A2(n7691), .ZN(n8525) );
  AND2_X1 U8434 ( .A1(n7694), .A2(n8526), .ZN(n8521) );
  OR2_X1 U8435 ( .A1(n8527), .A2(n7701), .ZN(n8526) );
  AND2_X1 U8436 ( .A1(n7667), .A2(n7703), .ZN(n8527) );
  INV_X1 U8437 ( .A(n7702), .ZN(n7694) );
  OR2_X1 U8438 ( .A1(n7662), .A2(n7698), .ZN(n7711) );
  XNOR2_X1 U8439 ( .A(n8530), .B(n8531), .ZN(n7708) );
  XNOR2_X1 U8440 ( .A(n8532), .B(n8533), .ZN(n8531) );
  OR2_X1 U8441 ( .A1(n7660), .A2(n7698), .ZN(n7724) );
  XOR2_X1 U8442 ( .A(n8535), .B(n8536), .Z(n7721) );
  XOR2_X1 U8443 ( .A(n8537), .B(n8538), .Z(n8536) );
  OR2_X1 U8444 ( .A1(n7658), .A2(n7698), .ZN(n7728) );
  XOR2_X1 U8445 ( .A(n8540), .B(n8541), .Z(n7725) );
  XOR2_X1 U8446 ( .A(n8542), .B(n8543), .Z(n8541) );
  OR2_X1 U8447 ( .A1(n7656), .A2(n7698), .ZN(n7732) );
  XOR2_X1 U8448 ( .A(n8545), .B(n8546), .Z(n7729) );
  XOR2_X1 U8449 ( .A(n8547), .B(n8548), .Z(n8546) );
  OR2_X1 U8450 ( .A1(n7654), .A2(n7698), .ZN(n7736) );
  XOR2_X1 U8451 ( .A(n8550), .B(n8551), .Z(n7733) );
  XOR2_X1 U8452 ( .A(n8552), .B(n8553), .Z(n8551) );
  OR2_X1 U8453 ( .A1(n7652), .A2(n7698), .ZN(n7740) );
  XOR2_X1 U8454 ( .A(n8555), .B(n8556), .Z(n7737) );
  XOR2_X1 U8455 ( .A(n8557), .B(n8558), .Z(n8556) );
  OR2_X1 U8456 ( .A1(n7650), .A2(n7698), .ZN(n7744) );
  XOR2_X1 U8457 ( .A(n8560), .B(n8561), .Z(n7741) );
  XOR2_X1 U8458 ( .A(n8562), .B(n8563), .Z(n8561) );
  OR2_X1 U8459 ( .A1(n7648), .A2(n7698), .ZN(n7748) );
  XOR2_X1 U8460 ( .A(n8565), .B(n8566), .Z(n7745) );
  XOR2_X1 U8461 ( .A(n8567), .B(n8568), .Z(n8566) );
  OR2_X1 U8462 ( .A1(n7646), .A2(n7698), .ZN(n7752) );
  XOR2_X1 U8463 ( .A(n8570), .B(n8571), .Z(n7749) );
  XOR2_X1 U8464 ( .A(n8572), .B(n8573), .Z(n8571) );
  OR2_X1 U8465 ( .A1(n7644), .A2(n7698), .ZN(n7756) );
  XOR2_X1 U8466 ( .A(n8575), .B(n8576), .Z(n7753) );
  XOR2_X1 U8467 ( .A(n8577), .B(n8578), .Z(n8576) );
  OR2_X1 U8468 ( .A1(n7642), .A2(n7698), .ZN(n7760) );
  XOR2_X1 U8469 ( .A(n8580), .B(n8581), .Z(n7757) );
  XOR2_X1 U8470 ( .A(n8582), .B(n8583), .Z(n8581) );
  OR2_X1 U8471 ( .A1(n7640), .A2(n7698), .ZN(n7766) );
  XOR2_X1 U8472 ( .A(n8585), .B(n8586), .Z(n7763) );
  XOR2_X1 U8473 ( .A(n8587), .B(n8588), .Z(n8586) );
  OR2_X1 U8474 ( .A1(n7638), .A2(n7698), .ZN(n7770) );
  XOR2_X1 U8475 ( .A(n8590), .B(n8591), .Z(n7767) );
  XOR2_X1 U8476 ( .A(n8592), .B(n8593), .Z(n8591) );
  OR2_X1 U8477 ( .A1(n7636), .A2(n7698), .ZN(n7774) );
  XOR2_X1 U8478 ( .A(n8595), .B(n8596), .Z(n7771) );
  XOR2_X1 U8479 ( .A(n8597), .B(n8598), .Z(n8596) );
  OR2_X1 U8480 ( .A1(n7634), .A2(n7698), .ZN(n7778) );
  XOR2_X1 U8481 ( .A(n8600), .B(n8601), .Z(n7775) );
  XOR2_X1 U8482 ( .A(n8602), .B(n8603), .Z(n8601) );
  OR2_X1 U8483 ( .A1(n7632), .A2(n7698), .ZN(n7782) );
  XOR2_X1 U8484 ( .A(n8605), .B(n8606), .Z(n7779) );
  XOR2_X1 U8485 ( .A(n8607), .B(n8608), .Z(n8606) );
  OR2_X1 U8486 ( .A1(n7630), .A2(n7698), .ZN(n7786) );
  XOR2_X1 U8487 ( .A(n8610), .B(n8611), .Z(n7783) );
  XOR2_X1 U8488 ( .A(n8612), .B(n8613), .Z(n8611) );
  OR2_X1 U8489 ( .A1(n7628), .A2(n7698), .ZN(n7790) );
  XOR2_X1 U8490 ( .A(n8615), .B(n8616), .Z(n7787) );
  XOR2_X1 U8491 ( .A(n8617), .B(n8618), .Z(n8616) );
  OR2_X1 U8492 ( .A1(n7626), .A2(n7698), .ZN(n7794) );
  XOR2_X1 U8493 ( .A(n8620), .B(n8621), .Z(n7791) );
  XOR2_X1 U8494 ( .A(n8622), .B(n8623), .Z(n8621) );
  OR2_X1 U8495 ( .A1(n7624), .A2(n7698), .ZN(n7798) );
  XOR2_X1 U8496 ( .A(n8625), .B(n8626), .Z(n7795) );
  XOR2_X1 U8497 ( .A(n8627), .B(n8628), .Z(n8626) );
  OR2_X1 U8498 ( .A1(n7622), .A2(n7698), .ZN(n7802) );
  XOR2_X1 U8499 ( .A(n8630), .B(n8631), .Z(n7799) );
  XOR2_X1 U8500 ( .A(n8632), .B(n8633), .Z(n8631) );
  OR2_X1 U8501 ( .A1(n7620), .A2(n7698), .ZN(n7815) );
  XOR2_X1 U8502 ( .A(n8635), .B(n8636), .Z(n7812) );
  XOR2_X1 U8503 ( .A(n8637), .B(n8638), .Z(n8636) );
  OR2_X1 U8504 ( .A1(n7618), .A2(n7698), .ZN(n7819) );
  XOR2_X1 U8505 ( .A(n8640), .B(n8641), .Z(n7816) );
  XOR2_X1 U8506 ( .A(n8642), .B(n8643), .Z(n8641) );
  OR2_X1 U8507 ( .A1(n7616), .A2(n7698), .ZN(n7823) );
  XOR2_X1 U8508 ( .A(n8645), .B(n8646), .Z(n7820) );
  XOR2_X1 U8509 ( .A(n8647), .B(n8648), .Z(n8646) );
  OR2_X1 U8510 ( .A1(n7614), .A2(n7698), .ZN(n7827) );
  XOR2_X1 U8511 ( .A(n8649), .B(n8650), .Z(n7824) );
  XOR2_X1 U8512 ( .A(n8651), .B(n8652), .Z(n8650) );
  OR2_X1 U8513 ( .A1(n7612), .A2(n7698), .ZN(n7831) );
  XOR2_X1 U8514 ( .A(n8653), .B(n8654), .Z(n7828) );
  XOR2_X1 U8515 ( .A(n8655), .B(n8656), .Z(n8654) );
  OR2_X1 U8516 ( .A1(n7610), .A2(n7698), .ZN(n7835) );
  XOR2_X1 U8517 ( .A(n8657), .B(n8658), .Z(n7832) );
  XOR2_X1 U8518 ( .A(n8659), .B(n8660), .Z(n8658) );
  OR2_X1 U8519 ( .A1(n7608), .A2(n7698), .ZN(n7839) );
  XOR2_X1 U8520 ( .A(n8661), .B(n8662), .Z(n7836) );
  XOR2_X1 U8521 ( .A(n8663), .B(n8664), .Z(n8662) );
  OR2_X1 U8522 ( .A1(n7960), .A2(n7698), .ZN(n7843) );
  INV_X1 U8523 ( .A(n7690), .ZN(n7698) );
  AND2_X1 U8524 ( .A1(n8665), .A2(n8666), .ZN(n7690) );
  INV_X1 U8525 ( .A(n8667), .ZN(n8666) );
  OR2_X1 U8526 ( .A1(c_31_), .A2(d_31_), .ZN(n8665) );
  XOR2_X1 U8527 ( .A(n8668), .B(n8669), .Z(n7840) );
  XOR2_X1 U8528 ( .A(n8670), .B(n8671), .Z(n8669) );
  XOR2_X1 U8529 ( .A(n8404), .B(n8405), .Z(n7849) );
  OR2_X1 U8530 ( .A1(n8672), .A2(n8673), .ZN(n8405) );
  AND2_X1 U8531 ( .A1(n8674), .A2(n8675), .ZN(n8673) );
  AND2_X1 U8532 ( .A1(n8676), .A2(n8677), .ZN(n8672) );
  OR2_X1 U8533 ( .A1(n8674), .A2(n8675), .ZN(n8677) );
  XOR2_X1 U8534 ( .A(n8414), .B(n8678), .Z(n8404) );
  XOR2_X1 U8535 ( .A(n8413), .B(n8412), .Z(n8678) );
  OR2_X1 U8536 ( .A1(n7960), .A2(n7667), .ZN(n8412) );
  OR2_X1 U8537 ( .A1(n8679), .A2(n8680), .ZN(n8413) );
  AND2_X1 U8538 ( .A1(n8681), .A2(n8682), .ZN(n8680) );
  AND2_X1 U8539 ( .A1(n8683), .A2(n8684), .ZN(n8679) );
  OR2_X1 U8540 ( .A1(n8681), .A2(n8682), .ZN(n8684) );
  XOR2_X1 U8541 ( .A(n8422), .B(n8685), .Z(n8414) );
  XOR2_X1 U8542 ( .A(n8421), .B(n8420), .Z(n8685) );
  OR2_X1 U8543 ( .A1(n8023), .A2(n8417), .ZN(n8420) );
  OR2_X1 U8544 ( .A1(n8686), .A2(n8687), .ZN(n8421) );
  AND2_X1 U8545 ( .A1(n8688), .A2(n8689), .ZN(n8687) );
  AND2_X1 U8546 ( .A1(n8690), .A2(n8691), .ZN(n8686) );
  OR2_X1 U8547 ( .A1(n8688), .A2(n8689), .ZN(n8691) );
  XOR2_X1 U8548 ( .A(n8692), .B(n8693), .Z(n8422) );
  XOR2_X1 U8549 ( .A(n8694), .B(n8695), .Z(n8693) );
  XNOR2_X1 U8550 ( .A(n8676), .B(n8696), .ZN(n7845) );
  XOR2_X1 U8551 ( .A(n8675), .B(n8674), .Z(n8696) );
  OR2_X1 U8552 ( .A1(n7702), .A2(n7664), .ZN(n8674) );
  OR2_X1 U8553 ( .A1(n8697), .A2(n8698), .ZN(n8675) );
  AND2_X1 U8554 ( .A1(n8668), .A2(n8671), .ZN(n8698) );
  AND2_X1 U8555 ( .A1(n8699), .A2(n8670), .ZN(n8697) );
  OR2_X1 U8556 ( .A1(n8700), .A2(n8701), .ZN(n8670) );
  AND2_X1 U8557 ( .A1(n8661), .A2(n8664), .ZN(n8701) );
  AND2_X1 U8558 ( .A1(n8702), .A2(n8663), .ZN(n8700) );
  OR2_X1 U8559 ( .A1(n8703), .A2(n8704), .ZN(n8663) );
  AND2_X1 U8560 ( .A1(n8657), .A2(n8660), .ZN(n8704) );
  AND2_X1 U8561 ( .A1(n8705), .A2(n8659), .ZN(n8703) );
  OR2_X1 U8562 ( .A1(n8706), .A2(n8707), .ZN(n8659) );
  AND2_X1 U8563 ( .A1(n8653), .A2(n8656), .ZN(n8707) );
  AND2_X1 U8564 ( .A1(n8708), .A2(n8655), .ZN(n8706) );
  OR2_X1 U8565 ( .A1(n8709), .A2(n8710), .ZN(n8655) );
  AND2_X1 U8566 ( .A1(n8649), .A2(n8652), .ZN(n8710) );
  AND2_X1 U8567 ( .A1(n8711), .A2(n8651), .ZN(n8709) );
  OR2_X1 U8568 ( .A1(n8712), .A2(n8713), .ZN(n8651) );
  AND2_X1 U8569 ( .A1(n8645), .A2(n8648), .ZN(n8713) );
  AND2_X1 U8570 ( .A1(n8714), .A2(n8647), .ZN(n8712) );
  OR2_X1 U8571 ( .A1(n8715), .A2(n8716), .ZN(n8647) );
  AND2_X1 U8572 ( .A1(n8640), .A2(n8643), .ZN(n8716) );
  AND2_X1 U8573 ( .A1(n8717), .A2(n8642), .ZN(n8715) );
  OR2_X1 U8574 ( .A1(n8718), .A2(n8719), .ZN(n8642) );
  AND2_X1 U8575 ( .A1(n8635), .A2(n8638), .ZN(n8719) );
  AND2_X1 U8576 ( .A1(n8720), .A2(n8637), .ZN(n8718) );
  OR2_X1 U8577 ( .A1(n8721), .A2(n8722), .ZN(n8637) );
  AND2_X1 U8578 ( .A1(n8630), .A2(n8633), .ZN(n8722) );
  AND2_X1 U8579 ( .A1(n8723), .A2(n8632), .ZN(n8721) );
  OR2_X1 U8580 ( .A1(n8724), .A2(n8725), .ZN(n8632) );
  AND2_X1 U8581 ( .A1(n8625), .A2(n8628), .ZN(n8725) );
  AND2_X1 U8582 ( .A1(n8726), .A2(n8627), .ZN(n8724) );
  OR2_X1 U8583 ( .A1(n8727), .A2(n8728), .ZN(n8627) );
  AND2_X1 U8584 ( .A1(n8620), .A2(n8623), .ZN(n8728) );
  AND2_X1 U8585 ( .A1(n8729), .A2(n8622), .ZN(n8727) );
  OR2_X1 U8586 ( .A1(n8730), .A2(n8731), .ZN(n8622) );
  AND2_X1 U8587 ( .A1(n8615), .A2(n8618), .ZN(n8731) );
  AND2_X1 U8588 ( .A1(n8732), .A2(n8617), .ZN(n8730) );
  OR2_X1 U8589 ( .A1(n8733), .A2(n8734), .ZN(n8617) );
  AND2_X1 U8590 ( .A1(n8610), .A2(n8613), .ZN(n8734) );
  AND2_X1 U8591 ( .A1(n8735), .A2(n8612), .ZN(n8733) );
  OR2_X1 U8592 ( .A1(n8736), .A2(n8737), .ZN(n8612) );
  AND2_X1 U8593 ( .A1(n8605), .A2(n8608), .ZN(n8737) );
  AND2_X1 U8594 ( .A1(n8738), .A2(n8607), .ZN(n8736) );
  OR2_X1 U8595 ( .A1(n8739), .A2(n8740), .ZN(n8607) );
  AND2_X1 U8596 ( .A1(n8600), .A2(n8603), .ZN(n8740) );
  AND2_X1 U8597 ( .A1(n8741), .A2(n8602), .ZN(n8739) );
  OR2_X1 U8598 ( .A1(n8742), .A2(n8743), .ZN(n8602) );
  AND2_X1 U8599 ( .A1(n8595), .A2(n8598), .ZN(n8743) );
  AND2_X1 U8600 ( .A1(n8744), .A2(n8597), .ZN(n8742) );
  OR2_X1 U8601 ( .A1(n8745), .A2(n8746), .ZN(n8597) );
  AND2_X1 U8602 ( .A1(n8590), .A2(n8593), .ZN(n8746) );
  AND2_X1 U8603 ( .A1(n8747), .A2(n8592), .ZN(n8745) );
  OR2_X1 U8604 ( .A1(n8748), .A2(n8749), .ZN(n8592) );
  AND2_X1 U8605 ( .A1(n8585), .A2(n8588), .ZN(n8749) );
  AND2_X1 U8606 ( .A1(n8750), .A2(n8587), .ZN(n8748) );
  OR2_X1 U8607 ( .A1(n8751), .A2(n8752), .ZN(n8587) );
  AND2_X1 U8608 ( .A1(n8580), .A2(n8583), .ZN(n8752) );
  AND2_X1 U8609 ( .A1(n8753), .A2(n8582), .ZN(n8751) );
  OR2_X1 U8610 ( .A1(n8754), .A2(n8755), .ZN(n8582) );
  AND2_X1 U8611 ( .A1(n8575), .A2(n8578), .ZN(n8755) );
  AND2_X1 U8612 ( .A1(n8756), .A2(n8577), .ZN(n8754) );
  OR2_X1 U8613 ( .A1(n8757), .A2(n8758), .ZN(n8577) );
  AND2_X1 U8614 ( .A1(n8570), .A2(n8573), .ZN(n8758) );
  AND2_X1 U8615 ( .A1(n8759), .A2(n8572), .ZN(n8757) );
  OR2_X1 U8616 ( .A1(n8760), .A2(n8761), .ZN(n8572) );
  AND2_X1 U8617 ( .A1(n8565), .A2(n8568), .ZN(n8761) );
  AND2_X1 U8618 ( .A1(n8762), .A2(n8567), .ZN(n8760) );
  OR2_X1 U8619 ( .A1(n8763), .A2(n8764), .ZN(n8567) );
  AND2_X1 U8620 ( .A1(n8560), .A2(n8563), .ZN(n8764) );
  AND2_X1 U8621 ( .A1(n8765), .A2(n8562), .ZN(n8763) );
  OR2_X1 U8622 ( .A1(n8766), .A2(n8767), .ZN(n8562) );
  AND2_X1 U8623 ( .A1(n8555), .A2(n8558), .ZN(n8767) );
  AND2_X1 U8624 ( .A1(n8768), .A2(n8557), .ZN(n8766) );
  OR2_X1 U8625 ( .A1(n8769), .A2(n8770), .ZN(n8557) );
  AND2_X1 U8626 ( .A1(n8550), .A2(n8553), .ZN(n8770) );
  AND2_X1 U8627 ( .A1(n8771), .A2(n8552), .ZN(n8769) );
  OR2_X1 U8628 ( .A1(n8772), .A2(n8773), .ZN(n8552) );
  AND2_X1 U8629 ( .A1(n8545), .A2(n8548), .ZN(n8773) );
  AND2_X1 U8630 ( .A1(n8774), .A2(n8547), .ZN(n8772) );
  OR2_X1 U8631 ( .A1(n8775), .A2(n8776), .ZN(n8547) );
  AND2_X1 U8632 ( .A1(n8540), .A2(n8543), .ZN(n8776) );
  AND2_X1 U8633 ( .A1(n8777), .A2(n8542), .ZN(n8775) );
  OR2_X1 U8634 ( .A1(n8778), .A2(n8779), .ZN(n8542) );
  AND2_X1 U8635 ( .A1(n8535), .A2(n8538), .ZN(n8779) );
  AND2_X1 U8636 ( .A1(n8780), .A2(n8537), .ZN(n8778) );
  OR2_X1 U8637 ( .A1(n8781), .A2(n8782), .ZN(n8537) );
  AND2_X1 U8638 ( .A1(n8530), .A2(n8533), .ZN(n8782) );
  AND2_X1 U8639 ( .A1(n8532), .A2(n8783), .ZN(n8781) );
  OR2_X1 U8640 ( .A1(n8533), .A2(n8530), .ZN(n8783) );
  OR2_X1 U8641 ( .A1(n7702), .A2(n7606), .ZN(n8530) );
  OR3_X1 U8642 ( .A1(n7702), .A2(n8519), .A3(n7667), .ZN(n8533) );
  INV_X1 U8643 ( .A(n8784), .ZN(n8532) );
  OR2_X1 U8644 ( .A1(n8785), .A2(n8786), .ZN(n8784) );
  AND2_X1 U8645 ( .A1(n8787), .A2(n8788), .ZN(n8786) );
  OR2_X1 U8646 ( .A1(n8789), .A2(n7697), .ZN(n8788) );
  AND2_X1 U8647 ( .A1(n7691), .A2(n8528), .ZN(n8789) );
  AND2_X1 U8648 ( .A1(n8523), .A2(n8790), .ZN(n8785) );
  OR2_X1 U8649 ( .A1(n8791), .A2(n7701), .ZN(n8790) );
  AND2_X1 U8650 ( .A1(n8417), .A2(n7703), .ZN(n8791) );
  INV_X1 U8651 ( .A(n8528), .ZN(n8523) );
  OR2_X1 U8652 ( .A1(n8538), .A2(n8535), .ZN(n8780) );
  XNOR2_X1 U8653 ( .A(n8792), .B(n8793), .ZN(n8535) );
  XNOR2_X1 U8654 ( .A(n8794), .B(n8795), .ZN(n8793) );
  OR2_X1 U8655 ( .A1(n7662), .A2(n7665), .ZN(n8538) );
  OR2_X1 U8656 ( .A1(n8543), .A2(n8540), .ZN(n8777) );
  XOR2_X1 U8657 ( .A(n8796), .B(n8797), .Z(n8540) );
  XOR2_X1 U8658 ( .A(n8798), .B(n8799), .Z(n8797) );
  OR2_X1 U8659 ( .A1(n7660), .A2(n7665), .ZN(n8543) );
  OR2_X1 U8660 ( .A1(n8548), .A2(n8545), .ZN(n8774) );
  XOR2_X1 U8661 ( .A(n8800), .B(n8801), .Z(n8545) );
  XOR2_X1 U8662 ( .A(n8802), .B(n8803), .Z(n8801) );
  OR2_X1 U8663 ( .A1(n7658), .A2(n7665), .ZN(n8548) );
  OR2_X1 U8664 ( .A1(n8553), .A2(n8550), .ZN(n8771) );
  XOR2_X1 U8665 ( .A(n8804), .B(n8805), .Z(n8550) );
  XOR2_X1 U8666 ( .A(n8806), .B(n8807), .Z(n8805) );
  OR2_X1 U8667 ( .A1(n7656), .A2(n7665), .ZN(n8553) );
  OR2_X1 U8668 ( .A1(n8558), .A2(n8555), .ZN(n8768) );
  XOR2_X1 U8669 ( .A(n8808), .B(n8809), .Z(n8555) );
  XOR2_X1 U8670 ( .A(n8810), .B(n8811), .Z(n8809) );
  OR2_X1 U8671 ( .A1(n7654), .A2(n7665), .ZN(n8558) );
  OR2_X1 U8672 ( .A1(n8563), .A2(n8560), .ZN(n8765) );
  XOR2_X1 U8673 ( .A(n8812), .B(n8813), .Z(n8560) );
  XOR2_X1 U8674 ( .A(n8814), .B(n8815), .Z(n8813) );
  OR2_X1 U8675 ( .A1(n7652), .A2(n7665), .ZN(n8563) );
  OR2_X1 U8676 ( .A1(n8568), .A2(n8565), .ZN(n8762) );
  XOR2_X1 U8677 ( .A(n8816), .B(n8817), .Z(n8565) );
  XOR2_X1 U8678 ( .A(n8818), .B(n8819), .Z(n8817) );
  OR2_X1 U8679 ( .A1(n7650), .A2(n7665), .ZN(n8568) );
  OR2_X1 U8680 ( .A1(n8573), .A2(n8570), .ZN(n8759) );
  XOR2_X1 U8681 ( .A(n8820), .B(n8821), .Z(n8570) );
  XOR2_X1 U8682 ( .A(n8822), .B(n8823), .Z(n8821) );
  OR2_X1 U8683 ( .A1(n7648), .A2(n7665), .ZN(n8573) );
  OR2_X1 U8684 ( .A1(n8578), .A2(n8575), .ZN(n8756) );
  XOR2_X1 U8685 ( .A(n8824), .B(n8825), .Z(n8575) );
  XOR2_X1 U8686 ( .A(n8826), .B(n8827), .Z(n8825) );
  OR2_X1 U8687 ( .A1(n7646), .A2(n7665), .ZN(n8578) );
  OR2_X1 U8688 ( .A1(n8583), .A2(n8580), .ZN(n8753) );
  XOR2_X1 U8689 ( .A(n8828), .B(n8829), .Z(n8580) );
  XOR2_X1 U8690 ( .A(n8830), .B(n8831), .Z(n8829) );
  OR2_X1 U8691 ( .A1(n7644), .A2(n7665), .ZN(n8583) );
  OR2_X1 U8692 ( .A1(n8588), .A2(n8585), .ZN(n8750) );
  XOR2_X1 U8693 ( .A(n8832), .B(n8833), .Z(n8585) );
  XOR2_X1 U8694 ( .A(n8834), .B(n8835), .Z(n8833) );
  OR2_X1 U8695 ( .A1(n7642), .A2(n7665), .ZN(n8588) );
  OR2_X1 U8696 ( .A1(n8593), .A2(n8590), .ZN(n8747) );
  XOR2_X1 U8697 ( .A(n8836), .B(n8837), .Z(n8590) );
  XOR2_X1 U8698 ( .A(n8838), .B(n8839), .Z(n8837) );
  OR2_X1 U8699 ( .A1(n7640), .A2(n7665), .ZN(n8593) );
  OR2_X1 U8700 ( .A1(n8598), .A2(n8595), .ZN(n8744) );
  XOR2_X1 U8701 ( .A(n8840), .B(n8841), .Z(n8595) );
  XOR2_X1 U8702 ( .A(n8842), .B(n8843), .Z(n8841) );
  OR2_X1 U8703 ( .A1(n7638), .A2(n7665), .ZN(n8598) );
  OR2_X1 U8704 ( .A1(n8603), .A2(n8600), .ZN(n8741) );
  XOR2_X1 U8705 ( .A(n8844), .B(n8845), .Z(n8600) );
  XOR2_X1 U8706 ( .A(n8846), .B(n8847), .Z(n8845) );
  OR2_X1 U8707 ( .A1(n7636), .A2(n7665), .ZN(n8603) );
  OR2_X1 U8708 ( .A1(n8608), .A2(n8605), .ZN(n8738) );
  XOR2_X1 U8709 ( .A(n8848), .B(n8849), .Z(n8605) );
  XOR2_X1 U8710 ( .A(n8850), .B(n8851), .Z(n8849) );
  OR2_X1 U8711 ( .A1(n7634), .A2(n7665), .ZN(n8608) );
  OR2_X1 U8712 ( .A1(n8613), .A2(n8610), .ZN(n8735) );
  XOR2_X1 U8713 ( .A(n8852), .B(n8853), .Z(n8610) );
  XOR2_X1 U8714 ( .A(n8854), .B(n8855), .Z(n8853) );
  OR2_X1 U8715 ( .A1(n7632), .A2(n7665), .ZN(n8613) );
  OR2_X1 U8716 ( .A1(n8618), .A2(n8615), .ZN(n8732) );
  XOR2_X1 U8717 ( .A(n8856), .B(n8857), .Z(n8615) );
  XOR2_X1 U8718 ( .A(n8858), .B(n8859), .Z(n8857) );
  OR2_X1 U8719 ( .A1(n7630), .A2(n7665), .ZN(n8618) );
  OR2_X1 U8720 ( .A1(n8623), .A2(n8620), .ZN(n8729) );
  XOR2_X1 U8721 ( .A(n8860), .B(n8861), .Z(n8620) );
  XOR2_X1 U8722 ( .A(n8862), .B(n8863), .Z(n8861) );
  OR2_X1 U8723 ( .A1(n7628), .A2(n7665), .ZN(n8623) );
  OR2_X1 U8724 ( .A1(n8628), .A2(n8625), .ZN(n8726) );
  XOR2_X1 U8725 ( .A(n8864), .B(n8865), .Z(n8625) );
  XOR2_X1 U8726 ( .A(n8866), .B(n8867), .Z(n8865) );
  OR2_X1 U8727 ( .A1(n7626), .A2(n7665), .ZN(n8628) );
  OR2_X1 U8728 ( .A1(n8633), .A2(n8630), .ZN(n8723) );
  XOR2_X1 U8729 ( .A(n8868), .B(n8869), .Z(n8630) );
  XOR2_X1 U8730 ( .A(n8870), .B(n8871), .Z(n8869) );
  OR2_X1 U8731 ( .A1(n7624), .A2(n7702), .ZN(n8633) );
  OR2_X1 U8732 ( .A1(n8638), .A2(n8635), .ZN(n8720) );
  XOR2_X1 U8733 ( .A(n8872), .B(n8873), .Z(n8635) );
  XOR2_X1 U8734 ( .A(n8874), .B(n8875), .Z(n8873) );
  OR2_X1 U8735 ( .A1(n7622), .A2(n7702), .ZN(n8638) );
  OR2_X1 U8736 ( .A1(n8643), .A2(n8640), .ZN(n8717) );
  XOR2_X1 U8737 ( .A(n8876), .B(n8877), .Z(n8640) );
  XOR2_X1 U8738 ( .A(n8878), .B(n8879), .Z(n8877) );
  OR2_X1 U8739 ( .A1(n7620), .A2(n7702), .ZN(n8643) );
  OR2_X1 U8740 ( .A1(n8648), .A2(n8645), .ZN(n8714) );
  XOR2_X1 U8741 ( .A(n8880), .B(n8881), .Z(n8645) );
  XOR2_X1 U8742 ( .A(n8882), .B(n8883), .Z(n8881) );
  OR2_X1 U8743 ( .A1(n7618), .A2(n7702), .ZN(n8648) );
  OR2_X1 U8744 ( .A1(n8652), .A2(n8649), .ZN(n8711) );
  XOR2_X1 U8745 ( .A(n8884), .B(n8885), .Z(n8649) );
  XOR2_X1 U8746 ( .A(n8886), .B(n8887), .Z(n8885) );
  OR2_X1 U8747 ( .A1(n7616), .A2(n7702), .ZN(n8652) );
  OR2_X1 U8748 ( .A1(n8656), .A2(n8653), .ZN(n8708) );
  XOR2_X1 U8749 ( .A(n8888), .B(n8889), .Z(n8653) );
  XOR2_X1 U8750 ( .A(n8890), .B(n8891), .Z(n8889) );
  OR2_X1 U8751 ( .A1(n7614), .A2(n7702), .ZN(n8656) );
  OR2_X1 U8752 ( .A1(n8660), .A2(n8657), .ZN(n8705) );
  XOR2_X1 U8753 ( .A(n8892), .B(n8893), .Z(n8657) );
  XOR2_X1 U8754 ( .A(n8894), .B(n8895), .Z(n8893) );
  OR2_X1 U8755 ( .A1(n7612), .A2(n7702), .ZN(n8660) );
  OR2_X1 U8756 ( .A1(n8664), .A2(n8661), .ZN(n8702) );
  XOR2_X1 U8757 ( .A(n8896), .B(n8897), .Z(n8661) );
  XOR2_X1 U8758 ( .A(n8898), .B(n8899), .Z(n8897) );
  OR2_X1 U8759 ( .A1(n7610), .A2(n7702), .ZN(n8664) );
  OR2_X1 U8760 ( .A1(n8671), .A2(n8668), .ZN(n8699) );
  XOR2_X1 U8761 ( .A(n8900), .B(n8901), .Z(n8668) );
  XOR2_X1 U8762 ( .A(n8902), .B(n8903), .Z(n8901) );
  OR2_X1 U8763 ( .A1(n8023), .A2(n7702), .ZN(n8671) );
  XNOR2_X1 U8764 ( .A(n8667), .B(n8904), .ZN(n7702) );
  XOR2_X1 U8765 ( .A(d_30_), .B(c_30_), .Z(n8904) );
  XOR2_X1 U8766 ( .A(n8683), .B(n8905), .Z(n8676) );
  XOR2_X1 U8767 ( .A(n8682), .B(n8681), .Z(n8905) );
  OR2_X1 U8768 ( .A1(n8023), .A2(n7667), .ZN(n8681) );
  OR2_X1 U8769 ( .A1(n8906), .A2(n8907), .ZN(n8682) );
  AND2_X1 U8770 ( .A1(n8903), .A2(n8902), .ZN(n8907) );
  AND2_X1 U8771 ( .A1(n8900), .A2(n8908), .ZN(n8906) );
  OR2_X1 U8772 ( .A1(n8903), .A2(n8902), .ZN(n8908) );
  OR2_X1 U8773 ( .A1(n7610), .A2(n7667), .ZN(n8902) );
  OR2_X1 U8774 ( .A1(n8909), .A2(n8910), .ZN(n8903) );
  AND2_X1 U8775 ( .A1(n8899), .A2(n8898), .ZN(n8910) );
  AND2_X1 U8776 ( .A1(n8896), .A2(n8911), .ZN(n8909) );
  OR2_X1 U8777 ( .A1(n8899), .A2(n8898), .ZN(n8911) );
  OR2_X1 U8778 ( .A1(n8912), .A2(n8913), .ZN(n8898) );
  AND2_X1 U8779 ( .A1(n8895), .A2(n8894), .ZN(n8913) );
  AND2_X1 U8780 ( .A1(n8892), .A2(n8914), .ZN(n8912) );
  OR2_X1 U8781 ( .A1(n8895), .A2(n8894), .ZN(n8914) );
  OR2_X1 U8782 ( .A1(n8915), .A2(n8916), .ZN(n8894) );
  AND2_X1 U8783 ( .A1(n8891), .A2(n8890), .ZN(n8916) );
  AND2_X1 U8784 ( .A1(n8888), .A2(n8917), .ZN(n8915) );
  OR2_X1 U8785 ( .A1(n8891), .A2(n8890), .ZN(n8917) );
  OR2_X1 U8786 ( .A1(n8918), .A2(n8919), .ZN(n8890) );
  AND2_X1 U8787 ( .A1(n8887), .A2(n8886), .ZN(n8919) );
  AND2_X1 U8788 ( .A1(n8884), .A2(n8920), .ZN(n8918) );
  OR2_X1 U8789 ( .A1(n8887), .A2(n8886), .ZN(n8920) );
  OR2_X1 U8790 ( .A1(n8921), .A2(n8922), .ZN(n8886) );
  AND2_X1 U8791 ( .A1(n8883), .A2(n8882), .ZN(n8922) );
  AND2_X1 U8792 ( .A1(n8880), .A2(n8923), .ZN(n8921) );
  OR2_X1 U8793 ( .A1(n8883), .A2(n8882), .ZN(n8923) );
  OR2_X1 U8794 ( .A1(n8924), .A2(n8925), .ZN(n8882) );
  AND2_X1 U8795 ( .A1(n8879), .A2(n8878), .ZN(n8925) );
  AND2_X1 U8796 ( .A1(n8876), .A2(n8926), .ZN(n8924) );
  OR2_X1 U8797 ( .A1(n8879), .A2(n8878), .ZN(n8926) );
  OR2_X1 U8798 ( .A1(n8927), .A2(n8928), .ZN(n8878) );
  AND2_X1 U8799 ( .A1(n8875), .A2(n8874), .ZN(n8928) );
  AND2_X1 U8800 ( .A1(n8872), .A2(n8929), .ZN(n8927) );
  OR2_X1 U8801 ( .A1(n8875), .A2(n8874), .ZN(n8929) );
  OR2_X1 U8802 ( .A1(n8930), .A2(n8931), .ZN(n8874) );
  AND2_X1 U8803 ( .A1(n8871), .A2(n8870), .ZN(n8931) );
  AND2_X1 U8804 ( .A1(n8868), .A2(n8932), .ZN(n8930) );
  OR2_X1 U8805 ( .A1(n8871), .A2(n8870), .ZN(n8932) );
  OR2_X1 U8806 ( .A1(n8933), .A2(n8934), .ZN(n8870) );
  AND2_X1 U8807 ( .A1(n8867), .A2(n8866), .ZN(n8934) );
  AND2_X1 U8808 ( .A1(n8864), .A2(n8935), .ZN(n8933) );
  OR2_X1 U8809 ( .A1(n8867), .A2(n8866), .ZN(n8935) );
  OR2_X1 U8810 ( .A1(n8936), .A2(n8937), .ZN(n8866) );
  AND2_X1 U8811 ( .A1(n8863), .A2(n8862), .ZN(n8937) );
  AND2_X1 U8812 ( .A1(n8860), .A2(n8938), .ZN(n8936) );
  OR2_X1 U8813 ( .A1(n8863), .A2(n8862), .ZN(n8938) );
  OR2_X1 U8814 ( .A1(n8939), .A2(n8940), .ZN(n8862) );
  AND2_X1 U8815 ( .A1(n8859), .A2(n8858), .ZN(n8940) );
  AND2_X1 U8816 ( .A1(n8856), .A2(n8941), .ZN(n8939) );
  OR2_X1 U8817 ( .A1(n8859), .A2(n8858), .ZN(n8941) );
  OR2_X1 U8818 ( .A1(n8942), .A2(n8943), .ZN(n8858) );
  AND2_X1 U8819 ( .A1(n8855), .A2(n8854), .ZN(n8943) );
  AND2_X1 U8820 ( .A1(n8852), .A2(n8944), .ZN(n8942) );
  OR2_X1 U8821 ( .A1(n8855), .A2(n8854), .ZN(n8944) );
  OR2_X1 U8822 ( .A1(n8945), .A2(n8946), .ZN(n8854) );
  AND2_X1 U8823 ( .A1(n8851), .A2(n8850), .ZN(n8946) );
  AND2_X1 U8824 ( .A1(n8848), .A2(n8947), .ZN(n8945) );
  OR2_X1 U8825 ( .A1(n8851), .A2(n8850), .ZN(n8947) );
  OR2_X1 U8826 ( .A1(n8948), .A2(n8949), .ZN(n8850) );
  AND2_X1 U8827 ( .A1(n8847), .A2(n8846), .ZN(n8949) );
  AND2_X1 U8828 ( .A1(n8844), .A2(n8950), .ZN(n8948) );
  OR2_X1 U8829 ( .A1(n8847), .A2(n8846), .ZN(n8950) );
  OR2_X1 U8830 ( .A1(n8951), .A2(n8952), .ZN(n8846) );
  AND2_X1 U8831 ( .A1(n8843), .A2(n8842), .ZN(n8952) );
  AND2_X1 U8832 ( .A1(n8840), .A2(n8953), .ZN(n8951) );
  OR2_X1 U8833 ( .A1(n8843), .A2(n8842), .ZN(n8953) );
  OR2_X1 U8834 ( .A1(n8954), .A2(n8955), .ZN(n8842) );
  AND2_X1 U8835 ( .A1(n8839), .A2(n8838), .ZN(n8955) );
  AND2_X1 U8836 ( .A1(n8836), .A2(n8956), .ZN(n8954) );
  OR2_X1 U8837 ( .A1(n8839), .A2(n8838), .ZN(n8956) );
  OR2_X1 U8838 ( .A1(n8957), .A2(n8958), .ZN(n8838) );
  AND2_X1 U8839 ( .A1(n8835), .A2(n8834), .ZN(n8958) );
  AND2_X1 U8840 ( .A1(n8832), .A2(n8959), .ZN(n8957) );
  OR2_X1 U8841 ( .A1(n8835), .A2(n8834), .ZN(n8959) );
  OR2_X1 U8842 ( .A1(n8960), .A2(n8961), .ZN(n8834) );
  AND2_X1 U8843 ( .A1(n8831), .A2(n8830), .ZN(n8961) );
  AND2_X1 U8844 ( .A1(n8828), .A2(n8962), .ZN(n8960) );
  OR2_X1 U8845 ( .A1(n8831), .A2(n8830), .ZN(n8962) );
  OR2_X1 U8846 ( .A1(n8963), .A2(n8964), .ZN(n8830) );
  AND2_X1 U8847 ( .A1(n8827), .A2(n8826), .ZN(n8964) );
  AND2_X1 U8848 ( .A1(n8824), .A2(n8965), .ZN(n8963) );
  OR2_X1 U8849 ( .A1(n8827), .A2(n8826), .ZN(n8965) );
  OR2_X1 U8850 ( .A1(n8966), .A2(n8967), .ZN(n8826) );
  AND2_X1 U8851 ( .A1(n8823), .A2(n8822), .ZN(n8967) );
  AND2_X1 U8852 ( .A1(n8820), .A2(n8968), .ZN(n8966) );
  OR2_X1 U8853 ( .A1(n8823), .A2(n8822), .ZN(n8968) );
  OR2_X1 U8854 ( .A1(n8969), .A2(n8970), .ZN(n8822) );
  AND2_X1 U8855 ( .A1(n8819), .A2(n8818), .ZN(n8970) );
  AND2_X1 U8856 ( .A1(n8816), .A2(n8971), .ZN(n8969) );
  OR2_X1 U8857 ( .A1(n8819), .A2(n8818), .ZN(n8971) );
  OR2_X1 U8858 ( .A1(n8972), .A2(n8973), .ZN(n8818) );
  AND2_X1 U8859 ( .A1(n8815), .A2(n8814), .ZN(n8973) );
  AND2_X1 U8860 ( .A1(n8812), .A2(n8974), .ZN(n8972) );
  OR2_X1 U8861 ( .A1(n8815), .A2(n8814), .ZN(n8974) );
  OR2_X1 U8862 ( .A1(n8975), .A2(n8976), .ZN(n8814) );
  AND2_X1 U8863 ( .A1(n8811), .A2(n8810), .ZN(n8976) );
  AND2_X1 U8864 ( .A1(n8808), .A2(n8977), .ZN(n8975) );
  OR2_X1 U8865 ( .A1(n8811), .A2(n8810), .ZN(n8977) );
  OR2_X1 U8866 ( .A1(n8978), .A2(n8979), .ZN(n8810) );
  AND2_X1 U8867 ( .A1(n8807), .A2(n8806), .ZN(n8979) );
  AND2_X1 U8868 ( .A1(n8804), .A2(n8980), .ZN(n8978) );
  OR2_X1 U8869 ( .A1(n8807), .A2(n8806), .ZN(n8980) );
  OR2_X1 U8870 ( .A1(n8981), .A2(n8982), .ZN(n8806) );
  AND2_X1 U8871 ( .A1(n8803), .A2(n8802), .ZN(n8982) );
  AND2_X1 U8872 ( .A1(n8800), .A2(n8983), .ZN(n8981) );
  OR2_X1 U8873 ( .A1(n8803), .A2(n8802), .ZN(n8983) );
  OR2_X1 U8874 ( .A1(n8984), .A2(n8985), .ZN(n8802) );
  AND2_X1 U8875 ( .A1(n8799), .A2(n8798), .ZN(n8985) );
  AND2_X1 U8876 ( .A1(n8796), .A2(n8986), .ZN(n8984) );
  OR2_X1 U8877 ( .A1(n8799), .A2(n8798), .ZN(n8986) );
  OR2_X1 U8878 ( .A1(n8987), .A2(n8988), .ZN(n8798) );
  AND2_X1 U8879 ( .A1(n8792), .A2(n8795), .ZN(n8988) );
  AND2_X1 U8880 ( .A1(n8794), .A2(n8989), .ZN(n8987) );
  OR2_X1 U8881 ( .A1(n8792), .A2(n8795), .ZN(n8989) );
  OR3_X1 U8882 ( .A1(n8417), .A2(n8519), .A3(n7667), .ZN(n8795) );
  OR2_X1 U8883 ( .A1(n8518), .A2(n7667), .ZN(n8792) );
  INV_X1 U8884 ( .A(n8990), .ZN(n8794) );
  OR2_X1 U8885 ( .A1(n8991), .A2(n8992), .ZN(n8990) );
  AND2_X1 U8886 ( .A1(n8993), .A2(n8994), .ZN(n8992) );
  OR2_X1 U8887 ( .A1(n8995), .A2(n7697), .ZN(n8994) );
  AND2_X1 U8888 ( .A1(n8417), .A2(n7691), .ZN(n8995) );
  AND2_X1 U8889 ( .A1(n8787), .A2(n8996), .ZN(n8991) );
  OR2_X1 U8890 ( .A1(n8997), .A2(n7701), .ZN(n8996) );
  AND2_X1 U8891 ( .A1(n8998), .A2(n7703), .ZN(n8997) );
  OR2_X1 U8892 ( .A1(n7662), .A2(n7667), .ZN(n8799) );
  XNOR2_X1 U8893 ( .A(n8999), .B(n9000), .ZN(n8796) );
  XNOR2_X1 U8894 ( .A(n9001), .B(n9002), .ZN(n9000) );
  OR2_X1 U8895 ( .A1(n7660), .A2(n7667), .ZN(n8803) );
  XOR2_X1 U8896 ( .A(n9003), .B(n9004), .Z(n8800) );
  XOR2_X1 U8897 ( .A(n9005), .B(n9006), .Z(n9004) );
  OR2_X1 U8898 ( .A1(n7658), .A2(n7667), .ZN(n8807) );
  XOR2_X1 U8899 ( .A(n9007), .B(n9008), .Z(n8804) );
  XOR2_X1 U8900 ( .A(n9009), .B(n9010), .Z(n9008) );
  OR2_X1 U8901 ( .A1(n7656), .A2(n7667), .ZN(n8811) );
  XOR2_X1 U8902 ( .A(n9011), .B(n9012), .Z(n8808) );
  XOR2_X1 U8903 ( .A(n9013), .B(n9014), .Z(n9012) );
  OR2_X1 U8904 ( .A1(n7654), .A2(n7667), .ZN(n8815) );
  XOR2_X1 U8905 ( .A(n9015), .B(n9016), .Z(n8812) );
  XOR2_X1 U8906 ( .A(n9017), .B(n9018), .Z(n9016) );
  OR2_X1 U8907 ( .A1(n7652), .A2(n7667), .ZN(n8819) );
  XOR2_X1 U8908 ( .A(n9019), .B(n9020), .Z(n8816) );
  XOR2_X1 U8909 ( .A(n9021), .B(n9022), .Z(n9020) );
  OR2_X1 U8910 ( .A1(n7650), .A2(n7667), .ZN(n8823) );
  XOR2_X1 U8911 ( .A(n9023), .B(n9024), .Z(n8820) );
  XOR2_X1 U8912 ( .A(n9025), .B(n9026), .Z(n9024) );
  OR2_X1 U8913 ( .A1(n7648), .A2(n7667), .ZN(n8827) );
  XOR2_X1 U8914 ( .A(n9027), .B(n9028), .Z(n8824) );
  XOR2_X1 U8915 ( .A(n9029), .B(n9030), .Z(n9028) );
  OR2_X1 U8916 ( .A1(n7646), .A2(n7667), .ZN(n8831) );
  XOR2_X1 U8917 ( .A(n9031), .B(n9032), .Z(n8828) );
  XOR2_X1 U8918 ( .A(n9033), .B(n9034), .Z(n9032) );
  OR2_X1 U8919 ( .A1(n7644), .A2(n7667), .ZN(n8835) );
  XOR2_X1 U8920 ( .A(n9035), .B(n9036), .Z(n8832) );
  XOR2_X1 U8921 ( .A(n9037), .B(n9038), .Z(n9036) );
  OR2_X1 U8922 ( .A1(n7642), .A2(n7667), .ZN(n8839) );
  XOR2_X1 U8923 ( .A(n9039), .B(n9040), .Z(n8836) );
  XOR2_X1 U8924 ( .A(n9041), .B(n9042), .Z(n9040) );
  OR2_X1 U8925 ( .A1(n7640), .A2(n7667), .ZN(n8843) );
  XOR2_X1 U8926 ( .A(n9043), .B(n9044), .Z(n8840) );
  XOR2_X1 U8927 ( .A(n9045), .B(n9046), .Z(n9044) );
  OR2_X1 U8928 ( .A1(n7638), .A2(n7667), .ZN(n8847) );
  XOR2_X1 U8929 ( .A(n9047), .B(n9048), .Z(n8844) );
  XOR2_X1 U8930 ( .A(n9049), .B(n9050), .Z(n9048) );
  OR2_X1 U8931 ( .A1(n7636), .A2(n7667), .ZN(n8851) );
  XOR2_X1 U8932 ( .A(n9051), .B(n9052), .Z(n8848) );
  XOR2_X1 U8933 ( .A(n9053), .B(n9054), .Z(n9052) );
  OR2_X1 U8934 ( .A1(n7634), .A2(n8528), .ZN(n8855) );
  XOR2_X1 U8935 ( .A(n9055), .B(n9056), .Z(n8852) );
  XOR2_X1 U8936 ( .A(n9057), .B(n9058), .Z(n9056) );
  OR2_X1 U8937 ( .A1(n7632), .A2(n8528), .ZN(n8859) );
  XOR2_X1 U8938 ( .A(n9059), .B(n9060), .Z(n8856) );
  XOR2_X1 U8939 ( .A(n9061), .B(n9062), .Z(n9060) );
  OR2_X1 U8940 ( .A1(n7630), .A2(n8528), .ZN(n8863) );
  XOR2_X1 U8941 ( .A(n9063), .B(n9064), .Z(n8860) );
  XOR2_X1 U8942 ( .A(n9065), .B(n9066), .Z(n9064) );
  OR2_X1 U8943 ( .A1(n7628), .A2(n8528), .ZN(n8867) );
  XOR2_X1 U8944 ( .A(n9067), .B(n9068), .Z(n8864) );
  XOR2_X1 U8945 ( .A(n9069), .B(n9070), .Z(n9068) );
  OR2_X1 U8946 ( .A1(n7626), .A2(n8528), .ZN(n8871) );
  XOR2_X1 U8947 ( .A(n9071), .B(n9072), .Z(n8868) );
  XOR2_X1 U8948 ( .A(n9073), .B(n9074), .Z(n9072) );
  OR2_X1 U8949 ( .A1(n7624), .A2(n8528), .ZN(n8875) );
  XOR2_X1 U8950 ( .A(n9075), .B(n9076), .Z(n8872) );
  XOR2_X1 U8951 ( .A(n9077), .B(n9078), .Z(n9076) );
  OR2_X1 U8952 ( .A1(n7622), .A2(n8528), .ZN(n8879) );
  XOR2_X1 U8953 ( .A(n9079), .B(n9080), .Z(n8876) );
  XOR2_X1 U8954 ( .A(n9081), .B(n9082), .Z(n9080) );
  OR2_X1 U8955 ( .A1(n7620), .A2(n8528), .ZN(n8883) );
  XOR2_X1 U8956 ( .A(n9083), .B(n9084), .Z(n8880) );
  XOR2_X1 U8957 ( .A(n9085), .B(n9086), .Z(n9084) );
  OR2_X1 U8958 ( .A1(n7618), .A2(n8528), .ZN(n8887) );
  XOR2_X1 U8959 ( .A(n9087), .B(n9088), .Z(n8884) );
  XOR2_X1 U8960 ( .A(n9089), .B(n9090), .Z(n9088) );
  OR2_X1 U8961 ( .A1(n7616), .A2(n8528), .ZN(n8891) );
  XOR2_X1 U8962 ( .A(n9091), .B(n9092), .Z(n8888) );
  XOR2_X1 U8963 ( .A(n9093), .B(n9094), .Z(n9092) );
  OR2_X1 U8964 ( .A1(n7614), .A2(n8528), .ZN(n8895) );
  XOR2_X1 U8965 ( .A(n9095), .B(n9096), .Z(n8892) );
  XOR2_X1 U8966 ( .A(n9097), .B(n9098), .Z(n9096) );
  OR2_X1 U8967 ( .A1(n7612), .A2(n8528), .ZN(n8899) );
  XOR2_X1 U8968 ( .A(n9099), .B(n9100), .Z(n8528) );
  XNOR2_X1 U8969 ( .A(n9101), .B(c_29_), .ZN(n9100) );
  XOR2_X1 U8970 ( .A(n9102), .B(n9103), .Z(n8896) );
  XOR2_X1 U8971 ( .A(n9104), .B(n9105), .Z(n9103) );
  XOR2_X1 U8972 ( .A(n9106), .B(n9107), .Z(n8900) );
  XOR2_X1 U8973 ( .A(n9108), .B(n9109), .Z(n9107) );
  XOR2_X1 U8974 ( .A(n8690), .B(n9110), .Z(n8683) );
  XOR2_X1 U8975 ( .A(n8689), .B(n8688), .Z(n9110) );
  OR2_X1 U8976 ( .A1(n9111), .A2(n9112), .ZN(n8688) );
  AND2_X1 U8977 ( .A1(n9109), .A2(n9108), .ZN(n9112) );
  AND2_X1 U8978 ( .A1(n9106), .A2(n9113), .ZN(n9111) );
  OR2_X1 U8979 ( .A1(n9109), .A2(n9108), .ZN(n9113) );
  OR2_X1 U8980 ( .A1(n9114), .A2(n9115), .ZN(n9108) );
  AND2_X1 U8981 ( .A1(n9105), .A2(n9104), .ZN(n9115) );
  AND2_X1 U8982 ( .A1(n9102), .A2(n9116), .ZN(n9114) );
  OR2_X1 U8983 ( .A1(n9105), .A2(n9104), .ZN(n9116) );
  OR2_X1 U8984 ( .A1(n9117), .A2(n9118), .ZN(n9104) );
  AND2_X1 U8985 ( .A1(n9098), .A2(n9097), .ZN(n9118) );
  AND2_X1 U8986 ( .A1(n9095), .A2(n9119), .ZN(n9117) );
  OR2_X1 U8987 ( .A1(n9098), .A2(n9097), .ZN(n9119) );
  OR2_X1 U8988 ( .A1(n9120), .A2(n9121), .ZN(n9097) );
  AND2_X1 U8989 ( .A1(n9094), .A2(n9093), .ZN(n9121) );
  AND2_X1 U8990 ( .A1(n9091), .A2(n9122), .ZN(n9120) );
  OR2_X1 U8991 ( .A1(n9094), .A2(n9093), .ZN(n9122) );
  OR2_X1 U8992 ( .A1(n9123), .A2(n9124), .ZN(n9093) );
  AND2_X1 U8993 ( .A1(n9090), .A2(n9089), .ZN(n9124) );
  AND2_X1 U8994 ( .A1(n9087), .A2(n9125), .ZN(n9123) );
  OR2_X1 U8995 ( .A1(n9090), .A2(n9089), .ZN(n9125) );
  OR2_X1 U8996 ( .A1(n9126), .A2(n9127), .ZN(n9089) );
  AND2_X1 U8997 ( .A1(n9086), .A2(n9085), .ZN(n9127) );
  AND2_X1 U8998 ( .A1(n9083), .A2(n9128), .ZN(n9126) );
  OR2_X1 U8999 ( .A1(n9086), .A2(n9085), .ZN(n9128) );
  OR2_X1 U9000 ( .A1(n9129), .A2(n9130), .ZN(n9085) );
  AND2_X1 U9001 ( .A1(n9082), .A2(n9081), .ZN(n9130) );
  AND2_X1 U9002 ( .A1(n9079), .A2(n9131), .ZN(n9129) );
  OR2_X1 U9003 ( .A1(n9082), .A2(n9081), .ZN(n9131) );
  OR2_X1 U9004 ( .A1(n9132), .A2(n9133), .ZN(n9081) );
  AND2_X1 U9005 ( .A1(n9078), .A2(n9077), .ZN(n9133) );
  AND2_X1 U9006 ( .A1(n9075), .A2(n9134), .ZN(n9132) );
  OR2_X1 U9007 ( .A1(n9078), .A2(n9077), .ZN(n9134) );
  OR2_X1 U9008 ( .A1(n9135), .A2(n9136), .ZN(n9077) );
  AND2_X1 U9009 ( .A1(n9074), .A2(n9073), .ZN(n9136) );
  AND2_X1 U9010 ( .A1(n9071), .A2(n9137), .ZN(n9135) );
  OR2_X1 U9011 ( .A1(n9074), .A2(n9073), .ZN(n9137) );
  OR2_X1 U9012 ( .A1(n9138), .A2(n9139), .ZN(n9073) );
  AND2_X1 U9013 ( .A1(n9070), .A2(n9069), .ZN(n9139) );
  AND2_X1 U9014 ( .A1(n9067), .A2(n9140), .ZN(n9138) );
  OR2_X1 U9015 ( .A1(n9070), .A2(n9069), .ZN(n9140) );
  OR2_X1 U9016 ( .A1(n9141), .A2(n9142), .ZN(n9069) );
  AND2_X1 U9017 ( .A1(n9066), .A2(n9065), .ZN(n9142) );
  AND2_X1 U9018 ( .A1(n9063), .A2(n9143), .ZN(n9141) );
  OR2_X1 U9019 ( .A1(n9066), .A2(n9065), .ZN(n9143) );
  OR2_X1 U9020 ( .A1(n9144), .A2(n9145), .ZN(n9065) );
  AND2_X1 U9021 ( .A1(n9062), .A2(n9061), .ZN(n9145) );
  AND2_X1 U9022 ( .A1(n9059), .A2(n9146), .ZN(n9144) );
  OR2_X1 U9023 ( .A1(n9062), .A2(n9061), .ZN(n9146) );
  OR2_X1 U9024 ( .A1(n9147), .A2(n9148), .ZN(n9061) );
  AND2_X1 U9025 ( .A1(n9058), .A2(n9057), .ZN(n9148) );
  AND2_X1 U9026 ( .A1(n9055), .A2(n9149), .ZN(n9147) );
  OR2_X1 U9027 ( .A1(n9058), .A2(n9057), .ZN(n9149) );
  OR2_X1 U9028 ( .A1(n9150), .A2(n9151), .ZN(n9057) );
  AND2_X1 U9029 ( .A1(n9054), .A2(n9053), .ZN(n9151) );
  AND2_X1 U9030 ( .A1(n9051), .A2(n9152), .ZN(n9150) );
  OR2_X1 U9031 ( .A1(n9054), .A2(n9053), .ZN(n9152) );
  OR2_X1 U9032 ( .A1(n9153), .A2(n9154), .ZN(n9053) );
  AND2_X1 U9033 ( .A1(n9050), .A2(n9049), .ZN(n9154) );
  AND2_X1 U9034 ( .A1(n9047), .A2(n9155), .ZN(n9153) );
  OR2_X1 U9035 ( .A1(n9050), .A2(n9049), .ZN(n9155) );
  OR2_X1 U9036 ( .A1(n9156), .A2(n9157), .ZN(n9049) );
  AND2_X1 U9037 ( .A1(n9046), .A2(n9045), .ZN(n9157) );
  AND2_X1 U9038 ( .A1(n9043), .A2(n9158), .ZN(n9156) );
  OR2_X1 U9039 ( .A1(n9046), .A2(n9045), .ZN(n9158) );
  OR2_X1 U9040 ( .A1(n9159), .A2(n9160), .ZN(n9045) );
  AND2_X1 U9041 ( .A1(n9042), .A2(n9041), .ZN(n9160) );
  AND2_X1 U9042 ( .A1(n9039), .A2(n9161), .ZN(n9159) );
  OR2_X1 U9043 ( .A1(n9042), .A2(n9041), .ZN(n9161) );
  OR2_X1 U9044 ( .A1(n9162), .A2(n9163), .ZN(n9041) );
  AND2_X1 U9045 ( .A1(n9038), .A2(n9037), .ZN(n9163) );
  AND2_X1 U9046 ( .A1(n9035), .A2(n9164), .ZN(n9162) );
  OR2_X1 U9047 ( .A1(n9038), .A2(n9037), .ZN(n9164) );
  OR2_X1 U9048 ( .A1(n9165), .A2(n9166), .ZN(n9037) );
  AND2_X1 U9049 ( .A1(n9034), .A2(n9033), .ZN(n9166) );
  AND2_X1 U9050 ( .A1(n9031), .A2(n9167), .ZN(n9165) );
  OR2_X1 U9051 ( .A1(n9034), .A2(n9033), .ZN(n9167) );
  OR2_X1 U9052 ( .A1(n9168), .A2(n9169), .ZN(n9033) );
  AND2_X1 U9053 ( .A1(n9030), .A2(n9029), .ZN(n9169) );
  AND2_X1 U9054 ( .A1(n9027), .A2(n9170), .ZN(n9168) );
  OR2_X1 U9055 ( .A1(n9030), .A2(n9029), .ZN(n9170) );
  OR2_X1 U9056 ( .A1(n9171), .A2(n9172), .ZN(n9029) );
  AND2_X1 U9057 ( .A1(n9026), .A2(n9025), .ZN(n9172) );
  AND2_X1 U9058 ( .A1(n9023), .A2(n9173), .ZN(n9171) );
  OR2_X1 U9059 ( .A1(n9026), .A2(n9025), .ZN(n9173) );
  OR2_X1 U9060 ( .A1(n9174), .A2(n9175), .ZN(n9025) );
  AND2_X1 U9061 ( .A1(n9022), .A2(n9021), .ZN(n9175) );
  AND2_X1 U9062 ( .A1(n9019), .A2(n9176), .ZN(n9174) );
  OR2_X1 U9063 ( .A1(n9022), .A2(n9021), .ZN(n9176) );
  OR2_X1 U9064 ( .A1(n9177), .A2(n9178), .ZN(n9021) );
  AND2_X1 U9065 ( .A1(n9018), .A2(n9017), .ZN(n9178) );
  AND2_X1 U9066 ( .A1(n9015), .A2(n9179), .ZN(n9177) );
  OR2_X1 U9067 ( .A1(n9018), .A2(n9017), .ZN(n9179) );
  OR2_X1 U9068 ( .A1(n9180), .A2(n9181), .ZN(n9017) );
  AND2_X1 U9069 ( .A1(n9014), .A2(n9013), .ZN(n9181) );
  AND2_X1 U9070 ( .A1(n9011), .A2(n9182), .ZN(n9180) );
  OR2_X1 U9071 ( .A1(n9014), .A2(n9013), .ZN(n9182) );
  OR2_X1 U9072 ( .A1(n9183), .A2(n9184), .ZN(n9013) );
  AND2_X1 U9073 ( .A1(n9010), .A2(n9009), .ZN(n9184) );
  AND2_X1 U9074 ( .A1(n9007), .A2(n9185), .ZN(n9183) );
  OR2_X1 U9075 ( .A1(n9010), .A2(n9009), .ZN(n9185) );
  OR2_X1 U9076 ( .A1(n9186), .A2(n9187), .ZN(n9009) );
  AND2_X1 U9077 ( .A1(n9006), .A2(n9005), .ZN(n9187) );
  AND2_X1 U9078 ( .A1(n9003), .A2(n9188), .ZN(n9186) );
  OR2_X1 U9079 ( .A1(n9006), .A2(n9005), .ZN(n9188) );
  OR2_X1 U9080 ( .A1(n9189), .A2(n9190), .ZN(n9005) );
  AND2_X1 U9081 ( .A1(n8999), .A2(n9002), .ZN(n9190) );
  AND2_X1 U9082 ( .A1(n9001), .A2(n9191), .ZN(n9189) );
  OR2_X1 U9083 ( .A1(n8999), .A2(n9002), .ZN(n9191) );
  OR3_X1 U9084 ( .A1(n8998), .A2(n8417), .A3(n8519), .ZN(n9002) );
  OR2_X1 U9085 ( .A1(n8417), .A2(n7606), .ZN(n8999) );
  INV_X1 U9086 ( .A(n9192), .ZN(n9001) );
  OR2_X1 U9087 ( .A1(n9193), .A2(n9194), .ZN(n9192) );
  AND2_X1 U9088 ( .A1(n9195), .A2(n9196), .ZN(n9194) );
  OR2_X1 U9089 ( .A1(n9197), .A2(n7697), .ZN(n9196) );
  AND2_X1 U9090 ( .A1(n8998), .A2(n7691), .ZN(n9197) );
  AND2_X1 U9091 ( .A1(n8993), .A2(n9198), .ZN(n9193) );
  OR2_X1 U9092 ( .A1(n9199), .A2(n7701), .ZN(n9198) );
  AND2_X1 U9093 ( .A1(n9200), .A2(n7703), .ZN(n9199) );
  OR2_X1 U9094 ( .A1(n7662), .A2(n8417), .ZN(n9006) );
  XNOR2_X1 U9095 ( .A(n9201), .B(n9202), .ZN(n9003) );
  XNOR2_X1 U9096 ( .A(n9203), .B(n9204), .ZN(n9202) );
  OR2_X1 U9097 ( .A1(n7660), .A2(n8417), .ZN(n9010) );
  XOR2_X1 U9098 ( .A(n9205), .B(n9206), .Z(n9007) );
  XOR2_X1 U9099 ( .A(n9207), .B(n9208), .Z(n9206) );
  OR2_X1 U9100 ( .A1(n7658), .A2(n8417), .ZN(n9014) );
  XOR2_X1 U9101 ( .A(n9209), .B(n9210), .Z(n9011) );
  XOR2_X1 U9102 ( .A(n9211), .B(n9212), .Z(n9210) );
  OR2_X1 U9103 ( .A1(n7656), .A2(n8417), .ZN(n9018) );
  XOR2_X1 U9104 ( .A(n9213), .B(n9214), .Z(n9015) );
  XOR2_X1 U9105 ( .A(n9215), .B(n9216), .Z(n9214) );
  OR2_X1 U9106 ( .A1(n7654), .A2(n8417), .ZN(n9022) );
  XOR2_X1 U9107 ( .A(n9217), .B(n9218), .Z(n9019) );
  XOR2_X1 U9108 ( .A(n9219), .B(n9220), .Z(n9218) );
  OR2_X1 U9109 ( .A1(n7652), .A2(n8417), .ZN(n9026) );
  XOR2_X1 U9110 ( .A(n9221), .B(n9222), .Z(n9023) );
  XOR2_X1 U9111 ( .A(n9223), .B(n9224), .Z(n9222) );
  OR2_X1 U9112 ( .A1(n7650), .A2(n8417), .ZN(n9030) );
  XOR2_X1 U9113 ( .A(n9225), .B(n9226), .Z(n9027) );
  XOR2_X1 U9114 ( .A(n9227), .B(n9228), .Z(n9226) );
  OR2_X1 U9115 ( .A1(n7648), .A2(n8417), .ZN(n9034) );
  XOR2_X1 U9116 ( .A(n9229), .B(n9230), .Z(n9031) );
  XOR2_X1 U9117 ( .A(n9231), .B(n9232), .Z(n9230) );
  OR2_X1 U9118 ( .A1(n7646), .A2(n8417), .ZN(n9038) );
  XOR2_X1 U9119 ( .A(n9233), .B(n9234), .Z(n9035) );
  XOR2_X1 U9120 ( .A(n9235), .B(n9236), .Z(n9234) );
  OR2_X1 U9121 ( .A1(n7644), .A2(n8417), .ZN(n9042) );
  XOR2_X1 U9122 ( .A(n9237), .B(n9238), .Z(n9039) );
  XOR2_X1 U9123 ( .A(n9239), .B(n9240), .Z(n9238) );
  OR2_X1 U9124 ( .A1(n7642), .A2(n8417), .ZN(n9046) );
  XOR2_X1 U9125 ( .A(n9241), .B(n9242), .Z(n9043) );
  XOR2_X1 U9126 ( .A(n9243), .B(n9244), .Z(n9242) );
  OR2_X1 U9127 ( .A1(n7640), .A2(n8417), .ZN(n9050) );
  XOR2_X1 U9128 ( .A(n9245), .B(n9246), .Z(n9047) );
  XOR2_X1 U9129 ( .A(n9247), .B(n9248), .Z(n9246) );
  OR2_X1 U9130 ( .A1(n7638), .A2(n8417), .ZN(n9054) );
  XOR2_X1 U9131 ( .A(n9249), .B(n9250), .Z(n9051) );
  XOR2_X1 U9132 ( .A(n9251), .B(n9252), .Z(n9250) );
  OR2_X1 U9133 ( .A1(n7636), .A2(n8417), .ZN(n9058) );
  XOR2_X1 U9134 ( .A(n9253), .B(n9254), .Z(n9055) );
  XOR2_X1 U9135 ( .A(n9255), .B(n9256), .Z(n9254) );
  OR2_X1 U9136 ( .A1(n7634), .A2(n8417), .ZN(n9062) );
  XOR2_X1 U9137 ( .A(n9257), .B(n9258), .Z(n9059) );
  XOR2_X1 U9138 ( .A(n9259), .B(n9260), .Z(n9258) );
  OR2_X1 U9139 ( .A1(n7632), .A2(n8417), .ZN(n9066) );
  XOR2_X1 U9140 ( .A(n9261), .B(n9262), .Z(n9063) );
  XOR2_X1 U9141 ( .A(n9263), .B(n9264), .Z(n9262) );
  OR2_X1 U9142 ( .A1(n7630), .A2(n8417), .ZN(n9070) );
  XOR2_X1 U9143 ( .A(n9265), .B(n9266), .Z(n9067) );
  XOR2_X1 U9144 ( .A(n9267), .B(n9268), .Z(n9266) );
  OR2_X1 U9145 ( .A1(n7628), .A2(n8417), .ZN(n9074) );
  XOR2_X1 U9146 ( .A(n9269), .B(n9270), .Z(n9071) );
  XOR2_X1 U9147 ( .A(n9271), .B(n9272), .Z(n9270) );
  OR2_X1 U9148 ( .A1(n7626), .A2(n8417), .ZN(n9078) );
  XOR2_X1 U9149 ( .A(n9273), .B(n9274), .Z(n9075) );
  XOR2_X1 U9150 ( .A(n9275), .B(n9276), .Z(n9274) );
  OR2_X1 U9151 ( .A1(n7624), .A2(n8417), .ZN(n9082) );
  XOR2_X1 U9152 ( .A(n9277), .B(n9278), .Z(n9079) );
  XOR2_X1 U9153 ( .A(n9279), .B(n9280), .Z(n9278) );
  OR2_X1 U9154 ( .A1(n7622), .A2(n8417), .ZN(n9086) );
  XOR2_X1 U9155 ( .A(n9281), .B(n9282), .Z(n9083) );
  XOR2_X1 U9156 ( .A(n9283), .B(n9284), .Z(n9282) );
  OR2_X1 U9157 ( .A1(n7620), .A2(n8417), .ZN(n9090) );
  XOR2_X1 U9158 ( .A(n9285), .B(n9286), .Z(n9087) );
  XOR2_X1 U9159 ( .A(n9287), .B(n9288), .Z(n9286) );
  OR2_X1 U9160 ( .A1(n7618), .A2(n8417), .ZN(n9094) );
  XOR2_X1 U9161 ( .A(n9289), .B(n9290), .Z(n9091) );
  XOR2_X1 U9162 ( .A(n9291), .B(n9292), .Z(n9290) );
  OR2_X1 U9163 ( .A1(n7616), .A2(n8417), .ZN(n9098) );
  XOR2_X1 U9164 ( .A(n9293), .B(n9294), .Z(n9095) );
  XOR2_X1 U9165 ( .A(n9295), .B(n9296), .Z(n9294) );
  OR2_X1 U9166 ( .A1(n7614), .A2(n8417), .ZN(n9105) );
  XOR2_X1 U9167 ( .A(n9297), .B(n9298), .Z(n9102) );
  XOR2_X1 U9168 ( .A(n9299), .B(n9300), .Z(n9298) );
  OR2_X1 U9169 ( .A1(n7612), .A2(n8417), .ZN(n9109) );
  XOR2_X1 U9170 ( .A(n9301), .B(n9302), .Z(n9106) );
  XOR2_X1 U9171 ( .A(n9303), .B(n9304), .Z(n9302) );
  OR2_X1 U9172 ( .A1(n7610), .A2(n8417), .ZN(n8689) );
  INV_X1 U9173 ( .A(n8787), .ZN(n8417) );
  XOR2_X1 U9174 ( .A(n9305), .B(n9306), .Z(n8787) );
  XNOR2_X1 U9175 ( .A(c_28_), .B(d_28_), .ZN(n9305) );
  XOR2_X1 U9176 ( .A(n9307), .B(n9308), .Z(n8690) );
  XOR2_X1 U9177 ( .A(n9309), .B(n9310), .Z(n9308) );
  AND2_X1 U9178 ( .A1(n8378), .A2(n8377), .ZN(n7871) );
  XNOR2_X1 U9179 ( .A(n8347), .B(n8349), .ZN(n8377) );
  OR2_X1 U9180 ( .A1(n9311), .A2(n9312), .ZN(n8349) );
  AND2_X1 U9181 ( .A1(n9313), .A2(n9314), .ZN(n9312) );
  AND2_X1 U9182 ( .A1(n9315), .A2(n9316), .ZN(n9311) );
  OR2_X1 U9183 ( .A1(n9313), .A2(n9314), .ZN(n9316) );
  XOR2_X1 U9184 ( .A(n8355), .B(n9317), .Z(n8347) );
  XOR2_X1 U9185 ( .A(n8354), .B(n8353), .Z(n9317) );
  OR2_X1 U9186 ( .A1(n9318), .A2(n7664), .ZN(n8353) );
  OR2_X1 U9187 ( .A1(n9319), .A2(n9320), .ZN(n8354) );
  AND2_X1 U9188 ( .A1(n9321), .A2(n9322), .ZN(n9320) );
  AND2_X1 U9189 ( .A1(n9323), .A2(n9324), .ZN(n9319) );
  OR2_X1 U9190 ( .A1(n9321), .A2(n9322), .ZN(n9324) );
  XNOR2_X1 U9191 ( .A(n9325), .B(n8363), .ZN(n8355) );
  XOR2_X1 U9192 ( .A(n8370), .B(n9326), .Z(n8363) );
  XOR2_X1 U9193 ( .A(n8369), .B(n8368), .Z(n9326) );
  OR2_X1 U9194 ( .A1(n8056), .A2(n8335), .ZN(n8368) );
  OR2_X1 U9195 ( .A1(n9327), .A2(n9328), .ZN(n8369) );
  AND2_X1 U9196 ( .A1(n9329), .A2(n9330), .ZN(n9328) );
  AND2_X1 U9197 ( .A1(n9331), .A2(n9332), .ZN(n9327) );
  OR2_X1 U9198 ( .A1(n9329), .A2(n9330), .ZN(n9332) );
  XOR2_X1 U9199 ( .A(n9333), .B(n9334), .Z(n8370) );
  XOR2_X1 U9200 ( .A(n9335), .B(n9336), .Z(n9334) );
  XNOR2_X1 U9201 ( .A(n8361), .B(n8362), .ZN(n9325) );
  OR2_X1 U9202 ( .A1(n8023), .A2(n8358), .ZN(n8362) );
  OR2_X1 U9203 ( .A1(n9337), .A2(n9338), .ZN(n8361) );
  AND2_X1 U9204 ( .A1(n9339), .A2(n9340), .ZN(n9338) );
  AND2_X1 U9205 ( .A1(n9341), .A2(n9342), .ZN(n9337) );
  OR2_X1 U9206 ( .A1(n9339), .A2(n9340), .ZN(n9342) );
  OR2_X1 U9207 ( .A1(n8384), .A2(n8385), .ZN(n8378) );
  OR2_X1 U9208 ( .A1(n9343), .A2(n9344), .ZN(n8385) );
  AND2_X1 U9209 ( .A1(n8397), .A2(n8400), .ZN(n9344) );
  AND2_X1 U9210 ( .A1(n9345), .A2(n8399), .ZN(n9343) );
  OR2_X1 U9211 ( .A1(n9346), .A2(n9347), .ZN(n8399) );
  AND2_X1 U9212 ( .A1(n8427), .A2(n8426), .ZN(n9347) );
  AND2_X1 U9213 ( .A1(n8424), .A2(n9348), .ZN(n9346) );
  OR2_X1 U9214 ( .A1(n8426), .A2(n8427), .ZN(n9348) );
  OR2_X1 U9215 ( .A1(n8023), .A2(n8998), .ZN(n8427) );
  OR2_X1 U9216 ( .A1(n9349), .A2(n9350), .ZN(n8426) );
  AND2_X1 U9217 ( .A1(n8695), .A2(n8694), .ZN(n9350) );
  AND2_X1 U9218 ( .A1(n8692), .A2(n9351), .ZN(n9349) );
  OR2_X1 U9219 ( .A1(n8694), .A2(n8695), .ZN(n9351) );
  OR2_X1 U9220 ( .A1(n9352), .A2(n9353), .ZN(n8695) );
  AND2_X1 U9221 ( .A1(n9310), .A2(n9309), .ZN(n9353) );
  AND2_X1 U9222 ( .A1(n9307), .A2(n9354), .ZN(n9352) );
  OR2_X1 U9223 ( .A1(n9309), .A2(n9310), .ZN(n9354) );
  OR2_X1 U9224 ( .A1(n7612), .A2(n8998), .ZN(n9310) );
  OR2_X1 U9225 ( .A1(n9355), .A2(n9356), .ZN(n9309) );
  AND2_X1 U9226 ( .A1(n9304), .A2(n9303), .ZN(n9356) );
  AND2_X1 U9227 ( .A1(n9301), .A2(n9357), .ZN(n9355) );
  OR2_X1 U9228 ( .A1(n9303), .A2(n9304), .ZN(n9357) );
  OR2_X1 U9229 ( .A1(n7614), .A2(n8998), .ZN(n9304) );
  OR2_X1 U9230 ( .A1(n9358), .A2(n9359), .ZN(n9303) );
  AND2_X1 U9231 ( .A1(n9300), .A2(n9299), .ZN(n9359) );
  AND2_X1 U9232 ( .A1(n9297), .A2(n9360), .ZN(n9358) );
  OR2_X1 U9233 ( .A1(n9299), .A2(n9300), .ZN(n9360) );
  OR2_X1 U9234 ( .A1(n7616), .A2(n8998), .ZN(n9300) );
  OR2_X1 U9235 ( .A1(n9361), .A2(n9362), .ZN(n9299) );
  AND2_X1 U9236 ( .A1(n9296), .A2(n9295), .ZN(n9362) );
  AND2_X1 U9237 ( .A1(n9293), .A2(n9363), .ZN(n9361) );
  OR2_X1 U9238 ( .A1(n9295), .A2(n9296), .ZN(n9363) );
  OR2_X1 U9239 ( .A1(n9364), .A2(n9365), .ZN(n9296) );
  AND2_X1 U9240 ( .A1(n9292), .A2(n9291), .ZN(n9365) );
  AND2_X1 U9241 ( .A1(n9289), .A2(n9366), .ZN(n9364) );
  OR2_X1 U9242 ( .A1(n9291), .A2(n9292), .ZN(n9366) );
  OR2_X1 U9243 ( .A1(n7620), .A2(n8998), .ZN(n9292) );
  OR2_X1 U9244 ( .A1(n9367), .A2(n9368), .ZN(n9291) );
  AND2_X1 U9245 ( .A1(n9288), .A2(n9287), .ZN(n9368) );
  AND2_X1 U9246 ( .A1(n9285), .A2(n9369), .ZN(n9367) );
  OR2_X1 U9247 ( .A1(n9287), .A2(n9288), .ZN(n9369) );
  OR2_X1 U9248 ( .A1(n7622), .A2(n8998), .ZN(n9288) );
  OR2_X1 U9249 ( .A1(n9370), .A2(n9371), .ZN(n9287) );
  AND2_X1 U9250 ( .A1(n9284), .A2(n9283), .ZN(n9371) );
  AND2_X1 U9251 ( .A1(n9281), .A2(n9372), .ZN(n9370) );
  OR2_X1 U9252 ( .A1(n9283), .A2(n9284), .ZN(n9372) );
  OR2_X1 U9253 ( .A1(n7624), .A2(n8998), .ZN(n9284) );
  OR2_X1 U9254 ( .A1(n9373), .A2(n9374), .ZN(n9283) );
  AND2_X1 U9255 ( .A1(n9280), .A2(n9279), .ZN(n9374) );
  AND2_X1 U9256 ( .A1(n9277), .A2(n9375), .ZN(n9373) );
  OR2_X1 U9257 ( .A1(n9279), .A2(n9280), .ZN(n9375) );
  OR2_X1 U9258 ( .A1(n7626), .A2(n8998), .ZN(n9280) );
  OR2_X1 U9259 ( .A1(n9376), .A2(n9377), .ZN(n9279) );
  AND2_X1 U9260 ( .A1(n9276), .A2(n9275), .ZN(n9377) );
  AND2_X1 U9261 ( .A1(n9273), .A2(n9378), .ZN(n9376) );
  OR2_X1 U9262 ( .A1(n9275), .A2(n9276), .ZN(n9378) );
  OR2_X1 U9263 ( .A1(n7628), .A2(n8998), .ZN(n9276) );
  OR2_X1 U9264 ( .A1(n9379), .A2(n9380), .ZN(n9275) );
  AND2_X1 U9265 ( .A1(n9272), .A2(n9271), .ZN(n9380) );
  AND2_X1 U9266 ( .A1(n9269), .A2(n9381), .ZN(n9379) );
  OR2_X1 U9267 ( .A1(n9271), .A2(n9272), .ZN(n9381) );
  OR2_X1 U9268 ( .A1(n7630), .A2(n8998), .ZN(n9272) );
  OR2_X1 U9269 ( .A1(n9382), .A2(n9383), .ZN(n9271) );
  AND2_X1 U9270 ( .A1(n9268), .A2(n9267), .ZN(n9383) );
  AND2_X1 U9271 ( .A1(n9265), .A2(n9384), .ZN(n9382) );
  OR2_X1 U9272 ( .A1(n9267), .A2(n9268), .ZN(n9384) );
  OR2_X1 U9273 ( .A1(n7632), .A2(n8998), .ZN(n9268) );
  OR2_X1 U9274 ( .A1(n9385), .A2(n9386), .ZN(n9267) );
  AND2_X1 U9275 ( .A1(n9264), .A2(n9263), .ZN(n9386) );
  AND2_X1 U9276 ( .A1(n9261), .A2(n9387), .ZN(n9385) );
  OR2_X1 U9277 ( .A1(n9263), .A2(n9264), .ZN(n9387) );
  OR2_X1 U9278 ( .A1(n7634), .A2(n8998), .ZN(n9264) );
  OR2_X1 U9279 ( .A1(n9388), .A2(n9389), .ZN(n9263) );
  AND2_X1 U9280 ( .A1(n9260), .A2(n9259), .ZN(n9389) );
  AND2_X1 U9281 ( .A1(n9257), .A2(n9390), .ZN(n9388) );
  OR2_X1 U9282 ( .A1(n9259), .A2(n9260), .ZN(n9390) );
  OR2_X1 U9283 ( .A1(n7636), .A2(n8998), .ZN(n9260) );
  OR2_X1 U9284 ( .A1(n9391), .A2(n9392), .ZN(n9259) );
  AND2_X1 U9285 ( .A1(n9256), .A2(n9255), .ZN(n9392) );
  AND2_X1 U9286 ( .A1(n9253), .A2(n9393), .ZN(n9391) );
  OR2_X1 U9287 ( .A1(n9255), .A2(n9256), .ZN(n9393) );
  OR2_X1 U9288 ( .A1(n7638), .A2(n8998), .ZN(n9256) );
  OR2_X1 U9289 ( .A1(n9394), .A2(n9395), .ZN(n9255) );
  AND2_X1 U9290 ( .A1(n9252), .A2(n9251), .ZN(n9395) );
  AND2_X1 U9291 ( .A1(n9249), .A2(n9396), .ZN(n9394) );
  OR2_X1 U9292 ( .A1(n9251), .A2(n9252), .ZN(n9396) );
  OR2_X1 U9293 ( .A1(n7640), .A2(n8998), .ZN(n9252) );
  OR2_X1 U9294 ( .A1(n9397), .A2(n9398), .ZN(n9251) );
  AND2_X1 U9295 ( .A1(n9248), .A2(n9247), .ZN(n9398) );
  AND2_X1 U9296 ( .A1(n9245), .A2(n9399), .ZN(n9397) );
  OR2_X1 U9297 ( .A1(n9247), .A2(n9248), .ZN(n9399) );
  OR2_X1 U9298 ( .A1(n7642), .A2(n8998), .ZN(n9248) );
  OR2_X1 U9299 ( .A1(n9400), .A2(n9401), .ZN(n9247) );
  AND2_X1 U9300 ( .A1(n9244), .A2(n9243), .ZN(n9401) );
  AND2_X1 U9301 ( .A1(n9241), .A2(n9402), .ZN(n9400) );
  OR2_X1 U9302 ( .A1(n9243), .A2(n9244), .ZN(n9402) );
  OR2_X1 U9303 ( .A1(n7644), .A2(n8998), .ZN(n9244) );
  OR2_X1 U9304 ( .A1(n9403), .A2(n9404), .ZN(n9243) );
  AND2_X1 U9305 ( .A1(n9240), .A2(n9239), .ZN(n9404) );
  AND2_X1 U9306 ( .A1(n9237), .A2(n9405), .ZN(n9403) );
  OR2_X1 U9307 ( .A1(n9239), .A2(n9240), .ZN(n9405) );
  OR2_X1 U9308 ( .A1(n7646), .A2(n8998), .ZN(n9240) );
  OR2_X1 U9309 ( .A1(n9406), .A2(n9407), .ZN(n9239) );
  AND2_X1 U9310 ( .A1(n9236), .A2(n9235), .ZN(n9407) );
  AND2_X1 U9311 ( .A1(n9233), .A2(n9408), .ZN(n9406) );
  OR2_X1 U9312 ( .A1(n9235), .A2(n9236), .ZN(n9408) );
  OR2_X1 U9313 ( .A1(n7648), .A2(n8998), .ZN(n9236) );
  OR2_X1 U9314 ( .A1(n9409), .A2(n9410), .ZN(n9235) );
  AND2_X1 U9315 ( .A1(n9232), .A2(n9231), .ZN(n9410) );
  AND2_X1 U9316 ( .A1(n9229), .A2(n9411), .ZN(n9409) );
  OR2_X1 U9317 ( .A1(n9231), .A2(n9232), .ZN(n9411) );
  OR2_X1 U9318 ( .A1(n7650), .A2(n8998), .ZN(n9232) );
  OR2_X1 U9319 ( .A1(n9412), .A2(n9413), .ZN(n9231) );
  AND2_X1 U9320 ( .A1(n9228), .A2(n9227), .ZN(n9413) );
  AND2_X1 U9321 ( .A1(n9225), .A2(n9414), .ZN(n9412) );
  OR2_X1 U9322 ( .A1(n9227), .A2(n9228), .ZN(n9414) );
  OR2_X1 U9323 ( .A1(n7652), .A2(n8998), .ZN(n9228) );
  OR2_X1 U9324 ( .A1(n9415), .A2(n9416), .ZN(n9227) );
  AND2_X1 U9325 ( .A1(n9224), .A2(n9223), .ZN(n9416) );
  AND2_X1 U9326 ( .A1(n9221), .A2(n9417), .ZN(n9415) );
  OR2_X1 U9327 ( .A1(n9223), .A2(n9224), .ZN(n9417) );
  OR2_X1 U9328 ( .A1(n7654), .A2(n8998), .ZN(n9224) );
  OR2_X1 U9329 ( .A1(n9418), .A2(n9419), .ZN(n9223) );
  AND2_X1 U9330 ( .A1(n9220), .A2(n9219), .ZN(n9419) );
  AND2_X1 U9331 ( .A1(n9217), .A2(n9420), .ZN(n9418) );
  OR2_X1 U9332 ( .A1(n9219), .A2(n9220), .ZN(n9420) );
  OR2_X1 U9333 ( .A1(n7656), .A2(n8998), .ZN(n9220) );
  OR2_X1 U9334 ( .A1(n9421), .A2(n9422), .ZN(n9219) );
  AND2_X1 U9335 ( .A1(n9216), .A2(n9215), .ZN(n9422) );
  AND2_X1 U9336 ( .A1(n9213), .A2(n9423), .ZN(n9421) );
  OR2_X1 U9337 ( .A1(n9215), .A2(n9216), .ZN(n9423) );
  OR2_X1 U9338 ( .A1(n7658), .A2(n8998), .ZN(n9216) );
  OR2_X1 U9339 ( .A1(n9424), .A2(n9425), .ZN(n9215) );
  AND2_X1 U9340 ( .A1(n9212), .A2(n9211), .ZN(n9425) );
  AND2_X1 U9341 ( .A1(n9209), .A2(n9426), .ZN(n9424) );
  OR2_X1 U9342 ( .A1(n9211), .A2(n9212), .ZN(n9426) );
  OR2_X1 U9343 ( .A1(n7660), .A2(n8998), .ZN(n9212) );
  OR2_X1 U9344 ( .A1(n9427), .A2(n9428), .ZN(n9211) );
  AND2_X1 U9345 ( .A1(n9208), .A2(n9207), .ZN(n9428) );
  AND2_X1 U9346 ( .A1(n9205), .A2(n9429), .ZN(n9427) );
  OR2_X1 U9347 ( .A1(n9207), .A2(n9208), .ZN(n9429) );
  OR2_X1 U9348 ( .A1(n7662), .A2(n8998), .ZN(n9208) );
  OR2_X1 U9349 ( .A1(n9430), .A2(n9431), .ZN(n9207) );
  AND2_X1 U9350 ( .A1(n9201), .A2(n9204), .ZN(n9431) );
  AND2_X1 U9351 ( .A1(n9203), .A2(n9432), .ZN(n9430) );
  OR2_X1 U9352 ( .A1(n9204), .A2(n9201), .ZN(n9432) );
  OR2_X1 U9353 ( .A1(n8998), .A2(n7606), .ZN(n9201) );
  OR3_X1 U9354 ( .A1(n9200), .A2(n8998), .A3(n8519), .ZN(n9204) );
  INV_X1 U9355 ( .A(n9433), .ZN(n9203) );
  OR2_X1 U9356 ( .A1(n9434), .A2(n9435), .ZN(n9433) );
  AND2_X1 U9357 ( .A1(n9436), .A2(n9437), .ZN(n9435) );
  OR2_X1 U9358 ( .A1(n9438), .A2(n7697), .ZN(n9437) );
  AND2_X1 U9359 ( .A1(n9200), .A2(n7691), .ZN(n9438) );
  AND2_X1 U9360 ( .A1(n9195), .A2(n9439), .ZN(n9434) );
  OR2_X1 U9361 ( .A1(n9440), .A2(n7701), .ZN(n9439) );
  AND2_X1 U9362 ( .A1(n9318), .A2(n7703), .ZN(n9440) );
  XNOR2_X1 U9363 ( .A(n9441), .B(n9442), .ZN(n9205) );
  XNOR2_X1 U9364 ( .A(n9443), .B(n9444), .ZN(n9442) );
  XOR2_X1 U9365 ( .A(n9445), .B(n9446), .Z(n9209) );
  XOR2_X1 U9366 ( .A(n9447), .B(n9448), .Z(n9446) );
  XOR2_X1 U9367 ( .A(n9449), .B(n9450), .Z(n9213) );
  XOR2_X1 U9368 ( .A(n9451), .B(n9452), .Z(n9450) );
  XOR2_X1 U9369 ( .A(n9453), .B(n9454), .Z(n9217) );
  XOR2_X1 U9370 ( .A(n9455), .B(n9456), .Z(n9454) );
  XOR2_X1 U9371 ( .A(n9457), .B(n9458), .Z(n9221) );
  XOR2_X1 U9372 ( .A(n9459), .B(n9460), .Z(n9458) );
  XOR2_X1 U9373 ( .A(n9461), .B(n9462), .Z(n9225) );
  XOR2_X1 U9374 ( .A(n9463), .B(n9464), .Z(n9462) );
  XOR2_X1 U9375 ( .A(n9465), .B(n9466), .Z(n9229) );
  XOR2_X1 U9376 ( .A(n9467), .B(n9468), .Z(n9466) );
  XOR2_X1 U9377 ( .A(n9469), .B(n9470), .Z(n9233) );
  XOR2_X1 U9378 ( .A(n9471), .B(n9472), .Z(n9470) );
  XOR2_X1 U9379 ( .A(n9473), .B(n9474), .Z(n9237) );
  XOR2_X1 U9380 ( .A(n9475), .B(n9476), .Z(n9474) );
  XOR2_X1 U9381 ( .A(n9477), .B(n9478), .Z(n9241) );
  XOR2_X1 U9382 ( .A(n9479), .B(n9480), .Z(n9478) );
  XOR2_X1 U9383 ( .A(n9481), .B(n9482), .Z(n9245) );
  XOR2_X1 U9384 ( .A(n9483), .B(n9484), .Z(n9482) );
  XOR2_X1 U9385 ( .A(n9485), .B(n9486), .Z(n9249) );
  XOR2_X1 U9386 ( .A(n9487), .B(n9488), .Z(n9486) );
  XOR2_X1 U9387 ( .A(n9489), .B(n9490), .Z(n9253) );
  XOR2_X1 U9388 ( .A(n9491), .B(n9492), .Z(n9490) );
  XOR2_X1 U9389 ( .A(n9493), .B(n9494), .Z(n9257) );
  XOR2_X1 U9390 ( .A(n9495), .B(n9496), .Z(n9494) );
  XOR2_X1 U9391 ( .A(n9497), .B(n9498), .Z(n9261) );
  XOR2_X1 U9392 ( .A(n9499), .B(n9500), .Z(n9498) );
  XOR2_X1 U9393 ( .A(n9501), .B(n9502), .Z(n9265) );
  XOR2_X1 U9394 ( .A(n9503), .B(n9504), .Z(n9502) );
  XOR2_X1 U9395 ( .A(n9505), .B(n9506), .Z(n9269) );
  XOR2_X1 U9396 ( .A(n9507), .B(n9508), .Z(n9506) );
  XOR2_X1 U9397 ( .A(n9509), .B(n9510), .Z(n9273) );
  XOR2_X1 U9398 ( .A(n9511), .B(n9512), .Z(n9510) );
  XOR2_X1 U9399 ( .A(n9513), .B(n9514), .Z(n9277) );
  XOR2_X1 U9400 ( .A(n9515), .B(n9516), .Z(n9514) );
  XOR2_X1 U9401 ( .A(n9517), .B(n9518), .Z(n9281) );
  XOR2_X1 U9402 ( .A(n9519), .B(n9520), .Z(n9518) );
  XOR2_X1 U9403 ( .A(n9521), .B(n9522), .Z(n9285) );
  XOR2_X1 U9404 ( .A(n9523), .B(n9524), .Z(n9522) );
  XOR2_X1 U9405 ( .A(n9525), .B(n9526), .Z(n9289) );
  XOR2_X1 U9406 ( .A(n9527), .B(n9528), .Z(n9526) );
  OR2_X1 U9407 ( .A1(n7618), .A2(n8998), .ZN(n9295) );
  XOR2_X1 U9408 ( .A(n9529), .B(n9530), .Z(n9293) );
  XOR2_X1 U9409 ( .A(n9531), .B(n9532), .Z(n9530) );
  XOR2_X1 U9410 ( .A(n9533), .B(n9534), .Z(n9297) );
  XOR2_X1 U9411 ( .A(n9535), .B(n9536), .Z(n9534) );
  XOR2_X1 U9412 ( .A(n9537), .B(n9538), .Z(n9301) );
  XOR2_X1 U9413 ( .A(n9539), .B(n9540), .Z(n9538) );
  XOR2_X1 U9414 ( .A(n9541), .B(n9542), .Z(n9307) );
  XOR2_X1 U9415 ( .A(n9543), .B(n9544), .Z(n9542) );
  OR2_X1 U9416 ( .A1(n8056), .A2(n8998), .ZN(n8694) );
  XOR2_X1 U9417 ( .A(n9545), .B(n9546), .Z(n8692) );
  XOR2_X1 U9418 ( .A(n9547), .B(n9548), .Z(n9546) );
  XOR2_X1 U9419 ( .A(n9549), .B(n9550), .Z(n8424) );
  XOR2_X1 U9420 ( .A(n9551), .B(n9552), .Z(n9550) );
  OR2_X1 U9421 ( .A1(n8397), .A2(n8400), .ZN(n9345) );
  OR2_X1 U9422 ( .A1(n8998), .A2(n7664), .ZN(n8400) );
  INV_X1 U9423 ( .A(n8993), .ZN(n8998) );
  XOR2_X1 U9424 ( .A(n9553), .B(n9554), .Z(n8993) );
  XNOR2_X1 U9425 ( .A(c_27_), .B(d_27_), .ZN(n9553) );
  XOR2_X1 U9426 ( .A(n9555), .B(n9556), .Z(n8397) );
  XOR2_X1 U9427 ( .A(n9557), .B(n9558), .Z(n9556) );
  XOR2_X1 U9428 ( .A(n9315), .B(n9559), .Z(n8384) );
  XOR2_X1 U9429 ( .A(n9314), .B(n9313), .Z(n9559) );
  OR2_X1 U9430 ( .A1(n9200), .A2(n7664), .ZN(n9313) );
  OR2_X1 U9431 ( .A1(n9560), .A2(n9561), .ZN(n9314) );
  AND2_X1 U9432 ( .A1(n9558), .A2(n9557), .ZN(n9561) );
  AND2_X1 U9433 ( .A1(n9555), .A2(n9562), .ZN(n9560) );
  OR2_X1 U9434 ( .A1(n9558), .A2(n9557), .ZN(n9562) );
  OR2_X1 U9435 ( .A1(n9563), .A2(n9564), .ZN(n9557) );
  AND2_X1 U9436 ( .A1(n9552), .A2(n9551), .ZN(n9564) );
  AND2_X1 U9437 ( .A1(n9549), .A2(n9565), .ZN(n9563) );
  OR2_X1 U9438 ( .A1(n9552), .A2(n9551), .ZN(n9565) );
  OR2_X1 U9439 ( .A1(n9566), .A2(n9567), .ZN(n9551) );
  AND2_X1 U9440 ( .A1(n9548), .A2(n9547), .ZN(n9567) );
  AND2_X1 U9441 ( .A1(n9545), .A2(n9568), .ZN(n9566) );
  OR2_X1 U9442 ( .A1(n9548), .A2(n9547), .ZN(n9568) );
  OR2_X1 U9443 ( .A1(n9569), .A2(n9570), .ZN(n9547) );
  AND2_X1 U9444 ( .A1(n9544), .A2(n9543), .ZN(n9570) );
  AND2_X1 U9445 ( .A1(n9541), .A2(n9571), .ZN(n9569) );
  OR2_X1 U9446 ( .A1(n9544), .A2(n9543), .ZN(n9571) );
  OR2_X1 U9447 ( .A1(n9572), .A2(n9573), .ZN(n9543) );
  AND2_X1 U9448 ( .A1(n9540), .A2(n9539), .ZN(n9573) );
  AND2_X1 U9449 ( .A1(n9537), .A2(n9574), .ZN(n9572) );
  OR2_X1 U9450 ( .A1(n9540), .A2(n9539), .ZN(n9574) );
  OR2_X1 U9451 ( .A1(n9575), .A2(n9576), .ZN(n9539) );
  AND2_X1 U9452 ( .A1(n9536), .A2(n9535), .ZN(n9576) );
  AND2_X1 U9453 ( .A1(n9533), .A2(n9577), .ZN(n9575) );
  OR2_X1 U9454 ( .A1(n9536), .A2(n9535), .ZN(n9577) );
  OR2_X1 U9455 ( .A1(n7618), .A2(n9200), .ZN(n9535) );
  OR2_X1 U9456 ( .A1(n9578), .A2(n9579), .ZN(n9536) );
  AND2_X1 U9457 ( .A1(n9532), .A2(n9531), .ZN(n9579) );
  AND2_X1 U9458 ( .A1(n9529), .A2(n9580), .ZN(n9578) );
  OR2_X1 U9459 ( .A1(n9532), .A2(n9531), .ZN(n9580) );
  OR2_X1 U9460 ( .A1(n9581), .A2(n9582), .ZN(n9531) );
  AND2_X1 U9461 ( .A1(n9528), .A2(n9527), .ZN(n9582) );
  AND2_X1 U9462 ( .A1(n9525), .A2(n9583), .ZN(n9581) );
  OR2_X1 U9463 ( .A1(n9528), .A2(n9527), .ZN(n9583) );
  OR2_X1 U9464 ( .A1(n9584), .A2(n9585), .ZN(n9527) );
  AND2_X1 U9465 ( .A1(n9524), .A2(n9523), .ZN(n9585) );
  AND2_X1 U9466 ( .A1(n9521), .A2(n9586), .ZN(n9584) );
  OR2_X1 U9467 ( .A1(n9524), .A2(n9523), .ZN(n9586) );
  OR2_X1 U9468 ( .A1(n9587), .A2(n9588), .ZN(n9523) );
  AND2_X1 U9469 ( .A1(n9520), .A2(n9519), .ZN(n9588) );
  AND2_X1 U9470 ( .A1(n9517), .A2(n9589), .ZN(n9587) );
  OR2_X1 U9471 ( .A1(n9520), .A2(n9519), .ZN(n9589) );
  OR2_X1 U9472 ( .A1(n9590), .A2(n9591), .ZN(n9519) );
  AND2_X1 U9473 ( .A1(n9516), .A2(n9515), .ZN(n9591) );
  AND2_X1 U9474 ( .A1(n9513), .A2(n9592), .ZN(n9590) );
  OR2_X1 U9475 ( .A1(n9516), .A2(n9515), .ZN(n9592) );
  OR2_X1 U9476 ( .A1(n9593), .A2(n9594), .ZN(n9515) );
  AND2_X1 U9477 ( .A1(n9512), .A2(n9511), .ZN(n9594) );
  AND2_X1 U9478 ( .A1(n9509), .A2(n9595), .ZN(n9593) );
  OR2_X1 U9479 ( .A1(n9512), .A2(n9511), .ZN(n9595) );
  OR2_X1 U9480 ( .A1(n9596), .A2(n9597), .ZN(n9511) );
  AND2_X1 U9481 ( .A1(n9508), .A2(n9507), .ZN(n9597) );
  AND2_X1 U9482 ( .A1(n9505), .A2(n9598), .ZN(n9596) );
  OR2_X1 U9483 ( .A1(n9508), .A2(n9507), .ZN(n9598) );
  OR2_X1 U9484 ( .A1(n9599), .A2(n9600), .ZN(n9507) );
  AND2_X1 U9485 ( .A1(n9504), .A2(n9503), .ZN(n9600) );
  AND2_X1 U9486 ( .A1(n9501), .A2(n9601), .ZN(n9599) );
  OR2_X1 U9487 ( .A1(n9504), .A2(n9503), .ZN(n9601) );
  OR2_X1 U9488 ( .A1(n9602), .A2(n9603), .ZN(n9503) );
  AND2_X1 U9489 ( .A1(n9500), .A2(n9499), .ZN(n9603) );
  AND2_X1 U9490 ( .A1(n9497), .A2(n9604), .ZN(n9602) );
  OR2_X1 U9491 ( .A1(n9500), .A2(n9499), .ZN(n9604) );
  OR2_X1 U9492 ( .A1(n9605), .A2(n9606), .ZN(n9499) );
  AND2_X1 U9493 ( .A1(n9496), .A2(n9495), .ZN(n9606) );
  AND2_X1 U9494 ( .A1(n9493), .A2(n9607), .ZN(n9605) );
  OR2_X1 U9495 ( .A1(n9496), .A2(n9495), .ZN(n9607) );
  OR2_X1 U9496 ( .A1(n9608), .A2(n9609), .ZN(n9495) );
  AND2_X1 U9497 ( .A1(n9492), .A2(n9491), .ZN(n9609) );
  AND2_X1 U9498 ( .A1(n9489), .A2(n9610), .ZN(n9608) );
  OR2_X1 U9499 ( .A1(n9492), .A2(n9491), .ZN(n9610) );
  OR2_X1 U9500 ( .A1(n9611), .A2(n9612), .ZN(n9491) );
  AND2_X1 U9501 ( .A1(n9488), .A2(n9487), .ZN(n9612) );
  AND2_X1 U9502 ( .A1(n9485), .A2(n9613), .ZN(n9611) );
  OR2_X1 U9503 ( .A1(n9488), .A2(n9487), .ZN(n9613) );
  OR2_X1 U9504 ( .A1(n9614), .A2(n9615), .ZN(n9487) );
  AND2_X1 U9505 ( .A1(n9484), .A2(n9483), .ZN(n9615) );
  AND2_X1 U9506 ( .A1(n9481), .A2(n9616), .ZN(n9614) );
  OR2_X1 U9507 ( .A1(n9484), .A2(n9483), .ZN(n9616) );
  OR2_X1 U9508 ( .A1(n9617), .A2(n9618), .ZN(n9483) );
  AND2_X1 U9509 ( .A1(n9480), .A2(n9479), .ZN(n9618) );
  AND2_X1 U9510 ( .A1(n9477), .A2(n9619), .ZN(n9617) );
  OR2_X1 U9511 ( .A1(n9480), .A2(n9479), .ZN(n9619) );
  OR2_X1 U9512 ( .A1(n9620), .A2(n9621), .ZN(n9479) );
  AND2_X1 U9513 ( .A1(n9476), .A2(n9475), .ZN(n9621) );
  AND2_X1 U9514 ( .A1(n9473), .A2(n9622), .ZN(n9620) );
  OR2_X1 U9515 ( .A1(n9476), .A2(n9475), .ZN(n9622) );
  OR2_X1 U9516 ( .A1(n9623), .A2(n9624), .ZN(n9475) );
  AND2_X1 U9517 ( .A1(n9472), .A2(n9471), .ZN(n9624) );
  AND2_X1 U9518 ( .A1(n9469), .A2(n9625), .ZN(n9623) );
  OR2_X1 U9519 ( .A1(n9472), .A2(n9471), .ZN(n9625) );
  OR2_X1 U9520 ( .A1(n9626), .A2(n9627), .ZN(n9471) );
  AND2_X1 U9521 ( .A1(n9468), .A2(n9467), .ZN(n9627) );
  AND2_X1 U9522 ( .A1(n9465), .A2(n9628), .ZN(n9626) );
  OR2_X1 U9523 ( .A1(n9468), .A2(n9467), .ZN(n9628) );
  OR2_X1 U9524 ( .A1(n9629), .A2(n9630), .ZN(n9467) );
  AND2_X1 U9525 ( .A1(n9464), .A2(n9463), .ZN(n9630) );
  AND2_X1 U9526 ( .A1(n9461), .A2(n9631), .ZN(n9629) );
  OR2_X1 U9527 ( .A1(n9464), .A2(n9463), .ZN(n9631) );
  OR2_X1 U9528 ( .A1(n9632), .A2(n9633), .ZN(n9463) );
  AND2_X1 U9529 ( .A1(n9460), .A2(n9459), .ZN(n9633) );
  AND2_X1 U9530 ( .A1(n9457), .A2(n9634), .ZN(n9632) );
  OR2_X1 U9531 ( .A1(n9460), .A2(n9459), .ZN(n9634) );
  OR2_X1 U9532 ( .A1(n9635), .A2(n9636), .ZN(n9459) );
  AND2_X1 U9533 ( .A1(n9456), .A2(n9455), .ZN(n9636) );
  AND2_X1 U9534 ( .A1(n9453), .A2(n9637), .ZN(n9635) );
  OR2_X1 U9535 ( .A1(n9456), .A2(n9455), .ZN(n9637) );
  OR2_X1 U9536 ( .A1(n9638), .A2(n9639), .ZN(n9455) );
  AND2_X1 U9537 ( .A1(n9452), .A2(n9451), .ZN(n9639) );
  AND2_X1 U9538 ( .A1(n9449), .A2(n9640), .ZN(n9638) );
  OR2_X1 U9539 ( .A1(n9452), .A2(n9451), .ZN(n9640) );
  OR2_X1 U9540 ( .A1(n9641), .A2(n9642), .ZN(n9451) );
  AND2_X1 U9541 ( .A1(n9448), .A2(n9447), .ZN(n9642) );
  AND2_X1 U9542 ( .A1(n9445), .A2(n9643), .ZN(n9641) );
  OR2_X1 U9543 ( .A1(n9448), .A2(n9447), .ZN(n9643) );
  OR2_X1 U9544 ( .A1(n9644), .A2(n9645), .ZN(n9447) );
  AND2_X1 U9545 ( .A1(n9441), .A2(n9444), .ZN(n9645) );
  AND2_X1 U9546 ( .A1(n9443), .A2(n9646), .ZN(n9644) );
  OR2_X1 U9547 ( .A1(n9441), .A2(n9444), .ZN(n9646) );
  OR3_X1 U9548 ( .A1(n9318), .A2(n9200), .A3(n8519), .ZN(n9444) );
  OR2_X1 U9549 ( .A1(n9200), .A2(n7606), .ZN(n9441) );
  INV_X1 U9550 ( .A(n9647), .ZN(n9443) );
  OR2_X1 U9551 ( .A1(n9648), .A2(n9649), .ZN(n9647) );
  AND2_X1 U9552 ( .A1(n9650), .A2(n9651), .ZN(n9649) );
  OR2_X1 U9553 ( .A1(n9652), .A2(n7697), .ZN(n9651) );
  AND2_X1 U9554 ( .A1(n9318), .A2(n7691), .ZN(n9652) );
  AND2_X1 U9555 ( .A1(n9436), .A2(n9653), .ZN(n9648) );
  OR2_X1 U9556 ( .A1(n9654), .A2(n7701), .ZN(n9653) );
  AND2_X1 U9557 ( .A1(n8358), .A2(n7703), .ZN(n9654) );
  OR2_X1 U9558 ( .A1(n7662), .A2(n9200), .ZN(n9448) );
  XNOR2_X1 U9559 ( .A(n9655), .B(n9656), .ZN(n9445) );
  XNOR2_X1 U9560 ( .A(n9657), .B(n9658), .ZN(n9656) );
  OR2_X1 U9561 ( .A1(n7660), .A2(n9200), .ZN(n9452) );
  XOR2_X1 U9562 ( .A(n9659), .B(n9660), .Z(n9449) );
  XOR2_X1 U9563 ( .A(n9661), .B(n9662), .Z(n9660) );
  OR2_X1 U9564 ( .A1(n7658), .A2(n9200), .ZN(n9456) );
  XOR2_X1 U9565 ( .A(n9663), .B(n9664), .Z(n9453) );
  XOR2_X1 U9566 ( .A(n9665), .B(n9666), .Z(n9664) );
  OR2_X1 U9567 ( .A1(n7656), .A2(n9200), .ZN(n9460) );
  XOR2_X1 U9568 ( .A(n9667), .B(n9668), .Z(n9457) );
  XOR2_X1 U9569 ( .A(n9669), .B(n9670), .Z(n9668) );
  OR2_X1 U9570 ( .A1(n7654), .A2(n9200), .ZN(n9464) );
  XOR2_X1 U9571 ( .A(n9671), .B(n9672), .Z(n9461) );
  XOR2_X1 U9572 ( .A(n9673), .B(n9674), .Z(n9672) );
  OR2_X1 U9573 ( .A1(n7652), .A2(n9200), .ZN(n9468) );
  XOR2_X1 U9574 ( .A(n9675), .B(n9676), .Z(n9465) );
  XOR2_X1 U9575 ( .A(n9677), .B(n9678), .Z(n9676) );
  OR2_X1 U9576 ( .A1(n7650), .A2(n9200), .ZN(n9472) );
  XOR2_X1 U9577 ( .A(n9679), .B(n9680), .Z(n9469) );
  XOR2_X1 U9578 ( .A(n9681), .B(n9682), .Z(n9680) );
  OR2_X1 U9579 ( .A1(n7648), .A2(n9200), .ZN(n9476) );
  XOR2_X1 U9580 ( .A(n9683), .B(n9684), .Z(n9473) );
  XOR2_X1 U9581 ( .A(n9685), .B(n9686), .Z(n9684) );
  OR2_X1 U9582 ( .A1(n7646), .A2(n9200), .ZN(n9480) );
  XOR2_X1 U9583 ( .A(n9687), .B(n9688), .Z(n9477) );
  XOR2_X1 U9584 ( .A(n9689), .B(n9690), .Z(n9688) );
  OR2_X1 U9585 ( .A1(n7644), .A2(n9200), .ZN(n9484) );
  XOR2_X1 U9586 ( .A(n9691), .B(n9692), .Z(n9481) );
  XOR2_X1 U9587 ( .A(n9693), .B(n9694), .Z(n9692) );
  OR2_X1 U9588 ( .A1(n7642), .A2(n9200), .ZN(n9488) );
  XOR2_X1 U9589 ( .A(n9695), .B(n9696), .Z(n9485) );
  XOR2_X1 U9590 ( .A(n9697), .B(n9698), .Z(n9696) );
  OR2_X1 U9591 ( .A1(n7640), .A2(n9200), .ZN(n9492) );
  XOR2_X1 U9592 ( .A(n9699), .B(n9700), .Z(n9489) );
  XOR2_X1 U9593 ( .A(n9701), .B(n9702), .Z(n9700) );
  OR2_X1 U9594 ( .A1(n7638), .A2(n9200), .ZN(n9496) );
  XOR2_X1 U9595 ( .A(n9703), .B(n9704), .Z(n9493) );
  XOR2_X1 U9596 ( .A(n9705), .B(n9706), .Z(n9704) );
  OR2_X1 U9597 ( .A1(n7636), .A2(n9200), .ZN(n9500) );
  XOR2_X1 U9598 ( .A(n9707), .B(n9708), .Z(n9497) );
  XOR2_X1 U9599 ( .A(n9709), .B(n9710), .Z(n9708) );
  OR2_X1 U9600 ( .A1(n7634), .A2(n9200), .ZN(n9504) );
  XOR2_X1 U9601 ( .A(n9711), .B(n9712), .Z(n9501) );
  XOR2_X1 U9602 ( .A(n9713), .B(n9714), .Z(n9712) );
  OR2_X1 U9603 ( .A1(n7632), .A2(n9200), .ZN(n9508) );
  XOR2_X1 U9604 ( .A(n9715), .B(n9716), .Z(n9505) );
  XOR2_X1 U9605 ( .A(n9717), .B(n9718), .Z(n9716) );
  OR2_X1 U9606 ( .A1(n7630), .A2(n9200), .ZN(n9512) );
  XOR2_X1 U9607 ( .A(n9719), .B(n9720), .Z(n9509) );
  XOR2_X1 U9608 ( .A(n9721), .B(n9722), .Z(n9720) );
  OR2_X1 U9609 ( .A1(n7628), .A2(n9200), .ZN(n9516) );
  XOR2_X1 U9610 ( .A(n9723), .B(n9724), .Z(n9513) );
  XOR2_X1 U9611 ( .A(n9725), .B(n9726), .Z(n9724) );
  OR2_X1 U9612 ( .A1(n7626), .A2(n9200), .ZN(n9520) );
  XOR2_X1 U9613 ( .A(n9727), .B(n9728), .Z(n9517) );
  XOR2_X1 U9614 ( .A(n9729), .B(n9730), .Z(n9728) );
  OR2_X1 U9615 ( .A1(n7624), .A2(n9200), .ZN(n9524) );
  XOR2_X1 U9616 ( .A(n9731), .B(n9732), .Z(n9521) );
  XOR2_X1 U9617 ( .A(n9733), .B(n9734), .Z(n9732) );
  OR2_X1 U9618 ( .A1(n7622), .A2(n9200), .ZN(n9528) );
  XOR2_X1 U9619 ( .A(n9735), .B(n9736), .Z(n9525) );
  XOR2_X1 U9620 ( .A(n9737), .B(n9738), .Z(n9736) );
  OR2_X1 U9621 ( .A1(n7620), .A2(n9200), .ZN(n9532) );
  XOR2_X1 U9622 ( .A(n9739), .B(n9740), .Z(n9529) );
  XOR2_X1 U9623 ( .A(n9741), .B(n9742), .Z(n9740) );
  XOR2_X1 U9624 ( .A(n9743), .B(n9744), .Z(n9533) );
  XOR2_X1 U9625 ( .A(n9745), .B(n9746), .Z(n9744) );
  OR2_X1 U9626 ( .A1(n7616), .A2(n9200), .ZN(n9540) );
  XOR2_X1 U9627 ( .A(n9747), .B(n9748), .Z(n9537) );
  XOR2_X1 U9628 ( .A(n9749), .B(n9750), .Z(n9748) );
  OR2_X1 U9629 ( .A1(n7614), .A2(n9200), .ZN(n9544) );
  XOR2_X1 U9630 ( .A(n9751), .B(n9752), .Z(n9541) );
  XOR2_X1 U9631 ( .A(n9753), .B(n9754), .Z(n9752) );
  OR2_X1 U9632 ( .A1(n7612), .A2(n9200), .ZN(n9548) );
  XOR2_X1 U9633 ( .A(n9755), .B(n9756), .Z(n9545) );
  XOR2_X1 U9634 ( .A(n9757), .B(n9758), .Z(n9756) );
  OR2_X1 U9635 ( .A1(n8056), .A2(n9200), .ZN(n9552) );
  XOR2_X1 U9636 ( .A(n9759), .B(n9760), .Z(n9549) );
  XOR2_X1 U9637 ( .A(n9761), .B(n9762), .Z(n9760) );
  OR2_X1 U9638 ( .A1(n8023), .A2(n9200), .ZN(n9558) );
  INV_X1 U9639 ( .A(n9195), .ZN(n9200) );
  XOR2_X1 U9640 ( .A(n9763), .B(n9764), .Z(n9195) );
  XNOR2_X1 U9641 ( .A(c_26_), .B(d_26_), .ZN(n9763) );
  XOR2_X1 U9642 ( .A(n9765), .B(n9766), .Z(n9555) );
  XOR2_X1 U9643 ( .A(n9767), .B(n9768), .Z(n9766) );
  XOR2_X1 U9644 ( .A(n9323), .B(n9769), .Z(n9315) );
  XOR2_X1 U9645 ( .A(n9322), .B(n9321), .Z(n9769) );
  OR2_X1 U9646 ( .A1(n8023), .A2(n9318), .ZN(n9321) );
  OR2_X1 U9647 ( .A1(n9770), .A2(n9771), .ZN(n9322) );
  AND2_X1 U9648 ( .A1(n9768), .A2(n9767), .ZN(n9771) );
  AND2_X1 U9649 ( .A1(n9765), .A2(n9772), .ZN(n9770) );
  OR2_X1 U9650 ( .A1(n9768), .A2(n9767), .ZN(n9772) );
  OR2_X1 U9651 ( .A1(n9773), .A2(n9774), .ZN(n9767) );
  AND2_X1 U9652 ( .A1(n9762), .A2(n9761), .ZN(n9774) );
  AND2_X1 U9653 ( .A1(n9759), .A2(n9775), .ZN(n9773) );
  OR2_X1 U9654 ( .A1(n9762), .A2(n9761), .ZN(n9775) );
  OR2_X1 U9655 ( .A1(n9776), .A2(n9777), .ZN(n9761) );
  AND2_X1 U9656 ( .A1(n9758), .A2(n9757), .ZN(n9777) );
  AND2_X1 U9657 ( .A1(n9755), .A2(n9778), .ZN(n9776) );
  OR2_X1 U9658 ( .A1(n9758), .A2(n9757), .ZN(n9778) );
  OR2_X1 U9659 ( .A1(n9779), .A2(n9780), .ZN(n9757) );
  AND2_X1 U9660 ( .A1(n9754), .A2(n9753), .ZN(n9780) );
  AND2_X1 U9661 ( .A1(n9751), .A2(n9781), .ZN(n9779) );
  OR2_X1 U9662 ( .A1(n9754), .A2(n9753), .ZN(n9781) );
  OR2_X1 U9663 ( .A1(n9782), .A2(n9783), .ZN(n9753) );
  AND2_X1 U9664 ( .A1(n9750), .A2(n9749), .ZN(n9783) );
  AND2_X1 U9665 ( .A1(n9747), .A2(n9784), .ZN(n9782) );
  OR2_X1 U9666 ( .A1(n9750), .A2(n9749), .ZN(n9784) );
  OR2_X1 U9667 ( .A1(n7618), .A2(n9318), .ZN(n9749) );
  OR2_X1 U9668 ( .A1(n9785), .A2(n9786), .ZN(n9750) );
  AND2_X1 U9669 ( .A1(n9746), .A2(n9745), .ZN(n9786) );
  AND2_X1 U9670 ( .A1(n9743), .A2(n9787), .ZN(n9785) );
  OR2_X1 U9671 ( .A1(n9746), .A2(n9745), .ZN(n9787) );
  OR2_X1 U9672 ( .A1(n9788), .A2(n9789), .ZN(n9745) );
  AND2_X1 U9673 ( .A1(n9742), .A2(n9741), .ZN(n9789) );
  AND2_X1 U9674 ( .A1(n9739), .A2(n9790), .ZN(n9788) );
  OR2_X1 U9675 ( .A1(n9742), .A2(n9741), .ZN(n9790) );
  OR2_X1 U9676 ( .A1(n9791), .A2(n9792), .ZN(n9741) );
  AND2_X1 U9677 ( .A1(n9738), .A2(n9737), .ZN(n9792) );
  AND2_X1 U9678 ( .A1(n9735), .A2(n9793), .ZN(n9791) );
  OR2_X1 U9679 ( .A1(n9738), .A2(n9737), .ZN(n9793) );
  OR2_X1 U9680 ( .A1(n9794), .A2(n9795), .ZN(n9737) );
  AND2_X1 U9681 ( .A1(n9734), .A2(n9733), .ZN(n9795) );
  AND2_X1 U9682 ( .A1(n9731), .A2(n9796), .ZN(n9794) );
  OR2_X1 U9683 ( .A1(n9734), .A2(n9733), .ZN(n9796) );
  OR2_X1 U9684 ( .A1(n7626), .A2(n9318), .ZN(n9733) );
  OR2_X1 U9685 ( .A1(n9797), .A2(n9798), .ZN(n9734) );
  AND2_X1 U9686 ( .A1(n9730), .A2(n9729), .ZN(n9798) );
  AND2_X1 U9687 ( .A1(n9727), .A2(n9799), .ZN(n9797) );
  OR2_X1 U9688 ( .A1(n9730), .A2(n9729), .ZN(n9799) );
  OR2_X1 U9689 ( .A1(n9800), .A2(n9801), .ZN(n9729) );
  AND2_X1 U9690 ( .A1(n9726), .A2(n9725), .ZN(n9801) );
  AND2_X1 U9691 ( .A1(n9723), .A2(n9802), .ZN(n9800) );
  OR2_X1 U9692 ( .A1(n9726), .A2(n9725), .ZN(n9802) );
  OR2_X1 U9693 ( .A1(n9803), .A2(n9804), .ZN(n9725) );
  AND2_X1 U9694 ( .A1(n9722), .A2(n9721), .ZN(n9804) );
  AND2_X1 U9695 ( .A1(n9719), .A2(n9805), .ZN(n9803) );
  OR2_X1 U9696 ( .A1(n9722), .A2(n9721), .ZN(n9805) );
  OR2_X1 U9697 ( .A1(n9806), .A2(n9807), .ZN(n9721) );
  AND2_X1 U9698 ( .A1(n9718), .A2(n9717), .ZN(n9807) );
  AND2_X1 U9699 ( .A1(n9715), .A2(n9808), .ZN(n9806) );
  OR2_X1 U9700 ( .A1(n9718), .A2(n9717), .ZN(n9808) );
  OR2_X1 U9701 ( .A1(n9809), .A2(n9810), .ZN(n9717) );
  AND2_X1 U9702 ( .A1(n9714), .A2(n9713), .ZN(n9810) );
  AND2_X1 U9703 ( .A1(n9711), .A2(n9811), .ZN(n9809) );
  OR2_X1 U9704 ( .A1(n9714), .A2(n9713), .ZN(n9811) );
  OR2_X1 U9705 ( .A1(n9812), .A2(n9813), .ZN(n9713) );
  AND2_X1 U9706 ( .A1(n9710), .A2(n9709), .ZN(n9813) );
  AND2_X1 U9707 ( .A1(n9707), .A2(n9814), .ZN(n9812) );
  OR2_X1 U9708 ( .A1(n9710), .A2(n9709), .ZN(n9814) );
  OR2_X1 U9709 ( .A1(n9815), .A2(n9816), .ZN(n9709) );
  AND2_X1 U9710 ( .A1(n9706), .A2(n9705), .ZN(n9816) );
  AND2_X1 U9711 ( .A1(n9703), .A2(n9817), .ZN(n9815) );
  OR2_X1 U9712 ( .A1(n9706), .A2(n9705), .ZN(n9817) );
  OR2_X1 U9713 ( .A1(n9818), .A2(n9819), .ZN(n9705) );
  AND2_X1 U9714 ( .A1(n9702), .A2(n9701), .ZN(n9819) );
  AND2_X1 U9715 ( .A1(n9699), .A2(n9820), .ZN(n9818) );
  OR2_X1 U9716 ( .A1(n9702), .A2(n9701), .ZN(n9820) );
  OR2_X1 U9717 ( .A1(n9821), .A2(n9822), .ZN(n9701) );
  AND2_X1 U9718 ( .A1(n9698), .A2(n9697), .ZN(n9822) );
  AND2_X1 U9719 ( .A1(n9695), .A2(n9823), .ZN(n9821) );
  OR2_X1 U9720 ( .A1(n9698), .A2(n9697), .ZN(n9823) );
  OR2_X1 U9721 ( .A1(n9824), .A2(n9825), .ZN(n9697) );
  AND2_X1 U9722 ( .A1(n9694), .A2(n9693), .ZN(n9825) );
  AND2_X1 U9723 ( .A1(n9691), .A2(n9826), .ZN(n9824) );
  OR2_X1 U9724 ( .A1(n9694), .A2(n9693), .ZN(n9826) );
  OR2_X1 U9725 ( .A1(n9827), .A2(n9828), .ZN(n9693) );
  AND2_X1 U9726 ( .A1(n9690), .A2(n9689), .ZN(n9828) );
  AND2_X1 U9727 ( .A1(n9687), .A2(n9829), .ZN(n9827) );
  OR2_X1 U9728 ( .A1(n9690), .A2(n9689), .ZN(n9829) );
  OR2_X1 U9729 ( .A1(n9830), .A2(n9831), .ZN(n9689) );
  AND2_X1 U9730 ( .A1(n9686), .A2(n9685), .ZN(n9831) );
  AND2_X1 U9731 ( .A1(n9683), .A2(n9832), .ZN(n9830) );
  OR2_X1 U9732 ( .A1(n9686), .A2(n9685), .ZN(n9832) );
  OR2_X1 U9733 ( .A1(n9833), .A2(n9834), .ZN(n9685) );
  AND2_X1 U9734 ( .A1(n9682), .A2(n9681), .ZN(n9834) );
  AND2_X1 U9735 ( .A1(n9679), .A2(n9835), .ZN(n9833) );
  OR2_X1 U9736 ( .A1(n9682), .A2(n9681), .ZN(n9835) );
  OR2_X1 U9737 ( .A1(n9836), .A2(n9837), .ZN(n9681) );
  AND2_X1 U9738 ( .A1(n9678), .A2(n9677), .ZN(n9837) );
  AND2_X1 U9739 ( .A1(n9675), .A2(n9838), .ZN(n9836) );
  OR2_X1 U9740 ( .A1(n9678), .A2(n9677), .ZN(n9838) );
  OR2_X1 U9741 ( .A1(n9839), .A2(n9840), .ZN(n9677) );
  AND2_X1 U9742 ( .A1(n9674), .A2(n9673), .ZN(n9840) );
  AND2_X1 U9743 ( .A1(n9671), .A2(n9841), .ZN(n9839) );
  OR2_X1 U9744 ( .A1(n9674), .A2(n9673), .ZN(n9841) );
  OR2_X1 U9745 ( .A1(n9842), .A2(n9843), .ZN(n9673) );
  AND2_X1 U9746 ( .A1(n9670), .A2(n9669), .ZN(n9843) );
  AND2_X1 U9747 ( .A1(n9667), .A2(n9844), .ZN(n9842) );
  OR2_X1 U9748 ( .A1(n9670), .A2(n9669), .ZN(n9844) );
  OR2_X1 U9749 ( .A1(n9845), .A2(n9846), .ZN(n9669) );
  AND2_X1 U9750 ( .A1(n9666), .A2(n9665), .ZN(n9846) );
  AND2_X1 U9751 ( .A1(n9663), .A2(n9847), .ZN(n9845) );
  OR2_X1 U9752 ( .A1(n9666), .A2(n9665), .ZN(n9847) );
  OR2_X1 U9753 ( .A1(n9848), .A2(n9849), .ZN(n9665) );
  AND2_X1 U9754 ( .A1(n9662), .A2(n9661), .ZN(n9849) );
  AND2_X1 U9755 ( .A1(n9659), .A2(n9850), .ZN(n9848) );
  OR2_X1 U9756 ( .A1(n9662), .A2(n9661), .ZN(n9850) );
  OR2_X1 U9757 ( .A1(n9851), .A2(n9852), .ZN(n9661) );
  AND2_X1 U9758 ( .A1(n9655), .A2(n9658), .ZN(n9852) );
  AND2_X1 U9759 ( .A1(n9657), .A2(n9853), .ZN(n9851) );
  OR2_X1 U9760 ( .A1(n9655), .A2(n9658), .ZN(n9853) );
  OR3_X1 U9761 ( .A1(n8358), .A2(n9318), .A3(n8519), .ZN(n9658) );
  OR2_X1 U9762 ( .A1(n9318), .A2(n7606), .ZN(n9655) );
  INV_X1 U9763 ( .A(n9854), .ZN(n9657) );
  OR2_X1 U9764 ( .A1(n9855), .A2(n9856), .ZN(n9854) );
  AND2_X1 U9765 ( .A1(n9857), .A2(n9858), .ZN(n9856) );
  OR2_X1 U9766 ( .A1(n9859), .A2(n7697), .ZN(n9858) );
  AND2_X1 U9767 ( .A1(n8358), .A2(n7691), .ZN(n9859) );
  AND2_X1 U9768 ( .A1(n9650), .A2(n9860), .ZN(n9855) );
  OR2_X1 U9769 ( .A1(n9861), .A2(n7701), .ZN(n9860) );
  AND2_X1 U9770 ( .A1(n8335), .A2(n7703), .ZN(n9861) );
  OR2_X1 U9771 ( .A1(n7662), .A2(n9318), .ZN(n9662) );
  XNOR2_X1 U9772 ( .A(n9862), .B(n9863), .ZN(n9659) );
  XNOR2_X1 U9773 ( .A(n9864), .B(n9865), .ZN(n9863) );
  OR2_X1 U9774 ( .A1(n7660), .A2(n9318), .ZN(n9666) );
  XOR2_X1 U9775 ( .A(n9866), .B(n9867), .Z(n9663) );
  XOR2_X1 U9776 ( .A(n9868), .B(n9869), .Z(n9867) );
  OR2_X1 U9777 ( .A1(n7658), .A2(n9318), .ZN(n9670) );
  XOR2_X1 U9778 ( .A(n9870), .B(n9871), .Z(n9667) );
  XOR2_X1 U9779 ( .A(n9872), .B(n9873), .Z(n9871) );
  OR2_X1 U9780 ( .A1(n7656), .A2(n9318), .ZN(n9674) );
  XOR2_X1 U9781 ( .A(n9874), .B(n9875), .Z(n9671) );
  XOR2_X1 U9782 ( .A(n9876), .B(n9877), .Z(n9875) );
  OR2_X1 U9783 ( .A1(n7654), .A2(n9318), .ZN(n9678) );
  XOR2_X1 U9784 ( .A(n9878), .B(n9879), .Z(n9675) );
  XOR2_X1 U9785 ( .A(n9880), .B(n9881), .Z(n9879) );
  OR2_X1 U9786 ( .A1(n7652), .A2(n9318), .ZN(n9682) );
  XOR2_X1 U9787 ( .A(n9882), .B(n9883), .Z(n9679) );
  XOR2_X1 U9788 ( .A(n9884), .B(n9885), .Z(n9883) );
  OR2_X1 U9789 ( .A1(n7650), .A2(n9318), .ZN(n9686) );
  XOR2_X1 U9790 ( .A(n9886), .B(n9887), .Z(n9683) );
  XOR2_X1 U9791 ( .A(n9888), .B(n9889), .Z(n9887) );
  OR2_X1 U9792 ( .A1(n7648), .A2(n9318), .ZN(n9690) );
  XOR2_X1 U9793 ( .A(n9890), .B(n9891), .Z(n9687) );
  XOR2_X1 U9794 ( .A(n9892), .B(n9893), .Z(n9891) );
  OR2_X1 U9795 ( .A1(n7646), .A2(n9318), .ZN(n9694) );
  XOR2_X1 U9796 ( .A(n9894), .B(n9895), .Z(n9691) );
  XOR2_X1 U9797 ( .A(n9896), .B(n9897), .Z(n9895) );
  OR2_X1 U9798 ( .A1(n7644), .A2(n9318), .ZN(n9698) );
  XOR2_X1 U9799 ( .A(n9898), .B(n9899), .Z(n9695) );
  XOR2_X1 U9800 ( .A(n9900), .B(n9901), .Z(n9899) );
  OR2_X1 U9801 ( .A1(n7642), .A2(n9318), .ZN(n9702) );
  XOR2_X1 U9802 ( .A(n9902), .B(n9903), .Z(n9699) );
  XOR2_X1 U9803 ( .A(n9904), .B(n9905), .Z(n9903) );
  OR2_X1 U9804 ( .A1(n7640), .A2(n9318), .ZN(n9706) );
  XOR2_X1 U9805 ( .A(n9906), .B(n9907), .Z(n9703) );
  XOR2_X1 U9806 ( .A(n9908), .B(n9909), .Z(n9907) );
  OR2_X1 U9807 ( .A1(n7638), .A2(n9318), .ZN(n9710) );
  XOR2_X1 U9808 ( .A(n9910), .B(n9911), .Z(n9707) );
  XOR2_X1 U9809 ( .A(n9912), .B(n9913), .Z(n9911) );
  OR2_X1 U9810 ( .A1(n7636), .A2(n9318), .ZN(n9714) );
  XOR2_X1 U9811 ( .A(n9914), .B(n9915), .Z(n9711) );
  XOR2_X1 U9812 ( .A(n9916), .B(n9917), .Z(n9915) );
  OR2_X1 U9813 ( .A1(n7634), .A2(n9318), .ZN(n9718) );
  XOR2_X1 U9814 ( .A(n9918), .B(n9919), .Z(n9715) );
  XOR2_X1 U9815 ( .A(n9920), .B(n9921), .Z(n9919) );
  OR2_X1 U9816 ( .A1(n7632), .A2(n9318), .ZN(n9722) );
  XOR2_X1 U9817 ( .A(n9922), .B(n9923), .Z(n9719) );
  XOR2_X1 U9818 ( .A(n9924), .B(n9925), .Z(n9923) );
  OR2_X1 U9819 ( .A1(n7630), .A2(n9318), .ZN(n9726) );
  XOR2_X1 U9820 ( .A(n9926), .B(n9927), .Z(n9723) );
  XOR2_X1 U9821 ( .A(n9928), .B(n9929), .Z(n9927) );
  OR2_X1 U9822 ( .A1(n7628), .A2(n9318), .ZN(n9730) );
  XOR2_X1 U9823 ( .A(n9930), .B(n9931), .Z(n9727) );
  XOR2_X1 U9824 ( .A(n9932), .B(n9933), .Z(n9931) );
  XOR2_X1 U9825 ( .A(n9934), .B(n9935), .Z(n9731) );
  XOR2_X1 U9826 ( .A(n9936), .B(n9937), .Z(n9935) );
  OR2_X1 U9827 ( .A1(n7624), .A2(n9318), .ZN(n9738) );
  XOR2_X1 U9828 ( .A(n9938), .B(n9939), .Z(n9735) );
  XOR2_X1 U9829 ( .A(n9940), .B(n9941), .Z(n9939) );
  OR2_X1 U9830 ( .A1(n7622), .A2(n9318), .ZN(n9742) );
  XOR2_X1 U9831 ( .A(n9942), .B(n9943), .Z(n9739) );
  XOR2_X1 U9832 ( .A(n9944), .B(n9945), .Z(n9943) );
  OR2_X1 U9833 ( .A1(n7620), .A2(n9318), .ZN(n9746) );
  XOR2_X1 U9834 ( .A(n9946), .B(n9947), .Z(n9743) );
  XOR2_X1 U9835 ( .A(n9948), .B(n9949), .Z(n9947) );
  XOR2_X1 U9836 ( .A(n9950), .B(n9951), .Z(n9747) );
  XOR2_X1 U9837 ( .A(n9952), .B(n9953), .Z(n9951) );
  OR2_X1 U9838 ( .A1(n7616), .A2(n9318), .ZN(n9754) );
  XOR2_X1 U9839 ( .A(n9954), .B(n9955), .Z(n9751) );
  XOR2_X1 U9840 ( .A(n9956), .B(n9957), .Z(n9955) );
  OR2_X1 U9841 ( .A1(n7614), .A2(n9318), .ZN(n9758) );
  XOR2_X1 U9842 ( .A(n9958), .B(n9959), .Z(n9755) );
  XOR2_X1 U9843 ( .A(n9960), .B(n9961), .Z(n9959) );
  OR2_X1 U9844 ( .A1(n8105), .A2(n9318), .ZN(n9762) );
  XOR2_X1 U9845 ( .A(n9962), .B(n9963), .Z(n9759) );
  XOR2_X1 U9846 ( .A(n9964), .B(n9965), .Z(n9963) );
  OR2_X1 U9847 ( .A1(n8056), .A2(n9318), .ZN(n9768) );
  INV_X1 U9848 ( .A(n9436), .ZN(n9318) );
  XOR2_X1 U9849 ( .A(n9966), .B(n9967), .Z(n9436) );
  XNOR2_X1 U9850 ( .A(c_25_), .B(d_25_), .ZN(n9966) );
  XOR2_X1 U9851 ( .A(n9968), .B(n9969), .Z(n9765) );
  XOR2_X1 U9852 ( .A(n9970), .B(n9971), .Z(n9969) );
  XOR2_X1 U9853 ( .A(n9341), .B(n9972), .Z(n9323) );
  XOR2_X1 U9854 ( .A(n9340), .B(n9339), .Z(n9972) );
  OR2_X1 U9855 ( .A1(n8056), .A2(n8358), .ZN(n9339) );
  OR2_X1 U9856 ( .A1(n9973), .A2(n9974), .ZN(n9340) );
  AND2_X1 U9857 ( .A1(n9971), .A2(n9970), .ZN(n9974) );
  AND2_X1 U9858 ( .A1(n9968), .A2(n9975), .ZN(n9973) );
  OR2_X1 U9859 ( .A1(n9971), .A2(n9970), .ZN(n9975) );
  OR2_X1 U9860 ( .A1(n8105), .A2(n8358), .ZN(n9970) );
  OR2_X1 U9861 ( .A1(n9976), .A2(n9977), .ZN(n9971) );
  AND2_X1 U9862 ( .A1(n9965), .A2(n9964), .ZN(n9977) );
  AND2_X1 U9863 ( .A1(n9962), .A2(n9978), .ZN(n9976) );
  OR2_X1 U9864 ( .A1(n9965), .A2(n9964), .ZN(n9978) );
  OR2_X1 U9865 ( .A1(n9979), .A2(n9980), .ZN(n9964) );
  AND2_X1 U9866 ( .A1(n9961), .A2(n9960), .ZN(n9980) );
  AND2_X1 U9867 ( .A1(n9958), .A2(n9981), .ZN(n9979) );
  OR2_X1 U9868 ( .A1(n9961), .A2(n9960), .ZN(n9981) );
  OR2_X1 U9869 ( .A1(n9982), .A2(n9983), .ZN(n9960) );
  AND2_X1 U9870 ( .A1(n9957), .A2(n9956), .ZN(n9983) );
  AND2_X1 U9871 ( .A1(n9954), .A2(n9984), .ZN(n9982) );
  OR2_X1 U9872 ( .A1(n9957), .A2(n9956), .ZN(n9984) );
  OR2_X1 U9873 ( .A1(n7618), .A2(n8358), .ZN(n9956) );
  OR2_X1 U9874 ( .A1(n9985), .A2(n9986), .ZN(n9957) );
  AND2_X1 U9875 ( .A1(n9953), .A2(n9952), .ZN(n9986) );
  AND2_X1 U9876 ( .A1(n9950), .A2(n9987), .ZN(n9985) );
  OR2_X1 U9877 ( .A1(n9953), .A2(n9952), .ZN(n9987) );
  OR2_X1 U9878 ( .A1(n9988), .A2(n9989), .ZN(n9952) );
  AND2_X1 U9879 ( .A1(n9949), .A2(n9948), .ZN(n9989) );
  AND2_X1 U9880 ( .A1(n9946), .A2(n9990), .ZN(n9988) );
  OR2_X1 U9881 ( .A1(n9949), .A2(n9948), .ZN(n9990) );
  OR2_X1 U9882 ( .A1(n9991), .A2(n9992), .ZN(n9948) );
  AND2_X1 U9883 ( .A1(n9945), .A2(n9944), .ZN(n9992) );
  AND2_X1 U9884 ( .A1(n9942), .A2(n9993), .ZN(n9991) );
  OR2_X1 U9885 ( .A1(n9945), .A2(n9944), .ZN(n9993) );
  OR2_X1 U9886 ( .A1(n9994), .A2(n9995), .ZN(n9944) );
  AND2_X1 U9887 ( .A1(n9941), .A2(n9940), .ZN(n9995) );
  AND2_X1 U9888 ( .A1(n9938), .A2(n9996), .ZN(n9994) );
  OR2_X1 U9889 ( .A1(n9941), .A2(n9940), .ZN(n9996) );
  OR2_X1 U9890 ( .A1(n7626), .A2(n8358), .ZN(n9940) );
  OR2_X1 U9891 ( .A1(n9997), .A2(n9998), .ZN(n9941) );
  AND2_X1 U9892 ( .A1(n9937), .A2(n9936), .ZN(n9998) );
  AND2_X1 U9893 ( .A1(n9934), .A2(n9999), .ZN(n9997) );
  OR2_X1 U9894 ( .A1(n9937), .A2(n9936), .ZN(n9999) );
  OR2_X1 U9895 ( .A1(n10000), .A2(n10001), .ZN(n9936) );
  AND2_X1 U9896 ( .A1(n9933), .A2(n9932), .ZN(n10001) );
  AND2_X1 U9897 ( .A1(n9930), .A2(n10002), .ZN(n10000) );
  OR2_X1 U9898 ( .A1(n9933), .A2(n9932), .ZN(n10002) );
  OR2_X1 U9899 ( .A1(n10003), .A2(n10004), .ZN(n9932) );
  AND2_X1 U9900 ( .A1(n9929), .A2(n9928), .ZN(n10004) );
  AND2_X1 U9901 ( .A1(n9926), .A2(n10005), .ZN(n10003) );
  OR2_X1 U9902 ( .A1(n9929), .A2(n9928), .ZN(n10005) );
  OR2_X1 U9903 ( .A1(n10006), .A2(n10007), .ZN(n9928) );
  AND2_X1 U9904 ( .A1(n9925), .A2(n9924), .ZN(n10007) );
  AND2_X1 U9905 ( .A1(n9922), .A2(n10008), .ZN(n10006) );
  OR2_X1 U9906 ( .A1(n9925), .A2(n9924), .ZN(n10008) );
  OR2_X1 U9907 ( .A1(n10009), .A2(n10010), .ZN(n9924) );
  AND2_X1 U9908 ( .A1(n9921), .A2(n9920), .ZN(n10010) );
  AND2_X1 U9909 ( .A1(n9918), .A2(n10011), .ZN(n10009) );
  OR2_X1 U9910 ( .A1(n9921), .A2(n9920), .ZN(n10011) );
  OR2_X1 U9911 ( .A1(n10012), .A2(n10013), .ZN(n9920) );
  AND2_X1 U9912 ( .A1(n9917), .A2(n9916), .ZN(n10013) );
  AND2_X1 U9913 ( .A1(n9914), .A2(n10014), .ZN(n10012) );
  OR2_X1 U9914 ( .A1(n9917), .A2(n9916), .ZN(n10014) );
  OR2_X1 U9915 ( .A1(n10015), .A2(n10016), .ZN(n9916) );
  AND2_X1 U9916 ( .A1(n9913), .A2(n9912), .ZN(n10016) );
  AND2_X1 U9917 ( .A1(n9910), .A2(n10017), .ZN(n10015) );
  OR2_X1 U9918 ( .A1(n9913), .A2(n9912), .ZN(n10017) );
  OR2_X1 U9919 ( .A1(n10018), .A2(n10019), .ZN(n9912) );
  AND2_X1 U9920 ( .A1(n9909), .A2(n9908), .ZN(n10019) );
  AND2_X1 U9921 ( .A1(n9906), .A2(n10020), .ZN(n10018) );
  OR2_X1 U9922 ( .A1(n9909), .A2(n9908), .ZN(n10020) );
  OR2_X1 U9923 ( .A1(n10021), .A2(n10022), .ZN(n9908) );
  AND2_X1 U9924 ( .A1(n9905), .A2(n9904), .ZN(n10022) );
  AND2_X1 U9925 ( .A1(n9902), .A2(n10023), .ZN(n10021) );
  OR2_X1 U9926 ( .A1(n9905), .A2(n9904), .ZN(n10023) );
  OR2_X1 U9927 ( .A1(n10024), .A2(n10025), .ZN(n9904) );
  AND2_X1 U9928 ( .A1(n9901), .A2(n9900), .ZN(n10025) );
  AND2_X1 U9929 ( .A1(n9898), .A2(n10026), .ZN(n10024) );
  OR2_X1 U9930 ( .A1(n9901), .A2(n9900), .ZN(n10026) );
  OR2_X1 U9931 ( .A1(n10027), .A2(n10028), .ZN(n9900) );
  AND2_X1 U9932 ( .A1(n9897), .A2(n9896), .ZN(n10028) );
  AND2_X1 U9933 ( .A1(n9894), .A2(n10029), .ZN(n10027) );
  OR2_X1 U9934 ( .A1(n9897), .A2(n9896), .ZN(n10029) );
  OR2_X1 U9935 ( .A1(n10030), .A2(n10031), .ZN(n9896) );
  AND2_X1 U9936 ( .A1(n9893), .A2(n9892), .ZN(n10031) );
  AND2_X1 U9937 ( .A1(n9890), .A2(n10032), .ZN(n10030) );
  OR2_X1 U9938 ( .A1(n9893), .A2(n9892), .ZN(n10032) );
  OR2_X1 U9939 ( .A1(n10033), .A2(n10034), .ZN(n9892) );
  AND2_X1 U9940 ( .A1(n9889), .A2(n9888), .ZN(n10034) );
  AND2_X1 U9941 ( .A1(n9886), .A2(n10035), .ZN(n10033) );
  OR2_X1 U9942 ( .A1(n9889), .A2(n9888), .ZN(n10035) );
  OR2_X1 U9943 ( .A1(n10036), .A2(n10037), .ZN(n9888) );
  AND2_X1 U9944 ( .A1(n9885), .A2(n9884), .ZN(n10037) );
  AND2_X1 U9945 ( .A1(n9882), .A2(n10038), .ZN(n10036) );
  OR2_X1 U9946 ( .A1(n9885), .A2(n9884), .ZN(n10038) );
  OR2_X1 U9947 ( .A1(n10039), .A2(n10040), .ZN(n9884) );
  AND2_X1 U9948 ( .A1(n9881), .A2(n9880), .ZN(n10040) );
  AND2_X1 U9949 ( .A1(n9878), .A2(n10041), .ZN(n10039) );
  OR2_X1 U9950 ( .A1(n9881), .A2(n9880), .ZN(n10041) );
  OR2_X1 U9951 ( .A1(n10042), .A2(n10043), .ZN(n9880) );
  AND2_X1 U9952 ( .A1(n9877), .A2(n9876), .ZN(n10043) );
  AND2_X1 U9953 ( .A1(n9874), .A2(n10044), .ZN(n10042) );
  OR2_X1 U9954 ( .A1(n9877), .A2(n9876), .ZN(n10044) );
  OR2_X1 U9955 ( .A1(n10045), .A2(n10046), .ZN(n9876) );
  AND2_X1 U9956 ( .A1(n9873), .A2(n9872), .ZN(n10046) );
  AND2_X1 U9957 ( .A1(n9870), .A2(n10047), .ZN(n10045) );
  OR2_X1 U9958 ( .A1(n9873), .A2(n9872), .ZN(n10047) );
  OR2_X1 U9959 ( .A1(n10048), .A2(n10049), .ZN(n9872) );
  AND2_X1 U9960 ( .A1(n9869), .A2(n9868), .ZN(n10049) );
  AND2_X1 U9961 ( .A1(n9866), .A2(n10050), .ZN(n10048) );
  OR2_X1 U9962 ( .A1(n9869), .A2(n9868), .ZN(n10050) );
  OR2_X1 U9963 ( .A1(n10051), .A2(n10052), .ZN(n9868) );
  AND2_X1 U9964 ( .A1(n9862), .A2(n9865), .ZN(n10052) );
  AND2_X1 U9965 ( .A1(n9864), .A2(n10053), .ZN(n10051) );
  OR2_X1 U9966 ( .A1(n9862), .A2(n9865), .ZN(n10053) );
  OR3_X1 U9967 ( .A1(n8335), .A2(n8358), .A3(n8519), .ZN(n9865) );
  OR2_X1 U9968 ( .A1(n8358), .A2(n7606), .ZN(n9862) );
  INV_X1 U9969 ( .A(n10054), .ZN(n9864) );
  OR2_X1 U9970 ( .A1(n10055), .A2(n10056), .ZN(n10054) );
  AND2_X1 U9971 ( .A1(n10057), .A2(n10058), .ZN(n10056) );
  OR2_X1 U9972 ( .A1(n10059), .A2(n7697), .ZN(n10058) );
  AND2_X1 U9973 ( .A1(n8335), .A2(n7691), .ZN(n10059) );
  AND2_X1 U9974 ( .A1(n9857), .A2(n10060), .ZN(n10055) );
  OR2_X1 U9975 ( .A1(n10061), .A2(n7701), .ZN(n10060) );
  AND2_X1 U9976 ( .A1(n10062), .A2(n7703), .ZN(n10061) );
  OR2_X1 U9977 ( .A1(n7662), .A2(n8358), .ZN(n9869) );
  XNOR2_X1 U9978 ( .A(n10063), .B(n10064), .ZN(n9866) );
  XNOR2_X1 U9979 ( .A(n10065), .B(n10066), .ZN(n10064) );
  OR2_X1 U9980 ( .A1(n7660), .A2(n8358), .ZN(n9873) );
  XOR2_X1 U9981 ( .A(n10067), .B(n10068), .Z(n9870) );
  XOR2_X1 U9982 ( .A(n10069), .B(n10070), .Z(n10068) );
  OR2_X1 U9983 ( .A1(n7658), .A2(n8358), .ZN(n9877) );
  XOR2_X1 U9984 ( .A(n10071), .B(n10072), .Z(n9874) );
  XOR2_X1 U9985 ( .A(n10073), .B(n10074), .Z(n10072) );
  OR2_X1 U9986 ( .A1(n7656), .A2(n8358), .ZN(n9881) );
  XOR2_X1 U9987 ( .A(n10075), .B(n10076), .Z(n9878) );
  XOR2_X1 U9988 ( .A(n10077), .B(n10078), .Z(n10076) );
  OR2_X1 U9989 ( .A1(n7654), .A2(n8358), .ZN(n9885) );
  XOR2_X1 U9990 ( .A(n10079), .B(n10080), .Z(n9882) );
  XOR2_X1 U9991 ( .A(n10081), .B(n10082), .Z(n10080) );
  OR2_X1 U9992 ( .A1(n7652), .A2(n8358), .ZN(n9889) );
  XOR2_X1 U9993 ( .A(n10083), .B(n10084), .Z(n9886) );
  XOR2_X1 U9994 ( .A(n10085), .B(n10086), .Z(n10084) );
  OR2_X1 U9995 ( .A1(n7650), .A2(n8358), .ZN(n9893) );
  XOR2_X1 U9996 ( .A(n10087), .B(n10088), .Z(n9890) );
  XOR2_X1 U9997 ( .A(n10089), .B(n10090), .Z(n10088) );
  OR2_X1 U9998 ( .A1(n7648), .A2(n8358), .ZN(n9897) );
  XOR2_X1 U9999 ( .A(n10091), .B(n10092), .Z(n9894) );
  XOR2_X1 U10000 ( .A(n10093), .B(n10094), .Z(n10092) );
  OR2_X1 U10001 ( .A1(n7646), .A2(n8358), .ZN(n9901) );
  XOR2_X1 U10002 ( .A(n10095), .B(n10096), .Z(n9898) );
  XOR2_X1 U10003 ( .A(n10097), .B(n10098), .Z(n10096) );
  OR2_X1 U10004 ( .A1(n7644), .A2(n8358), .ZN(n9905) );
  XOR2_X1 U10005 ( .A(n10099), .B(n10100), .Z(n9902) );
  XOR2_X1 U10006 ( .A(n10101), .B(n10102), .Z(n10100) );
  OR2_X1 U10007 ( .A1(n7642), .A2(n8358), .ZN(n9909) );
  XOR2_X1 U10008 ( .A(n10103), .B(n10104), .Z(n9906) );
  XOR2_X1 U10009 ( .A(n10105), .B(n10106), .Z(n10104) );
  OR2_X1 U10010 ( .A1(n7640), .A2(n8358), .ZN(n9913) );
  XOR2_X1 U10011 ( .A(n10107), .B(n10108), .Z(n9910) );
  XOR2_X1 U10012 ( .A(n10109), .B(n10110), .Z(n10108) );
  OR2_X1 U10013 ( .A1(n7638), .A2(n8358), .ZN(n9917) );
  XOR2_X1 U10014 ( .A(n10111), .B(n10112), .Z(n9914) );
  XOR2_X1 U10015 ( .A(n10113), .B(n10114), .Z(n10112) );
  OR2_X1 U10016 ( .A1(n7636), .A2(n8358), .ZN(n9921) );
  XOR2_X1 U10017 ( .A(n10115), .B(n10116), .Z(n9918) );
  XOR2_X1 U10018 ( .A(n10117), .B(n10118), .Z(n10116) );
  OR2_X1 U10019 ( .A1(n7634), .A2(n8358), .ZN(n9925) );
  XOR2_X1 U10020 ( .A(n10119), .B(n10120), .Z(n9922) );
  XOR2_X1 U10021 ( .A(n10121), .B(n10122), .Z(n10120) );
  OR2_X1 U10022 ( .A1(n7632), .A2(n8358), .ZN(n9929) );
  XOR2_X1 U10023 ( .A(n10123), .B(n10124), .Z(n9926) );
  XOR2_X1 U10024 ( .A(n10125), .B(n10126), .Z(n10124) );
  OR2_X1 U10025 ( .A1(n7630), .A2(n8358), .ZN(n9933) );
  XOR2_X1 U10026 ( .A(n10127), .B(n10128), .Z(n9930) );
  XOR2_X1 U10027 ( .A(n10129), .B(n10130), .Z(n10128) );
  OR2_X1 U10028 ( .A1(n7628), .A2(n8358), .ZN(n9937) );
  XOR2_X1 U10029 ( .A(n10131), .B(n10132), .Z(n9934) );
  XOR2_X1 U10030 ( .A(n10133), .B(n10134), .Z(n10132) );
  XOR2_X1 U10031 ( .A(n10135), .B(n10136), .Z(n9938) );
  XOR2_X1 U10032 ( .A(n10137), .B(n10138), .Z(n10136) );
  OR2_X1 U10033 ( .A1(n7624), .A2(n8358), .ZN(n9945) );
  XOR2_X1 U10034 ( .A(n10139), .B(n10140), .Z(n9942) );
  XOR2_X1 U10035 ( .A(n10141), .B(n10142), .Z(n10140) );
  OR2_X1 U10036 ( .A1(n7622), .A2(n8358), .ZN(n9949) );
  XOR2_X1 U10037 ( .A(n10143), .B(n10144), .Z(n9946) );
  XOR2_X1 U10038 ( .A(n10145), .B(n10146), .Z(n10144) );
  OR2_X1 U10039 ( .A1(n7620), .A2(n8358), .ZN(n9953) );
  XOR2_X1 U10040 ( .A(n10147), .B(n10148), .Z(n9950) );
  XOR2_X1 U10041 ( .A(n10149), .B(n10150), .Z(n10148) );
  XOR2_X1 U10042 ( .A(n10151), .B(n10152), .Z(n9954) );
  XOR2_X1 U10043 ( .A(n10153), .B(n10154), .Z(n10152) );
  OR2_X1 U10044 ( .A1(n7616), .A2(n8358), .ZN(n9961) );
  XOR2_X1 U10045 ( .A(n10155), .B(n10156), .Z(n9958) );
  XOR2_X1 U10046 ( .A(n10157), .B(n10158), .Z(n10156) );
  OR2_X1 U10047 ( .A1(n8152), .A2(n8358), .ZN(n9965) );
  INV_X1 U10048 ( .A(n9650), .ZN(n8358) );
  XOR2_X1 U10049 ( .A(n10159), .B(n10160), .Z(n9650) );
  XNOR2_X1 U10050 ( .A(c_24_), .B(d_24_), .ZN(n10159) );
  XOR2_X1 U10051 ( .A(n10161), .B(n10162), .Z(n9962) );
  XOR2_X1 U10052 ( .A(n10163), .B(n10164), .Z(n10162) );
  XOR2_X1 U10053 ( .A(n10165), .B(n10166), .Z(n9968) );
  XOR2_X1 U10054 ( .A(n10167), .B(n10168), .Z(n10166) );
  XOR2_X1 U10055 ( .A(n9331), .B(n10169), .Z(n9341) );
  XOR2_X1 U10056 ( .A(n9330), .B(n9329), .Z(n10169) );
  OR2_X1 U10057 ( .A1(n8105), .A2(n8335), .ZN(n9329) );
  OR2_X1 U10058 ( .A1(n10170), .A2(n10171), .ZN(n9330) );
  AND2_X1 U10059 ( .A1(n10168), .A2(n10167), .ZN(n10171) );
  AND2_X1 U10060 ( .A1(n10165), .A2(n10172), .ZN(n10170) );
  OR2_X1 U10061 ( .A1(n10168), .A2(n10167), .ZN(n10172) );
  OR2_X1 U10062 ( .A1(n10173), .A2(n10174), .ZN(n10167) );
  AND2_X1 U10063 ( .A1(n10164), .A2(n10163), .ZN(n10174) );
  AND2_X1 U10064 ( .A1(n10161), .A2(n10175), .ZN(n10173) );
  OR2_X1 U10065 ( .A1(n10164), .A2(n10163), .ZN(n10175) );
  OR2_X1 U10066 ( .A1(n10176), .A2(n10177), .ZN(n10163) );
  AND2_X1 U10067 ( .A1(n10158), .A2(n10157), .ZN(n10177) );
  AND2_X1 U10068 ( .A1(n10155), .A2(n10178), .ZN(n10176) );
  OR2_X1 U10069 ( .A1(n10158), .A2(n10157), .ZN(n10178) );
  OR2_X1 U10070 ( .A1(n7618), .A2(n8335), .ZN(n10157) );
  OR2_X1 U10071 ( .A1(n10179), .A2(n10180), .ZN(n10158) );
  AND2_X1 U10072 ( .A1(n10154), .A2(n10153), .ZN(n10180) );
  AND2_X1 U10073 ( .A1(n10151), .A2(n10181), .ZN(n10179) );
  OR2_X1 U10074 ( .A1(n10154), .A2(n10153), .ZN(n10181) );
  OR2_X1 U10075 ( .A1(n10182), .A2(n10183), .ZN(n10153) );
  AND2_X1 U10076 ( .A1(n10150), .A2(n10149), .ZN(n10183) );
  AND2_X1 U10077 ( .A1(n10147), .A2(n10184), .ZN(n10182) );
  OR2_X1 U10078 ( .A1(n10150), .A2(n10149), .ZN(n10184) );
  OR2_X1 U10079 ( .A1(n10185), .A2(n10186), .ZN(n10149) );
  AND2_X1 U10080 ( .A1(n10146), .A2(n10145), .ZN(n10186) );
  AND2_X1 U10081 ( .A1(n10143), .A2(n10187), .ZN(n10185) );
  OR2_X1 U10082 ( .A1(n10146), .A2(n10145), .ZN(n10187) );
  OR2_X1 U10083 ( .A1(n10188), .A2(n10189), .ZN(n10145) );
  AND2_X1 U10084 ( .A1(n10142), .A2(n10141), .ZN(n10189) );
  AND2_X1 U10085 ( .A1(n10139), .A2(n10190), .ZN(n10188) );
  OR2_X1 U10086 ( .A1(n10142), .A2(n10141), .ZN(n10190) );
  OR2_X1 U10087 ( .A1(n7626), .A2(n8335), .ZN(n10141) );
  OR2_X1 U10088 ( .A1(n10191), .A2(n10192), .ZN(n10142) );
  AND2_X1 U10089 ( .A1(n10138), .A2(n10137), .ZN(n10192) );
  AND2_X1 U10090 ( .A1(n10135), .A2(n10193), .ZN(n10191) );
  OR2_X1 U10091 ( .A1(n10138), .A2(n10137), .ZN(n10193) );
  OR2_X1 U10092 ( .A1(n10194), .A2(n10195), .ZN(n10137) );
  AND2_X1 U10093 ( .A1(n10134), .A2(n10133), .ZN(n10195) );
  AND2_X1 U10094 ( .A1(n10131), .A2(n10196), .ZN(n10194) );
  OR2_X1 U10095 ( .A1(n10134), .A2(n10133), .ZN(n10196) );
  OR2_X1 U10096 ( .A1(n10197), .A2(n10198), .ZN(n10133) );
  AND2_X1 U10097 ( .A1(n10130), .A2(n10129), .ZN(n10198) );
  AND2_X1 U10098 ( .A1(n10127), .A2(n10199), .ZN(n10197) );
  OR2_X1 U10099 ( .A1(n10130), .A2(n10129), .ZN(n10199) );
  OR2_X1 U10100 ( .A1(n10200), .A2(n10201), .ZN(n10129) );
  AND2_X1 U10101 ( .A1(n10126), .A2(n10125), .ZN(n10201) );
  AND2_X1 U10102 ( .A1(n10123), .A2(n10202), .ZN(n10200) );
  OR2_X1 U10103 ( .A1(n10126), .A2(n10125), .ZN(n10202) );
  OR2_X1 U10104 ( .A1(n7634), .A2(n8335), .ZN(n10125) );
  OR2_X1 U10105 ( .A1(n10203), .A2(n10204), .ZN(n10126) );
  AND2_X1 U10106 ( .A1(n10122), .A2(n10121), .ZN(n10204) );
  AND2_X1 U10107 ( .A1(n10119), .A2(n10205), .ZN(n10203) );
  OR2_X1 U10108 ( .A1(n10122), .A2(n10121), .ZN(n10205) );
  OR2_X1 U10109 ( .A1(n10206), .A2(n10207), .ZN(n10121) );
  AND2_X1 U10110 ( .A1(n10118), .A2(n10117), .ZN(n10207) );
  AND2_X1 U10111 ( .A1(n10115), .A2(n10208), .ZN(n10206) );
  OR2_X1 U10112 ( .A1(n10118), .A2(n10117), .ZN(n10208) );
  OR2_X1 U10113 ( .A1(n10209), .A2(n10210), .ZN(n10117) );
  AND2_X1 U10114 ( .A1(n10114), .A2(n10113), .ZN(n10210) );
  AND2_X1 U10115 ( .A1(n10111), .A2(n10211), .ZN(n10209) );
  OR2_X1 U10116 ( .A1(n10114), .A2(n10113), .ZN(n10211) );
  OR2_X1 U10117 ( .A1(n10212), .A2(n10213), .ZN(n10113) );
  AND2_X1 U10118 ( .A1(n10110), .A2(n10109), .ZN(n10213) );
  AND2_X1 U10119 ( .A1(n10107), .A2(n10214), .ZN(n10212) );
  OR2_X1 U10120 ( .A1(n10110), .A2(n10109), .ZN(n10214) );
  OR2_X1 U10121 ( .A1(n10215), .A2(n10216), .ZN(n10109) );
  AND2_X1 U10122 ( .A1(n10106), .A2(n10105), .ZN(n10216) );
  AND2_X1 U10123 ( .A1(n10103), .A2(n10217), .ZN(n10215) );
  OR2_X1 U10124 ( .A1(n10106), .A2(n10105), .ZN(n10217) );
  OR2_X1 U10125 ( .A1(n10218), .A2(n10219), .ZN(n10105) );
  AND2_X1 U10126 ( .A1(n10102), .A2(n10101), .ZN(n10219) );
  AND2_X1 U10127 ( .A1(n10099), .A2(n10220), .ZN(n10218) );
  OR2_X1 U10128 ( .A1(n10102), .A2(n10101), .ZN(n10220) );
  OR2_X1 U10129 ( .A1(n10221), .A2(n10222), .ZN(n10101) );
  AND2_X1 U10130 ( .A1(n10098), .A2(n10097), .ZN(n10222) );
  AND2_X1 U10131 ( .A1(n10095), .A2(n10223), .ZN(n10221) );
  OR2_X1 U10132 ( .A1(n10098), .A2(n10097), .ZN(n10223) );
  OR2_X1 U10133 ( .A1(n10224), .A2(n10225), .ZN(n10097) );
  AND2_X1 U10134 ( .A1(n10094), .A2(n10093), .ZN(n10225) );
  AND2_X1 U10135 ( .A1(n10091), .A2(n10226), .ZN(n10224) );
  OR2_X1 U10136 ( .A1(n10094), .A2(n10093), .ZN(n10226) );
  OR2_X1 U10137 ( .A1(n10227), .A2(n10228), .ZN(n10093) );
  AND2_X1 U10138 ( .A1(n10090), .A2(n10089), .ZN(n10228) );
  AND2_X1 U10139 ( .A1(n10087), .A2(n10229), .ZN(n10227) );
  OR2_X1 U10140 ( .A1(n10090), .A2(n10089), .ZN(n10229) );
  OR2_X1 U10141 ( .A1(n10230), .A2(n10231), .ZN(n10089) );
  AND2_X1 U10142 ( .A1(n10086), .A2(n10085), .ZN(n10231) );
  AND2_X1 U10143 ( .A1(n10083), .A2(n10232), .ZN(n10230) );
  OR2_X1 U10144 ( .A1(n10086), .A2(n10085), .ZN(n10232) );
  OR2_X1 U10145 ( .A1(n10233), .A2(n10234), .ZN(n10085) );
  AND2_X1 U10146 ( .A1(n10082), .A2(n10081), .ZN(n10234) );
  AND2_X1 U10147 ( .A1(n10079), .A2(n10235), .ZN(n10233) );
  OR2_X1 U10148 ( .A1(n10082), .A2(n10081), .ZN(n10235) );
  OR2_X1 U10149 ( .A1(n10236), .A2(n10237), .ZN(n10081) );
  AND2_X1 U10150 ( .A1(n10078), .A2(n10077), .ZN(n10237) );
  AND2_X1 U10151 ( .A1(n10075), .A2(n10238), .ZN(n10236) );
  OR2_X1 U10152 ( .A1(n10078), .A2(n10077), .ZN(n10238) );
  OR2_X1 U10153 ( .A1(n10239), .A2(n10240), .ZN(n10077) );
  AND2_X1 U10154 ( .A1(n10074), .A2(n10073), .ZN(n10240) );
  AND2_X1 U10155 ( .A1(n10071), .A2(n10241), .ZN(n10239) );
  OR2_X1 U10156 ( .A1(n10074), .A2(n10073), .ZN(n10241) );
  OR2_X1 U10157 ( .A1(n10242), .A2(n10243), .ZN(n10073) );
  AND2_X1 U10158 ( .A1(n10070), .A2(n10069), .ZN(n10243) );
  AND2_X1 U10159 ( .A1(n10067), .A2(n10244), .ZN(n10242) );
  OR2_X1 U10160 ( .A1(n10070), .A2(n10069), .ZN(n10244) );
  OR2_X1 U10161 ( .A1(n10245), .A2(n10246), .ZN(n10069) );
  AND2_X1 U10162 ( .A1(n10063), .A2(n10066), .ZN(n10246) );
  AND2_X1 U10163 ( .A1(n10065), .A2(n10247), .ZN(n10245) );
  OR2_X1 U10164 ( .A1(n10063), .A2(n10066), .ZN(n10247) );
  OR3_X1 U10165 ( .A1(n10062), .A2(n8335), .A3(n8519), .ZN(n10066) );
  OR2_X1 U10166 ( .A1(n8335), .A2(n7606), .ZN(n10063) );
  INV_X1 U10167 ( .A(n10248), .ZN(n10065) );
  OR2_X1 U10168 ( .A1(n10249), .A2(n10250), .ZN(n10248) );
  AND2_X1 U10169 ( .A1(n10251), .A2(n10252), .ZN(n10250) );
  OR2_X1 U10170 ( .A1(n10253), .A2(n7697), .ZN(n10252) );
  AND2_X1 U10171 ( .A1(n10062), .A2(n7691), .ZN(n10253) );
  AND2_X1 U10172 ( .A1(n10057), .A2(n10254), .ZN(n10249) );
  OR2_X1 U10173 ( .A1(n10255), .A2(n7701), .ZN(n10254) );
  AND2_X1 U10174 ( .A1(n10256), .A2(n7703), .ZN(n10255) );
  OR2_X1 U10175 ( .A1(n7662), .A2(n8335), .ZN(n10070) );
  XNOR2_X1 U10176 ( .A(n10257), .B(n10258), .ZN(n10067) );
  XNOR2_X1 U10177 ( .A(n10259), .B(n10260), .ZN(n10258) );
  OR2_X1 U10178 ( .A1(n7660), .A2(n8335), .ZN(n10074) );
  XOR2_X1 U10179 ( .A(n10261), .B(n10262), .Z(n10071) );
  XOR2_X1 U10180 ( .A(n10263), .B(n10264), .Z(n10262) );
  OR2_X1 U10181 ( .A1(n7658), .A2(n8335), .ZN(n10078) );
  XOR2_X1 U10182 ( .A(n10265), .B(n10266), .Z(n10075) );
  XOR2_X1 U10183 ( .A(n10267), .B(n10268), .Z(n10266) );
  OR2_X1 U10184 ( .A1(n7656), .A2(n8335), .ZN(n10082) );
  XOR2_X1 U10185 ( .A(n10269), .B(n10270), .Z(n10079) );
  XOR2_X1 U10186 ( .A(n10271), .B(n10272), .Z(n10270) );
  OR2_X1 U10187 ( .A1(n7654), .A2(n8335), .ZN(n10086) );
  XOR2_X1 U10188 ( .A(n10273), .B(n10274), .Z(n10083) );
  XOR2_X1 U10189 ( .A(n10275), .B(n10276), .Z(n10274) );
  OR2_X1 U10190 ( .A1(n7652), .A2(n8335), .ZN(n10090) );
  XOR2_X1 U10191 ( .A(n10277), .B(n10278), .Z(n10087) );
  XOR2_X1 U10192 ( .A(n10279), .B(n10280), .Z(n10278) );
  OR2_X1 U10193 ( .A1(n7650), .A2(n8335), .ZN(n10094) );
  XOR2_X1 U10194 ( .A(n10281), .B(n10282), .Z(n10091) );
  XOR2_X1 U10195 ( .A(n10283), .B(n10284), .Z(n10282) );
  OR2_X1 U10196 ( .A1(n7648), .A2(n8335), .ZN(n10098) );
  XOR2_X1 U10197 ( .A(n10285), .B(n10286), .Z(n10095) );
  XOR2_X1 U10198 ( .A(n10287), .B(n10288), .Z(n10286) );
  OR2_X1 U10199 ( .A1(n7646), .A2(n8335), .ZN(n10102) );
  XOR2_X1 U10200 ( .A(n10289), .B(n10290), .Z(n10099) );
  XOR2_X1 U10201 ( .A(n10291), .B(n10292), .Z(n10290) );
  OR2_X1 U10202 ( .A1(n7644), .A2(n8335), .ZN(n10106) );
  XOR2_X1 U10203 ( .A(n10293), .B(n10294), .Z(n10103) );
  XOR2_X1 U10204 ( .A(n10295), .B(n10296), .Z(n10294) );
  OR2_X1 U10205 ( .A1(n7642), .A2(n8335), .ZN(n10110) );
  XOR2_X1 U10206 ( .A(n10297), .B(n10298), .Z(n10107) );
  XOR2_X1 U10207 ( .A(n10299), .B(n10300), .Z(n10298) );
  OR2_X1 U10208 ( .A1(n7640), .A2(n8335), .ZN(n10114) );
  XOR2_X1 U10209 ( .A(n10301), .B(n10302), .Z(n10111) );
  XOR2_X1 U10210 ( .A(n10303), .B(n10304), .Z(n10302) );
  OR2_X1 U10211 ( .A1(n7638), .A2(n8335), .ZN(n10118) );
  XOR2_X1 U10212 ( .A(n10305), .B(n10306), .Z(n10115) );
  XOR2_X1 U10213 ( .A(n10307), .B(n10308), .Z(n10306) );
  OR2_X1 U10214 ( .A1(n7636), .A2(n8335), .ZN(n10122) );
  XOR2_X1 U10215 ( .A(n10309), .B(n10310), .Z(n10119) );
  XOR2_X1 U10216 ( .A(n10311), .B(n10312), .Z(n10310) );
  XOR2_X1 U10217 ( .A(n10313), .B(n10314), .Z(n10123) );
  XOR2_X1 U10218 ( .A(n10315), .B(n10316), .Z(n10314) );
  OR2_X1 U10219 ( .A1(n7632), .A2(n8335), .ZN(n10130) );
  XOR2_X1 U10220 ( .A(n10317), .B(n10318), .Z(n10127) );
  XOR2_X1 U10221 ( .A(n10319), .B(n10320), .Z(n10318) );
  OR2_X1 U10222 ( .A1(n7630), .A2(n8335), .ZN(n10134) );
  XOR2_X1 U10223 ( .A(n10321), .B(n10322), .Z(n10131) );
  XOR2_X1 U10224 ( .A(n10323), .B(n10324), .Z(n10322) );
  OR2_X1 U10225 ( .A1(n7628), .A2(n8335), .ZN(n10138) );
  XOR2_X1 U10226 ( .A(n10325), .B(n10326), .Z(n10135) );
  XOR2_X1 U10227 ( .A(n10327), .B(n10328), .Z(n10326) );
  XOR2_X1 U10228 ( .A(n10329), .B(n10330), .Z(n10139) );
  XOR2_X1 U10229 ( .A(n10331), .B(n10332), .Z(n10330) );
  OR2_X1 U10230 ( .A1(n7624), .A2(n8335), .ZN(n10146) );
  XOR2_X1 U10231 ( .A(n10333), .B(n10334), .Z(n10143) );
  XOR2_X1 U10232 ( .A(n10335), .B(n10336), .Z(n10334) );
  OR2_X1 U10233 ( .A1(n7622), .A2(n8335), .ZN(n10150) );
  XOR2_X1 U10234 ( .A(n10337), .B(n10338), .Z(n10147) );
  XOR2_X1 U10235 ( .A(n10339), .B(n10340), .Z(n10338) );
  OR2_X1 U10236 ( .A1(n7620), .A2(n8335), .ZN(n10154) );
  XOR2_X1 U10237 ( .A(n10341), .B(n10342), .Z(n10151) );
  XOR2_X1 U10238 ( .A(n10343), .B(n10344), .Z(n10342) );
  XOR2_X1 U10239 ( .A(n10345), .B(n10346), .Z(n10155) );
  XOR2_X1 U10240 ( .A(n10347), .B(n10348), .Z(n10346) );
  OR2_X1 U10241 ( .A1(n8644), .A2(n8335), .ZN(n10164) );
  XOR2_X1 U10242 ( .A(n10349), .B(n10350), .Z(n10161) );
  XOR2_X1 U10243 ( .A(n10351), .B(n10352), .Z(n10350) );
  OR2_X1 U10244 ( .A1(n8152), .A2(n8335), .ZN(n10168) );
  INV_X1 U10245 ( .A(n9857), .ZN(n8335) );
  XOR2_X1 U10246 ( .A(n10353), .B(n10354), .Z(n9857) );
  XNOR2_X1 U10247 ( .A(c_23_), .B(d_23_), .ZN(n10353) );
  XOR2_X1 U10248 ( .A(n10355), .B(n10356), .Z(n10165) );
  XOR2_X1 U10249 ( .A(n10357), .B(n10358), .Z(n10356) );
  XOR2_X1 U10250 ( .A(n10359), .B(n10360), .Z(n9331) );
  XOR2_X1 U10251 ( .A(n10361), .B(n10362), .Z(n10360) );
  INV_X1 U10252 ( .A(n10363), .ZN(n7895) );
  OR2_X1 U10253 ( .A1(n10364), .A2(n8301), .ZN(n10363) );
  XOR2_X1 U10254 ( .A(n8262), .B(n8264), .Z(n8301) );
  OR2_X1 U10255 ( .A1(n10365), .A2(n10366), .ZN(n8264) );
  AND2_X1 U10256 ( .A1(n10367), .A2(n10368), .ZN(n10366) );
  AND2_X1 U10257 ( .A1(n10369), .A2(n10370), .ZN(n10365) );
  OR2_X1 U10258 ( .A1(n10367), .A2(n10368), .ZN(n10370) );
  XOR2_X1 U10259 ( .A(n8270), .B(n10371), .Z(n8262) );
  XOR2_X1 U10260 ( .A(n8269), .B(n8268), .Z(n10371) );
  OR2_X1 U10261 ( .A1(n10372), .A2(n7664), .ZN(n8268) );
  OR2_X1 U10262 ( .A1(n10373), .A2(n10374), .ZN(n8269) );
  AND2_X1 U10263 ( .A1(n10375), .A2(n10376), .ZN(n10374) );
  AND2_X1 U10264 ( .A1(n10377), .A2(n10378), .ZN(n10373) );
  OR2_X1 U10265 ( .A1(n10375), .A2(n10376), .ZN(n10378) );
  XOR2_X1 U10266 ( .A(n8278), .B(n10379), .Z(n8270) );
  XOR2_X1 U10267 ( .A(n8277), .B(n8276), .Z(n10379) );
  OR2_X1 U10268 ( .A1(n8023), .A2(n8273), .ZN(n8276) );
  OR2_X1 U10269 ( .A1(n10380), .A2(n10381), .ZN(n8277) );
  AND2_X1 U10270 ( .A1(n10382), .A2(n10383), .ZN(n10381) );
  AND2_X1 U10271 ( .A1(n10384), .A2(n10385), .ZN(n10380) );
  OR2_X1 U10272 ( .A1(n10382), .A2(n10383), .ZN(n10385) );
  XOR2_X1 U10273 ( .A(n8285), .B(n10386), .Z(n8278) );
  XOR2_X1 U10274 ( .A(n8284), .B(n8283), .Z(n10386) );
  OR2_X1 U10275 ( .A1(n8056), .A2(n8243), .ZN(n8283) );
  OR2_X1 U10276 ( .A1(n10387), .A2(n10388), .ZN(n8284) );
  AND2_X1 U10277 ( .A1(n10389), .A2(n10390), .ZN(n10388) );
  AND2_X1 U10278 ( .A1(n10391), .A2(n10392), .ZN(n10387) );
  OR2_X1 U10279 ( .A1(n10389), .A2(n10390), .ZN(n10392) );
  XOR2_X1 U10280 ( .A(n8292), .B(n10393), .Z(n8285) );
  XOR2_X1 U10281 ( .A(n8291), .B(n8290), .Z(n10393) );
  OR2_X1 U10282 ( .A1(n8105), .A2(n8220), .ZN(n8290) );
  OR2_X1 U10283 ( .A1(n10394), .A2(n10395), .ZN(n8291) );
  AND2_X1 U10284 ( .A1(n10396), .A2(n10397), .ZN(n10395) );
  AND2_X1 U10285 ( .A1(n10398), .A2(n10399), .ZN(n10394) );
  OR2_X1 U10286 ( .A1(n10396), .A2(n10397), .ZN(n10399) );
  XOR2_X1 U10287 ( .A(n10400), .B(n10401), .Z(n8292) );
  XOR2_X1 U10288 ( .A(n10402), .B(n10403), .Z(n10401) );
  AND2_X1 U10289 ( .A1(n8302), .A2(n8300), .ZN(n10364) );
  XNOR2_X1 U10290 ( .A(n10369), .B(n10404), .ZN(n8300) );
  XOR2_X1 U10291 ( .A(n10368), .B(n10367), .Z(n10404) );
  OR2_X1 U10292 ( .A1(n10256), .A2(n7664), .ZN(n10367) );
  OR2_X1 U10293 ( .A1(n10405), .A2(n10406), .ZN(n10368) );
  AND2_X1 U10294 ( .A1(n10407), .A2(n10408), .ZN(n10406) );
  AND2_X1 U10295 ( .A1(n10409), .A2(n10410), .ZN(n10405) );
  OR2_X1 U10296 ( .A1(n10407), .A2(n10408), .ZN(n10410) );
  XOR2_X1 U10297 ( .A(n10377), .B(n10411), .Z(n10369) );
  XOR2_X1 U10298 ( .A(n10376), .B(n10375), .Z(n10411) );
  OR2_X1 U10299 ( .A1(n8023), .A2(n10372), .ZN(n10375) );
  OR2_X1 U10300 ( .A1(n10412), .A2(n10413), .ZN(n10376) );
  AND2_X1 U10301 ( .A1(n10414), .A2(n10415), .ZN(n10413) );
  AND2_X1 U10302 ( .A1(n10416), .A2(n10417), .ZN(n10412) );
  OR2_X1 U10303 ( .A1(n10414), .A2(n10415), .ZN(n10417) );
  XOR2_X1 U10304 ( .A(n10384), .B(n10418), .Z(n10377) );
  XOR2_X1 U10305 ( .A(n10383), .B(n10382), .Z(n10418) );
  OR2_X1 U10306 ( .A1(n8056), .A2(n8273), .ZN(n10382) );
  OR2_X1 U10307 ( .A1(n10419), .A2(n10420), .ZN(n10383) );
  AND2_X1 U10308 ( .A1(n10421), .A2(n10422), .ZN(n10420) );
  AND2_X1 U10309 ( .A1(n10423), .A2(n10424), .ZN(n10419) );
  OR2_X1 U10310 ( .A1(n10421), .A2(n10422), .ZN(n10424) );
  XOR2_X1 U10311 ( .A(n10391), .B(n10425), .Z(n10384) );
  XOR2_X1 U10312 ( .A(n10390), .B(n10389), .Z(n10425) );
  OR2_X1 U10313 ( .A1(n8105), .A2(n8243), .ZN(n10389) );
  OR2_X1 U10314 ( .A1(n10426), .A2(n10427), .ZN(n10390) );
  AND2_X1 U10315 ( .A1(n10428), .A2(n10429), .ZN(n10427) );
  AND2_X1 U10316 ( .A1(n10430), .A2(n10431), .ZN(n10426) );
  OR2_X1 U10317 ( .A1(n10428), .A2(n10429), .ZN(n10431) );
  XOR2_X1 U10318 ( .A(n10398), .B(n10432), .Z(n10391) );
  XOR2_X1 U10319 ( .A(n10397), .B(n10396), .Z(n10432) );
  OR2_X1 U10320 ( .A1(n8152), .A2(n8220), .ZN(n10396) );
  OR2_X1 U10321 ( .A1(n10433), .A2(n10434), .ZN(n10397) );
  AND2_X1 U10322 ( .A1(n10435), .A2(n10436), .ZN(n10434) );
  AND2_X1 U10323 ( .A1(n10437), .A2(n10438), .ZN(n10433) );
  OR2_X1 U10324 ( .A1(n10435), .A2(n10436), .ZN(n10438) );
  XOR2_X1 U10325 ( .A(n10439), .B(n10440), .Z(n10398) );
  XOR2_X1 U10326 ( .A(n10441), .B(n10442), .Z(n10440) );
  INV_X1 U10327 ( .A(n10443), .ZN(n8302) );
  OR2_X1 U10328 ( .A1(n10444), .A2(n10445), .ZN(n10443) );
  AND2_X1 U10329 ( .A1(n8322), .A2(n8321), .ZN(n10445) );
  AND2_X1 U10330 ( .A1(n8319), .A2(n10446), .ZN(n10444) );
  OR2_X1 U10331 ( .A1(n8321), .A2(n8322), .ZN(n10446) );
  OR2_X1 U10332 ( .A1(n10062), .A2(n7664), .ZN(n8322) );
  OR2_X1 U10333 ( .A1(n10447), .A2(n10448), .ZN(n8321) );
  AND2_X1 U10334 ( .A1(n8345), .A2(n8344), .ZN(n10448) );
  AND2_X1 U10335 ( .A1(n8342), .A2(n10449), .ZN(n10447) );
  OR2_X1 U10336 ( .A1(n8344), .A2(n8345), .ZN(n10449) );
  OR2_X1 U10337 ( .A1(n8023), .A2(n10062), .ZN(n8345) );
  OR2_X1 U10338 ( .A1(n10450), .A2(n10451), .ZN(n8344) );
  AND2_X1 U10339 ( .A1(n8375), .A2(n8374), .ZN(n10451) );
  AND2_X1 U10340 ( .A1(n8372), .A2(n10452), .ZN(n10450) );
  OR2_X1 U10341 ( .A1(n8374), .A2(n8375), .ZN(n10452) );
  OR2_X1 U10342 ( .A1(n8056), .A2(n10062), .ZN(n8375) );
  OR2_X1 U10343 ( .A1(n10453), .A2(n10454), .ZN(n8374) );
  AND2_X1 U10344 ( .A1(n9336), .A2(n9335), .ZN(n10454) );
  AND2_X1 U10345 ( .A1(n9333), .A2(n10455), .ZN(n10453) );
  OR2_X1 U10346 ( .A1(n9335), .A2(n9336), .ZN(n10455) );
  OR2_X1 U10347 ( .A1(n8105), .A2(n10062), .ZN(n9336) );
  OR2_X1 U10348 ( .A1(n10456), .A2(n10457), .ZN(n9335) );
  AND2_X1 U10349 ( .A1(n10362), .A2(n10361), .ZN(n10457) );
  AND2_X1 U10350 ( .A1(n10359), .A2(n10458), .ZN(n10456) );
  OR2_X1 U10351 ( .A1(n10361), .A2(n10362), .ZN(n10458) );
  OR2_X1 U10352 ( .A1(n8152), .A2(n10062), .ZN(n10362) );
  OR2_X1 U10353 ( .A1(n10459), .A2(n10460), .ZN(n10361) );
  AND2_X1 U10354 ( .A1(n10358), .A2(n10357), .ZN(n10460) );
  AND2_X1 U10355 ( .A1(n10355), .A2(n10461), .ZN(n10459) );
  OR2_X1 U10356 ( .A1(n10357), .A2(n10358), .ZN(n10461) );
  OR2_X1 U10357 ( .A1(n8644), .A2(n10062), .ZN(n10358) );
  OR2_X1 U10358 ( .A1(n10462), .A2(n10463), .ZN(n10357) );
  AND2_X1 U10359 ( .A1(n10352), .A2(n10351), .ZN(n10463) );
  AND2_X1 U10360 ( .A1(n10349), .A2(n10464), .ZN(n10462) );
  OR2_X1 U10361 ( .A1(n10351), .A2(n10352), .ZN(n10464) );
  OR2_X1 U10362 ( .A1(n8639), .A2(n10062), .ZN(n10352) );
  OR2_X1 U10363 ( .A1(n10465), .A2(n10466), .ZN(n10351) );
  AND2_X1 U10364 ( .A1(n10348), .A2(n10347), .ZN(n10466) );
  AND2_X1 U10365 ( .A1(n10345), .A2(n10467), .ZN(n10465) );
  OR2_X1 U10366 ( .A1(n10347), .A2(n10348), .ZN(n10467) );
  OR2_X1 U10367 ( .A1(n7620), .A2(n10062), .ZN(n10348) );
  OR2_X1 U10368 ( .A1(n10468), .A2(n10469), .ZN(n10347) );
  AND2_X1 U10369 ( .A1(n10344), .A2(n10343), .ZN(n10469) );
  AND2_X1 U10370 ( .A1(n10341), .A2(n10470), .ZN(n10468) );
  OR2_X1 U10371 ( .A1(n10343), .A2(n10344), .ZN(n10470) );
  OR2_X1 U10372 ( .A1(n7622), .A2(n10062), .ZN(n10344) );
  OR2_X1 U10373 ( .A1(n10471), .A2(n10472), .ZN(n10343) );
  AND2_X1 U10374 ( .A1(n10340), .A2(n10339), .ZN(n10472) );
  AND2_X1 U10375 ( .A1(n10337), .A2(n10473), .ZN(n10471) );
  OR2_X1 U10376 ( .A1(n10339), .A2(n10340), .ZN(n10473) );
  OR2_X1 U10377 ( .A1(n7624), .A2(n10062), .ZN(n10340) );
  OR2_X1 U10378 ( .A1(n10474), .A2(n10475), .ZN(n10339) );
  AND2_X1 U10379 ( .A1(n10336), .A2(n10335), .ZN(n10475) );
  AND2_X1 U10380 ( .A1(n10333), .A2(n10476), .ZN(n10474) );
  OR2_X1 U10381 ( .A1(n10335), .A2(n10336), .ZN(n10476) );
  OR2_X1 U10382 ( .A1(n7626), .A2(n10062), .ZN(n10336) );
  OR2_X1 U10383 ( .A1(n10477), .A2(n10478), .ZN(n10335) );
  AND2_X1 U10384 ( .A1(n10332), .A2(n10331), .ZN(n10478) );
  AND2_X1 U10385 ( .A1(n10329), .A2(n10479), .ZN(n10477) );
  OR2_X1 U10386 ( .A1(n10331), .A2(n10332), .ZN(n10479) );
  OR2_X1 U10387 ( .A1(n7628), .A2(n10062), .ZN(n10332) );
  OR2_X1 U10388 ( .A1(n10480), .A2(n10481), .ZN(n10331) );
  AND2_X1 U10389 ( .A1(n10328), .A2(n10327), .ZN(n10481) );
  AND2_X1 U10390 ( .A1(n10325), .A2(n10482), .ZN(n10480) );
  OR2_X1 U10391 ( .A1(n10327), .A2(n10328), .ZN(n10482) );
  OR2_X1 U10392 ( .A1(n7630), .A2(n10062), .ZN(n10328) );
  OR2_X1 U10393 ( .A1(n10483), .A2(n10484), .ZN(n10327) );
  AND2_X1 U10394 ( .A1(n10324), .A2(n10323), .ZN(n10484) );
  AND2_X1 U10395 ( .A1(n10321), .A2(n10485), .ZN(n10483) );
  OR2_X1 U10396 ( .A1(n10323), .A2(n10324), .ZN(n10485) );
  OR2_X1 U10397 ( .A1(n7632), .A2(n10062), .ZN(n10324) );
  OR2_X1 U10398 ( .A1(n10486), .A2(n10487), .ZN(n10323) );
  AND2_X1 U10399 ( .A1(n10320), .A2(n10319), .ZN(n10487) );
  AND2_X1 U10400 ( .A1(n10317), .A2(n10488), .ZN(n10486) );
  OR2_X1 U10401 ( .A1(n10319), .A2(n10320), .ZN(n10488) );
  OR2_X1 U10402 ( .A1(n7634), .A2(n10062), .ZN(n10320) );
  OR2_X1 U10403 ( .A1(n10489), .A2(n10490), .ZN(n10319) );
  AND2_X1 U10404 ( .A1(n10316), .A2(n10315), .ZN(n10490) );
  AND2_X1 U10405 ( .A1(n10313), .A2(n10491), .ZN(n10489) );
  OR2_X1 U10406 ( .A1(n10315), .A2(n10316), .ZN(n10491) );
  OR2_X1 U10407 ( .A1(n7636), .A2(n10062), .ZN(n10316) );
  OR2_X1 U10408 ( .A1(n10492), .A2(n10493), .ZN(n10315) );
  AND2_X1 U10409 ( .A1(n10312), .A2(n10311), .ZN(n10493) );
  AND2_X1 U10410 ( .A1(n10309), .A2(n10494), .ZN(n10492) );
  OR2_X1 U10411 ( .A1(n10311), .A2(n10312), .ZN(n10494) );
  OR2_X1 U10412 ( .A1(n7638), .A2(n10062), .ZN(n10312) );
  OR2_X1 U10413 ( .A1(n10495), .A2(n10496), .ZN(n10311) );
  AND2_X1 U10414 ( .A1(n10308), .A2(n10307), .ZN(n10496) );
  AND2_X1 U10415 ( .A1(n10305), .A2(n10497), .ZN(n10495) );
  OR2_X1 U10416 ( .A1(n10307), .A2(n10308), .ZN(n10497) );
  OR2_X1 U10417 ( .A1(n7640), .A2(n10062), .ZN(n10308) );
  OR2_X1 U10418 ( .A1(n10498), .A2(n10499), .ZN(n10307) );
  AND2_X1 U10419 ( .A1(n10304), .A2(n10303), .ZN(n10499) );
  AND2_X1 U10420 ( .A1(n10301), .A2(n10500), .ZN(n10498) );
  OR2_X1 U10421 ( .A1(n10303), .A2(n10304), .ZN(n10500) );
  OR2_X1 U10422 ( .A1(n7642), .A2(n10062), .ZN(n10304) );
  OR2_X1 U10423 ( .A1(n10501), .A2(n10502), .ZN(n10303) );
  AND2_X1 U10424 ( .A1(n10300), .A2(n10299), .ZN(n10502) );
  AND2_X1 U10425 ( .A1(n10297), .A2(n10503), .ZN(n10501) );
  OR2_X1 U10426 ( .A1(n10299), .A2(n10300), .ZN(n10503) );
  OR2_X1 U10427 ( .A1(n7644), .A2(n10062), .ZN(n10300) );
  OR2_X1 U10428 ( .A1(n10504), .A2(n10505), .ZN(n10299) );
  AND2_X1 U10429 ( .A1(n10296), .A2(n10295), .ZN(n10505) );
  AND2_X1 U10430 ( .A1(n10293), .A2(n10506), .ZN(n10504) );
  OR2_X1 U10431 ( .A1(n10295), .A2(n10296), .ZN(n10506) );
  OR2_X1 U10432 ( .A1(n7646), .A2(n10062), .ZN(n10296) );
  OR2_X1 U10433 ( .A1(n10507), .A2(n10508), .ZN(n10295) );
  AND2_X1 U10434 ( .A1(n10292), .A2(n10291), .ZN(n10508) );
  AND2_X1 U10435 ( .A1(n10289), .A2(n10509), .ZN(n10507) );
  OR2_X1 U10436 ( .A1(n10291), .A2(n10292), .ZN(n10509) );
  OR2_X1 U10437 ( .A1(n7648), .A2(n10062), .ZN(n10292) );
  OR2_X1 U10438 ( .A1(n10510), .A2(n10511), .ZN(n10291) );
  AND2_X1 U10439 ( .A1(n10288), .A2(n10287), .ZN(n10511) );
  AND2_X1 U10440 ( .A1(n10285), .A2(n10512), .ZN(n10510) );
  OR2_X1 U10441 ( .A1(n10287), .A2(n10288), .ZN(n10512) );
  OR2_X1 U10442 ( .A1(n7650), .A2(n10062), .ZN(n10288) );
  OR2_X1 U10443 ( .A1(n10513), .A2(n10514), .ZN(n10287) );
  AND2_X1 U10444 ( .A1(n10284), .A2(n10283), .ZN(n10514) );
  AND2_X1 U10445 ( .A1(n10281), .A2(n10515), .ZN(n10513) );
  OR2_X1 U10446 ( .A1(n10283), .A2(n10284), .ZN(n10515) );
  OR2_X1 U10447 ( .A1(n7652), .A2(n10062), .ZN(n10284) );
  OR2_X1 U10448 ( .A1(n10516), .A2(n10517), .ZN(n10283) );
  AND2_X1 U10449 ( .A1(n10280), .A2(n10279), .ZN(n10517) );
  AND2_X1 U10450 ( .A1(n10277), .A2(n10518), .ZN(n10516) );
  OR2_X1 U10451 ( .A1(n10279), .A2(n10280), .ZN(n10518) );
  OR2_X1 U10452 ( .A1(n7654), .A2(n10062), .ZN(n10280) );
  OR2_X1 U10453 ( .A1(n10519), .A2(n10520), .ZN(n10279) );
  AND2_X1 U10454 ( .A1(n10276), .A2(n10275), .ZN(n10520) );
  AND2_X1 U10455 ( .A1(n10273), .A2(n10521), .ZN(n10519) );
  OR2_X1 U10456 ( .A1(n10275), .A2(n10276), .ZN(n10521) );
  OR2_X1 U10457 ( .A1(n7656), .A2(n10062), .ZN(n10276) );
  OR2_X1 U10458 ( .A1(n10522), .A2(n10523), .ZN(n10275) );
  AND2_X1 U10459 ( .A1(n10272), .A2(n10271), .ZN(n10523) );
  AND2_X1 U10460 ( .A1(n10269), .A2(n10524), .ZN(n10522) );
  OR2_X1 U10461 ( .A1(n10271), .A2(n10272), .ZN(n10524) );
  OR2_X1 U10462 ( .A1(n7658), .A2(n10062), .ZN(n10272) );
  OR2_X1 U10463 ( .A1(n10525), .A2(n10526), .ZN(n10271) );
  AND2_X1 U10464 ( .A1(n10268), .A2(n10267), .ZN(n10526) );
  AND2_X1 U10465 ( .A1(n10265), .A2(n10527), .ZN(n10525) );
  OR2_X1 U10466 ( .A1(n10267), .A2(n10268), .ZN(n10527) );
  OR2_X1 U10467 ( .A1(n7660), .A2(n10062), .ZN(n10268) );
  OR2_X1 U10468 ( .A1(n10528), .A2(n10529), .ZN(n10267) );
  AND2_X1 U10469 ( .A1(n10264), .A2(n10263), .ZN(n10529) );
  AND2_X1 U10470 ( .A1(n10261), .A2(n10530), .ZN(n10528) );
  OR2_X1 U10471 ( .A1(n10263), .A2(n10264), .ZN(n10530) );
  OR2_X1 U10472 ( .A1(n7662), .A2(n10062), .ZN(n10264) );
  OR2_X1 U10473 ( .A1(n10531), .A2(n10532), .ZN(n10263) );
  AND2_X1 U10474 ( .A1(n10257), .A2(n10260), .ZN(n10532) );
  AND2_X1 U10475 ( .A1(n10259), .A2(n10533), .ZN(n10531) );
  OR2_X1 U10476 ( .A1(n10260), .A2(n10257), .ZN(n10533) );
  OR2_X1 U10477 ( .A1(n10062), .A2(n7606), .ZN(n10257) );
  OR3_X1 U10478 ( .A1(n10256), .A2(n10062), .A3(n8519), .ZN(n10260) );
  INV_X1 U10479 ( .A(n10057), .ZN(n10062) );
  XOR2_X1 U10480 ( .A(n10534), .B(n10535), .Z(n10057) );
  XNOR2_X1 U10481 ( .A(c_22_), .B(d_22_), .ZN(n10534) );
  INV_X1 U10482 ( .A(n10536), .ZN(n10259) );
  OR2_X1 U10483 ( .A1(n10537), .A2(n10538), .ZN(n10536) );
  AND2_X1 U10484 ( .A1(n10539), .A2(n10540), .ZN(n10538) );
  OR2_X1 U10485 ( .A1(n10541), .A2(n7697), .ZN(n10540) );
  AND2_X1 U10486 ( .A1(n10256), .A2(n7691), .ZN(n10541) );
  AND2_X1 U10487 ( .A1(n10251), .A2(n10542), .ZN(n10537) );
  OR2_X1 U10488 ( .A1(n10543), .A2(n7701), .ZN(n10542) );
  AND2_X1 U10489 ( .A1(n10372), .A2(n7703), .ZN(n10543) );
  XNOR2_X1 U10490 ( .A(n10544), .B(n10545), .ZN(n10261) );
  XNOR2_X1 U10491 ( .A(n10546), .B(n10547), .ZN(n10545) );
  XOR2_X1 U10492 ( .A(n10548), .B(n10549), .Z(n10265) );
  XOR2_X1 U10493 ( .A(n10550), .B(n10551), .Z(n10549) );
  XOR2_X1 U10494 ( .A(n10552), .B(n10553), .Z(n10269) );
  XOR2_X1 U10495 ( .A(n10554), .B(n10555), .Z(n10553) );
  XOR2_X1 U10496 ( .A(n10556), .B(n10557), .Z(n10273) );
  XOR2_X1 U10497 ( .A(n10558), .B(n10559), .Z(n10557) );
  XOR2_X1 U10498 ( .A(n10560), .B(n10561), .Z(n10277) );
  XOR2_X1 U10499 ( .A(n10562), .B(n10563), .Z(n10561) );
  XOR2_X1 U10500 ( .A(n10564), .B(n10565), .Z(n10281) );
  XOR2_X1 U10501 ( .A(n10566), .B(n10567), .Z(n10565) );
  XOR2_X1 U10502 ( .A(n10568), .B(n10569), .Z(n10285) );
  XOR2_X1 U10503 ( .A(n10570), .B(n10571), .Z(n10569) );
  XOR2_X1 U10504 ( .A(n10572), .B(n10573), .Z(n10289) );
  XOR2_X1 U10505 ( .A(n10574), .B(n10575), .Z(n10573) );
  XOR2_X1 U10506 ( .A(n10576), .B(n10577), .Z(n10293) );
  XOR2_X1 U10507 ( .A(n10578), .B(n10579), .Z(n10577) );
  XOR2_X1 U10508 ( .A(n10580), .B(n10581), .Z(n10297) );
  XOR2_X1 U10509 ( .A(n10582), .B(n10583), .Z(n10581) );
  XOR2_X1 U10510 ( .A(n10584), .B(n10585), .Z(n10301) );
  XOR2_X1 U10511 ( .A(n10586), .B(n10587), .Z(n10585) );
  XOR2_X1 U10512 ( .A(n10588), .B(n10589), .Z(n10305) );
  XOR2_X1 U10513 ( .A(n10590), .B(n10591), .Z(n10589) );
  XOR2_X1 U10514 ( .A(n10592), .B(n10593), .Z(n10309) );
  XOR2_X1 U10515 ( .A(n10594), .B(n10595), .Z(n10593) );
  XOR2_X1 U10516 ( .A(n10596), .B(n10597), .Z(n10313) );
  XOR2_X1 U10517 ( .A(n10598), .B(n10599), .Z(n10597) );
  XOR2_X1 U10518 ( .A(n10600), .B(n10601), .Z(n10317) );
  XOR2_X1 U10519 ( .A(n10602), .B(n10603), .Z(n10601) );
  XOR2_X1 U10520 ( .A(n10604), .B(n10605), .Z(n10321) );
  XOR2_X1 U10521 ( .A(n10606), .B(n10607), .Z(n10605) );
  XOR2_X1 U10522 ( .A(n10608), .B(n10609), .Z(n10325) );
  XOR2_X1 U10523 ( .A(n10610), .B(n10611), .Z(n10609) );
  XOR2_X1 U10524 ( .A(n10612), .B(n10613), .Z(n10329) );
  XOR2_X1 U10525 ( .A(n10614), .B(n10615), .Z(n10613) );
  XOR2_X1 U10526 ( .A(n10616), .B(n10617), .Z(n10333) );
  XOR2_X1 U10527 ( .A(n10618), .B(n10619), .Z(n10617) );
  XOR2_X1 U10528 ( .A(n10620), .B(n10621), .Z(n10337) );
  XOR2_X1 U10529 ( .A(n10622), .B(n10623), .Z(n10621) );
  XOR2_X1 U10530 ( .A(n10624), .B(n10625), .Z(n10341) );
  XOR2_X1 U10531 ( .A(n10626), .B(n10627), .Z(n10625) );
  XOR2_X1 U10532 ( .A(n10628), .B(n10629), .Z(n10345) );
  XOR2_X1 U10533 ( .A(n10630), .B(n10631), .Z(n10629) );
  XOR2_X1 U10534 ( .A(n10632), .B(n10633), .Z(n10349) );
  XOR2_X1 U10535 ( .A(n10634), .B(n10635), .Z(n10633) );
  XOR2_X1 U10536 ( .A(n10636), .B(n10637), .Z(n10355) );
  XOR2_X1 U10537 ( .A(n10638), .B(n10639), .Z(n10637) );
  XOR2_X1 U10538 ( .A(n10640), .B(n10641), .Z(n10359) );
  XOR2_X1 U10539 ( .A(n10642), .B(n10643), .Z(n10641) );
  XOR2_X1 U10540 ( .A(n10644), .B(n10645), .Z(n9333) );
  XOR2_X1 U10541 ( .A(n10646), .B(n10647), .Z(n10645) );
  XOR2_X1 U10542 ( .A(n10648), .B(n10649), .Z(n8372) );
  XOR2_X1 U10543 ( .A(n10650), .B(n10651), .Z(n10649) );
  XOR2_X1 U10544 ( .A(n10652), .B(n10653), .Z(n8342) );
  XOR2_X1 U10545 ( .A(n10654), .B(n10655), .Z(n10653) );
  XOR2_X1 U10546 ( .A(n10409), .B(n10656), .Z(n8319) );
  XOR2_X1 U10547 ( .A(n10408), .B(n10407), .Z(n10656) );
  OR2_X1 U10548 ( .A1(n8023), .A2(n10256), .ZN(n10407) );
  OR2_X1 U10549 ( .A1(n10657), .A2(n10658), .ZN(n10408) );
  AND2_X1 U10550 ( .A1(n10655), .A2(n10654), .ZN(n10658) );
  AND2_X1 U10551 ( .A1(n10652), .A2(n10659), .ZN(n10657) );
  OR2_X1 U10552 ( .A1(n10655), .A2(n10654), .ZN(n10659) );
  OR2_X1 U10553 ( .A1(n10660), .A2(n10661), .ZN(n10654) );
  AND2_X1 U10554 ( .A1(n10651), .A2(n10650), .ZN(n10661) );
  AND2_X1 U10555 ( .A1(n10648), .A2(n10662), .ZN(n10660) );
  OR2_X1 U10556 ( .A1(n10651), .A2(n10650), .ZN(n10662) );
  OR2_X1 U10557 ( .A1(n10663), .A2(n10664), .ZN(n10650) );
  AND2_X1 U10558 ( .A1(n10647), .A2(n10646), .ZN(n10664) );
  AND2_X1 U10559 ( .A1(n10644), .A2(n10665), .ZN(n10663) );
  OR2_X1 U10560 ( .A1(n10647), .A2(n10646), .ZN(n10665) );
  OR2_X1 U10561 ( .A1(n10666), .A2(n10667), .ZN(n10646) );
  AND2_X1 U10562 ( .A1(n10643), .A2(n10642), .ZN(n10667) );
  AND2_X1 U10563 ( .A1(n10640), .A2(n10668), .ZN(n10666) );
  OR2_X1 U10564 ( .A1(n10643), .A2(n10642), .ZN(n10668) );
  OR2_X1 U10565 ( .A1(n10669), .A2(n10670), .ZN(n10642) );
  AND2_X1 U10566 ( .A1(n10639), .A2(n10638), .ZN(n10670) );
  AND2_X1 U10567 ( .A1(n10636), .A2(n10671), .ZN(n10669) );
  OR2_X1 U10568 ( .A1(n10639), .A2(n10638), .ZN(n10671) );
  OR2_X1 U10569 ( .A1(n10672), .A2(n10673), .ZN(n10638) );
  AND2_X1 U10570 ( .A1(n10635), .A2(n10634), .ZN(n10673) );
  AND2_X1 U10571 ( .A1(n10632), .A2(n10674), .ZN(n10672) );
  OR2_X1 U10572 ( .A1(n10635), .A2(n10634), .ZN(n10674) );
  OR2_X1 U10573 ( .A1(n10675), .A2(n10676), .ZN(n10634) );
  AND2_X1 U10574 ( .A1(n10631), .A2(n10630), .ZN(n10676) );
  AND2_X1 U10575 ( .A1(n10628), .A2(n10677), .ZN(n10675) );
  OR2_X1 U10576 ( .A1(n10631), .A2(n10630), .ZN(n10677) );
  OR2_X1 U10577 ( .A1(n10678), .A2(n10679), .ZN(n10630) );
  AND2_X1 U10578 ( .A1(n10627), .A2(n10626), .ZN(n10679) );
  AND2_X1 U10579 ( .A1(n10624), .A2(n10680), .ZN(n10678) );
  OR2_X1 U10580 ( .A1(n10627), .A2(n10626), .ZN(n10680) );
  OR2_X1 U10581 ( .A1(n10681), .A2(n10682), .ZN(n10626) );
  AND2_X1 U10582 ( .A1(n10623), .A2(n10622), .ZN(n10682) );
  AND2_X1 U10583 ( .A1(n10620), .A2(n10683), .ZN(n10681) );
  OR2_X1 U10584 ( .A1(n10623), .A2(n10622), .ZN(n10683) );
  OR2_X1 U10585 ( .A1(n10684), .A2(n10685), .ZN(n10622) );
  AND2_X1 U10586 ( .A1(n10619), .A2(n10618), .ZN(n10685) );
  AND2_X1 U10587 ( .A1(n10616), .A2(n10686), .ZN(n10684) );
  OR2_X1 U10588 ( .A1(n10619), .A2(n10618), .ZN(n10686) );
  OR2_X1 U10589 ( .A1(n10687), .A2(n10688), .ZN(n10618) );
  AND2_X1 U10590 ( .A1(n10615), .A2(n10614), .ZN(n10688) );
  AND2_X1 U10591 ( .A1(n10612), .A2(n10689), .ZN(n10687) );
  OR2_X1 U10592 ( .A1(n10615), .A2(n10614), .ZN(n10689) );
  OR2_X1 U10593 ( .A1(n10690), .A2(n10691), .ZN(n10614) );
  AND2_X1 U10594 ( .A1(n10611), .A2(n10610), .ZN(n10691) );
  AND2_X1 U10595 ( .A1(n10608), .A2(n10692), .ZN(n10690) );
  OR2_X1 U10596 ( .A1(n10611), .A2(n10610), .ZN(n10692) );
  OR2_X1 U10597 ( .A1(n10693), .A2(n10694), .ZN(n10610) );
  AND2_X1 U10598 ( .A1(n10607), .A2(n10606), .ZN(n10694) );
  AND2_X1 U10599 ( .A1(n10604), .A2(n10695), .ZN(n10693) );
  OR2_X1 U10600 ( .A1(n10607), .A2(n10606), .ZN(n10695) );
  OR2_X1 U10601 ( .A1(n10696), .A2(n10697), .ZN(n10606) );
  AND2_X1 U10602 ( .A1(n10603), .A2(n10602), .ZN(n10697) );
  AND2_X1 U10603 ( .A1(n10600), .A2(n10698), .ZN(n10696) );
  OR2_X1 U10604 ( .A1(n10603), .A2(n10602), .ZN(n10698) );
  OR2_X1 U10605 ( .A1(n10699), .A2(n10700), .ZN(n10602) );
  AND2_X1 U10606 ( .A1(n10599), .A2(n10598), .ZN(n10700) );
  AND2_X1 U10607 ( .A1(n10596), .A2(n10701), .ZN(n10699) );
  OR2_X1 U10608 ( .A1(n10599), .A2(n10598), .ZN(n10701) );
  OR2_X1 U10609 ( .A1(n10702), .A2(n10703), .ZN(n10598) );
  AND2_X1 U10610 ( .A1(n10595), .A2(n10594), .ZN(n10703) );
  AND2_X1 U10611 ( .A1(n10592), .A2(n10704), .ZN(n10702) );
  OR2_X1 U10612 ( .A1(n10595), .A2(n10594), .ZN(n10704) );
  OR2_X1 U10613 ( .A1(n10705), .A2(n10706), .ZN(n10594) );
  AND2_X1 U10614 ( .A1(n10591), .A2(n10590), .ZN(n10706) );
  AND2_X1 U10615 ( .A1(n10588), .A2(n10707), .ZN(n10705) );
  OR2_X1 U10616 ( .A1(n10591), .A2(n10590), .ZN(n10707) );
  OR2_X1 U10617 ( .A1(n10708), .A2(n10709), .ZN(n10590) );
  AND2_X1 U10618 ( .A1(n10587), .A2(n10586), .ZN(n10709) );
  AND2_X1 U10619 ( .A1(n10584), .A2(n10710), .ZN(n10708) );
  OR2_X1 U10620 ( .A1(n10587), .A2(n10586), .ZN(n10710) );
  OR2_X1 U10621 ( .A1(n10711), .A2(n10712), .ZN(n10586) );
  AND2_X1 U10622 ( .A1(n10583), .A2(n10582), .ZN(n10712) );
  AND2_X1 U10623 ( .A1(n10580), .A2(n10713), .ZN(n10711) );
  OR2_X1 U10624 ( .A1(n10583), .A2(n10582), .ZN(n10713) );
  OR2_X1 U10625 ( .A1(n10714), .A2(n10715), .ZN(n10582) );
  AND2_X1 U10626 ( .A1(n10579), .A2(n10578), .ZN(n10715) );
  AND2_X1 U10627 ( .A1(n10576), .A2(n10716), .ZN(n10714) );
  OR2_X1 U10628 ( .A1(n10579), .A2(n10578), .ZN(n10716) );
  OR2_X1 U10629 ( .A1(n10717), .A2(n10718), .ZN(n10578) );
  AND2_X1 U10630 ( .A1(n10575), .A2(n10574), .ZN(n10718) );
  AND2_X1 U10631 ( .A1(n10572), .A2(n10719), .ZN(n10717) );
  OR2_X1 U10632 ( .A1(n10575), .A2(n10574), .ZN(n10719) );
  OR2_X1 U10633 ( .A1(n10720), .A2(n10721), .ZN(n10574) );
  AND2_X1 U10634 ( .A1(n10571), .A2(n10570), .ZN(n10721) );
  AND2_X1 U10635 ( .A1(n10568), .A2(n10722), .ZN(n10720) );
  OR2_X1 U10636 ( .A1(n10571), .A2(n10570), .ZN(n10722) );
  OR2_X1 U10637 ( .A1(n10723), .A2(n10724), .ZN(n10570) );
  AND2_X1 U10638 ( .A1(n10567), .A2(n10566), .ZN(n10724) );
  AND2_X1 U10639 ( .A1(n10564), .A2(n10725), .ZN(n10723) );
  OR2_X1 U10640 ( .A1(n10567), .A2(n10566), .ZN(n10725) );
  OR2_X1 U10641 ( .A1(n10726), .A2(n10727), .ZN(n10566) );
  AND2_X1 U10642 ( .A1(n10563), .A2(n10562), .ZN(n10727) );
  AND2_X1 U10643 ( .A1(n10560), .A2(n10728), .ZN(n10726) );
  OR2_X1 U10644 ( .A1(n10563), .A2(n10562), .ZN(n10728) );
  OR2_X1 U10645 ( .A1(n10729), .A2(n10730), .ZN(n10562) );
  AND2_X1 U10646 ( .A1(n10559), .A2(n10558), .ZN(n10730) );
  AND2_X1 U10647 ( .A1(n10556), .A2(n10731), .ZN(n10729) );
  OR2_X1 U10648 ( .A1(n10559), .A2(n10558), .ZN(n10731) );
  OR2_X1 U10649 ( .A1(n10732), .A2(n10733), .ZN(n10558) );
  AND2_X1 U10650 ( .A1(n10555), .A2(n10554), .ZN(n10733) );
  AND2_X1 U10651 ( .A1(n10552), .A2(n10734), .ZN(n10732) );
  OR2_X1 U10652 ( .A1(n10555), .A2(n10554), .ZN(n10734) );
  OR2_X1 U10653 ( .A1(n10735), .A2(n10736), .ZN(n10554) );
  AND2_X1 U10654 ( .A1(n10551), .A2(n10550), .ZN(n10736) );
  AND2_X1 U10655 ( .A1(n10548), .A2(n10737), .ZN(n10735) );
  OR2_X1 U10656 ( .A1(n10551), .A2(n10550), .ZN(n10737) );
  OR2_X1 U10657 ( .A1(n10738), .A2(n10739), .ZN(n10550) );
  AND2_X1 U10658 ( .A1(n10544), .A2(n10547), .ZN(n10739) );
  AND2_X1 U10659 ( .A1(n10546), .A2(n10740), .ZN(n10738) );
  OR2_X1 U10660 ( .A1(n10544), .A2(n10547), .ZN(n10740) );
  OR3_X1 U10661 ( .A1(n10372), .A2(n10256), .A3(n8519), .ZN(n10547) );
  OR2_X1 U10662 ( .A1(n10256), .A2(n7606), .ZN(n10544) );
  INV_X1 U10663 ( .A(n10741), .ZN(n10546) );
  OR2_X1 U10664 ( .A1(n10742), .A2(n10743), .ZN(n10741) );
  AND2_X1 U10665 ( .A1(n10744), .A2(n10745), .ZN(n10743) );
  OR2_X1 U10666 ( .A1(n10746), .A2(n7697), .ZN(n10745) );
  AND2_X1 U10667 ( .A1(n10372), .A2(n7691), .ZN(n10746) );
  AND2_X1 U10668 ( .A1(n10539), .A2(n10747), .ZN(n10742) );
  OR2_X1 U10669 ( .A1(n10748), .A2(n7701), .ZN(n10747) );
  AND2_X1 U10670 ( .A1(n8273), .A2(n7703), .ZN(n10748) );
  OR2_X1 U10671 ( .A1(n7662), .A2(n10256), .ZN(n10551) );
  XNOR2_X1 U10672 ( .A(n10749), .B(n10750), .ZN(n10548) );
  XNOR2_X1 U10673 ( .A(n10751), .B(n10752), .ZN(n10750) );
  OR2_X1 U10674 ( .A1(n7660), .A2(n10256), .ZN(n10555) );
  XOR2_X1 U10675 ( .A(n10753), .B(n10754), .Z(n10552) );
  XOR2_X1 U10676 ( .A(n10755), .B(n10756), .Z(n10754) );
  OR2_X1 U10677 ( .A1(n7658), .A2(n10256), .ZN(n10559) );
  XOR2_X1 U10678 ( .A(n10757), .B(n10758), .Z(n10556) );
  XOR2_X1 U10679 ( .A(n10759), .B(n10760), .Z(n10758) );
  OR2_X1 U10680 ( .A1(n7656), .A2(n10256), .ZN(n10563) );
  XOR2_X1 U10681 ( .A(n10761), .B(n10762), .Z(n10560) );
  XOR2_X1 U10682 ( .A(n10763), .B(n10764), .Z(n10762) );
  OR2_X1 U10683 ( .A1(n7654), .A2(n10256), .ZN(n10567) );
  XOR2_X1 U10684 ( .A(n10765), .B(n10766), .Z(n10564) );
  XOR2_X1 U10685 ( .A(n10767), .B(n10768), .Z(n10766) );
  OR2_X1 U10686 ( .A1(n7652), .A2(n10256), .ZN(n10571) );
  XOR2_X1 U10687 ( .A(n10769), .B(n10770), .Z(n10568) );
  XOR2_X1 U10688 ( .A(n10771), .B(n10772), .Z(n10770) );
  OR2_X1 U10689 ( .A1(n7650), .A2(n10256), .ZN(n10575) );
  XOR2_X1 U10690 ( .A(n10773), .B(n10774), .Z(n10572) );
  XOR2_X1 U10691 ( .A(n10775), .B(n10776), .Z(n10774) );
  OR2_X1 U10692 ( .A1(n7648), .A2(n10256), .ZN(n10579) );
  XOR2_X1 U10693 ( .A(n10777), .B(n10778), .Z(n10576) );
  XOR2_X1 U10694 ( .A(n10779), .B(n10780), .Z(n10778) );
  OR2_X1 U10695 ( .A1(n7646), .A2(n10256), .ZN(n10583) );
  XOR2_X1 U10696 ( .A(n10781), .B(n10782), .Z(n10580) );
  XOR2_X1 U10697 ( .A(n10783), .B(n10784), .Z(n10782) );
  OR2_X1 U10698 ( .A1(n7644), .A2(n10256), .ZN(n10587) );
  XOR2_X1 U10699 ( .A(n10785), .B(n10786), .Z(n10584) );
  XOR2_X1 U10700 ( .A(n10787), .B(n10788), .Z(n10786) );
  OR2_X1 U10701 ( .A1(n7642), .A2(n10256), .ZN(n10591) );
  XOR2_X1 U10702 ( .A(n10789), .B(n10790), .Z(n10588) );
  XOR2_X1 U10703 ( .A(n10791), .B(n10792), .Z(n10790) );
  OR2_X1 U10704 ( .A1(n7640), .A2(n10256), .ZN(n10595) );
  XOR2_X1 U10705 ( .A(n10793), .B(n10794), .Z(n10592) );
  XOR2_X1 U10706 ( .A(n10795), .B(n10796), .Z(n10794) );
  OR2_X1 U10707 ( .A1(n7638), .A2(n10256), .ZN(n10599) );
  XOR2_X1 U10708 ( .A(n10797), .B(n10798), .Z(n10596) );
  XOR2_X1 U10709 ( .A(n10799), .B(n10800), .Z(n10798) );
  OR2_X1 U10710 ( .A1(n7636), .A2(n10256), .ZN(n10603) );
  XOR2_X1 U10711 ( .A(n10801), .B(n10802), .Z(n10600) );
  XOR2_X1 U10712 ( .A(n10803), .B(n10804), .Z(n10802) );
  OR2_X1 U10713 ( .A1(n7634), .A2(n10256), .ZN(n10607) );
  XOR2_X1 U10714 ( .A(n10805), .B(n10806), .Z(n10604) );
  XOR2_X1 U10715 ( .A(n10807), .B(n10808), .Z(n10806) );
  OR2_X1 U10716 ( .A1(n7632), .A2(n10256), .ZN(n10611) );
  XOR2_X1 U10717 ( .A(n10809), .B(n10810), .Z(n10608) );
  XOR2_X1 U10718 ( .A(n10811), .B(n10812), .Z(n10810) );
  OR2_X1 U10719 ( .A1(n7630), .A2(n10256), .ZN(n10615) );
  XOR2_X1 U10720 ( .A(n10813), .B(n10814), .Z(n10612) );
  XOR2_X1 U10721 ( .A(n10815), .B(n10816), .Z(n10814) );
  OR2_X1 U10722 ( .A1(n7628), .A2(n10256), .ZN(n10619) );
  XOR2_X1 U10723 ( .A(n10817), .B(n10818), .Z(n10616) );
  XOR2_X1 U10724 ( .A(n10819), .B(n10820), .Z(n10818) );
  OR2_X1 U10725 ( .A1(n7626), .A2(n10256), .ZN(n10623) );
  XOR2_X1 U10726 ( .A(n10821), .B(n10822), .Z(n10620) );
  XOR2_X1 U10727 ( .A(n10823), .B(n10824), .Z(n10822) );
  OR2_X1 U10728 ( .A1(n7624), .A2(n10256), .ZN(n10627) );
  XOR2_X1 U10729 ( .A(n10825), .B(n10826), .Z(n10624) );
  XOR2_X1 U10730 ( .A(n10827), .B(n10828), .Z(n10826) );
  OR2_X1 U10731 ( .A1(n7622), .A2(n10256), .ZN(n10631) );
  XOR2_X1 U10732 ( .A(n10829), .B(n10830), .Z(n10628) );
  XOR2_X1 U10733 ( .A(n10831), .B(n10832), .Z(n10830) );
  OR2_X1 U10734 ( .A1(n8634), .A2(n10256), .ZN(n10635) );
  XOR2_X1 U10735 ( .A(n10833), .B(n10834), .Z(n10632) );
  XOR2_X1 U10736 ( .A(n10835), .B(n10836), .Z(n10834) );
  OR2_X1 U10737 ( .A1(n8639), .A2(n10256), .ZN(n10639) );
  XOR2_X1 U10738 ( .A(n10837), .B(n10838), .Z(n10636) );
  XOR2_X1 U10739 ( .A(n10839), .B(n10840), .Z(n10838) );
  OR2_X1 U10740 ( .A1(n8644), .A2(n10256), .ZN(n10643) );
  XOR2_X1 U10741 ( .A(n10841), .B(n10842), .Z(n10640) );
  XOR2_X1 U10742 ( .A(n10843), .B(n10844), .Z(n10842) );
  OR2_X1 U10743 ( .A1(n8152), .A2(n10256), .ZN(n10647) );
  XOR2_X1 U10744 ( .A(n10845), .B(n10846), .Z(n10644) );
  XOR2_X1 U10745 ( .A(n10847), .B(n10848), .Z(n10846) );
  OR2_X1 U10746 ( .A1(n8105), .A2(n10256), .ZN(n10651) );
  XOR2_X1 U10747 ( .A(n10849), .B(n10850), .Z(n10648) );
  XOR2_X1 U10748 ( .A(n10851), .B(n10852), .Z(n10850) );
  OR2_X1 U10749 ( .A1(n8056), .A2(n10256), .ZN(n10655) );
  INV_X1 U10750 ( .A(n10251), .ZN(n10256) );
  XOR2_X1 U10751 ( .A(n10853), .B(n10854), .Z(n10251) );
  XNOR2_X1 U10752 ( .A(c_21_), .B(d_21_), .ZN(n10853) );
  XOR2_X1 U10753 ( .A(n10855), .B(n10856), .Z(n10652) );
  XOR2_X1 U10754 ( .A(n10857), .B(n10858), .Z(n10856) );
  XOR2_X1 U10755 ( .A(n10416), .B(n10859), .Z(n10409) );
  XOR2_X1 U10756 ( .A(n10415), .B(n10414), .Z(n10859) );
  OR2_X1 U10757 ( .A1(n8056), .A2(n10372), .ZN(n10414) );
  OR2_X1 U10758 ( .A1(n10860), .A2(n10861), .ZN(n10415) );
  AND2_X1 U10759 ( .A1(n10858), .A2(n10857), .ZN(n10861) );
  AND2_X1 U10760 ( .A1(n10855), .A2(n10862), .ZN(n10860) );
  OR2_X1 U10761 ( .A1(n10858), .A2(n10857), .ZN(n10862) );
  OR2_X1 U10762 ( .A1(n10863), .A2(n10864), .ZN(n10857) );
  AND2_X1 U10763 ( .A1(n10852), .A2(n10851), .ZN(n10864) );
  AND2_X1 U10764 ( .A1(n10849), .A2(n10865), .ZN(n10863) );
  OR2_X1 U10765 ( .A1(n10852), .A2(n10851), .ZN(n10865) );
  OR2_X1 U10766 ( .A1(n10866), .A2(n10867), .ZN(n10851) );
  AND2_X1 U10767 ( .A1(n10848), .A2(n10847), .ZN(n10867) );
  AND2_X1 U10768 ( .A1(n10845), .A2(n10868), .ZN(n10866) );
  OR2_X1 U10769 ( .A1(n10848), .A2(n10847), .ZN(n10868) );
  OR2_X1 U10770 ( .A1(n10869), .A2(n10870), .ZN(n10847) );
  AND2_X1 U10771 ( .A1(n10844), .A2(n10843), .ZN(n10870) );
  AND2_X1 U10772 ( .A1(n10841), .A2(n10871), .ZN(n10869) );
  OR2_X1 U10773 ( .A1(n10844), .A2(n10843), .ZN(n10871) );
  OR2_X1 U10774 ( .A1(n10872), .A2(n10873), .ZN(n10843) );
  AND2_X1 U10775 ( .A1(n10840), .A2(n10839), .ZN(n10873) );
  AND2_X1 U10776 ( .A1(n10837), .A2(n10874), .ZN(n10872) );
  OR2_X1 U10777 ( .A1(n10840), .A2(n10839), .ZN(n10874) );
  OR2_X1 U10778 ( .A1(n10875), .A2(n10876), .ZN(n10839) );
  AND2_X1 U10779 ( .A1(n10836), .A2(n10835), .ZN(n10876) );
  AND2_X1 U10780 ( .A1(n10833), .A2(n10877), .ZN(n10875) );
  OR2_X1 U10781 ( .A1(n10836), .A2(n10835), .ZN(n10877) );
  OR2_X1 U10782 ( .A1(n10878), .A2(n10879), .ZN(n10835) );
  AND2_X1 U10783 ( .A1(n10832), .A2(n10831), .ZN(n10879) );
  AND2_X1 U10784 ( .A1(n10829), .A2(n10880), .ZN(n10878) );
  OR2_X1 U10785 ( .A1(n10832), .A2(n10831), .ZN(n10880) );
  OR2_X1 U10786 ( .A1(n10881), .A2(n10882), .ZN(n10831) );
  AND2_X1 U10787 ( .A1(n10828), .A2(n10827), .ZN(n10882) );
  AND2_X1 U10788 ( .A1(n10825), .A2(n10883), .ZN(n10881) );
  OR2_X1 U10789 ( .A1(n10828), .A2(n10827), .ZN(n10883) );
  OR2_X1 U10790 ( .A1(n10884), .A2(n10885), .ZN(n10827) );
  AND2_X1 U10791 ( .A1(n10824), .A2(n10823), .ZN(n10885) );
  AND2_X1 U10792 ( .A1(n10821), .A2(n10886), .ZN(n10884) );
  OR2_X1 U10793 ( .A1(n10824), .A2(n10823), .ZN(n10886) );
  OR2_X1 U10794 ( .A1(n10887), .A2(n10888), .ZN(n10823) );
  AND2_X1 U10795 ( .A1(n10820), .A2(n10819), .ZN(n10888) );
  AND2_X1 U10796 ( .A1(n10817), .A2(n10889), .ZN(n10887) );
  OR2_X1 U10797 ( .A1(n10820), .A2(n10819), .ZN(n10889) );
  OR2_X1 U10798 ( .A1(n10890), .A2(n10891), .ZN(n10819) );
  AND2_X1 U10799 ( .A1(n10816), .A2(n10815), .ZN(n10891) );
  AND2_X1 U10800 ( .A1(n10813), .A2(n10892), .ZN(n10890) );
  OR2_X1 U10801 ( .A1(n10816), .A2(n10815), .ZN(n10892) );
  OR2_X1 U10802 ( .A1(n10893), .A2(n10894), .ZN(n10815) );
  AND2_X1 U10803 ( .A1(n10812), .A2(n10811), .ZN(n10894) );
  AND2_X1 U10804 ( .A1(n10809), .A2(n10895), .ZN(n10893) );
  OR2_X1 U10805 ( .A1(n10812), .A2(n10811), .ZN(n10895) );
  OR2_X1 U10806 ( .A1(n10896), .A2(n10897), .ZN(n10811) );
  AND2_X1 U10807 ( .A1(n10808), .A2(n10807), .ZN(n10897) );
  AND2_X1 U10808 ( .A1(n10805), .A2(n10898), .ZN(n10896) );
  OR2_X1 U10809 ( .A1(n10808), .A2(n10807), .ZN(n10898) );
  OR2_X1 U10810 ( .A1(n10899), .A2(n10900), .ZN(n10807) );
  AND2_X1 U10811 ( .A1(n10804), .A2(n10803), .ZN(n10900) );
  AND2_X1 U10812 ( .A1(n10801), .A2(n10901), .ZN(n10899) );
  OR2_X1 U10813 ( .A1(n10804), .A2(n10803), .ZN(n10901) );
  OR2_X1 U10814 ( .A1(n10902), .A2(n10903), .ZN(n10803) );
  AND2_X1 U10815 ( .A1(n10800), .A2(n10799), .ZN(n10903) );
  AND2_X1 U10816 ( .A1(n10797), .A2(n10904), .ZN(n10902) );
  OR2_X1 U10817 ( .A1(n10800), .A2(n10799), .ZN(n10904) );
  OR2_X1 U10818 ( .A1(n10905), .A2(n10906), .ZN(n10799) );
  AND2_X1 U10819 ( .A1(n10796), .A2(n10795), .ZN(n10906) );
  AND2_X1 U10820 ( .A1(n10793), .A2(n10907), .ZN(n10905) );
  OR2_X1 U10821 ( .A1(n10796), .A2(n10795), .ZN(n10907) );
  OR2_X1 U10822 ( .A1(n10908), .A2(n10909), .ZN(n10795) );
  AND2_X1 U10823 ( .A1(n10792), .A2(n10791), .ZN(n10909) );
  AND2_X1 U10824 ( .A1(n10789), .A2(n10910), .ZN(n10908) );
  OR2_X1 U10825 ( .A1(n10792), .A2(n10791), .ZN(n10910) );
  OR2_X1 U10826 ( .A1(n10911), .A2(n10912), .ZN(n10791) );
  AND2_X1 U10827 ( .A1(n10788), .A2(n10787), .ZN(n10912) );
  AND2_X1 U10828 ( .A1(n10785), .A2(n10913), .ZN(n10911) );
  OR2_X1 U10829 ( .A1(n10788), .A2(n10787), .ZN(n10913) );
  OR2_X1 U10830 ( .A1(n10914), .A2(n10915), .ZN(n10787) );
  AND2_X1 U10831 ( .A1(n10784), .A2(n10783), .ZN(n10915) );
  AND2_X1 U10832 ( .A1(n10781), .A2(n10916), .ZN(n10914) );
  OR2_X1 U10833 ( .A1(n10784), .A2(n10783), .ZN(n10916) );
  OR2_X1 U10834 ( .A1(n10917), .A2(n10918), .ZN(n10783) );
  AND2_X1 U10835 ( .A1(n10780), .A2(n10779), .ZN(n10918) );
  AND2_X1 U10836 ( .A1(n10777), .A2(n10919), .ZN(n10917) );
  OR2_X1 U10837 ( .A1(n10780), .A2(n10779), .ZN(n10919) );
  OR2_X1 U10838 ( .A1(n10920), .A2(n10921), .ZN(n10779) );
  AND2_X1 U10839 ( .A1(n10776), .A2(n10775), .ZN(n10921) );
  AND2_X1 U10840 ( .A1(n10773), .A2(n10922), .ZN(n10920) );
  OR2_X1 U10841 ( .A1(n10776), .A2(n10775), .ZN(n10922) );
  OR2_X1 U10842 ( .A1(n10923), .A2(n10924), .ZN(n10775) );
  AND2_X1 U10843 ( .A1(n10772), .A2(n10771), .ZN(n10924) );
  AND2_X1 U10844 ( .A1(n10769), .A2(n10925), .ZN(n10923) );
  OR2_X1 U10845 ( .A1(n10772), .A2(n10771), .ZN(n10925) );
  OR2_X1 U10846 ( .A1(n10926), .A2(n10927), .ZN(n10771) );
  AND2_X1 U10847 ( .A1(n10768), .A2(n10767), .ZN(n10927) );
  AND2_X1 U10848 ( .A1(n10765), .A2(n10928), .ZN(n10926) );
  OR2_X1 U10849 ( .A1(n10768), .A2(n10767), .ZN(n10928) );
  OR2_X1 U10850 ( .A1(n10929), .A2(n10930), .ZN(n10767) );
  AND2_X1 U10851 ( .A1(n10764), .A2(n10763), .ZN(n10930) );
  AND2_X1 U10852 ( .A1(n10761), .A2(n10931), .ZN(n10929) );
  OR2_X1 U10853 ( .A1(n10764), .A2(n10763), .ZN(n10931) );
  OR2_X1 U10854 ( .A1(n10932), .A2(n10933), .ZN(n10763) );
  AND2_X1 U10855 ( .A1(n10760), .A2(n10759), .ZN(n10933) );
  AND2_X1 U10856 ( .A1(n10757), .A2(n10934), .ZN(n10932) );
  OR2_X1 U10857 ( .A1(n10760), .A2(n10759), .ZN(n10934) );
  OR2_X1 U10858 ( .A1(n10935), .A2(n10936), .ZN(n10759) );
  AND2_X1 U10859 ( .A1(n10756), .A2(n10755), .ZN(n10936) );
  AND2_X1 U10860 ( .A1(n10753), .A2(n10937), .ZN(n10935) );
  OR2_X1 U10861 ( .A1(n10756), .A2(n10755), .ZN(n10937) );
  OR2_X1 U10862 ( .A1(n10938), .A2(n10939), .ZN(n10755) );
  AND2_X1 U10863 ( .A1(n10749), .A2(n10752), .ZN(n10939) );
  AND2_X1 U10864 ( .A1(n10751), .A2(n10940), .ZN(n10938) );
  OR2_X1 U10865 ( .A1(n10749), .A2(n10752), .ZN(n10940) );
  OR3_X1 U10866 ( .A1(n8273), .A2(n10372), .A3(n8519), .ZN(n10752) );
  OR2_X1 U10867 ( .A1(n10372), .A2(n7606), .ZN(n10749) );
  INV_X1 U10868 ( .A(n10941), .ZN(n10751) );
  OR2_X1 U10869 ( .A1(n10942), .A2(n10943), .ZN(n10941) );
  AND2_X1 U10870 ( .A1(n10944), .A2(n10945), .ZN(n10943) );
  OR2_X1 U10871 ( .A1(n10946), .A2(n7697), .ZN(n10945) );
  AND2_X1 U10872 ( .A1(n8273), .A2(n7691), .ZN(n10946) );
  AND2_X1 U10873 ( .A1(n10744), .A2(n10947), .ZN(n10942) );
  OR2_X1 U10874 ( .A1(n10948), .A2(n7701), .ZN(n10947) );
  AND2_X1 U10875 ( .A1(n8243), .A2(n7703), .ZN(n10948) );
  OR2_X1 U10876 ( .A1(n7662), .A2(n10372), .ZN(n10756) );
  XNOR2_X1 U10877 ( .A(n10949), .B(n10950), .ZN(n10753) );
  XNOR2_X1 U10878 ( .A(n10951), .B(n10952), .ZN(n10950) );
  OR2_X1 U10879 ( .A1(n7660), .A2(n10372), .ZN(n10760) );
  XOR2_X1 U10880 ( .A(n10953), .B(n10954), .Z(n10757) );
  XOR2_X1 U10881 ( .A(n10955), .B(n10956), .Z(n10954) );
  OR2_X1 U10882 ( .A1(n7658), .A2(n10372), .ZN(n10764) );
  XOR2_X1 U10883 ( .A(n10957), .B(n10958), .Z(n10761) );
  XOR2_X1 U10884 ( .A(n10959), .B(n10960), .Z(n10958) );
  OR2_X1 U10885 ( .A1(n7656), .A2(n10372), .ZN(n10768) );
  XOR2_X1 U10886 ( .A(n10961), .B(n10962), .Z(n10765) );
  XOR2_X1 U10887 ( .A(n10963), .B(n10964), .Z(n10962) );
  OR2_X1 U10888 ( .A1(n7654), .A2(n10372), .ZN(n10772) );
  XOR2_X1 U10889 ( .A(n10965), .B(n10966), .Z(n10769) );
  XOR2_X1 U10890 ( .A(n10967), .B(n10968), .Z(n10966) );
  OR2_X1 U10891 ( .A1(n7652), .A2(n10372), .ZN(n10776) );
  XOR2_X1 U10892 ( .A(n10969), .B(n10970), .Z(n10773) );
  XOR2_X1 U10893 ( .A(n10971), .B(n10972), .Z(n10970) );
  OR2_X1 U10894 ( .A1(n7650), .A2(n10372), .ZN(n10780) );
  XOR2_X1 U10895 ( .A(n10973), .B(n10974), .Z(n10777) );
  XOR2_X1 U10896 ( .A(n10975), .B(n10976), .Z(n10974) );
  OR2_X1 U10897 ( .A1(n7648), .A2(n10372), .ZN(n10784) );
  XOR2_X1 U10898 ( .A(n10977), .B(n10978), .Z(n10781) );
  XOR2_X1 U10899 ( .A(n10979), .B(n10980), .Z(n10978) );
  OR2_X1 U10900 ( .A1(n7646), .A2(n10372), .ZN(n10788) );
  XOR2_X1 U10901 ( .A(n10981), .B(n10982), .Z(n10785) );
  XOR2_X1 U10902 ( .A(n10983), .B(n10984), .Z(n10982) );
  OR2_X1 U10903 ( .A1(n7644), .A2(n10372), .ZN(n10792) );
  XOR2_X1 U10904 ( .A(n10985), .B(n10986), .Z(n10789) );
  XOR2_X1 U10905 ( .A(n10987), .B(n10988), .Z(n10986) );
  OR2_X1 U10906 ( .A1(n7642), .A2(n10372), .ZN(n10796) );
  XOR2_X1 U10907 ( .A(n10989), .B(n10990), .Z(n10793) );
  XOR2_X1 U10908 ( .A(n10991), .B(n10992), .Z(n10990) );
  OR2_X1 U10909 ( .A1(n7640), .A2(n10372), .ZN(n10800) );
  XOR2_X1 U10910 ( .A(n10993), .B(n10994), .Z(n10797) );
  XOR2_X1 U10911 ( .A(n10995), .B(n10996), .Z(n10994) );
  OR2_X1 U10912 ( .A1(n7638), .A2(n10372), .ZN(n10804) );
  XOR2_X1 U10913 ( .A(n10997), .B(n10998), .Z(n10801) );
  XOR2_X1 U10914 ( .A(n10999), .B(n11000), .Z(n10998) );
  OR2_X1 U10915 ( .A1(n7636), .A2(n10372), .ZN(n10808) );
  XOR2_X1 U10916 ( .A(n11001), .B(n11002), .Z(n10805) );
  XOR2_X1 U10917 ( .A(n11003), .B(n11004), .Z(n11002) );
  OR2_X1 U10918 ( .A1(n7634), .A2(n10372), .ZN(n10812) );
  XOR2_X1 U10919 ( .A(n11005), .B(n11006), .Z(n10809) );
  XOR2_X1 U10920 ( .A(n11007), .B(n11008), .Z(n11006) );
  OR2_X1 U10921 ( .A1(n7632), .A2(n10372), .ZN(n10816) );
  XOR2_X1 U10922 ( .A(n11009), .B(n11010), .Z(n10813) );
  XOR2_X1 U10923 ( .A(n11011), .B(n11012), .Z(n11010) );
  OR2_X1 U10924 ( .A1(n7630), .A2(n10372), .ZN(n10820) );
  XOR2_X1 U10925 ( .A(n11013), .B(n11014), .Z(n10817) );
  XOR2_X1 U10926 ( .A(n11015), .B(n11016), .Z(n11014) );
  OR2_X1 U10927 ( .A1(n7628), .A2(n10372), .ZN(n10824) );
  XOR2_X1 U10928 ( .A(n11017), .B(n11018), .Z(n10821) );
  XOR2_X1 U10929 ( .A(n11019), .B(n11020), .Z(n11018) );
  OR2_X1 U10930 ( .A1(n7626), .A2(n10372), .ZN(n10828) );
  XOR2_X1 U10931 ( .A(n11021), .B(n11022), .Z(n10825) );
  XOR2_X1 U10932 ( .A(n11023), .B(n11024), .Z(n11022) );
  OR2_X1 U10933 ( .A1(n7624), .A2(n10372), .ZN(n10832) );
  XOR2_X1 U10934 ( .A(n11025), .B(n11026), .Z(n10829) );
  XOR2_X1 U10935 ( .A(n11027), .B(n11028), .Z(n11026) );
  OR2_X1 U10936 ( .A1(n8629), .A2(n10372), .ZN(n10836) );
  XOR2_X1 U10937 ( .A(n11029), .B(n11030), .Z(n10833) );
  XOR2_X1 U10938 ( .A(n11031), .B(n11032), .Z(n11030) );
  OR2_X1 U10939 ( .A1(n8634), .A2(n10372), .ZN(n10840) );
  XOR2_X1 U10940 ( .A(n11033), .B(n11034), .Z(n10837) );
  XOR2_X1 U10941 ( .A(n11035), .B(n11036), .Z(n11034) );
  OR2_X1 U10942 ( .A1(n8639), .A2(n10372), .ZN(n10844) );
  XOR2_X1 U10943 ( .A(n11037), .B(n11038), .Z(n10841) );
  XOR2_X1 U10944 ( .A(n11039), .B(n11040), .Z(n11038) );
  OR2_X1 U10945 ( .A1(n8644), .A2(n10372), .ZN(n10848) );
  XOR2_X1 U10946 ( .A(n11041), .B(n11042), .Z(n10845) );
  XOR2_X1 U10947 ( .A(n11043), .B(n11044), .Z(n11042) );
  OR2_X1 U10948 ( .A1(n8152), .A2(n10372), .ZN(n10852) );
  XOR2_X1 U10949 ( .A(n11045), .B(n11046), .Z(n10849) );
  XOR2_X1 U10950 ( .A(n11047), .B(n11048), .Z(n11046) );
  OR2_X1 U10951 ( .A1(n8105), .A2(n10372), .ZN(n10858) );
  INV_X1 U10952 ( .A(n10539), .ZN(n10372) );
  XOR2_X1 U10953 ( .A(n11049), .B(n11050), .Z(n10539) );
  XNOR2_X1 U10954 ( .A(c_20_), .B(d_20_), .ZN(n11049) );
  XOR2_X1 U10955 ( .A(n11051), .B(n11052), .Z(n10855) );
  XOR2_X1 U10956 ( .A(n11053), .B(n11054), .Z(n11052) );
  XOR2_X1 U10957 ( .A(n10423), .B(n11055), .Z(n10416) );
  XOR2_X1 U10958 ( .A(n10422), .B(n10421), .Z(n11055) );
  OR2_X1 U10959 ( .A1(n8105), .A2(n8273), .ZN(n10421) );
  OR2_X1 U10960 ( .A1(n11056), .A2(n11057), .ZN(n10422) );
  AND2_X1 U10961 ( .A1(n11054), .A2(n11053), .ZN(n11057) );
  AND2_X1 U10962 ( .A1(n11051), .A2(n11058), .ZN(n11056) );
  OR2_X1 U10963 ( .A1(n11054), .A2(n11053), .ZN(n11058) );
  OR2_X1 U10964 ( .A1(n11059), .A2(n11060), .ZN(n11053) );
  AND2_X1 U10965 ( .A1(n11048), .A2(n11047), .ZN(n11060) );
  AND2_X1 U10966 ( .A1(n11045), .A2(n11061), .ZN(n11059) );
  OR2_X1 U10967 ( .A1(n11048), .A2(n11047), .ZN(n11061) );
  OR2_X1 U10968 ( .A1(n11062), .A2(n11063), .ZN(n11047) );
  AND2_X1 U10969 ( .A1(n11044), .A2(n11043), .ZN(n11063) );
  AND2_X1 U10970 ( .A1(n11041), .A2(n11064), .ZN(n11062) );
  OR2_X1 U10971 ( .A1(n11044), .A2(n11043), .ZN(n11064) );
  OR2_X1 U10972 ( .A1(n11065), .A2(n11066), .ZN(n11043) );
  AND2_X1 U10973 ( .A1(n11040), .A2(n11039), .ZN(n11066) );
  AND2_X1 U10974 ( .A1(n11037), .A2(n11067), .ZN(n11065) );
  OR2_X1 U10975 ( .A1(n11040), .A2(n11039), .ZN(n11067) );
  OR2_X1 U10976 ( .A1(n11068), .A2(n11069), .ZN(n11039) );
  AND2_X1 U10977 ( .A1(n11036), .A2(n11035), .ZN(n11069) );
  AND2_X1 U10978 ( .A1(n11033), .A2(n11070), .ZN(n11068) );
  OR2_X1 U10979 ( .A1(n11036), .A2(n11035), .ZN(n11070) );
  OR2_X1 U10980 ( .A1(n11071), .A2(n11072), .ZN(n11035) );
  AND2_X1 U10981 ( .A1(n11032), .A2(n11031), .ZN(n11072) );
  AND2_X1 U10982 ( .A1(n11029), .A2(n11073), .ZN(n11071) );
  OR2_X1 U10983 ( .A1(n11032), .A2(n11031), .ZN(n11073) );
  OR2_X1 U10984 ( .A1(n11074), .A2(n11075), .ZN(n11031) );
  AND2_X1 U10985 ( .A1(n11028), .A2(n11027), .ZN(n11075) );
  AND2_X1 U10986 ( .A1(n11025), .A2(n11076), .ZN(n11074) );
  OR2_X1 U10987 ( .A1(n11028), .A2(n11027), .ZN(n11076) );
  OR2_X1 U10988 ( .A1(n11077), .A2(n11078), .ZN(n11027) );
  AND2_X1 U10989 ( .A1(n11024), .A2(n11023), .ZN(n11078) );
  AND2_X1 U10990 ( .A1(n11021), .A2(n11079), .ZN(n11077) );
  OR2_X1 U10991 ( .A1(n11024), .A2(n11023), .ZN(n11079) );
  OR2_X1 U10992 ( .A1(n11080), .A2(n11081), .ZN(n11023) );
  AND2_X1 U10993 ( .A1(n11020), .A2(n11019), .ZN(n11081) );
  AND2_X1 U10994 ( .A1(n11017), .A2(n11082), .ZN(n11080) );
  OR2_X1 U10995 ( .A1(n11020), .A2(n11019), .ZN(n11082) );
  OR2_X1 U10996 ( .A1(n11083), .A2(n11084), .ZN(n11019) );
  AND2_X1 U10997 ( .A1(n11016), .A2(n11015), .ZN(n11084) );
  AND2_X1 U10998 ( .A1(n11013), .A2(n11085), .ZN(n11083) );
  OR2_X1 U10999 ( .A1(n11016), .A2(n11015), .ZN(n11085) );
  OR2_X1 U11000 ( .A1(n11086), .A2(n11087), .ZN(n11015) );
  AND2_X1 U11001 ( .A1(n11012), .A2(n11011), .ZN(n11087) );
  AND2_X1 U11002 ( .A1(n11009), .A2(n11088), .ZN(n11086) );
  OR2_X1 U11003 ( .A1(n11012), .A2(n11011), .ZN(n11088) );
  OR2_X1 U11004 ( .A1(n11089), .A2(n11090), .ZN(n11011) );
  AND2_X1 U11005 ( .A1(n11008), .A2(n11007), .ZN(n11090) );
  AND2_X1 U11006 ( .A1(n11005), .A2(n11091), .ZN(n11089) );
  OR2_X1 U11007 ( .A1(n11008), .A2(n11007), .ZN(n11091) );
  OR2_X1 U11008 ( .A1(n11092), .A2(n11093), .ZN(n11007) );
  AND2_X1 U11009 ( .A1(n11004), .A2(n11003), .ZN(n11093) );
  AND2_X1 U11010 ( .A1(n11001), .A2(n11094), .ZN(n11092) );
  OR2_X1 U11011 ( .A1(n11004), .A2(n11003), .ZN(n11094) );
  OR2_X1 U11012 ( .A1(n11095), .A2(n11096), .ZN(n11003) );
  AND2_X1 U11013 ( .A1(n11000), .A2(n10999), .ZN(n11096) );
  AND2_X1 U11014 ( .A1(n10997), .A2(n11097), .ZN(n11095) );
  OR2_X1 U11015 ( .A1(n11000), .A2(n10999), .ZN(n11097) );
  OR2_X1 U11016 ( .A1(n11098), .A2(n11099), .ZN(n10999) );
  AND2_X1 U11017 ( .A1(n10996), .A2(n10995), .ZN(n11099) );
  AND2_X1 U11018 ( .A1(n10993), .A2(n11100), .ZN(n11098) );
  OR2_X1 U11019 ( .A1(n10996), .A2(n10995), .ZN(n11100) );
  OR2_X1 U11020 ( .A1(n11101), .A2(n11102), .ZN(n10995) );
  AND2_X1 U11021 ( .A1(n10992), .A2(n10991), .ZN(n11102) );
  AND2_X1 U11022 ( .A1(n10989), .A2(n11103), .ZN(n11101) );
  OR2_X1 U11023 ( .A1(n10992), .A2(n10991), .ZN(n11103) );
  OR2_X1 U11024 ( .A1(n11104), .A2(n11105), .ZN(n10991) );
  AND2_X1 U11025 ( .A1(n10988), .A2(n10987), .ZN(n11105) );
  AND2_X1 U11026 ( .A1(n10985), .A2(n11106), .ZN(n11104) );
  OR2_X1 U11027 ( .A1(n10988), .A2(n10987), .ZN(n11106) );
  OR2_X1 U11028 ( .A1(n11107), .A2(n11108), .ZN(n10987) );
  AND2_X1 U11029 ( .A1(n10984), .A2(n10983), .ZN(n11108) );
  AND2_X1 U11030 ( .A1(n10981), .A2(n11109), .ZN(n11107) );
  OR2_X1 U11031 ( .A1(n10984), .A2(n10983), .ZN(n11109) );
  OR2_X1 U11032 ( .A1(n11110), .A2(n11111), .ZN(n10983) );
  AND2_X1 U11033 ( .A1(n10980), .A2(n10979), .ZN(n11111) );
  AND2_X1 U11034 ( .A1(n10977), .A2(n11112), .ZN(n11110) );
  OR2_X1 U11035 ( .A1(n10980), .A2(n10979), .ZN(n11112) );
  OR2_X1 U11036 ( .A1(n11113), .A2(n11114), .ZN(n10979) );
  AND2_X1 U11037 ( .A1(n10976), .A2(n10975), .ZN(n11114) );
  AND2_X1 U11038 ( .A1(n10973), .A2(n11115), .ZN(n11113) );
  OR2_X1 U11039 ( .A1(n10976), .A2(n10975), .ZN(n11115) );
  OR2_X1 U11040 ( .A1(n11116), .A2(n11117), .ZN(n10975) );
  AND2_X1 U11041 ( .A1(n10972), .A2(n10971), .ZN(n11117) );
  AND2_X1 U11042 ( .A1(n10969), .A2(n11118), .ZN(n11116) );
  OR2_X1 U11043 ( .A1(n10972), .A2(n10971), .ZN(n11118) );
  OR2_X1 U11044 ( .A1(n11119), .A2(n11120), .ZN(n10971) );
  AND2_X1 U11045 ( .A1(n10968), .A2(n10967), .ZN(n11120) );
  AND2_X1 U11046 ( .A1(n10965), .A2(n11121), .ZN(n11119) );
  OR2_X1 U11047 ( .A1(n10968), .A2(n10967), .ZN(n11121) );
  OR2_X1 U11048 ( .A1(n11122), .A2(n11123), .ZN(n10967) );
  AND2_X1 U11049 ( .A1(n10964), .A2(n10963), .ZN(n11123) );
  AND2_X1 U11050 ( .A1(n10961), .A2(n11124), .ZN(n11122) );
  OR2_X1 U11051 ( .A1(n10964), .A2(n10963), .ZN(n11124) );
  OR2_X1 U11052 ( .A1(n11125), .A2(n11126), .ZN(n10963) );
  AND2_X1 U11053 ( .A1(n10960), .A2(n10959), .ZN(n11126) );
  AND2_X1 U11054 ( .A1(n10957), .A2(n11127), .ZN(n11125) );
  OR2_X1 U11055 ( .A1(n10960), .A2(n10959), .ZN(n11127) );
  OR2_X1 U11056 ( .A1(n11128), .A2(n11129), .ZN(n10959) );
  AND2_X1 U11057 ( .A1(n10956), .A2(n10955), .ZN(n11129) );
  AND2_X1 U11058 ( .A1(n10953), .A2(n11130), .ZN(n11128) );
  OR2_X1 U11059 ( .A1(n10956), .A2(n10955), .ZN(n11130) );
  OR2_X1 U11060 ( .A1(n11131), .A2(n11132), .ZN(n10955) );
  AND2_X1 U11061 ( .A1(n10949), .A2(n10952), .ZN(n11132) );
  AND2_X1 U11062 ( .A1(n10951), .A2(n11133), .ZN(n11131) );
  OR2_X1 U11063 ( .A1(n10949), .A2(n10952), .ZN(n11133) );
  OR3_X1 U11064 ( .A1(n8243), .A2(n8273), .A3(n8519), .ZN(n10952) );
  OR2_X1 U11065 ( .A1(n8273), .A2(n7606), .ZN(n10949) );
  INV_X1 U11066 ( .A(n11134), .ZN(n10951) );
  OR2_X1 U11067 ( .A1(n11135), .A2(n11136), .ZN(n11134) );
  AND2_X1 U11068 ( .A1(n11137), .A2(n11138), .ZN(n11136) );
  OR2_X1 U11069 ( .A1(n11139), .A2(n7697), .ZN(n11138) );
  AND2_X1 U11070 ( .A1(n8243), .A2(n7691), .ZN(n11139) );
  AND2_X1 U11071 ( .A1(n10944), .A2(n11140), .ZN(n11135) );
  OR2_X1 U11072 ( .A1(n11141), .A2(n7701), .ZN(n11140) );
  AND2_X1 U11073 ( .A1(n8220), .A2(n7703), .ZN(n11141) );
  OR2_X1 U11074 ( .A1(n7662), .A2(n8273), .ZN(n10956) );
  XNOR2_X1 U11075 ( .A(n11142), .B(n11143), .ZN(n10953) );
  XNOR2_X1 U11076 ( .A(n11144), .B(n11145), .ZN(n11143) );
  OR2_X1 U11077 ( .A1(n7660), .A2(n8273), .ZN(n10960) );
  XOR2_X1 U11078 ( .A(n11146), .B(n11147), .Z(n10957) );
  XOR2_X1 U11079 ( .A(n11148), .B(n11149), .Z(n11147) );
  OR2_X1 U11080 ( .A1(n7658), .A2(n8273), .ZN(n10964) );
  XOR2_X1 U11081 ( .A(n11150), .B(n11151), .Z(n10961) );
  XOR2_X1 U11082 ( .A(n11152), .B(n11153), .Z(n11151) );
  OR2_X1 U11083 ( .A1(n7656), .A2(n8273), .ZN(n10968) );
  XOR2_X1 U11084 ( .A(n11154), .B(n11155), .Z(n10965) );
  XOR2_X1 U11085 ( .A(n11156), .B(n11157), .Z(n11155) );
  OR2_X1 U11086 ( .A1(n7654), .A2(n8273), .ZN(n10972) );
  XOR2_X1 U11087 ( .A(n11158), .B(n11159), .Z(n10969) );
  XOR2_X1 U11088 ( .A(n11160), .B(n11161), .Z(n11159) );
  OR2_X1 U11089 ( .A1(n7652), .A2(n8273), .ZN(n10976) );
  XOR2_X1 U11090 ( .A(n11162), .B(n11163), .Z(n10973) );
  XOR2_X1 U11091 ( .A(n11164), .B(n11165), .Z(n11163) );
  OR2_X1 U11092 ( .A1(n7650), .A2(n8273), .ZN(n10980) );
  XOR2_X1 U11093 ( .A(n11166), .B(n11167), .Z(n10977) );
  XOR2_X1 U11094 ( .A(n11168), .B(n11169), .Z(n11167) );
  OR2_X1 U11095 ( .A1(n7648), .A2(n8273), .ZN(n10984) );
  XOR2_X1 U11096 ( .A(n11170), .B(n11171), .Z(n10981) );
  XOR2_X1 U11097 ( .A(n11172), .B(n11173), .Z(n11171) );
  OR2_X1 U11098 ( .A1(n7646), .A2(n8273), .ZN(n10988) );
  XOR2_X1 U11099 ( .A(n11174), .B(n11175), .Z(n10985) );
  XOR2_X1 U11100 ( .A(n11176), .B(n11177), .Z(n11175) );
  OR2_X1 U11101 ( .A1(n7644), .A2(n8273), .ZN(n10992) );
  XOR2_X1 U11102 ( .A(n11178), .B(n11179), .Z(n10989) );
  XOR2_X1 U11103 ( .A(n11180), .B(n11181), .Z(n11179) );
  OR2_X1 U11104 ( .A1(n7642), .A2(n8273), .ZN(n10996) );
  XOR2_X1 U11105 ( .A(n11182), .B(n11183), .Z(n10993) );
  XOR2_X1 U11106 ( .A(n11184), .B(n11185), .Z(n11183) );
  OR2_X1 U11107 ( .A1(n7640), .A2(n8273), .ZN(n11000) );
  XOR2_X1 U11108 ( .A(n11186), .B(n11187), .Z(n10997) );
  XOR2_X1 U11109 ( .A(n11188), .B(n11189), .Z(n11187) );
  OR2_X1 U11110 ( .A1(n7638), .A2(n8273), .ZN(n11004) );
  XOR2_X1 U11111 ( .A(n11190), .B(n11191), .Z(n11001) );
  XOR2_X1 U11112 ( .A(n11192), .B(n11193), .Z(n11191) );
  OR2_X1 U11113 ( .A1(n7636), .A2(n8273), .ZN(n11008) );
  XOR2_X1 U11114 ( .A(n11194), .B(n11195), .Z(n11005) );
  XOR2_X1 U11115 ( .A(n11196), .B(n11197), .Z(n11195) );
  OR2_X1 U11116 ( .A1(n7634), .A2(n8273), .ZN(n11012) );
  XOR2_X1 U11117 ( .A(n11198), .B(n11199), .Z(n11009) );
  XOR2_X1 U11118 ( .A(n11200), .B(n11201), .Z(n11199) );
  OR2_X1 U11119 ( .A1(n7632), .A2(n8273), .ZN(n11016) );
  XOR2_X1 U11120 ( .A(n11202), .B(n11203), .Z(n11013) );
  XOR2_X1 U11121 ( .A(n11204), .B(n11205), .Z(n11203) );
  OR2_X1 U11122 ( .A1(n7630), .A2(n8273), .ZN(n11020) );
  XOR2_X1 U11123 ( .A(n11206), .B(n11207), .Z(n11017) );
  XOR2_X1 U11124 ( .A(n11208), .B(n11209), .Z(n11207) );
  OR2_X1 U11125 ( .A1(n7628), .A2(n8273), .ZN(n11024) );
  XOR2_X1 U11126 ( .A(n11210), .B(n11211), .Z(n11021) );
  XOR2_X1 U11127 ( .A(n11212), .B(n11213), .Z(n11211) );
  OR2_X1 U11128 ( .A1(n7626), .A2(n8273), .ZN(n11028) );
  XOR2_X1 U11129 ( .A(n11214), .B(n11215), .Z(n11025) );
  XOR2_X1 U11130 ( .A(n11216), .B(n11217), .Z(n11215) );
  OR2_X1 U11131 ( .A1(n8624), .A2(n8273), .ZN(n11032) );
  XOR2_X1 U11132 ( .A(n11218), .B(n11219), .Z(n11029) );
  XOR2_X1 U11133 ( .A(n11220), .B(n11221), .Z(n11219) );
  OR2_X1 U11134 ( .A1(n8629), .A2(n8273), .ZN(n11036) );
  XOR2_X1 U11135 ( .A(n11222), .B(n11223), .Z(n11033) );
  XOR2_X1 U11136 ( .A(n11224), .B(n11225), .Z(n11223) );
  OR2_X1 U11137 ( .A1(n8634), .A2(n8273), .ZN(n11040) );
  XOR2_X1 U11138 ( .A(n11226), .B(n11227), .Z(n11037) );
  XOR2_X1 U11139 ( .A(n11228), .B(n11229), .Z(n11227) );
  OR2_X1 U11140 ( .A1(n8639), .A2(n8273), .ZN(n11044) );
  XOR2_X1 U11141 ( .A(n11230), .B(n11231), .Z(n11041) );
  XOR2_X1 U11142 ( .A(n11232), .B(n11233), .Z(n11231) );
  OR2_X1 U11143 ( .A1(n8644), .A2(n8273), .ZN(n11048) );
  XOR2_X1 U11144 ( .A(n11234), .B(n11235), .Z(n11045) );
  XOR2_X1 U11145 ( .A(n11236), .B(n11237), .Z(n11235) );
  OR2_X1 U11146 ( .A1(n8152), .A2(n8273), .ZN(n11054) );
  INV_X1 U11147 ( .A(n10744), .ZN(n8273) );
  XOR2_X1 U11148 ( .A(n11238), .B(n11239), .Z(n10744) );
  XNOR2_X1 U11149 ( .A(c_19_), .B(d_19_), .ZN(n11238) );
  XOR2_X1 U11150 ( .A(n11240), .B(n11241), .Z(n11051) );
  XOR2_X1 U11151 ( .A(n11242), .B(n11243), .Z(n11241) );
  XOR2_X1 U11152 ( .A(n10430), .B(n11244), .Z(n10423) );
  XOR2_X1 U11153 ( .A(n10429), .B(n10428), .Z(n11244) );
  OR2_X1 U11154 ( .A1(n8152), .A2(n8243), .ZN(n10428) );
  OR2_X1 U11155 ( .A1(n11245), .A2(n11246), .ZN(n10429) );
  AND2_X1 U11156 ( .A1(n11243), .A2(n11242), .ZN(n11246) );
  AND2_X1 U11157 ( .A1(n11240), .A2(n11247), .ZN(n11245) );
  OR2_X1 U11158 ( .A1(n11243), .A2(n11242), .ZN(n11247) );
  OR2_X1 U11159 ( .A1(n11248), .A2(n11249), .ZN(n11242) );
  AND2_X1 U11160 ( .A1(n11237), .A2(n11236), .ZN(n11249) );
  AND2_X1 U11161 ( .A1(n11234), .A2(n11250), .ZN(n11248) );
  OR2_X1 U11162 ( .A1(n11237), .A2(n11236), .ZN(n11250) );
  OR2_X1 U11163 ( .A1(n11251), .A2(n11252), .ZN(n11236) );
  AND2_X1 U11164 ( .A1(n11233), .A2(n11232), .ZN(n11252) );
  AND2_X1 U11165 ( .A1(n11230), .A2(n11253), .ZN(n11251) );
  OR2_X1 U11166 ( .A1(n11233), .A2(n11232), .ZN(n11253) );
  OR2_X1 U11167 ( .A1(n11254), .A2(n11255), .ZN(n11232) );
  AND2_X1 U11168 ( .A1(n11229), .A2(n11228), .ZN(n11255) );
  AND2_X1 U11169 ( .A1(n11226), .A2(n11256), .ZN(n11254) );
  OR2_X1 U11170 ( .A1(n11229), .A2(n11228), .ZN(n11256) );
  OR2_X1 U11171 ( .A1(n11257), .A2(n11258), .ZN(n11228) );
  AND2_X1 U11172 ( .A1(n11225), .A2(n11224), .ZN(n11258) );
  AND2_X1 U11173 ( .A1(n11222), .A2(n11259), .ZN(n11257) );
  OR2_X1 U11174 ( .A1(n11225), .A2(n11224), .ZN(n11259) );
  OR2_X1 U11175 ( .A1(n11260), .A2(n11261), .ZN(n11224) );
  AND2_X1 U11176 ( .A1(n11221), .A2(n11220), .ZN(n11261) );
  AND2_X1 U11177 ( .A1(n11218), .A2(n11262), .ZN(n11260) );
  OR2_X1 U11178 ( .A1(n11221), .A2(n11220), .ZN(n11262) );
  OR2_X1 U11179 ( .A1(n11263), .A2(n11264), .ZN(n11220) );
  AND2_X1 U11180 ( .A1(n11217), .A2(n11216), .ZN(n11264) );
  AND2_X1 U11181 ( .A1(n11214), .A2(n11265), .ZN(n11263) );
  OR2_X1 U11182 ( .A1(n11217), .A2(n11216), .ZN(n11265) );
  OR2_X1 U11183 ( .A1(n11266), .A2(n11267), .ZN(n11216) );
  AND2_X1 U11184 ( .A1(n11213), .A2(n11212), .ZN(n11267) );
  AND2_X1 U11185 ( .A1(n11210), .A2(n11268), .ZN(n11266) );
  OR2_X1 U11186 ( .A1(n11213), .A2(n11212), .ZN(n11268) );
  OR2_X1 U11187 ( .A1(n11269), .A2(n11270), .ZN(n11212) );
  AND2_X1 U11188 ( .A1(n11209), .A2(n11208), .ZN(n11270) );
  AND2_X1 U11189 ( .A1(n11206), .A2(n11271), .ZN(n11269) );
  OR2_X1 U11190 ( .A1(n11209), .A2(n11208), .ZN(n11271) );
  OR2_X1 U11191 ( .A1(n11272), .A2(n11273), .ZN(n11208) );
  AND2_X1 U11192 ( .A1(n11205), .A2(n11204), .ZN(n11273) );
  AND2_X1 U11193 ( .A1(n11202), .A2(n11274), .ZN(n11272) );
  OR2_X1 U11194 ( .A1(n11205), .A2(n11204), .ZN(n11274) );
  OR2_X1 U11195 ( .A1(n11275), .A2(n11276), .ZN(n11204) );
  AND2_X1 U11196 ( .A1(n11201), .A2(n11200), .ZN(n11276) );
  AND2_X1 U11197 ( .A1(n11198), .A2(n11277), .ZN(n11275) );
  OR2_X1 U11198 ( .A1(n11201), .A2(n11200), .ZN(n11277) );
  OR2_X1 U11199 ( .A1(n11278), .A2(n11279), .ZN(n11200) );
  AND2_X1 U11200 ( .A1(n11197), .A2(n11196), .ZN(n11279) );
  AND2_X1 U11201 ( .A1(n11194), .A2(n11280), .ZN(n11278) );
  OR2_X1 U11202 ( .A1(n11197), .A2(n11196), .ZN(n11280) );
  OR2_X1 U11203 ( .A1(n11281), .A2(n11282), .ZN(n11196) );
  AND2_X1 U11204 ( .A1(n11193), .A2(n11192), .ZN(n11282) );
  AND2_X1 U11205 ( .A1(n11190), .A2(n11283), .ZN(n11281) );
  OR2_X1 U11206 ( .A1(n11193), .A2(n11192), .ZN(n11283) );
  OR2_X1 U11207 ( .A1(n11284), .A2(n11285), .ZN(n11192) );
  AND2_X1 U11208 ( .A1(n11189), .A2(n11188), .ZN(n11285) );
  AND2_X1 U11209 ( .A1(n11186), .A2(n11286), .ZN(n11284) );
  OR2_X1 U11210 ( .A1(n11189), .A2(n11188), .ZN(n11286) );
  OR2_X1 U11211 ( .A1(n11287), .A2(n11288), .ZN(n11188) );
  AND2_X1 U11212 ( .A1(n11185), .A2(n11184), .ZN(n11288) );
  AND2_X1 U11213 ( .A1(n11182), .A2(n11289), .ZN(n11287) );
  OR2_X1 U11214 ( .A1(n11185), .A2(n11184), .ZN(n11289) );
  OR2_X1 U11215 ( .A1(n11290), .A2(n11291), .ZN(n11184) );
  AND2_X1 U11216 ( .A1(n11181), .A2(n11180), .ZN(n11291) );
  AND2_X1 U11217 ( .A1(n11178), .A2(n11292), .ZN(n11290) );
  OR2_X1 U11218 ( .A1(n11181), .A2(n11180), .ZN(n11292) );
  OR2_X1 U11219 ( .A1(n11293), .A2(n11294), .ZN(n11180) );
  AND2_X1 U11220 ( .A1(n11177), .A2(n11176), .ZN(n11294) );
  AND2_X1 U11221 ( .A1(n11174), .A2(n11295), .ZN(n11293) );
  OR2_X1 U11222 ( .A1(n11177), .A2(n11176), .ZN(n11295) );
  OR2_X1 U11223 ( .A1(n11296), .A2(n11297), .ZN(n11176) );
  AND2_X1 U11224 ( .A1(n11173), .A2(n11172), .ZN(n11297) );
  AND2_X1 U11225 ( .A1(n11170), .A2(n11298), .ZN(n11296) );
  OR2_X1 U11226 ( .A1(n11173), .A2(n11172), .ZN(n11298) );
  OR2_X1 U11227 ( .A1(n11299), .A2(n11300), .ZN(n11172) );
  AND2_X1 U11228 ( .A1(n11169), .A2(n11168), .ZN(n11300) );
  AND2_X1 U11229 ( .A1(n11166), .A2(n11301), .ZN(n11299) );
  OR2_X1 U11230 ( .A1(n11169), .A2(n11168), .ZN(n11301) );
  OR2_X1 U11231 ( .A1(n11302), .A2(n11303), .ZN(n11168) );
  AND2_X1 U11232 ( .A1(n11165), .A2(n11164), .ZN(n11303) );
  AND2_X1 U11233 ( .A1(n11162), .A2(n11304), .ZN(n11302) );
  OR2_X1 U11234 ( .A1(n11165), .A2(n11164), .ZN(n11304) );
  OR2_X1 U11235 ( .A1(n11305), .A2(n11306), .ZN(n11164) );
  AND2_X1 U11236 ( .A1(n11161), .A2(n11160), .ZN(n11306) );
  AND2_X1 U11237 ( .A1(n11158), .A2(n11307), .ZN(n11305) );
  OR2_X1 U11238 ( .A1(n11161), .A2(n11160), .ZN(n11307) );
  OR2_X1 U11239 ( .A1(n11308), .A2(n11309), .ZN(n11160) );
  AND2_X1 U11240 ( .A1(n11157), .A2(n11156), .ZN(n11309) );
  AND2_X1 U11241 ( .A1(n11154), .A2(n11310), .ZN(n11308) );
  OR2_X1 U11242 ( .A1(n11157), .A2(n11156), .ZN(n11310) );
  OR2_X1 U11243 ( .A1(n11311), .A2(n11312), .ZN(n11156) );
  AND2_X1 U11244 ( .A1(n11153), .A2(n11152), .ZN(n11312) );
  AND2_X1 U11245 ( .A1(n11150), .A2(n11313), .ZN(n11311) );
  OR2_X1 U11246 ( .A1(n11153), .A2(n11152), .ZN(n11313) );
  OR2_X1 U11247 ( .A1(n11314), .A2(n11315), .ZN(n11152) );
  AND2_X1 U11248 ( .A1(n11149), .A2(n11148), .ZN(n11315) );
  AND2_X1 U11249 ( .A1(n11146), .A2(n11316), .ZN(n11314) );
  OR2_X1 U11250 ( .A1(n11149), .A2(n11148), .ZN(n11316) );
  OR2_X1 U11251 ( .A1(n11317), .A2(n11318), .ZN(n11148) );
  AND2_X1 U11252 ( .A1(n11142), .A2(n11145), .ZN(n11318) );
  AND2_X1 U11253 ( .A1(n11144), .A2(n11319), .ZN(n11317) );
  OR2_X1 U11254 ( .A1(n11142), .A2(n11145), .ZN(n11319) );
  OR3_X1 U11255 ( .A1(n8220), .A2(n8243), .A3(n8519), .ZN(n11145) );
  OR2_X1 U11256 ( .A1(n8243), .A2(n7606), .ZN(n11142) );
  INV_X1 U11257 ( .A(n11320), .ZN(n11144) );
  OR2_X1 U11258 ( .A1(n11321), .A2(n11322), .ZN(n11320) );
  AND2_X1 U11259 ( .A1(n11323), .A2(n11324), .ZN(n11322) );
  OR2_X1 U11260 ( .A1(n11325), .A2(n7697), .ZN(n11324) );
  AND2_X1 U11261 ( .A1(n8220), .A2(n7691), .ZN(n11325) );
  AND2_X1 U11262 ( .A1(n11137), .A2(n11326), .ZN(n11321) );
  OR2_X1 U11263 ( .A1(n11327), .A2(n7701), .ZN(n11326) );
  AND2_X1 U11264 ( .A1(n11328), .A2(n7703), .ZN(n11327) );
  OR2_X1 U11265 ( .A1(n7662), .A2(n8243), .ZN(n11149) );
  XNOR2_X1 U11266 ( .A(n11329), .B(n11330), .ZN(n11146) );
  XNOR2_X1 U11267 ( .A(n11331), .B(n11332), .ZN(n11330) );
  OR2_X1 U11268 ( .A1(n7660), .A2(n8243), .ZN(n11153) );
  XOR2_X1 U11269 ( .A(n11333), .B(n11334), .Z(n11150) );
  XOR2_X1 U11270 ( .A(n11335), .B(n11336), .Z(n11334) );
  OR2_X1 U11271 ( .A1(n7658), .A2(n8243), .ZN(n11157) );
  XOR2_X1 U11272 ( .A(n11337), .B(n11338), .Z(n11154) );
  XOR2_X1 U11273 ( .A(n11339), .B(n11340), .Z(n11338) );
  OR2_X1 U11274 ( .A1(n7656), .A2(n8243), .ZN(n11161) );
  XOR2_X1 U11275 ( .A(n11341), .B(n11342), .Z(n11158) );
  XOR2_X1 U11276 ( .A(n11343), .B(n11344), .Z(n11342) );
  OR2_X1 U11277 ( .A1(n7654), .A2(n8243), .ZN(n11165) );
  XOR2_X1 U11278 ( .A(n11345), .B(n11346), .Z(n11162) );
  XOR2_X1 U11279 ( .A(n11347), .B(n11348), .Z(n11346) );
  OR2_X1 U11280 ( .A1(n7652), .A2(n8243), .ZN(n11169) );
  XOR2_X1 U11281 ( .A(n11349), .B(n11350), .Z(n11166) );
  XOR2_X1 U11282 ( .A(n11351), .B(n11352), .Z(n11350) );
  OR2_X1 U11283 ( .A1(n7650), .A2(n8243), .ZN(n11173) );
  XOR2_X1 U11284 ( .A(n11353), .B(n11354), .Z(n11170) );
  XOR2_X1 U11285 ( .A(n11355), .B(n11356), .Z(n11354) );
  OR2_X1 U11286 ( .A1(n7648), .A2(n8243), .ZN(n11177) );
  XOR2_X1 U11287 ( .A(n11357), .B(n11358), .Z(n11174) );
  XOR2_X1 U11288 ( .A(n11359), .B(n11360), .Z(n11358) );
  OR2_X1 U11289 ( .A1(n7646), .A2(n8243), .ZN(n11181) );
  XOR2_X1 U11290 ( .A(n11361), .B(n11362), .Z(n11178) );
  XOR2_X1 U11291 ( .A(n11363), .B(n11364), .Z(n11362) );
  OR2_X1 U11292 ( .A1(n7644), .A2(n8243), .ZN(n11185) );
  XOR2_X1 U11293 ( .A(n11365), .B(n11366), .Z(n11182) );
  XOR2_X1 U11294 ( .A(n11367), .B(n11368), .Z(n11366) );
  OR2_X1 U11295 ( .A1(n7642), .A2(n8243), .ZN(n11189) );
  XOR2_X1 U11296 ( .A(n11369), .B(n11370), .Z(n11186) );
  XOR2_X1 U11297 ( .A(n11371), .B(n11372), .Z(n11370) );
  OR2_X1 U11298 ( .A1(n7640), .A2(n8243), .ZN(n11193) );
  XOR2_X1 U11299 ( .A(n11373), .B(n11374), .Z(n11190) );
  XOR2_X1 U11300 ( .A(n11375), .B(n11376), .Z(n11374) );
  OR2_X1 U11301 ( .A1(n7638), .A2(n8243), .ZN(n11197) );
  XOR2_X1 U11302 ( .A(n11377), .B(n11378), .Z(n11194) );
  XOR2_X1 U11303 ( .A(n11379), .B(n11380), .Z(n11378) );
  OR2_X1 U11304 ( .A1(n7636), .A2(n8243), .ZN(n11201) );
  XOR2_X1 U11305 ( .A(n11381), .B(n11382), .Z(n11198) );
  XOR2_X1 U11306 ( .A(n11383), .B(n11384), .Z(n11382) );
  OR2_X1 U11307 ( .A1(n7634), .A2(n8243), .ZN(n11205) );
  XOR2_X1 U11308 ( .A(n11385), .B(n11386), .Z(n11202) );
  XOR2_X1 U11309 ( .A(n11387), .B(n11388), .Z(n11386) );
  OR2_X1 U11310 ( .A1(n7632), .A2(n8243), .ZN(n11209) );
  XOR2_X1 U11311 ( .A(n11389), .B(n11390), .Z(n11206) );
  XOR2_X1 U11312 ( .A(n11391), .B(n11392), .Z(n11390) );
  OR2_X1 U11313 ( .A1(n7630), .A2(n8243), .ZN(n11213) );
  XOR2_X1 U11314 ( .A(n11393), .B(n11394), .Z(n11210) );
  XOR2_X1 U11315 ( .A(n11395), .B(n11396), .Z(n11394) );
  OR2_X1 U11316 ( .A1(n7628), .A2(n8243), .ZN(n11217) );
  XOR2_X1 U11317 ( .A(n11397), .B(n11398), .Z(n11214) );
  XOR2_X1 U11318 ( .A(n11399), .B(n11400), .Z(n11398) );
  OR2_X1 U11319 ( .A1(n8619), .A2(n8243), .ZN(n11221) );
  XOR2_X1 U11320 ( .A(n11401), .B(n11402), .Z(n11218) );
  XOR2_X1 U11321 ( .A(n11403), .B(n11404), .Z(n11402) );
  OR2_X1 U11322 ( .A1(n8624), .A2(n8243), .ZN(n11225) );
  XOR2_X1 U11323 ( .A(n11405), .B(n11406), .Z(n11222) );
  XOR2_X1 U11324 ( .A(n11407), .B(n11408), .Z(n11406) );
  OR2_X1 U11325 ( .A1(n8629), .A2(n8243), .ZN(n11229) );
  XOR2_X1 U11326 ( .A(n11409), .B(n11410), .Z(n11226) );
  XOR2_X1 U11327 ( .A(n11411), .B(n11412), .Z(n11410) );
  OR2_X1 U11328 ( .A1(n8634), .A2(n8243), .ZN(n11233) );
  XOR2_X1 U11329 ( .A(n11413), .B(n11414), .Z(n11230) );
  XOR2_X1 U11330 ( .A(n11415), .B(n11416), .Z(n11414) );
  OR2_X1 U11331 ( .A1(n8639), .A2(n8243), .ZN(n11237) );
  XOR2_X1 U11332 ( .A(n11417), .B(n11418), .Z(n11234) );
  XOR2_X1 U11333 ( .A(n11419), .B(n11420), .Z(n11418) );
  OR2_X1 U11334 ( .A1(n8644), .A2(n8243), .ZN(n11243) );
  INV_X1 U11335 ( .A(n10944), .ZN(n8243) );
  XOR2_X1 U11336 ( .A(n11421), .B(n11422), .Z(n10944) );
  XNOR2_X1 U11337 ( .A(c_18_), .B(d_18_), .ZN(n11421) );
  XOR2_X1 U11338 ( .A(n11423), .B(n11424), .Z(n11240) );
  XOR2_X1 U11339 ( .A(n11425), .B(n11426), .Z(n11424) );
  XOR2_X1 U11340 ( .A(n10437), .B(n11427), .Z(n10430) );
  XOR2_X1 U11341 ( .A(n10436), .B(n10435), .Z(n11427) );
  OR2_X1 U11342 ( .A1(n8644), .A2(n8220), .ZN(n10435) );
  OR2_X1 U11343 ( .A1(n11428), .A2(n11429), .ZN(n10436) );
  AND2_X1 U11344 ( .A1(n11426), .A2(n11425), .ZN(n11429) );
  AND2_X1 U11345 ( .A1(n11423), .A2(n11430), .ZN(n11428) );
  OR2_X1 U11346 ( .A1(n11426), .A2(n11425), .ZN(n11430) );
  OR2_X1 U11347 ( .A1(n11431), .A2(n11432), .ZN(n11425) );
  AND2_X1 U11348 ( .A1(n11420), .A2(n11419), .ZN(n11432) );
  AND2_X1 U11349 ( .A1(n11417), .A2(n11433), .ZN(n11431) );
  OR2_X1 U11350 ( .A1(n11420), .A2(n11419), .ZN(n11433) );
  OR2_X1 U11351 ( .A1(n11434), .A2(n11435), .ZN(n11419) );
  AND2_X1 U11352 ( .A1(n11416), .A2(n11415), .ZN(n11435) );
  AND2_X1 U11353 ( .A1(n11413), .A2(n11436), .ZN(n11434) );
  OR2_X1 U11354 ( .A1(n11416), .A2(n11415), .ZN(n11436) );
  OR2_X1 U11355 ( .A1(n11437), .A2(n11438), .ZN(n11415) );
  AND2_X1 U11356 ( .A1(n11412), .A2(n11411), .ZN(n11438) );
  AND2_X1 U11357 ( .A1(n11409), .A2(n11439), .ZN(n11437) );
  OR2_X1 U11358 ( .A1(n11412), .A2(n11411), .ZN(n11439) );
  OR2_X1 U11359 ( .A1(n11440), .A2(n11441), .ZN(n11411) );
  AND2_X1 U11360 ( .A1(n11408), .A2(n11407), .ZN(n11441) );
  AND2_X1 U11361 ( .A1(n11405), .A2(n11442), .ZN(n11440) );
  OR2_X1 U11362 ( .A1(n11408), .A2(n11407), .ZN(n11442) );
  OR2_X1 U11363 ( .A1(n11443), .A2(n11444), .ZN(n11407) );
  AND2_X1 U11364 ( .A1(n11404), .A2(n11403), .ZN(n11444) );
  AND2_X1 U11365 ( .A1(n11401), .A2(n11445), .ZN(n11443) );
  OR2_X1 U11366 ( .A1(n11404), .A2(n11403), .ZN(n11445) );
  OR2_X1 U11367 ( .A1(n11446), .A2(n11447), .ZN(n11403) );
  AND2_X1 U11368 ( .A1(n11400), .A2(n11399), .ZN(n11447) );
  AND2_X1 U11369 ( .A1(n11397), .A2(n11448), .ZN(n11446) );
  OR2_X1 U11370 ( .A1(n11400), .A2(n11399), .ZN(n11448) );
  OR2_X1 U11371 ( .A1(n11449), .A2(n11450), .ZN(n11399) );
  AND2_X1 U11372 ( .A1(n11396), .A2(n11395), .ZN(n11450) );
  AND2_X1 U11373 ( .A1(n11393), .A2(n11451), .ZN(n11449) );
  OR2_X1 U11374 ( .A1(n11396), .A2(n11395), .ZN(n11451) );
  OR2_X1 U11375 ( .A1(n11452), .A2(n11453), .ZN(n11395) );
  AND2_X1 U11376 ( .A1(n11392), .A2(n11391), .ZN(n11453) );
  AND2_X1 U11377 ( .A1(n11389), .A2(n11454), .ZN(n11452) );
  OR2_X1 U11378 ( .A1(n11392), .A2(n11391), .ZN(n11454) );
  OR2_X1 U11379 ( .A1(n11455), .A2(n11456), .ZN(n11391) );
  AND2_X1 U11380 ( .A1(n11388), .A2(n11387), .ZN(n11456) );
  AND2_X1 U11381 ( .A1(n11385), .A2(n11457), .ZN(n11455) );
  OR2_X1 U11382 ( .A1(n11388), .A2(n11387), .ZN(n11457) );
  OR2_X1 U11383 ( .A1(n11458), .A2(n11459), .ZN(n11387) );
  AND2_X1 U11384 ( .A1(n11384), .A2(n11383), .ZN(n11459) );
  AND2_X1 U11385 ( .A1(n11381), .A2(n11460), .ZN(n11458) );
  OR2_X1 U11386 ( .A1(n11384), .A2(n11383), .ZN(n11460) );
  OR2_X1 U11387 ( .A1(n11461), .A2(n11462), .ZN(n11383) );
  AND2_X1 U11388 ( .A1(n11380), .A2(n11379), .ZN(n11462) );
  AND2_X1 U11389 ( .A1(n11377), .A2(n11463), .ZN(n11461) );
  OR2_X1 U11390 ( .A1(n11380), .A2(n11379), .ZN(n11463) );
  OR2_X1 U11391 ( .A1(n11464), .A2(n11465), .ZN(n11379) );
  AND2_X1 U11392 ( .A1(n11376), .A2(n11375), .ZN(n11465) );
  AND2_X1 U11393 ( .A1(n11373), .A2(n11466), .ZN(n11464) );
  OR2_X1 U11394 ( .A1(n11376), .A2(n11375), .ZN(n11466) );
  OR2_X1 U11395 ( .A1(n11467), .A2(n11468), .ZN(n11375) );
  AND2_X1 U11396 ( .A1(n11372), .A2(n11371), .ZN(n11468) );
  AND2_X1 U11397 ( .A1(n11369), .A2(n11469), .ZN(n11467) );
  OR2_X1 U11398 ( .A1(n11372), .A2(n11371), .ZN(n11469) );
  OR2_X1 U11399 ( .A1(n11470), .A2(n11471), .ZN(n11371) );
  AND2_X1 U11400 ( .A1(n11368), .A2(n11367), .ZN(n11471) );
  AND2_X1 U11401 ( .A1(n11365), .A2(n11472), .ZN(n11470) );
  OR2_X1 U11402 ( .A1(n11368), .A2(n11367), .ZN(n11472) );
  OR2_X1 U11403 ( .A1(n11473), .A2(n11474), .ZN(n11367) );
  AND2_X1 U11404 ( .A1(n11364), .A2(n11363), .ZN(n11474) );
  AND2_X1 U11405 ( .A1(n11361), .A2(n11475), .ZN(n11473) );
  OR2_X1 U11406 ( .A1(n11364), .A2(n11363), .ZN(n11475) );
  OR2_X1 U11407 ( .A1(n11476), .A2(n11477), .ZN(n11363) );
  AND2_X1 U11408 ( .A1(n11360), .A2(n11359), .ZN(n11477) );
  AND2_X1 U11409 ( .A1(n11357), .A2(n11478), .ZN(n11476) );
  OR2_X1 U11410 ( .A1(n11360), .A2(n11359), .ZN(n11478) );
  OR2_X1 U11411 ( .A1(n11479), .A2(n11480), .ZN(n11359) );
  AND2_X1 U11412 ( .A1(n11356), .A2(n11355), .ZN(n11480) );
  AND2_X1 U11413 ( .A1(n11353), .A2(n11481), .ZN(n11479) );
  OR2_X1 U11414 ( .A1(n11356), .A2(n11355), .ZN(n11481) );
  OR2_X1 U11415 ( .A1(n11482), .A2(n11483), .ZN(n11355) );
  AND2_X1 U11416 ( .A1(n11352), .A2(n11351), .ZN(n11483) );
  AND2_X1 U11417 ( .A1(n11349), .A2(n11484), .ZN(n11482) );
  OR2_X1 U11418 ( .A1(n11352), .A2(n11351), .ZN(n11484) );
  OR2_X1 U11419 ( .A1(n11485), .A2(n11486), .ZN(n11351) );
  AND2_X1 U11420 ( .A1(n11348), .A2(n11347), .ZN(n11486) );
  AND2_X1 U11421 ( .A1(n11345), .A2(n11487), .ZN(n11485) );
  OR2_X1 U11422 ( .A1(n11348), .A2(n11347), .ZN(n11487) );
  OR2_X1 U11423 ( .A1(n11488), .A2(n11489), .ZN(n11347) );
  AND2_X1 U11424 ( .A1(n11344), .A2(n11343), .ZN(n11489) );
  AND2_X1 U11425 ( .A1(n11341), .A2(n11490), .ZN(n11488) );
  OR2_X1 U11426 ( .A1(n11344), .A2(n11343), .ZN(n11490) );
  OR2_X1 U11427 ( .A1(n11491), .A2(n11492), .ZN(n11343) );
  AND2_X1 U11428 ( .A1(n11340), .A2(n11339), .ZN(n11492) );
  AND2_X1 U11429 ( .A1(n11337), .A2(n11493), .ZN(n11491) );
  OR2_X1 U11430 ( .A1(n11340), .A2(n11339), .ZN(n11493) );
  OR2_X1 U11431 ( .A1(n11494), .A2(n11495), .ZN(n11339) );
  AND2_X1 U11432 ( .A1(n11336), .A2(n11335), .ZN(n11495) );
  AND2_X1 U11433 ( .A1(n11333), .A2(n11496), .ZN(n11494) );
  OR2_X1 U11434 ( .A1(n11336), .A2(n11335), .ZN(n11496) );
  OR2_X1 U11435 ( .A1(n11497), .A2(n11498), .ZN(n11335) );
  AND2_X1 U11436 ( .A1(n11329), .A2(n11332), .ZN(n11498) );
  AND2_X1 U11437 ( .A1(n11331), .A2(n11499), .ZN(n11497) );
  OR2_X1 U11438 ( .A1(n11329), .A2(n11332), .ZN(n11499) );
  OR3_X1 U11439 ( .A1(n11328), .A2(n8220), .A3(n8519), .ZN(n11332) );
  OR2_X1 U11440 ( .A1(n8220), .A2(n7606), .ZN(n11329) );
  INV_X1 U11441 ( .A(n11500), .ZN(n11331) );
  OR2_X1 U11442 ( .A1(n11501), .A2(n11502), .ZN(n11500) );
  AND2_X1 U11443 ( .A1(n11503), .A2(n11504), .ZN(n11502) );
  OR2_X1 U11444 ( .A1(n11505), .A2(n7697), .ZN(n11504) );
  AND2_X1 U11445 ( .A1(n11328), .A2(n7691), .ZN(n11505) );
  AND2_X1 U11446 ( .A1(n11323), .A2(n11506), .ZN(n11501) );
  OR2_X1 U11447 ( .A1(n11507), .A2(n7701), .ZN(n11506) );
  AND2_X1 U11448 ( .A1(n11508), .A2(n7703), .ZN(n11507) );
  OR2_X1 U11449 ( .A1(n7662), .A2(n8220), .ZN(n11336) );
  XNOR2_X1 U11450 ( .A(n11509), .B(n11510), .ZN(n11333) );
  XNOR2_X1 U11451 ( .A(n11511), .B(n11512), .ZN(n11510) );
  OR2_X1 U11452 ( .A1(n7660), .A2(n8220), .ZN(n11340) );
  XOR2_X1 U11453 ( .A(n11513), .B(n11514), .Z(n11337) );
  XOR2_X1 U11454 ( .A(n11515), .B(n11516), .Z(n11514) );
  OR2_X1 U11455 ( .A1(n7658), .A2(n8220), .ZN(n11344) );
  XOR2_X1 U11456 ( .A(n11517), .B(n11518), .Z(n11341) );
  XOR2_X1 U11457 ( .A(n11519), .B(n11520), .Z(n11518) );
  OR2_X1 U11458 ( .A1(n7656), .A2(n8220), .ZN(n11348) );
  XOR2_X1 U11459 ( .A(n11521), .B(n11522), .Z(n11345) );
  XOR2_X1 U11460 ( .A(n11523), .B(n11524), .Z(n11522) );
  OR2_X1 U11461 ( .A1(n7654), .A2(n8220), .ZN(n11352) );
  XOR2_X1 U11462 ( .A(n11525), .B(n11526), .Z(n11349) );
  XOR2_X1 U11463 ( .A(n11527), .B(n11528), .Z(n11526) );
  OR2_X1 U11464 ( .A1(n7652), .A2(n8220), .ZN(n11356) );
  XOR2_X1 U11465 ( .A(n11529), .B(n11530), .Z(n11353) );
  XOR2_X1 U11466 ( .A(n11531), .B(n11532), .Z(n11530) );
  OR2_X1 U11467 ( .A1(n7650), .A2(n8220), .ZN(n11360) );
  XOR2_X1 U11468 ( .A(n11533), .B(n11534), .Z(n11357) );
  XOR2_X1 U11469 ( .A(n11535), .B(n11536), .Z(n11534) );
  OR2_X1 U11470 ( .A1(n7648), .A2(n8220), .ZN(n11364) );
  XOR2_X1 U11471 ( .A(n11537), .B(n11538), .Z(n11361) );
  XOR2_X1 U11472 ( .A(n11539), .B(n11540), .Z(n11538) );
  OR2_X1 U11473 ( .A1(n7646), .A2(n8220), .ZN(n11368) );
  XOR2_X1 U11474 ( .A(n11541), .B(n11542), .Z(n11365) );
  XOR2_X1 U11475 ( .A(n11543), .B(n11544), .Z(n11542) );
  OR2_X1 U11476 ( .A1(n7644), .A2(n8220), .ZN(n11372) );
  XOR2_X1 U11477 ( .A(n11545), .B(n11546), .Z(n11369) );
  XOR2_X1 U11478 ( .A(n11547), .B(n11548), .Z(n11546) );
  OR2_X1 U11479 ( .A1(n7642), .A2(n8220), .ZN(n11376) );
  XOR2_X1 U11480 ( .A(n11549), .B(n11550), .Z(n11373) );
  XOR2_X1 U11481 ( .A(n11551), .B(n11552), .Z(n11550) );
  OR2_X1 U11482 ( .A1(n7640), .A2(n8220), .ZN(n11380) );
  XOR2_X1 U11483 ( .A(n11553), .B(n11554), .Z(n11377) );
  XOR2_X1 U11484 ( .A(n11555), .B(n11556), .Z(n11554) );
  OR2_X1 U11485 ( .A1(n7638), .A2(n8220), .ZN(n11384) );
  XOR2_X1 U11486 ( .A(n11557), .B(n11558), .Z(n11381) );
  XOR2_X1 U11487 ( .A(n11559), .B(n11560), .Z(n11558) );
  OR2_X1 U11488 ( .A1(n7636), .A2(n8220), .ZN(n11388) );
  XOR2_X1 U11489 ( .A(n11561), .B(n11562), .Z(n11385) );
  XOR2_X1 U11490 ( .A(n11563), .B(n11564), .Z(n11562) );
  OR2_X1 U11491 ( .A1(n7634), .A2(n8220), .ZN(n11392) );
  XOR2_X1 U11492 ( .A(n11565), .B(n11566), .Z(n11389) );
  XOR2_X1 U11493 ( .A(n11567), .B(n11568), .Z(n11566) );
  OR2_X1 U11494 ( .A1(n7632), .A2(n8220), .ZN(n11396) );
  XOR2_X1 U11495 ( .A(n11569), .B(n11570), .Z(n11393) );
  XOR2_X1 U11496 ( .A(n11571), .B(n11572), .Z(n11570) );
  OR2_X1 U11497 ( .A1(n7630), .A2(n8220), .ZN(n11400) );
  XOR2_X1 U11498 ( .A(n11573), .B(n11574), .Z(n11397) );
  XOR2_X1 U11499 ( .A(n11575), .B(n11576), .Z(n11574) );
  OR2_X1 U11500 ( .A1(n8614), .A2(n8220), .ZN(n11404) );
  XOR2_X1 U11501 ( .A(n11577), .B(n11578), .Z(n11401) );
  XOR2_X1 U11502 ( .A(n11579), .B(n11580), .Z(n11578) );
  OR2_X1 U11503 ( .A1(n8619), .A2(n8220), .ZN(n11408) );
  XOR2_X1 U11504 ( .A(n11581), .B(n11582), .Z(n11405) );
  XOR2_X1 U11505 ( .A(n11583), .B(n11584), .Z(n11582) );
  OR2_X1 U11506 ( .A1(n8624), .A2(n8220), .ZN(n11412) );
  XOR2_X1 U11507 ( .A(n11585), .B(n11586), .Z(n11409) );
  XOR2_X1 U11508 ( .A(n11587), .B(n11588), .Z(n11586) );
  OR2_X1 U11509 ( .A1(n8629), .A2(n8220), .ZN(n11416) );
  XOR2_X1 U11510 ( .A(n11589), .B(n11590), .Z(n11413) );
  XOR2_X1 U11511 ( .A(n11591), .B(n11592), .Z(n11590) );
  OR2_X1 U11512 ( .A1(n8634), .A2(n8220), .ZN(n11420) );
  XOR2_X1 U11513 ( .A(n11593), .B(n11594), .Z(n11417) );
  XOR2_X1 U11514 ( .A(n11595), .B(n11596), .Z(n11594) );
  OR2_X1 U11515 ( .A1(n8639), .A2(n8220), .ZN(n11426) );
  INV_X1 U11516 ( .A(n11137), .ZN(n8220) );
  XOR2_X1 U11517 ( .A(n11597), .B(n11598), .Z(n11137) );
  XNOR2_X1 U11518 ( .A(c_17_), .B(d_17_), .ZN(n11597) );
  XOR2_X1 U11519 ( .A(n11599), .B(n11600), .Z(n11423) );
  XOR2_X1 U11520 ( .A(n11601), .B(n11602), .Z(n11600) );
  XOR2_X1 U11521 ( .A(n11603), .B(n11604), .Z(n10437) );
  XOR2_X1 U11522 ( .A(n11605), .B(n11606), .Z(n11604) );
  OR2_X1 U11523 ( .A1(n8185), .A2(n8184), .ZN(n7933) );
  OR2_X1 U11524 ( .A1(n11607), .A2(n7937), .ZN(n8184) );
  INV_X1 U11525 ( .A(n11608), .ZN(n7937) );
  OR2_X1 U11526 ( .A1(n11609), .A2(n11610), .ZN(n11608) );
  AND2_X1 U11527 ( .A1(n11609), .A2(n11610), .ZN(n11607) );
  OR2_X1 U11528 ( .A1(n11611), .A2(n11612), .ZN(n11610) );
  AND2_X1 U11529 ( .A1(n11613), .A2(n11614), .ZN(n11612) );
  AND2_X1 U11530 ( .A1(n11615), .A2(n11616), .ZN(n11611) );
  OR2_X1 U11531 ( .A1(n11613), .A2(n11614), .ZN(n11616) );
  XOR2_X1 U11532 ( .A(n11617), .B(n11618), .Z(n11609) );
  XOR2_X1 U11533 ( .A(n11619), .B(n11620), .Z(n11618) );
  OR2_X1 U11534 ( .A1(n8191), .A2(n8192), .ZN(n8185) );
  OR2_X1 U11535 ( .A1(n11621), .A2(n11622), .ZN(n8192) );
  AND2_X1 U11536 ( .A1(n8207), .A2(n8206), .ZN(n11622) );
  AND2_X1 U11537 ( .A1(n8205), .A2(n11623), .ZN(n11621) );
  OR2_X1 U11538 ( .A1(n8207), .A2(n8206), .ZN(n11623) );
  OR2_X1 U11539 ( .A1(n11624), .A2(n11625), .ZN(n8206) );
  AND2_X1 U11540 ( .A1(n8230), .A2(n8229), .ZN(n11625) );
  AND2_X1 U11541 ( .A1(n8228), .A2(n11626), .ZN(n11624) );
  OR2_X1 U11542 ( .A1(n8230), .A2(n8229), .ZN(n11626) );
  OR2_X1 U11543 ( .A1(n11627), .A2(n11628), .ZN(n8229) );
  AND2_X1 U11544 ( .A1(n8260), .A2(n8259), .ZN(n11628) );
  AND2_X1 U11545 ( .A1(n8257), .A2(n11629), .ZN(n11627) );
  OR2_X1 U11546 ( .A1(n8260), .A2(n8259), .ZN(n11629) );
  OR2_X1 U11547 ( .A1(n11630), .A2(n11631), .ZN(n8259) );
  AND2_X1 U11548 ( .A1(n8297), .A2(n8296), .ZN(n11631) );
  AND2_X1 U11549 ( .A1(n8294), .A2(n11632), .ZN(n11630) );
  OR2_X1 U11550 ( .A1(n8297), .A2(n8296), .ZN(n11632) );
  OR2_X1 U11551 ( .A1(n11633), .A2(n11634), .ZN(n8296) );
  AND2_X1 U11552 ( .A1(n10403), .A2(n10402), .ZN(n11634) );
  AND2_X1 U11553 ( .A1(n10400), .A2(n11635), .ZN(n11633) );
  OR2_X1 U11554 ( .A1(n10403), .A2(n10402), .ZN(n11635) );
  OR2_X1 U11555 ( .A1(n11636), .A2(n11637), .ZN(n10402) );
  AND2_X1 U11556 ( .A1(n10442), .A2(n10441), .ZN(n11637) );
  AND2_X1 U11557 ( .A1(n10439), .A2(n11638), .ZN(n11636) );
  OR2_X1 U11558 ( .A1(n10442), .A2(n10441), .ZN(n11638) );
  OR2_X1 U11559 ( .A1(n11639), .A2(n11640), .ZN(n10441) );
  AND2_X1 U11560 ( .A1(n11606), .A2(n11605), .ZN(n11640) );
  AND2_X1 U11561 ( .A1(n11603), .A2(n11641), .ZN(n11639) );
  OR2_X1 U11562 ( .A1(n11606), .A2(n11605), .ZN(n11641) );
  OR2_X1 U11563 ( .A1(n11642), .A2(n11643), .ZN(n11605) );
  AND2_X1 U11564 ( .A1(n11602), .A2(n11601), .ZN(n11643) );
  AND2_X1 U11565 ( .A1(n11599), .A2(n11644), .ZN(n11642) );
  OR2_X1 U11566 ( .A1(n11602), .A2(n11601), .ZN(n11644) );
  OR2_X1 U11567 ( .A1(n11645), .A2(n11646), .ZN(n11601) );
  AND2_X1 U11568 ( .A1(n11596), .A2(n11595), .ZN(n11646) );
  AND2_X1 U11569 ( .A1(n11593), .A2(n11647), .ZN(n11645) );
  OR2_X1 U11570 ( .A1(n11596), .A2(n11595), .ZN(n11647) );
  OR2_X1 U11571 ( .A1(n11648), .A2(n11649), .ZN(n11595) );
  AND2_X1 U11572 ( .A1(n11592), .A2(n11591), .ZN(n11649) );
  AND2_X1 U11573 ( .A1(n11589), .A2(n11650), .ZN(n11648) );
  OR2_X1 U11574 ( .A1(n11592), .A2(n11591), .ZN(n11650) );
  OR2_X1 U11575 ( .A1(n11651), .A2(n11652), .ZN(n11591) );
  AND2_X1 U11576 ( .A1(n11588), .A2(n11587), .ZN(n11652) );
  AND2_X1 U11577 ( .A1(n11585), .A2(n11653), .ZN(n11651) );
  OR2_X1 U11578 ( .A1(n11588), .A2(n11587), .ZN(n11653) );
  OR2_X1 U11579 ( .A1(n11654), .A2(n11655), .ZN(n11587) );
  AND2_X1 U11580 ( .A1(n11584), .A2(n11583), .ZN(n11655) );
  AND2_X1 U11581 ( .A1(n11581), .A2(n11656), .ZN(n11654) );
  OR2_X1 U11582 ( .A1(n11584), .A2(n11583), .ZN(n11656) );
  OR2_X1 U11583 ( .A1(n11657), .A2(n11658), .ZN(n11583) );
  AND2_X1 U11584 ( .A1(n11580), .A2(n11579), .ZN(n11658) );
  AND2_X1 U11585 ( .A1(n11577), .A2(n11659), .ZN(n11657) );
  OR2_X1 U11586 ( .A1(n11580), .A2(n11579), .ZN(n11659) );
  OR2_X1 U11587 ( .A1(n11660), .A2(n11661), .ZN(n11579) );
  AND2_X1 U11588 ( .A1(n11576), .A2(n11575), .ZN(n11661) );
  AND2_X1 U11589 ( .A1(n11573), .A2(n11662), .ZN(n11660) );
  OR2_X1 U11590 ( .A1(n11576), .A2(n11575), .ZN(n11662) );
  OR2_X1 U11591 ( .A1(n11663), .A2(n11664), .ZN(n11575) );
  AND2_X1 U11592 ( .A1(n11572), .A2(n11571), .ZN(n11664) );
  AND2_X1 U11593 ( .A1(n11569), .A2(n11665), .ZN(n11663) );
  OR2_X1 U11594 ( .A1(n11572), .A2(n11571), .ZN(n11665) );
  OR2_X1 U11595 ( .A1(n11666), .A2(n11667), .ZN(n11571) );
  AND2_X1 U11596 ( .A1(n11568), .A2(n11567), .ZN(n11667) );
  AND2_X1 U11597 ( .A1(n11565), .A2(n11668), .ZN(n11666) );
  OR2_X1 U11598 ( .A1(n11568), .A2(n11567), .ZN(n11668) );
  OR2_X1 U11599 ( .A1(n11669), .A2(n11670), .ZN(n11567) );
  AND2_X1 U11600 ( .A1(n11564), .A2(n11563), .ZN(n11670) );
  AND2_X1 U11601 ( .A1(n11561), .A2(n11671), .ZN(n11669) );
  OR2_X1 U11602 ( .A1(n11564), .A2(n11563), .ZN(n11671) );
  OR2_X1 U11603 ( .A1(n11672), .A2(n11673), .ZN(n11563) );
  AND2_X1 U11604 ( .A1(n11560), .A2(n11559), .ZN(n11673) );
  AND2_X1 U11605 ( .A1(n11557), .A2(n11674), .ZN(n11672) );
  OR2_X1 U11606 ( .A1(n11560), .A2(n11559), .ZN(n11674) );
  OR2_X1 U11607 ( .A1(n11675), .A2(n11676), .ZN(n11559) );
  AND2_X1 U11608 ( .A1(n11556), .A2(n11555), .ZN(n11676) );
  AND2_X1 U11609 ( .A1(n11553), .A2(n11677), .ZN(n11675) );
  OR2_X1 U11610 ( .A1(n11556), .A2(n11555), .ZN(n11677) );
  OR2_X1 U11611 ( .A1(n11678), .A2(n11679), .ZN(n11555) );
  AND2_X1 U11612 ( .A1(n11552), .A2(n11551), .ZN(n11679) );
  AND2_X1 U11613 ( .A1(n11549), .A2(n11680), .ZN(n11678) );
  OR2_X1 U11614 ( .A1(n11552), .A2(n11551), .ZN(n11680) );
  OR2_X1 U11615 ( .A1(n11681), .A2(n11682), .ZN(n11551) );
  AND2_X1 U11616 ( .A1(n11548), .A2(n11547), .ZN(n11682) );
  AND2_X1 U11617 ( .A1(n11545), .A2(n11683), .ZN(n11681) );
  OR2_X1 U11618 ( .A1(n11548), .A2(n11547), .ZN(n11683) );
  OR2_X1 U11619 ( .A1(n11684), .A2(n11685), .ZN(n11547) );
  AND2_X1 U11620 ( .A1(n11544), .A2(n11543), .ZN(n11685) );
  AND2_X1 U11621 ( .A1(n11541), .A2(n11686), .ZN(n11684) );
  OR2_X1 U11622 ( .A1(n11544), .A2(n11543), .ZN(n11686) );
  OR2_X1 U11623 ( .A1(n11687), .A2(n11688), .ZN(n11543) );
  AND2_X1 U11624 ( .A1(n11540), .A2(n11539), .ZN(n11688) );
  AND2_X1 U11625 ( .A1(n11537), .A2(n11689), .ZN(n11687) );
  OR2_X1 U11626 ( .A1(n11540), .A2(n11539), .ZN(n11689) );
  OR2_X1 U11627 ( .A1(n11690), .A2(n11691), .ZN(n11539) );
  AND2_X1 U11628 ( .A1(n11536), .A2(n11535), .ZN(n11691) );
  AND2_X1 U11629 ( .A1(n11533), .A2(n11692), .ZN(n11690) );
  OR2_X1 U11630 ( .A1(n11536), .A2(n11535), .ZN(n11692) );
  OR2_X1 U11631 ( .A1(n11693), .A2(n11694), .ZN(n11535) );
  AND2_X1 U11632 ( .A1(n11532), .A2(n11531), .ZN(n11694) );
  AND2_X1 U11633 ( .A1(n11529), .A2(n11695), .ZN(n11693) );
  OR2_X1 U11634 ( .A1(n11532), .A2(n11531), .ZN(n11695) );
  OR2_X1 U11635 ( .A1(n11696), .A2(n11697), .ZN(n11531) );
  AND2_X1 U11636 ( .A1(n11528), .A2(n11527), .ZN(n11697) );
  AND2_X1 U11637 ( .A1(n11525), .A2(n11698), .ZN(n11696) );
  OR2_X1 U11638 ( .A1(n11528), .A2(n11527), .ZN(n11698) );
  OR2_X1 U11639 ( .A1(n11699), .A2(n11700), .ZN(n11527) );
  AND2_X1 U11640 ( .A1(n11524), .A2(n11523), .ZN(n11700) );
  AND2_X1 U11641 ( .A1(n11521), .A2(n11701), .ZN(n11699) );
  OR2_X1 U11642 ( .A1(n11524), .A2(n11523), .ZN(n11701) );
  OR2_X1 U11643 ( .A1(n11702), .A2(n11703), .ZN(n11523) );
  AND2_X1 U11644 ( .A1(n11520), .A2(n11519), .ZN(n11703) );
  AND2_X1 U11645 ( .A1(n11517), .A2(n11704), .ZN(n11702) );
  OR2_X1 U11646 ( .A1(n11520), .A2(n11519), .ZN(n11704) );
  OR2_X1 U11647 ( .A1(n11705), .A2(n11706), .ZN(n11519) );
  AND2_X1 U11648 ( .A1(n11516), .A2(n11515), .ZN(n11706) );
  AND2_X1 U11649 ( .A1(n11513), .A2(n11707), .ZN(n11705) );
  OR2_X1 U11650 ( .A1(n11516), .A2(n11515), .ZN(n11707) );
  OR2_X1 U11651 ( .A1(n11708), .A2(n11709), .ZN(n11515) );
  AND2_X1 U11652 ( .A1(n11509), .A2(n11512), .ZN(n11709) );
  AND2_X1 U11653 ( .A1(n11511), .A2(n11710), .ZN(n11708) );
  OR2_X1 U11654 ( .A1(n11509), .A2(n11512), .ZN(n11710) );
  OR3_X1 U11655 ( .A1(n11508), .A2(n11328), .A3(n8519), .ZN(n11512) );
  OR2_X1 U11656 ( .A1(n11328), .A2(n7606), .ZN(n11509) );
  INV_X1 U11657 ( .A(n11711), .ZN(n11511) );
  OR2_X1 U11658 ( .A1(n11712), .A2(n11713), .ZN(n11711) );
  AND2_X1 U11659 ( .A1(n11714), .A2(n11715), .ZN(n11713) );
  OR2_X1 U11660 ( .A1(n11716), .A2(n7697), .ZN(n11715) );
  AND2_X1 U11661 ( .A1(n11508), .A2(n7691), .ZN(n11716) );
  AND2_X1 U11662 ( .A1(n11503), .A2(n11717), .ZN(n11712) );
  OR2_X1 U11663 ( .A1(n11718), .A2(n7701), .ZN(n11717) );
  AND2_X1 U11664 ( .A1(n11719), .A2(n7703), .ZN(n11718) );
  OR2_X1 U11665 ( .A1(n7662), .A2(n11328), .ZN(n11516) );
  XNOR2_X1 U11666 ( .A(n11720), .B(n11721), .ZN(n11513) );
  XNOR2_X1 U11667 ( .A(n11722), .B(n11723), .ZN(n11721) );
  OR2_X1 U11668 ( .A1(n7660), .A2(n11328), .ZN(n11520) );
  XOR2_X1 U11669 ( .A(n11724), .B(n11725), .Z(n11517) );
  XOR2_X1 U11670 ( .A(n11726), .B(n11727), .Z(n11725) );
  OR2_X1 U11671 ( .A1(n7658), .A2(n11328), .ZN(n11524) );
  XOR2_X1 U11672 ( .A(n11728), .B(n11729), .Z(n11521) );
  XOR2_X1 U11673 ( .A(n11730), .B(n11731), .Z(n11729) );
  OR2_X1 U11674 ( .A1(n7656), .A2(n11328), .ZN(n11528) );
  XOR2_X1 U11675 ( .A(n11732), .B(n11733), .Z(n11525) );
  XOR2_X1 U11676 ( .A(n11734), .B(n11735), .Z(n11733) );
  OR2_X1 U11677 ( .A1(n7654), .A2(n11328), .ZN(n11532) );
  XOR2_X1 U11678 ( .A(n11736), .B(n11737), .Z(n11529) );
  XOR2_X1 U11679 ( .A(n11738), .B(n11739), .Z(n11737) );
  OR2_X1 U11680 ( .A1(n7652), .A2(n11328), .ZN(n11536) );
  XOR2_X1 U11681 ( .A(n11740), .B(n11741), .Z(n11533) );
  XOR2_X1 U11682 ( .A(n11742), .B(n11743), .Z(n11741) );
  OR2_X1 U11683 ( .A1(n7650), .A2(n11328), .ZN(n11540) );
  XOR2_X1 U11684 ( .A(n11744), .B(n11745), .Z(n11537) );
  XOR2_X1 U11685 ( .A(n11746), .B(n11747), .Z(n11745) );
  OR2_X1 U11686 ( .A1(n7648), .A2(n11328), .ZN(n11544) );
  XOR2_X1 U11687 ( .A(n11748), .B(n11749), .Z(n11541) );
  XOR2_X1 U11688 ( .A(n11750), .B(n11751), .Z(n11749) );
  OR2_X1 U11689 ( .A1(n7646), .A2(n11328), .ZN(n11548) );
  XOR2_X1 U11690 ( .A(n11752), .B(n11753), .Z(n11545) );
  XOR2_X1 U11691 ( .A(n11754), .B(n11755), .Z(n11753) );
  OR2_X1 U11692 ( .A1(n7644), .A2(n11328), .ZN(n11552) );
  XOR2_X1 U11693 ( .A(n11756), .B(n11757), .Z(n11549) );
  XOR2_X1 U11694 ( .A(n11758), .B(n11759), .Z(n11757) );
  OR2_X1 U11695 ( .A1(n7642), .A2(n11328), .ZN(n11556) );
  XOR2_X1 U11696 ( .A(n11760), .B(n11761), .Z(n11553) );
  XOR2_X1 U11697 ( .A(n11762), .B(n11763), .Z(n11761) );
  OR2_X1 U11698 ( .A1(n7640), .A2(n11328), .ZN(n11560) );
  XOR2_X1 U11699 ( .A(n11764), .B(n11765), .Z(n11557) );
  XOR2_X1 U11700 ( .A(n11766), .B(n11767), .Z(n11765) );
  OR2_X1 U11701 ( .A1(n7638), .A2(n11328), .ZN(n11564) );
  XOR2_X1 U11702 ( .A(n11768), .B(n11769), .Z(n11561) );
  XOR2_X1 U11703 ( .A(n11770), .B(n11771), .Z(n11769) );
  OR2_X1 U11704 ( .A1(n7636), .A2(n11328), .ZN(n11568) );
  XOR2_X1 U11705 ( .A(n11772), .B(n11773), .Z(n11565) );
  XOR2_X1 U11706 ( .A(n11774), .B(n11775), .Z(n11773) );
  OR2_X1 U11707 ( .A1(n7634), .A2(n11328), .ZN(n11572) );
  XOR2_X1 U11708 ( .A(n11776), .B(n11777), .Z(n11569) );
  XOR2_X1 U11709 ( .A(n11778), .B(n11779), .Z(n11777) );
  OR2_X1 U11710 ( .A1(n7632), .A2(n11328), .ZN(n11576) );
  XOR2_X1 U11711 ( .A(n11780), .B(n11781), .Z(n11573) );
  XOR2_X1 U11712 ( .A(n11782), .B(n11783), .Z(n11781) );
  OR2_X1 U11713 ( .A1(n8609), .A2(n11328), .ZN(n11580) );
  XOR2_X1 U11714 ( .A(n11784), .B(n11785), .Z(n11577) );
  XOR2_X1 U11715 ( .A(n11786), .B(n11787), .Z(n11785) );
  OR2_X1 U11716 ( .A1(n8614), .A2(n11328), .ZN(n11584) );
  XOR2_X1 U11717 ( .A(n11788), .B(n11789), .Z(n11581) );
  XOR2_X1 U11718 ( .A(n11790), .B(n11791), .Z(n11789) );
  OR2_X1 U11719 ( .A1(n8619), .A2(n11328), .ZN(n11588) );
  XOR2_X1 U11720 ( .A(n11792), .B(n11793), .Z(n11585) );
  XOR2_X1 U11721 ( .A(n11794), .B(n11795), .Z(n11793) );
  OR2_X1 U11722 ( .A1(n8624), .A2(n11328), .ZN(n11592) );
  XOR2_X1 U11723 ( .A(n11796), .B(n11797), .Z(n11589) );
  XOR2_X1 U11724 ( .A(n11798), .B(n11799), .Z(n11797) );
  OR2_X1 U11725 ( .A1(n8629), .A2(n11328), .ZN(n11596) );
  XOR2_X1 U11726 ( .A(n11800), .B(n11801), .Z(n11593) );
  XOR2_X1 U11727 ( .A(n11802), .B(n11803), .Z(n11801) );
  OR2_X1 U11728 ( .A1(n8634), .A2(n11328), .ZN(n11602) );
  XOR2_X1 U11729 ( .A(n11804), .B(n11805), .Z(n11599) );
  XOR2_X1 U11730 ( .A(n11806), .B(n11807), .Z(n11805) );
  OR2_X1 U11731 ( .A1(n8639), .A2(n11328), .ZN(n11606) );
  XOR2_X1 U11732 ( .A(n11808), .B(n11809), .Z(n11603) );
  XOR2_X1 U11733 ( .A(n11810), .B(n11811), .Z(n11809) );
  OR2_X1 U11734 ( .A1(n8644), .A2(n11328), .ZN(n10442) );
  XOR2_X1 U11735 ( .A(n11812), .B(n11813), .Z(n10439) );
  XOR2_X1 U11736 ( .A(n11814), .B(n11815), .Z(n11813) );
  OR2_X1 U11737 ( .A1(n8152), .A2(n11328), .ZN(n10403) );
  XNOR2_X1 U11738 ( .A(n11816), .B(n11817), .ZN(n10400) );
  XNOR2_X1 U11739 ( .A(n11818), .B(n11819), .ZN(n11816) );
  OR2_X1 U11740 ( .A1(n8105), .A2(n11328), .ZN(n8297) );
  XNOR2_X1 U11741 ( .A(n11820), .B(n11821), .ZN(n8294) );
  XNOR2_X1 U11742 ( .A(n11822), .B(n11823), .ZN(n11820) );
  OR2_X1 U11743 ( .A1(n8056), .A2(n11328), .ZN(n8260) );
  XNOR2_X1 U11744 ( .A(n11824), .B(n11825), .ZN(n8257) );
  XNOR2_X1 U11745 ( .A(n11826), .B(n11827), .ZN(n11824) );
  OR2_X1 U11746 ( .A1(n8023), .A2(n11328), .ZN(n8230) );
  XOR2_X1 U11747 ( .A(n11828), .B(n11829), .Z(n8228) );
  XOR2_X1 U11748 ( .A(n11830), .B(n11831), .Z(n11829) );
  OR2_X1 U11749 ( .A1(n11328), .A2(n7664), .ZN(n8207) );
  INV_X1 U11750 ( .A(n11323), .ZN(n11328) );
  XOR2_X1 U11751 ( .A(n11832), .B(n11833), .Z(n11323) );
  XNOR2_X1 U11752 ( .A(c_16_), .B(d_16_), .ZN(n11832) );
  XOR2_X1 U11753 ( .A(n11834), .B(n11835), .Z(n8205) );
  XOR2_X1 U11754 ( .A(n11836), .B(n11837), .Z(n11835) );
  XOR2_X1 U11755 ( .A(n11615), .B(n11838), .Z(n8191) );
  XOR2_X1 U11756 ( .A(n11614), .B(n11613), .Z(n11838) );
  OR2_X1 U11757 ( .A1(n11508), .A2(n7664), .ZN(n11613) );
  OR2_X1 U11758 ( .A1(n11839), .A2(n11840), .ZN(n11614) );
  AND2_X1 U11759 ( .A1(n11837), .A2(n11836), .ZN(n11840) );
  AND2_X1 U11760 ( .A1(n11834), .A2(n11841), .ZN(n11839) );
  OR2_X1 U11761 ( .A1(n11837), .A2(n11836), .ZN(n11841) );
  OR2_X1 U11762 ( .A1(n11842), .A2(n11843), .ZN(n11836) );
  AND2_X1 U11763 ( .A1(n11831), .A2(n11830), .ZN(n11843) );
  AND2_X1 U11764 ( .A1(n11828), .A2(n11844), .ZN(n11842) );
  OR2_X1 U11765 ( .A1(n11831), .A2(n11830), .ZN(n11844) );
  OR2_X1 U11766 ( .A1(n11845), .A2(n11846), .ZN(n11830) );
  AND2_X1 U11767 ( .A1(n11827), .A2(n11826), .ZN(n11846) );
  AND2_X1 U11768 ( .A1(n11825), .A2(n11847), .ZN(n11845) );
  OR2_X1 U11769 ( .A1(n11827), .A2(n11826), .ZN(n11847) );
  OR2_X1 U11770 ( .A1(n11848), .A2(n11849), .ZN(n11826) );
  AND2_X1 U11771 ( .A1(n11823), .A2(n11822), .ZN(n11849) );
  AND2_X1 U11772 ( .A1(n11821), .A2(n11850), .ZN(n11848) );
  OR2_X1 U11773 ( .A1(n11823), .A2(n11822), .ZN(n11850) );
  OR2_X1 U11774 ( .A1(n11851), .A2(n11852), .ZN(n11822) );
  AND2_X1 U11775 ( .A1(n11819), .A2(n11818), .ZN(n11852) );
  AND2_X1 U11776 ( .A1(n11817), .A2(n11853), .ZN(n11851) );
  OR2_X1 U11777 ( .A1(n11819), .A2(n11818), .ZN(n11853) );
  OR2_X1 U11778 ( .A1(n11854), .A2(n11855), .ZN(n11818) );
  AND2_X1 U11779 ( .A1(n11815), .A2(n11814), .ZN(n11855) );
  AND2_X1 U11780 ( .A1(n11812), .A2(n11856), .ZN(n11854) );
  OR2_X1 U11781 ( .A1(n11815), .A2(n11814), .ZN(n11856) );
  OR2_X1 U11782 ( .A1(n11857), .A2(n11858), .ZN(n11814) );
  AND2_X1 U11783 ( .A1(n11811), .A2(n11810), .ZN(n11858) );
  AND2_X1 U11784 ( .A1(n11808), .A2(n11859), .ZN(n11857) );
  OR2_X1 U11785 ( .A1(n11811), .A2(n11810), .ZN(n11859) );
  OR2_X1 U11786 ( .A1(n11860), .A2(n11861), .ZN(n11810) );
  AND2_X1 U11787 ( .A1(n11807), .A2(n11806), .ZN(n11861) );
  AND2_X1 U11788 ( .A1(n11804), .A2(n11862), .ZN(n11860) );
  OR2_X1 U11789 ( .A1(n11807), .A2(n11806), .ZN(n11862) );
  OR2_X1 U11790 ( .A1(n11863), .A2(n11864), .ZN(n11806) );
  AND2_X1 U11791 ( .A1(n11803), .A2(n11802), .ZN(n11864) );
  AND2_X1 U11792 ( .A1(n11800), .A2(n11865), .ZN(n11863) );
  OR2_X1 U11793 ( .A1(n11803), .A2(n11802), .ZN(n11865) );
  OR2_X1 U11794 ( .A1(n11866), .A2(n11867), .ZN(n11802) );
  AND2_X1 U11795 ( .A1(n11799), .A2(n11798), .ZN(n11867) );
  AND2_X1 U11796 ( .A1(n11796), .A2(n11868), .ZN(n11866) );
  OR2_X1 U11797 ( .A1(n11799), .A2(n11798), .ZN(n11868) );
  OR2_X1 U11798 ( .A1(n11869), .A2(n11870), .ZN(n11798) );
  AND2_X1 U11799 ( .A1(n11795), .A2(n11794), .ZN(n11870) );
  AND2_X1 U11800 ( .A1(n11792), .A2(n11871), .ZN(n11869) );
  OR2_X1 U11801 ( .A1(n11795), .A2(n11794), .ZN(n11871) );
  OR2_X1 U11802 ( .A1(n11872), .A2(n11873), .ZN(n11794) );
  AND2_X1 U11803 ( .A1(n11791), .A2(n11790), .ZN(n11873) );
  AND2_X1 U11804 ( .A1(n11788), .A2(n11874), .ZN(n11872) );
  OR2_X1 U11805 ( .A1(n11791), .A2(n11790), .ZN(n11874) );
  OR2_X1 U11806 ( .A1(n11875), .A2(n11876), .ZN(n11790) );
  AND2_X1 U11807 ( .A1(n11787), .A2(n11786), .ZN(n11876) );
  AND2_X1 U11808 ( .A1(n11784), .A2(n11877), .ZN(n11875) );
  OR2_X1 U11809 ( .A1(n11787), .A2(n11786), .ZN(n11877) );
  OR2_X1 U11810 ( .A1(n11878), .A2(n11879), .ZN(n11786) );
  AND2_X1 U11811 ( .A1(n11783), .A2(n11782), .ZN(n11879) );
  AND2_X1 U11812 ( .A1(n11780), .A2(n11880), .ZN(n11878) );
  OR2_X1 U11813 ( .A1(n11783), .A2(n11782), .ZN(n11880) );
  OR2_X1 U11814 ( .A1(n11881), .A2(n11882), .ZN(n11782) );
  AND2_X1 U11815 ( .A1(n11779), .A2(n11778), .ZN(n11882) );
  AND2_X1 U11816 ( .A1(n11776), .A2(n11883), .ZN(n11881) );
  OR2_X1 U11817 ( .A1(n11779), .A2(n11778), .ZN(n11883) );
  OR2_X1 U11818 ( .A1(n11884), .A2(n11885), .ZN(n11778) );
  AND2_X1 U11819 ( .A1(n11775), .A2(n11774), .ZN(n11885) );
  AND2_X1 U11820 ( .A1(n11772), .A2(n11886), .ZN(n11884) );
  OR2_X1 U11821 ( .A1(n11775), .A2(n11774), .ZN(n11886) );
  OR2_X1 U11822 ( .A1(n11887), .A2(n11888), .ZN(n11774) );
  AND2_X1 U11823 ( .A1(n11771), .A2(n11770), .ZN(n11888) );
  AND2_X1 U11824 ( .A1(n11768), .A2(n11889), .ZN(n11887) );
  OR2_X1 U11825 ( .A1(n11771), .A2(n11770), .ZN(n11889) );
  OR2_X1 U11826 ( .A1(n11890), .A2(n11891), .ZN(n11770) );
  AND2_X1 U11827 ( .A1(n11767), .A2(n11766), .ZN(n11891) );
  AND2_X1 U11828 ( .A1(n11764), .A2(n11892), .ZN(n11890) );
  OR2_X1 U11829 ( .A1(n11767), .A2(n11766), .ZN(n11892) );
  OR2_X1 U11830 ( .A1(n11893), .A2(n11894), .ZN(n11766) );
  AND2_X1 U11831 ( .A1(n11763), .A2(n11762), .ZN(n11894) );
  AND2_X1 U11832 ( .A1(n11760), .A2(n11895), .ZN(n11893) );
  OR2_X1 U11833 ( .A1(n11763), .A2(n11762), .ZN(n11895) );
  OR2_X1 U11834 ( .A1(n11896), .A2(n11897), .ZN(n11762) );
  AND2_X1 U11835 ( .A1(n11759), .A2(n11758), .ZN(n11897) );
  AND2_X1 U11836 ( .A1(n11756), .A2(n11898), .ZN(n11896) );
  OR2_X1 U11837 ( .A1(n11759), .A2(n11758), .ZN(n11898) );
  OR2_X1 U11838 ( .A1(n11899), .A2(n11900), .ZN(n11758) );
  AND2_X1 U11839 ( .A1(n11755), .A2(n11754), .ZN(n11900) );
  AND2_X1 U11840 ( .A1(n11752), .A2(n11901), .ZN(n11899) );
  OR2_X1 U11841 ( .A1(n11755), .A2(n11754), .ZN(n11901) );
  OR2_X1 U11842 ( .A1(n11902), .A2(n11903), .ZN(n11754) );
  AND2_X1 U11843 ( .A1(n11751), .A2(n11750), .ZN(n11903) );
  AND2_X1 U11844 ( .A1(n11748), .A2(n11904), .ZN(n11902) );
  OR2_X1 U11845 ( .A1(n11751), .A2(n11750), .ZN(n11904) );
  OR2_X1 U11846 ( .A1(n11905), .A2(n11906), .ZN(n11750) );
  AND2_X1 U11847 ( .A1(n11747), .A2(n11746), .ZN(n11906) );
  AND2_X1 U11848 ( .A1(n11744), .A2(n11907), .ZN(n11905) );
  OR2_X1 U11849 ( .A1(n11747), .A2(n11746), .ZN(n11907) );
  OR2_X1 U11850 ( .A1(n11908), .A2(n11909), .ZN(n11746) );
  AND2_X1 U11851 ( .A1(n11743), .A2(n11742), .ZN(n11909) );
  AND2_X1 U11852 ( .A1(n11740), .A2(n11910), .ZN(n11908) );
  OR2_X1 U11853 ( .A1(n11743), .A2(n11742), .ZN(n11910) );
  OR2_X1 U11854 ( .A1(n11911), .A2(n11912), .ZN(n11742) );
  AND2_X1 U11855 ( .A1(n11739), .A2(n11738), .ZN(n11912) );
  AND2_X1 U11856 ( .A1(n11736), .A2(n11913), .ZN(n11911) );
  OR2_X1 U11857 ( .A1(n11739), .A2(n11738), .ZN(n11913) );
  OR2_X1 U11858 ( .A1(n11914), .A2(n11915), .ZN(n11738) );
  AND2_X1 U11859 ( .A1(n11735), .A2(n11734), .ZN(n11915) );
  AND2_X1 U11860 ( .A1(n11732), .A2(n11916), .ZN(n11914) );
  OR2_X1 U11861 ( .A1(n11735), .A2(n11734), .ZN(n11916) );
  OR2_X1 U11862 ( .A1(n11917), .A2(n11918), .ZN(n11734) );
  AND2_X1 U11863 ( .A1(n11731), .A2(n11730), .ZN(n11918) );
  AND2_X1 U11864 ( .A1(n11728), .A2(n11919), .ZN(n11917) );
  OR2_X1 U11865 ( .A1(n11731), .A2(n11730), .ZN(n11919) );
  OR2_X1 U11866 ( .A1(n11920), .A2(n11921), .ZN(n11730) );
  AND2_X1 U11867 ( .A1(n11727), .A2(n11726), .ZN(n11921) );
  AND2_X1 U11868 ( .A1(n11724), .A2(n11922), .ZN(n11920) );
  OR2_X1 U11869 ( .A1(n11727), .A2(n11726), .ZN(n11922) );
  OR2_X1 U11870 ( .A1(n11923), .A2(n11924), .ZN(n11726) );
  AND2_X1 U11871 ( .A1(n11720), .A2(n11723), .ZN(n11924) );
  AND2_X1 U11872 ( .A1(n11722), .A2(n11925), .ZN(n11923) );
  OR2_X1 U11873 ( .A1(n11720), .A2(n11723), .ZN(n11925) );
  OR3_X1 U11874 ( .A1(n11719), .A2(n11508), .A3(n8519), .ZN(n11723) );
  OR2_X1 U11875 ( .A1(n11508), .A2(n7606), .ZN(n11720) );
  INV_X1 U11876 ( .A(n11926), .ZN(n11722) );
  OR2_X1 U11877 ( .A1(n11927), .A2(n11928), .ZN(n11926) );
  AND2_X1 U11878 ( .A1(n11929), .A2(n11930), .ZN(n11928) );
  OR2_X1 U11879 ( .A1(n11931), .A2(n7697), .ZN(n11930) );
  AND2_X1 U11880 ( .A1(n7691), .A2(n11719), .ZN(n11931) );
  AND2_X1 U11881 ( .A1(n11714), .A2(n11932), .ZN(n11927) );
  OR2_X1 U11882 ( .A1(n11933), .A2(n7701), .ZN(n11932) );
  AND2_X1 U11883 ( .A1(n11934), .A2(n7703), .ZN(n11933) );
  OR2_X1 U11884 ( .A1(n8529), .A2(n11508), .ZN(n11727) );
  XNOR2_X1 U11885 ( .A(n11935), .B(n11936), .ZN(n11724) );
  XNOR2_X1 U11886 ( .A(n11937), .B(n11938), .ZN(n11936) );
  OR2_X1 U11887 ( .A1(n8534), .A2(n11508), .ZN(n11731) );
  XOR2_X1 U11888 ( .A(n11939), .B(n11940), .Z(n11728) );
  XOR2_X1 U11889 ( .A(n11941), .B(n11942), .Z(n11940) );
  OR2_X1 U11890 ( .A1(n8539), .A2(n11508), .ZN(n11735) );
  XOR2_X1 U11891 ( .A(n11943), .B(n11944), .Z(n11732) );
  XOR2_X1 U11892 ( .A(n11945), .B(n11946), .Z(n11944) );
  OR2_X1 U11893 ( .A1(n8544), .A2(n11508), .ZN(n11739) );
  XOR2_X1 U11894 ( .A(n11947), .B(n11948), .Z(n11736) );
  XOR2_X1 U11895 ( .A(n11949), .B(n11950), .Z(n11948) );
  OR2_X1 U11896 ( .A1(n8549), .A2(n11508), .ZN(n11743) );
  XOR2_X1 U11897 ( .A(n11951), .B(n11952), .Z(n11740) );
  XOR2_X1 U11898 ( .A(n11953), .B(n11954), .Z(n11952) );
  OR2_X1 U11899 ( .A1(n8554), .A2(n11508), .ZN(n11747) );
  XOR2_X1 U11900 ( .A(n11955), .B(n11956), .Z(n11744) );
  XOR2_X1 U11901 ( .A(n11957), .B(n11958), .Z(n11956) );
  OR2_X1 U11902 ( .A1(n8559), .A2(n11508), .ZN(n11751) );
  XOR2_X1 U11903 ( .A(n11959), .B(n11960), .Z(n11748) );
  XOR2_X1 U11904 ( .A(n11961), .B(n11962), .Z(n11960) );
  OR2_X1 U11905 ( .A1(n8564), .A2(n11508), .ZN(n11755) );
  XOR2_X1 U11906 ( .A(n11963), .B(n11964), .Z(n11752) );
  XOR2_X1 U11907 ( .A(n11965), .B(n11966), .Z(n11964) );
  OR2_X1 U11908 ( .A1(n8569), .A2(n11508), .ZN(n11759) );
  XOR2_X1 U11909 ( .A(n11967), .B(n11968), .Z(n11756) );
  XOR2_X1 U11910 ( .A(n11969), .B(n11970), .Z(n11968) );
  OR2_X1 U11911 ( .A1(n8574), .A2(n11508), .ZN(n11763) );
  XOR2_X1 U11912 ( .A(n11971), .B(n11972), .Z(n11760) );
  XOR2_X1 U11913 ( .A(n11973), .B(n11974), .Z(n11972) );
  OR2_X1 U11914 ( .A1(n8579), .A2(n11508), .ZN(n11767) );
  XOR2_X1 U11915 ( .A(n11975), .B(n11976), .Z(n11764) );
  XOR2_X1 U11916 ( .A(n11977), .B(n11978), .Z(n11976) );
  OR2_X1 U11917 ( .A1(n8584), .A2(n11508), .ZN(n11771) );
  XOR2_X1 U11918 ( .A(n11979), .B(n11980), .Z(n11768) );
  XOR2_X1 U11919 ( .A(n11981), .B(n11982), .Z(n11980) );
  OR2_X1 U11920 ( .A1(n8589), .A2(n11508), .ZN(n11775) );
  XOR2_X1 U11921 ( .A(n11983), .B(n11984), .Z(n11772) );
  XOR2_X1 U11922 ( .A(n11985), .B(n11986), .Z(n11984) );
  OR2_X1 U11923 ( .A1(n8594), .A2(n11508), .ZN(n11779) );
  XOR2_X1 U11924 ( .A(n11987), .B(n11988), .Z(n11776) );
  XOR2_X1 U11925 ( .A(n11989), .B(n11990), .Z(n11988) );
  OR2_X1 U11926 ( .A1(n8599), .A2(n11508), .ZN(n11783) );
  XOR2_X1 U11927 ( .A(n11991), .B(n11992), .Z(n11780) );
  XOR2_X1 U11928 ( .A(n11993), .B(n11994), .Z(n11992) );
  OR2_X1 U11929 ( .A1(n8604), .A2(n11508), .ZN(n11787) );
  XOR2_X1 U11930 ( .A(n11995), .B(n11996), .Z(n11784) );
  XOR2_X1 U11931 ( .A(n11997), .B(n11998), .Z(n11996) );
  OR2_X1 U11932 ( .A1(n8609), .A2(n11508), .ZN(n11791) );
  XOR2_X1 U11933 ( .A(n11999), .B(n12000), .Z(n11788) );
  XOR2_X1 U11934 ( .A(n12001), .B(n12002), .Z(n12000) );
  OR2_X1 U11935 ( .A1(n8614), .A2(n11508), .ZN(n11795) );
  XOR2_X1 U11936 ( .A(n12003), .B(n12004), .Z(n11792) );
  XOR2_X1 U11937 ( .A(n12005), .B(n12006), .Z(n12004) );
  OR2_X1 U11938 ( .A1(n8619), .A2(n11508), .ZN(n11799) );
  XOR2_X1 U11939 ( .A(n12007), .B(n12008), .Z(n11796) );
  XOR2_X1 U11940 ( .A(n12009), .B(n12010), .Z(n12008) );
  OR2_X1 U11941 ( .A1(n8624), .A2(n11508), .ZN(n11803) );
  XOR2_X1 U11942 ( .A(n12011), .B(n12012), .Z(n11800) );
  XOR2_X1 U11943 ( .A(n12013), .B(n12014), .Z(n12012) );
  OR2_X1 U11944 ( .A1(n8629), .A2(n11508), .ZN(n11807) );
  XOR2_X1 U11945 ( .A(n12015), .B(n12016), .Z(n11804) );
  XOR2_X1 U11946 ( .A(n12017), .B(n12018), .Z(n12016) );
  OR2_X1 U11947 ( .A1(n8634), .A2(n11508), .ZN(n11811) );
  XOR2_X1 U11948 ( .A(n12019), .B(n12020), .Z(n11808) );
  XOR2_X1 U11949 ( .A(n12021), .B(n12022), .Z(n12020) );
  OR2_X1 U11950 ( .A1(n8639), .A2(n11508), .ZN(n11815) );
  XOR2_X1 U11951 ( .A(n12023), .B(n12024), .Z(n11812) );
  XOR2_X1 U11952 ( .A(n12025), .B(n12026), .Z(n12024) );
  OR2_X1 U11953 ( .A1(n8644), .A2(n11508), .ZN(n11819) );
  XNOR2_X1 U11954 ( .A(n12027), .B(n12028), .ZN(n11817) );
  XNOR2_X1 U11955 ( .A(n12029), .B(n12030), .ZN(n12027) );
  OR2_X1 U11956 ( .A1(n8152), .A2(n11508), .ZN(n11823) );
  XNOR2_X1 U11957 ( .A(n12031), .B(n12032), .ZN(n11821) );
  XNOR2_X1 U11958 ( .A(n12033), .B(n12034), .ZN(n12031) );
  OR2_X1 U11959 ( .A1(n8105), .A2(n11508), .ZN(n11827) );
  XNOR2_X1 U11960 ( .A(n12035), .B(n12036), .ZN(n11825) );
  XNOR2_X1 U11961 ( .A(n12037), .B(n12038), .ZN(n12035) );
  OR2_X1 U11962 ( .A1(n8056), .A2(n11508), .ZN(n11831) );
  XNOR2_X1 U11963 ( .A(n12039), .B(n12040), .ZN(n11828) );
  XNOR2_X1 U11964 ( .A(n12041), .B(n12042), .ZN(n12039) );
  OR2_X1 U11965 ( .A1(n8023), .A2(n11508), .ZN(n11837) );
  INV_X1 U11966 ( .A(n11503), .ZN(n11508) );
  XOR2_X1 U11967 ( .A(n12043), .B(n12044), .Z(n11503) );
  XNOR2_X1 U11968 ( .A(c_15_), .B(d_15_), .ZN(n12043) );
  XNOR2_X1 U11969 ( .A(n12045), .B(n12046), .ZN(n11834) );
  XNOR2_X1 U11970 ( .A(n12047), .B(n12048), .ZN(n12045) );
  XOR2_X1 U11971 ( .A(n12049), .B(n12050), .Z(n11615) );
  XOR2_X1 U11972 ( .A(n12051), .B(n12052), .Z(n12050) );
  AND2_X1 U11973 ( .A1(n12053), .A2(n8179), .ZN(n7939) );
  OR2_X1 U11974 ( .A1(n12054), .A2(n12055), .ZN(n8179) );
  INV_X1 U11975 ( .A(n12056), .ZN(n12053) );
  AND2_X1 U11976 ( .A1(n12054), .A2(n12055), .ZN(n12056) );
  OR2_X1 U11977 ( .A1(n12057), .A2(n12058), .ZN(n12055) );
  AND2_X1 U11978 ( .A1(n11620), .A2(n11619), .ZN(n12058) );
  AND2_X1 U11979 ( .A1(n11617), .A2(n12059), .ZN(n12057) );
  OR2_X1 U11980 ( .A1(n11619), .A2(n11620), .ZN(n12059) );
  OR2_X1 U11981 ( .A1(n11719), .A2(n7960), .ZN(n11620) );
  OR2_X1 U11982 ( .A1(n12060), .A2(n12061), .ZN(n11619) );
  AND2_X1 U11983 ( .A1(n12052), .A2(n12051), .ZN(n12061) );
  AND2_X1 U11984 ( .A1(n12049), .A2(n12062), .ZN(n12060) );
  OR2_X1 U11985 ( .A1(n12051), .A2(n12052), .ZN(n12062) );
  OR2_X1 U11986 ( .A1(n8023), .A2(n11719), .ZN(n12052) );
  OR2_X1 U11987 ( .A1(n12063), .A2(n12064), .ZN(n12051) );
  AND2_X1 U11988 ( .A1(n12048), .A2(n12047), .ZN(n12064) );
  AND2_X1 U11989 ( .A1(n12046), .A2(n12065), .ZN(n12063) );
  OR2_X1 U11990 ( .A1(n12047), .A2(n12048), .ZN(n12065) );
  OR2_X1 U11991 ( .A1(n8056), .A2(n11719), .ZN(n12048) );
  OR2_X1 U11992 ( .A1(n12066), .A2(n12067), .ZN(n12047) );
  AND2_X1 U11993 ( .A1(n12042), .A2(n12041), .ZN(n12067) );
  AND2_X1 U11994 ( .A1(n12040), .A2(n12068), .ZN(n12066) );
  OR2_X1 U11995 ( .A1(n12041), .A2(n12042), .ZN(n12068) );
  OR2_X1 U11996 ( .A1(n8105), .A2(n11719), .ZN(n12042) );
  OR2_X1 U11997 ( .A1(n12069), .A2(n12070), .ZN(n12041) );
  AND2_X1 U11998 ( .A1(n12038), .A2(n12037), .ZN(n12070) );
  AND2_X1 U11999 ( .A1(n12036), .A2(n12071), .ZN(n12069) );
  OR2_X1 U12000 ( .A1(n12037), .A2(n12038), .ZN(n12071) );
  OR2_X1 U12001 ( .A1(n8152), .A2(n11719), .ZN(n12038) );
  OR2_X1 U12002 ( .A1(n12072), .A2(n12073), .ZN(n12037) );
  AND2_X1 U12003 ( .A1(n12034), .A2(n12033), .ZN(n12073) );
  AND2_X1 U12004 ( .A1(n12032), .A2(n12074), .ZN(n12072) );
  OR2_X1 U12005 ( .A1(n12033), .A2(n12034), .ZN(n12074) );
  OR2_X1 U12006 ( .A1(n8644), .A2(n11719), .ZN(n12034) );
  OR2_X1 U12007 ( .A1(n12075), .A2(n12076), .ZN(n12033) );
  AND2_X1 U12008 ( .A1(n12030), .A2(n12029), .ZN(n12076) );
  AND2_X1 U12009 ( .A1(n12028), .A2(n12077), .ZN(n12075) );
  OR2_X1 U12010 ( .A1(n12029), .A2(n12030), .ZN(n12077) );
  OR2_X1 U12011 ( .A1(n8639), .A2(n11719), .ZN(n12030) );
  OR2_X1 U12012 ( .A1(n12078), .A2(n12079), .ZN(n12029) );
  AND2_X1 U12013 ( .A1(n12026), .A2(n12025), .ZN(n12079) );
  AND2_X1 U12014 ( .A1(n12023), .A2(n12080), .ZN(n12078) );
  OR2_X1 U12015 ( .A1(n12025), .A2(n12026), .ZN(n12080) );
  OR2_X1 U12016 ( .A1(n8634), .A2(n11719), .ZN(n12026) );
  OR2_X1 U12017 ( .A1(n12081), .A2(n12082), .ZN(n12025) );
  AND2_X1 U12018 ( .A1(n12022), .A2(n12021), .ZN(n12082) );
  AND2_X1 U12019 ( .A1(n12019), .A2(n12083), .ZN(n12081) );
  OR2_X1 U12020 ( .A1(n12021), .A2(n12022), .ZN(n12083) );
  OR2_X1 U12021 ( .A1(n8629), .A2(n11719), .ZN(n12022) );
  OR2_X1 U12022 ( .A1(n12084), .A2(n12085), .ZN(n12021) );
  AND2_X1 U12023 ( .A1(n12018), .A2(n12017), .ZN(n12085) );
  AND2_X1 U12024 ( .A1(n12015), .A2(n12086), .ZN(n12084) );
  OR2_X1 U12025 ( .A1(n12017), .A2(n12018), .ZN(n12086) );
  OR2_X1 U12026 ( .A1(n8624), .A2(n11719), .ZN(n12018) );
  OR2_X1 U12027 ( .A1(n12087), .A2(n12088), .ZN(n12017) );
  AND2_X1 U12028 ( .A1(n12014), .A2(n12013), .ZN(n12088) );
  AND2_X1 U12029 ( .A1(n12011), .A2(n12089), .ZN(n12087) );
  OR2_X1 U12030 ( .A1(n12013), .A2(n12014), .ZN(n12089) );
  OR2_X1 U12031 ( .A1(n8619), .A2(n11719), .ZN(n12014) );
  OR2_X1 U12032 ( .A1(n12090), .A2(n12091), .ZN(n12013) );
  AND2_X1 U12033 ( .A1(n12010), .A2(n12009), .ZN(n12091) );
  AND2_X1 U12034 ( .A1(n12007), .A2(n12092), .ZN(n12090) );
  OR2_X1 U12035 ( .A1(n12009), .A2(n12010), .ZN(n12092) );
  OR2_X1 U12036 ( .A1(n8614), .A2(n11719), .ZN(n12010) );
  OR2_X1 U12037 ( .A1(n12093), .A2(n12094), .ZN(n12009) );
  AND2_X1 U12038 ( .A1(n12006), .A2(n12005), .ZN(n12094) );
  AND2_X1 U12039 ( .A1(n12003), .A2(n12095), .ZN(n12093) );
  OR2_X1 U12040 ( .A1(n12005), .A2(n12006), .ZN(n12095) );
  OR2_X1 U12041 ( .A1(n8609), .A2(n11719), .ZN(n12006) );
  OR2_X1 U12042 ( .A1(n12096), .A2(n12097), .ZN(n12005) );
  AND2_X1 U12043 ( .A1(n12002), .A2(n12001), .ZN(n12097) );
  AND2_X1 U12044 ( .A1(n11999), .A2(n12098), .ZN(n12096) );
  OR2_X1 U12045 ( .A1(n12001), .A2(n12002), .ZN(n12098) );
  OR2_X1 U12046 ( .A1(n8604), .A2(n11719), .ZN(n12002) );
  OR2_X1 U12047 ( .A1(n12099), .A2(n12100), .ZN(n12001) );
  AND2_X1 U12048 ( .A1(n11998), .A2(n11997), .ZN(n12100) );
  AND2_X1 U12049 ( .A1(n11995), .A2(n12101), .ZN(n12099) );
  OR2_X1 U12050 ( .A1(n11997), .A2(n11998), .ZN(n12101) );
  OR2_X1 U12051 ( .A1(n8599), .A2(n11719), .ZN(n11998) );
  OR2_X1 U12052 ( .A1(n12102), .A2(n12103), .ZN(n11997) );
  AND2_X1 U12053 ( .A1(n11994), .A2(n11993), .ZN(n12103) );
  AND2_X1 U12054 ( .A1(n11991), .A2(n12104), .ZN(n12102) );
  OR2_X1 U12055 ( .A1(n11993), .A2(n11994), .ZN(n12104) );
  OR2_X1 U12056 ( .A1(n8594), .A2(n11719), .ZN(n11994) );
  OR2_X1 U12057 ( .A1(n12105), .A2(n12106), .ZN(n11993) );
  AND2_X1 U12058 ( .A1(n11990), .A2(n11989), .ZN(n12106) );
  AND2_X1 U12059 ( .A1(n11987), .A2(n12107), .ZN(n12105) );
  OR2_X1 U12060 ( .A1(n11989), .A2(n11990), .ZN(n12107) );
  OR2_X1 U12061 ( .A1(n8589), .A2(n11719), .ZN(n11990) );
  OR2_X1 U12062 ( .A1(n12108), .A2(n12109), .ZN(n11989) );
  AND2_X1 U12063 ( .A1(n11986), .A2(n11985), .ZN(n12109) );
  AND2_X1 U12064 ( .A1(n11983), .A2(n12110), .ZN(n12108) );
  OR2_X1 U12065 ( .A1(n11985), .A2(n11986), .ZN(n12110) );
  OR2_X1 U12066 ( .A1(n8584), .A2(n11719), .ZN(n11986) );
  OR2_X1 U12067 ( .A1(n12111), .A2(n12112), .ZN(n11985) );
  AND2_X1 U12068 ( .A1(n11982), .A2(n11981), .ZN(n12112) );
  AND2_X1 U12069 ( .A1(n11979), .A2(n12113), .ZN(n12111) );
  OR2_X1 U12070 ( .A1(n11981), .A2(n11982), .ZN(n12113) );
  OR2_X1 U12071 ( .A1(n8579), .A2(n11719), .ZN(n11982) );
  OR2_X1 U12072 ( .A1(n12114), .A2(n12115), .ZN(n11981) );
  AND2_X1 U12073 ( .A1(n11978), .A2(n11977), .ZN(n12115) );
  AND2_X1 U12074 ( .A1(n11975), .A2(n12116), .ZN(n12114) );
  OR2_X1 U12075 ( .A1(n11977), .A2(n11978), .ZN(n12116) );
  OR2_X1 U12076 ( .A1(n8574), .A2(n11719), .ZN(n11978) );
  OR2_X1 U12077 ( .A1(n12117), .A2(n12118), .ZN(n11977) );
  AND2_X1 U12078 ( .A1(n11974), .A2(n11973), .ZN(n12118) );
  AND2_X1 U12079 ( .A1(n11971), .A2(n12119), .ZN(n12117) );
  OR2_X1 U12080 ( .A1(n11973), .A2(n11974), .ZN(n12119) );
  OR2_X1 U12081 ( .A1(n8569), .A2(n11719), .ZN(n11974) );
  OR2_X1 U12082 ( .A1(n12120), .A2(n12121), .ZN(n11973) );
  AND2_X1 U12083 ( .A1(n11970), .A2(n11969), .ZN(n12121) );
  AND2_X1 U12084 ( .A1(n11967), .A2(n12122), .ZN(n12120) );
  OR2_X1 U12085 ( .A1(n11969), .A2(n11970), .ZN(n12122) );
  OR2_X1 U12086 ( .A1(n8564), .A2(n11719), .ZN(n11970) );
  OR2_X1 U12087 ( .A1(n12123), .A2(n12124), .ZN(n11969) );
  AND2_X1 U12088 ( .A1(n11966), .A2(n11965), .ZN(n12124) );
  AND2_X1 U12089 ( .A1(n11963), .A2(n12125), .ZN(n12123) );
  OR2_X1 U12090 ( .A1(n11965), .A2(n11966), .ZN(n12125) );
  OR2_X1 U12091 ( .A1(n8559), .A2(n11719), .ZN(n11966) );
  OR2_X1 U12092 ( .A1(n12126), .A2(n12127), .ZN(n11965) );
  AND2_X1 U12093 ( .A1(n11962), .A2(n11961), .ZN(n12127) );
  AND2_X1 U12094 ( .A1(n11959), .A2(n12128), .ZN(n12126) );
  OR2_X1 U12095 ( .A1(n11961), .A2(n11962), .ZN(n12128) );
  OR2_X1 U12096 ( .A1(n8554), .A2(n11719), .ZN(n11962) );
  OR2_X1 U12097 ( .A1(n12129), .A2(n12130), .ZN(n11961) );
  AND2_X1 U12098 ( .A1(n11958), .A2(n11957), .ZN(n12130) );
  AND2_X1 U12099 ( .A1(n11955), .A2(n12131), .ZN(n12129) );
  OR2_X1 U12100 ( .A1(n11957), .A2(n11958), .ZN(n12131) );
  OR2_X1 U12101 ( .A1(n8549), .A2(n11719), .ZN(n11958) );
  OR2_X1 U12102 ( .A1(n12132), .A2(n12133), .ZN(n11957) );
  AND2_X1 U12103 ( .A1(n11954), .A2(n11953), .ZN(n12133) );
  AND2_X1 U12104 ( .A1(n11951), .A2(n12134), .ZN(n12132) );
  OR2_X1 U12105 ( .A1(n11953), .A2(n11954), .ZN(n12134) );
  OR2_X1 U12106 ( .A1(n8544), .A2(n11719), .ZN(n11954) );
  OR2_X1 U12107 ( .A1(n12135), .A2(n12136), .ZN(n11953) );
  AND2_X1 U12108 ( .A1(n11950), .A2(n11949), .ZN(n12136) );
  AND2_X1 U12109 ( .A1(n11947), .A2(n12137), .ZN(n12135) );
  OR2_X1 U12110 ( .A1(n11949), .A2(n11950), .ZN(n12137) );
  OR2_X1 U12111 ( .A1(n8539), .A2(n11719), .ZN(n11950) );
  OR2_X1 U12112 ( .A1(n12138), .A2(n12139), .ZN(n11949) );
  AND2_X1 U12113 ( .A1(n11946), .A2(n11945), .ZN(n12139) );
  AND2_X1 U12114 ( .A1(n11943), .A2(n12140), .ZN(n12138) );
  OR2_X1 U12115 ( .A1(n11945), .A2(n11946), .ZN(n12140) );
  OR2_X1 U12116 ( .A1(n8534), .A2(n11719), .ZN(n11946) );
  OR2_X1 U12117 ( .A1(n12141), .A2(n12142), .ZN(n11945) );
  AND2_X1 U12118 ( .A1(n11942), .A2(n11941), .ZN(n12142) );
  AND2_X1 U12119 ( .A1(n11939), .A2(n12143), .ZN(n12141) );
  OR2_X1 U12120 ( .A1(n11941), .A2(n11942), .ZN(n12143) );
  OR2_X1 U12121 ( .A1(n8529), .A2(n11719), .ZN(n11942) );
  OR2_X1 U12122 ( .A1(n12144), .A2(n12145), .ZN(n11941) );
  AND2_X1 U12123 ( .A1(n11935), .A2(n11938), .ZN(n12145) );
  AND2_X1 U12124 ( .A1(n11937), .A2(n12146), .ZN(n12144) );
  OR2_X1 U12125 ( .A1(n11938), .A2(n11935), .ZN(n12146) );
  OR2_X1 U12126 ( .A1(n11719), .A2(n7606), .ZN(n11935) );
  OR3_X1 U12127 ( .A1(n11934), .A2(n11719), .A3(n8519), .ZN(n11938) );
  INV_X1 U12128 ( .A(n11714), .ZN(n11719) );
  XOR2_X1 U12129 ( .A(n12147), .B(n12148), .Z(n11714) );
  XNOR2_X1 U12130 ( .A(c_14_), .B(d_14_), .ZN(n12147) );
  INV_X1 U12131 ( .A(n12149), .ZN(n11937) );
  OR2_X1 U12132 ( .A1(n12150), .A2(n12151), .ZN(n12149) );
  AND2_X1 U12133 ( .A1(n12152), .A2(n12153), .ZN(n12151) );
  OR2_X1 U12134 ( .A1(n12154), .A2(n7697), .ZN(n12153) );
  AND2_X1 U12135 ( .A1(n7691), .A2(n11934), .ZN(n12154) );
  AND2_X1 U12136 ( .A1(n11929), .A2(n12155), .ZN(n12150) );
  OR2_X1 U12137 ( .A1(n12156), .A2(n7701), .ZN(n12155) );
  AND2_X1 U12138 ( .A1(n12157), .A2(n7703), .ZN(n12156) );
  XNOR2_X1 U12139 ( .A(n12158), .B(n12159), .ZN(n11939) );
  XNOR2_X1 U12140 ( .A(n12160), .B(n12161), .ZN(n12159) );
  XOR2_X1 U12141 ( .A(n12162), .B(n12163), .Z(n11943) );
  XOR2_X1 U12142 ( .A(n12164), .B(n12165), .Z(n12163) );
  XOR2_X1 U12143 ( .A(n12166), .B(n12167), .Z(n11947) );
  XOR2_X1 U12144 ( .A(n12168), .B(n12169), .Z(n12167) );
  XOR2_X1 U12145 ( .A(n12170), .B(n12171), .Z(n11951) );
  XOR2_X1 U12146 ( .A(n12172), .B(n12173), .Z(n12171) );
  XOR2_X1 U12147 ( .A(n12174), .B(n12175), .Z(n11955) );
  XOR2_X1 U12148 ( .A(n12176), .B(n12177), .Z(n12175) );
  XOR2_X1 U12149 ( .A(n12178), .B(n12179), .Z(n11959) );
  XOR2_X1 U12150 ( .A(n12180), .B(n12181), .Z(n12179) );
  XOR2_X1 U12151 ( .A(n12182), .B(n12183), .Z(n11963) );
  XOR2_X1 U12152 ( .A(n12184), .B(n12185), .Z(n12183) );
  XOR2_X1 U12153 ( .A(n12186), .B(n12187), .Z(n11967) );
  XOR2_X1 U12154 ( .A(n12188), .B(n12189), .Z(n12187) );
  XOR2_X1 U12155 ( .A(n12190), .B(n12191), .Z(n11971) );
  XOR2_X1 U12156 ( .A(n12192), .B(n12193), .Z(n12191) );
  XOR2_X1 U12157 ( .A(n12194), .B(n12195), .Z(n11975) );
  XOR2_X1 U12158 ( .A(n12196), .B(n12197), .Z(n12195) );
  XOR2_X1 U12159 ( .A(n12198), .B(n12199), .Z(n11979) );
  XOR2_X1 U12160 ( .A(n12200), .B(n12201), .Z(n12199) );
  XOR2_X1 U12161 ( .A(n12202), .B(n12203), .Z(n11983) );
  XOR2_X1 U12162 ( .A(n12204), .B(n12205), .Z(n12203) );
  XOR2_X1 U12163 ( .A(n12206), .B(n12207), .Z(n11987) );
  XOR2_X1 U12164 ( .A(n12208), .B(n12209), .Z(n12207) );
  XOR2_X1 U12165 ( .A(n12210), .B(n12211), .Z(n11991) );
  XOR2_X1 U12166 ( .A(n12212), .B(n12213), .Z(n12211) );
  XOR2_X1 U12167 ( .A(n12214), .B(n12215), .Z(n11995) );
  XOR2_X1 U12168 ( .A(n12216), .B(n12217), .Z(n12215) );
  XOR2_X1 U12169 ( .A(n12218), .B(n12219), .Z(n11999) );
  XOR2_X1 U12170 ( .A(n12220), .B(n12221), .Z(n12219) );
  XOR2_X1 U12171 ( .A(n12222), .B(n12223), .Z(n12003) );
  XOR2_X1 U12172 ( .A(n12224), .B(n12225), .Z(n12223) );
  XOR2_X1 U12173 ( .A(n12226), .B(n12227), .Z(n12007) );
  XOR2_X1 U12174 ( .A(n12228), .B(n12229), .Z(n12227) );
  XOR2_X1 U12175 ( .A(n12230), .B(n12231), .Z(n12011) );
  XOR2_X1 U12176 ( .A(n12232), .B(n12233), .Z(n12231) );
  XOR2_X1 U12177 ( .A(n12234), .B(n12235), .Z(n12015) );
  XOR2_X1 U12178 ( .A(n12236), .B(n12237), .Z(n12235) );
  XOR2_X1 U12179 ( .A(n12238), .B(n12239), .Z(n12019) );
  XOR2_X1 U12180 ( .A(n12240), .B(n12241), .Z(n12239) );
  XNOR2_X1 U12181 ( .A(n12242), .B(n12243), .ZN(n12023) );
  XNOR2_X1 U12182 ( .A(n12244), .B(n12245), .ZN(n12242) );
  XNOR2_X1 U12183 ( .A(n12246), .B(n12247), .ZN(n12028) );
  XNOR2_X1 U12184 ( .A(n12248), .B(n12249), .ZN(n12246) );
  XNOR2_X1 U12185 ( .A(n12250), .B(n12251), .ZN(n12032) );
  XNOR2_X1 U12186 ( .A(n12252), .B(n12253), .ZN(n12250) );
  XNOR2_X1 U12187 ( .A(n12254), .B(n12255), .ZN(n12036) );
  XNOR2_X1 U12188 ( .A(n12256), .B(n12257), .ZN(n12254) );
  XNOR2_X1 U12189 ( .A(n12258), .B(n12259), .ZN(n12040) );
  XNOR2_X1 U12190 ( .A(n12260), .B(n12261), .ZN(n12258) );
  XOR2_X1 U12191 ( .A(n12262), .B(n12263), .Z(n12046) );
  XOR2_X1 U12192 ( .A(n12264), .B(n12265), .Z(n12263) );
  XOR2_X1 U12193 ( .A(n12266), .B(n12267), .Z(n12049) );
  XOR2_X1 U12194 ( .A(n12268), .B(n12269), .Z(n12267) );
  XOR2_X1 U12195 ( .A(n12270), .B(n12271), .Z(n11617) );
  XOR2_X1 U12196 ( .A(n12272), .B(n12273), .Z(n12271) );
  XOR2_X1 U12197 ( .A(n12274), .B(n12275), .Z(n12054) );
  XOR2_X1 U12198 ( .A(n12276), .B(n12277), .Z(n12275) );
  INV_X1 U12199 ( .A(n7943), .ZN(n8178) );
  OR2_X1 U12200 ( .A1(n12278), .A2(n8175), .ZN(n7943) );
  INV_X1 U12201 ( .A(n7945), .ZN(n8175) );
  OR2_X1 U12202 ( .A1(n12279), .A2(n12280), .ZN(n7945) );
  AND2_X1 U12203 ( .A1(n12279), .A2(n12280), .ZN(n12278) );
  OR2_X1 U12204 ( .A1(n12281), .A2(n12282), .ZN(n12280) );
  AND2_X1 U12205 ( .A1(n12277), .A2(n12276), .ZN(n12282) );
  AND2_X1 U12206 ( .A1(n12274), .A2(n12283), .ZN(n12281) );
  OR2_X1 U12207 ( .A1(n12276), .A2(n12277), .ZN(n12283) );
  OR2_X1 U12208 ( .A1(n11934), .A2(n7960), .ZN(n12277) );
  OR2_X1 U12209 ( .A1(n12284), .A2(n12285), .ZN(n12276) );
  AND2_X1 U12210 ( .A1(n12273), .A2(n12272), .ZN(n12285) );
  AND2_X1 U12211 ( .A1(n12270), .A2(n12286), .ZN(n12284) );
  OR2_X1 U12212 ( .A1(n12272), .A2(n12273), .ZN(n12286) );
  OR2_X1 U12213 ( .A1(n11934), .A2(n7608), .ZN(n12273) );
  OR2_X1 U12214 ( .A1(n12287), .A2(n12288), .ZN(n12272) );
  AND2_X1 U12215 ( .A1(n12269), .A2(n12268), .ZN(n12288) );
  AND2_X1 U12216 ( .A1(n12266), .A2(n12289), .ZN(n12287) );
  OR2_X1 U12217 ( .A1(n12268), .A2(n12269), .ZN(n12289) );
  OR2_X1 U12218 ( .A1(n8056), .A2(n11934), .ZN(n12269) );
  OR2_X1 U12219 ( .A1(n12290), .A2(n12291), .ZN(n12268) );
  AND2_X1 U12220 ( .A1(n12265), .A2(n12264), .ZN(n12291) );
  AND2_X1 U12221 ( .A1(n12262), .A2(n12292), .ZN(n12290) );
  OR2_X1 U12222 ( .A1(n12264), .A2(n12265), .ZN(n12292) );
  OR2_X1 U12223 ( .A1(n8105), .A2(n11934), .ZN(n12265) );
  OR2_X1 U12224 ( .A1(n12293), .A2(n12294), .ZN(n12264) );
  AND2_X1 U12225 ( .A1(n12261), .A2(n12260), .ZN(n12294) );
  AND2_X1 U12226 ( .A1(n12259), .A2(n12295), .ZN(n12293) );
  OR2_X1 U12227 ( .A1(n12260), .A2(n12261), .ZN(n12295) );
  OR2_X1 U12228 ( .A1(n8152), .A2(n11934), .ZN(n12261) );
  OR2_X1 U12229 ( .A1(n12296), .A2(n12297), .ZN(n12260) );
  AND2_X1 U12230 ( .A1(n12257), .A2(n12256), .ZN(n12297) );
  AND2_X1 U12231 ( .A1(n12255), .A2(n12298), .ZN(n12296) );
  OR2_X1 U12232 ( .A1(n12256), .A2(n12257), .ZN(n12298) );
  OR2_X1 U12233 ( .A1(n8644), .A2(n11934), .ZN(n12257) );
  OR2_X1 U12234 ( .A1(n12299), .A2(n12300), .ZN(n12256) );
  AND2_X1 U12235 ( .A1(n12253), .A2(n12252), .ZN(n12300) );
  AND2_X1 U12236 ( .A1(n12251), .A2(n12301), .ZN(n12299) );
  OR2_X1 U12237 ( .A1(n12252), .A2(n12253), .ZN(n12301) );
  OR2_X1 U12238 ( .A1(n8639), .A2(n11934), .ZN(n12253) );
  OR2_X1 U12239 ( .A1(n12302), .A2(n12303), .ZN(n12252) );
  AND2_X1 U12240 ( .A1(n12249), .A2(n12248), .ZN(n12303) );
  AND2_X1 U12241 ( .A1(n12247), .A2(n12304), .ZN(n12302) );
  OR2_X1 U12242 ( .A1(n12248), .A2(n12249), .ZN(n12304) );
  OR2_X1 U12243 ( .A1(n8634), .A2(n11934), .ZN(n12249) );
  OR2_X1 U12244 ( .A1(n12305), .A2(n12306), .ZN(n12248) );
  AND2_X1 U12245 ( .A1(n12245), .A2(n12244), .ZN(n12306) );
  AND2_X1 U12246 ( .A1(n12243), .A2(n12307), .ZN(n12305) );
  OR2_X1 U12247 ( .A1(n12244), .A2(n12245), .ZN(n12307) );
  OR2_X1 U12248 ( .A1(n8629), .A2(n11934), .ZN(n12245) );
  OR2_X1 U12249 ( .A1(n12308), .A2(n12309), .ZN(n12244) );
  AND2_X1 U12250 ( .A1(n12241), .A2(n12240), .ZN(n12309) );
  AND2_X1 U12251 ( .A1(n12238), .A2(n12310), .ZN(n12308) );
  OR2_X1 U12252 ( .A1(n12240), .A2(n12241), .ZN(n12310) );
  OR2_X1 U12253 ( .A1(n8624), .A2(n11934), .ZN(n12241) );
  OR2_X1 U12254 ( .A1(n12311), .A2(n12312), .ZN(n12240) );
  AND2_X1 U12255 ( .A1(n12237), .A2(n12236), .ZN(n12312) );
  AND2_X1 U12256 ( .A1(n12234), .A2(n12313), .ZN(n12311) );
  OR2_X1 U12257 ( .A1(n12236), .A2(n12237), .ZN(n12313) );
  OR2_X1 U12258 ( .A1(n8619), .A2(n11934), .ZN(n12237) );
  OR2_X1 U12259 ( .A1(n12314), .A2(n12315), .ZN(n12236) );
  AND2_X1 U12260 ( .A1(n12233), .A2(n12232), .ZN(n12315) );
  AND2_X1 U12261 ( .A1(n12230), .A2(n12316), .ZN(n12314) );
  OR2_X1 U12262 ( .A1(n12232), .A2(n12233), .ZN(n12316) );
  OR2_X1 U12263 ( .A1(n8614), .A2(n11934), .ZN(n12233) );
  OR2_X1 U12264 ( .A1(n12317), .A2(n12318), .ZN(n12232) );
  AND2_X1 U12265 ( .A1(n12229), .A2(n12228), .ZN(n12318) );
  AND2_X1 U12266 ( .A1(n12226), .A2(n12319), .ZN(n12317) );
  OR2_X1 U12267 ( .A1(n12228), .A2(n12229), .ZN(n12319) );
  OR2_X1 U12268 ( .A1(n8609), .A2(n11934), .ZN(n12229) );
  OR2_X1 U12269 ( .A1(n12320), .A2(n12321), .ZN(n12228) );
  AND2_X1 U12270 ( .A1(n12225), .A2(n12224), .ZN(n12321) );
  AND2_X1 U12271 ( .A1(n12222), .A2(n12322), .ZN(n12320) );
  OR2_X1 U12272 ( .A1(n12224), .A2(n12225), .ZN(n12322) );
  OR2_X1 U12273 ( .A1(n8604), .A2(n11934), .ZN(n12225) );
  OR2_X1 U12274 ( .A1(n12323), .A2(n12324), .ZN(n12224) );
  AND2_X1 U12275 ( .A1(n12221), .A2(n12220), .ZN(n12324) );
  AND2_X1 U12276 ( .A1(n12218), .A2(n12325), .ZN(n12323) );
  OR2_X1 U12277 ( .A1(n12220), .A2(n12221), .ZN(n12325) );
  OR2_X1 U12278 ( .A1(n8599), .A2(n11934), .ZN(n12221) );
  OR2_X1 U12279 ( .A1(n12326), .A2(n12327), .ZN(n12220) );
  AND2_X1 U12280 ( .A1(n12217), .A2(n12216), .ZN(n12327) );
  AND2_X1 U12281 ( .A1(n12214), .A2(n12328), .ZN(n12326) );
  OR2_X1 U12282 ( .A1(n12216), .A2(n12217), .ZN(n12328) );
  OR2_X1 U12283 ( .A1(n8594), .A2(n11934), .ZN(n12217) );
  OR2_X1 U12284 ( .A1(n12329), .A2(n12330), .ZN(n12216) );
  AND2_X1 U12285 ( .A1(n12213), .A2(n12212), .ZN(n12330) );
  AND2_X1 U12286 ( .A1(n12210), .A2(n12331), .ZN(n12329) );
  OR2_X1 U12287 ( .A1(n12212), .A2(n12213), .ZN(n12331) );
  OR2_X1 U12288 ( .A1(n8589), .A2(n11934), .ZN(n12213) );
  OR2_X1 U12289 ( .A1(n12332), .A2(n12333), .ZN(n12212) );
  AND2_X1 U12290 ( .A1(n12209), .A2(n12208), .ZN(n12333) );
  AND2_X1 U12291 ( .A1(n12206), .A2(n12334), .ZN(n12332) );
  OR2_X1 U12292 ( .A1(n12208), .A2(n12209), .ZN(n12334) );
  OR2_X1 U12293 ( .A1(n8584), .A2(n11934), .ZN(n12209) );
  OR2_X1 U12294 ( .A1(n12335), .A2(n12336), .ZN(n12208) );
  AND2_X1 U12295 ( .A1(n12205), .A2(n12204), .ZN(n12336) );
  AND2_X1 U12296 ( .A1(n12202), .A2(n12337), .ZN(n12335) );
  OR2_X1 U12297 ( .A1(n12204), .A2(n12205), .ZN(n12337) );
  OR2_X1 U12298 ( .A1(n8579), .A2(n11934), .ZN(n12205) );
  OR2_X1 U12299 ( .A1(n12338), .A2(n12339), .ZN(n12204) );
  AND2_X1 U12300 ( .A1(n12201), .A2(n12200), .ZN(n12339) );
  AND2_X1 U12301 ( .A1(n12198), .A2(n12340), .ZN(n12338) );
  OR2_X1 U12302 ( .A1(n12200), .A2(n12201), .ZN(n12340) );
  OR2_X1 U12303 ( .A1(n8574), .A2(n11934), .ZN(n12201) );
  OR2_X1 U12304 ( .A1(n12341), .A2(n12342), .ZN(n12200) );
  AND2_X1 U12305 ( .A1(n12197), .A2(n12196), .ZN(n12342) );
  AND2_X1 U12306 ( .A1(n12194), .A2(n12343), .ZN(n12341) );
  OR2_X1 U12307 ( .A1(n12196), .A2(n12197), .ZN(n12343) );
  OR2_X1 U12308 ( .A1(n8569), .A2(n11934), .ZN(n12197) );
  OR2_X1 U12309 ( .A1(n12344), .A2(n12345), .ZN(n12196) );
  AND2_X1 U12310 ( .A1(n12193), .A2(n12192), .ZN(n12345) );
  AND2_X1 U12311 ( .A1(n12190), .A2(n12346), .ZN(n12344) );
  OR2_X1 U12312 ( .A1(n12192), .A2(n12193), .ZN(n12346) );
  OR2_X1 U12313 ( .A1(n8564), .A2(n11934), .ZN(n12193) );
  OR2_X1 U12314 ( .A1(n12347), .A2(n12348), .ZN(n12192) );
  AND2_X1 U12315 ( .A1(n12189), .A2(n12188), .ZN(n12348) );
  AND2_X1 U12316 ( .A1(n12186), .A2(n12349), .ZN(n12347) );
  OR2_X1 U12317 ( .A1(n12188), .A2(n12189), .ZN(n12349) );
  OR2_X1 U12318 ( .A1(n8559), .A2(n11934), .ZN(n12189) );
  OR2_X1 U12319 ( .A1(n12350), .A2(n12351), .ZN(n12188) );
  AND2_X1 U12320 ( .A1(n12185), .A2(n12184), .ZN(n12351) );
  AND2_X1 U12321 ( .A1(n12182), .A2(n12352), .ZN(n12350) );
  OR2_X1 U12322 ( .A1(n12184), .A2(n12185), .ZN(n12352) );
  OR2_X1 U12323 ( .A1(n8554), .A2(n11934), .ZN(n12185) );
  OR2_X1 U12324 ( .A1(n12353), .A2(n12354), .ZN(n12184) );
  AND2_X1 U12325 ( .A1(n12181), .A2(n12180), .ZN(n12354) );
  AND2_X1 U12326 ( .A1(n12178), .A2(n12355), .ZN(n12353) );
  OR2_X1 U12327 ( .A1(n12180), .A2(n12181), .ZN(n12355) );
  OR2_X1 U12328 ( .A1(n8549), .A2(n11934), .ZN(n12181) );
  OR2_X1 U12329 ( .A1(n12356), .A2(n12357), .ZN(n12180) );
  AND2_X1 U12330 ( .A1(n12177), .A2(n12176), .ZN(n12357) );
  AND2_X1 U12331 ( .A1(n12174), .A2(n12358), .ZN(n12356) );
  OR2_X1 U12332 ( .A1(n12176), .A2(n12177), .ZN(n12358) );
  OR2_X1 U12333 ( .A1(n8544), .A2(n11934), .ZN(n12177) );
  OR2_X1 U12334 ( .A1(n12359), .A2(n12360), .ZN(n12176) );
  AND2_X1 U12335 ( .A1(n12173), .A2(n12172), .ZN(n12360) );
  AND2_X1 U12336 ( .A1(n12170), .A2(n12361), .ZN(n12359) );
  OR2_X1 U12337 ( .A1(n12172), .A2(n12173), .ZN(n12361) );
  OR2_X1 U12338 ( .A1(n8539), .A2(n11934), .ZN(n12173) );
  OR2_X1 U12339 ( .A1(n12362), .A2(n12363), .ZN(n12172) );
  AND2_X1 U12340 ( .A1(n12169), .A2(n12168), .ZN(n12363) );
  AND2_X1 U12341 ( .A1(n12166), .A2(n12364), .ZN(n12362) );
  OR2_X1 U12342 ( .A1(n12168), .A2(n12169), .ZN(n12364) );
  OR2_X1 U12343 ( .A1(n8534), .A2(n11934), .ZN(n12169) );
  OR2_X1 U12344 ( .A1(n12365), .A2(n12366), .ZN(n12168) );
  AND2_X1 U12345 ( .A1(n12165), .A2(n12164), .ZN(n12366) );
  AND2_X1 U12346 ( .A1(n12162), .A2(n12367), .ZN(n12365) );
  OR2_X1 U12347 ( .A1(n12164), .A2(n12165), .ZN(n12367) );
  OR2_X1 U12348 ( .A1(n8529), .A2(n11934), .ZN(n12165) );
  OR2_X1 U12349 ( .A1(n12368), .A2(n12369), .ZN(n12164) );
  AND2_X1 U12350 ( .A1(n12158), .A2(n12161), .ZN(n12369) );
  AND2_X1 U12351 ( .A1(n12160), .A2(n12370), .ZN(n12368) );
  OR2_X1 U12352 ( .A1(n12161), .A2(n12158), .ZN(n12370) );
  OR2_X1 U12353 ( .A1(n11934), .A2(n7606), .ZN(n12158) );
  OR3_X1 U12354 ( .A1(n12157), .A2(n11934), .A3(n8519), .ZN(n12161) );
  INV_X1 U12355 ( .A(n11929), .ZN(n11934) );
  XOR2_X1 U12356 ( .A(n12371), .B(n12372), .Z(n11929) );
  XNOR2_X1 U12357 ( .A(c_13_), .B(d_13_), .ZN(n12371) );
  INV_X1 U12358 ( .A(n12373), .ZN(n12160) );
  OR2_X1 U12359 ( .A1(n12374), .A2(n12375), .ZN(n12373) );
  AND2_X1 U12360 ( .A1(n12376), .A2(n12377), .ZN(n12375) );
  OR2_X1 U12361 ( .A1(n12378), .A2(n7697), .ZN(n12377) );
  AND2_X1 U12362 ( .A1(n12157), .A2(n7691), .ZN(n12378) );
  AND2_X1 U12363 ( .A1(n12152), .A2(n12379), .ZN(n12374) );
  OR2_X1 U12364 ( .A1(n12380), .A2(n7701), .ZN(n12379) );
  AND2_X1 U12365 ( .A1(n12381), .A2(n7703), .ZN(n12380) );
  XNOR2_X1 U12366 ( .A(n12382), .B(n12383), .ZN(n12162) );
  XNOR2_X1 U12367 ( .A(n12384), .B(n12385), .ZN(n12383) );
  XOR2_X1 U12368 ( .A(n12386), .B(n12387), .Z(n12166) );
  XOR2_X1 U12369 ( .A(n12388), .B(n12389), .Z(n12387) );
  XOR2_X1 U12370 ( .A(n12390), .B(n12391), .Z(n12170) );
  XOR2_X1 U12371 ( .A(n12392), .B(n12393), .Z(n12391) );
  XOR2_X1 U12372 ( .A(n12394), .B(n12395), .Z(n12174) );
  XOR2_X1 U12373 ( .A(n12396), .B(n12397), .Z(n12395) );
  XOR2_X1 U12374 ( .A(n12398), .B(n12399), .Z(n12178) );
  XOR2_X1 U12375 ( .A(n12400), .B(n12401), .Z(n12399) );
  XOR2_X1 U12376 ( .A(n12402), .B(n12403), .Z(n12182) );
  XOR2_X1 U12377 ( .A(n12404), .B(n12405), .Z(n12403) );
  XOR2_X1 U12378 ( .A(n12406), .B(n12407), .Z(n12186) );
  XOR2_X1 U12379 ( .A(n12408), .B(n12409), .Z(n12407) );
  XOR2_X1 U12380 ( .A(n12410), .B(n12411), .Z(n12190) );
  XOR2_X1 U12381 ( .A(n12412), .B(n12413), .Z(n12411) );
  XOR2_X1 U12382 ( .A(n12414), .B(n12415), .Z(n12194) );
  XOR2_X1 U12383 ( .A(n12416), .B(n12417), .Z(n12415) );
  XOR2_X1 U12384 ( .A(n12418), .B(n12419), .Z(n12198) );
  XOR2_X1 U12385 ( .A(n12420), .B(n12421), .Z(n12419) );
  XOR2_X1 U12386 ( .A(n12422), .B(n12423), .Z(n12202) );
  XOR2_X1 U12387 ( .A(n12424), .B(n12425), .Z(n12423) );
  XOR2_X1 U12388 ( .A(n12426), .B(n12427), .Z(n12206) );
  XOR2_X1 U12389 ( .A(n12428), .B(n12429), .Z(n12427) );
  XOR2_X1 U12390 ( .A(n12430), .B(n12431), .Z(n12210) );
  XOR2_X1 U12391 ( .A(n12432), .B(n12433), .Z(n12431) );
  XOR2_X1 U12392 ( .A(n12434), .B(n12435), .Z(n12214) );
  XOR2_X1 U12393 ( .A(n12436), .B(n12437), .Z(n12435) );
  XOR2_X1 U12394 ( .A(n12438), .B(n12439), .Z(n12218) );
  XOR2_X1 U12395 ( .A(n12440), .B(n12441), .Z(n12439) );
  XOR2_X1 U12396 ( .A(n12442), .B(n12443), .Z(n12222) );
  XOR2_X1 U12397 ( .A(n12444), .B(n12445), .Z(n12443) );
  XOR2_X1 U12398 ( .A(n12446), .B(n12447), .Z(n12226) );
  XOR2_X1 U12399 ( .A(n12448), .B(n12449), .Z(n12447) );
  XOR2_X1 U12400 ( .A(n12450), .B(n12451), .Z(n12230) );
  XOR2_X1 U12401 ( .A(n12452), .B(n12453), .Z(n12451) );
  XOR2_X1 U12402 ( .A(n12454), .B(n12455), .Z(n12234) );
  XOR2_X1 U12403 ( .A(n12456), .B(n12457), .Z(n12455) );
  XNOR2_X1 U12404 ( .A(n12458), .B(n12459), .ZN(n12238) );
  XNOR2_X1 U12405 ( .A(n12460), .B(n12461), .ZN(n12458) );
  XNOR2_X1 U12406 ( .A(n12462), .B(n12463), .ZN(n12243) );
  XNOR2_X1 U12407 ( .A(n12464), .B(n12465), .ZN(n12462) );
  XNOR2_X1 U12408 ( .A(n12466), .B(n12467), .ZN(n12247) );
  XNOR2_X1 U12409 ( .A(n12468), .B(n12469), .ZN(n12466) );
  XNOR2_X1 U12410 ( .A(n12470), .B(n12471), .ZN(n12251) );
  XNOR2_X1 U12411 ( .A(n12472), .B(n12473), .ZN(n12470) );
  XOR2_X1 U12412 ( .A(n12474), .B(n12475), .Z(n12255) );
  XOR2_X1 U12413 ( .A(n12476), .B(n12477), .Z(n12475) );
  XOR2_X1 U12414 ( .A(n12478), .B(n12479), .Z(n12259) );
  XOR2_X1 U12415 ( .A(n12480), .B(n12481), .Z(n12479) );
  XOR2_X1 U12416 ( .A(n12482), .B(n12483), .Z(n12262) );
  XOR2_X1 U12417 ( .A(n12484), .B(n12485), .Z(n12483) );
  XOR2_X1 U12418 ( .A(n12486), .B(n12487), .Z(n12266) );
  XOR2_X1 U12419 ( .A(n12488), .B(n12489), .Z(n12487) );
  XOR2_X1 U12420 ( .A(n12490), .B(n12491), .Z(n12270) );
  XOR2_X1 U12421 ( .A(n12492), .B(n12493), .Z(n12491) );
  XOR2_X1 U12422 ( .A(n12494), .B(n12495), .Z(n12274) );
  XOR2_X1 U12423 ( .A(n12496), .B(n12497), .Z(n12495) );
  XOR2_X1 U12424 ( .A(n12498), .B(n12499), .Z(n12279) );
  XOR2_X1 U12425 ( .A(n12500), .B(n12501), .Z(n12499) );
  AND2_X1 U12426 ( .A1(n12502), .A2(n7949), .ZN(n7947) );
  OR2_X1 U12427 ( .A1(n12503), .A2(n12504), .ZN(n7949) );
  INV_X1 U12428 ( .A(n12505), .ZN(n12502) );
  AND2_X1 U12429 ( .A1(n12503), .A2(n12504), .ZN(n12505) );
  OR2_X1 U12430 ( .A1(n12506), .A2(n12507), .ZN(n12504) );
  AND2_X1 U12431 ( .A1(n12501), .A2(n12500), .ZN(n12507) );
  AND2_X1 U12432 ( .A1(n12498), .A2(n12508), .ZN(n12506) );
  OR2_X1 U12433 ( .A1(n12500), .A2(n12501), .ZN(n12508) );
  OR2_X1 U12434 ( .A1(n12157), .A2(n7960), .ZN(n12501) );
  OR2_X1 U12435 ( .A1(n12509), .A2(n12510), .ZN(n12500) );
  AND2_X1 U12436 ( .A1(n12497), .A2(n12496), .ZN(n12510) );
  AND2_X1 U12437 ( .A1(n12494), .A2(n12511), .ZN(n12509) );
  OR2_X1 U12438 ( .A1(n12496), .A2(n12497), .ZN(n12511) );
  OR2_X1 U12439 ( .A1(n12157), .A2(n7608), .ZN(n12497) );
  OR2_X1 U12440 ( .A1(n12512), .A2(n12513), .ZN(n12496) );
  AND2_X1 U12441 ( .A1(n12493), .A2(n12492), .ZN(n12513) );
  AND2_X1 U12442 ( .A1(n12490), .A2(n12514), .ZN(n12512) );
  OR2_X1 U12443 ( .A1(n12492), .A2(n12493), .ZN(n12514) );
  OR2_X1 U12444 ( .A1(n12157), .A2(n7610), .ZN(n12493) );
  OR2_X1 U12445 ( .A1(n12515), .A2(n12516), .ZN(n12492) );
  AND2_X1 U12446 ( .A1(n12489), .A2(n12488), .ZN(n12516) );
  AND2_X1 U12447 ( .A1(n12486), .A2(n12517), .ZN(n12515) );
  OR2_X1 U12448 ( .A1(n12488), .A2(n12489), .ZN(n12517) );
  OR2_X1 U12449 ( .A1(n8105), .A2(n12157), .ZN(n12489) );
  OR2_X1 U12450 ( .A1(n12518), .A2(n12519), .ZN(n12488) );
  AND2_X1 U12451 ( .A1(n12485), .A2(n12484), .ZN(n12519) );
  AND2_X1 U12452 ( .A1(n12482), .A2(n12520), .ZN(n12518) );
  OR2_X1 U12453 ( .A1(n12484), .A2(n12485), .ZN(n12520) );
  OR2_X1 U12454 ( .A1(n8152), .A2(n12157), .ZN(n12485) );
  OR2_X1 U12455 ( .A1(n12521), .A2(n12522), .ZN(n12484) );
  AND2_X1 U12456 ( .A1(n12481), .A2(n12480), .ZN(n12522) );
  AND2_X1 U12457 ( .A1(n12478), .A2(n12523), .ZN(n12521) );
  OR2_X1 U12458 ( .A1(n12480), .A2(n12481), .ZN(n12523) );
  OR2_X1 U12459 ( .A1(n8644), .A2(n12157), .ZN(n12481) );
  OR2_X1 U12460 ( .A1(n12524), .A2(n12525), .ZN(n12480) );
  AND2_X1 U12461 ( .A1(n12477), .A2(n12476), .ZN(n12525) );
  AND2_X1 U12462 ( .A1(n12474), .A2(n12526), .ZN(n12524) );
  OR2_X1 U12463 ( .A1(n12476), .A2(n12477), .ZN(n12526) );
  OR2_X1 U12464 ( .A1(n8639), .A2(n12157), .ZN(n12477) );
  OR2_X1 U12465 ( .A1(n12527), .A2(n12528), .ZN(n12476) );
  AND2_X1 U12466 ( .A1(n12473), .A2(n12472), .ZN(n12528) );
  AND2_X1 U12467 ( .A1(n12471), .A2(n12529), .ZN(n12527) );
  OR2_X1 U12468 ( .A1(n12472), .A2(n12473), .ZN(n12529) );
  OR2_X1 U12469 ( .A1(n8634), .A2(n12157), .ZN(n12473) );
  OR2_X1 U12470 ( .A1(n12530), .A2(n12531), .ZN(n12472) );
  AND2_X1 U12471 ( .A1(n12469), .A2(n12468), .ZN(n12531) );
  AND2_X1 U12472 ( .A1(n12467), .A2(n12532), .ZN(n12530) );
  OR2_X1 U12473 ( .A1(n12468), .A2(n12469), .ZN(n12532) );
  OR2_X1 U12474 ( .A1(n8629), .A2(n12157), .ZN(n12469) );
  OR2_X1 U12475 ( .A1(n12533), .A2(n12534), .ZN(n12468) );
  AND2_X1 U12476 ( .A1(n12465), .A2(n12464), .ZN(n12534) );
  AND2_X1 U12477 ( .A1(n12463), .A2(n12535), .ZN(n12533) );
  OR2_X1 U12478 ( .A1(n12464), .A2(n12465), .ZN(n12535) );
  OR2_X1 U12479 ( .A1(n8624), .A2(n12157), .ZN(n12465) );
  OR2_X1 U12480 ( .A1(n12536), .A2(n12537), .ZN(n12464) );
  AND2_X1 U12481 ( .A1(n12461), .A2(n12460), .ZN(n12537) );
  AND2_X1 U12482 ( .A1(n12459), .A2(n12538), .ZN(n12536) );
  OR2_X1 U12483 ( .A1(n12460), .A2(n12461), .ZN(n12538) );
  OR2_X1 U12484 ( .A1(n8619), .A2(n12157), .ZN(n12461) );
  OR2_X1 U12485 ( .A1(n12539), .A2(n12540), .ZN(n12460) );
  AND2_X1 U12486 ( .A1(n12457), .A2(n12456), .ZN(n12540) );
  AND2_X1 U12487 ( .A1(n12454), .A2(n12541), .ZN(n12539) );
  OR2_X1 U12488 ( .A1(n12456), .A2(n12457), .ZN(n12541) );
  OR2_X1 U12489 ( .A1(n8614), .A2(n12157), .ZN(n12457) );
  OR2_X1 U12490 ( .A1(n12542), .A2(n12543), .ZN(n12456) );
  AND2_X1 U12491 ( .A1(n12453), .A2(n12452), .ZN(n12543) );
  AND2_X1 U12492 ( .A1(n12450), .A2(n12544), .ZN(n12542) );
  OR2_X1 U12493 ( .A1(n12452), .A2(n12453), .ZN(n12544) );
  OR2_X1 U12494 ( .A1(n8609), .A2(n12157), .ZN(n12453) );
  OR2_X1 U12495 ( .A1(n12545), .A2(n12546), .ZN(n12452) );
  AND2_X1 U12496 ( .A1(n12449), .A2(n12448), .ZN(n12546) );
  AND2_X1 U12497 ( .A1(n12446), .A2(n12547), .ZN(n12545) );
  OR2_X1 U12498 ( .A1(n12448), .A2(n12449), .ZN(n12547) );
  OR2_X1 U12499 ( .A1(n8604), .A2(n12157), .ZN(n12449) );
  OR2_X1 U12500 ( .A1(n12548), .A2(n12549), .ZN(n12448) );
  AND2_X1 U12501 ( .A1(n12445), .A2(n12444), .ZN(n12549) );
  AND2_X1 U12502 ( .A1(n12442), .A2(n12550), .ZN(n12548) );
  OR2_X1 U12503 ( .A1(n12444), .A2(n12445), .ZN(n12550) );
  OR2_X1 U12504 ( .A1(n8599), .A2(n12157), .ZN(n12445) );
  OR2_X1 U12505 ( .A1(n12551), .A2(n12552), .ZN(n12444) );
  AND2_X1 U12506 ( .A1(n12441), .A2(n12440), .ZN(n12552) );
  AND2_X1 U12507 ( .A1(n12438), .A2(n12553), .ZN(n12551) );
  OR2_X1 U12508 ( .A1(n12440), .A2(n12441), .ZN(n12553) );
  OR2_X1 U12509 ( .A1(n8594), .A2(n12157), .ZN(n12441) );
  OR2_X1 U12510 ( .A1(n12554), .A2(n12555), .ZN(n12440) );
  AND2_X1 U12511 ( .A1(n12437), .A2(n12436), .ZN(n12555) );
  AND2_X1 U12512 ( .A1(n12434), .A2(n12556), .ZN(n12554) );
  OR2_X1 U12513 ( .A1(n12436), .A2(n12437), .ZN(n12556) );
  OR2_X1 U12514 ( .A1(n8589), .A2(n12157), .ZN(n12437) );
  OR2_X1 U12515 ( .A1(n12557), .A2(n12558), .ZN(n12436) );
  AND2_X1 U12516 ( .A1(n12433), .A2(n12432), .ZN(n12558) );
  AND2_X1 U12517 ( .A1(n12430), .A2(n12559), .ZN(n12557) );
  OR2_X1 U12518 ( .A1(n12432), .A2(n12433), .ZN(n12559) );
  OR2_X1 U12519 ( .A1(n8584), .A2(n12157), .ZN(n12433) );
  OR2_X1 U12520 ( .A1(n12560), .A2(n12561), .ZN(n12432) );
  AND2_X1 U12521 ( .A1(n12429), .A2(n12428), .ZN(n12561) );
  AND2_X1 U12522 ( .A1(n12426), .A2(n12562), .ZN(n12560) );
  OR2_X1 U12523 ( .A1(n12428), .A2(n12429), .ZN(n12562) );
  OR2_X1 U12524 ( .A1(n8579), .A2(n12157), .ZN(n12429) );
  OR2_X1 U12525 ( .A1(n12563), .A2(n12564), .ZN(n12428) );
  AND2_X1 U12526 ( .A1(n12425), .A2(n12424), .ZN(n12564) );
  AND2_X1 U12527 ( .A1(n12422), .A2(n12565), .ZN(n12563) );
  OR2_X1 U12528 ( .A1(n12424), .A2(n12425), .ZN(n12565) );
  OR2_X1 U12529 ( .A1(n8574), .A2(n12157), .ZN(n12425) );
  OR2_X1 U12530 ( .A1(n12566), .A2(n12567), .ZN(n12424) );
  AND2_X1 U12531 ( .A1(n12421), .A2(n12420), .ZN(n12567) );
  AND2_X1 U12532 ( .A1(n12418), .A2(n12568), .ZN(n12566) );
  OR2_X1 U12533 ( .A1(n12420), .A2(n12421), .ZN(n12568) );
  OR2_X1 U12534 ( .A1(n8569), .A2(n12157), .ZN(n12421) );
  OR2_X1 U12535 ( .A1(n12569), .A2(n12570), .ZN(n12420) );
  AND2_X1 U12536 ( .A1(n12417), .A2(n12416), .ZN(n12570) );
  AND2_X1 U12537 ( .A1(n12414), .A2(n12571), .ZN(n12569) );
  OR2_X1 U12538 ( .A1(n12416), .A2(n12417), .ZN(n12571) );
  OR2_X1 U12539 ( .A1(n8564), .A2(n12157), .ZN(n12417) );
  OR2_X1 U12540 ( .A1(n12572), .A2(n12573), .ZN(n12416) );
  AND2_X1 U12541 ( .A1(n12413), .A2(n12412), .ZN(n12573) );
  AND2_X1 U12542 ( .A1(n12410), .A2(n12574), .ZN(n12572) );
  OR2_X1 U12543 ( .A1(n12412), .A2(n12413), .ZN(n12574) );
  OR2_X1 U12544 ( .A1(n8559), .A2(n12157), .ZN(n12413) );
  OR2_X1 U12545 ( .A1(n12575), .A2(n12576), .ZN(n12412) );
  AND2_X1 U12546 ( .A1(n12409), .A2(n12408), .ZN(n12576) );
  AND2_X1 U12547 ( .A1(n12406), .A2(n12577), .ZN(n12575) );
  OR2_X1 U12548 ( .A1(n12408), .A2(n12409), .ZN(n12577) );
  OR2_X1 U12549 ( .A1(n8554), .A2(n12157), .ZN(n12409) );
  OR2_X1 U12550 ( .A1(n12578), .A2(n12579), .ZN(n12408) );
  AND2_X1 U12551 ( .A1(n12405), .A2(n12404), .ZN(n12579) );
  AND2_X1 U12552 ( .A1(n12402), .A2(n12580), .ZN(n12578) );
  OR2_X1 U12553 ( .A1(n12404), .A2(n12405), .ZN(n12580) );
  OR2_X1 U12554 ( .A1(n8549), .A2(n12157), .ZN(n12405) );
  OR2_X1 U12555 ( .A1(n12581), .A2(n12582), .ZN(n12404) );
  AND2_X1 U12556 ( .A1(n12401), .A2(n12400), .ZN(n12582) );
  AND2_X1 U12557 ( .A1(n12398), .A2(n12583), .ZN(n12581) );
  OR2_X1 U12558 ( .A1(n12400), .A2(n12401), .ZN(n12583) );
  OR2_X1 U12559 ( .A1(n8544), .A2(n12157), .ZN(n12401) );
  OR2_X1 U12560 ( .A1(n12584), .A2(n12585), .ZN(n12400) );
  AND2_X1 U12561 ( .A1(n12397), .A2(n12396), .ZN(n12585) );
  AND2_X1 U12562 ( .A1(n12394), .A2(n12586), .ZN(n12584) );
  OR2_X1 U12563 ( .A1(n12396), .A2(n12397), .ZN(n12586) );
  OR2_X1 U12564 ( .A1(n8539), .A2(n12157), .ZN(n12397) );
  OR2_X1 U12565 ( .A1(n12587), .A2(n12588), .ZN(n12396) );
  AND2_X1 U12566 ( .A1(n12393), .A2(n12392), .ZN(n12588) );
  AND2_X1 U12567 ( .A1(n12390), .A2(n12589), .ZN(n12587) );
  OR2_X1 U12568 ( .A1(n12392), .A2(n12393), .ZN(n12589) );
  OR2_X1 U12569 ( .A1(n8534), .A2(n12157), .ZN(n12393) );
  OR2_X1 U12570 ( .A1(n12590), .A2(n12591), .ZN(n12392) );
  AND2_X1 U12571 ( .A1(n12389), .A2(n12388), .ZN(n12591) );
  AND2_X1 U12572 ( .A1(n12386), .A2(n12592), .ZN(n12590) );
  OR2_X1 U12573 ( .A1(n12388), .A2(n12389), .ZN(n12592) );
  OR2_X1 U12574 ( .A1(n8529), .A2(n12157), .ZN(n12389) );
  OR2_X1 U12575 ( .A1(n12593), .A2(n12594), .ZN(n12388) );
  AND2_X1 U12576 ( .A1(n12382), .A2(n12385), .ZN(n12594) );
  AND2_X1 U12577 ( .A1(n12384), .A2(n12595), .ZN(n12593) );
  OR2_X1 U12578 ( .A1(n12385), .A2(n12382), .ZN(n12595) );
  OR2_X1 U12579 ( .A1(n12157), .A2(n8518), .ZN(n12382) );
  OR3_X1 U12580 ( .A1(n12381), .A2(n12157), .A3(n8519), .ZN(n12385) );
  INV_X1 U12581 ( .A(n12152), .ZN(n12157) );
  XOR2_X1 U12582 ( .A(n12596), .B(n12597), .Z(n12152) );
  XNOR2_X1 U12583 ( .A(c_12_), .B(d_12_), .ZN(n12596) );
  INV_X1 U12584 ( .A(n12598), .ZN(n12384) );
  OR2_X1 U12585 ( .A1(n12599), .A2(n12600), .ZN(n12598) );
  AND2_X1 U12586 ( .A1(n12601), .A2(n12602), .ZN(n12600) );
  OR2_X1 U12587 ( .A1(n12603), .A2(n7697), .ZN(n12602) );
  AND2_X1 U12588 ( .A1(n12381), .A2(n7691), .ZN(n12603) );
  AND2_X1 U12589 ( .A1(n12376), .A2(n12604), .ZN(n12599) );
  OR2_X1 U12590 ( .A1(n12605), .A2(n7701), .ZN(n12604) );
  AND2_X1 U12591 ( .A1(n12606), .A2(n7703), .ZN(n12605) );
  XNOR2_X1 U12592 ( .A(n12607), .B(n12608), .ZN(n12386) );
  XNOR2_X1 U12593 ( .A(n12609), .B(n12610), .ZN(n12608) );
  XOR2_X1 U12594 ( .A(n12611), .B(n12612), .Z(n12390) );
  XOR2_X1 U12595 ( .A(n12613), .B(n12614), .Z(n12612) );
  XOR2_X1 U12596 ( .A(n12615), .B(n12616), .Z(n12394) );
  XOR2_X1 U12597 ( .A(n12617), .B(n12618), .Z(n12616) );
  XOR2_X1 U12598 ( .A(n12619), .B(n12620), .Z(n12398) );
  XOR2_X1 U12599 ( .A(n12621), .B(n12622), .Z(n12620) );
  XOR2_X1 U12600 ( .A(n12623), .B(n12624), .Z(n12402) );
  XOR2_X1 U12601 ( .A(n12625), .B(n12626), .Z(n12624) );
  XOR2_X1 U12602 ( .A(n12627), .B(n12628), .Z(n12406) );
  XOR2_X1 U12603 ( .A(n12629), .B(n12630), .Z(n12628) );
  XOR2_X1 U12604 ( .A(n12631), .B(n12632), .Z(n12410) );
  XOR2_X1 U12605 ( .A(n12633), .B(n12634), .Z(n12632) );
  XOR2_X1 U12606 ( .A(n12635), .B(n12636), .Z(n12414) );
  XOR2_X1 U12607 ( .A(n12637), .B(n12638), .Z(n12636) );
  XOR2_X1 U12608 ( .A(n12639), .B(n12640), .Z(n12418) );
  XOR2_X1 U12609 ( .A(n12641), .B(n12642), .Z(n12640) );
  XOR2_X1 U12610 ( .A(n12643), .B(n12644), .Z(n12422) );
  XOR2_X1 U12611 ( .A(n12645), .B(n12646), .Z(n12644) );
  XOR2_X1 U12612 ( .A(n12647), .B(n12648), .Z(n12426) );
  XOR2_X1 U12613 ( .A(n12649), .B(n12650), .Z(n12648) );
  XOR2_X1 U12614 ( .A(n12651), .B(n12652), .Z(n12430) );
  XOR2_X1 U12615 ( .A(n12653), .B(n12654), .Z(n12652) );
  XOR2_X1 U12616 ( .A(n12655), .B(n12656), .Z(n12434) );
  XOR2_X1 U12617 ( .A(n12657), .B(n12658), .Z(n12656) );
  XOR2_X1 U12618 ( .A(n12659), .B(n12660), .Z(n12438) );
  XOR2_X1 U12619 ( .A(n12661), .B(n12662), .Z(n12660) );
  XOR2_X1 U12620 ( .A(n12663), .B(n12664), .Z(n12442) );
  XOR2_X1 U12621 ( .A(n12665), .B(n12666), .Z(n12664) );
  XOR2_X1 U12622 ( .A(n12667), .B(n12668), .Z(n12446) );
  XOR2_X1 U12623 ( .A(n12669), .B(n12670), .Z(n12668) );
  XOR2_X1 U12624 ( .A(n12671), .B(n12672), .Z(n12450) );
  XOR2_X1 U12625 ( .A(n12673), .B(n12674), .Z(n12672) );
  XNOR2_X1 U12626 ( .A(n12675), .B(n12676), .ZN(n12454) );
  XNOR2_X1 U12627 ( .A(n12677), .B(n12678), .ZN(n12675) );
  XNOR2_X1 U12628 ( .A(n12679), .B(n12680), .ZN(n12459) );
  XNOR2_X1 U12629 ( .A(n12681), .B(n12682), .ZN(n12679) );
  XNOR2_X1 U12630 ( .A(n12683), .B(n12684), .ZN(n12463) );
  XNOR2_X1 U12631 ( .A(n12685), .B(n12686), .ZN(n12683) );
  XNOR2_X1 U12632 ( .A(n12687), .B(n12688), .ZN(n12467) );
  XNOR2_X1 U12633 ( .A(n12689), .B(n12690), .ZN(n12687) );
  XOR2_X1 U12634 ( .A(n12691), .B(n12692), .Z(n12471) );
  XOR2_X1 U12635 ( .A(n12693), .B(n12694), .Z(n12692) );
  XOR2_X1 U12636 ( .A(n12695), .B(n12696), .Z(n12474) );
  XOR2_X1 U12637 ( .A(n12697), .B(n12698), .Z(n12696) );
  XOR2_X1 U12638 ( .A(n12699), .B(n12700), .Z(n12478) );
  XOR2_X1 U12639 ( .A(n12701), .B(n12702), .Z(n12700) );
  XOR2_X1 U12640 ( .A(n12703), .B(n12704), .Z(n12482) );
  XOR2_X1 U12641 ( .A(n12705), .B(n12706), .Z(n12704) );
  XOR2_X1 U12642 ( .A(n12707), .B(n12708), .Z(n12486) );
  XOR2_X1 U12643 ( .A(n12709), .B(n12710), .Z(n12708) );
  XOR2_X1 U12644 ( .A(n12711), .B(n12712), .Z(n12490) );
  XOR2_X1 U12645 ( .A(n12713), .B(n12714), .Z(n12712) );
  XOR2_X1 U12646 ( .A(n12715), .B(n12716), .Z(n12494) );
  XOR2_X1 U12647 ( .A(n12717), .B(n12718), .Z(n12716) );
  XOR2_X1 U12648 ( .A(n12719), .B(n12720), .Z(n12498) );
  XOR2_X1 U12649 ( .A(n12721), .B(n12722), .Z(n12720) );
  XOR2_X1 U12650 ( .A(n12723), .B(n12724), .Z(n12503) );
  XOR2_X1 U12651 ( .A(n12725), .B(n12726), .Z(n12724) );
  AND2_X1 U12652 ( .A1(n12727), .A2(n8169), .ZN(n7951) );
  OR2_X1 U12653 ( .A1(n12728), .A2(n12729), .ZN(n8169) );
  INV_X1 U12654 ( .A(n12730), .ZN(n12727) );
  AND2_X1 U12655 ( .A1(n12728), .A2(n12729), .ZN(n12730) );
  OR2_X1 U12656 ( .A1(n12731), .A2(n12732), .ZN(n12729) );
  AND2_X1 U12657 ( .A1(n12726), .A2(n12725), .ZN(n12732) );
  AND2_X1 U12658 ( .A1(n12723), .A2(n12733), .ZN(n12731) );
  OR2_X1 U12659 ( .A1(n12725), .A2(n12726), .ZN(n12733) );
  OR2_X1 U12660 ( .A1(n12381), .A2(n7960), .ZN(n12726) );
  OR2_X1 U12661 ( .A1(n12734), .A2(n12735), .ZN(n12725) );
  AND2_X1 U12662 ( .A1(n12722), .A2(n12721), .ZN(n12735) );
  AND2_X1 U12663 ( .A1(n12719), .A2(n12736), .ZN(n12734) );
  OR2_X1 U12664 ( .A1(n12721), .A2(n12722), .ZN(n12736) );
  OR2_X1 U12665 ( .A1(n12381), .A2(n7608), .ZN(n12722) );
  OR2_X1 U12666 ( .A1(n12737), .A2(n12738), .ZN(n12721) );
  AND2_X1 U12667 ( .A1(n12718), .A2(n12717), .ZN(n12738) );
  AND2_X1 U12668 ( .A1(n12715), .A2(n12739), .ZN(n12737) );
  OR2_X1 U12669 ( .A1(n12717), .A2(n12718), .ZN(n12739) );
  OR2_X1 U12670 ( .A1(n12381), .A2(n7610), .ZN(n12718) );
  OR2_X1 U12671 ( .A1(n12740), .A2(n12741), .ZN(n12717) );
  AND2_X1 U12672 ( .A1(n12714), .A2(n12713), .ZN(n12741) );
  AND2_X1 U12673 ( .A1(n12711), .A2(n12742), .ZN(n12740) );
  OR2_X1 U12674 ( .A1(n12713), .A2(n12714), .ZN(n12742) );
  OR2_X1 U12675 ( .A1(n12381), .A2(n7612), .ZN(n12714) );
  OR2_X1 U12676 ( .A1(n12743), .A2(n12744), .ZN(n12713) );
  AND2_X1 U12677 ( .A1(n12710), .A2(n12709), .ZN(n12744) );
  AND2_X1 U12678 ( .A1(n12707), .A2(n12745), .ZN(n12743) );
  OR2_X1 U12679 ( .A1(n12709), .A2(n12710), .ZN(n12745) );
  OR2_X1 U12680 ( .A1(n8152), .A2(n12381), .ZN(n12710) );
  OR2_X1 U12681 ( .A1(n12746), .A2(n12747), .ZN(n12709) );
  AND2_X1 U12682 ( .A1(n12706), .A2(n12705), .ZN(n12747) );
  AND2_X1 U12683 ( .A1(n12703), .A2(n12748), .ZN(n12746) );
  OR2_X1 U12684 ( .A1(n12705), .A2(n12706), .ZN(n12748) );
  OR2_X1 U12685 ( .A1(n8644), .A2(n12381), .ZN(n12706) );
  OR2_X1 U12686 ( .A1(n12749), .A2(n12750), .ZN(n12705) );
  AND2_X1 U12687 ( .A1(n12702), .A2(n12701), .ZN(n12750) );
  AND2_X1 U12688 ( .A1(n12699), .A2(n12751), .ZN(n12749) );
  OR2_X1 U12689 ( .A1(n12701), .A2(n12702), .ZN(n12751) );
  OR2_X1 U12690 ( .A1(n8639), .A2(n12381), .ZN(n12702) );
  OR2_X1 U12691 ( .A1(n12752), .A2(n12753), .ZN(n12701) );
  AND2_X1 U12692 ( .A1(n12698), .A2(n12697), .ZN(n12753) );
  AND2_X1 U12693 ( .A1(n12695), .A2(n12754), .ZN(n12752) );
  OR2_X1 U12694 ( .A1(n12697), .A2(n12698), .ZN(n12754) );
  OR2_X1 U12695 ( .A1(n8634), .A2(n12381), .ZN(n12698) );
  OR2_X1 U12696 ( .A1(n12755), .A2(n12756), .ZN(n12697) );
  AND2_X1 U12697 ( .A1(n12694), .A2(n12693), .ZN(n12756) );
  AND2_X1 U12698 ( .A1(n12691), .A2(n12757), .ZN(n12755) );
  OR2_X1 U12699 ( .A1(n12693), .A2(n12694), .ZN(n12757) );
  OR2_X1 U12700 ( .A1(n8629), .A2(n12381), .ZN(n12694) );
  OR2_X1 U12701 ( .A1(n12758), .A2(n12759), .ZN(n12693) );
  AND2_X1 U12702 ( .A1(n12690), .A2(n12689), .ZN(n12759) );
  AND2_X1 U12703 ( .A1(n12688), .A2(n12760), .ZN(n12758) );
  OR2_X1 U12704 ( .A1(n12689), .A2(n12690), .ZN(n12760) );
  OR2_X1 U12705 ( .A1(n8624), .A2(n12381), .ZN(n12690) );
  OR2_X1 U12706 ( .A1(n12761), .A2(n12762), .ZN(n12689) );
  AND2_X1 U12707 ( .A1(n12686), .A2(n12685), .ZN(n12762) );
  AND2_X1 U12708 ( .A1(n12684), .A2(n12763), .ZN(n12761) );
  OR2_X1 U12709 ( .A1(n12685), .A2(n12686), .ZN(n12763) );
  OR2_X1 U12710 ( .A1(n8619), .A2(n12381), .ZN(n12686) );
  OR2_X1 U12711 ( .A1(n12764), .A2(n12765), .ZN(n12685) );
  AND2_X1 U12712 ( .A1(n12682), .A2(n12681), .ZN(n12765) );
  AND2_X1 U12713 ( .A1(n12680), .A2(n12766), .ZN(n12764) );
  OR2_X1 U12714 ( .A1(n12681), .A2(n12682), .ZN(n12766) );
  OR2_X1 U12715 ( .A1(n8614), .A2(n12381), .ZN(n12682) );
  OR2_X1 U12716 ( .A1(n12767), .A2(n12768), .ZN(n12681) );
  AND2_X1 U12717 ( .A1(n12678), .A2(n12677), .ZN(n12768) );
  AND2_X1 U12718 ( .A1(n12676), .A2(n12769), .ZN(n12767) );
  OR2_X1 U12719 ( .A1(n12677), .A2(n12678), .ZN(n12769) );
  OR2_X1 U12720 ( .A1(n8609), .A2(n12381), .ZN(n12678) );
  OR2_X1 U12721 ( .A1(n12770), .A2(n12771), .ZN(n12677) );
  AND2_X1 U12722 ( .A1(n12674), .A2(n12673), .ZN(n12771) );
  AND2_X1 U12723 ( .A1(n12671), .A2(n12772), .ZN(n12770) );
  OR2_X1 U12724 ( .A1(n12673), .A2(n12674), .ZN(n12772) );
  OR2_X1 U12725 ( .A1(n8604), .A2(n12381), .ZN(n12674) );
  OR2_X1 U12726 ( .A1(n12773), .A2(n12774), .ZN(n12673) );
  AND2_X1 U12727 ( .A1(n12670), .A2(n12669), .ZN(n12774) );
  AND2_X1 U12728 ( .A1(n12667), .A2(n12775), .ZN(n12773) );
  OR2_X1 U12729 ( .A1(n12669), .A2(n12670), .ZN(n12775) );
  OR2_X1 U12730 ( .A1(n8599), .A2(n12381), .ZN(n12670) );
  OR2_X1 U12731 ( .A1(n12776), .A2(n12777), .ZN(n12669) );
  AND2_X1 U12732 ( .A1(n12666), .A2(n12665), .ZN(n12777) );
  AND2_X1 U12733 ( .A1(n12663), .A2(n12778), .ZN(n12776) );
  OR2_X1 U12734 ( .A1(n12665), .A2(n12666), .ZN(n12778) );
  OR2_X1 U12735 ( .A1(n8594), .A2(n12381), .ZN(n12666) );
  OR2_X1 U12736 ( .A1(n12779), .A2(n12780), .ZN(n12665) );
  AND2_X1 U12737 ( .A1(n12662), .A2(n12661), .ZN(n12780) );
  AND2_X1 U12738 ( .A1(n12659), .A2(n12781), .ZN(n12779) );
  OR2_X1 U12739 ( .A1(n12661), .A2(n12662), .ZN(n12781) );
  OR2_X1 U12740 ( .A1(n8589), .A2(n12381), .ZN(n12662) );
  OR2_X1 U12741 ( .A1(n12782), .A2(n12783), .ZN(n12661) );
  AND2_X1 U12742 ( .A1(n12658), .A2(n12657), .ZN(n12783) );
  AND2_X1 U12743 ( .A1(n12655), .A2(n12784), .ZN(n12782) );
  OR2_X1 U12744 ( .A1(n12657), .A2(n12658), .ZN(n12784) );
  OR2_X1 U12745 ( .A1(n8584), .A2(n12381), .ZN(n12658) );
  OR2_X1 U12746 ( .A1(n12785), .A2(n12786), .ZN(n12657) );
  AND2_X1 U12747 ( .A1(n12654), .A2(n12653), .ZN(n12786) );
  AND2_X1 U12748 ( .A1(n12651), .A2(n12787), .ZN(n12785) );
  OR2_X1 U12749 ( .A1(n12653), .A2(n12654), .ZN(n12787) );
  OR2_X1 U12750 ( .A1(n8579), .A2(n12381), .ZN(n12654) );
  OR2_X1 U12751 ( .A1(n12788), .A2(n12789), .ZN(n12653) );
  AND2_X1 U12752 ( .A1(n12650), .A2(n12649), .ZN(n12789) );
  AND2_X1 U12753 ( .A1(n12647), .A2(n12790), .ZN(n12788) );
  OR2_X1 U12754 ( .A1(n12649), .A2(n12650), .ZN(n12790) );
  OR2_X1 U12755 ( .A1(n8574), .A2(n12381), .ZN(n12650) );
  OR2_X1 U12756 ( .A1(n12791), .A2(n12792), .ZN(n12649) );
  AND2_X1 U12757 ( .A1(n12646), .A2(n12645), .ZN(n12792) );
  AND2_X1 U12758 ( .A1(n12643), .A2(n12793), .ZN(n12791) );
  OR2_X1 U12759 ( .A1(n12645), .A2(n12646), .ZN(n12793) );
  OR2_X1 U12760 ( .A1(n8569), .A2(n12381), .ZN(n12646) );
  OR2_X1 U12761 ( .A1(n12794), .A2(n12795), .ZN(n12645) );
  AND2_X1 U12762 ( .A1(n12642), .A2(n12641), .ZN(n12795) );
  AND2_X1 U12763 ( .A1(n12639), .A2(n12796), .ZN(n12794) );
  OR2_X1 U12764 ( .A1(n12641), .A2(n12642), .ZN(n12796) );
  OR2_X1 U12765 ( .A1(n8564), .A2(n12381), .ZN(n12642) );
  OR2_X1 U12766 ( .A1(n12797), .A2(n12798), .ZN(n12641) );
  AND2_X1 U12767 ( .A1(n12638), .A2(n12637), .ZN(n12798) );
  AND2_X1 U12768 ( .A1(n12635), .A2(n12799), .ZN(n12797) );
  OR2_X1 U12769 ( .A1(n12637), .A2(n12638), .ZN(n12799) );
  OR2_X1 U12770 ( .A1(n8559), .A2(n12381), .ZN(n12638) );
  OR2_X1 U12771 ( .A1(n12800), .A2(n12801), .ZN(n12637) );
  AND2_X1 U12772 ( .A1(n12634), .A2(n12633), .ZN(n12801) );
  AND2_X1 U12773 ( .A1(n12631), .A2(n12802), .ZN(n12800) );
  OR2_X1 U12774 ( .A1(n12633), .A2(n12634), .ZN(n12802) );
  OR2_X1 U12775 ( .A1(n8554), .A2(n12381), .ZN(n12634) );
  OR2_X1 U12776 ( .A1(n12803), .A2(n12804), .ZN(n12633) );
  AND2_X1 U12777 ( .A1(n12630), .A2(n12629), .ZN(n12804) );
  AND2_X1 U12778 ( .A1(n12627), .A2(n12805), .ZN(n12803) );
  OR2_X1 U12779 ( .A1(n12629), .A2(n12630), .ZN(n12805) );
  OR2_X1 U12780 ( .A1(n8549), .A2(n12381), .ZN(n12630) );
  OR2_X1 U12781 ( .A1(n12806), .A2(n12807), .ZN(n12629) );
  AND2_X1 U12782 ( .A1(n12626), .A2(n12625), .ZN(n12807) );
  AND2_X1 U12783 ( .A1(n12623), .A2(n12808), .ZN(n12806) );
  OR2_X1 U12784 ( .A1(n12625), .A2(n12626), .ZN(n12808) );
  OR2_X1 U12785 ( .A1(n8544), .A2(n12381), .ZN(n12626) );
  OR2_X1 U12786 ( .A1(n12809), .A2(n12810), .ZN(n12625) );
  AND2_X1 U12787 ( .A1(n12622), .A2(n12621), .ZN(n12810) );
  AND2_X1 U12788 ( .A1(n12619), .A2(n12811), .ZN(n12809) );
  OR2_X1 U12789 ( .A1(n12621), .A2(n12622), .ZN(n12811) );
  OR2_X1 U12790 ( .A1(n8539), .A2(n12381), .ZN(n12622) );
  OR2_X1 U12791 ( .A1(n12812), .A2(n12813), .ZN(n12621) );
  AND2_X1 U12792 ( .A1(n12618), .A2(n12617), .ZN(n12813) );
  AND2_X1 U12793 ( .A1(n12615), .A2(n12814), .ZN(n12812) );
  OR2_X1 U12794 ( .A1(n12617), .A2(n12618), .ZN(n12814) );
  OR2_X1 U12795 ( .A1(n8534), .A2(n12381), .ZN(n12618) );
  OR2_X1 U12796 ( .A1(n12815), .A2(n12816), .ZN(n12617) );
  AND2_X1 U12797 ( .A1(n12614), .A2(n12613), .ZN(n12816) );
  AND2_X1 U12798 ( .A1(n12611), .A2(n12817), .ZN(n12815) );
  OR2_X1 U12799 ( .A1(n12613), .A2(n12614), .ZN(n12817) );
  OR2_X1 U12800 ( .A1(n8529), .A2(n12381), .ZN(n12614) );
  OR2_X1 U12801 ( .A1(n12818), .A2(n12819), .ZN(n12613) );
  AND2_X1 U12802 ( .A1(n12607), .A2(n12610), .ZN(n12819) );
  AND2_X1 U12803 ( .A1(n12609), .A2(n12820), .ZN(n12818) );
  OR2_X1 U12804 ( .A1(n12610), .A2(n12607), .ZN(n12820) );
  OR2_X1 U12805 ( .A1(n12381), .A2(n8518), .ZN(n12607) );
  OR3_X1 U12806 ( .A1(n12606), .A2(n12381), .A3(n8519), .ZN(n12610) );
  INV_X1 U12807 ( .A(n12376), .ZN(n12381) );
  XOR2_X1 U12808 ( .A(n12821), .B(n12822), .Z(n12376) );
  XNOR2_X1 U12809 ( .A(c_11_), .B(d_11_), .ZN(n12821) );
  INV_X1 U12810 ( .A(n12823), .ZN(n12609) );
  OR2_X1 U12811 ( .A1(n12824), .A2(n12825), .ZN(n12823) );
  AND2_X1 U12812 ( .A1(n12826), .A2(n12827), .ZN(n12825) );
  OR2_X1 U12813 ( .A1(n12828), .A2(n7697), .ZN(n12827) );
  AND2_X1 U12814 ( .A1(n12606), .A2(n7691), .ZN(n12828) );
  AND2_X1 U12815 ( .A1(n12601), .A2(n12829), .ZN(n12824) );
  OR2_X1 U12816 ( .A1(n12830), .A2(n7701), .ZN(n12829) );
  AND2_X1 U12817 ( .A1(n12831), .A2(n7703), .ZN(n12830) );
  XNOR2_X1 U12818 ( .A(n12832), .B(n12833), .ZN(n12611) );
  XNOR2_X1 U12819 ( .A(n12834), .B(n12835), .ZN(n12833) );
  XOR2_X1 U12820 ( .A(n12836), .B(n12837), .Z(n12615) );
  XOR2_X1 U12821 ( .A(n12838), .B(n12839), .Z(n12837) );
  XOR2_X1 U12822 ( .A(n12840), .B(n12841), .Z(n12619) );
  XOR2_X1 U12823 ( .A(n12842), .B(n12843), .Z(n12841) );
  XOR2_X1 U12824 ( .A(n12844), .B(n12845), .Z(n12623) );
  XOR2_X1 U12825 ( .A(n12846), .B(n12847), .Z(n12845) );
  XOR2_X1 U12826 ( .A(n12848), .B(n12849), .Z(n12627) );
  XOR2_X1 U12827 ( .A(n12850), .B(n12851), .Z(n12849) );
  XOR2_X1 U12828 ( .A(n12852), .B(n12853), .Z(n12631) );
  XOR2_X1 U12829 ( .A(n12854), .B(n12855), .Z(n12853) );
  XOR2_X1 U12830 ( .A(n12856), .B(n12857), .Z(n12635) );
  XOR2_X1 U12831 ( .A(n12858), .B(n12859), .Z(n12857) );
  XOR2_X1 U12832 ( .A(n12860), .B(n12861), .Z(n12639) );
  XOR2_X1 U12833 ( .A(n12862), .B(n12863), .Z(n12861) );
  XOR2_X1 U12834 ( .A(n12864), .B(n12865), .Z(n12643) );
  XOR2_X1 U12835 ( .A(n12866), .B(n12867), .Z(n12865) );
  XOR2_X1 U12836 ( .A(n12868), .B(n12869), .Z(n12647) );
  XOR2_X1 U12837 ( .A(n12870), .B(n12871), .Z(n12869) );
  XOR2_X1 U12838 ( .A(n12872), .B(n12873), .Z(n12651) );
  XOR2_X1 U12839 ( .A(n12874), .B(n12875), .Z(n12873) );
  XOR2_X1 U12840 ( .A(n12876), .B(n12877), .Z(n12655) );
  XOR2_X1 U12841 ( .A(n12878), .B(n12879), .Z(n12877) );
  XOR2_X1 U12842 ( .A(n12880), .B(n12881), .Z(n12659) );
  XOR2_X1 U12843 ( .A(n12882), .B(n12883), .Z(n12881) );
  XOR2_X1 U12844 ( .A(n12884), .B(n12885), .Z(n12663) );
  XOR2_X1 U12845 ( .A(n12886), .B(n12887), .Z(n12885) );
  XOR2_X1 U12846 ( .A(n12888), .B(n12889), .Z(n12667) );
  XOR2_X1 U12847 ( .A(n12890), .B(n12891), .Z(n12889) );
  XNOR2_X1 U12848 ( .A(n12892), .B(n12893), .ZN(n12671) );
  XNOR2_X1 U12849 ( .A(n12894), .B(n12895), .ZN(n12892) );
  XNOR2_X1 U12850 ( .A(n12896), .B(n12897), .ZN(n12676) );
  XNOR2_X1 U12851 ( .A(n12898), .B(n12899), .ZN(n12896) );
  XNOR2_X1 U12852 ( .A(n12900), .B(n12901), .ZN(n12680) );
  XNOR2_X1 U12853 ( .A(n12902), .B(n12903), .ZN(n12900) );
  XOR2_X1 U12854 ( .A(n12904), .B(n12905), .Z(n12684) );
  XOR2_X1 U12855 ( .A(n12906), .B(n12907), .Z(n12905) );
  XOR2_X1 U12856 ( .A(n12908), .B(n12909), .Z(n12688) );
  XOR2_X1 U12857 ( .A(n12910), .B(n12911), .Z(n12909) );
  XOR2_X1 U12858 ( .A(n12912), .B(n12913), .Z(n12691) );
  XOR2_X1 U12859 ( .A(n12914), .B(n12915), .Z(n12913) );
  XOR2_X1 U12860 ( .A(n12916), .B(n12917), .Z(n12695) );
  XOR2_X1 U12861 ( .A(n12918), .B(n12919), .Z(n12917) );
  XOR2_X1 U12862 ( .A(n12920), .B(n12921), .Z(n12699) );
  XOR2_X1 U12863 ( .A(n12922), .B(n12923), .Z(n12921) );
  XOR2_X1 U12864 ( .A(n12924), .B(n12925), .Z(n12703) );
  XOR2_X1 U12865 ( .A(n12926), .B(n12927), .Z(n12925) );
  XOR2_X1 U12866 ( .A(n12928), .B(n12929), .Z(n12707) );
  XOR2_X1 U12867 ( .A(n12930), .B(n12931), .Z(n12929) );
  XOR2_X1 U12868 ( .A(n12932), .B(n12933), .Z(n12711) );
  XOR2_X1 U12869 ( .A(n12934), .B(n12935), .Z(n12933) );
  XOR2_X1 U12870 ( .A(n12936), .B(n12937), .Z(n12715) );
  XOR2_X1 U12871 ( .A(n12938), .B(n12939), .Z(n12937) );
  XOR2_X1 U12872 ( .A(n12940), .B(n12941), .Z(n12719) );
  XOR2_X1 U12873 ( .A(n12942), .B(n12943), .Z(n12941) );
  XOR2_X1 U12874 ( .A(n12944), .B(n12945), .Z(n12723) );
  XOR2_X1 U12875 ( .A(n12946), .B(n12947), .Z(n12945) );
  XOR2_X1 U12876 ( .A(n12948), .B(n12949), .Z(n12728) );
  XOR2_X1 U12877 ( .A(n12950), .B(n12951), .Z(n12949) );
  XNOR2_X1 U12878 ( .A(n7675), .B(n8166), .ZN(n7953) );
  OR2_X1 U12879 ( .A1(n12952), .A2(n12953), .ZN(n8166) );
  AND2_X1 U12880 ( .A1(n12951), .A2(n12950), .ZN(n12953) );
  AND2_X1 U12881 ( .A1(n12948), .A2(n12954), .ZN(n12952) );
  OR2_X1 U12882 ( .A1(n12950), .A2(n12951), .ZN(n12954) );
  OR2_X1 U12883 ( .A1(n12606), .A2(n7960), .ZN(n12951) );
  OR2_X1 U12884 ( .A1(n12955), .A2(n12956), .ZN(n12950) );
  AND2_X1 U12885 ( .A1(n12947), .A2(n12946), .ZN(n12956) );
  AND2_X1 U12886 ( .A1(n12944), .A2(n12957), .ZN(n12955) );
  OR2_X1 U12887 ( .A1(n12946), .A2(n12947), .ZN(n12957) );
  OR2_X1 U12888 ( .A1(n12606), .A2(n7608), .ZN(n12947) );
  OR2_X1 U12889 ( .A1(n12958), .A2(n12959), .ZN(n12946) );
  AND2_X1 U12890 ( .A1(n12943), .A2(n12942), .ZN(n12959) );
  AND2_X1 U12891 ( .A1(n12940), .A2(n12960), .ZN(n12958) );
  OR2_X1 U12892 ( .A1(n12942), .A2(n12943), .ZN(n12960) );
  OR2_X1 U12893 ( .A1(n12606), .A2(n7610), .ZN(n12943) );
  OR2_X1 U12894 ( .A1(n12961), .A2(n12962), .ZN(n12942) );
  AND2_X1 U12895 ( .A1(n12939), .A2(n12938), .ZN(n12962) );
  AND2_X1 U12896 ( .A1(n12936), .A2(n12963), .ZN(n12961) );
  OR2_X1 U12897 ( .A1(n12938), .A2(n12939), .ZN(n12963) );
  OR2_X1 U12898 ( .A1(n12606), .A2(n7612), .ZN(n12939) );
  OR2_X1 U12899 ( .A1(n12964), .A2(n12965), .ZN(n12938) );
  AND2_X1 U12900 ( .A1(n12935), .A2(n12934), .ZN(n12965) );
  AND2_X1 U12901 ( .A1(n12932), .A2(n12966), .ZN(n12964) );
  OR2_X1 U12902 ( .A1(n12934), .A2(n12935), .ZN(n12966) );
  OR2_X1 U12903 ( .A1(n12606), .A2(n7614), .ZN(n12935) );
  OR2_X1 U12904 ( .A1(n12967), .A2(n12968), .ZN(n12934) );
  AND2_X1 U12905 ( .A1(n12931), .A2(n12930), .ZN(n12968) );
  AND2_X1 U12906 ( .A1(n12928), .A2(n12969), .ZN(n12967) );
  OR2_X1 U12907 ( .A1(n12930), .A2(n12931), .ZN(n12969) );
  OR2_X1 U12908 ( .A1(n8644), .A2(n12606), .ZN(n12931) );
  OR2_X1 U12909 ( .A1(n12970), .A2(n12971), .ZN(n12930) );
  AND2_X1 U12910 ( .A1(n12927), .A2(n12926), .ZN(n12971) );
  AND2_X1 U12911 ( .A1(n12924), .A2(n12972), .ZN(n12970) );
  OR2_X1 U12912 ( .A1(n12926), .A2(n12927), .ZN(n12972) );
  OR2_X1 U12913 ( .A1(n8639), .A2(n12606), .ZN(n12927) );
  OR2_X1 U12914 ( .A1(n12973), .A2(n12974), .ZN(n12926) );
  AND2_X1 U12915 ( .A1(n12923), .A2(n12922), .ZN(n12974) );
  AND2_X1 U12916 ( .A1(n12920), .A2(n12975), .ZN(n12973) );
  OR2_X1 U12917 ( .A1(n12922), .A2(n12923), .ZN(n12975) );
  OR2_X1 U12918 ( .A1(n8634), .A2(n12606), .ZN(n12923) );
  OR2_X1 U12919 ( .A1(n12976), .A2(n12977), .ZN(n12922) );
  AND2_X1 U12920 ( .A1(n12919), .A2(n12918), .ZN(n12977) );
  AND2_X1 U12921 ( .A1(n12916), .A2(n12978), .ZN(n12976) );
  OR2_X1 U12922 ( .A1(n12918), .A2(n12919), .ZN(n12978) );
  OR2_X1 U12923 ( .A1(n8629), .A2(n12606), .ZN(n12919) );
  OR2_X1 U12924 ( .A1(n12979), .A2(n12980), .ZN(n12918) );
  AND2_X1 U12925 ( .A1(n12915), .A2(n12914), .ZN(n12980) );
  AND2_X1 U12926 ( .A1(n12912), .A2(n12981), .ZN(n12979) );
  OR2_X1 U12927 ( .A1(n12914), .A2(n12915), .ZN(n12981) );
  OR2_X1 U12928 ( .A1(n8624), .A2(n12606), .ZN(n12915) );
  OR2_X1 U12929 ( .A1(n12982), .A2(n12983), .ZN(n12914) );
  AND2_X1 U12930 ( .A1(n12911), .A2(n12910), .ZN(n12983) );
  AND2_X1 U12931 ( .A1(n12908), .A2(n12984), .ZN(n12982) );
  OR2_X1 U12932 ( .A1(n12910), .A2(n12911), .ZN(n12984) );
  OR2_X1 U12933 ( .A1(n8619), .A2(n12606), .ZN(n12911) );
  OR2_X1 U12934 ( .A1(n12985), .A2(n12986), .ZN(n12910) );
  AND2_X1 U12935 ( .A1(n12907), .A2(n12906), .ZN(n12986) );
  AND2_X1 U12936 ( .A1(n12904), .A2(n12987), .ZN(n12985) );
  OR2_X1 U12937 ( .A1(n12906), .A2(n12907), .ZN(n12987) );
  OR2_X1 U12938 ( .A1(n8614), .A2(n12606), .ZN(n12907) );
  OR2_X1 U12939 ( .A1(n12988), .A2(n12989), .ZN(n12906) );
  AND2_X1 U12940 ( .A1(n12903), .A2(n12902), .ZN(n12989) );
  AND2_X1 U12941 ( .A1(n12901), .A2(n12990), .ZN(n12988) );
  OR2_X1 U12942 ( .A1(n12902), .A2(n12903), .ZN(n12990) );
  OR2_X1 U12943 ( .A1(n8609), .A2(n12606), .ZN(n12903) );
  OR2_X1 U12944 ( .A1(n12991), .A2(n12992), .ZN(n12902) );
  AND2_X1 U12945 ( .A1(n12899), .A2(n12898), .ZN(n12992) );
  AND2_X1 U12946 ( .A1(n12897), .A2(n12993), .ZN(n12991) );
  OR2_X1 U12947 ( .A1(n12898), .A2(n12899), .ZN(n12993) );
  OR2_X1 U12948 ( .A1(n8604), .A2(n12606), .ZN(n12899) );
  OR2_X1 U12949 ( .A1(n12994), .A2(n12995), .ZN(n12898) );
  AND2_X1 U12950 ( .A1(n12895), .A2(n12894), .ZN(n12995) );
  AND2_X1 U12951 ( .A1(n12893), .A2(n12996), .ZN(n12994) );
  OR2_X1 U12952 ( .A1(n12894), .A2(n12895), .ZN(n12996) );
  OR2_X1 U12953 ( .A1(n8599), .A2(n12606), .ZN(n12895) );
  OR2_X1 U12954 ( .A1(n12997), .A2(n12998), .ZN(n12894) );
  AND2_X1 U12955 ( .A1(n12891), .A2(n12890), .ZN(n12998) );
  AND2_X1 U12956 ( .A1(n12888), .A2(n12999), .ZN(n12997) );
  OR2_X1 U12957 ( .A1(n12890), .A2(n12891), .ZN(n12999) );
  OR2_X1 U12958 ( .A1(n8594), .A2(n12606), .ZN(n12891) );
  OR2_X1 U12959 ( .A1(n13000), .A2(n13001), .ZN(n12890) );
  AND2_X1 U12960 ( .A1(n12887), .A2(n12886), .ZN(n13001) );
  AND2_X1 U12961 ( .A1(n12884), .A2(n13002), .ZN(n13000) );
  OR2_X1 U12962 ( .A1(n12886), .A2(n12887), .ZN(n13002) );
  OR2_X1 U12963 ( .A1(n8589), .A2(n12606), .ZN(n12887) );
  OR2_X1 U12964 ( .A1(n13003), .A2(n13004), .ZN(n12886) );
  AND2_X1 U12965 ( .A1(n12883), .A2(n12882), .ZN(n13004) );
  AND2_X1 U12966 ( .A1(n12880), .A2(n13005), .ZN(n13003) );
  OR2_X1 U12967 ( .A1(n12882), .A2(n12883), .ZN(n13005) );
  OR2_X1 U12968 ( .A1(n8584), .A2(n12606), .ZN(n12883) );
  OR2_X1 U12969 ( .A1(n13006), .A2(n13007), .ZN(n12882) );
  AND2_X1 U12970 ( .A1(n12879), .A2(n12878), .ZN(n13007) );
  AND2_X1 U12971 ( .A1(n12876), .A2(n13008), .ZN(n13006) );
  OR2_X1 U12972 ( .A1(n12878), .A2(n12879), .ZN(n13008) );
  OR2_X1 U12973 ( .A1(n8579), .A2(n12606), .ZN(n12879) );
  OR2_X1 U12974 ( .A1(n13009), .A2(n13010), .ZN(n12878) );
  AND2_X1 U12975 ( .A1(n12872), .A2(n12875), .ZN(n13010) );
  AND2_X1 U12976 ( .A1(n13011), .A2(n12874), .ZN(n13009) );
  OR2_X1 U12977 ( .A1(n13012), .A2(n13013), .ZN(n12874) );
  AND2_X1 U12978 ( .A1(n12871), .A2(n12870), .ZN(n13013) );
  AND2_X1 U12979 ( .A1(n12868), .A2(n13014), .ZN(n13012) );
  OR2_X1 U12980 ( .A1(n12870), .A2(n12871), .ZN(n13014) );
  OR2_X1 U12981 ( .A1(n8569), .A2(n12606), .ZN(n12871) );
  OR2_X1 U12982 ( .A1(n13015), .A2(n13016), .ZN(n12870) );
  AND2_X1 U12983 ( .A1(n12864), .A2(n12867), .ZN(n13016) );
  AND2_X1 U12984 ( .A1(n13017), .A2(n12866), .ZN(n13015) );
  OR2_X1 U12985 ( .A1(n13018), .A2(n13019), .ZN(n12866) );
  AND2_X1 U12986 ( .A1(n12860), .A2(n12863), .ZN(n13019) );
  AND2_X1 U12987 ( .A1(n13020), .A2(n12862), .ZN(n13018) );
  OR2_X1 U12988 ( .A1(n13021), .A2(n13022), .ZN(n12862) );
  AND2_X1 U12989 ( .A1(n12856), .A2(n12859), .ZN(n13022) );
  AND2_X1 U12990 ( .A1(n13023), .A2(n12858), .ZN(n13021) );
  OR2_X1 U12991 ( .A1(n13024), .A2(n13025), .ZN(n12858) );
  AND2_X1 U12992 ( .A1(n12852), .A2(n12855), .ZN(n13025) );
  AND2_X1 U12993 ( .A1(n13026), .A2(n12854), .ZN(n13024) );
  OR2_X1 U12994 ( .A1(n13027), .A2(n13028), .ZN(n12854) );
  AND2_X1 U12995 ( .A1(n12848), .A2(n12851), .ZN(n13028) );
  AND2_X1 U12996 ( .A1(n13029), .A2(n12850), .ZN(n13027) );
  OR2_X1 U12997 ( .A1(n13030), .A2(n13031), .ZN(n12850) );
  AND2_X1 U12998 ( .A1(n12844), .A2(n12847), .ZN(n13031) );
  AND2_X1 U12999 ( .A1(n13032), .A2(n12846), .ZN(n13030) );
  OR2_X1 U13000 ( .A1(n13033), .A2(n13034), .ZN(n12846) );
  AND2_X1 U13001 ( .A1(n12840), .A2(n12843), .ZN(n13034) );
  AND2_X1 U13002 ( .A1(n13035), .A2(n12842), .ZN(n13033) );
  OR2_X1 U13003 ( .A1(n13036), .A2(n13037), .ZN(n12842) );
  AND2_X1 U13004 ( .A1(n12836), .A2(n12839), .ZN(n13037) );
  AND2_X1 U13005 ( .A1(n13038), .A2(n12838), .ZN(n13036) );
  OR2_X1 U13006 ( .A1(n13039), .A2(n13040), .ZN(n12838) );
  AND2_X1 U13007 ( .A1(n12832), .A2(n12835), .ZN(n13040) );
  AND2_X1 U13008 ( .A1(n12834), .A2(n13041), .ZN(n13039) );
  OR2_X1 U13009 ( .A1(n12835), .A2(n12832), .ZN(n13041) );
  OR2_X1 U13010 ( .A1(n12606), .A2(n8518), .ZN(n12832) );
  OR3_X1 U13011 ( .A1(n12831), .A2(n12606), .A3(n8519), .ZN(n12835) );
  INV_X1 U13012 ( .A(n13042), .ZN(n12834) );
  OR2_X1 U13013 ( .A1(n13043), .A2(n13044), .ZN(n13042) );
  AND2_X1 U13014 ( .A1(n13045), .A2(n13046), .ZN(n13044) );
  OR2_X1 U13015 ( .A1(n13047), .A2(n7697), .ZN(n13046) );
  AND2_X1 U13016 ( .A1(n12831), .A2(n7691), .ZN(n13047) );
  AND2_X1 U13017 ( .A1(n12826), .A2(n13048), .ZN(n13043) );
  OR2_X1 U13018 ( .A1(n13049), .A2(n7701), .ZN(n13048) );
  AND2_X1 U13019 ( .A1(n13050), .A2(n7703), .ZN(n13049) );
  OR2_X1 U13020 ( .A1(n12839), .A2(n12836), .ZN(n13038) );
  XNOR2_X1 U13021 ( .A(n13051), .B(n13052), .ZN(n12836) );
  XNOR2_X1 U13022 ( .A(n13053), .B(n13054), .ZN(n13052) );
  OR2_X1 U13023 ( .A1(n8529), .A2(n12606), .ZN(n12839) );
  OR2_X1 U13024 ( .A1(n12843), .A2(n12840), .ZN(n13035) );
  XOR2_X1 U13025 ( .A(n13055), .B(n13056), .Z(n12840) );
  XOR2_X1 U13026 ( .A(n13057), .B(n13058), .Z(n13056) );
  OR2_X1 U13027 ( .A1(n8534), .A2(n12606), .ZN(n12843) );
  OR2_X1 U13028 ( .A1(n12847), .A2(n12844), .ZN(n13032) );
  XOR2_X1 U13029 ( .A(n13059), .B(n13060), .Z(n12844) );
  XOR2_X1 U13030 ( .A(n13061), .B(n13062), .Z(n13060) );
  OR2_X1 U13031 ( .A1(n8539), .A2(n12606), .ZN(n12847) );
  OR2_X1 U13032 ( .A1(n12851), .A2(n12848), .ZN(n13029) );
  XOR2_X1 U13033 ( .A(n13063), .B(n13064), .Z(n12848) );
  XOR2_X1 U13034 ( .A(n13065), .B(n13066), .Z(n13064) );
  OR2_X1 U13035 ( .A1(n8544), .A2(n12606), .ZN(n12851) );
  OR2_X1 U13036 ( .A1(n12855), .A2(n12852), .ZN(n13026) );
  XOR2_X1 U13037 ( .A(n13067), .B(n13068), .Z(n12852) );
  XOR2_X1 U13038 ( .A(n13069), .B(n13070), .Z(n13068) );
  OR2_X1 U13039 ( .A1(n8549), .A2(n12606), .ZN(n12855) );
  OR2_X1 U13040 ( .A1(n12859), .A2(n12856), .ZN(n13023) );
  XOR2_X1 U13041 ( .A(n13071), .B(n13072), .Z(n12856) );
  XOR2_X1 U13042 ( .A(n13073), .B(n13074), .Z(n13072) );
  OR2_X1 U13043 ( .A1(n8554), .A2(n12606), .ZN(n12859) );
  OR2_X1 U13044 ( .A1(n12863), .A2(n12860), .ZN(n13020) );
  XOR2_X1 U13045 ( .A(n13075), .B(n13076), .Z(n12860) );
  XOR2_X1 U13046 ( .A(n13077), .B(n13078), .Z(n13076) );
  OR2_X1 U13047 ( .A1(n8559), .A2(n12606), .ZN(n12863) );
  OR2_X1 U13048 ( .A1(n12867), .A2(n12864), .ZN(n13017) );
  XOR2_X1 U13049 ( .A(n13079), .B(n13080), .Z(n12864) );
  XOR2_X1 U13050 ( .A(n13081), .B(n13082), .Z(n13080) );
  OR2_X1 U13051 ( .A1(n8564), .A2(n12606), .ZN(n12867) );
  XOR2_X1 U13052 ( .A(n13083), .B(n13084), .Z(n12868) );
  XOR2_X1 U13053 ( .A(n13085), .B(n13086), .Z(n13084) );
  OR2_X1 U13054 ( .A1(n12875), .A2(n12872), .ZN(n13011) );
  XOR2_X1 U13055 ( .A(n13087), .B(n13088), .Z(n12872) );
  XOR2_X1 U13056 ( .A(n13089), .B(n13090), .Z(n13088) );
  OR2_X1 U13057 ( .A1(n8574), .A2(n12606), .ZN(n12875) );
  INV_X1 U13058 ( .A(n12601), .ZN(n12606) );
  XOR2_X1 U13059 ( .A(n13091), .B(n13092), .Z(n12601) );
  XNOR2_X1 U13060 ( .A(c_10_), .B(d_10_), .ZN(n13091) );
  XOR2_X1 U13061 ( .A(n13093), .B(n13094), .Z(n12876) );
  XOR2_X1 U13062 ( .A(n13095), .B(n13096), .Z(n13094) );
  XOR2_X1 U13063 ( .A(n13097), .B(n13098), .Z(n12880) );
  XOR2_X1 U13064 ( .A(n13099), .B(n13100), .Z(n13098) );
  XOR2_X1 U13065 ( .A(n13101), .B(n13102), .Z(n12884) );
  XOR2_X1 U13066 ( .A(n13103), .B(n13104), .Z(n13102) );
  XNOR2_X1 U13067 ( .A(n13105), .B(n13106), .ZN(n12888) );
  XNOR2_X1 U13068 ( .A(n13107), .B(n13108), .ZN(n13105) );
  XNOR2_X1 U13069 ( .A(n13109), .B(n13110), .ZN(n12893) );
  XNOR2_X1 U13070 ( .A(n13111), .B(n13112), .ZN(n13109) );
  XNOR2_X1 U13071 ( .A(n13113), .B(n13114), .ZN(n12897) );
  XNOR2_X1 U13072 ( .A(n13115), .B(n13116), .ZN(n13113) );
  XOR2_X1 U13073 ( .A(n13117), .B(n13118), .Z(n12901) );
  XOR2_X1 U13074 ( .A(n13119), .B(n13120), .Z(n13118) );
  XOR2_X1 U13075 ( .A(n13121), .B(n13122), .Z(n12904) );
  XOR2_X1 U13076 ( .A(n13123), .B(n13124), .Z(n13122) );
  XOR2_X1 U13077 ( .A(n13125), .B(n13126), .Z(n12908) );
  XOR2_X1 U13078 ( .A(n13127), .B(n13128), .Z(n13126) );
  XOR2_X1 U13079 ( .A(n13129), .B(n13130), .Z(n12912) );
  XOR2_X1 U13080 ( .A(n13131), .B(n13132), .Z(n13130) );
  XOR2_X1 U13081 ( .A(n13133), .B(n13134), .Z(n12916) );
  XOR2_X1 U13082 ( .A(n13135), .B(n13136), .Z(n13134) );
  XOR2_X1 U13083 ( .A(n13137), .B(n13138), .Z(n12920) );
  XOR2_X1 U13084 ( .A(n13139), .B(n13140), .Z(n13138) );
  XOR2_X1 U13085 ( .A(n13141), .B(n13142), .Z(n12924) );
  XOR2_X1 U13086 ( .A(n13143), .B(n13144), .Z(n13142) );
  XOR2_X1 U13087 ( .A(n13145), .B(n13146), .Z(n12928) );
  XOR2_X1 U13088 ( .A(n13147), .B(n13148), .Z(n13146) );
  XOR2_X1 U13089 ( .A(n13149), .B(n13150), .Z(n12932) );
  XOR2_X1 U13090 ( .A(n13151), .B(n13152), .Z(n13150) );
  XOR2_X1 U13091 ( .A(n13153), .B(n13154), .Z(n12936) );
  XOR2_X1 U13092 ( .A(n13155), .B(n13156), .Z(n13154) );
  XOR2_X1 U13093 ( .A(n13157), .B(n13158), .Z(n12940) );
  XOR2_X1 U13094 ( .A(n13159), .B(n13160), .Z(n13158) );
  XOR2_X1 U13095 ( .A(n13161), .B(n13162), .Z(n12944) );
  XOR2_X1 U13096 ( .A(n13163), .B(n13164), .Z(n13162) );
  XOR2_X1 U13097 ( .A(n13165), .B(n13166), .Z(n12948) );
  XOR2_X1 U13098 ( .A(n13167), .B(n13168), .Z(n13166) );
  XNOR2_X1 U13099 ( .A(n13169), .B(n13170), .ZN(n7675) );
  XOR2_X1 U13100 ( .A(n13171), .B(n13172), .Z(n13170) );
  INV_X1 U13101 ( .A(n13173), .ZN(n7672) );
  OR2_X1 U13102 ( .A1(n13174), .A2(n8164), .ZN(n13173) );
  INV_X1 U13103 ( .A(n13175), .ZN(n8164) );
  OR2_X1 U13104 ( .A1(n13176), .A2(n13177), .ZN(n13175) );
  AND2_X1 U13105 ( .A1(n13176), .A2(n13177), .ZN(n13174) );
  OR2_X1 U13106 ( .A1(n13178), .A2(n13179), .ZN(n13177) );
  AND2_X1 U13107 ( .A1(n13172), .A2(n13171), .ZN(n13179) );
  AND2_X1 U13108 ( .A1(n13169), .A2(n13180), .ZN(n13178) );
  OR2_X1 U13109 ( .A1(n13171), .A2(n13172), .ZN(n13180) );
  OR2_X1 U13110 ( .A1(n12831), .A2(n7960), .ZN(n13172) );
  OR2_X1 U13111 ( .A1(n13181), .A2(n13182), .ZN(n13171) );
  AND2_X1 U13112 ( .A1(n13168), .A2(n13167), .ZN(n13182) );
  AND2_X1 U13113 ( .A1(n13165), .A2(n13183), .ZN(n13181) );
  OR2_X1 U13114 ( .A1(n13167), .A2(n13168), .ZN(n13183) );
  OR2_X1 U13115 ( .A1(n12831), .A2(n7608), .ZN(n13168) );
  OR2_X1 U13116 ( .A1(n13184), .A2(n13185), .ZN(n13167) );
  AND2_X1 U13117 ( .A1(n13164), .A2(n13163), .ZN(n13185) );
  AND2_X1 U13118 ( .A1(n13161), .A2(n13186), .ZN(n13184) );
  OR2_X1 U13119 ( .A1(n13163), .A2(n13164), .ZN(n13186) );
  OR2_X1 U13120 ( .A1(n12831), .A2(n7610), .ZN(n13164) );
  OR2_X1 U13121 ( .A1(n13187), .A2(n13188), .ZN(n13163) );
  AND2_X1 U13122 ( .A1(n13160), .A2(n13159), .ZN(n13188) );
  AND2_X1 U13123 ( .A1(n13157), .A2(n13189), .ZN(n13187) );
  OR2_X1 U13124 ( .A1(n13159), .A2(n13160), .ZN(n13189) );
  OR2_X1 U13125 ( .A1(n12831), .A2(n7612), .ZN(n13160) );
  OR2_X1 U13126 ( .A1(n13190), .A2(n13191), .ZN(n13159) );
  AND2_X1 U13127 ( .A1(n13156), .A2(n13155), .ZN(n13191) );
  AND2_X1 U13128 ( .A1(n13153), .A2(n13192), .ZN(n13190) );
  OR2_X1 U13129 ( .A1(n13155), .A2(n13156), .ZN(n13192) );
  OR2_X1 U13130 ( .A1(n12831), .A2(n7614), .ZN(n13156) );
  OR2_X1 U13131 ( .A1(n13193), .A2(n13194), .ZN(n13155) );
  AND2_X1 U13132 ( .A1(n13152), .A2(n13151), .ZN(n13194) );
  AND2_X1 U13133 ( .A1(n13149), .A2(n13195), .ZN(n13193) );
  OR2_X1 U13134 ( .A1(n13151), .A2(n13152), .ZN(n13195) );
  OR2_X1 U13135 ( .A1(n12831), .A2(n7616), .ZN(n13152) );
  OR2_X1 U13136 ( .A1(n13196), .A2(n13197), .ZN(n13151) );
  AND2_X1 U13137 ( .A1(n13148), .A2(n13147), .ZN(n13197) );
  AND2_X1 U13138 ( .A1(n13145), .A2(n13198), .ZN(n13196) );
  OR2_X1 U13139 ( .A1(n13147), .A2(n13148), .ZN(n13198) );
  OR2_X1 U13140 ( .A1(n8639), .A2(n12831), .ZN(n13148) );
  OR2_X1 U13141 ( .A1(n13199), .A2(n13200), .ZN(n13147) );
  AND2_X1 U13142 ( .A1(n13144), .A2(n13143), .ZN(n13200) );
  AND2_X1 U13143 ( .A1(n13141), .A2(n13201), .ZN(n13199) );
  OR2_X1 U13144 ( .A1(n13143), .A2(n13144), .ZN(n13201) );
  OR2_X1 U13145 ( .A1(n8634), .A2(n12831), .ZN(n13144) );
  OR2_X1 U13146 ( .A1(n13202), .A2(n13203), .ZN(n13143) );
  AND2_X1 U13147 ( .A1(n13140), .A2(n13139), .ZN(n13203) );
  AND2_X1 U13148 ( .A1(n13137), .A2(n13204), .ZN(n13202) );
  OR2_X1 U13149 ( .A1(n13139), .A2(n13140), .ZN(n13204) );
  OR2_X1 U13150 ( .A1(n8629), .A2(n12831), .ZN(n13140) );
  OR2_X1 U13151 ( .A1(n13205), .A2(n13206), .ZN(n13139) );
  AND2_X1 U13152 ( .A1(n13136), .A2(n13135), .ZN(n13206) );
  AND2_X1 U13153 ( .A1(n13133), .A2(n13207), .ZN(n13205) );
  OR2_X1 U13154 ( .A1(n13135), .A2(n13136), .ZN(n13207) );
  OR2_X1 U13155 ( .A1(n8624), .A2(n12831), .ZN(n13136) );
  OR2_X1 U13156 ( .A1(n13208), .A2(n13209), .ZN(n13135) );
  AND2_X1 U13157 ( .A1(n13132), .A2(n13131), .ZN(n13209) );
  AND2_X1 U13158 ( .A1(n13129), .A2(n13210), .ZN(n13208) );
  OR2_X1 U13159 ( .A1(n13131), .A2(n13132), .ZN(n13210) );
  OR2_X1 U13160 ( .A1(n8619), .A2(n12831), .ZN(n13132) );
  OR2_X1 U13161 ( .A1(n13211), .A2(n13212), .ZN(n13131) );
  AND2_X1 U13162 ( .A1(n13128), .A2(n13127), .ZN(n13212) );
  AND2_X1 U13163 ( .A1(n13125), .A2(n13213), .ZN(n13211) );
  OR2_X1 U13164 ( .A1(n13127), .A2(n13128), .ZN(n13213) );
  OR2_X1 U13165 ( .A1(n8614), .A2(n12831), .ZN(n13128) );
  OR2_X1 U13166 ( .A1(n13214), .A2(n13215), .ZN(n13127) );
  AND2_X1 U13167 ( .A1(n13124), .A2(n13123), .ZN(n13215) );
  AND2_X1 U13168 ( .A1(n13121), .A2(n13216), .ZN(n13214) );
  OR2_X1 U13169 ( .A1(n13123), .A2(n13124), .ZN(n13216) );
  OR2_X1 U13170 ( .A1(n8609), .A2(n12831), .ZN(n13124) );
  OR2_X1 U13171 ( .A1(n13217), .A2(n13218), .ZN(n13123) );
  AND2_X1 U13172 ( .A1(n13120), .A2(n13119), .ZN(n13218) );
  AND2_X1 U13173 ( .A1(n13117), .A2(n13219), .ZN(n13217) );
  OR2_X1 U13174 ( .A1(n13119), .A2(n13120), .ZN(n13219) );
  OR2_X1 U13175 ( .A1(n8604), .A2(n12831), .ZN(n13120) );
  OR2_X1 U13176 ( .A1(n13220), .A2(n13221), .ZN(n13119) );
  AND2_X1 U13177 ( .A1(n13116), .A2(n13115), .ZN(n13221) );
  AND2_X1 U13178 ( .A1(n13114), .A2(n13222), .ZN(n13220) );
  OR2_X1 U13179 ( .A1(n13115), .A2(n13116), .ZN(n13222) );
  OR2_X1 U13180 ( .A1(n8599), .A2(n12831), .ZN(n13116) );
  OR2_X1 U13181 ( .A1(n13223), .A2(n13224), .ZN(n13115) );
  AND2_X1 U13182 ( .A1(n13112), .A2(n13111), .ZN(n13224) );
  AND2_X1 U13183 ( .A1(n13110), .A2(n13225), .ZN(n13223) );
  OR2_X1 U13184 ( .A1(n13111), .A2(n13112), .ZN(n13225) );
  OR2_X1 U13185 ( .A1(n8594), .A2(n12831), .ZN(n13112) );
  OR2_X1 U13186 ( .A1(n13226), .A2(n13227), .ZN(n13111) );
  AND2_X1 U13187 ( .A1(n13108), .A2(n13107), .ZN(n13227) );
  AND2_X1 U13188 ( .A1(n13106), .A2(n13228), .ZN(n13226) );
  OR2_X1 U13189 ( .A1(n13107), .A2(n13108), .ZN(n13228) );
  OR2_X1 U13190 ( .A1(n8589), .A2(n12831), .ZN(n13108) );
  OR2_X1 U13191 ( .A1(n13229), .A2(n13230), .ZN(n13107) );
  AND2_X1 U13192 ( .A1(n13104), .A2(n13103), .ZN(n13230) );
  AND2_X1 U13193 ( .A1(n13101), .A2(n13231), .ZN(n13229) );
  OR2_X1 U13194 ( .A1(n13103), .A2(n13104), .ZN(n13231) );
  OR2_X1 U13195 ( .A1(n8584), .A2(n12831), .ZN(n13104) );
  OR2_X1 U13196 ( .A1(n13232), .A2(n13233), .ZN(n13103) );
  AND2_X1 U13197 ( .A1(n13100), .A2(n13099), .ZN(n13233) );
  AND2_X1 U13198 ( .A1(n13097), .A2(n13234), .ZN(n13232) );
  OR2_X1 U13199 ( .A1(n13099), .A2(n13100), .ZN(n13234) );
  OR2_X1 U13200 ( .A1(n8579), .A2(n12831), .ZN(n13100) );
  OR2_X1 U13201 ( .A1(n13235), .A2(n13236), .ZN(n13099) );
  AND2_X1 U13202 ( .A1(n13096), .A2(n13095), .ZN(n13236) );
  AND2_X1 U13203 ( .A1(n13093), .A2(n13237), .ZN(n13235) );
  OR2_X1 U13204 ( .A1(n13095), .A2(n13096), .ZN(n13237) );
  OR2_X1 U13205 ( .A1(n8574), .A2(n12831), .ZN(n13096) );
  OR2_X1 U13206 ( .A1(n13238), .A2(n13239), .ZN(n13095) );
  AND2_X1 U13207 ( .A1(n13087), .A2(n13090), .ZN(n13239) );
  AND2_X1 U13208 ( .A1(n13240), .A2(n13089), .ZN(n13238) );
  OR2_X1 U13209 ( .A1(n13241), .A2(n13242), .ZN(n13089) );
  AND2_X1 U13210 ( .A1(n13086), .A2(n13085), .ZN(n13242) );
  AND2_X1 U13211 ( .A1(n13083), .A2(n13243), .ZN(n13241) );
  OR2_X1 U13212 ( .A1(n13085), .A2(n13086), .ZN(n13243) );
  OR2_X1 U13213 ( .A1(n8564), .A2(n12831), .ZN(n13086) );
  OR2_X1 U13214 ( .A1(n13244), .A2(n13245), .ZN(n13085) );
  AND2_X1 U13215 ( .A1(n13079), .A2(n13082), .ZN(n13245) );
  AND2_X1 U13216 ( .A1(n13246), .A2(n13081), .ZN(n13244) );
  OR2_X1 U13217 ( .A1(n13247), .A2(n13248), .ZN(n13081) );
  AND2_X1 U13218 ( .A1(n13075), .A2(n13078), .ZN(n13248) );
  AND2_X1 U13219 ( .A1(n13249), .A2(n13077), .ZN(n13247) );
  OR2_X1 U13220 ( .A1(n13250), .A2(n13251), .ZN(n13077) );
  AND2_X1 U13221 ( .A1(n13071), .A2(n13074), .ZN(n13251) );
  AND2_X1 U13222 ( .A1(n13252), .A2(n13073), .ZN(n13250) );
  OR2_X1 U13223 ( .A1(n13253), .A2(n13254), .ZN(n13073) );
  AND2_X1 U13224 ( .A1(n13067), .A2(n13070), .ZN(n13254) );
  AND2_X1 U13225 ( .A1(n13255), .A2(n13069), .ZN(n13253) );
  OR2_X1 U13226 ( .A1(n13256), .A2(n13257), .ZN(n13069) );
  AND2_X1 U13227 ( .A1(n13063), .A2(n13066), .ZN(n13257) );
  AND2_X1 U13228 ( .A1(n13258), .A2(n13065), .ZN(n13256) );
  OR2_X1 U13229 ( .A1(n13259), .A2(n13260), .ZN(n13065) );
  AND2_X1 U13230 ( .A1(n13059), .A2(n13062), .ZN(n13260) );
  AND2_X1 U13231 ( .A1(n13261), .A2(n13061), .ZN(n13259) );
  OR2_X1 U13232 ( .A1(n13262), .A2(n13263), .ZN(n13061) );
  AND2_X1 U13233 ( .A1(n13055), .A2(n13058), .ZN(n13263) );
  AND2_X1 U13234 ( .A1(n13264), .A2(n13057), .ZN(n13262) );
  OR2_X1 U13235 ( .A1(n13265), .A2(n13266), .ZN(n13057) );
  AND2_X1 U13236 ( .A1(n13051), .A2(n13054), .ZN(n13266) );
  AND2_X1 U13237 ( .A1(n13053), .A2(n13267), .ZN(n13265) );
  OR2_X1 U13238 ( .A1(n13054), .A2(n13051), .ZN(n13267) );
  OR2_X1 U13239 ( .A1(n12831), .A2(n8518), .ZN(n13051) );
  OR3_X1 U13240 ( .A1(n13050), .A2(n12831), .A3(n8519), .ZN(n13054) );
  INV_X1 U13241 ( .A(n13268), .ZN(n13053) );
  OR2_X1 U13242 ( .A1(n13269), .A2(n13270), .ZN(n13268) );
  AND2_X1 U13243 ( .A1(n13271), .A2(n13272), .ZN(n13270) );
  OR2_X1 U13244 ( .A1(n13273), .A2(n7697), .ZN(n13272) );
  AND2_X1 U13245 ( .A1(n13050), .A2(n7691), .ZN(n13273) );
  AND2_X1 U13246 ( .A1(n13045), .A2(n13274), .ZN(n13269) );
  OR2_X1 U13247 ( .A1(n13275), .A2(n7701), .ZN(n13274) );
  AND2_X1 U13248 ( .A1(n8123), .A2(n7703), .ZN(n13275) );
  OR2_X1 U13249 ( .A1(n13058), .A2(n13055), .ZN(n13264) );
  XNOR2_X1 U13250 ( .A(n13276), .B(n13277), .ZN(n13055) );
  XNOR2_X1 U13251 ( .A(n13278), .B(n13279), .ZN(n13277) );
  OR2_X1 U13252 ( .A1(n8529), .A2(n12831), .ZN(n13058) );
  OR2_X1 U13253 ( .A1(n13062), .A2(n13059), .ZN(n13261) );
  XOR2_X1 U13254 ( .A(n13280), .B(n13281), .Z(n13059) );
  XOR2_X1 U13255 ( .A(n13282), .B(n13283), .Z(n13281) );
  OR2_X1 U13256 ( .A1(n8534), .A2(n12831), .ZN(n13062) );
  OR2_X1 U13257 ( .A1(n13066), .A2(n13063), .ZN(n13258) );
  XOR2_X1 U13258 ( .A(n13284), .B(n13285), .Z(n13063) );
  XOR2_X1 U13259 ( .A(n13286), .B(n13287), .Z(n13285) );
  OR2_X1 U13260 ( .A1(n8539), .A2(n12831), .ZN(n13066) );
  OR2_X1 U13261 ( .A1(n13070), .A2(n13067), .ZN(n13255) );
  XOR2_X1 U13262 ( .A(n13288), .B(n13289), .Z(n13067) );
  XOR2_X1 U13263 ( .A(n13290), .B(n13291), .Z(n13289) );
  OR2_X1 U13264 ( .A1(n8544), .A2(n12831), .ZN(n13070) );
  OR2_X1 U13265 ( .A1(n13074), .A2(n13071), .ZN(n13252) );
  XOR2_X1 U13266 ( .A(n13292), .B(n13293), .Z(n13071) );
  XOR2_X1 U13267 ( .A(n13294), .B(n13295), .Z(n13293) );
  OR2_X1 U13268 ( .A1(n8549), .A2(n12831), .ZN(n13074) );
  OR2_X1 U13269 ( .A1(n13078), .A2(n13075), .ZN(n13249) );
  XOR2_X1 U13270 ( .A(n13296), .B(n13297), .Z(n13075) );
  XOR2_X1 U13271 ( .A(n13298), .B(n13299), .Z(n13297) );
  OR2_X1 U13272 ( .A1(n8554), .A2(n12831), .ZN(n13078) );
  OR2_X1 U13273 ( .A1(n13082), .A2(n13079), .ZN(n13246) );
  XOR2_X1 U13274 ( .A(n13300), .B(n13301), .Z(n13079) );
  XOR2_X1 U13275 ( .A(n13302), .B(n13303), .Z(n13301) );
  OR2_X1 U13276 ( .A1(n8559), .A2(n12831), .ZN(n13082) );
  XOR2_X1 U13277 ( .A(n13304), .B(n13305), .Z(n13083) );
  XOR2_X1 U13278 ( .A(n13306), .B(n13307), .Z(n13305) );
  OR2_X1 U13279 ( .A1(n13090), .A2(n13087), .ZN(n13240) );
  XOR2_X1 U13280 ( .A(n13308), .B(n13309), .Z(n13087) );
  XOR2_X1 U13281 ( .A(n13310), .B(n13311), .Z(n13309) );
  OR2_X1 U13282 ( .A1(n8569), .A2(n12831), .ZN(n13090) );
  INV_X1 U13283 ( .A(n12826), .ZN(n12831) );
  XOR2_X1 U13284 ( .A(n13312), .B(n13313), .Z(n12826) );
  XNOR2_X1 U13285 ( .A(c_9_), .B(d_9_), .ZN(n13312) );
  XOR2_X1 U13286 ( .A(n13314), .B(n13315), .Z(n13093) );
  XOR2_X1 U13287 ( .A(n13316), .B(n13317), .Z(n13315) );
  XOR2_X1 U13288 ( .A(n13318), .B(n13319), .Z(n13097) );
  XOR2_X1 U13289 ( .A(n13320), .B(n13321), .Z(n13319) );
  XOR2_X1 U13290 ( .A(n13322), .B(n13323), .Z(n13101) );
  XOR2_X1 U13291 ( .A(n13324), .B(n13325), .Z(n13323) );
  XNOR2_X1 U13292 ( .A(n13326), .B(n13327), .ZN(n13106) );
  XNOR2_X1 U13293 ( .A(n13328), .B(n13329), .ZN(n13326) );
  XNOR2_X1 U13294 ( .A(n13330), .B(n13331), .ZN(n13110) );
  XNOR2_X1 U13295 ( .A(n13332), .B(n13333), .ZN(n13330) );
  XOR2_X1 U13296 ( .A(n13334), .B(n13335), .Z(n13114) );
  XOR2_X1 U13297 ( .A(n13336), .B(n13337), .Z(n13335) );
  XOR2_X1 U13298 ( .A(n13338), .B(n13339), .Z(n13117) );
  XOR2_X1 U13299 ( .A(n13340), .B(n13341), .Z(n13339) );
  XOR2_X1 U13300 ( .A(n13342), .B(n13343), .Z(n13121) );
  XOR2_X1 U13301 ( .A(n13344), .B(n13345), .Z(n13343) );
  XOR2_X1 U13302 ( .A(n13346), .B(n13347), .Z(n13125) );
  XOR2_X1 U13303 ( .A(n13348), .B(n13349), .Z(n13347) );
  XOR2_X1 U13304 ( .A(n13350), .B(n13351), .Z(n13129) );
  XOR2_X1 U13305 ( .A(n13352), .B(n13353), .Z(n13351) );
  XOR2_X1 U13306 ( .A(n13354), .B(n13355), .Z(n13133) );
  XOR2_X1 U13307 ( .A(n13356), .B(n13357), .Z(n13355) );
  XOR2_X1 U13308 ( .A(n13358), .B(n13359), .Z(n13137) );
  XOR2_X1 U13309 ( .A(n13360), .B(n13361), .Z(n13359) );
  XOR2_X1 U13310 ( .A(n13362), .B(n13363), .Z(n13141) );
  XOR2_X1 U13311 ( .A(n13364), .B(n13365), .Z(n13363) );
  XOR2_X1 U13312 ( .A(n13366), .B(n13367), .Z(n13145) );
  XOR2_X1 U13313 ( .A(n13368), .B(n13369), .Z(n13367) );
  XOR2_X1 U13314 ( .A(n13370), .B(n13371), .Z(n13149) );
  XOR2_X1 U13315 ( .A(n13372), .B(n13373), .Z(n13371) );
  XOR2_X1 U13316 ( .A(n13374), .B(n13375), .Z(n13153) );
  XOR2_X1 U13317 ( .A(n13376), .B(n13377), .Z(n13375) );
  XOR2_X1 U13318 ( .A(n13378), .B(n13379), .Z(n13157) );
  XOR2_X1 U13319 ( .A(n13380), .B(n13381), .Z(n13379) );
  XOR2_X1 U13320 ( .A(n13382), .B(n13383), .Z(n13161) );
  XOR2_X1 U13321 ( .A(n13384), .B(n13385), .Z(n13383) );
  XOR2_X1 U13322 ( .A(n13386), .B(n13387), .Z(n13165) );
  XOR2_X1 U13323 ( .A(n13388), .B(n13389), .Z(n13387) );
  XOR2_X1 U13324 ( .A(n13390), .B(n13391), .Z(n13169) );
  XOR2_X1 U13325 ( .A(n13392), .B(n13393), .Z(n13391) );
  XOR2_X1 U13326 ( .A(n8120), .B(n13394), .Z(n13176) );
  XOR2_X1 U13327 ( .A(n8119), .B(n8118), .Z(n13394) );
  OR2_X1 U13328 ( .A1(n13050), .A2(n7960), .ZN(n8118) );
  OR2_X1 U13329 ( .A1(n13395), .A2(n13396), .ZN(n8119) );
  AND2_X1 U13330 ( .A1(n13393), .A2(n13392), .ZN(n13396) );
  AND2_X1 U13331 ( .A1(n13390), .A2(n13397), .ZN(n13395) );
  OR2_X1 U13332 ( .A1(n13392), .A2(n13393), .ZN(n13397) );
  OR2_X1 U13333 ( .A1(n13050), .A2(n7608), .ZN(n13393) );
  OR2_X1 U13334 ( .A1(n13398), .A2(n13399), .ZN(n13392) );
  AND2_X1 U13335 ( .A1(n13389), .A2(n13388), .ZN(n13399) );
  AND2_X1 U13336 ( .A1(n13386), .A2(n13400), .ZN(n13398) );
  OR2_X1 U13337 ( .A1(n13388), .A2(n13389), .ZN(n13400) );
  OR2_X1 U13338 ( .A1(n13050), .A2(n7610), .ZN(n13389) );
  OR2_X1 U13339 ( .A1(n13401), .A2(n13402), .ZN(n13388) );
  AND2_X1 U13340 ( .A1(n13385), .A2(n13384), .ZN(n13402) );
  AND2_X1 U13341 ( .A1(n13382), .A2(n13403), .ZN(n13401) );
  OR2_X1 U13342 ( .A1(n13384), .A2(n13385), .ZN(n13403) );
  OR2_X1 U13343 ( .A1(n13050), .A2(n7612), .ZN(n13385) );
  OR2_X1 U13344 ( .A1(n13404), .A2(n13405), .ZN(n13384) );
  AND2_X1 U13345 ( .A1(n13381), .A2(n13380), .ZN(n13405) );
  AND2_X1 U13346 ( .A1(n13378), .A2(n13406), .ZN(n13404) );
  OR2_X1 U13347 ( .A1(n13380), .A2(n13381), .ZN(n13406) );
  OR2_X1 U13348 ( .A1(n13050), .A2(n7614), .ZN(n13381) );
  OR2_X1 U13349 ( .A1(n13407), .A2(n13408), .ZN(n13380) );
  AND2_X1 U13350 ( .A1(n13377), .A2(n13376), .ZN(n13408) );
  AND2_X1 U13351 ( .A1(n13374), .A2(n13409), .ZN(n13407) );
  OR2_X1 U13352 ( .A1(n13376), .A2(n13377), .ZN(n13409) );
  OR2_X1 U13353 ( .A1(n13050), .A2(n7616), .ZN(n13377) );
  OR2_X1 U13354 ( .A1(n13410), .A2(n13411), .ZN(n13376) );
  AND2_X1 U13355 ( .A1(n13373), .A2(n13372), .ZN(n13411) );
  AND2_X1 U13356 ( .A1(n13370), .A2(n13412), .ZN(n13410) );
  OR2_X1 U13357 ( .A1(n13372), .A2(n13373), .ZN(n13412) );
  OR2_X1 U13358 ( .A1(n13050), .A2(n7618), .ZN(n13373) );
  OR2_X1 U13359 ( .A1(n13413), .A2(n13414), .ZN(n13372) );
  AND2_X1 U13360 ( .A1(n13369), .A2(n13368), .ZN(n13414) );
  AND2_X1 U13361 ( .A1(n13366), .A2(n13415), .ZN(n13413) );
  OR2_X1 U13362 ( .A1(n13368), .A2(n13369), .ZN(n13415) );
  OR2_X1 U13363 ( .A1(n8634), .A2(n13050), .ZN(n13369) );
  OR2_X1 U13364 ( .A1(n13416), .A2(n13417), .ZN(n13368) );
  AND2_X1 U13365 ( .A1(n13365), .A2(n13364), .ZN(n13417) );
  AND2_X1 U13366 ( .A1(n13362), .A2(n13418), .ZN(n13416) );
  OR2_X1 U13367 ( .A1(n13364), .A2(n13365), .ZN(n13418) );
  OR2_X1 U13368 ( .A1(n8629), .A2(n13050), .ZN(n13365) );
  OR2_X1 U13369 ( .A1(n13419), .A2(n13420), .ZN(n13364) );
  AND2_X1 U13370 ( .A1(n13361), .A2(n13360), .ZN(n13420) );
  AND2_X1 U13371 ( .A1(n13358), .A2(n13421), .ZN(n13419) );
  OR2_X1 U13372 ( .A1(n13360), .A2(n13361), .ZN(n13421) );
  OR2_X1 U13373 ( .A1(n8624), .A2(n13050), .ZN(n13361) );
  OR2_X1 U13374 ( .A1(n13422), .A2(n13423), .ZN(n13360) );
  AND2_X1 U13375 ( .A1(n13357), .A2(n13356), .ZN(n13423) );
  AND2_X1 U13376 ( .A1(n13354), .A2(n13424), .ZN(n13422) );
  OR2_X1 U13377 ( .A1(n13356), .A2(n13357), .ZN(n13424) );
  OR2_X1 U13378 ( .A1(n8619), .A2(n13050), .ZN(n13357) );
  OR2_X1 U13379 ( .A1(n13425), .A2(n13426), .ZN(n13356) );
  AND2_X1 U13380 ( .A1(n13353), .A2(n13352), .ZN(n13426) );
  AND2_X1 U13381 ( .A1(n13350), .A2(n13427), .ZN(n13425) );
  OR2_X1 U13382 ( .A1(n13352), .A2(n13353), .ZN(n13427) );
  OR2_X1 U13383 ( .A1(n8614), .A2(n13050), .ZN(n13353) );
  OR2_X1 U13384 ( .A1(n13428), .A2(n13429), .ZN(n13352) );
  AND2_X1 U13385 ( .A1(n13349), .A2(n13348), .ZN(n13429) );
  AND2_X1 U13386 ( .A1(n13346), .A2(n13430), .ZN(n13428) );
  OR2_X1 U13387 ( .A1(n13348), .A2(n13349), .ZN(n13430) );
  OR2_X1 U13388 ( .A1(n8609), .A2(n13050), .ZN(n13349) );
  OR2_X1 U13389 ( .A1(n13431), .A2(n13432), .ZN(n13348) );
  AND2_X1 U13390 ( .A1(n13345), .A2(n13344), .ZN(n13432) );
  AND2_X1 U13391 ( .A1(n13342), .A2(n13433), .ZN(n13431) );
  OR2_X1 U13392 ( .A1(n13344), .A2(n13345), .ZN(n13433) );
  OR2_X1 U13393 ( .A1(n8604), .A2(n13050), .ZN(n13345) );
  OR2_X1 U13394 ( .A1(n13434), .A2(n13435), .ZN(n13344) );
  AND2_X1 U13395 ( .A1(n13341), .A2(n13340), .ZN(n13435) );
  AND2_X1 U13396 ( .A1(n13338), .A2(n13436), .ZN(n13434) );
  OR2_X1 U13397 ( .A1(n13340), .A2(n13341), .ZN(n13436) );
  OR2_X1 U13398 ( .A1(n8599), .A2(n13050), .ZN(n13341) );
  OR2_X1 U13399 ( .A1(n13437), .A2(n13438), .ZN(n13340) );
  AND2_X1 U13400 ( .A1(n13337), .A2(n13336), .ZN(n13438) );
  AND2_X1 U13401 ( .A1(n13334), .A2(n13439), .ZN(n13437) );
  OR2_X1 U13402 ( .A1(n13336), .A2(n13337), .ZN(n13439) );
  OR2_X1 U13403 ( .A1(n8594), .A2(n13050), .ZN(n13337) );
  OR2_X1 U13404 ( .A1(n13440), .A2(n13441), .ZN(n13336) );
  AND2_X1 U13405 ( .A1(n13333), .A2(n13332), .ZN(n13441) );
  AND2_X1 U13406 ( .A1(n13331), .A2(n13442), .ZN(n13440) );
  OR2_X1 U13407 ( .A1(n13332), .A2(n13333), .ZN(n13442) );
  OR2_X1 U13408 ( .A1(n8589), .A2(n13050), .ZN(n13333) );
  OR2_X1 U13409 ( .A1(n13443), .A2(n13444), .ZN(n13332) );
  AND2_X1 U13410 ( .A1(n13329), .A2(n13328), .ZN(n13444) );
  AND2_X1 U13411 ( .A1(n13327), .A2(n13445), .ZN(n13443) );
  OR2_X1 U13412 ( .A1(n13328), .A2(n13329), .ZN(n13445) );
  OR2_X1 U13413 ( .A1(n8584), .A2(n13050), .ZN(n13329) );
  OR2_X1 U13414 ( .A1(n13446), .A2(n13447), .ZN(n13328) );
  AND2_X1 U13415 ( .A1(n13325), .A2(n13324), .ZN(n13447) );
  AND2_X1 U13416 ( .A1(n13322), .A2(n13448), .ZN(n13446) );
  OR2_X1 U13417 ( .A1(n13324), .A2(n13325), .ZN(n13448) );
  OR2_X1 U13418 ( .A1(n8579), .A2(n13050), .ZN(n13325) );
  OR2_X1 U13419 ( .A1(n13449), .A2(n13450), .ZN(n13324) );
  AND2_X1 U13420 ( .A1(n13321), .A2(n13320), .ZN(n13450) );
  AND2_X1 U13421 ( .A1(n13318), .A2(n13451), .ZN(n13449) );
  OR2_X1 U13422 ( .A1(n13320), .A2(n13321), .ZN(n13451) );
  OR2_X1 U13423 ( .A1(n8574), .A2(n13050), .ZN(n13321) );
  OR2_X1 U13424 ( .A1(n13452), .A2(n13453), .ZN(n13320) );
  AND2_X1 U13425 ( .A1(n13317), .A2(n13316), .ZN(n13453) );
  AND2_X1 U13426 ( .A1(n13314), .A2(n13454), .ZN(n13452) );
  OR2_X1 U13427 ( .A1(n13316), .A2(n13317), .ZN(n13454) );
  OR2_X1 U13428 ( .A1(n8569), .A2(n13050), .ZN(n13317) );
  OR2_X1 U13429 ( .A1(n13455), .A2(n13456), .ZN(n13316) );
  AND2_X1 U13430 ( .A1(n13308), .A2(n13311), .ZN(n13456) );
  AND2_X1 U13431 ( .A1(n13457), .A2(n13310), .ZN(n13455) );
  OR2_X1 U13432 ( .A1(n13458), .A2(n13459), .ZN(n13310) );
  AND2_X1 U13433 ( .A1(n13307), .A2(n13306), .ZN(n13459) );
  AND2_X1 U13434 ( .A1(n13304), .A2(n13460), .ZN(n13458) );
  OR2_X1 U13435 ( .A1(n13306), .A2(n13307), .ZN(n13460) );
  OR2_X1 U13436 ( .A1(n8559), .A2(n13050), .ZN(n13307) );
  OR2_X1 U13437 ( .A1(n13461), .A2(n13462), .ZN(n13306) );
  AND2_X1 U13438 ( .A1(n13300), .A2(n13303), .ZN(n13462) );
  AND2_X1 U13439 ( .A1(n13463), .A2(n13302), .ZN(n13461) );
  OR2_X1 U13440 ( .A1(n13464), .A2(n13465), .ZN(n13302) );
  AND2_X1 U13441 ( .A1(n13296), .A2(n13299), .ZN(n13465) );
  AND2_X1 U13442 ( .A1(n13466), .A2(n13298), .ZN(n13464) );
  OR2_X1 U13443 ( .A1(n13467), .A2(n13468), .ZN(n13298) );
  AND2_X1 U13444 ( .A1(n13292), .A2(n13295), .ZN(n13468) );
  AND2_X1 U13445 ( .A1(n13469), .A2(n13294), .ZN(n13467) );
  OR2_X1 U13446 ( .A1(n13470), .A2(n13471), .ZN(n13294) );
  AND2_X1 U13447 ( .A1(n13288), .A2(n13291), .ZN(n13471) );
  AND2_X1 U13448 ( .A1(n13472), .A2(n13290), .ZN(n13470) );
  OR2_X1 U13449 ( .A1(n13473), .A2(n13474), .ZN(n13290) );
  AND2_X1 U13450 ( .A1(n13284), .A2(n13287), .ZN(n13474) );
  AND2_X1 U13451 ( .A1(n13475), .A2(n13286), .ZN(n13473) );
  OR2_X1 U13452 ( .A1(n13476), .A2(n13477), .ZN(n13286) );
  AND2_X1 U13453 ( .A1(n13280), .A2(n13283), .ZN(n13477) );
  AND2_X1 U13454 ( .A1(n13478), .A2(n13282), .ZN(n13476) );
  OR2_X1 U13455 ( .A1(n13479), .A2(n13480), .ZN(n13282) );
  AND2_X1 U13456 ( .A1(n13276), .A2(n13279), .ZN(n13480) );
  AND2_X1 U13457 ( .A1(n13278), .A2(n13481), .ZN(n13479) );
  OR2_X1 U13458 ( .A1(n13279), .A2(n13276), .ZN(n13481) );
  OR2_X1 U13459 ( .A1(n13050), .A2(n8518), .ZN(n13276) );
  OR3_X1 U13460 ( .A1(n8123), .A2(n13050), .A3(n8519), .ZN(n13279) );
  INV_X1 U13461 ( .A(n13482), .ZN(n13278) );
  OR2_X1 U13462 ( .A1(n13483), .A2(n13484), .ZN(n13482) );
  AND2_X1 U13463 ( .A1(n13485), .A2(n13486), .ZN(n13484) );
  OR2_X1 U13464 ( .A1(n13487), .A2(n7697), .ZN(n13486) );
  AND2_X1 U13465 ( .A1(n8123), .A2(n7691), .ZN(n13487) );
  AND2_X1 U13466 ( .A1(n13271), .A2(n13488), .ZN(n13483) );
  OR2_X1 U13467 ( .A1(n13489), .A2(n7701), .ZN(n13488) );
  AND2_X1 U13468 ( .A1(n8083), .A2(n7703), .ZN(n13489) );
  OR2_X1 U13469 ( .A1(n13283), .A2(n13280), .ZN(n13478) );
  XNOR2_X1 U13470 ( .A(n13490), .B(n13491), .ZN(n13280) );
  XNOR2_X1 U13471 ( .A(n13492), .B(n13493), .ZN(n13491) );
  OR2_X1 U13472 ( .A1(n8529), .A2(n13050), .ZN(n13283) );
  OR2_X1 U13473 ( .A1(n13287), .A2(n13284), .ZN(n13475) );
  XOR2_X1 U13474 ( .A(n13494), .B(n13495), .Z(n13284) );
  XOR2_X1 U13475 ( .A(n13496), .B(n13497), .Z(n13495) );
  OR2_X1 U13476 ( .A1(n8534), .A2(n13050), .ZN(n13287) );
  OR2_X1 U13477 ( .A1(n13291), .A2(n13288), .ZN(n13472) );
  XOR2_X1 U13478 ( .A(n13498), .B(n13499), .Z(n13288) );
  XOR2_X1 U13479 ( .A(n13500), .B(n13501), .Z(n13499) );
  OR2_X1 U13480 ( .A1(n8539), .A2(n13050), .ZN(n13291) );
  OR2_X1 U13481 ( .A1(n13295), .A2(n13292), .ZN(n13469) );
  XOR2_X1 U13482 ( .A(n13502), .B(n13503), .Z(n13292) );
  XOR2_X1 U13483 ( .A(n13504), .B(n13505), .Z(n13503) );
  OR2_X1 U13484 ( .A1(n8544), .A2(n13050), .ZN(n13295) );
  OR2_X1 U13485 ( .A1(n13299), .A2(n13296), .ZN(n13466) );
  XOR2_X1 U13486 ( .A(n13506), .B(n13507), .Z(n13296) );
  XOR2_X1 U13487 ( .A(n13508), .B(n13509), .Z(n13507) );
  OR2_X1 U13488 ( .A1(n8549), .A2(n13050), .ZN(n13299) );
  OR2_X1 U13489 ( .A1(n13303), .A2(n13300), .ZN(n13463) );
  XOR2_X1 U13490 ( .A(n13510), .B(n13511), .Z(n13300) );
  XOR2_X1 U13491 ( .A(n13512), .B(n13513), .Z(n13511) );
  OR2_X1 U13492 ( .A1(n8554), .A2(n13050), .ZN(n13303) );
  XOR2_X1 U13493 ( .A(n13514), .B(n13515), .Z(n13304) );
  XOR2_X1 U13494 ( .A(n13516), .B(n13517), .Z(n13515) );
  OR2_X1 U13495 ( .A1(n13311), .A2(n13308), .ZN(n13457) );
  XOR2_X1 U13496 ( .A(n13518), .B(n13519), .Z(n13308) );
  XOR2_X1 U13497 ( .A(n13520), .B(n13521), .Z(n13519) );
  OR2_X1 U13498 ( .A1(n8564), .A2(n13050), .ZN(n13311) );
  INV_X1 U13499 ( .A(n13045), .ZN(n13050) );
  XOR2_X1 U13500 ( .A(n13522), .B(n13523), .Z(n13045) );
  XNOR2_X1 U13501 ( .A(c_8_), .B(d_8_), .ZN(n13522) );
  XOR2_X1 U13502 ( .A(n13524), .B(n13525), .Z(n13314) );
  XOR2_X1 U13503 ( .A(n13526), .B(n13527), .Z(n13525) );
  XOR2_X1 U13504 ( .A(n13528), .B(n13529), .Z(n13318) );
  XOR2_X1 U13505 ( .A(n13530), .B(n13531), .Z(n13529) );
  XNOR2_X1 U13506 ( .A(n13532), .B(n13533), .ZN(n13322) );
  XNOR2_X1 U13507 ( .A(n13534), .B(n13535), .ZN(n13532) );
  XOR2_X1 U13508 ( .A(n13536), .B(n13537), .Z(n13327) );
  XOR2_X1 U13509 ( .A(n13538), .B(n13539), .Z(n13537) );
  XOR2_X1 U13510 ( .A(n13540), .B(n13541), .Z(n13331) );
  XOR2_X1 U13511 ( .A(n13542), .B(n13543), .Z(n13541) );
  XOR2_X1 U13512 ( .A(n13544), .B(n13545), .Z(n13334) );
  XOR2_X1 U13513 ( .A(n13546), .B(n13547), .Z(n13545) );
  XOR2_X1 U13514 ( .A(n13548), .B(n13549), .Z(n13338) );
  XOR2_X1 U13515 ( .A(n13550), .B(n13551), .Z(n13549) );
  XOR2_X1 U13516 ( .A(n13552), .B(n13553), .Z(n13342) );
  XOR2_X1 U13517 ( .A(n13554), .B(n13555), .Z(n13553) );
  XOR2_X1 U13518 ( .A(n13556), .B(n13557), .Z(n13346) );
  XOR2_X1 U13519 ( .A(n13558), .B(n13559), .Z(n13557) );
  XOR2_X1 U13520 ( .A(n13560), .B(n13561), .Z(n13350) );
  XOR2_X1 U13521 ( .A(n13562), .B(n13563), .Z(n13561) );
  XOR2_X1 U13522 ( .A(n13564), .B(n13565), .Z(n13354) );
  XOR2_X1 U13523 ( .A(n13566), .B(n13567), .Z(n13565) );
  XOR2_X1 U13524 ( .A(n13568), .B(n13569), .Z(n13358) );
  XOR2_X1 U13525 ( .A(n13570), .B(n13571), .Z(n13569) );
  XOR2_X1 U13526 ( .A(n13572), .B(n13573), .Z(n13362) );
  XOR2_X1 U13527 ( .A(n13574), .B(n13575), .Z(n13573) );
  XOR2_X1 U13528 ( .A(n13576), .B(n13577), .Z(n13366) );
  XOR2_X1 U13529 ( .A(n13578), .B(n13579), .Z(n13577) );
  XOR2_X1 U13530 ( .A(n13580), .B(n13581), .Z(n13370) );
  XOR2_X1 U13531 ( .A(n13582), .B(n13583), .Z(n13581) );
  XOR2_X1 U13532 ( .A(n13584), .B(n13585), .Z(n13374) );
  XOR2_X1 U13533 ( .A(n13586), .B(n13587), .Z(n13585) );
  XOR2_X1 U13534 ( .A(n13588), .B(n13589), .Z(n13378) );
  XOR2_X1 U13535 ( .A(n13590), .B(n13591), .Z(n13589) );
  XOR2_X1 U13536 ( .A(n13592), .B(n13593), .Z(n13382) );
  XOR2_X1 U13537 ( .A(n13594), .B(n13595), .Z(n13593) );
  XOR2_X1 U13538 ( .A(n13596), .B(n13597), .Z(n13386) );
  XOR2_X1 U13539 ( .A(n13598), .B(n13599), .Z(n13597) );
  XOR2_X1 U13540 ( .A(n13600), .B(n13601), .Z(n13390) );
  XOR2_X1 U13541 ( .A(n13602), .B(n13603), .Z(n13601) );
  XOR2_X1 U13542 ( .A(n8128), .B(n13604), .Z(n8120) );
  XOR2_X1 U13543 ( .A(n8127), .B(n8126), .Z(n13604) );
  OR2_X1 U13544 ( .A1(n8123), .A2(n7608), .ZN(n8126) );
  OR2_X1 U13545 ( .A1(n13605), .A2(n13606), .ZN(n8127) );
  AND2_X1 U13546 ( .A1(n13603), .A2(n13602), .ZN(n13606) );
  AND2_X1 U13547 ( .A1(n13600), .A2(n13607), .ZN(n13605) );
  OR2_X1 U13548 ( .A1(n13602), .A2(n13603), .ZN(n13607) );
  OR2_X1 U13549 ( .A1(n8123), .A2(n7610), .ZN(n13603) );
  OR2_X1 U13550 ( .A1(n13608), .A2(n13609), .ZN(n13602) );
  AND2_X1 U13551 ( .A1(n13599), .A2(n13598), .ZN(n13609) );
  AND2_X1 U13552 ( .A1(n13596), .A2(n13610), .ZN(n13608) );
  OR2_X1 U13553 ( .A1(n13598), .A2(n13599), .ZN(n13610) );
  OR2_X1 U13554 ( .A1(n8123), .A2(n7612), .ZN(n13599) );
  OR2_X1 U13555 ( .A1(n13611), .A2(n13612), .ZN(n13598) );
  AND2_X1 U13556 ( .A1(n13595), .A2(n13594), .ZN(n13612) );
  AND2_X1 U13557 ( .A1(n13592), .A2(n13613), .ZN(n13611) );
  OR2_X1 U13558 ( .A1(n13594), .A2(n13595), .ZN(n13613) );
  OR2_X1 U13559 ( .A1(n8123), .A2(n7614), .ZN(n13595) );
  OR2_X1 U13560 ( .A1(n13614), .A2(n13615), .ZN(n13594) );
  AND2_X1 U13561 ( .A1(n13591), .A2(n13590), .ZN(n13615) );
  AND2_X1 U13562 ( .A1(n13588), .A2(n13616), .ZN(n13614) );
  OR2_X1 U13563 ( .A1(n13590), .A2(n13591), .ZN(n13616) );
  OR2_X1 U13564 ( .A1(n8123), .A2(n7616), .ZN(n13591) );
  OR2_X1 U13565 ( .A1(n13617), .A2(n13618), .ZN(n13590) );
  AND2_X1 U13566 ( .A1(n13587), .A2(n13586), .ZN(n13618) );
  AND2_X1 U13567 ( .A1(n13584), .A2(n13619), .ZN(n13617) );
  OR2_X1 U13568 ( .A1(n13586), .A2(n13587), .ZN(n13619) );
  OR2_X1 U13569 ( .A1(n8123), .A2(n7618), .ZN(n13587) );
  OR2_X1 U13570 ( .A1(n13620), .A2(n13621), .ZN(n13586) );
  AND2_X1 U13571 ( .A1(n13583), .A2(n13582), .ZN(n13621) );
  AND2_X1 U13572 ( .A1(n13580), .A2(n13622), .ZN(n13620) );
  OR2_X1 U13573 ( .A1(n13582), .A2(n13583), .ZN(n13622) );
  OR2_X1 U13574 ( .A1(n8123), .A2(n7620), .ZN(n13583) );
  OR2_X1 U13575 ( .A1(n13623), .A2(n13624), .ZN(n13582) );
  AND2_X1 U13576 ( .A1(n13579), .A2(n13578), .ZN(n13624) );
  AND2_X1 U13577 ( .A1(n13576), .A2(n13625), .ZN(n13623) );
  OR2_X1 U13578 ( .A1(n13578), .A2(n13579), .ZN(n13625) );
  OR2_X1 U13579 ( .A1(n8629), .A2(n8123), .ZN(n13579) );
  OR2_X1 U13580 ( .A1(n13626), .A2(n13627), .ZN(n13578) );
  AND2_X1 U13581 ( .A1(n13575), .A2(n13574), .ZN(n13627) );
  AND2_X1 U13582 ( .A1(n13572), .A2(n13628), .ZN(n13626) );
  OR2_X1 U13583 ( .A1(n13574), .A2(n13575), .ZN(n13628) );
  OR2_X1 U13584 ( .A1(n8624), .A2(n8123), .ZN(n13575) );
  OR2_X1 U13585 ( .A1(n13629), .A2(n13630), .ZN(n13574) );
  AND2_X1 U13586 ( .A1(n13571), .A2(n13570), .ZN(n13630) );
  AND2_X1 U13587 ( .A1(n13568), .A2(n13631), .ZN(n13629) );
  OR2_X1 U13588 ( .A1(n13570), .A2(n13571), .ZN(n13631) );
  OR2_X1 U13589 ( .A1(n8619), .A2(n8123), .ZN(n13571) );
  OR2_X1 U13590 ( .A1(n13632), .A2(n13633), .ZN(n13570) );
  AND2_X1 U13591 ( .A1(n13567), .A2(n13566), .ZN(n13633) );
  AND2_X1 U13592 ( .A1(n13564), .A2(n13634), .ZN(n13632) );
  OR2_X1 U13593 ( .A1(n13566), .A2(n13567), .ZN(n13634) );
  OR2_X1 U13594 ( .A1(n8614), .A2(n8123), .ZN(n13567) );
  OR2_X1 U13595 ( .A1(n13635), .A2(n13636), .ZN(n13566) );
  AND2_X1 U13596 ( .A1(n13563), .A2(n13562), .ZN(n13636) );
  AND2_X1 U13597 ( .A1(n13560), .A2(n13637), .ZN(n13635) );
  OR2_X1 U13598 ( .A1(n13562), .A2(n13563), .ZN(n13637) );
  OR2_X1 U13599 ( .A1(n8609), .A2(n8123), .ZN(n13563) );
  OR2_X1 U13600 ( .A1(n13638), .A2(n13639), .ZN(n13562) );
  AND2_X1 U13601 ( .A1(n13559), .A2(n13558), .ZN(n13639) );
  AND2_X1 U13602 ( .A1(n13556), .A2(n13640), .ZN(n13638) );
  OR2_X1 U13603 ( .A1(n13558), .A2(n13559), .ZN(n13640) );
  OR2_X1 U13604 ( .A1(n8604), .A2(n8123), .ZN(n13559) );
  OR2_X1 U13605 ( .A1(n13641), .A2(n13642), .ZN(n13558) );
  AND2_X1 U13606 ( .A1(n13555), .A2(n13554), .ZN(n13642) );
  AND2_X1 U13607 ( .A1(n13552), .A2(n13643), .ZN(n13641) );
  OR2_X1 U13608 ( .A1(n13554), .A2(n13555), .ZN(n13643) );
  OR2_X1 U13609 ( .A1(n8599), .A2(n8123), .ZN(n13555) );
  OR2_X1 U13610 ( .A1(n13644), .A2(n13645), .ZN(n13554) );
  AND2_X1 U13611 ( .A1(n13551), .A2(n13550), .ZN(n13645) );
  AND2_X1 U13612 ( .A1(n13548), .A2(n13646), .ZN(n13644) );
  OR2_X1 U13613 ( .A1(n13550), .A2(n13551), .ZN(n13646) );
  OR2_X1 U13614 ( .A1(n8594), .A2(n8123), .ZN(n13551) );
  OR2_X1 U13615 ( .A1(n13647), .A2(n13648), .ZN(n13550) );
  AND2_X1 U13616 ( .A1(n13547), .A2(n13546), .ZN(n13648) );
  AND2_X1 U13617 ( .A1(n13544), .A2(n13649), .ZN(n13647) );
  OR2_X1 U13618 ( .A1(n13546), .A2(n13547), .ZN(n13649) );
  OR2_X1 U13619 ( .A1(n8589), .A2(n8123), .ZN(n13547) );
  OR2_X1 U13620 ( .A1(n13650), .A2(n13651), .ZN(n13546) );
  AND2_X1 U13621 ( .A1(n13543), .A2(n13542), .ZN(n13651) );
  AND2_X1 U13622 ( .A1(n13540), .A2(n13652), .ZN(n13650) );
  OR2_X1 U13623 ( .A1(n13542), .A2(n13543), .ZN(n13652) );
  OR2_X1 U13624 ( .A1(n8584), .A2(n8123), .ZN(n13543) );
  OR2_X1 U13625 ( .A1(n13653), .A2(n13654), .ZN(n13542) );
  AND2_X1 U13626 ( .A1(n13539), .A2(n13538), .ZN(n13654) );
  AND2_X1 U13627 ( .A1(n13536), .A2(n13655), .ZN(n13653) );
  OR2_X1 U13628 ( .A1(n13538), .A2(n13539), .ZN(n13655) );
  OR2_X1 U13629 ( .A1(n8579), .A2(n8123), .ZN(n13539) );
  OR2_X1 U13630 ( .A1(n13656), .A2(n13657), .ZN(n13538) );
  AND2_X1 U13631 ( .A1(n13535), .A2(n13534), .ZN(n13657) );
  AND2_X1 U13632 ( .A1(n13533), .A2(n13658), .ZN(n13656) );
  OR2_X1 U13633 ( .A1(n13534), .A2(n13535), .ZN(n13658) );
  OR2_X1 U13634 ( .A1(n8574), .A2(n8123), .ZN(n13535) );
  OR2_X1 U13635 ( .A1(n13659), .A2(n13660), .ZN(n13534) );
  AND2_X1 U13636 ( .A1(n13531), .A2(n13530), .ZN(n13660) );
  AND2_X1 U13637 ( .A1(n13528), .A2(n13661), .ZN(n13659) );
  OR2_X1 U13638 ( .A1(n13530), .A2(n13531), .ZN(n13661) );
  OR2_X1 U13639 ( .A1(n8569), .A2(n8123), .ZN(n13531) );
  OR2_X1 U13640 ( .A1(n13662), .A2(n13663), .ZN(n13530) );
  AND2_X1 U13641 ( .A1(n13527), .A2(n13526), .ZN(n13663) );
  AND2_X1 U13642 ( .A1(n13524), .A2(n13664), .ZN(n13662) );
  OR2_X1 U13643 ( .A1(n13526), .A2(n13527), .ZN(n13664) );
  OR2_X1 U13644 ( .A1(n8564), .A2(n8123), .ZN(n13527) );
  OR2_X1 U13645 ( .A1(n13665), .A2(n13666), .ZN(n13526) );
  AND2_X1 U13646 ( .A1(n13518), .A2(n13521), .ZN(n13666) );
  AND2_X1 U13647 ( .A1(n13667), .A2(n13520), .ZN(n13665) );
  OR2_X1 U13648 ( .A1(n13668), .A2(n13669), .ZN(n13520) );
  AND2_X1 U13649 ( .A1(n13517), .A2(n13516), .ZN(n13669) );
  AND2_X1 U13650 ( .A1(n13514), .A2(n13670), .ZN(n13668) );
  OR2_X1 U13651 ( .A1(n13516), .A2(n13517), .ZN(n13670) );
  OR2_X1 U13652 ( .A1(n8554), .A2(n8123), .ZN(n13517) );
  OR2_X1 U13653 ( .A1(n13671), .A2(n13672), .ZN(n13516) );
  AND2_X1 U13654 ( .A1(n13510), .A2(n13513), .ZN(n13672) );
  AND2_X1 U13655 ( .A1(n13673), .A2(n13512), .ZN(n13671) );
  OR2_X1 U13656 ( .A1(n13674), .A2(n13675), .ZN(n13512) );
  AND2_X1 U13657 ( .A1(n13506), .A2(n13509), .ZN(n13675) );
  AND2_X1 U13658 ( .A1(n13676), .A2(n13508), .ZN(n13674) );
  OR2_X1 U13659 ( .A1(n13677), .A2(n13678), .ZN(n13508) );
  AND2_X1 U13660 ( .A1(n13502), .A2(n13505), .ZN(n13678) );
  AND2_X1 U13661 ( .A1(n13679), .A2(n13504), .ZN(n13677) );
  OR2_X1 U13662 ( .A1(n13680), .A2(n13681), .ZN(n13504) );
  AND2_X1 U13663 ( .A1(n13498), .A2(n13501), .ZN(n13681) );
  AND2_X1 U13664 ( .A1(n13682), .A2(n13500), .ZN(n13680) );
  OR2_X1 U13665 ( .A1(n13683), .A2(n13684), .ZN(n13500) );
  AND2_X1 U13666 ( .A1(n13494), .A2(n13497), .ZN(n13684) );
  AND2_X1 U13667 ( .A1(n13685), .A2(n13496), .ZN(n13683) );
  OR2_X1 U13668 ( .A1(n13686), .A2(n13687), .ZN(n13496) );
  AND2_X1 U13669 ( .A1(n13490), .A2(n13493), .ZN(n13687) );
  AND2_X1 U13670 ( .A1(n13492), .A2(n13688), .ZN(n13686) );
  OR2_X1 U13671 ( .A1(n13493), .A2(n13490), .ZN(n13688) );
  OR2_X1 U13672 ( .A1(n8123), .A2(n8518), .ZN(n13490) );
  OR3_X1 U13673 ( .A1(n8083), .A2(n8123), .A3(n8519), .ZN(n13493) );
  INV_X1 U13674 ( .A(n13689), .ZN(n13492) );
  OR2_X1 U13675 ( .A1(n13690), .A2(n13691), .ZN(n13689) );
  AND2_X1 U13676 ( .A1(n13692), .A2(n13693), .ZN(n13691) );
  OR2_X1 U13677 ( .A1(n13694), .A2(n7697), .ZN(n13693) );
  AND2_X1 U13678 ( .A1(n8083), .A2(n7691), .ZN(n13694) );
  AND2_X1 U13679 ( .A1(n13485), .A2(n13695), .ZN(n13690) );
  OR2_X1 U13680 ( .A1(n13696), .A2(n7701), .ZN(n13695) );
  AND2_X1 U13681 ( .A1(n8041), .A2(n7703), .ZN(n13696) );
  OR2_X1 U13682 ( .A1(n13497), .A2(n13494), .ZN(n13685) );
  XNOR2_X1 U13683 ( .A(n13697), .B(n13698), .ZN(n13494) );
  XNOR2_X1 U13684 ( .A(n13699), .B(n13700), .ZN(n13698) );
  OR2_X1 U13685 ( .A1(n8529), .A2(n8123), .ZN(n13497) );
  OR2_X1 U13686 ( .A1(n13501), .A2(n13498), .ZN(n13682) );
  XOR2_X1 U13687 ( .A(n13701), .B(n13702), .Z(n13498) );
  XOR2_X1 U13688 ( .A(n13703), .B(n13704), .Z(n13702) );
  OR2_X1 U13689 ( .A1(n8534), .A2(n8123), .ZN(n13501) );
  OR2_X1 U13690 ( .A1(n13505), .A2(n13502), .ZN(n13679) );
  XOR2_X1 U13691 ( .A(n13705), .B(n13706), .Z(n13502) );
  XOR2_X1 U13692 ( .A(n13707), .B(n13708), .Z(n13706) );
  OR2_X1 U13693 ( .A1(n8539), .A2(n8123), .ZN(n13505) );
  OR2_X1 U13694 ( .A1(n13509), .A2(n13506), .ZN(n13676) );
  XOR2_X1 U13695 ( .A(n13709), .B(n13710), .Z(n13506) );
  XOR2_X1 U13696 ( .A(n13711), .B(n13712), .Z(n13710) );
  OR2_X1 U13697 ( .A1(n8544), .A2(n8123), .ZN(n13509) );
  OR2_X1 U13698 ( .A1(n13513), .A2(n13510), .ZN(n13673) );
  XOR2_X1 U13699 ( .A(n13713), .B(n13714), .Z(n13510) );
  XOR2_X1 U13700 ( .A(n13715), .B(n13716), .Z(n13714) );
  OR2_X1 U13701 ( .A1(n8549), .A2(n8123), .ZN(n13513) );
  XOR2_X1 U13702 ( .A(n13717), .B(n13718), .Z(n13514) );
  XOR2_X1 U13703 ( .A(n13719), .B(n13720), .Z(n13718) );
  OR2_X1 U13704 ( .A1(n13521), .A2(n13518), .ZN(n13667) );
  XOR2_X1 U13705 ( .A(n13721), .B(n13722), .Z(n13518) );
  XOR2_X1 U13706 ( .A(n13723), .B(n13724), .Z(n13722) );
  OR2_X1 U13707 ( .A1(n8559), .A2(n8123), .ZN(n13521) );
  INV_X1 U13708 ( .A(n13271), .ZN(n8123) );
  XOR2_X1 U13709 ( .A(n13725), .B(n13726), .Z(n13271) );
  XNOR2_X1 U13710 ( .A(c_7_), .B(d_7_), .ZN(n13725) );
  XOR2_X1 U13711 ( .A(n13727), .B(n13728), .Z(n13524) );
  XOR2_X1 U13712 ( .A(n13729), .B(n13730), .Z(n13728) );
  XOR2_X1 U13713 ( .A(n13731), .B(n13732), .Z(n13528) );
  XOR2_X1 U13714 ( .A(n13733), .B(n13734), .Z(n13732) );
  XOR2_X1 U13715 ( .A(n13735), .B(n13736), .Z(n13533) );
  XOR2_X1 U13716 ( .A(n13737), .B(n13738), .Z(n13736) );
  XOR2_X1 U13717 ( .A(n13739), .B(n13740), .Z(n13536) );
  XOR2_X1 U13718 ( .A(n13741), .B(n13742), .Z(n13740) );
  XOR2_X1 U13719 ( .A(n13743), .B(n13744), .Z(n13540) );
  XOR2_X1 U13720 ( .A(n13745), .B(n13746), .Z(n13744) );
  XOR2_X1 U13721 ( .A(n13747), .B(n13748), .Z(n13544) );
  XOR2_X1 U13722 ( .A(n13749), .B(n13750), .Z(n13748) );
  XOR2_X1 U13723 ( .A(n13751), .B(n13752), .Z(n13548) );
  XOR2_X1 U13724 ( .A(n13753), .B(n13754), .Z(n13752) );
  XOR2_X1 U13725 ( .A(n13755), .B(n13756), .Z(n13552) );
  XOR2_X1 U13726 ( .A(n13757), .B(n13758), .Z(n13756) );
  XOR2_X1 U13727 ( .A(n13759), .B(n13760), .Z(n13556) );
  XOR2_X1 U13728 ( .A(n13761), .B(n13762), .Z(n13760) );
  XOR2_X1 U13729 ( .A(n13763), .B(n13764), .Z(n13560) );
  XOR2_X1 U13730 ( .A(n13765), .B(n13766), .Z(n13764) );
  XOR2_X1 U13731 ( .A(n13767), .B(n13768), .Z(n13564) );
  XOR2_X1 U13732 ( .A(n13769), .B(n13770), .Z(n13768) );
  XOR2_X1 U13733 ( .A(n13771), .B(n13772), .Z(n13568) );
  XOR2_X1 U13734 ( .A(n13773), .B(n13774), .Z(n13772) );
  XOR2_X1 U13735 ( .A(n13775), .B(n13776), .Z(n13572) );
  XOR2_X1 U13736 ( .A(n13777), .B(n13778), .Z(n13776) );
  XOR2_X1 U13737 ( .A(n13779), .B(n13780), .Z(n13576) );
  XOR2_X1 U13738 ( .A(n13781), .B(n13782), .Z(n13780) );
  XOR2_X1 U13739 ( .A(n13783), .B(n13784), .Z(n13580) );
  XOR2_X1 U13740 ( .A(n13785), .B(n13786), .Z(n13784) );
  XOR2_X1 U13741 ( .A(n13787), .B(n13788), .Z(n13584) );
  XOR2_X1 U13742 ( .A(n13789), .B(n13790), .Z(n13788) );
  XOR2_X1 U13743 ( .A(n13791), .B(n13792), .Z(n13588) );
  XOR2_X1 U13744 ( .A(n13793), .B(n13794), .Z(n13792) );
  XOR2_X1 U13745 ( .A(n13795), .B(n13796), .Z(n13592) );
  XOR2_X1 U13746 ( .A(n13797), .B(n13798), .Z(n13796) );
  XOR2_X1 U13747 ( .A(n13799), .B(n13800), .Z(n13596) );
  XOR2_X1 U13748 ( .A(n13801), .B(n13802), .Z(n13800) );
  XOR2_X1 U13749 ( .A(n13803), .B(n13804), .Z(n13600) );
  XOR2_X1 U13750 ( .A(n13805), .B(n13806), .Z(n13804) );
  XOR2_X1 U13751 ( .A(n8135), .B(n13807), .Z(n8128) );
  XOR2_X1 U13752 ( .A(n8134), .B(n8133), .Z(n13807) );
  OR2_X1 U13753 ( .A1(n8083), .A2(n7610), .ZN(n8133) );
  OR2_X1 U13754 ( .A1(n13808), .A2(n13809), .ZN(n8134) );
  AND2_X1 U13755 ( .A1(n13806), .A2(n13805), .ZN(n13809) );
  AND2_X1 U13756 ( .A1(n13803), .A2(n13810), .ZN(n13808) );
  OR2_X1 U13757 ( .A1(n13805), .A2(n13806), .ZN(n13810) );
  OR2_X1 U13758 ( .A1(n8083), .A2(n7612), .ZN(n13806) );
  OR2_X1 U13759 ( .A1(n13811), .A2(n13812), .ZN(n13805) );
  AND2_X1 U13760 ( .A1(n13802), .A2(n13801), .ZN(n13812) );
  AND2_X1 U13761 ( .A1(n13799), .A2(n13813), .ZN(n13811) );
  OR2_X1 U13762 ( .A1(n13801), .A2(n13802), .ZN(n13813) );
  OR2_X1 U13763 ( .A1(n8083), .A2(n7614), .ZN(n13802) );
  OR2_X1 U13764 ( .A1(n13814), .A2(n13815), .ZN(n13801) );
  AND2_X1 U13765 ( .A1(n13798), .A2(n13797), .ZN(n13815) );
  AND2_X1 U13766 ( .A1(n13795), .A2(n13816), .ZN(n13814) );
  OR2_X1 U13767 ( .A1(n13797), .A2(n13798), .ZN(n13816) );
  OR2_X1 U13768 ( .A1(n8083), .A2(n7616), .ZN(n13798) );
  OR2_X1 U13769 ( .A1(n13817), .A2(n13818), .ZN(n13797) );
  AND2_X1 U13770 ( .A1(n13794), .A2(n13793), .ZN(n13818) );
  AND2_X1 U13771 ( .A1(n13791), .A2(n13819), .ZN(n13817) );
  OR2_X1 U13772 ( .A1(n13793), .A2(n13794), .ZN(n13819) );
  OR2_X1 U13773 ( .A1(n8083), .A2(n7618), .ZN(n13794) );
  OR2_X1 U13774 ( .A1(n13820), .A2(n13821), .ZN(n13793) );
  AND2_X1 U13775 ( .A1(n13790), .A2(n13789), .ZN(n13821) );
  AND2_X1 U13776 ( .A1(n13787), .A2(n13822), .ZN(n13820) );
  OR2_X1 U13777 ( .A1(n13789), .A2(n13790), .ZN(n13822) );
  OR2_X1 U13778 ( .A1(n8083), .A2(n7620), .ZN(n13790) );
  OR2_X1 U13779 ( .A1(n13823), .A2(n13824), .ZN(n13789) );
  AND2_X1 U13780 ( .A1(n13786), .A2(n13785), .ZN(n13824) );
  AND2_X1 U13781 ( .A1(n13783), .A2(n13825), .ZN(n13823) );
  OR2_X1 U13782 ( .A1(n13785), .A2(n13786), .ZN(n13825) );
  OR2_X1 U13783 ( .A1(n8083), .A2(n7622), .ZN(n13786) );
  OR2_X1 U13784 ( .A1(n13826), .A2(n13827), .ZN(n13785) );
  AND2_X1 U13785 ( .A1(n13782), .A2(n13781), .ZN(n13827) );
  AND2_X1 U13786 ( .A1(n13779), .A2(n13828), .ZN(n13826) );
  OR2_X1 U13787 ( .A1(n13781), .A2(n13782), .ZN(n13828) );
  OR2_X1 U13788 ( .A1(n8624), .A2(n8083), .ZN(n13782) );
  OR2_X1 U13789 ( .A1(n13829), .A2(n13830), .ZN(n13781) );
  AND2_X1 U13790 ( .A1(n13778), .A2(n13777), .ZN(n13830) );
  AND2_X1 U13791 ( .A1(n13775), .A2(n13831), .ZN(n13829) );
  OR2_X1 U13792 ( .A1(n13777), .A2(n13778), .ZN(n13831) );
  OR2_X1 U13793 ( .A1(n8619), .A2(n8083), .ZN(n13778) );
  OR2_X1 U13794 ( .A1(n13832), .A2(n13833), .ZN(n13777) );
  AND2_X1 U13795 ( .A1(n13774), .A2(n13773), .ZN(n13833) );
  AND2_X1 U13796 ( .A1(n13771), .A2(n13834), .ZN(n13832) );
  OR2_X1 U13797 ( .A1(n13773), .A2(n13774), .ZN(n13834) );
  OR2_X1 U13798 ( .A1(n8614), .A2(n8083), .ZN(n13774) );
  OR2_X1 U13799 ( .A1(n13835), .A2(n13836), .ZN(n13773) );
  AND2_X1 U13800 ( .A1(n13770), .A2(n13769), .ZN(n13836) );
  AND2_X1 U13801 ( .A1(n13767), .A2(n13837), .ZN(n13835) );
  OR2_X1 U13802 ( .A1(n13769), .A2(n13770), .ZN(n13837) );
  OR2_X1 U13803 ( .A1(n8609), .A2(n8083), .ZN(n13770) );
  OR2_X1 U13804 ( .A1(n13838), .A2(n13839), .ZN(n13769) );
  AND2_X1 U13805 ( .A1(n13766), .A2(n13765), .ZN(n13839) );
  AND2_X1 U13806 ( .A1(n13763), .A2(n13840), .ZN(n13838) );
  OR2_X1 U13807 ( .A1(n13765), .A2(n13766), .ZN(n13840) );
  OR2_X1 U13808 ( .A1(n8604), .A2(n8083), .ZN(n13766) );
  OR2_X1 U13809 ( .A1(n13841), .A2(n13842), .ZN(n13765) );
  AND2_X1 U13810 ( .A1(n13762), .A2(n13761), .ZN(n13842) );
  AND2_X1 U13811 ( .A1(n13759), .A2(n13843), .ZN(n13841) );
  OR2_X1 U13812 ( .A1(n13761), .A2(n13762), .ZN(n13843) );
  OR2_X1 U13813 ( .A1(n8599), .A2(n8083), .ZN(n13762) );
  OR2_X1 U13814 ( .A1(n13844), .A2(n13845), .ZN(n13761) );
  AND2_X1 U13815 ( .A1(n13758), .A2(n13757), .ZN(n13845) );
  AND2_X1 U13816 ( .A1(n13755), .A2(n13846), .ZN(n13844) );
  OR2_X1 U13817 ( .A1(n13757), .A2(n13758), .ZN(n13846) );
  OR2_X1 U13818 ( .A1(n8594), .A2(n8083), .ZN(n13758) );
  OR2_X1 U13819 ( .A1(n13847), .A2(n13848), .ZN(n13757) );
  AND2_X1 U13820 ( .A1(n13754), .A2(n13753), .ZN(n13848) );
  AND2_X1 U13821 ( .A1(n13751), .A2(n13849), .ZN(n13847) );
  OR2_X1 U13822 ( .A1(n13753), .A2(n13754), .ZN(n13849) );
  OR2_X1 U13823 ( .A1(n8589), .A2(n8083), .ZN(n13754) );
  OR2_X1 U13824 ( .A1(n13850), .A2(n13851), .ZN(n13753) );
  AND2_X1 U13825 ( .A1(n13750), .A2(n13749), .ZN(n13851) );
  AND2_X1 U13826 ( .A1(n13747), .A2(n13852), .ZN(n13850) );
  OR2_X1 U13827 ( .A1(n13749), .A2(n13750), .ZN(n13852) );
  OR2_X1 U13828 ( .A1(n8584), .A2(n8083), .ZN(n13750) );
  OR2_X1 U13829 ( .A1(n13853), .A2(n13854), .ZN(n13749) );
  AND2_X1 U13830 ( .A1(n13746), .A2(n13745), .ZN(n13854) );
  AND2_X1 U13831 ( .A1(n13743), .A2(n13855), .ZN(n13853) );
  OR2_X1 U13832 ( .A1(n13745), .A2(n13746), .ZN(n13855) );
  OR2_X1 U13833 ( .A1(n8579), .A2(n8083), .ZN(n13746) );
  OR2_X1 U13834 ( .A1(n13856), .A2(n13857), .ZN(n13745) );
  AND2_X1 U13835 ( .A1(n13742), .A2(n13741), .ZN(n13857) );
  AND2_X1 U13836 ( .A1(n13739), .A2(n13858), .ZN(n13856) );
  OR2_X1 U13837 ( .A1(n13741), .A2(n13742), .ZN(n13858) );
  OR2_X1 U13838 ( .A1(n8574), .A2(n8083), .ZN(n13742) );
  OR2_X1 U13839 ( .A1(n13859), .A2(n13860), .ZN(n13741) );
  AND2_X1 U13840 ( .A1(n13738), .A2(n13737), .ZN(n13860) );
  AND2_X1 U13841 ( .A1(n13735), .A2(n13861), .ZN(n13859) );
  OR2_X1 U13842 ( .A1(n13737), .A2(n13738), .ZN(n13861) );
  OR2_X1 U13843 ( .A1(n8569), .A2(n8083), .ZN(n13738) );
  OR2_X1 U13844 ( .A1(n13862), .A2(n13863), .ZN(n13737) );
  AND2_X1 U13845 ( .A1(n13734), .A2(n13733), .ZN(n13863) );
  AND2_X1 U13846 ( .A1(n13731), .A2(n13864), .ZN(n13862) );
  OR2_X1 U13847 ( .A1(n13733), .A2(n13734), .ZN(n13864) );
  OR2_X1 U13848 ( .A1(n8564), .A2(n8083), .ZN(n13734) );
  OR2_X1 U13849 ( .A1(n13865), .A2(n13866), .ZN(n13733) );
  AND2_X1 U13850 ( .A1(n13730), .A2(n13729), .ZN(n13866) );
  AND2_X1 U13851 ( .A1(n13727), .A2(n13867), .ZN(n13865) );
  OR2_X1 U13852 ( .A1(n13729), .A2(n13730), .ZN(n13867) );
  OR2_X1 U13853 ( .A1(n8559), .A2(n8083), .ZN(n13730) );
  OR2_X1 U13854 ( .A1(n13868), .A2(n13869), .ZN(n13729) );
  AND2_X1 U13855 ( .A1(n13721), .A2(n13724), .ZN(n13869) );
  AND2_X1 U13856 ( .A1(n13870), .A2(n13723), .ZN(n13868) );
  OR2_X1 U13857 ( .A1(n13871), .A2(n13872), .ZN(n13723) );
  AND2_X1 U13858 ( .A1(n13720), .A2(n13719), .ZN(n13872) );
  AND2_X1 U13859 ( .A1(n13717), .A2(n13873), .ZN(n13871) );
  OR2_X1 U13860 ( .A1(n13719), .A2(n13720), .ZN(n13873) );
  OR2_X1 U13861 ( .A1(n8549), .A2(n8083), .ZN(n13720) );
  OR2_X1 U13862 ( .A1(n13874), .A2(n13875), .ZN(n13719) );
  AND2_X1 U13863 ( .A1(n13713), .A2(n13716), .ZN(n13875) );
  AND2_X1 U13864 ( .A1(n13876), .A2(n13715), .ZN(n13874) );
  OR2_X1 U13865 ( .A1(n13877), .A2(n13878), .ZN(n13715) );
  AND2_X1 U13866 ( .A1(n13709), .A2(n13712), .ZN(n13878) );
  AND2_X1 U13867 ( .A1(n13879), .A2(n13711), .ZN(n13877) );
  OR2_X1 U13868 ( .A1(n13880), .A2(n13881), .ZN(n13711) );
  AND2_X1 U13869 ( .A1(n13705), .A2(n13708), .ZN(n13881) );
  AND2_X1 U13870 ( .A1(n13882), .A2(n13707), .ZN(n13880) );
  OR2_X1 U13871 ( .A1(n13883), .A2(n13884), .ZN(n13707) );
  AND2_X1 U13872 ( .A1(n13701), .A2(n13704), .ZN(n13884) );
  AND2_X1 U13873 ( .A1(n13885), .A2(n13703), .ZN(n13883) );
  OR2_X1 U13874 ( .A1(n13886), .A2(n13887), .ZN(n13703) );
  AND2_X1 U13875 ( .A1(n13697), .A2(n13700), .ZN(n13887) );
  AND2_X1 U13876 ( .A1(n13699), .A2(n13888), .ZN(n13886) );
  OR2_X1 U13877 ( .A1(n13700), .A2(n13697), .ZN(n13888) );
  OR2_X1 U13878 ( .A1(n8083), .A2(n8518), .ZN(n13697) );
  OR3_X1 U13879 ( .A1(n8041), .A2(n8083), .A3(n8519), .ZN(n13700) );
  INV_X1 U13880 ( .A(n13889), .ZN(n13699) );
  OR2_X1 U13881 ( .A1(n13890), .A2(n13891), .ZN(n13889) );
  AND2_X1 U13882 ( .A1(n13892), .A2(n13893), .ZN(n13891) );
  OR2_X1 U13883 ( .A1(n13894), .A2(n7697), .ZN(n13893) );
  AND2_X1 U13884 ( .A1(n8041), .A2(n7691), .ZN(n13894) );
  AND2_X1 U13885 ( .A1(n13692), .A2(n13895), .ZN(n13890) );
  OR2_X1 U13886 ( .A1(n13896), .A2(n7701), .ZN(n13895) );
  AND2_X1 U13887 ( .A1(n8015), .A2(n7703), .ZN(n13896) );
  OR2_X1 U13888 ( .A1(n13704), .A2(n13701), .ZN(n13885) );
  XNOR2_X1 U13889 ( .A(n13897), .B(n13898), .ZN(n13701) );
  XNOR2_X1 U13890 ( .A(n13899), .B(n13900), .ZN(n13898) );
  OR2_X1 U13891 ( .A1(n8529), .A2(n8083), .ZN(n13704) );
  OR2_X1 U13892 ( .A1(n13708), .A2(n13705), .ZN(n13882) );
  XOR2_X1 U13893 ( .A(n13901), .B(n13902), .Z(n13705) );
  XOR2_X1 U13894 ( .A(n13903), .B(n13904), .Z(n13902) );
  OR2_X1 U13895 ( .A1(n8534), .A2(n8083), .ZN(n13708) );
  OR2_X1 U13896 ( .A1(n13712), .A2(n13709), .ZN(n13879) );
  XOR2_X1 U13897 ( .A(n13905), .B(n13906), .Z(n13709) );
  XOR2_X1 U13898 ( .A(n13907), .B(n13908), .Z(n13906) );
  OR2_X1 U13899 ( .A1(n8539), .A2(n8083), .ZN(n13712) );
  OR2_X1 U13900 ( .A1(n13716), .A2(n13713), .ZN(n13876) );
  XOR2_X1 U13901 ( .A(n13909), .B(n13910), .Z(n13713) );
  XOR2_X1 U13902 ( .A(n13911), .B(n13912), .Z(n13910) );
  OR2_X1 U13903 ( .A1(n8544), .A2(n8083), .ZN(n13716) );
  XOR2_X1 U13904 ( .A(n13913), .B(n13914), .Z(n13717) );
  XOR2_X1 U13905 ( .A(n13915), .B(n13916), .Z(n13914) );
  OR2_X1 U13906 ( .A1(n13724), .A2(n13721), .ZN(n13870) );
  XOR2_X1 U13907 ( .A(n13917), .B(n13918), .Z(n13721) );
  XOR2_X1 U13908 ( .A(n13919), .B(n13920), .Z(n13918) );
  OR2_X1 U13909 ( .A1(n8554), .A2(n8083), .ZN(n13724) );
  INV_X1 U13910 ( .A(n13485), .ZN(n8083) );
  XOR2_X1 U13911 ( .A(n13921), .B(n13922), .Z(n13485) );
  XNOR2_X1 U13912 ( .A(c_6_), .B(d_6_), .ZN(n13921) );
  XOR2_X1 U13913 ( .A(n13923), .B(n13924), .Z(n13727) );
  XOR2_X1 U13914 ( .A(n13925), .B(n13926), .Z(n13924) );
  XOR2_X1 U13915 ( .A(n13927), .B(n13928), .Z(n13731) );
  XOR2_X1 U13916 ( .A(n13929), .B(n13930), .Z(n13928) );
  XOR2_X1 U13917 ( .A(n13931), .B(n13932), .Z(n13735) );
  XOR2_X1 U13918 ( .A(n13933), .B(n13934), .Z(n13932) );
  XOR2_X1 U13919 ( .A(n13935), .B(n13936), .Z(n13739) );
  XOR2_X1 U13920 ( .A(n13937), .B(n13938), .Z(n13936) );
  XOR2_X1 U13921 ( .A(n13939), .B(n13940), .Z(n13743) );
  XOR2_X1 U13922 ( .A(n13941), .B(n13942), .Z(n13940) );
  XOR2_X1 U13923 ( .A(n13943), .B(n13944), .Z(n13747) );
  XOR2_X1 U13924 ( .A(n13945), .B(n13946), .Z(n13944) );
  XOR2_X1 U13925 ( .A(n13947), .B(n13948), .Z(n13751) );
  XOR2_X1 U13926 ( .A(n13949), .B(n13950), .Z(n13948) );
  XOR2_X1 U13927 ( .A(n13951), .B(n13952), .Z(n13755) );
  XOR2_X1 U13928 ( .A(n13953), .B(n13954), .Z(n13952) );
  XOR2_X1 U13929 ( .A(n13955), .B(n13956), .Z(n13759) );
  XOR2_X1 U13930 ( .A(n13957), .B(n13958), .Z(n13956) );
  XOR2_X1 U13931 ( .A(n13959), .B(n13960), .Z(n13763) );
  XOR2_X1 U13932 ( .A(n13961), .B(n13962), .Z(n13960) );
  XOR2_X1 U13933 ( .A(n13963), .B(n13964), .Z(n13767) );
  XOR2_X1 U13934 ( .A(n13965), .B(n13966), .Z(n13964) );
  XOR2_X1 U13935 ( .A(n13967), .B(n13968), .Z(n13771) );
  XOR2_X1 U13936 ( .A(n13969), .B(n13970), .Z(n13968) );
  XOR2_X1 U13937 ( .A(n13971), .B(n13972), .Z(n13775) );
  XOR2_X1 U13938 ( .A(n13973), .B(n13974), .Z(n13972) );
  XOR2_X1 U13939 ( .A(n13975), .B(n13976), .Z(n13779) );
  XOR2_X1 U13940 ( .A(n13977), .B(n13978), .Z(n13976) );
  XOR2_X1 U13941 ( .A(n13979), .B(n13980), .Z(n13783) );
  XOR2_X1 U13942 ( .A(n13981), .B(n13982), .Z(n13980) );
  XOR2_X1 U13943 ( .A(n13983), .B(n13984), .Z(n13787) );
  XOR2_X1 U13944 ( .A(n13985), .B(n13986), .Z(n13984) );
  XOR2_X1 U13945 ( .A(n13987), .B(n13988), .Z(n13791) );
  XOR2_X1 U13946 ( .A(n13989), .B(n13990), .Z(n13988) );
  XOR2_X1 U13947 ( .A(n13991), .B(n13992), .Z(n13795) );
  XOR2_X1 U13948 ( .A(n13993), .B(n13994), .Z(n13992) );
  XOR2_X1 U13949 ( .A(n13995), .B(n13996), .Z(n13799) );
  XOR2_X1 U13950 ( .A(n13997), .B(n13998), .Z(n13996) );
  XOR2_X1 U13951 ( .A(n13999), .B(n14000), .Z(n13803) );
  XOR2_X1 U13952 ( .A(n14001), .B(n14002), .Z(n14000) );
  XOR2_X1 U13953 ( .A(n8142), .B(n14003), .Z(n8135) );
  XOR2_X1 U13954 ( .A(n8141), .B(n8140), .Z(n14003) );
  OR2_X1 U13955 ( .A1(n8041), .A2(n7612), .ZN(n8140) );
  OR2_X1 U13956 ( .A1(n14004), .A2(n14005), .ZN(n8141) );
  AND2_X1 U13957 ( .A1(n14002), .A2(n14001), .ZN(n14005) );
  AND2_X1 U13958 ( .A1(n13999), .A2(n14006), .ZN(n14004) );
  OR2_X1 U13959 ( .A1(n14001), .A2(n14002), .ZN(n14006) );
  OR2_X1 U13960 ( .A1(n8041), .A2(n7614), .ZN(n14002) );
  OR2_X1 U13961 ( .A1(n14007), .A2(n14008), .ZN(n14001) );
  AND2_X1 U13962 ( .A1(n13998), .A2(n13997), .ZN(n14008) );
  AND2_X1 U13963 ( .A1(n13995), .A2(n14009), .ZN(n14007) );
  OR2_X1 U13964 ( .A1(n13997), .A2(n13998), .ZN(n14009) );
  OR2_X1 U13965 ( .A1(n8041), .A2(n7616), .ZN(n13998) );
  OR2_X1 U13966 ( .A1(n14010), .A2(n14011), .ZN(n13997) );
  AND2_X1 U13967 ( .A1(n13994), .A2(n13993), .ZN(n14011) );
  AND2_X1 U13968 ( .A1(n13991), .A2(n14012), .ZN(n14010) );
  OR2_X1 U13969 ( .A1(n13993), .A2(n13994), .ZN(n14012) );
  OR2_X1 U13970 ( .A1(n8041), .A2(n7618), .ZN(n13994) );
  OR2_X1 U13971 ( .A1(n14013), .A2(n14014), .ZN(n13993) );
  AND2_X1 U13972 ( .A1(n13990), .A2(n13989), .ZN(n14014) );
  AND2_X1 U13973 ( .A1(n13987), .A2(n14015), .ZN(n14013) );
  OR2_X1 U13974 ( .A1(n13989), .A2(n13990), .ZN(n14015) );
  OR2_X1 U13975 ( .A1(n8041), .A2(n7620), .ZN(n13990) );
  OR2_X1 U13976 ( .A1(n14016), .A2(n14017), .ZN(n13989) );
  AND2_X1 U13977 ( .A1(n13986), .A2(n13985), .ZN(n14017) );
  AND2_X1 U13978 ( .A1(n13983), .A2(n14018), .ZN(n14016) );
  OR2_X1 U13979 ( .A1(n13985), .A2(n13986), .ZN(n14018) );
  OR2_X1 U13980 ( .A1(n8041), .A2(n7622), .ZN(n13986) );
  OR2_X1 U13981 ( .A1(n14019), .A2(n14020), .ZN(n13985) );
  AND2_X1 U13982 ( .A1(n13982), .A2(n13981), .ZN(n14020) );
  AND2_X1 U13983 ( .A1(n13979), .A2(n14021), .ZN(n14019) );
  OR2_X1 U13984 ( .A1(n13981), .A2(n13982), .ZN(n14021) );
  OR2_X1 U13985 ( .A1(n8041), .A2(n7624), .ZN(n13982) );
  OR2_X1 U13986 ( .A1(n14022), .A2(n14023), .ZN(n13981) );
  AND2_X1 U13987 ( .A1(n13978), .A2(n13977), .ZN(n14023) );
  AND2_X1 U13988 ( .A1(n13975), .A2(n14024), .ZN(n14022) );
  OR2_X1 U13989 ( .A1(n13977), .A2(n13978), .ZN(n14024) );
  OR2_X1 U13990 ( .A1(n8619), .A2(n8041), .ZN(n13978) );
  OR2_X1 U13991 ( .A1(n14025), .A2(n14026), .ZN(n13977) );
  AND2_X1 U13992 ( .A1(n13974), .A2(n13973), .ZN(n14026) );
  AND2_X1 U13993 ( .A1(n13971), .A2(n14027), .ZN(n14025) );
  OR2_X1 U13994 ( .A1(n13973), .A2(n13974), .ZN(n14027) );
  OR2_X1 U13995 ( .A1(n8614), .A2(n8041), .ZN(n13974) );
  OR2_X1 U13996 ( .A1(n14028), .A2(n14029), .ZN(n13973) );
  AND2_X1 U13997 ( .A1(n13970), .A2(n13969), .ZN(n14029) );
  AND2_X1 U13998 ( .A1(n13967), .A2(n14030), .ZN(n14028) );
  OR2_X1 U13999 ( .A1(n13969), .A2(n13970), .ZN(n14030) );
  OR2_X1 U14000 ( .A1(n8609), .A2(n8041), .ZN(n13970) );
  OR2_X1 U14001 ( .A1(n14031), .A2(n14032), .ZN(n13969) );
  AND2_X1 U14002 ( .A1(n13966), .A2(n13965), .ZN(n14032) );
  AND2_X1 U14003 ( .A1(n13963), .A2(n14033), .ZN(n14031) );
  OR2_X1 U14004 ( .A1(n13965), .A2(n13966), .ZN(n14033) );
  OR2_X1 U14005 ( .A1(n8604), .A2(n8041), .ZN(n13966) );
  OR2_X1 U14006 ( .A1(n14034), .A2(n14035), .ZN(n13965) );
  AND2_X1 U14007 ( .A1(n13962), .A2(n13961), .ZN(n14035) );
  AND2_X1 U14008 ( .A1(n13959), .A2(n14036), .ZN(n14034) );
  OR2_X1 U14009 ( .A1(n13961), .A2(n13962), .ZN(n14036) );
  OR2_X1 U14010 ( .A1(n8599), .A2(n8041), .ZN(n13962) );
  OR2_X1 U14011 ( .A1(n14037), .A2(n14038), .ZN(n13961) );
  AND2_X1 U14012 ( .A1(n13958), .A2(n13957), .ZN(n14038) );
  AND2_X1 U14013 ( .A1(n13955), .A2(n14039), .ZN(n14037) );
  OR2_X1 U14014 ( .A1(n13957), .A2(n13958), .ZN(n14039) );
  OR2_X1 U14015 ( .A1(n8594), .A2(n8041), .ZN(n13958) );
  OR2_X1 U14016 ( .A1(n14040), .A2(n14041), .ZN(n13957) );
  AND2_X1 U14017 ( .A1(n13954), .A2(n13953), .ZN(n14041) );
  AND2_X1 U14018 ( .A1(n13951), .A2(n14042), .ZN(n14040) );
  OR2_X1 U14019 ( .A1(n13953), .A2(n13954), .ZN(n14042) );
  OR2_X1 U14020 ( .A1(n8589), .A2(n8041), .ZN(n13954) );
  OR2_X1 U14021 ( .A1(n14043), .A2(n14044), .ZN(n13953) );
  AND2_X1 U14022 ( .A1(n13950), .A2(n13949), .ZN(n14044) );
  AND2_X1 U14023 ( .A1(n13947), .A2(n14045), .ZN(n14043) );
  OR2_X1 U14024 ( .A1(n13949), .A2(n13950), .ZN(n14045) );
  OR2_X1 U14025 ( .A1(n8584), .A2(n8041), .ZN(n13950) );
  OR2_X1 U14026 ( .A1(n14046), .A2(n14047), .ZN(n13949) );
  AND2_X1 U14027 ( .A1(n13946), .A2(n13945), .ZN(n14047) );
  AND2_X1 U14028 ( .A1(n13943), .A2(n14048), .ZN(n14046) );
  OR2_X1 U14029 ( .A1(n13945), .A2(n13946), .ZN(n14048) );
  OR2_X1 U14030 ( .A1(n8579), .A2(n8041), .ZN(n13946) );
  OR2_X1 U14031 ( .A1(n14049), .A2(n14050), .ZN(n13945) );
  AND2_X1 U14032 ( .A1(n13942), .A2(n13941), .ZN(n14050) );
  AND2_X1 U14033 ( .A1(n13939), .A2(n14051), .ZN(n14049) );
  OR2_X1 U14034 ( .A1(n13941), .A2(n13942), .ZN(n14051) );
  OR2_X1 U14035 ( .A1(n8574), .A2(n8041), .ZN(n13942) );
  OR2_X1 U14036 ( .A1(n14052), .A2(n14053), .ZN(n13941) );
  AND2_X1 U14037 ( .A1(n13938), .A2(n13937), .ZN(n14053) );
  AND2_X1 U14038 ( .A1(n13935), .A2(n14054), .ZN(n14052) );
  OR2_X1 U14039 ( .A1(n13937), .A2(n13938), .ZN(n14054) );
  OR2_X1 U14040 ( .A1(n8569), .A2(n8041), .ZN(n13938) );
  OR2_X1 U14041 ( .A1(n14055), .A2(n14056), .ZN(n13937) );
  AND2_X1 U14042 ( .A1(n13934), .A2(n13933), .ZN(n14056) );
  AND2_X1 U14043 ( .A1(n13931), .A2(n14057), .ZN(n14055) );
  OR2_X1 U14044 ( .A1(n13933), .A2(n13934), .ZN(n14057) );
  OR2_X1 U14045 ( .A1(n8564), .A2(n8041), .ZN(n13934) );
  OR2_X1 U14046 ( .A1(n14058), .A2(n14059), .ZN(n13933) );
  AND2_X1 U14047 ( .A1(n13930), .A2(n13929), .ZN(n14059) );
  AND2_X1 U14048 ( .A1(n13927), .A2(n14060), .ZN(n14058) );
  OR2_X1 U14049 ( .A1(n13929), .A2(n13930), .ZN(n14060) );
  OR2_X1 U14050 ( .A1(n8559), .A2(n8041), .ZN(n13930) );
  OR2_X1 U14051 ( .A1(n14061), .A2(n14062), .ZN(n13929) );
  AND2_X1 U14052 ( .A1(n13926), .A2(n13925), .ZN(n14062) );
  AND2_X1 U14053 ( .A1(n13923), .A2(n14063), .ZN(n14061) );
  OR2_X1 U14054 ( .A1(n13925), .A2(n13926), .ZN(n14063) );
  OR2_X1 U14055 ( .A1(n8554), .A2(n8041), .ZN(n13926) );
  OR2_X1 U14056 ( .A1(n14064), .A2(n14065), .ZN(n13925) );
  AND2_X1 U14057 ( .A1(n13917), .A2(n13920), .ZN(n14065) );
  AND2_X1 U14058 ( .A1(n14066), .A2(n13919), .ZN(n14064) );
  OR2_X1 U14059 ( .A1(n14067), .A2(n14068), .ZN(n13919) );
  AND2_X1 U14060 ( .A1(n13916), .A2(n13915), .ZN(n14068) );
  AND2_X1 U14061 ( .A1(n13913), .A2(n14069), .ZN(n14067) );
  OR2_X1 U14062 ( .A1(n13915), .A2(n13916), .ZN(n14069) );
  OR2_X1 U14063 ( .A1(n8544), .A2(n8041), .ZN(n13916) );
  OR2_X1 U14064 ( .A1(n14070), .A2(n14071), .ZN(n13915) );
  AND2_X1 U14065 ( .A1(n13909), .A2(n13912), .ZN(n14071) );
  AND2_X1 U14066 ( .A1(n14072), .A2(n13911), .ZN(n14070) );
  OR2_X1 U14067 ( .A1(n14073), .A2(n14074), .ZN(n13911) );
  AND2_X1 U14068 ( .A1(n13905), .A2(n13908), .ZN(n14074) );
  AND2_X1 U14069 ( .A1(n14075), .A2(n13907), .ZN(n14073) );
  OR2_X1 U14070 ( .A1(n14076), .A2(n14077), .ZN(n13907) );
  AND2_X1 U14071 ( .A1(n13901), .A2(n13904), .ZN(n14077) );
  AND2_X1 U14072 ( .A1(n14078), .A2(n13903), .ZN(n14076) );
  OR2_X1 U14073 ( .A1(n14079), .A2(n14080), .ZN(n13903) );
  AND2_X1 U14074 ( .A1(n13897), .A2(n13900), .ZN(n14080) );
  AND2_X1 U14075 ( .A1(n13899), .A2(n14081), .ZN(n14079) );
  OR2_X1 U14076 ( .A1(n13900), .A2(n13897), .ZN(n14081) );
  OR2_X1 U14077 ( .A1(n8041), .A2(n8518), .ZN(n13897) );
  OR3_X1 U14078 ( .A1(n8015), .A2(n8041), .A3(n8519), .ZN(n13900) );
  INV_X1 U14079 ( .A(n14082), .ZN(n13899) );
  OR2_X1 U14080 ( .A1(n14083), .A2(n14084), .ZN(n14082) );
  AND2_X1 U14081 ( .A1(n14085), .A2(n14086), .ZN(n14084) );
  OR2_X1 U14082 ( .A1(n14087), .A2(n7697), .ZN(n14086) );
  AND2_X1 U14083 ( .A1(n8015), .A2(n7691), .ZN(n14087) );
  AND2_X1 U14084 ( .A1(n13892), .A2(n14088), .ZN(n14083) );
  OR2_X1 U14085 ( .A1(n14089), .A2(n7701), .ZN(n14088) );
  AND2_X1 U14086 ( .A1(n7988), .A2(n7703), .ZN(n14089) );
  OR2_X1 U14087 ( .A1(n13904), .A2(n13901), .ZN(n14078) );
  XNOR2_X1 U14088 ( .A(n14090), .B(n14091), .ZN(n13901) );
  XNOR2_X1 U14089 ( .A(n14092), .B(n14093), .ZN(n14091) );
  OR2_X1 U14090 ( .A1(n8529), .A2(n8041), .ZN(n13904) );
  OR2_X1 U14091 ( .A1(n13908), .A2(n13905), .ZN(n14075) );
  XOR2_X1 U14092 ( .A(n14094), .B(n14095), .Z(n13905) );
  XOR2_X1 U14093 ( .A(n14096), .B(n14097), .Z(n14095) );
  OR2_X1 U14094 ( .A1(n8534), .A2(n8041), .ZN(n13908) );
  OR2_X1 U14095 ( .A1(n13912), .A2(n13909), .ZN(n14072) );
  XOR2_X1 U14096 ( .A(n14098), .B(n14099), .Z(n13909) );
  XOR2_X1 U14097 ( .A(n14100), .B(n14101), .Z(n14099) );
  OR2_X1 U14098 ( .A1(n8539), .A2(n8041), .ZN(n13912) );
  XOR2_X1 U14099 ( .A(n14102), .B(n14103), .Z(n13913) );
  XOR2_X1 U14100 ( .A(n14104), .B(n14105), .Z(n14103) );
  OR2_X1 U14101 ( .A1(n13920), .A2(n13917), .ZN(n14066) );
  XOR2_X1 U14102 ( .A(n14106), .B(n14107), .Z(n13917) );
  XOR2_X1 U14103 ( .A(n14108), .B(n14109), .Z(n14107) );
  OR2_X1 U14104 ( .A1(n8549), .A2(n8041), .ZN(n13920) );
  INV_X1 U14105 ( .A(n13692), .ZN(n8041) );
  XOR2_X1 U14106 ( .A(n14110), .B(n14111), .Z(n13692) );
  XNOR2_X1 U14107 ( .A(c_5_), .B(d_5_), .ZN(n14110) );
  XOR2_X1 U14108 ( .A(n14112), .B(n14113), .Z(n13923) );
  XOR2_X1 U14109 ( .A(n14114), .B(n14115), .Z(n14113) );
  XOR2_X1 U14110 ( .A(n14116), .B(n14117), .Z(n13927) );
  XOR2_X1 U14111 ( .A(n14118), .B(n14119), .Z(n14117) );
  XOR2_X1 U14112 ( .A(n14120), .B(n14121), .Z(n13931) );
  XOR2_X1 U14113 ( .A(n14122), .B(n14123), .Z(n14121) );
  XOR2_X1 U14114 ( .A(n14124), .B(n14125), .Z(n13935) );
  XOR2_X1 U14115 ( .A(n14126), .B(n14127), .Z(n14125) );
  XOR2_X1 U14116 ( .A(n14128), .B(n14129), .Z(n13939) );
  XOR2_X1 U14117 ( .A(n14130), .B(n14131), .Z(n14129) );
  XOR2_X1 U14118 ( .A(n14132), .B(n14133), .Z(n13943) );
  XOR2_X1 U14119 ( .A(n14134), .B(n14135), .Z(n14133) );
  XOR2_X1 U14120 ( .A(n14136), .B(n14137), .Z(n13947) );
  XOR2_X1 U14121 ( .A(n14138), .B(n14139), .Z(n14137) );
  XOR2_X1 U14122 ( .A(n14140), .B(n14141), .Z(n13951) );
  XOR2_X1 U14123 ( .A(n14142), .B(n14143), .Z(n14141) );
  XOR2_X1 U14124 ( .A(n14144), .B(n14145), .Z(n13955) );
  XOR2_X1 U14125 ( .A(n14146), .B(n14147), .Z(n14145) );
  XOR2_X1 U14126 ( .A(n14148), .B(n14149), .Z(n13959) );
  XOR2_X1 U14127 ( .A(n14150), .B(n14151), .Z(n14149) );
  XOR2_X1 U14128 ( .A(n14152), .B(n14153), .Z(n13963) );
  XOR2_X1 U14129 ( .A(n14154), .B(n14155), .Z(n14153) );
  XOR2_X1 U14130 ( .A(n14156), .B(n14157), .Z(n13967) );
  XOR2_X1 U14131 ( .A(n14158), .B(n14159), .Z(n14157) );
  XOR2_X1 U14132 ( .A(n14160), .B(n14161), .Z(n13971) );
  XOR2_X1 U14133 ( .A(n14162), .B(n14163), .Z(n14161) );
  XOR2_X1 U14134 ( .A(n14164), .B(n14165), .Z(n13975) );
  XOR2_X1 U14135 ( .A(n14166), .B(n14167), .Z(n14165) );
  XOR2_X1 U14136 ( .A(n14168), .B(n14169), .Z(n13979) );
  XOR2_X1 U14137 ( .A(n14170), .B(n14171), .Z(n14169) );
  XOR2_X1 U14138 ( .A(n14172), .B(n14173), .Z(n13983) );
  XOR2_X1 U14139 ( .A(n14174), .B(n14175), .Z(n14173) );
  XOR2_X1 U14140 ( .A(n14176), .B(n14177), .Z(n13987) );
  XOR2_X1 U14141 ( .A(n14178), .B(n14179), .Z(n14177) );
  XOR2_X1 U14142 ( .A(n14180), .B(n14181), .Z(n13991) );
  XOR2_X1 U14143 ( .A(n14182), .B(n14183), .Z(n14181) );
  XOR2_X1 U14144 ( .A(n14184), .B(n14185), .Z(n13995) );
  XOR2_X1 U14145 ( .A(n14186), .B(n14187), .Z(n14185) );
  XOR2_X1 U14146 ( .A(n14188), .B(n14189), .Z(n13999) );
  XOR2_X1 U14147 ( .A(n14190), .B(n14191), .Z(n14189) );
  XOR2_X1 U14148 ( .A(n8149), .B(n14192), .Z(n8142) );
  XOR2_X1 U14149 ( .A(n8148), .B(n8147), .Z(n14192) );
  OR2_X1 U14150 ( .A1(n8015), .A2(n7614), .ZN(n8147) );
  OR2_X1 U14151 ( .A1(n14193), .A2(n14194), .ZN(n8148) );
  AND2_X1 U14152 ( .A1(n14191), .A2(n14190), .ZN(n14194) );
  AND2_X1 U14153 ( .A1(n14188), .A2(n14195), .ZN(n14193) );
  OR2_X1 U14154 ( .A1(n14190), .A2(n14191), .ZN(n14195) );
  OR2_X1 U14155 ( .A1(n8015), .A2(n7616), .ZN(n14191) );
  OR2_X1 U14156 ( .A1(n14196), .A2(n14197), .ZN(n14190) );
  AND2_X1 U14157 ( .A1(n14187), .A2(n14186), .ZN(n14197) );
  AND2_X1 U14158 ( .A1(n14184), .A2(n14198), .ZN(n14196) );
  OR2_X1 U14159 ( .A1(n14186), .A2(n14187), .ZN(n14198) );
  OR2_X1 U14160 ( .A1(n8015), .A2(n7618), .ZN(n14187) );
  OR2_X1 U14161 ( .A1(n14199), .A2(n14200), .ZN(n14186) );
  AND2_X1 U14162 ( .A1(n14183), .A2(n14182), .ZN(n14200) );
  AND2_X1 U14163 ( .A1(n14180), .A2(n14201), .ZN(n14199) );
  OR2_X1 U14164 ( .A1(n14182), .A2(n14183), .ZN(n14201) );
  OR2_X1 U14165 ( .A1(n8015), .A2(n7620), .ZN(n14183) );
  OR2_X1 U14166 ( .A1(n14202), .A2(n14203), .ZN(n14182) );
  AND2_X1 U14167 ( .A1(n14179), .A2(n14178), .ZN(n14203) );
  AND2_X1 U14168 ( .A1(n14176), .A2(n14204), .ZN(n14202) );
  OR2_X1 U14169 ( .A1(n14178), .A2(n14179), .ZN(n14204) );
  OR2_X1 U14170 ( .A1(n8015), .A2(n7622), .ZN(n14179) );
  OR2_X1 U14171 ( .A1(n14205), .A2(n14206), .ZN(n14178) );
  AND2_X1 U14172 ( .A1(n14175), .A2(n14174), .ZN(n14206) );
  AND2_X1 U14173 ( .A1(n14172), .A2(n14207), .ZN(n14205) );
  OR2_X1 U14174 ( .A1(n14174), .A2(n14175), .ZN(n14207) );
  OR2_X1 U14175 ( .A1(n8015), .A2(n7624), .ZN(n14175) );
  OR2_X1 U14176 ( .A1(n14208), .A2(n14209), .ZN(n14174) );
  AND2_X1 U14177 ( .A1(n14171), .A2(n14170), .ZN(n14209) );
  AND2_X1 U14178 ( .A1(n14168), .A2(n14210), .ZN(n14208) );
  OR2_X1 U14179 ( .A1(n14170), .A2(n14171), .ZN(n14210) );
  OR2_X1 U14180 ( .A1(n8015), .A2(n7626), .ZN(n14171) );
  OR2_X1 U14181 ( .A1(n14211), .A2(n14212), .ZN(n14170) );
  AND2_X1 U14182 ( .A1(n14167), .A2(n14166), .ZN(n14212) );
  AND2_X1 U14183 ( .A1(n14164), .A2(n14213), .ZN(n14211) );
  OR2_X1 U14184 ( .A1(n14166), .A2(n14167), .ZN(n14213) );
  OR2_X1 U14185 ( .A1(n8614), .A2(n8015), .ZN(n14167) );
  OR2_X1 U14186 ( .A1(n14214), .A2(n14215), .ZN(n14166) );
  AND2_X1 U14187 ( .A1(n14163), .A2(n14162), .ZN(n14215) );
  AND2_X1 U14188 ( .A1(n14160), .A2(n14216), .ZN(n14214) );
  OR2_X1 U14189 ( .A1(n14162), .A2(n14163), .ZN(n14216) );
  OR2_X1 U14190 ( .A1(n8609), .A2(n8015), .ZN(n14163) );
  OR2_X1 U14191 ( .A1(n14217), .A2(n14218), .ZN(n14162) );
  AND2_X1 U14192 ( .A1(n14159), .A2(n14158), .ZN(n14218) );
  AND2_X1 U14193 ( .A1(n14156), .A2(n14219), .ZN(n14217) );
  OR2_X1 U14194 ( .A1(n14158), .A2(n14159), .ZN(n14219) );
  OR2_X1 U14195 ( .A1(n8604), .A2(n8015), .ZN(n14159) );
  OR2_X1 U14196 ( .A1(n14220), .A2(n14221), .ZN(n14158) );
  AND2_X1 U14197 ( .A1(n14155), .A2(n14154), .ZN(n14221) );
  AND2_X1 U14198 ( .A1(n14152), .A2(n14222), .ZN(n14220) );
  OR2_X1 U14199 ( .A1(n14154), .A2(n14155), .ZN(n14222) );
  OR2_X1 U14200 ( .A1(n8599), .A2(n8015), .ZN(n14155) );
  OR2_X1 U14201 ( .A1(n14223), .A2(n14224), .ZN(n14154) );
  AND2_X1 U14202 ( .A1(n14151), .A2(n14150), .ZN(n14224) );
  AND2_X1 U14203 ( .A1(n14148), .A2(n14225), .ZN(n14223) );
  OR2_X1 U14204 ( .A1(n14150), .A2(n14151), .ZN(n14225) );
  OR2_X1 U14205 ( .A1(n8594), .A2(n8015), .ZN(n14151) );
  OR2_X1 U14206 ( .A1(n14226), .A2(n14227), .ZN(n14150) );
  AND2_X1 U14207 ( .A1(n14147), .A2(n14146), .ZN(n14227) );
  AND2_X1 U14208 ( .A1(n14144), .A2(n14228), .ZN(n14226) );
  OR2_X1 U14209 ( .A1(n14146), .A2(n14147), .ZN(n14228) );
  OR2_X1 U14210 ( .A1(n8589), .A2(n8015), .ZN(n14147) );
  OR2_X1 U14211 ( .A1(n14229), .A2(n14230), .ZN(n14146) );
  AND2_X1 U14212 ( .A1(n14143), .A2(n14142), .ZN(n14230) );
  AND2_X1 U14213 ( .A1(n14140), .A2(n14231), .ZN(n14229) );
  OR2_X1 U14214 ( .A1(n14142), .A2(n14143), .ZN(n14231) );
  OR2_X1 U14215 ( .A1(n8584), .A2(n8015), .ZN(n14143) );
  OR2_X1 U14216 ( .A1(n14232), .A2(n14233), .ZN(n14142) );
  AND2_X1 U14217 ( .A1(n14139), .A2(n14138), .ZN(n14233) );
  AND2_X1 U14218 ( .A1(n14136), .A2(n14234), .ZN(n14232) );
  OR2_X1 U14219 ( .A1(n14138), .A2(n14139), .ZN(n14234) );
  OR2_X1 U14220 ( .A1(n8579), .A2(n8015), .ZN(n14139) );
  OR2_X1 U14221 ( .A1(n14235), .A2(n14236), .ZN(n14138) );
  AND2_X1 U14222 ( .A1(n14135), .A2(n14134), .ZN(n14236) );
  AND2_X1 U14223 ( .A1(n14132), .A2(n14237), .ZN(n14235) );
  OR2_X1 U14224 ( .A1(n14134), .A2(n14135), .ZN(n14237) );
  OR2_X1 U14225 ( .A1(n8574), .A2(n8015), .ZN(n14135) );
  OR2_X1 U14226 ( .A1(n14238), .A2(n14239), .ZN(n14134) );
  AND2_X1 U14227 ( .A1(n14131), .A2(n14130), .ZN(n14239) );
  AND2_X1 U14228 ( .A1(n14128), .A2(n14240), .ZN(n14238) );
  OR2_X1 U14229 ( .A1(n14130), .A2(n14131), .ZN(n14240) );
  OR2_X1 U14230 ( .A1(n8569), .A2(n8015), .ZN(n14131) );
  OR2_X1 U14231 ( .A1(n14241), .A2(n14242), .ZN(n14130) );
  AND2_X1 U14232 ( .A1(n14127), .A2(n14126), .ZN(n14242) );
  AND2_X1 U14233 ( .A1(n14124), .A2(n14243), .ZN(n14241) );
  OR2_X1 U14234 ( .A1(n14126), .A2(n14127), .ZN(n14243) );
  OR2_X1 U14235 ( .A1(n8564), .A2(n8015), .ZN(n14127) );
  OR2_X1 U14236 ( .A1(n14244), .A2(n14245), .ZN(n14126) );
  AND2_X1 U14237 ( .A1(n14123), .A2(n14122), .ZN(n14245) );
  AND2_X1 U14238 ( .A1(n14120), .A2(n14246), .ZN(n14244) );
  OR2_X1 U14239 ( .A1(n14122), .A2(n14123), .ZN(n14246) );
  OR2_X1 U14240 ( .A1(n8559), .A2(n8015), .ZN(n14123) );
  OR2_X1 U14241 ( .A1(n14247), .A2(n14248), .ZN(n14122) );
  AND2_X1 U14242 ( .A1(n14119), .A2(n14118), .ZN(n14248) );
  AND2_X1 U14243 ( .A1(n14116), .A2(n14249), .ZN(n14247) );
  OR2_X1 U14244 ( .A1(n14118), .A2(n14119), .ZN(n14249) );
  OR2_X1 U14245 ( .A1(n8554), .A2(n8015), .ZN(n14119) );
  OR2_X1 U14246 ( .A1(n14250), .A2(n14251), .ZN(n14118) );
  AND2_X1 U14247 ( .A1(n14115), .A2(n14114), .ZN(n14251) );
  AND2_X1 U14248 ( .A1(n14112), .A2(n14252), .ZN(n14250) );
  OR2_X1 U14249 ( .A1(n14114), .A2(n14115), .ZN(n14252) );
  OR2_X1 U14250 ( .A1(n8549), .A2(n8015), .ZN(n14115) );
  OR2_X1 U14251 ( .A1(n14253), .A2(n14254), .ZN(n14114) );
  AND2_X1 U14252 ( .A1(n14106), .A2(n14109), .ZN(n14254) );
  AND2_X1 U14253 ( .A1(n14255), .A2(n14108), .ZN(n14253) );
  OR2_X1 U14254 ( .A1(n14256), .A2(n14257), .ZN(n14108) );
  AND2_X1 U14255 ( .A1(n14105), .A2(n14104), .ZN(n14257) );
  AND2_X1 U14256 ( .A1(n14102), .A2(n14258), .ZN(n14256) );
  OR2_X1 U14257 ( .A1(n14104), .A2(n14105), .ZN(n14258) );
  OR2_X1 U14258 ( .A1(n8539), .A2(n8015), .ZN(n14105) );
  OR2_X1 U14259 ( .A1(n14259), .A2(n14260), .ZN(n14104) );
  AND2_X1 U14260 ( .A1(n14098), .A2(n14101), .ZN(n14260) );
  AND2_X1 U14261 ( .A1(n14261), .A2(n14100), .ZN(n14259) );
  OR2_X1 U14262 ( .A1(n14262), .A2(n14263), .ZN(n14100) );
  AND2_X1 U14263 ( .A1(n14094), .A2(n14097), .ZN(n14263) );
  AND2_X1 U14264 ( .A1(n14264), .A2(n14096), .ZN(n14262) );
  OR2_X1 U14265 ( .A1(n14265), .A2(n14266), .ZN(n14096) );
  AND2_X1 U14266 ( .A1(n14090), .A2(n14093), .ZN(n14266) );
  AND2_X1 U14267 ( .A1(n14092), .A2(n14267), .ZN(n14265) );
  OR2_X1 U14268 ( .A1(n14093), .A2(n14090), .ZN(n14267) );
  OR2_X1 U14269 ( .A1(n8015), .A2(n8518), .ZN(n14090) );
  OR3_X1 U14270 ( .A1(n7988), .A2(n8015), .A3(n8519), .ZN(n14093) );
  INV_X1 U14271 ( .A(n14268), .ZN(n14092) );
  OR2_X1 U14272 ( .A1(n14269), .A2(n14270), .ZN(n14268) );
  AND2_X1 U14273 ( .A1(n14271), .A2(n14272), .ZN(n14270) );
  OR2_X1 U14274 ( .A1(n14273), .A2(n7697), .ZN(n14272) );
  AND2_X1 U14275 ( .A1(n7988), .A2(n7691), .ZN(n14273) );
  AND2_X1 U14276 ( .A1(n14085), .A2(n14274), .ZN(n14269) );
  OR2_X1 U14277 ( .A1(n14275), .A2(n7701), .ZN(n14274) );
  AND2_X1 U14278 ( .A1(n14276), .A2(n7703), .ZN(n14275) );
  OR2_X1 U14279 ( .A1(n14097), .A2(n14094), .ZN(n14264) );
  XNOR2_X1 U14280 ( .A(n14277), .B(n14278), .ZN(n14094) );
  XNOR2_X1 U14281 ( .A(n14279), .B(n14280), .ZN(n14278) );
  OR2_X1 U14282 ( .A1(n8529), .A2(n8015), .ZN(n14097) );
  OR2_X1 U14283 ( .A1(n14101), .A2(n14098), .ZN(n14261) );
  XOR2_X1 U14284 ( .A(n14281), .B(n14282), .Z(n14098) );
  XOR2_X1 U14285 ( .A(n14283), .B(n14284), .Z(n14282) );
  OR2_X1 U14286 ( .A1(n8534), .A2(n8015), .ZN(n14101) );
  XOR2_X1 U14287 ( .A(n14285), .B(n14286), .Z(n14102) );
  XOR2_X1 U14288 ( .A(n14287), .B(n14288), .Z(n14286) );
  OR2_X1 U14289 ( .A1(n14109), .A2(n14106), .ZN(n14255) );
  XOR2_X1 U14290 ( .A(n14289), .B(n14290), .Z(n14106) );
  XOR2_X1 U14291 ( .A(n14291), .B(n14292), .Z(n14290) );
  OR2_X1 U14292 ( .A1(n8544), .A2(n8015), .ZN(n14109) );
  INV_X1 U14293 ( .A(n13892), .ZN(n8015) );
  XOR2_X1 U14294 ( .A(n14293), .B(n14294), .Z(n13892) );
  XNOR2_X1 U14295 ( .A(c_4_), .B(d_4_), .ZN(n14293) );
  XOR2_X1 U14296 ( .A(n14295), .B(n14296), .Z(n14112) );
  XOR2_X1 U14297 ( .A(n14297), .B(n14298), .Z(n14296) );
  XOR2_X1 U14298 ( .A(n14299), .B(n14300), .Z(n14116) );
  XOR2_X1 U14299 ( .A(n14301), .B(n14302), .Z(n14300) );
  XOR2_X1 U14300 ( .A(n14303), .B(n14304), .Z(n14120) );
  XOR2_X1 U14301 ( .A(n14305), .B(n14306), .Z(n14304) );
  XOR2_X1 U14302 ( .A(n14307), .B(n14308), .Z(n14124) );
  XOR2_X1 U14303 ( .A(n14309), .B(n14310), .Z(n14308) );
  XOR2_X1 U14304 ( .A(n14311), .B(n14312), .Z(n14128) );
  XOR2_X1 U14305 ( .A(n14313), .B(n14314), .Z(n14312) );
  XOR2_X1 U14306 ( .A(n14315), .B(n14316), .Z(n14132) );
  XOR2_X1 U14307 ( .A(n14317), .B(n14318), .Z(n14316) );
  XOR2_X1 U14308 ( .A(n14319), .B(n14320), .Z(n14136) );
  XOR2_X1 U14309 ( .A(n14321), .B(n14322), .Z(n14320) );
  XOR2_X1 U14310 ( .A(n14323), .B(n14324), .Z(n14140) );
  XOR2_X1 U14311 ( .A(n14325), .B(n14326), .Z(n14324) );
  XOR2_X1 U14312 ( .A(n14327), .B(n14328), .Z(n14144) );
  XOR2_X1 U14313 ( .A(n14329), .B(n14330), .Z(n14328) );
  XOR2_X1 U14314 ( .A(n14331), .B(n14332), .Z(n14148) );
  XOR2_X1 U14315 ( .A(n14333), .B(n14334), .Z(n14332) );
  XOR2_X1 U14316 ( .A(n14335), .B(n14336), .Z(n14152) );
  XOR2_X1 U14317 ( .A(n14337), .B(n14338), .Z(n14336) );
  XOR2_X1 U14318 ( .A(n14339), .B(n14340), .Z(n14156) );
  XOR2_X1 U14319 ( .A(n14341), .B(n14342), .Z(n14340) );
  XOR2_X1 U14320 ( .A(n14343), .B(n14344), .Z(n14160) );
  XOR2_X1 U14321 ( .A(n14345), .B(n14346), .Z(n14344) );
  XOR2_X1 U14322 ( .A(n14347), .B(n14348), .Z(n14164) );
  XOR2_X1 U14323 ( .A(n14349), .B(n14350), .Z(n14348) );
  XOR2_X1 U14324 ( .A(n14351), .B(n14352), .Z(n14168) );
  XOR2_X1 U14325 ( .A(n14353), .B(n14354), .Z(n14352) );
  XOR2_X1 U14326 ( .A(n14355), .B(n14356), .Z(n14172) );
  XOR2_X1 U14327 ( .A(n14357), .B(n14358), .Z(n14356) );
  XOR2_X1 U14328 ( .A(n14359), .B(n14360), .Z(n14176) );
  XOR2_X1 U14329 ( .A(n14361), .B(n14362), .Z(n14360) );
  XOR2_X1 U14330 ( .A(n14363), .B(n14364), .Z(n14180) );
  XOR2_X1 U14331 ( .A(n14365), .B(n14366), .Z(n14364) );
  XOR2_X1 U14332 ( .A(n14367), .B(n14368), .Z(n14184) );
  XOR2_X1 U14333 ( .A(n14369), .B(n14370), .Z(n14368) );
  XOR2_X1 U14334 ( .A(n14371), .B(n14372), .Z(n14188) );
  XOR2_X1 U14335 ( .A(n14373), .B(n14374), .Z(n14372) );
  XOR2_X1 U14336 ( .A(n8157), .B(n14375), .Z(n8149) );
  XOR2_X1 U14337 ( .A(n8156), .B(n8155), .Z(n14375) );
  OR2_X1 U14338 ( .A1(n7988), .A2(n7616), .ZN(n8155) );
  OR2_X1 U14339 ( .A1(n14376), .A2(n14377), .ZN(n8156) );
  AND2_X1 U14340 ( .A1(n14374), .A2(n14373), .ZN(n14377) );
  AND2_X1 U14341 ( .A1(n14371), .A2(n14378), .ZN(n14376) );
  OR2_X1 U14342 ( .A1(n14373), .A2(n14374), .ZN(n14378) );
  OR2_X1 U14343 ( .A1(n7988), .A2(n7618), .ZN(n14374) );
  OR2_X1 U14344 ( .A1(n14379), .A2(n14380), .ZN(n14373) );
  AND2_X1 U14345 ( .A1(n14370), .A2(n14369), .ZN(n14380) );
  AND2_X1 U14346 ( .A1(n14367), .A2(n14381), .ZN(n14379) );
  OR2_X1 U14347 ( .A1(n14369), .A2(n14370), .ZN(n14381) );
  OR2_X1 U14348 ( .A1(n7988), .A2(n7620), .ZN(n14370) );
  OR2_X1 U14349 ( .A1(n14382), .A2(n14383), .ZN(n14369) );
  AND2_X1 U14350 ( .A1(n14366), .A2(n14365), .ZN(n14383) );
  AND2_X1 U14351 ( .A1(n14363), .A2(n14384), .ZN(n14382) );
  OR2_X1 U14352 ( .A1(n14365), .A2(n14366), .ZN(n14384) );
  OR2_X1 U14353 ( .A1(n7988), .A2(n7622), .ZN(n14366) );
  OR2_X1 U14354 ( .A1(n14385), .A2(n14386), .ZN(n14365) );
  AND2_X1 U14355 ( .A1(n14362), .A2(n14361), .ZN(n14386) );
  AND2_X1 U14356 ( .A1(n14359), .A2(n14387), .ZN(n14385) );
  OR2_X1 U14357 ( .A1(n14361), .A2(n14362), .ZN(n14387) );
  OR2_X1 U14358 ( .A1(n7988), .A2(n7624), .ZN(n14362) );
  OR2_X1 U14359 ( .A1(n14388), .A2(n14389), .ZN(n14361) );
  AND2_X1 U14360 ( .A1(n14358), .A2(n14357), .ZN(n14389) );
  AND2_X1 U14361 ( .A1(n14355), .A2(n14390), .ZN(n14388) );
  OR2_X1 U14362 ( .A1(n14357), .A2(n14358), .ZN(n14390) );
  OR2_X1 U14363 ( .A1(n7988), .A2(n7626), .ZN(n14358) );
  OR2_X1 U14364 ( .A1(n14391), .A2(n14392), .ZN(n14357) );
  AND2_X1 U14365 ( .A1(n14354), .A2(n14353), .ZN(n14392) );
  AND2_X1 U14366 ( .A1(n14351), .A2(n14393), .ZN(n14391) );
  OR2_X1 U14367 ( .A1(n14353), .A2(n14354), .ZN(n14393) );
  OR2_X1 U14368 ( .A1(n7988), .A2(n7628), .ZN(n14354) );
  OR2_X1 U14369 ( .A1(n14394), .A2(n14395), .ZN(n14353) );
  AND2_X1 U14370 ( .A1(n14350), .A2(n14349), .ZN(n14395) );
  AND2_X1 U14371 ( .A1(n14347), .A2(n14396), .ZN(n14394) );
  OR2_X1 U14372 ( .A1(n14349), .A2(n14350), .ZN(n14396) );
  OR2_X1 U14373 ( .A1(n8609), .A2(n7988), .ZN(n14350) );
  OR2_X1 U14374 ( .A1(n14397), .A2(n14398), .ZN(n14349) );
  AND2_X1 U14375 ( .A1(n14346), .A2(n14345), .ZN(n14398) );
  AND2_X1 U14376 ( .A1(n14343), .A2(n14399), .ZN(n14397) );
  OR2_X1 U14377 ( .A1(n14345), .A2(n14346), .ZN(n14399) );
  OR2_X1 U14378 ( .A1(n8604), .A2(n7988), .ZN(n14346) );
  OR2_X1 U14379 ( .A1(n14400), .A2(n14401), .ZN(n14345) );
  AND2_X1 U14380 ( .A1(n14342), .A2(n14341), .ZN(n14401) );
  AND2_X1 U14381 ( .A1(n14339), .A2(n14402), .ZN(n14400) );
  OR2_X1 U14382 ( .A1(n14341), .A2(n14342), .ZN(n14402) );
  OR2_X1 U14383 ( .A1(n8599), .A2(n7988), .ZN(n14342) );
  OR2_X1 U14384 ( .A1(n14403), .A2(n14404), .ZN(n14341) );
  AND2_X1 U14385 ( .A1(n14338), .A2(n14337), .ZN(n14404) );
  AND2_X1 U14386 ( .A1(n14335), .A2(n14405), .ZN(n14403) );
  OR2_X1 U14387 ( .A1(n14337), .A2(n14338), .ZN(n14405) );
  OR2_X1 U14388 ( .A1(n8594), .A2(n7988), .ZN(n14338) );
  OR2_X1 U14389 ( .A1(n14406), .A2(n14407), .ZN(n14337) );
  AND2_X1 U14390 ( .A1(n14334), .A2(n14333), .ZN(n14407) );
  AND2_X1 U14391 ( .A1(n14331), .A2(n14408), .ZN(n14406) );
  OR2_X1 U14392 ( .A1(n14333), .A2(n14334), .ZN(n14408) );
  OR2_X1 U14393 ( .A1(n8589), .A2(n7988), .ZN(n14334) );
  OR2_X1 U14394 ( .A1(n14409), .A2(n14410), .ZN(n14333) );
  AND2_X1 U14395 ( .A1(n14330), .A2(n14329), .ZN(n14410) );
  AND2_X1 U14396 ( .A1(n14327), .A2(n14411), .ZN(n14409) );
  OR2_X1 U14397 ( .A1(n14329), .A2(n14330), .ZN(n14411) );
  OR2_X1 U14398 ( .A1(n8584), .A2(n7988), .ZN(n14330) );
  OR2_X1 U14399 ( .A1(n14412), .A2(n14413), .ZN(n14329) );
  AND2_X1 U14400 ( .A1(n14326), .A2(n14325), .ZN(n14413) );
  AND2_X1 U14401 ( .A1(n14323), .A2(n14414), .ZN(n14412) );
  OR2_X1 U14402 ( .A1(n14325), .A2(n14326), .ZN(n14414) );
  OR2_X1 U14403 ( .A1(n8579), .A2(n7988), .ZN(n14326) );
  OR2_X1 U14404 ( .A1(n14415), .A2(n14416), .ZN(n14325) );
  AND2_X1 U14405 ( .A1(n14322), .A2(n14321), .ZN(n14416) );
  AND2_X1 U14406 ( .A1(n14319), .A2(n14417), .ZN(n14415) );
  OR2_X1 U14407 ( .A1(n14321), .A2(n14322), .ZN(n14417) );
  OR2_X1 U14408 ( .A1(n8574), .A2(n7988), .ZN(n14322) );
  OR2_X1 U14409 ( .A1(n14418), .A2(n14419), .ZN(n14321) );
  AND2_X1 U14410 ( .A1(n14318), .A2(n14317), .ZN(n14419) );
  AND2_X1 U14411 ( .A1(n14315), .A2(n14420), .ZN(n14418) );
  OR2_X1 U14412 ( .A1(n14317), .A2(n14318), .ZN(n14420) );
  OR2_X1 U14413 ( .A1(n8569), .A2(n7988), .ZN(n14318) );
  OR2_X1 U14414 ( .A1(n14421), .A2(n14422), .ZN(n14317) );
  AND2_X1 U14415 ( .A1(n14314), .A2(n14313), .ZN(n14422) );
  AND2_X1 U14416 ( .A1(n14311), .A2(n14423), .ZN(n14421) );
  OR2_X1 U14417 ( .A1(n14313), .A2(n14314), .ZN(n14423) );
  OR2_X1 U14418 ( .A1(n8564), .A2(n7988), .ZN(n14314) );
  OR2_X1 U14419 ( .A1(n14424), .A2(n14425), .ZN(n14313) );
  AND2_X1 U14420 ( .A1(n14310), .A2(n14309), .ZN(n14425) );
  AND2_X1 U14421 ( .A1(n14307), .A2(n14426), .ZN(n14424) );
  OR2_X1 U14422 ( .A1(n14309), .A2(n14310), .ZN(n14426) );
  OR2_X1 U14423 ( .A1(n8559), .A2(n7988), .ZN(n14310) );
  OR2_X1 U14424 ( .A1(n14427), .A2(n14428), .ZN(n14309) );
  AND2_X1 U14425 ( .A1(n14306), .A2(n14305), .ZN(n14428) );
  AND2_X1 U14426 ( .A1(n14303), .A2(n14429), .ZN(n14427) );
  OR2_X1 U14427 ( .A1(n14305), .A2(n14306), .ZN(n14429) );
  OR2_X1 U14428 ( .A1(n8554), .A2(n7988), .ZN(n14306) );
  OR2_X1 U14429 ( .A1(n14430), .A2(n14431), .ZN(n14305) );
  AND2_X1 U14430 ( .A1(n14302), .A2(n14301), .ZN(n14431) );
  AND2_X1 U14431 ( .A1(n14299), .A2(n14432), .ZN(n14430) );
  OR2_X1 U14432 ( .A1(n14301), .A2(n14302), .ZN(n14432) );
  OR2_X1 U14433 ( .A1(n8549), .A2(n7988), .ZN(n14302) );
  OR2_X1 U14434 ( .A1(n14433), .A2(n14434), .ZN(n14301) );
  AND2_X1 U14435 ( .A1(n14298), .A2(n14297), .ZN(n14434) );
  AND2_X1 U14436 ( .A1(n14295), .A2(n14435), .ZN(n14433) );
  OR2_X1 U14437 ( .A1(n14297), .A2(n14298), .ZN(n14435) );
  OR2_X1 U14438 ( .A1(n8544), .A2(n7988), .ZN(n14298) );
  OR2_X1 U14439 ( .A1(n14436), .A2(n14437), .ZN(n14297) );
  AND2_X1 U14440 ( .A1(n14289), .A2(n14292), .ZN(n14437) );
  AND2_X1 U14441 ( .A1(n14438), .A2(n14291), .ZN(n14436) );
  OR2_X1 U14442 ( .A1(n14439), .A2(n14440), .ZN(n14291) );
  AND2_X1 U14443 ( .A1(n14288), .A2(n14287), .ZN(n14440) );
  AND2_X1 U14444 ( .A1(n14285), .A2(n14441), .ZN(n14439) );
  OR2_X1 U14445 ( .A1(n14287), .A2(n14288), .ZN(n14441) );
  OR2_X1 U14446 ( .A1(n8534), .A2(n7988), .ZN(n14288) );
  OR2_X1 U14447 ( .A1(n14442), .A2(n14443), .ZN(n14287) );
  AND2_X1 U14448 ( .A1(n14281), .A2(n14284), .ZN(n14443) );
  AND2_X1 U14449 ( .A1(n14444), .A2(n14283), .ZN(n14442) );
  OR2_X1 U14450 ( .A1(n14445), .A2(n14446), .ZN(n14283) );
  AND2_X1 U14451 ( .A1(n14277), .A2(n14280), .ZN(n14446) );
  AND2_X1 U14452 ( .A1(n14279), .A2(n14447), .ZN(n14445) );
  OR2_X1 U14453 ( .A1(n14280), .A2(n14277), .ZN(n14447) );
  OR2_X1 U14454 ( .A1(n7988), .A2(n8518), .ZN(n14277) );
  OR3_X1 U14455 ( .A1(n14276), .A2(n7988), .A3(n8519), .ZN(n14280) );
  INV_X1 U14456 ( .A(n14448), .ZN(n14279) );
  OR2_X1 U14457 ( .A1(n14449), .A2(n14450), .ZN(n14448) );
  AND2_X1 U14458 ( .A1(n14451), .A2(n14452), .ZN(n14450) );
  OR2_X1 U14459 ( .A1(n14453), .A2(n7697), .ZN(n14452) );
  AND2_X1 U14460 ( .A1(n14276), .A2(n7691), .ZN(n14453) );
  AND2_X1 U14461 ( .A1(n14271), .A2(n14454), .ZN(n14449) );
  OR2_X1 U14462 ( .A1(n14455), .A2(n7701), .ZN(n14454) );
  AND2_X1 U14463 ( .A1(n14456), .A2(n7703), .ZN(n14455) );
  OR2_X1 U14464 ( .A1(n14284), .A2(n14281), .ZN(n14444) );
  XNOR2_X1 U14465 ( .A(n14457), .B(n14458), .ZN(n14281) );
  XNOR2_X1 U14466 ( .A(n14459), .B(n14460), .ZN(n14458) );
  OR2_X1 U14467 ( .A1(n8529), .A2(n7988), .ZN(n14284) );
  XNOR2_X1 U14468 ( .A(n14461), .B(n14462), .ZN(n14285) );
  XNOR2_X1 U14469 ( .A(n14463), .B(n14464), .ZN(n14461) );
  OR2_X1 U14470 ( .A1(n14292), .A2(n14289), .ZN(n14438) );
  XOR2_X1 U14471 ( .A(n14465), .B(n14466), .Z(n14289) );
  XOR2_X1 U14472 ( .A(n14467), .B(n14468), .Z(n14466) );
  OR2_X1 U14473 ( .A1(n8539), .A2(n7988), .ZN(n14292) );
  INV_X1 U14474 ( .A(n14085), .ZN(n7988) );
  XOR2_X1 U14475 ( .A(n14469), .B(n14470), .Z(n14085) );
  XNOR2_X1 U14476 ( .A(c_3_), .B(d_3_), .ZN(n14469) );
  XOR2_X1 U14477 ( .A(n14471), .B(n14472), .Z(n14295) );
  XOR2_X1 U14478 ( .A(n14473), .B(n14474), .Z(n14472) );
  XOR2_X1 U14479 ( .A(n14475), .B(n14476), .Z(n14299) );
  XOR2_X1 U14480 ( .A(n14477), .B(n14478), .Z(n14476) );
  XOR2_X1 U14481 ( .A(n14479), .B(n14480), .Z(n14303) );
  XOR2_X1 U14482 ( .A(n14481), .B(n14482), .Z(n14480) );
  XOR2_X1 U14483 ( .A(n14483), .B(n14484), .Z(n14307) );
  XOR2_X1 U14484 ( .A(n14485), .B(n14486), .Z(n14484) );
  XOR2_X1 U14485 ( .A(n14487), .B(n14488), .Z(n14311) );
  XOR2_X1 U14486 ( .A(n14489), .B(n14490), .Z(n14488) );
  XOR2_X1 U14487 ( .A(n14491), .B(n14492), .Z(n14315) );
  XOR2_X1 U14488 ( .A(n14493), .B(n14494), .Z(n14492) );
  XOR2_X1 U14489 ( .A(n14495), .B(n14496), .Z(n14319) );
  XOR2_X1 U14490 ( .A(n14497), .B(n14498), .Z(n14496) );
  XOR2_X1 U14491 ( .A(n14499), .B(n14500), .Z(n14323) );
  XOR2_X1 U14492 ( .A(n14501), .B(n14502), .Z(n14500) );
  XOR2_X1 U14493 ( .A(n14503), .B(n14504), .Z(n14327) );
  XOR2_X1 U14494 ( .A(n14505), .B(n14506), .Z(n14504) );
  XOR2_X1 U14495 ( .A(n14507), .B(n14508), .Z(n14331) );
  XOR2_X1 U14496 ( .A(n14509), .B(n14510), .Z(n14508) );
  XOR2_X1 U14497 ( .A(n14511), .B(n14512), .Z(n14335) );
  XOR2_X1 U14498 ( .A(n14513), .B(n14514), .Z(n14512) );
  XOR2_X1 U14499 ( .A(n14515), .B(n14516), .Z(n14339) );
  XOR2_X1 U14500 ( .A(n14517), .B(n14518), .Z(n14516) );
  XOR2_X1 U14501 ( .A(n14519), .B(n14520), .Z(n14343) );
  XOR2_X1 U14502 ( .A(n14521), .B(n14522), .Z(n14520) );
  XOR2_X1 U14503 ( .A(n14523), .B(n14524), .Z(n14347) );
  XOR2_X1 U14504 ( .A(n14525), .B(n14526), .Z(n14524) );
  XOR2_X1 U14505 ( .A(n14527), .B(n14528), .Z(n14351) );
  XOR2_X1 U14506 ( .A(n14529), .B(n14530), .Z(n14528) );
  XOR2_X1 U14507 ( .A(n14531), .B(n14532), .Z(n14355) );
  XOR2_X1 U14508 ( .A(n14533), .B(n14534), .Z(n14532) );
  XOR2_X1 U14509 ( .A(n14535), .B(n14536), .Z(n14359) );
  XOR2_X1 U14510 ( .A(n14537), .B(n14538), .Z(n14536) );
  XOR2_X1 U14511 ( .A(n14539), .B(n14540), .Z(n14363) );
  XOR2_X1 U14512 ( .A(n14541), .B(n14542), .Z(n14540) );
  XOR2_X1 U14513 ( .A(n14543), .B(n14544), .Z(n14367) );
  XOR2_X1 U14514 ( .A(n14545), .B(n14546), .Z(n14544) );
  XOR2_X1 U14515 ( .A(n14547), .B(n14548), .Z(n14371) );
  XOR2_X1 U14516 ( .A(n14549), .B(n14550), .Z(n14548) );
  XOR2_X1 U14517 ( .A(n14551), .B(n14552), .Z(n8157) );
  XOR2_X1 U14518 ( .A(n14553), .B(n14554), .Z(n14552) );
  AND3_X1 U14519 ( .A1(n7909), .A2(n7907), .A3(n7908), .ZN(n7910) );
  INV_X1 U14520 ( .A(n7961), .ZN(n7908) );
  OR2_X1 U14521 ( .A1(n14555), .A2(n14556), .ZN(n7961) );
  AND2_X1 U14522 ( .A1(n7980), .A2(n7979), .ZN(n14556) );
  AND2_X1 U14523 ( .A1(n7977), .A2(n14557), .ZN(n14555) );
  OR2_X1 U14524 ( .A1(n7979), .A2(n7980), .ZN(n14557) );
  OR2_X1 U14525 ( .A1(n14276), .A2(n7960), .ZN(n7980) );
  OR2_X1 U14526 ( .A1(n14558), .A2(n14559), .ZN(n7979) );
  AND2_X1 U14527 ( .A1(n7998), .A2(n7997), .ZN(n14559) );
  AND2_X1 U14528 ( .A1(n7995), .A2(n14560), .ZN(n14558) );
  OR2_X1 U14529 ( .A1(n7997), .A2(n7998), .ZN(n14560) );
  OR2_X1 U14530 ( .A1(n14276), .A2(n7608), .ZN(n7998) );
  OR2_X1 U14531 ( .A1(n14561), .A2(n14562), .ZN(n7997) );
  AND2_X1 U14532 ( .A1(n8033), .A2(n8032), .ZN(n14562) );
  AND2_X1 U14533 ( .A1(n8030), .A2(n14563), .ZN(n14561) );
  OR2_X1 U14534 ( .A1(n8032), .A2(n8033), .ZN(n14563) );
  OR2_X1 U14535 ( .A1(n14276), .A2(n7610), .ZN(n8033) );
  OR2_X1 U14536 ( .A1(n14564), .A2(n14565), .ZN(n8032) );
  AND2_X1 U14537 ( .A1(n8066), .A2(n8065), .ZN(n14565) );
  AND2_X1 U14538 ( .A1(n8063), .A2(n14566), .ZN(n14564) );
  OR2_X1 U14539 ( .A1(n8065), .A2(n8066), .ZN(n14566) );
  OR2_X1 U14540 ( .A1(n14276), .A2(n7612), .ZN(n8066) );
  OR2_X1 U14541 ( .A1(n14567), .A2(n14568), .ZN(n8065) );
  AND2_X1 U14542 ( .A1(n8115), .A2(n8114), .ZN(n14568) );
  AND2_X1 U14543 ( .A1(n8112), .A2(n14569), .ZN(n14567) );
  OR2_X1 U14544 ( .A1(n8114), .A2(n8115), .ZN(n14569) );
  OR2_X1 U14545 ( .A1(n14276), .A2(n7614), .ZN(n8115) );
  OR2_X1 U14546 ( .A1(n14570), .A2(n14571), .ZN(n8114) );
  AND2_X1 U14547 ( .A1(n8162), .A2(n8161), .ZN(n14571) );
  AND2_X1 U14548 ( .A1(n8159), .A2(n14572), .ZN(n14570) );
  OR2_X1 U14549 ( .A1(n8161), .A2(n8162), .ZN(n14572) );
  OR2_X1 U14550 ( .A1(n14276), .A2(n7616), .ZN(n8162) );
  OR2_X1 U14551 ( .A1(n14573), .A2(n14574), .ZN(n8161) );
  AND2_X1 U14552 ( .A1(n14554), .A2(n14553), .ZN(n14574) );
  AND2_X1 U14553 ( .A1(n14551), .A2(n14575), .ZN(n14573) );
  OR2_X1 U14554 ( .A1(n14553), .A2(n14554), .ZN(n14575) );
  OR2_X1 U14555 ( .A1(n14276), .A2(n7618), .ZN(n14554) );
  OR2_X1 U14556 ( .A1(n14576), .A2(n14577), .ZN(n14553) );
  AND2_X1 U14557 ( .A1(n14550), .A2(n14549), .ZN(n14577) );
  AND2_X1 U14558 ( .A1(n14547), .A2(n14578), .ZN(n14576) );
  OR2_X1 U14559 ( .A1(n14549), .A2(n14550), .ZN(n14578) );
  OR2_X1 U14560 ( .A1(n14276), .A2(n7620), .ZN(n14550) );
  OR2_X1 U14561 ( .A1(n14579), .A2(n14580), .ZN(n14549) );
  AND2_X1 U14562 ( .A1(n14546), .A2(n14545), .ZN(n14580) );
  AND2_X1 U14563 ( .A1(n14543), .A2(n14581), .ZN(n14579) );
  OR2_X1 U14564 ( .A1(n14545), .A2(n14546), .ZN(n14581) );
  OR2_X1 U14565 ( .A1(n14276), .A2(n7622), .ZN(n14546) );
  OR2_X1 U14566 ( .A1(n14582), .A2(n14583), .ZN(n14545) );
  AND2_X1 U14567 ( .A1(n14542), .A2(n14541), .ZN(n14583) );
  AND2_X1 U14568 ( .A1(n14539), .A2(n14584), .ZN(n14582) );
  OR2_X1 U14569 ( .A1(n14541), .A2(n14542), .ZN(n14584) );
  OR2_X1 U14570 ( .A1(n14276), .A2(n7624), .ZN(n14542) );
  OR2_X1 U14571 ( .A1(n14585), .A2(n14586), .ZN(n14541) );
  AND2_X1 U14572 ( .A1(n14538), .A2(n14537), .ZN(n14586) );
  AND2_X1 U14573 ( .A1(n14535), .A2(n14587), .ZN(n14585) );
  OR2_X1 U14574 ( .A1(n14537), .A2(n14538), .ZN(n14587) );
  OR2_X1 U14575 ( .A1(n14276), .A2(n7626), .ZN(n14538) );
  OR2_X1 U14576 ( .A1(n14588), .A2(n14589), .ZN(n14537) );
  AND2_X1 U14577 ( .A1(n14534), .A2(n14533), .ZN(n14589) );
  AND2_X1 U14578 ( .A1(n14531), .A2(n14590), .ZN(n14588) );
  OR2_X1 U14579 ( .A1(n14533), .A2(n14534), .ZN(n14590) );
  OR2_X1 U14580 ( .A1(n14276), .A2(n7628), .ZN(n14534) );
  OR2_X1 U14581 ( .A1(n14591), .A2(n14592), .ZN(n14533) );
  AND2_X1 U14582 ( .A1(n14530), .A2(n14529), .ZN(n14592) );
  AND2_X1 U14583 ( .A1(n14527), .A2(n14593), .ZN(n14591) );
  OR2_X1 U14584 ( .A1(n14529), .A2(n14530), .ZN(n14593) );
  OR2_X1 U14585 ( .A1(n14276), .A2(n7630), .ZN(n14530) );
  OR2_X1 U14586 ( .A1(n14594), .A2(n14595), .ZN(n14529) );
  AND2_X1 U14587 ( .A1(n14526), .A2(n14525), .ZN(n14595) );
  AND2_X1 U14588 ( .A1(n14523), .A2(n14596), .ZN(n14594) );
  OR2_X1 U14589 ( .A1(n14525), .A2(n14526), .ZN(n14596) );
  OR2_X1 U14590 ( .A1(n8604), .A2(n14276), .ZN(n14526) );
  OR2_X1 U14591 ( .A1(n14597), .A2(n14598), .ZN(n14525) );
  AND2_X1 U14592 ( .A1(n14522), .A2(n14521), .ZN(n14598) );
  AND2_X1 U14593 ( .A1(n14519), .A2(n14599), .ZN(n14597) );
  OR2_X1 U14594 ( .A1(n14521), .A2(n14522), .ZN(n14599) );
  OR2_X1 U14595 ( .A1(n8599), .A2(n14276), .ZN(n14522) );
  OR2_X1 U14596 ( .A1(n14600), .A2(n14601), .ZN(n14521) );
  AND2_X1 U14597 ( .A1(n14518), .A2(n14517), .ZN(n14601) );
  AND2_X1 U14598 ( .A1(n14515), .A2(n14602), .ZN(n14600) );
  OR2_X1 U14599 ( .A1(n14517), .A2(n14518), .ZN(n14602) );
  OR2_X1 U14600 ( .A1(n8594), .A2(n14276), .ZN(n14518) );
  OR2_X1 U14601 ( .A1(n14603), .A2(n14604), .ZN(n14517) );
  AND2_X1 U14602 ( .A1(n14514), .A2(n14513), .ZN(n14604) );
  AND2_X1 U14603 ( .A1(n14511), .A2(n14605), .ZN(n14603) );
  OR2_X1 U14604 ( .A1(n14513), .A2(n14514), .ZN(n14605) );
  OR2_X1 U14605 ( .A1(n8589), .A2(n14276), .ZN(n14514) );
  OR2_X1 U14606 ( .A1(n14606), .A2(n14607), .ZN(n14513) );
  AND2_X1 U14607 ( .A1(n14510), .A2(n14509), .ZN(n14607) );
  AND2_X1 U14608 ( .A1(n14507), .A2(n14608), .ZN(n14606) );
  OR2_X1 U14609 ( .A1(n14509), .A2(n14510), .ZN(n14608) );
  OR2_X1 U14610 ( .A1(n8584), .A2(n14276), .ZN(n14510) );
  OR2_X1 U14611 ( .A1(n14609), .A2(n14610), .ZN(n14509) );
  AND2_X1 U14612 ( .A1(n14506), .A2(n14505), .ZN(n14610) );
  AND2_X1 U14613 ( .A1(n14503), .A2(n14611), .ZN(n14609) );
  OR2_X1 U14614 ( .A1(n14505), .A2(n14506), .ZN(n14611) );
  OR2_X1 U14615 ( .A1(n8579), .A2(n14276), .ZN(n14506) );
  OR2_X1 U14616 ( .A1(n14612), .A2(n14613), .ZN(n14505) );
  AND2_X1 U14617 ( .A1(n14502), .A2(n14501), .ZN(n14613) );
  AND2_X1 U14618 ( .A1(n14499), .A2(n14614), .ZN(n14612) );
  OR2_X1 U14619 ( .A1(n14501), .A2(n14502), .ZN(n14614) );
  OR2_X1 U14620 ( .A1(n8574), .A2(n14276), .ZN(n14502) );
  OR2_X1 U14621 ( .A1(n14615), .A2(n14616), .ZN(n14501) );
  AND2_X1 U14622 ( .A1(n14498), .A2(n14497), .ZN(n14616) );
  AND2_X1 U14623 ( .A1(n14495), .A2(n14617), .ZN(n14615) );
  OR2_X1 U14624 ( .A1(n14497), .A2(n14498), .ZN(n14617) );
  OR2_X1 U14625 ( .A1(n8569), .A2(n14276), .ZN(n14498) );
  OR2_X1 U14626 ( .A1(n14618), .A2(n14619), .ZN(n14497) );
  AND2_X1 U14627 ( .A1(n14494), .A2(n14493), .ZN(n14619) );
  AND2_X1 U14628 ( .A1(n14491), .A2(n14620), .ZN(n14618) );
  OR2_X1 U14629 ( .A1(n14493), .A2(n14494), .ZN(n14620) );
  OR2_X1 U14630 ( .A1(n8564), .A2(n14276), .ZN(n14494) );
  OR2_X1 U14631 ( .A1(n14621), .A2(n14622), .ZN(n14493) );
  AND2_X1 U14632 ( .A1(n14490), .A2(n14489), .ZN(n14622) );
  AND2_X1 U14633 ( .A1(n14487), .A2(n14623), .ZN(n14621) );
  OR2_X1 U14634 ( .A1(n14489), .A2(n14490), .ZN(n14623) );
  OR2_X1 U14635 ( .A1(n8559), .A2(n14276), .ZN(n14490) );
  OR2_X1 U14636 ( .A1(n14624), .A2(n14625), .ZN(n14489) );
  AND2_X1 U14637 ( .A1(n14486), .A2(n14485), .ZN(n14625) );
  AND2_X1 U14638 ( .A1(n14483), .A2(n14626), .ZN(n14624) );
  OR2_X1 U14639 ( .A1(n14485), .A2(n14486), .ZN(n14626) );
  OR2_X1 U14640 ( .A1(n8554), .A2(n14276), .ZN(n14486) );
  OR2_X1 U14641 ( .A1(n14627), .A2(n14628), .ZN(n14485) );
  AND2_X1 U14642 ( .A1(n14482), .A2(n14481), .ZN(n14628) );
  AND2_X1 U14643 ( .A1(n14479), .A2(n14629), .ZN(n14627) );
  OR2_X1 U14644 ( .A1(n14481), .A2(n14482), .ZN(n14629) );
  OR2_X1 U14645 ( .A1(n8549), .A2(n14276), .ZN(n14482) );
  OR2_X1 U14646 ( .A1(n14630), .A2(n14631), .ZN(n14481) );
  AND2_X1 U14647 ( .A1(n14478), .A2(n14477), .ZN(n14631) );
  AND2_X1 U14648 ( .A1(n14475), .A2(n14632), .ZN(n14630) );
  OR2_X1 U14649 ( .A1(n14477), .A2(n14478), .ZN(n14632) );
  OR2_X1 U14650 ( .A1(n8544), .A2(n14276), .ZN(n14478) );
  OR2_X1 U14651 ( .A1(n14633), .A2(n14634), .ZN(n14477) );
  AND2_X1 U14652 ( .A1(n14474), .A2(n14473), .ZN(n14634) );
  AND2_X1 U14653 ( .A1(n14471), .A2(n14635), .ZN(n14633) );
  OR2_X1 U14654 ( .A1(n14473), .A2(n14474), .ZN(n14635) );
  OR2_X1 U14655 ( .A1(n8539), .A2(n14276), .ZN(n14474) );
  OR2_X1 U14656 ( .A1(n14636), .A2(n14637), .ZN(n14473) );
  AND2_X1 U14657 ( .A1(n14465), .A2(n14468), .ZN(n14637) );
  AND2_X1 U14658 ( .A1(n14638), .A2(n14467), .ZN(n14636) );
  OR2_X1 U14659 ( .A1(n14639), .A2(n14640), .ZN(n14467) );
  AND2_X1 U14660 ( .A1(n14464), .A2(n14463), .ZN(n14640) );
  AND2_X1 U14661 ( .A1(n14462), .A2(n14641), .ZN(n14639) );
  OR2_X1 U14662 ( .A1(n14463), .A2(n14464), .ZN(n14641) );
  OR2_X1 U14663 ( .A1(n8529), .A2(n14276), .ZN(n14464) );
  OR2_X1 U14664 ( .A1(n14642), .A2(n14643), .ZN(n14463) );
  AND2_X1 U14665 ( .A1(n14457), .A2(n14460), .ZN(n14643) );
  AND2_X1 U14666 ( .A1(n14459), .A2(n14644), .ZN(n14642) );
  OR2_X1 U14667 ( .A1(n14460), .A2(n14457), .ZN(n14644) );
  OR2_X1 U14668 ( .A1(n14276), .A2(n8518), .ZN(n14457) );
  OR3_X1 U14669 ( .A1(n14456), .A2(n14276), .A3(n8519), .ZN(n14460) );
  INV_X1 U14670 ( .A(n14645), .ZN(n14459) );
  OR2_X1 U14671 ( .A1(n14646), .A2(n14647), .ZN(n14645) );
  AND2_X1 U14672 ( .A1(n14451), .A2(n14648), .ZN(n14647) );
  OR2_X1 U14673 ( .A1(n14649), .A2(n7701), .ZN(n14648) );
  AND2_X1 U14674 ( .A1(n14650), .A2(n7703), .ZN(n7701) );
  AND2_X1 U14675 ( .A1(n7703), .A2(n14651), .ZN(n14649) );
  INV_X1 U14676 ( .A(n14652), .ZN(n7703) );
  AND2_X1 U14677 ( .A1(n14653), .A2(n14654), .ZN(n14646) );
  OR2_X1 U14678 ( .A1(n14655), .A2(n7697), .ZN(n14654) );
  AND2_X1 U14679 ( .A1(n7691), .A2(n14652), .ZN(n7697) );
  AND2_X1 U14680 ( .A1(n14456), .A2(n7691), .ZN(n14655) );
  INV_X1 U14681 ( .A(n14651), .ZN(n14653) );
  XNOR2_X1 U14682 ( .A(n14656), .B(n14657), .ZN(n14462) );
  OR2_X1 U14683 ( .A1(n14658), .A2(n14659), .ZN(n14656) );
  INV_X1 U14684 ( .A(n14660), .ZN(n14659) );
  AND2_X1 U14685 ( .A1(n14661), .A2(n14662), .ZN(n14658) );
  OR2_X1 U14686 ( .A1(n14652), .A2(n7666), .ZN(n14661) );
  OR2_X1 U14687 ( .A1(n14468), .A2(n14465), .ZN(n14638) );
  XNOR2_X1 U14688 ( .A(n14663), .B(n14664), .ZN(n14465) );
  XNOR2_X1 U14689 ( .A(n14665), .B(n14666), .ZN(n14664) );
  OR2_X1 U14690 ( .A1(n8534), .A2(n14276), .ZN(n14468) );
  INV_X1 U14691 ( .A(n14271), .ZN(n14276) );
  XOR2_X1 U14692 ( .A(n14667), .B(n14668), .Z(n14271) );
  XNOR2_X1 U14693 ( .A(c_2_), .B(d_2_), .ZN(n14667) );
  XOR2_X1 U14694 ( .A(n14669), .B(n14670), .Z(n14471) );
  XOR2_X1 U14695 ( .A(n14671), .B(n14672), .Z(n14670) );
  XNOR2_X1 U14696 ( .A(n14673), .B(n14674), .ZN(n14475) );
  XNOR2_X1 U14697 ( .A(n14675), .B(n14676), .ZN(n14673) );
  XNOR2_X1 U14698 ( .A(n14677), .B(n14678), .ZN(n14479) );
  XNOR2_X1 U14699 ( .A(n14679), .B(n14680), .ZN(n14677) );
  XNOR2_X1 U14700 ( .A(n14681), .B(n14682), .ZN(n14483) );
  XNOR2_X1 U14701 ( .A(n14683), .B(n14684), .ZN(n14681) );
  XNOR2_X1 U14702 ( .A(n14685), .B(n14686), .ZN(n14487) );
  XNOR2_X1 U14703 ( .A(n14687), .B(n14688), .ZN(n14685) );
  XNOR2_X1 U14704 ( .A(n14689), .B(n14690), .ZN(n14491) );
  XNOR2_X1 U14705 ( .A(n14691), .B(n14692), .ZN(n14689) );
  XNOR2_X1 U14706 ( .A(n14693), .B(n14694), .ZN(n14495) );
  XNOR2_X1 U14707 ( .A(n14695), .B(n14696), .ZN(n14693) );
  XNOR2_X1 U14708 ( .A(n14697), .B(n14698), .ZN(n14499) );
  XNOR2_X1 U14709 ( .A(n14699), .B(n14700), .ZN(n14697) );
  XNOR2_X1 U14710 ( .A(n14701), .B(n14702), .ZN(n14503) );
  XNOR2_X1 U14711 ( .A(n14703), .B(n14704), .ZN(n14701) );
  XNOR2_X1 U14712 ( .A(n14705), .B(n14706), .ZN(n14507) );
  XNOR2_X1 U14713 ( .A(n14707), .B(n14708), .ZN(n14705) );
  XNOR2_X1 U14714 ( .A(n14709), .B(n14710), .ZN(n14511) );
  XNOR2_X1 U14715 ( .A(n14711), .B(n14712), .ZN(n14709) );
  XNOR2_X1 U14716 ( .A(n14713), .B(n14714), .ZN(n14515) );
  XNOR2_X1 U14717 ( .A(n14715), .B(n14716), .ZN(n14713) );
  XNOR2_X1 U14718 ( .A(n14717), .B(n14718), .ZN(n14519) );
  XNOR2_X1 U14719 ( .A(n14719), .B(n14720), .ZN(n14717) );
  XNOR2_X1 U14720 ( .A(n14721), .B(n14722), .ZN(n14523) );
  XNOR2_X1 U14721 ( .A(n14723), .B(n14724), .ZN(n14721) );
  XNOR2_X1 U14722 ( .A(n14725), .B(n14726), .ZN(n14527) );
  XNOR2_X1 U14723 ( .A(n14727), .B(n14728), .ZN(n14725) );
  XNOR2_X1 U14724 ( .A(n14729), .B(n14730), .ZN(n14531) );
  XNOR2_X1 U14725 ( .A(n14731), .B(n14732), .ZN(n14729) );
  XNOR2_X1 U14726 ( .A(n14733), .B(n14734), .ZN(n14535) );
  XNOR2_X1 U14727 ( .A(n14735), .B(n14736), .ZN(n14733) );
  XNOR2_X1 U14728 ( .A(n14737), .B(n14738), .ZN(n14539) );
  XNOR2_X1 U14729 ( .A(n14739), .B(n14740), .ZN(n14737) );
  XNOR2_X1 U14730 ( .A(n14741), .B(n14742), .ZN(n14543) );
  XNOR2_X1 U14731 ( .A(n14743), .B(n14744), .ZN(n14741) );
  XOR2_X1 U14732 ( .A(n14745), .B(n14746), .Z(n14547) );
  XOR2_X1 U14733 ( .A(n14747), .B(n14748), .Z(n14746) );
  XOR2_X1 U14734 ( .A(n14749), .B(n14750), .Z(n14551) );
  XOR2_X1 U14735 ( .A(n14751), .B(n14752), .Z(n14750) );
  XOR2_X1 U14736 ( .A(n14753), .B(n14754), .Z(n8159) );
  XOR2_X1 U14737 ( .A(n14755), .B(n14756), .Z(n14754) );
  XOR2_X1 U14738 ( .A(n14757), .B(n14758), .Z(n8112) );
  XOR2_X1 U14739 ( .A(n14759), .B(n14760), .Z(n14758) );
  XOR2_X1 U14740 ( .A(n14761), .B(n14762), .Z(n8063) );
  XOR2_X1 U14741 ( .A(n14763), .B(n14764), .Z(n14762) );
  XOR2_X1 U14742 ( .A(n14765), .B(n14766), .Z(n8030) );
  XOR2_X1 U14743 ( .A(n14767), .B(n14768), .Z(n14766) );
  XOR2_X1 U14744 ( .A(n14769), .B(n14770), .Z(n7995) );
  XOR2_X1 U14745 ( .A(n14771), .B(n14772), .Z(n14770) );
  XOR2_X1 U14746 ( .A(n14773), .B(n14774), .Z(n7977) );
  XOR2_X1 U14747 ( .A(n14775), .B(n14776), .Z(n14774) );
  XOR2_X1 U14748 ( .A(n14777), .B(n7959), .Z(n7907) );
  OR2_X1 U14749 ( .A1(n14778), .A2(n14779), .ZN(n7959) );
  AND2_X1 U14750 ( .A1(n14780), .A2(n14781), .ZN(n14779) );
  AND2_X1 U14751 ( .A1(n14782), .A2(n14783), .ZN(n14778) );
  OR2_X1 U14752 ( .A1(n14781), .A2(n14780), .ZN(n14782) );
  OR2_X1 U14753 ( .A1(n14651), .A2(n7960), .ZN(n14777) );
  XOR2_X1 U14754 ( .A(n14784), .B(n14780), .Z(n7909) );
  OR2_X1 U14755 ( .A1(n14785), .A2(n14786), .ZN(n14780) );
  AND2_X1 U14756 ( .A1(n14773), .A2(n14775), .ZN(n14786) );
  AND2_X1 U14757 ( .A1(n14787), .A2(n14776), .ZN(n14785) );
  OR2_X1 U14758 ( .A1(n14456), .A2(n7608), .ZN(n14776) );
  OR2_X1 U14759 ( .A1(n14775), .A2(n14773), .ZN(n14787) );
  OR2_X1 U14760 ( .A1(n8056), .A2(n7666), .ZN(n14773) );
  OR2_X1 U14761 ( .A1(n14788), .A2(n14789), .ZN(n14775) );
  AND2_X1 U14762 ( .A1(n14769), .A2(n14771), .ZN(n14789) );
  AND2_X1 U14763 ( .A1(n14790), .A2(n14772), .ZN(n14788) );
  OR2_X1 U14764 ( .A1(n8105), .A2(n7666), .ZN(n14772) );
  OR2_X1 U14765 ( .A1(n14771), .A2(n14769), .ZN(n14790) );
  OR2_X1 U14766 ( .A1(n14456), .A2(n7610), .ZN(n14769) );
  XNOR2_X1 U14767 ( .A(n14791), .B(n14792), .ZN(n8056) );
  XNOR2_X1 U14768 ( .A(a_2_), .B(b_2_), .ZN(n14791) );
  OR2_X1 U14769 ( .A1(n14793), .A2(n14794), .ZN(n14771) );
  AND2_X1 U14770 ( .A1(n14765), .A2(n14767), .ZN(n14794) );
  AND2_X1 U14771 ( .A1(n14795), .A2(n14768), .ZN(n14793) );
  OR2_X1 U14772 ( .A1(n8152), .A2(n7666), .ZN(n14768) );
  OR2_X1 U14773 ( .A1(n14767), .A2(n14765), .ZN(n14795) );
  OR2_X1 U14774 ( .A1(n14456), .A2(n7612), .ZN(n14765) );
  XNOR2_X1 U14775 ( .A(n14796), .B(n14797), .ZN(n8105) );
  XNOR2_X1 U14776 ( .A(a_3_), .B(b_3_), .ZN(n14796) );
  OR2_X1 U14777 ( .A1(n14798), .A2(n14799), .ZN(n14767) );
  AND2_X1 U14778 ( .A1(n14761), .A2(n14763), .ZN(n14799) );
  AND2_X1 U14779 ( .A1(n14800), .A2(n14764), .ZN(n14798) );
  OR2_X1 U14780 ( .A1(n8644), .A2(n7666), .ZN(n14764) );
  OR2_X1 U14781 ( .A1(n14763), .A2(n14761), .ZN(n14800) );
  OR2_X1 U14782 ( .A1(n14456), .A2(n7614), .ZN(n14761) );
  XNOR2_X1 U14783 ( .A(n14801), .B(n14802), .ZN(n8152) );
  XNOR2_X1 U14784 ( .A(a_4_), .B(b_4_), .ZN(n14801) );
  OR2_X1 U14785 ( .A1(n14803), .A2(n14804), .ZN(n14763) );
  AND2_X1 U14786 ( .A1(n14757), .A2(n14759), .ZN(n14804) );
  AND2_X1 U14787 ( .A1(n14805), .A2(n14760), .ZN(n14803) );
  OR2_X1 U14788 ( .A1(n8639), .A2(n7666), .ZN(n14760) );
  OR2_X1 U14789 ( .A1(n14759), .A2(n14757), .ZN(n14805) );
  OR2_X1 U14790 ( .A1(n14456), .A2(n7616), .ZN(n14757) );
  XNOR2_X1 U14791 ( .A(n14806), .B(n14807), .ZN(n8644) );
  XNOR2_X1 U14792 ( .A(a_5_), .B(b_5_), .ZN(n14806) );
  OR2_X1 U14793 ( .A1(n14808), .A2(n14809), .ZN(n14759) );
  AND2_X1 U14794 ( .A1(n14753), .A2(n14755), .ZN(n14809) );
  AND2_X1 U14795 ( .A1(n14810), .A2(n14756), .ZN(n14808) );
  OR2_X1 U14796 ( .A1(n8634), .A2(n7666), .ZN(n14756) );
  OR2_X1 U14797 ( .A1(n14755), .A2(n14753), .ZN(n14810) );
  OR2_X1 U14798 ( .A1(n14456), .A2(n7618), .ZN(n14753) );
  XNOR2_X1 U14799 ( .A(n14811), .B(n14812), .ZN(n8639) );
  XNOR2_X1 U14800 ( .A(a_6_), .B(b_6_), .ZN(n14811) );
  OR2_X1 U14801 ( .A1(n14813), .A2(n14814), .ZN(n14755) );
  AND2_X1 U14802 ( .A1(n14749), .A2(n14751), .ZN(n14814) );
  AND2_X1 U14803 ( .A1(n14815), .A2(n14752), .ZN(n14813) );
  OR2_X1 U14804 ( .A1(n8629), .A2(n7666), .ZN(n14752) );
  OR2_X1 U14805 ( .A1(n14751), .A2(n14749), .ZN(n14815) );
  OR2_X1 U14806 ( .A1(n14456), .A2(n7620), .ZN(n14749) );
  XNOR2_X1 U14807 ( .A(n14816), .B(n14817), .ZN(n8634) );
  XNOR2_X1 U14808 ( .A(a_7_), .B(b_7_), .ZN(n14816) );
  OR2_X1 U14809 ( .A1(n14818), .A2(n14819), .ZN(n14751) );
  AND2_X1 U14810 ( .A1(n14745), .A2(n14747), .ZN(n14819) );
  AND2_X1 U14811 ( .A1(n14820), .A2(n14748), .ZN(n14818) );
  OR2_X1 U14812 ( .A1(n8624), .A2(n7666), .ZN(n14748) );
  OR2_X1 U14813 ( .A1(n14747), .A2(n14745), .ZN(n14820) );
  OR2_X1 U14814 ( .A1(n14456), .A2(n7622), .ZN(n14745) );
  XNOR2_X1 U14815 ( .A(n14821), .B(n14822), .ZN(n8629) );
  XNOR2_X1 U14816 ( .A(a_8_), .B(b_8_), .ZN(n14821) );
  OR2_X1 U14817 ( .A1(n14823), .A2(n14824), .ZN(n14747) );
  AND2_X1 U14818 ( .A1(n14742), .A2(n14744), .ZN(n14824) );
  AND2_X1 U14819 ( .A1(n14825), .A2(n14743), .ZN(n14823) );
  OR2_X1 U14820 ( .A1(n8619), .A2(n7666), .ZN(n14743) );
  OR2_X1 U14821 ( .A1(n14744), .A2(n14742), .ZN(n14825) );
  OR2_X1 U14822 ( .A1(n14456), .A2(n7624), .ZN(n14742) );
  XNOR2_X1 U14823 ( .A(n14826), .B(n14827), .ZN(n8624) );
  XNOR2_X1 U14824 ( .A(a_9_), .B(b_9_), .ZN(n14826) );
  OR2_X1 U14825 ( .A1(n14828), .A2(n14829), .ZN(n14744) );
  AND2_X1 U14826 ( .A1(n14738), .A2(n14740), .ZN(n14829) );
  AND2_X1 U14827 ( .A1(n14830), .A2(n14739), .ZN(n14828) );
  OR2_X1 U14828 ( .A1(n8614), .A2(n7666), .ZN(n14739) );
  OR2_X1 U14829 ( .A1(n14740), .A2(n14738), .ZN(n14830) );
  OR2_X1 U14830 ( .A1(n14456), .A2(n7626), .ZN(n14738) );
  XNOR2_X1 U14831 ( .A(n14831), .B(n14832), .ZN(n8619) );
  XNOR2_X1 U14832 ( .A(a_10_), .B(b_10_), .ZN(n14831) );
  OR2_X1 U14833 ( .A1(n14833), .A2(n14834), .ZN(n14740) );
  AND2_X1 U14834 ( .A1(n14734), .A2(n14736), .ZN(n14834) );
  AND2_X1 U14835 ( .A1(n14835), .A2(n14735), .ZN(n14833) );
  OR2_X1 U14836 ( .A1(n8609), .A2(n7666), .ZN(n14735) );
  OR2_X1 U14837 ( .A1(n14736), .A2(n14734), .ZN(n14835) );
  OR2_X1 U14838 ( .A1(n14456), .A2(n7628), .ZN(n14734) );
  XNOR2_X1 U14839 ( .A(n14836), .B(n14837), .ZN(n8614) );
  XNOR2_X1 U14840 ( .A(a_11_), .B(b_11_), .ZN(n14836) );
  OR2_X1 U14841 ( .A1(n14838), .A2(n14839), .ZN(n14736) );
  AND2_X1 U14842 ( .A1(n14730), .A2(n14732), .ZN(n14839) );
  AND2_X1 U14843 ( .A1(n14840), .A2(n14731), .ZN(n14838) );
  OR2_X1 U14844 ( .A1(n8604), .A2(n7666), .ZN(n14731) );
  OR2_X1 U14845 ( .A1(n14732), .A2(n14730), .ZN(n14840) );
  OR2_X1 U14846 ( .A1(n14456), .A2(n7630), .ZN(n14730) );
  XNOR2_X1 U14847 ( .A(n14841), .B(n14842), .ZN(n8609) );
  XNOR2_X1 U14848 ( .A(a_12_), .B(b_12_), .ZN(n14841) );
  OR2_X1 U14849 ( .A1(n14843), .A2(n14844), .ZN(n14732) );
  AND2_X1 U14850 ( .A1(n14726), .A2(n14728), .ZN(n14844) );
  AND2_X1 U14851 ( .A1(n14845), .A2(n14727), .ZN(n14843) );
  OR2_X1 U14852 ( .A1(n8599), .A2(n7666), .ZN(n14727) );
  OR2_X1 U14853 ( .A1(n14728), .A2(n14726), .ZN(n14845) );
  OR2_X1 U14854 ( .A1(n14456), .A2(n7632), .ZN(n14726) );
  XNOR2_X1 U14855 ( .A(n14846), .B(n14847), .ZN(n8604) );
  XNOR2_X1 U14856 ( .A(a_13_), .B(b_13_), .ZN(n14846) );
  OR2_X1 U14857 ( .A1(n14848), .A2(n14849), .ZN(n14728) );
  AND2_X1 U14858 ( .A1(n14722), .A2(n14724), .ZN(n14849) );
  AND2_X1 U14859 ( .A1(n14850), .A2(n14723), .ZN(n14848) );
  OR2_X1 U14860 ( .A1(n8594), .A2(n7666), .ZN(n14723) );
  OR2_X1 U14861 ( .A1(n14724), .A2(n14722), .ZN(n14850) );
  OR2_X1 U14862 ( .A1(n14456), .A2(n7634), .ZN(n14722) );
  XNOR2_X1 U14863 ( .A(n14851), .B(n14852), .ZN(n8599) );
  XNOR2_X1 U14864 ( .A(a_14_), .B(b_14_), .ZN(n14851) );
  OR2_X1 U14865 ( .A1(n14853), .A2(n14854), .ZN(n14724) );
  AND2_X1 U14866 ( .A1(n14718), .A2(n14720), .ZN(n14854) );
  AND2_X1 U14867 ( .A1(n14855), .A2(n14719), .ZN(n14853) );
  OR2_X1 U14868 ( .A1(n8589), .A2(n7666), .ZN(n14719) );
  OR2_X1 U14869 ( .A1(n14720), .A2(n14718), .ZN(n14855) );
  OR2_X1 U14870 ( .A1(n14456), .A2(n7636), .ZN(n14718) );
  XNOR2_X1 U14871 ( .A(n14856), .B(n14857), .ZN(n8594) );
  XNOR2_X1 U14872 ( .A(a_15_), .B(b_15_), .ZN(n14856) );
  OR2_X1 U14873 ( .A1(n14858), .A2(n14859), .ZN(n14720) );
  AND2_X1 U14874 ( .A1(n14714), .A2(n14716), .ZN(n14859) );
  AND2_X1 U14875 ( .A1(n14860), .A2(n14715), .ZN(n14858) );
  OR2_X1 U14876 ( .A1(n8584), .A2(n7666), .ZN(n14715) );
  OR2_X1 U14877 ( .A1(n14716), .A2(n14714), .ZN(n14860) );
  OR2_X1 U14878 ( .A1(n14456), .A2(n7638), .ZN(n14714) );
  XNOR2_X1 U14879 ( .A(n14861), .B(n14862), .ZN(n8589) );
  XNOR2_X1 U14880 ( .A(a_16_), .B(b_16_), .ZN(n14861) );
  OR2_X1 U14881 ( .A1(n14863), .A2(n14864), .ZN(n14716) );
  AND2_X1 U14882 ( .A1(n14710), .A2(n14712), .ZN(n14864) );
  AND2_X1 U14883 ( .A1(n14865), .A2(n14711), .ZN(n14863) );
  OR2_X1 U14884 ( .A1(n8579), .A2(n7666), .ZN(n14711) );
  OR2_X1 U14885 ( .A1(n14712), .A2(n14710), .ZN(n14865) );
  OR2_X1 U14886 ( .A1(n14456), .A2(n7640), .ZN(n14710) );
  XNOR2_X1 U14887 ( .A(n14866), .B(n14867), .ZN(n8584) );
  XNOR2_X1 U14888 ( .A(a_17_), .B(b_17_), .ZN(n14866) );
  OR2_X1 U14889 ( .A1(n14868), .A2(n14869), .ZN(n14712) );
  AND2_X1 U14890 ( .A1(n14706), .A2(n14708), .ZN(n14869) );
  AND2_X1 U14891 ( .A1(n14870), .A2(n14707), .ZN(n14868) );
  OR2_X1 U14892 ( .A1(n8574), .A2(n7666), .ZN(n14707) );
  OR2_X1 U14893 ( .A1(n14708), .A2(n14706), .ZN(n14870) );
  OR2_X1 U14894 ( .A1(n14456), .A2(n7642), .ZN(n14706) );
  XNOR2_X1 U14895 ( .A(n14871), .B(n14872), .ZN(n8579) );
  XNOR2_X1 U14896 ( .A(a_18_), .B(b_18_), .ZN(n14871) );
  OR2_X1 U14897 ( .A1(n14873), .A2(n14874), .ZN(n14708) );
  AND2_X1 U14898 ( .A1(n14702), .A2(n14704), .ZN(n14874) );
  AND2_X1 U14899 ( .A1(n14875), .A2(n14703), .ZN(n14873) );
  OR2_X1 U14900 ( .A1(n8569), .A2(n14651), .ZN(n14703) );
  OR2_X1 U14901 ( .A1(n14704), .A2(n14702), .ZN(n14875) );
  OR2_X1 U14902 ( .A1(n14456), .A2(n7644), .ZN(n14702) );
  XNOR2_X1 U14903 ( .A(n14876), .B(n14877), .ZN(n8574) );
  XNOR2_X1 U14904 ( .A(a_19_), .B(b_19_), .ZN(n14876) );
  OR2_X1 U14905 ( .A1(n14878), .A2(n14879), .ZN(n14704) );
  AND2_X1 U14906 ( .A1(n14698), .A2(n14700), .ZN(n14879) );
  AND2_X1 U14907 ( .A1(n14880), .A2(n14699), .ZN(n14878) );
  OR2_X1 U14908 ( .A1(n8564), .A2(n14651), .ZN(n14699) );
  OR2_X1 U14909 ( .A1(n14700), .A2(n14698), .ZN(n14880) );
  OR2_X1 U14910 ( .A1(n14456), .A2(n7646), .ZN(n14698) );
  XNOR2_X1 U14911 ( .A(n14881), .B(n14882), .ZN(n8569) );
  XNOR2_X1 U14912 ( .A(a_20_), .B(b_20_), .ZN(n14881) );
  OR2_X1 U14913 ( .A1(n14883), .A2(n14884), .ZN(n14700) );
  AND2_X1 U14914 ( .A1(n14694), .A2(n14696), .ZN(n14884) );
  AND2_X1 U14915 ( .A1(n14885), .A2(n14695), .ZN(n14883) );
  OR2_X1 U14916 ( .A1(n8559), .A2(n14651), .ZN(n14695) );
  OR2_X1 U14917 ( .A1(n14696), .A2(n14694), .ZN(n14885) );
  OR2_X1 U14918 ( .A1(n14456), .A2(n7648), .ZN(n14694) );
  XNOR2_X1 U14919 ( .A(n14886), .B(n14887), .ZN(n8564) );
  XNOR2_X1 U14920 ( .A(a_21_), .B(b_21_), .ZN(n14886) );
  OR2_X1 U14921 ( .A1(n14888), .A2(n14889), .ZN(n14696) );
  AND2_X1 U14922 ( .A1(n14690), .A2(n14692), .ZN(n14889) );
  AND2_X1 U14923 ( .A1(n14890), .A2(n14691), .ZN(n14888) );
  OR2_X1 U14924 ( .A1(n8554), .A2(n14651), .ZN(n14691) );
  OR2_X1 U14925 ( .A1(n14692), .A2(n14690), .ZN(n14890) );
  OR2_X1 U14926 ( .A1(n14456), .A2(n7650), .ZN(n14690) );
  XNOR2_X1 U14927 ( .A(n14891), .B(n14892), .ZN(n8559) );
  XNOR2_X1 U14928 ( .A(a_22_), .B(b_22_), .ZN(n14891) );
  OR2_X1 U14929 ( .A1(n14893), .A2(n14894), .ZN(n14692) );
  AND2_X1 U14930 ( .A1(n14686), .A2(n14688), .ZN(n14894) );
  AND2_X1 U14931 ( .A1(n14895), .A2(n14687), .ZN(n14893) );
  OR2_X1 U14932 ( .A1(n8549), .A2(n14651), .ZN(n14687) );
  OR2_X1 U14933 ( .A1(n14688), .A2(n14686), .ZN(n14895) );
  OR2_X1 U14934 ( .A1(n14456), .A2(n7652), .ZN(n14686) );
  XNOR2_X1 U14935 ( .A(n14896), .B(n14897), .ZN(n8554) );
  XNOR2_X1 U14936 ( .A(a_23_), .B(b_23_), .ZN(n14896) );
  OR2_X1 U14937 ( .A1(n14898), .A2(n14899), .ZN(n14688) );
  AND2_X1 U14938 ( .A1(n14682), .A2(n14684), .ZN(n14899) );
  AND2_X1 U14939 ( .A1(n14900), .A2(n14683), .ZN(n14898) );
  OR2_X1 U14940 ( .A1(n8544), .A2(n14651), .ZN(n14683) );
  OR2_X1 U14941 ( .A1(n14684), .A2(n14682), .ZN(n14900) );
  OR2_X1 U14942 ( .A1(n14456), .A2(n7654), .ZN(n14682) );
  XNOR2_X1 U14943 ( .A(n14901), .B(n14902), .ZN(n8549) );
  XNOR2_X1 U14944 ( .A(a_24_), .B(b_24_), .ZN(n14901) );
  OR2_X1 U14945 ( .A1(n14903), .A2(n14904), .ZN(n14684) );
  AND2_X1 U14946 ( .A1(n14678), .A2(n14680), .ZN(n14904) );
  AND2_X1 U14947 ( .A1(n14905), .A2(n14679), .ZN(n14903) );
  OR2_X1 U14948 ( .A1(n8539), .A2(n14651), .ZN(n14679) );
  OR2_X1 U14949 ( .A1(n14680), .A2(n14678), .ZN(n14905) );
  OR2_X1 U14950 ( .A1(n14456), .A2(n7656), .ZN(n14678) );
  XNOR2_X1 U14951 ( .A(n14906), .B(n14907), .ZN(n8544) );
  XNOR2_X1 U14952 ( .A(a_25_), .B(b_25_), .ZN(n14906) );
  OR2_X1 U14953 ( .A1(n14908), .A2(n14909), .ZN(n14680) );
  AND2_X1 U14954 ( .A1(n14674), .A2(n14676), .ZN(n14909) );
  AND2_X1 U14955 ( .A1(n14910), .A2(n14675), .ZN(n14908) );
  OR2_X1 U14956 ( .A1(n8534), .A2(n14651), .ZN(n14675) );
  OR2_X1 U14957 ( .A1(n14676), .A2(n14674), .ZN(n14910) );
  OR2_X1 U14958 ( .A1(n14456), .A2(n7658), .ZN(n14674) );
  XNOR2_X1 U14959 ( .A(n14911), .B(n14912), .ZN(n8539) );
  XNOR2_X1 U14960 ( .A(a_26_), .B(b_26_), .ZN(n14911) );
  OR2_X1 U14961 ( .A1(n14913), .A2(n14914), .ZN(n14676) );
  AND2_X1 U14962 ( .A1(n14669), .A2(n14672), .ZN(n14914) );
  AND2_X1 U14963 ( .A1(n14915), .A2(n14671), .ZN(n14913) );
  OR2_X1 U14964 ( .A1(n8529), .A2(n14651), .ZN(n14671) );
  OR2_X1 U14965 ( .A1(n14672), .A2(n14669), .ZN(n14915) );
  OR2_X1 U14966 ( .A1(n14456), .A2(n7660), .ZN(n14669) );
  XNOR2_X1 U14967 ( .A(n14916), .B(n14917), .ZN(n8534) );
  XNOR2_X1 U14968 ( .A(a_27_), .B(b_27_), .ZN(n14916) );
  OR2_X1 U14969 ( .A1(n14918), .A2(n14919), .ZN(n14672) );
  AND2_X1 U14970 ( .A1(n14663), .A2(n14666), .ZN(n14919) );
  AND2_X1 U14971 ( .A1(n14665), .A2(n14920), .ZN(n14918) );
  OR2_X1 U14972 ( .A1(n14666), .A2(n14663), .ZN(n14920) );
  OR2_X1 U14973 ( .A1(n14456), .A2(n7662), .ZN(n14663) );
  XNOR2_X1 U14974 ( .A(n14921), .B(n14922), .ZN(n8529) );
  XNOR2_X1 U14975 ( .A(a_28_), .B(b_28_), .ZN(n14921) );
  OR2_X1 U14976 ( .A1(n8518), .A2(n14651), .ZN(n14666) );
  AND2_X1 U14977 ( .A1(n14660), .A2(n14657), .ZN(n14665) );
  OR3_X1 U14978 ( .A1(n14456), .A2(n8519), .A3(n7666), .ZN(n14657) );
  OR2_X1 U14979 ( .A1(n14652), .A2(n14650), .ZN(n8519) );
  INV_X1 U14980 ( .A(n7691), .ZN(n14650) );
  AND2_X1 U14981 ( .A1(n14923), .A2(n14924), .ZN(n7691) );
  OR2_X1 U14982 ( .A1(b_31_), .A2(a_31_), .ZN(n14924) );
  OR3_X1 U14983 ( .A1(n14652), .A2(n7666), .A3(n14662), .ZN(n14660) );
  OR2_X1 U14984 ( .A1(n14456), .A2(n8518), .ZN(n14662) );
  XNOR2_X1 U14985 ( .A(n14925), .B(n14926), .ZN(n8518) );
  XNOR2_X1 U14986 ( .A(n14927), .B(a_29_), .ZN(n14926) );
  XOR2_X1 U14987 ( .A(n14923), .B(n14928), .Z(n14652) );
  XOR2_X1 U14988 ( .A(b_30_), .B(a_30_), .Z(n14928) );
  INV_X1 U14989 ( .A(n14929), .ZN(n14923) );
  XNOR2_X1 U14990 ( .A(n14781), .B(n14783), .ZN(n14784) );
  OR2_X1 U14991 ( .A1(n14456), .A2(n7960), .ZN(n14783) );
  XNOR2_X1 U14992 ( .A(n14930), .B(n14931), .ZN(n7960) );
  XOR2_X1 U14993 ( .A(b_0_), .B(a_0_), .Z(n14931) );
  OR2_X1 U14994 ( .A1(n14932), .A2(n14933), .ZN(n14930) );
  AND2_X1 U14995 ( .A1(n14934), .A2(a_1_), .ZN(n14933) );
  AND2_X1 U14996 ( .A1(b_1_), .A2(n14935), .ZN(n14932) );
  OR2_X1 U14997 ( .A1(n14934), .A2(a_1_), .ZN(n14935) );
  INV_X1 U14998 ( .A(n14936), .ZN(n14934) );
  INV_X1 U14999 ( .A(n14451), .ZN(n14456) );
  XOR2_X1 U15000 ( .A(n14937), .B(n14938), .Z(n14451) );
  XNOR2_X1 U15001 ( .A(c_1_), .B(d_1_), .ZN(n14937) );
  OR2_X1 U15002 ( .A1(n8023), .A2(n14651), .ZN(n14781) );
  XNOR2_X1 U15003 ( .A(n14939), .B(n14940), .ZN(n14651) );
  XOR2_X1 U15004 ( .A(d_0_), .B(c_0_), .Z(n14940) );
  OR2_X1 U15005 ( .A1(n14941), .A2(n14942), .ZN(n14939) );
  AND2_X1 U15006 ( .A1(n14943), .A2(c_1_), .ZN(n14942) );
  AND2_X1 U15007 ( .A1(d_1_), .A2(n14944), .ZN(n14941) );
  OR2_X1 U15008 ( .A1(n14943), .A2(c_1_), .ZN(n14944) );
  INV_X1 U15009 ( .A(n14938), .ZN(n14943) );
  OR2_X1 U15010 ( .A1(n14945), .A2(n14946), .ZN(n14938) );
  AND2_X1 U15011 ( .A1(n14668), .A2(n14947), .ZN(n14946) );
  AND2_X1 U15012 ( .A1(n14948), .A2(n14949), .ZN(n14945) );
  INV_X1 U15013 ( .A(d_2_), .ZN(n14949) );
  OR2_X1 U15014 ( .A1(n14947), .A2(n14668), .ZN(n14948) );
  OR2_X1 U15015 ( .A1(n14950), .A2(n14951), .ZN(n14668) );
  AND2_X1 U15016 ( .A1(n14470), .A2(n14952), .ZN(n14951) );
  AND2_X1 U15017 ( .A1(n14953), .A2(n14954), .ZN(n14950) );
  INV_X1 U15018 ( .A(d_3_), .ZN(n14954) );
  OR2_X1 U15019 ( .A1(n14952), .A2(n14470), .ZN(n14953) );
  OR2_X1 U15020 ( .A1(n14955), .A2(n14956), .ZN(n14470) );
  AND2_X1 U15021 ( .A1(n14294), .A2(n14957), .ZN(n14956) );
  AND2_X1 U15022 ( .A1(n14958), .A2(n14959), .ZN(n14955) );
  INV_X1 U15023 ( .A(d_4_), .ZN(n14959) );
  OR2_X1 U15024 ( .A1(n14957), .A2(n14294), .ZN(n14958) );
  OR2_X1 U15025 ( .A1(n14960), .A2(n14961), .ZN(n14294) );
  AND2_X1 U15026 ( .A1(n14111), .A2(n14962), .ZN(n14961) );
  AND2_X1 U15027 ( .A1(n14963), .A2(n14964), .ZN(n14960) );
  INV_X1 U15028 ( .A(d_5_), .ZN(n14964) );
  OR2_X1 U15029 ( .A1(n14962), .A2(n14111), .ZN(n14963) );
  OR2_X1 U15030 ( .A1(n14965), .A2(n14966), .ZN(n14111) );
  AND2_X1 U15031 ( .A1(n13922), .A2(n14967), .ZN(n14966) );
  AND2_X1 U15032 ( .A1(n14968), .A2(n14969), .ZN(n14965) );
  INV_X1 U15033 ( .A(d_6_), .ZN(n14969) );
  OR2_X1 U15034 ( .A1(n14967), .A2(n13922), .ZN(n14968) );
  OR2_X1 U15035 ( .A1(n14970), .A2(n14971), .ZN(n13922) );
  AND2_X1 U15036 ( .A1(n13726), .A2(n14972), .ZN(n14971) );
  AND2_X1 U15037 ( .A1(n14973), .A2(n14974), .ZN(n14970) );
  INV_X1 U15038 ( .A(d_7_), .ZN(n14974) );
  OR2_X1 U15039 ( .A1(n14972), .A2(n13726), .ZN(n14973) );
  OR2_X1 U15040 ( .A1(n14975), .A2(n14976), .ZN(n13726) );
  AND2_X1 U15041 ( .A1(n13523), .A2(n14977), .ZN(n14976) );
  AND2_X1 U15042 ( .A1(n14978), .A2(n14979), .ZN(n14975) );
  INV_X1 U15043 ( .A(d_8_), .ZN(n14979) );
  OR2_X1 U15044 ( .A1(n14977), .A2(n13523), .ZN(n14978) );
  OR2_X1 U15045 ( .A1(n14980), .A2(n14981), .ZN(n13523) );
  AND2_X1 U15046 ( .A1(n13313), .A2(n14982), .ZN(n14981) );
  AND2_X1 U15047 ( .A1(n14983), .A2(n14984), .ZN(n14980) );
  INV_X1 U15048 ( .A(d_9_), .ZN(n14984) );
  OR2_X1 U15049 ( .A1(n14982), .A2(n13313), .ZN(n14983) );
  OR2_X1 U15050 ( .A1(n14985), .A2(n14986), .ZN(n13313) );
  AND2_X1 U15051 ( .A1(n13092), .A2(n14987), .ZN(n14986) );
  AND2_X1 U15052 ( .A1(n14988), .A2(n14989), .ZN(n14985) );
  INV_X1 U15053 ( .A(d_10_), .ZN(n14989) );
  OR2_X1 U15054 ( .A1(n14987), .A2(n13092), .ZN(n14988) );
  OR2_X1 U15055 ( .A1(n14990), .A2(n14991), .ZN(n13092) );
  AND2_X1 U15056 ( .A1(n12822), .A2(n14992), .ZN(n14991) );
  AND2_X1 U15057 ( .A1(n14993), .A2(n14994), .ZN(n14990) );
  INV_X1 U15058 ( .A(d_11_), .ZN(n14994) );
  OR2_X1 U15059 ( .A1(n14992), .A2(n12822), .ZN(n14993) );
  OR2_X1 U15060 ( .A1(n14995), .A2(n14996), .ZN(n12822) );
  AND2_X1 U15061 ( .A1(n12597), .A2(n14997), .ZN(n14996) );
  AND2_X1 U15062 ( .A1(n14998), .A2(n14999), .ZN(n14995) );
  INV_X1 U15063 ( .A(d_12_), .ZN(n14999) );
  OR2_X1 U15064 ( .A1(n14997), .A2(n12597), .ZN(n14998) );
  OR2_X1 U15065 ( .A1(n15000), .A2(n15001), .ZN(n12597) );
  AND2_X1 U15066 ( .A1(n12372), .A2(n15002), .ZN(n15001) );
  AND2_X1 U15067 ( .A1(n15003), .A2(n15004), .ZN(n15000) );
  INV_X1 U15068 ( .A(d_13_), .ZN(n15004) );
  OR2_X1 U15069 ( .A1(n15002), .A2(n12372), .ZN(n15003) );
  OR2_X1 U15070 ( .A1(n15005), .A2(n15006), .ZN(n12372) );
  AND2_X1 U15071 ( .A1(n12148), .A2(n15007), .ZN(n15006) );
  AND2_X1 U15072 ( .A1(n15008), .A2(n15009), .ZN(n15005) );
  INV_X1 U15073 ( .A(d_14_), .ZN(n15009) );
  OR2_X1 U15074 ( .A1(n12148), .A2(n15007), .ZN(n15008) );
  INV_X1 U15075 ( .A(c_14_), .ZN(n15007) );
  OR2_X1 U15076 ( .A1(n15010), .A2(n15011), .ZN(n12148) );
  AND2_X1 U15077 ( .A1(n12044), .A2(n15012), .ZN(n15011) );
  AND2_X1 U15078 ( .A1(n15013), .A2(n15014), .ZN(n15010) );
  INV_X1 U15079 ( .A(d_15_), .ZN(n15014) );
  OR2_X1 U15080 ( .A1(n12044), .A2(n15012), .ZN(n15013) );
  INV_X1 U15081 ( .A(c_15_), .ZN(n15012) );
  OR2_X1 U15082 ( .A1(n15015), .A2(n15016), .ZN(n12044) );
  AND2_X1 U15083 ( .A1(n11833), .A2(n15017), .ZN(n15016) );
  AND2_X1 U15084 ( .A1(n15018), .A2(n15019), .ZN(n15015) );
  INV_X1 U15085 ( .A(d_16_), .ZN(n15019) );
  OR2_X1 U15086 ( .A1(n11833), .A2(n15017), .ZN(n15018) );
  INV_X1 U15087 ( .A(c_16_), .ZN(n15017) );
  OR2_X1 U15088 ( .A1(n15020), .A2(n15021), .ZN(n11833) );
  AND2_X1 U15089 ( .A1(n11598), .A2(n15022), .ZN(n15021) );
  AND2_X1 U15090 ( .A1(n15023), .A2(n15024), .ZN(n15020) );
  INV_X1 U15091 ( .A(d_17_), .ZN(n15024) );
  OR2_X1 U15092 ( .A1(n11598), .A2(n15022), .ZN(n15023) );
  INV_X1 U15093 ( .A(c_17_), .ZN(n15022) );
  OR2_X1 U15094 ( .A1(n15025), .A2(n15026), .ZN(n11598) );
  AND2_X1 U15095 ( .A1(n11422), .A2(n15027), .ZN(n15026) );
  AND2_X1 U15096 ( .A1(n15028), .A2(n15029), .ZN(n15025) );
  INV_X1 U15097 ( .A(d_18_), .ZN(n15029) );
  OR2_X1 U15098 ( .A1(n11422), .A2(n15027), .ZN(n15028) );
  INV_X1 U15099 ( .A(c_18_), .ZN(n15027) );
  OR2_X1 U15100 ( .A1(n15030), .A2(n15031), .ZN(n11422) );
  AND2_X1 U15101 ( .A1(n11239), .A2(n15032), .ZN(n15031) );
  AND2_X1 U15102 ( .A1(n15033), .A2(n15034), .ZN(n15030) );
  INV_X1 U15103 ( .A(d_19_), .ZN(n15034) );
  OR2_X1 U15104 ( .A1(n11239), .A2(n15032), .ZN(n15033) );
  INV_X1 U15105 ( .A(c_19_), .ZN(n15032) );
  OR2_X1 U15106 ( .A1(n15035), .A2(n15036), .ZN(n11239) );
  AND2_X1 U15107 ( .A1(n11050), .A2(n15037), .ZN(n15036) );
  AND2_X1 U15108 ( .A1(n15038), .A2(n15039), .ZN(n15035) );
  INV_X1 U15109 ( .A(d_20_), .ZN(n15039) );
  OR2_X1 U15110 ( .A1(n11050), .A2(n15037), .ZN(n15038) );
  INV_X1 U15111 ( .A(c_20_), .ZN(n15037) );
  OR2_X1 U15112 ( .A1(n15040), .A2(n15041), .ZN(n11050) );
  AND2_X1 U15113 ( .A1(n10854), .A2(n15042), .ZN(n15041) );
  AND2_X1 U15114 ( .A1(n15043), .A2(n15044), .ZN(n15040) );
  INV_X1 U15115 ( .A(d_21_), .ZN(n15044) );
  OR2_X1 U15116 ( .A1(n10854), .A2(n15042), .ZN(n15043) );
  INV_X1 U15117 ( .A(c_21_), .ZN(n15042) );
  OR2_X1 U15118 ( .A1(n15045), .A2(n15046), .ZN(n10854) );
  AND2_X1 U15119 ( .A1(n10535), .A2(n15047), .ZN(n15046) );
  AND2_X1 U15120 ( .A1(n15048), .A2(n15049), .ZN(n15045) );
  INV_X1 U15121 ( .A(d_22_), .ZN(n15049) );
  OR2_X1 U15122 ( .A1(n10535), .A2(n15047), .ZN(n15048) );
  INV_X1 U15123 ( .A(c_22_), .ZN(n15047) );
  OR2_X1 U15124 ( .A1(n15050), .A2(n15051), .ZN(n10535) );
  AND2_X1 U15125 ( .A1(n10354), .A2(n15052), .ZN(n15051) );
  AND2_X1 U15126 ( .A1(n15053), .A2(n15054), .ZN(n15050) );
  INV_X1 U15127 ( .A(d_23_), .ZN(n15054) );
  OR2_X1 U15128 ( .A1(n10354), .A2(n15052), .ZN(n15053) );
  INV_X1 U15129 ( .A(c_23_), .ZN(n15052) );
  OR2_X1 U15130 ( .A1(n15055), .A2(n15056), .ZN(n10354) );
  AND2_X1 U15131 ( .A1(n10160), .A2(n15057), .ZN(n15056) );
  AND2_X1 U15132 ( .A1(n15058), .A2(n15059), .ZN(n15055) );
  INV_X1 U15133 ( .A(d_24_), .ZN(n15059) );
  OR2_X1 U15134 ( .A1(n10160), .A2(n15057), .ZN(n15058) );
  INV_X1 U15135 ( .A(c_24_), .ZN(n15057) );
  OR2_X1 U15136 ( .A1(n15060), .A2(n15061), .ZN(n10160) );
  AND2_X1 U15137 ( .A1(n9967), .A2(n15062), .ZN(n15061) );
  AND2_X1 U15138 ( .A1(n15063), .A2(n15064), .ZN(n15060) );
  INV_X1 U15139 ( .A(d_25_), .ZN(n15064) );
  OR2_X1 U15140 ( .A1(n9967), .A2(n15062), .ZN(n15063) );
  INV_X1 U15141 ( .A(c_25_), .ZN(n15062) );
  OR2_X1 U15142 ( .A1(n15065), .A2(n15066), .ZN(n9967) );
  AND2_X1 U15143 ( .A1(n9764), .A2(n15067), .ZN(n15066) );
  AND2_X1 U15144 ( .A1(n15068), .A2(n15069), .ZN(n15065) );
  INV_X1 U15145 ( .A(d_26_), .ZN(n15069) );
  OR2_X1 U15146 ( .A1(n9764), .A2(n15067), .ZN(n15068) );
  INV_X1 U15147 ( .A(c_26_), .ZN(n15067) );
  OR2_X1 U15148 ( .A1(n15070), .A2(n15071), .ZN(n9764) );
  AND2_X1 U15149 ( .A1(n9554), .A2(n15072), .ZN(n15071) );
  AND2_X1 U15150 ( .A1(n15073), .A2(n15074), .ZN(n15070) );
  INV_X1 U15151 ( .A(d_27_), .ZN(n15074) );
  OR2_X1 U15152 ( .A1(n9554), .A2(n15072), .ZN(n15073) );
  INV_X1 U15153 ( .A(c_27_), .ZN(n15072) );
  OR2_X1 U15154 ( .A1(n15075), .A2(n15076), .ZN(n9554) );
  AND2_X1 U15155 ( .A1(n9306), .A2(n15077), .ZN(n15076) );
  AND2_X1 U15156 ( .A1(n15078), .A2(n15079), .ZN(n15075) );
  INV_X1 U15157 ( .A(d_28_), .ZN(n15079) );
  OR2_X1 U15158 ( .A1(n9306), .A2(n15077), .ZN(n15078) );
  INV_X1 U15159 ( .A(c_28_), .ZN(n15077) );
  OR2_X1 U15160 ( .A1(n15080), .A2(n15081), .ZN(n9306) );
  AND2_X1 U15161 ( .A1(n9099), .A2(n15082), .ZN(n15081) );
  AND2_X1 U15162 ( .A1(n15083), .A2(n9101), .ZN(n15080) );
  INV_X1 U15163 ( .A(d_29_), .ZN(n9101) );
  OR2_X1 U15164 ( .A1(n9099), .A2(n15082), .ZN(n15083) );
  INV_X1 U15165 ( .A(c_29_), .ZN(n15082) );
  INV_X1 U15166 ( .A(n15084), .ZN(n9099) );
  OR2_X1 U15167 ( .A1(n15085), .A2(n15086), .ZN(n15084) );
  AND2_X1 U15168 ( .A1(c_30_), .A2(n8667), .ZN(n15086) );
  AND2_X1 U15169 ( .A1(d_30_), .A2(n15087), .ZN(n15085) );
  OR2_X1 U15170 ( .A1(n8667), .A2(c_30_), .ZN(n15087) );
  AND2_X1 U15171 ( .A1(c_31_), .A2(d_31_), .ZN(n8667) );
  INV_X1 U15172 ( .A(c_13_), .ZN(n15002) );
  INV_X1 U15173 ( .A(c_12_), .ZN(n14997) );
  INV_X1 U15174 ( .A(c_11_), .ZN(n14992) );
  INV_X1 U15175 ( .A(c_10_), .ZN(n14987) );
  INV_X1 U15176 ( .A(c_9_), .ZN(n14982) );
  INV_X1 U15177 ( .A(c_8_), .ZN(n14977) );
  INV_X1 U15178 ( .A(c_7_), .ZN(n14972) );
  INV_X1 U15179 ( .A(c_6_), .ZN(n14967) );
  INV_X1 U15180 ( .A(c_5_), .ZN(n14962) );
  INV_X1 U15181 ( .A(c_4_), .ZN(n14957) );
  INV_X1 U15182 ( .A(c_3_), .ZN(n14952) );
  INV_X1 U15183 ( .A(c_2_), .ZN(n14947) );
  XNOR2_X1 U15184 ( .A(n15088), .B(n14936), .ZN(n8023) );
  OR2_X1 U15185 ( .A1(n15089), .A2(n15090), .ZN(n14936) );
  AND2_X1 U15186 ( .A1(n14792), .A2(n15091), .ZN(n15090) );
  AND2_X1 U15187 ( .A1(n15092), .A2(n15093), .ZN(n15089) );
  INV_X1 U15188 ( .A(b_2_), .ZN(n15093) );
  OR2_X1 U15189 ( .A1(n15091), .A2(n14792), .ZN(n15092) );
  OR2_X1 U15190 ( .A1(n15094), .A2(n15095), .ZN(n14792) );
  AND2_X1 U15191 ( .A1(n14797), .A2(n15096), .ZN(n15095) );
  AND2_X1 U15192 ( .A1(n15097), .A2(n15098), .ZN(n15094) );
  INV_X1 U15193 ( .A(b_3_), .ZN(n15098) );
  OR2_X1 U15194 ( .A1(n15096), .A2(n14797), .ZN(n15097) );
  OR2_X1 U15195 ( .A1(n15099), .A2(n15100), .ZN(n14797) );
  AND2_X1 U15196 ( .A1(n14802), .A2(n15101), .ZN(n15100) );
  AND2_X1 U15197 ( .A1(n15102), .A2(n15103), .ZN(n15099) );
  INV_X1 U15198 ( .A(b_4_), .ZN(n15103) );
  OR2_X1 U15199 ( .A1(n15101), .A2(n14802), .ZN(n15102) );
  OR2_X1 U15200 ( .A1(n15104), .A2(n15105), .ZN(n14802) );
  AND2_X1 U15201 ( .A1(n14807), .A2(n15106), .ZN(n15105) );
  AND2_X1 U15202 ( .A1(n15107), .A2(n15108), .ZN(n15104) );
  INV_X1 U15203 ( .A(b_5_), .ZN(n15108) );
  OR2_X1 U15204 ( .A1(n15106), .A2(n14807), .ZN(n15107) );
  OR2_X1 U15205 ( .A1(n15109), .A2(n15110), .ZN(n14807) );
  AND2_X1 U15206 ( .A1(n14812), .A2(n15111), .ZN(n15110) );
  AND2_X1 U15207 ( .A1(n15112), .A2(n15113), .ZN(n15109) );
  INV_X1 U15208 ( .A(b_6_), .ZN(n15113) );
  OR2_X1 U15209 ( .A1(n15111), .A2(n14812), .ZN(n15112) );
  OR2_X1 U15210 ( .A1(n15114), .A2(n15115), .ZN(n14812) );
  AND2_X1 U15211 ( .A1(n14817), .A2(n15116), .ZN(n15115) );
  AND2_X1 U15212 ( .A1(n15117), .A2(n15118), .ZN(n15114) );
  INV_X1 U15213 ( .A(b_7_), .ZN(n15118) );
  OR2_X1 U15214 ( .A1(n15116), .A2(n14817), .ZN(n15117) );
  OR2_X1 U15215 ( .A1(n15119), .A2(n15120), .ZN(n14817) );
  AND2_X1 U15216 ( .A1(n14822), .A2(n15121), .ZN(n15120) );
  AND2_X1 U15217 ( .A1(n15122), .A2(n15123), .ZN(n15119) );
  INV_X1 U15218 ( .A(b_8_), .ZN(n15123) );
  OR2_X1 U15219 ( .A1(n15121), .A2(n14822), .ZN(n15122) );
  OR2_X1 U15220 ( .A1(n15124), .A2(n15125), .ZN(n14822) );
  AND2_X1 U15221 ( .A1(n14827), .A2(n15126), .ZN(n15125) );
  AND2_X1 U15222 ( .A1(n15127), .A2(n15128), .ZN(n15124) );
  INV_X1 U15223 ( .A(b_9_), .ZN(n15128) );
  OR2_X1 U15224 ( .A1(n15126), .A2(n14827), .ZN(n15127) );
  OR2_X1 U15225 ( .A1(n15129), .A2(n15130), .ZN(n14827) );
  AND2_X1 U15226 ( .A1(n14832), .A2(n15131), .ZN(n15130) );
  AND2_X1 U15227 ( .A1(n15132), .A2(n15133), .ZN(n15129) );
  INV_X1 U15228 ( .A(b_10_), .ZN(n15133) );
  OR2_X1 U15229 ( .A1(n15131), .A2(n14832), .ZN(n15132) );
  OR2_X1 U15230 ( .A1(n15134), .A2(n15135), .ZN(n14832) );
  AND2_X1 U15231 ( .A1(n14837), .A2(n15136), .ZN(n15135) );
  AND2_X1 U15232 ( .A1(n15137), .A2(n15138), .ZN(n15134) );
  INV_X1 U15233 ( .A(b_11_), .ZN(n15138) );
  OR2_X1 U15234 ( .A1(n15136), .A2(n14837), .ZN(n15137) );
  OR2_X1 U15235 ( .A1(n15139), .A2(n15140), .ZN(n14837) );
  AND2_X1 U15236 ( .A1(n14842), .A2(n15141), .ZN(n15140) );
  AND2_X1 U15237 ( .A1(n15142), .A2(n15143), .ZN(n15139) );
  INV_X1 U15238 ( .A(b_12_), .ZN(n15143) );
  OR2_X1 U15239 ( .A1(n15141), .A2(n14842), .ZN(n15142) );
  OR2_X1 U15240 ( .A1(n15144), .A2(n15145), .ZN(n14842) );
  AND2_X1 U15241 ( .A1(n14847), .A2(n15146), .ZN(n15145) );
  AND2_X1 U15242 ( .A1(n15147), .A2(n15148), .ZN(n15144) );
  INV_X1 U15243 ( .A(b_13_), .ZN(n15148) );
  OR2_X1 U15244 ( .A1(n15146), .A2(n14847), .ZN(n15147) );
  OR2_X1 U15245 ( .A1(n15149), .A2(n15150), .ZN(n14847) );
  AND2_X1 U15246 ( .A1(n14852), .A2(n15151), .ZN(n15150) );
  AND2_X1 U15247 ( .A1(n15152), .A2(n15153), .ZN(n15149) );
  INV_X1 U15248 ( .A(b_14_), .ZN(n15153) );
  OR2_X1 U15249 ( .A1(n15151), .A2(n14852), .ZN(n15152) );
  OR2_X1 U15250 ( .A1(n15154), .A2(n15155), .ZN(n14852) );
  AND2_X1 U15251 ( .A1(n14857), .A2(n15156), .ZN(n15155) );
  AND2_X1 U15252 ( .A1(n15157), .A2(n15158), .ZN(n15154) );
  INV_X1 U15253 ( .A(b_15_), .ZN(n15158) );
  OR2_X1 U15254 ( .A1(n15156), .A2(n14857), .ZN(n15157) );
  OR2_X1 U15255 ( .A1(n15159), .A2(n15160), .ZN(n14857) );
  AND2_X1 U15256 ( .A1(n14862), .A2(n15161), .ZN(n15160) );
  AND2_X1 U15257 ( .A1(n15162), .A2(n15163), .ZN(n15159) );
  INV_X1 U15258 ( .A(b_16_), .ZN(n15163) );
  OR2_X1 U15259 ( .A1(n15161), .A2(n14862), .ZN(n15162) );
  OR2_X1 U15260 ( .A1(n15164), .A2(n15165), .ZN(n14862) );
  AND2_X1 U15261 ( .A1(n14867), .A2(n15166), .ZN(n15165) );
  AND2_X1 U15262 ( .A1(n15167), .A2(n15168), .ZN(n15164) );
  INV_X1 U15263 ( .A(b_17_), .ZN(n15168) );
  OR2_X1 U15264 ( .A1(n15166), .A2(n14867), .ZN(n15167) );
  OR2_X1 U15265 ( .A1(n15169), .A2(n15170), .ZN(n14867) );
  AND2_X1 U15266 ( .A1(n14872), .A2(n15171), .ZN(n15170) );
  AND2_X1 U15267 ( .A1(n15172), .A2(n15173), .ZN(n15169) );
  INV_X1 U15268 ( .A(b_18_), .ZN(n15173) );
  OR2_X1 U15269 ( .A1(n15171), .A2(n14872), .ZN(n15172) );
  OR2_X1 U15270 ( .A1(n15174), .A2(n15175), .ZN(n14872) );
  AND2_X1 U15271 ( .A1(n14877), .A2(n15176), .ZN(n15175) );
  AND2_X1 U15272 ( .A1(n15177), .A2(n15178), .ZN(n15174) );
  INV_X1 U15273 ( .A(b_19_), .ZN(n15178) );
  OR2_X1 U15274 ( .A1(n15176), .A2(n14877), .ZN(n15177) );
  OR2_X1 U15275 ( .A1(n15179), .A2(n15180), .ZN(n14877) );
  AND2_X1 U15276 ( .A1(n14882), .A2(n15181), .ZN(n15180) );
  AND2_X1 U15277 ( .A1(n15182), .A2(n15183), .ZN(n15179) );
  INV_X1 U15278 ( .A(b_20_), .ZN(n15183) );
  OR2_X1 U15279 ( .A1(n15181), .A2(n14882), .ZN(n15182) );
  OR2_X1 U15280 ( .A1(n15184), .A2(n15185), .ZN(n14882) );
  AND2_X1 U15281 ( .A1(n14887), .A2(n15186), .ZN(n15185) );
  AND2_X1 U15282 ( .A1(n15187), .A2(n15188), .ZN(n15184) );
  INV_X1 U15283 ( .A(b_21_), .ZN(n15188) );
  OR2_X1 U15284 ( .A1(n15186), .A2(n14887), .ZN(n15187) );
  OR2_X1 U15285 ( .A1(n15189), .A2(n15190), .ZN(n14887) );
  AND2_X1 U15286 ( .A1(n14892), .A2(n15191), .ZN(n15190) );
  AND2_X1 U15287 ( .A1(n15192), .A2(n15193), .ZN(n15189) );
  INV_X1 U15288 ( .A(b_22_), .ZN(n15193) );
  OR2_X1 U15289 ( .A1(n15191), .A2(n14892), .ZN(n15192) );
  OR2_X1 U15290 ( .A1(n15194), .A2(n15195), .ZN(n14892) );
  AND2_X1 U15291 ( .A1(n14897), .A2(n15196), .ZN(n15195) );
  AND2_X1 U15292 ( .A1(n15197), .A2(n15198), .ZN(n15194) );
  INV_X1 U15293 ( .A(b_23_), .ZN(n15198) );
  OR2_X1 U15294 ( .A1(n15196), .A2(n14897), .ZN(n15197) );
  OR2_X1 U15295 ( .A1(n15199), .A2(n15200), .ZN(n14897) );
  AND2_X1 U15296 ( .A1(n14902), .A2(n15201), .ZN(n15200) );
  AND2_X1 U15297 ( .A1(n15202), .A2(n15203), .ZN(n15199) );
  INV_X1 U15298 ( .A(b_24_), .ZN(n15203) );
  OR2_X1 U15299 ( .A1(n15201), .A2(n14902), .ZN(n15202) );
  OR2_X1 U15300 ( .A1(n15204), .A2(n15205), .ZN(n14902) );
  AND2_X1 U15301 ( .A1(n14907), .A2(n15206), .ZN(n15205) );
  AND2_X1 U15302 ( .A1(n15207), .A2(n15208), .ZN(n15204) );
  INV_X1 U15303 ( .A(b_25_), .ZN(n15208) );
  OR2_X1 U15304 ( .A1(n15206), .A2(n14907), .ZN(n15207) );
  OR2_X1 U15305 ( .A1(n15209), .A2(n15210), .ZN(n14907) );
  AND2_X1 U15306 ( .A1(n14912), .A2(n15211), .ZN(n15210) );
  AND2_X1 U15307 ( .A1(n15212), .A2(n15213), .ZN(n15209) );
  INV_X1 U15308 ( .A(b_26_), .ZN(n15213) );
  OR2_X1 U15309 ( .A1(n15211), .A2(n14912), .ZN(n15212) );
  OR2_X1 U15310 ( .A1(n15214), .A2(n15215), .ZN(n14912) );
  AND2_X1 U15311 ( .A1(n14917), .A2(n15216), .ZN(n15215) );
  AND2_X1 U15312 ( .A1(n15217), .A2(n15218), .ZN(n15214) );
  INV_X1 U15313 ( .A(b_27_), .ZN(n15218) );
  OR2_X1 U15314 ( .A1(n15216), .A2(n14917), .ZN(n15217) );
  OR2_X1 U15315 ( .A1(n15219), .A2(n15220), .ZN(n14917) );
  AND2_X1 U15316 ( .A1(n14922), .A2(n15221), .ZN(n15220) );
  AND2_X1 U15317 ( .A1(n15222), .A2(n15223), .ZN(n15219) );
  INV_X1 U15318 ( .A(b_28_), .ZN(n15223) );
  OR2_X1 U15319 ( .A1(n15221), .A2(n14922), .ZN(n15222) );
  OR2_X1 U15320 ( .A1(n15224), .A2(n15225), .ZN(n14922) );
  AND2_X1 U15321 ( .A1(n15226), .A2(n15227), .ZN(n15225) );
  AND2_X1 U15322 ( .A1(n15228), .A2(n14927), .ZN(n15224) );
  INV_X1 U15323 ( .A(b_29_), .ZN(n14927) );
  OR2_X1 U15324 ( .A1(n15226), .A2(n15227), .ZN(n15228) );
  INV_X1 U15325 ( .A(a_29_), .ZN(n15227) );
  INV_X1 U15326 ( .A(n14925), .ZN(n15226) );
  OR2_X1 U15327 ( .A1(n15229), .A2(n15230), .ZN(n14925) );
  AND2_X1 U15328 ( .A1(n14929), .A2(a_30_), .ZN(n15230) );
  AND2_X1 U15329 ( .A1(b_30_), .A2(n15231), .ZN(n15229) );
  OR2_X1 U15330 ( .A1(n14929), .A2(a_30_), .ZN(n15231) );
  AND2_X1 U15331 ( .A1(a_31_), .A2(b_31_), .ZN(n14929) );
  INV_X1 U15332 ( .A(a_28_), .ZN(n15221) );
  INV_X1 U15333 ( .A(a_27_), .ZN(n15216) );
  INV_X1 U15334 ( .A(a_26_), .ZN(n15211) );
  INV_X1 U15335 ( .A(a_25_), .ZN(n15206) );
  INV_X1 U15336 ( .A(a_24_), .ZN(n15201) );
  INV_X1 U15337 ( .A(a_23_), .ZN(n15196) );
  INV_X1 U15338 ( .A(a_22_), .ZN(n15191) );
  INV_X1 U15339 ( .A(a_21_), .ZN(n15186) );
  INV_X1 U15340 ( .A(a_20_), .ZN(n15181) );
  INV_X1 U15341 ( .A(a_19_), .ZN(n15176) );
  INV_X1 U15342 ( .A(a_18_), .ZN(n15171) );
  INV_X1 U15343 ( .A(a_17_), .ZN(n15166) );
  INV_X1 U15344 ( .A(a_16_), .ZN(n15161) );
  INV_X1 U15345 ( .A(a_15_), .ZN(n15156) );
  INV_X1 U15346 ( .A(a_14_), .ZN(n15151) );
  INV_X1 U15347 ( .A(a_13_), .ZN(n15146) );
  INV_X1 U15348 ( .A(a_12_), .ZN(n15141) );
  INV_X1 U15349 ( .A(a_11_), .ZN(n15136) );
  INV_X1 U15350 ( .A(a_10_), .ZN(n15131) );
  INV_X1 U15351 ( .A(a_9_), .ZN(n15126) );
  INV_X1 U15352 ( .A(a_8_), .ZN(n15121) );
  INV_X1 U15353 ( .A(a_7_), .ZN(n15116) );
  INV_X1 U15354 ( .A(a_6_), .ZN(n15111) );
  INV_X1 U15355 ( .A(a_5_), .ZN(n15106) );
  INV_X1 U15356 ( .A(a_4_), .ZN(n15101) );
  INV_X1 U15357 ( .A(a_3_), .ZN(n15096) );
  INV_X1 U15358 ( .A(a_2_), .ZN(n15091) );
  XNOR2_X1 U15359 ( .A(a_1_), .B(b_1_), .ZN(n15088) );
endmodule

