module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n1359_, new_n595_, new_n1233_, new_n445_, new_n1009_, new_n238_, new_n479_, new_n1105_, new_n1215_, new_n1448_, new_n608_, new_n501_, new_n1157_, new_n1442_, new_n1345_, new_n421_, new_n777_, new_n1433_, new_n1517_, new_n1575_, new_n1472_, new_n1048_, new_n885_, new_n439_, new_n1532_, new_n283_, new_n223_, new_n390_, new_n743_, new_n1327_, new_n241_, new_n1535_, new_n566_, new_n641_, new_n339_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n1351_, new_n556_, new_n636_, new_n691_, new_n1024_, new_n670_, new_n456_, new_n1125_, new_n1590_, new_n246_, new_n911_, new_n679_, new_n937_, new_n667_, new_n367_, new_n1237_, new_n1568_, new_n728_, new_n1479_, new_n1071_, new_n1294_, new_n214_, new_n894_, new_n853_, new_n695_, new_n660_, new_n1311_, new_n526_, new_n908_, new_n552_, new_n678_, new_n342_, new_n706_, new_n649_, new_n1119_, new_n1213_, new_n752_, new_n1524_, new_n1045_, new_n1305_, new_n500_, new_n1163_, new_n786_, new_n317_, new_n1188_, new_n1415_, new_n1390_, new_n721_, new_n504_, new_n1414_, new_n742_, new_n892_, new_n1368_, new_n234_, new_n472_, new_n873_, new_n1167_, new_n1530_, new_n1300_, new_n1490_, new_n774_, new_n792_, new_n1620_, new_n953_, new_n257_, new_n481_, new_n1265_, new_n1073_, new_n1110_, new_n1580_, new_n449_, new_n580_, new_n639_, new_n484_, new_n766_, new_n272_, new_n282_, new_n1262_, new_n1212_, new_n1059_, new_n634_, new_n1332_, new_n1447_, new_n635_, new_n685_, new_n326_, new_n648_, new_n903_, new_n1595_, new_n983_, new_n822_, new_n1406_, new_n1082_, new_n1018_, new_n606_, new_n796_, new_n1054_, new_n655_, new_n1288_, new_n630_, new_n385_, new_n1049_, new_n1330_, new_n694_, new_n461_, new_n1323_, new_n297_, new_n565_, new_n1196_, new_n1366_, new_n511_, new_n303_, new_n1640_, new_n325_, new_n1285_, new_n1031_, new_n1216_, new_n1632_, new_n1281_, new_n629_, new_n1214_, new_n883_, new_n1005_, new_n999_, new_n321_, new_n1647_, new_n324_, new_n960_, new_n1377_, new_n1522_, new_n549_, new_n491_, new_n676_, new_n995_, new_n1035_, new_n271_, new_n674_, new_n274_, new_n991_, new_n1362_, new_n1404_, new_n1443_, new_n1484_, new_n1512_, new_n497_, new_n816_, new_n1355_, new_n568_, new_n420_, new_n876_, new_n423_, new_n498_, new_n496_, new_n1217_, new_n1046_, new_n1182_, new_n708_, new_n206_, new_n1463_, new_n429_, new_n1222_, new_n353_, new_n734_, new_n912_, new_n1424_, new_n1062_, new_n680_, new_n981_, new_n506_, new_n872_, new_n1527_, new_n1275_, new_n1277_, new_n1198_, new_n1428_, new_n1440_, new_n656_, new_n1127_, new_n388_, new_n1028_, new_n1168_, new_n483_, new_n1004_, new_n1152_, new_n1558_, new_n299_, new_n394_, new_n935_, new_n657_, new_n1150_, new_n652_, new_n582_, new_n363_, new_n1266_, new_n1113_, new_n785_, new_n1501_, new_n441_, new_n477_, new_n664_, new_n600_, new_n280_, new_n1041_, new_n1657_, new_n1562_, new_n426_, new_n1036_, new_n235_, new_n398_, new_n1576_, new_n301_, new_n1333_, new_n1132_, new_n395_, new_n383_, new_n343_, new_n854_, new_n458_, new_n1106_, new_n207_, new_n267_, new_n1395_, new_n473_, new_n1624_, new_n1147_, new_n1373_, new_n1229_, new_n1422_, new_n1523_, new_n1468_, new_n969_, new_n334_, new_n331_, new_n1234_, new_n835_, new_n1360_, new_n378_, new_n1574_, new_n1614_, new_n621_, new_n1423_, new_n1637_, new_n244_, new_n705_, new_n943_, new_n874_, new_n402_, new_n1321_, new_n1209_, new_n335_, new_n347_, new_n659_, new_n700_, new_n1419_, new_n921_, new_n346_, new_n396_, new_n1315_, new_n1003_, new_n696_, new_n208_, new_n1507_, new_n1439_, new_n1658_, new_n1365_, new_n1239_, new_n528_, new_n952_, new_n729_, new_n1111_, new_n1413_, new_n1218_, new_n1385_, new_n1346_, new_n1201_, new_n559_, new_n1282_, new_n1630_, new_n762_, new_n1349_, new_n1193_, new_n1547_, new_n1437_, new_n1598_, new_n1187_, new_n1205_, new_n1154_, new_n1253_, new_n1546_, new_n295_, new_n1453_, new_n1256_, new_n628_, new_n1513_, new_n409_, new_n1090_, new_n745_, new_n1489_, new_n553_, new_n1114_, new_n1084_, new_n1061_, new_n668_, new_n333_, new_n290_, new_n834_, new_n1573_, new_n369_, new_n1032_, new_n867_, new_n954_, new_n1591_, new_n1626_, new_n276_, new_n1545_, new_n901_, new_n688_, new_n1255_, new_n410_, new_n985_, new_n851_, new_n1518_, new_n932_, new_n878_, new_n543_, new_n886_, new_n371_, new_n509_, new_n202_, new_n296_, new_n661_, new_n797_, new_n232_, new_n1358_, new_n724_, new_n1070_, new_n1416_, new_n1109_, new_n261_, new_n672_, new_n1496_, new_n1269_, new_n616_, new_n1653_, new_n529_, new_n323_, new_n914_, new_n884_, new_n938_, new_n362_, new_n1600_, new_n1592_, new_n809_, new_n1631_, new_n1142_, new_n1623_, new_n604_, new_n1461_, new_n1104_, new_n1511_, new_n571_, new_n1504_, new_n758_, new_n460_, new_n1267_, new_n328_, new_n268_, new_n1466_, new_n1516_, new_n1299_, new_n380_, new_n1477_, new_n1079_, new_n861_, new_n1564_, new_n1656_, new_n1252_, new_n352_, new_n1553_, new_n931_, new_n575_, new_n1493_, new_n562_, new_n1593_, new_n944_, new_n1542_, new_n1064_, new_n1065_, new_n1118_, new_n1645_, new_n493_, new_n547_, new_n1480_, new_n264_, new_n379_, new_n273_, new_n224_, new_n586_, new_n963_, new_n1481_, new_n1325_, new_n993_, new_n1625_, new_n1357_, new_n1191_, new_n824_, new_n1628_, new_n717_, new_n1455_, new_n403_, new_n868_, new_n1242_, new_n475_, new_n237_, new_n858_, new_n1612_, new_n1384_, new_n1343_, new_n936_, new_n1459_, new_n1434_, new_n1438_, new_n1016_, new_n411_, new_n673_, new_n1144_, new_n1465_, new_n666_, new_n1290_, new_n407_, new_n1519_, new_n1407_, new_n879_, new_n1417_, new_n736_, new_n513_, new_n558_, new_n219_, new_n382_, new_n313_, new_n1370_, new_n239_, new_n718_, new_n1310_, new_n1398_, new_n1126_, new_n546_, new_n612_, new_n1015_, new_n919_, new_n302_, new_n755_, new_n1040_, new_n1635_, new_n1509_, new_n1559_, new_n544_, new_n615_, new_n722_, new_n856_, new_n415_, new_n1324_, new_n1293_, new_n537_, new_n1336_, new_n345_, new_n499_, new_n533_, new_n255_, new_n1130_, new_n795_, new_n459_, new_n1122_, new_n1185_, new_n1240_, new_n1510_, new_n354_, new_n1174_, new_n968_, new_n1655_, new_n1464_, new_n613_, new_n1508_, new_n337_, new_n1195_, new_n417_, new_n658_, new_n837_, new_n591_, new_n801_, new_n1458_, new_n631_, new_n453_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n1521_, new_n1334_, new_n531_, new_n593_, new_n1543_, new_n974_, new_n1565_, new_n252_, new_n1248_, new_n751_, new_n1038_, new_n372_, new_n852_, new_n1454_, new_n1474_, new_n1328_, new_n978_, new_n1308_, new_n408_, new_n1430_, new_n470_, new_n213_, new_n769_, new_n433_, new_n871_, new_n1450_, new_n992_, new_n1098_, new_n265_, new_n732_, new_n689_, new_n933_, new_n584_, new_n815_, new_n1608_, new_n1492_, new_n1367_, new_n1619_, new_n278_, new_n304_, new_n1052_, new_n1425_, new_n857_, new_n1379_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n269_, new_n512_, new_n1471_, new_n1220_, new_n989_, new_n1117_, new_n1421_, new_n644_, new_n1594_, new_n836_, new_n1116_, new_n904_, new_n1392_, new_n1276_, new_n1444_, new_n913_, new_n327_, new_n681_, new_n594_, new_n561_, new_n495_, new_n927_, new_n431_, new_n1206_, new_n1427_, new_n818_, new_n881_, new_n1268_, new_n1376_, new_n1381_, new_n1566_, new_n1534_, new_n684_, new_n640_, new_n1274_, new_n754_, new_n653_, new_n905_, new_n377_, new_n1258_, new_n1539_, new_n1643_, new_n375_, new_n962_, new_n760_, new_n627_, new_n1391_, new_n1436_, new_n567_, new_n1353_, new_n1033_, new_n576_, new_n831_, new_n791_, new_n1153_, new_n357_, new_n1339_, new_n320_, new_n984_, new_n780_, new_n1183_, new_n245_, new_n643_, new_n1316_, new_n1194_, new_n1338_, new_n1460_, new_n1230_, new_n1602_, new_n1027_, new_n348_, new_n610_, new_n1369_, new_n843_, new_n322_, new_n703_, new_n698_, new_n1639_, new_n1165_, new_n1401_, new_n1259_, new_n226_, new_n1208_, new_n697_, new_n1099_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n1235_, new_n1320_, new_n540_, new_n1149_, new_n1066_, new_n434_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n686_, new_n293_, new_n934_, new_n1567_, new_n1651_, new_n770_, new_n1389_, new_n1400_, new_n757_, new_n1225_, new_n521_, new_n793_, new_n406_, new_n1597_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n1616_, new_n1089_, new_n1192_, new_n405_, new_n942_, new_n614_, new_n895_, new_n958_, new_n976_, new_n699_, new_n236_, new_n1405_, new_n1249_, new_n1354_, new_n955_, new_n847_, new_n250_, new_n888_, new_n1505_, new_n288_, new_n798_, new_n1180_, new_n817_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1410_, new_n941_, new_n738_, new_n827_, new_n1356_, new_n1363_, new_n1317_, new_n366_, new_n779_, new_n1232_, new_n1025_, new_n365_, new_n859_, new_n1211_, new_n1412_, new_n1207_, new_n1374_, new_n601_, new_n842_, new_n1552_, new_n1057_, new_n1644_, new_n682_, new_n1075_, new_n812_, new_n1563_, new_n266_, new_n821_, new_n542_, new_n548_, new_n669_, new_n1397_, new_n220_, new_n1402_, new_n1313_, new_n1172_, new_n419_, new_n624_, new_n534_, new_n1131_, new_n819_, new_n637_, new_n1603_, new_n451_, new_n489_, new_n804_, new_n1342_, new_n424_, new_n602_, new_n1210_, new_n1060_, new_n1303_, new_n240_, new_n413_, new_n1544_, new_n1382_, new_n442_, new_n677_, new_n1487_, new_n1646_, new_n642_, new_n211_, new_n1418_, new_n462_, new_n603_, new_n564_, new_n1528_, new_n761_, new_n840_, new_n735_, new_n1283_, new_n898_, new_n799_, new_n1304_, new_n1537_, new_n946_, new_n344_, new_n287_, new_n1108_, new_n1469_, new_n862_, new_n1606_, new_n427_, new_n532_, new_n393_, new_n418_, new_n746_, new_n1221_, new_n292_, new_n1585_, new_n1587_, new_n1264_, new_n215_, new_n626_, new_n1473_, new_n959_, new_n990_, new_n1629_, new_n716_, new_n701_, new_n1238_, new_n1058_, new_n1162_, new_n212_, new_n1278_, new_n902_, new_n364_, new_n832_, new_n414_, new_n1250_, new_n315_, new_n1482_, new_n1050_, new_n554_, new_n230_, new_n1151_, new_n844_, new_n1302_, new_n281_, new_n430_, new_n482_, new_n849_, new_n1203_, new_n855_, new_n1037_, new_n589_, new_n248_, new_n350_, new_n759_, new_n1083_, new_n1297_, new_n829_, new_n1257_, new_n1306_, new_n988_, new_n478_, new_n1307_, new_n1228_, new_n710_, new_n1486_, new_n361_, new_n764_, new_n906_, new_n683_, new_n1409_, new_n1429_, new_n463_, new_n1372_, new_n510_, new_n351_, new_n1184_, new_n1292_, new_n1426_, new_n517_, new_n609_, new_n530_, new_n890_, new_n318_, new_n1006_, new_n622_, new_n702_, new_n833_, new_n1560_, new_n715_, new_n811_, new_n1445_, new_n1371_, new_n443_, new_n1086_, new_n763_, new_n1622_, new_n1138_, new_n486_, new_n970_, new_n466_, new_n262_, new_n1618_, new_n1652_, new_n218_, new_n1170_, new_n845_, new_n768_, new_n773_, new_n305_, new_n1452_, new_n1051_, new_n899_, new_n1053_, new_n1540_, new_n1611_, new_n205_, new_n492_, new_n1200_, new_n1533_, new_n650_, new_n750_, new_n887_, new_n254_, new_n355_, new_n926_, new_n432_, new_n925_, new_n875_, new_n256_, new_n1226_, new_n778_, new_n452_, new_n381_, new_n1483_, new_n1219_, new_n920_, new_n1121_, new_n1495_, new_n1341_, new_n820_, new_n1386_, new_n771_, new_n979_, new_n508_, new_n1435_, new_n714_, new_n1280_, new_n1007_, new_n1613_, new_n1241_, new_n882_, new_n1145_, new_n929_, new_n986_, new_n1159_, new_n314_, new_n1584_, new_n1337_, new_n216_, new_n1348_, new_n917_, new_n1555_, new_n1636_, new_n1322_, new_n1133_, new_n1177_, new_n646_, new_n538_, new_n1026_, new_n541_, new_n210_, new_n447_, new_n1388_, new_n1550_, new_n790_, new_n1081_, new_n311_, new_n587_, new_n1247_, new_n1411_, new_n465_, new_n783_, new_n1380_, new_n739_, new_n263_, new_n341_, new_n996_, new_n1601_, new_n1318_, new_n846_, new_n915_, new_n488_, new_n524_, new_n349_, new_n848_, new_n277_, new_n1245_, new_n663_, new_n1499_, new_n1497_, new_n579_, new_n286_, new_n1375_, new_n1254_, new_n438_, new_n1344_, new_n939_, new_n1393_, new_n632_, new_n1335_, new_n1364_, new_n671_, new_n965_, new_n1514_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n1202_, new_n1526_, new_n397_, new_n1446_, new_n975_, new_n1199_, new_n399_, new_n1581_, new_n596_, new_n945_, new_n870_, new_n805_, new_n1403_, new_n1115_, new_n1383_, new_n1231_, new_n948_, new_n1520_, new_n1055_, new_n1431_, new_n838_, new_n1609_, new_n923_, new_n233_, new_n469_, new_n391_, new_n437_, new_n1085_, new_n1633_, new_n1607_, new_n359_, new_n794_, new_n457_, new_n1301_, new_n1128_, new_n1582_, new_n1002_, new_n1169_, new_n448_, new_n384_, new_n900_, new_n1329_, new_n1161_, new_n1648_, new_n924_, new_n775_, new_n454_, new_n1034_, new_n1124_, new_n1000_, new_n308_, new_n633_, new_n784_, new_n1273_, new_n1396_, new_n1491_, new_n1554_, new_n258_, new_n860_, new_n306_, new_n494_, new_n291_, new_n309_, new_n1160_, new_n259_, new_n654_, new_n1456_, new_n713_, new_n880_, new_n1102_, new_n227_, new_n690_, new_n416_, new_n1043_, new_n222_, new_n744_, new_n400_, new_n1175_, new_n1136_, new_n1272_, new_n693_, new_n1287_, new_n1485_, new_n505_, new_n619_, new_n471_, new_n967_, new_n577_, new_n374_, new_n1135_, new_n376_, new_n1538_, new_n1579_, new_n1289_, new_n1561_, new_n1271_, new_n1251_, new_n747_, new_n749_, new_n1091_, new_n1095_, new_n310_, new_n275_, new_n998_, new_n1056_, new_n1331_, new_n1094_, new_n1621_, new_n839_, new_n1030_, new_n485_, new_n578_, new_n525_, new_n918_, new_n1586_, new_n940_, new_n810_, new_n808_, new_n1284_, new_n1572_, new_n907_, new_n665_, new_n800_, new_n897_, new_n1012_, new_n1387_, new_n719_, new_n869_, new_n1178_, new_n1525_, new_n270_, new_n570_, new_n598_, new_n893_, new_n520_, new_n1347_, new_n1001_, new_n253_, new_n825_, new_n1627_, new_n557_, new_n260_, new_n1642_, new_n251_, new_n300_, new_n1503_, new_n507_, new_n741_, new_n806_, new_n605_, new_n1224_, new_n1074_, new_n748_, new_n1137_, new_n1286_, new_n1551_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n1141_, new_n1650_, new_n807_, new_n1326_, new_n592_, new_n726_, new_n1263_, new_n1123_, new_n231_, new_n1080_, new_n583_, new_n617_, new_n1279_, new_n1467_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n916_, new_n428_, new_n487_, new_n675_, new_n1155_, new_n360_, new_n1186_, new_n1261_, new_n225_, new_n1246_, new_n1488_, new_n922_, new_n387_, new_n476_, new_n987_, new_n1641_, new_n949_, new_n221_, new_n450_, new_n1394_, new_n243_, new_n1179_, new_n298_, new_n1088_, new_n1148_, new_n1146_, new_n569_, new_n555_, new_n468_, new_n977_, new_n782_, new_n444_, new_n392_, new_n518_, new_n950_, new_n737_, new_n1022_, new_n340_, new_n285_, new_n692_, new_n502_, new_n209_, new_n623_, new_n446_, new_n316_, new_n203_, new_n590_, new_n826_, new_n789_, new_n1476_, new_n515_, new_n332_, new_n972_, new_n1634_, new_n1067_, new_n891_, new_n516_, new_n1227_, new_n1352_, new_n733_, new_n1021_, new_n1076_, new_n585_, new_n1350_, new_n312_, new_n535_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n1244_, new_n307_, new_n1378_, new_n1478_, new_n1093_, new_n597_, new_n1451_, new_n1092_, new_n1143_, new_n1072_, new_n1190_, new_n1097_, new_n1069_, new_n651_, new_n1164_, new_n1296_, new_n435_, new_n1309_, new_n1010_, new_n776_, new_n687_, new_n1029_, new_n370_, new_n1649_, new_n1654_, new_n638_, new_n523_, new_n909_, new_n1571_, new_n217_, new_n788_, new_n841_, new_n1457_, new_n1204_, new_n1610_, new_n1470_, new_n1112_, new_n711_, new_n1156_, new_n731_, new_n599_, new_n930_, new_n1475_, new_n1604_, new_n1260_, new_n973_, new_n412_, new_n607_, new_n1529_, new_n1541_, new_n645_, new_n1087_, new_n1096_, new_n723_, new_n1599_, new_n756_, new_n823_, new_n1549_, new_n1577_, new_n574_, new_n1500_, new_n928_, new_n1548_, new_n1578_, new_n319_, new_n1008_, new_n338_, new_n1615_, new_n707_, new_n740_, new_n957_, new_n1047_, new_n787_, new_n1134_, new_n336_, new_n1291_, new_n247_, new_n539_, new_n803_, new_n330_, new_n1270_, new_n727_, new_n1531_, new_n294_, new_n1589_, new_n1295_, new_n1173_, new_n704_, new_n1432_, new_n1570_, new_n1189_, new_n1197_, new_n1312_, new_n1502_, new_n474_, new_n1223_, new_n1129_, new_n1013_, new_n467_, new_n404_, new_n1243_, new_n1077_, new_n490_, new_n560_, new_n1100_, new_n865_, new_n358_, new_n877_, new_n1506_, new_n1583_, new_n545_, new_n228_, new_n611_, new_n289_, new_n1011_, new_n425_, new_n896_, new_n802_, new_n1236_, new_n866_, new_n1556_, new_n947_, new_n994_, new_n982_, new_n1449_, new_n964_, new_n1078_, new_n551_, new_n1408_, new_n279_, new_n455_, new_n1569_, new_n618_, new_n1140_, new_n1042_, new_n863_, new_n828_, new_n980_, new_n1605_, new_n464_, new_n1498_, new_n204_, new_n1588_, new_n573_, new_n765_, new_n1314_, new_n1103_;

not g0000 ( new_n202_, keyIn_0_55 );
not g0001 ( new_n203_, keyIn_0_43 );
not g0002 ( new_n204_, keyIn_0_10 );
not g0003 ( new_n205_, N85 );
and g0004 ( new_n206_, new_n205_, N81 );
not g0005 ( new_n207_, N81 );
and g0006 ( new_n208_, new_n207_, N85 );
or g0007 ( new_n209_, new_n206_, new_n208_ );
and g0008 ( new_n210_, new_n209_, new_n204_ );
not g0009 ( new_n211_, new_n210_ );
or g0010 ( new_n212_, new_n209_, new_n204_ );
and g0011 ( new_n213_, new_n211_, new_n212_ );
not g0012 ( new_n214_, new_n213_ );
not g0013 ( new_n215_, N93 );
and g0014 ( new_n216_, new_n215_, N89 );
not g0015 ( new_n217_, N89 );
and g0016 ( new_n218_, new_n217_, N93 );
or g0017 ( new_n219_, new_n216_, new_n218_ );
not g0018 ( new_n220_, new_n219_ );
and g0019 ( new_n221_, new_n220_, keyIn_0_11 );
not g0020 ( new_n222_, new_n221_ );
or g0021 ( new_n223_, new_n220_, keyIn_0_11 );
and g0022 ( new_n224_, new_n222_, new_n223_ );
and g0023 ( new_n225_, new_n214_, new_n224_ );
not g0024 ( new_n226_, new_n225_ );
or g0025 ( new_n227_, new_n214_, new_n224_ );
and g0026 ( new_n228_, new_n226_, new_n227_ );
not g0027 ( new_n229_, new_n228_ );
and g0028 ( new_n230_, new_n229_, keyIn_0_33 );
not g0029 ( new_n231_, new_n230_ );
or g0030 ( new_n232_, new_n229_, keyIn_0_33 );
and g0031 ( new_n233_, new_n231_, new_n232_ );
not g0032 ( new_n234_, new_n233_ );
not g0033 ( new_n235_, keyIn_0_32 );
not g0034 ( new_n236_, N69 );
and g0035 ( new_n237_, new_n236_, N65 );
not g0036 ( new_n238_, N65 );
and g0037 ( new_n239_, new_n238_, N69 );
or g0038 ( new_n240_, new_n237_, new_n239_ );
and g0039 ( new_n241_, new_n240_, keyIn_0_8 );
not g0040 ( new_n242_, new_n241_ );
or g0041 ( new_n243_, new_n240_, keyIn_0_8 );
and g0042 ( new_n244_, new_n242_, new_n243_ );
not g0043 ( new_n245_, new_n244_ );
not g0044 ( new_n246_, keyIn_0_9 );
not g0045 ( new_n247_, N77 );
and g0046 ( new_n248_, new_n247_, N73 );
not g0047 ( new_n249_, N73 );
and g0048 ( new_n250_, new_n249_, N77 );
or g0049 ( new_n251_, new_n248_, new_n250_ );
and g0050 ( new_n252_, new_n251_, new_n246_ );
not g0051 ( new_n253_, new_n252_ );
or g0052 ( new_n254_, new_n251_, new_n246_ );
and g0053 ( new_n255_, new_n253_, new_n254_ );
not g0054 ( new_n256_, new_n255_ );
and g0055 ( new_n257_, new_n245_, new_n256_ );
and g0056 ( new_n258_, new_n244_, new_n255_ );
or g0057 ( new_n259_, new_n257_, new_n258_ );
and g0058 ( new_n260_, new_n259_, new_n235_ );
not g0059 ( new_n261_, new_n260_ );
or g0060 ( new_n262_, new_n259_, new_n235_ );
and g0061 ( new_n263_, new_n261_, new_n262_ );
not g0062 ( new_n264_, new_n263_ );
and g0063 ( new_n265_, new_n234_, new_n264_ );
and g0064 ( new_n266_, new_n233_, new_n263_ );
or g0065 ( new_n267_, new_n265_, new_n266_ );
and g0066 ( new_n268_, new_n267_, new_n203_ );
not g0067 ( new_n269_, new_n268_ );
or g0068 ( new_n270_, new_n267_, new_n203_ );
and g0069 ( new_n271_, new_n269_, new_n270_ );
and g0070 ( new_n272_, N129, N137 );
not g0071 ( new_n273_, new_n272_ );
and g0072 ( new_n274_, new_n271_, new_n273_ );
not g0073 ( new_n275_, new_n274_ );
or g0074 ( new_n276_, new_n271_, new_n273_ );
and g0075 ( new_n277_, new_n275_, new_n276_ );
not g0076 ( new_n278_, new_n277_ );
and g0077 ( new_n279_, new_n278_, keyIn_0_47 );
not g0078 ( new_n280_, new_n279_ );
or g0079 ( new_n281_, new_n278_, keyIn_0_47 );
and g0080 ( new_n282_, new_n280_, new_n281_ );
not g0081 ( new_n283_, N49 );
and g0082 ( new_n284_, new_n283_, N33 );
not g0083 ( new_n285_, N33 );
and g0084 ( new_n286_, new_n285_, N49 );
or g0085 ( new_n287_, new_n284_, new_n286_ );
not g0086 ( new_n288_, new_n287_ );
not g0087 ( new_n289_, N17 );
and g0088 ( new_n290_, new_n289_, N1 );
not g0089 ( new_n291_, N1 );
and g0090 ( new_n292_, new_n291_, N17 );
or g0091 ( new_n293_, new_n290_, new_n292_ );
and g0092 ( new_n294_, new_n288_, new_n293_ );
not g0093 ( new_n295_, new_n294_ );
or g0094 ( new_n296_, new_n288_, new_n293_ );
and g0095 ( new_n297_, new_n295_, new_n296_ );
or g0096 ( new_n298_, new_n282_, new_n297_ );
not g0097 ( new_n299_, new_n298_ );
and g0098 ( new_n300_, new_n282_, new_n297_ );
or g0099 ( new_n301_, new_n299_, new_n300_ );
or g0100 ( new_n302_, new_n301_, new_n202_ );
not g0101 ( new_n303_, new_n300_ );
and g0102 ( new_n304_, new_n303_, new_n298_ );
or g0103 ( new_n305_, new_n304_, keyIn_0_55 );
and g0104 ( new_n306_, new_n302_, new_n305_ );
not g0105 ( new_n307_, new_n306_ );
not g0106 ( new_n308_, keyIn_0_57 );
not g0107 ( new_n309_, keyIn_0_49 );
and g0108 ( new_n310_, N131, N137 );
not g0109 ( new_n311_, N101 );
and g0110 ( new_n312_, new_n311_, N97 );
not g0111 ( new_n313_, N97 );
and g0112 ( new_n314_, new_n313_, N101 );
or g0113 ( new_n315_, new_n312_, new_n314_ );
and g0114 ( new_n316_, new_n315_, keyIn_0_12 );
not g0115 ( new_n317_, new_n316_ );
or g0116 ( new_n318_, new_n315_, keyIn_0_12 );
and g0117 ( new_n319_, new_n317_, new_n318_ );
not g0118 ( new_n320_, new_n319_ );
not g0119 ( new_n321_, keyIn_0_13 );
not g0120 ( new_n322_, N109 );
and g0121 ( new_n323_, new_n322_, N105 );
not g0122 ( new_n324_, N105 );
and g0123 ( new_n325_, new_n324_, N109 );
or g0124 ( new_n326_, new_n323_, new_n325_ );
and g0125 ( new_n327_, new_n326_, new_n321_ );
not g0126 ( new_n328_, new_n327_ );
or g0127 ( new_n329_, new_n326_, new_n321_ );
and g0128 ( new_n330_, new_n328_, new_n329_ );
not g0129 ( new_n331_, new_n330_ );
and g0130 ( new_n332_, new_n320_, new_n331_ );
and g0131 ( new_n333_, new_n319_, new_n330_ );
or g0132 ( new_n334_, new_n332_, new_n333_ );
and g0133 ( new_n335_, new_n334_, keyIn_0_34 );
not g0134 ( new_n336_, new_n335_ );
or g0135 ( new_n337_, new_n334_, keyIn_0_34 );
and g0136 ( new_n338_, new_n336_, new_n337_ );
and g0137 ( new_n339_, new_n264_, new_n338_ );
not g0138 ( new_n340_, new_n338_ );
and g0139 ( new_n341_, new_n340_, new_n263_ );
or g0140 ( new_n342_, new_n339_, new_n341_ );
and g0141 ( new_n343_, new_n342_, keyIn_0_45 );
not g0142 ( new_n344_, new_n343_ );
or g0143 ( new_n345_, new_n342_, keyIn_0_45 );
and g0144 ( new_n346_, new_n344_, new_n345_ );
not g0145 ( new_n347_, new_n346_ );
and g0146 ( new_n348_, new_n347_, keyIn_0_16 );
not g0147 ( new_n349_, new_n348_ );
or g0148 ( new_n350_, new_n347_, keyIn_0_16 );
and g0149 ( new_n351_, new_n349_, new_n350_ );
and g0150 ( new_n352_, new_n351_, new_n310_ );
not g0151 ( new_n353_, new_n352_ );
or g0152 ( new_n354_, new_n351_, new_n310_ );
and g0153 ( new_n355_, new_n353_, new_n354_ );
or g0154 ( new_n356_, new_n355_, new_n309_ );
and g0155 ( new_n357_, new_n355_, new_n309_ );
not g0156 ( new_n358_, new_n357_ );
and g0157 ( new_n359_, new_n358_, new_n356_ );
not g0158 ( new_n360_, N25 );
and g0159 ( new_n361_, new_n360_, N9 );
not g0160 ( new_n362_, N9 );
and g0161 ( new_n363_, new_n362_, N25 );
or g0162 ( new_n364_, new_n361_, new_n363_ );
and g0163 ( new_n365_, new_n364_, keyIn_0_21 );
not g0164 ( new_n366_, new_n365_ );
or g0165 ( new_n367_, new_n364_, keyIn_0_21 );
and g0166 ( new_n368_, new_n366_, new_n367_ );
not g0167 ( new_n369_, new_n368_ );
not g0168 ( new_n370_, N57 );
and g0169 ( new_n371_, new_n370_, N41 );
not g0170 ( new_n372_, N41 );
and g0171 ( new_n373_, new_n372_, N57 );
or g0172 ( new_n374_, new_n371_, new_n373_ );
and g0173 ( new_n375_, new_n374_, keyIn_0_22 );
not g0174 ( new_n376_, new_n375_ );
or g0175 ( new_n377_, new_n374_, keyIn_0_22 );
and g0176 ( new_n378_, new_n376_, new_n377_ );
and g0177 ( new_n379_, new_n369_, new_n378_ );
not g0178 ( new_n380_, new_n379_ );
or g0179 ( new_n381_, new_n369_, new_n378_ );
and g0180 ( new_n382_, new_n380_, new_n381_ );
not g0181 ( new_n383_, new_n382_ );
and g0182 ( new_n384_, new_n383_, keyIn_0_36 );
not g0183 ( new_n385_, new_n384_ );
or g0184 ( new_n386_, new_n383_, keyIn_0_36 );
and g0185 ( new_n387_, new_n385_, new_n386_ );
or g0186 ( new_n388_, new_n359_, new_n387_ );
not g0187 ( new_n389_, new_n356_ );
or g0188 ( new_n390_, new_n389_, new_n357_ );
not g0189 ( new_n391_, new_n387_ );
or g0190 ( new_n392_, new_n390_, new_n391_ );
and g0191 ( new_n393_, new_n392_, new_n388_ );
and g0192 ( new_n394_, new_n393_, new_n308_ );
and g0193 ( new_n395_, new_n390_, new_n391_ );
and g0194 ( new_n396_, new_n359_, new_n387_ );
or g0195 ( new_n397_, new_n395_, new_n396_ );
and g0196 ( new_n398_, new_n397_, keyIn_0_57 );
or g0197 ( new_n399_, new_n398_, new_n394_ );
and g0198 ( new_n400_, new_n399_, keyIn_0_63 );
not g0199 ( new_n401_, new_n400_ );
or g0200 ( new_n402_, new_n399_, keyIn_0_63 );
not g0201 ( new_n403_, keyIn_0_56 );
not g0202 ( new_n404_, keyIn_0_48 );
not g0203 ( new_n405_, keyIn_0_35 );
not g0204 ( new_n406_, keyIn_0_14 );
not g0205 ( new_n407_, N117 );
and g0206 ( new_n408_, new_n407_, N113 );
not g0207 ( new_n409_, N113 );
and g0208 ( new_n410_, new_n409_, N117 );
or g0209 ( new_n411_, new_n408_, new_n410_ );
and g0210 ( new_n412_, new_n411_, new_n406_ );
not g0211 ( new_n413_, new_n412_ );
or g0212 ( new_n414_, new_n411_, new_n406_ );
and g0213 ( new_n415_, new_n413_, new_n414_ );
not g0214 ( new_n416_, new_n415_ );
not g0215 ( new_n417_, keyIn_0_15 );
not g0216 ( new_n418_, N125 );
and g0217 ( new_n419_, new_n418_, N121 );
not g0218 ( new_n420_, N121 );
and g0219 ( new_n421_, new_n420_, N125 );
or g0220 ( new_n422_, new_n419_, new_n421_ );
and g0221 ( new_n423_, new_n422_, new_n417_ );
not g0222 ( new_n424_, new_n423_ );
or g0223 ( new_n425_, new_n422_, new_n417_ );
and g0224 ( new_n426_, new_n424_, new_n425_ );
not g0225 ( new_n427_, new_n426_ );
and g0226 ( new_n428_, new_n416_, new_n427_ );
and g0227 ( new_n429_, new_n415_, new_n426_ );
or g0228 ( new_n430_, new_n428_, new_n429_ );
and g0229 ( new_n431_, new_n430_, new_n405_ );
not g0230 ( new_n432_, new_n431_ );
or g0231 ( new_n433_, new_n430_, new_n405_ );
and g0232 ( new_n434_, new_n432_, new_n433_ );
and g0233 ( new_n435_, new_n340_, new_n434_ );
not g0234 ( new_n436_, new_n434_ );
and g0235 ( new_n437_, new_n436_, new_n338_ );
or g0236 ( new_n438_, new_n435_, new_n437_ );
and g0237 ( new_n439_, new_n438_, keyIn_0_44 );
not g0238 ( new_n440_, new_n439_ );
or g0239 ( new_n441_, new_n438_, keyIn_0_44 );
and g0240 ( new_n442_, new_n440_, new_n441_ );
and g0241 ( new_n443_, N130, N137 );
not g0242 ( new_n444_, new_n443_ );
and g0243 ( new_n445_, new_n442_, new_n444_ );
not g0244 ( new_n446_, new_n445_ );
or g0245 ( new_n447_, new_n442_, new_n444_ );
and g0246 ( new_n448_, new_n446_, new_n447_ );
or g0247 ( new_n449_, new_n448_, new_n404_ );
and g0248 ( new_n450_, new_n448_, new_n404_ );
not g0249 ( new_n451_, new_n450_ );
and g0250 ( new_n452_, new_n451_, new_n449_ );
not g0251 ( new_n453_, N53 );
and g0252 ( new_n454_, new_n453_, N37 );
not g0253 ( new_n455_, N37 );
and g0254 ( new_n456_, new_n455_, N53 );
or g0255 ( new_n457_, new_n454_, new_n456_ );
not g0256 ( new_n458_, new_n457_ );
not g0257 ( new_n459_, N21 );
and g0258 ( new_n460_, new_n459_, N5 );
not g0259 ( new_n461_, N5 );
and g0260 ( new_n462_, new_n461_, N21 );
or g0261 ( new_n463_, new_n460_, new_n462_ );
and g0262 ( new_n464_, new_n458_, new_n463_ );
not g0263 ( new_n465_, new_n464_ );
or g0264 ( new_n466_, new_n458_, new_n463_ );
and g0265 ( new_n467_, new_n465_, new_n466_ );
or g0266 ( new_n468_, new_n452_, new_n467_ );
and g0267 ( new_n469_, new_n452_, new_n467_ );
not g0268 ( new_n470_, new_n469_ );
and g0269 ( new_n471_, new_n470_, new_n468_ );
not g0270 ( new_n472_, new_n471_ );
and g0271 ( new_n473_, new_n472_, new_n403_ );
and g0272 ( new_n474_, new_n471_, keyIn_0_56 );
or g0273 ( new_n475_, new_n473_, new_n474_ );
not g0274 ( new_n476_, new_n475_ );
or g0275 ( new_n477_, new_n306_, new_n476_ );
not g0276 ( new_n478_, keyIn_0_50 );
not g0277 ( new_n479_, keyIn_0_46 );
and g0278 ( new_n480_, new_n234_, new_n436_ );
and g0279 ( new_n481_, new_n233_, new_n434_ );
or g0280 ( new_n482_, new_n480_, new_n481_ );
and g0281 ( new_n483_, new_n482_, new_n479_ );
not g0282 ( new_n484_, new_n483_ );
or g0283 ( new_n485_, new_n482_, new_n479_ );
and g0284 ( new_n486_, new_n484_, new_n485_ );
and g0285 ( new_n487_, N132, N137 );
and g0286 ( new_n488_, new_n486_, new_n487_ );
not g0287 ( new_n489_, new_n488_ );
or g0288 ( new_n490_, new_n486_, new_n487_ );
and g0289 ( new_n491_, new_n489_, new_n490_ );
not g0290 ( new_n492_, new_n491_ );
and g0291 ( new_n493_, new_n492_, new_n478_ );
and g0292 ( new_n494_, new_n491_, keyIn_0_50 );
or g0293 ( new_n495_, new_n493_, new_n494_ );
not g0294 ( new_n496_, new_n495_ );
not g0295 ( new_n497_, keyIn_0_23 );
not g0296 ( new_n498_, N29 );
and g0297 ( new_n499_, new_n498_, N13 );
not g0298 ( new_n500_, N13 );
and g0299 ( new_n501_, new_n500_, N29 );
or g0300 ( new_n502_, new_n499_, new_n501_ );
and g0301 ( new_n503_, new_n502_, new_n497_ );
not g0302 ( new_n504_, new_n503_ );
or g0303 ( new_n505_, new_n502_, new_n497_ );
and g0304 ( new_n506_, new_n504_, new_n505_ );
not g0305 ( new_n507_, new_n506_ );
not g0306 ( new_n508_, N61 );
and g0307 ( new_n509_, new_n508_, N45 );
not g0308 ( new_n510_, N45 );
and g0309 ( new_n511_, new_n510_, N61 );
or g0310 ( new_n512_, new_n509_, new_n511_ );
not g0311 ( new_n513_, new_n512_ );
and g0312 ( new_n514_, new_n507_, new_n513_ );
and g0313 ( new_n515_, new_n506_, new_n512_ );
or g0314 ( new_n516_, new_n514_, new_n515_ );
and g0315 ( new_n517_, new_n496_, new_n516_ );
not g0316 ( new_n518_, new_n517_ );
or g0317 ( new_n519_, new_n496_, new_n516_ );
and g0318 ( new_n520_, new_n518_, new_n519_ );
and g0319 ( new_n521_, new_n520_, keyIn_0_58 );
not g0320 ( new_n522_, keyIn_0_58 );
not g0321 ( new_n523_, new_n520_ );
and g0322 ( new_n524_, new_n523_, new_n522_ );
or g0323 ( new_n525_, new_n524_, new_n521_ );
or g0324 ( new_n526_, new_n477_, new_n525_ );
not g0325 ( new_n527_, new_n526_ );
and g0326 ( new_n528_, new_n527_, new_n402_ );
and g0327 ( new_n529_, new_n528_, new_n401_ );
or g0328 ( new_n530_, new_n397_, keyIn_0_57 );
or g0329 ( new_n531_, new_n393_, new_n308_ );
and g0330 ( new_n532_, new_n530_, new_n531_ );
not g0331 ( new_n533_, new_n521_ );
or g0332 ( new_n534_, new_n520_, keyIn_0_58 );
and g0333 ( new_n535_, new_n533_, new_n534_ );
and g0334 ( new_n536_, new_n535_, new_n475_ );
and g0335 ( new_n537_, new_n532_, new_n536_ );
not g0336 ( new_n538_, new_n537_ );
or g0337 ( new_n539_, new_n532_, new_n536_ );
or g0338 ( new_n540_, new_n535_, new_n475_ );
and g0339 ( new_n541_, new_n540_, new_n306_ );
and g0340 ( new_n542_, new_n539_, new_n541_ );
and g0341 ( new_n543_, new_n542_, new_n538_ );
or g0342 ( new_n544_, new_n529_, new_n543_ );
not g0343 ( new_n545_, keyIn_0_52 );
not g0344 ( new_n546_, keyIn_0_40 );
not g0345 ( new_n547_, keyIn_0_30 );
and g0346 ( new_n548_, new_n455_, N33 );
and g0347 ( new_n549_, new_n285_, N37 );
or g0348 ( new_n550_, new_n548_, new_n549_ );
and g0349 ( new_n551_, new_n550_, keyIn_0_4 );
not g0350 ( new_n552_, keyIn_0_4 );
or g0351 ( new_n553_, new_n285_, N37 );
or g0352 ( new_n554_, new_n455_, N33 );
and g0353 ( new_n555_, new_n553_, new_n554_ );
and g0354 ( new_n556_, new_n555_, new_n552_ );
or g0355 ( new_n557_, new_n551_, new_n556_ );
and g0356 ( new_n558_, new_n510_, N41 );
and g0357 ( new_n559_, new_n372_, N45 );
or g0358 ( new_n560_, new_n558_, new_n559_ );
and g0359 ( new_n561_, new_n560_, keyIn_0_5 );
not g0360 ( new_n562_, keyIn_0_5 );
or g0361 ( new_n563_, new_n372_, N45 );
or g0362 ( new_n564_, new_n510_, N41 );
and g0363 ( new_n565_, new_n563_, new_n564_ );
and g0364 ( new_n566_, new_n565_, new_n562_ );
or g0365 ( new_n567_, new_n561_, new_n566_ );
and g0366 ( new_n568_, new_n557_, new_n567_ );
or g0367 ( new_n569_, new_n555_, new_n552_ );
or g0368 ( new_n570_, new_n550_, keyIn_0_4 );
and g0369 ( new_n571_, new_n570_, new_n569_ );
or g0370 ( new_n572_, new_n565_, new_n562_ );
or g0371 ( new_n573_, new_n560_, keyIn_0_5 );
and g0372 ( new_n574_, new_n573_, new_n572_ );
and g0373 ( new_n575_, new_n571_, new_n574_ );
or g0374 ( new_n576_, new_n568_, new_n575_ );
and g0375 ( new_n577_, new_n576_, new_n547_ );
or g0376 ( new_n578_, new_n571_, new_n574_ );
or g0377 ( new_n579_, new_n557_, new_n567_ );
and g0378 ( new_n580_, new_n579_, new_n578_ );
and g0379 ( new_n581_, new_n580_, keyIn_0_30 );
or g0380 ( new_n582_, new_n577_, new_n581_ );
not g0381 ( new_n583_, keyIn_0_31 );
not g0382 ( new_n584_, keyIn_0_6 );
and g0383 ( new_n585_, new_n453_, N49 );
and g0384 ( new_n586_, new_n283_, N53 );
or g0385 ( new_n587_, new_n585_, new_n586_ );
and g0386 ( new_n588_, new_n587_, new_n584_ );
or g0387 ( new_n589_, new_n283_, N53 );
or g0388 ( new_n590_, new_n453_, N49 );
and g0389 ( new_n591_, new_n589_, new_n590_ );
and g0390 ( new_n592_, new_n591_, keyIn_0_6 );
or g0391 ( new_n593_, new_n588_, new_n592_ );
and g0392 ( new_n594_, new_n508_, N57 );
and g0393 ( new_n595_, new_n370_, N61 );
or g0394 ( new_n596_, new_n594_, new_n595_ );
and g0395 ( new_n597_, new_n596_, keyIn_0_7 );
not g0396 ( new_n598_, keyIn_0_7 );
or g0397 ( new_n599_, new_n370_, N61 );
or g0398 ( new_n600_, new_n508_, N57 );
and g0399 ( new_n601_, new_n599_, new_n600_ );
and g0400 ( new_n602_, new_n601_, new_n598_ );
or g0401 ( new_n603_, new_n597_, new_n602_ );
and g0402 ( new_n604_, new_n593_, new_n603_ );
or g0403 ( new_n605_, new_n591_, keyIn_0_6 );
or g0404 ( new_n606_, new_n587_, new_n584_ );
and g0405 ( new_n607_, new_n606_, new_n605_ );
or g0406 ( new_n608_, new_n601_, new_n598_ );
or g0407 ( new_n609_, new_n596_, keyIn_0_7 );
and g0408 ( new_n610_, new_n609_, new_n608_ );
and g0409 ( new_n611_, new_n607_, new_n610_ );
or g0410 ( new_n612_, new_n604_, new_n611_ );
and g0411 ( new_n613_, new_n612_, new_n583_ );
or g0412 ( new_n614_, new_n607_, new_n610_ );
or g0413 ( new_n615_, new_n593_, new_n603_ );
and g0414 ( new_n616_, new_n615_, new_n614_ );
and g0415 ( new_n617_, new_n616_, keyIn_0_31 );
or g0416 ( new_n618_, new_n613_, new_n617_ );
or g0417 ( new_n619_, new_n582_, new_n618_ );
or g0418 ( new_n620_, new_n580_, keyIn_0_30 );
or g0419 ( new_n621_, new_n576_, new_n547_ );
and g0420 ( new_n622_, new_n620_, new_n621_ );
or g0421 ( new_n623_, new_n616_, keyIn_0_31 );
or g0422 ( new_n624_, new_n612_, new_n583_ );
and g0423 ( new_n625_, new_n623_, new_n624_ );
or g0424 ( new_n626_, new_n622_, new_n625_ );
and g0425 ( new_n627_, new_n619_, new_n626_ );
and g0426 ( new_n628_, new_n627_, new_n546_ );
and g0427 ( new_n629_, new_n622_, new_n625_ );
and g0428 ( new_n630_, new_n582_, new_n618_ );
or g0429 ( new_n631_, new_n630_, new_n629_ );
and g0430 ( new_n632_, new_n631_, keyIn_0_40 );
or g0431 ( new_n633_, new_n628_, new_n632_ );
not g0432 ( new_n634_, keyIn_0_18 );
and g0433 ( new_n635_, N134, N137 );
or g0434 ( new_n636_, new_n635_, new_n634_ );
and g0435 ( new_n637_, new_n635_, new_n634_ );
not g0436 ( new_n638_, new_n637_ );
and g0437 ( new_n639_, new_n638_, new_n636_ );
not g0438 ( new_n640_, new_n639_ );
or g0439 ( new_n641_, new_n633_, new_n640_ );
or g0440 ( new_n642_, new_n631_, keyIn_0_40 );
or g0441 ( new_n643_, new_n627_, new_n546_ );
and g0442 ( new_n644_, new_n643_, new_n642_ );
or g0443 ( new_n645_, new_n644_, new_n639_ );
and g0444 ( new_n646_, new_n641_, new_n645_ );
and g0445 ( new_n647_, new_n646_, new_n545_ );
and g0446 ( new_n648_, new_n644_, new_n639_ );
and g0447 ( new_n649_, new_n633_, new_n640_ );
or g0448 ( new_n650_, new_n649_, new_n648_ );
and g0449 ( new_n651_, new_n650_, keyIn_0_52 );
or g0450 ( new_n652_, new_n651_, new_n647_ );
not g0451 ( new_n653_, keyIn_0_37 );
and g0452 ( new_n654_, new_n205_, N69 );
and g0453 ( new_n655_, new_n236_, N85 );
or g0454 ( new_n656_, new_n654_, new_n655_ );
and g0455 ( new_n657_, new_n656_, keyIn_0_24 );
not g0456 ( new_n658_, new_n657_ );
or g0457 ( new_n659_, new_n656_, keyIn_0_24 );
and g0458 ( new_n660_, new_n658_, new_n659_ );
not g0459 ( new_n661_, new_n660_ );
and g0460 ( new_n662_, new_n407_, N101 );
and g0461 ( new_n663_, new_n311_, N117 );
or g0462 ( new_n664_, new_n662_, new_n663_ );
and g0463 ( new_n665_, new_n664_, keyIn_0_25 );
not g0464 ( new_n666_, new_n665_ );
or g0465 ( new_n667_, new_n664_, keyIn_0_25 );
and g0466 ( new_n668_, new_n666_, new_n667_ );
not g0467 ( new_n669_, new_n668_ );
and g0468 ( new_n670_, new_n661_, new_n669_ );
and g0469 ( new_n671_, new_n660_, new_n668_ );
or g0470 ( new_n672_, new_n670_, new_n671_ );
and g0471 ( new_n673_, new_n672_, new_n653_ );
not g0472 ( new_n674_, new_n673_ );
or g0473 ( new_n675_, new_n672_, new_n653_ );
and g0474 ( new_n676_, new_n674_, new_n675_ );
and g0475 ( new_n677_, new_n652_, new_n676_ );
or g0476 ( new_n678_, new_n650_, keyIn_0_52 );
or g0477 ( new_n679_, new_n646_, new_n545_ );
and g0478 ( new_n680_, new_n678_, new_n679_ );
not g0479 ( new_n681_, new_n676_ );
and g0480 ( new_n682_, new_n680_, new_n681_ );
or g0481 ( new_n683_, new_n677_, new_n682_ );
and g0482 ( new_n684_, new_n683_, keyIn_0_60 );
not g0483 ( new_n685_, keyIn_0_60 );
or g0484 ( new_n686_, new_n680_, new_n681_ );
or g0485 ( new_n687_, new_n652_, new_n676_ );
and g0486 ( new_n688_, new_n687_, new_n686_ );
and g0487 ( new_n689_, new_n688_, new_n685_ );
or g0488 ( new_n690_, new_n684_, new_n689_ );
not g0489 ( new_n691_, keyIn_0_2 );
and g0490 ( new_n692_, new_n459_, N17 );
and g0491 ( new_n693_, new_n289_, N21 );
or g0492 ( new_n694_, new_n692_, new_n693_ );
and g0493 ( new_n695_, new_n694_, new_n691_ );
or g0494 ( new_n696_, new_n289_, N21 );
or g0495 ( new_n697_, new_n459_, N17 );
and g0496 ( new_n698_, new_n696_, new_n697_ );
and g0497 ( new_n699_, new_n698_, keyIn_0_2 );
or g0498 ( new_n700_, new_n695_, new_n699_ );
and g0499 ( new_n701_, new_n498_, N25 );
and g0500 ( new_n702_, new_n360_, N29 );
or g0501 ( new_n703_, new_n701_, new_n702_ );
or g0502 ( new_n704_, new_n703_, keyIn_0_3 );
not g0503 ( new_n705_, keyIn_0_3 );
or g0504 ( new_n706_, new_n360_, N29 );
or g0505 ( new_n707_, new_n498_, N25 );
and g0506 ( new_n708_, new_n706_, new_n707_ );
or g0507 ( new_n709_, new_n708_, new_n705_ );
and g0508 ( new_n710_, new_n704_, new_n709_ );
and g0509 ( new_n711_, new_n700_, new_n710_ );
or g0510 ( new_n712_, new_n698_, keyIn_0_2 );
or g0511 ( new_n713_, new_n694_, new_n691_ );
and g0512 ( new_n714_, new_n713_, new_n712_ );
and g0513 ( new_n715_, new_n708_, new_n705_ );
and g0514 ( new_n716_, new_n703_, keyIn_0_3 );
or g0515 ( new_n717_, new_n716_, new_n715_ );
and g0516 ( new_n718_, new_n717_, new_n714_ );
or g0517 ( new_n719_, new_n711_, new_n718_ );
and g0518 ( new_n720_, new_n719_, keyIn_0_29 );
not g0519 ( new_n721_, keyIn_0_29 );
or g0520 ( new_n722_, new_n717_, new_n714_ );
or g0521 ( new_n723_, new_n700_, new_n710_ );
and g0522 ( new_n724_, new_n722_, new_n723_ );
and g0523 ( new_n725_, new_n724_, new_n721_ );
or g0524 ( new_n726_, new_n720_, new_n725_ );
and g0525 ( new_n727_, new_n726_, new_n625_ );
or g0526 ( new_n728_, new_n724_, new_n721_ );
or g0527 ( new_n729_, new_n719_, keyIn_0_29 );
and g0528 ( new_n730_, new_n728_, new_n729_ );
and g0529 ( new_n731_, new_n618_, new_n730_ );
or g0530 ( new_n732_, new_n727_, new_n731_ );
and g0531 ( new_n733_, new_n732_, keyIn_0_42 );
not g0532 ( new_n734_, keyIn_0_42 );
or g0533 ( new_n735_, new_n618_, new_n730_ );
or g0534 ( new_n736_, new_n726_, new_n625_ );
and g0535 ( new_n737_, new_n735_, new_n736_ );
and g0536 ( new_n738_, new_n737_, new_n734_ );
or g0537 ( new_n739_, new_n733_, new_n738_ );
not g0538 ( new_n740_, keyIn_0_20 );
and g0539 ( new_n741_, N136, N137 );
or g0540 ( new_n742_, new_n741_, new_n740_ );
and g0541 ( new_n743_, new_n741_, new_n740_ );
not g0542 ( new_n744_, new_n743_ );
and g0543 ( new_n745_, new_n744_, new_n742_ );
not g0544 ( new_n746_, new_n745_ );
or g0545 ( new_n747_, new_n739_, new_n746_ );
or g0546 ( new_n748_, new_n737_, new_n734_ );
or g0547 ( new_n749_, new_n732_, keyIn_0_42 );
and g0548 ( new_n750_, new_n749_, new_n748_ );
or g0549 ( new_n751_, new_n750_, new_n745_ );
and g0550 ( new_n752_, new_n747_, new_n751_ );
and g0551 ( new_n753_, new_n752_, keyIn_0_54 );
not g0552 ( new_n754_, keyIn_0_54 );
and g0553 ( new_n755_, new_n750_, new_n745_ );
and g0554 ( new_n756_, new_n739_, new_n746_ );
or g0555 ( new_n757_, new_n756_, new_n755_ );
and g0556 ( new_n758_, new_n757_, new_n754_ );
or g0557 ( new_n759_, new_n758_, new_n753_ );
and g0558 ( new_n760_, new_n418_, N109 );
and g0559 ( new_n761_, new_n322_, N125 );
or g0560 ( new_n762_, new_n760_, new_n761_ );
not g0561 ( new_n763_, new_n762_ );
and g0562 ( new_n764_, new_n215_, N77 );
and g0563 ( new_n765_, new_n247_, N93 );
or g0564 ( new_n766_, new_n764_, new_n765_ );
and g0565 ( new_n767_, new_n763_, new_n766_ );
not g0566 ( new_n768_, new_n767_ );
or g0567 ( new_n769_, new_n763_, new_n766_ );
and g0568 ( new_n770_, new_n768_, new_n769_ );
not g0569 ( new_n771_, new_n770_ );
and g0570 ( new_n772_, new_n759_, new_n771_ );
or g0571 ( new_n773_, new_n757_, new_n754_ );
or g0572 ( new_n774_, new_n752_, keyIn_0_54 );
and g0573 ( new_n775_, new_n773_, new_n774_ );
and g0574 ( new_n776_, new_n775_, new_n770_ );
or g0575 ( new_n777_, new_n772_, new_n776_ );
or g0576 ( new_n778_, new_n777_, keyIn_0_62 );
not g0577 ( new_n779_, keyIn_0_62 );
or g0578 ( new_n780_, new_n775_, new_n770_ );
or g0579 ( new_n781_, new_n759_, new_n771_ );
and g0580 ( new_n782_, new_n781_, new_n780_ );
or g0581 ( new_n783_, new_n782_, new_n779_ );
and g0582 ( new_n784_, new_n778_, new_n783_ );
and g0583 ( new_n785_, new_n690_, new_n784_ );
not g0584 ( new_n786_, keyIn_0_53 );
and g0585 ( new_n787_, new_n461_, N1 );
and g0586 ( new_n788_, new_n291_, N5 );
or g0587 ( new_n789_, new_n787_, new_n788_ );
and g0588 ( new_n790_, new_n789_, keyIn_0_0 );
not g0589 ( new_n791_, keyIn_0_0 );
or g0590 ( new_n792_, new_n291_, N5 );
or g0591 ( new_n793_, new_n461_, N1 );
and g0592 ( new_n794_, new_n792_, new_n793_ );
and g0593 ( new_n795_, new_n794_, new_n791_ );
or g0594 ( new_n796_, new_n790_, new_n795_ );
and g0595 ( new_n797_, new_n500_, N9 );
and g0596 ( new_n798_, new_n362_, N13 );
or g0597 ( new_n799_, new_n797_, new_n798_ );
or g0598 ( new_n800_, new_n799_, keyIn_0_1 );
not g0599 ( new_n801_, keyIn_0_1 );
or g0600 ( new_n802_, new_n362_, N13 );
or g0601 ( new_n803_, new_n500_, N9 );
and g0602 ( new_n804_, new_n802_, new_n803_ );
or g0603 ( new_n805_, new_n804_, new_n801_ );
and g0604 ( new_n806_, new_n800_, new_n805_ );
and g0605 ( new_n807_, new_n796_, new_n806_ );
or g0606 ( new_n808_, new_n794_, new_n791_ );
or g0607 ( new_n809_, new_n789_, keyIn_0_0 );
and g0608 ( new_n810_, new_n809_, new_n808_ );
and g0609 ( new_n811_, new_n804_, new_n801_ );
and g0610 ( new_n812_, new_n799_, keyIn_0_1 );
or g0611 ( new_n813_, new_n812_, new_n811_ );
and g0612 ( new_n814_, new_n813_, new_n810_ );
or g0613 ( new_n815_, new_n807_, new_n814_ );
and g0614 ( new_n816_, new_n815_, keyIn_0_28 );
not g0615 ( new_n817_, keyIn_0_28 );
or g0616 ( new_n818_, new_n813_, new_n810_ );
or g0617 ( new_n819_, new_n796_, new_n806_ );
and g0618 ( new_n820_, new_n818_, new_n819_ );
and g0619 ( new_n821_, new_n820_, new_n817_ );
or g0620 ( new_n822_, new_n816_, new_n821_ );
and g0621 ( new_n823_, new_n822_, new_n622_ );
or g0622 ( new_n824_, new_n820_, new_n817_ );
or g0623 ( new_n825_, new_n815_, keyIn_0_28 );
and g0624 ( new_n826_, new_n824_, new_n825_ );
and g0625 ( new_n827_, new_n582_, new_n826_ );
or g0626 ( new_n828_, new_n823_, new_n827_ );
and g0627 ( new_n829_, new_n828_, keyIn_0_41 );
not g0628 ( new_n830_, keyIn_0_41 );
or g0629 ( new_n831_, new_n582_, new_n826_ );
or g0630 ( new_n832_, new_n822_, new_n622_ );
and g0631 ( new_n833_, new_n831_, new_n832_ );
and g0632 ( new_n834_, new_n833_, new_n830_ );
or g0633 ( new_n835_, new_n829_, new_n834_ );
not g0634 ( new_n836_, keyIn_0_19 );
and g0635 ( new_n837_, N135, N137 );
or g0636 ( new_n838_, new_n837_, new_n836_ );
and g0637 ( new_n839_, new_n837_, new_n836_ );
not g0638 ( new_n840_, new_n839_ );
and g0639 ( new_n841_, new_n840_, new_n838_ );
not g0640 ( new_n842_, new_n841_ );
or g0641 ( new_n843_, new_n835_, new_n842_ );
or g0642 ( new_n844_, new_n833_, new_n830_ );
or g0643 ( new_n845_, new_n828_, keyIn_0_41 );
and g0644 ( new_n846_, new_n845_, new_n844_ );
or g0645 ( new_n847_, new_n846_, new_n841_ );
and g0646 ( new_n848_, new_n843_, new_n847_ );
and g0647 ( new_n849_, new_n848_, new_n786_ );
and g0648 ( new_n850_, new_n846_, new_n841_ );
and g0649 ( new_n851_, new_n835_, new_n842_ );
or g0650 ( new_n852_, new_n851_, new_n850_ );
and g0651 ( new_n853_, new_n852_, keyIn_0_53 );
or g0652 ( new_n854_, new_n853_, new_n849_ );
not g0653 ( new_n855_, keyIn_0_26 );
and g0654 ( new_n856_, new_n217_, N73 );
and g0655 ( new_n857_, new_n249_, N89 );
or g0656 ( new_n858_, new_n856_, new_n857_ );
and g0657 ( new_n859_, new_n858_, new_n855_ );
not g0658 ( new_n860_, new_n859_ );
or g0659 ( new_n861_, new_n858_, new_n855_ );
and g0660 ( new_n862_, new_n860_, new_n861_ );
not g0661 ( new_n863_, new_n862_ );
not g0662 ( new_n864_, keyIn_0_27 );
and g0663 ( new_n865_, new_n420_, N105 );
and g0664 ( new_n866_, new_n324_, N121 );
or g0665 ( new_n867_, new_n865_, new_n866_ );
and g0666 ( new_n868_, new_n867_, new_n864_ );
not g0667 ( new_n869_, new_n868_ );
or g0668 ( new_n870_, new_n867_, new_n864_ );
and g0669 ( new_n871_, new_n869_, new_n870_ );
not g0670 ( new_n872_, new_n871_ );
and g0671 ( new_n873_, new_n863_, new_n872_ );
and g0672 ( new_n874_, new_n862_, new_n871_ );
or g0673 ( new_n875_, new_n873_, new_n874_ );
and g0674 ( new_n876_, new_n875_, keyIn_0_38 );
not g0675 ( new_n877_, new_n876_ );
or g0676 ( new_n878_, new_n875_, keyIn_0_38 );
and g0677 ( new_n879_, new_n877_, new_n878_ );
not g0678 ( new_n880_, new_n879_ );
and g0679 ( new_n881_, new_n854_, new_n880_ );
or g0680 ( new_n882_, new_n852_, keyIn_0_53 );
or g0681 ( new_n883_, new_n848_, new_n786_ );
and g0682 ( new_n884_, new_n882_, new_n883_ );
and g0683 ( new_n885_, new_n884_, new_n879_ );
or g0684 ( new_n886_, new_n881_, new_n885_ );
or g0685 ( new_n887_, new_n886_, keyIn_0_61 );
not g0686 ( new_n888_, keyIn_0_61 );
or g0687 ( new_n889_, new_n884_, new_n879_ );
or g0688 ( new_n890_, new_n854_, new_n880_ );
and g0689 ( new_n891_, new_n890_, new_n889_ );
or g0690 ( new_n892_, new_n891_, new_n888_ );
and g0691 ( new_n893_, new_n887_, new_n892_ );
and g0692 ( new_n894_, new_n785_, new_n893_ );
not g0693 ( new_n895_, keyIn_0_59 );
not g0694 ( new_n896_, keyIn_0_51 );
not g0695 ( new_n897_, keyIn_0_39 );
and g0696 ( new_n898_, new_n730_, new_n826_ );
and g0697 ( new_n899_, new_n726_, new_n822_ );
or g0698 ( new_n900_, new_n899_, new_n898_ );
or g0699 ( new_n901_, new_n900_, new_n897_ );
or g0700 ( new_n902_, new_n726_, new_n822_ );
or g0701 ( new_n903_, new_n730_, new_n826_ );
and g0702 ( new_n904_, new_n902_, new_n903_ );
or g0703 ( new_n905_, new_n904_, keyIn_0_39 );
and g0704 ( new_n906_, new_n905_, new_n901_ );
not g0705 ( new_n907_, keyIn_0_17 );
and g0706 ( new_n908_, N133, N137 );
or g0707 ( new_n909_, new_n908_, new_n907_ );
and g0708 ( new_n910_, new_n908_, new_n907_ );
not g0709 ( new_n911_, new_n910_ );
and g0710 ( new_n912_, new_n911_, new_n909_ );
and g0711 ( new_n913_, new_n906_, new_n912_ );
and g0712 ( new_n914_, new_n904_, keyIn_0_39 );
and g0713 ( new_n915_, new_n900_, new_n897_ );
or g0714 ( new_n916_, new_n914_, new_n915_ );
not g0715 ( new_n917_, new_n912_ );
and g0716 ( new_n918_, new_n916_, new_n917_ );
or g0717 ( new_n919_, new_n918_, new_n913_ );
and g0718 ( new_n920_, new_n919_, new_n896_ );
or g0719 ( new_n921_, new_n916_, new_n917_ );
or g0720 ( new_n922_, new_n906_, new_n912_ );
and g0721 ( new_n923_, new_n921_, new_n922_ );
and g0722 ( new_n924_, new_n923_, keyIn_0_51 );
or g0723 ( new_n925_, new_n920_, new_n924_ );
and g0724 ( new_n926_, new_n409_, N97 );
and g0725 ( new_n927_, new_n313_, N113 );
or g0726 ( new_n928_, new_n926_, new_n927_ );
not g0727 ( new_n929_, new_n928_ );
and g0728 ( new_n930_, new_n207_, N65 );
and g0729 ( new_n931_, new_n238_, N81 );
or g0730 ( new_n932_, new_n930_, new_n931_ );
and g0731 ( new_n933_, new_n929_, new_n932_ );
not g0732 ( new_n934_, new_n933_ );
or g0733 ( new_n935_, new_n929_, new_n932_ );
and g0734 ( new_n936_, new_n934_, new_n935_ );
not g0735 ( new_n937_, new_n936_ );
and g0736 ( new_n938_, new_n925_, new_n937_ );
or g0737 ( new_n939_, new_n923_, keyIn_0_51 );
or g0738 ( new_n940_, new_n919_, new_n896_ );
and g0739 ( new_n941_, new_n940_, new_n939_ );
and g0740 ( new_n942_, new_n941_, new_n936_ );
or g0741 ( new_n943_, new_n938_, new_n942_ );
or g0742 ( new_n944_, new_n943_, new_n895_ );
or g0743 ( new_n945_, new_n941_, new_n936_ );
or g0744 ( new_n946_, new_n925_, new_n937_ );
and g0745 ( new_n947_, new_n946_, new_n945_ );
or g0746 ( new_n948_, new_n947_, keyIn_0_59 );
and g0747 ( new_n949_, new_n944_, new_n948_ );
and g0748 ( new_n950_, new_n894_, new_n949_ );
and g0749 ( new_n951_, new_n544_, new_n950_ );
and g0750 ( new_n952_, new_n951_, new_n307_ );
not g0751 ( new_n953_, new_n952_ );
and g0752 ( new_n954_, new_n953_, N1 );
and g0753 ( new_n955_, new_n952_, new_n291_ );
or g0754 ( N724, new_n954_, new_n955_ );
and g0755 ( new_n957_, new_n951_, new_n476_ );
not g0756 ( new_n958_, new_n957_ );
and g0757 ( new_n959_, new_n958_, N5 );
and g0758 ( new_n960_, new_n957_, new_n461_ );
or g0759 ( N725, new_n959_, new_n960_ );
and g0760 ( new_n962_, new_n951_, new_n399_ );
not g0761 ( new_n963_, new_n962_ );
and g0762 ( new_n964_, new_n963_, N9 );
and g0763 ( new_n965_, new_n962_, new_n362_ );
or g0764 ( N726, new_n964_, new_n965_ );
and g0765 ( new_n967_, new_n951_, new_n525_ );
not g0766 ( new_n968_, new_n967_ );
and g0767 ( new_n969_, new_n968_, N13 );
and g0768 ( new_n970_, new_n967_, new_n500_ );
or g0769 ( N727, new_n969_, new_n970_ );
not g0770 ( new_n972_, keyIn_0_63 );
and g0771 ( new_n973_, new_n532_, new_n972_ );
or g0772 ( new_n974_, new_n973_, new_n526_ );
or g0773 ( new_n975_, new_n974_, new_n400_ );
or g0774 ( new_n976_, new_n525_, new_n476_ );
and g0775 ( new_n977_, new_n399_, new_n976_ );
and g0776 ( new_n978_, new_n525_, new_n476_ );
or g0777 ( new_n979_, new_n978_, new_n307_ );
or g0778 ( new_n980_, new_n977_, new_n979_ );
or g0779 ( new_n981_, new_n980_, new_n537_ );
and g0780 ( new_n982_, new_n981_, new_n975_ );
and g0781 ( new_n983_, new_n782_, new_n779_ );
and g0782 ( new_n984_, new_n777_, keyIn_0_62 );
or g0783 ( new_n985_, new_n984_, new_n983_ );
and g0784 ( new_n986_, new_n891_, new_n888_ );
and g0785 ( new_n987_, new_n886_, keyIn_0_61 );
or g0786 ( new_n988_, new_n987_, new_n986_ );
and g0787 ( new_n989_, new_n985_, new_n988_ );
and g0788 ( new_n990_, new_n690_, new_n949_ );
and g0789 ( new_n991_, new_n989_, new_n990_ );
not g0790 ( new_n992_, new_n991_ );
or g0791 ( new_n993_, new_n982_, new_n992_ );
and g0792 ( new_n994_, new_n993_, keyIn_0_76 );
not g0793 ( new_n995_, keyIn_0_76 );
and g0794 ( new_n996_, new_n544_, new_n991_ );
and g0795 ( new_n997_, new_n996_, new_n995_ );
or g0796 ( new_n998_, new_n994_, new_n997_ );
or g0797 ( new_n999_, new_n998_, new_n306_ );
and g0798 ( new_n1000_, new_n999_, keyIn_0_82 );
not g0799 ( new_n1001_, keyIn_0_82 );
or g0800 ( new_n1002_, new_n996_, new_n995_ );
or g0801 ( new_n1003_, new_n993_, keyIn_0_76 );
and g0802 ( new_n1004_, new_n1003_, new_n1002_ );
and g0803 ( new_n1005_, new_n1004_, new_n307_ );
and g0804 ( new_n1006_, new_n1005_, new_n1001_ );
or g0805 ( new_n1007_, new_n1000_, new_n1006_ );
and g0806 ( new_n1008_, new_n1007_, new_n289_ );
or g0807 ( new_n1009_, new_n1005_, new_n1001_ );
or g0808 ( new_n1010_, new_n999_, keyIn_0_82 );
and g0809 ( new_n1011_, new_n1010_, new_n1009_ );
and g0810 ( new_n1012_, new_n1011_, N17 );
or g0811 ( new_n1013_, new_n1008_, new_n1012_ );
or g0812 ( new_n1014_, new_n1013_, keyIn_0_105 );
not g0813 ( new_n1015_, keyIn_0_105 );
or g0814 ( new_n1016_, new_n1011_, N17 );
or g0815 ( new_n1017_, new_n1007_, new_n289_ );
and g0816 ( new_n1018_, new_n1017_, new_n1016_ );
or g0817 ( new_n1019_, new_n1018_, new_n1015_ );
and g0818 ( N728, new_n1014_, new_n1019_ );
not g0819 ( new_n1021_, keyIn_0_106 );
not g0820 ( new_n1022_, keyIn_0_83 );
or g0821 ( new_n1023_, new_n998_, new_n475_ );
and g0822 ( new_n1024_, new_n1023_, new_n1022_ );
and g0823 ( new_n1025_, new_n1004_, new_n476_ );
and g0824 ( new_n1026_, new_n1025_, keyIn_0_83 );
or g0825 ( new_n1027_, new_n1024_, new_n1026_ );
and g0826 ( new_n1028_, new_n1027_, N21 );
or g0827 ( new_n1029_, new_n1025_, keyIn_0_83 );
or g0828 ( new_n1030_, new_n1023_, new_n1022_ );
and g0829 ( new_n1031_, new_n1030_, new_n1029_ );
and g0830 ( new_n1032_, new_n1031_, new_n459_ );
or g0831 ( new_n1033_, new_n1028_, new_n1032_ );
or g0832 ( new_n1034_, new_n1033_, new_n1021_ );
or g0833 ( new_n1035_, new_n1031_, new_n459_ );
or g0834 ( new_n1036_, new_n1027_, N21 );
and g0835 ( new_n1037_, new_n1036_, new_n1035_ );
or g0836 ( new_n1038_, new_n1037_, keyIn_0_106 );
and g0837 ( N729, new_n1034_, new_n1038_ );
and g0838 ( new_n1040_, new_n1004_, new_n399_ );
not g0839 ( new_n1041_, new_n1040_ );
and g0840 ( new_n1042_, new_n1041_, N25 );
and g0841 ( new_n1043_, new_n1040_, new_n360_ );
or g0842 ( N730, new_n1042_, new_n1043_ );
not g0843 ( new_n1045_, keyIn_0_107 );
not g0844 ( new_n1046_, keyIn_0_84 );
or g0845 ( new_n1047_, new_n998_, new_n535_ );
and g0846 ( new_n1048_, new_n1047_, new_n1046_ );
and g0847 ( new_n1049_, new_n1004_, new_n525_ );
and g0848 ( new_n1050_, new_n1049_, keyIn_0_84 );
or g0849 ( new_n1051_, new_n1048_, new_n1050_ );
and g0850 ( new_n1052_, new_n1051_, new_n498_ );
or g0851 ( new_n1053_, new_n1049_, keyIn_0_84 );
or g0852 ( new_n1054_, new_n1047_, new_n1046_ );
and g0853 ( new_n1055_, new_n1054_, new_n1053_ );
and g0854 ( new_n1056_, new_n1055_, N29 );
or g0855 ( new_n1057_, new_n1052_, new_n1056_ );
or g0856 ( new_n1058_, new_n1057_, new_n1045_ );
or g0857 ( new_n1059_, new_n1055_, N29 );
or g0858 ( new_n1060_, new_n1051_, new_n498_ );
and g0859 ( new_n1061_, new_n1060_, new_n1059_ );
or g0860 ( new_n1062_, new_n1061_, keyIn_0_107 );
and g0861 ( N731, new_n1058_, new_n1062_ );
not g0862 ( new_n1064_, keyIn_0_85 );
or g0863 ( new_n1065_, new_n688_, new_n685_ );
or g0864 ( new_n1066_, new_n683_, keyIn_0_60 );
and g0865 ( new_n1067_, new_n1066_, new_n1065_ );
and g0866 ( new_n1068_, new_n947_, keyIn_0_59 );
and g0867 ( new_n1069_, new_n943_, new_n895_ );
or g0868 ( new_n1070_, new_n1069_, new_n1068_ );
and g0869 ( new_n1071_, new_n784_, new_n893_ );
and g0870 ( new_n1072_, new_n1071_, new_n1070_ );
and g0871 ( new_n1073_, new_n1072_, new_n1067_ );
not g0872 ( new_n1074_, new_n1073_ );
or g0873 ( new_n1075_, new_n982_, new_n1074_ );
and g0874 ( new_n1076_, new_n1075_, keyIn_0_77 );
not g0875 ( new_n1077_, keyIn_0_77 );
and g0876 ( new_n1078_, new_n544_, new_n1073_ );
and g0877 ( new_n1079_, new_n1078_, new_n1077_ );
or g0878 ( new_n1080_, new_n1076_, new_n1079_ );
or g0879 ( new_n1081_, new_n1080_, new_n306_ );
and g0880 ( new_n1082_, new_n1081_, new_n1064_ );
or g0881 ( new_n1083_, new_n1078_, new_n1077_ );
or g0882 ( new_n1084_, new_n1075_, keyIn_0_77 );
and g0883 ( new_n1085_, new_n1084_, new_n1083_ );
and g0884 ( new_n1086_, new_n1085_, new_n307_ );
and g0885 ( new_n1087_, new_n1086_, keyIn_0_85 );
or g0886 ( new_n1088_, new_n1082_, new_n1087_ );
and g0887 ( new_n1089_, new_n1088_, N33 );
or g0888 ( new_n1090_, new_n1086_, keyIn_0_85 );
or g0889 ( new_n1091_, new_n1081_, new_n1064_ );
and g0890 ( new_n1092_, new_n1091_, new_n1090_ );
and g0891 ( new_n1093_, new_n1092_, new_n285_ );
or g0892 ( new_n1094_, new_n1089_, new_n1093_ );
or g0893 ( new_n1095_, new_n1094_, keyIn_0_108 );
not g0894 ( new_n1096_, keyIn_0_108 );
or g0895 ( new_n1097_, new_n1092_, new_n285_ );
or g0896 ( new_n1098_, new_n1088_, N33 );
and g0897 ( new_n1099_, new_n1098_, new_n1097_ );
or g0898 ( new_n1100_, new_n1099_, new_n1096_ );
and g0899 ( N732, new_n1095_, new_n1100_ );
not g0900 ( new_n1102_, keyIn_0_109 );
or g0901 ( new_n1103_, new_n1080_, new_n475_ );
and g0902 ( new_n1104_, new_n1103_, keyIn_0_86 );
not g0903 ( new_n1105_, keyIn_0_86 );
and g0904 ( new_n1106_, new_n1085_, new_n476_ );
and g0905 ( new_n1107_, new_n1106_, new_n1105_ );
or g0906 ( new_n1108_, new_n1104_, new_n1107_ );
and g0907 ( new_n1109_, new_n1108_, N37 );
or g0908 ( new_n1110_, new_n1106_, new_n1105_ );
or g0909 ( new_n1111_, new_n1103_, keyIn_0_86 );
and g0910 ( new_n1112_, new_n1111_, new_n1110_ );
and g0911 ( new_n1113_, new_n1112_, new_n455_ );
or g0912 ( new_n1114_, new_n1109_, new_n1113_ );
or g0913 ( new_n1115_, new_n1114_, new_n1102_ );
or g0914 ( new_n1116_, new_n1112_, new_n455_ );
or g0915 ( new_n1117_, new_n1108_, N37 );
and g0916 ( new_n1118_, new_n1117_, new_n1116_ );
or g0917 ( new_n1119_, new_n1118_, keyIn_0_109 );
and g0918 ( N733, new_n1115_, new_n1119_ );
not g0919 ( new_n1121_, keyIn_0_110 );
or g0920 ( new_n1122_, new_n1080_, new_n532_ );
and g0921 ( new_n1123_, new_n1122_, keyIn_0_87 );
not g0922 ( new_n1124_, keyIn_0_87 );
and g0923 ( new_n1125_, new_n1085_, new_n399_ );
and g0924 ( new_n1126_, new_n1125_, new_n1124_ );
or g0925 ( new_n1127_, new_n1123_, new_n1126_ );
and g0926 ( new_n1128_, new_n1127_, new_n372_ );
or g0927 ( new_n1129_, new_n1125_, new_n1124_ );
or g0928 ( new_n1130_, new_n1122_, keyIn_0_87 );
and g0929 ( new_n1131_, new_n1130_, new_n1129_ );
and g0930 ( new_n1132_, new_n1131_, N41 );
or g0931 ( new_n1133_, new_n1128_, new_n1132_ );
and g0932 ( new_n1134_, new_n1133_, new_n1121_ );
or g0933 ( new_n1135_, new_n1131_, N41 );
or g0934 ( new_n1136_, new_n1127_, new_n372_ );
and g0935 ( new_n1137_, new_n1136_, new_n1135_ );
and g0936 ( new_n1138_, new_n1137_, keyIn_0_110 );
or g0937 ( N734, new_n1134_, new_n1138_ );
or g0938 ( new_n1140_, new_n1080_, new_n535_ );
and g0939 ( new_n1141_, new_n1140_, keyIn_0_88 );
not g0940 ( new_n1142_, keyIn_0_88 );
and g0941 ( new_n1143_, new_n1085_, new_n525_ );
and g0942 ( new_n1144_, new_n1143_, new_n1142_ );
or g0943 ( new_n1145_, new_n1141_, new_n1144_ );
and g0944 ( new_n1146_, new_n1145_, new_n510_ );
or g0945 ( new_n1147_, new_n1143_, new_n1142_ );
or g0946 ( new_n1148_, new_n1140_, keyIn_0_88 );
and g0947 ( new_n1149_, new_n1148_, new_n1147_ );
and g0948 ( new_n1150_, new_n1149_, N45 );
or g0949 ( new_n1151_, new_n1146_, new_n1150_ );
or g0950 ( new_n1152_, new_n1151_, keyIn_0_111 );
not g0951 ( new_n1153_, keyIn_0_111 );
or g0952 ( new_n1154_, new_n1149_, N45 );
or g0953 ( new_n1155_, new_n1145_, new_n510_ );
and g0954 ( new_n1156_, new_n1155_, new_n1154_ );
or g0955 ( new_n1157_, new_n1156_, new_n1153_ );
and g0956 ( N735, new_n1152_, new_n1157_ );
and g0957 ( new_n1159_, new_n1070_, new_n1067_ );
and g0958 ( new_n1160_, new_n989_, new_n1159_ );
and g0959 ( new_n1161_, new_n544_, new_n1160_ );
and g0960 ( new_n1162_, new_n1161_, new_n307_ );
not g0961 ( new_n1163_, new_n1162_ );
and g0962 ( new_n1164_, new_n1163_, N49 );
and g0963 ( new_n1165_, new_n1162_, new_n283_ );
or g0964 ( N736, new_n1164_, new_n1165_ );
and g0965 ( new_n1167_, new_n1161_, new_n476_ );
not g0966 ( new_n1168_, new_n1167_ );
and g0967 ( new_n1169_, new_n1168_, N53 );
and g0968 ( new_n1170_, new_n1167_, new_n453_ );
or g0969 ( N737, new_n1169_, new_n1170_ );
and g0970 ( new_n1172_, new_n1161_, new_n399_ );
not g0971 ( new_n1173_, new_n1172_ );
and g0972 ( new_n1174_, new_n1173_, N57 );
and g0973 ( new_n1175_, new_n1172_, new_n370_ );
or g0974 ( N738, new_n1174_, new_n1175_ );
and g0975 ( new_n1177_, new_n1161_, new_n525_ );
not g0976 ( new_n1178_, new_n1177_ );
and g0977 ( new_n1179_, new_n1178_, N61 );
and g0978 ( new_n1180_, new_n1177_, new_n508_ );
or g0979 ( N739, new_n1179_, new_n1180_ );
not g0980 ( new_n1182_, keyIn_0_112 );
not g0981 ( new_n1183_, keyIn_0_78 );
or g0982 ( new_n1184_, new_n1067_, new_n784_ );
or g0983 ( new_n1185_, new_n1184_, new_n949_ );
and g0984 ( new_n1186_, new_n893_, keyIn_0_64 );
not g0985 ( new_n1187_, keyIn_0_64 );
and g0986 ( new_n1188_, new_n988_, new_n1187_ );
or g0987 ( new_n1189_, new_n1188_, new_n1186_ );
or g0988 ( new_n1190_, new_n1185_, new_n1189_ );
and g0989 ( new_n1191_, new_n1190_, keyIn_0_71 );
not g0990 ( new_n1192_, keyIn_0_71 );
and g0991 ( new_n1193_, new_n690_, new_n985_ );
and g0992 ( new_n1194_, new_n1193_, new_n1070_ );
not g0993 ( new_n1195_, new_n1186_ );
or g0994 ( new_n1196_, new_n893_, keyIn_0_64 );
and g0995 ( new_n1197_, new_n1195_, new_n1196_ );
and g0996 ( new_n1198_, new_n1197_, new_n1194_ );
and g0997 ( new_n1199_, new_n1198_, new_n1192_ );
or g0998 ( new_n1200_, new_n1199_, new_n1191_ );
not g0999 ( new_n1201_, keyIn_0_73 );
not g1000 ( new_n1202_, keyIn_0_65 );
and g1001 ( new_n1203_, new_n893_, new_n1202_ );
and g1002 ( new_n1204_, new_n988_, keyIn_0_65 );
or g1003 ( new_n1205_, new_n1204_, new_n1203_ );
and g1004 ( new_n1206_, new_n1159_, new_n784_ );
and g1005 ( new_n1207_, new_n1205_, new_n1206_ );
or g1006 ( new_n1208_, new_n1207_, new_n1201_ );
and g1007 ( new_n1209_, new_n1207_, new_n1201_ );
not g1008 ( new_n1210_, new_n1209_ );
and g1009 ( new_n1211_, new_n1210_, new_n1208_ );
and g1010 ( new_n1212_, new_n1211_, new_n1200_ );
not g1011 ( new_n1213_, keyIn_0_74 );
not g1012 ( new_n1214_, keyIn_0_66 );
and g1013 ( new_n1215_, new_n893_, new_n1214_ );
and g1014 ( new_n1216_, new_n988_, keyIn_0_66 );
or g1015 ( new_n1217_, new_n1216_, new_n1215_ );
and g1016 ( new_n1218_, new_n785_, new_n949_ );
and g1017 ( new_n1219_, new_n1217_, new_n1218_ );
and g1018 ( new_n1220_, new_n1219_, new_n1213_ );
or g1019 ( new_n1221_, new_n988_, keyIn_0_66 );
or g1020 ( new_n1222_, new_n893_, new_n1214_ );
and g1021 ( new_n1223_, new_n1221_, new_n1222_ );
or g1022 ( new_n1224_, new_n985_, new_n1067_ );
or g1023 ( new_n1225_, new_n1224_, new_n1070_ );
or g1024 ( new_n1226_, new_n1225_, new_n1223_ );
and g1025 ( new_n1227_, new_n1226_, keyIn_0_74 );
or g1026 ( new_n1228_, new_n1227_, new_n1220_ );
not g1027 ( new_n1229_, keyIn_0_72 );
and g1028 ( new_n1230_, new_n1072_, new_n690_ );
or g1029 ( new_n1231_, new_n1230_, new_n1229_ );
and g1030 ( new_n1232_, new_n1070_, new_n1229_ );
and g1031 ( new_n1233_, new_n894_, new_n1232_ );
not g1032 ( new_n1234_, new_n1233_ );
and g1033 ( new_n1235_, new_n1231_, new_n1234_ );
not g1034 ( new_n1236_, new_n1235_ );
and g1035 ( new_n1237_, new_n1236_, new_n1228_ );
and g1036 ( new_n1238_, new_n1212_, new_n1237_ );
and g1037 ( new_n1239_, new_n1238_, keyIn_0_75 );
not g1038 ( new_n1240_, keyIn_0_75 );
or g1039 ( new_n1241_, new_n1198_, new_n1192_ );
or g1040 ( new_n1242_, new_n1190_, keyIn_0_71 );
and g1041 ( new_n1243_, new_n1241_, new_n1242_ );
or g1042 ( new_n1244_, new_n988_, keyIn_0_65 );
or g1043 ( new_n1245_, new_n893_, new_n1202_ );
and g1044 ( new_n1246_, new_n1244_, new_n1245_ );
or g1045 ( new_n1247_, new_n690_, new_n949_ );
or g1046 ( new_n1248_, new_n1247_, new_n985_ );
or g1047 ( new_n1249_, new_n1248_, new_n1246_ );
and g1048 ( new_n1250_, new_n1249_, keyIn_0_73 );
or g1049 ( new_n1251_, new_n1250_, new_n1209_ );
or g1050 ( new_n1252_, new_n1243_, new_n1251_ );
or g1051 ( new_n1253_, new_n1226_, keyIn_0_74 );
or g1052 ( new_n1254_, new_n1219_, new_n1213_ );
and g1053 ( new_n1255_, new_n1253_, new_n1254_ );
or g1054 ( new_n1256_, new_n1255_, new_n1235_ );
or g1055 ( new_n1257_, new_n1252_, new_n1256_ );
and g1056 ( new_n1258_, new_n1257_, new_n1240_ );
or g1057 ( new_n1259_, new_n1258_, new_n1239_ );
not g1058 ( new_n1260_, keyIn_0_67 );
and g1059 ( new_n1261_, new_n475_, new_n1260_ );
not g1060 ( new_n1262_, new_n1261_ );
and g1061 ( new_n1263_, new_n476_, keyIn_0_67 );
not g1062 ( new_n1264_, new_n1263_ );
and g1063 ( new_n1265_, new_n307_, new_n535_ );
and g1064 ( new_n1266_, new_n1265_, new_n1264_ );
and g1065 ( new_n1267_, new_n1266_, new_n1262_ );
and g1066 ( new_n1268_, new_n1267_, new_n399_ );
and g1067 ( new_n1269_, new_n1259_, new_n1268_ );
and g1068 ( new_n1270_, new_n1269_, new_n1183_ );
or g1069 ( new_n1271_, new_n1257_, new_n1240_ );
or g1070 ( new_n1272_, new_n1238_, keyIn_0_75 );
and g1071 ( new_n1273_, new_n1271_, new_n1272_ );
not g1072 ( new_n1274_, new_n1268_ );
or g1073 ( new_n1275_, new_n1273_, new_n1274_ );
and g1074 ( new_n1276_, new_n1275_, keyIn_0_78 );
or g1075 ( new_n1277_, new_n1276_, new_n1070_ );
or g1076 ( new_n1278_, new_n1277_, new_n1270_ );
and g1077 ( new_n1279_, new_n1278_, keyIn_0_89 );
not g1078 ( new_n1280_, keyIn_0_89 );
not g1079 ( new_n1281_, new_n1270_ );
or g1080 ( new_n1282_, new_n1269_, new_n1183_ );
and g1081 ( new_n1283_, new_n1282_, new_n949_ );
and g1082 ( new_n1284_, new_n1283_, new_n1281_ );
and g1083 ( new_n1285_, new_n1284_, new_n1280_ );
or g1084 ( new_n1286_, new_n1279_, new_n1285_ );
and g1085 ( new_n1287_, new_n1286_, new_n238_ );
or g1086 ( new_n1288_, new_n1284_, new_n1280_ );
or g1087 ( new_n1289_, new_n1278_, keyIn_0_89 );
and g1088 ( new_n1290_, new_n1289_, new_n1288_ );
and g1089 ( new_n1291_, new_n1290_, N65 );
or g1090 ( new_n1292_, new_n1287_, new_n1291_ );
and g1091 ( new_n1293_, new_n1292_, new_n1182_ );
or g1092 ( new_n1294_, new_n1290_, N65 );
or g1093 ( new_n1295_, new_n1286_, new_n238_ );
and g1094 ( new_n1296_, new_n1294_, new_n1295_ );
and g1095 ( new_n1297_, new_n1296_, keyIn_0_112 );
or g1096 ( N740, new_n1293_, new_n1297_ );
not g1097 ( new_n1299_, keyIn_0_113 );
not g1098 ( new_n1300_, keyIn_0_90 );
or g1099 ( new_n1301_, new_n1276_, new_n690_ );
or g1100 ( new_n1302_, new_n1301_, new_n1270_ );
and g1101 ( new_n1303_, new_n1302_, new_n1300_ );
and g1102 ( new_n1304_, new_n1282_, new_n1067_ );
and g1103 ( new_n1305_, new_n1304_, new_n1281_ );
and g1104 ( new_n1306_, new_n1305_, keyIn_0_90 );
or g1105 ( new_n1307_, new_n1303_, new_n1306_ );
and g1106 ( new_n1308_, new_n1307_, new_n236_ );
or g1107 ( new_n1309_, new_n1305_, keyIn_0_90 );
or g1108 ( new_n1310_, new_n1302_, new_n1300_ );
and g1109 ( new_n1311_, new_n1310_, new_n1309_ );
and g1110 ( new_n1312_, new_n1311_, N69 );
or g1111 ( new_n1313_, new_n1308_, new_n1312_ );
or g1112 ( new_n1314_, new_n1313_, new_n1299_ );
or g1113 ( new_n1315_, new_n1311_, N69 );
or g1114 ( new_n1316_, new_n1307_, new_n236_ );
and g1115 ( new_n1317_, new_n1315_, new_n1316_ );
or g1116 ( new_n1318_, new_n1317_, keyIn_0_113 );
and g1117 ( N741, new_n1314_, new_n1318_ );
not g1118 ( new_n1320_, keyIn_0_91 );
or g1119 ( new_n1321_, new_n1276_, new_n988_ );
or g1120 ( new_n1322_, new_n1321_, new_n1270_ );
and g1121 ( new_n1323_, new_n1322_, new_n1320_ );
and g1122 ( new_n1324_, new_n1282_, new_n893_ );
and g1123 ( new_n1325_, new_n1324_, new_n1281_ );
and g1124 ( new_n1326_, new_n1325_, keyIn_0_91 );
or g1125 ( new_n1327_, new_n1323_, new_n1326_ );
and g1126 ( new_n1328_, new_n1327_, new_n249_ );
or g1127 ( new_n1329_, new_n1325_, keyIn_0_91 );
or g1128 ( new_n1330_, new_n1322_, new_n1320_ );
and g1129 ( new_n1331_, new_n1330_, new_n1329_ );
and g1130 ( new_n1332_, new_n1331_, N73 );
or g1131 ( new_n1333_, new_n1328_, new_n1332_ );
and g1132 ( new_n1334_, new_n1333_, keyIn_0_114 );
not g1133 ( new_n1335_, keyIn_0_114 );
or g1134 ( new_n1336_, new_n1331_, N73 );
or g1135 ( new_n1337_, new_n1327_, new_n249_ );
and g1136 ( new_n1338_, new_n1336_, new_n1337_ );
and g1137 ( new_n1339_, new_n1338_, new_n1335_ );
or g1138 ( N742, new_n1334_, new_n1339_ );
or g1139 ( new_n1341_, new_n1276_, new_n784_ );
or g1140 ( new_n1342_, new_n1341_, new_n1270_ );
and g1141 ( new_n1343_, new_n1342_, keyIn_0_92 );
not g1142 ( new_n1344_, keyIn_0_92 );
and g1143 ( new_n1345_, new_n1282_, new_n985_ );
and g1144 ( new_n1346_, new_n1345_, new_n1281_ );
and g1145 ( new_n1347_, new_n1346_, new_n1344_ );
or g1146 ( new_n1348_, new_n1343_, new_n1347_ );
and g1147 ( new_n1349_, new_n1348_, new_n247_ );
or g1148 ( new_n1350_, new_n1346_, new_n1344_ );
or g1149 ( new_n1351_, new_n1342_, keyIn_0_92 );
and g1150 ( new_n1352_, new_n1351_, new_n1350_ );
and g1151 ( new_n1353_, new_n1352_, N77 );
or g1152 ( new_n1354_, new_n1349_, new_n1353_ );
and g1153 ( new_n1355_, new_n1354_, keyIn_0_115 );
not g1154 ( new_n1356_, keyIn_0_115 );
or g1155 ( new_n1357_, new_n1352_, N77 );
or g1156 ( new_n1358_, new_n1348_, new_n247_ );
and g1157 ( new_n1359_, new_n1357_, new_n1358_ );
and g1158 ( new_n1360_, new_n1359_, new_n1356_ );
or g1159 ( N743, new_n1355_, new_n1360_ );
not g1160 ( new_n1362_, keyIn_0_116 );
not g1161 ( new_n1363_, keyIn_0_93 );
not g1162 ( new_n1364_, keyIn_0_68 );
and g1163 ( new_n1365_, new_n399_, new_n1364_ );
not g1164 ( new_n1366_, new_n1365_ );
and g1165 ( new_n1367_, new_n532_, keyIn_0_68 );
not g1166 ( new_n1368_, new_n1367_ );
not g1167 ( new_n1369_, new_n477_ );
and g1168 ( new_n1370_, new_n1369_, new_n525_ );
and g1169 ( new_n1371_, new_n1368_, new_n1370_ );
and g1170 ( new_n1372_, new_n1371_, new_n1366_ );
and g1171 ( new_n1373_, new_n1259_, new_n1372_ );
and g1172 ( new_n1374_, new_n1373_, keyIn_0_79 );
not g1173 ( new_n1375_, keyIn_0_79 );
not g1174 ( new_n1376_, new_n1372_ );
or g1175 ( new_n1377_, new_n1273_, new_n1376_ );
and g1176 ( new_n1378_, new_n1377_, new_n1375_ );
or g1177 ( new_n1379_, new_n1378_, new_n1070_ );
or g1178 ( new_n1380_, new_n1379_, new_n1374_ );
and g1179 ( new_n1381_, new_n1380_, new_n1363_ );
not g1180 ( new_n1382_, new_n1374_ );
or g1181 ( new_n1383_, new_n1373_, keyIn_0_79 );
and g1182 ( new_n1384_, new_n1383_, new_n949_ );
and g1183 ( new_n1385_, new_n1384_, new_n1382_ );
and g1184 ( new_n1386_, new_n1385_, keyIn_0_93 );
or g1185 ( new_n1387_, new_n1381_, new_n1386_ );
and g1186 ( new_n1388_, new_n1387_, new_n207_ );
or g1187 ( new_n1389_, new_n1385_, keyIn_0_93 );
or g1188 ( new_n1390_, new_n1380_, new_n1363_ );
and g1189 ( new_n1391_, new_n1390_, new_n1389_ );
and g1190 ( new_n1392_, new_n1391_, N81 );
or g1191 ( new_n1393_, new_n1388_, new_n1392_ );
or g1192 ( new_n1394_, new_n1393_, new_n1362_ );
or g1193 ( new_n1395_, new_n1391_, N81 );
or g1194 ( new_n1396_, new_n1387_, new_n207_ );
and g1195 ( new_n1397_, new_n1395_, new_n1396_ );
or g1196 ( new_n1398_, new_n1397_, keyIn_0_116 );
and g1197 ( N744, new_n1394_, new_n1398_ );
not g1198 ( new_n1400_, keyIn_0_117 );
or g1199 ( new_n1401_, new_n1378_, new_n690_ );
or g1200 ( new_n1402_, new_n1401_, new_n1374_ );
and g1201 ( new_n1403_, new_n1402_, keyIn_0_94 );
not g1202 ( new_n1404_, keyIn_0_94 );
and g1203 ( new_n1405_, new_n1383_, new_n1067_ );
and g1204 ( new_n1406_, new_n1405_, new_n1382_ );
and g1205 ( new_n1407_, new_n1406_, new_n1404_ );
or g1206 ( new_n1408_, new_n1403_, new_n1407_ );
and g1207 ( new_n1409_, new_n1408_, new_n205_ );
or g1208 ( new_n1410_, new_n1406_, new_n1404_ );
or g1209 ( new_n1411_, new_n1402_, keyIn_0_94 );
and g1210 ( new_n1412_, new_n1411_, new_n1410_ );
and g1211 ( new_n1413_, new_n1412_, N85 );
or g1212 ( new_n1414_, new_n1409_, new_n1413_ );
or g1213 ( new_n1415_, new_n1414_, new_n1400_ );
or g1214 ( new_n1416_, new_n1412_, N85 );
or g1215 ( new_n1417_, new_n1408_, new_n205_ );
and g1216 ( new_n1418_, new_n1416_, new_n1417_ );
or g1217 ( new_n1419_, new_n1418_, keyIn_0_117 );
and g1218 ( N745, new_n1415_, new_n1419_ );
not g1219 ( new_n1421_, keyIn_0_118 );
or g1220 ( new_n1422_, new_n1378_, new_n988_ );
or g1221 ( new_n1423_, new_n1422_, new_n1374_ );
and g1222 ( new_n1424_, new_n1423_, keyIn_0_95 );
not g1223 ( new_n1425_, keyIn_0_95 );
and g1224 ( new_n1426_, new_n1383_, new_n893_ );
and g1225 ( new_n1427_, new_n1426_, new_n1382_ );
and g1226 ( new_n1428_, new_n1427_, new_n1425_ );
or g1227 ( new_n1429_, new_n1424_, new_n1428_ );
and g1228 ( new_n1430_, new_n1429_, N89 );
or g1229 ( new_n1431_, new_n1427_, new_n1425_ );
or g1230 ( new_n1432_, new_n1423_, keyIn_0_95 );
and g1231 ( new_n1433_, new_n1432_, new_n1431_ );
and g1232 ( new_n1434_, new_n1433_, new_n217_ );
or g1233 ( new_n1435_, new_n1430_, new_n1434_ );
or g1234 ( new_n1436_, new_n1435_, new_n1421_ );
or g1235 ( new_n1437_, new_n1433_, new_n217_ );
or g1236 ( new_n1438_, new_n1429_, N89 );
and g1237 ( new_n1439_, new_n1437_, new_n1438_ );
or g1238 ( new_n1440_, new_n1439_, keyIn_0_118 );
and g1239 ( N746, new_n1436_, new_n1440_ );
or g1240 ( new_n1442_, new_n1378_, new_n784_ );
or g1241 ( new_n1443_, new_n1442_, new_n1374_ );
and g1242 ( new_n1444_, new_n1443_, keyIn_0_96 );
not g1243 ( new_n1445_, keyIn_0_96 );
and g1244 ( new_n1446_, new_n1383_, new_n985_ );
and g1245 ( new_n1447_, new_n1446_, new_n1382_ );
and g1246 ( new_n1448_, new_n1447_, new_n1445_ );
or g1247 ( new_n1449_, new_n1444_, new_n1448_ );
and g1248 ( new_n1450_, new_n1449_, N93 );
or g1249 ( new_n1451_, new_n1447_, new_n1445_ );
or g1250 ( new_n1452_, new_n1443_, keyIn_0_96 );
and g1251 ( new_n1453_, new_n1452_, new_n1451_ );
and g1252 ( new_n1454_, new_n1453_, new_n215_ );
or g1253 ( new_n1455_, new_n1450_, new_n1454_ );
and g1254 ( new_n1456_, new_n1455_, keyIn_0_119 );
not g1255 ( new_n1457_, keyIn_0_119 );
or g1256 ( new_n1458_, new_n1453_, new_n215_ );
or g1257 ( new_n1459_, new_n1449_, N93 );
and g1258 ( new_n1460_, new_n1458_, new_n1459_ );
and g1259 ( new_n1461_, new_n1460_, new_n1457_ );
or g1260 ( N747, new_n1456_, new_n1461_ );
not g1261 ( new_n1463_, keyIn_0_97 );
not g1262 ( new_n1464_, keyIn_0_80 );
and g1263 ( new_n1465_, new_n306_, new_n476_ );
and g1264 ( new_n1466_, new_n1465_, new_n535_ );
and g1265 ( new_n1467_, new_n1466_, new_n399_ );
and g1266 ( new_n1468_, new_n1259_, new_n1467_ );
and g1267 ( new_n1469_, new_n1468_, new_n1464_ );
not g1268 ( new_n1470_, new_n1467_ );
or g1269 ( new_n1471_, new_n1273_, new_n1470_ );
and g1270 ( new_n1472_, new_n1471_, keyIn_0_80 );
or g1271 ( new_n1473_, new_n1472_, new_n1070_ );
or g1272 ( new_n1474_, new_n1473_, new_n1469_ );
and g1273 ( new_n1475_, new_n1474_, new_n1463_ );
not g1274 ( new_n1476_, new_n1469_ );
or g1275 ( new_n1477_, new_n1468_, new_n1464_ );
and g1276 ( new_n1478_, new_n1477_, new_n949_ );
and g1277 ( new_n1479_, new_n1478_, new_n1476_ );
and g1278 ( new_n1480_, new_n1479_, keyIn_0_97 );
or g1279 ( new_n1481_, new_n1475_, new_n1480_ );
and g1280 ( new_n1482_, new_n1481_, N97 );
or g1281 ( new_n1483_, new_n1479_, keyIn_0_97 );
or g1282 ( new_n1484_, new_n1474_, new_n1463_ );
and g1283 ( new_n1485_, new_n1484_, new_n1483_ );
and g1284 ( new_n1486_, new_n1485_, new_n313_ );
or g1285 ( new_n1487_, new_n1482_, new_n1486_ );
and g1286 ( new_n1488_, new_n1487_, keyIn_0_120 );
not g1287 ( new_n1489_, keyIn_0_120 );
or g1288 ( new_n1490_, new_n1485_, new_n313_ );
or g1289 ( new_n1491_, new_n1481_, N97 );
and g1290 ( new_n1492_, new_n1490_, new_n1491_ );
and g1291 ( new_n1493_, new_n1492_, new_n1489_ );
or g1292 ( N748, new_n1488_, new_n1493_ );
not g1293 ( new_n1495_, keyIn_0_121 );
or g1294 ( new_n1496_, new_n1472_, new_n690_ );
or g1295 ( new_n1497_, new_n1496_, new_n1469_ );
and g1296 ( new_n1498_, new_n1497_, keyIn_0_98 );
not g1297 ( new_n1499_, keyIn_0_98 );
and g1298 ( new_n1500_, new_n1477_, new_n1067_ );
and g1299 ( new_n1501_, new_n1500_, new_n1476_ );
and g1300 ( new_n1502_, new_n1501_, new_n1499_ );
or g1301 ( new_n1503_, new_n1498_, new_n1502_ );
and g1302 ( new_n1504_, new_n1503_, new_n311_ );
or g1303 ( new_n1505_, new_n1501_, new_n1499_ );
or g1304 ( new_n1506_, new_n1497_, keyIn_0_98 );
and g1305 ( new_n1507_, new_n1506_, new_n1505_ );
and g1306 ( new_n1508_, new_n1507_, N101 );
or g1307 ( new_n1509_, new_n1504_, new_n1508_ );
or g1308 ( new_n1510_, new_n1509_, new_n1495_ );
or g1309 ( new_n1511_, new_n1507_, N101 );
or g1310 ( new_n1512_, new_n1503_, new_n311_ );
and g1311 ( new_n1513_, new_n1511_, new_n1512_ );
or g1312 ( new_n1514_, new_n1513_, keyIn_0_121 );
and g1313 ( N749, new_n1510_, new_n1514_ );
not g1314 ( new_n1516_, keyIn_0_99 );
or g1315 ( new_n1517_, new_n1472_, new_n988_ );
or g1316 ( new_n1518_, new_n1517_, new_n1469_ );
and g1317 ( new_n1519_, new_n1518_, new_n1516_ );
and g1318 ( new_n1520_, new_n1477_, new_n893_ );
and g1319 ( new_n1521_, new_n1520_, new_n1476_ );
and g1320 ( new_n1522_, new_n1521_, keyIn_0_99 );
or g1321 ( new_n1523_, new_n1519_, new_n1522_ );
and g1322 ( new_n1524_, new_n1523_, N105 );
or g1323 ( new_n1525_, new_n1521_, keyIn_0_99 );
or g1324 ( new_n1526_, new_n1518_, new_n1516_ );
and g1325 ( new_n1527_, new_n1526_, new_n1525_ );
and g1326 ( new_n1528_, new_n1527_, new_n324_ );
or g1327 ( new_n1529_, new_n1524_, new_n1528_ );
or g1328 ( new_n1530_, new_n1529_, keyIn_0_122 );
not g1329 ( new_n1531_, keyIn_0_122 );
or g1330 ( new_n1532_, new_n1527_, new_n324_ );
or g1331 ( new_n1533_, new_n1523_, N105 );
and g1332 ( new_n1534_, new_n1532_, new_n1533_ );
or g1333 ( new_n1535_, new_n1534_, new_n1531_ );
and g1334 ( N750, new_n1530_, new_n1535_ );
not g1335 ( new_n1537_, keyIn_0_123 );
not g1336 ( new_n1538_, keyIn_0_100 );
or g1337 ( new_n1539_, new_n1472_, new_n784_ );
or g1338 ( new_n1540_, new_n1539_, new_n1469_ );
and g1339 ( new_n1541_, new_n1540_, new_n1538_ );
and g1340 ( new_n1542_, new_n1477_, new_n985_ );
and g1341 ( new_n1543_, new_n1542_, new_n1476_ );
and g1342 ( new_n1544_, new_n1543_, keyIn_0_100 );
or g1343 ( new_n1545_, new_n1541_, new_n1544_ );
and g1344 ( new_n1546_, new_n1545_, N109 );
or g1345 ( new_n1547_, new_n1543_, keyIn_0_100 );
or g1346 ( new_n1548_, new_n1540_, new_n1538_ );
and g1347 ( new_n1549_, new_n1548_, new_n1547_ );
and g1348 ( new_n1550_, new_n1549_, new_n322_ );
or g1349 ( new_n1551_, new_n1546_, new_n1550_ );
or g1350 ( new_n1552_, new_n1551_, new_n1537_ );
or g1351 ( new_n1553_, new_n1549_, new_n322_ );
or g1352 ( new_n1554_, new_n1545_, N109 );
and g1353 ( new_n1555_, new_n1553_, new_n1554_ );
or g1354 ( new_n1556_, new_n1555_, keyIn_0_123 );
and g1355 ( N751, new_n1552_, new_n1556_ );
not g1356 ( new_n1558_, keyIn_0_101 );
not g1357 ( new_n1559_, keyIn_0_81 );
and g1358 ( new_n1560_, new_n399_, keyIn_0_70 );
not g1359 ( new_n1561_, new_n1560_ );
or g1360 ( new_n1562_, new_n399_, keyIn_0_70 );
and g1361 ( new_n1563_, new_n1561_, new_n1562_ );
not g1362 ( new_n1564_, keyIn_0_69 );
and g1363 ( new_n1565_, new_n306_, new_n1564_ );
and g1364 ( new_n1566_, new_n307_, keyIn_0_69 );
or g1365 ( new_n1567_, new_n1566_, new_n540_ );
or g1366 ( new_n1568_, new_n1567_, new_n1565_ );
or g1367 ( new_n1569_, new_n1563_, new_n1568_ );
not g1368 ( new_n1570_, new_n1569_ );
and g1369 ( new_n1571_, new_n1259_, new_n1570_ );
and g1370 ( new_n1572_, new_n1571_, new_n1559_ );
or g1371 ( new_n1573_, new_n1273_, new_n1569_ );
and g1372 ( new_n1574_, new_n1573_, keyIn_0_81 );
or g1373 ( new_n1575_, new_n1574_, new_n1070_ );
or g1374 ( new_n1576_, new_n1575_, new_n1572_ );
and g1375 ( new_n1577_, new_n1576_, new_n1558_ );
not g1376 ( new_n1578_, new_n1572_ );
or g1377 ( new_n1579_, new_n1571_, new_n1559_ );
and g1378 ( new_n1580_, new_n1579_, new_n949_ );
and g1379 ( new_n1581_, new_n1580_, new_n1578_ );
and g1380 ( new_n1582_, new_n1581_, keyIn_0_101 );
or g1381 ( new_n1583_, new_n1577_, new_n1582_ );
and g1382 ( new_n1584_, new_n1583_, new_n409_ );
or g1383 ( new_n1585_, new_n1581_, keyIn_0_101 );
or g1384 ( new_n1586_, new_n1576_, new_n1558_ );
and g1385 ( new_n1587_, new_n1586_, new_n1585_ );
and g1386 ( new_n1588_, new_n1587_, N113 );
or g1387 ( new_n1589_, new_n1584_, new_n1588_ );
or g1388 ( new_n1590_, new_n1589_, keyIn_0_124 );
not g1389 ( new_n1591_, keyIn_0_124 );
or g1390 ( new_n1592_, new_n1587_, N113 );
or g1391 ( new_n1593_, new_n1583_, new_n409_ );
and g1392 ( new_n1594_, new_n1592_, new_n1593_ );
or g1393 ( new_n1595_, new_n1594_, new_n1591_ );
and g1394 ( N752, new_n1590_, new_n1595_ );
or g1395 ( new_n1597_, new_n1574_, new_n690_ );
or g1396 ( new_n1598_, new_n1597_, new_n1572_ );
and g1397 ( new_n1599_, new_n1598_, keyIn_0_102 );
not g1398 ( new_n1600_, keyIn_0_102 );
and g1399 ( new_n1601_, new_n1579_, new_n1067_ );
and g1400 ( new_n1602_, new_n1601_, new_n1578_ );
and g1401 ( new_n1603_, new_n1602_, new_n1600_ );
or g1402 ( new_n1604_, new_n1599_, new_n1603_ );
and g1403 ( new_n1605_, new_n1604_, N117 );
or g1404 ( new_n1606_, new_n1602_, new_n1600_ );
or g1405 ( new_n1607_, new_n1598_, keyIn_0_102 );
and g1406 ( new_n1608_, new_n1607_, new_n1606_ );
and g1407 ( new_n1609_, new_n1608_, new_n407_ );
or g1408 ( new_n1610_, new_n1605_, new_n1609_ );
and g1409 ( new_n1611_, new_n1610_, keyIn_0_125 );
not g1410 ( new_n1612_, keyIn_0_125 );
or g1411 ( new_n1613_, new_n1608_, new_n407_ );
or g1412 ( new_n1614_, new_n1604_, N117 );
and g1413 ( new_n1615_, new_n1613_, new_n1614_ );
and g1414 ( new_n1616_, new_n1615_, new_n1612_ );
or g1415 ( N753, new_n1611_, new_n1616_ );
not g1416 ( new_n1618_, keyIn_0_126 );
or g1417 ( new_n1619_, new_n1574_, new_n988_ );
or g1418 ( new_n1620_, new_n1619_, new_n1572_ );
and g1419 ( new_n1621_, new_n1620_, keyIn_0_103 );
not g1420 ( new_n1622_, keyIn_0_103 );
and g1421 ( new_n1623_, new_n1579_, new_n893_ );
and g1422 ( new_n1624_, new_n1623_, new_n1578_ );
and g1423 ( new_n1625_, new_n1624_, new_n1622_ );
or g1424 ( new_n1626_, new_n1621_, new_n1625_ );
and g1425 ( new_n1627_, new_n1626_, new_n420_ );
or g1426 ( new_n1628_, new_n1624_, new_n1622_ );
or g1427 ( new_n1629_, new_n1620_, keyIn_0_103 );
and g1428 ( new_n1630_, new_n1629_, new_n1628_ );
and g1429 ( new_n1631_, new_n1630_, N121 );
or g1430 ( new_n1632_, new_n1627_, new_n1631_ );
and g1431 ( new_n1633_, new_n1632_, new_n1618_ );
or g1432 ( new_n1634_, new_n1630_, N121 );
or g1433 ( new_n1635_, new_n1626_, new_n420_ );
and g1434 ( new_n1636_, new_n1634_, new_n1635_ );
and g1435 ( new_n1637_, new_n1636_, keyIn_0_126 );
or g1436 ( N754, new_n1633_, new_n1637_ );
not g1437 ( new_n1639_, keyIn_0_127 );
or g1438 ( new_n1640_, new_n1574_, new_n784_ );
or g1439 ( new_n1641_, new_n1640_, new_n1572_ );
and g1440 ( new_n1642_, new_n1641_, keyIn_0_104 );
not g1441 ( new_n1643_, keyIn_0_104 );
and g1442 ( new_n1644_, new_n1579_, new_n985_ );
and g1443 ( new_n1645_, new_n1644_, new_n1578_ );
and g1444 ( new_n1646_, new_n1645_, new_n1643_ );
or g1445 ( new_n1647_, new_n1642_, new_n1646_ );
and g1446 ( new_n1648_, new_n1647_, N125 );
or g1447 ( new_n1649_, new_n1645_, new_n1643_ );
or g1448 ( new_n1650_, new_n1641_, keyIn_0_104 );
and g1449 ( new_n1651_, new_n1650_, new_n1649_ );
and g1450 ( new_n1652_, new_n1651_, new_n418_ );
or g1451 ( new_n1653_, new_n1648_, new_n1652_ );
or g1452 ( new_n1654_, new_n1653_, new_n1639_ );
or g1453 ( new_n1655_, new_n1651_, new_n418_ );
or g1454 ( new_n1656_, new_n1647_, N125 );
and g1455 ( new_n1657_, new_n1655_, new_n1656_ );
or g1456 ( new_n1658_, new_n1657_, keyIn_0_127 );
and g1457 ( N755, new_n1654_, new_n1658_ );
endmodule