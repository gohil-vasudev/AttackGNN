module locked_c3540 (  G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698, G2897, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,  G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698, G2897, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n143_, new_n144_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1251_, new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1281_, new_n1282_, new_n1283_, new_n1284_;
  NOR2_X1 g0000 ( .A1(G58), .A2(G68), .ZN(new_n137_) );
  INV_X1 g0001 ( .A(new_n137_), .ZN(new_n138_) );
  INV_X1 g0002 ( .A(G50), .ZN(new_n139_) );
  INV_X1 g0003 ( .A(G77), .ZN(new_n140_) );
  NAND2_X1 g0004 ( .A1(new_n139_), .A2(new_n140_), .ZN(new_n141_) );
  NOR2_X1 g0005 ( .A1(new_n138_), .A2(new_n141_), .ZN(G353) );
  NOR2_X1 g0006 ( .A1(G97), .A2(G107), .ZN(new_n143_) );
  INV_X1 g0007 ( .A(new_n143_), .ZN(new_n144_) );
  NAND2_X1 g0008 ( .A1(new_n144_), .A2(G87), .ZN(G355) );
  INV_X1 g0009 ( .A(KEYINPUT49), .ZN(new_n146_) );
  NAND2_X1 g0010 ( .A1(G68), .A2(G238), .ZN(new_n147_) );
  NAND2_X1 g0011 ( .A1(G77), .A2(G244), .ZN(new_n148_) );
  NAND2_X1 g0012 ( .A1(G50), .A2(G226), .ZN(new_n149_) );
  NAND2_X1 g0013 ( .A1(G58), .A2(G232), .ZN(new_n150_) );
  NAND4_X1 g0014 ( .A1(new_n147_), .A2(new_n148_), .A3(new_n149_), .A4(new_n150_), .ZN(new_n151_) );
  NAND2_X1 g0015 ( .A1(new_n151_), .A2(new_n146_), .ZN(new_n152_) );
  NOR2_X1 g0016 ( .A1(new_n151_), .A2(new_n146_), .ZN(new_n153_) );
  NAND2_X1 g0017 ( .A1(G87), .A2(G250), .ZN(new_n154_) );
  NAND2_X1 g0018 ( .A1(G116), .A2(G270), .ZN(new_n155_) );
  NAND2_X1 g0019 ( .A1(G97), .A2(G257), .ZN(new_n156_) );
  NAND3_X1 g0020 ( .A1(new_n154_), .A2(new_n155_), .A3(new_n156_), .ZN(new_n157_) );
  NAND3_X1 g0021 ( .A1(G107), .A2(G264), .A3(KEYINPUT50), .ZN(new_n158_) );
  INV_X1 g0022 ( .A(KEYINPUT50), .ZN(new_n159_) );
  NAND2_X1 g0023 ( .A1(G107), .A2(G264), .ZN(new_n160_) );
  NAND2_X1 g0024 ( .A1(new_n160_), .A2(new_n159_), .ZN(new_n161_) );
  NAND2_X1 g0025 ( .A1(new_n161_), .A2(new_n158_), .ZN(new_n162_) );
  NOR3_X1 g0026 ( .A1(new_n153_), .A2(new_n157_), .A3(new_n162_), .ZN(new_n163_) );
  NAND2_X1 g0027 ( .A1(new_n163_), .A2(new_n152_), .ZN(new_n164_) );
  NAND2_X1 g0028 ( .A1(G1), .A2(G20), .ZN(new_n165_) );
  NAND2_X1 g0029 ( .A1(new_n164_), .A2(new_n165_), .ZN(new_n166_) );
  INV_X1 g0030 ( .A(KEYINPUT2), .ZN(new_n167_) );
  NAND2_X1 g0031 ( .A1(G1), .A2(G13), .ZN(new_n168_) );
  NAND2_X1 g0032 ( .A1(new_n168_), .A2(new_n167_), .ZN(new_n169_) );
  NAND3_X1 g0033 ( .A1(G1), .A2(G13), .A3(KEYINPUT2), .ZN(new_n170_) );
  NAND2_X1 g0034 ( .A1(new_n169_), .A2(new_n170_), .ZN(new_n171_) );
  NAND2_X1 g0035 ( .A1(new_n171_), .A2(G20), .ZN(new_n172_) );
  INV_X1 g0036 ( .A(new_n172_), .ZN(new_n173_) );
  NOR2_X1 g0037 ( .A1(new_n137_), .A2(new_n139_), .ZN(new_n174_) );
  NAND2_X1 g0038 ( .A1(new_n173_), .A2(new_n174_), .ZN(new_n175_) );
  NOR2_X1 g0039 ( .A1(new_n165_), .A2(G13), .ZN(new_n176_) );
  INV_X1 g0040 ( .A(G257), .ZN(new_n177_) );
  INV_X1 g0041 ( .A(G264), .ZN(new_n178_) );
  NAND2_X1 g0042 ( .A1(new_n177_), .A2(new_n178_), .ZN(new_n179_) );
  NAND3_X1 g0043 ( .A1(new_n176_), .A2(G250), .A3(new_n179_), .ZN(new_n180_) );
  NAND3_X1 g0044 ( .A1(new_n166_), .A2(new_n175_), .A3(new_n180_), .ZN(new_n181_) );
  INV_X1 g0045 ( .A(new_n181_), .ZN(G361) );
  INV_X1 g0046 ( .A(G238), .ZN(new_n183_) );
  NOR2_X1 g0047 ( .A1(G232), .A2(G244), .ZN(new_n184_) );
  INV_X1 g0048 ( .A(new_n184_), .ZN(new_n185_) );
  NAND2_X1 g0049 ( .A1(G232), .A2(G244), .ZN(new_n186_) );
  NAND2_X1 g0050 ( .A1(new_n185_), .A2(new_n186_), .ZN(new_n187_) );
  NAND2_X1 g0051 ( .A1(new_n187_), .A2(G226), .ZN(new_n188_) );
  INV_X1 g0052 ( .A(new_n188_), .ZN(new_n189_) );
  NOR2_X1 g0053 ( .A1(new_n187_), .A2(G226), .ZN(new_n190_) );
  NOR2_X1 g0054 ( .A1(new_n189_), .A2(new_n190_), .ZN(new_n191_) );
  INV_X1 g0055 ( .A(new_n191_), .ZN(new_n192_) );
  NAND2_X1 g0056 ( .A1(new_n192_), .A2(new_n183_), .ZN(new_n193_) );
  NAND2_X1 g0057 ( .A1(new_n191_), .A2(G238), .ZN(new_n194_) );
  INV_X1 g0058 ( .A(G270), .ZN(new_n195_) );
  NAND2_X1 g0059 ( .A1(new_n178_), .A2(new_n195_), .ZN(new_n196_) );
  NAND2_X1 g0060 ( .A1(G264), .A2(G270), .ZN(new_n197_) );
  NAND2_X1 g0061 ( .A1(new_n196_), .A2(new_n197_), .ZN(new_n198_) );
  INV_X1 g0062 ( .A(G250), .ZN(new_n199_) );
  NAND2_X1 g0063 ( .A1(new_n199_), .A2(new_n177_), .ZN(new_n200_) );
  NAND2_X1 g0064 ( .A1(G250), .A2(G257), .ZN(new_n201_) );
  NAND2_X1 g0065 ( .A1(new_n200_), .A2(new_n201_), .ZN(new_n202_) );
  NAND2_X1 g0066 ( .A1(new_n198_), .A2(new_n202_), .ZN(new_n203_) );
  NAND4_X1 g0067 ( .A1(new_n196_), .A2(new_n200_), .A3(new_n197_), .A4(new_n201_), .ZN(new_n204_) );
  NAND2_X1 g0068 ( .A1(new_n203_), .A2(new_n204_), .ZN(new_n205_) );
  NAND3_X1 g0069 ( .A1(new_n193_), .A2(new_n194_), .A3(new_n205_), .ZN(new_n206_) );
  NAND2_X1 g0070 ( .A1(new_n193_), .A2(new_n194_), .ZN(new_n207_) );
  NAND3_X1 g0071 ( .A1(new_n207_), .A2(new_n203_), .A3(new_n204_), .ZN(new_n208_) );
  NAND2_X1 g0072 ( .A1(new_n208_), .A2(new_n206_), .ZN(G358) );
  INV_X1 g0073 ( .A(KEYINPUT51), .ZN(new_n210_) );
  NAND2_X1 g0074 ( .A1(G97), .A2(G107), .ZN(new_n211_) );
  NAND2_X1 g0075 ( .A1(new_n144_), .A2(new_n211_), .ZN(new_n212_) );
  INV_X1 g0076 ( .A(new_n212_), .ZN(new_n213_) );
  NAND2_X1 g0077 ( .A1(new_n213_), .A2(new_n210_), .ZN(new_n214_) );
  NAND2_X1 g0078 ( .A1(new_n212_), .A2(KEYINPUT51), .ZN(new_n215_) );
  NAND2_X1 g0079 ( .A1(new_n214_), .A2(new_n215_), .ZN(new_n216_) );
  INV_X1 g0080 ( .A(G87), .ZN(new_n217_) );
  NOR2_X1 g0081 ( .A1(new_n217_), .A2(G116), .ZN(new_n218_) );
  INV_X1 g0082 ( .A(G116), .ZN(new_n219_) );
  NOR2_X1 g0083 ( .A1(new_n219_), .A2(G87), .ZN(new_n220_) );
  NOR2_X1 g0084 ( .A1(new_n218_), .A2(new_n220_), .ZN(new_n221_) );
  INV_X1 g0085 ( .A(new_n221_), .ZN(new_n222_) );
  NAND2_X1 g0086 ( .A1(new_n216_), .A2(new_n222_), .ZN(new_n223_) );
  NAND3_X1 g0087 ( .A1(new_n214_), .A2(new_n215_), .A3(new_n221_), .ZN(new_n224_) );
  NAND2_X1 g0088 ( .A1(new_n223_), .A2(new_n224_), .ZN(new_n225_) );
  NAND2_X1 g0089 ( .A1(G58), .A2(G68), .ZN(new_n226_) );
  NAND2_X1 g0090 ( .A1(new_n138_), .A2(new_n226_), .ZN(new_n227_) );
  NAND2_X1 g0091 ( .A1(G50), .A2(G77), .ZN(new_n228_) );
  NAND2_X1 g0092 ( .A1(new_n141_), .A2(new_n228_), .ZN(new_n229_) );
  NAND2_X1 g0093 ( .A1(new_n227_), .A2(new_n229_), .ZN(new_n230_) );
  NAND4_X1 g0094 ( .A1(new_n138_), .A2(new_n141_), .A3(new_n226_), .A4(new_n228_), .ZN(new_n231_) );
  NAND2_X1 g0095 ( .A1(new_n230_), .A2(new_n231_), .ZN(new_n232_) );
  NAND2_X1 g0096 ( .A1(new_n225_), .A2(new_n232_), .ZN(new_n233_) );
  NAND4_X1 g0097 ( .A1(new_n223_), .A2(new_n224_), .A3(new_n230_), .A4(new_n231_), .ZN(new_n234_) );
  NAND2_X1 g0098 ( .A1(new_n233_), .A2(new_n234_), .ZN(G351) );
  INV_X1 g0099 ( .A(KEYINPUT4), .ZN(new_n236_) );
  NAND4_X1 g0100 ( .A1(G1), .A2(G20), .A3(G33), .A4(KEYINPUT3), .ZN(new_n237_) );
  INV_X1 g0101 ( .A(KEYINPUT3), .ZN(new_n238_) );
  NAND3_X1 g0102 ( .A1(G1), .A2(G20), .A3(G33), .ZN(new_n239_) );
  NAND2_X1 g0103 ( .A1(new_n239_), .A2(new_n238_), .ZN(new_n240_) );
  NAND2_X1 g0104 ( .A1(new_n240_), .A2(new_n237_), .ZN(new_n241_) );
  NAND3_X1 g0105 ( .A1(new_n241_), .A2(new_n169_), .A3(new_n170_), .ZN(new_n242_) );
  NAND3_X1 g0106 ( .A1(new_n242_), .A2(G20), .A3(new_n236_), .ZN(new_n243_) );
  NAND2_X1 g0107 ( .A1(new_n242_), .A2(G20), .ZN(new_n244_) );
  NAND2_X1 g0108 ( .A1(new_n244_), .A2(KEYINPUT4), .ZN(new_n245_) );
  NAND2_X1 g0109 ( .A1(new_n245_), .A2(new_n243_), .ZN(new_n246_) );
  INV_X1 g0110 ( .A(new_n246_), .ZN(new_n247_) );
  NAND2_X1 g0111 ( .A1(new_n247_), .A2(new_n227_), .ZN(new_n248_) );
  INV_X1 g0112 ( .A(new_n242_), .ZN(new_n249_) );
  INV_X1 g0113 ( .A(G1), .ZN(new_n250_) );
  NAND2_X1 g0114 ( .A1(new_n250_), .A2(G20), .ZN(new_n251_) );
  NAND3_X1 g0115 ( .A1(new_n249_), .A2(G58), .A3(new_n251_), .ZN(new_n252_) );
  INV_X1 g0116 ( .A(new_n252_), .ZN(new_n253_) );
  INV_X1 g0117 ( .A(G20), .ZN(new_n254_) );
  INV_X1 g0118 ( .A(G33), .ZN(new_n255_) );
  NAND2_X1 g0119 ( .A1(new_n171_), .A2(new_n255_), .ZN(new_n256_) );
  INV_X1 g0120 ( .A(new_n256_), .ZN(new_n257_) );
  NAND2_X1 g0121 ( .A1(new_n257_), .A2(new_n254_), .ZN(new_n258_) );
  INV_X1 g0122 ( .A(new_n258_), .ZN(new_n259_) );
  NAND2_X1 g0123 ( .A1(new_n259_), .A2(G159), .ZN(new_n260_) );
  NOR2_X1 g0124 ( .A1(new_n255_), .A2(G20), .ZN(new_n261_) );
  NAND2_X1 g0125 ( .A1(new_n171_), .A2(new_n261_), .ZN(new_n262_) );
  INV_X1 g0126 ( .A(new_n262_), .ZN(new_n263_) );
  NAND2_X1 g0127 ( .A1(new_n263_), .A2(G68), .ZN(new_n264_) );
  INV_X1 g0128 ( .A(G58), .ZN(new_n265_) );
  NAND3_X1 g0129 ( .A1(new_n250_), .A2(G13), .A3(G20), .ZN(new_n266_) );
  INV_X1 g0130 ( .A(new_n266_), .ZN(new_n267_) );
  NAND2_X1 g0131 ( .A1(new_n267_), .A2(new_n265_), .ZN(new_n268_) );
  NAND3_X1 g0132 ( .A1(new_n260_), .A2(new_n264_), .A3(new_n268_), .ZN(new_n269_) );
  NOR2_X1 g0133 ( .A1(new_n269_), .A2(new_n253_), .ZN(new_n270_) );
  NAND2_X1 g0134 ( .A1(new_n270_), .A2(new_n248_), .ZN(new_n271_) );
  NAND2_X1 g0135 ( .A1(new_n271_), .A2(KEYINPUT30), .ZN(new_n272_) );
  INV_X1 g0136 ( .A(KEYINPUT30), .ZN(new_n273_) );
  NAND3_X1 g0137 ( .A1(new_n270_), .A2(new_n248_), .A3(new_n273_), .ZN(new_n274_) );
  NAND2_X1 g0138 ( .A1(new_n272_), .A2(new_n274_), .ZN(new_n275_) );
  INV_X1 g0139 ( .A(KEYINPUT32), .ZN(new_n276_) );
  NAND4_X1 g0140 ( .A1(new_n257_), .A2(G226), .A3(G1698), .A4(new_n276_), .ZN(new_n277_) );
  NAND3_X1 g0141 ( .A1(new_n257_), .A2(G226), .A3(G1698), .ZN(new_n278_) );
  NAND2_X1 g0142 ( .A1(new_n278_), .A2(KEYINPUT32), .ZN(new_n279_) );
  NAND2_X1 g0143 ( .A1(new_n279_), .A2(new_n277_), .ZN(new_n280_) );
  INV_X1 g0144 ( .A(G1698), .ZN(new_n281_) );
  NAND2_X1 g0145 ( .A1(new_n257_), .A2(new_n281_), .ZN(new_n282_) );
  INV_X1 g0146 ( .A(new_n282_), .ZN(new_n283_) );
  NAND2_X1 g0147 ( .A1(new_n283_), .A2(G223), .ZN(new_n284_) );
  NAND2_X1 g0148 ( .A1(new_n280_), .A2(new_n284_), .ZN(new_n285_) );
  NAND2_X1 g0149 ( .A1(new_n285_), .A2(KEYINPUT33), .ZN(new_n286_) );
  INV_X1 g0150 ( .A(KEYINPUT33), .ZN(new_n287_) );
  NAND3_X1 g0151 ( .A1(new_n280_), .A2(new_n287_), .A3(new_n284_), .ZN(new_n288_) );
  NAND2_X1 g0152 ( .A1(new_n286_), .A2(new_n288_), .ZN(new_n289_) );
  INV_X1 g0153 ( .A(G41), .ZN(new_n290_) );
  INV_X1 g0154 ( .A(G45), .ZN(new_n291_) );
  NAND2_X1 g0155 ( .A1(new_n290_), .A2(new_n291_), .ZN(new_n292_) );
  NAND3_X1 g0156 ( .A1(new_n292_), .A2(new_n250_), .A3(G274), .ZN(new_n293_) );
  NOR2_X1 g0157 ( .A1(new_n255_), .A2(G41), .ZN(new_n294_) );
  NAND2_X1 g0158 ( .A1(new_n171_), .A2(new_n294_), .ZN(new_n295_) );
  INV_X1 g0159 ( .A(new_n295_), .ZN(new_n296_) );
  NAND2_X1 g0160 ( .A1(new_n296_), .A2(G87), .ZN(new_n297_) );
  NAND2_X1 g0161 ( .A1(new_n297_), .A2(KEYINPUT31), .ZN(new_n298_) );
  INV_X1 g0162 ( .A(KEYINPUT31), .ZN(new_n299_) );
  NAND3_X1 g0163 ( .A1(new_n296_), .A2(G87), .A3(new_n299_), .ZN(new_n300_) );
  NAND2_X1 g0164 ( .A1(new_n292_), .A2(new_n250_), .ZN(new_n301_) );
  NAND2_X1 g0165 ( .A1(G33), .A2(G41), .ZN(new_n302_) );
  NAND2_X1 g0166 ( .A1(new_n171_), .A2(new_n302_), .ZN(new_n303_) );
  NAND2_X1 g0167 ( .A1(new_n303_), .A2(new_n301_), .ZN(new_n304_) );
  INV_X1 g0168 ( .A(new_n304_), .ZN(new_n305_) );
  NAND2_X1 g0169 ( .A1(new_n305_), .A2(G232), .ZN(new_n306_) );
  NAND4_X1 g0170 ( .A1(new_n298_), .A2(new_n306_), .A3(new_n293_), .A4(new_n300_), .ZN(new_n307_) );
  INV_X1 g0171 ( .A(new_n307_), .ZN(new_n308_) );
  NAND3_X1 g0172 ( .A1(new_n289_), .A2(G179), .A3(new_n308_), .ZN(new_n309_) );
  NAND2_X1 g0173 ( .A1(new_n309_), .A2(KEYINPUT34), .ZN(new_n310_) );
  INV_X1 g0174 ( .A(KEYINPUT34), .ZN(new_n311_) );
  NAND4_X1 g0175 ( .A1(new_n289_), .A2(G179), .A3(new_n311_), .A4(new_n308_), .ZN(new_n312_) );
  NAND2_X1 g0176 ( .A1(new_n310_), .A2(new_n312_), .ZN(new_n313_) );
  NAND2_X1 g0177 ( .A1(new_n289_), .A2(new_n308_), .ZN(new_n314_) );
  NAND2_X1 g0178 ( .A1(new_n314_), .A2(G169), .ZN(new_n315_) );
  NAND2_X1 g0179 ( .A1(new_n313_), .A2(new_n315_), .ZN(new_n316_) );
  NAND2_X1 g0180 ( .A1(new_n316_), .A2(new_n275_), .ZN(new_n317_) );
  INV_X1 g0181 ( .A(new_n317_), .ZN(new_n318_) );
  NAND4_X1 g0182 ( .A1(new_n171_), .A2(new_n255_), .A3(G238), .A4(G1698), .ZN(new_n319_) );
  INV_X1 g0183 ( .A(new_n319_), .ZN(new_n320_) );
  NAND2_X1 g0184 ( .A1(new_n320_), .A2(KEYINPUT6), .ZN(new_n321_) );
  INV_X1 g0185 ( .A(KEYINPUT6), .ZN(new_n322_) );
  NAND2_X1 g0186 ( .A1(new_n319_), .A2(new_n322_), .ZN(new_n323_) );
  NAND3_X1 g0187 ( .A1(new_n257_), .A2(G232), .A3(new_n281_), .ZN(new_n324_) );
  NAND3_X1 g0188 ( .A1(new_n171_), .A2(G107), .A3(new_n294_), .ZN(new_n325_) );
  NAND2_X1 g0189 ( .A1(new_n325_), .A2(new_n293_), .ZN(new_n326_) );
  INV_X1 g0190 ( .A(new_n326_), .ZN(new_n327_) );
  NAND4_X1 g0191 ( .A1(new_n321_), .A2(new_n324_), .A3(new_n327_), .A4(new_n323_), .ZN(new_n328_) );
  NAND2_X1 g0192 ( .A1(new_n328_), .A2(KEYINPUT7), .ZN(new_n329_) );
  INV_X1 g0193 ( .A(KEYINPUT7), .ZN(new_n330_) );
  NAND2_X1 g0194 ( .A1(new_n324_), .A2(new_n327_), .ZN(new_n331_) );
  INV_X1 g0195 ( .A(new_n331_), .ZN(new_n332_) );
  NAND4_X1 g0196 ( .A1(new_n332_), .A2(new_n330_), .A3(new_n321_), .A4(new_n323_), .ZN(new_n333_) );
  NAND2_X1 g0197 ( .A1(new_n333_), .A2(new_n329_), .ZN(new_n334_) );
  NAND2_X1 g0198 ( .A1(new_n305_), .A2(G244), .ZN(new_n335_) );
  NAND3_X1 g0199 ( .A1(new_n334_), .A2(G179), .A3(new_n335_), .ZN(new_n336_) );
  NAND2_X1 g0200 ( .A1(new_n334_), .A2(new_n335_), .ZN(new_n337_) );
  NAND2_X1 g0201 ( .A1(new_n337_), .A2(G169), .ZN(new_n338_) );
  NAND2_X1 g0202 ( .A1(new_n338_), .A2(new_n336_), .ZN(new_n339_) );
  NAND2_X1 g0203 ( .A1(new_n249_), .A2(new_n251_), .ZN(new_n340_) );
  NAND2_X1 g0204 ( .A1(new_n246_), .A2(new_n340_), .ZN(new_n341_) );
  NAND2_X1 g0205 ( .A1(new_n341_), .A2(G77), .ZN(new_n342_) );
  NAND2_X1 g0206 ( .A1(new_n259_), .A2(G58), .ZN(new_n343_) );
  NAND2_X1 g0207 ( .A1(new_n263_), .A2(G87), .ZN(new_n344_) );
  NAND2_X1 g0208 ( .A1(new_n267_), .A2(new_n140_), .ZN(new_n345_) );
  NAND3_X1 g0209 ( .A1(new_n343_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_) );
  INV_X1 g0210 ( .A(new_n346_), .ZN(new_n347_) );
  NAND2_X1 g0211 ( .A1(new_n342_), .A2(new_n347_), .ZN(new_n348_) );
  NAND2_X1 g0212 ( .A1(new_n339_), .A2(new_n348_), .ZN(new_n349_) );
  NAND2_X1 g0213 ( .A1(new_n337_), .A2(G200), .ZN(new_n350_) );
  NAND3_X1 g0214 ( .A1(new_n334_), .A2(G190), .A3(new_n335_), .ZN(new_n351_) );
  NAND4_X1 g0215 ( .A1(new_n350_), .A2(new_n342_), .A3(new_n347_), .A4(new_n351_), .ZN(new_n352_) );
  NAND2_X1 g0216 ( .A1(new_n349_), .A2(new_n352_), .ZN(new_n353_) );
  INV_X1 g0217 ( .A(new_n353_), .ZN(new_n354_) );
  INV_X1 g0218 ( .A(KEYINPUT35), .ZN(new_n355_) );
  NAND2_X1 g0219 ( .A1(new_n314_), .A2(G200), .ZN(new_n356_) );
  NAND2_X1 g0220 ( .A1(new_n356_), .A2(new_n355_), .ZN(new_n357_) );
  NAND3_X1 g0221 ( .A1(new_n314_), .A2(G200), .A3(KEYINPUT35), .ZN(new_n358_) );
  NAND2_X1 g0222 ( .A1(new_n357_), .A2(new_n358_), .ZN(new_n359_) );
  NAND3_X1 g0223 ( .A1(new_n289_), .A2(G190), .A3(new_n308_), .ZN(new_n360_) );
  NAND4_X1 g0224 ( .A1(new_n359_), .A2(new_n272_), .A3(new_n274_), .A4(new_n360_), .ZN(new_n361_) );
  NAND2_X1 g0225 ( .A1(new_n341_), .A2(G50), .ZN(new_n362_) );
  NAND2_X1 g0226 ( .A1(new_n247_), .A2(new_n138_), .ZN(new_n363_) );
  NAND2_X1 g0227 ( .A1(new_n259_), .A2(G150), .ZN(new_n364_) );
  NAND2_X1 g0228 ( .A1(new_n263_), .A2(G58), .ZN(new_n365_) );
  NAND2_X1 g0229 ( .A1(new_n267_), .A2(new_n139_), .ZN(new_n366_) );
  NAND4_X1 g0230 ( .A1(new_n363_), .A2(new_n364_), .A3(new_n365_), .A4(new_n366_), .ZN(new_n367_) );
  INV_X1 g0231 ( .A(new_n367_), .ZN(new_n368_) );
  NAND2_X1 g0232 ( .A1(new_n368_), .A2(new_n362_), .ZN(new_n369_) );
  INV_X1 g0233 ( .A(G179), .ZN(new_n370_) );
  NAND2_X1 g0234 ( .A1(new_n283_), .A2(G222), .ZN(new_n371_) );
  NAND2_X1 g0235 ( .A1(new_n371_), .A2(KEYINPUT36), .ZN(new_n372_) );
  INV_X1 g0236 ( .A(KEYINPUT36), .ZN(new_n373_) );
  NAND3_X1 g0237 ( .A1(new_n283_), .A2(G222), .A3(new_n373_), .ZN(new_n374_) );
  NAND2_X1 g0238 ( .A1(new_n372_), .A2(new_n374_), .ZN(new_n375_) );
  NAND2_X1 g0239 ( .A1(new_n305_), .A2(G226), .ZN(new_n376_) );
  INV_X1 g0240 ( .A(new_n376_), .ZN(new_n377_) );
  NAND3_X1 g0241 ( .A1(new_n257_), .A2(G223), .A3(G1698), .ZN(new_n378_) );
  NAND2_X1 g0242 ( .A1(new_n296_), .A2(G77), .ZN(new_n379_) );
  NAND3_X1 g0243 ( .A1(new_n378_), .A2(new_n293_), .A3(new_n379_), .ZN(new_n380_) );
  NOR2_X1 g0244 ( .A1(new_n377_), .A2(new_n380_), .ZN(new_n381_) );
  NAND2_X1 g0245 ( .A1(new_n375_), .A2(new_n381_), .ZN(new_n382_) );
  INV_X1 g0246 ( .A(new_n382_), .ZN(new_n383_) );
  NAND2_X1 g0247 ( .A1(new_n383_), .A2(new_n370_), .ZN(new_n384_) );
  INV_X1 g0248 ( .A(G169), .ZN(new_n385_) );
  NAND2_X1 g0249 ( .A1(new_n382_), .A2(new_n385_), .ZN(new_n386_) );
  NAND3_X1 g0250 ( .A1(new_n369_), .A2(new_n384_), .A3(new_n386_), .ZN(new_n387_) );
  NAND2_X1 g0251 ( .A1(new_n383_), .A2(G190), .ZN(new_n388_) );
  NAND2_X1 g0252 ( .A1(new_n382_), .A2(G200), .ZN(new_n389_) );
  NAND4_X1 g0253 ( .A1(new_n388_), .A2(new_n362_), .A3(new_n368_), .A4(new_n389_), .ZN(new_n390_) );
  NAND2_X1 g0254 ( .A1(new_n387_), .A2(new_n390_), .ZN(new_n391_) );
  NAND2_X1 g0255 ( .A1(new_n391_), .A2(KEYINPUT37), .ZN(new_n392_) );
  INV_X1 g0256 ( .A(KEYINPUT37), .ZN(new_n393_) );
  NAND3_X1 g0257 ( .A1(new_n387_), .A2(new_n390_), .A3(new_n393_), .ZN(new_n394_) );
  NAND2_X1 g0258 ( .A1(new_n392_), .A2(new_n394_), .ZN(new_n395_) );
  NAND3_X1 g0259 ( .A1(new_n303_), .A2(G238), .A3(new_n301_), .ZN(new_n396_) );
  INV_X1 g0260 ( .A(new_n396_), .ZN(new_n397_) );
  NAND3_X1 g0261 ( .A1(new_n171_), .A2(G97), .A3(new_n294_), .ZN(new_n398_) );
  NAND2_X1 g0262 ( .A1(new_n398_), .A2(new_n293_), .ZN(new_n399_) );
  NAND4_X1 g0263 ( .A1(new_n171_), .A2(new_n255_), .A3(G232), .A4(G1698), .ZN(new_n400_) );
  NAND4_X1 g0264 ( .A1(new_n171_), .A2(new_n255_), .A3(G226), .A4(new_n281_), .ZN(new_n401_) );
  NAND2_X1 g0265 ( .A1(new_n400_), .A2(new_n401_), .ZN(new_n402_) );
  NOR3_X1 g0266 ( .A1(new_n397_), .A2(new_n402_), .A3(new_n399_), .ZN(new_n403_) );
  NAND2_X1 g0267 ( .A1(new_n403_), .A2(G190), .ZN(new_n404_) );
  NAND2_X1 g0268 ( .A1(new_n404_), .A2(KEYINPUT28), .ZN(new_n405_) );
  INV_X1 g0269 ( .A(KEYINPUT28), .ZN(new_n406_) );
  NAND3_X1 g0270 ( .A1(new_n403_), .A2(G190), .A3(new_n406_), .ZN(new_n407_) );
  NAND2_X1 g0271 ( .A1(new_n405_), .A2(new_n407_), .ZN(new_n408_) );
  INV_X1 g0272 ( .A(G68), .ZN(new_n409_) );
  NAND2_X1 g0273 ( .A1(new_n246_), .A2(new_n266_), .ZN(new_n410_) );
  NAND2_X1 g0274 ( .A1(new_n410_), .A2(new_n409_), .ZN(new_n411_) );
  NAND3_X1 g0275 ( .A1(new_n249_), .A2(G68), .A3(new_n251_), .ZN(new_n412_) );
  INV_X1 g0276 ( .A(new_n412_), .ZN(new_n413_) );
  NAND2_X1 g0277 ( .A1(new_n259_), .A2(G50), .ZN(new_n414_) );
  NAND2_X1 g0278 ( .A1(new_n263_), .A2(G77), .ZN(new_n415_) );
  NAND2_X1 g0279 ( .A1(new_n414_), .A2(new_n415_), .ZN(new_n416_) );
  NOR2_X1 g0280 ( .A1(new_n416_), .A2(new_n413_), .ZN(new_n417_) );
  INV_X1 g0281 ( .A(new_n399_), .ZN(new_n418_) );
  NAND4_X1 g0282 ( .A1(new_n418_), .A2(new_n396_), .A3(new_n400_), .A4(new_n401_), .ZN(new_n419_) );
  NAND2_X1 g0283 ( .A1(new_n419_), .A2(G200), .ZN(new_n420_) );
  NAND2_X1 g0284 ( .A1(new_n420_), .A2(KEYINPUT27), .ZN(new_n421_) );
  INV_X1 g0285 ( .A(KEYINPUT27), .ZN(new_n422_) );
  NAND3_X1 g0286 ( .A1(new_n419_), .A2(G200), .A3(new_n422_), .ZN(new_n423_) );
  NAND2_X1 g0287 ( .A1(new_n421_), .A2(new_n423_), .ZN(new_n424_) );
  INV_X1 g0288 ( .A(new_n424_), .ZN(new_n425_) );
  NAND4_X1 g0289 ( .A1(new_n425_), .A2(new_n408_), .A3(new_n411_), .A4(new_n417_), .ZN(new_n426_) );
  INV_X1 g0290 ( .A(new_n426_), .ZN(new_n427_) );
  NAND2_X1 g0291 ( .A1(new_n417_), .A2(new_n411_), .ZN(new_n428_) );
  NOR2_X1 g0292 ( .A1(new_n419_), .A2(G179), .ZN(new_n429_) );
  NOR2_X1 g0293 ( .A1(new_n403_), .A2(G169), .ZN(new_n430_) );
  NOR2_X1 g0294 ( .A1(new_n430_), .A2(new_n429_), .ZN(new_n431_) );
  NAND2_X1 g0295 ( .A1(new_n428_), .A2(new_n431_), .ZN(new_n432_) );
  INV_X1 g0296 ( .A(new_n432_), .ZN(new_n433_) );
  NOR2_X1 g0297 ( .A1(new_n427_), .A2(new_n433_), .ZN(new_n434_) );
  NAND4_X1 g0298 ( .A1(new_n395_), .A2(new_n354_), .A3(new_n361_), .A4(new_n434_), .ZN(new_n435_) );
  NOR2_X1 g0299 ( .A1(new_n435_), .A2(new_n318_), .ZN(new_n436_) );
  INV_X1 g0300 ( .A(new_n436_), .ZN(new_n437_) );
  INV_X1 g0301 ( .A(KEYINPUT0), .ZN(new_n438_) );
  INV_X1 g0302 ( .A(G107), .ZN(new_n439_) );
  NAND2_X1 g0303 ( .A1(new_n410_), .A2(new_n439_), .ZN(new_n440_) );
  INV_X1 g0304 ( .A(KEYINPUT16), .ZN(new_n441_) );
  NAND4_X1 g0305 ( .A1(new_n171_), .A2(G116), .A3(new_n441_), .A4(new_n261_), .ZN(new_n442_) );
  NAND3_X1 g0306 ( .A1(new_n171_), .A2(G116), .A3(new_n261_), .ZN(new_n443_) );
  NAND2_X1 g0307 ( .A1(new_n443_), .A2(KEYINPUT16), .ZN(new_n444_) );
  NAND2_X1 g0308 ( .A1(new_n444_), .A2(new_n442_), .ZN(new_n445_) );
  INV_X1 g0309 ( .A(new_n171_), .ZN(new_n446_) );
  NAND2_X1 g0310 ( .A1(new_n250_), .A2(G33), .ZN(new_n447_) );
  NAND2_X1 g0311 ( .A1(new_n266_), .A2(new_n447_), .ZN(new_n448_) );
  INV_X1 g0312 ( .A(new_n448_), .ZN(new_n449_) );
  NAND4_X1 g0313 ( .A1(new_n446_), .A2(new_n449_), .A3(G107), .A4(new_n241_), .ZN(new_n450_) );
  NAND3_X1 g0314 ( .A1(new_n445_), .A2(KEYINPUT17), .A3(new_n450_), .ZN(new_n451_) );
  INV_X1 g0315 ( .A(KEYINPUT17), .ZN(new_n452_) );
  NAND2_X1 g0316 ( .A1(new_n445_), .A2(new_n450_), .ZN(new_n453_) );
  NAND2_X1 g0317 ( .A1(new_n453_), .A2(new_n452_), .ZN(new_n454_) );
  NAND2_X1 g0318 ( .A1(new_n259_), .A2(G87), .ZN(new_n455_) );
  NAND4_X1 g0319 ( .A1(new_n440_), .A2(new_n451_), .A3(new_n454_), .A4(new_n455_), .ZN(new_n456_) );
  INV_X1 g0320 ( .A(KEYINPUT15), .ZN(new_n457_) );
  NOR3_X1 g0321 ( .A1(new_n291_), .A2(G1), .A3(G41), .ZN(new_n458_) );
  NAND2_X1 g0322 ( .A1(new_n458_), .A2(G274), .ZN(new_n459_) );
  INV_X1 g0323 ( .A(KEYINPUT14), .ZN(new_n460_) );
  NAND3_X1 g0324 ( .A1(new_n290_), .A2(G33), .A3(G294), .ZN(new_n461_) );
  INV_X1 g0325 ( .A(new_n461_), .ZN(new_n462_) );
  NAND2_X1 g0326 ( .A1(new_n171_), .A2(new_n462_), .ZN(new_n463_) );
  NAND2_X1 g0327 ( .A1(new_n463_), .A2(new_n460_), .ZN(new_n464_) );
  NAND3_X1 g0328 ( .A1(new_n171_), .A2(KEYINPUT14), .A3(new_n462_), .ZN(new_n465_) );
  NOR2_X1 g0329 ( .A1(new_n458_), .A2(new_n178_), .ZN(new_n466_) );
  NAND2_X1 g0330 ( .A1(new_n303_), .A2(new_n466_), .ZN(new_n467_) );
  NAND4_X1 g0331 ( .A1(new_n464_), .A2(new_n467_), .A3(new_n459_), .A4(new_n465_), .ZN(new_n468_) );
  NAND4_X1 g0332 ( .A1(new_n171_), .A2(new_n255_), .A3(G250), .A4(new_n281_), .ZN(new_n469_) );
  NAND4_X1 g0333 ( .A1(new_n171_), .A2(new_n255_), .A3(G257), .A4(G1698), .ZN(new_n470_) );
  NAND2_X1 g0334 ( .A1(new_n469_), .A2(new_n470_), .ZN(new_n471_) );
  NOR3_X1 g0335 ( .A1(new_n468_), .A2(G179), .A3(new_n471_), .ZN(new_n472_) );
  NOR2_X1 g0336 ( .A1(new_n472_), .A2(new_n457_), .ZN(new_n473_) );
  NOR4_X1 g0337 ( .A1(new_n468_), .A2(G179), .A3(KEYINPUT15), .A4(new_n471_), .ZN(new_n474_) );
  NOR2_X1 g0338 ( .A1(new_n468_), .A2(new_n471_), .ZN(new_n475_) );
  NOR2_X1 g0339 ( .A1(new_n475_), .A2(G169), .ZN(new_n476_) );
  NOR3_X1 g0340 ( .A1(new_n473_), .A2(new_n476_), .A3(new_n474_), .ZN(new_n477_) );
  NAND2_X1 g0341 ( .A1(new_n477_), .A2(new_n456_), .ZN(new_n478_) );
  NAND3_X1 g0342 ( .A1(new_n454_), .A2(new_n451_), .A3(new_n455_), .ZN(new_n479_) );
  INV_X1 g0343 ( .A(new_n479_), .ZN(new_n480_) );
  INV_X1 g0344 ( .A(new_n475_), .ZN(new_n481_) );
  NAND2_X1 g0345 ( .A1(new_n481_), .A2(G200), .ZN(new_n482_) );
  NAND2_X1 g0346 ( .A1(new_n475_), .A2(G190), .ZN(new_n483_) );
  NAND4_X1 g0347 ( .A1(new_n480_), .A2(new_n440_), .A3(new_n482_), .A4(new_n483_), .ZN(new_n484_) );
  NAND2_X1 g0348 ( .A1(new_n478_), .A2(new_n484_), .ZN(new_n485_) );
  NAND2_X1 g0349 ( .A1(new_n485_), .A2(new_n438_), .ZN(new_n486_) );
  NAND3_X1 g0350 ( .A1(new_n478_), .A2(KEYINPUT0), .A3(new_n484_), .ZN(new_n487_) );
  NAND2_X1 g0351 ( .A1(new_n486_), .A2(new_n487_), .ZN(new_n488_) );
  NAND2_X1 g0352 ( .A1(new_n283_), .A2(G244), .ZN(new_n489_) );
  NAND3_X1 g0353 ( .A1(new_n257_), .A2(G250), .A3(G1698), .ZN(new_n490_) );
  NAND2_X1 g0354 ( .A1(new_n296_), .A2(G283), .ZN(new_n491_) );
  NAND2_X1 g0355 ( .A1(new_n491_), .A2(new_n459_), .ZN(new_n492_) );
  INV_X1 g0356 ( .A(new_n492_), .ZN(new_n493_) );
  NAND4_X1 g0357 ( .A1(new_n489_), .A2(new_n493_), .A3(KEYINPUT12), .A4(new_n490_), .ZN(new_n494_) );
  INV_X1 g0358 ( .A(KEYINPUT12), .ZN(new_n495_) );
  NAND3_X1 g0359 ( .A1(new_n489_), .A2(new_n493_), .A3(new_n490_), .ZN(new_n496_) );
  NAND2_X1 g0360 ( .A1(new_n496_), .A2(new_n495_), .ZN(new_n497_) );
  NAND2_X1 g0361 ( .A1(new_n497_), .A2(new_n494_), .ZN(new_n498_) );
  INV_X1 g0362 ( .A(new_n458_), .ZN(new_n499_) );
  NAND3_X1 g0363 ( .A1(new_n303_), .A2(G257), .A3(new_n499_), .ZN(new_n500_) );
  NAND2_X1 g0364 ( .A1(new_n498_), .A2(new_n500_), .ZN(new_n501_) );
  NAND2_X1 g0365 ( .A1(new_n501_), .A2(new_n385_), .ZN(new_n502_) );
  NAND3_X1 g0366 ( .A1(new_n498_), .A2(new_n370_), .A3(new_n500_), .ZN(new_n503_) );
  NAND2_X1 g0367 ( .A1(new_n247_), .A2(new_n212_), .ZN(new_n504_) );
  NAND2_X1 g0368 ( .A1(new_n263_), .A2(G107), .ZN(new_n505_) );
  INV_X1 g0369 ( .A(G97), .ZN(new_n506_) );
  NAND2_X1 g0370 ( .A1(new_n267_), .A2(new_n506_), .ZN(new_n507_) );
  NAND3_X1 g0371 ( .A1(new_n505_), .A2(KEYINPUT13), .A3(new_n507_), .ZN(new_n508_) );
  NAND2_X1 g0372 ( .A1(new_n259_), .A2(G77), .ZN(new_n509_) );
  NAND2_X1 g0373 ( .A1(new_n509_), .A2(new_n508_), .ZN(new_n510_) );
  INV_X1 g0374 ( .A(KEYINPUT13), .ZN(new_n511_) );
  NAND2_X1 g0375 ( .A1(new_n505_), .A2(new_n507_), .ZN(new_n512_) );
  NAND2_X1 g0376 ( .A1(new_n512_), .A2(new_n511_), .ZN(new_n513_) );
  NOR2_X1 g0377 ( .A1(new_n242_), .A2(new_n448_), .ZN(new_n514_) );
  NAND2_X1 g0378 ( .A1(new_n514_), .A2(G97), .ZN(new_n515_) );
  NAND2_X1 g0379 ( .A1(new_n513_), .A2(new_n515_), .ZN(new_n516_) );
  NOR2_X1 g0380 ( .A1(new_n516_), .A2(new_n510_), .ZN(new_n517_) );
  NAND2_X1 g0381 ( .A1(new_n517_), .A2(new_n504_), .ZN(new_n518_) );
  NAND3_X1 g0382 ( .A1(new_n502_), .A2(new_n503_), .A3(new_n518_), .ZN(new_n519_) );
  NAND3_X1 g0383 ( .A1(new_n498_), .A2(G190), .A3(new_n500_), .ZN(new_n520_) );
  NAND2_X1 g0384 ( .A1(new_n501_), .A2(G200), .ZN(new_n521_) );
  NAND4_X1 g0385 ( .A1(new_n521_), .A2(new_n504_), .A3(new_n517_), .A4(new_n520_), .ZN(new_n522_) );
  NAND2_X1 g0386 ( .A1(new_n522_), .A2(new_n519_), .ZN(new_n523_) );
  INV_X1 g0387 ( .A(new_n523_), .ZN(new_n524_) );
  INV_X1 g0388 ( .A(new_n514_), .ZN(new_n525_) );
  NAND2_X1 g0389 ( .A1(new_n246_), .A2(new_n525_), .ZN(new_n526_) );
  NAND2_X1 g0390 ( .A1(new_n526_), .A2(G116), .ZN(new_n527_) );
  NAND2_X1 g0391 ( .A1(new_n259_), .A2(G97), .ZN(new_n528_) );
  NAND2_X1 g0392 ( .A1(new_n263_), .A2(G283), .ZN(new_n529_) );
  NAND2_X1 g0393 ( .A1(new_n267_), .A2(new_n219_), .ZN(new_n530_) );
  NAND3_X1 g0394 ( .A1(new_n528_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_) );
  INV_X1 g0395 ( .A(new_n531_), .ZN(new_n532_) );
  NAND2_X1 g0396 ( .A1(new_n527_), .A2(new_n532_), .ZN(new_n533_) );
  NAND4_X1 g0397 ( .A1(new_n171_), .A2(new_n255_), .A3(G257), .A4(new_n281_), .ZN(new_n534_) );
  NAND3_X1 g0398 ( .A1(new_n171_), .A2(G303), .A3(new_n294_), .ZN(new_n535_) );
  NAND3_X1 g0399 ( .A1(new_n534_), .A2(new_n459_), .A3(new_n535_), .ZN(new_n536_) );
  INV_X1 g0400 ( .A(new_n536_), .ZN(new_n537_) );
  INV_X1 g0401 ( .A(KEYINPUT10), .ZN(new_n538_) );
  NAND3_X1 g0402 ( .A1(new_n303_), .A2(G270), .A3(new_n499_), .ZN(new_n539_) );
  NAND2_X1 g0403 ( .A1(new_n539_), .A2(new_n538_), .ZN(new_n540_) );
  NAND3_X1 g0404 ( .A1(new_n257_), .A2(G264), .A3(G1698), .ZN(new_n541_) );
  NAND4_X1 g0405 ( .A1(new_n303_), .A2(G270), .A3(KEYINPUT10), .A4(new_n499_), .ZN(new_n542_) );
  NAND2_X1 g0406 ( .A1(new_n541_), .A2(new_n542_), .ZN(new_n543_) );
  INV_X1 g0407 ( .A(new_n543_), .ZN(new_n544_) );
  NAND4_X1 g0408 ( .A1(new_n544_), .A2(G179), .A3(new_n537_), .A4(new_n540_), .ZN(new_n545_) );
  NAND4_X1 g0409 ( .A1(new_n537_), .A2(new_n540_), .A3(new_n541_), .A4(new_n542_), .ZN(new_n546_) );
  NAND2_X1 g0410 ( .A1(new_n546_), .A2(G169), .ZN(new_n547_) );
  NAND2_X1 g0411 ( .A1(new_n545_), .A2(new_n547_), .ZN(new_n548_) );
  NAND2_X1 g0412 ( .A1(new_n533_), .A2(new_n548_), .ZN(new_n549_) );
  NAND4_X1 g0413 ( .A1(new_n544_), .A2(G190), .A3(new_n537_), .A4(new_n540_), .ZN(new_n550_) );
  NAND2_X1 g0414 ( .A1(new_n546_), .A2(G200), .ZN(new_n551_) );
  NAND4_X1 g0415 ( .A1(new_n527_), .A2(new_n532_), .A3(new_n550_), .A4(new_n551_), .ZN(new_n552_) );
  NAND2_X1 g0416 ( .A1(new_n549_), .A2(new_n552_), .ZN(new_n553_) );
  NAND2_X1 g0417 ( .A1(new_n553_), .A2(KEYINPUT11), .ZN(new_n554_) );
  INV_X1 g0418 ( .A(KEYINPUT11), .ZN(new_n555_) );
  NAND3_X1 g0419 ( .A1(new_n549_), .A2(new_n555_), .A3(new_n552_), .ZN(new_n556_) );
  NAND2_X1 g0420 ( .A1(new_n554_), .A2(new_n556_), .ZN(new_n557_) );
  INV_X1 g0421 ( .A(KEYINPUT9), .ZN(new_n558_) );
  NAND2_X1 g0422 ( .A1(new_n514_), .A2(G87), .ZN(new_n559_) );
  NAND2_X1 g0423 ( .A1(new_n246_), .A2(new_n559_), .ZN(new_n560_) );
  NAND2_X1 g0424 ( .A1(new_n143_), .A2(new_n217_), .ZN(new_n561_) );
  NAND3_X1 g0425 ( .A1(new_n560_), .A2(new_n558_), .A3(new_n561_), .ZN(new_n562_) );
  NAND2_X1 g0426 ( .A1(new_n560_), .A2(new_n561_), .ZN(new_n563_) );
  NAND2_X1 g0427 ( .A1(new_n563_), .A2(KEYINPUT9), .ZN(new_n564_) );
  NAND2_X1 g0428 ( .A1(new_n259_), .A2(G68), .ZN(new_n565_) );
  NAND2_X1 g0429 ( .A1(new_n263_), .A2(G97), .ZN(new_n566_) );
  NAND2_X1 g0430 ( .A1(new_n267_), .A2(new_n217_), .ZN(new_n567_) );
  NAND3_X1 g0431 ( .A1(new_n565_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_) );
  INV_X1 g0432 ( .A(new_n568_), .ZN(new_n569_) );
  NAND3_X1 g0433 ( .A1(new_n564_), .A2(new_n562_), .A3(new_n569_), .ZN(new_n570_) );
  NAND4_X1 g0434 ( .A1(new_n171_), .A2(new_n255_), .A3(G238), .A4(new_n281_), .ZN(new_n571_) );
  NAND4_X1 g0435 ( .A1(new_n171_), .A2(new_n255_), .A3(G244), .A4(G1698), .ZN(new_n572_) );
  NAND2_X1 g0436 ( .A1(new_n571_), .A2(new_n572_), .ZN(new_n573_) );
  NAND2_X1 g0437 ( .A1(new_n573_), .A2(KEYINPUT8), .ZN(new_n574_) );
  INV_X1 g0438 ( .A(KEYINPUT8), .ZN(new_n575_) );
  NAND3_X1 g0439 ( .A1(new_n571_), .A2(new_n572_), .A3(new_n575_), .ZN(new_n576_) );
  NAND3_X1 g0440 ( .A1(new_n171_), .A2(G116), .A3(new_n294_), .ZN(new_n577_) );
  NAND2_X1 g0441 ( .A1(new_n250_), .A2(G45), .ZN(new_n578_) );
  NAND3_X1 g0442 ( .A1(new_n303_), .A2(G250), .A3(new_n578_), .ZN(new_n579_) );
  NAND3_X1 g0443 ( .A1(new_n250_), .A2(G45), .A3(G274), .ZN(new_n580_) );
  NAND3_X1 g0444 ( .A1(new_n579_), .A2(new_n577_), .A3(new_n580_), .ZN(new_n581_) );
  INV_X1 g0445 ( .A(new_n581_), .ZN(new_n582_) );
  NAND3_X1 g0446 ( .A1(new_n582_), .A2(new_n574_), .A3(new_n576_), .ZN(new_n583_) );
  NAND2_X1 g0447 ( .A1(new_n583_), .A2(G169), .ZN(new_n584_) );
  INV_X1 g0448 ( .A(new_n583_), .ZN(new_n585_) );
  NAND2_X1 g0449 ( .A1(new_n585_), .A2(G179), .ZN(new_n586_) );
  NAND2_X1 g0450 ( .A1(new_n586_), .A2(new_n584_), .ZN(new_n587_) );
  NAND2_X1 g0451 ( .A1(new_n570_), .A2(new_n587_), .ZN(new_n588_) );
  NAND2_X1 g0452 ( .A1(new_n583_), .A2(G200), .ZN(new_n589_) );
  NAND4_X1 g0453 ( .A1(new_n582_), .A2(G190), .A3(new_n574_), .A4(new_n576_), .ZN(new_n590_) );
  NAND2_X1 g0454 ( .A1(new_n589_), .A2(new_n590_), .ZN(new_n591_) );
  INV_X1 g0455 ( .A(new_n591_), .ZN(new_n592_) );
  NAND4_X1 g0456 ( .A1(new_n592_), .A2(new_n562_), .A3(new_n564_), .A4(new_n569_), .ZN(new_n593_) );
  NAND2_X1 g0457 ( .A1(new_n588_), .A2(new_n593_), .ZN(new_n594_) );
  INV_X1 g0458 ( .A(new_n594_), .ZN(new_n595_) );
  NAND2_X1 g0459 ( .A1(new_n595_), .A2(new_n557_), .ZN(new_n596_) );
  INV_X1 g0460 ( .A(new_n596_), .ZN(new_n597_) );
  NAND3_X1 g0461 ( .A1(new_n597_), .A2(new_n488_), .A3(new_n524_), .ZN(new_n598_) );
  NOR2_X1 g0462 ( .A1(new_n437_), .A2(new_n598_), .ZN(G372) );
  INV_X1 g0463 ( .A(new_n549_), .ZN(new_n600_) );
  NAND2_X1 g0464 ( .A1(new_n488_), .A2(new_n600_), .ZN(new_n601_) );
  NAND2_X1 g0465 ( .A1(new_n601_), .A2(new_n478_), .ZN(new_n602_) );
  NAND2_X1 g0466 ( .A1(new_n602_), .A2(new_n524_), .ZN(new_n603_) );
  NAND3_X1 g0467 ( .A1(new_n603_), .A2(new_n519_), .A3(new_n588_), .ZN(new_n604_) );
  NAND2_X1 g0468 ( .A1(new_n604_), .A2(new_n593_), .ZN(new_n605_) );
  INV_X1 g0469 ( .A(new_n605_), .ZN(new_n606_) );
  NAND2_X1 g0470 ( .A1(new_n606_), .A2(new_n436_), .ZN(new_n607_) );
  NAND3_X1 g0471 ( .A1(new_n434_), .A2(new_n339_), .A3(new_n348_), .ZN(new_n608_) );
  NAND2_X1 g0472 ( .A1(new_n608_), .A2(new_n432_), .ZN(new_n609_) );
  NAND2_X1 g0473 ( .A1(new_n609_), .A2(new_n361_), .ZN(new_n610_) );
  NAND2_X1 g0474 ( .A1(new_n610_), .A2(new_n317_), .ZN(new_n611_) );
  NAND2_X1 g0475 ( .A1(new_n611_), .A2(new_n395_), .ZN(new_n612_) );
  NAND2_X1 g0476 ( .A1(new_n612_), .A2(new_n387_), .ZN(new_n613_) );
  INV_X1 g0477 ( .A(new_n613_), .ZN(new_n614_) );
  NAND2_X1 g0478 ( .A1(new_n607_), .A2(new_n614_), .ZN(G369) );
  INV_X1 g0479 ( .A(G343), .ZN(new_n616_) );
  NAND4_X1 g0480 ( .A1(new_n250_), .A2(new_n254_), .A3(G13), .A4(G213), .ZN(new_n617_) );
  NOR2_X1 g0481 ( .A1(new_n617_), .A2(new_n616_), .ZN(new_n618_) );
  NAND2_X1 g0482 ( .A1(new_n533_), .A2(new_n618_), .ZN(new_n619_) );
  NAND2_X1 g0483 ( .A1(new_n557_), .A2(new_n619_), .ZN(new_n620_) );
  NAND2_X1 g0484 ( .A1(new_n600_), .A2(new_n618_), .ZN(new_n621_) );
  NAND2_X1 g0485 ( .A1(new_n620_), .A2(new_n621_), .ZN(new_n622_) );
  NAND2_X1 g0486 ( .A1(new_n622_), .A2(G330), .ZN(new_n623_) );
  NAND2_X1 g0487 ( .A1(new_n456_), .A2(new_n618_), .ZN(new_n624_) );
  NAND2_X1 g0488 ( .A1(new_n488_), .A2(new_n624_), .ZN(new_n625_) );
  NAND3_X1 g0489 ( .A1(new_n477_), .A2(new_n456_), .A3(new_n618_), .ZN(new_n626_) );
  NAND2_X1 g0490 ( .A1(new_n625_), .A2(new_n626_), .ZN(new_n627_) );
  INV_X1 g0491 ( .A(new_n627_), .ZN(new_n628_) );
  NOR2_X1 g0492 ( .A1(new_n628_), .A2(new_n623_), .ZN(new_n629_) );
  INV_X1 g0493 ( .A(new_n629_), .ZN(new_n630_) );
  INV_X1 g0494 ( .A(new_n618_), .ZN(new_n631_) );
  NAND2_X1 g0495 ( .A1(new_n602_), .A2(new_n631_), .ZN(new_n632_) );
  NAND2_X1 g0496 ( .A1(new_n630_), .A2(new_n632_), .ZN(G399) );
  NAND2_X1 g0497 ( .A1(new_n606_), .A2(new_n631_), .ZN(new_n634_) );
  NAND4_X1 g0498 ( .A1(new_n597_), .A2(new_n488_), .A3(new_n524_), .A4(new_n631_), .ZN(new_n635_) );
  INV_X1 g0499 ( .A(new_n545_), .ZN(new_n636_) );
  INV_X1 g0500 ( .A(KEYINPUT18), .ZN(new_n637_) );
  NAND3_X1 g0501 ( .A1(new_n498_), .A2(new_n500_), .A3(new_n585_), .ZN(new_n638_) );
  NAND2_X1 g0502 ( .A1(new_n638_), .A2(new_n637_), .ZN(new_n639_) );
  NAND4_X1 g0503 ( .A1(new_n498_), .A2(KEYINPUT18), .A3(new_n500_), .A4(new_n585_), .ZN(new_n640_) );
  NAND2_X1 g0504 ( .A1(new_n639_), .A2(new_n640_), .ZN(new_n641_) );
  NAND3_X1 g0505 ( .A1(new_n641_), .A2(new_n475_), .A3(new_n636_), .ZN(new_n642_) );
  NOR2_X1 g0506 ( .A1(new_n475_), .A2(G179), .ZN(new_n643_) );
  NAND4_X1 g0507 ( .A1(new_n501_), .A2(new_n546_), .A3(new_n583_), .A4(new_n643_), .ZN(new_n644_) );
  NAND2_X1 g0508 ( .A1(new_n642_), .A2(new_n644_), .ZN(new_n645_) );
  NAND2_X1 g0509 ( .A1(new_n645_), .A2(new_n618_), .ZN(new_n646_) );
  NAND2_X1 g0510 ( .A1(new_n635_), .A2(new_n646_), .ZN(new_n647_) );
  NAND2_X1 g0511 ( .A1(new_n647_), .A2(G330), .ZN(new_n648_) );
  NAND2_X1 g0512 ( .A1(new_n634_), .A2(new_n648_), .ZN(new_n649_) );
  NAND2_X1 g0513 ( .A1(new_n649_), .A2(new_n250_), .ZN(new_n650_) );
  NOR2_X1 g0514 ( .A1(new_n561_), .A2(G116), .ZN(new_n651_) );
  INV_X1 g0515 ( .A(new_n176_), .ZN(new_n652_) );
  NOR2_X1 g0516 ( .A1(new_n652_), .A2(G41), .ZN(new_n653_) );
  INV_X1 g0517 ( .A(new_n653_), .ZN(new_n654_) );
  NAND3_X1 g0518 ( .A1(new_n654_), .A2(G1), .A3(new_n651_), .ZN(new_n655_) );
  NAND2_X1 g0519 ( .A1(new_n653_), .A2(new_n174_), .ZN(new_n656_) );
  NAND3_X1 g0520 ( .A1(new_n650_), .A2(new_n655_), .A3(new_n656_), .ZN(G364) );
  INV_X1 g0521 ( .A(new_n622_), .ZN(new_n658_) );
  NOR2_X1 g0522 ( .A1(G13), .A2(G33), .ZN(new_n659_) );
  INV_X1 g0523 ( .A(new_n659_), .ZN(new_n660_) );
  NOR2_X1 g0524 ( .A1(new_n660_), .A2(G20), .ZN(new_n661_) );
  NAND3_X1 g0525 ( .A1(new_n658_), .A2(KEYINPUT62), .A3(new_n661_), .ZN(new_n662_) );
  INV_X1 g0526 ( .A(KEYINPUT62), .ZN(new_n663_) );
  NAND2_X1 g0527 ( .A1(new_n658_), .A2(new_n661_), .ZN(new_n664_) );
  NAND2_X1 g0528 ( .A1(new_n664_), .A2(new_n663_), .ZN(new_n665_) );
  NAND3_X1 g0529 ( .A1(new_n176_), .A2(G33), .A3(KEYINPUT24), .ZN(new_n666_) );
  INV_X1 g0530 ( .A(KEYINPUT24), .ZN(new_n667_) );
  NAND2_X1 g0531 ( .A1(new_n176_), .A2(G33), .ZN(new_n668_) );
  NAND2_X1 g0532 ( .A1(new_n668_), .A2(new_n667_), .ZN(new_n669_) );
  NAND2_X1 g0533 ( .A1(new_n669_), .A2(new_n666_), .ZN(new_n670_) );
  NAND2_X1 g0534 ( .A1(new_n232_), .A2(G45), .ZN(new_n671_) );
  NAND2_X1 g0535 ( .A1(new_n174_), .A2(new_n291_), .ZN(new_n672_) );
  NAND3_X1 g0536 ( .A1(new_n671_), .A2(new_n670_), .A3(new_n672_), .ZN(new_n673_) );
  NAND3_X1 g0537 ( .A1(new_n652_), .A2(new_n219_), .A3(KEYINPUT60), .ZN(new_n674_) );
  NAND2_X1 g0538 ( .A1(G355), .A2(new_n659_), .ZN(new_n675_) );
  INV_X1 g0539 ( .A(KEYINPUT60), .ZN(new_n676_) );
  NAND2_X1 g0540 ( .A1(new_n652_), .A2(new_n219_), .ZN(new_n677_) );
  NAND2_X1 g0541 ( .A1(new_n677_), .A2(new_n676_), .ZN(new_n678_) );
  NAND4_X1 g0542 ( .A1(new_n673_), .A2(new_n674_), .A3(new_n675_), .A4(new_n678_), .ZN(new_n679_) );
  INV_X1 g0543 ( .A(new_n661_), .ZN(new_n680_) );
  NAND2_X1 g0544 ( .A1(new_n385_), .A2(G20), .ZN(new_n681_) );
  NAND2_X1 g0545 ( .A1(new_n171_), .A2(new_n681_), .ZN(new_n682_) );
  NAND2_X1 g0546 ( .A1(new_n680_), .A2(new_n682_), .ZN(new_n683_) );
  INV_X1 g0547 ( .A(new_n683_), .ZN(new_n684_) );
  NAND2_X1 g0548 ( .A1(new_n679_), .A2(new_n684_), .ZN(new_n685_) );
  INV_X1 g0549 ( .A(new_n685_), .ZN(new_n686_) );
  INV_X1 g0550 ( .A(G190), .ZN(new_n687_) );
  NOR2_X1 g0551 ( .A1(new_n687_), .A2(G200), .ZN(new_n688_) );
  NAND2_X1 g0552 ( .A1(new_n688_), .A2(new_n370_), .ZN(new_n689_) );
  NAND2_X1 g0553 ( .A1(new_n689_), .A2(G20), .ZN(new_n690_) );
  INV_X1 g0554 ( .A(new_n690_), .ZN(new_n691_) );
  NOR2_X1 g0555 ( .A1(new_n691_), .A2(new_n506_), .ZN(new_n692_) );
  INV_X1 g0556 ( .A(G200), .ZN(new_n693_) );
  NAND2_X1 g0557 ( .A1(G20), .A2(G179), .ZN(new_n694_) );
  NOR3_X1 g0558 ( .A1(new_n694_), .A2(new_n693_), .A3(G190), .ZN(new_n695_) );
  INV_X1 g0559 ( .A(new_n695_), .ZN(new_n696_) );
  NOR2_X1 g0560 ( .A1(new_n696_), .A2(new_n409_), .ZN(new_n697_) );
  NOR2_X1 g0561 ( .A1(new_n254_), .A2(G179), .ZN(new_n698_) );
  NAND3_X1 g0562 ( .A1(new_n698_), .A2(new_n687_), .A3(new_n693_), .ZN(new_n699_) );
  INV_X1 g0563 ( .A(new_n699_), .ZN(new_n700_) );
  NAND2_X1 g0564 ( .A1(new_n700_), .A2(G159), .ZN(new_n701_) );
  NOR3_X1 g0565 ( .A1(new_n694_), .A2(G190), .A3(G200), .ZN(new_n702_) );
  INV_X1 g0566 ( .A(new_n702_), .ZN(new_n703_) );
  NOR2_X1 g0567 ( .A1(new_n703_), .A2(new_n140_), .ZN(new_n704_) );
  INV_X1 g0568 ( .A(new_n704_), .ZN(new_n705_) );
  NAND2_X1 g0569 ( .A1(new_n705_), .A2(new_n701_), .ZN(new_n706_) );
  NOR3_X1 g0570 ( .A1(new_n706_), .A2(new_n692_), .A3(new_n697_), .ZN(new_n707_) );
  NAND2_X1 g0571 ( .A1(new_n707_), .A2(KEYINPUT61), .ZN(new_n708_) );
  INV_X1 g0572 ( .A(KEYINPUT61), .ZN(new_n709_) );
  INV_X1 g0573 ( .A(new_n707_), .ZN(new_n710_) );
  NAND2_X1 g0574 ( .A1(new_n710_), .A2(new_n709_), .ZN(new_n711_) );
  INV_X1 g0575 ( .A(new_n682_), .ZN(new_n712_) );
  NAND2_X1 g0576 ( .A1(new_n712_), .A2(new_n255_), .ZN(new_n713_) );
  NAND3_X1 g0577 ( .A1(new_n698_), .A2(new_n687_), .A3(G200), .ZN(new_n714_) );
  NOR2_X1 g0578 ( .A1(new_n714_), .A2(new_n439_), .ZN(new_n715_) );
  NAND2_X1 g0579 ( .A1(G190), .A2(G200), .ZN(new_n716_) );
  INV_X1 g0580 ( .A(new_n716_), .ZN(new_n717_) );
  NAND2_X1 g0581 ( .A1(new_n698_), .A2(new_n717_), .ZN(new_n718_) );
  INV_X1 g0582 ( .A(new_n718_), .ZN(new_n719_) );
  NAND2_X1 g0583 ( .A1(new_n719_), .A2(G87), .ZN(new_n720_) );
  INV_X1 g0584 ( .A(new_n694_), .ZN(new_n721_) );
  NAND2_X1 g0585 ( .A1(new_n688_), .A2(new_n721_), .ZN(new_n722_) );
  INV_X1 g0586 ( .A(new_n722_), .ZN(new_n723_) );
  NAND2_X1 g0587 ( .A1(new_n723_), .A2(G58), .ZN(new_n724_) );
  NOR2_X1 g0588 ( .A1(new_n694_), .A2(new_n716_), .ZN(new_n725_) );
  NAND2_X1 g0589 ( .A1(new_n725_), .A2(G50), .ZN(new_n726_) );
  NAND3_X1 g0590 ( .A1(new_n720_), .A2(new_n724_), .A3(new_n726_), .ZN(new_n727_) );
  NOR3_X1 g0591 ( .A1(new_n727_), .A2(new_n713_), .A3(new_n715_), .ZN(new_n728_) );
  NAND3_X1 g0592 ( .A1(new_n711_), .A2(new_n708_), .A3(new_n728_), .ZN(new_n729_) );
  INV_X1 g0593 ( .A(new_n714_), .ZN(new_n730_) );
  NAND2_X1 g0594 ( .A1(new_n730_), .A2(G283), .ZN(new_n731_) );
  NAND2_X1 g0595 ( .A1(new_n700_), .A2(G329), .ZN(new_n732_) );
  NAND2_X1 g0596 ( .A1(new_n702_), .A2(G311), .ZN(new_n733_) );
  NAND2_X1 g0597 ( .A1(new_n712_), .A2(G33), .ZN(new_n734_) );
  NAND2_X1 g0598 ( .A1(new_n719_), .A2(G303), .ZN(new_n735_) );
  NAND2_X1 g0599 ( .A1(new_n723_), .A2(G322), .ZN(new_n736_) );
  NAND2_X1 g0600 ( .A1(new_n725_), .A2(G326), .ZN(new_n737_) );
  NAND3_X1 g0601 ( .A1(new_n735_), .A2(new_n736_), .A3(new_n737_), .ZN(new_n738_) );
  INV_X1 g0602 ( .A(G294), .ZN(new_n739_) );
  NOR2_X1 g0603 ( .A1(new_n691_), .A2(new_n739_), .ZN(new_n740_) );
  INV_X1 g0604 ( .A(G317), .ZN(new_n741_) );
  NOR2_X1 g0605 ( .A1(new_n696_), .A2(new_n741_), .ZN(new_n742_) );
  NOR4_X1 g0606 ( .A1(new_n738_), .A2(new_n740_), .A3(new_n734_), .A4(new_n742_), .ZN(new_n743_) );
  NAND4_X1 g0607 ( .A1(new_n743_), .A2(new_n731_), .A3(new_n732_), .A4(new_n733_), .ZN(new_n744_) );
  INV_X1 g0608 ( .A(KEYINPUT1), .ZN(new_n745_) );
  NAND3_X1 g0609 ( .A1(new_n254_), .A2(G13), .A3(G45), .ZN(new_n746_) );
  NAND2_X1 g0610 ( .A1(new_n746_), .A2(G1), .ZN(new_n747_) );
  NAND2_X1 g0611 ( .A1(new_n747_), .A2(new_n745_), .ZN(new_n748_) );
  NAND3_X1 g0612 ( .A1(new_n746_), .A2(G1), .A3(KEYINPUT1), .ZN(new_n749_) );
  NAND2_X1 g0613 ( .A1(new_n748_), .A2(new_n749_), .ZN(new_n750_) );
  INV_X1 g0614 ( .A(new_n750_), .ZN(new_n751_) );
  NAND2_X1 g0615 ( .A1(new_n751_), .A2(new_n654_), .ZN(new_n752_) );
  INV_X1 g0616 ( .A(new_n752_), .ZN(new_n753_) );
  NAND3_X1 g0617 ( .A1(new_n729_), .A2(new_n744_), .A3(new_n753_), .ZN(new_n754_) );
  NOR2_X1 g0618 ( .A1(new_n754_), .A2(new_n686_), .ZN(new_n755_) );
  NAND3_X1 g0619 ( .A1(new_n665_), .A2(new_n662_), .A3(new_n755_), .ZN(new_n756_) );
  INV_X1 g0620 ( .A(G330), .ZN(new_n757_) );
  NAND2_X1 g0621 ( .A1(new_n658_), .A2(new_n757_), .ZN(new_n758_) );
  NAND3_X1 g0622 ( .A1(new_n758_), .A2(new_n623_), .A3(new_n752_), .ZN(new_n759_) );
  NAND2_X1 g0623 ( .A1(new_n756_), .A2(new_n759_), .ZN(G396) );
  INV_X1 g0624 ( .A(new_n649_), .ZN(new_n761_) );
  INV_X1 g0625 ( .A(KEYINPUT5), .ZN(new_n762_) );
  NAND2_X1 g0626 ( .A1(new_n348_), .A2(new_n618_), .ZN(new_n763_) );
  NAND2_X1 g0627 ( .A1(new_n763_), .A2(new_n762_), .ZN(new_n764_) );
  NAND3_X1 g0628 ( .A1(new_n348_), .A2(KEYINPUT5), .A3(new_n618_), .ZN(new_n765_) );
  NAND2_X1 g0629 ( .A1(new_n764_), .A2(new_n765_), .ZN(new_n766_) );
  NAND3_X1 g0630 ( .A1(new_n349_), .A2(new_n766_), .A3(new_n352_), .ZN(new_n767_) );
  NAND3_X1 g0631 ( .A1(new_n339_), .A2(new_n765_), .A3(new_n764_), .ZN(new_n768_) );
  NAND2_X1 g0632 ( .A1(new_n767_), .A2(new_n768_), .ZN(new_n769_) );
  NAND2_X1 g0633 ( .A1(new_n761_), .A2(new_n769_), .ZN(new_n770_) );
  INV_X1 g0634 ( .A(new_n769_), .ZN(new_n771_) );
  NAND2_X1 g0635 ( .A1(new_n649_), .A2(new_n771_), .ZN(new_n772_) );
  NAND2_X1 g0636 ( .A1(new_n770_), .A2(new_n772_), .ZN(new_n773_) );
  NAND2_X1 g0637 ( .A1(new_n773_), .A2(new_n752_), .ZN(new_n774_) );
  NAND2_X1 g0638 ( .A1(new_n771_), .A2(new_n659_), .ZN(new_n775_) );
  NAND2_X1 g0639 ( .A1(new_n730_), .A2(G68), .ZN(new_n776_) );
  NAND2_X1 g0640 ( .A1(new_n695_), .A2(G150), .ZN(new_n777_) );
  NAND2_X1 g0641 ( .A1(new_n723_), .A2(G143), .ZN(new_n778_) );
  NAND2_X1 g0642 ( .A1(new_n700_), .A2(G132), .ZN(new_n779_) );
  NOR2_X1 g0643 ( .A1(new_n779_), .A2(KEYINPUT19), .ZN(new_n780_) );
  INV_X1 g0644 ( .A(new_n713_), .ZN(new_n781_) );
  NAND2_X1 g0645 ( .A1(new_n779_), .A2(KEYINPUT19), .ZN(new_n782_) );
  NAND2_X1 g0646 ( .A1(new_n781_), .A2(new_n782_), .ZN(new_n783_) );
  NOR2_X1 g0647 ( .A1(new_n783_), .A2(new_n780_), .ZN(new_n784_) );
  NAND4_X1 g0648 ( .A1(new_n784_), .A2(new_n776_), .A3(new_n777_), .A4(new_n778_), .ZN(new_n785_) );
  NAND2_X1 g0649 ( .A1(new_n702_), .A2(G159), .ZN(new_n786_) );
  NAND2_X1 g0650 ( .A1(new_n690_), .A2(G58), .ZN(new_n787_) );
  NAND2_X1 g0651 ( .A1(new_n719_), .A2(G50), .ZN(new_n788_) );
  NAND2_X1 g0652 ( .A1(new_n725_), .A2(G137), .ZN(new_n789_) );
  NAND4_X1 g0653 ( .A1(new_n787_), .A2(new_n788_), .A3(new_n786_), .A4(new_n789_), .ZN(new_n790_) );
  NOR2_X1 g0654 ( .A1(new_n790_), .A2(KEYINPUT20), .ZN(new_n791_) );
  NAND2_X1 g0655 ( .A1(new_n790_), .A2(KEYINPUT20), .ZN(new_n792_) );
  INV_X1 g0656 ( .A(new_n792_), .ZN(new_n793_) );
  NOR3_X1 g0657 ( .A1(new_n785_), .A2(new_n791_), .A3(new_n793_), .ZN(new_n794_) );
  NAND2_X1 g0658 ( .A1(new_n702_), .A2(G116), .ZN(new_n795_) );
  NAND2_X1 g0659 ( .A1(new_n795_), .A2(KEYINPUT21), .ZN(new_n796_) );
  NOR2_X1 g0660 ( .A1(new_n795_), .A2(KEYINPUT21), .ZN(new_n797_) );
  NAND2_X1 g0661 ( .A1(new_n719_), .A2(G107), .ZN(new_n798_) );
  NAND2_X1 g0662 ( .A1(new_n723_), .A2(G294), .ZN(new_n799_) );
  NAND2_X1 g0663 ( .A1(new_n725_), .A2(G303), .ZN(new_n800_) );
  NAND4_X1 g0664 ( .A1(new_n798_), .A2(new_n799_), .A3(G33), .A4(new_n800_), .ZN(new_n801_) );
  NOR2_X1 g0665 ( .A1(new_n801_), .A2(new_n797_), .ZN(new_n802_) );
  INV_X1 g0666 ( .A(KEYINPUT22), .ZN(new_n803_) );
  NAND3_X1 g0667 ( .A1(new_n730_), .A2(G87), .A3(new_n803_), .ZN(new_n804_) );
  NAND2_X1 g0668 ( .A1(new_n730_), .A2(G87), .ZN(new_n805_) );
  NAND2_X1 g0669 ( .A1(new_n805_), .A2(KEYINPUT22), .ZN(new_n806_) );
  NAND2_X1 g0670 ( .A1(new_n806_), .A2(new_n804_), .ZN(new_n807_) );
  INV_X1 g0671 ( .A(G311), .ZN(new_n808_) );
  NOR2_X1 g0672 ( .A1(new_n699_), .A2(new_n808_), .ZN(new_n809_) );
  INV_X1 g0673 ( .A(G283), .ZN(new_n810_) );
  NOR2_X1 g0674 ( .A1(new_n696_), .A2(new_n810_), .ZN(new_n811_) );
  NOR4_X1 g0675 ( .A1(new_n692_), .A2(new_n682_), .A3(new_n809_), .A4(new_n811_), .ZN(new_n812_) );
  NAND4_X1 g0676 ( .A1(new_n812_), .A2(new_n796_), .A3(new_n802_), .A4(new_n807_), .ZN(new_n813_) );
  NAND2_X1 g0677 ( .A1(new_n682_), .A2(new_n660_), .ZN(new_n814_) );
  INV_X1 g0678 ( .A(new_n814_), .ZN(new_n815_) );
  NAND2_X1 g0679 ( .A1(new_n815_), .A2(new_n140_), .ZN(new_n816_) );
  NAND3_X1 g0680 ( .A1(new_n813_), .A2(new_n753_), .A3(new_n816_), .ZN(new_n817_) );
  NOR2_X1 g0681 ( .A1(new_n794_), .A2(new_n817_), .ZN(new_n818_) );
  NAND2_X1 g0682 ( .A1(new_n775_), .A2(new_n818_), .ZN(new_n819_) );
  NAND2_X1 g0683 ( .A1(new_n774_), .A2(new_n819_), .ZN(G384) );
  INV_X1 g0684 ( .A(new_n648_), .ZN(new_n821_) );
  NAND2_X1 g0685 ( .A1(new_n318_), .A2(new_n617_), .ZN(new_n822_) );
  NAND3_X1 g0686 ( .A1(new_n604_), .A2(new_n352_), .A3(new_n593_), .ZN(new_n823_) );
  NAND2_X1 g0687 ( .A1(new_n823_), .A2(new_n349_), .ZN(new_n824_) );
  INV_X1 g0688 ( .A(KEYINPUT29), .ZN(new_n825_) );
  NAND2_X1 g0689 ( .A1(new_n428_), .A2(new_n618_), .ZN(new_n826_) );
  NAND3_X1 g0690 ( .A1(new_n426_), .A2(new_n432_), .A3(new_n826_), .ZN(new_n827_) );
  NAND2_X1 g0691 ( .A1(new_n433_), .A2(new_n618_), .ZN(new_n828_) );
  NAND2_X1 g0692 ( .A1(new_n827_), .A2(new_n828_), .ZN(new_n829_) );
  NAND2_X1 g0693 ( .A1(new_n829_), .A2(new_n825_), .ZN(new_n830_) );
  NAND3_X1 g0694 ( .A1(new_n827_), .A2(KEYINPUT29), .A3(new_n828_), .ZN(new_n831_) );
  NAND2_X1 g0695 ( .A1(new_n830_), .A2(new_n831_), .ZN(new_n832_) );
  NAND3_X1 g0696 ( .A1(new_n824_), .A2(new_n631_), .A3(new_n832_), .ZN(new_n833_) );
  NAND2_X1 g0697 ( .A1(new_n433_), .A2(new_n631_), .ZN(new_n834_) );
  NAND2_X1 g0698 ( .A1(new_n833_), .A2(new_n834_), .ZN(new_n835_) );
  INV_X1 g0699 ( .A(new_n617_), .ZN(new_n836_) );
  NAND2_X1 g0700 ( .A1(new_n275_), .A2(new_n836_), .ZN(new_n837_) );
  NAND2_X1 g0701 ( .A1(new_n361_), .A2(new_n837_), .ZN(new_n838_) );
  NAND2_X1 g0702 ( .A1(new_n838_), .A2(new_n317_), .ZN(new_n839_) );
  NAND2_X1 g0703 ( .A1(new_n839_), .A2(new_n822_), .ZN(new_n840_) );
  INV_X1 g0704 ( .A(new_n840_), .ZN(new_n841_) );
  NAND2_X1 g0705 ( .A1(new_n835_), .A2(new_n841_), .ZN(new_n842_) );
  NAND4_X1 g0706 ( .A1(new_n436_), .A2(new_n604_), .A3(new_n593_), .A4(new_n631_), .ZN(new_n843_) );
  NAND4_X1 g0707 ( .A1(new_n842_), .A2(new_n614_), .A3(new_n822_), .A4(new_n843_), .ZN(new_n844_) );
  NAND2_X1 g0708 ( .A1(new_n842_), .A2(new_n822_), .ZN(new_n845_) );
  NAND2_X1 g0709 ( .A1(new_n614_), .A2(new_n843_), .ZN(new_n846_) );
  NAND2_X1 g0710 ( .A1(new_n845_), .A2(new_n846_), .ZN(new_n847_) );
  NAND2_X1 g0711 ( .A1(new_n832_), .A2(new_n769_), .ZN(new_n848_) );
  NOR2_X1 g0712 ( .A1(new_n840_), .A2(new_n848_), .ZN(new_n849_) );
  INV_X1 g0713 ( .A(new_n849_), .ZN(new_n850_) );
  NAND2_X1 g0714 ( .A1(new_n850_), .A2(new_n436_), .ZN(new_n851_) );
  NAND2_X1 g0715 ( .A1(new_n849_), .A2(new_n437_), .ZN(new_n852_) );
  NAND2_X1 g0716 ( .A1(new_n851_), .A2(new_n852_), .ZN(new_n853_) );
  NAND4_X1 g0717 ( .A1(new_n847_), .A2(new_n821_), .A3(new_n844_), .A4(new_n853_), .ZN(new_n854_) );
  NAND2_X1 g0718 ( .A1(new_n847_), .A2(new_n844_), .ZN(new_n855_) );
  NAND2_X1 g0719 ( .A1(new_n853_), .A2(new_n821_), .ZN(new_n856_) );
  NAND2_X1 g0720 ( .A1(new_n855_), .A2(new_n856_), .ZN(new_n857_) );
  NAND3_X1 g0721 ( .A1(new_n857_), .A2(new_n172_), .A3(new_n854_), .ZN(new_n858_) );
  INV_X1 g0722 ( .A(G13), .ZN(new_n859_) );
  NAND2_X1 g0723 ( .A1(new_n859_), .A2(G1), .ZN(new_n860_) );
  NAND2_X1 g0724 ( .A1(new_n858_), .A2(new_n860_), .ZN(new_n861_) );
  NAND3_X1 g0725 ( .A1(G50), .A2(G58), .A3(G68), .ZN(new_n862_) );
  NAND2_X1 g0726 ( .A1(G50), .A2(G58), .ZN(new_n863_) );
  NAND2_X1 g0727 ( .A1(new_n863_), .A2(new_n409_), .ZN(new_n864_) );
  NAND2_X1 g0728 ( .A1(new_n140_), .A2(G50), .ZN(new_n865_) );
  NAND3_X1 g0729 ( .A1(new_n864_), .A2(new_n862_), .A3(new_n865_), .ZN(new_n866_) );
  NAND3_X1 g0730 ( .A1(new_n866_), .A2(G1), .A3(new_n859_), .ZN(new_n867_) );
  NAND2_X1 g0731 ( .A1(new_n861_), .A2(new_n867_), .ZN(new_n868_) );
  NAND3_X1 g0732 ( .A1(new_n173_), .A2(G116), .A3(new_n213_), .ZN(new_n869_) );
  NAND2_X1 g0733 ( .A1(new_n868_), .A2(new_n869_), .ZN(G367) );
  INV_X1 g0734 ( .A(KEYINPUT53), .ZN(new_n871_) );
  NAND2_X1 g0735 ( .A1(new_n603_), .A2(new_n519_), .ZN(new_n872_) );
  NAND2_X1 g0736 ( .A1(new_n872_), .A2(new_n594_), .ZN(new_n873_) );
  NAND3_X1 g0737 ( .A1(new_n603_), .A2(new_n519_), .A3(new_n595_), .ZN(new_n874_) );
  NAND2_X1 g0738 ( .A1(new_n873_), .A2(new_n874_), .ZN(new_n875_) );
  NAND2_X1 g0739 ( .A1(new_n875_), .A2(new_n631_), .ZN(new_n876_) );
  NAND2_X1 g0740 ( .A1(new_n593_), .A2(new_n618_), .ZN(new_n877_) );
  NAND3_X1 g0741 ( .A1(new_n876_), .A2(new_n871_), .A3(new_n877_), .ZN(new_n878_) );
  NAND2_X1 g0742 ( .A1(new_n876_), .A2(new_n877_), .ZN(new_n879_) );
  NAND2_X1 g0743 ( .A1(new_n879_), .A2(KEYINPUT53), .ZN(new_n880_) );
  NAND4_X1 g0744 ( .A1(new_n570_), .A2(new_n584_), .A3(new_n586_), .A4(new_n618_), .ZN(new_n881_) );
  NAND3_X1 g0745 ( .A1(new_n880_), .A2(new_n878_), .A3(new_n881_), .ZN(new_n882_) );
  NAND2_X1 g0746 ( .A1(new_n518_), .A2(new_n618_), .ZN(new_n883_) );
  NAND2_X1 g0747 ( .A1(new_n524_), .A2(new_n883_), .ZN(new_n884_) );
  NAND4_X1 g0748 ( .A1(new_n502_), .A2(new_n503_), .A3(new_n518_), .A4(new_n618_), .ZN(new_n885_) );
  NAND2_X1 g0749 ( .A1(new_n884_), .A2(new_n885_), .ZN(new_n886_) );
  NAND2_X1 g0750 ( .A1(new_n629_), .A2(new_n886_), .ZN(new_n887_) );
  INV_X1 g0751 ( .A(new_n887_), .ZN(new_n888_) );
  NAND2_X1 g0752 ( .A1(new_n882_), .A2(new_n888_), .ZN(new_n889_) );
  NAND4_X1 g0753 ( .A1(new_n880_), .A2(new_n878_), .A3(new_n881_), .A4(new_n887_), .ZN(new_n890_) );
  NAND2_X1 g0754 ( .A1(new_n889_), .A2(new_n890_), .ZN(new_n891_) );
  INV_X1 g0755 ( .A(KEYINPUT52), .ZN(new_n892_) );
  NAND2_X1 g0756 ( .A1(new_n632_), .A2(new_n883_), .ZN(new_n893_) );
  NAND2_X1 g0757 ( .A1(new_n893_), .A2(new_n523_), .ZN(new_n894_) );
  NAND3_X1 g0758 ( .A1(new_n632_), .A2(new_n524_), .A3(new_n883_), .ZN(new_n895_) );
  NAND2_X1 g0759 ( .A1(new_n894_), .A2(new_n895_), .ZN(new_n896_) );
  NAND2_X1 g0760 ( .A1(new_n896_), .A2(new_n630_), .ZN(new_n897_) );
  NAND3_X1 g0761 ( .A1(new_n894_), .A2(new_n629_), .A3(new_n895_), .ZN(new_n898_) );
  NAND2_X1 g0762 ( .A1(new_n897_), .A2(new_n898_), .ZN(new_n899_) );
  NAND2_X1 g0763 ( .A1(new_n600_), .A2(new_n631_), .ZN(new_n900_) );
  NAND3_X1 g0764 ( .A1(new_n488_), .A2(new_n624_), .A3(new_n900_), .ZN(new_n901_) );
  NAND2_X1 g0765 ( .A1(new_n900_), .A2(new_n624_), .ZN(new_n902_) );
  NAND3_X1 g0766 ( .A1(new_n902_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n903_) );
  NAND2_X1 g0767 ( .A1(new_n901_), .A2(new_n903_), .ZN(new_n904_) );
  NAND2_X1 g0768 ( .A1(new_n623_), .A2(new_n904_), .ZN(new_n905_) );
  NAND4_X1 g0769 ( .A1(new_n622_), .A2(new_n901_), .A3(G330), .A4(new_n903_), .ZN(new_n906_) );
  NAND2_X1 g0770 ( .A1(new_n905_), .A2(new_n906_), .ZN(new_n907_) );
  NAND3_X1 g0771 ( .A1(new_n899_), .A2(new_n892_), .A3(new_n907_), .ZN(new_n908_) );
  NAND2_X1 g0772 ( .A1(new_n899_), .A2(new_n907_), .ZN(new_n909_) );
  NAND2_X1 g0773 ( .A1(new_n909_), .A2(KEYINPUT52), .ZN(new_n910_) );
  NAND2_X1 g0774 ( .A1(new_n910_), .A2(new_n908_), .ZN(new_n911_) );
  NAND3_X1 g0775 ( .A1(new_n634_), .A2(new_n648_), .A3(new_n751_), .ZN(new_n912_) );
  INV_X1 g0776 ( .A(new_n912_), .ZN(new_n913_) );
  NAND2_X1 g0777 ( .A1(new_n911_), .A2(new_n913_), .ZN(new_n914_) );
  NAND3_X1 g0778 ( .A1(new_n891_), .A2(new_n752_), .A3(new_n914_), .ZN(new_n915_) );
  NAND2_X1 g0779 ( .A1(new_n594_), .A2(new_n661_), .ZN(new_n916_) );
  INV_X1 g0780 ( .A(new_n734_), .ZN(new_n917_) );
  NOR2_X1 g0781 ( .A1(new_n699_), .A2(new_n741_), .ZN(new_n918_) );
  NOR2_X1 g0782 ( .A1(new_n714_), .A2(new_n506_), .ZN(new_n919_) );
  NOR2_X1 g0783 ( .A1(new_n703_), .A2(new_n810_), .ZN(new_n920_) );
  NOR2_X1 g0784 ( .A1(new_n696_), .A2(new_n739_), .ZN(new_n921_) );
  NOR4_X1 g0785 ( .A1(new_n920_), .A2(new_n921_), .A3(new_n918_), .A4(new_n919_), .ZN(new_n922_) );
  INV_X1 g0786 ( .A(KEYINPUT54), .ZN(new_n923_) );
  NAND3_X1 g0787 ( .A1(new_n725_), .A2(G311), .A3(new_n923_), .ZN(new_n924_) );
  NAND2_X1 g0788 ( .A1(new_n725_), .A2(G311), .ZN(new_n925_) );
  NAND2_X1 g0789 ( .A1(new_n925_), .A2(KEYINPUT54), .ZN(new_n926_) );
  NAND2_X1 g0790 ( .A1(new_n926_), .A2(new_n924_), .ZN(new_n927_) );
  NOR2_X1 g0791 ( .A1(new_n691_), .A2(new_n439_), .ZN(new_n928_) );
  NOR2_X1 g0792 ( .A1(new_n718_), .A2(new_n219_), .ZN(new_n929_) );
  INV_X1 g0793 ( .A(G303), .ZN(new_n930_) );
  NOR2_X1 g0794 ( .A1(new_n722_), .A2(new_n930_), .ZN(new_n931_) );
  NOR3_X1 g0795 ( .A1(new_n928_), .A2(new_n929_), .A3(new_n931_), .ZN(new_n932_) );
  NAND4_X1 g0796 ( .A1(new_n932_), .A2(new_n922_), .A3(new_n917_), .A4(new_n927_), .ZN(new_n933_) );
  NOR2_X1 g0797 ( .A1(new_n691_), .A2(new_n409_), .ZN(new_n934_) );
  NOR2_X1 g0798 ( .A1(new_n714_), .A2(new_n140_), .ZN(new_n935_) );
  NOR2_X1 g0799 ( .A1(new_n703_), .A2(new_n139_), .ZN(new_n936_) );
  NOR3_X1 g0800 ( .A1(new_n934_), .A2(new_n935_), .A3(new_n936_), .ZN(new_n937_) );
  NAND2_X1 g0801 ( .A1(new_n719_), .A2(G58), .ZN(new_n938_) );
  NAND2_X1 g0802 ( .A1(new_n723_), .A2(G150), .ZN(new_n939_) );
  NAND2_X1 g0803 ( .A1(new_n725_), .A2(G143), .ZN(new_n940_) );
  NAND3_X1 g0804 ( .A1(new_n938_), .A2(new_n939_), .A3(new_n940_), .ZN(new_n941_) );
  NAND2_X1 g0805 ( .A1(new_n700_), .A2(G137), .ZN(new_n942_) );
  NAND2_X1 g0806 ( .A1(new_n695_), .A2(G159), .ZN(new_n943_) );
  NAND2_X1 g0807 ( .A1(new_n942_), .A2(new_n943_), .ZN(new_n944_) );
  NOR2_X1 g0808 ( .A1(new_n941_), .A2(new_n944_), .ZN(new_n945_) );
  NAND3_X1 g0809 ( .A1(new_n937_), .A2(new_n945_), .A3(new_n781_), .ZN(new_n946_) );
  NAND2_X1 g0810 ( .A1(new_n670_), .A2(new_n205_), .ZN(new_n947_) );
  NAND2_X1 g0811 ( .A1(new_n652_), .A2(G87), .ZN(new_n948_) );
  NAND3_X1 g0812 ( .A1(new_n947_), .A2(new_n684_), .A3(new_n948_), .ZN(new_n949_) );
  NAND4_X1 g0813 ( .A1(new_n933_), .A2(new_n753_), .A3(new_n946_), .A4(new_n949_), .ZN(new_n950_) );
  INV_X1 g0814 ( .A(new_n950_), .ZN(new_n951_) );
  NAND2_X1 g0815 ( .A1(new_n916_), .A2(new_n951_), .ZN(new_n952_) );
  NAND2_X1 g0816 ( .A1(new_n915_), .A2(new_n952_), .ZN(new_n953_) );
  NAND2_X1 g0817 ( .A1(new_n953_), .A2(KEYINPUT55), .ZN(new_n954_) );
  INV_X1 g0818 ( .A(KEYINPUT55), .ZN(new_n955_) );
  NAND3_X1 g0819 ( .A1(new_n915_), .A2(new_n955_), .A3(new_n952_), .ZN(new_n956_) );
  NAND2_X1 g0820 ( .A1(new_n954_), .A2(new_n956_), .ZN(new_n957_) );
  INV_X1 g0821 ( .A(new_n957_), .ZN(G387) );
  NAND3_X1 g0822 ( .A1(new_n912_), .A2(new_n752_), .A3(new_n907_), .ZN(new_n959_) );
  NAND4_X1 g0823 ( .A1(new_n761_), .A2(new_n653_), .A3(new_n905_), .A4(new_n906_), .ZN(new_n960_) );
  NAND2_X1 g0824 ( .A1(new_n628_), .A2(new_n661_), .ZN(new_n961_) );
  NAND2_X1 g0825 ( .A1(new_n207_), .A2(G45), .ZN(new_n962_) );
  INV_X1 g0826 ( .A(KEYINPUT23), .ZN(new_n963_) );
  NAND2_X1 g0827 ( .A1(G68), .A2(G77), .ZN(new_n964_) );
  NAND4_X1 g0828 ( .A1(new_n651_), .A2(new_n139_), .A3(G58), .A4(new_n964_), .ZN(new_n965_) );
  NAND2_X1 g0829 ( .A1(new_n965_), .A2(new_n291_), .ZN(new_n966_) );
  NAND2_X1 g0830 ( .A1(new_n966_), .A2(new_n963_), .ZN(new_n967_) );
  NAND3_X1 g0831 ( .A1(new_n965_), .A2(new_n291_), .A3(KEYINPUT23), .ZN(new_n968_) );
  NAND2_X1 g0832 ( .A1(new_n967_), .A2(new_n968_), .ZN(new_n969_) );
  NAND2_X1 g0833 ( .A1(new_n962_), .A2(new_n969_), .ZN(new_n970_) );
  NAND2_X1 g0834 ( .A1(new_n970_), .A2(new_n670_), .ZN(new_n971_) );
  INV_X1 g0835 ( .A(new_n651_), .ZN(new_n972_) );
  NAND2_X1 g0836 ( .A1(new_n972_), .A2(new_n659_), .ZN(new_n973_) );
  NAND2_X1 g0837 ( .A1(new_n652_), .A2(new_n439_), .ZN(new_n974_) );
  NAND3_X1 g0838 ( .A1(new_n971_), .A2(new_n973_), .A3(new_n974_), .ZN(new_n975_) );
  NAND2_X1 g0839 ( .A1(new_n975_), .A2(new_n684_), .ZN(new_n976_) );
  NAND2_X1 g0840 ( .A1(new_n695_), .A2(G311), .ZN(new_n977_) );
  NAND2_X1 g0841 ( .A1(new_n690_), .A2(G283), .ZN(new_n978_) );
  NAND2_X1 g0842 ( .A1(new_n700_), .A2(G326), .ZN(new_n979_) );
  NAND3_X1 g0843 ( .A1(new_n979_), .A2(new_n978_), .A3(new_n977_), .ZN(new_n980_) );
  NAND2_X1 g0844 ( .A1(new_n702_), .A2(G303), .ZN(new_n981_) );
  NAND2_X1 g0845 ( .A1(new_n723_), .A2(G317), .ZN(new_n982_) );
  NAND3_X1 g0846 ( .A1(new_n917_), .A2(new_n981_), .A3(new_n982_), .ZN(new_n983_) );
  INV_X1 g0847 ( .A(KEYINPUT26), .ZN(new_n984_) );
  NAND2_X1 g0848 ( .A1(new_n719_), .A2(G294), .ZN(new_n985_) );
  NAND2_X1 g0849 ( .A1(new_n725_), .A2(G322), .ZN(new_n986_) );
  NAND2_X1 g0850 ( .A1(new_n985_), .A2(new_n986_), .ZN(new_n987_) );
  NAND2_X1 g0851 ( .A1(new_n987_), .A2(new_n984_), .ZN(new_n988_) );
  NAND3_X1 g0852 ( .A1(new_n985_), .A2(KEYINPUT26), .A3(new_n986_), .ZN(new_n989_) );
  NAND2_X1 g0853 ( .A1(new_n988_), .A2(new_n989_), .ZN(new_n990_) );
  NAND3_X1 g0854 ( .A1(new_n730_), .A2(G116), .A3(KEYINPUT25), .ZN(new_n991_) );
  INV_X1 g0855 ( .A(KEYINPUT25), .ZN(new_n992_) );
  NAND2_X1 g0856 ( .A1(new_n730_), .A2(G116), .ZN(new_n993_) );
  NAND2_X1 g0857 ( .A1(new_n993_), .A2(new_n992_), .ZN(new_n994_) );
  NAND2_X1 g0858 ( .A1(new_n994_), .A2(new_n991_), .ZN(new_n995_) );
  NAND2_X1 g0859 ( .A1(new_n990_), .A2(new_n995_), .ZN(new_n996_) );
  NOR3_X1 g0860 ( .A1(new_n996_), .A2(new_n980_), .A3(new_n983_), .ZN(new_n997_) );
  NOR2_X1 g0861 ( .A1(new_n691_), .A2(new_n217_), .ZN(new_n998_) );
  INV_X1 g0862 ( .A(new_n998_), .ZN(new_n999_) );
  NAND2_X1 g0863 ( .A1(new_n700_), .A2(G150), .ZN(new_n1000_) );
  NAND2_X1 g0864 ( .A1(new_n695_), .A2(G58), .ZN(new_n1001_) );
  NAND2_X1 g0865 ( .A1(new_n723_), .A2(G50), .ZN(new_n1002_) );
  NOR2_X1 g0866 ( .A1(new_n718_), .A2(new_n140_), .ZN(new_n1003_) );
  INV_X1 g0867 ( .A(new_n1003_), .ZN(new_n1004_) );
  NAND2_X1 g0868 ( .A1(new_n725_), .A2(G159), .ZN(new_n1005_) );
  NAND3_X1 g0869 ( .A1(new_n1004_), .A2(new_n1002_), .A3(new_n1005_), .ZN(new_n1006_) );
  NOR2_X1 g0870 ( .A1(new_n703_), .A2(new_n409_), .ZN(new_n1007_) );
  NOR4_X1 g0871 ( .A1(new_n1006_), .A2(new_n713_), .A3(new_n919_), .A4(new_n1007_), .ZN(new_n1008_) );
  NAND4_X1 g0872 ( .A1(new_n1008_), .A2(new_n999_), .A3(new_n1000_), .A4(new_n1001_), .ZN(new_n1009_) );
  NAND2_X1 g0873 ( .A1(new_n1009_), .A2(new_n753_), .ZN(new_n1010_) );
  NOR2_X1 g0874 ( .A1(new_n1010_), .A2(new_n997_), .ZN(new_n1011_) );
  NAND3_X1 g0875 ( .A1(new_n961_), .A2(new_n976_), .A3(new_n1011_), .ZN(new_n1012_) );
  NAND2_X1 g0876 ( .A1(new_n960_), .A2(new_n1012_), .ZN(new_n1013_) );
  INV_X1 g0877 ( .A(new_n1013_), .ZN(new_n1014_) );
  NAND2_X1 g0878 ( .A1(new_n1014_), .A2(new_n959_), .ZN(G393) );
  NAND2_X1 g0879 ( .A1(new_n761_), .A2(new_n907_), .ZN(new_n1016_) );
  NAND3_X1 g0880 ( .A1(new_n1016_), .A2(new_n897_), .A3(new_n898_), .ZN(new_n1017_) );
  NAND3_X1 g0881 ( .A1(new_n1017_), .A2(new_n911_), .A3(new_n653_), .ZN(new_n1018_) );
  NAND3_X1 g0882 ( .A1(new_n912_), .A2(new_n752_), .A3(new_n899_), .ZN(new_n1019_) );
  NAND3_X1 g0883 ( .A1(new_n884_), .A2(new_n661_), .A3(new_n885_), .ZN(new_n1020_) );
  INV_X1 g0884 ( .A(KEYINPUT58), .ZN(new_n1021_) );
  NOR2_X1 g0885 ( .A1(new_n722_), .A2(new_n808_), .ZN(new_n1022_) );
  NAND2_X1 g0886 ( .A1(new_n690_), .A2(G116), .ZN(new_n1023_) );
  NAND2_X1 g0887 ( .A1(new_n700_), .A2(G322), .ZN(new_n1024_) );
  NAND2_X1 g0888 ( .A1(new_n695_), .A2(G303), .ZN(new_n1025_) );
  NAND2_X1 g0889 ( .A1(new_n702_), .A2(G294), .ZN(new_n1026_) );
  NAND4_X1 g0890 ( .A1(new_n1024_), .A2(new_n1023_), .A3(new_n1025_), .A4(new_n1026_), .ZN(new_n1027_) );
  NOR4_X1 g0891 ( .A1(new_n1027_), .A2(new_n255_), .A3(new_n715_), .A4(new_n1022_), .ZN(new_n1028_) );
  NAND2_X1 g0892 ( .A1(new_n1028_), .A2(new_n1021_), .ZN(new_n1029_) );
  INV_X1 g0893 ( .A(new_n1028_), .ZN(new_n1030_) );
  NAND2_X1 g0894 ( .A1(new_n1030_), .A2(KEYINPUT58), .ZN(new_n1031_) );
  NAND2_X1 g0895 ( .A1(new_n719_), .A2(G283), .ZN(new_n1032_) );
  NAND2_X1 g0896 ( .A1(new_n725_), .A2(G317), .ZN(new_n1033_) );
  NAND2_X1 g0897 ( .A1(new_n1032_), .A2(new_n1033_), .ZN(new_n1034_) );
  NAND2_X1 g0898 ( .A1(new_n1034_), .A2(KEYINPUT59), .ZN(new_n1035_) );
  INV_X1 g0899 ( .A(KEYINPUT59), .ZN(new_n1036_) );
  NAND3_X1 g0900 ( .A1(new_n1032_), .A2(new_n1036_), .A3(new_n1033_), .ZN(new_n1037_) );
  NAND2_X1 g0901 ( .A1(new_n1035_), .A2(new_n1037_), .ZN(new_n1038_) );
  NAND3_X1 g0902 ( .A1(new_n1031_), .A2(new_n1029_), .A3(new_n1038_), .ZN(new_n1039_) );
  NAND2_X1 g0903 ( .A1(new_n700_), .A2(G143), .ZN(new_n1040_) );
  NAND2_X1 g0904 ( .A1(new_n723_), .A2(G159), .ZN(new_n1041_) );
  NAND3_X1 g0905 ( .A1(new_n1040_), .A2(new_n255_), .A3(new_n1041_), .ZN(new_n1042_) );
  NAND2_X1 g0906 ( .A1(new_n695_), .A2(G50), .ZN(new_n1043_) );
  NAND2_X1 g0907 ( .A1(new_n702_), .A2(G58), .ZN(new_n1044_) );
  NAND2_X1 g0908 ( .A1(new_n690_), .A2(G77), .ZN(new_n1045_) );
  NAND3_X1 g0909 ( .A1(new_n1045_), .A2(new_n1043_), .A3(new_n1044_), .ZN(new_n1046_) );
  NOR2_X1 g0910 ( .A1(new_n1042_), .A2(new_n1046_), .ZN(new_n1047_) );
  INV_X1 g0911 ( .A(KEYINPUT57), .ZN(new_n1048_) );
  INV_X1 g0912 ( .A(KEYINPUT56), .ZN(new_n1049_) );
  NAND3_X1 g0913 ( .A1(new_n725_), .A2(G150), .A3(new_n1049_), .ZN(new_n1050_) );
  NAND2_X1 g0914 ( .A1(new_n725_), .A2(G150), .ZN(new_n1051_) );
  NAND2_X1 g0915 ( .A1(new_n1051_), .A2(KEYINPUT56), .ZN(new_n1052_) );
  NAND2_X1 g0916 ( .A1(new_n1052_), .A2(new_n1050_), .ZN(new_n1053_) );
  NAND2_X1 g0917 ( .A1(new_n719_), .A2(G68), .ZN(new_n1054_) );
  NAND2_X1 g0918 ( .A1(new_n1053_), .A2(new_n1054_), .ZN(new_n1055_) );
  NAND2_X1 g0919 ( .A1(new_n1055_), .A2(new_n1048_), .ZN(new_n1056_) );
  NAND3_X1 g0920 ( .A1(new_n1053_), .A2(KEYINPUT57), .A3(new_n1054_), .ZN(new_n1057_) );
  NAND4_X1 g0921 ( .A1(new_n1047_), .A2(new_n1056_), .A3(new_n807_), .A4(new_n1057_), .ZN(new_n1058_) );
  NAND2_X1 g0922 ( .A1(new_n1039_), .A2(new_n1058_), .ZN(new_n1059_) );
  NAND2_X1 g0923 ( .A1(new_n1059_), .A2(new_n712_), .ZN(new_n1060_) );
  NAND2_X1 g0924 ( .A1(new_n225_), .A2(new_n670_), .ZN(new_n1061_) );
  NAND2_X1 g0925 ( .A1(new_n652_), .A2(G97), .ZN(new_n1062_) );
  NAND3_X1 g0926 ( .A1(new_n1061_), .A2(new_n684_), .A3(new_n1062_), .ZN(new_n1063_) );
  NAND4_X1 g0927 ( .A1(new_n1020_), .A2(new_n753_), .A3(new_n1060_), .A4(new_n1063_), .ZN(new_n1064_) );
  NAND2_X1 g0928 ( .A1(new_n1019_), .A2(new_n1064_), .ZN(new_n1065_) );
  INV_X1 g0929 ( .A(new_n1065_), .ZN(new_n1066_) );
  NAND2_X1 g0930 ( .A1(new_n1018_), .A2(new_n1066_), .ZN(G390) );
  INV_X1 g0931 ( .A(KEYINPUT39), .ZN(new_n1068_) );
  INV_X1 g0932 ( .A(new_n848_), .ZN(new_n1069_) );
  NAND4_X1 g0933 ( .A1(new_n647_), .A2(new_n1069_), .A3(G330), .A4(new_n1068_), .ZN(new_n1070_) );
  NAND3_X1 g0934 ( .A1(new_n647_), .A2(new_n1069_), .A3(G330), .ZN(new_n1071_) );
  NAND2_X1 g0935 ( .A1(new_n1071_), .A2(KEYINPUT39), .ZN(new_n1072_) );
  NAND2_X1 g0936 ( .A1(new_n1072_), .A2(new_n1070_), .ZN(new_n1073_) );
  INV_X1 g0937 ( .A(new_n1073_), .ZN(new_n1074_) );
  INV_X1 g0938 ( .A(KEYINPUT40), .ZN(new_n1075_) );
  NAND2_X1 g0939 ( .A1(new_n841_), .A2(new_n1075_), .ZN(new_n1076_) );
  NAND2_X1 g0940 ( .A1(new_n840_), .A2(KEYINPUT40), .ZN(new_n1077_) );
  NAND2_X1 g0941 ( .A1(new_n1076_), .A2(new_n1077_), .ZN(new_n1078_) );
  INV_X1 g0942 ( .A(new_n1078_), .ZN(new_n1079_) );
  NAND4_X1 g0943 ( .A1(new_n833_), .A2(new_n1074_), .A3(new_n1079_), .A4(new_n834_), .ZN(new_n1080_) );
  NAND3_X1 g0944 ( .A1(new_n833_), .A2(new_n1074_), .A3(new_n834_), .ZN(new_n1081_) );
  NAND2_X1 g0945 ( .A1(new_n1081_), .A2(new_n1078_), .ZN(new_n1082_) );
  NAND2_X1 g0946 ( .A1(new_n1082_), .A2(new_n1080_), .ZN(new_n1083_) );
  NAND2_X1 g0947 ( .A1(new_n824_), .A2(new_n631_), .ZN(new_n1084_) );
  NAND2_X1 g0948 ( .A1(new_n821_), .A2(new_n769_), .ZN(new_n1085_) );
  NAND3_X1 g0949 ( .A1(new_n1084_), .A2(new_n832_), .A3(new_n1085_), .ZN(new_n1086_) );
  INV_X1 g0950 ( .A(new_n832_), .ZN(new_n1087_) );
  NAND2_X1 g0951 ( .A1(new_n1084_), .A2(new_n1085_), .ZN(new_n1088_) );
  NAND2_X1 g0952 ( .A1(new_n1088_), .A2(new_n1087_), .ZN(new_n1089_) );
  NAND2_X1 g0953 ( .A1(new_n1089_), .A2(new_n1086_), .ZN(new_n1090_) );
  NAND3_X1 g0954 ( .A1(new_n436_), .A2(G330), .A3(new_n647_), .ZN(new_n1091_) );
  NAND3_X1 g0955 ( .A1(new_n614_), .A2(new_n843_), .A3(new_n1091_), .ZN(new_n1092_) );
  NAND2_X1 g0956 ( .A1(new_n1092_), .A2(KEYINPUT38), .ZN(new_n1093_) );
  INV_X1 g0957 ( .A(KEYINPUT38), .ZN(new_n1094_) );
  NAND4_X1 g0958 ( .A1(new_n614_), .A2(new_n843_), .A3(new_n1094_), .A4(new_n1091_), .ZN(new_n1095_) );
  NAND2_X1 g0959 ( .A1(new_n1093_), .A2(new_n1095_), .ZN(new_n1096_) );
  INV_X1 g0960 ( .A(new_n1096_), .ZN(new_n1097_) );
  NAND3_X1 g0961 ( .A1(new_n1083_), .A2(new_n1090_), .A3(new_n1097_), .ZN(new_n1098_) );
  NAND2_X1 g0962 ( .A1(new_n1090_), .A2(new_n1097_), .ZN(new_n1099_) );
  NAND3_X1 g0963 ( .A1(new_n1099_), .A2(new_n1080_), .A3(new_n1082_), .ZN(new_n1100_) );
  NAND3_X1 g0964 ( .A1(new_n1100_), .A2(new_n653_), .A3(new_n1098_), .ZN(new_n1101_) );
  NAND2_X1 g0965 ( .A1(new_n1083_), .A2(new_n750_), .ZN(new_n1102_) );
  NAND2_X1 g0966 ( .A1(new_n840_), .A2(new_n659_), .ZN(new_n1103_) );
  NAND2_X1 g0967 ( .A1(new_n695_), .A2(G137), .ZN(new_n1104_) );
  NAND2_X1 g0968 ( .A1(new_n690_), .A2(G159), .ZN(new_n1105_) );
  NAND2_X1 g0969 ( .A1(new_n700_), .A2(G125), .ZN(new_n1106_) );
  NAND3_X1 g0970 ( .A1(new_n1106_), .A2(new_n1105_), .A3(new_n1104_), .ZN(new_n1107_) );
  NAND2_X1 g0971 ( .A1(new_n723_), .A2(G132), .ZN(new_n1108_) );
  NAND2_X1 g0972 ( .A1(new_n719_), .A2(G150), .ZN(new_n1109_) );
  NAND2_X1 g0973 ( .A1(new_n725_), .A2(G128), .ZN(new_n1110_) );
  NAND3_X1 g0974 ( .A1(new_n1108_), .A2(new_n1109_), .A3(new_n1110_), .ZN(new_n1111_) );
  NAND2_X1 g0975 ( .A1(new_n730_), .A2(G50), .ZN(new_n1112_) );
  NAND2_X1 g0976 ( .A1(new_n702_), .A2(G143), .ZN(new_n1113_) );
  NAND2_X1 g0977 ( .A1(new_n1112_), .A2(new_n1113_), .ZN(new_n1114_) );
  NOR4_X1 g0978 ( .A1(new_n1107_), .A2(new_n1111_), .A3(new_n1114_), .A4(new_n713_), .ZN(new_n1115_) );
  INV_X1 g0979 ( .A(KEYINPUT47), .ZN(new_n1116_) );
  NAND3_X1 g0980 ( .A1(new_n723_), .A2(G116), .A3(new_n1116_), .ZN(new_n1117_) );
  NAND2_X1 g0981 ( .A1(new_n723_), .A2(G116), .ZN(new_n1118_) );
  NAND2_X1 g0982 ( .A1(new_n1118_), .A2(KEYINPUT47), .ZN(new_n1119_) );
  NAND2_X1 g0983 ( .A1(new_n695_), .A2(G107), .ZN(new_n1120_) );
  NAND4_X1 g0984 ( .A1(new_n1119_), .A2(new_n1045_), .A3(new_n1117_), .A4(new_n1120_), .ZN(new_n1121_) );
  NAND2_X1 g0985 ( .A1(new_n725_), .A2(G283), .ZN(new_n1122_) );
  NAND4_X1 g0986 ( .A1(new_n917_), .A2(new_n720_), .A3(new_n776_), .A4(new_n1122_), .ZN(new_n1123_) );
  NAND2_X1 g0987 ( .A1(new_n700_), .A2(G294), .ZN(new_n1124_) );
  NAND2_X1 g0988 ( .A1(new_n702_), .A2(G97), .ZN(new_n1125_) );
  NAND2_X1 g0989 ( .A1(new_n1124_), .A2(new_n1125_), .ZN(new_n1126_) );
  NAND2_X1 g0990 ( .A1(new_n1126_), .A2(KEYINPUT48), .ZN(new_n1127_) );
  INV_X1 g0991 ( .A(KEYINPUT48), .ZN(new_n1128_) );
  NAND3_X1 g0992 ( .A1(new_n1124_), .A2(new_n1128_), .A3(new_n1125_), .ZN(new_n1129_) );
  NAND2_X1 g0993 ( .A1(new_n1127_), .A2(new_n1129_), .ZN(new_n1130_) );
  NOR3_X1 g0994 ( .A1(new_n1123_), .A2(new_n1130_), .A3(new_n1121_), .ZN(new_n1131_) );
  NAND2_X1 g0995 ( .A1(new_n815_), .A2(new_n265_), .ZN(new_n1132_) );
  NAND2_X1 g0996 ( .A1(new_n753_), .A2(new_n1132_), .ZN(new_n1133_) );
  NOR3_X1 g0997 ( .A1(new_n1131_), .A2(new_n1115_), .A3(new_n1133_), .ZN(new_n1134_) );
  NAND2_X1 g0998 ( .A1(new_n1103_), .A2(new_n1134_), .ZN(new_n1135_) );
  NAND2_X1 g0999 ( .A1(new_n1102_), .A2(new_n1135_), .ZN(new_n1136_) );
  INV_X1 g1000 ( .A(new_n1136_), .ZN(new_n1137_) );
  NAND2_X1 g1001 ( .A1(new_n1101_), .A2(new_n1137_), .ZN(G378) );
  NAND3_X1 g1002 ( .A1(new_n1083_), .A2(KEYINPUT41), .A3(new_n1090_), .ZN(new_n1139_) );
  INV_X1 g1003 ( .A(KEYINPUT41), .ZN(new_n1140_) );
  NAND2_X1 g1004 ( .A1(new_n1083_), .A2(new_n1090_), .ZN(new_n1141_) );
  NAND2_X1 g1005 ( .A1(new_n1141_), .A2(new_n1140_), .ZN(new_n1142_) );
  NAND2_X1 g1006 ( .A1(new_n1142_), .A2(new_n1139_), .ZN(new_n1143_) );
  NAND2_X1 g1007 ( .A1(new_n1097_), .A2(new_n751_), .ZN(new_n1144_) );
  INV_X1 g1008 ( .A(new_n1144_), .ZN(new_n1145_) );
  NAND2_X1 g1009 ( .A1(new_n1143_), .A2(new_n1145_), .ZN(new_n1146_) );
  NAND2_X1 g1010 ( .A1(new_n821_), .A2(new_n849_), .ZN(new_n1147_) );
  NAND3_X1 g1011 ( .A1(new_n842_), .A2(new_n822_), .A3(new_n1147_), .ZN(new_n1148_) );
  NAND2_X1 g1012 ( .A1(new_n369_), .A2(new_n836_), .ZN(new_n1149_) );
  NAND2_X1 g1013 ( .A1(new_n395_), .A2(new_n1149_), .ZN(new_n1150_) );
  NAND4_X1 g1014 ( .A1(new_n369_), .A2(new_n384_), .A3(new_n386_), .A4(new_n836_), .ZN(new_n1151_) );
  NAND2_X1 g1015 ( .A1(new_n1150_), .A2(new_n1151_), .ZN(new_n1152_) );
  NAND2_X1 g1016 ( .A1(new_n1148_), .A2(new_n1152_), .ZN(new_n1153_) );
  INV_X1 g1017 ( .A(new_n1153_), .ZN(new_n1154_) );
  INV_X1 g1018 ( .A(new_n1152_), .ZN(new_n1155_) );
  NAND4_X1 g1019 ( .A1(new_n842_), .A2(new_n822_), .A3(new_n1147_), .A4(new_n1155_), .ZN(new_n1156_) );
  INV_X1 g1020 ( .A(new_n1156_), .ZN(new_n1157_) );
  NOR3_X1 g1021 ( .A1(new_n1154_), .A2(new_n753_), .A3(new_n1157_), .ZN(new_n1158_) );
  NAND2_X1 g1022 ( .A1(new_n1146_), .A2(new_n1158_), .ZN(new_n1159_) );
  NAND2_X1 g1023 ( .A1(new_n1155_), .A2(new_n659_), .ZN(new_n1160_) );
  NAND3_X1 g1024 ( .A1(new_n702_), .A2(G137), .A3(KEYINPUT43), .ZN(new_n1161_) );
  INV_X1 g1025 ( .A(KEYINPUT43), .ZN(new_n1162_) );
  NAND2_X1 g1026 ( .A1(new_n702_), .A2(G137), .ZN(new_n1163_) );
  NAND2_X1 g1027 ( .A1(new_n1163_), .A2(new_n1162_), .ZN(new_n1164_) );
  NAND2_X1 g1028 ( .A1(new_n1164_), .A2(new_n1161_), .ZN(new_n1165_) );
  NAND2_X1 g1029 ( .A1(new_n723_), .A2(G128), .ZN(new_n1166_) );
  NAND2_X1 g1030 ( .A1(new_n719_), .A2(G143), .ZN(new_n1167_) );
  NAND2_X1 g1031 ( .A1(new_n725_), .A2(G125), .ZN(new_n1168_) );
  NAND3_X1 g1032 ( .A1(new_n1166_), .A2(new_n1167_), .A3(new_n1168_), .ZN(new_n1169_) );
  NAND2_X1 g1033 ( .A1(new_n690_), .A2(G150), .ZN(new_n1170_) );
  NAND2_X1 g1034 ( .A1(new_n700_), .A2(G124), .ZN(new_n1171_) );
  NAND2_X1 g1035 ( .A1(new_n1171_), .A2(new_n1170_), .ZN(new_n1172_) );
  NOR2_X1 g1036 ( .A1(new_n1169_), .A2(new_n1172_), .ZN(new_n1173_) );
  NAND2_X1 g1037 ( .A1(new_n730_), .A2(G159), .ZN(new_n1174_) );
  NAND2_X1 g1038 ( .A1(new_n695_), .A2(G132), .ZN(new_n1175_) );
  NAND2_X1 g1039 ( .A1(new_n1174_), .A2(new_n1175_), .ZN(new_n1176_) );
  NAND2_X1 g1040 ( .A1(new_n1176_), .A2(KEYINPUT44), .ZN(new_n1177_) );
  INV_X1 g1041 ( .A(KEYINPUT44), .ZN(new_n1178_) );
  NAND3_X1 g1042 ( .A1(new_n1174_), .A2(new_n1178_), .A3(new_n1175_), .ZN(new_n1179_) );
  NAND4_X1 g1043 ( .A1(new_n1173_), .A2(new_n1177_), .A3(new_n1165_), .A4(new_n1179_), .ZN(new_n1180_) );
  NAND2_X1 g1044 ( .A1(new_n1180_), .A2(new_n255_), .ZN(new_n1181_) );
  NOR2_X1 g1045 ( .A1(new_n714_), .A2(new_n265_), .ZN(new_n1182_) );
  INV_X1 g1046 ( .A(KEYINPUT42), .ZN(new_n1183_) );
  NOR3_X1 g1047 ( .A1(new_n722_), .A2(new_n439_), .A3(new_n1183_), .ZN(new_n1184_) );
  NOR2_X1 g1048 ( .A1(new_n722_), .A2(new_n439_), .ZN(new_n1185_) );
  NOR2_X1 g1049 ( .A1(new_n1185_), .A2(KEYINPUT42), .ZN(new_n1186_) );
  NOR2_X1 g1050 ( .A1(new_n703_), .A2(new_n217_), .ZN(new_n1187_) );
  NOR4_X1 g1051 ( .A1(new_n1186_), .A2(new_n1187_), .A3(new_n1184_), .A4(new_n1182_), .ZN(new_n1188_) );
  INV_X1 g1052 ( .A(new_n725_), .ZN(new_n1189_) );
  NOR2_X1 g1053 ( .A1(new_n1189_), .A2(new_n219_), .ZN(new_n1190_) );
  NOR3_X1 g1054 ( .A1(new_n934_), .A2(new_n1003_), .A3(new_n1190_), .ZN(new_n1191_) );
  NAND2_X1 g1055 ( .A1(new_n700_), .A2(G283), .ZN(new_n1192_) );
  NAND2_X1 g1056 ( .A1(new_n695_), .A2(G97), .ZN(new_n1193_) );
  NAND4_X1 g1057 ( .A1(new_n1188_), .A2(new_n1191_), .A3(new_n1192_), .A4(new_n1193_), .ZN(new_n1194_) );
  NAND2_X1 g1058 ( .A1(new_n1194_), .A2(G33), .ZN(new_n1195_) );
  NAND4_X1 g1059 ( .A1(new_n1195_), .A2(new_n290_), .A3(new_n1181_), .A4(new_n712_), .ZN(new_n1196_) );
  NAND2_X1 g1060 ( .A1(new_n712_), .A2(new_n290_), .ZN(new_n1197_) );
  NAND3_X1 g1061 ( .A1(new_n1197_), .A2(new_n139_), .A3(new_n660_), .ZN(new_n1198_) );
  NAND4_X1 g1062 ( .A1(new_n1160_), .A2(new_n753_), .A3(new_n1196_), .A4(new_n1198_), .ZN(new_n1199_) );
  NAND2_X1 g1063 ( .A1(new_n1159_), .A2(new_n1199_), .ZN(G375) );
  INV_X1 g1064 ( .A(KEYINPUT46), .ZN(new_n1201_) );
  NAND3_X1 g1065 ( .A1(new_n1096_), .A2(new_n1086_), .A3(new_n1089_), .ZN(new_n1202_) );
  NAND2_X1 g1066 ( .A1(new_n1099_), .A2(new_n1202_), .ZN(new_n1203_) );
  NAND2_X1 g1067 ( .A1(new_n1203_), .A2(new_n1201_), .ZN(new_n1204_) );
  NAND3_X1 g1068 ( .A1(new_n1099_), .A2(KEYINPUT46), .A3(new_n1202_), .ZN(new_n1205_) );
  NAND2_X1 g1069 ( .A1(new_n1204_), .A2(new_n1205_), .ZN(new_n1206_) );
  NAND2_X1 g1070 ( .A1(new_n1206_), .A2(new_n653_), .ZN(new_n1207_) );
  NAND2_X1 g1071 ( .A1(new_n1090_), .A2(new_n750_), .ZN(new_n1208_) );
  NAND2_X1 g1072 ( .A1(new_n1087_), .A2(new_n659_), .ZN(new_n1209_) );
  NAND2_X1 g1073 ( .A1(new_n690_), .A2(G50), .ZN(new_n1210_) );
  NAND2_X1 g1074 ( .A1(new_n700_), .A2(G128), .ZN(new_n1211_) );
  NAND2_X1 g1075 ( .A1(new_n702_), .A2(G150), .ZN(new_n1212_) );
  NAND2_X1 g1076 ( .A1(new_n723_), .A2(G137), .ZN(new_n1213_) );
  NAND2_X1 g1077 ( .A1(new_n719_), .A2(G159), .ZN(new_n1214_) );
  NAND2_X1 g1078 ( .A1(new_n725_), .A2(G132), .ZN(new_n1215_) );
  NAND3_X1 g1079 ( .A1(new_n1213_), .A2(new_n1214_), .A3(new_n1215_), .ZN(new_n1216_) );
  INV_X1 g1080 ( .A(G143), .ZN(new_n1217_) );
  NOR2_X1 g1081 ( .A1(new_n696_), .A2(new_n1217_), .ZN(new_n1218_) );
  NOR4_X1 g1082 ( .A1(new_n1216_), .A2(new_n713_), .A3(new_n1182_), .A4(new_n1218_), .ZN(new_n1219_) );
  NAND4_X1 g1083 ( .A1(new_n1219_), .A2(new_n1210_), .A3(new_n1211_), .A4(new_n1212_), .ZN(new_n1220_) );
  NOR2_X1 g1084 ( .A1(new_n696_), .A2(new_n219_), .ZN(new_n1221_) );
  NOR2_X1 g1085 ( .A1(new_n699_), .A2(new_n930_), .ZN(new_n1222_) );
  NOR2_X1 g1086 ( .A1(new_n703_), .A2(new_n439_), .ZN(new_n1223_) );
  NOR3_X1 g1087 ( .A1(new_n1221_), .A2(new_n1223_), .A3(new_n1222_), .ZN(new_n1224_) );
  NOR2_X1 g1088 ( .A1(new_n722_), .A2(new_n810_), .ZN(new_n1225_) );
  NAND2_X1 g1089 ( .A1(new_n719_), .A2(G97), .ZN(new_n1226_) );
  NAND2_X1 g1090 ( .A1(new_n725_), .A2(G294), .ZN(new_n1227_) );
  NAND2_X1 g1091 ( .A1(new_n1226_), .A2(new_n1227_), .ZN(new_n1228_) );
  NOR4_X1 g1092 ( .A1(new_n998_), .A2(new_n1228_), .A3(new_n935_), .A4(new_n1225_), .ZN(new_n1229_) );
  NAND3_X1 g1093 ( .A1(new_n1229_), .A2(new_n917_), .A3(new_n1224_), .ZN(new_n1230_) );
  NAND2_X1 g1094 ( .A1(new_n815_), .A2(new_n409_), .ZN(new_n1231_) );
  INV_X1 g1095 ( .A(new_n1231_), .ZN(new_n1232_) );
  NOR2_X1 g1096 ( .A1(new_n1232_), .A2(new_n752_), .ZN(new_n1233_) );
  NAND3_X1 g1097 ( .A1(new_n1220_), .A2(new_n1230_), .A3(new_n1233_), .ZN(new_n1234_) );
  NAND2_X1 g1098 ( .A1(new_n1234_), .A2(KEYINPUT45), .ZN(new_n1235_) );
  INV_X1 g1099 ( .A(KEYINPUT45), .ZN(new_n1236_) );
  NAND4_X1 g1100 ( .A1(new_n1220_), .A2(new_n1236_), .A3(new_n1230_), .A4(new_n1233_), .ZN(new_n1237_) );
  NAND2_X1 g1101 ( .A1(new_n1235_), .A2(new_n1237_), .ZN(new_n1238_) );
  NAND2_X1 g1102 ( .A1(new_n1209_), .A2(new_n1238_), .ZN(new_n1239_) );
  NAND2_X1 g1103 ( .A1(new_n1208_), .A2(new_n1239_), .ZN(new_n1240_) );
  INV_X1 g1104 ( .A(new_n1240_), .ZN(new_n1241_) );
  NAND2_X1 g1105 ( .A1(new_n1207_), .A2(new_n1241_), .ZN(G381) );
  INV_X1 g1106 ( .A(G378), .ZN(new_n1243_) );
  NAND3_X1 g1107 ( .A1(new_n1159_), .A2(new_n1243_), .A3(new_n1199_), .ZN(new_n1244_) );
  INV_X1 g1108 ( .A(new_n1244_), .ZN(new_n1245_) );
  INV_X1 g1109 ( .A(G396), .ZN(new_n1246_) );
  NAND3_X1 g1110 ( .A1(new_n1018_), .A2(new_n1246_), .A3(new_n1066_), .ZN(new_n1247_) );
  NAND4_X1 g1111 ( .A1(new_n1014_), .A2(new_n774_), .A3(new_n819_), .A4(new_n959_), .ZN(new_n1248_) );
  NOR4_X1 g1112 ( .A1(G387), .A2(G381), .A3(new_n1247_), .A4(new_n1248_), .ZN(new_n1249_) );
  NAND2_X1 g1113 ( .A1(new_n1249_), .A2(new_n1245_), .ZN(G407) );
  NAND2_X1 g1114 ( .A1(new_n1245_), .A2(new_n616_), .ZN(new_n1251_) );
  NAND3_X1 g1115 ( .A1(G407), .A2(G213), .A3(new_n1251_), .ZN(G409) );
  NAND2_X1 g1116 ( .A1(G375), .A2(G378), .ZN(new_n1253_) );
  NAND2_X1 g1117 ( .A1(new_n616_), .A2(G213), .ZN(new_n1254_) );
  NAND3_X1 g1118 ( .A1(new_n1253_), .A2(new_n1244_), .A3(new_n1254_), .ZN(new_n1255_) );
  NAND3_X1 g1119 ( .A1(new_n616_), .A2(G213), .A3(G2897), .ZN(new_n1256_) );
  NAND2_X1 g1120 ( .A1(new_n1256_), .A2(KEYINPUT63), .ZN(new_n1257_) );
  INV_X1 g1121 ( .A(KEYINPUT63), .ZN(new_n1258_) );
  NAND4_X1 g1122 ( .A1(new_n616_), .A2(new_n1258_), .A3(G213), .A4(G2897), .ZN(new_n1259_) );
  NAND2_X1 g1123 ( .A1(new_n1257_), .A2(new_n1259_), .ZN(new_n1260_) );
  INV_X1 g1124 ( .A(new_n1260_), .ZN(new_n1261_) );
  NAND2_X1 g1125 ( .A1(G390), .A2(G396), .ZN(new_n1262_) );
  NAND2_X1 g1126 ( .A1(new_n1262_), .A2(new_n1247_), .ZN(new_n1263_) );
  INV_X1 g1127 ( .A(new_n1263_), .ZN(new_n1264_) );
  NAND2_X1 g1128 ( .A1(G381), .A2(new_n1264_), .ZN(new_n1265_) );
  NAND3_X1 g1129 ( .A1(new_n1207_), .A2(new_n1263_), .A3(new_n1241_), .ZN(new_n1266_) );
  NAND2_X1 g1130 ( .A1(G393), .A2(G384), .ZN(new_n1267_) );
  NAND2_X1 g1131 ( .A1(new_n1267_), .A2(new_n1248_), .ZN(new_n1268_) );
  INV_X1 g1132 ( .A(new_n1268_), .ZN(new_n1269_) );
  NAND2_X1 g1133 ( .A1(new_n957_), .A2(new_n1269_), .ZN(new_n1270_) );
  NAND3_X1 g1134 ( .A1(new_n954_), .A2(new_n956_), .A3(new_n1268_), .ZN(new_n1271_) );
  NAND4_X1 g1135 ( .A1(new_n1265_), .A2(new_n1270_), .A3(new_n1266_), .A4(new_n1271_), .ZN(new_n1272_) );
  NAND2_X1 g1136 ( .A1(new_n1265_), .A2(new_n1266_), .ZN(new_n1273_) );
  NAND2_X1 g1137 ( .A1(new_n1270_), .A2(new_n1271_), .ZN(new_n1274_) );
  NAND2_X1 g1138 ( .A1(new_n1273_), .A2(new_n1274_), .ZN(new_n1275_) );
  NAND4_X1 g1139 ( .A1(new_n1275_), .A2(new_n1255_), .A3(new_n1261_), .A4(new_n1272_), .ZN(new_n1276_) );
  NAND2_X1 g1140 ( .A1(new_n1255_), .A2(new_n1261_), .ZN(new_n1277_) );
  NAND2_X1 g1141 ( .A1(new_n1275_), .A2(new_n1272_), .ZN(new_n1278_) );
  NAND2_X1 g1142 ( .A1(new_n1278_), .A2(new_n1277_), .ZN(new_n1279_) );
  NAND2_X1 g1143 ( .A1(new_n1279_), .A2(new_n1276_), .ZN(G405) );
  NAND2_X1 g1144 ( .A1(new_n1253_), .A2(new_n1244_), .ZN(new_n1281_) );
  NAND3_X1 g1145 ( .A1(new_n1275_), .A2(new_n1281_), .A3(new_n1272_), .ZN(new_n1282_) );
  INV_X1 g1146 ( .A(new_n1281_), .ZN(new_n1283_) );
  NAND2_X1 g1147 ( .A1(new_n1278_), .A2(new_n1283_), .ZN(new_n1284_) );
  NAND2_X1 g1148 ( .A1(new_n1284_), .A2(new_n1282_), .ZN(G402) );
endmodule


