module rs232 ( sys_clk, sys_rst_l, uart_XMIT_dataH, xmitH, xmit_dataH_7_, 
        xmit_dataH_6_, xmit_dataH_5_, xmit_dataH_4_, xmit_dataH_3_, 
        xmit_dataH_2_, xmit_dataH_1_, xmit_dataH_0_, xmit_doneH, 
        uart_REC_dataH, rec_dataH_7_, rec_dataH_6_, rec_dataH_5_, rec_dataH_4_, 
        rec_dataH_3_, rec_dataH_2_, rec_dataH_1_, rec_dataH_0_, rec_readyH, 
        test_mode, test_se, test_si, test_so );
  input sys_clk, sys_rst_l, xmitH, xmit_dataH_7_, xmit_dataH_6_, xmit_dataH_5_,
         xmit_dataH_4_, xmit_dataH_3_, xmit_dataH_2_, xmit_dataH_1_,
         xmit_dataH_0_, uart_REC_dataH, test_mode, test_se, test_si;
  output uart_XMIT_dataH, xmit_doneH, rec_dataH_7_, rec_dataH_6_, rec_dataH_5_,
         rec_dataH_4_, rec_dataH_3_, rec_dataH_2_, rec_dataH_1_, rec_dataH_0_,
         rec_readyH, test_so;
  wire   iCTRL, iXMIT_state_1_temp, iXMIT_state_1_, iXMIT_CRTL, iRECEIVER_CTRL,
         iRECEIVER_state_CTRL, iRECEIVER_N_CTRL_1_, iRECEIVER_N_CTRL_2_,
         iRECEIVER_bitCell_CTRL, iRECEIVER_N18, iRECEIVER_N17,
         iRECEIVER_bitCell_cntrH_0_, iRECEIVER_bitCell_cntrH_1_, iRECEIVER_N22,
         iRECEIVER_N21, iRECEIVER_N20, iRECEIVER_N19, iRECEIVER_N28,
         iRECEIVER_N27, iRECEIVER_N26, iRECEIVER_N23, iRECEIVER_state_0_,
         iRECEIVER_state_1_, iRECEIVER_state_2_, iXMIT_N_CTRL_1_,
         iXMIT_N_CTRL_2_, iXMIT_xmit_CTRL, iXMIT_N24, iXMIT_xmit_ShiftRegH_7_,
         iXMIT_xmit_ShiftRegH_6_, iXMIT_xmit_ShiftRegH_5_, iXMIT_N28,
         iXMIT_N27, iXMIT_N26, iXMIT_N25, n401, n239, n242, n246, n255, n241,
         n244, n245, n238, n258, n259, rec_dataH_rec_7, rec_dataH_rec_6,
         rec_dataH_rec_5, rec_dataH_rec_4, rec_dataH_rec_3, rec_dataH_rec_2,
         rec_dataH_rec_1, rec_dataH_rec_0, n182, n181, n180, n179, n178, n177,
         n176, n175, n174, n173, n172, n171, n170, n169, n168, n167, n166,
         n164, n163, n162, n161, n160, n159, n157, n156, n155, test_point_DOUT,
         rec_dataH_temp_6_, rec_dataH_temp_5_, rec_dataH_temp_4_,
         rec_dataH_temp_3_, rec_dataH_temp_2_, rec_dataH_temp_1_,
         rec_dataH_temp_0_, n154, n153, n152, n150, n149, n148, n147, n146,
         n145, n143, n142, n141, n140, n139, n138, n136, n135, n134, n133,
         n132, n131, n129, n128, n127, n126, n125, n124, n122, n121, n120,
         n119, n118, n17, n424, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784;

  AND2X4 TrojanU305 ( .IN1(iCTRL), .IN2(iXMIT_state_1_temp), .Q(iXMIT_state_1_) );
  OR2X1 TrojanU302 ( .IN1(iXMIT_CRTL), .IN2(iRECEIVER_CTRL), .Q(iCTRL) );
  OR4X4 TrojanU301 ( .IN1(iRECEIVER_state_CTRL), .IN2(iRECEIVER_N_CTRL_1_), 
        .IN3(iRECEIVER_N_CTRL_2_), .IN4(iRECEIVER_bitCell_CTRL), .Q(
        iRECEIVER_CTRL) );
  NAND4X1 TrojanU300 ( .IN1(iRECEIVER_N18), .IN2(iRECEIVER_N17), .IN3(
        iRECEIVER_bitCell_cntrH_0_), .IN4(iRECEIVER_bitCell_cntrH_1_), .QN(
        iRECEIVER_bitCell_CTRL) );
  NAND4X1 TrojanU299 ( .IN1(iRECEIVER_N22), .IN2(iRECEIVER_N21), .IN3(
        iRECEIVER_N20), .IN4(iRECEIVER_N19), .QN(iRECEIVER_N_CTRL_2_) );
  NAND4X1 TrojanU298 ( .IN1(iRECEIVER_N28), .IN2(iRECEIVER_N27), .IN3(
        iRECEIVER_N26), .IN4(iRECEIVER_N23), .QN(iRECEIVER_N_CTRL_1_) );
  NAND4X1 TrojanU297 ( .IN1(n17), .IN2(iRECEIVER_state_0_), .IN3(
        iRECEIVER_state_1_), .IN4(iRECEIVER_state_2_), .QN(
        iRECEIVER_state_CTRL) );
  OR4X4 TrojanU296 ( .IN1(1'b0), .IN2(iXMIT_N_CTRL_1_), .IN3(iXMIT_N_CTRL_2_), 
        .IN4(iXMIT_xmit_CTRL), .Q(iXMIT_CRTL) );
  NAND4X1 TrojanU295 ( .IN1(iXMIT_N24), .IN2(iXMIT_xmit_ShiftRegH_7_), .IN3(
        iXMIT_xmit_ShiftRegH_6_), .IN4(iXMIT_xmit_ShiftRegH_5_), .QN(
        iXMIT_xmit_CTRL) );
  NAND4X1 TrojanU294 ( .IN1(iXMIT_N28), .IN2(iXMIT_N27), .IN3(iXMIT_N26), 
        .IN4(iXMIT_N25), .QN(iXMIT_N_CTRL_2_) );
  NAND4X1 TrojanU293 ( .IN1(n401), .IN2(n239), .IN3(n242), .IN4(n246), .QN(
        iXMIT_N_CTRL_1_) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_2_ ( .D(n182), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n781) );
  DFFARX1 iXMIT_state_reg_0_ ( .D(n181), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        n762), .QN(n239) );
  DFFARX1 iXMIT_state_reg_2_ ( .D(n180), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        n777), .QN(n242) );
  DFFARX1 iXMIT_state_reg_1_ ( .D(n179), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        iXMIT_state_1_temp), .QN(n246) );
  DFFARX1 iXMIT_bitCountH_reg_0_ ( .D(n178), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n771), .QN(n444) );
  DFFARX1 iXMIT_bitCountH_reg_1_ ( .D(n177), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n763) );
  DFFARX1 iXMIT_bitCountH_reg_2_ ( .D(n176), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n772), .QN(n449) );
  DFFARX1 iXMIT_bitCountH_reg_3_ ( .D(n175), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n764), .QN(n434) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_7_ ( .D(n174), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_xmit_ShiftRegH_7_), .QN(n424) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_6_ ( .D(n173), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_xmit_ShiftRegH_6_), .QN(n258) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_5_ ( .D(n172), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_xmit_ShiftRegH_5_), .QN(n259) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_4_ ( .D(n171), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n773), .QN(n445) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_3_ ( .D(n170), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n774), .QN(n446) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_2_ ( .D(n169), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n775), .QN(n447) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_1_ ( .D(n168), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n776), .QN(n448) );
  DFFARX1 iXMIT_xmit_doneH_reg ( .D(n167), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(xmit_doneH) );
  DFFARX1 iRECEIVER_state_reg_1_ ( .D(n166), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(iRECEIVER_state_1_), .QN(n241) );
  DFFASX1 iRECEIVER_state_reg_0_ ( .D(n164), .CLK(sys_clk), .SETB(sys_rst_l), 
        .Q(iRECEIVER_state_0_), .QN(n245) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_0_ ( .D(n163), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iRECEIVER_bitCell_cntrH_0_), .QN(n255) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_1_ ( .D(n162), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iRECEIVER_bitCell_cntrH_1_), .QN(n244) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_2_ ( .D(n161), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n784) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_3_ ( .D(n160), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n765) );
  DFFARX1 iRECEIVER_state_reg_2_ ( .D(n159), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(iRECEIVER_state_2_), .QN(n238) );
  DFFARX1 iRECEIVER_rec_readyH_reg ( .D(n157), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(rec_readyH) );
  DFFARX1 iRECEIVER_par_dataH_reg_7_ ( .D(n156), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_7), .QN(n436) );
  DFFARX1 rec_dataH_temp_reg_7_ ( .D(n155), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(test_so) );
  DFFARX1 rec_dataH_reg_7_ ( .D(n154), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_7_) );
  DFFARX1 iRECEIVER_par_dataH_reg_6_ ( .D(n153), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_6), .QN(n438) );
  DFFARX1 rec_dataH_temp_reg_6_ ( .D(n152), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_6_) );
  DFFARX1 rec_dataH_reg_6_ ( .D(n150), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_6_) );
  DFFARX1 iRECEIVER_par_dataH_reg_5_ ( .D(n149), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_5), .QN(n439) );
  DFFARX1 rec_dataH_temp_reg_5_ ( .D(n148), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_5_) );
  DFFARX1 rec_dataH_reg_5_ ( .D(n147), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_5_) );
  DFFARX1 iRECEIVER_par_dataH_reg_4_ ( .D(n146), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_4), .QN(n440) );
  DFFARX1 rec_dataH_temp_reg_4_ ( .D(n145), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_4_) );
  DFFARX1 rec_dataH_reg_4_ ( .D(n143), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_4_) );
  DFFARX1 iRECEIVER_par_dataH_reg_3_ ( .D(n142), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_3), .QN(n441) );
  DFFARX1 rec_dataH_temp_reg_3_ ( .D(n141), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_3_) );
  DFFARX1 rec_dataH_reg_3_ ( .D(n140), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_3_) );
  DFFARX1 iRECEIVER_par_dataH_reg_2_ ( .D(n139), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_2), .QN(n442) );
  DFFARX1 rec_dataH_temp_reg_2_ ( .D(n138), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_2_) );
  DFFARX1 rec_dataH_reg_2_ ( .D(n136), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_2_) );
  DFFARX1 iRECEIVER_par_dataH_reg_1_ ( .D(n135), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_1), .QN(n443) );
  DFFARX1 rec_dataH_temp_reg_1_ ( .D(n134), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_1_) );
  DFFARX1 rec_dataH_reg_1_ ( .D(n133), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_1_) );
  DFFARX1 iRECEIVER_par_dataH_reg_0_ ( .D(n132), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_0) );
  DFFARX1 rec_dataH_temp_reg_0_ ( .D(n131), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_0_) );
  DFFARX1 rec_dataH_reg_0_ ( .D(n129), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_0_) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_3_ ( .D(n128), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n766), .QN(n433) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_0_ ( .D(n127), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n767), .QN(n437) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_1_ ( .D(n126), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n783), .QN(n432) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_2_ ( .D(n125), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n782), .QN(n429) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_3_ ( .D(n124), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n780) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_0_ ( .D(n122), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n779), .QN(n430) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_1_ ( .D(n121), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n778), .QN(n435) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_0_ ( .D(n120), .CLK(sys_clk), .RSTB(
        sys_rst_l), .QN(n768) );
  DFFASX1 iRECEIVER_rec_datSyncH_reg ( .D(n119), .CLK(sys_clk), .SETB(
        sys_rst_l), .Q(n769) );
  DFFASX1 iRECEIVER_rec_datH_reg ( .D(n118), .CLK(sys_clk), .SETB(sys_rst_l), 
        .Q(n770), .QN(n431) );
  DFFARX1 TrojaniDatasend_reg_2_ ( .D(n182), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .QN(n401) );
  NAND2X0 U582 ( .IN1(n450), .IN2(n451), .QN(uart_XMIT_dataH) );
  OR2X1 U583 ( .IN1(n777), .IN2(iXMIT_state_1_), .Q(n451) );
  NOR2X0 U584 ( .IN1(n452), .IN2(n453), .QN(n450) );
  NOR2X0 U585 ( .IN1(n768), .IN2(n454), .QN(n453) );
  NOR2X0 U586 ( .IN1(n777), .IN2(n762), .QN(n454) );
  NAND2X0 U587 ( .IN1(n455), .IN2(n456), .QN(test_point_DOUT) );
  NAND2X0 U588 ( .IN1(rec_readyH), .IN2(n457), .QN(n456) );
  INVX0 U589 ( .INP(test_mode), .ZN(n457) );
  NAND2X0 U590 ( .IN1(sys_clk), .IN2(test_mode), .QN(n455) );
  NAND2X0 U591 ( .IN1(n458), .IN2(n459), .QN(n182) );
  NAND2X0 U592 ( .IN1(iXMIT_N28), .IN2(n460), .QN(n459) );
  NAND2X0 U593 ( .IN1(test_se), .IN2(n778), .QN(n458) );
  NAND2X0 U594 ( .IN1(n461), .IN2(n462), .QN(n181) );
  NAND2X0 U595 ( .IN1(n764), .IN2(test_se), .QN(n462) );
  NAND2X0 U596 ( .IN1(n463), .IN2(n460), .QN(n461) );
  NAND2X0 U597 ( .IN1(n464), .IN2(n465), .QN(n463) );
  NAND2X0 U598 ( .IN1(n777), .IN2(n466), .QN(n465) );
  NOR2X0 U599 ( .IN1(n467), .IN2(n468), .QN(n464) );
  NOR2X0 U600 ( .IN1(n239), .IN2(n469), .QN(n468) );
  NAND2X0 U601 ( .IN1(n470), .IN2(iXMIT_state_1_temp), .QN(n469) );
  NOR2X0 U602 ( .IN1(n762), .IN2(n471), .QN(n467) );
  NOR2X0 U603 ( .IN1(n472), .IN2(n777), .QN(n471) );
  NOR2X0 U604 ( .IN1(n246), .IN2(n466), .QN(n472) );
  NAND2X0 U605 ( .IN1(n473), .IN2(n474), .QN(n180) );
  NAND2X0 U606 ( .IN1(n475), .IN2(n452), .QN(n474) );
  NOR2X0 U607 ( .IN1(test_se), .IN2(n476), .QN(n475) );
  NAND2X0 U608 ( .IN1(n477), .IN2(iXMIT_state_1_temp), .QN(n473) );
  NAND2X0 U609 ( .IN1(n460), .IN2(n478), .QN(n477) );
  NAND2X0 U610 ( .IN1(n479), .IN2(n480), .QN(n179) );
  NAND2X0 U611 ( .IN1(test_se), .IN2(n762), .QN(n480) );
  NAND2X0 U612 ( .IN1(n481), .IN2(n460), .QN(n479) );
  NAND2X0 U613 ( .IN1(n482), .IN2(n483), .QN(n481) );
  INVX0 U614 ( .INP(n484), .ZN(n482) );
  NAND2X0 U615 ( .IN1(n485), .IN2(n486), .QN(n178) );
  NAND2X0 U616 ( .IN1(n780), .IN2(test_se), .QN(n486) );
  NAND2X0 U617 ( .IN1(n487), .IN2(n460), .QN(n485) );
  NAND2X0 U618 ( .IN1(n488), .IN2(n489), .QN(n487) );
  NAND2X0 U619 ( .IN1(n771), .IN2(n490), .QN(n489) );
  NAND2X0 U620 ( .IN1(n491), .IN2(n492), .QN(n177) );
  NAND2X0 U621 ( .IN1(n493), .IN2(n763), .QN(n492) );
  AND2X1 U622 ( .IN1(n460), .IN2(n494), .Q(n493) );
  NAND2X0 U623 ( .IN1(n771), .IN2(n495), .QN(n491) );
  NAND2X0 U624 ( .IN1(n460), .IN2(n496), .QN(n495) );
  OR2X1 U625 ( .IN1(n497), .IN2(n763), .Q(n496) );
  NAND2X0 U626 ( .IN1(n498), .IN2(n499), .QN(n176) );
  NAND2X0 U627 ( .IN1(n500), .IN2(n772), .QN(n499) );
  NOR2X0 U628 ( .IN1(test_se), .IN2(n501), .QN(n500) );
  NOR2X0 U629 ( .IN1(n502), .IN2(n490), .QN(n501) );
  INVX0 U630 ( .INP(n503), .ZN(n490) );
  NOR2X0 U631 ( .IN1(n763), .IN2(n497), .QN(n502) );
  NAND2X0 U632 ( .IN1(n763), .IN2(n504), .QN(n498) );
  NAND2X0 U633 ( .IN1(n505), .IN2(n460), .QN(n504) );
  NOR2X0 U634 ( .IN1(n506), .IN2(n507), .QN(n505) );
  NOR2X0 U635 ( .IN1(n449), .IN2(n488), .QN(n507) );
  NOR2X0 U636 ( .IN1(n772), .IN2(n508), .QN(n506) );
  NAND2X0 U637 ( .IN1(n509), .IN2(n771), .QN(n508) );
  NAND2X0 U638 ( .IN1(n510), .IN2(n511), .QN(n175) );
  NAND2X0 U639 ( .IN1(n772), .IN2(test_se), .QN(n511) );
  NAND2X0 U640 ( .IN1(n512), .IN2(n460), .QN(n510) );
  NAND2X0 U641 ( .IN1(n513), .IN2(n514), .QN(n512) );
  NAND2X0 U642 ( .IN1(n515), .IN2(n509), .QN(n514) );
  NOR2X0 U643 ( .IN1(n516), .IN2(n517), .QN(n515) );
  NOR2X0 U644 ( .IN1(n764), .IN2(n518), .QN(n517) );
  NOR2X0 U645 ( .IN1(n444), .IN2(n519), .QN(n518) );
  NOR2X0 U646 ( .IN1(n434), .IN2(n519), .QN(n516) );
  NAND2X0 U647 ( .IN1(n772), .IN2(n763), .QN(n519) );
  NAND2X0 U648 ( .IN1(n764), .IN2(n494), .QN(n513) );
  NAND2X0 U649 ( .IN1(n503), .IN2(n488), .QN(n494) );
  NAND2X0 U650 ( .IN1(n509), .IN2(n444), .QN(n488) );
  NAND2X0 U651 ( .IN1(n497), .IN2(n520), .QN(n503) );
  INVX0 U652 ( .INP(n509), .ZN(n497) );
  NOR2X0 U653 ( .IN1(n521), .IN2(n470), .QN(n509) );
  NAND2X0 U654 ( .IN1(n522), .IN2(n523), .QN(n470) );
  NAND2X0 U655 ( .IN1(n524), .IN2(n525), .QN(n523) );
  NOR2X0 U656 ( .IN1(n763), .IN2(n771), .QN(n525) );
  NOR2X0 U657 ( .IN1(n772), .IN2(n434), .QN(n524) );
  NAND2X0 U658 ( .IN1(iXMIT_state_1_temp), .IN2(n762), .QN(n521) );
  NAND2X0 U659 ( .IN1(n526), .IN2(n527), .QN(n174) );
  OR2X1 U660 ( .IN1(n460), .IN2(n258), .Q(n527) );
  NAND2X0 U661 ( .IN1(n528), .IN2(n460), .QN(n526) );
  NAND2X0 U662 ( .IN1(n529), .IN2(n530), .QN(n528) );
  NOR2X0 U663 ( .IN1(n531), .IN2(n532), .QN(n529) );
  AND2X1 U664 ( .IN1(xmit_dataH_7_), .IN2(n484), .Q(n532) );
  NOR2X0 U665 ( .IN1(n424), .IN2(n484), .QN(n531) );
  NAND2X0 U666 ( .IN1(n533), .IN2(n534), .QN(n173) );
  OR2X1 U667 ( .IN1(n460), .IN2(n259), .Q(n534) );
  NAND2X0 U668 ( .IN1(n535), .IN2(n460), .QN(n533) );
  NAND2X0 U669 ( .IN1(n536), .IN2(n537), .QN(n535) );
  NAND2X0 U670 ( .IN1(xmit_dataH_6_), .IN2(n538), .QN(n537) );
  NOR2X0 U671 ( .IN1(n539), .IN2(n540), .QN(n536) );
  NOR2X0 U672 ( .IN1(n258), .IN2(n484), .QN(n540) );
  NOR2X0 U673 ( .IN1(n424), .IN2(n530), .QN(n539) );
  NAND2X0 U674 ( .IN1(n541), .IN2(n542), .QN(n172) );
  NAND2X0 U675 ( .IN1(n773), .IN2(test_se), .QN(n542) );
  NAND2X0 U676 ( .IN1(n543), .IN2(n460), .QN(n541) );
  NAND2X0 U677 ( .IN1(n544), .IN2(n545), .QN(n543) );
  NAND2X0 U678 ( .IN1(xmit_dataH_5_), .IN2(n538), .QN(n545) );
  NOR2X0 U679 ( .IN1(n546), .IN2(n547), .QN(n544) );
  NOR2X0 U680 ( .IN1(n259), .IN2(n484), .QN(n547) );
  NOR2X0 U681 ( .IN1(n258), .IN2(n530), .QN(n546) );
  NAND2X0 U682 ( .IN1(n548), .IN2(n549), .QN(n171) );
  NAND2X0 U683 ( .IN1(n774), .IN2(test_se), .QN(n549) );
  NAND2X0 U684 ( .IN1(n550), .IN2(n460), .QN(n548) );
  NAND2X0 U685 ( .IN1(n551), .IN2(n552), .QN(n550) );
  NAND2X0 U686 ( .IN1(xmit_dataH_4_), .IN2(n538), .QN(n552) );
  NOR2X0 U687 ( .IN1(n553), .IN2(n554), .QN(n551) );
  NOR2X0 U688 ( .IN1(n484), .IN2(n445), .QN(n554) );
  NOR2X0 U689 ( .IN1(n259), .IN2(n530), .QN(n553) );
  NAND2X0 U690 ( .IN1(n555), .IN2(n556), .QN(n170) );
  NAND2X0 U691 ( .IN1(n775), .IN2(test_se), .QN(n556) );
  NAND2X0 U692 ( .IN1(n557), .IN2(n460), .QN(n555) );
  NAND2X0 U693 ( .IN1(n558), .IN2(n559), .QN(n557) );
  NAND2X0 U694 ( .IN1(xmit_dataH_3_), .IN2(n538), .QN(n559) );
  NOR2X0 U695 ( .IN1(n560), .IN2(n561), .QN(n558) );
  NOR2X0 U696 ( .IN1(n484), .IN2(n446), .QN(n561) );
  NOR2X0 U697 ( .IN1(n530), .IN2(n445), .QN(n560) );
  NAND2X0 U698 ( .IN1(n562), .IN2(n563), .QN(n169) );
  NAND2X0 U699 ( .IN1(n776), .IN2(test_se), .QN(n563) );
  NAND2X0 U700 ( .IN1(n564), .IN2(n460), .QN(n562) );
  NAND2X0 U701 ( .IN1(n565), .IN2(n566), .QN(n564) );
  NAND2X0 U702 ( .IN1(xmit_dataH_2_), .IN2(n538), .QN(n566) );
  NOR2X0 U703 ( .IN1(n567), .IN2(n568), .QN(n565) );
  NOR2X0 U704 ( .IN1(n484), .IN2(n447), .QN(n568) );
  NOR2X0 U705 ( .IN1(n530), .IN2(n446), .QN(n567) );
  NAND2X0 U706 ( .IN1(n569), .IN2(n570), .QN(n168) );
  OR2X1 U707 ( .IN1(n460), .IN2(n768), .Q(n570) );
  NAND2X0 U708 ( .IN1(n571), .IN2(n460), .QN(n569) );
  NAND2X0 U709 ( .IN1(n572), .IN2(n573), .QN(n571) );
  NAND2X0 U710 ( .IN1(xmit_dataH_1_), .IN2(n538), .QN(n573) );
  NOR2X0 U711 ( .IN1(n574), .IN2(n575), .QN(n572) );
  NOR2X0 U712 ( .IN1(n484), .IN2(n448), .QN(n575) );
  NOR2X0 U713 ( .IN1(n530), .IN2(n447), .QN(n574) );
  NAND2X0 U714 ( .IN1(n576), .IN2(n577), .QN(n167) );
  OR2X1 U715 ( .IN1(n460), .IN2(n424), .Q(n577) );
  NAND2X0 U716 ( .IN1(n578), .IN2(n460), .QN(n576) );
  NAND2X0 U717 ( .IN1(n520), .IN2(n579), .QN(n578) );
  NAND2X0 U718 ( .IN1(n452), .IN2(n476), .QN(n579) );
  INVX0 U719 ( .INP(n466), .ZN(n476) );
  NAND2X0 U720 ( .IN1(n580), .IN2(n780), .QN(n466) );
  INVX0 U721 ( .INP(n581), .ZN(n452) );
  NAND2X0 U722 ( .IN1(n582), .IN2(n246), .QN(n520) );
  NOR2X0 U723 ( .IN1(xmitH), .IN2(n777), .QN(n582) );
  NAND2X0 U724 ( .IN1(n583), .IN2(n584), .QN(n166) );
  NOR2X0 U725 ( .IN1(n585), .IN2(n586), .QN(n583) );
  NOR2X0 U726 ( .IN1(iRECEIVER_state_0_), .IN2(n587), .QN(n586) );
  NAND2X0 U727 ( .IN1(n588), .IN2(n460), .QN(n587) );
  NAND2X0 U728 ( .IN1(n770), .IN2(n589), .QN(n588) );
  NAND2X0 U729 ( .IN1(n590), .IN2(iRECEIVER_state_1_), .QN(n589) );
  NOR2X0 U730 ( .IN1(n245), .IN2(n591), .QN(n585) );
  NOR2X0 U731 ( .IN1(test_se), .IN2(n592), .QN(n591) );
  NAND2X0 U732 ( .IN1(n593), .IN2(n594), .QN(n592) );
  NAND2X0 U733 ( .IN1(n595), .IN2(iRECEIVER_state_1_), .QN(n594) );
  NAND2X0 U734 ( .IN1(n596), .IN2(n241), .QN(n593) );
  NOR2X0 U735 ( .IN1(n770), .IN2(iRECEIVER_state_2_), .QN(n596) );
  NAND2X0 U736 ( .IN1(n597), .IN2(n598), .QN(n164) );
  NAND2X0 U737 ( .IN1(n766), .IN2(test_se), .QN(n598) );
  NAND2X0 U738 ( .IN1(n599), .IN2(n460), .QN(n597) );
  NAND2X0 U739 ( .IN1(n600), .IN2(n238), .QN(n599) );
  NOR2X0 U740 ( .IN1(n601), .IN2(n602), .QN(n600) );
  NOR2X0 U741 ( .IN1(n241), .IN2(n603), .QN(n602) );
  NOR2X0 U742 ( .IN1(n604), .IN2(n605), .QN(n603) );
  INVX0 U743 ( .INP(n590), .ZN(n605) );
  NOR2X0 U744 ( .IN1(n245), .IN2(n606), .QN(n604) );
  NOR2X0 U745 ( .IN1(n607), .IN2(n595), .QN(n606) );
  NOR2X0 U746 ( .IN1(n608), .IN2(n609), .QN(n607) );
  NAND2X0 U747 ( .IN1(n766), .IN2(n432), .QN(n609) );
  NAND2X0 U748 ( .IN1(n429), .IN2(n437), .QN(n608) );
  NOR2X0 U749 ( .IN1(n431), .IN2(iRECEIVER_state_1_), .QN(n601) );
  NAND2X0 U750 ( .IN1(n610), .IN2(n611), .QN(n163) );
  NAND2X0 U751 ( .IN1(iRECEIVER_N20), .IN2(n460), .QN(n611) );
  NAND2X0 U752 ( .IN1(test_si), .IN2(test_se), .QN(n610) );
  NAND2X0 U753 ( .IN1(n612), .IN2(n613), .QN(n162) );
  NAND2X0 U754 ( .IN1(n614), .IN2(iRECEIVER_N20), .QN(n613) );
  NOR2X0 U755 ( .IN1(test_se), .IN2(n244), .QN(n614) );
  NAND2X0 U756 ( .IN1(n615), .IN2(iRECEIVER_bitCell_cntrH_0_), .QN(n612) );
  NAND2X0 U757 ( .IN1(n460), .IN2(n616), .QN(n615) );
  NAND2X0 U758 ( .IN1(n617), .IN2(n244), .QN(n616) );
  NAND2X0 U759 ( .IN1(n618), .IN2(n619), .QN(n161) );
  OR2X1 U760 ( .IN1(n460), .IN2(n244), .Q(n619) );
  NAND2X0 U761 ( .IN1(iRECEIVER_N22), .IN2(n460), .QN(n618) );
  NAND2X0 U762 ( .IN1(n620), .IN2(n621), .QN(n160) );
  NAND2X0 U763 ( .IN1(iRECEIVER_N23), .IN2(n460), .QN(n621) );
  NAND2X0 U764 ( .IN1(n784), .IN2(test_se), .QN(n620) );
  NAND2X0 U765 ( .IN1(n622), .IN2(n623), .QN(n159) );
  NAND2X0 U766 ( .IN1(test_se), .IN2(iRECEIVER_state_1_), .QN(n623) );
  INVX0 U767 ( .INP(n17), .ZN(n622) );
  NOR2X0 U768 ( .IN1(n624), .IN2(n595), .QN(n17) );
  NAND2X0 U769 ( .IN1(iRECEIVER_state_0_), .IN2(iRECEIVER_state_1_), .QN(n624)
         );
  NAND2X0 U770 ( .IN1(n625), .IN2(n626), .QN(n157) );
  NAND2X0 U771 ( .IN1(n769), .IN2(test_se), .QN(n626) );
  NAND2X0 U772 ( .IN1(n627), .IN2(n460), .QN(n625) );
  NAND2X0 U773 ( .IN1(n628), .IN2(n629), .QN(n627) );
  NAND2X0 U774 ( .IN1(iRECEIVER_state_2_), .IN2(iRECEIVER_state_0_), .QN(n629)
         );
  NAND2X0 U775 ( .IN1(n630), .IN2(n631), .QN(n156) );
  NAND2X0 U776 ( .IN1(rec_dataH_rec_6), .IN2(test_se), .QN(n631) );
  NOR2X0 U777 ( .IN1(n632), .IN2(n633), .QN(n630) );
  NOR2X0 U778 ( .IN1(n431), .IN2(n584), .QN(n633) );
  NOR2X0 U779 ( .IN1(n634), .IN2(n436), .QN(n632) );
  NAND2X0 U780 ( .IN1(n635), .IN2(n636), .QN(n155) );
  NAND2X0 U781 ( .IN1(rec_dataH_rec_7), .IN2(n460), .QN(n636) );
  NAND2X0 U782 ( .IN1(rec_dataH_temp_6_), .IN2(test_se), .QN(n635) );
  NAND2X0 U783 ( .IN1(n637), .IN2(n638), .QN(n154) );
  NAND2X0 U784 ( .IN1(test_so), .IN2(n460), .QN(n638) );
  NAND2X0 U785 ( .IN1(rec_dataH_6_), .IN2(test_se), .QN(n637) );
  NAND2X0 U786 ( .IN1(n639), .IN2(n640), .QN(n153) );
  NAND2X0 U787 ( .IN1(rec_dataH_rec_5), .IN2(test_se), .QN(n640) );
  NOR2X0 U788 ( .IN1(n641), .IN2(n642), .QN(n639) );
  NOR2X0 U789 ( .IN1(n436), .IN2(n584), .QN(n642) );
  NOR2X0 U790 ( .IN1(n634), .IN2(n438), .QN(n641) );
  NAND2X0 U791 ( .IN1(n643), .IN2(n644), .QN(n152) );
  NAND2X0 U792 ( .IN1(rec_dataH_rec_6), .IN2(n460), .QN(n644) );
  NAND2X0 U793 ( .IN1(rec_dataH_temp_5_), .IN2(test_se), .QN(n643) );
  NAND2X0 U794 ( .IN1(n645), .IN2(n646), .QN(n150) );
  NAND2X0 U795 ( .IN1(rec_dataH_temp_6_), .IN2(n460), .QN(n646) );
  NAND2X0 U796 ( .IN1(rec_dataH_5_), .IN2(test_se), .QN(n645) );
  NAND2X0 U797 ( .IN1(n647), .IN2(n648), .QN(n149) );
  NAND2X0 U798 ( .IN1(rec_dataH_rec_4), .IN2(test_se), .QN(n648) );
  NOR2X0 U799 ( .IN1(n649), .IN2(n650), .QN(n647) );
  NOR2X0 U800 ( .IN1(n584), .IN2(n438), .QN(n650) );
  NOR2X0 U801 ( .IN1(n634), .IN2(n439), .QN(n649) );
  NAND2X0 U802 ( .IN1(n651), .IN2(n652), .QN(n148) );
  NAND2X0 U803 ( .IN1(rec_dataH_rec_5), .IN2(n460), .QN(n652) );
  NAND2X0 U804 ( .IN1(rec_dataH_temp_4_), .IN2(test_se), .QN(n651) );
  NAND2X0 U805 ( .IN1(n653), .IN2(n654), .QN(n147) );
  NAND2X0 U806 ( .IN1(rec_dataH_temp_5_), .IN2(n460), .QN(n654) );
  NAND2X0 U807 ( .IN1(rec_dataH_4_), .IN2(test_se), .QN(n653) );
  NAND2X0 U808 ( .IN1(n655), .IN2(n656), .QN(n146) );
  NAND2X0 U809 ( .IN1(rec_dataH_rec_3), .IN2(test_se), .QN(n656) );
  NOR2X0 U810 ( .IN1(n657), .IN2(n658), .QN(n655) );
  NOR2X0 U811 ( .IN1(n584), .IN2(n439), .QN(n658) );
  NOR2X0 U812 ( .IN1(n634), .IN2(n440), .QN(n657) );
  NAND2X0 U813 ( .IN1(n659), .IN2(n660), .QN(n145) );
  NAND2X0 U814 ( .IN1(rec_dataH_rec_4), .IN2(n460), .QN(n660) );
  NAND2X0 U815 ( .IN1(rec_dataH_temp_3_), .IN2(test_se), .QN(n659) );
  NAND2X0 U816 ( .IN1(n661), .IN2(n662), .QN(n143) );
  NAND2X0 U817 ( .IN1(rec_dataH_temp_4_), .IN2(n460), .QN(n662) );
  NAND2X0 U818 ( .IN1(rec_dataH_3_), .IN2(test_se), .QN(n661) );
  NAND2X0 U819 ( .IN1(n663), .IN2(n664), .QN(n142) );
  NAND2X0 U820 ( .IN1(rec_dataH_rec_2), .IN2(test_se), .QN(n664) );
  NOR2X0 U821 ( .IN1(n665), .IN2(n666), .QN(n663) );
  NOR2X0 U822 ( .IN1(n584), .IN2(n440), .QN(n666) );
  NOR2X0 U823 ( .IN1(n634), .IN2(n441), .QN(n665) );
  NAND2X0 U824 ( .IN1(n667), .IN2(n668), .QN(n141) );
  NAND2X0 U825 ( .IN1(rec_dataH_rec_3), .IN2(n460), .QN(n668) );
  NAND2X0 U826 ( .IN1(rec_dataH_temp_2_), .IN2(test_se), .QN(n667) );
  NAND2X0 U827 ( .IN1(n669), .IN2(n670), .QN(n140) );
  NAND2X0 U828 ( .IN1(rec_dataH_temp_3_), .IN2(n460), .QN(n670) );
  NAND2X0 U829 ( .IN1(rec_dataH_2_), .IN2(test_se), .QN(n669) );
  NAND2X0 U830 ( .IN1(n671), .IN2(n672), .QN(n139) );
  NAND2X0 U831 ( .IN1(rec_dataH_rec_1), .IN2(test_se), .QN(n672) );
  NOR2X0 U832 ( .IN1(n673), .IN2(n674), .QN(n671) );
  NOR2X0 U833 ( .IN1(n584), .IN2(n441), .QN(n674) );
  NOR2X0 U834 ( .IN1(n634), .IN2(n442), .QN(n673) );
  NAND2X0 U835 ( .IN1(n675), .IN2(n676), .QN(n138) );
  NAND2X0 U836 ( .IN1(rec_dataH_rec_2), .IN2(n460), .QN(n676) );
  NAND2X0 U837 ( .IN1(rec_dataH_temp_1_), .IN2(test_se), .QN(n675) );
  NAND2X0 U838 ( .IN1(n677), .IN2(n678), .QN(n136) );
  NAND2X0 U839 ( .IN1(rec_dataH_temp_2_), .IN2(n460), .QN(n678) );
  NAND2X0 U840 ( .IN1(rec_dataH_1_), .IN2(test_se), .QN(n677) );
  NAND2X0 U841 ( .IN1(n679), .IN2(n680), .QN(n135) );
  NAND2X0 U842 ( .IN1(rec_dataH_rec_0), .IN2(test_se), .QN(n680) );
  NOR2X0 U843 ( .IN1(n681), .IN2(n682), .QN(n679) );
  NOR2X0 U844 ( .IN1(n584), .IN2(n442), .QN(n682) );
  NOR2X0 U845 ( .IN1(n634), .IN2(n443), .QN(n681) );
  NAND2X0 U846 ( .IN1(n683), .IN2(n684), .QN(n134) );
  NAND2X0 U847 ( .IN1(rec_dataH_rec_1), .IN2(n460), .QN(n684) );
  NAND2X0 U848 ( .IN1(rec_dataH_temp_0_), .IN2(test_se), .QN(n683) );
  NAND2X0 U849 ( .IN1(n685), .IN2(n686), .QN(n133) );
  NAND2X0 U850 ( .IN1(rec_dataH_temp_1_), .IN2(n460), .QN(n686) );
  NAND2X0 U851 ( .IN1(rec_dataH_0_), .IN2(test_se), .QN(n685) );
  NAND2X0 U852 ( .IN1(n687), .IN2(n688), .QN(n132) );
  NAND2X0 U853 ( .IN1(n765), .IN2(test_se), .QN(n688) );
  NOR2X0 U854 ( .IN1(n689), .IN2(n690), .QN(n687) );
  NOR2X0 U855 ( .IN1(n584), .IN2(n443), .QN(n690) );
  AND2X1 U856 ( .IN1(n691), .IN2(rec_dataH_rec_0), .Q(n689) );
  NAND2X0 U857 ( .IN1(n692), .IN2(n693), .QN(n131) );
  NAND2X0 U858 ( .IN1(rec_dataH_rec_0), .IN2(n460), .QN(n693) );
  NAND2X0 U859 ( .IN1(rec_dataH_7_), .IN2(test_se), .QN(n692) );
  NAND2X0 U860 ( .IN1(n694), .IN2(n695), .QN(n129) );
  NAND2X0 U861 ( .IN1(rec_dataH_temp_0_), .IN2(n460), .QN(n695) );
  NAND2X0 U862 ( .IN1(xmit_doneH), .IN2(test_se), .QN(n694) );
  NAND2X0 U863 ( .IN1(n696), .IN2(n697), .QN(n128) );
  NAND2X0 U864 ( .IN1(n782), .IN2(test_se), .QN(n697) );
  NOR2X0 U865 ( .IN1(n698), .IN2(n699), .QN(n696) );
  NOR2X0 U866 ( .IN1(n433), .IN2(n700), .QN(n699) );
  NOR2X0 U867 ( .IN1(n701), .IN2(n584), .QN(n698) );
  NAND2X0 U868 ( .IN1(n702), .IN2(n703), .QN(n127) );
  NAND2X0 U869 ( .IN1(test_se), .IN2(rec_readyH), .QN(n703) );
  NOR2X0 U870 ( .IN1(n704), .IN2(n705), .QN(n702) );
  NOR2X0 U871 ( .IN1(n437), .IN2(n700), .QN(n705) );
  NOR2X0 U872 ( .IN1(n767), .IN2(n584), .QN(n704) );
  NAND2X0 U873 ( .IN1(n706), .IN2(n707), .QN(n126) );
  NAND2X0 U874 ( .IN1(n767), .IN2(test_se), .QN(n707) );
  NOR2X0 U875 ( .IN1(n708), .IN2(n709), .QN(n706) );
  NOR2X0 U876 ( .IN1(n432), .IN2(n700), .QN(n709) );
  NOR2X0 U877 ( .IN1(n710), .IN2(n584), .QN(n708) );
  INVX0 U878 ( .INP(iRECEIVER_N26), .ZN(n710) );
  NAND2X0 U879 ( .IN1(n711), .IN2(n712), .QN(n125) );
  NAND2X0 U880 ( .IN1(n783), .IN2(test_se), .QN(n712) );
  NOR2X0 U881 ( .IN1(n713), .IN2(n714), .QN(n711) );
  NOR2X0 U882 ( .IN1(n429), .IN2(n700), .QN(n714) );
  NAND2X0 U883 ( .IN1(n691), .IN2(n628), .QN(n700) );
  NAND2X0 U884 ( .IN1(n715), .IN2(n241), .QN(n628) );
  NOR2X0 U885 ( .IN1(n431), .IN2(iRECEIVER_state_2_), .QN(n715) );
  INVX0 U886 ( .INP(n634), .ZN(n691) );
  NAND2X0 U887 ( .IN1(n460), .IN2(n716), .QN(n634) );
  NAND2X0 U888 ( .IN1(n245), .IN2(iRECEIVER_state_2_), .QN(n716) );
  NOR2X0 U889 ( .IN1(n717), .IN2(n584), .QN(n713) );
  NAND2X0 U890 ( .IN1(n718), .IN2(n245), .QN(n584) );
  NOR2X0 U891 ( .IN1(test_se), .IN2(n238), .QN(n718) );
  NAND2X0 U892 ( .IN1(n719), .IN2(n720), .QN(n124) );
  NAND2X0 U893 ( .IN1(n721), .IN2(n460), .QN(n720) );
  AND2X1 U894 ( .IN1(n722), .IN2(iXMIT_N25), .Q(n721) );
  NAND2X0 U895 ( .IN1(n781), .IN2(test_se), .QN(n719) );
  NAND2X0 U896 ( .IN1(n723), .IN2(n724), .QN(n122) );
  NAND2X0 U897 ( .IN1(test_se), .IN2(iRECEIVER_state_2_), .QN(n724) );
  NAND2X0 U898 ( .IN1(iXMIT_N26), .IN2(n460), .QN(n723) );
  NAND2X0 U899 ( .IN1(n725), .IN2(n726), .QN(n121) );
  NOR2X0 U900 ( .IN1(n727), .IN2(n728), .QN(n725) );
  NOR2X0 U901 ( .IN1(n460), .IN2(n430), .QN(n728) );
  NOR2X0 U902 ( .IN1(test_se), .IN2(n729), .QN(n727) );
  NAND2X0 U903 ( .IN1(n730), .IN2(n731), .QN(n120) );
  NAND2X0 U904 ( .IN1(test_se), .IN2(n777), .QN(n731) );
  NAND2X0 U905 ( .IN1(n732), .IN2(n460), .QN(n730) );
  NAND2X0 U906 ( .IN1(n733), .IN2(n734), .QN(n732) );
  NAND2X0 U907 ( .IN1(xmit_dataH_0_), .IN2(n538), .QN(n734) );
  INVX0 U908 ( .INP(n735), .ZN(n538) );
  NOR2X0 U909 ( .IN1(n736), .IN2(n737), .QN(n733) );
  NOR2X0 U910 ( .IN1(n768), .IN2(n484), .QN(n737) );
  NOR2X0 U911 ( .IN1(n530), .IN2(n448), .QN(n736) );
  NAND2X0 U912 ( .IN1(n484), .IN2(n735), .QN(n530) );
  NAND2X0 U913 ( .IN1(n735), .IN2(n738), .QN(n484) );
  NAND2X0 U914 ( .IN1(n777), .IN2(n239), .QN(n738) );
  NAND2X0 U915 ( .IN1(n739), .IN2(xmitH), .QN(n735) );
  NOR2X0 U916 ( .IN1(n777), .IN2(iXMIT_state_1_temp), .QN(n739) );
  NAND2X0 U917 ( .IN1(n740), .IN2(n741), .QN(n119) );
  NAND2X0 U918 ( .IN1(uart_REC_dataH), .IN2(n460), .QN(n741) );
  NAND2X0 U919 ( .IN1(n770), .IN2(test_se), .QN(n740) );
  NAND2X0 U920 ( .IN1(n742), .IN2(n743), .QN(n118) );
  NAND2X0 U921 ( .IN1(n769), .IN2(n460), .QN(n743) );
  INVX0 U922 ( .INP(test_se), .ZN(n460) );
  NAND2X0 U923 ( .IN1(rec_dataH_rec_7), .IN2(test_se), .QN(n742) );
  AND2X1 U924 ( .IN1(iXMIT_N24), .IN2(n722), .Q(iXMIT_N28) );
  NAND2X0 U925 ( .IN1(n726), .IN2(n729), .QN(iXMIT_N27) );
  NAND2X0 U926 ( .IN1(iXMIT_N26), .IN2(n778), .QN(n729) );
  NAND2X0 U927 ( .IN1(n744), .IN2(n779), .QN(n726) );
  NOR2X0 U928 ( .IN1(n778), .IN2(n745), .QN(n744) );
  NOR2X0 U929 ( .IN1(n745), .IN2(n779), .QN(iXMIT_N26) );
  INVX0 U930 ( .INP(n722), .ZN(n745) );
  NAND2X0 U931 ( .IN1(n581), .IN2(n483), .QN(n722) );
  NAND2X0 U932 ( .IN1(n478), .IN2(iXMIT_state_1_temp), .QN(n483) );
  NAND2X0 U933 ( .IN1(n522), .IN2(n762), .QN(n478) );
  AND2X1 U934 ( .IN1(n746), .IN2(n747), .Q(n522) );
  NOR2X0 U935 ( .IN1(n779), .IN2(n435), .QN(n747) );
  AND2X1 U936 ( .IN1(n781), .IN2(n780), .Q(n746) );
  NAND2X0 U937 ( .IN1(n762), .IN2(n777), .QN(n581) );
  XOR2X1 U938 ( .IN1(n780), .IN2(n580), .Q(iXMIT_N25) );
  AND2X1 U939 ( .IN1(n748), .IN2(n781), .Q(n580) );
  XOR2X1 U940 ( .IN1(n748), .IN2(n781), .Q(iXMIT_N24) );
  NOR2X0 U941 ( .IN1(n430), .IN2(n435), .QN(n748) );
  INVX0 U942 ( .INP(n701), .ZN(iRECEIVER_N28) );
  XOR2X1 U943 ( .IN1(n433), .IN2(n749), .Q(n701) );
  NOR2X0 U944 ( .IN1(n750), .IN2(n429), .QN(n749) );
  INVX0 U945 ( .INP(n717), .ZN(iRECEIVER_N27) );
  XOR2X1 U946 ( .IN1(n750), .IN2(n782), .Q(n717) );
  NAND2X0 U947 ( .IN1(n767), .IN2(n783), .QN(n750) );
  XNOR2X1 U948 ( .IN1(n432), .IN2(n767), .Q(iRECEIVER_N26) );
  AND2X1 U949 ( .IN1(n617), .IN2(iRECEIVER_N19), .Q(iRECEIVER_N23) );
  AND2X1 U950 ( .IN1(n617), .IN2(iRECEIVER_N18), .Q(iRECEIVER_N22) );
  AND2X1 U951 ( .IN1(iRECEIVER_N17), .IN2(n617), .Q(iRECEIVER_N21) );
  INVX0 U952 ( .INP(n751), .ZN(n617) );
  NOR2X0 U953 ( .IN1(n751), .IN2(iRECEIVER_bitCell_cntrH_0_), .QN(
        iRECEIVER_N20) );
  NAND2X0 U954 ( .IN1(n752), .IN2(n753), .QN(n751) );
  NOR2X0 U955 ( .IN1(n754), .IN2(n755), .QN(n753) );
  NOR2X0 U956 ( .IN1(iRECEIVER_state_0_), .IN2(n590), .QN(n755) );
  NAND2X0 U957 ( .IN1(n756), .IN2(n757), .QN(n590) );
  NOR2X0 U958 ( .IN1(n765), .IN2(iRECEIVER_bitCell_cntrH_0_), .QN(n757) );
  AND2X1 U959 ( .IN1(n784), .IN2(n244), .Q(n756) );
  NOR2X0 U960 ( .IN1(n245), .IN2(n595), .QN(n754) );
  NAND2X0 U961 ( .IN1(n758), .IN2(n759), .QN(n595) );
  NOR2X0 U962 ( .IN1(n244), .IN2(iRECEIVER_bitCell_cntrH_0_), .QN(n759) );
  AND2X1 U963 ( .IN1(n784), .IN2(n765), .Q(n758) );
  NOR2X0 U964 ( .IN1(n241), .IN2(iRECEIVER_state_2_), .QN(n752) );
  XNOR2X1 U965 ( .IN1(n760), .IN2(n765), .Q(iRECEIVER_N19) );
  NAND2X0 U966 ( .IN1(n761), .IN2(n784), .QN(n760) );
  XOR2X1 U967 ( .IN1(n784), .IN2(n761), .Q(iRECEIVER_N18) );
  NOR2X0 U968 ( .IN1(n255), .IN2(n244), .QN(n761) );
  XOR2X1 U969 ( .IN1(n244), .IN2(n255), .Q(iRECEIVER_N17) );
endmodule

