module locked_c1908 (  G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,  G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n123_, new_n124_, new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_, new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_, new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n389_, new_n390_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n418_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n430_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n481_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_;
  INV_X1 g000 ( .A(KEYINPUT22), .ZN(new_n123_) );
  INV_X1 g001 ( .A(G902), .ZN(new_n124_) );
  INV_X1 g002 ( .A(KEYINPUT8), .ZN(new_n125_) );
  INV_X1 g003 ( .A(G953), .ZN(new_n126_) );
  NAND2_X1 g004 ( .A1(new_n126_), .A2(G234), .ZN(new_n127_) );
  NAND2_X1 g005 ( .A1(new_n127_), .A2(new_n125_), .ZN(new_n128_) );
  NAND3_X1 g006 ( .A1(new_n126_), .A2(G234), .A3(KEYINPUT8), .ZN(new_n129_) );
  NAND2_X1 g007 ( .A1(new_n128_), .A2(new_n129_), .ZN(new_n130_) );
  NAND2_X1 g008 ( .A1(new_n130_), .A2(G217), .ZN(new_n131_) );
  XOR2_X1 g009 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(new_n132_) );
  INV_X1 g010 ( .A(new_n132_), .ZN(new_n133_) );
  NAND2_X1 g011 ( .A1(new_n131_), .A2(new_n133_), .ZN(new_n134_) );
  NAND3_X1 g012 ( .A1(new_n130_), .A2(G217), .A3(new_n132_), .ZN(new_n135_) );
  NAND2_X1 g013 ( .A1(new_n134_), .A2(new_n135_), .ZN(new_n136_) );
  NAND2_X1 g014 ( .A1(new_n136_), .A2(G116), .ZN(new_n137_) );
  INV_X1 g015 ( .A(G116), .ZN(new_n138_) );
  NAND3_X1 g016 ( .A1(new_n134_), .A2(new_n138_), .A3(new_n135_), .ZN(new_n139_) );
  NAND2_X1 g017 ( .A1(new_n137_), .A2(new_n139_), .ZN(new_n140_) );
  INV_X1 g018 ( .A(G107), .ZN(new_n141_) );
  NAND2_X1 g019 ( .A1(G128), .A2(G143), .ZN(new_n142_) );
  INV_X1 g020 ( .A(G128), .ZN(new_n143_) );
  INV_X1 g021 ( .A(G143), .ZN(new_n144_) );
  NAND2_X1 g022 ( .A1(new_n143_), .A2(new_n144_), .ZN(new_n145_) );
  NAND2_X1 g023 ( .A1(new_n145_), .A2(new_n142_), .ZN(new_n146_) );
  XNOR2_X1 g024 ( .A(new_n146_), .B(new_n141_), .ZN(new_n147_) );
  INV_X1 g025 ( .A(new_n147_), .ZN(new_n148_) );
  NAND2_X1 g026 ( .A1(new_n140_), .A2(new_n148_), .ZN(new_n149_) );
  NAND3_X1 g027 ( .A1(new_n137_), .A2(new_n139_), .A3(new_n147_), .ZN(new_n150_) );
  NAND2_X1 g028 ( .A1(new_n149_), .A2(new_n150_), .ZN(new_n151_) );
  XOR2_X1 g029 ( .A(G122), .B(G134), .Z(new_n152_) );
  INV_X1 g030 ( .A(new_n152_), .ZN(new_n153_) );
  NAND2_X1 g031 ( .A1(new_n151_), .A2(new_n153_), .ZN(new_n154_) );
  NAND3_X1 g032 ( .A1(new_n149_), .A2(new_n150_), .A3(new_n152_), .ZN(new_n155_) );
  NAND4_X1 g033 ( .A1(new_n154_), .A2(G478), .A3(new_n124_), .A4(new_n155_), .ZN(new_n156_) );
  INV_X1 g034 ( .A(G478), .ZN(new_n157_) );
  NAND3_X1 g035 ( .A1(new_n154_), .A2(new_n124_), .A3(new_n155_), .ZN(new_n158_) );
  NAND2_X1 g036 ( .A1(new_n158_), .A2(new_n157_), .ZN(new_n159_) );
  NAND2_X1 g037 ( .A1(new_n159_), .A2(new_n156_), .ZN(new_n160_) );
  XNOR2_X1 g038 ( .A(G113), .B(G122), .ZN(new_n161_) );
  INV_X1 g039 ( .A(new_n161_), .ZN(new_n162_) );
  XNOR2_X1 g040 ( .A(G140), .B(KEYINPUT11), .ZN(new_n163_) );
  NAND2_X1 g041 ( .A1(new_n162_), .A2(new_n163_), .ZN(new_n164_) );
  INV_X1 g042 ( .A(new_n163_), .ZN(new_n165_) );
  NAND2_X1 g043 ( .A1(new_n165_), .A2(new_n161_), .ZN(new_n166_) );
  NAND2_X1 g044 ( .A1(new_n164_), .A2(new_n166_), .ZN(new_n167_) );
  XOR2_X1 g045 ( .A(G125), .B(KEYINPUT10), .Z(new_n168_) );
  NAND2_X1 g046 ( .A1(new_n167_), .A2(new_n168_), .ZN(new_n169_) );
  XNOR2_X1 g047 ( .A(G125), .B(KEYINPUT10), .ZN(new_n170_) );
  NAND3_X1 g048 ( .A1(new_n164_), .A2(new_n166_), .A3(new_n170_), .ZN(new_n171_) );
  NAND2_X1 g049 ( .A1(new_n169_), .A2(new_n171_), .ZN(new_n172_) );
  XNOR2_X1 g050 ( .A(G104), .B(G143), .ZN(new_n173_) );
  INV_X1 g051 ( .A(new_n173_), .ZN(new_n174_) );
  NAND2_X1 g052 ( .A1(new_n172_), .A2(new_n174_), .ZN(new_n175_) );
  NAND3_X1 g053 ( .A1(new_n169_), .A2(new_n171_), .A3(new_n173_), .ZN(new_n176_) );
  NAND2_X1 g054 ( .A1(new_n175_), .A2(new_n176_), .ZN(new_n177_) );
  NAND2_X1 g055 ( .A1(G131), .A2(G146), .ZN(new_n178_) );
  INV_X1 g056 ( .A(G131), .ZN(new_n179_) );
  INV_X1 g057 ( .A(G146), .ZN(new_n180_) );
  NAND2_X1 g058 ( .A1(new_n179_), .A2(new_n180_), .ZN(new_n181_) );
  NAND2_X1 g059 ( .A1(new_n181_), .A2(new_n178_), .ZN(new_n182_) );
  XNOR2_X1 g060 ( .A(new_n182_), .B(KEYINPUT12), .ZN(new_n183_) );
  NOR2_X1 g061 ( .A1(G237), .A2(G953), .ZN(new_n184_) );
  NAND2_X1 g062 ( .A1(new_n184_), .A2(G214), .ZN(new_n185_) );
  XNOR2_X1 g063 ( .A(new_n183_), .B(new_n185_), .ZN(new_n186_) );
  INV_X1 g064 ( .A(new_n186_), .ZN(new_n187_) );
  NAND2_X1 g065 ( .A1(new_n177_), .A2(new_n187_), .ZN(new_n188_) );
  NAND3_X1 g066 ( .A1(new_n175_), .A2(new_n176_), .A3(new_n186_), .ZN(new_n189_) );
  NAND2_X1 g067 ( .A1(new_n188_), .A2(new_n189_), .ZN(new_n190_) );
  NAND2_X1 g068 ( .A1(new_n190_), .A2(new_n124_), .ZN(new_n191_) );
  XOR2_X1 g069 ( .A(G475), .B(KEYINPUT13), .Z(new_n192_) );
  INV_X1 g070 ( .A(new_n192_), .ZN(new_n193_) );
  NAND2_X1 g071 ( .A1(new_n191_), .A2(new_n193_), .ZN(new_n194_) );
  NAND3_X1 g072 ( .A1(new_n190_), .A2(new_n124_), .A3(new_n192_), .ZN(new_n195_) );
  NAND2_X1 g073 ( .A1(new_n194_), .A2(new_n195_), .ZN(new_n196_) );
  NAND2_X1 g074 ( .A1(new_n160_), .A2(new_n196_), .ZN(new_n197_) );
  INV_X1 g075 ( .A(new_n197_), .ZN(new_n198_) );
  XNOR2_X1 g076 ( .A(G902), .B(KEYINPUT15), .ZN(new_n199_) );
  NAND2_X1 g077 ( .A1(new_n199_), .A2(G234), .ZN(new_n200_) );
  XNOR2_X1 g078 ( .A(new_n200_), .B(KEYINPUT20), .ZN(new_n201_) );
  NAND2_X1 g079 ( .A1(new_n201_), .A2(G221), .ZN(new_n202_) );
  XOR2_X1 g080 ( .A(new_n202_), .B(KEYINPUT21), .Z(new_n203_) );
  NAND2_X1 g081 ( .A1(new_n198_), .A2(new_n203_), .ZN(new_n204_) );
  INV_X1 g082 ( .A(new_n204_), .ZN(new_n205_) );
  INV_X1 g083 ( .A(KEYINPUT0), .ZN(new_n206_) );
  INV_X1 g084 ( .A(G101), .ZN(new_n207_) );
  NAND2_X1 g085 ( .A1(new_n146_), .A2(KEYINPUT4), .ZN(new_n208_) );
  INV_X1 g086 ( .A(KEYINPUT4), .ZN(new_n209_) );
  NAND3_X1 g087 ( .A1(new_n145_), .A2(new_n209_), .A3(new_n142_), .ZN(new_n210_) );
  NAND2_X1 g088 ( .A1(new_n208_), .A2(new_n210_), .ZN(new_n211_) );
  NAND2_X1 g089 ( .A1(new_n211_), .A2(new_n207_), .ZN(new_n212_) );
  NAND3_X1 g090 ( .A1(new_n208_), .A2(G101), .A3(new_n210_), .ZN(new_n213_) );
  NAND2_X1 g091 ( .A1(new_n212_), .A2(new_n213_), .ZN(new_n214_) );
  XNOR2_X1 g092 ( .A(G104), .B(G110), .ZN(new_n215_) );
  XNOR2_X1 g093 ( .A(new_n215_), .B(G107), .ZN(new_n216_) );
  INV_X1 g094 ( .A(new_n216_), .ZN(new_n217_) );
  NAND2_X1 g095 ( .A1(new_n214_), .A2(new_n217_), .ZN(new_n218_) );
  NAND3_X1 g096 ( .A1(new_n212_), .A2(new_n213_), .A3(new_n216_), .ZN(new_n219_) );
  XOR2_X1 g097 ( .A(G125), .B(G146), .Z(new_n220_) );
  INV_X1 g098 ( .A(new_n220_), .ZN(new_n221_) );
  NAND2_X1 g099 ( .A1(new_n126_), .A2(G224), .ZN(new_n222_) );
  INV_X1 g100 ( .A(new_n222_), .ZN(new_n223_) );
  INV_X1 g101 ( .A(KEYINPUT18), .ZN(new_n224_) );
  NAND2_X1 g102 ( .A1(new_n224_), .A2(KEYINPUT17), .ZN(new_n225_) );
  INV_X1 g103 ( .A(KEYINPUT17), .ZN(new_n226_) );
  NAND2_X1 g104 ( .A1(new_n226_), .A2(KEYINPUT18), .ZN(new_n227_) );
  NAND2_X1 g105 ( .A1(new_n225_), .A2(new_n227_), .ZN(new_n228_) );
  NAND2_X1 g106 ( .A1(new_n228_), .A2(new_n223_), .ZN(new_n229_) );
  NAND3_X1 g107 ( .A1(new_n222_), .A2(new_n225_), .A3(new_n227_), .ZN(new_n230_) );
  NAND3_X1 g108 ( .A1(new_n221_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_) );
  NAND2_X1 g109 ( .A1(new_n229_), .A2(new_n230_), .ZN(new_n232_) );
  NAND2_X1 g110 ( .A1(new_n232_), .A2(new_n220_), .ZN(new_n233_) );
  NAND2_X1 g111 ( .A1(G119), .A2(KEYINPUT3), .ZN(new_n234_) );
  INV_X1 g112 ( .A(G119), .ZN(new_n235_) );
  INV_X1 g113 ( .A(KEYINPUT3), .ZN(new_n236_) );
  NAND2_X1 g114 ( .A1(new_n235_), .A2(new_n236_), .ZN(new_n237_) );
  NAND2_X1 g115 ( .A1(new_n237_), .A2(new_n234_), .ZN(new_n238_) );
  NAND2_X1 g116 ( .A1(new_n138_), .A2(G113), .ZN(new_n239_) );
  INV_X1 g117 ( .A(G113), .ZN(new_n240_) );
  NAND2_X1 g118 ( .A1(new_n240_), .A2(G116), .ZN(new_n241_) );
  NAND2_X1 g119 ( .A1(new_n239_), .A2(new_n241_), .ZN(new_n242_) );
  NAND2_X1 g120 ( .A1(new_n242_), .A2(new_n238_), .ZN(new_n243_) );
  NAND4_X1 g121 ( .A1(new_n237_), .A2(new_n239_), .A3(new_n241_), .A4(new_n234_), .ZN(new_n244_) );
  NAND2_X1 g122 ( .A1(new_n243_), .A2(new_n244_), .ZN(new_n245_) );
  XNOR2_X1 g123 ( .A(G122), .B(KEYINPUT16), .ZN(new_n246_) );
  NAND2_X1 g124 ( .A1(new_n245_), .A2(new_n246_), .ZN(new_n247_) );
  INV_X1 g125 ( .A(new_n246_), .ZN(new_n248_) );
  NAND3_X1 g126 ( .A1(new_n243_), .A2(new_n244_), .A3(new_n248_), .ZN(new_n249_) );
  NAND2_X1 g127 ( .A1(new_n247_), .A2(new_n249_), .ZN(new_n250_) );
  NAND3_X1 g128 ( .A1(new_n250_), .A2(new_n231_), .A3(new_n233_), .ZN(new_n251_) );
  NAND3_X1 g129 ( .A1(new_n243_), .A2(new_n244_), .A3(new_n248_), .ZN(new_n252_) );
  NAND3_X1 g130 ( .A1(new_n222_), .A2(new_n225_), .A3(new_n227_), .ZN(new_n253_) );
  NAND3_X1 g131 ( .A1(new_n221_), .A2(new_n229_), .A3(new_n253_), .ZN(new_n254_) );
  NAND2_X1 g132 ( .A1(new_n233_), .A2(new_n254_), .ZN(new_n255_) );
  NAND3_X1 g133 ( .A1(new_n255_), .A2(new_n247_), .A3(new_n252_), .ZN(new_n256_) );
  NAND4_X1 g134 ( .A1(new_n251_), .A2(new_n256_), .A3(new_n218_), .A4(new_n219_), .ZN(new_n257_) );
  NAND2_X1 g135 ( .A1(new_n218_), .A2(new_n219_), .ZN(new_n258_) );
  NAND2_X1 g136 ( .A1(new_n233_), .A2(new_n231_), .ZN(new_n259_) );
  NAND3_X1 g137 ( .A1(new_n259_), .A2(new_n247_), .A3(new_n249_), .ZN(new_n260_) );
  NAND2_X1 g138 ( .A1(new_n247_), .A2(new_n252_), .ZN(new_n261_) );
  NAND3_X1 g139 ( .A1(new_n261_), .A2(new_n233_), .A3(new_n254_), .ZN(new_n262_) );
  NAND2_X1 g140 ( .A1(new_n262_), .A2(new_n260_), .ZN(new_n263_) );
  NAND2_X1 g141 ( .A1(new_n263_), .A2(new_n258_), .ZN(new_n264_) );
  NAND2_X1 g142 ( .A1(new_n264_), .A2(new_n257_), .ZN(new_n265_) );
  NAND2_X1 g143 ( .A1(new_n265_), .A2(new_n199_), .ZN(new_n266_) );
  NOR2_X1 g144 ( .A1(G237), .A2(G902), .ZN(new_n267_) );
  INV_X1 g145 ( .A(new_n267_), .ZN(new_n268_) );
  NAND2_X1 g146 ( .A1(new_n268_), .A2(G210), .ZN(new_n269_) );
  INV_X1 g147 ( .A(new_n269_), .ZN(new_n270_) );
  NAND2_X1 g148 ( .A1(new_n266_), .A2(new_n270_), .ZN(new_n271_) );
  NAND3_X1 g149 ( .A1(new_n265_), .A2(new_n199_), .A3(new_n269_), .ZN(new_n272_) );
  NAND2_X1 g150 ( .A1(new_n271_), .A2(new_n272_), .ZN(new_n273_) );
  NAND2_X1 g151 ( .A1(new_n268_), .A2(G214), .ZN(new_n274_) );
  NAND2_X1 g152 ( .A1(new_n273_), .A2(new_n274_), .ZN(new_n275_) );
  NAND2_X1 g153 ( .A1(new_n275_), .A2(KEYINPUT19), .ZN(new_n276_) );
  INV_X1 g154 ( .A(KEYINPUT19), .ZN(new_n277_) );
  NAND3_X1 g155 ( .A1(new_n273_), .A2(new_n277_), .A3(new_n274_), .ZN(new_n278_) );
  NAND2_X1 g156 ( .A1(new_n276_), .A2(new_n278_), .ZN(new_n279_) );
  INV_X1 g157 ( .A(G898), .ZN(new_n280_) );
  NAND2_X1 g158 ( .A1(G234), .A2(G237), .ZN(new_n281_) );
  XNOR2_X1 g159 ( .A(new_n281_), .B(KEYINPUT14), .ZN(new_n282_) );
  NAND2_X1 g160 ( .A1(new_n282_), .A2(G902), .ZN(new_n283_) );
  INV_X1 g161 ( .A(new_n283_), .ZN(new_n284_) );
  NAND3_X1 g162 ( .A1(new_n284_), .A2(new_n280_), .A3(G953), .ZN(new_n285_) );
  NAND2_X1 g163 ( .A1(new_n282_), .A2(G952), .ZN(new_n286_) );
  INV_X1 g164 ( .A(new_n286_), .ZN(new_n287_) );
  NAND2_X1 g165 ( .A1(new_n287_), .A2(new_n126_), .ZN(new_n288_) );
  NAND2_X1 g166 ( .A1(new_n285_), .A2(new_n288_), .ZN(new_n289_) );
  NAND3_X1 g167 ( .A1(new_n279_), .A2(new_n206_), .A3(new_n289_), .ZN(new_n290_) );
  NAND2_X1 g168 ( .A1(new_n279_), .A2(new_n289_), .ZN(new_n291_) );
  NAND2_X1 g169 ( .A1(new_n291_), .A2(KEYINPUT0), .ZN(new_n292_) );
  NAND3_X1 g170 ( .A1(new_n292_), .A2(new_n205_), .A3(new_n290_), .ZN(new_n293_) );
  NAND2_X1 g171 ( .A1(new_n293_), .A2(new_n123_), .ZN(new_n294_) );
  NAND4_X1 g172 ( .A1(new_n292_), .A2(KEYINPUT22), .A3(new_n205_), .A4(new_n290_), .ZN(new_n295_) );
  NAND2_X1 g173 ( .A1(new_n294_), .A2(new_n295_), .ZN(new_n296_) );
  INV_X1 g174 ( .A(KEYINPUT1), .ZN(new_n297_) );
  XNOR2_X1 g175 ( .A(G137), .B(G140), .ZN(new_n298_) );
  INV_X1 g176 ( .A(new_n298_), .ZN(new_n299_) );
  NAND2_X1 g177 ( .A1(new_n182_), .A2(G134), .ZN(new_n300_) );
  INV_X1 g178 ( .A(G134), .ZN(new_n301_) );
  NAND3_X1 g179 ( .A1(new_n181_), .A2(new_n301_), .A3(new_n178_), .ZN(new_n302_) );
  NAND3_X1 g180 ( .A1(new_n300_), .A2(new_n299_), .A3(new_n302_), .ZN(new_n303_) );
  NAND2_X1 g181 ( .A1(new_n300_), .A2(new_n302_), .ZN(new_n304_) );
  NAND2_X1 g182 ( .A1(new_n304_), .A2(new_n298_), .ZN(new_n305_) );
  NAND2_X1 g183 ( .A1(new_n305_), .A2(new_n303_), .ZN(new_n306_) );
  NAND3_X1 g184 ( .A1(new_n306_), .A2(G227), .A3(new_n126_), .ZN(new_n307_) );
  NAND2_X1 g185 ( .A1(new_n126_), .A2(G227), .ZN(new_n308_) );
  NAND3_X1 g186 ( .A1(new_n305_), .A2(new_n303_), .A3(new_n308_), .ZN(new_n309_) );
  NAND4_X1 g187 ( .A1(new_n307_), .A2(new_n218_), .A3(new_n219_), .A4(new_n309_), .ZN(new_n310_) );
  NAND2_X1 g188 ( .A1(new_n307_), .A2(new_n309_), .ZN(new_n311_) );
  NAND2_X1 g189 ( .A1(new_n311_), .A2(new_n258_), .ZN(new_n312_) );
  NAND4_X1 g190 ( .A1(new_n312_), .A2(G469), .A3(new_n124_), .A4(new_n310_), .ZN(new_n313_) );
  INV_X1 g191 ( .A(G469), .ZN(new_n314_) );
  NAND3_X1 g192 ( .A1(new_n312_), .A2(new_n124_), .A3(new_n310_), .ZN(new_n315_) );
  NAND2_X1 g193 ( .A1(new_n315_), .A2(new_n314_), .ZN(new_n316_) );
  NAND2_X1 g194 ( .A1(new_n316_), .A2(new_n313_), .ZN(new_n317_) );
  XNOR2_X1 g195 ( .A(new_n317_), .B(new_n297_), .ZN(new_n318_) );
  INV_X1 g196 ( .A(new_n318_), .ZN(new_n319_) );
  INV_X1 g197 ( .A(G472), .ZN(new_n320_) );
  NAND2_X1 g198 ( .A1(G137), .A2(KEYINPUT5), .ZN(new_n321_) );
  INV_X1 g199 ( .A(G137), .ZN(new_n322_) );
  INV_X1 g200 ( .A(KEYINPUT5), .ZN(new_n323_) );
  NAND2_X1 g201 ( .A1(new_n322_), .A2(new_n323_), .ZN(new_n324_) );
  NAND2_X1 g202 ( .A1(new_n324_), .A2(new_n321_), .ZN(new_n325_) );
  NAND2_X1 g203 ( .A1(new_n184_), .A2(G210), .ZN(new_n326_) );
  NAND2_X1 g204 ( .A1(new_n325_), .A2(new_n326_), .ZN(new_n327_) );
  NAND4_X1 g205 ( .A1(new_n324_), .A2(G210), .A3(new_n184_), .A4(new_n321_), .ZN(new_n328_) );
  NAND2_X1 g206 ( .A1(new_n327_), .A2(new_n328_), .ZN(new_n329_) );
  NAND2_X1 g207 ( .A1(new_n245_), .A2(new_n329_), .ZN(new_n330_) );
  NAND4_X1 g208 ( .A1(new_n243_), .A2(new_n327_), .A3(new_n244_), .A4(new_n328_), .ZN(new_n331_) );
  NAND2_X1 g209 ( .A1(new_n330_), .A2(new_n331_), .ZN(new_n332_) );
  NAND2_X1 g210 ( .A1(new_n332_), .A2(new_n304_), .ZN(new_n333_) );
  NAND4_X1 g211 ( .A1(new_n330_), .A2(new_n300_), .A3(new_n302_), .A4(new_n331_), .ZN(new_n334_) );
  NAND2_X1 g212 ( .A1(new_n333_), .A2(new_n334_), .ZN(new_n335_) );
  NAND2_X1 g213 ( .A1(new_n335_), .A2(new_n214_), .ZN(new_n336_) );
  NAND4_X1 g214 ( .A1(new_n333_), .A2(new_n212_), .A3(new_n213_), .A4(new_n334_), .ZN(new_n337_) );
  NAND4_X1 g215 ( .A1(new_n336_), .A2(new_n320_), .A3(new_n124_), .A4(new_n337_), .ZN(new_n338_) );
  NAND3_X1 g216 ( .A1(new_n336_), .A2(new_n124_), .A3(new_n337_), .ZN(new_n339_) );
  NAND2_X1 g217 ( .A1(new_n339_), .A2(G472), .ZN(new_n340_) );
  NAND2_X1 g218 ( .A1(new_n340_), .A2(new_n338_), .ZN(new_n341_) );
  XNOR2_X1 g219 ( .A(new_n341_), .B(KEYINPUT6), .ZN(new_n342_) );
  NAND2_X1 g220 ( .A1(new_n201_), .A2(G217), .ZN(new_n343_) );
  XNOR2_X1 g221 ( .A(new_n168_), .B(new_n298_), .ZN(new_n344_) );
  XNOR2_X1 g222 ( .A(G119), .B(G146), .ZN(new_n345_) );
  XNOR2_X1 g223 ( .A(G110), .B(G128), .ZN(new_n346_) );
  NAND2_X1 g224 ( .A1(new_n345_), .A2(new_n346_), .ZN(new_n347_) );
  INV_X1 g225 ( .A(new_n345_), .ZN(new_n348_) );
  INV_X1 g226 ( .A(new_n346_), .ZN(new_n349_) );
  NAND2_X1 g227 ( .A1(new_n348_), .A2(new_n349_), .ZN(new_n350_) );
  NAND2_X1 g228 ( .A1(new_n350_), .A2(new_n347_), .ZN(new_n351_) );
  NAND2_X1 g229 ( .A1(new_n344_), .A2(new_n351_), .ZN(new_n352_) );
  XNOR2_X1 g230 ( .A(new_n170_), .B(new_n298_), .ZN(new_n353_) );
  NAND3_X1 g231 ( .A1(new_n353_), .A2(new_n347_), .A3(new_n350_), .ZN(new_n354_) );
  NAND2_X1 g232 ( .A1(new_n352_), .A2(new_n354_), .ZN(new_n355_) );
  NAND2_X1 g233 ( .A1(new_n130_), .A2(G221), .ZN(new_n356_) );
  XNOR2_X1 g234 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(new_n357_) );
  XOR2_X1 g235 ( .A(new_n356_), .B(new_n357_), .Z(new_n358_) );
  NAND2_X1 g236 ( .A1(new_n355_), .A2(new_n358_), .ZN(new_n359_) );
  XNOR2_X1 g237 ( .A(new_n356_), .B(new_n357_), .ZN(new_n360_) );
  NAND3_X1 g238 ( .A1(new_n360_), .A2(new_n352_), .A3(new_n354_), .ZN(new_n361_) );
  NAND4_X1 g239 ( .A1(new_n359_), .A2(new_n124_), .A3(new_n343_), .A4(new_n361_), .ZN(new_n362_) );
  NAND3_X1 g240 ( .A1(new_n359_), .A2(new_n124_), .A3(new_n361_), .ZN(new_n363_) );
  NAND3_X1 g241 ( .A1(new_n363_), .A2(G217), .A3(new_n201_), .ZN(new_n364_) );
  NAND3_X1 g242 ( .A1(new_n364_), .A2(KEYINPUT25), .A3(new_n362_), .ZN(new_n365_) );
  INV_X1 g243 ( .A(KEYINPUT25), .ZN(new_n366_) );
  NAND2_X1 g244 ( .A1(new_n364_), .A2(new_n362_), .ZN(new_n367_) );
  NAND2_X1 g245 ( .A1(new_n367_), .A2(new_n366_), .ZN(new_n368_) );
  NAND2_X1 g246 ( .A1(new_n368_), .A2(new_n365_), .ZN(new_n369_) );
  INV_X1 g247 ( .A(new_n369_), .ZN(new_n370_) );
  NAND4_X1 g248 ( .A1(new_n296_), .A2(new_n319_), .A3(new_n342_), .A4(new_n370_), .ZN(new_n371_) );
  XNOR2_X1 g249 ( .A(new_n371_), .B(G101), .ZN(G3) );
  NAND3_X1 g250 ( .A1(new_n368_), .A2(new_n203_), .A3(new_n365_), .ZN(new_n373_) );
  NOR3_X1 g251 ( .A1(new_n373_), .A2(new_n317_), .A3(new_n341_), .ZN(new_n374_) );
  NAND3_X1 g252 ( .A1(new_n292_), .A2(new_n290_), .A3(new_n374_), .ZN(new_n375_) );
  INV_X1 g253 ( .A(new_n375_), .ZN(new_n376_) );
  INV_X1 g254 ( .A(new_n196_), .ZN(new_n377_) );
  NAND2_X1 g255 ( .A1(new_n377_), .A2(new_n160_), .ZN(new_n378_) );
  INV_X1 g256 ( .A(new_n378_), .ZN(new_n379_) );
  NAND2_X1 g257 ( .A1(new_n376_), .A2(new_n379_), .ZN(new_n380_) );
  XNOR2_X1 g258 ( .A(new_n380_), .B(G104), .ZN(G6) );
  INV_X1 g259 ( .A(new_n160_), .ZN(new_n382_) );
  NAND2_X1 g260 ( .A1(new_n382_), .A2(new_n196_), .ZN(new_n383_) );
  INV_X1 g261 ( .A(new_n383_), .ZN(new_n384_) );
  NAND2_X1 g262 ( .A1(new_n376_), .A2(new_n384_), .ZN(new_n385_) );
  XNOR2_X1 g263 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(new_n386_) );
  XNOR2_X1 g264 ( .A(new_n385_), .B(new_n386_), .ZN(new_n387_) );
  XNOR2_X1 g265 ( .A(new_n387_), .B(new_n141_), .ZN(G9) );
  INV_X1 g266 ( .A(new_n341_), .ZN(new_n389_) );
  NAND4_X1 g267 ( .A1(new_n296_), .A2(new_n319_), .A3(new_n389_), .A4(new_n369_), .ZN(new_n390_) );
  XNOR2_X1 g268 ( .A(new_n390_), .B(G110), .ZN(G12) );
  INV_X1 g269 ( .A(new_n279_), .ZN(new_n392_) );
  INV_X1 g270 ( .A(new_n317_), .ZN(new_n393_) );
  INV_X1 g271 ( .A(KEYINPUT28), .ZN(new_n394_) );
  INV_X1 g272 ( .A(G900), .ZN(new_n395_) );
  NAND3_X1 g273 ( .A1(new_n284_), .A2(new_n395_), .A3(G953), .ZN(new_n396_) );
  NAND2_X1 g274 ( .A1(new_n396_), .A2(new_n288_), .ZN(new_n397_) );
  NAND2_X1 g275 ( .A1(new_n203_), .A2(new_n397_), .ZN(new_n398_) );
  INV_X1 g276 ( .A(new_n398_), .ZN(new_n399_) );
  NAND4_X1 g277 ( .A1(new_n369_), .A2(new_n394_), .A3(new_n341_), .A4(new_n399_), .ZN(new_n400_) );
  NAND3_X1 g278 ( .A1(new_n369_), .A2(new_n341_), .A3(new_n399_), .ZN(new_n401_) );
  NAND2_X1 g279 ( .A1(new_n401_), .A2(KEYINPUT28), .ZN(new_n402_) );
  NAND3_X1 g280 ( .A1(new_n402_), .A2(new_n393_), .A3(new_n400_), .ZN(new_n403_) );
  NOR2_X1 g281 ( .A1(new_n403_), .A2(new_n392_), .ZN(new_n404_) );
  NAND2_X1 g282 ( .A1(new_n404_), .A2(new_n384_), .ZN(new_n405_) );
  XOR2_X1 g283 ( .A(G128), .B(KEYINPUT29), .Z(new_n406_) );
  XNOR2_X1 g284 ( .A(new_n405_), .B(new_n406_), .ZN(G30) );
  INV_X1 g285 ( .A(KEYINPUT30), .ZN(new_n408_) );
  NAND2_X1 g286 ( .A1(new_n341_), .A2(new_n274_), .ZN(new_n409_) );
  NAND2_X1 g287 ( .A1(new_n409_), .A2(new_n408_), .ZN(new_n410_) );
  NAND3_X1 g288 ( .A1(new_n341_), .A2(KEYINPUT30), .A3(new_n274_), .ZN(new_n411_) );
  NAND2_X1 g289 ( .A1(new_n410_), .A2(new_n411_), .ZN(new_n412_) );
  INV_X1 g290 ( .A(new_n397_), .ZN(new_n413_) );
  NOR3_X1 g291 ( .A1(new_n373_), .A2(new_n317_), .A3(new_n413_), .ZN(new_n414_) );
  NOR2_X1 g292 ( .A1(new_n160_), .A2(new_n196_), .ZN(new_n415_) );
  NAND4_X1 g293 ( .A1(new_n414_), .A2(new_n412_), .A3(new_n415_), .A4(new_n273_), .ZN(new_n416_) );
  XNOR2_X1 g294 ( .A(new_n416_), .B(G143), .ZN(G45) );
  NAND2_X1 g295 ( .A1(new_n404_), .A2(new_n379_), .ZN(new_n418_) );
  XNOR2_X1 g296 ( .A(new_n418_), .B(G146), .ZN(G48) );
  INV_X1 g297 ( .A(KEYINPUT31), .ZN(new_n420_) );
  INV_X1 g298 ( .A(new_n373_), .ZN(new_n421_) );
  NAND3_X1 g299 ( .A1(new_n318_), .A2(new_n341_), .A3(new_n421_), .ZN(new_n422_) );
  INV_X1 g300 ( .A(new_n422_), .ZN(new_n423_) );
  NAND4_X1 g301 ( .A1(new_n292_), .A2(new_n420_), .A3(new_n290_), .A4(new_n423_), .ZN(new_n424_) );
  NAND3_X1 g302 ( .A1(new_n292_), .A2(new_n290_), .A3(new_n423_), .ZN(new_n425_) );
  NAND2_X1 g303 ( .A1(new_n425_), .A2(KEYINPUT31), .ZN(new_n426_) );
  NAND2_X1 g304 ( .A1(new_n426_), .A2(new_n424_), .ZN(new_n427_) );
  NAND2_X1 g305 ( .A1(new_n427_), .A2(new_n379_), .ZN(new_n428_) );
  XNOR2_X1 g306 ( .A(new_n428_), .B(G113), .ZN(G15) );
  NAND2_X1 g307 ( .A1(new_n427_), .A2(new_n384_), .ZN(new_n430_) );
  XNOR2_X1 g308 ( .A(new_n430_), .B(G116), .ZN(G18) );
  INV_X1 g309 ( .A(KEYINPUT6), .ZN(new_n432_) );
  XNOR2_X1 g310 ( .A(new_n341_), .B(new_n432_), .ZN(new_n433_) );
  NOR3_X1 g311 ( .A1(new_n319_), .A2(new_n433_), .A3(new_n370_), .ZN(new_n434_) );
  NAND2_X1 g312 ( .A1(new_n296_), .A2(new_n434_), .ZN(new_n435_) );
  NAND2_X1 g313 ( .A1(new_n435_), .A2(KEYINPUT32), .ZN(new_n436_) );
  INV_X1 g314 ( .A(KEYINPUT32), .ZN(new_n437_) );
  NAND3_X1 g315 ( .A1(new_n296_), .A2(new_n437_), .A3(new_n434_), .ZN(new_n438_) );
  NAND2_X1 g316 ( .A1(new_n436_), .A2(new_n438_), .ZN(new_n439_) );
  XNOR2_X1 g317 ( .A(new_n439_), .B(G119), .ZN(G21) );
  INV_X1 g318 ( .A(KEYINPUT35), .ZN(new_n441_) );
  INV_X1 g319 ( .A(KEYINPUT33), .ZN(new_n442_) );
  NAND4_X1 g320 ( .A1(new_n318_), .A2(new_n433_), .A3(new_n442_), .A4(new_n421_), .ZN(new_n443_) );
  NAND3_X1 g321 ( .A1(new_n318_), .A2(new_n433_), .A3(new_n421_), .ZN(new_n444_) );
  NAND2_X1 g322 ( .A1(new_n444_), .A2(KEYINPUT33), .ZN(new_n445_) );
  NAND2_X1 g323 ( .A1(new_n445_), .A2(new_n443_), .ZN(new_n446_) );
  NAND4_X1 g324 ( .A1(new_n446_), .A2(new_n292_), .A3(KEYINPUT34), .A4(new_n290_), .ZN(new_n447_) );
  INV_X1 g325 ( .A(KEYINPUT34), .ZN(new_n448_) );
  NAND3_X1 g326 ( .A1(new_n446_), .A2(new_n292_), .A3(new_n290_), .ZN(new_n449_) );
  NAND2_X1 g327 ( .A1(new_n449_), .A2(new_n448_), .ZN(new_n450_) );
  NAND2_X1 g328 ( .A1(new_n450_), .A2(new_n447_), .ZN(new_n451_) );
  NAND2_X1 g329 ( .A1(new_n451_), .A2(new_n415_), .ZN(new_n452_) );
  NAND2_X1 g330 ( .A1(new_n452_), .A2(new_n441_), .ZN(new_n453_) );
  NAND3_X1 g331 ( .A1(new_n451_), .A2(KEYINPUT35), .A3(new_n415_), .ZN(new_n454_) );
  NAND2_X1 g332 ( .A1(new_n453_), .A2(new_n454_), .ZN(new_n455_) );
  XNOR2_X1 g333 ( .A(new_n455_), .B(G122), .ZN(G24) );
  INV_X1 g334 ( .A(KEYINPUT36), .ZN(new_n457_) );
  NAND4_X1 g335 ( .A1(new_n379_), .A2(new_n433_), .A3(new_n369_), .A4(new_n399_), .ZN(new_n458_) );
  NOR2_X1 g336 ( .A1(new_n458_), .A2(new_n275_), .ZN(new_n459_) );
  NAND2_X1 g337 ( .A1(new_n459_), .A2(new_n457_), .ZN(new_n460_) );
  NOR2_X1 g338 ( .A1(new_n459_), .A2(new_n457_), .ZN(new_n461_) );
  NOR2_X1 g339 ( .A1(new_n461_), .A2(new_n319_), .ZN(new_n462_) );
  NAND2_X1 g340 ( .A1(new_n462_), .A2(new_n460_), .ZN(new_n463_) );
  XNOR2_X1 g341 ( .A(new_n463_), .B(G125), .ZN(new_n464_) );
  XOR2_X1 g342 ( .A(new_n464_), .B(KEYINPUT37), .Z(G27) );
  NAND2_X1 g343 ( .A1(new_n273_), .A2(KEYINPUT38), .ZN(new_n466_) );
  INV_X1 g344 ( .A(KEYINPUT38), .ZN(new_n467_) );
  NAND3_X1 g345 ( .A1(new_n271_), .A2(new_n467_), .A3(new_n272_), .ZN(new_n468_) );
  NAND4_X1 g346 ( .A1(new_n414_), .A2(new_n412_), .A3(new_n466_), .A4(new_n468_), .ZN(new_n469_) );
  NAND2_X1 g347 ( .A1(new_n469_), .A2(KEYINPUT39), .ZN(new_n470_) );
  INV_X1 g348 ( .A(KEYINPUT39), .ZN(new_n471_) );
  XNOR2_X1 g349 ( .A(new_n273_), .B(new_n467_), .ZN(new_n472_) );
  NAND4_X1 g350 ( .A1(new_n472_), .A2(new_n471_), .A3(new_n414_), .A4(new_n412_), .ZN(new_n473_) );
  NAND2_X1 g351 ( .A1(new_n470_), .A2(new_n473_), .ZN(new_n474_) );
  NAND2_X1 g352 ( .A1(new_n474_), .A2(new_n379_), .ZN(new_n475_) );
  NAND2_X1 g353 ( .A1(new_n475_), .A2(KEYINPUT40), .ZN(new_n476_) );
  INV_X1 g354 ( .A(KEYINPUT40), .ZN(new_n477_) );
  NAND3_X1 g355 ( .A1(new_n474_), .A2(new_n477_), .A3(new_n379_), .ZN(new_n478_) );
  NAND2_X1 g356 ( .A1(new_n476_), .A2(new_n478_), .ZN(new_n479_) );
  XNOR2_X1 g357 ( .A(new_n479_), .B(G131), .ZN(G33) );
  NAND2_X1 g358 ( .A1(new_n474_), .A2(new_n384_), .ZN(new_n481_) );
  XNOR2_X1 g359 ( .A(new_n481_), .B(G134), .ZN(G36) );
  INV_X1 g360 ( .A(new_n403_), .ZN(new_n483_) );
  INV_X1 g361 ( .A(KEYINPUT41), .ZN(new_n484_) );
  NAND4_X1 g362 ( .A1(new_n472_), .A2(new_n198_), .A3(new_n484_), .A4(new_n274_), .ZN(new_n485_) );
  NAND3_X1 g363 ( .A1(new_n472_), .A2(new_n198_), .A3(new_n274_), .ZN(new_n486_) );
  NAND2_X1 g364 ( .A1(new_n486_), .A2(KEYINPUT41), .ZN(new_n487_) );
  NAND2_X1 g365 ( .A1(new_n487_), .A2(new_n485_), .ZN(new_n488_) );
  NAND2_X1 g366 ( .A1(new_n488_), .A2(new_n483_), .ZN(new_n489_) );
  NAND2_X1 g367 ( .A1(new_n489_), .A2(KEYINPUT42), .ZN(new_n490_) );
  INV_X1 g368 ( .A(KEYINPUT42), .ZN(new_n491_) );
  NAND3_X1 g369 ( .A1(new_n488_), .A2(new_n491_), .A3(new_n483_), .ZN(new_n492_) );
  NAND2_X1 g370 ( .A1(new_n490_), .A2(new_n492_), .ZN(new_n493_) );
  XNOR2_X1 g371 ( .A(new_n493_), .B(G137), .ZN(G39) );
  INV_X1 g372 ( .A(new_n274_), .ZN(new_n495_) );
  NOR3_X1 g373 ( .A1(new_n458_), .A2(new_n495_), .A3(new_n318_), .ZN(new_n496_) );
  NAND2_X1 g374 ( .A1(new_n496_), .A2(KEYINPUT43), .ZN(new_n497_) );
  NOR2_X1 g375 ( .A1(new_n496_), .A2(KEYINPUT43), .ZN(new_n498_) );
  NOR2_X1 g376 ( .A1(new_n498_), .A2(new_n273_), .ZN(new_n499_) );
  NAND2_X1 g377 ( .A1(new_n499_), .A2(new_n497_), .ZN(new_n500_) );
  XNOR2_X1 g378 ( .A(new_n500_), .B(G140), .ZN(G42) );
  INV_X1 g379 ( .A(KEYINPUT2), .ZN(new_n502_) );
  INV_X1 g380 ( .A(KEYINPUT48), .ZN(new_n503_) );
  NAND3_X1 g381 ( .A1(new_n493_), .A2(new_n479_), .A3(KEYINPUT46), .ZN(new_n504_) );
  INV_X1 g382 ( .A(KEYINPUT46), .ZN(new_n505_) );
  NAND2_X1 g383 ( .A1(new_n493_), .A2(new_n479_), .ZN(new_n506_) );
  NAND2_X1 g384 ( .A1(new_n506_), .A2(new_n505_), .ZN(new_n507_) );
  NAND2_X1 g385 ( .A1(new_n507_), .A2(new_n504_), .ZN(new_n508_) );
  NAND2_X1 g386 ( .A1(new_n463_), .A2(new_n416_), .ZN(new_n509_) );
  NAND2_X1 g387 ( .A1(new_n383_), .A2(new_n378_), .ZN(new_n510_) );
  NAND2_X1 g388 ( .A1(new_n404_), .A2(new_n510_), .ZN(new_n511_) );
  XNOR2_X1 g389 ( .A(new_n511_), .B(KEYINPUT47), .ZN(new_n512_) );
  NOR2_X1 g390 ( .A1(new_n509_), .A2(new_n512_), .ZN(new_n513_) );
  NAND3_X1 g391 ( .A1(new_n508_), .A2(new_n503_), .A3(new_n513_), .ZN(new_n514_) );
  NAND2_X1 g392 ( .A1(new_n508_), .A2(new_n513_), .ZN(new_n515_) );
  NAND2_X1 g393 ( .A1(new_n515_), .A2(KEYINPUT48), .ZN(new_n516_) );
  NAND2_X1 g394 ( .A1(new_n500_), .A2(new_n481_), .ZN(new_n517_) );
  INV_X1 g395 ( .A(new_n517_), .ZN(new_n518_) );
  NAND3_X1 g396 ( .A1(new_n516_), .A2(new_n514_), .A3(new_n518_), .ZN(new_n519_) );
  INV_X1 g397 ( .A(new_n519_), .ZN(new_n520_) );
  INV_X1 g398 ( .A(KEYINPUT44), .ZN(new_n521_) );
  NAND4_X1 g399 ( .A1(new_n455_), .A2(new_n439_), .A3(new_n521_), .A4(new_n390_), .ZN(new_n522_) );
  NAND2_X1 g400 ( .A1(new_n439_), .A2(new_n390_), .ZN(new_n523_) );
  NAND2_X1 g401 ( .A1(new_n523_), .A2(KEYINPUT44), .ZN(new_n524_) );
  NAND3_X1 g402 ( .A1(new_n453_), .A2(KEYINPUT44), .A3(new_n454_), .ZN(new_n525_) );
  NAND3_X1 g403 ( .A1(new_n426_), .A2(new_n375_), .A3(new_n424_), .ZN(new_n526_) );
  NAND2_X1 g404 ( .A1(new_n526_), .A2(new_n510_), .ZN(new_n527_) );
  NAND2_X1 g405 ( .A1(new_n371_), .A2(new_n527_), .ZN(new_n528_) );
  INV_X1 g406 ( .A(new_n528_), .ZN(new_n529_) );
  NAND2_X1 g407 ( .A1(new_n525_), .A2(new_n529_), .ZN(new_n530_) );
  INV_X1 g408 ( .A(new_n530_), .ZN(new_n531_) );
  NAND4_X1 g409 ( .A1(new_n531_), .A2(new_n524_), .A3(KEYINPUT45), .A4(new_n522_), .ZN(new_n532_) );
  INV_X1 g410 ( .A(KEYINPUT45), .ZN(new_n533_) );
  NAND3_X1 g411 ( .A1(new_n531_), .A2(new_n524_), .A3(new_n522_), .ZN(new_n534_) );
  NAND2_X1 g412 ( .A1(new_n534_), .A2(new_n533_), .ZN(new_n535_) );
  NAND3_X1 g413 ( .A1(new_n520_), .A2(new_n532_), .A3(new_n535_), .ZN(new_n536_) );
  NAND2_X1 g414 ( .A1(new_n536_), .A2(new_n502_), .ZN(new_n537_) );
  NAND4_X1 g415 ( .A1(new_n520_), .A2(new_n535_), .A3(KEYINPUT2), .A4(new_n532_), .ZN(new_n538_) );
  NAND2_X1 g416 ( .A1(new_n537_), .A2(new_n538_), .ZN(new_n539_) );
  NAND3_X1 g417 ( .A1(new_n319_), .A2(KEYINPUT50), .A3(new_n373_), .ZN(new_n540_) );
  INV_X1 g418 ( .A(KEYINPUT50), .ZN(new_n541_) );
  NAND2_X1 g419 ( .A1(new_n319_), .A2(new_n373_), .ZN(new_n542_) );
  NAND2_X1 g420 ( .A1(new_n542_), .A2(new_n541_), .ZN(new_n543_) );
  INV_X1 g421 ( .A(new_n203_), .ZN(new_n544_) );
  NAND2_X1 g422 ( .A1(new_n369_), .A2(new_n544_), .ZN(new_n545_) );
  XOR2_X1 g423 ( .A(new_n545_), .B(KEYINPUT49), .Z(new_n546_) );
  NAND4_X1 g424 ( .A1(new_n546_), .A2(new_n543_), .A3(new_n389_), .A4(new_n540_), .ZN(new_n547_) );
  NAND2_X1 g425 ( .A1(new_n547_), .A2(new_n422_), .ZN(new_n548_) );
  NAND2_X1 g426 ( .A1(new_n548_), .A2(KEYINPUT51), .ZN(new_n549_) );
  INV_X1 g427 ( .A(KEYINPUT51), .ZN(new_n550_) );
  NAND3_X1 g428 ( .A1(new_n547_), .A2(new_n550_), .A3(new_n422_), .ZN(new_n551_) );
  NAND3_X1 g429 ( .A1(new_n549_), .A2(new_n488_), .A3(new_n551_), .ZN(new_n552_) );
  NAND3_X1 g430 ( .A1(new_n510_), .A2(new_n274_), .A3(new_n472_), .ZN(new_n553_) );
  INV_X1 g431 ( .A(new_n472_), .ZN(new_n554_) );
  NAND2_X1 g432 ( .A1(new_n554_), .A2(new_n495_), .ZN(new_n555_) );
  NAND2_X1 g433 ( .A1(new_n555_), .A2(new_n198_), .ZN(new_n556_) );
  NAND2_X1 g434 ( .A1(new_n556_), .A2(new_n553_), .ZN(new_n557_) );
  NAND2_X1 g435 ( .A1(new_n557_), .A2(new_n446_), .ZN(new_n558_) );
  NAND3_X1 g436 ( .A1(new_n552_), .A2(KEYINPUT52), .A3(new_n558_), .ZN(new_n559_) );
  INV_X1 g437 ( .A(KEYINPUT52), .ZN(new_n560_) );
  NAND2_X1 g438 ( .A1(new_n552_), .A2(new_n558_), .ZN(new_n561_) );
  NAND2_X1 g439 ( .A1(new_n561_), .A2(new_n560_), .ZN(new_n562_) );
  NAND3_X1 g440 ( .A1(new_n562_), .A2(new_n287_), .A3(new_n559_), .ZN(new_n563_) );
  NAND2_X1 g441 ( .A1(new_n488_), .A2(new_n446_), .ZN(new_n564_) );
  NAND4_X1 g442 ( .A1(new_n539_), .A2(new_n126_), .A3(new_n563_), .A4(new_n564_), .ZN(new_n565_) );
  XOR2_X1 g443 ( .A(new_n565_), .B(KEYINPUT53), .Z(G75) );
  INV_X1 g444 ( .A(KEYINPUT56), .ZN(new_n567_) );
  INV_X1 g445 ( .A(new_n199_), .ZN(new_n568_) );
  XNOR2_X1 g446 ( .A(new_n536_), .B(KEYINPUT2), .ZN(new_n569_) );
  XNOR2_X1 g447 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(new_n570_) );
  XNOR2_X1 g448 ( .A(new_n265_), .B(new_n570_), .ZN(new_n571_) );
  INV_X1 g449 ( .A(new_n571_), .ZN(new_n572_) );
  NAND4_X1 g450 ( .A1(new_n569_), .A2(G210), .A3(new_n568_), .A4(new_n572_), .ZN(new_n573_) );
  NAND4_X1 g451 ( .A1(new_n537_), .A2(G210), .A3(new_n568_), .A4(new_n538_), .ZN(new_n574_) );
  NAND2_X1 g452 ( .A1(new_n574_), .A2(new_n571_), .ZN(new_n575_) );
  NOR2_X1 g453 ( .A1(new_n126_), .A2(G952), .ZN(new_n576_) );
  INV_X1 g454 ( .A(new_n576_), .ZN(new_n577_) );
  NAND3_X1 g455 ( .A1(new_n573_), .A2(new_n575_), .A3(new_n577_), .ZN(new_n578_) );
  XNOR2_X1 g456 ( .A(new_n578_), .B(new_n567_), .ZN(G51) );
  NAND2_X1 g457 ( .A1(new_n312_), .A2(new_n310_), .ZN(new_n580_) );
  XOR2_X1 g458 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(new_n581_) );
  NAND4_X1 g459 ( .A1(new_n537_), .A2(G469), .A3(new_n568_), .A4(new_n538_), .ZN(new_n582_) );
  NOR2_X1 g460 ( .A1(new_n582_), .A2(new_n581_), .ZN(new_n583_) );
  NAND2_X1 g461 ( .A1(new_n582_), .A2(new_n581_), .ZN(new_n584_) );
  INV_X1 g462 ( .A(new_n584_), .ZN(new_n585_) );
  NOR3_X1 g463 ( .A1(new_n585_), .A2(new_n580_), .A3(new_n583_), .ZN(new_n586_) );
  INV_X1 g464 ( .A(new_n580_), .ZN(new_n587_) );
  INV_X1 g465 ( .A(new_n581_), .ZN(new_n588_) );
  XNOR2_X1 g466 ( .A(new_n582_), .B(new_n588_), .ZN(new_n589_) );
  NOR2_X1 g467 ( .A1(new_n589_), .A2(new_n587_), .ZN(new_n590_) );
  NOR3_X1 g468 ( .A1(new_n590_), .A2(new_n586_), .A3(new_n576_), .ZN(G54) );
  INV_X1 g469 ( .A(KEYINPUT60), .ZN(new_n592_) );
  XNOR2_X1 g470 ( .A(new_n190_), .B(KEYINPUT59), .ZN(new_n593_) );
  INV_X1 g471 ( .A(new_n593_), .ZN(new_n594_) );
  NAND4_X1 g472 ( .A1(new_n569_), .A2(G475), .A3(new_n568_), .A4(new_n594_), .ZN(new_n595_) );
  NAND4_X1 g473 ( .A1(new_n537_), .A2(G475), .A3(new_n568_), .A4(new_n538_), .ZN(new_n596_) );
  NAND2_X1 g474 ( .A1(new_n596_), .A2(new_n593_), .ZN(new_n597_) );
  NAND3_X1 g475 ( .A1(new_n595_), .A2(new_n577_), .A3(new_n597_), .ZN(new_n598_) );
  XNOR2_X1 g476 ( .A(new_n598_), .B(new_n592_), .ZN(G60) );
  NAND2_X1 g477 ( .A1(new_n154_), .A2(new_n155_), .ZN(new_n600_) );
  NAND3_X1 g478 ( .A1(new_n569_), .A2(G478), .A3(new_n568_), .ZN(new_n601_) );
  NOR2_X1 g479 ( .A1(new_n601_), .A2(new_n600_), .ZN(new_n602_) );
  NAND2_X1 g480 ( .A1(new_n601_), .A2(new_n600_), .ZN(new_n603_) );
  INV_X1 g481 ( .A(new_n603_), .ZN(new_n604_) );
  NOR3_X1 g482 ( .A1(new_n604_), .A2(new_n602_), .A3(new_n576_), .ZN(G63) );
  NAND2_X1 g483 ( .A1(new_n359_), .A2(new_n361_), .ZN(new_n606_) );
  NAND3_X1 g484 ( .A1(new_n569_), .A2(G217), .A3(new_n568_), .ZN(new_n607_) );
  NOR2_X1 g485 ( .A1(new_n607_), .A2(new_n606_), .ZN(new_n608_) );
  NAND2_X1 g486 ( .A1(new_n607_), .A2(new_n606_), .ZN(new_n609_) );
  INV_X1 g487 ( .A(new_n609_), .ZN(new_n610_) );
  NOR3_X1 g488 ( .A1(new_n610_), .A2(new_n608_), .A3(new_n576_), .ZN(G66) );
  NAND3_X1 g489 ( .A1(new_n535_), .A2(new_n126_), .A3(new_n532_), .ZN(new_n612_) );
  NAND3_X1 g490 ( .A1(G224), .A2(G953), .A3(KEYINPUT61), .ZN(new_n613_) );
  INV_X1 g491 ( .A(KEYINPUT61), .ZN(new_n614_) );
  NAND2_X1 g492 ( .A1(G224), .A2(G953), .ZN(new_n615_) );
  NAND2_X1 g493 ( .A1(new_n615_), .A2(new_n614_), .ZN(new_n616_) );
  NAND3_X1 g494 ( .A1(new_n616_), .A2(G898), .A3(new_n613_), .ZN(new_n617_) );
  NAND2_X1 g495 ( .A1(new_n612_), .A2(new_n617_), .ZN(new_n618_) );
  NAND2_X1 g496 ( .A1(new_n280_), .A2(G953), .ZN(new_n619_) );
  XNOR2_X1 g497 ( .A(new_n216_), .B(new_n207_), .ZN(new_n620_) );
  NAND2_X1 g498 ( .A1(new_n620_), .A2(new_n250_), .ZN(new_n621_) );
  INV_X1 g499 ( .A(new_n620_), .ZN(new_n622_) );
  NAND3_X1 g500 ( .A1(new_n622_), .A2(new_n247_), .A3(new_n249_), .ZN(new_n623_) );
  NAND3_X1 g501 ( .A1(new_n623_), .A2(new_n619_), .A3(new_n621_), .ZN(new_n624_) );
  XOR2_X1 g502 ( .A(new_n618_), .B(new_n624_), .Z(G69) );
  XNOR2_X1 g503 ( .A(new_n211_), .B(new_n168_), .ZN(new_n626_) );
  XNOR2_X1 g504 ( .A(new_n626_), .B(new_n306_), .ZN(new_n627_) );
  XNOR2_X1 g505 ( .A(new_n519_), .B(new_n627_), .ZN(new_n628_) );
  NAND2_X1 g506 ( .A1(new_n628_), .A2(new_n126_), .ZN(new_n629_) );
  XNOR2_X1 g507 ( .A(new_n627_), .B(G227), .ZN(new_n630_) );
  NAND2_X1 g508 ( .A1(new_n630_), .A2(G900), .ZN(new_n631_) );
  NAND2_X1 g509 ( .A1(new_n631_), .A2(G953), .ZN(new_n632_) );
  NAND2_X1 g510 ( .A1(new_n629_), .A2(new_n632_), .ZN(G72) );
  NAND2_X1 g511 ( .A1(new_n336_), .A2(new_n337_), .ZN(new_n634_) );
  XNOR2_X1 g512 ( .A(new_n634_), .B(KEYINPUT62), .ZN(new_n635_) );
  INV_X1 g513 ( .A(new_n635_), .ZN(new_n636_) );
  NAND4_X1 g514 ( .A1(new_n569_), .A2(G472), .A3(new_n568_), .A4(new_n636_), .ZN(new_n637_) );
  NAND4_X1 g515 ( .A1(new_n537_), .A2(G472), .A3(new_n568_), .A4(new_n538_), .ZN(new_n638_) );
  NAND2_X1 g516 ( .A1(new_n638_), .A2(new_n635_), .ZN(new_n639_) );
  NAND3_X1 g517 ( .A1(new_n637_), .A2(new_n577_), .A3(new_n639_), .ZN(new_n640_) );
  XNOR2_X1 g518 ( .A(new_n640_), .B(KEYINPUT63), .ZN(G57) );
endmodule


