module locked_c2670 (  G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,  G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397, G329, G231, G308, G225  );
  input  G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire new_n359_, new_n360_, new_n361_, new_n362_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n385_, new_n386_, new_n389_, new_n390_, new_n391_, new_n392_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n401_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n416_, new_n417_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n574_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n632_, new_n633_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n642_, new_n643_, new_n644_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_;
  AND2_X1 g0000 ( .A1(G44), .A2(KEYINPUT3), .ZN(new_n359_) );
  INV_X1 g0001 ( .A(new_n359_), .ZN(new_n360_) );
  OR2_X1 g0002 ( .A1(G44), .A2(KEYINPUT3), .ZN(new_n361_) );
  AND2_X1 g0003 ( .A1(new_n360_), .A2(new_n361_), .ZN(new_n362_) );
  INV_X1 g0004 ( .A(new_n362_), .ZN(G218) );
  INV_X1 g0005 ( .A(G132), .ZN(G219) );
  INV_X1 g0006 ( .A(G82), .ZN(G220) );
  INV_X1 g0007 ( .A(G96), .ZN(G221) );
  INV_X1 g0008 ( .A(G69), .ZN(G235) );
  INV_X1 g0009 ( .A(G120), .ZN(G236) );
  INV_X1 g0010 ( .A(G57), .ZN(G237) );
  INV_X1 g0011 ( .A(G108), .ZN(G238) );
  INV_X1 g0012 ( .A(G2072), .ZN(new_n371_) );
  INV_X1 g0013 ( .A(KEYINPUT21), .ZN(new_n372_) );
  INV_X1 g0014 ( .A(KEYINPUT20), .ZN(new_n373_) );
  AND2_X1 g0015 ( .A1(G2078), .A2(G2084), .ZN(new_n374_) );
  AND2_X1 g0016 ( .A1(new_n374_), .A2(new_n373_), .ZN(new_n375_) );
  INV_X1 g0017 ( .A(new_n375_), .ZN(new_n376_) );
  OR2_X1 g0018 ( .A1(new_n374_), .A2(new_n373_), .ZN(new_n377_) );
  AND2_X1 g0019 ( .A1(new_n377_), .A2(G2090), .ZN(new_n378_) );
  AND2_X1 g0020 ( .A1(new_n378_), .A2(new_n376_), .ZN(new_n379_) );
  AND2_X1 g0021 ( .A1(new_n379_), .A2(new_n372_), .ZN(new_n380_) );
  INV_X1 g0022 ( .A(new_n380_), .ZN(new_n381_) );
  OR2_X1 g0023 ( .A1(new_n379_), .A2(new_n372_), .ZN(new_n382_) );
  AND2_X1 g0024 ( .A1(new_n381_), .A2(new_n382_), .ZN(new_n383_) );
  OR2_X1 g0025 ( .A1(new_n383_), .A2(new_n371_), .ZN(G158) );
  AND2_X1 g0026 ( .A1(G2), .A2(G15), .ZN(new_n385_) );
  AND2_X1 g0027 ( .A1(new_n385_), .A2(G661), .ZN(new_n386_) );
  INV_X1 g0028 ( .A(new_n386_), .ZN(G259) );
  AND2_X1 g0029 ( .A1(G94), .A2(G452), .ZN(G173) );
  AND2_X1 g0030 ( .A1(G7), .A2(G661), .ZN(new_n389_) );
  AND2_X1 g0031 ( .A1(new_n389_), .A2(KEYINPUT10), .ZN(new_n390_) );
  INV_X1 g0032 ( .A(new_n390_), .ZN(new_n391_) );
  OR2_X1 g0033 ( .A1(new_n389_), .A2(KEYINPUT10), .ZN(new_n392_) );
  AND2_X1 g0034 ( .A1(new_n391_), .A2(new_n392_), .ZN(G223) );
  INV_X1 g0035 ( .A(G567), .ZN(new_n394_) );
  OR2_X1 g0036 ( .A1(G223), .A2(new_n394_), .ZN(new_n395_) );
  INV_X1 g0037 ( .A(new_n395_), .ZN(new_n396_) );
  AND2_X1 g0038 ( .A1(new_n396_), .A2(KEYINPUT11), .ZN(new_n397_) );
  INV_X1 g0039 ( .A(KEYINPUT11), .ZN(new_n398_) );
  AND2_X1 g0040 ( .A1(new_n395_), .A2(new_n398_), .ZN(new_n399_) );
  OR2_X1 g0041 ( .A1(new_n397_), .A2(new_n399_), .ZN(G234) );
  INV_X1 g0042 ( .A(G2106), .ZN(new_n401_) );
  OR2_X1 g0043 ( .A1(G223), .A2(new_n401_), .ZN(G217) );
  AND2_X1 g0044 ( .A1(G82), .A2(G132), .ZN(new_n403_) );
  AND2_X1 g0045 ( .A1(new_n403_), .A2(KEYINPUT22), .ZN(new_n404_) );
  INV_X1 g0046 ( .A(new_n404_), .ZN(new_n405_) );
  OR2_X1 g0047 ( .A1(new_n403_), .A2(KEYINPUT22), .ZN(new_n406_) );
  AND2_X1 g0048 ( .A1(new_n405_), .A2(new_n406_), .ZN(new_n407_) );
  INV_X1 g0049 ( .A(new_n407_), .ZN(new_n408_) );
  AND2_X1 g0050 ( .A1(new_n362_), .A2(G96), .ZN(new_n409_) );
  AND2_X1 g0051 ( .A1(new_n408_), .A2(new_n409_), .ZN(new_n410_) );
  AND2_X1 g0052 ( .A1(G57), .A2(G69), .ZN(new_n411_) );
  AND2_X1 g0053 ( .A1(G108), .A2(G120), .ZN(new_n412_) );
  AND2_X1 g0054 ( .A1(new_n411_), .A2(new_n412_), .ZN(new_n413_) );
  AND2_X1 g0055 ( .A1(new_n410_), .A2(new_n413_), .ZN(G325) );
  INV_X1 g0056 ( .A(G325), .ZN(G261) );
  OR2_X1 g0057 ( .A1(new_n410_), .A2(new_n401_), .ZN(new_n416_) );
  OR2_X1 g0058 ( .A1(new_n413_), .A2(new_n394_), .ZN(new_n417_) );
  AND2_X1 g0059 ( .A1(new_n416_), .A2(new_n417_), .ZN(G319) );
  INV_X1 g0060 ( .A(G137), .ZN(new_n419_) );
  INV_X1 g0061 ( .A(G2104), .ZN(new_n420_) );
  INV_X1 g0062 ( .A(G2105), .ZN(new_n421_) );
  AND2_X1 g0063 ( .A1(new_n420_), .A2(new_n421_), .ZN(new_n422_) );
  AND2_X1 g0064 ( .A1(new_n422_), .A2(KEYINPUT17), .ZN(new_n423_) );
  INV_X1 g0065 ( .A(KEYINPUT17), .ZN(new_n424_) );
  OR2_X1 g0066 ( .A1(G2104), .A2(G2105), .ZN(new_n425_) );
  AND2_X1 g0067 ( .A1(new_n425_), .A2(new_n424_), .ZN(new_n426_) );
  OR2_X1 g0068 ( .A1(new_n423_), .A2(new_n426_), .ZN(new_n427_) );
  OR2_X1 g0069 ( .A1(new_n427_), .A2(new_n419_), .ZN(new_n428_) );
  AND2_X1 g0070 ( .A1(G101), .A2(G2104), .ZN(new_n429_) );
  AND2_X1 g0071 ( .A1(new_n429_), .A2(new_n421_), .ZN(new_n430_) );
  OR2_X1 g0072 ( .A1(new_n430_), .A2(KEYINPUT23), .ZN(new_n431_) );
  INV_X1 g0073 ( .A(new_n431_), .ZN(new_n432_) );
  AND2_X1 g0074 ( .A1(new_n430_), .A2(KEYINPUT23), .ZN(new_n433_) );
  OR2_X1 g0075 ( .A1(new_n432_), .A2(new_n433_), .ZN(new_n434_) );
  AND2_X1 g0076 ( .A1(new_n428_), .A2(new_n434_), .ZN(new_n435_) );
  AND2_X1 g0077 ( .A1(G2104), .A2(G2105), .ZN(new_n436_) );
  AND2_X1 g0078 ( .A1(new_n436_), .A2(G113), .ZN(new_n437_) );
  AND2_X1 g0079 ( .A1(new_n420_), .A2(G2105), .ZN(new_n438_) );
  AND2_X1 g0080 ( .A1(new_n438_), .A2(G125), .ZN(new_n439_) );
  OR2_X1 g0081 ( .A1(new_n439_), .A2(new_n437_), .ZN(new_n440_) );
  INV_X1 g0082 ( .A(new_n440_), .ZN(new_n441_) );
  AND2_X1 g0083 ( .A1(new_n435_), .A2(new_n441_), .ZN(G160) );
  AND2_X1 g0084 ( .A1(new_n438_), .A2(G124), .ZN(new_n443_) );
  INV_X1 g0085 ( .A(new_n443_), .ZN(new_n444_) );
  AND2_X1 g0086 ( .A1(new_n444_), .A2(KEYINPUT44), .ZN(new_n445_) );
  INV_X1 g0087 ( .A(new_n445_), .ZN(new_n446_) );
  OR2_X1 g0088 ( .A1(new_n444_), .A2(KEYINPUT44), .ZN(new_n447_) );
  AND2_X1 g0089 ( .A1(new_n446_), .A2(new_n447_), .ZN(new_n448_) );
  OR2_X1 g0090 ( .A1(new_n425_), .A2(new_n424_), .ZN(new_n449_) );
  OR2_X1 g0091 ( .A1(new_n422_), .A2(KEYINPUT17), .ZN(new_n450_) );
  AND2_X1 g0092 ( .A1(new_n450_), .A2(new_n449_), .ZN(new_n451_) );
  AND2_X1 g0093 ( .A1(new_n451_), .A2(G136), .ZN(new_n452_) );
  AND2_X1 g0094 ( .A1(new_n421_), .A2(G2104), .ZN(new_n453_) );
  AND2_X1 g0095 ( .A1(new_n453_), .A2(G100), .ZN(new_n454_) );
  AND2_X1 g0096 ( .A1(new_n436_), .A2(G112), .ZN(new_n455_) );
  OR2_X1 g0097 ( .A1(new_n454_), .A2(new_n455_), .ZN(new_n456_) );
  OR2_X1 g0098 ( .A1(new_n452_), .A2(new_n456_), .ZN(new_n457_) );
  OR2_X1 g0099 ( .A1(new_n457_), .A2(new_n448_), .ZN(new_n458_) );
  INV_X1 g0100 ( .A(new_n458_), .ZN(G162) );
  AND2_X1 g0101 ( .A1(new_n451_), .A2(G138), .ZN(new_n460_) );
  AND2_X1 g0102 ( .A1(new_n453_), .A2(G102), .ZN(new_n461_) );
  AND2_X1 g0103 ( .A1(new_n436_), .A2(G114), .ZN(new_n462_) );
  AND2_X1 g0104 ( .A1(new_n438_), .A2(G126), .ZN(new_n463_) );
  OR2_X1 g0105 ( .A1(new_n463_), .A2(new_n462_), .ZN(new_n464_) );
  OR2_X1 g0106 ( .A1(new_n464_), .A2(new_n461_), .ZN(new_n465_) );
  OR2_X1 g0107 ( .A1(new_n465_), .A2(new_n460_), .ZN(new_n466_) );
  INV_X1 g0108 ( .A(new_n466_), .ZN(G164) );
  AND2_X1 g0109 ( .A1(G543), .A2(KEYINPUT0), .ZN(new_n468_) );
  INV_X1 g0110 ( .A(new_n468_), .ZN(new_n469_) );
  OR2_X1 g0111 ( .A1(G543), .A2(KEYINPUT0), .ZN(new_n470_) );
  AND2_X1 g0112 ( .A1(new_n469_), .A2(new_n470_), .ZN(new_n471_) );
  OR2_X1 g0113 ( .A1(new_n471_), .A2(G651), .ZN(new_n472_) );
  INV_X1 g0114 ( .A(new_n472_), .ZN(new_n473_) );
  AND2_X1 g0115 ( .A1(new_n473_), .A2(G50), .ZN(new_n474_) );
  INV_X1 g0116 ( .A(G543), .ZN(new_n475_) );
  INV_X1 g0117 ( .A(G651), .ZN(new_n476_) );
  AND2_X1 g0118 ( .A1(new_n475_), .A2(new_n476_), .ZN(new_n477_) );
  AND2_X1 g0119 ( .A1(new_n477_), .A2(G88), .ZN(new_n478_) );
  OR2_X1 g0120 ( .A1(new_n474_), .A2(new_n478_), .ZN(new_n479_) );
  INV_X1 g0121 ( .A(KEYINPUT0), .ZN(new_n480_) );
  AND2_X1 g0122 ( .A1(new_n475_), .A2(new_n480_), .ZN(new_n481_) );
  OR2_X1 g0123 ( .A1(new_n481_), .A2(new_n468_), .ZN(new_n482_) );
  AND2_X1 g0124 ( .A1(new_n482_), .A2(G651), .ZN(new_n483_) );
  AND2_X1 g0125 ( .A1(new_n483_), .A2(G75), .ZN(new_n484_) );
  OR2_X1 g0126 ( .A1(new_n476_), .A2(G543), .ZN(new_n485_) );
  AND2_X1 g0127 ( .A1(new_n485_), .A2(KEYINPUT1), .ZN(new_n486_) );
  INV_X1 g0128 ( .A(KEYINPUT1), .ZN(new_n487_) );
  AND2_X1 g0129 ( .A1(new_n475_), .A2(G651), .ZN(new_n488_) );
  AND2_X1 g0130 ( .A1(new_n488_), .A2(new_n487_), .ZN(new_n489_) );
  OR2_X1 g0131 ( .A1(new_n486_), .A2(new_n489_), .ZN(new_n490_) );
  AND2_X1 g0132 ( .A1(new_n490_), .A2(G62), .ZN(new_n491_) );
  OR2_X1 g0133 ( .A1(new_n491_), .A2(new_n484_), .ZN(new_n492_) );
  OR2_X1 g0134 ( .A1(new_n479_), .A2(new_n492_), .ZN(G303) );
  INV_X1 g0135 ( .A(G303), .ZN(G166) );
  INV_X1 g0136 ( .A(KEYINPUT7), .ZN(new_n495_) );
  AND2_X1 g0137 ( .A1(new_n477_), .A2(G89), .ZN(new_n496_) );
  INV_X1 g0138 ( .A(new_n496_), .ZN(new_n497_) );
  AND2_X1 g0139 ( .A1(new_n497_), .A2(KEYINPUT4), .ZN(new_n498_) );
  INV_X1 g0140 ( .A(new_n498_), .ZN(new_n499_) );
  OR2_X1 g0141 ( .A1(new_n497_), .A2(KEYINPUT4), .ZN(new_n500_) );
  AND2_X1 g0142 ( .A1(new_n499_), .A2(new_n500_), .ZN(new_n501_) );
  AND2_X1 g0143 ( .A1(new_n483_), .A2(G76), .ZN(new_n502_) );
  OR2_X1 g0144 ( .A1(new_n501_), .A2(new_n502_), .ZN(new_n503_) );
  AND2_X1 g0145 ( .A1(new_n503_), .A2(KEYINPUT5), .ZN(new_n504_) );
  INV_X1 g0146 ( .A(new_n504_), .ZN(new_n505_) );
  OR2_X1 g0147 ( .A1(new_n503_), .A2(KEYINPUT5), .ZN(new_n506_) );
  AND2_X1 g0148 ( .A1(new_n505_), .A2(new_n506_), .ZN(new_n507_) );
  INV_X1 g0149 ( .A(KEYINPUT6), .ZN(new_n508_) );
  AND2_X1 g0150 ( .A1(new_n473_), .A2(G51), .ZN(new_n509_) );
  AND2_X1 g0151 ( .A1(new_n490_), .A2(G63), .ZN(new_n510_) );
  OR2_X1 g0152 ( .A1(new_n509_), .A2(new_n510_), .ZN(new_n511_) );
  AND2_X1 g0153 ( .A1(new_n511_), .A2(new_n508_), .ZN(new_n512_) );
  INV_X1 g0154 ( .A(new_n512_), .ZN(new_n513_) );
  OR2_X1 g0155 ( .A1(new_n511_), .A2(new_n508_), .ZN(new_n514_) );
  AND2_X1 g0156 ( .A1(new_n513_), .A2(new_n514_), .ZN(new_n515_) );
  OR2_X1 g0157 ( .A1(new_n507_), .A2(new_n515_), .ZN(new_n516_) );
  AND2_X1 g0158 ( .A1(new_n516_), .A2(new_n495_), .ZN(new_n517_) );
  INV_X1 g0159 ( .A(new_n517_), .ZN(new_n518_) );
  OR2_X1 g0160 ( .A1(new_n516_), .A2(new_n495_), .ZN(new_n519_) );
  AND2_X1 g0161 ( .A1(new_n518_), .A2(new_n519_), .ZN(G168) );
  AND2_X1 g0162 ( .A1(new_n483_), .A2(G77), .ZN(new_n521_) );
  AND2_X1 g0163 ( .A1(new_n477_), .A2(G90), .ZN(new_n522_) );
  OR2_X1 g0164 ( .A1(new_n521_), .A2(new_n522_), .ZN(new_n523_) );
  INV_X1 g0165 ( .A(new_n523_), .ZN(new_n524_) );
  AND2_X1 g0166 ( .A1(new_n524_), .A2(KEYINPUT9), .ZN(new_n525_) );
  INV_X1 g0167 ( .A(new_n525_), .ZN(new_n526_) );
  OR2_X1 g0168 ( .A1(new_n524_), .A2(KEYINPUT9), .ZN(new_n527_) );
  AND2_X1 g0169 ( .A1(new_n473_), .A2(G52), .ZN(new_n528_) );
  AND2_X1 g0170 ( .A1(new_n490_), .A2(G64), .ZN(new_n529_) );
  OR2_X1 g0171 ( .A1(new_n528_), .A2(new_n529_), .ZN(new_n530_) );
  INV_X1 g0172 ( .A(new_n530_), .ZN(new_n531_) );
  AND2_X1 g0173 ( .A1(new_n527_), .A2(new_n531_), .ZN(new_n532_) );
  AND2_X1 g0174 ( .A1(new_n532_), .A2(new_n526_), .ZN(G171) );
  INV_X1 g0175 ( .A(G860), .ZN(new_n534_) );
  INV_X1 g0176 ( .A(KEYINPUT14), .ZN(new_n535_) );
  AND2_X1 g0177 ( .A1(new_n490_), .A2(G56), .ZN(new_n536_) );
  INV_X1 g0178 ( .A(new_n536_), .ZN(new_n537_) );
  OR2_X1 g0179 ( .A1(new_n537_), .A2(new_n535_), .ZN(new_n538_) );
  OR2_X1 g0180 ( .A1(new_n536_), .A2(KEYINPUT14), .ZN(new_n539_) );
  INV_X1 g0181 ( .A(G43), .ZN(new_n540_) );
  OR2_X1 g0182 ( .A1(new_n472_), .A2(new_n540_), .ZN(new_n541_) );
  AND2_X1 g0183 ( .A1(new_n539_), .A2(new_n541_), .ZN(new_n542_) );
  AND2_X1 g0184 ( .A1(new_n542_), .A2(new_n538_), .ZN(new_n543_) );
  INV_X1 g0185 ( .A(KEYINPUT13), .ZN(new_n544_) );
  INV_X1 g0186 ( .A(KEYINPUT12), .ZN(new_n545_) );
  AND2_X1 g0187 ( .A1(new_n477_), .A2(G81), .ZN(new_n546_) );
  OR2_X1 g0188 ( .A1(new_n546_), .A2(new_n545_), .ZN(new_n547_) );
  INV_X1 g0189 ( .A(G81), .ZN(new_n548_) );
  OR2_X1 g0190 ( .A1(G543), .A2(G651), .ZN(new_n549_) );
  OR2_X1 g0191 ( .A1(new_n549_), .A2(new_n548_), .ZN(new_n550_) );
  OR2_X1 g0192 ( .A1(new_n550_), .A2(KEYINPUT12), .ZN(new_n551_) );
  AND2_X1 g0193 ( .A1(new_n547_), .A2(new_n551_), .ZN(new_n552_) );
  AND2_X1 g0194 ( .A1(new_n483_), .A2(G68), .ZN(new_n553_) );
  OR2_X1 g0195 ( .A1(new_n552_), .A2(new_n553_), .ZN(new_n554_) );
  OR2_X1 g0196 ( .A1(new_n554_), .A2(new_n544_), .ZN(new_n555_) );
  AND2_X1 g0197 ( .A1(new_n550_), .A2(KEYINPUT12), .ZN(new_n556_) );
  AND2_X1 g0198 ( .A1(new_n546_), .A2(new_n545_), .ZN(new_n557_) );
  OR2_X1 g0199 ( .A1(new_n557_), .A2(new_n556_), .ZN(new_n558_) );
  INV_X1 g0200 ( .A(G68), .ZN(new_n559_) );
  OR2_X1 g0201 ( .A1(new_n471_), .A2(new_n476_), .ZN(new_n560_) );
  OR2_X1 g0202 ( .A1(new_n560_), .A2(new_n559_), .ZN(new_n561_) );
  AND2_X1 g0203 ( .A1(new_n561_), .A2(new_n558_), .ZN(new_n562_) );
  OR2_X1 g0204 ( .A1(new_n562_), .A2(KEYINPUT13), .ZN(new_n563_) );
  AND2_X1 g0205 ( .A1(new_n555_), .A2(new_n563_), .ZN(new_n564_) );
  AND2_X1 g0206 ( .A1(new_n564_), .A2(new_n543_), .ZN(new_n565_) );
  INV_X1 g0207 ( .A(new_n565_), .ZN(new_n566_) );
  OR2_X1 g0208 ( .A1(new_n566_), .A2(new_n534_), .ZN(G153) );
  INV_X1 g0209 ( .A(G36), .ZN(new_n568_) );
  INV_X1 g0210 ( .A(G319), .ZN(new_n569_) );
  AND2_X1 g0211 ( .A1(G483), .A2(G661), .ZN(new_n570_) );
  INV_X1 g0212 ( .A(new_n570_), .ZN(new_n571_) );
  OR2_X1 g0213 ( .A1(new_n569_), .A2(new_n571_), .ZN(new_n572_) );
  OR2_X1 g0214 ( .A1(new_n572_), .A2(new_n568_), .ZN(G176) );
  AND2_X1 g0215 ( .A1(G1), .A2(G3), .ZN(new_n574_) );
  OR2_X1 g0216 ( .A1(new_n572_), .A2(new_n574_), .ZN(G188) );
  AND2_X1 g0217 ( .A1(new_n473_), .A2(G53), .ZN(new_n576_) );
  AND2_X1 g0218 ( .A1(new_n477_), .A2(G91), .ZN(new_n577_) );
  OR2_X1 g0219 ( .A1(new_n576_), .A2(new_n577_), .ZN(new_n578_) );
  AND2_X1 g0220 ( .A1(new_n483_), .A2(G78), .ZN(new_n579_) );
  AND2_X1 g0221 ( .A1(new_n490_), .A2(G65), .ZN(new_n580_) );
  OR2_X1 g0222 ( .A1(new_n580_), .A2(new_n579_), .ZN(new_n581_) );
  OR2_X1 g0223 ( .A1(new_n578_), .A2(new_n581_), .ZN(G299) );
  INV_X1 g0224 ( .A(G171), .ZN(G301) );
  INV_X1 g0225 ( .A(G168), .ZN(new_n584_) );
  AND2_X1 g0226 ( .A1(new_n584_), .A2(KEYINPUT8), .ZN(new_n585_) );
  INV_X1 g0227 ( .A(new_n585_), .ZN(new_n586_) );
  OR2_X1 g0228 ( .A1(new_n584_), .A2(KEYINPUT8), .ZN(new_n587_) );
  AND2_X1 g0229 ( .A1(new_n586_), .A2(new_n587_), .ZN(new_n588_) );
  INV_X1 g0230 ( .A(new_n588_), .ZN(G286) );
  AND2_X1 g0231 ( .A1(new_n473_), .A2(G49), .ZN(new_n590_) );
  AND2_X1 g0232 ( .A1(new_n471_), .A2(G87), .ZN(new_n591_) );
  AND2_X1 g0233 ( .A1(G74), .A2(G651), .ZN(new_n592_) );
  OR2_X1 g0234 ( .A1(new_n490_), .A2(new_n592_), .ZN(new_n593_) );
  OR2_X1 g0235 ( .A1(new_n593_), .A2(new_n591_), .ZN(new_n594_) );
  OR2_X1 g0236 ( .A1(new_n594_), .A2(new_n590_), .ZN(G288) );
  AND2_X1 g0237 ( .A1(new_n483_), .A2(G73), .ZN(new_n596_) );
  INV_X1 g0238 ( .A(new_n596_), .ZN(new_n597_) );
  AND2_X1 g0239 ( .A1(new_n597_), .A2(KEYINPUT2), .ZN(new_n598_) );
  INV_X1 g0240 ( .A(new_n598_), .ZN(new_n599_) );
  OR2_X1 g0241 ( .A1(new_n597_), .A2(KEYINPUT2), .ZN(new_n600_) );
  AND2_X1 g0242 ( .A1(new_n599_), .A2(new_n600_), .ZN(new_n601_) );
  AND2_X1 g0243 ( .A1(new_n490_), .A2(G61), .ZN(new_n602_) );
  AND2_X1 g0244 ( .A1(new_n473_), .A2(G48), .ZN(new_n603_) );
  AND2_X1 g0245 ( .A1(new_n477_), .A2(G86), .ZN(new_n604_) );
  OR2_X1 g0246 ( .A1(new_n603_), .A2(new_n604_), .ZN(new_n605_) );
  OR2_X1 g0247 ( .A1(new_n605_), .A2(new_n602_), .ZN(new_n606_) );
  OR2_X1 g0248 ( .A1(new_n601_), .A2(new_n606_), .ZN(G305) );
  AND2_X1 g0249 ( .A1(new_n473_), .A2(G47), .ZN(new_n608_) );
  AND2_X1 g0250 ( .A1(new_n477_), .A2(G85), .ZN(new_n609_) );
  OR2_X1 g0251 ( .A1(new_n608_), .A2(new_n609_), .ZN(new_n610_) );
  AND2_X1 g0252 ( .A1(new_n483_), .A2(G72), .ZN(new_n611_) );
  AND2_X1 g0253 ( .A1(new_n490_), .A2(G60), .ZN(new_n612_) );
  OR2_X1 g0254 ( .A1(new_n612_), .A2(new_n611_), .ZN(new_n613_) );
  OR2_X1 g0255 ( .A1(new_n610_), .A2(new_n613_), .ZN(G290) );
  INV_X1 g0256 ( .A(G868), .ZN(new_n615_) );
  INV_X1 g0257 ( .A(KEYINPUT15), .ZN(new_n616_) );
  AND2_X1 g0258 ( .A1(new_n473_), .A2(G54), .ZN(new_n617_) );
  AND2_X1 g0259 ( .A1(new_n477_), .A2(G92), .ZN(new_n618_) );
  OR2_X1 g0260 ( .A1(new_n617_), .A2(new_n618_), .ZN(new_n619_) );
  AND2_X1 g0261 ( .A1(new_n483_), .A2(G79), .ZN(new_n620_) );
  AND2_X1 g0262 ( .A1(new_n490_), .A2(G66), .ZN(new_n621_) );
  OR2_X1 g0263 ( .A1(new_n621_), .A2(new_n620_), .ZN(new_n622_) );
  OR2_X1 g0264 ( .A1(new_n619_), .A2(new_n622_), .ZN(new_n623_) );
  AND2_X1 g0265 ( .A1(new_n623_), .A2(new_n616_), .ZN(new_n624_) );
  INV_X1 g0266 ( .A(new_n624_), .ZN(new_n625_) );
  OR2_X1 g0267 ( .A1(new_n623_), .A2(new_n616_), .ZN(new_n626_) );
  AND2_X1 g0268 ( .A1(new_n625_), .A2(new_n626_), .ZN(new_n627_) );
  INV_X1 g0269 ( .A(new_n627_), .ZN(new_n628_) );
  AND2_X1 g0270 ( .A1(new_n628_), .A2(new_n615_), .ZN(new_n629_) );
  AND2_X1 g0271 ( .A1(G301), .A2(G868), .ZN(new_n630_) );
  OR2_X1 g0272 ( .A1(new_n629_), .A2(new_n630_), .ZN(G284) );
  OR2_X1 g0273 ( .A1(G286), .A2(new_n615_), .ZN(new_n632_) );
  OR2_X1 g0274 ( .A1(G299), .A2(G868), .ZN(new_n633_) );
  AND2_X1 g0275 ( .A1(new_n632_), .A2(new_n633_), .ZN(G297) );
  INV_X1 g0276 ( .A(KEYINPUT16), .ZN(new_n635_) );
  AND2_X1 g0277 ( .A1(new_n534_), .A2(G559), .ZN(new_n636_) );
  OR2_X1 g0278 ( .A1(new_n628_), .A2(new_n636_), .ZN(new_n637_) );
  INV_X1 g0279 ( .A(new_n637_), .ZN(new_n638_) );
  AND2_X1 g0280 ( .A1(new_n638_), .A2(new_n635_), .ZN(new_n639_) );
  AND2_X1 g0281 ( .A1(new_n637_), .A2(KEYINPUT16), .ZN(new_n640_) );
  OR2_X1 g0282 ( .A1(new_n639_), .A2(new_n640_), .ZN(G148) );
  OR2_X1 g0283 ( .A1(new_n615_), .A2(G559), .ZN(new_n642_) );
  OR2_X1 g0284 ( .A1(new_n628_), .A2(new_n642_), .ZN(new_n643_) );
  OR2_X1 g0285 ( .A1(new_n566_), .A2(G868), .ZN(new_n644_) );
  AND2_X1 g0286 ( .A1(new_n643_), .A2(new_n644_), .ZN(G282) );
  INV_X1 g0287 ( .A(G2096), .ZN(new_n646_) );
  AND2_X1 g0288 ( .A1(new_n438_), .A2(G123), .ZN(new_n647_) );
  INV_X1 g0289 ( .A(new_n647_), .ZN(new_n648_) );
  AND2_X1 g0290 ( .A1(new_n648_), .A2(KEYINPUT18), .ZN(new_n649_) );
  INV_X1 g0291 ( .A(new_n649_), .ZN(new_n650_) );
  OR2_X1 g0292 ( .A1(new_n648_), .A2(KEYINPUT18), .ZN(new_n651_) );
  AND2_X1 g0293 ( .A1(new_n650_), .A2(new_n651_), .ZN(new_n652_) );
  AND2_X1 g0294 ( .A1(new_n451_), .A2(G135), .ZN(new_n653_) );
  AND2_X1 g0295 ( .A1(new_n453_), .A2(G99), .ZN(new_n654_) );
  AND2_X1 g0296 ( .A1(new_n436_), .A2(G111), .ZN(new_n655_) );
  OR2_X1 g0297 ( .A1(new_n654_), .A2(new_n655_), .ZN(new_n656_) );
  OR2_X1 g0298 ( .A1(new_n653_), .A2(new_n656_), .ZN(new_n657_) );
  OR2_X1 g0299 ( .A1(new_n657_), .A2(new_n652_), .ZN(new_n658_) );
  INV_X1 g0300 ( .A(new_n658_), .ZN(new_n659_) );
  AND2_X1 g0301 ( .A1(new_n659_), .A2(new_n646_), .ZN(new_n660_) );
  AND2_X1 g0302 ( .A1(new_n658_), .A2(G2096), .ZN(new_n661_) );
  OR2_X1 g0303 ( .A1(new_n661_), .A2(G2100), .ZN(new_n662_) );
  OR2_X1 g0304 ( .A1(new_n662_), .A2(new_n660_), .ZN(G156) );
  INV_X1 g0305 ( .A(G2454), .ZN(new_n664_) );
  AND2_X1 g0306 ( .A1(new_n664_), .A2(G2430), .ZN(new_n665_) );
  INV_X1 g0307 ( .A(new_n665_), .ZN(new_n666_) );
  OR2_X1 g0308 ( .A1(new_n664_), .A2(G2430), .ZN(new_n667_) );
  AND2_X1 g0309 ( .A1(new_n666_), .A2(new_n667_), .ZN(new_n668_) );
  INV_X1 g0310 ( .A(new_n668_), .ZN(new_n669_) );
  INV_X1 g0311 ( .A(G1341), .ZN(new_n670_) );
  INV_X1 g0312 ( .A(G1348), .ZN(new_n671_) );
  AND2_X1 g0313 ( .A1(new_n670_), .A2(new_n671_), .ZN(new_n672_) );
  AND2_X1 g0314 ( .A1(G1341), .A2(G1348), .ZN(new_n673_) );
  OR2_X1 g0315 ( .A1(new_n672_), .A2(new_n673_), .ZN(new_n674_) );
  AND2_X1 g0316 ( .A1(new_n669_), .A2(new_n674_), .ZN(new_n675_) );
  INV_X1 g0317 ( .A(new_n675_), .ZN(new_n676_) );
  OR2_X1 g0318 ( .A1(new_n669_), .A2(new_n674_), .ZN(new_n677_) );
  AND2_X1 g0319 ( .A1(new_n676_), .A2(new_n677_), .ZN(new_n678_) );
  INV_X1 g0320 ( .A(new_n678_), .ZN(new_n679_) );
  AND2_X1 g0321 ( .A1(G2435), .A2(G2438), .ZN(new_n680_) );
  INV_X1 g0322 ( .A(new_n680_), .ZN(new_n681_) );
  OR2_X1 g0323 ( .A1(G2435), .A2(G2438), .ZN(new_n682_) );
  AND2_X1 g0324 ( .A1(new_n681_), .A2(new_n682_), .ZN(new_n683_) );
  INV_X1 g0325 ( .A(new_n683_), .ZN(new_n684_) );
  AND2_X1 g0326 ( .A1(new_n679_), .A2(new_n684_), .ZN(new_n685_) );
  AND2_X1 g0327 ( .A1(new_n678_), .A2(new_n683_), .ZN(new_n686_) );
  OR2_X1 g0328 ( .A1(new_n685_), .A2(new_n686_), .ZN(new_n687_) );
  INV_X1 g0329 ( .A(G2451), .ZN(new_n688_) );
  AND2_X1 g0330 ( .A1(new_n688_), .A2(G2446), .ZN(new_n689_) );
  INV_X1 g0331 ( .A(new_n689_), .ZN(new_n690_) );
  OR2_X1 g0332 ( .A1(new_n688_), .A2(G2446), .ZN(new_n691_) );
  AND2_X1 g0333 ( .A1(new_n690_), .A2(new_n691_), .ZN(new_n692_) );
  INV_X1 g0334 ( .A(new_n692_), .ZN(new_n693_) );
  AND2_X1 g0335 ( .A1(G2427), .A2(G2443), .ZN(new_n694_) );
  INV_X1 g0336 ( .A(new_n694_), .ZN(new_n695_) );
  OR2_X1 g0337 ( .A1(G2427), .A2(G2443), .ZN(new_n696_) );
  AND2_X1 g0338 ( .A1(new_n695_), .A2(new_n696_), .ZN(new_n697_) );
  INV_X1 g0339 ( .A(new_n697_), .ZN(new_n698_) );
  AND2_X1 g0340 ( .A1(new_n693_), .A2(new_n698_), .ZN(new_n699_) );
  AND2_X1 g0341 ( .A1(new_n692_), .A2(new_n697_), .ZN(new_n700_) );
  OR2_X1 g0342 ( .A1(new_n699_), .A2(new_n700_), .ZN(new_n701_) );
  AND2_X1 g0343 ( .A1(new_n687_), .A2(new_n701_), .ZN(new_n702_) );
  INV_X1 g0344 ( .A(new_n702_), .ZN(new_n703_) );
  OR2_X1 g0345 ( .A1(new_n687_), .A2(new_n701_), .ZN(new_n704_) );
  AND2_X1 g0346 ( .A1(new_n703_), .A2(new_n704_), .ZN(new_n705_) );
  INV_X1 g0347 ( .A(new_n705_), .ZN(new_n706_) );
  AND2_X1 g0348 ( .A1(new_n706_), .A2(G14), .ZN(G401) );
  INV_X1 g0349 ( .A(KEYINPUT42), .ZN(new_n708_) );
  AND2_X1 g0350 ( .A1(new_n708_), .A2(G2090), .ZN(new_n709_) );
  INV_X1 g0351 ( .A(G2090), .ZN(new_n710_) );
  AND2_X1 g0352 ( .A1(new_n710_), .A2(KEYINPUT42), .ZN(new_n711_) );
  OR2_X1 g0353 ( .A1(new_n709_), .A2(new_n711_), .ZN(new_n712_) );
  INV_X1 g0354 ( .A(G2067), .ZN(new_n713_) );
  AND2_X1 g0355 ( .A1(new_n713_), .A2(new_n371_), .ZN(new_n714_) );
  AND2_X1 g0356 ( .A1(G2067), .A2(G2072), .ZN(new_n715_) );
  OR2_X1 g0357 ( .A1(new_n714_), .A2(new_n715_), .ZN(new_n716_) );
  AND2_X1 g0358 ( .A1(new_n712_), .A2(new_n716_), .ZN(new_n717_) );
  INV_X1 g0359 ( .A(new_n717_), .ZN(new_n718_) );
  OR2_X1 g0360 ( .A1(new_n712_), .A2(new_n716_), .ZN(new_n719_) );
  AND2_X1 g0361 ( .A1(new_n718_), .A2(new_n719_), .ZN(new_n720_) );
  INV_X1 g0362 ( .A(new_n720_), .ZN(new_n721_) );
  AND2_X1 g0363 ( .A1(G2096), .A2(G2100), .ZN(new_n722_) );
  INV_X1 g0364 ( .A(new_n722_), .ZN(new_n723_) );
  OR2_X1 g0365 ( .A1(G2096), .A2(G2100), .ZN(new_n724_) );
  AND2_X1 g0366 ( .A1(new_n723_), .A2(new_n724_), .ZN(new_n725_) );
  INV_X1 g0367 ( .A(new_n725_), .ZN(new_n726_) );
  AND2_X1 g0368 ( .A1(G2678), .A2(KEYINPUT43), .ZN(new_n727_) );
  INV_X1 g0369 ( .A(new_n727_), .ZN(new_n728_) );
  OR2_X1 g0370 ( .A1(G2678), .A2(KEYINPUT43), .ZN(new_n729_) );
  AND2_X1 g0371 ( .A1(new_n728_), .A2(new_n729_), .ZN(new_n730_) );
  INV_X1 g0372 ( .A(new_n730_), .ZN(new_n731_) );
  AND2_X1 g0373 ( .A1(new_n726_), .A2(new_n731_), .ZN(new_n732_) );
  AND2_X1 g0374 ( .A1(new_n725_), .A2(new_n730_), .ZN(new_n733_) );
  OR2_X1 g0375 ( .A1(new_n732_), .A2(new_n733_), .ZN(new_n734_) );
  AND2_X1 g0376 ( .A1(new_n721_), .A2(new_n734_), .ZN(new_n735_) );
  INV_X1 g0377 ( .A(new_n735_), .ZN(new_n736_) );
  OR2_X1 g0378 ( .A1(new_n721_), .A2(new_n734_), .ZN(new_n737_) );
  AND2_X1 g0379 ( .A1(new_n736_), .A2(new_n737_), .ZN(new_n738_) );
  INV_X1 g0380 ( .A(new_n738_), .ZN(new_n739_) );
  INV_X1 g0381 ( .A(G2078), .ZN(new_n740_) );
  INV_X1 g0382 ( .A(G2084), .ZN(new_n741_) );
  AND2_X1 g0383 ( .A1(new_n740_), .A2(new_n741_), .ZN(new_n742_) );
  OR2_X1 g0384 ( .A1(new_n742_), .A2(new_n374_), .ZN(new_n743_) );
  AND2_X1 g0385 ( .A1(new_n739_), .A2(new_n743_), .ZN(new_n744_) );
  INV_X1 g0386 ( .A(new_n744_), .ZN(new_n745_) );
  OR2_X1 g0387 ( .A1(new_n739_), .A2(new_n743_), .ZN(new_n746_) );
  AND2_X1 g0388 ( .A1(new_n745_), .A2(new_n746_), .ZN(new_n747_) );
  INV_X1 g0389 ( .A(new_n747_), .ZN(G227) );
  INV_X1 g0390 ( .A(G1981), .ZN(new_n749_) );
  AND2_X1 g0391 ( .A1(new_n749_), .A2(G1976), .ZN(new_n750_) );
  INV_X1 g0392 ( .A(G1976), .ZN(new_n751_) );
  AND2_X1 g0393 ( .A1(new_n751_), .A2(G1981), .ZN(new_n752_) );
  OR2_X1 g0394 ( .A1(new_n750_), .A2(new_n752_), .ZN(new_n753_) );
  INV_X1 g0395 ( .A(G1956), .ZN(new_n754_) );
  INV_X1 g0396 ( .A(G1966), .ZN(new_n755_) );
  AND2_X1 g0397 ( .A1(new_n754_), .A2(new_n755_), .ZN(new_n756_) );
  AND2_X1 g0398 ( .A1(G1956), .A2(G1966), .ZN(new_n757_) );
  OR2_X1 g0399 ( .A1(new_n756_), .A2(new_n757_), .ZN(new_n758_) );
  AND2_X1 g0400 ( .A1(new_n753_), .A2(new_n758_), .ZN(new_n759_) );
  INV_X1 g0401 ( .A(new_n759_), .ZN(new_n760_) );
  OR2_X1 g0402 ( .A1(new_n753_), .A2(new_n758_), .ZN(new_n761_) );
  AND2_X1 g0403 ( .A1(new_n760_), .A2(new_n761_), .ZN(new_n762_) );
  INV_X1 g0404 ( .A(new_n762_), .ZN(new_n763_) );
  AND2_X1 g0405 ( .A1(new_n763_), .A2(G2474), .ZN(new_n764_) );
  INV_X1 g0406 ( .A(new_n764_), .ZN(new_n765_) );
  OR2_X1 g0407 ( .A1(new_n763_), .A2(G2474), .ZN(new_n766_) );
  AND2_X1 g0408 ( .A1(new_n765_), .A2(new_n766_), .ZN(new_n767_) );
  INV_X1 g0409 ( .A(new_n767_), .ZN(new_n768_) );
  INV_X1 g0410 ( .A(G1996), .ZN(new_n769_) );
  AND2_X1 g0411 ( .A1(new_n769_), .A2(G1991), .ZN(new_n770_) );
  INV_X1 g0412 ( .A(G1991), .ZN(new_n771_) );
  AND2_X1 g0413 ( .A1(new_n771_), .A2(G1996), .ZN(new_n772_) );
  OR2_X1 g0414 ( .A1(new_n770_), .A2(new_n772_), .ZN(new_n773_) );
  AND2_X1 g0415 ( .A1(new_n768_), .A2(new_n773_), .ZN(new_n774_) );
  INV_X1 g0416 ( .A(new_n774_), .ZN(new_n775_) );
  OR2_X1 g0417 ( .A1(new_n768_), .A2(new_n773_), .ZN(new_n776_) );
  AND2_X1 g0418 ( .A1(new_n775_), .A2(new_n776_), .ZN(new_n777_) );
  INV_X1 g0419 ( .A(new_n777_), .ZN(new_n778_) );
  INV_X1 g0420 ( .A(KEYINPUT41), .ZN(new_n779_) );
  AND2_X1 g0421 ( .A1(new_n779_), .A2(G1971), .ZN(new_n780_) );
  INV_X1 g0422 ( .A(G1971), .ZN(new_n781_) );
  AND2_X1 g0423 ( .A1(new_n781_), .A2(KEYINPUT41), .ZN(new_n782_) );
  OR2_X1 g0424 ( .A1(new_n780_), .A2(new_n782_), .ZN(new_n783_) );
  INV_X1 g0425 ( .A(G1961), .ZN(new_n784_) );
  INV_X1 g0426 ( .A(G1986), .ZN(new_n785_) );
  AND2_X1 g0427 ( .A1(new_n784_), .A2(new_n785_), .ZN(new_n786_) );
  AND2_X1 g0428 ( .A1(G1961), .A2(G1986), .ZN(new_n787_) );
  OR2_X1 g0429 ( .A1(new_n786_), .A2(new_n787_), .ZN(new_n788_) );
  AND2_X1 g0430 ( .A1(new_n783_), .A2(new_n788_), .ZN(new_n789_) );
  INV_X1 g0431 ( .A(new_n789_), .ZN(new_n790_) );
  OR2_X1 g0432 ( .A1(new_n783_), .A2(new_n788_), .ZN(new_n791_) );
  AND2_X1 g0433 ( .A1(new_n790_), .A2(new_n791_), .ZN(new_n792_) );
  INV_X1 g0434 ( .A(new_n792_), .ZN(new_n793_) );
  AND2_X1 g0435 ( .A1(new_n778_), .A2(new_n793_), .ZN(new_n794_) );
  AND2_X1 g0436 ( .A1(new_n777_), .A2(new_n792_), .ZN(new_n795_) );
  OR2_X1 g0437 ( .A1(new_n794_), .A2(new_n795_), .ZN(G229) );
  INV_X1 g0438 ( .A(G29), .ZN(new_n797_) );
  INV_X1 g0439 ( .A(KEYINPUT52), .ZN(new_n798_) );
  INV_X1 g0440 ( .A(KEYINPUT50), .ZN(new_n799_) );
  INV_X1 g0441 ( .A(KEYINPUT47), .ZN(new_n800_) );
  AND2_X1 g0442 ( .A1(new_n438_), .A2(G127), .ZN(new_n801_) );
  AND2_X1 g0443 ( .A1(new_n436_), .A2(G115), .ZN(new_n802_) );
  OR2_X1 g0444 ( .A1(new_n801_), .A2(new_n802_), .ZN(new_n803_) );
  AND2_X1 g0445 ( .A1(new_n803_), .A2(new_n800_), .ZN(new_n804_) );
  AND2_X1 g0446 ( .A1(new_n453_), .A2(G103), .ZN(new_n805_) );
  OR2_X1 g0447 ( .A1(new_n804_), .A2(new_n805_), .ZN(new_n806_) );
  INV_X1 g0448 ( .A(new_n806_), .ZN(new_n807_) );
  AND2_X1 g0449 ( .A1(new_n451_), .A2(G139), .ZN(new_n808_) );
  INV_X1 g0450 ( .A(new_n808_), .ZN(new_n809_) );
  OR2_X1 g0451 ( .A1(new_n803_), .A2(new_n800_), .ZN(new_n810_) );
  AND2_X1 g0452 ( .A1(new_n809_), .A2(new_n810_), .ZN(new_n811_) );
  AND2_X1 g0453 ( .A1(new_n807_), .A2(new_n811_), .ZN(new_n812_) );
  AND2_X1 g0454 ( .A1(new_n812_), .A2(new_n371_), .ZN(new_n813_) );
  INV_X1 g0455 ( .A(new_n812_), .ZN(new_n814_) );
  AND2_X1 g0456 ( .A1(new_n814_), .A2(G2072), .ZN(new_n815_) );
  AND2_X1 g0457 ( .A1(G164), .A2(new_n740_), .ZN(new_n816_) );
  AND2_X1 g0458 ( .A1(new_n466_), .A2(G2078), .ZN(new_n817_) );
  OR2_X1 g0459 ( .A1(new_n816_), .A2(new_n817_), .ZN(new_n818_) );
  OR2_X1 g0460 ( .A1(new_n815_), .A2(new_n818_), .ZN(new_n819_) );
  OR2_X1 g0461 ( .A1(new_n819_), .A2(new_n813_), .ZN(new_n820_) );
  INV_X1 g0462 ( .A(new_n820_), .ZN(new_n821_) );
  AND2_X1 g0463 ( .A1(new_n821_), .A2(new_n799_), .ZN(new_n822_) );
  AND2_X1 g0464 ( .A1(new_n820_), .A2(KEYINPUT50), .ZN(new_n823_) );
  INV_X1 g0465 ( .A(KEYINPUT51), .ZN(new_n824_) );
  AND2_X1 g0466 ( .A1(new_n451_), .A2(G141), .ZN(new_n825_) );
  INV_X1 g0467 ( .A(KEYINPUT38), .ZN(new_n826_) );
  AND2_X1 g0468 ( .A1(new_n453_), .A2(G105), .ZN(new_n827_) );
  INV_X1 g0469 ( .A(new_n827_), .ZN(new_n828_) );
  AND2_X1 g0470 ( .A1(new_n828_), .A2(new_n826_), .ZN(new_n829_) );
  AND2_X1 g0471 ( .A1(new_n827_), .A2(KEYINPUT38), .ZN(new_n830_) );
  AND2_X1 g0472 ( .A1(new_n438_), .A2(G129), .ZN(new_n831_) );
  AND2_X1 g0473 ( .A1(new_n436_), .A2(G117), .ZN(new_n832_) );
  OR2_X1 g0474 ( .A1(new_n831_), .A2(new_n832_), .ZN(new_n833_) );
  OR2_X1 g0475 ( .A1(new_n833_), .A2(new_n830_), .ZN(new_n834_) );
  OR2_X1 g0476 ( .A1(new_n834_), .A2(new_n829_), .ZN(new_n835_) );
  OR2_X1 g0477 ( .A1(new_n835_), .A2(new_n825_), .ZN(new_n836_) );
  INV_X1 g0478 ( .A(new_n836_), .ZN(new_n837_) );
  AND2_X1 g0479 ( .A1(new_n837_), .A2(new_n769_), .ZN(new_n838_) );
  AND2_X1 g0480 ( .A1(G162), .A2(new_n710_), .ZN(new_n839_) );
  AND2_X1 g0481 ( .A1(new_n458_), .A2(G2090), .ZN(new_n840_) );
  OR2_X1 g0482 ( .A1(new_n839_), .A2(new_n840_), .ZN(new_n841_) );
  OR2_X1 g0483 ( .A1(new_n841_), .A2(new_n838_), .ZN(new_n842_) );
  AND2_X1 g0484 ( .A1(new_n842_), .A2(new_n824_), .ZN(new_n843_) );
  OR2_X1 g0485 ( .A1(new_n823_), .A2(new_n843_), .ZN(new_n844_) );
  OR2_X1 g0486 ( .A1(new_n844_), .A2(new_n822_), .ZN(new_n845_) );
  INV_X1 g0487 ( .A(new_n845_), .ZN(new_n846_) );
  INV_X1 g0488 ( .A(KEYINPUT34), .ZN(new_n847_) );
  AND2_X1 g0489 ( .A1(new_n451_), .A2(G140), .ZN(new_n848_) );
  AND2_X1 g0490 ( .A1(new_n453_), .A2(G104), .ZN(new_n849_) );
  OR2_X1 g0491 ( .A1(new_n848_), .A2(new_n849_), .ZN(new_n850_) );
  INV_X1 g0492 ( .A(new_n850_), .ZN(new_n851_) );
  AND2_X1 g0493 ( .A1(new_n851_), .A2(new_n847_), .ZN(new_n852_) );
  AND2_X1 g0494 ( .A1(new_n850_), .A2(KEYINPUT34), .ZN(new_n853_) );
  AND2_X1 g0495 ( .A1(new_n438_), .A2(G128), .ZN(new_n854_) );
  AND2_X1 g0496 ( .A1(new_n436_), .A2(G116), .ZN(new_n855_) );
  OR2_X1 g0497 ( .A1(new_n854_), .A2(new_n855_), .ZN(new_n856_) );
  AND2_X1 g0498 ( .A1(new_n856_), .A2(KEYINPUT35), .ZN(new_n857_) );
  INV_X1 g0499 ( .A(new_n857_), .ZN(new_n858_) );
  OR2_X1 g0500 ( .A1(new_n856_), .A2(KEYINPUT35), .ZN(new_n859_) );
  AND2_X1 g0501 ( .A1(new_n858_), .A2(new_n859_), .ZN(new_n860_) );
  OR2_X1 g0502 ( .A1(new_n853_), .A2(new_n860_), .ZN(new_n861_) );
  OR2_X1 g0503 ( .A1(new_n861_), .A2(new_n852_), .ZN(new_n862_) );
  AND2_X1 g0504 ( .A1(new_n862_), .A2(KEYINPUT36), .ZN(new_n863_) );
  INV_X1 g0505 ( .A(new_n863_), .ZN(new_n864_) );
  OR2_X1 g0506 ( .A1(new_n862_), .A2(KEYINPUT36), .ZN(new_n865_) );
  AND2_X1 g0507 ( .A1(new_n864_), .A2(new_n865_), .ZN(new_n866_) );
  INV_X1 g0508 ( .A(new_n866_), .ZN(new_n867_) );
  AND2_X1 g0509 ( .A1(new_n713_), .A2(KEYINPUT37), .ZN(new_n868_) );
  INV_X1 g0510 ( .A(new_n868_), .ZN(new_n869_) );
  OR2_X1 g0511 ( .A1(new_n713_), .A2(KEYINPUT37), .ZN(new_n870_) );
  AND2_X1 g0512 ( .A1(new_n869_), .A2(new_n870_), .ZN(new_n871_) );
  INV_X1 g0513 ( .A(new_n871_), .ZN(new_n872_) );
  AND2_X1 g0514 ( .A1(new_n867_), .A2(new_n872_), .ZN(new_n873_) );
  INV_X1 g0515 ( .A(new_n873_), .ZN(new_n874_) );
  AND2_X1 g0516 ( .A1(new_n866_), .A2(new_n871_), .ZN(new_n875_) );
  INV_X1 g0517 ( .A(new_n875_), .ZN(new_n876_) );
  OR2_X1 g0518 ( .A1(new_n842_), .A2(new_n824_), .ZN(new_n877_) );
  INV_X1 g0519 ( .A(G160), .ZN(new_n878_) );
  AND2_X1 g0520 ( .A1(new_n878_), .A2(new_n741_), .ZN(new_n879_) );
  AND2_X1 g0521 ( .A1(G160), .A2(G2084), .ZN(new_n880_) );
  OR2_X1 g0522 ( .A1(new_n879_), .A2(new_n880_), .ZN(new_n881_) );
  AND2_X1 g0523 ( .A1(new_n836_), .A2(G1996), .ZN(new_n882_) );
  AND2_X1 g0524 ( .A1(new_n451_), .A2(G131), .ZN(new_n883_) );
  AND2_X1 g0525 ( .A1(new_n438_), .A2(G119), .ZN(new_n884_) );
  AND2_X1 g0526 ( .A1(new_n453_), .A2(G95), .ZN(new_n885_) );
  AND2_X1 g0527 ( .A1(new_n436_), .A2(G107), .ZN(new_n886_) );
  OR2_X1 g0528 ( .A1(new_n885_), .A2(new_n886_), .ZN(new_n887_) );
  OR2_X1 g0529 ( .A1(new_n887_), .A2(new_n884_), .ZN(new_n888_) );
  OR2_X1 g0530 ( .A1(new_n888_), .A2(new_n883_), .ZN(new_n889_) );
  AND2_X1 g0531 ( .A1(new_n889_), .A2(G1991), .ZN(new_n890_) );
  OR2_X1 g0532 ( .A1(new_n882_), .A2(new_n890_), .ZN(new_n891_) );
  INV_X1 g0533 ( .A(new_n891_), .ZN(new_n892_) );
  INV_X1 g0534 ( .A(new_n889_), .ZN(new_n893_) );
  AND2_X1 g0535 ( .A1(new_n893_), .A2(new_n771_), .ZN(new_n894_) );
  INV_X1 g0536 ( .A(new_n894_), .ZN(new_n895_) );
  AND2_X1 g0537 ( .A1(new_n895_), .A2(new_n658_), .ZN(new_n896_) );
  AND2_X1 g0538 ( .A1(new_n892_), .A2(new_n896_), .ZN(new_n897_) );
  AND2_X1 g0539 ( .A1(new_n897_), .A2(new_n881_), .ZN(new_n898_) );
  AND2_X1 g0540 ( .A1(new_n877_), .A2(new_n898_), .ZN(new_n899_) );
  AND2_X1 g0541 ( .A1(new_n876_), .A2(new_n899_), .ZN(new_n900_) );
  AND2_X1 g0542 ( .A1(new_n900_), .A2(new_n874_), .ZN(new_n901_) );
  AND2_X1 g0543 ( .A1(new_n901_), .A2(new_n846_), .ZN(new_n902_) );
  OR2_X1 g0544 ( .A1(new_n902_), .A2(new_n798_), .ZN(new_n903_) );
  AND2_X1 g0545 ( .A1(new_n902_), .A2(new_n798_), .ZN(new_n904_) );
  OR2_X1 g0546 ( .A1(new_n904_), .A2(KEYINPUT55), .ZN(new_n905_) );
  INV_X1 g0547 ( .A(new_n905_), .ZN(new_n906_) );
  AND2_X1 g0548 ( .A1(new_n906_), .A2(new_n903_), .ZN(new_n907_) );
  OR2_X1 g0549 ( .A1(new_n907_), .A2(new_n797_), .ZN(new_n908_) );
  AND2_X1 g0550 ( .A1(new_n584_), .A2(new_n755_), .ZN(new_n909_) );
  AND2_X1 g0551 ( .A1(G168), .A2(G1966), .ZN(new_n910_) );
  OR2_X1 g0552 ( .A1(new_n909_), .A2(new_n910_), .ZN(new_n911_) );
  INV_X1 g0553 ( .A(G305), .ZN(new_n912_) );
  AND2_X1 g0554 ( .A1(new_n912_), .A2(new_n749_), .ZN(new_n913_) );
  AND2_X1 g0555 ( .A1(G305), .A2(G1981), .ZN(new_n914_) );
  OR2_X1 g0556 ( .A1(new_n913_), .A2(new_n914_), .ZN(new_n915_) );
  INV_X1 g0557 ( .A(new_n915_), .ZN(new_n916_) );
  AND2_X1 g0558 ( .A1(new_n911_), .A2(new_n916_), .ZN(new_n917_) );
  INV_X1 g0559 ( .A(new_n917_), .ZN(new_n918_) );
  AND2_X1 g0560 ( .A1(new_n918_), .A2(KEYINPUT57), .ZN(new_n919_) );
  INV_X1 g0561 ( .A(new_n919_), .ZN(new_n920_) );
  OR2_X1 g0562 ( .A1(new_n918_), .A2(KEYINPUT57), .ZN(new_n921_) );
  AND2_X1 g0563 ( .A1(new_n920_), .A2(new_n921_), .ZN(new_n922_) );
  INV_X1 g0564 ( .A(new_n922_), .ZN(new_n923_) );
  AND2_X1 g0565 ( .A1(G301), .A2(new_n784_), .ZN(new_n924_) );
  AND2_X1 g0566 ( .A1(G171), .A2(G1961), .ZN(new_n925_) );
  OR2_X1 g0567 ( .A1(new_n924_), .A2(new_n925_), .ZN(new_n926_) );
  AND2_X1 g0568 ( .A1(G166), .A2(new_n781_), .ZN(new_n927_) );
  INV_X1 g0569 ( .A(G288), .ZN(new_n928_) );
  AND2_X1 g0570 ( .A1(new_n928_), .A2(new_n751_), .ZN(new_n929_) );
  OR2_X1 g0571 ( .A1(new_n927_), .A2(new_n929_), .ZN(new_n930_) );
  AND2_X1 g0572 ( .A1(G303), .A2(G1971), .ZN(new_n931_) );
  AND2_X1 g0573 ( .A1(G288), .A2(G1976), .ZN(new_n932_) );
  OR2_X1 g0574 ( .A1(new_n931_), .A2(new_n932_), .ZN(new_n933_) );
  OR2_X1 g0575 ( .A1(new_n930_), .A2(new_n933_), .ZN(new_n934_) );
  INV_X1 g0576 ( .A(new_n934_), .ZN(new_n935_) );
  INV_X1 g0577 ( .A(G290), .ZN(new_n936_) );
  AND2_X1 g0578 ( .A1(new_n936_), .A2(new_n785_), .ZN(new_n937_) );
  AND2_X1 g0579 ( .A1(G290), .A2(G1986), .ZN(new_n938_) );
  OR2_X1 g0580 ( .A1(new_n937_), .A2(new_n938_), .ZN(new_n939_) );
  INV_X1 g0581 ( .A(new_n939_), .ZN(new_n940_) );
  INV_X1 g0582 ( .A(G299), .ZN(new_n941_) );
  AND2_X1 g0583 ( .A1(new_n941_), .A2(G1956), .ZN(new_n942_) );
  AND2_X1 g0584 ( .A1(G299), .A2(new_n754_), .ZN(new_n943_) );
  OR2_X1 g0585 ( .A1(new_n942_), .A2(new_n943_), .ZN(new_n944_) );
  AND2_X1 g0586 ( .A1(new_n940_), .A2(new_n944_), .ZN(new_n945_) );
  AND2_X1 g0587 ( .A1(new_n935_), .A2(new_n945_), .ZN(new_n946_) );
  AND2_X1 g0588 ( .A1(new_n946_), .A2(new_n926_), .ZN(new_n947_) );
  AND2_X1 g0589 ( .A1(new_n628_), .A2(new_n671_), .ZN(new_n948_) );
  AND2_X1 g0590 ( .A1(new_n627_), .A2(G1348), .ZN(new_n949_) );
  OR2_X1 g0591 ( .A1(new_n948_), .A2(new_n949_), .ZN(new_n950_) );
  AND2_X1 g0592 ( .A1(new_n566_), .A2(new_n670_), .ZN(new_n951_) );
  AND2_X1 g0593 ( .A1(new_n565_), .A2(G1341), .ZN(new_n952_) );
  OR2_X1 g0594 ( .A1(new_n951_), .A2(new_n952_), .ZN(new_n953_) );
  AND2_X1 g0595 ( .A1(new_n950_), .A2(new_n953_), .ZN(new_n954_) );
  AND2_X1 g0596 ( .A1(new_n947_), .A2(new_n954_), .ZN(new_n955_) );
  AND2_X1 g0597 ( .A1(new_n923_), .A2(new_n955_), .ZN(new_n956_) );
  AND2_X1 g0598 ( .A1(G16), .A2(KEYINPUT56), .ZN(new_n957_) );
  INV_X1 g0599 ( .A(new_n957_), .ZN(new_n958_) );
  OR2_X1 g0600 ( .A1(G16), .A2(KEYINPUT56), .ZN(new_n959_) );
  AND2_X1 g0601 ( .A1(new_n958_), .A2(new_n959_), .ZN(new_n960_) );
  OR2_X1 g0602 ( .A1(new_n956_), .A2(new_n960_), .ZN(new_n961_) );
  INV_X1 g0603 ( .A(KEYINPUT55), .ZN(new_n962_) );
  AND2_X1 g0604 ( .A1(G33), .A2(G2072), .ZN(new_n963_) );
  INV_X1 g0605 ( .A(new_n963_), .ZN(new_n964_) );
  AND2_X1 g0606 ( .A1(new_n964_), .A2(G28), .ZN(new_n965_) );
  OR2_X1 g0607 ( .A1(G33), .A2(G2072), .ZN(new_n966_) );
  AND2_X1 g0608 ( .A1(G26), .A2(G2067), .ZN(new_n967_) );
  INV_X1 g0609 ( .A(new_n967_), .ZN(new_n968_) );
  AND2_X1 g0610 ( .A1(new_n968_), .A2(new_n966_), .ZN(new_n969_) );
  AND2_X1 g0611 ( .A1(G25), .A2(G1991), .ZN(new_n970_) );
  INV_X1 g0612 ( .A(new_n970_), .ZN(new_n971_) );
  OR2_X1 g0613 ( .A1(G25), .A2(G1991), .ZN(new_n972_) );
  AND2_X1 g0614 ( .A1(new_n971_), .A2(new_n972_), .ZN(new_n973_) );
  AND2_X1 g0615 ( .A1(new_n969_), .A2(new_n973_), .ZN(new_n974_) );
  AND2_X1 g0616 ( .A1(new_n974_), .A2(new_n965_), .ZN(new_n975_) );
  INV_X1 g0617 ( .A(G27), .ZN(new_n976_) );
  AND2_X1 g0618 ( .A1(G2078), .A2(KEYINPUT25), .ZN(new_n977_) );
  INV_X1 g0619 ( .A(new_n977_), .ZN(new_n978_) );
  OR2_X1 g0620 ( .A1(G2078), .A2(KEYINPUT25), .ZN(new_n979_) );
  AND2_X1 g0621 ( .A1(new_n978_), .A2(new_n979_), .ZN(new_n980_) );
  INV_X1 g0622 ( .A(new_n980_), .ZN(new_n981_) );
  OR2_X1 g0623 ( .A1(new_n981_), .A2(new_n976_), .ZN(new_n982_) );
  OR2_X1 g0624 ( .A1(new_n980_), .A2(G27), .ZN(new_n983_) );
  AND2_X1 g0625 ( .A1(G32), .A2(G1996), .ZN(new_n984_) );
  INV_X1 g0626 ( .A(new_n984_), .ZN(new_n985_) );
  OR2_X1 g0627 ( .A1(G32), .A2(G1996), .ZN(new_n986_) );
  OR2_X1 g0628 ( .A1(G26), .A2(G2067), .ZN(new_n987_) );
  AND2_X1 g0629 ( .A1(new_n986_), .A2(new_n987_), .ZN(new_n988_) );
  AND2_X1 g0630 ( .A1(new_n988_), .A2(new_n985_), .ZN(new_n989_) );
  AND2_X1 g0631 ( .A1(new_n983_), .A2(new_n989_), .ZN(new_n990_) );
  AND2_X1 g0632 ( .A1(new_n990_), .A2(new_n982_), .ZN(new_n991_) );
  AND2_X1 g0633 ( .A1(new_n991_), .A2(new_n975_), .ZN(new_n992_) );
  AND2_X1 g0634 ( .A1(new_n992_), .A2(KEYINPUT53), .ZN(new_n993_) );
  INV_X1 g0635 ( .A(new_n993_), .ZN(new_n994_) );
  OR2_X1 g0636 ( .A1(new_n992_), .A2(KEYINPUT53), .ZN(new_n995_) );
  INV_X1 g0637 ( .A(G34), .ZN(new_n996_) );
  INV_X1 g0638 ( .A(KEYINPUT54), .ZN(new_n997_) );
  AND2_X1 g0639 ( .A1(new_n997_), .A2(G2084), .ZN(new_n998_) );
  AND2_X1 g0640 ( .A1(new_n741_), .A2(KEYINPUT54), .ZN(new_n999_) );
  OR2_X1 g0641 ( .A1(new_n998_), .A2(new_n999_), .ZN(new_n1000_) );
  INV_X1 g0642 ( .A(new_n1000_), .ZN(new_n1001_) );
  AND2_X1 g0643 ( .A1(new_n1001_), .A2(new_n996_), .ZN(new_n1002_) );
  AND2_X1 g0644 ( .A1(new_n1000_), .A2(G34), .ZN(new_n1003_) );
  OR2_X1 g0645 ( .A1(new_n1002_), .A2(new_n1003_), .ZN(new_n1004_) );
  AND2_X1 g0646 ( .A1(new_n710_), .A2(G35), .ZN(new_n1005_) );
  INV_X1 g0647 ( .A(G35), .ZN(new_n1006_) );
  AND2_X1 g0648 ( .A1(new_n1006_), .A2(G2090), .ZN(new_n1007_) );
  OR2_X1 g0649 ( .A1(new_n1005_), .A2(new_n1007_), .ZN(new_n1008_) );
  AND2_X1 g0650 ( .A1(new_n1004_), .A2(new_n1008_), .ZN(new_n1009_) );
  AND2_X1 g0651 ( .A1(new_n995_), .A2(new_n1009_), .ZN(new_n1010_) );
  AND2_X1 g0652 ( .A1(new_n1010_), .A2(new_n994_), .ZN(new_n1011_) );
  AND2_X1 g0653 ( .A1(new_n1011_), .A2(new_n962_), .ZN(new_n1012_) );
  INV_X1 g0654 ( .A(new_n1012_), .ZN(new_n1013_) );
  OR2_X1 g0655 ( .A1(new_n1011_), .A2(new_n962_), .ZN(new_n1014_) );
  AND2_X1 g0656 ( .A1(new_n1014_), .A2(new_n797_), .ZN(new_n1015_) );
  AND2_X1 g0657 ( .A1(new_n1015_), .A2(new_n1013_), .ZN(new_n1016_) );
  INV_X1 g0658 ( .A(new_n1016_), .ZN(new_n1017_) );
  INV_X1 g0659 ( .A(KEYINPUT61), .ZN(new_n1018_) );
  INV_X1 g0660 ( .A(KEYINPUT60), .ZN(new_n1019_) );
  AND2_X1 g0661 ( .A1(G1348), .A2(KEYINPUT59), .ZN(new_n1020_) );
  INV_X1 g0662 ( .A(new_n1020_), .ZN(new_n1021_) );
  OR2_X1 g0663 ( .A1(G1348), .A2(KEYINPUT59), .ZN(new_n1022_) );
  AND2_X1 g0664 ( .A1(new_n1021_), .A2(new_n1022_), .ZN(new_n1023_) );
  INV_X1 g0665 ( .A(new_n1023_), .ZN(new_n1024_) );
  AND2_X1 g0666 ( .A1(new_n1024_), .A2(G4), .ZN(new_n1025_) );
  INV_X1 g0667 ( .A(new_n1025_), .ZN(new_n1026_) );
  OR2_X1 g0668 ( .A1(new_n1024_), .A2(G4), .ZN(new_n1027_) );
  AND2_X1 g0669 ( .A1(new_n1026_), .A2(new_n1027_), .ZN(new_n1028_) );
  INV_X1 g0670 ( .A(new_n1028_), .ZN(new_n1029_) );
  AND2_X1 g0671 ( .A1(new_n749_), .A2(G6), .ZN(new_n1030_) );
  INV_X1 g0672 ( .A(new_n1030_), .ZN(new_n1031_) );
  OR2_X1 g0673 ( .A1(new_n749_), .A2(G6), .ZN(new_n1032_) );
  AND2_X1 g0674 ( .A1(new_n1031_), .A2(new_n1032_), .ZN(new_n1033_) );
  INV_X1 g0675 ( .A(new_n1033_), .ZN(new_n1034_) );
  AND2_X1 g0676 ( .A1(new_n670_), .A2(G19), .ZN(new_n1035_) );
  INV_X1 g0677 ( .A(new_n1035_), .ZN(new_n1036_) );
  OR2_X1 g0678 ( .A1(new_n670_), .A2(G19), .ZN(new_n1037_) );
  AND2_X1 g0679 ( .A1(new_n1036_), .A2(new_n1037_), .ZN(new_n1038_) );
  INV_X1 g0680 ( .A(new_n1038_), .ZN(new_n1039_) );
  AND2_X1 g0681 ( .A1(G20), .A2(G1956), .ZN(new_n1040_) );
  INV_X1 g0682 ( .A(new_n1040_), .ZN(new_n1041_) );
  OR2_X1 g0683 ( .A1(G20), .A2(G1956), .ZN(new_n1042_) );
  AND2_X1 g0684 ( .A1(new_n1041_), .A2(new_n1042_), .ZN(new_n1043_) );
  AND2_X1 g0685 ( .A1(new_n1039_), .A2(new_n1043_), .ZN(new_n1044_) );
  AND2_X1 g0686 ( .A1(new_n1044_), .A2(new_n1034_), .ZN(new_n1045_) );
  AND2_X1 g0687 ( .A1(new_n1029_), .A2(new_n1045_), .ZN(new_n1046_) );
  INV_X1 g0688 ( .A(new_n1046_), .ZN(new_n1047_) );
  AND2_X1 g0689 ( .A1(new_n1047_), .A2(new_n1019_), .ZN(new_n1048_) );
  AND2_X1 g0690 ( .A1(new_n1046_), .A2(KEYINPUT60), .ZN(new_n1049_) );
  OR2_X1 g0691 ( .A1(new_n1048_), .A2(new_n1049_), .ZN(new_n1050_) );
  INV_X1 g0692 ( .A(KEYINPUT58), .ZN(new_n1051_) );
  AND2_X1 g0693 ( .A1(new_n785_), .A2(G24), .ZN(new_n1052_) );
  INV_X1 g0694 ( .A(G24), .ZN(new_n1053_) );
  AND2_X1 g0695 ( .A1(new_n1053_), .A2(G1986), .ZN(new_n1054_) );
  OR2_X1 g0696 ( .A1(new_n1052_), .A2(new_n1054_), .ZN(new_n1055_) );
  AND2_X1 g0697 ( .A1(G23), .A2(G1976), .ZN(new_n1056_) );
  INV_X1 g0698 ( .A(new_n1056_), .ZN(new_n1057_) );
  OR2_X1 g0699 ( .A1(G23), .A2(G1976), .ZN(new_n1058_) );
  AND2_X1 g0700 ( .A1(new_n1057_), .A2(new_n1058_), .ZN(new_n1059_) );
  AND2_X1 g0701 ( .A1(G22), .A2(G1971), .ZN(new_n1060_) );
  INV_X1 g0702 ( .A(new_n1060_), .ZN(new_n1061_) );
  OR2_X1 g0703 ( .A1(G22), .A2(G1971), .ZN(new_n1062_) );
  AND2_X1 g0704 ( .A1(new_n1061_), .A2(new_n1062_), .ZN(new_n1063_) );
  AND2_X1 g0705 ( .A1(new_n1059_), .A2(new_n1063_), .ZN(new_n1064_) );
  AND2_X1 g0706 ( .A1(new_n1064_), .A2(new_n1055_), .ZN(new_n1065_) );
  AND2_X1 g0707 ( .A1(new_n1065_), .A2(new_n1051_), .ZN(new_n1066_) );
  INV_X1 g0708 ( .A(new_n1066_), .ZN(new_n1067_) );
  OR2_X1 g0709 ( .A1(new_n1065_), .A2(new_n1051_), .ZN(new_n1068_) );
  AND2_X1 g0710 ( .A1(G21), .A2(G1966), .ZN(new_n1069_) );
  INV_X1 g0711 ( .A(new_n1069_), .ZN(new_n1070_) );
  AND2_X1 g0712 ( .A1(G5), .A2(G1961), .ZN(new_n1071_) );
  INV_X1 g0713 ( .A(new_n1071_), .ZN(new_n1072_) );
  AND2_X1 g0714 ( .A1(new_n1070_), .A2(new_n1072_), .ZN(new_n1073_) );
  OR2_X1 g0715 ( .A1(G5), .A2(G1961), .ZN(new_n1074_) );
  OR2_X1 g0716 ( .A1(G21), .A2(G1966), .ZN(new_n1075_) );
  AND2_X1 g0717 ( .A1(new_n1074_), .A2(new_n1075_), .ZN(new_n1076_) );
  AND2_X1 g0718 ( .A1(new_n1073_), .A2(new_n1076_), .ZN(new_n1077_) );
  AND2_X1 g0719 ( .A1(new_n1068_), .A2(new_n1077_), .ZN(new_n1078_) );
  AND2_X1 g0720 ( .A1(new_n1078_), .A2(new_n1067_), .ZN(new_n1079_) );
  AND2_X1 g0721 ( .A1(new_n1050_), .A2(new_n1079_), .ZN(new_n1080_) );
  AND2_X1 g0722 ( .A1(new_n1080_), .A2(new_n1018_), .ZN(new_n1081_) );
  INV_X1 g0723 ( .A(new_n1081_), .ZN(new_n1082_) );
  INV_X1 g0724 ( .A(G16), .ZN(new_n1083_) );
  OR2_X1 g0725 ( .A1(new_n1080_), .A2(new_n1018_), .ZN(new_n1084_) );
  AND2_X1 g0726 ( .A1(new_n1084_), .A2(new_n1083_), .ZN(new_n1085_) );
  AND2_X1 g0727 ( .A1(new_n1085_), .A2(new_n1082_), .ZN(new_n1086_) );
  INV_X1 g0728 ( .A(new_n1086_), .ZN(new_n1087_) );
  AND2_X1 g0729 ( .A1(new_n1087_), .A2(G11), .ZN(new_n1088_) );
  AND2_X1 g0730 ( .A1(new_n1088_), .A2(new_n1017_), .ZN(new_n1089_) );
  AND2_X1 g0731 ( .A1(new_n961_), .A2(new_n1089_), .ZN(new_n1090_) );
  AND2_X1 g0732 ( .A1(new_n1090_), .A2(new_n908_), .ZN(new_n1091_) );
  INV_X1 g0733 ( .A(new_n1091_), .ZN(new_n1092_) );
  AND2_X1 g0734 ( .A1(new_n1092_), .A2(KEYINPUT62), .ZN(new_n1093_) );
  INV_X1 g0735 ( .A(new_n1093_), .ZN(new_n1094_) );
  OR2_X1 g0736 ( .A1(new_n1092_), .A2(KEYINPUT62), .ZN(new_n1095_) );
  AND2_X1 g0737 ( .A1(new_n1094_), .A2(new_n1095_), .ZN(G311) );
  INV_X1 g0738 ( .A(G311), .ZN(G150) );
  AND2_X1 g0739 ( .A1(new_n627_), .A2(G559), .ZN(new_n1098_) );
  INV_X1 g0740 ( .A(new_n1098_), .ZN(new_n1099_) );
  AND2_X1 g0741 ( .A1(new_n1099_), .A2(new_n566_), .ZN(new_n1100_) );
  AND2_X1 g0742 ( .A1(new_n1098_), .A2(new_n565_), .ZN(new_n1101_) );
  OR2_X1 g0743 ( .A1(new_n1101_), .A2(G860), .ZN(new_n1102_) );
  OR2_X1 g0744 ( .A1(new_n1102_), .A2(new_n1100_), .ZN(new_n1103_) );
  INV_X1 g0745 ( .A(new_n1103_), .ZN(new_n1104_) );
  AND2_X1 g0746 ( .A1(new_n473_), .A2(G55), .ZN(new_n1105_) );
  AND2_X1 g0747 ( .A1(new_n477_), .A2(G93), .ZN(new_n1106_) );
  OR2_X1 g0748 ( .A1(new_n1105_), .A2(new_n1106_), .ZN(new_n1107_) );
  AND2_X1 g0749 ( .A1(new_n483_), .A2(G80), .ZN(new_n1108_) );
  AND2_X1 g0750 ( .A1(new_n490_), .A2(G67), .ZN(new_n1109_) );
  OR2_X1 g0751 ( .A1(new_n1109_), .A2(new_n1108_), .ZN(new_n1110_) );
  OR2_X1 g0752 ( .A1(new_n1107_), .A2(new_n1110_), .ZN(new_n1111_) );
  INV_X1 g0753 ( .A(new_n1111_), .ZN(new_n1112_) );
  AND2_X1 g0754 ( .A1(new_n1104_), .A2(new_n1112_), .ZN(new_n1113_) );
  AND2_X1 g0755 ( .A1(new_n1103_), .A2(new_n1111_), .ZN(new_n1114_) );
  OR2_X1 g0756 ( .A1(new_n1113_), .A2(new_n1114_), .ZN(G145) );
  AND2_X1 g0757 ( .A1(new_n451_), .A2(G142), .ZN(new_n1116_) );
  AND2_X1 g0758 ( .A1(new_n453_), .A2(G106), .ZN(new_n1117_) );
  OR2_X1 g0759 ( .A1(new_n1116_), .A2(new_n1117_), .ZN(new_n1118_) );
  INV_X1 g0760 ( .A(new_n1118_), .ZN(new_n1119_) );
  AND2_X1 g0761 ( .A1(new_n1119_), .A2(KEYINPUT45), .ZN(new_n1120_) );
  INV_X1 g0762 ( .A(new_n1120_), .ZN(new_n1121_) );
  OR2_X1 g0763 ( .A1(new_n1119_), .A2(KEYINPUT45), .ZN(new_n1122_) );
  AND2_X1 g0764 ( .A1(new_n438_), .A2(G130), .ZN(new_n1123_) );
  AND2_X1 g0765 ( .A1(new_n436_), .A2(G118), .ZN(new_n1124_) );
  OR2_X1 g0766 ( .A1(new_n1123_), .A2(new_n1124_), .ZN(new_n1125_) );
  INV_X1 g0767 ( .A(new_n1125_), .ZN(new_n1126_) );
  AND2_X1 g0768 ( .A1(new_n1122_), .A2(new_n1126_), .ZN(new_n1127_) );
  AND2_X1 g0769 ( .A1(new_n1127_), .A2(new_n1121_), .ZN(new_n1128_) );
  AND2_X1 g0770 ( .A1(new_n1128_), .A2(new_n836_), .ZN(new_n1129_) );
  INV_X1 g0771 ( .A(new_n1129_), .ZN(new_n1130_) );
  OR2_X1 g0772 ( .A1(new_n1128_), .A2(new_n836_), .ZN(new_n1131_) );
  AND2_X1 g0773 ( .A1(new_n1130_), .A2(new_n1131_), .ZN(new_n1132_) );
  INV_X1 g0774 ( .A(new_n1132_), .ZN(new_n1133_) );
  AND2_X1 g0775 ( .A1(new_n1133_), .A2(G162), .ZN(new_n1134_) );
  AND2_X1 g0776 ( .A1(new_n1132_), .A2(new_n458_), .ZN(new_n1135_) );
  OR2_X1 g0777 ( .A1(new_n1134_), .A2(new_n1135_), .ZN(new_n1136_) );
  AND2_X1 g0778 ( .A1(new_n814_), .A2(new_n878_), .ZN(new_n1137_) );
  AND2_X1 g0779 ( .A1(new_n812_), .A2(G160), .ZN(new_n1138_) );
  OR2_X1 g0780 ( .A1(new_n1137_), .A2(new_n1138_), .ZN(new_n1139_) );
  AND2_X1 g0781 ( .A1(new_n867_), .A2(new_n1139_), .ZN(new_n1140_) );
  INV_X1 g0782 ( .A(new_n1140_), .ZN(new_n1141_) );
  OR2_X1 g0783 ( .A1(new_n867_), .A2(new_n1139_), .ZN(new_n1142_) );
  AND2_X1 g0784 ( .A1(new_n1141_), .A2(new_n1142_), .ZN(new_n1143_) );
  INV_X1 g0785 ( .A(new_n1143_), .ZN(new_n1144_) );
  AND2_X1 g0786 ( .A1(new_n1144_), .A2(new_n1136_), .ZN(new_n1145_) );
  INV_X1 g0787 ( .A(new_n1145_), .ZN(new_n1146_) );
  OR2_X1 g0788 ( .A1(new_n1144_), .A2(new_n1136_), .ZN(new_n1147_) );
  AND2_X1 g0789 ( .A1(new_n1146_), .A2(new_n1147_), .ZN(new_n1148_) );
  AND2_X1 g0790 ( .A1(new_n659_), .A2(new_n889_), .ZN(new_n1149_) );
  AND2_X1 g0791 ( .A1(new_n658_), .A2(new_n893_), .ZN(new_n1150_) );
  OR2_X1 g0792 ( .A1(new_n1149_), .A2(new_n1150_), .ZN(new_n1151_) );
  AND2_X1 g0793 ( .A1(KEYINPUT48), .A2(KEYINPUT46), .ZN(new_n1152_) );
  INV_X1 g0794 ( .A(new_n1152_), .ZN(new_n1153_) );
  OR2_X1 g0795 ( .A1(KEYINPUT48), .A2(KEYINPUT46), .ZN(new_n1154_) );
  AND2_X1 g0796 ( .A1(new_n1153_), .A2(new_n1154_), .ZN(new_n1155_) );
  INV_X1 g0797 ( .A(new_n1155_), .ZN(new_n1156_) );
  AND2_X1 g0798 ( .A1(new_n1151_), .A2(new_n1156_), .ZN(new_n1157_) );
  INV_X1 g0799 ( .A(new_n1157_), .ZN(new_n1158_) );
  OR2_X1 g0800 ( .A1(new_n1151_), .A2(new_n1156_), .ZN(new_n1159_) );
  AND2_X1 g0801 ( .A1(new_n1158_), .A2(new_n1159_), .ZN(new_n1160_) );
  INV_X1 g0802 ( .A(new_n1160_), .ZN(new_n1161_) );
  AND2_X1 g0803 ( .A1(new_n1161_), .A2(new_n466_), .ZN(new_n1162_) );
  AND2_X1 g0804 ( .A1(new_n1160_), .A2(G164), .ZN(new_n1163_) );
  OR2_X1 g0805 ( .A1(new_n1162_), .A2(new_n1163_), .ZN(new_n1164_) );
  INV_X1 g0806 ( .A(new_n1164_), .ZN(new_n1165_) );
  AND2_X1 g0807 ( .A1(new_n1148_), .A2(new_n1165_), .ZN(new_n1166_) );
  INV_X1 g0808 ( .A(new_n1166_), .ZN(new_n1167_) );
  INV_X1 g0809 ( .A(G37), .ZN(new_n1168_) );
  OR2_X1 g0810 ( .A1(new_n1148_), .A2(new_n1165_), .ZN(new_n1169_) );
  AND2_X1 g0811 ( .A1(new_n1169_), .A2(new_n1168_), .ZN(new_n1170_) );
  AND2_X1 g0812 ( .A1(new_n1170_), .A2(new_n1167_), .ZN(G395) );
  AND2_X1 g0813 ( .A1(new_n566_), .A2(G290), .ZN(new_n1172_) );
  AND2_X1 g0814 ( .A1(new_n565_), .A2(new_n936_), .ZN(new_n1173_) );
  OR2_X1 g0815 ( .A1(new_n1172_), .A2(new_n1173_), .ZN(new_n1174_) );
  AND2_X1 g0816 ( .A1(new_n1174_), .A2(new_n928_), .ZN(new_n1175_) );
  INV_X1 g0817 ( .A(new_n1175_), .ZN(new_n1176_) );
  OR2_X1 g0818 ( .A1(new_n1174_), .A2(new_n928_), .ZN(new_n1177_) );
  AND2_X1 g0819 ( .A1(new_n1176_), .A2(new_n1177_), .ZN(new_n1178_) );
  INV_X1 g0820 ( .A(new_n1178_), .ZN(new_n1179_) );
  AND2_X1 g0821 ( .A1(new_n941_), .A2(KEYINPUT19), .ZN(new_n1180_) );
  INV_X1 g0822 ( .A(new_n1180_), .ZN(new_n1181_) );
  OR2_X1 g0823 ( .A1(new_n941_), .A2(KEYINPUT19), .ZN(new_n1182_) );
  AND2_X1 g0824 ( .A1(new_n1181_), .A2(new_n1182_), .ZN(new_n1183_) );
  INV_X1 g0825 ( .A(new_n1183_), .ZN(new_n1184_) );
  AND2_X1 g0826 ( .A1(new_n1184_), .A2(G305), .ZN(new_n1185_) );
  AND2_X1 g0827 ( .A1(new_n1183_), .A2(new_n912_), .ZN(new_n1186_) );
  OR2_X1 g0828 ( .A1(new_n1185_), .A2(new_n1186_), .ZN(new_n1187_) );
  AND2_X1 g0829 ( .A1(new_n1179_), .A2(new_n1187_), .ZN(new_n1188_) );
  INV_X1 g0830 ( .A(new_n1188_), .ZN(new_n1189_) );
  OR2_X1 g0831 ( .A1(new_n1179_), .A2(new_n1187_), .ZN(new_n1190_) );
  AND2_X1 g0832 ( .A1(new_n1189_), .A2(new_n1190_), .ZN(new_n1191_) );
  INV_X1 g0833 ( .A(new_n1191_), .ZN(new_n1192_) );
  AND2_X1 g0834 ( .A1(G166), .A2(new_n1112_), .ZN(new_n1193_) );
  AND2_X1 g0835 ( .A1(G303), .A2(new_n1111_), .ZN(new_n1194_) );
  OR2_X1 g0836 ( .A1(new_n1193_), .A2(new_n1194_), .ZN(new_n1195_) );
  AND2_X1 g0837 ( .A1(new_n1192_), .A2(new_n1195_), .ZN(new_n1196_) );
  INV_X1 g0838 ( .A(new_n1196_), .ZN(new_n1197_) );
  OR2_X1 g0839 ( .A1(new_n1192_), .A2(new_n1195_), .ZN(new_n1198_) );
  AND2_X1 g0840 ( .A1(new_n1197_), .A2(new_n1198_), .ZN(new_n1199_) );
  INV_X1 g0841 ( .A(new_n1199_), .ZN(new_n1200_) );
  AND2_X1 g0842 ( .A1(new_n1200_), .A2(new_n1098_), .ZN(new_n1201_) );
  AND2_X1 g0843 ( .A1(new_n1199_), .A2(new_n1099_), .ZN(new_n1202_) );
  OR2_X1 g0844 ( .A1(new_n1201_), .A2(new_n1202_), .ZN(new_n1203_) );
  AND2_X1 g0845 ( .A1(new_n1203_), .A2(G868), .ZN(new_n1204_) );
  AND2_X1 g0846 ( .A1(new_n1111_), .A2(new_n615_), .ZN(new_n1205_) );
  OR2_X1 g0847 ( .A1(new_n1204_), .A2(new_n1205_), .ZN(G295) );
  AND2_X1 g0848 ( .A1(new_n588_), .A2(new_n628_), .ZN(new_n1207_) );
  AND2_X1 g0849 ( .A1(G286), .A2(new_n627_), .ZN(new_n1208_) );
  OR2_X1 g0850 ( .A1(new_n1208_), .A2(new_n1207_), .ZN(new_n1209_) );
  AND2_X1 g0851 ( .A1(new_n1200_), .A2(new_n1209_), .ZN(new_n1210_) );
  INV_X1 g0852 ( .A(new_n1210_), .ZN(new_n1211_) );
  OR2_X1 g0853 ( .A1(new_n1200_), .A2(new_n1209_), .ZN(new_n1212_) );
  AND2_X1 g0854 ( .A1(new_n1211_), .A2(new_n1212_), .ZN(new_n1213_) );
  AND2_X1 g0855 ( .A1(new_n1213_), .A2(G301), .ZN(new_n1214_) );
  INV_X1 g0856 ( .A(new_n1214_), .ZN(new_n1215_) );
  OR2_X1 g0857 ( .A1(new_n1213_), .A2(G301), .ZN(new_n1216_) );
  AND2_X1 g0858 ( .A1(new_n1216_), .A2(new_n1168_), .ZN(new_n1217_) );
  AND2_X1 g0859 ( .A1(new_n1217_), .A2(new_n1215_), .ZN(G397) );
  INV_X1 g0860 ( .A(G8), .ZN(new_n1219_) );
  INV_X1 g0861 ( .A(KEYINPUT26), .ZN(new_n1220_) );
  INV_X1 g0862 ( .A(G1384), .ZN(new_n1221_) );
  AND2_X1 g0863 ( .A1(new_n466_), .A2(new_n1221_), .ZN(new_n1222_) );
  AND2_X1 g0864 ( .A1(new_n441_), .A2(G40), .ZN(new_n1223_) );
  AND2_X1 g0865 ( .A1(new_n435_), .A2(new_n1223_), .ZN(new_n1224_) );
  AND2_X1 g0866 ( .A1(new_n1222_), .A2(new_n1224_), .ZN(new_n1225_) );
  AND2_X1 g0867 ( .A1(new_n1225_), .A2(G1996), .ZN(new_n1226_) );
  INV_X1 g0868 ( .A(new_n1226_), .ZN(new_n1227_) );
  OR2_X1 g0869 ( .A1(new_n1227_), .A2(new_n1220_), .ZN(new_n1228_) );
  OR2_X1 g0870 ( .A1(new_n1226_), .A2(KEYINPUT26), .ZN(new_n1229_) );
  OR2_X1 g0871 ( .A1(new_n1225_), .A2(new_n670_), .ZN(new_n1230_) );
  AND2_X1 g0872 ( .A1(new_n565_), .A2(new_n1230_), .ZN(new_n1231_) );
  AND2_X1 g0873 ( .A1(new_n1231_), .A2(new_n1229_), .ZN(new_n1232_) );
  AND2_X1 g0874 ( .A1(new_n1232_), .A2(new_n1228_), .ZN(new_n1233_) );
  AND2_X1 g0875 ( .A1(new_n1233_), .A2(new_n627_), .ZN(new_n1234_) );
  INV_X1 g0876 ( .A(new_n1225_), .ZN(new_n1235_) );
  AND2_X1 g0877 ( .A1(new_n1235_), .A2(G1348), .ZN(new_n1236_) );
  AND2_X1 g0878 ( .A1(new_n1225_), .A2(G2067), .ZN(new_n1237_) );
  OR2_X1 g0879 ( .A1(new_n1236_), .A2(new_n1237_), .ZN(new_n1238_) );
  INV_X1 g0880 ( .A(new_n1238_), .ZN(new_n1239_) );
  OR2_X1 g0881 ( .A1(new_n1234_), .A2(new_n1239_), .ZN(new_n1240_) );
  OR2_X1 g0882 ( .A1(new_n1233_), .A2(new_n627_), .ZN(new_n1241_) );
  AND2_X1 g0883 ( .A1(new_n1240_), .A2(new_n1241_), .ZN(new_n1242_) );
  INV_X1 g0884 ( .A(KEYINPUT27), .ZN(new_n1243_) );
  AND2_X1 g0885 ( .A1(new_n1225_), .A2(G2072), .ZN(new_n1244_) );
  AND2_X1 g0886 ( .A1(new_n1244_), .A2(new_n1243_), .ZN(new_n1245_) );
  INV_X1 g0887 ( .A(new_n1245_), .ZN(new_n1246_) );
  OR2_X1 g0888 ( .A1(new_n1244_), .A2(new_n1243_), .ZN(new_n1247_) );
  AND2_X1 g0889 ( .A1(new_n1235_), .A2(G1956), .ZN(new_n1248_) );
  INV_X1 g0890 ( .A(new_n1248_), .ZN(new_n1249_) );
  AND2_X1 g0891 ( .A1(new_n1247_), .A2(new_n1249_), .ZN(new_n1250_) );
  AND2_X1 g0892 ( .A1(new_n1250_), .A2(new_n1246_), .ZN(new_n1251_) );
  AND2_X1 g0893 ( .A1(new_n1251_), .A2(new_n941_), .ZN(new_n1252_) );
  OR2_X1 g0894 ( .A1(new_n1242_), .A2(new_n1252_), .ZN(new_n1253_) );
  OR2_X1 g0895 ( .A1(new_n1251_), .A2(new_n941_), .ZN(new_n1254_) );
  AND2_X1 g0896 ( .A1(new_n1254_), .A2(KEYINPUT28), .ZN(new_n1255_) );
  INV_X1 g0897 ( .A(new_n1255_), .ZN(new_n1256_) );
  OR2_X1 g0898 ( .A1(new_n1254_), .A2(KEYINPUT28), .ZN(new_n1257_) );
  AND2_X1 g0899 ( .A1(new_n1256_), .A2(new_n1257_), .ZN(new_n1258_) );
  INV_X1 g0900 ( .A(new_n1258_), .ZN(new_n1259_) );
  AND2_X1 g0901 ( .A1(new_n1253_), .A2(new_n1259_), .ZN(new_n1260_) );
  AND2_X1 g0902 ( .A1(new_n1260_), .A2(KEYINPUT29), .ZN(new_n1261_) );
  INV_X1 g0903 ( .A(new_n1261_), .ZN(new_n1262_) );
  OR2_X1 g0904 ( .A1(new_n1260_), .A2(KEYINPUT29), .ZN(new_n1263_) );
  AND2_X1 g0905 ( .A1(new_n1262_), .A2(new_n1263_), .ZN(new_n1264_) );
  AND2_X1 g0906 ( .A1(new_n1235_), .A2(new_n784_), .ZN(new_n1265_) );
  AND2_X1 g0907 ( .A1(new_n1225_), .A2(new_n981_), .ZN(new_n1266_) );
  OR2_X1 g0908 ( .A1(new_n1265_), .A2(new_n1266_), .ZN(new_n1267_) );
  AND2_X1 g0909 ( .A1(new_n1267_), .A2(G171), .ZN(new_n1268_) );
  OR2_X1 g0910 ( .A1(new_n1264_), .A2(new_n1268_), .ZN(new_n1269_) );
  INV_X1 g0911 ( .A(KEYINPUT31), .ZN(new_n1270_) );
  INV_X1 g0912 ( .A(KEYINPUT30), .ZN(new_n1271_) );
  AND2_X1 g0913 ( .A1(new_n1235_), .A2(G8), .ZN(new_n1272_) );
  AND2_X1 g0914 ( .A1(new_n1272_), .A2(new_n755_), .ZN(new_n1273_) );
  INV_X1 g0915 ( .A(new_n1273_), .ZN(new_n1274_) );
  AND2_X1 g0916 ( .A1(new_n1225_), .A2(new_n741_), .ZN(new_n1275_) );
  INV_X1 g0917 ( .A(new_n1275_), .ZN(new_n1276_) );
  AND2_X1 g0918 ( .A1(new_n1276_), .A2(G8), .ZN(new_n1277_) );
  AND2_X1 g0919 ( .A1(new_n1274_), .A2(new_n1277_), .ZN(new_n1278_) );
  AND2_X1 g0920 ( .A1(new_n1278_), .A2(new_n1271_), .ZN(new_n1279_) );
  INV_X1 g0921 ( .A(new_n1279_), .ZN(new_n1280_) );
  OR2_X1 g0922 ( .A1(new_n1278_), .A2(new_n1271_), .ZN(new_n1281_) );
  AND2_X1 g0923 ( .A1(new_n584_), .A2(new_n1281_), .ZN(new_n1282_) );
  AND2_X1 g0924 ( .A1(new_n1282_), .A2(new_n1280_), .ZN(new_n1283_) );
  INV_X1 g0925 ( .A(new_n1283_), .ZN(new_n1284_) );
  OR2_X1 g0926 ( .A1(new_n1267_), .A2(G171), .ZN(new_n1285_) );
  AND2_X1 g0927 ( .A1(new_n1284_), .A2(new_n1285_), .ZN(new_n1286_) );
  AND2_X1 g0928 ( .A1(new_n1286_), .A2(new_n1270_), .ZN(new_n1287_) );
  INV_X1 g0929 ( .A(new_n1287_), .ZN(new_n1288_) );
  OR2_X1 g0930 ( .A1(new_n1286_), .A2(new_n1270_), .ZN(new_n1289_) );
  AND2_X1 g0931 ( .A1(new_n1288_), .A2(new_n1289_), .ZN(new_n1290_) );
  INV_X1 g0932 ( .A(new_n1290_), .ZN(new_n1291_) );
  AND2_X1 g0933 ( .A1(new_n1269_), .A2(new_n1291_), .ZN(new_n1292_) );
  OR2_X1 g0934 ( .A1(new_n1292_), .A2(new_n588_), .ZN(new_n1293_) );
  AND2_X1 g0935 ( .A1(new_n1272_), .A2(new_n781_), .ZN(new_n1294_) );
  AND2_X1 g0936 ( .A1(new_n1225_), .A2(new_n710_), .ZN(new_n1295_) );
  OR2_X1 g0937 ( .A1(new_n1295_), .A2(G166), .ZN(new_n1296_) );
  OR2_X1 g0938 ( .A1(new_n1294_), .A2(new_n1296_), .ZN(new_n1297_) );
  AND2_X1 g0939 ( .A1(new_n1293_), .A2(new_n1297_), .ZN(new_n1298_) );
  OR2_X1 g0940 ( .A1(new_n1298_), .A2(new_n1219_), .ZN(new_n1299_) );
  AND2_X1 g0941 ( .A1(new_n1299_), .A2(KEYINPUT32), .ZN(new_n1300_) );
  INV_X1 g0942 ( .A(KEYINPUT32), .ZN(new_n1301_) );
  INV_X1 g0943 ( .A(KEYINPUT29), .ZN(new_n1302_) );
  INV_X1 g0944 ( .A(new_n1260_), .ZN(new_n1303_) );
  AND2_X1 g0945 ( .A1(new_n1303_), .A2(new_n1302_), .ZN(new_n1304_) );
  OR2_X1 g0946 ( .A1(new_n1304_), .A2(new_n1261_), .ZN(new_n1305_) );
  INV_X1 g0947 ( .A(new_n1268_), .ZN(new_n1306_) );
  AND2_X1 g0948 ( .A1(new_n1305_), .A2(new_n1306_), .ZN(new_n1307_) );
  OR2_X1 g0949 ( .A1(new_n1307_), .A2(new_n1290_), .ZN(new_n1308_) );
  AND2_X1 g0950 ( .A1(new_n1308_), .A2(G286), .ZN(new_n1309_) );
  INV_X1 g0951 ( .A(new_n1297_), .ZN(new_n1310_) );
  OR2_X1 g0952 ( .A1(new_n1309_), .A2(new_n1310_), .ZN(new_n1311_) );
  AND2_X1 g0953 ( .A1(new_n1311_), .A2(G8), .ZN(new_n1312_) );
  AND2_X1 g0954 ( .A1(new_n1312_), .A2(new_n1301_), .ZN(new_n1313_) );
  OR2_X1 g0955 ( .A1(new_n1300_), .A2(new_n1313_), .ZN(new_n1314_) );
  AND2_X1 g0956 ( .A1(new_n1275_), .A2(G8), .ZN(new_n1315_) );
  OR2_X1 g0957 ( .A1(new_n1273_), .A2(new_n1315_), .ZN(new_n1316_) );
  OR2_X1 g0958 ( .A1(new_n1292_), .A2(new_n1316_), .ZN(new_n1317_) );
  AND2_X1 g0959 ( .A1(new_n1314_), .A2(new_n1317_), .ZN(new_n1318_) );
  OR2_X1 g0960 ( .A1(new_n1318_), .A2(new_n930_), .ZN(new_n1319_) );
  INV_X1 g0961 ( .A(new_n1272_), .ZN(new_n1320_) );
  OR2_X1 g0962 ( .A1(new_n1320_), .A2(new_n932_), .ZN(new_n1321_) );
  INV_X1 g0963 ( .A(new_n1321_), .ZN(new_n1322_) );
  AND2_X1 g0964 ( .A1(new_n1319_), .A2(new_n1322_), .ZN(new_n1323_) );
  OR2_X1 g0965 ( .A1(new_n1323_), .A2(KEYINPUT33), .ZN(new_n1324_) );
  AND2_X1 g0966 ( .A1(new_n929_), .A2(KEYINPUT33), .ZN(new_n1325_) );
  AND2_X1 g0967 ( .A1(new_n1325_), .A2(new_n1272_), .ZN(new_n1326_) );
  OR2_X1 g0968 ( .A1(new_n915_), .A2(new_n1326_), .ZN(new_n1327_) );
  INV_X1 g0969 ( .A(new_n1327_), .ZN(new_n1328_) );
  AND2_X1 g0970 ( .A1(new_n1324_), .A2(new_n1328_), .ZN(new_n1329_) );
  AND2_X1 g0971 ( .A1(new_n710_), .A2(G8), .ZN(new_n1330_) );
  AND2_X1 g0972 ( .A1(G166), .A2(new_n1330_), .ZN(new_n1331_) );
  OR2_X1 g0973 ( .A1(new_n1318_), .A2(new_n1331_), .ZN(new_n1332_) );
  AND2_X1 g0974 ( .A1(new_n1332_), .A2(new_n1320_), .ZN(new_n1333_) );
  INV_X1 g0975 ( .A(new_n913_), .ZN(new_n1334_) );
  AND2_X1 g0976 ( .A1(new_n1334_), .A2(KEYINPUT24), .ZN(new_n1335_) );
  INV_X1 g0977 ( .A(new_n1335_), .ZN(new_n1336_) );
  OR2_X1 g0978 ( .A1(new_n1334_), .A2(KEYINPUT24), .ZN(new_n1337_) );
  AND2_X1 g0979 ( .A1(new_n1337_), .A2(new_n1272_), .ZN(new_n1338_) );
  AND2_X1 g0980 ( .A1(new_n1338_), .A2(new_n1336_), .ZN(new_n1339_) );
  OR2_X1 g0981 ( .A1(new_n1333_), .A2(new_n1339_), .ZN(new_n1340_) );
  OR2_X1 g0982 ( .A1(new_n1329_), .A2(new_n1340_), .ZN(new_n1341_) );
  INV_X1 g0983 ( .A(new_n1222_), .ZN(new_n1342_) );
  AND2_X1 g0984 ( .A1(new_n1342_), .A2(new_n1224_), .ZN(new_n1343_) );
  AND2_X1 g0985 ( .A1(new_n873_), .A2(new_n1343_), .ZN(new_n1344_) );
  AND2_X1 g0986 ( .A1(new_n939_), .A2(new_n1343_), .ZN(new_n1345_) );
  AND2_X1 g0987 ( .A1(new_n891_), .A2(new_n1343_), .ZN(new_n1346_) );
  OR2_X1 g0988 ( .A1(new_n1345_), .A2(new_n1346_), .ZN(new_n1347_) );
  OR2_X1 g0989 ( .A1(new_n1344_), .A2(new_n1347_), .ZN(new_n1348_) );
  INV_X1 g0990 ( .A(new_n1348_), .ZN(new_n1349_) );
  AND2_X1 g0991 ( .A1(new_n1341_), .A2(new_n1349_), .ZN(new_n1350_) );
  INV_X1 g0992 ( .A(KEYINPUT39), .ZN(new_n1351_) );
  INV_X1 g0993 ( .A(new_n1346_), .ZN(new_n1352_) );
  OR2_X1 g0994 ( .A1(new_n937_), .A2(new_n894_), .ZN(new_n1353_) );
  AND2_X1 g0995 ( .A1(new_n1352_), .A2(new_n1353_), .ZN(new_n1354_) );
  OR2_X1 g0996 ( .A1(new_n1354_), .A2(new_n838_), .ZN(new_n1355_) );
  INV_X1 g0997 ( .A(new_n1355_), .ZN(new_n1356_) );
  AND2_X1 g0998 ( .A1(new_n1356_), .A2(new_n1351_), .ZN(new_n1357_) );
  AND2_X1 g0999 ( .A1(new_n1355_), .A2(KEYINPUT39), .ZN(new_n1358_) );
  OR2_X1 g1000 ( .A1(new_n1344_), .A2(new_n1358_), .ZN(new_n1359_) );
  OR2_X1 g1001 ( .A1(new_n1359_), .A2(new_n1357_), .ZN(new_n1360_) );
  AND2_X1 g1002 ( .A1(new_n1360_), .A2(new_n876_), .ZN(new_n1361_) );
  INV_X1 g1003 ( .A(new_n1361_), .ZN(new_n1362_) );
  AND2_X1 g1004 ( .A1(new_n1362_), .A2(new_n1343_), .ZN(new_n1363_) );
  OR2_X1 g1005 ( .A1(new_n1350_), .A2(new_n1363_), .ZN(new_n1364_) );
  AND2_X1 g1006 ( .A1(new_n1364_), .A2(KEYINPUT40), .ZN(new_n1365_) );
  INV_X1 g1007 ( .A(KEYINPUT40), .ZN(new_n1366_) );
  INV_X1 g1008 ( .A(KEYINPUT33), .ZN(new_n1367_) );
  INV_X1 g1009 ( .A(new_n930_), .ZN(new_n1368_) );
  OR2_X1 g1010 ( .A1(new_n1312_), .A2(new_n1301_), .ZN(new_n1369_) );
  OR2_X1 g1011 ( .A1(new_n1299_), .A2(KEYINPUT32), .ZN(new_n1370_) );
  AND2_X1 g1012 ( .A1(new_n1369_), .A2(new_n1370_), .ZN(new_n1371_) );
  INV_X1 g1013 ( .A(new_n1317_), .ZN(new_n1372_) );
  OR2_X1 g1014 ( .A1(new_n1371_), .A2(new_n1372_), .ZN(new_n1373_) );
  AND2_X1 g1015 ( .A1(new_n1373_), .A2(new_n1368_), .ZN(new_n1374_) );
  OR2_X1 g1016 ( .A1(new_n1374_), .A2(new_n1321_), .ZN(new_n1375_) );
  AND2_X1 g1017 ( .A1(new_n1375_), .A2(new_n1367_), .ZN(new_n1376_) );
  OR2_X1 g1018 ( .A1(new_n1376_), .A2(new_n1327_), .ZN(new_n1377_) );
  INV_X1 g1019 ( .A(new_n1340_), .ZN(new_n1378_) );
  AND2_X1 g1020 ( .A1(new_n1377_), .A2(new_n1378_), .ZN(new_n1379_) );
  OR2_X1 g1021 ( .A1(new_n1379_), .A2(new_n1348_), .ZN(new_n1380_) );
  INV_X1 g1022 ( .A(new_n1363_), .ZN(new_n1381_) );
  AND2_X1 g1023 ( .A1(new_n1380_), .A2(new_n1381_), .ZN(new_n1382_) );
  AND2_X1 g1024 ( .A1(new_n1382_), .A2(new_n1366_), .ZN(new_n1383_) );
  OR2_X1 g1025 ( .A1(new_n1365_), .A2(new_n1383_), .ZN(G329) );
  INV_X1 g1026 ( .A(G397), .ZN(new_n1386_) );
  INV_X1 g1027 ( .A(G395), .ZN(new_n1387_) );
  INV_X1 g1028 ( .A(KEYINPUT49), .ZN(new_n1388_) );
  OR2_X1 g1029 ( .A1(G229), .A2(G227), .ZN(new_n1389_) );
  AND2_X1 g1030 ( .A1(new_n1389_), .A2(new_n1388_), .ZN(new_n1390_) );
  INV_X1 g1031 ( .A(new_n1390_), .ZN(new_n1391_) );
  OR2_X1 g1032 ( .A1(new_n1389_), .A2(new_n1388_), .ZN(new_n1392_) );
  OR2_X1 g1033 ( .A1(G401), .A2(new_n569_), .ZN(new_n1393_) );
  INV_X1 g1034 ( .A(new_n1393_), .ZN(new_n1394_) );
  AND2_X1 g1035 ( .A1(new_n1392_), .A2(new_n1394_), .ZN(new_n1395_) );
  AND2_X1 g1036 ( .A1(new_n1395_), .A2(new_n1391_), .ZN(new_n1396_) );
  AND2_X1 g1037 ( .A1(new_n1387_), .A2(new_n1396_), .ZN(new_n1397_) );
  AND2_X1 g1038 ( .A1(new_n1386_), .A2(new_n1397_), .ZN(G308) );
  INV_X1 g1039 ( .A(G308), .ZN(G225) );
  assign   G231 = 1'b0;
  BUF_X1 g1040 ( .A(G452), .Z(G350) );
  BUF_X1 g1041 ( .A(G452), .Z(G335) );
  BUF_X1 g1042 ( .A(G452), .Z(G409) );
  BUF_X1 g1043 ( .A(G1083), .Z(G369) );
  BUF_X1 g1044 ( .A(G1083), .Z(G367) );
  BUF_X1 g1045 ( .A(G2066), .Z(G411) );
  BUF_X1 g1046 ( .A(G2066), .Z(G337) );
  BUF_X1 g1047 ( .A(G2066), .Z(G384) );
  BUF_X1 g1048 ( .A(G452), .Z(G391) );
  OR2_X1 g1049 ( .A1(new_n629_), .A2(new_n630_), .ZN(G321) );
  AND2_X1 g1050 ( .A1(new_n632_), .A2(new_n633_), .ZN(G280) );
  AND2_X1 g1051 ( .A1(new_n643_), .A2(new_n644_), .ZN(G323) );
  OR2_X1 g1052 ( .A1(new_n1204_), .A2(new_n1205_), .ZN(G331) );
endmodule


