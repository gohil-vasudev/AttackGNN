module s35932 ( CK, CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_10, CRC_OUT_1_11, 
        CRC_OUT_1_12, CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, 
        CRC_OUT_1_17, CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_2, CRC_OUT_1_20, 
        CRC_OUT_1_21, CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, 
        CRC_OUT_1_26, CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_3, 
        CRC_OUT_1_30, CRC_OUT_1_31, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, 
        CRC_OUT_1_7, CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_2_0, CRC_OUT_2_1, 
        CRC_OUT_2_10, CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, 
        CRC_OUT_2_15, CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, 
        CRC_OUT_2_2, CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, 
        CRC_OUT_2_24, CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, 
        CRC_OUT_2_29, CRC_OUT_2_3, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_2_4, 
        CRC_OUT_2_5, CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, 
        CRC_OUT_3_0, CRC_OUT_3_1, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, 
        CRC_OUT_3_13, CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, 
        CRC_OUT_3_18, CRC_OUT_3_19, CRC_OUT_3_2, CRC_OUT_3_20, CRC_OUT_3_21, 
        CRC_OUT_3_22, CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, 
        CRC_OUT_3_27, CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_3, CRC_OUT_3_30, 
        CRC_OUT_3_31, CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, 
        CRC_OUT_3_8, CRC_OUT_3_9, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_10, 
        CRC_OUT_4_11, CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, 
        CRC_OUT_4_16, CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_2, 
        CRC_OUT_4_20, CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, 
        CRC_OUT_4_25, CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, 
        CRC_OUT_4_3, CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_4_4, CRC_OUT_4_5, 
        CRC_OUT_4_6, CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_5_0, 
        CRC_OUT_5_1, CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, 
        CRC_OUT_5_14, CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, 
        CRC_OUT_5_19, CRC_OUT_5_2, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, 
        CRC_OUT_5_23, CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, 
        CRC_OUT_5_28, CRC_OUT_5_29, CRC_OUT_5_3, CRC_OUT_5_30, CRC_OUT_5_31, 
        CRC_OUT_5_4, CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, 
        CRC_OUT_5_9, CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_10, CRC_OUT_6_11, 
        CRC_OUT_6_12, CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, 
        CRC_OUT_6_17, CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_2, CRC_OUT_6_20, 
        CRC_OUT_6_21, CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, 
        CRC_OUT_6_26, CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_3, 
        CRC_OUT_6_30, CRC_OUT_6_31, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, 
        CRC_OUT_6_7, CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_7_0, CRC_OUT_7_1, 
        CRC_OUT_7_10, CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, 
        CRC_OUT_7_15, CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, 
        CRC_OUT_7_2, CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, 
        CRC_OUT_7_24, CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, 
        CRC_OUT_7_29, CRC_OUT_7_3, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_7_4, 
        CRC_OUT_7_5, CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, 
        CRC_OUT_8_0, CRC_OUT_8_1, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, 
        CRC_OUT_8_13, CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, 
        CRC_OUT_8_18, CRC_OUT_8_19, CRC_OUT_8_2, CRC_OUT_8_20, CRC_OUT_8_21, 
        CRC_OUT_8_22, CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, 
        CRC_OUT_8_27, CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_3, CRC_OUT_8_30, 
        CRC_OUT_8_31, CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, 
        CRC_OUT_8_8, CRC_OUT_8_9, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_10, 
        CRC_OUT_9_11, CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, 
        CRC_OUT_9_16, CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_2, 
        CRC_OUT_9_20, CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, 
        CRC_OUT_9_25, CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, 
        CRC_OUT_9_3, CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_9_4, CRC_OUT_9_5, 
        CRC_OUT_9_6, CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, DATA_0_0, DATA_0_1, 
        DATA_0_10, DATA_0_11, DATA_0_12, DATA_0_13, DATA_0_14, DATA_0_15, 
        DATA_0_16, DATA_0_17, DATA_0_18, DATA_0_19, DATA_0_2, DATA_0_20, 
        DATA_0_21, DATA_0_22, DATA_0_23, DATA_0_24, DATA_0_25, DATA_0_26, 
        DATA_0_27, DATA_0_28, DATA_0_29, DATA_0_3, DATA_0_30, DATA_0_31, 
        DATA_0_4, DATA_0_5, DATA_0_6, DATA_0_7, DATA_0_8, DATA_0_9, DATA_9_0, 
        DATA_9_1, DATA_9_10, DATA_9_11, DATA_9_12, DATA_9_13, DATA_9_14, 
        DATA_9_15, DATA_9_16, DATA_9_17, DATA_9_18, DATA_9_19, DATA_9_2, 
        DATA_9_20, DATA_9_21, DATA_9_22, DATA_9_23, DATA_9_24, DATA_9_25, 
        DATA_9_26, DATA_9_27, DATA_9_28, DATA_9_29, DATA_9_3, DATA_9_30, 
        DATA_9_31, DATA_9_4, DATA_9_5, DATA_9_6, DATA_9_7, DATA_9_8, DATA_9_9, 
        RESET, TM0, TM1, test_se, test_si1, test_so1, test_si2, test_so2, 
        test_si3, test_so3, test_si4, test_so4, test_si5, test_so5, test_si6, 
        test_so6, test_si7, test_so7, test_si8, test_so8, test_si9, test_so9, 
        test_si10, test_so10, test_si11, test_so11, test_si12, test_so12, 
        test_si13, test_so13, test_si14, test_so14, test_si15, test_so15, 
        test_si16, test_so16, test_si17, test_so17, test_si18, test_so18, 
        test_si19, test_so19, test_si20, test_so20, test_si21, test_so21, 
        test_si22, test_so22, test_si23, test_so23, test_si24, test_so24, 
        test_si25, test_so25, test_si26, test_so26, test_si27, test_so27, 
        test_si28, test_so28, test_si29, test_so29, test_si30, test_so30, 
        test_si31, test_so31, test_si32, test_so32, test_si33, test_so33, 
        test_si34, test_so34, test_si35, test_so35, test_si36, test_so36, 
        test_si37, test_so37, test_si38, test_so38, test_si39, test_so39, 
        test_si40, test_so40, test_si41, test_so41, test_si42, test_so42, 
        test_si43, test_so43, test_si44, test_so44, test_si45, test_so45, 
        test_si46, test_so46, test_si47, test_so47, test_si48, test_so48, 
        test_si49, test_so49, test_si50, test_so50, test_si51, test_so51, 
        test_si52, test_so52, test_si53, test_so53, test_si54, test_so54, 
        test_si55, test_so55, test_si56, test_so56, test_si57, test_so57, 
        test_si58, test_so58, test_si59, test_so59, test_si60, test_so60, 
        test_si61, test_so61, test_si62, test_so62, test_si63, test_so63, 
        test_si64, test_so64, test_si65, test_so65, test_si66, test_so66, 
        test_si67, test_so67, test_si68, test_so68, test_si69, test_so69, 
        test_si70, test_so70, test_si71, test_so71, test_si72, test_so72, 
        test_si73, test_so73, test_si74, test_so74, test_si75, test_so75, 
        test_si76, test_so76, test_si77, test_so77, test_si78, test_so78, 
        test_si79, test_so79, test_si80, test_so80, test_si81, test_so81, 
        test_si82, test_so82, test_si83, test_so83, test_si84, test_so84, 
        test_si85, test_so85, test_si86, test_so86, test_si87, test_so87, 
        test_si88, test_so88, test_si89, test_so89, test_si90, test_so90, 
        test_si91, test_so91, test_si92, test_so92, test_si93, test_so93, 
        test_si94, test_so94, test_si95, test_so95, test_si96, test_so96, 
        test_si97, test_so97, test_si98, test_so98, test_si99, test_so99, 
        test_si100, test_so100 );
  input CK, DATA_0_0, DATA_0_1, DATA_0_10, DATA_0_11, DATA_0_12, DATA_0_13,
         DATA_0_14, DATA_0_15, DATA_0_16, DATA_0_17, DATA_0_18, DATA_0_19,
         DATA_0_2, DATA_0_20, DATA_0_21, DATA_0_22, DATA_0_23, DATA_0_24,
         DATA_0_25, DATA_0_26, DATA_0_27, DATA_0_28, DATA_0_29, DATA_0_3,
         DATA_0_30, DATA_0_31, DATA_0_4, DATA_0_5, DATA_0_6, DATA_0_7,
         DATA_0_8, DATA_0_9, RESET, TM0, TM1, test_se, test_si1, test_si2,
         test_si3, test_si4, test_si5, test_si6, test_si7, test_si8, test_si9,
         test_si10, test_si11, test_si12, test_si13, test_si14, test_si15,
         test_si16, test_si17, test_si18, test_si19, test_si20, test_si21,
         test_si22, test_si23, test_si24, test_si25, test_si26, test_si27,
         test_si28, test_si29, test_si30, test_si31, test_si32, test_si33,
         test_si34, test_si35, test_si36, test_si37, test_si38, test_si39,
         test_si40, test_si41, test_si42, test_si43, test_si44, test_si45,
         test_si46, test_si47, test_si48, test_si49, test_si50, test_si51,
         test_si52, test_si53, test_si54, test_si55, test_si56, test_si57,
         test_si58, test_si59, test_si60, test_si61, test_si62, test_si63,
         test_si64, test_si65, test_si66, test_si67, test_si68, test_si69,
         test_si70, test_si71, test_si72, test_si73, test_si74, test_si75,
         test_si76, test_si77, test_si78, test_si79, test_si80, test_si81,
         test_si82, test_si83, test_si84, test_si85, test_si86, test_si87,
         test_si88, test_si89, test_si90, test_si91, test_si92, test_si93,
         test_si94, test_si95, test_si96, test_si97, test_si98, test_si99,
         test_si100;
  output CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_10, CRC_OUT_1_11, CRC_OUT_1_12,
         CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, CRC_OUT_1_17,
         CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_2, CRC_OUT_1_20, CRC_OUT_1_21,
         CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, CRC_OUT_1_26,
         CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_3, CRC_OUT_1_30,
         CRC_OUT_1_31, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, CRC_OUT_1_7,
         CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_2_0, CRC_OUT_2_1, CRC_OUT_2_10,
         CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, CRC_OUT_2_15,
         CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, CRC_OUT_2_2,
         CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, CRC_OUT_2_24,
         CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, CRC_OUT_2_29,
         CRC_OUT_2_3, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_2_4, CRC_OUT_2_5,
         CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, CRC_OUT_3_0,
         CRC_OUT_3_1, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, CRC_OUT_3_13,
         CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, CRC_OUT_3_18,
         CRC_OUT_3_19, CRC_OUT_3_2, CRC_OUT_3_20, CRC_OUT_3_21, CRC_OUT_3_22,
         CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, CRC_OUT_3_27,
         CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_3, CRC_OUT_3_30, CRC_OUT_3_31,
         CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, CRC_OUT_3_8,
         CRC_OUT_3_9, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_10, CRC_OUT_4_11,
         CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, CRC_OUT_4_16,
         CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_2, CRC_OUT_4_20,
         CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, CRC_OUT_4_25,
         CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, CRC_OUT_4_3,
         CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_4_4, CRC_OUT_4_5, CRC_OUT_4_6,
         CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_5_0, CRC_OUT_5_1,
         CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, CRC_OUT_5_14,
         CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, CRC_OUT_5_19,
         CRC_OUT_5_2, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, CRC_OUT_5_23,
         CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, CRC_OUT_5_28,
         CRC_OUT_5_29, CRC_OUT_5_3, CRC_OUT_5_30, CRC_OUT_5_31, CRC_OUT_5_4,
         CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, CRC_OUT_5_9,
         CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_10, CRC_OUT_6_11, CRC_OUT_6_12,
         CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, CRC_OUT_6_17,
         CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_2, CRC_OUT_6_20, CRC_OUT_6_21,
         CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, CRC_OUT_6_26,
         CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_3, CRC_OUT_6_30,
         CRC_OUT_6_31, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, CRC_OUT_6_7,
         CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_7_0, CRC_OUT_7_1, CRC_OUT_7_10,
         CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, CRC_OUT_7_15,
         CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, CRC_OUT_7_2,
         CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, CRC_OUT_7_24,
         CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, CRC_OUT_7_29,
         CRC_OUT_7_3, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_7_4, CRC_OUT_7_5,
         CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, CRC_OUT_8_0,
         CRC_OUT_8_1, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, CRC_OUT_8_13,
         CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, CRC_OUT_8_18,
         CRC_OUT_8_19, CRC_OUT_8_2, CRC_OUT_8_20, CRC_OUT_8_21, CRC_OUT_8_22,
         CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, CRC_OUT_8_27,
         CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_3, CRC_OUT_8_30, CRC_OUT_8_31,
         CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, CRC_OUT_8_8,
         CRC_OUT_8_9, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_10, CRC_OUT_9_11,
         CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, CRC_OUT_9_16,
         CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_2, CRC_OUT_9_20,
         CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, CRC_OUT_9_25,
         CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, CRC_OUT_9_3,
         CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_9_4, CRC_OUT_9_5, CRC_OUT_9_6,
         CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, DATA_9_0, DATA_9_1, DATA_9_10,
         DATA_9_11, DATA_9_12, DATA_9_13, DATA_9_14, DATA_9_15, DATA_9_16,
         DATA_9_17, DATA_9_18, DATA_9_19, DATA_9_2, DATA_9_20, DATA_9_21,
         DATA_9_22, DATA_9_23, DATA_9_24, DATA_9_25, DATA_9_26, DATA_9_27,
         DATA_9_28, DATA_9_29, DATA_9_3, DATA_9_30, DATA_9_31, DATA_9_4,
         DATA_9_5, DATA_9_6, DATA_9_7, DATA_9_8, DATA_9_9, test_so1, test_so2,
         test_so3, test_so4, test_so5, test_so6, test_so7, test_so8, test_so9,
         test_so10, test_so11, test_so12, test_so13, test_so14, test_so15,
         test_so16, test_so17, test_so18, test_so19, test_so20, test_so21,
         test_so22, test_so23, test_so24, test_so25, test_so26, test_so27,
         test_so28, test_so29, test_so30, test_so31, test_so32, test_so33,
         test_so34, test_so35, test_so36, test_so37, test_so38, test_so39,
         test_so40, test_so41, test_so42, test_so43, test_so44, test_so45,
         test_so46, test_so47, test_so48, test_so49, test_so50, test_so51,
         test_so52, test_so53, test_so54, test_so55, test_so56, test_so57,
         test_so58, test_so59, test_so60, test_so61, test_so62, test_so63,
         test_so64, test_so65, test_so66, test_so67, test_so68, test_so69,
         test_so70, test_so71, test_so72, test_so73, test_so74, test_so75,
         test_so76, test_so77, test_so78, test_so79, test_so80, test_so81,
         test_so82, test_so83, test_so84, test_so85, test_so86, test_so87,
         test_so88, test_so89, test_so90, test_so91, test_so92, test_so93,
         test_so94, test_so95, test_so96, test_so97, test_so98, test_so99,
         test_so100;
  wire   test_so9, test_so10, test_so20, test_so21, test_so31, test_so32,
         test_so42, test_so43, test_so53, test_so54, test_so65, test_so66,
         test_so76, test_so77, test_so87, test_so88, test_so99, test_so100,
         WX484, WX485, WX486, WX487, WX488, WX489, WX490, WX491, WX492, WX493,
         WX494, WX495, WX496, WX497, WX498, WX499, WX500, WX501, WX502, WX503,
         WX504, WX505, WX506, WX507, WX508, WX509, WX510, WX511, WX512, WX513,
         WX514, WX515, WX516, WX517, WX518, WX520, WX521, WX522, WX523, WX524,
         WX525, WX526, WX527, WX528, WX529, WX530, WX531, WX532, WX533, WX534,
         WX535, WX536, WX537, WX538, WX539, WX540, WX541, WX542, WX543, WX544,
         WX545, WX546, WX547, WX644, WX645, n3529, WX646, WX647, n3527, WX648,
         WX649, n3525, WX650, WX652, WX653, n3521, WX654, WX655, n3519, WX656,
         WX657, n3517, WX658, WX659, n3515, WX660, WX661, n3513, WX662, WX663,
         n3511, WX664, WX665, n3509, WX666, WX667, n3507, WX668, WX669, n3505,
         WX670, WX671, n3503, WX672, WX673, n3501, WX674, WX675, n3499, WX676,
         WX677, n3497, WX678, WX679, n3495, WX680, WX681, n3493, WX682, WX683,
         n3491, WX684, WX685, n3489, WX686, WX688, WX689, n3485, WX690, WX691,
         n3483, WX692, WX693, n3481, WX694, WX695, n3479, WX696, WX697, n3477,
         WX698, WX699, n3475, WX700, WX701, n3473, WX702, WX703, n3471, WX704,
         WX705, n3469, WX706, WX707, n3467, WX708, WX709, WX710, WX711, WX712,
         WX713, WX714, WX715, WX716, WX717, WX718, WX719, WX720, WX721, WX722,
         WX724, WX725, WX726, WX727, WX728, WX729, WX730, WX731, WX732, WX733,
         WX734, WX735, WX736, WX737, WX738, WX739, WX740, WX741, WX742, WX743,
         WX744, WX745, WX746, WX747, WX748, WX749, WX750, WX751, WX752, WX753,
         WX754, WX755, WX756, WX757, WX758, WX760, WX761, WX762, WX763, WX764,
         WX765, WX766, WX767, WX768, WX769, WX770, WX771, WX772, WX773, WX774,
         WX775, WX776, WX777, WX778, WX779, WX780, WX781, WX782, WX783, WX784,
         WX785, WX786, WX787, WX788, WX789, WX790, WX791, WX792, WX793, WX794,
         WX796, WX797, WX798, WX799, WX800, WX801, WX802, WX803, WX804, WX805,
         WX806, WX807, WX808, WX809, WX810, WX811, WX812, WX813, WX814, WX815,
         WX816, WX817, WX818, WX819, WX820, WX821, WX822, WX823, WX824, WX825,
         WX826, WX827, WX828, WX829, WX830, WX832, WX833, WX834, WX835, WX836,
         WX837, WX838, WX839, WX840, WX841, WX842, WX843, WX844, WX845, WX846,
         WX847, WX848, WX849, WX850, WX851, WX852, WX853, WX854, WX855, WX856,
         WX857, WX858, WX859, WX860, WX861, WX862, WX863, WX864, WX865, WX866,
         WX868, WX869, WX870, WX871, WX872, WX873, WX874, WX875, WX876, WX877,
         WX878, WX879, WX880, WX881, WX882, WX883, WX884, WX885, WX886, WX887,
         WX888, WX889, WX890, WX891, WX892, WX893, WX894, WX895, WX896, WX897,
         WX898, WX899, WX1264, DFF_160_n1, WX1266, WX1268, DFF_162_n1, WX1270,
         DFF_163_n1, WX1272, DFF_164_n1, WX1274, DFF_165_n1, WX1276,
         DFF_166_n1, WX1278, DFF_167_n1, WX1280, DFF_168_n1, WX1282,
         DFF_169_n1, WX1284, DFF_170_n1, WX1286, DFF_171_n1, WX1288,
         DFF_172_n1, WX1290, DFF_173_n1, WX1292, DFF_174_n1, WX1294,
         DFF_175_n1, WX1296, DFF_176_n1, WX1298, DFF_177_n1, WX1300,
         DFF_178_n1, WX1302, WX1304, DFF_180_n1, WX1306, DFF_181_n1, WX1308,
         DFF_182_n1, WX1310, DFF_183_n1, WX1312, DFF_184_n1, WX1314,
         DFF_185_n1, WX1316, DFF_186_n1, WX1318, DFF_187_n1, WX1320,
         DFF_188_n1, WX1322, DFF_189_n1, WX1324, DFF_190_n1, WX1326,
         DFF_191_n1, WX1778, n8702, n8701, n8700, n8699, n8696, n8695, n8694,
         n8693, n8692, n8691, n8690, n8689, n8688, n8687, n8686, n8685, n8684,
         n8683, n8682, n8681, n8680, n8677, n8676, n8675, n8674, n8673, n8672,
         n8671, WX1839, n8670, WX1937, n8669, WX1939, n8668, WX1941, n8667,
         WX1943, n8666, WX1945, n8665, WX1947, n8664, WX1949, n8663, WX1951,
         n8662, WX1953, n8661, WX1955, WX1957, n8658, WX1959, n8657, WX1961,
         n8656, WX1963, n8655, WX1965, n8654, WX1967, n8653, WX1969, WX1970,
         WX1971, WX1972, WX1973, WX1974, WX1975, WX1976, WX1977, WX1978,
         WX1979, WX1980, WX1981, WX1982, WX1983, WX1984, WX1985, WX1986,
         WX1987, WX1988, WX1989, WX1990, WX1991, WX1993, WX1994, WX1995,
         WX1996, WX1997, WX1998, WX1999, WX2000, WX2001, WX2002, WX2003,
         WX2004, WX2005, WX2006, WX2007, WX2008, WX2009, WX2010, WX2011,
         WX2012, WX2013, WX2014, WX2015, WX2016, WX2017, WX2018, WX2019,
         WX2020, WX2021, WX2022, WX2023, WX2024, WX2025, WX2026, WX2027,
         WX2029, WX2030, WX2031, WX2032, WX2033, WX2034, WX2035, WX2036,
         WX2037, WX2038, WX2039, WX2040, WX2041, WX2042, WX2043, WX2044,
         WX2045, WX2046, WX2047, WX2048, WX2049, WX2050, WX2051, WX2052,
         WX2053, WX2054, WX2055, WX2056, WX2057, WX2058, WX2059, WX2060,
         WX2061, WX2062, WX2063, WX2065, WX2066, WX2067, WX2068, WX2069,
         WX2070, WX2071, WX2072, WX2073, WX2074, WX2075, WX2076, WX2077,
         WX2078, WX2079, WX2080, WX2081, WX2082, WX2083, WX2084, WX2085,
         WX2086, WX2087, WX2088, WX2089, WX2090, WX2091, WX2092, WX2093,
         WX2094, WX2095, WX2096, WX2097, WX2098, WX2099, WX2101, WX2102,
         WX2103, WX2104, WX2105, WX2106, WX2107, WX2108, WX2109, WX2110,
         WX2111, WX2112, WX2113, WX2114, WX2115, WX2116, WX2117, WX2118,
         WX2119, WX2120, WX2121, WX2122, WX2123, WX2124, WX2125, WX2126,
         WX2127, WX2128, WX2129, WX2130, WX2131, WX2132, WX2133, WX2134,
         WX2135, WX2137, WX2138, WX2139, WX2140, WX2141, WX2142, WX2143,
         WX2144, WX2145, WX2146, WX2147, WX2148, WX2149, WX2150, WX2151,
         WX2152, WX2153, WX2154, WX2155, WX2156, WX2157, WX2158, WX2159,
         WX2160, WX2161, WX2162, WX2163, WX2164, WX2165, WX2166, WX2167,
         WX2168, WX2169, WX2170, WX2171, WX2173, WX2174, WX2175, WX2176,
         WX2177, WX2178, WX2179, WX2180, WX2181, WX2182, WX2183, WX2184,
         WX2185, WX2186, WX2187, WX2188, WX2189, WX2190, WX2191, WX2192,
         WX2557, DFF_352_n1, WX2559, DFF_353_n1, WX2561, DFF_354_n1, WX2563,
         DFF_355_n1, WX2565, DFF_356_n1, WX2567, DFF_357_n1, WX2569,
         DFF_358_n1, WX2571, WX2573, DFF_360_n1, WX2575, DFF_361_n1, WX2577,
         DFF_362_n1, WX2579, DFF_363_n1, WX2581, DFF_364_n1, WX2583,
         DFF_365_n1, WX2585, DFF_366_n1, WX2587, DFF_367_n1, WX2589,
         DFF_368_n1, WX2591, DFF_369_n1, WX2593, DFF_370_n1, WX2595,
         DFF_371_n1, WX2597, DFF_372_n1, WX2599, DFF_373_n1, WX2601,
         DFF_374_n1, WX2603, DFF_375_n1, WX2605, DFF_376_n1, WX2607, WX2609,
         DFF_378_n1, WX2611, DFF_379_n1, WX2613, DFF_380_n1, WX2615,
         DFF_381_n1, WX2617, DFF_382_n1, WX2619, DFF_383_n1, WX3071, n8644,
         n8643, n8642, n8641, n8640, n8639, n8638, n8637, n8636, n8635, n8632,
         n8631, n8630, n8629, n8628, n8627, n8626, n8625, n8624, n8623, n8622,
         n8621, n8620, n8619, n8618, n8617, n8616, n8613, WX3132, n8612,
         WX3230, n8611, WX3232, n8610, WX3234, n8609, WX3236, n8608, WX3238,
         n8607, WX3240, n8606, WX3242, n8605, WX3244, n8604, WX3246, n8603,
         WX3248, n8602, WX3250, n8601, WX3252, n8600, WX3254, n8599, WX3256,
         n8598, WX3258, n8597, WX3260, WX3262, WX3263, WX3264, WX3265, WX3266,
         WX3267, WX3268, WX3269, WX3270, WX3271, WX3272, WX3273, WX3274,
         WX3275, WX3276, WX3277, WX3278, WX3279, WX3280, WX3281, WX3282,
         WX3283, WX3284, WX3285, WX3286, WX3287, WX3288, WX3289, WX3290,
         WX3291, WX3292, WX3293, WX3294, WX3295, WX3296, WX3298, WX3299,
         WX3300, WX3301, WX3302, WX3303, WX3304, WX3305, WX3306, WX3307,
         WX3308, WX3309, WX3310, WX3311, WX3312, WX3313, WX3314, WX3315,
         WX3316, WX3317, WX3318, WX3319, WX3320, WX3321, WX3322, WX3323,
         WX3324, WX3325, WX3326, WX3327, WX3328, WX3329, WX3330, WX3331,
         WX3332, WX3334, WX3335, WX3336, WX3337, WX3338, WX3339, WX3340,
         WX3341, WX3342, WX3343, WX3344, WX3345, WX3346, WX3347, WX3348,
         WX3349, WX3350, WX3351, WX3352, WX3353, WX3354, WX3355, WX3356,
         WX3357, WX3358, WX3359, WX3360, WX3361, WX3362, WX3363, WX3364,
         WX3365, WX3366, WX3367, WX3368, WX3370, WX3371, WX3372, WX3373,
         WX3374, WX3375, WX3376, WX3377, WX3378, WX3379, WX3380, WX3381,
         WX3382, WX3383, WX3384, WX3385, WX3386, WX3387, WX3388, WX3389,
         WX3390, WX3391, WX3392, WX3393, WX3394, WX3395, WX3396, WX3397,
         WX3398, WX3399, WX3400, WX3401, WX3402, WX3403, WX3404, WX3406,
         WX3407, WX3408, WX3409, WX3410, WX3411, WX3412, WX3413, WX3414,
         WX3415, WX3416, WX3417, WX3418, WX3419, WX3420, WX3421, WX3422,
         WX3423, WX3424, WX3425, WX3426, WX3427, WX3428, WX3429, WX3430,
         WX3431, WX3432, WX3433, WX3434, WX3435, WX3436, WX3437, WX3438,
         WX3440, WX3441, WX3442, WX3443, WX3444, WX3445, WX3446, WX3447,
         WX3448, WX3449, WX3450, WX3451, WX3452, WX3453, WX3454, WX3455,
         WX3456, WX3457, WX3458, WX3459, WX3460, WX3461, WX3462, WX3463,
         WX3464, WX3465, WX3466, WX3467, WX3468, WX3469, WX3470, WX3471,
         WX3472, WX3474, WX3475, WX3476, WX3477, WX3478, WX3479, WX3480,
         WX3481, WX3482, WX3483, WX3484, WX3485, WX3850, DFF_544_n1, WX3852,
         DFF_545_n1, WX3854, DFF_546_n1, WX3856, DFF_547_n1, WX3858,
         DFF_548_n1, WX3860, DFF_549_n1, WX3862, DFF_550_n1, WX3864,
         DFF_551_n1, WX3866, DFF_552_n1, WX3868, DFF_553_n1, WX3870, WX3872,
         DFF_555_n1, WX3874, DFF_556_n1, WX3876, DFF_557_n1, WX3878,
         DFF_558_n1, WX3880, DFF_559_n1, WX3882, DFF_560_n1, WX3884,
         DFF_561_n1, WX3886, DFF_562_n1, WX3888, DFF_563_n1, WX3890,
         DFF_564_n1, WX3892, DFF_565_n1, WX3894, DFF_566_n1, WX3896,
         DFF_567_n1, WX3898, DFF_568_n1, WX3900, DFF_569_n1, WX3902,
         DFF_570_n1, WX3904, WX3906, DFF_572_n1, WX3908, DFF_573_n1, WX3910,
         DFF_574_n1, WX3912, DFF_575_n1, WX4364, n8586, n8585, n8584, n8583,
         n8582, n8581, n8580, n8579, n8578, n8577, n8576, n8573, n8572, n8571,
         n8570, n8569, n8568, n8567, n8566, n8565, n8564, n8563, n8562, n8561,
         n8560, n8559, n8558, n8555, WX4425, n8554, WX4523, n8553, WX4525,
         n8552, WX4527, n8551, WX4529, n8550, WX4531, n8549, WX4533, n8548,
         WX4535, n8547, WX4537, n8546, WX4539, n8545, WX4541, n8544, WX4543,
         n8543, WX4545, n8542, WX4547, n8541, WX4549, n8540, WX4551, WX4553,
         n8537, WX4555, WX4556, WX4557, WX4558, WX4559, WX4560, WX4561, WX4562,
         WX4563, WX4564, WX4565, WX4566, WX4567, WX4568, WX4569, WX4570,
         WX4571, WX4572, WX4573, WX4574, WX4575, WX4576, WX4577, WX4578,
         WX4579, WX4580, WX4581, WX4582, WX4583, WX4584, WX4585, WX4587,
         WX4588, WX4589, WX4590, WX4591, WX4592, WX4593, WX4594, WX4595,
         WX4596, WX4597, WX4598, WX4599, WX4600, WX4601, WX4602, WX4603,
         WX4604, WX4605, WX4606, WX4607, WX4608, WX4609, WX4610, WX4611,
         WX4612, WX4613, WX4614, WX4615, WX4616, WX4617, WX4618, WX4619,
         WX4621, WX4622, WX4623, WX4624, WX4625, WX4626, WX4627, WX4628,
         WX4629, WX4630, WX4631, WX4632, WX4633, WX4634, WX4635, WX4636,
         WX4637, WX4638, WX4639, WX4640, WX4641, WX4642, WX4643, WX4644,
         WX4645, WX4646, WX4647, WX4648, WX4649, WX4650, WX4651, WX4652,
         WX4653, WX4655, WX4656, WX4657, WX4658, WX4659, WX4660, WX4661,
         WX4662, WX4663, WX4664, WX4665, WX4666, WX4667, WX4668, WX4669,
         WX4670, WX4671, WX4672, WX4673, WX4674, WX4675, WX4676, WX4677,
         WX4678, WX4679, WX4680, WX4681, WX4682, WX4683, WX4684, WX4685,
         WX4686, WX4687, WX4689, WX4690, WX4691, WX4692, WX4693, WX4694,
         WX4695, WX4696, WX4697, WX4698, WX4699, WX4700, WX4701, WX4702,
         WX4703, WX4704, WX4705, WX4706, WX4707, WX4708, WX4709, WX4710,
         WX4711, WX4712, WX4713, WX4714, WX4715, WX4716, WX4717, WX4718,
         WX4719, WX4720, WX4721, WX4723, WX4724, WX4725, WX4726, WX4727,
         WX4728, WX4729, WX4730, WX4731, WX4732, WX4733, WX4734, WX4735,
         WX4736, WX4737, WX4738, WX4739, WX4740, WX4741, WX4742, WX4743,
         WX4744, WX4745, WX4746, WX4747, WX4748, WX4749, WX4750, WX4751,
         WX4752, WX4753, WX4754, WX4755, WX4757, WX4758, WX4759, WX4760,
         WX4761, WX4762, WX4763, WX4764, WX4765, WX4766, WX4767, WX4768,
         WX4769, WX4770, WX4771, WX4772, WX4773, WX4774, WX4775, WX4776,
         WX4777, WX4778, WX5143, DFF_736_n1, WX5145, DFF_737_n1, WX5147,
         DFF_738_n1, WX5149, DFF_739_n1, WX5151, DFF_740_n1, WX5153, WX5155,
         DFF_742_n1, WX5157, DFF_743_n1, WX5159, DFF_744_n1, WX5161,
         DFF_745_n1, WX5163, DFF_746_n1, WX5165, DFF_747_n1, WX5167,
         DFF_748_n1, WX5169, DFF_749_n1, WX5171, DFF_750_n1, WX5173,
         DFF_751_n1, WX5175, DFF_752_n1, WX5177, DFF_753_n1, WX5179,
         DFF_754_n1, WX5181, DFF_755_n1, WX5183, DFF_756_n1, WX5185,
         DFF_757_n1, WX5187, WX5189, DFF_759_n1, WX5191, DFF_760_n1, WX5193,
         DFF_761_n1, WX5195, DFF_762_n1, WX5197, DFF_763_n1, WX5199,
         DFF_764_n1, WX5201, DFF_765_n1, WX5203, DFF_766_n1, WX5205,
         DFF_767_n1, WX5657, n8528, n8527, n8526, n8525, n8524, n8523, n8520,
         n8519, n8518, n8517, n8516, n8515, n8514, n8513, n8512, n8511, n8510,
         n8509, n8508, n8507, n8506, n8505, n8502, n8501, n8500, n8499, n8498,
         n8497, WX5718, n8496, WX5816, n8495, WX5818, n8494, WX5820, n8493,
         WX5822, n8492, WX5824, n8491, WX5826, n8490, WX5828, n8489, WX5830,
         n8488, WX5832, n8487, WX5834, WX5836, n8484, WX5838, n8483, WX5840,
         n8482, WX5842, n8481, WX5844, n8480, WX5846, n8479, WX5848, WX5849,
         WX5850, WX5851, WX5852, WX5853, WX5854, WX5855, WX5856, WX5857,
         WX5858, WX5859, WX5860, WX5861, WX5862, WX5863, WX5864, WX5865,
         WX5866, WX5867, WX5868, WX5870, WX5871, WX5872, WX5873, WX5874,
         WX5875, WX5876, WX5877, WX5878, WX5879, WX5880, WX5881, WX5882,
         WX5883, WX5884, WX5885, WX5886, WX5887, WX5888, WX5889, WX5890,
         WX5891, WX5892, WX5893, WX5894, WX5895, WX5896, WX5897, WX5898,
         WX5899, WX5900, WX5901, WX5902, WX5904, WX5905, WX5906, WX5907,
         WX5908, WX5909, WX5910, WX5911, WX5912, WX5913, WX5914, WX5915,
         WX5916, WX5917, WX5918, WX5919, WX5920, WX5921, WX5922, WX5923,
         WX5924, WX5925, WX5926, WX5927, WX5928, WX5929, WX5930, WX5931,
         WX5932, WX5933, WX5934, WX5935, WX5936, WX5938, WX5939, WX5940,
         WX5941, WX5942, WX5943, WX5944, WX5945, WX5946, WX5947, WX5948,
         WX5949, WX5950, WX5951, WX5952, WX5953, WX5954, WX5955, WX5956,
         WX5957, WX5958, WX5959, WX5960, WX5961, WX5962, WX5963, WX5964,
         WX5965, WX5966, WX5967, WX5968, WX5969, WX5970, WX5972, WX5973,
         WX5974, WX5975, WX5976, WX5977, WX5978, WX5979, WX5980, WX5981,
         WX5982, WX5983, WX5984, WX5985, WX5986, WX5987, WX5988, WX5989,
         WX5990, WX5991, WX5992, WX5993, WX5994, WX5995, WX5996, WX5997,
         WX5998, WX5999, WX6000, WX6001, WX6002, WX6003, WX6004, WX6006,
         WX6007, WX6008, WX6009, WX6010, WX6011, WX6012, WX6013, WX6014,
         WX6015, WX6016, WX6017, WX6018, WX6019, WX6020, WX6021, WX6022,
         WX6023, WX6024, WX6025, WX6026, WX6027, WX6028, WX6029, WX6030,
         WX6031, WX6032, WX6033, WX6034, WX6035, WX6036, WX6037, WX6038,
         WX6040, WX6041, WX6042, WX6043, WX6044, WX6045, WX6046, WX6047,
         WX6048, WX6049, WX6050, WX6051, WX6052, WX6053, WX6054, WX6055,
         WX6056, WX6057, WX6058, WX6059, WX6060, WX6061, WX6062, WX6063,
         WX6064, WX6065, WX6066, WX6067, WX6068, WX6069, WX6070, WX6071,
         WX6436, WX6438, DFF_929_n1, WX6440, DFF_930_n1, WX6442, DFF_931_n1,
         WX6444, DFF_932_n1, WX6446, DFF_933_n1, WX6448, DFF_934_n1, WX6450,
         DFF_935_n1, WX6452, DFF_936_n1, WX6454, DFF_937_n1, WX6456,
         DFF_938_n1, WX6458, DFF_939_n1, WX6460, DFF_940_n1, WX6462,
         DFF_941_n1, WX6464, DFF_942_n1, WX6466, DFF_943_n1, WX6468,
         DFF_944_n1, WX6470, WX6472, DFF_946_n1, WX6474, DFF_947_n1, WX6476,
         DFF_948_n1, WX6478, DFF_949_n1, WX6480, DFF_950_n1, WX6482,
         DFF_951_n1, WX6484, DFF_952_n1, WX6486, DFF_953_n1, WX6488,
         DFF_954_n1, WX6490, DFF_955_n1, WX6492, DFF_956_n1, WX6494,
         DFF_957_n1, WX6496, DFF_958_n1, WX6498, DFF_959_n1, WX6950, n8470,
         n8467, n8466, n8465, n8464, n8463, n8462, n8461, n8460, n8459, n8458,
         n8457, n8456, n8455, n8454, n8453, n8452, n8449, n8448, n8447, n8446,
         n8445, n8444, n8443, n8442, n8441, n8440, n8439, WX7011, n8438,
         WX7109, n8437, WX7111, n8436, WX7113, n8435, WX7115, n8434, WX7117,
         WX7119, n8431, WX7121, n8430, WX7123, n8429, WX7125, n8428, WX7127,
         n8427, WX7129, n8426, WX7131, n8425, WX7133, n8424, WX7135, n8423,
         WX7137, n8422, WX7139, n8421, WX7141, WX7142, WX7143, WX7144, WX7145,
         WX7146, WX7147, WX7148, WX7149, WX7150, WX7151, WX7153, WX7154,
         WX7155, WX7156, WX7157, WX7158, WX7159, WX7160, WX7161, WX7162,
         WX7163, WX7164, WX7165, WX7166, WX7167, WX7168, WX7169, WX7170,
         WX7171, WX7172, WX7173, WX7174, WX7175, WX7176, WX7177, WX7178,
         WX7179, WX7180, WX7181, WX7182, WX7183, WX7184, WX7185, WX7187,
         WX7188, WX7189, WX7190, WX7191, WX7192, WX7193, WX7194, WX7195,
         WX7196, WX7197, WX7198, WX7199, WX7200, WX7201, WX7202, WX7203,
         WX7204, WX7205, WX7206, WX7207, WX7208, WX7209, WX7210, WX7211,
         WX7212, WX7213, WX7214, WX7215, WX7216, WX7217, WX7218, WX7219,
         WX7221, WX7222, WX7223, WX7224, WX7225, WX7226, WX7227, WX7228,
         WX7229, WX7230, WX7231, WX7232, WX7233, WX7234, WX7235, WX7236,
         WX7237, WX7238, WX7239, WX7240, WX7241, WX7242, WX7243, WX7244,
         WX7245, WX7246, WX7247, WX7248, WX7249, WX7250, WX7251, WX7252,
         WX7253, WX7255, WX7256, WX7257, WX7258, WX7259, WX7260, WX7261,
         WX7262, WX7263, WX7264, WX7265, WX7266, WX7267, WX7268, WX7269,
         WX7270, WX7271, WX7272, WX7273, WX7274, WX7275, WX7276, WX7277,
         WX7278, WX7279, WX7280, WX7281, WX7282, WX7283, WX7284, WX7285,
         WX7286, WX7287, WX7289, WX7290, WX7291, WX7292, WX7293, WX7294,
         WX7295, WX7296, WX7297, WX7298, WX7299, WX7300, WX7301, WX7302,
         WX7303, WX7304, WX7305, WX7306, WX7307, WX7308, WX7309, WX7310,
         WX7311, WX7312, WX7313, WX7314, WX7315, WX7316, WX7317, WX7318,
         WX7319, WX7320, WX7321, WX7323, WX7324, WX7325, WX7326, WX7327,
         WX7328, WX7329, WX7330, WX7331, WX7332, WX7333, WX7334, WX7335,
         WX7336, WX7337, WX7338, WX7339, WX7340, WX7341, WX7342, WX7343,
         WX7344, WX7345, WX7346, WX7347, WX7348, WX7349, WX7350, WX7351,
         WX7352, WX7353, WX7354, WX7355, WX7357, WX7358, WX7359, WX7360,
         WX7361, WX7362, WX7363, WX7364, WX7729, DFF_1120_n1, WX7731,
         DFF_1121_n1, WX7733, DFF_1122_n1, WX7735, DFF_1123_n1, WX7737,
         DFF_1124_n1, WX7739, DFF_1125_n1, WX7741, DFF_1126_n1, WX7743,
         DFF_1127_n1, WX7745, DFF_1128_n1, WX7747, DFF_1129_n1, WX7749,
         DFF_1130_n1, WX7751, DFF_1131_n1, WX7753, WX7755, DFF_1133_n1, WX7757,
         DFF_1134_n1, WX7759, DFF_1135_n1, WX7761, DFF_1136_n1, WX7763,
         DFF_1137_n1, WX7765, DFF_1138_n1, WX7767, DFF_1139_n1, WX7769,
         DFF_1140_n1, WX7771, DFF_1141_n1, WX7773, DFF_1142_n1, WX7775,
         DFF_1143_n1, WX7777, DFF_1144_n1, WX7779, DFF_1145_n1, WX7781,
         DFF_1146_n1, WX7783, DFF_1147_n1, WX7785, DFF_1148_n1, WX7787, WX7789,
         DFF_1150_n1, WX7791, DFF_1151_n1, WX8243, n8411, n8410, n8409, n8408,
         n8407, n8406, n8405, n8404, n8403, n8402, n8401, n8400, n8399, n8396,
         n8395, n8394, n8393, n8392, n8391, n8390, n8389, n8388, n8387, n8386,
         n8385, n8384, n8383, n8382, n8381, WX8304, WX8402, n8378, WX8404,
         n8377, WX8406, n8376, WX8408, n8375, WX8410, n8374, WX8412, n8373,
         WX8414, n8372, WX8416, n8371, WX8418, n8370, WX8420, n8369, WX8422,
         n8368, WX8424, n8367, WX8426, n8366, WX8428, n8365, WX8430, n8364,
         WX8432, n8363, WX8434, WX8436, WX8437, WX8438, WX8439, WX8440, WX8441,
         WX8442, WX8443, WX8444, WX8445, WX8446, WX8447, WX8448, WX8449,
         WX8450, WX8451, WX8452, WX8453, WX8454, WX8455, WX8456, WX8457,
         WX8458, WX8459, WX8460, WX8461, WX8462, WX8463, WX8464, WX8465,
         WX8466, WX8467, WX8468, WX8470, WX8471, WX8472, WX8473, WX8474,
         WX8475, WX8476, WX8477, WX8478, WX8479, WX8480, WX8481, WX8482,
         WX8483, WX8484, WX8485, WX8486, WX8487, WX8488, WX8489, WX8490,
         WX8491, WX8492, WX8493, WX8494, WX8495, WX8496, WX8497, WX8498,
         WX8499, WX8500, WX8501, WX8502, WX8504, WX8505, WX8506, WX8507,
         WX8508, WX8509, WX8510, WX8511, WX8512, WX8513, WX8514, WX8515,
         WX8516, WX8517, WX8518, WX8519, WX8520, WX8521, WX8522, WX8523,
         WX8524, WX8525, WX8526, WX8527, WX8528, WX8529, WX8530, WX8531,
         WX8532, WX8533, WX8534, WX8535, WX8536, WX8538, WX8539, WX8540,
         WX8541, WX8542, WX8543, WX8544, WX8545, WX8546, WX8547, WX8548,
         WX8549, WX8550, WX8551, WX8552, WX8553, WX8554, WX8555, WX8556,
         WX8557, WX8558, WX8559, WX8560, WX8561, WX8562, WX8563, WX8564,
         WX8565, WX8566, WX8567, WX8568, WX8569, WX8570, WX8572, WX8573,
         WX8574, WX8575, WX8576, WX8577, WX8578, WX8579, WX8580, WX8581,
         WX8582, WX8583, WX8584, WX8585, WX8586, WX8587, WX8588, WX8589,
         WX8590, WX8591, WX8592, WX8593, WX8594, WX8595, WX8596, WX8597,
         WX8598, WX8599, WX8600, WX8601, WX8602, WX8603, WX8604, WX8606,
         WX8607, WX8608, WX8609, WX8610, WX8611, WX8612, WX8613, WX8614,
         WX8615, WX8616, WX8617, WX8618, WX8619, WX8620, WX8621, WX8622,
         WX8623, WX8624, WX8625, WX8626, WX8627, WX8628, WX8629, WX8630,
         WX8631, WX8632, WX8633, WX8634, WX8635, WX8636, WX8637, WX8638,
         WX8640, WX8641, WX8642, WX8643, WX8644, WX8645, WX8646, WX8647,
         WX8648, WX8649, WX8650, WX8651, WX8652, WX8653, WX8654, WX8655,
         WX8656, WX8657, WX9022, DFF_1312_n1, WX9024, DFF_1313_n1, WX9026,
         DFF_1314_n1, WX9028, DFF_1315_n1, WX9030, DFF_1316_n1, WX9032,
         DFF_1317_n1, WX9034, DFF_1318_n1, WX9036, WX9038, DFF_1320_n1, WX9040,
         DFF_1321_n1, WX9042, DFF_1322_n1, WX9044, DFF_1323_n1, WX9046,
         DFF_1324_n1, WX9048, DFF_1325_n1, WX9050, DFF_1326_n1, WX9052,
         DFF_1327_n1, WX9054, DFF_1328_n1, WX9056, DFF_1329_n1, WX9058,
         DFF_1330_n1, WX9060, DFF_1331_n1, WX9062, DFF_1332_n1, WX9064,
         DFF_1333_n1, WX9066, DFF_1334_n1, WX9068, DFF_1335_n1, WX9070, WX9072,
         DFF_1337_n1, WX9074, DFF_1338_n1, WX9076, DFF_1339_n1, WX9078,
         DFF_1340_n1, WX9080, DFF_1341_n1, WX9082, DFF_1342_n1, WX9084,
         DFF_1343_n1, WX9536, n8353, n8352, n8351, n8350, n8349, n8348, n8347,
         n8346, n8343, n8342, n8341, n8340, n8339, n8338, n8337, n8336, n8335,
         n8334, n8333, n8332, n8331, n8330, n8329, n8328, n8325, n8324, n8323,
         n8322, WX9597, n8321, WX9695, n8320, WX9697, n8319, WX9699, n8318,
         WX9701, n8317, WX9703, n8316, WX9705, n8315, WX9707, n8314, WX9709,
         n8313, WX9711, n8312, WX9713, n8311, WX9715, n8310, WX9717, WX9719,
         n8307, WX9721, n8306, WX9723, n8305, WX9725, n8304, WX9727, WX9728,
         WX9729, WX9730, WX9731, WX9732, WX9733, WX9734, WX9735, WX9736,
         WX9737, WX9738, WX9739, WX9740, WX9741, WX9742, WX9743, WX9744,
         WX9745, WX9746, WX9747, WX9748, WX9749, WX9750, WX9751, WX9753,
         WX9754, WX9755, WX9756, WX9757, WX9758, WX9759, WX9760, WX9761,
         WX9762, WX9763, WX9764, WX9765, WX9766, WX9767, WX9768, WX9769,
         WX9770, WX9771, WX9772, WX9773, WX9774, WX9775, WX9776, WX9777,
         WX9778, WX9779, WX9780, WX9781, WX9782, WX9783, WX9784, WX9785,
         WX9787, WX9788, WX9789, WX9790, WX9791, WX9792, WX9793, WX9794,
         WX9795, WX9796, WX9797, WX9798, WX9799, WX9800, WX9801, WX9802,
         WX9803, WX9804, WX9805, WX9806, WX9807, WX9808, WX9809, WX9810,
         WX9811, WX9812, WX9813, WX9814, WX9815, WX9816, WX9817, WX9818,
         WX9819, WX9821, WX9822, WX9823, WX9824, WX9825, WX9826, WX9827,
         WX9828, WX9829, WX9830, WX9831, WX9832, WX9833, WX9834, WX9835,
         WX9836, WX9837, WX9838, WX9839, WX9840, WX9841, WX9842, WX9843,
         WX9844, WX9845, WX9846, WX9847, WX9848, WX9849, WX9850, WX9851,
         WX9852, WX9853, WX9855, WX9856, WX9857, WX9858, WX9859, WX9860,
         WX9861, WX9862, WX9863, WX9864, WX9865, WX9866, WX9867, WX9868,
         WX9869, WX9870, WX9871, WX9872, WX9873, WX9874, WX9875, WX9876,
         WX9877, WX9878, WX9879, WX9880, WX9881, WX9882, WX9883, WX9884,
         WX9885, WX9886, WX9887, WX9889, WX9890, WX9891, WX9892, WX9893,
         WX9894, WX9895, WX9896, WX9897, WX9898, WX9899, WX9900, WX9901,
         WX9902, WX9903, WX9904, WX9905, WX9906, WX9907, WX9908, WX9909,
         WX9910, WX9911, WX9912, WX9913, WX9914, WX9915, WX9916, WX9917,
         WX9918, WX9919, WX9920, WX9921, WX9923, WX9924, WX9925, WX9926,
         WX9927, WX9928, WX9929, WX9930, WX9931, WX9932, WX9933, WX9934,
         WX9935, WX9936, WX9937, WX9938, WX9939, WX9940, WX9941, WX9942,
         WX9943, WX9944, WX9945, WX9946, WX9947, WX9948, WX9949, WX9950,
         WX10315, DFF_1504_n1, WX10317, DFF_1505_n1, WX10319, WX10321,
         DFF_1507_n1, WX10323, DFF_1508_n1, WX10325, DFF_1509_n1, WX10327,
         DFF_1510_n1, WX10329, DFF_1511_n1, WX10331, DFF_1512_n1, WX10333,
         DFF_1513_n1, WX10335, DFF_1514_n1, WX10337, DFF_1515_n1, WX10339,
         DFF_1516_n1, WX10341, DFF_1517_n1, WX10343, DFF_1518_n1, WX10345,
         DFF_1519_n1, WX10347, DFF_1520_n1, WX10349, DFF_1521_n1, WX10351,
         DFF_1522_n1, WX10353, WX10355, DFF_1524_n1, WX10357, DFF_1525_n1,
         WX10359, DFF_1526_n1, WX10361, DFF_1527_n1, WX10363, DFF_1528_n1,
         WX10365, DFF_1529_n1, WX10367, DFF_1530_n1, WX10369, DFF_1531_n1,
         WX10371, DFF_1532_n1, WX10373, DFF_1533_n1, WX10375, DFF_1534_n1,
         WX10377, DFF_1535_n1, WX10828, WX10829, WX10830, n8295, WX10832,
         n8294, WX10834, n8293, WX10836, WX10838, n8290, WX10840, n8289,
         WX10842, n8288, WX10844, n8287, WX10846, n8286, WX10848, n8285,
         WX10850, n8284, WX10852, n8283, WX10854, n8282, WX10856, n8281,
         WX10858, n8280, WX10860, n8279, WX10862, n8278, WX10864, n8277,
         WX10866, n8276, WX10868, n8275, WX10870, WX10872, n8272, WX10874,
         n8271, WX10876, n8270, WX10878, n8269, WX10880, n8268, WX10882, n8267,
         WX10884, n8266, WX10886, n8265, WX10888, n8264, WX10890, n8263,
         WX10988, n8262, WX10990, n8261, WX10992, n8260, WX10994, n8259,
         WX10996, n8258, WX10998, n8257, WX11000, WX11002, n8254, WX11004,
         n8253, WX11006, n8252, WX11008, n8251, WX11010, n8250, WX11012, n8249,
         WX11014, n8248, WX11016, n8247, WX11018, n8246, WX11020, WX11021,
         WX11022, WX11023, WX11024, WX11025, WX11026, WX11027, WX11028,
         WX11029, WX11030, WX11031, WX11032, WX11033, WX11034, WX11036,
         WX11037, WX11038, WX11039, WX11040, WX11041, WX11042, WX11043,
         WX11044, WX11045, WX11046, WX11047, WX11048, WX11049, WX11050,
         WX11051, WX11052, WX11053, WX11054, WX11055, WX11056, WX11057,
         WX11058, WX11059, WX11060, WX11061, WX11062, WX11063, WX11064,
         WX11065, WX11066, WX11067, WX11068, WX11070, WX11071, WX11072,
         WX11073, WX11074, WX11075, WX11076, WX11077, WX11078, WX11079,
         WX11080, WX11081, WX11082, WX11083, WX11084, WX11085, WX11086,
         WX11087, WX11088, WX11089, WX11090, WX11091, WX11092, WX11093,
         WX11094, WX11095, WX11096, WX11097, WX11098, WX11099, WX11100,
         WX11101, WX11102, WX11104, WX11105, WX11106, WX11107, WX11108,
         WX11109, WX11110, WX11111, WX11112, WX11113, WX11114, WX11115,
         WX11116, WX11117, WX11118, WX11119, WX11120, WX11121, WX11122,
         WX11123, WX11124, WX11125, WX11126, WX11127, WX11128, WX11129,
         WX11130, WX11131, WX11132, WX11133, WX11134, WX11135, WX11136,
         WX11138, WX11139, WX11140, WX11141, WX11142, WX11143, WX11144,
         WX11145, WX11146, WX11147, WX11148, WX11149, WX11150, WX11151,
         WX11152, WX11153, WX11154, WX11155, WX11156, WX11155_Tj_Payload,
         test_se_Trojan, WX11157, WX11158, WX11159, WX11160, WX11161, WX11162,
         WX11163, WX11164, WX11165, WX11166, WX11167, WX11168, WX11169,
         WX11170, WX11172, WX11173, WX11174, WX11175, WX11176, WX11177,
         WX11178, WX11179, WX11180, WX11181, WX11182, WX11183, WX11184,
         WX11185, WX11186, WX11187, WX11188, WX11189, WX11190, WX11191,
         WX11192, WX11193, WX11194, WX11195, WX11196, WX11197, WX11198,
         WX11199, WX11200, WX11201, WX11202, WX11203, WX11204, WX11206,
         WX11207, WX11208, WX11209, WX11210, WX11211, WX11212, WX11213,
         WX11214, WX11215, WX11216, WX11217, WX11218, WX11219, WX11220,
         WX11221, WX11222, WX11223, WX11224, WX11225, WX11226, WX11227,
         WX11228, WX11229, WX11230, WX11231, WX11232, WX11233, WX11234,
         WX11235, WX11236, WX11237, WX11238, WX11240, WX11241, WX11242,
         WX11243, WX11608, DFF_1696_n1, WX11610, DFF_1697_n1, WX11612,
         DFF_1698_n1, WX11614, DFF_1699_n1, WX11616, DFF_1700_n1, WX11618,
         DFF_1701_n1, WX11620, DFF_1702_n1, WX11622, DFF_1703_n1, WX11624,
         DFF_1704_n1, WX11626, DFF_1705_n1, WX11628, DFF_1706_n1, WX11630,
         DFF_1707_n1, WX11632, DFF_1708_n1, WX11634, DFF_1709_n1, WX11636,
         WX11638, DFF_1711_n1, WX11640, DFF_1712_n1, WX11642, DFF_1713_n1,
         WX11644, DFF_1714_n1, WX11646, DFF_1715_n1, WX11648, DFF_1716_n1,
         WX11650, DFF_1717_n1, WX11652, DFF_1718_n1, WX11654, DFF_1719_n1,
         WX11656, DFF_1720_n1, WX11658, DFF_1721_n1, WX11660, DFF_1722_n1,
         WX11662, DFF_1723_n1, WX11664, DFF_1724_n1, WX11666, DFF_1725_n1,
         WX11668, DFF_1726_n1, WX11670, n2245, n2153, n3278, n2152, Tj_OUT1,
         Tj_OUT2, Tj_OUT3, Tj_OUT4, Tj_OUT1234, Tj_OUT5, Tj_OUT6, Tj_OUT7,
         Tj_OUT8, Tj_OUT5678, test_se_NOT, Tj_Trigger, Trojan_SE, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n225, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3697, n3699, n3701, n3703, n3706, n3709, n3712, n3714, n3716, n3718,
         n3720, n3722, n3724, n3726, n3729, n3732, n3734, n3736, n3738, n3740,
         n3742, n3744, n3746, n3748, n3750, n3752, n3754, n3756, n3758, n3760,
         n3762, n3764, n3766, n3768, n3770, n3772, n3774, n3776, n3779, n3782,
         n3785, n3787, n3789, n3791, n3793, n3795, n3798, n3801, n3804, n3806,
         n3808, n3810, n3812, n3814, n3817, n3820, n3823, n3825, n3827, n3829,
         n3831, n3833, n3835, n3837, n3839, n3841, n3844, n3846, n3848, n3850,
         n3852, n3854, n3856, n3858, n3860, n3862, n3864, n3866, n3869, n3872,
         n3874, n3876, n3878, n3880, n3882, n3884, n3886, n3889, n3891, n3893,
         n3896, n3898, n3900, n3903, n3905, n3907, n3910, n3912, n3914, n3916,
         n3918, n3920, n3922, n3924, n3926, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8255, n8256, n8273,
         n8274, n8291, n8292, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8308, n8309, n8326, n8327, n8344, n8345, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8379, n8380, n8397, n8398,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8432,
         n8433, n8450, n8451, n8468, n8469, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8485, n8486, n8503, n8504, n8521, n8522, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8538, n8539, n8556,
         n8557, n8574, n8575, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8614, n8615, n8633, n8634, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8659, n8660, n8678, n8679, n8697,
         n8698, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, U3558_n1,
         U3871_n1, U3991_n1, U5716_n1, U5717_n1, U5718_n1, U5719_n1, U5720_n1,
         U5721_n1, U5722_n1, U5723_n1, U5724_n1, U5725_n1, U5726_n1, U5727_n1,
         U5728_n1, U5729_n1, U5730_n1, U5731_n1, U5732_n1, U5733_n1, U5734_n1,
         U5735_n1, U5736_n1, U5737_n1, U5738_n1, U5739_n1, U5740_n1, U5741_n1,
         U5742_n1, U5743_n1, U5744_n1, U5745_n1, U5746_n1, U5747_n1, U5748_n1,
         U5749_n1, U5750_n1, U5751_n1, U5752_n1, U5753_n1, U5754_n1, U5755_n1,
         U5756_n1, U5757_n1, U5758_n1, U5759_n1, U5760_n1, U5761_n1, U5762_n1,
         U5763_n1, U5764_n1, U5765_n1, U5766_n1, U5767_n1, U5768_n1, U5769_n1,
         U5770_n1, U5771_n1, U5772_n1, U5773_n1, U5774_n1, U5775_n1, U5776_n1,
         U5777_n1, U5778_n1, U5779_n1, U5780_n1, U5781_n1, U5782_n1, U5783_n1,
         U5784_n1, U5785_n1, U5786_n1, U5787_n1, U5788_n1, U5789_n1, U5790_n1,
         U5791_n1, U5792_n1, U5793_n1, U5794_n1, U5795_n1, U5796_n1, U5797_n1,
         U5798_n1, U5799_n1, U5800_n1, U5801_n1, U5802_n1, U5803_n1, U5804_n1,
         U5805_n1, U5806_n1, U5807_n1, U5808_n1, U5809_n1, U5810_n1, U5811_n1,
         U5812_n1, U5813_n1, U5814_n1, U5815_n1, U5816_n1, U5817_n1, U5818_n1,
         U5819_n1, U5820_n1, U5821_n1, U5822_n1, U5823_n1, U5824_n1, U5825_n1,
         U5826_n1, U5827_n1, U5828_n1, U5829_n1, U5830_n1, U5831_n1, U5832_n1,
         U5833_n1, U5834_n1, U5835_n1, U5836_n1, U5837_n1, U5838_n1, U5839_n1,
         U5840_n1, U5841_n1, U5842_n1, U5843_n1, U5844_n1, U5845_n1, U5846_n1,
         U5847_n1, U5848_n1, U5849_n1, U5850_n1, U5851_n1, U5852_n1, U5853_n1,
         U5854_n1, U5855_n1, U5856_n1, U5857_n1, U5858_n1, U5859_n1, U5860_n1,
         U5861_n1, U5862_n1, U5863_n1, U5864_n1, U5865_n1, U5866_n1, U5867_n1,
         U5868_n1, U5869_n1, U5870_n1, U5871_n1, U5872_n1, U5873_n1, U5874_n1,
         U5875_n1, U5876_n1, U5877_n1, U5878_n1, U5879_n1, U5880_n1, U5881_n1,
         U5882_n1, U5883_n1, U5884_n1, U5885_n1, U5886_n1, U5887_n1, U5888_n1,
         U5889_n1, U5890_n1, U5891_n1, U5892_n1, U5893_n1, U5894_n1, U5895_n1,
         U5896_n1, U5897_n1, U5898_n1, U5899_n1, U5900_n1, U5901_n1, U5902_n1,
         U5903_n1, U5904_n1, U5905_n1, U5906_n1, U5907_n1, U5908_n1, U5909_n1,
         U5910_n1, U5911_n1, U5912_n1, U5913_n1, U5914_n1, U5915_n1, U5916_n1,
         U5917_n1, U5918_n1, U5919_n1, U5920_n1, U5921_n1, U5922_n1, U5923_n1,
         U5924_n1, U5925_n1, U5926_n1, U5927_n1, U5928_n1, U5929_n1, U5930_n1,
         U5931_n1, U5932_n1, U5933_n1, U5934_n1, U5935_n1, U5936_n1, U5937_n1,
         U5938_n1, U5939_n1, U5940_n1, U5941_n1, U5942_n1, U5943_n1, U5944_n1,
         U5945_n1, U5946_n1, U5947_n1, U5948_n1, U5949_n1, U5950_n1, U5951_n1,
         U5952_n1, U5953_n1, U5954_n1, U5955_n1, U5956_n1, U5957_n1, U5958_n1,
         U5959_n1, U5960_n1, U5961_n1, U5962_n1, U5963_n1, U5964_n1, U5965_n1,
         U5966_n1, U5967_n1, U5968_n1, U5969_n1, U5970_n1, U5971_n1, U5972_n1,
         U5973_n1, U5974_n1, U5975_n1, U5976_n1, U5977_n1, U5978_n1, U5979_n1,
         U5980_n1, U5981_n1, U5982_n1, U5983_n1, U5984_n1, U5985_n1, U5986_n1,
         U5987_n1, U5988_n1, U5989_n1, U5990_n1, U5991_n1, U5992_n1, U5993_n1,
         U5994_n1, U5995_n1, U5996_n1, U5997_n1, U5998_n1, U5999_n1, U6000_n1,
         U6001_n1, U6002_n1, U6003_n1, U6004_n1, U6005_n1, U6006_n1, U6007_n1,
         U6008_n1, U6009_n1, U6010_n1, U6011_n1, U6012_n1, U6013_n1, U6014_n1,
         U6015_n1, U6016_n1, U6017_n1, U6018_n1, U6019_n1, U6020_n1, U6021_n1,
         U6022_n1, U6023_n1, U6024_n1, U6025_n1, U6026_n1, U6027_n1, U6028_n1,
         U6029_n1, U6030_n1, U6031_n1, U6032_n1, U6033_n1, U6034_n1, U6035_n1,
         U6036_n1, U6037_n1, U6038_n1, U6039_n1, U6040_n1, U6041_n1, U6042_n1,
         U6043_n1, U6044_n1, U6045_n1, U6046_n1, U6047_n1, U6048_n1, U6049_n1,
         U6050_n1, U6051_n1, U6052_n1, U6053_n1, U6054_n1, U6055_n1, U6056_n1,
         U6057_n1, U6058_n1, U6059_n1, U6060_n1, U6061_n1, U6062_n1, U6063_n1,
         U6064_n1, U6065_n1, U6066_n1, U6067_n1, U6068_n1, U6069_n1, U6070_n1,
         U6071_n1, U6072_n1, U6073_n1, U6074_n1, U6075_n1, U6076_n1, U6077_n1,
         U6078_n1, U6079_n1, U6080_n1, U6081_n1, U6082_n1, U6083_n1, U6084_n1,
         U6085_n1, U6086_n1, U6087_n1, U6088_n1, U6089_n1, U6090_n1, U6091_n1,
         U6092_n1, U6093_n1, U6094_n1, U6095_n1, U6096_n1, U6097_n1, U6098_n1,
         U6099_n1, U6100_n1, U6101_n1, U6102_n1, U6103_n1, U6104_n1, U6105_n1,
         U6106_n1, U6107_n1, U6108_n1, U6109_n1, U6110_n1, U6111_n1, U6112_n1,
         U6113_n1, U6114_n1, U6115_n1, U6116_n1, U6117_n1, U6118_n1, U6119_n1,
         U6120_n1, U6121_n1, U6122_n1, U6123_n1, U6124_n1, U6125_n1, U6126_n1,
         U6127_n1, U6128_n1, U6129_n1, U6130_n1, U6131_n1, U6132_n1, U6133_n1,
         U6134_n1, U6135_n1, U6136_n1, U6137_n1, U6138_n1, U6139_n1, U6140_n1,
         U6141_n1, U6142_n1, U6143_n1, U6144_n1, U6145_n1, U6146_n1, U6147_n1,
         U6148_n1, U6149_n1, U6150_n1, U6151_n1, U6152_n1, U6153_n1, U6154_n1,
         U6155_n1, U6156_n1, U6157_n1, U6158_n1, U6159_n1, U6160_n1, U6161_n1,
         U6162_n1, U6163_n1, U6164_n1, U6165_n1, U6166_n1, U6167_n1, U6168_n1,
         U6169_n1, U6170_n1, U6171_n1, U6172_n1, U6173_n1, U6174_n1, U6175_n1,
         U6176_n1, U6177_n1, U6178_n1, U6179_n1, U6180_n1, U6181_n1, U6182_n1,
         U6183_n1, U6184_n1, U6185_n1, U6186_n1, U6187_n1, U6188_n1, U6189_n1,
         U6190_n1, U6191_n1, U6192_n1, U6193_n1, U6194_n1, U6195_n1, U6196_n1,
         U6197_n1, U6198_n1, U6199_n1, U6200_n1, U6201_n1, U6202_n1, U6203_n1,
         U6204_n1, U6205_n1, U6206_n1, U6207_n1, U6208_n1, U6209_n1, U6210_n1,
         U6211_n1, U6212_n1, U6213_n1, U6214_n1, U6215_n1, U6216_n1, U6217_n1,
         U6218_n1, U6219_n1, U6220_n1, U6221_n1, U6222_n1, U6223_n1, U6224_n1,
         U6225_n1, U6226_n1, U6227_n1, U6228_n1, U6229_n1, U6230_n1, U6231_n1,
         U6232_n1, U6233_n1, U6234_n1, U6235_n1, U6236_n1, U6237_n1, U6238_n1,
         U6239_n1, U6240_n1, U6241_n1, U6242_n1, U6243_n1, U6244_n1, U6245_n1,
         U6246_n1, U6247_n1, U6248_n1, U6249_n1, U6250_n1, U6251_n1, U6252_n1,
         U6253_n1, U6254_n1, U6255_n1, U6256_n1, U6257_n1, U6258_n1, U6259_n1,
         U6260_n1, U6261_n1, U6262_n1, U6263_n1, U6264_n1, U6265_n1, U6266_n1,
         U6267_n1, U6268_n1, U6269_n1, U6270_n1, U6271_n1, U6272_n1, U6273_n1,
         U6274_n1, U6275_n1, U6276_n1, U6277_n1, U6278_n1, U6279_n1, U6280_n1,
         U6281_n1, U6282_n1, U6283_n1, U6284_n1, U6285_n1, U6286_n1, U6287_n1,
         U6288_n1, U6289_n1, U6290_n1, U6291_n1, U6292_n1, U6293_n1, U6294_n1,
         U6295_n1, U6296_n1, U6297_n1, U6298_n1, U6299_n1, U6300_n1, U6301_n1,
         U6302_n1, U6303_n1, U6304_n1, U6305_n1, U6306_n1, U6307_n1, U6308_n1,
         U6309_n1, U6310_n1, U6311_n1, U6312_n1, U6313_n1, U6314_n1, U6315_n1,
         U6316_n1, U6317_n1, U6318_n1, U6319_n1, U6320_n1, U6321_n1, U6322_n1,
         U6323_n1, U6324_n1, U6325_n1, U6326_n1, U6327_n1, U6328_n1, U6329_n1,
         U6330_n1, U6331_n1, U6332_n1, U6333_n1, U6334_n1, U6335_n1, U6336_n1,
         U6337_n1, U6338_n1, U6339_n1, U6340_n1, U6341_n1, U6342_n1, U6343_n1,
         U6344_n1, U6345_n1, U6346_n1, U6347_n1, U6348_n1, U6349_n1, U6350_n1,
         U6351_n1, U6352_n1, U6353_n1, U6354_n1, U6355_n1, U6356_n1, U6357_n1,
         U6358_n1, U6359_n1, U6360_n1, U6361_n1, U6362_n1, U6363_n1, U6364_n1,
         U6365_n1, U6366_n1, U6367_n1, U6368_n1, U6369_n1, U6370_n1, U6371_n1,
         U6372_n1, U6373_n1, U6374_n1, U6375_n1, U6376_n1, U6377_n1, U6378_n1,
         U6379_n1, U6380_n1, U6381_n1, U6382_n1, U6383_n1, U6384_n1, U6385_n1,
         U6386_n1, U6387_n1, U6388_n1, U6389_n1, U6390_n1, U6391_n1, U6392_n1,
         U6393_n1, U6394_n1, U6395_n1, U6396_n1, U6397_n1, U6398_n1, U6399_n1,
         U6400_n1, U6401_n1, U6402_n1, U6403_n1, U6404_n1, U6405_n1, U6406_n1,
         U6407_n1, U6408_n1, U6409_n1, U6410_n1, U6411_n1, U6412_n1, U6413_n1,
         U6414_n1, U6415_n1, U6416_n1, U6417_n1, U6418_n1, U6419_n1, U6420_n1,
         U6421_n1, U6422_n1, U6423_n1, U6424_n1, U6425_n1, U6426_n1, U6427_n1,
         U6428_n1, U6429_n1, U6430_n1, U6431_n1, U6432_n1, U6433_n1, U6434_n1,
         U6435_n1, U6436_n1, U6437_n1, U6438_n1, U6439_n1, U6440_n1, U6441_n1,
         U6442_n1, U6443_n1, U6444_n1, U6445_n1, U6446_n1, U6447_n1, U6448_n1,
         U6449_n1, U6450_n1, U6451_n1, U6452_n1, U6453_n1, U6454_n1, U6455_n1,
         U6456_n1, U6457_n1, U6458_n1, U6459_n1, U6460_n1, U6461_n1, U6462_n1,
         U6463_n1, U6464_n1, U6465_n1, U6466_n1, U6467_n1, U6468_n1, U6469_n1,
         U6470_n1, U6471_n1, U6472_n1, U6473_n1, U6474_n1, U6475_n1, U6476_n1,
         U6477_n1, U6478_n1, U6479_n1, U6480_n1, U6481_n1, U6482_n1;
  assign CRC_OUT_9_1 = test_so9;
  assign CRC_OUT_9_19 = test_so10;
  assign CRC_OUT_8_7 = test_so20;
  assign CRC_OUT_8_25 = test_so21;
  assign CRC_OUT_7_10 = test_so31;
  assign CRC_OUT_7_27 = test_so32;
  assign CRC_OUT_6_5 = test_so42;
  assign CRC_OUT_6_22 = test_so43;
  assign CRC_OUT_5_0 = test_so53;
  assign CRC_OUT_5_17 = test_so54;
  assign CRC_OUT_4_12 = test_so65;
  assign CRC_OUT_4_29 = test_so66;
  assign CRC_OUT_3_7 = test_so76;
  assign CRC_OUT_3_24 = test_so77;
  assign CRC_OUT_2_2 = test_so87;
  assign CRC_OUT_2_19 = test_so88;
  assign CRC_OUT_1_14 = test_so99;
  assign CRC_OUT_1_31 = test_so100;

  SDFFX1 DFF_0_Q_reg ( .D(WX484), .SI(test_si1), .SE(n4627), .CLK(n4946), .Q(
        WX485), .QN(n3930) );
  SDFFX1 DFF_1_Q_reg ( .D(WX486), .SI(WX485), .SE(n4622), .CLK(n4948), .Q(
        WX487) );
  SDFFX1 DFF_2_Q_reg ( .D(WX488), .SI(WX487), .SE(n4622), .CLK(n4948), .Q(
        WX489) );
  SDFFX1 DFF_3_Q_reg ( .D(WX490), .SI(WX489), .SE(n4622), .CLK(n4948), .Q(
        WX491) );
  SDFFX1 DFF_4_Q_reg ( .D(WX492), .SI(WX491), .SE(n4622), .CLK(n4948), .Q(
        WX493) );
  SDFFX1 DFF_5_Q_reg ( .D(WX494), .SI(WX493), .SE(n4623), .CLK(n4948), .Q(
        WX495) );
  SDFFX1 DFF_6_Q_reg ( .D(WX496), .SI(WX495), .SE(n4623), .CLK(n4948), .Q(
        WX497) );
  SDFFX1 DFF_7_Q_reg ( .D(WX498), .SI(WX497), .SE(n4623), .CLK(n4948), .Q(
        WX499) );
  SDFFX1 DFF_8_Q_reg ( .D(WX500), .SI(WX499), .SE(n4623), .CLK(n4948), .Q(
        WX501) );
  SDFFX1 DFF_9_Q_reg ( .D(WX502), .SI(WX501), .SE(n4623), .CLK(n4947), .Q(
        WX503) );
  SDFFX1 DFF_10_Q_reg ( .D(WX504), .SI(WX503), .SE(n4623), .CLK(n4947), .Q(
        WX505) );
  SDFFX1 DFF_11_Q_reg ( .D(WX506), .SI(WX505), .SE(n4624), .CLK(n4947), .Q(
        WX507) );
  SDFFX1 DFF_12_Q_reg ( .D(WX508), .SI(WX507), .SE(n4624), .CLK(n4947), .Q(
        WX509) );
  SDFFX1 DFF_13_Q_reg ( .D(WX510), .SI(WX509), .SE(n4624), .CLK(n4947), .Q(
        WX511) );
  SDFFX1 DFF_14_Q_reg ( .D(WX512), .SI(WX511), .SE(n4624), .CLK(n4947), .Q(
        WX513) );
  SDFFX1 DFF_15_Q_reg ( .D(WX514), .SI(WX513), .SE(n4624), .CLK(n4947), .Q(
        WX515) );
  SDFFX1 DFF_16_Q_reg ( .D(WX516), .SI(WX515), .SE(n4624), .CLK(n4947), .Q(
        WX517) );
  SDFFX1 DFF_17_Q_reg ( .D(WX518), .SI(WX517), .SE(n4625), .CLK(n4947), .Q(
        test_so1) );
  SDFFX1 DFF_18_Q_reg ( .D(WX520), .SI(test_si2), .SE(n4625), .CLK(n4947), .Q(
        WX521) );
  SDFFX1 DFF_19_Q_reg ( .D(WX522), .SI(WX521), .SE(n4625), .CLK(n4947), .Q(
        WX523) );
  SDFFX1 DFF_20_Q_reg ( .D(WX524), .SI(WX523), .SE(n4625), .CLK(n4947), .Q(
        WX525) );
  SDFFX1 DFF_21_Q_reg ( .D(WX526), .SI(WX525), .SE(n4625), .CLK(n4946), .Q(
        WX527) );
  SDFFX1 DFF_22_Q_reg ( .D(WX528), .SI(WX527), .SE(n4625), .CLK(n4946), .Q(
        WX529) );
  SDFFX1 DFF_23_Q_reg ( .D(WX530), .SI(WX529), .SE(n4626), .CLK(n4946), .Q(
        WX531) );
  SDFFX1 DFF_24_Q_reg ( .D(WX532), .SI(WX531), .SE(n4626), .CLK(n4946), .Q(
        WX533) );
  SDFFX1 DFF_25_Q_reg ( .D(WX534), .SI(WX533), .SE(n4626), .CLK(n4946), .Q(
        WX535) );
  SDFFX1 DFF_26_Q_reg ( .D(WX536), .SI(WX535), .SE(n4626), .CLK(n4946), .Q(
        WX537) );
  SDFFX1 DFF_27_Q_reg ( .D(WX538), .SI(WX537), .SE(n4626), .CLK(n4946), .Q(
        WX539) );
  SDFFX1 DFF_28_Q_reg ( .D(WX540), .SI(WX539), .SE(n4626), .CLK(n4946), .Q(
        WX541) );
  SDFFX1 DFF_29_Q_reg ( .D(WX542), .SI(WX541), .SE(n4627), .CLK(n4946), .Q(
        WX543) );
  SDFFX1 DFF_30_Q_reg ( .D(WX544), .SI(WX543), .SE(n4627), .CLK(n4946), .Q(
        WX545) );
  SDFFX1 DFF_31_Q_reg ( .D(WX546), .SI(WX545), .SE(n4627), .CLK(n4946), .Q(
        WX547) );
  SDFFX1 DFF_32_Q_reg ( .D(WX644), .SI(WX547), .SE(n4622), .CLK(n4948), .Q(
        WX645), .QN(n3529) );
  SDFFX1 DFF_33_Q_reg ( .D(WX646), .SI(WX645), .SE(n4622), .CLK(n4948), .Q(
        WX647), .QN(n3527) );
  SDFFX1 DFF_34_Q_reg ( .D(WX648), .SI(WX647), .SE(n4621), .CLK(n4948), .Q(
        WX649), .QN(n3525) );
  SDFFX1 DFF_35_Q_reg ( .D(WX650), .SI(WX649), .SE(n4621), .CLK(n4948), .Q(
        test_so2) );
  SDFFX1 DFF_36_Q_reg ( .D(WX652), .SI(test_si3), .SE(n4621), .CLK(n4949), .Q(
        WX653), .QN(n3521) );
  SDFFX1 DFF_37_Q_reg ( .D(WX654), .SI(WX653), .SE(n4621), .CLK(n4949), .Q(
        WX655), .QN(n3519) );
  SDFFX1 DFF_38_Q_reg ( .D(WX656), .SI(WX655), .SE(n4620), .CLK(n4949), .Q(
        WX657), .QN(n3517) );
  SDFFX1 DFF_39_Q_reg ( .D(WX658), .SI(WX657), .SE(n4620), .CLK(n4949), .Q(
        WX659), .QN(n3515) );
  SDFFX1 DFF_40_Q_reg ( .D(WX660), .SI(WX659), .SE(n4620), .CLK(n4949), .Q(
        WX661), .QN(n3513) );
  SDFFX1 DFF_41_Q_reg ( .D(WX662), .SI(WX661), .SE(n4619), .CLK(n4949), .Q(
        WX663), .QN(n3511) );
  SDFFX1 DFF_42_Q_reg ( .D(WX664), .SI(WX663), .SE(n4619), .CLK(n4950), .Q(
        WX665), .QN(n3509) );
  SDFFX1 DFF_43_Q_reg ( .D(WX666), .SI(WX665), .SE(n4619), .CLK(n4950), .Q(
        WX667), .QN(n3507) );
  SDFFX1 DFF_44_Q_reg ( .D(WX668), .SI(WX667), .SE(n4618), .CLK(n4950), .Q(
        WX669), .QN(n3505) );
  SDFFX1 DFF_45_Q_reg ( .D(WX670), .SI(WX669), .SE(n4618), .CLK(n4950), .Q(
        WX671), .QN(n3503) );
  SDFFX1 DFF_46_Q_reg ( .D(WX672), .SI(WX671), .SE(n4617), .CLK(n4950), .Q(
        WX673), .QN(n3501) );
  SDFFX1 DFF_47_Q_reg ( .D(WX674), .SI(WX673), .SE(n4617), .CLK(n4951), .Q(
        WX675), .QN(n3499) );
  SDFFX1 DFF_48_Q_reg ( .D(WX676), .SI(WX675), .SE(n4616), .CLK(n4951), .Q(
        WX677), .QN(n3497) );
  SDFFX1 DFF_49_Q_reg ( .D(WX678), .SI(WX677), .SE(n4616), .CLK(n4951), .Q(
        WX679), .QN(n3495) );
  SDFFX1 DFF_50_Q_reg ( .D(WX680), .SI(WX679), .SE(n4615), .CLK(n4952), .Q(
        WX681), .QN(n3493) );
  SDFFX1 DFF_51_Q_reg ( .D(WX682), .SI(WX681), .SE(n4614), .CLK(n4952), .Q(
        WX683), .QN(n3491) );
  SDFFX1 DFF_52_Q_reg ( .D(WX684), .SI(WX683), .SE(n4614), .CLK(n4952), .Q(
        WX685), .QN(n3489) );
  SDFFX1 DFF_53_Q_reg ( .D(WX686), .SI(WX685), .SE(n4613), .CLK(n4953), .Q(
        test_so3) );
  SDFFX1 DFF_54_Q_reg ( .D(WX688), .SI(test_si4), .SE(n4342), .CLK(n5089), .Q(
        WX689), .QN(n3485) );
  SDFFX1 DFF_55_Q_reg ( .D(WX690), .SI(WX689), .SE(n4611), .CLK(n4953), .Q(
        WX691), .QN(n3483) );
  SDFFX1 DFF_56_Q_reg ( .D(WX692), .SI(WX691), .SE(n4611), .CLK(n4954), .Q(
        WX693), .QN(n3481) );
  SDFFX1 DFF_57_Q_reg ( .D(WX694), .SI(WX693), .SE(n4610), .CLK(n4954), .Q(
        WX695), .QN(n3479) );
  SDFFX1 DFF_58_Q_reg ( .D(WX696), .SI(WX695), .SE(n4610), .CLK(n4954), .Q(
        WX697), .QN(n3477) );
  SDFFX1 DFF_59_Q_reg ( .D(WX698), .SI(WX697), .SE(n4609), .CLK(n4955), .Q(
        WX699), .QN(n3475) );
  SDFFX1 DFF_60_Q_reg ( .D(WX700), .SI(WX699), .SE(n4608), .CLK(n4955), .Q(
        WX701), .QN(n3473) );
  SDFFX1 DFF_61_Q_reg ( .D(WX702), .SI(WX701), .SE(n4608), .CLK(n4955), .Q(
        WX703), .QN(n3471) );
  SDFFX1 DFF_62_Q_reg ( .D(WX704), .SI(WX703), .SE(n4607), .CLK(n4956), .Q(
        WX705), .QN(n3469) );
  SDFFX1 DFF_63_Q_reg ( .D(WX706), .SI(WX705), .SE(n4606), .CLK(n4956), .Q(
        WX707), .QN(n3467) );
  SDFFX1 DFF_64_Q_reg ( .D(WX708), .SI(WX707), .SE(n4606), .CLK(n4956), .Q(
        WX709) );
  SDFFX1 DFF_65_Q_reg ( .D(WX710), .SI(WX709), .SE(n4605), .CLK(n4956), .Q(
        WX711), .QN(n4180) );
  SDFFX1 DFF_66_Q_reg ( .D(WX712), .SI(WX711), .SE(n4605), .CLK(n4957), .Q(
        WX713), .QN(n9087) );
  SDFFX1 DFF_67_Q_reg ( .D(WX714), .SI(WX713), .SE(n4621), .CLK(n4949), .Q(
        WX715), .QN(n4189) );
  SDFFX1 DFF_68_Q_reg ( .D(WX716), .SI(WX715), .SE(n4621), .CLK(n4949), .Q(
        WX717), .QN(n9088) );
  SDFFX1 DFF_69_Q_reg ( .D(WX718), .SI(WX717), .SE(n4620), .CLK(n4949), .Q(
        WX719), .QN(n9089) );
  SDFFX1 DFF_70_Q_reg ( .D(WX720), .SI(WX719), .SE(n4620), .CLK(n4949), .Q(
        WX721), .QN(n9090) );
  SDFFX1 DFF_71_Q_reg ( .D(WX722), .SI(WX721), .SE(n4620), .CLK(n4949), .Q(
        test_so4) );
  SDFFX1 DFF_72_Q_reg ( .D(WX724), .SI(test_si5), .SE(n4619), .CLK(n4949), .Q(
        WX725), .QN(n9091) );
  SDFFX1 DFF_73_Q_reg ( .D(WX726), .SI(WX725), .SE(n4619), .CLK(n4950), .Q(
        WX727), .QN(n4206) );
  SDFFX1 DFF_74_Q_reg ( .D(WX728), .SI(WX727), .SE(n4619), .CLK(n4950), .Q(
        WX729), .QN(n4210) );
  SDFFX1 DFF_75_Q_reg ( .D(WX730), .SI(WX729), .SE(n4618), .CLK(n4950), .Q(
        WX731) );
  SDFFX1 DFF_76_Q_reg ( .D(WX732), .SI(WX731), .SE(n4618), .CLK(n4950), .Q(
        WX733), .QN(n9092) );
  SDFFX1 DFF_77_Q_reg ( .D(WX734), .SI(WX733), .SE(n4618), .CLK(n4950), .Q(
        WX735), .QN(n9093) );
  SDFFX1 DFF_78_Q_reg ( .D(WX736), .SI(WX735), .SE(n4617), .CLK(n4951), .Q(
        WX737), .QN(n9094) );
  SDFFX1 DFF_79_Q_reg ( .D(WX738), .SI(WX737), .SE(n4617), .CLK(n4951), .Q(
        WX739) );
  SDFFX1 DFF_80_Q_reg ( .D(WX740), .SI(WX739), .SE(n4616), .CLK(n4951), .Q(
        WX741), .QN(n4208) );
  SDFFX1 DFF_81_Q_reg ( .D(WX742), .SI(WX741), .SE(n4615), .CLK(n4951), .Q(
        WX743), .QN(n9095) );
  SDFFX1 DFF_82_Q_reg ( .D(WX744), .SI(WX743), .SE(n4615), .CLK(n4952), .Q(
        WX745), .QN(n9096) );
  SDFFX1 DFF_83_Q_reg ( .D(WX746), .SI(WX745), .SE(n4614), .CLK(n4952), .Q(
        WX747), .QN(n9097) );
  SDFFX1 DFF_84_Q_reg ( .D(WX748), .SI(WX747), .SE(n4613), .CLK(n4952), .Q(
        WX749), .QN(n9098) );
  SDFFX1 DFF_85_Q_reg ( .D(WX750), .SI(WX749), .SE(n4613), .CLK(n4953), .Q(
        WX751), .QN(n4194) );
  SDFFX1 DFF_86_Q_reg ( .D(WX752), .SI(WX751), .SE(n4612), .CLK(n4953), .Q(
        WX753) );
  SDFFX1 DFF_87_Q_reg ( .D(WX754), .SI(WX753), .SE(n4612), .CLK(n4953), .Q(
        WX755), .QN(n9082) );
  SDFFX1 DFF_88_Q_reg ( .D(WX756), .SI(WX755), .SE(n4611), .CLK(n4954), .Q(
        WX757), .QN(n4218) );
  SDFFX1 DFF_89_Q_reg ( .D(WX758), .SI(WX757), .SE(n4610), .CLK(n4954), .Q(
        test_so5) );
  SDFFX1 DFF_90_Q_reg ( .D(WX760), .SI(test_si6), .SE(n4610), .CLK(n4954), .Q(
        WX761), .QN(n9083) );
  SDFFX1 DFF_91_Q_reg ( .D(WX762), .SI(WX761), .SE(n4609), .CLK(n4955), .Q(
        WX763), .QN(n9084) );
  SDFFX1 DFF_92_Q_reg ( .D(WX764), .SI(WX763), .SE(n4608), .CLK(n4955), .Q(
        WX765), .QN(n9086) );
  SDFFX1 DFF_93_Q_reg ( .D(WX766), .SI(WX765), .SE(n4608), .CLK(n4955), .Q(
        WX767) );
  SDFFX1 DFF_94_Q_reg ( .D(WX768), .SI(WX767), .SE(n4607), .CLK(n4956), .Q(
        WX769), .QN(n9099) );
  SDFFX1 DFF_95_Q_reg ( .D(WX770), .SI(WX769), .SE(n4606), .CLK(n4956), .Q(
        WX771), .QN(n4221) );
  SDFFX1 DFF_96_Q_reg ( .D(WX772), .SI(WX771), .SE(n4606), .CLK(n4956), .Q(
        WX773), .QN(n9085) );
  SDFFX1 DFF_97_Q_reg ( .D(WX774), .SI(WX773), .SE(n4605), .CLK(n4957), .Q(
        WX775) );
  SDFFX1 DFF_98_Q_reg ( .D(WX776), .SI(WX775), .SE(n4605), .CLK(n4957), .Q(
        WX777) );
  SDFFX1 DFF_99_Q_reg ( .D(WX778), .SI(WX777), .SE(n4604), .CLK(n4957), .Q(
        WX779) );
  SDFFX1 DFF_100_Q_reg ( .D(WX780), .SI(WX779), .SE(n4604), .CLK(n4957), .Q(
        WX781) );
  SDFFX1 DFF_101_Q_reg ( .D(WX782), .SI(WX781), .SE(n4604), .CLK(n4957), .Q(
        WX783) );
  SDFFX1 DFF_102_Q_reg ( .D(WX784), .SI(WX783), .SE(n4603), .CLK(n4957), .Q(
        WX785) );
  SDFFX1 DFF_103_Q_reg ( .D(WX786), .SI(WX785), .SE(n4603), .CLK(n4958), .Q(
        WX787) );
  SDFFX1 DFF_104_Q_reg ( .D(WX788), .SI(WX787), .SE(n4603), .CLK(n4958), .Q(
        WX789) );
  SDFFX1 DFF_105_Q_reg ( .D(WX790), .SI(WX789), .SE(n4602), .CLK(n4958), .Q(
        WX791) );
  SDFFX1 DFF_106_Q_reg ( .D(WX792), .SI(WX791), .SE(n4602), .CLK(n4958), .Q(
        WX793) );
  SDFFX1 DFF_107_Q_reg ( .D(WX794), .SI(WX793), .SE(n4602), .CLK(n4958), .Q(
        test_so6) );
  SDFFX1 DFF_108_Q_reg ( .D(WX796), .SI(test_si7), .SE(n4618), .CLK(n4950), 
        .Q(WX797) );
  SDFFX1 DFF_109_Q_reg ( .D(WX798), .SI(WX797), .SE(n4617), .CLK(n4950), .Q(
        WX799) );
  SDFFX1 DFF_110_Q_reg ( .D(WX800), .SI(WX799), .SE(n4617), .CLK(n4951), .Q(
        WX801) );
  SDFFX1 DFF_111_Q_reg ( .D(WX802), .SI(WX801), .SE(n4616), .CLK(n4951), .Q(
        WX803), .QN(n4202) );
  SDFFX1 DFF_112_Q_reg ( .D(WX804), .SI(WX803), .SE(n4616), .CLK(n4951), .Q(
        WX805) );
  SDFFX1 DFF_113_Q_reg ( .D(WX806), .SI(WX805), .SE(n4615), .CLK(n4951), .Q(
        WX807) );
  SDFFX1 DFF_114_Q_reg ( .D(WX808), .SI(WX807), .SE(n4615), .CLK(n4952), .Q(
        WX809) );
  SDFFX1 DFF_115_Q_reg ( .D(WX810), .SI(WX809), .SE(n4614), .CLK(n4952), .Q(
        WX811) );
  SDFFX1 DFF_116_Q_reg ( .D(WX812), .SI(WX811), .SE(n4613), .CLK(n4952), .Q(
        WX813) );
  SDFFX1 DFF_117_Q_reg ( .D(WX814), .SI(WX813), .SE(n4613), .CLK(n4953), .Q(
        WX815) );
  SDFFX1 DFF_118_Q_reg ( .D(WX816), .SI(WX815), .SE(n4612), .CLK(n4953), .Q(
        WX817), .QN(n9081) );
  SDFFX1 DFF_119_Q_reg ( .D(WX818), .SI(WX817), .SE(n4612), .CLK(n4953), .Q(
        WX819) );
  SDFFX1 DFF_120_Q_reg ( .D(WX820), .SI(WX819), .SE(n4611), .CLK(n4954), .Q(
        WX821) );
  SDFFX1 DFF_121_Q_reg ( .D(WX822), .SI(WX821), .SE(n4610), .CLK(n4954), .Q(
        WX823) );
  SDFFX1 DFF_122_Q_reg ( .D(WX824), .SI(WX823), .SE(n4609), .CLK(n4954), .Q(
        WX825) );
  SDFFX1 DFF_123_Q_reg ( .D(WX826), .SI(WX825), .SE(n4609), .CLK(n4955), .Q(
        WX827) );
  SDFFX1 DFF_124_Q_reg ( .D(WX828), .SI(WX827), .SE(n4608), .CLK(n4955), .Q(
        WX829) );
  SDFFX1 DFF_125_Q_reg ( .D(WX830), .SI(WX829), .SE(n4607), .CLK(n4955), .Q(
        test_so7) );
  SDFFX1 DFF_126_Q_reg ( .D(WX832), .SI(test_si8), .SE(n4607), .CLK(n4956), 
        .Q(WX833) );
  SDFFX1 DFF_127_Q_reg ( .D(WX834), .SI(WX833), .SE(n4606), .CLK(n4956), .Q(
        WX835) );
  SDFFX1 DFF_128_Q_reg ( .D(WX836), .SI(WX835), .SE(n4605), .CLK(n4956), .Q(
        WX837), .QN(n4215) );
  SDFFX1 DFF_129_Q_reg ( .D(WX838), .SI(WX837), .SE(n4605), .CLK(n4957), .Q(
        WX839), .QN(n4181) );
  SDFFX1 DFF_130_Q_reg ( .D(WX840), .SI(WX839), .SE(n4604), .CLK(n4957), .Q(
        WX841), .QN(n4184) );
  SDFFX1 DFF_131_Q_reg ( .D(WX842), .SI(WX841), .SE(n4604), .CLK(n4957), .Q(
        WX843), .QN(n4188) );
  SDFFX1 DFF_132_Q_reg ( .D(WX844), .SI(WX843), .SE(n4604), .CLK(n4957), .Q(
        WX845), .QN(n4191) );
  SDFFX1 DFF_133_Q_reg ( .D(WX846), .SI(WX845), .SE(n4603), .CLK(n4957), .Q(
        WX847), .QN(n4192) );
  SDFFX1 DFF_134_Q_reg ( .D(WX848), .SI(WX847), .SE(n4603), .CLK(n4958), .Q(
        WX849), .QN(n4196) );
  SDFFX1 DFF_135_Q_reg ( .D(WX850), .SI(WX849), .SE(n4603), .CLK(n4958), .Q(
        WX851), .QN(n4199) );
  SDFFX1 DFF_136_Q_reg ( .D(WX852), .SI(WX851), .SE(n4602), .CLK(n4958), .Q(
        WX853), .QN(n4201) );
  SDFFX1 DFF_137_Q_reg ( .D(WX854), .SI(WX853), .SE(n4602), .CLK(n4958), .Q(
        WX855), .QN(n4207) );
  SDFFX1 DFF_138_Q_reg ( .D(WX856), .SI(WX855), .SE(n4602), .CLK(n4958), .Q(
        WX857), .QN(n4211) );
  SDFFX1 DFF_139_Q_reg ( .D(WX858), .SI(WX857), .SE(n4601), .CLK(n4958), .Q(
        WX859), .QN(n4213) );
  SDFFX1 DFF_140_Q_reg ( .D(WX860), .SI(WX859), .SE(n4601), .CLK(n4958), .Q(
        WX861), .QN(n4183) );
  SDFFX1 DFF_141_Q_reg ( .D(WX862), .SI(WX861), .SE(n4601), .CLK(n4959), .Q(
        WX863), .QN(n4190) );
  SDFFX1 DFF_142_Q_reg ( .D(WX864), .SI(WX863), .SE(n4601), .CLK(n4959), .Q(
        WX865), .QN(n4195) );
  SDFFX1 DFF_143_Q_reg ( .D(WX866), .SI(WX865), .SE(n4601), .CLK(n4959), .Q(
        test_so8) );
  SDFFX1 DFF_144_Q_reg ( .D(WX868), .SI(test_si9), .SE(n4616), .CLK(n4951), 
        .Q(WX869), .QN(n4209) );
  SDFFX1 DFF_145_Q_reg ( .D(WX870), .SI(WX869), .SE(n4615), .CLK(n4952), .Q(
        WX871), .QN(n4216) );
  SDFFX1 DFF_146_Q_reg ( .D(WX872), .SI(WX871), .SE(n4614), .CLK(n4952), .Q(
        WX873), .QN(n4185) );
  SDFFX1 DFF_147_Q_reg ( .D(WX874), .SI(WX873), .SE(n4614), .CLK(n4952), .Q(
        WX875), .QN(n4197) );
  SDFFX1 DFF_148_Q_reg ( .D(WX876), .SI(WX875), .SE(n4613), .CLK(n4953), .Q(
        WX877), .QN(n4220) );
  SDFFX1 DFF_149_Q_reg ( .D(WX878), .SI(WX877), .SE(n4612), .CLK(n4953), .Q(
        WX879), .QN(n4193) );
  SDFFX1 DFF_150_Q_reg ( .D(WX880), .SI(WX879), .SE(n4612), .CLK(n4953), .Q(
        WX881), .QN(n4198) );
  SDFFX1 DFF_151_Q_reg ( .D(WX882), .SI(WX881), .SE(n4611), .CLK(n4953), .Q(
        WX883), .QN(n4203) );
  SDFFX1 DFF_152_Q_reg ( .D(WX884), .SI(WX883), .SE(n4611), .CLK(n4954), .Q(
        WX885), .QN(n4219) );
  SDFFX1 DFF_153_Q_reg ( .D(WX886), .SI(WX885), .SE(n4610), .CLK(n4954), .Q(
        WX887), .QN(n4212) );
  SDFFX1 DFF_154_Q_reg ( .D(WX888), .SI(WX887), .SE(n4609), .CLK(n4954), .Q(
        WX889), .QN(n4204) );
  SDFFX1 DFF_155_Q_reg ( .D(WX890), .SI(WX889), .SE(n4609), .CLK(n4955), .Q(
        WX891), .QN(n4205) );
  SDFFX1 DFF_156_Q_reg ( .D(WX892), .SI(WX891), .SE(n4608), .CLK(n4955), .Q(
        WX893), .QN(n4182) );
  SDFFX1 DFF_157_Q_reg ( .D(WX894), .SI(WX893), .SE(n4607), .CLK(n4955), .Q(
        WX895), .QN(n4217) );
  SDFFX1 DFF_158_Q_reg ( .D(WX896), .SI(WX895), .SE(n4607), .CLK(n4956), .Q(
        WX897), .QN(n4186) );
  SDFFX1 DFF_159_Q_reg ( .D(WX898), .SI(WX897), .SE(n4606), .CLK(n4956), .Q(
        WX899), .QN(n4222) );
  SDFFX1 DFF_160_Q_reg ( .D(WX1264), .SI(WX899), .SE(n4344), .CLK(n5088), .Q(
        CRC_OUT_9_0), .QN(DFF_160_n1) );
  SDFFX1 DFF_161_Q_reg ( .D(WX1266), .SI(CRC_OUT_9_0), .SE(n4344), .CLK(n5088), 
        .Q(test_so9) );
  SDFFX1 DFF_162_Q_reg ( .D(WX1268), .SI(test_si10), .SE(n4344), .CLK(n5088), 
        .Q(CRC_OUT_9_2), .QN(DFF_162_n1) );
  SDFFX1 DFF_163_Q_reg ( .D(WX1270), .SI(CRC_OUT_9_2), .SE(n4343), .CLK(n5088), 
        .Q(CRC_OUT_9_3), .QN(DFF_163_n1) );
  SDFFX1 DFF_164_Q_reg ( .D(WX1272), .SI(CRC_OUT_9_3), .SE(n4343), .CLK(n5088), 
        .Q(CRC_OUT_9_4), .QN(DFF_164_n1) );
  SDFFX1 DFF_165_Q_reg ( .D(WX1274), .SI(CRC_OUT_9_4), .SE(n4343), .CLK(n5088), 
        .Q(CRC_OUT_9_5), .QN(DFF_165_n1) );
  SDFFX1 DFF_166_Q_reg ( .D(WX1276), .SI(CRC_OUT_9_5), .SE(n4343), .CLK(n5088), 
        .Q(CRC_OUT_9_6), .QN(DFF_166_n1) );
  SDFFX1 DFF_167_Q_reg ( .D(WX1278), .SI(CRC_OUT_9_6), .SE(n4343), .CLK(n5088), 
        .Q(CRC_OUT_9_7), .QN(DFF_167_n1) );
  SDFFX1 DFF_168_Q_reg ( .D(WX1280), .SI(CRC_OUT_9_7), .SE(n4343), .CLK(n5088), 
        .Q(CRC_OUT_9_8), .QN(DFF_168_n1) );
  SDFFX1 DFF_169_Q_reg ( .D(WX1282), .SI(CRC_OUT_9_8), .SE(n4342), .CLK(n5089), 
        .Q(CRC_OUT_9_9), .QN(DFF_169_n1) );
  SDFFX1 DFF_170_Q_reg ( .D(WX1284), .SI(CRC_OUT_9_9), .SE(n4342), .CLK(n5089), 
        .Q(CRC_OUT_9_10), .QN(DFF_170_n1) );
  SDFFX1 DFF_171_Q_reg ( .D(WX1286), .SI(CRC_OUT_9_10), .SE(n4342), .CLK(n5089), .Q(CRC_OUT_9_11), .QN(DFF_171_n1) );
  SDFFX1 DFF_172_Q_reg ( .D(WX1288), .SI(CRC_OUT_9_11), .SE(n4342), .CLK(n5089), .Q(CRC_OUT_9_12), .QN(DFF_172_n1) );
  SDFFX1 DFF_173_Q_reg ( .D(WX1290), .SI(CRC_OUT_9_12), .SE(n4342), .CLK(n5089), .Q(CRC_OUT_9_13), .QN(DFF_173_n1) );
  SDFFX1 DFF_174_Q_reg ( .D(WX1292), .SI(CRC_OUT_9_13), .SE(n4341), .CLK(n5089), .Q(CRC_OUT_9_14), .QN(DFF_174_n1) );
  SDFFX1 DFF_175_Q_reg ( .D(WX1294), .SI(CRC_OUT_9_14), .SE(n4341), .CLK(n5089), .Q(CRC_OUT_9_15), .QN(DFF_175_n1) );
  SDFFX1 DFF_176_Q_reg ( .D(WX1296), .SI(CRC_OUT_9_15), .SE(n4341), .CLK(n5089), .Q(CRC_OUT_9_16), .QN(DFF_176_n1) );
  SDFFX1 DFF_177_Q_reg ( .D(WX1298), .SI(CRC_OUT_9_16), .SE(n4341), .CLK(n5089), .Q(CRC_OUT_9_17), .QN(DFF_177_n1) );
  SDFFX1 DFF_178_Q_reg ( .D(WX1300), .SI(CRC_OUT_9_17), .SE(n4341), .CLK(n5089), .Q(CRC_OUT_9_18), .QN(DFF_178_n1) );
  SDFFX1 DFF_179_Q_reg ( .D(WX1302), .SI(CRC_OUT_9_18), .SE(n4341), .CLK(n5089), .Q(test_so10) );
  SDFFX1 DFF_180_Q_reg ( .D(WX1304), .SI(test_si11), .SE(n4601), .CLK(n4959), 
        .Q(CRC_OUT_9_20), .QN(DFF_180_n1) );
  SDFFX1 DFF_181_Q_reg ( .D(WX1306), .SI(CRC_OUT_9_20), .SE(n4600), .CLK(n4959), .Q(CRC_OUT_9_21), .QN(DFF_181_n1) );
  SDFFX1 DFF_182_Q_reg ( .D(WX1308), .SI(CRC_OUT_9_21), .SE(n4600), .CLK(n4959), .Q(CRC_OUT_9_22), .QN(DFF_182_n1) );
  SDFFX1 DFF_183_Q_reg ( .D(WX1310), .SI(CRC_OUT_9_22), .SE(n4600), .CLK(n4959), .Q(CRC_OUT_9_23), .QN(DFF_183_n1) );
  SDFFX1 DFF_184_Q_reg ( .D(WX1312), .SI(CRC_OUT_9_23), .SE(n4600), .CLK(n4959), .Q(CRC_OUT_9_24), .QN(DFF_184_n1) );
  SDFFX1 DFF_185_Q_reg ( .D(WX1314), .SI(CRC_OUT_9_24), .SE(n4600), .CLK(n4959), .Q(CRC_OUT_9_25), .QN(DFF_185_n1) );
  SDFFX1 DFF_186_Q_reg ( .D(WX1316), .SI(CRC_OUT_9_25), .SE(n4600), .CLK(n4959), .Q(CRC_OUT_9_26), .QN(DFF_186_n1) );
  SDFFX1 DFF_187_Q_reg ( .D(WX1318), .SI(CRC_OUT_9_26), .SE(n4599), .CLK(n4959), .Q(CRC_OUT_9_27), .QN(DFF_187_n1) );
  SDFFX1 DFF_188_Q_reg ( .D(WX1320), .SI(CRC_OUT_9_27), .SE(n4599), .CLK(n4959), .Q(CRC_OUT_9_28), .QN(DFF_188_n1) );
  SDFFX1 DFF_189_Q_reg ( .D(WX1322), .SI(CRC_OUT_9_28), .SE(n4599), .CLK(n4960), .Q(CRC_OUT_9_29), .QN(DFF_189_n1) );
  SDFFX1 DFF_190_Q_reg ( .D(WX1324), .SI(CRC_OUT_9_29), .SE(n4599), .CLK(n4960), .Q(CRC_OUT_9_30), .QN(DFF_190_n1) );
  SDFFX1 DFF_191_Q_reg ( .D(WX1326), .SI(CRC_OUT_9_30), .SE(n4599), .CLK(n4960), .Q(CRC_OUT_9_31), .QN(DFF_191_n1) );
  SDFFX1 DFF_192_Q_reg ( .D(n2), .SI(CRC_OUT_9_31), .SE(n4599), .CLK(n4960), 
        .Q(WX1778), .QN(n3938) );
  SDFFX1 DFF_193_Q_reg ( .D(n3), .SI(WX1778), .SE(n4593), .CLK(n4962), .Q(
        n8702) );
  SDFFX1 DFF_194_Q_reg ( .D(n4), .SI(n8702), .SE(n4594), .CLK(n4962), .Q(n8701) );
  SDFFX1 DFF_195_Q_reg ( .D(n5), .SI(n8701), .SE(n4594), .CLK(n4962), .Q(n8700) );
  SDFFX1 DFF_196_Q_reg ( .D(n6), .SI(n8700), .SE(n4594), .CLK(n4962), .Q(n8699) );
  SDFFX1 DFF_197_Q_reg ( .D(n7), .SI(n8699), .SE(n4594), .CLK(n4962), .Q(
        test_so11) );
  SDFFX1 DFF_198_Q_reg ( .D(n8), .SI(test_si12), .SE(n4594), .CLK(n4962), .Q(
        n8696) );
  SDFFX1 DFF_199_Q_reg ( .D(n9), .SI(n8696), .SE(n4594), .CLK(n4962), .Q(n8695) );
  SDFFX1 DFF_200_Q_reg ( .D(n10), .SI(n8695), .SE(n4595), .CLK(n4962), .Q(
        n8694) );
  SDFFX1 DFF_201_Q_reg ( .D(n11), .SI(n8694), .SE(n4595), .CLK(n4962), .Q(
        n8693) );
  SDFFX1 DFF_202_Q_reg ( .D(n12), .SI(n8693), .SE(n4595), .CLK(n4962), .Q(
        n8692) );
  SDFFX1 DFF_203_Q_reg ( .D(n13), .SI(n8692), .SE(n4595), .CLK(n4962), .Q(
        n8691) );
  SDFFX1 DFF_204_Q_reg ( .D(n14), .SI(n8691), .SE(n4595), .CLK(n4961), .Q(
        n8690) );
  SDFFX1 DFF_205_Q_reg ( .D(n15), .SI(n8690), .SE(n4595), .CLK(n4961), .Q(
        n8689) );
  SDFFX1 DFF_206_Q_reg ( .D(n16), .SI(n8689), .SE(n4596), .CLK(n4961), .Q(
        n8688) );
  SDFFX1 DFF_207_Q_reg ( .D(n17), .SI(n8688), .SE(n4596), .CLK(n4961), .Q(
        n8687) );
  SDFFX1 DFF_208_Q_reg ( .D(n18), .SI(n8687), .SE(n4596), .CLK(n4961), .Q(
        n8686) );
  SDFFX1 DFF_209_Q_reg ( .D(n19), .SI(n8686), .SE(n4596), .CLK(n4961), .Q(
        n8685) );
  SDFFX1 DFF_210_Q_reg ( .D(n20), .SI(n8685), .SE(n4596), .CLK(n4961), .Q(
        n8684) );
  SDFFX1 DFF_211_Q_reg ( .D(n21), .SI(n8684), .SE(n4596), .CLK(n4961), .Q(
        n8683) );
  SDFFX1 DFF_212_Q_reg ( .D(n22), .SI(n8683), .SE(n4597), .CLK(n4961), .Q(
        n8682) );
  SDFFX1 DFF_213_Q_reg ( .D(n23), .SI(n8682), .SE(n4597), .CLK(n4961), .Q(
        n8681) );
  SDFFX1 DFF_214_Q_reg ( .D(n24), .SI(n8681), .SE(n4597), .CLK(n4961), .Q(
        n8680) );
  SDFFX1 DFF_215_Q_reg ( .D(n25), .SI(n8680), .SE(n4597), .CLK(n4961), .Q(
        test_so12) );
  SDFFX1 DFF_216_Q_reg ( .D(n26), .SI(test_si13), .SE(n4597), .CLK(n4960), .Q(
        n8677) );
  SDFFX1 DFF_217_Q_reg ( .D(n27), .SI(n8677), .SE(n4597), .CLK(n4960), .Q(
        n8676) );
  SDFFX1 DFF_218_Q_reg ( .D(n28), .SI(n8676), .SE(n4598), .CLK(n4960), .Q(
        n8675) );
  SDFFX1 DFF_219_Q_reg ( .D(n29), .SI(n8675), .SE(n4598), .CLK(n4960), .Q(
        n8674) );
  SDFFX1 DFF_220_Q_reg ( .D(n30), .SI(n8674), .SE(n4598), .CLK(n4960), .Q(
        n8673) );
  SDFFX1 DFF_221_Q_reg ( .D(n31), .SI(n8673), .SE(n4598), .CLK(n4960), .Q(
        n8672) );
  SDFFX1 DFF_222_Q_reg ( .D(n32), .SI(n8672), .SE(n4598), .CLK(n4960), .Q(
        n8671) );
  SDFFX1 DFF_223_Q_reg ( .D(WX1839), .SI(n8671), .SE(n4598), .CLK(n4960), .Q(
        n8670) );
  SDFFX1 DFF_224_Q_reg ( .D(WX1937), .SI(n8670), .SE(n4593), .CLK(n4962), .Q(
        n8669), .QN(n9045) );
  SDFFX1 DFF_225_Q_reg ( .D(WX1939), .SI(n8669), .SE(n4592), .CLK(n4963), .Q(
        n8668), .QN(n9040) );
  SDFFX1 DFF_226_Q_reg ( .D(WX1941), .SI(n8668), .SE(n4592), .CLK(n4963), .Q(
        n8667), .QN(n9038) );
  SDFFX1 DFF_227_Q_reg ( .D(WX1943), .SI(n8667), .SE(n4351), .CLK(n5084), .Q(
        n8666), .QN(n9036) );
  SDFFX1 DFF_228_Q_reg ( .D(WX1945), .SI(n8666), .SE(n4591), .CLK(n4964), .Q(
        n8665), .QN(n9034) );
  SDFFX1 DFF_229_Q_reg ( .D(WX1947), .SI(n8665), .SE(n4591), .CLK(n4964), .Q(
        n8664), .QN(n9030) );
  SDFFX1 DFF_230_Q_reg ( .D(WX1949), .SI(n8664), .SE(n4590), .CLK(n4964), .Q(
        n8663), .QN(n9028) );
  SDFFX1 DFF_231_Q_reg ( .D(WX1951), .SI(n8663), .SE(n4589), .CLK(n4964), .Q(
        n8662), .QN(n9026) );
  SDFFX1 DFF_232_Q_reg ( .D(WX1953), .SI(n8662), .SE(n4588), .CLK(n4965), .Q(
        n8661), .QN(n9024) );
  SDFFX1 DFF_233_Q_reg ( .D(WX1955), .SI(n8661), .SE(n4588), .CLK(n4965), .Q(
        test_so13) );
  SDFFX1 DFF_234_Q_reg ( .D(WX1957), .SI(test_si14), .SE(n4587), .CLK(n4966), 
        .Q(n8658), .QN(n9021) );
  SDFFX1 DFF_235_Q_reg ( .D(WX1959), .SI(n8658), .SE(n4587), .CLK(n4966), .Q(
        n8657), .QN(n9019) );
  SDFFX1 DFF_236_Q_reg ( .D(WX1961), .SI(n8657), .SE(n4586), .CLK(n4966), .Q(
        n8656), .QN(n9017) );
  SDFFX1 DFF_237_Q_reg ( .D(WX1963), .SI(n8656), .SE(n4585), .CLK(n4966), .Q(
        n8655), .QN(n9013) );
  SDFFX1 DFF_238_Q_reg ( .D(WX1965), .SI(n8655), .SE(n4351), .CLK(n5084), .Q(
        n8654), .QN(n9011) );
  SDFFX1 DFF_239_Q_reg ( .D(WX1967), .SI(n8654), .SE(n4351), .CLK(n5084), .Q(
        n8653), .QN(n9010) );
  SDFFX1 DFF_240_Q_reg ( .D(WX1969), .SI(n8653), .SE(n4584), .CLK(n4967), .Q(
        WX1970) );
  SDFFX1 DFF_241_Q_reg ( .D(WX1971), .SI(WX1970), .SE(n4584), .CLK(n4967), .Q(
        WX1972) );
  SDFFX1 DFF_242_Q_reg ( .D(WX1973), .SI(WX1972), .SE(n4583), .CLK(n4967), .Q(
        WX1974) );
  SDFFX1 DFF_243_Q_reg ( .D(WX1975), .SI(WX1974), .SE(n4583), .CLK(n4967), .Q(
        WX1976) );
  SDFFX1 DFF_244_Q_reg ( .D(WX1977), .SI(WX1976), .SE(n4583), .CLK(n4968), .Q(
        WX1978) );
  SDFFX1 DFF_245_Q_reg ( .D(WX1979), .SI(WX1978), .SE(n4583), .CLK(n4968), .Q(
        WX1980) );
  SDFFX1 DFF_246_Q_reg ( .D(WX1981), .SI(WX1980), .SE(n4583), .CLK(n4968), .Q(
        WX1982) );
  SDFFX1 DFF_247_Q_reg ( .D(WX1983), .SI(WX1982), .SE(n4583), .CLK(n4968), .Q(
        WX1984) );
  SDFFX1 DFF_248_Q_reg ( .D(WX1985), .SI(WX1984), .SE(n4582), .CLK(n4968), .Q(
        WX1986) );
  SDFFX1 DFF_249_Q_reg ( .D(WX1987), .SI(WX1986), .SE(n4582), .CLK(n4968), .Q(
        WX1988) );
  SDFFX1 DFF_250_Q_reg ( .D(WX1989), .SI(WX1988), .SE(n4582), .CLK(n4968), .Q(
        WX1990) );
  SDFFX1 DFF_251_Q_reg ( .D(WX1991), .SI(WX1990), .SE(n4582), .CLK(n4968), .Q(
        test_so14) );
  SDFFX1 DFF_252_Q_reg ( .D(WX1993), .SI(test_si15), .SE(n4581), .CLK(n4968), 
        .Q(WX1994) );
  SDFFX1 DFF_253_Q_reg ( .D(WX1995), .SI(WX1994), .SE(n4581), .CLK(n4968), .Q(
        WX1996) );
  SDFFX1 DFF_254_Q_reg ( .D(WX1997), .SI(WX1996), .SE(n4581), .CLK(n4969), .Q(
        WX1998) );
  SDFFX1 DFF_255_Q_reg ( .D(WX1999), .SI(WX1998), .SE(n4581), .CLK(n4969), .Q(
        WX2000) );
  SDFFX1 DFF_256_Q_reg ( .D(WX2001), .SI(WX2000), .SE(n4593), .CLK(n4963), .Q(
        WX2002), .QN(n3589) );
  SDFFX1 DFF_257_Q_reg ( .D(WX2003), .SI(WX2002), .SE(n4593), .CLK(n4963), .Q(
        WX2004), .QN(n3695) );
  SDFFX1 DFF_258_Q_reg ( .D(WX2005), .SI(WX2004), .SE(n4592), .CLK(n4963), .Q(
        WX2006), .QN(n3694) );
  SDFFX1 DFF_259_Q_reg ( .D(WX2007), .SI(WX2006), .SE(n4592), .CLK(n4963), .Q(
        WX2008) );
  SDFFX1 DFF_260_Q_reg ( .D(WX2009), .SI(WX2008), .SE(n4591), .CLK(n4963), .Q(
        WX2010), .QN(n3692) );
  SDFFX1 DFF_261_Q_reg ( .D(WX2011), .SI(WX2010), .SE(n4591), .CLK(n4964), .Q(
        WX2012), .QN(n3691) );
  SDFFX1 DFF_262_Q_reg ( .D(WX2013), .SI(WX2012), .SE(n4590), .CLK(n4964), .Q(
        WX2014), .QN(n3690) );
  SDFFX1 DFF_263_Q_reg ( .D(WX2015), .SI(WX2014), .SE(n4589), .CLK(n4964), .Q(
        WX2016), .QN(n3689) );
  SDFFX1 DFF_264_Q_reg ( .D(WX2017), .SI(WX2016), .SE(n4589), .CLK(n4965), .Q(
        WX2018), .QN(n3688) );
  SDFFX1 DFF_265_Q_reg ( .D(WX2019), .SI(WX2018), .SE(n4588), .CLK(n4965), .Q(
        WX2020) );
  SDFFX1 DFF_266_Q_reg ( .D(WX2021), .SI(WX2020), .SE(n4587), .CLK(n4965), .Q(
        WX2022), .QN(n3686) );
  SDFFX1 DFF_267_Q_reg ( .D(WX2023), .SI(WX2022), .SE(n4587), .CLK(n4966), .Q(
        WX2024), .QN(n3685) );
  SDFFX1 DFF_268_Q_reg ( .D(WX2025), .SI(WX2024), .SE(n4586), .CLK(n4966), .Q(
        WX2026), .QN(n3684) );
  SDFFX1 DFF_269_Q_reg ( .D(WX2027), .SI(WX2026), .SE(n4585), .CLK(n4966), .Q(
        test_so15), .QN(n9014) );
  SDFFX1 DFF_270_Q_reg ( .D(WX2029), .SI(test_si16), .SE(n4351), .CLK(n5084), 
        .Q(WX2030), .QN(n3683) );
  SDFFX1 DFF_271_Q_reg ( .D(WX2031), .SI(WX2030), .SE(n4351), .CLK(n5084), .Q(
        WX2032), .QN(n3682) );
  SDFFX1 DFF_272_Q_reg ( .D(WX2033), .SI(WX2032), .SE(n4351), .CLK(n5084), .Q(
        WX2034), .QN(n9008) );
  SDFFX1 DFF_273_Q_reg ( .D(WX2035), .SI(WX2034), .SE(n4350), .CLK(n5085), .Q(
        WX2036), .QN(n9006) );
  SDFFX1 DFF_274_Q_reg ( .D(WX2037), .SI(WX2036), .SE(n4350), .CLK(n5085), .Q(
        WX2038), .QN(n9004) );
  SDFFX1 DFF_275_Q_reg ( .D(WX2039), .SI(WX2038), .SE(n4349), .CLK(n5085), .Q(
        WX2040), .QN(n9002) );
  SDFFX1 DFF_276_Q_reg ( .D(WX2041), .SI(WX2040), .SE(n4349), .CLK(n5085), .Q(
        WX2042), .QN(n9000) );
  SDFFX1 DFF_277_Q_reg ( .D(WX2043), .SI(WX2042), .SE(n4348), .CLK(n5086), .Q(
        WX2044), .QN(n8998) );
  SDFFX1 DFF_278_Q_reg ( .D(WX2045), .SI(WX2044), .SE(n4348), .CLK(n5086), .Q(
        WX2046), .QN(n8996) );
  SDFFX1 DFF_279_Q_reg ( .D(WX2047), .SI(WX2046), .SE(n4347), .CLK(n5086), .Q(
        WX2048), .QN(n8994) );
  SDFFX1 DFF_280_Q_reg ( .D(WX2049), .SI(WX2048), .SE(n4347), .CLK(n5086), .Q(
        WX2050), .QN(n8992) );
  SDFFX1 DFF_281_Q_reg ( .D(WX2051), .SI(WX2050), .SE(n4346), .CLK(n5087), .Q(
        WX2052), .QN(n8990) );
  SDFFX1 DFF_282_Q_reg ( .D(WX2053), .SI(WX2052), .SE(n4346), .CLK(n5087), .Q(
        WX2054), .QN(n8988) );
  SDFFX1 DFF_283_Q_reg ( .D(WX2055), .SI(WX2054), .SE(n4582), .CLK(n4968), .Q(
        WX2056), .QN(n8986) );
  SDFFX1 DFF_284_Q_reg ( .D(WX2057), .SI(WX2056), .SE(n4582), .CLK(n4968), .Q(
        WX2058), .QN(n8984) );
  SDFFX1 DFF_285_Q_reg ( .D(WX2059), .SI(WX2058), .SE(n4581), .CLK(n4969), .Q(
        WX2060), .QN(n8982) );
  SDFFX1 DFF_286_Q_reg ( .D(WX2061), .SI(WX2060), .SE(n4581), .CLK(n4969), .Q(
        WX2062), .QN(n8980) );
  SDFFX1 DFF_287_Q_reg ( .D(WX2063), .SI(WX2062), .SE(n4580), .CLK(n4969), .Q(
        test_so16) );
  SDFFX1 DFF_288_Q_reg ( .D(WX2065), .SI(test_si17), .SE(n4593), .CLK(n4963), 
        .Q(WX2066) );
  SDFFX1 DFF_289_Q_reg ( .D(WX2067), .SI(WX2066), .SE(n4593), .CLK(n4963), .Q(
        WX2068) );
  SDFFX1 DFF_290_Q_reg ( .D(WX2069), .SI(WX2068), .SE(n4592), .CLK(n4963), .Q(
        WX2070) );
  SDFFX1 DFF_291_Q_reg ( .D(WX2071), .SI(WX2070), .SE(n4592), .CLK(n4963), .Q(
        WX2072), .QN(n3693) );
  SDFFX1 DFF_292_Q_reg ( .D(WX2073), .SI(WX2072), .SE(n4591), .CLK(n4963), .Q(
        WX2074) );
  SDFFX1 DFF_293_Q_reg ( .D(WX2075), .SI(WX2074), .SE(n4590), .CLK(n4964), .Q(
        WX2076) );
  SDFFX1 DFF_294_Q_reg ( .D(WX2077), .SI(WX2076), .SE(n4590), .CLK(n4964), .Q(
        WX2078) );
  SDFFX1 DFF_295_Q_reg ( .D(WX2079), .SI(WX2078), .SE(n4589), .CLK(n4965), .Q(
        WX2080) );
  SDFFX1 DFF_296_Q_reg ( .D(WX2081), .SI(WX2080), .SE(n4589), .CLK(n4965), .Q(
        WX2082) );
  SDFFX1 DFF_297_Q_reg ( .D(WX2083), .SI(WX2082), .SE(n4588), .CLK(n4965), .Q(
        WX2084), .QN(n3687) );
  SDFFX1 DFF_298_Q_reg ( .D(WX2085), .SI(WX2084), .SE(n4587), .CLK(n4965), .Q(
        WX2086) );
  SDFFX1 DFF_299_Q_reg ( .D(WX2087), .SI(WX2086), .SE(n4586), .CLK(n4966), .Q(
        WX2088) );
  SDFFX1 DFF_300_Q_reg ( .D(WX2089), .SI(WX2088), .SE(n4586), .CLK(n4966), .Q(
        WX2090) );
  SDFFX1 DFF_301_Q_reg ( .D(WX2091), .SI(WX2090), .SE(n4585), .CLK(n4967), .Q(
        WX2092), .QN(n9015) );
  SDFFX1 DFF_302_Q_reg ( .D(WX2093), .SI(WX2092), .SE(n4585), .CLK(n4967), .Q(
        WX2094) );
  SDFFX1 DFF_303_Q_reg ( .D(WX2095), .SI(WX2094), .SE(n4584), .CLK(n4967), .Q(
        WX2096) );
  SDFFX1 DFF_304_Q_reg ( .D(WX2097), .SI(WX2096), .SE(n4584), .CLK(n4967), .Q(
        WX2098), .QN(n3929) );
  SDFFX1 DFF_305_Q_reg ( .D(WX2099), .SI(WX2098), .SE(n4350), .CLK(n5085), .Q(
        test_so17) );
  SDFFX1 DFF_306_Q_reg ( .D(WX2101), .SI(test_si18), .SE(n4350), .CLK(n5085), 
        .Q(WX2102), .QN(n3926) );
  SDFFX1 DFF_307_Q_reg ( .D(WX2103), .SI(WX2102), .SE(n4349), .CLK(n5085), .Q(
        WX2104), .QN(n3924) );
  SDFFX1 DFF_308_Q_reg ( .D(WX2105), .SI(WX2104), .SE(n4349), .CLK(n5085), .Q(
        WX2106), .QN(n3922) );
  SDFFX1 DFF_309_Q_reg ( .D(WX2107), .SI(WX2106), .SE(n4348), .CLK(n5086), .Q(
        WX2108), .QN(n3920) );
  SDFFX1 DFF_310_Q_reg ( .D(WX2109), .SI(WX2108), .SE(n4348), .CLK(n5086), .Q(
        WX2110), .QN(n3918) );
  SDFFX1 DFF_311_Q_reg ( .D(WX2111), .SI(WX2110), .SE(n4347), .CLK(n5086), .Q(
        WX2112), .QN(n3916) );
  SDFFX1 DFF_312_Q_reg ( .D(WX2113), .SI(WX2112), .SE(n4347), .CLK(n5086), .Q(
        WX2114), .QN(n3914) );
  SDFFX1 DFF_313_Q_reg ( .D(WX2115), .SI(WX2114), .SE(n4346), .CLK(n5087), .Q(
        WX2116), .QN(n3912) );
  SDFFX1 DFF_314_Q_reg ( .D(WX2117), .SI(WX2116), .SE(n4346), .CLK(n5087), .Q(
        WX2118), .QN(n3910) );
  SDFFX1 DFF_315_Q_reg ( .D(WX2119), .SI(WX2118), .SE(n4345), .CLK(n5087), .Q(
        WX2120) );
  SDFFX1 DFF_316_Q_reg ( .D(WX2121), .SI(WX2120), .SE(n4345), .CLK(n5087), .Q(
        WX2122), .QN(n3907) );
  SDFFX1 DFF_317_Q_reg ( .D(WX2123), .SI(WX2122), .SE(n4345), .CLK(n5087), .Q(
        WX2124), .QN(n3905) );
  SDFFX1 DFF_318_Q_reg ( .D(WX2125), .SI(WX2124), .SE(n4344), .CLK(n5088), .Q(
        WX2126), .QN(n3903) );
  SDFFX1 DFF_319_Q_reg ( .D(WX2127), .SI(WX2126), .SE(n4580), .CLK(n4969), .Q(
        WX2128), .QN(n8978) );
  SDFFX1 DFF_320_Q_reg ( .D(WX2129), .SI(WX2128), .SE(n4580), .CLK(n4969), .Q(
        WX2130), .QN(n4154) );
  SDFFX1 DFF_321_Q_reg ( .D(WX2131), .SI(WX2130), .SE(n4580), .CLK(n4969), .Q(
        WX2132), .QN(n4155) );
  SDFFX1 DFF_322_Q_reg ( .D(WX2133), .SI(WX2132), .SE(n4580), .CLK(n4969), .Q(
        WX2134), .QN(n4156) );
  SDFFX1 DFF_323_Q_reg ( .D(WX2135), .SI(WX2134), .SE(n4580), .CLK(n4969), .Q(
        test_so18) );
  SDFFX1 DFF_324_Q_reg ( .D(WX2137), .SI(test_si19), .SE(n4591), .CLK(n4964), 
        .Q(WX2138), .QN(n4157) );
  SDFFX1 DFF_325_Q_reg ( .D(WX2139), .SI(WX2138), .SE(n4590), .CLK(n4964), .Q(
        WX2140), .QN(n4158) );
  SDFFX1 DFF_326_Q_reg ( .D(WX2141), .SI(WX2140), .SE(n4590), .CLK(n4964), .Q(
        WX2142), .QN(n4159) );
  SDFFX1 DFF_327_Q_reg ( .D(WX2143), .SI(WX2142), .SE(n4589), .CLK(n4965), .Q(
        WX2144), .QN(n4160) );
  SDFFX1 DFF_328_Q_reg ( .D(WX2145), .SI(WX2144), .SE(n4588), .CLK(n4965), .Q(
        WX2146), .QN(n4161) );
  SDFFX1 DFF_329_Q_reg ( .D(WX2147), .SI(WX2146), .SE(n4588), .CLK(n4965), .Q(
        WX2148), .QN(n4162) );
  SDFFX1 DFF_330_Q_reg ( .D(WX2149), .SI(WX2148), .SE(n4587), .CLK(n4966), .Q(
        WX2150), .QN(n4163) );
  SDFFX1 DFF_331_Q_reg ( .D(WX2151), .SI(WX2150), .SE(n4586), .CLK(n4966), .Q(
        WX2152), .QN(n4164) );
  SDFFX1 DFF_332_Q_reg ( .D(WX2153), .SI(WX2152), .SE(n4586), .CLK(n4966), .Q(
        WX2154), .QN(n4165) );
  SDFFX1 DFF_333_Q_reg ( .D(WX2155), .SI(WX2154), .SE(n4585), .CLK(n4967), .Q(
        WX2156), .QN(n4166) );
  SDFFX1 DFF_334_Q_reg ( .D(WX2157), .SI(WX2156), .SE(n4585), .CLK(n4967), .Q(
        WX2158), .QN(n4167) );
  SDFFX1 DFF_335_Q_reg ( .D(WX2159), .SI(WX2158), .SE(n4584), .CLK(n4967), .Q(
        WX2160), .QN(n3957) );
  SDFFX1 DFF_336_Q_reg ( .D(WX2161), .SI(WX2160), .SE(n4584), .CLK(n4967), .Q(
        WX2162), .QN(n4168) );
  SDFFX1 DFF_337_Q_reg ( .D(WX2163), .SI(WX2162), .SE(n4350), .CLK(n5085), .Q(
        WX2164), .QN(n4169) );
  SDFFX1 DFF_338_Q_reg ( .D(WX2165), .SI(WX2164), .SE(n4350), .CLK(n5085), .Q(
        WX2166), .QN(n4170) );
  SDFFX1 DFF_339_Q_reg ( .D(WX2167), .SI(WX2166), .SE(n4349), .CLK(n5085), .Q(
        WX2168), .QN(n4171) );
  SDFFX1 DFF_340_Q_reg ( .D(WX2169), .SI(WX2168), .SE(n4349), .CLK(n5085), .Q(
        WX2170), .QN(n3958) );
  SDFFX1 DFF_341_Q_reg ( .D(WX2171), .SI(WX2170), .SE(n4348), .CLK(n5086), .Q(
        test_so19) );
  SDFFX1 DFF_342_Q_reg ( .D(WX2173), .SI(test_si20), .SE(n4348), .CLK(n5086), 
        .Q(WX2174), .QN(n4172) );
  SDFFX1 DFF_343_Q_reg ( .D(WX2175), .SI(WX2174), .SE(n4347), .CLK(n5086), .Q(
        WX2176), .QN(n4173) );
  SDFFX1 DFF_344_Q_reg ( .D(WX2177), .SI(WX2176), .SE(n4347), .CLK(n5086), .Q(
        WX2178), .QN(n4174) );
  SDFFX1 DFF_345_Q_reg ( .D(WX2179), .SI(WX2178), .SE(n4346), .CLK(n5087), .Q(
        WX2180), .QN(n4175) );
  SDFFX1 DFF_346_Q_reg ( .D(WX2181), .SI(WX2180), .SE(n4346), .CLK(n5087), .Q(
        WX2182), .QN(n4176) );
  SDFFX1 DFF_347_Q_reg ( .D(WX2183), .SI(WX2182), .SE(n4345), .CLK(n5087), .Q(
        WX2184), .QN(n3959) );
  SDFFX1 DFF_348_Q_reg ( .D(WX2185), .SI(WX2184), .SE(n4345), .CLK(n5087), .Q(
        WX2186), .QN(n4177) );
  SDFFX1 DFF_349_Q_reg ( .D(WX2187), .SI(WX2186), .SE(n4345), .CLK(n5087), .Q(
        WX2188), .QN(n4178) );
  SDFFX1 DFF_350_Q_reg ( .D(WX2189), .SI(WX2188), .SE(n4344), .CLK(n5088), .Q(
        WX2190), .QN(n4179) );
  SDFFX1 DFF_351_Q_reg ( .D(WX2191), .SI(WX2190), .SE(n4344), .CLK(n5088), .Q(
        WX2192), .QN(n3967) );
  SDFFX1 DFF_352_Q_reg ( .D(WX2557), .SI(WX2192), .SE(n4357), .CLK(n5081), .Q(
        CRC_OUT_8_0), .QN(DFF_352_n1) );
  SDFFX1 DFF_353_Q_reg ( .D(WX2559), .SI(CRC_OUT_8_0), .SE(n4356), .CLK(n5082), 
        .Q(CRC_OUT_8_1), .QN(DFF_353_n1) );
  SDFFX1 DFF_354_Q_reg ( .D(WX2561), .SI(CRC_OUT_8_1), .SE(n4356), .CLK(n5082), 
        .Q(CRC_OUT_8_2), .QN(DFF_354_n1) );
  SDFFX1 DFF_355_Q_reg ( .D(WX2563), .SI(CRC_OUT_8_2), .SE(n4356), .CLK(n5082), 
        .Q(CRC_OUT_8_3), .QN(DFF_355_n1) );
  SDFFX1 DFF_356_Q_reg ( .D(WX2565), .SI(CRC_OUT_8_3), .SE(n4356), .CLK(n5082), 
        .Q(CRC_OUT_8_4), .QN(DFF_356_n1) );
  SDFFX1 DFF_357_Q_reg ( .D(WX2567), .SI(CRC_OUT_8_4), .SE(n4356), .CLK(n5082), 
        .Q(CRC_OUT_8_5), .QN(DFF_357_n1) );
  SDFFX1 DFF_358_Q_reg ( .D(WX2569), .SI(CRC_OUT_8_5), .SE(n4356), .CLK(n5082), 
        .Q(CRC_OUT_8_6), .QN(DFF_358_n1) );
  SDFFX1 DFF_359_Q_reg ( .D(WX2571), .SI(CRC_OUT_8_6), .SE(n4355), .CLK(n5082), 
        .Q(test_so20) );
  SDFFX1 DFF_360_Q_reg ( .D(WX2573), .SI(test_si21), .SE(n4355), .CLK(n5082), 
        .Q(CRC_OUT_8_8), .QN(DFF_360_n1) );
  SDFFX1 DFF_361_Q_reg ( .D(WX2575), .SI(CRC_OUT_8_8), .SE(n4355), .CLK(n5082), 
        .Q(CRC_OUT_8_9), .QN(DFF_361_n1) );
  SDFFX1 DFF_362_Q_reg ( .D(WX2577), .SI(CRC_OUT_8_9), .SE(n4355), .CLK(n5082), 
        .Q(CRC_OUT_8_10), .QN(DFF_362_n1) );
  SDFFX1 DFF_363_Q_reg ( .D(WX2579), .SI(CRC_OUT_8_10), .SE(n4355), .CLK(n5082), .Q(CRC_OUT_8_11), .QN(DFF_363_n1) );
  SDFFX1 DFF_364_Q_reg ( .D(WX2581), .SI(CRC_OUT_8_11), .SE(n4355), .CLK(n5082), .Q(CRC_OUT_8_12), .QN(DFF_364_n1) );
  SDFFX1 DFF_365_Q_reg ( .D(WX2583), .SI(CRC_OUT_8_12), .SE(n4354), .CLK(n5083), .Q(CRC_OUT_8_13), .QN(DFF_365_n1) );
  SDFFX1 DFF_366_Q_reg ( .D(WX2585), .SI(CRC_OUT_8_13), .SE(n4354), .CLK(n5083), .Q(CRC_OUT_8_14), .QN(DFF_366_n1) );
  SDFFX1 DFF_367_Q_reg ( .D(WX2587), .SI(CRC_OUT_8_14), .SE(n4354), .CLK(n5083), .Q(CRC_OUT_8_15), .QN(DFF_367_n1) );
  SDFFX1 DFF_368_Q_reg ( .D(WX2589), .SI(CRC_OUT_8_15), .SE(n4354), .CLK(n5083), .Q(CRC_OUT_8_16), .QN(DFF_368_n1) );
  SDFFX1 DFF_369_Q_reg ( .D(WX2591), .SI(CRC_OUT_8_16), .SE(n4354), .CLK(n5083), .Q(CRC_OUT_8_17), .QN(DFF_369_n1) );
  SDFFX1 DFF_370_Q_reg ( .D(WX2593), .SI(CRC_OUT_8_17), .SE(n4354), .CLK(n5083), .Q(CRC_OUT_8_18), .QN(DFF_370_n1) );
  SDFFX1 DFF_371_Q_reg ( .D(WX2595), .SI(CRC_OUT_8_18), .SE(n4353), .CLK(n5083), .Q(CRC_OUT_8_19), .QN(DFF_371_n1) );
  SDFFX1 DFF_372_Q_reg ( .D(WX2597), .SI(CRC_OUT_8_19), .SE(n4353), .CLK(n5083), .Q(CRC_OUT_8_20), .QN(DFF_372_n1) );
  SDFFX1 DFF_373_Q_reg ( .D(WX2599), .SI(CRC_OUT_8_20), .SE(n4353), .CLK(n5083), .Q(CRC_OUT_8_21), .QN(DFF_373_n1) );
  SDFFX1 DFF_374_Q_reg ( .D(WX2601), .SI(CRC_OUT_8_21), .SE(n4353), .CLK(n5083), .Q(CRC_OUT_8_22), .QN(DFF_374_n1) );
  SDFFX1 DFF_375_Q_reg ( .D(WX2603), .SI(CRC_OUT_8_22), .SE(n4353), .CLK(n5083), .Q(CRC_OUT_8_23), .QN(DFF_375_n1) );
  SDFFX1 DFF_376_Q_reg ( .D(WX2605), .SI(CRC_OUT_8_23), .SE(n4353), .CLK(n5083), .Q(CRC_OUT_8_24), .QN(DFF_376_n1) );
  SDFFX1 DFF_377_Q_reg ( .D(WX2607), .SI(CRC_OUT_8_24), .SE(n4352), .CLK(n5084), .Q(test_so21) );
  SDFFX1 DFF_378_Q_reg ( .D(WX2609), .SI(test_si22), .SE(n4352), .CLK(n5084), 
        .Q(CRC_OUT_8_26), .QN(DFF_378_n1) );
  SDFFX1 DFF_379_Q_reg ( .D(WX2611), .SI(CRC_OUT_8_26), .SE(n4352), .CLK(n5084), .Q(CRC_OUT_8_27), .QN(DFF_379_n1) );
  SDFFX1 DFF_380_Q_reg ( .D(WX2613), .SI(CRC_OUT_8_27), .SE(n4352), .CLK(n5084), .Q(CRC_OUT_8_28), .QN(DFF_380_n1) );
  SDFFX1 DFF_381_Q_reg ( .D(WX2615), .SI(CRC_OUT_8_28), .SE(n4352), .CLK(n5084), .Q(CRC_OUT_8_29), .QN(DFF_381_n1) );
  SDFFX1 DFF_382_Q_reg ( .D(WX2617), .SI(CRC_OUT_8_29), .SE(n4352), .CLK(n5084), .Q(CRC_OUT_8_30), .QN(DFF_382_n1) );
  SDFFX1 DFF_383_Q_reg ( .D(WX2619), .SI(CRC_OUT_8_30), .SE(n4579), .CLK(n4969), .Q(CRC_OUT_8_31), .QN(DFF_383_n1) );
  SDFFX1 DFF_384_Q_reg ( .D(n33), .SI(CRC_OUT_8_31), .SE(n4579), .CLK(n4969), 
        .Q(WX3071), .QN(n3937) );
  SDFFX1 DFF_385_Q_reg ( .D(n34), .SI(WX3071), .SE(n4574), .CLK(n4972), .Q(
        n8644) );
  SDFFX1 DFF_386_Q_reg ( .D(n35), .SI(n8644), .SE(n4574), .CLK(n4972), .Q(
        n8643) );
  SDFFX1 DFF_387_Q_reg ( .D(n36), .SI(n8643), .SE(n4574), .CLK(n4972), .Q(
        n8642) );
  SDFFX1 DFF_388_Q_reg ( .D(n37), .SI(n8642), .SE(n4575), .CLK(n4972), .Q(
        n8641) );
  SDFFX1 DFF_389_Q_reg ( .D(n38), .SI(n8641), .SE(n4575), .CLK(n4972), .Q(
        n8640) );
  SDFFX1 DFF_390_Q_reg ( .D(n39), .SI(n8640), .SE(n4575), .CLK(n4972), .Q(
        n8639) );
  SDFFX1 DFF_391_Q_reg ( .D(n40), .SI(n8639), .SE(n4575), .CLK(n4972), .Q(
        n8638) );
  SDFFX1 DFF_392_Q_reg ( .D(n41), .SI(n8638), .SE(n4575), .CLK(n4971), .Q(
        n8637) );
  SDFFX1 DFF_393_Q_reg ( .D(n42), .SI(n8637), .SE(n4575), .CLK(n4971), .Q(
        n8636) );
  SDFFX1 DFF_394_Q_reg ( .D(n43), .SI(n8636), .SE(n4576), .CLK(n4971), .Q(
        n8635) );
  SDFFX1 DFF_395_Q_reg ( .D(n44), .SI(n8635), .SE(n4576), .CLK(n4971), .Q(
        test_so22) );
  SDFFX1 DFF_396_Q_reg ( .D(n45), .SI(test_si23), .SE(n4576), .CLK(n4971), .Q(
        n8632) );
  SDFFX1 DFF_397_Q_reg ( .D(n46), .SI(n8632), .SE(n4576), .CLK(n4971), .Q(
        n8631) );
  SDFFX1 DFF_398_Q_reg ( .D(n47), .SI(n8631), .SE(n4576), .CLK(n4971), .Q(
        n8630) );
  SDFFX1 DFF_399_Q_reg ( .D(n48), .SI(n8630), .SE(n4576), .CLK(n4971), .Q(
        n8629) );
  SDFFX1 DFF_400_Q_reg ( .D(n49), .SI(n8629), .SE(n4577), .CLK(n4971), .Q(
        n8628) );
  SDFFX1 DFF_401_Q_reg ( .D(n50), .SI(n8628), .SE(n4577), .CLK(n4971), .Q(
        n8627) );
  SDFFX1 DFF_402_Q_reg ( .D(n51), .SI(n8627), .SE(n4577), .CLK(n4971), .Q(
        n8626) );
  SDFFX1 DFF_403_Q_reg ( .D(n52), .SI(n8626), .SE(n4577), .CLK(n4971), .Q(
        n8625) );
  SDFFX1 DFF_404_Q_reg ( .D(n53), .SI(n8625), .SE(n4577), .CLK(n4970), .Q(
        n8624) );
  SDFFX1 DFF_405_Q_reg ( .D(n54), .SI(n8624), .SE(n4577), .CLK(n4970), .Q(
        n8623) );
  SDFFX1 DFF_406_Q_reg ( .D(n55), .SI(n8623), .SE(n4578), .CLK(n4970), .Q(
        n8622) );
  SDFFX1 DFF_407_Q_reg ( .D(n56), .SI(n8622), .SE(n4578), .CLK(n4970), .Q(
        n8621) );
  SDFFX1 DFF_408_Q_reg ( .D(n57), .SI(n8621), .SE(n4578), .CLK(n4970), .Q(
        n8620) );
  SDFFX1 DFF_409_Q_reg ( .D(n58), .SI(n8620), .SE(n4578), .CLK(n4970), .Q(
        n8619) );
  SDFFX1 DFF_410_Q_reg ( .D(n59), .SI(n8619), .SE(n4578), .CLK(n4970), .Q(
        n8618) );
  SDFFX1 DFF_411_Q_reg ( .D(n60), .SI(n8618), .SE(n4578), .CLK(n4970), .Q(
        n8617) );
  SDFFX1 DFF_412_Q_reg ( .D(n61), .SI(n8617), .SE(n4579), .CLK(n4970), .Q(
        n8616) );
  SDFFX1 DFF_413_Q_reg ( .D(n62), .SI(n8616), .SE(n4579), .CLK(n4970), .Q(
        test_so23) );
  SDFFX1 DFF_414_Q_reg ( .D(n63), .SI(test_si24), .SE(n4579), .CLK(n4970), .Q(
        n8613) );
  SDFFX1 DFF_415_Q_reg ( .D(WX3132), .SI(n8613), .SE(n4579), .CLK(n4970), .Q(
        n8612) );
  SDFFX1 DFF_416_Q_reg ( .D(WX3230), .SI(n8612), .SE(n4574), .CLK(n4972), .Q(
        n8611), .QN(n9044) );
  SDFFX1 DFF_417_Q_reg ( .D(WX3232), .SI(n8611), .SE(n4573), .CLK(n4972), .Q(
        n8610), .QN(n9041) );
  SDFFX1 DFF_418_Q_reg ( .D(WX3234), .SI(n8610), .SE(n4573), .CLK(n4972), .Q(
        n8609), .QN(n9039) );
  SDFFX1 DFF_419_Q_reg ( .D(WX3236), .SI(n8609), .SE(n4573), .CLK(n4973), .Q(
        n8608), .QN(n9037) );
  SDFFX1 DFF_420_Q_reg ( .D(WX3238), .SI(n8608), .SE(n4573), .CLK(n4973), .Q(
        n8607), .QN(n9035) );
  SDFFX1 DFF_421_Q_reg ( .D(WX3240), .SI(n8607), .SE(n4572), .CLK(n4973), .Q(
        n8606), .QN(n9031) );
  SDFFX1 DFF_422_Q_reg ( .D(WX3242), .SI(n8606), .SE(n4572), .CLK(n4973), .Q(
        n8605), .QN(n9029) );
  SDFFX1 DFF_423_Q_reg ( .D(WX3244), .SI(n8605), .SE(n4571), .CLK(n4974), .Q(
        n8604), .QN(n9027) );
  SDFFX1 DFF_424_Q_reg ( .D(WX3246), .SI(n8604), .SE(n4571), .CLK(n4974), .Q(
        n8603), .QN(n9025) );
  SDFFX1 DFF_425_Q_reg ( .D(WX3248), .SI(n8603), .SE(n4570), .CLK(n4974), .Q(
        n8602), .QN(n9023) );
  SDFFX1 DFF_426_Q_reg ( .D(WX3250), .SI(n8602), .SE(n4570), .CLK(n4974), .Q(
        n8601), .QN(n9022) );
  SDFFX1 DFF_427_Q_reg ( .D(WX3252), .SI(n8601), .SE(n4569), .CLK(n4975), .Q(
        n8600), .QN(n9020) );
  SDFFX1 DFF_428_Q_reg ( .D(WX3254), .SI(n8600), .SE(n4568), .CLK(n4975), .Q(
        n8599), .QN(n9018) );
  SDFFX1 DFF_429_Q_reg ( .D(WX3256), .SI(n8599), .SE(n4567), .CLK(n4975), .Q(
        n8598), .QN(n9016) );
  SDFFX1 DFF_430_Q_reg ( .D(WX3258), .SI(n8598), .SE(n4567), .CLK(n4976), .Q(
        n8597), .QN(n9012) );
  SDFFX1 DFF_431_Q_reg ( .D(WX3260), .SI(n8597), .SE(n4357), .CLK(n5081), .Q(
        test_so24) );
  SDFFX1 DFF_432_Q_reg ( .D(WX3262), .SI(test_si25), .SE(n4565), .CLK(n4976), 
        .Q(WX3263) );
  SDFFX1 DFF_433_Q_reg ( .D(WX3264), .SI(WX3263), .SE(n4565), .CLK(n4976), .Q(
        WX3265) );
  SDFFX1 DFF_434_Q_reg ( .D(WX3266), .SI(WX3265), .SE(n4565), .CLK(n4977), .Q(
        WX3267) );
  SDFFX1 DFF_435_Q_reg ( .D(WX3268), .SI(WX3267), .SE(n4564), .CLK(n4977), .Q(
        WX3269) );
  SDFFX1 DFF_436_Q_reg ( .D(WX3270), .SI(WX3269), .SE(n4563), .CLK(n4977), .Q(
        WX3271) );
  SDFFX1 DFF_437_Q_reg ( .D(WX3272), .SI(WX3271), .SE(n4563), .CLK(n4978), .Q(
        WX3273) );
  SDFFX1 DFF_438_Q_reg ( .D(WX3274), .SI(WX3273), .SE(n4562), .CLK(n4978), .Q(
        WX3275) );
  SDFFX1 DFF_439_Q_reg ( .D(WX3276), .SI(WX3275), .SE(n4561), .CLK(n4978), .Q(
        WX3277) );
  SDFFX1 DFF_440_Q_reg ( .D(WX3278), .SI(WX3277), .SE(n4561), .CLK(n4979), .Q(
        WX3279) );
  SDFFX1 DFF_441_Q_reg ( .D(WX3280), .SI(WX3279), .SE(n4560), .CLK(n4979), .Q(
        WX3281) );
  SDFFX1 DFF_442_Q_reg ( .D(WX3282), .SI(WX3281), .SE(n4559), .CLK(n4979), .Q(
        WX3283) );
  SDFFX1 DFF_443_Q_reg ( .D(WX3284), .SI(WX3283), .SE(n4559), .CLK(n4980), .Q(
        WX3285) );
  SDFFX1 DFF_444_Q_reg ( .D(WX3286), .SI(WX3285), .SE(n4558), .CLK(n4980), .Q(
        WX3287) );
  SDFFX1 DFF_445_Q_reg ( .D(WX3288), .SI(WX3287), .SE(n4557), .CLK(n4980), .Q(
        WX3289) );
  SDFFX1 DFF_446_Q_reg ( .D(WX3290), .SI(WX3289), .SE(n4557), .CLK(n4981), .Q(
        WX3291) );
  SDFFX1 DFF_447_Q_reg ( .D(WX3292), .SI(WX3291), .SE(n4556), .CLK(n4981), .Q(
        WX3293) );
  SDFFX1 DFF_448_Q_reg ( .D(WX3294), .SI(WX3293), .SE(n4574), .CLK(n4972), .Q(
        WX3295), .QN(n3588) );
  SDFFX1 DFF_449_Q_reg ( .D(WX3296), .SI(WX3295), .SE(n4574), .CLK(n4972), .Q(
        test_so25), .QN(n9042) );
  SDFFX1 DFF_450_Q_reg ( .D(WX3298), .SI(test_si26), .SE(n4573), .CLK(n4973), 
        .Q(WX3299), .QN(n3681) );
  SDFFX1 DFF_451_Q_reg ( .D(WX3300), .SI(WX3299), .SE(n4573), .CLK(n4973), .Q(
        WX3301), .QN(n3680) );
  SDFFX1 DFF_452_Q_reg ( .D(WX3302), .SI(WX3301), .SE(n4572), .CLK(n4973), .Q(
        WX3303), .QN(n3679) );
  SDFFX1 DFF_453_Q_reg ( .D(WX3304), .SI(WX3303), .SE(n4572), .CLK(n4973), .Q(
        WX3305), .QN(n9033) );
  SDFFX1 DFF_454_Q_reg ( .D(WX3306), .SI(WX3305), .SE(n4572), .CLK(n4973), .Q(
        WX3307), .QN(n3678) );
  SDFFX1 DFF_455_Q_reg ( .D(WX3308), .SI(WX3307), .SE(n4571), .CLK(n4973), .Q(
        WX3309), .QN(n3677) );
  SDFFX1 DFF_456_Q_reg ( .D(WX3310), .SI(WX3309), .SE(n4571), .CLK(n4974), .Q(
        WX3311) );
  SDFFX1 DFF_457_Q_reg ( .D(WX3312), .SI(WX3311), .SE(n4570), .CLK(n4974), .Q(
        WX3313), .QN(n3675) );
  SDFFX1 DFF_458_Q_reg ( .D(WX3314), .SI(WX3313), .SE(n4570), .CLK(n4974), .Q(
        WX3315), .QN(n3674) );
  SDFFX1 DFF_459_Q_reg ( .D(WX3316), .SI(WX3315), .SE(n4569), .CLK(n4975), .Q(
        WX3317), .QN(n3673) );
  SDFFX1 DFF_460_Q_reg ( .D(WX3318), .SI(WX3317), .SE(n4568), .CLK(n4975), .Q(
        WX3319), .QN(n3672) );
  SDFFX1 DFF_461_Q_reg ( .D(WX3320), .SI(WX3319), .SE(n4568), .CLK(n4975), .Q(
        WX3321), .QN(n3671) );
  SDFFX1 DFF_462_Q_reg ( .D(WX3322), .SI(WX3321), .SE(n4567), .CLK(n4976), .Q(
        WX3323), .QN(n3670) );
  SDFFX1 DFF_463_Q_reg ( .D(WX3324), .SI(WX3323), .SE(n4566), .CLK(n4976), .Q(
        WX3325) );
  SDFFX1 DFF_464_Q_reg ( .D(WX3326), .SI(WX3325), .SE(n4566), .CLK(n4976), .Q(
        WX3327), .QN(n9009) );
  SDFFX1 DFF_465_Q_reg ( .D(WX3328), .SI(WX3327), .SE(n4565), .CLK(n4977), .Q(
        WX3329), .QN(n9007) );
  SDFFX1 DFF_466_Q_reg ( .D(WX3330), .SI(WX3329), .SE(n4564), .CLK(n4977), .Q(
        WX3331), .QN(n9005) );
  SDFFX1 DFF_467_Q_reg ( .D(WX3332), .SI(WX3331), .SE(n4564), .CLK(n4977), .Q(
        test_so26) );
  SDFFX1 DFF_468_Q_reg ( .D(WX3334), .SI(test_si27), .SE(n4563), .CLK(n4978), 
        .Q(WX3335), .QN(n9001) );
  SDFFX1 DFF_469_Q_reg ( .D(WX3336), .SI(WX3335), .SE(n4562), .CLK(n4978), .Q(
        WX3337), .QN(n8999) );
  SDFFX1 DFF_470_Q_reg ( .D(WX3338), .SI(WX3337), .SE(n4562), .CLK(n4978), .Q(
        WX3339), .QN(n8997) );
  SDFFX1 DFF_471_Q_reg ( .D(WX3340), .SI(WX3339), .SE(n4561), .CLK(n4979), .Q(
        WX3341), .QN(n8995) );
  SDFFX1 DFF_472_Q_reg ( .D(WX3342), .SI(WX3341), .SE(n4560), .CLK(n4979), .Q(
        WX3343), .QN(n8993) );
  SDFFX1 DFF_473_Q_reg ( .D(WX3344), .SI(WX3343), .SE(n4560), .CLK(n4979), .Q(
        WX3345), .QN(n8991) );
  SDFFX1 DFF_474_Q_reg ( .D(WX3346), .SI(WX3345), .SE(n4559), .CLK(n4980), .Q(
        WX3347), .QN(n8989) );
  SDFFX1 DFF_475_Q_reg ( .D(WX3348), .SI(WX3347), .SE(n4558), .CLK(n4980), .Q(
        WX3349), .QN(n8987) );
  SDFFX1 DFF_476_Q_reg ( .D(WX3350), .SI(WX3349), .SE(n4558), .CLK(n4980), .Q(
        WX3351), .QN(n8985) );
  SDFFX1 DFF_477_Q_reg ( .D(WX3352), .SI(WX3351), .SE(n4557), .CLK(n4981), .Q(
        WX3353), .QN(n8983) );
  SDFFX1 DFF_478_Q_reg ( .D(WX3354), .SI(WX3353), .SE(n4556), .CLK(n4981), .Q(
        WX3355), .QN(n8981) );
  SDFFX1 DFF_479_Q_reg ( .D(WX3356), .SI(WX3355), .SE(n4556), .CLK(n4981), .Q(
        WX3357), .QN(n8979) );
  SDFFX1 DFF_480_Q_reg ( .D(WX3358), .SI(WX3357), .SE(n4555), .CLK(n4981), .Q(
        WX3359) );
  SDFFX1 DFF_481_Q_reg ( .D(WX3360), .SI(WX3359), .SE(n4555), .CLK(n4982), .Q(
        WX3361), .QN(n9043) );
  SDFFX1 DFF_482_Q_reg ( .D(WX3362), .SI(WX3361), .SE(n4555), .CLK(n4982), .Q(
        WX3363) );
  SDFFX1 DFF_483_Q_reg ( .D(WX3364), .SI(WX3363), .SE(n4554), .CLK(n4982), .Q(
        WX3365) );
  SDFFX1 DFF_484_Q_reg ( .D(WX3366), .SI(WX3365), .SE(n4554), .CLK(n4982), .Q(
        WX3367) );
  SDFFX1 DFF_485_Q_reg ( .D(WX3368), .SI(WX3367), .SE(n4554), .CLK(n4982), .Q(
        test_so27), .QN(n9032) );
  SDFFX1 DFF_486_Q_reg ( .D(WX3370), .SI(test_si28), .SE(n4572), .CLK(n4973), 
        .Q(WX3371) );
  SDFFX1 DFF_487_Q_reg ( .D(WX3372), .SI(WX3371), .SE(n4571), .CLK(n4973), .Q(
        WX3373) );
  SDFFX1 DFF_488_Q_reg ( .D(WX3374), .SI(WX3373), .SE(n4571), .CLK(n4974), .Q(
        WX3375), .QN(n3676) );
  SDFFX1 DFF_489_Q_reg ( .D(WX3376), .SI(WX3375), .SE(n4570), .CLK(n4974), .Q(
        WX3377) );
  SDFFX1 DFF_490_Q_reg ( .D(WX3378), .SI(WX3377), .SE(n4569), .CLK(n4974), .Q(
        WX3379) );
  SDFFX1 DFF_491_Q_reg ( .D(WX3380), .SI(WX3379), .SE(n4569), .CLK(n4975), .Q(
        WX3381) );
  SDFFX1 DFF_492_Q_reg ( .D(WX3382), .SI(WX3381), .SE(n4568), .CLK(n4975), .Q(
        WX3383) );
  SDFFX1 DFF_493_Q_reg ( .D(WX3384), .SI(WX3383), .SE(n4568), .CLK(n4975), .Q(
        WX3385) );
  SDFFX1 DFF_494_Q_reg ( .D(WX3386), .SI(WX3385), .SE(n4567), .CLK(n4976), .Q(
        WX3387) );
  SDFFX1 DFF_495_Q_reg ( .D(WX3388), .SI(WX3387), .SE(n4566), .CLK(n4976), .Q(
        WX3389), .QN(n3669) );
  SDFFX1 DFF_496_Q_reg ( .D(WX3390), .SI(WX3389), .SE(n4566), .CLK(n4976), .Q(
        WX3391), .QN(n3900) );
  SDFFX1 DFF_497_Q_reg ( .D(WX3392), .SI(WX3391), .SE(n4565), .CLK(n4977), .Q(
        WX3393), .QN(n3898) );
  SDFFX1 DFF_498_Q_reg ( .D(WX3394), .SI(WX3393), .SE(n4564), .CLK(n4977), .Q(
        WX3395), .QN(n3896) );
  SDFFX1 DFF_499_Q_reg ( .D(WX3396), .SI(WX3395), .SE(n4564), .CLK(n4977), .Q(
        WX3397), .QN(n9003) );
  SDFFX1 DFF_500_Q_reg ( .D(WX3398), .SI(WX3397), .SE(n4563), .CLK(n4978), .Q(
        WX3399), .QN(n3893) );
  SDFFX1 DFF_501_Q_reg ( .D(WX3400), .SI(WX3399), .SE(n4562), .CLK(n4978), .Q(
        WX3401), .QN(n3891) );
  SDFFX1 DFF_502_Q_reg ( .D(WX3402), .SI(WX3401), .SE(n4562), .CLK(n4978), .Q(
        WX3403), .QN(n3889) );
  SDFFX1 DFF_503_Q_reg ( .D(WX3404), .SI(WX3403), .SE(n4561), .CLK(n4979), .Q(
        test_so28) );
  SDFFX1 DFF_504_Q_reg ( .D(WX3406), .SI(test_si29), .SE(n4560), .CLK(n4979), 
        .Q(WX3407), .QN(n3886) );
  SDFFX1 DFF_505_Q_reg ( .D(WX3408), .SI(WX3407), .SE(n4560), .CLK(n4979), .Q(
        WX3409), .QN(n3884) );
  SDFFX1 DFF_506_Q_reg ( .D(WX3410), .SI(WX3409), .SE(n4559), .CLK(n4980), .Q(
        WX3411), .QN(n3882) );
  SDFFX1 DFF_507_Q_reg ( .D(WX3412), .SI(WX3411), .SE(n4558), .CLK(n4980), .Q(
        WX3413), .QN(n3880) );
  SDFFX1 DFF_508_Q_reg ( .D(WX3414), .SI(WX3413), .SE(n4558), .CLK(n4980), .Q(
        WX3415), .QN(n3878) );
  SDFFX1 DFF_509_Q_reg ( .D(WX3416), .SI(WX3415), .SE(n4557), .CLK(n4981), .Q(
        WX3417), .QN(n3876) );
  SDFFX1 DFF_510_Q_reg ( .D(WX3418), .SI(WX3417), .SE(n4556), .CLK(n4981), .Q(
        WX3419), .QN(n3874) );
  SDFFX1 DFF_511_Q_reg ( .D(WX3420), .SI(WX3419), .SE(n4556), .CLK(n4981), .Q(
        WX3421), .QN(n3872) );
  SDFFX1 DFF_512_Q_reg ( .D(WX3422), .SI(WX3421), .SE(n4555), .CLK(n4982), .Q(
        WX3423), .QN(n4128) );
  SDFFX1 DFF_513_Q_reg ( .D(WX3424), .SI(WX3423), .SE(n4555), .CLK(n4982), .Q(
        WX3425), .QN(n4129) );
  SDFFX1 DFF_514_Q_reg ( .D(WX3426), .SI(WX3425), .SE(n4554), .CLK(n4982), .Q(
        WX3427), .QN(n4130) );
  SDFFX1 DFF_515_Q_reg ( .D(WX3428), .SI(WX3427), .SE(n4554), .CLK(n4982), .Q(
        WX3429), .QN(n4131) );
  SDFFX1 DFF_516_Q_reg ( .D(WX3430), .SI(WX3429), .SE(n4554), .CLK(n4982), .Q(
        WX3431), .QN(n4132) );
  SDFFX1 DFF_517_Q_reg ( .D(WX3432), .SI(WX3431), .SE(n4553), .CLK(n4982), .Q(
        WX3433), .QN(n4133) );
  SDFFX1 DFF_518_Q_reg ( .D(WX3434), .SI(WX3433), .SE(n4553), .CLK(n4982), .Q(
        WX3435), .QN(n4134) );
  SDFFX1 DFF_519_Q_reg ( .D(WX3436), .SI(WX3435), .SE(n4553), .CLK(n4983), .Q(
        WX3437), .QN(n4135) );
  SDFFX1 DFF_520_Q_reg ( .D(WX3438), .SI(WX3437), .SE(n4553), .CLK(n4983), .Q(
        test_so29) );
  SDFFX1 DFF_521_Q_reg ( .D(WX3440), .SI(test_si30), .SE(n4570), .CLK(n4974), 
        .Q(WX3441), .QN(n4136) );
  SDFFX1 DFF_522_Q_reg ( .D(WX3442), .SI(WX3441), .SE(n4569), .CLK(n4974), .Q(
        WX3443), .QN(n4137) );
  SDFFX1 DFF_523_Q_reg ( .D(WX3444), .SI(WX3443), .SE(n4569), .CLK(n4975), .Q(
        WX3445), .QN(n4138) );
  SDFFX1 DFF_524_Q_reg ( .D(WX3446), .SI(WX3445), .SE(n4568), .CLK(n4975), .Q(
        WX3447), .QN(n4139) );
  SDFFX1 DFF_525_Q_reg ( .D(WX3448), .SI(WX3447), .SE(n4567), .CLK(n4975), .Q(
        WX3449), .QN(n4140) );
  SDFFX1 DFF_526_Q_reg ( .D(WX3450), .SI(WX3449), .SE(n4567), .CLK(n4976), .Q(
        WX3451), .QN(n4141) );
  SDFFX1 DFF_527_Q_reg ( .D(WX3452), .SI(WX3451), .SE(n4566), .CLK(n4976), .Q(
        WX3453), .QN(n3954) );
  SDFFX1 DFF_528_Q_reg ( .D(WX3454), .SI(WX3453), .SE(n4566), .CLK(n4976), .Q(
        WX3455), .QN(n4142) );
  SDFFX1 DFF_529_Q_reg ( .D(WX3456), .SI(WX3455), .SE(n4565), .CLK(n4977), .Q(
        WX3457), .QN(n4143) );
  SDFFX1 DFF_530_Q_reg ( .D(WX3458), .SI(WX3457), .SE(n4564), .CLK(n4977), .Q(
        WX3459), .QN(n4144) );
  SDFFX1 DFF_531_Q_reg ( .D(WX3460), .SI(WX3459), .SE(n4563), .CLK(n4977), .Q(
        WX3461), .QN(n4145) );
  SDFFX1 DFF_532_Q_reg ( .D(WX3462), .SI(WX3461), .SE(n4563), .CLK(n4978), .Q(
        WX3463), .QN(n3955) );
  SDFFX1 DFF_533_Q_reg ( .D(WX3464), .SI(WX3463), .SE(n4562), .CLK(n4978), .Q(
        WX3465), .QN(n4146) );
  SDFFX1 DFF_534_Q_reg ( .D(WX3466), .SI(WX3465), .SE(n4561), .CLK(n4978), .Q(
        WX3467), .QN(n4147) );
  SDFFX1 DFF_535_Q_reg ( .D(WX3468), .SI(WX3467), .SE(n4561), .CLK(n4979), .Q(
        WX3469), .QN(n4148) );
  SDFFX1 DFF_536_Q_reg ( .D(WX3470), .SI(WX3469), .SE(n4560), .CLK(n4979), .Q(
        WX3471), .QN(n4149) );
  SDFFX1 DFF_537_Q_reg ( .D(WX3472), .SI(WX3471), .SE(n4559), .CLK(n4979), .Q(
        test_so30) );
  SDFFX1 DFF_538_Q_reg ( .D(WX3474), .SI(test_si31), .SE(n4559), .CLK(n4980), 
        .Q(WX3475), .QN(n4150) );
  SDFFX1 DFF_539_Q_reg ( .D(WX3476), .SI(WX3475), .SE(n4558), .CLK(n4980), .Q(
        WX3477), .QN(n3956) );
  SDFFX1 DFF_540_Q_reg ( .D(WX3478), .SI(WX3477), .SE(n4557), .CLK(n4980), .Q(
        WX3479), .QN(n4151) );
  SDFFX1 DFF_541_Q_reg ( .D(WX3480), .SI(WX3479), .SE(n4557), .CLK(n4981), .Q(
        WX3481), .QN(n4152) );
  SDFFX1 DFF_542_Q_reg ( .D(WX3482), .SI(WX3481), .SE(n4556), .CLK(n4981), .Q(
        WX3483), .QN(n4153) );
  SDFFX1 DFF_543_Q_reg ( .D(WX3484), .SI(WX3483), .SE(n4555), .CLK(n4981), .Q(
        WX3485), .QN(n3966) );
  SDFFX1 DFF_544_Q_reg ( .D(WX3850), .SI(WX3485), .SE(n4361), .CLK(n5079), .Q(
        CRC_OUT_7_0), .QN(DFF_544_n1) );
  SDFFX1 DFF_545_Q_reg ( .D(WX3852), .SI(CRC_OUT_7_0), .SE(n4361), .CLK(n5079), 
        .Q(CRC_OUT_7_1), .QN(DFF_545_n1) );
  SDFFX1 DFF_546_Q_reg ( .D(WX3854), .SI(CRC_OUT_7_1), .SE(n4361), .CLK(n5079), 
        .Q(CRC_OUT_7_2), .QN(DFF_546_n1) );
  SDFFX1 DFF_547_Q_reg ( .D(WX3856), .SI(CRC_OUT_7_2), .SE(n4361), .CLK(n5079), 
        .Q(CRC_OUT_7_3), .QN(DFF_547_n1) );
  SDFFX1 DFF_548_Q_reg ( .D(WX3858), .SI(CRC_OUT_7_3), .SE(n4360), .CLK(n5080), 
        .Q(CRC_OUT_7_4), .QN(DFF_548_n1) );
  SDFFX1 DFF_549_Q_reg ( .D(WX3860), .SI(CRC_OUT_7_4), .SE(n4360), .CLK(n5080), 
        .Q(CRC_OUT_7_5), .QN(DFF_549_n1) );
  SDFFX1 DFF_550_Q_reg ( .D(WX3862), .SI(CRC_OUT_7_5), .SE(n4360), .CLK(n5080), 
        .Q(CRC_OUT_7_6), .QN(DFF_550_n1) );
  SDFFX1 DFF_551_Q_reg ( .D(WX3864), .SI(CRC_OUT_7_6), .SE(n4360), .CLK(n5080), 
        .Q(CRC_OUT_7_7), .QN(DFF_551_n1) );
  SDFFX1 DFF_552_Q_reg ( .D(WX3866), .SI(CRC_OUT_7_7), .SE(n4360), .CLK(n5080), 
        .Q(CRC_OUT_7_8), .QN(DFF_552_n1) );
  SDFFX1 DFF_553_Q_reg ( .D(WX3868), .SI(CRC_OUT_7_8), .SE(n4360), .CLK(n5080), 
        .Q(CRC_OUT_7_9), .QN(DFF_553_n1) );
  SDFFX1 DFF_554_Q_reg ( .D(WX3870), .SI(CRC_OUT_7_9), .SE(n4359), .CLK(n5080), 
        .Q(test_so31) );
  SDFFX1 DFF_555_Q_reg ( .D(WX3872), .SI(test_si32), .SE(n4359), .CLK(n5080), 
        .Q(CRC_OUT_7_11), .QN(DFF_555_n1) );
  SDFFX1 DFF_556_Q_reg ( .D(WX3874), .SI(CRC_OUT_7_11), .SE(n4359), .CLK(n5080), .Q(CRC_OUT_7_12), .QN(DFF_556_n1) );
  SDFFX1 DFF_557_Q_reg ( .D(WX3876), .SI(CRC_OUT_7_12), .SE(n4359), .CLK(n5080), .Q(CRC_OUT_7_13), .QN(DFF_557_n1) );
  SDFFX1 DFF_558_Q_reg ( .D(WX3878), .SI(CRC_OUT_7_13), .SE(n4359), .CLK(n5080), .Q(CRC_OUT_7_14), .QN(DFF_558_n1) );
  SDFFX1 DFF_559_Q_reg ( .D(WX3880), .SI(CRC_OUT_7_14), .SE(n4359), .CLK(n5080), .Q(CRC_OUT_7_15), .QN(DFF_559_n1) );
  SDFFX1 DFF_560_Q_reg ( .D(WX3882), .SI(CRC_OUT_7_15), .SE(n4358), .CLK(n5081), .Q(CRC_OUT_7_16), .QN(DFF_560_n1) );
  SDFFX1 DFF_561_Q_reg ( .D(WX3884), .SI(CRC_OUT_7_16), .SE(n4358), .CLK(n5081), .Q(CRC_OUT_7_17), .QN(DFF_561_n1) );
  SDFFX1 DFF_562_Q_reg ( .D(WX3886), .SI(CRC_OUT_7_17), .SE(n4358), .CLK(n5081), .Q(CRC_OUT_7_18), .QN(DFF_562_n1) );
  SDFFX1 DFF_563_Q_reg ( .D(WX3888), .SI(CRC_OUT_7_18), .SE(n4358), .CLK(n5081), .Q(CRC_OUT_7_19), .QN(DFF_563_n1) );
  SDFFX1 DFF_564_Q_reg ( .D(WX3890), .SI(CRC_OUT_7_19), .SE(n4358), .CLK(n5081), .Q(CRC_OUT_7_20), .QN(DFF_564_n1) );
  SDFFX1 DFF_565_Q_reg ( .D(WX3892), .SI(CRC_OUT_7_20), .SE(n4358), .CLK(n5081), .Q(CRC_OUT_7_21), .QN(DFF_565_n1) );
  SDFFX1 DFF_566_Q_reg ( .D(WX3894), .SI(CRC_OUT_7_21), .SE(n4357), .CLK(n5081), .Q(CRC_OUT_7_22), .QN(DFF_566_n1) );
  SDFFX1 DFF_567_Q_reg ( .D(WX3896), .SI(CRC_OUT_7_22), .SE(n4357), .CLK(n5081), .Q(CRC_OUT_7_23), .QN(DFF_567_n1) );
  SDFFX1 DFF_568_Q_reg ( .D(WX3898), .SI(CRC_OUT_7_23), .SE(n4357), .CLK(n5081), .Q(CRC_OUT_7_24), .QN(DFF_568_n1) );
  SDFFX1 DFF_569_Q_reg ( .D(WX3900), .SI(CRC_OUT_7_24), .SE(n4357), .CLK(n5081), .Q(CRC_OUT_7_25), .QN(DFF_569_n1) );
  SDFFX1 DFF_570_Q_reg ( .D(WX3902), .SI(CRC_OUT_7_25), .SE(n4553), .CLK(n4983), .Q(CRC_OUT_7_26), .QN(DFF_570_n1) );
  SDFFX1 DFF_571_Q_reg ( .D(WX3904), .SI(CRC_OUT_7_26), .SE(n4553), .CLK(n4983), .Q(test_so32) );
  SDFFX1 DFF_572_Q_reg ( .D(WX3906), .SI(test_si33), .SE(n4552), .CLK(n4983), 
        .Q(CRC_OUT_7_28), .QN(DFF_572_n1) );
  SDFFX1 DFF_573_Q_reg ( .D(WX3908), .SI(CRC_OUT_7_28), .SE(n4552), .CLK(n4983), .Q(CRC_OUT_7_29), .QN(DFF_573_n1) );
  SDFFX1 DFF_574_Q_reg ( .D(WX3910), .SI(CRC_OUT_7_29), .SE(n4552), .CLK(n4983), .Q(CRC_OUT_7_30), .QN(DFF_574_n1) );
  SDFFX1 DFF_575_Q_reg ( .D(WX3912), .SI(CRC_OUT_7_30), .SE(n4552), .CLK(n4983), .Q(CRC_OUT_7_31), .QN(DFF_575_n1) );
  SDFFX1 DFF_576_Q_reg ( .D(n64), .SI(CRC_OUT_7_31), .SE(n4552), .CLK(n4983), 
        .Q(WX4364), .QN(n3936) );
  SDFFX1 DFF_577_Q_reg ( .D(n65), .SI(WX4364), .SE(n4547), .CLK(n4986), .Q(
        n8586) );
  SDFFX1 DFF_578_Q_reg ( .D(n66), .SI(n8586), .SE(n4547), .CLK(n4986), .Q(
        n8585) );
  SDFFX1 DFF_579_Q_reg ( .D(n67), .SI(n8585), .SE(n4547), .CLK(n4986), .Q(
        n8584) );
  SDFFX1 DFF_580_Q_reg ( .D(n68), .SI(n8584), .SE(n4547), .CLK(n4986), .Q(
        n8583) );
  SDFFX1 DFF_581_Q_reg ( .D(n69), .SI(n8583), .SE(n4547), .CLK(n4985), .Q(
        n8582) );
  SDFFX1 DFF_582_Q_reg ( .D(n70), .SI(n8582), .SE(n4547), .CLK(n4985), .Q(
        n8581) );
  SDFFX1 DFF_583_Q_reg ( .D(n71), .SI(n8581), .SE(n4548), .CLK(n4985), .Q(
        n8580) );
  SDFFX1 DFF_584_Q_reg ( .D(n72), .SI(n8580), .SE(n4548), .CLK(n4985), .Q(
        n8579) );
  SDFFX1 DFF_585_Q_reg ( .D(n73), .SI(n8579), .SE(n4548), .CLK(n4985), .Q(
        n8578) );
  SDFFX1 DFF_586_Q_reg ( .D(n74), .SI(n8578), .SE(n4548), .CLK(n4985), .Q(
        n8577) );
  SDFFX1 DFF_587_Q_reg ( .D(n75), .SI(n8577), .SE(n4548), .CLK(n4985), .Q(
        n8576) );
  SDFFX1 DFF_588_Q_reg ( .D(n76), .SI(n8576), .SE(n4548), .CLK(n4985), .Q(
        test_so33) );
  SDFFX1 DFF_589_Q_reg ( .D(n77), .SI(test_si34), .SE(n4549), .CLK(n4985), .Q(
        n8573) );
  SDFFX1 DFF_590_Q_reg ( .D(n78), .SI(n8573), .SE(n4549), .CLK(n4985), .Q(
        n8572) );
  SDFFX1 DFF_591_Q_reg ( .D(n79), .SI(n8572), .SE(n4549), .CLK(n4985), .Q(
        n8571) );
  SDFFX1 DFF_592_Q_reg ( .D(n80), .SI(n8571), .SE(n4549), .CLK(n4985), .Q(
        n8570) );
  SDFFX1 DFF_593_Q_reg ( .D(n81), .SI(n8570), .SE(n4549), .CLK(n4984), .Q(
        n8569) );
  SDFFX1 DFF_594_Q_reg ( .D(n82), .SI(n8569), .SE(n4549), .CLK(n4984), .Q(
        n8568) );
  SDFFX1 DFF_595_Q_reg ( .D(n83), .SI(n8568), .SE(n4550), .CLK(n4984), .Q(
        n8567) );
  SDFFX1 DFF_596_Q_reg ( .D(n84), .SI(n8567), .SE(n4550), .CLK(n4984), .Q(
        n8566) );
  SDFFX1 DFF_597_Q_reg ( .D(n85), .SI(n8566), .SE(n4550), .CLK(n4984), .Q(
        n8565) );
  SDFFX1 DFF_598_Q_reg ( .D(n86), .SI(n8565), .SE(n4550), .CLK(n4984), .Q(
        n8564) );
  SDFFX1 DFF_599_Q_reg ( .D(n87), .SI(n8564), .SE(n4550), .CLK(n4984), .Q(
        n8563) );
  SDFFX1 DFF_600_Q_reg ( .D(n88), .SI(n8563), .SE(n4550), .CLK(n4984), .Q(
        n8562) );
  SDFFX1 DFF_601_Q_reg ( .D(n89), .SI(n8562), .SE(n4551), .CLK(n4984), .Q(
        n8561) );
  SDFFX1 DFF_602_Q_reg ( .D(n90), .SI(n8561), .SE(n4551), .CLK(n4984), .Q(
        n8560) );
  SDFFX1 DFF_603_Q_reg ( .D(n91), .SI(n8560), .SE(n4551), .CLK(n4984), .Q(
        n8559) );
  SDFFX1 DFF_604_Q_reg ( .D(n92), .SI(n8559), .SE(n4551), .CLK(n4984), .Q(
        n8558) );
  SDFFX1 DFF_605_Q_reg ( .D(n93), .SI(n8558), .SE(n4551), .CLK(n4983), .Q(
        test_so34) );
  SDFFX1 DFF_606_Q_reg ( .D(n94), .SI(test_si35), .SE(n4551), .CLK(n4983), .Q(
        n8555) );
  SDFFX1 DFF_607_Q_reg ( .D(WX4425), .SI(n8555), .SE(n4552), .CLK(n4983), .Q(
        n8554) );
  SDFFX1 DFF_608_Q_reg ( .D(WX4523), .SI(n8554), .SE(n4546), .CLK(n4986), .Q(
        n8553), .QN(n8977) );
  SDFFX1 DFF_609_Q_reg ( .D(WX4525), .SI(n8553), .SE(n4546), .CLK(n4986), .Q(
        n8552), .QN(n8974) );
  SDFFX1 DFF_610_Q_reg ( .D(WX4527), .SI(n8552), .SE(n4546), .CLK(n4986), .Q(
        n8551), .QN(n8973) );
  SDFFX1 DFF_611_Q_reg ( .D(WX4529), .SI(n8551), .SE(n4361), .CLK(n5079), .Q(
        n8550), .QN(n8972) );
  SDFFX1 DFF_612_Q_reg ( .D(WX4531), .SI(n8550), .SE(n4544), .CLK(n4987), .Q(
        n8549), .QN(n8971) );
  SDFFX1 DFF_613_Q_reg ( .D(WX4533), .SI(n8549), .SE(n4544), .CLK(n4987), .Q(
        n8548), .QN(n8970) );
  SDFFX1 DFF_614_Q_reg ( .D(WX4535), .SI(n8548), .SE(n4543), .CLK(n4988), .Q(
        n8547), .QN(n8969) );
  SDFFX1 DFF_615_Q_reg ( .D(WX4537), .SI(n8547), .SE(n4543), .CLK(n4988), .Q(
        n8546), .QN(n8968) );
  SDFFX1 DFF_616_Q_reg ( .D(WX4539), .SI(n8546), .SE(n4542), .CLK(n4988), .Q(
        n8545), .QN(n8967) );
  SDFFX1 DFF_617_Q_reg ( .D(WX4541), .SI(n8545), .SE(n4542), .CLK(n4988), .Q(
        n8544), .QN(n8966) );
  SDFFX1 DFF_618_Q_reg ( .D(WX4543), .SI(n8544), .SE(n4540), .CLK(n4989), .Q(
        n8543), .QN(n8965) );
  SDFFX1 DFF_619_Q_reg ( .D(WX4545), .SI(n8543), .SE(n4540), .CLK(n4989), .Q(
        n8542), .QN(n8964) );
  SDFFX1 DFF_620_Q_reg ( .D(WX4547), .SI(n8542), .SE(n4539), .CLK(n4990), .Q(
        n8541), .QN(n8963) );
  SDFFX1 DFF_621_Q_reg ( .D(WX4549), .SI(n8541), .SE(n4539), .CLK(n4990), .Q(
        n8540), .QN(n8962) );
  SDFFX1 DFF_622_Q_reg ( .D(WX4551), .SI(n8540), .SE(n4361), .CLK(n5079), .Q(
        test_so35) );
  SDFFX1 DFF_623_Q_reg ( .D(WX4553), .SI(test_si36), .SE(n4537), .CLK(n4990), 
        .Q(n8537), .QN(n8961) );
  SDFFX1 DFF_624_Q_reg ( .D(WX4555), .SI(n8537), .SE(n4537), .CLK(n4991), .Q(
        WX4556) );
  SDFFX1 DFF_625_Q_reg ( .D(WX4557), .SI(WX4556), .SE(n4536), .CLK(n4991), .Q(
        WX4558) );
  SDFFX1 DFF_626_Q_reg ( .D(WX4559), .SI(WX4558), .SE(n4536), .CLK(n4991), .Q(
        WX4560) );
  SDFFX1 DFF_627_Q_reg ( .D(WX4561), .SI(WX4560), .SE(n4535), .CLK(n4992), .Q(
        WX4562) );
  SDFFX1 DFF_628_Q_reg ( .D(WX4563), .SI(WX4562), .SE(n4534), .CLK(n4992), .Q(
        WX4564) );
  SDFFX1 DFF_629_Q_reg ( .D(WX4565), .SI(WX4564), .SE(n4534), .CLK(n4992), .Q(
        WX4566) );
  SDFFX1 DFF_630_Q_reg ( .D(WX4567), .SI(WX4566), .SE(n4533), .CLK(n4993), .Q(
        WX4568) );
  SDFFX1 DFF_631_Q_reg ( .D(WX4569), .SI(WX4568), .SE(n4532), .CLK(n4993), .Q(
        WX4570) );
  SDFFX1 DFF_632_Q_reg ( .D(WX4571), .SI(WX4570), .SE(n4532), .CLK(n4993), .Q(
        WX4572) );
  SDFFX1 DFF_633_Q_reg ( .D(WX4573), .SI(WX4572), .SE(n4531), .CLK(n4994), .Q(
        WX4574) );
  SDFFX1 DFF_634_Q_reg ( .D(WX4575), .SI(WX4574), .SE(n4530), .CLK(n4994), .Q(
        WX4576) );
  SDFFX1 DFF_635_Q_reg ( .D(WX4577), .SI(WX4576), .SE(n4530), .CLK(n4994), .Q(
        WX4578) );
  SDFFX1 DFF_636_Q_reg ( .D(WX4579), .SI(WX4578), .SE(n4529), .CLK(n4995), .Q(
        WX4580) );
  SDFFX1 DFF_637_Q_reg ( .D(WX4581), .SI(WX4580), .SE(n4528), .CLK(n4995), .Q(
        WX4582) );
  SDFFX1 DFF_638_Q_reg ( .D(WX4583), .SI(WX4582), .SE(n4528), .CLK(n4995), .Q(
        WX4584) );
  SDFFX1 DFF_639_Q_reg ( .D(WX4585), .SI(WX4584), .SE(n4527), .CLK(n4996), .Q(
        test_so36) );
  SDFFX1 DFF_640_Q_reg ( .D(WX4587), .SI(test_si37), .SE(n4546), .CLK(n4986), 
        .Q(WX4588), .QN(n3587) );
  SDFFX1 DFF_641_Q_reg ( .D(WX4589), .SI(WX4588), .SE(n4546), .CLK(n4986), .Q(
        WX4590), .QN(n8976) );
  SDFFX1 DFF_642_Q_reg ( .D(WX4591), .SI(WX4590), .SE(n4546), .CLK(n4986), .Q(
        WX4592), .QN(n3668) );
  SDFFX1 DFF_643_Q_reg ( .D(WX4593), .SI(WX4592), .SE(n4545), .CLK(n4986), .Q(
        WX4594) );
  SDFFX1 DFF_644_Q_reg ( .D(WX4595), .SI(WX4594), .SE(n4545), .CLK(n4987), .Q(
        WX4596), .QN(n3666) );
  SDFFX1 DFF_645_Q_reg ( .D(WX4597), .SI(WX4596), .SE(n4544), .CLK(n4987), .Q(
        WX4598), .QN(n3665) );
  SDFFX1 DFF_646_Q_reg ( .D(WX4599), .SI(WX4598), .SE(n4544), .CLK(n4987), .Q(
        WX4600), .QN(n3664) );
  SDFFX1 DFF_647_Q_reg ( .D(WX4601), .SI(WX4600), .SE(n4543), .CLK(n4988), .Q(
        WX4602), .QN(n3663) );
  SDFFX1 DFF_648_Q_reg ( .D(WX4603), .SI(WX4602), .SE(n4542), .CLK(n4988), .Q(
        WX4604), .QN(n3662) );
  SDFFX1 DFF_649_Q_reg ( .D(WX4605), .SI(WX4604), .SE(n4541), .CLK(n4988), .Q(
        WX4606), .QN(n3661) );
  SDFFX1 DFF_650_Q_reg ( .D(WX4607), .SI(WX4606), .SE(n4541), .CLK(n4989), .Q(
        WX4608), .QN(n3660) );
  SDFFX1 DFF_651_Q_reg ( .D(WX4609), .SI(WX4608), .SE(n4540), .CLK(n4989), .Q(
        WX4610), .QN(n3659) );
  SDFFX1 DFF_652_Q_reg ( .D(WX4611), .SI(WX4610), .SE(n4540), .CLK(n4989), .Q(
        WX4612), .QN(n3658) );
  SDFFX1 DFF_653_Q_reg ( .D(WX4613), .SI(WX4612), .SE(n4539), .CLK(n4990), .Q(
        WX4614), .QN(n3657) );
  SDFFX1 DFF_654_Q_reg ( .D(WX4615), .SI(WX4614), .SE(n4538), .CLK(n4990), .Q(
        WX4616) );
  SDFFX1 DFF_655_Q_reg ( .D(WX4617), .SI(WX4616), .SE(n4538), .CLK(n4990), .Q(
        WX4618), .QN(n3655) );
  SDFFX1 DFF_656_Q_reg ( .D(WX4619), .SI(WX4618), .SE(n4537), .CLK(n4991), .Q(
        test_so37) );
  SDFFX1 DFF_657_Q_reg ( .D(WX4621), .SI(test_si38), .SE(n4536), .CLK(n4991), 
        .Q(WX4622), .QN(n8959) );
  SDFFX1 DFF_658_Q_reg ( .D(WX4623), .SI(WX4622), .SE(n4536), .CLK(n4991), .Q(
        WX4624), .QN(n8958) );
  SDFFX1 DFF_659_Q_reg ( .D(WX4625), .SI(WX4624), .SE(n4535), .CLK(n4992), .Q(
        WX4626), .QN(n8957) );
  SDFFX1 DFF_660_Q_reg ( .D(WX4627), .SI(WX4626), .SE(n4534), .CLK(n4992), .Q(
        WX4628), .QN(n8956) );
  SDFFX1 DFF_661_Q_reg ( .D(WX4629), .SI(WX4628), .SE(n4534), .CLK(n4992), .Q(
        WX4630), .QN(n8955) );
  SDFFX1 DFF_662_Q_reg ( .D(WX4631), .SI(WX4630), .SE(n4533), .CLK(n4993), .Q(
        WX4632), .QN(n8954) );
  SDFFX1 DFF_663_Q_reg ( .D(WX4633), .SI(WX4632), .SE(n4532), .CLK(n4993), .Q(
        WX4634), .QN(n8953) );
  SDFFX1 DFF_664_Q_reg ( .D(WX4635), .SI(WX4634), .SE(n4532), .CLK(n4993), .Q(
        WX4636), .QN(n8952) );
  SDFFX1 DFF_665_Q_reg ( .D(WX4637), .SI(WX4636), .SE(n4531), .CLK(n4994), .Q(
        WX4638), .QN(n8951) );
  SDFFX1 DFF_666_Q_reg ( .D(WX4639), .SI(WX4638), .SE(n4530), .CLK(n4994), .Q(
        WX4640), .QN(n8950) );
  SDFFX1 DFF_667_Q_reg ( .D(WX4641), .SI(WX4640), .SE(n4530), .CLK(n4994), .Q(
        WX4642), .QN(n8949) );
  SDFFX1 DFF_668_Q_reg ( .D(WX4643), .SI(WX4642), .SE(n4529), .CLK(n4995), .Q(
        WX4644), .QN(n8948) );
  SDFFX1 DFF_669_Q_reg ( .D(WX4645), .SI(WX4644), .SE(n4528), .CLK(n4995), .Q(
        WX4646), .QN(n8947) );
  SDFFX1 DFF_670_Q_reg ( .D(WX4647), .SI(WX4646), .SE(n4528), .CLK(n4995), .Q(
        WX4648), .QN(n8946) );
  SDFFX1 DFF_671_Q_reg ( .D(WX4649), .SI(WX4648), .SE(n4527), .CLK(n4996), .Q(
        WX4650), .QN(n8945) );
  SDFFX1 DFF_672_Q_reg ( .D(WX4651), .SI(WX4650), .SE(n4526), .CLK(n4996), .Q(
        WX4652) );
  SDFFX1 DFF_673_Q_reg ( .D(WX4653), .SI(WX4652), .SE(n4526), .CLK(n4996), .Q(
        test_so38), .QN(n8975) );
  SDFFX1 DFF_674_Q_reg ( .D(WX4655), .SI(test_si39), .SE(n4545), .CLK(n4986), 
        .Q(WX4656) );
  SDFFX1 DFF_675_Q_reg ( .D(WX4657), .SI(WX4656), .SE(n4545), .CLK(n4987), .Q(
        WX4658), .QN(n3667) );
  SDFFX1 DFF_676_Q_reg ( .D(WX4659), .SI(WX4658), .SE(n4545), .CLK(n4987), .Q(
        WX4660) );
  SDFFX1 DFF_677_Q_reg ( .D(WX4661), .SI(WX4660), .SE(n4544), .CLK(n4987), .Q(
        WX4662) );
  SDFFX1 DFF_678_Q_reg ( .D(WX4663), .SI(WX4662), .SE(n4543), .CLK(n4987), .Q(
        WX4664) );
  SDFFX1 DFF_679_Q_reg ( .D(WX4665), .SI(WX4664), .SE(n4543), .CLK(n4988), .Q(
        WX4666) );
  SDFFX1 DFF_680_Q_reg ( .D(WX4667), .SI(WX4666), .SE(n4542), .CLK(n4988), .Q(
        WX4668) );
  SDFFX1 DFF_681_Q_reg ( .D(WX4669), .SI(WX4668), .SE(n4541), .CLK(n4988), .Q(
        WX4670) );
  SDFFX1 DFF_682_Q_reg ( .D(WX4671), .SI(WX4670), .SE(n4541), .CLK(n4989), .Q(
        WX4672) );
  SDFFX1 DFF_683_Q_reg ( .D(WX4673), .SI(WX4672), .SE(n4540), .CLK(n4989), .Q(
        WX4674) );
  SDFFX1 DFF_684_Q_reg ( .D(WX4675), .SI(WX4674), .SE(n4539), .CLK(n4989), .Q(
        WX4676) );
  SDFFX1 DFF_685_Q_reg ( .D(WX4677), .SI(WX4676), .SE(n4539), .CLK(n4990), .Q(
        WX4678) );
  SDFFX1 DFF_686_Q_reg ( .D(WX4679), .SI(WX4678), .SE(n4538), .CLK(n4990), .Q(
        WX4680), .QN(n3656) );
  SDFFX1 DFF_687_Q_reg ( .D(WX4681), .SI(WX4680), .SE(n4538), .CLK(n4990), .Q(
        WX4682) );
  SDFFX1 DFF_688_Q_reg ( .D(WX4683), .SI(WX4682), .SE(n4537), .CLK(n4991), .Q(
        WX4684), .QN(n8960) );
  SDFFX1 DFF_689_Q_reg ( .D(WX4685), .SI(WX4684), .SE(n4536), .CLK(n4991), .Q(
        WX4686), .QN(n3869) );
  SDFFX1 DFF_690_Q_reg ( .D(WX4687), .SI(WX4686), .SE(n4535), .CLK(n4991), .Q(
        test_so39) );
  SDFFX1 DFF_691_Q_reg ( .D(WX4689), .SI(test_si40), .SE(n4535), .CLK(n4992), 
        .Q(WX4690), .QN(n3866) );
  SDFFX1 DFF_692_Q_reg ( .D(WX4691), .SI(WX4690), .SE(n4534), .CLK(n4992), .Q(
        WX4692), .QN(n3864) );
  SDFFX1 DFF_693_Q_reg ( .D(WX4693), .SI(WX4692), .SE(n4533), .CLK(n4992), .Q(
        WX4694), .QN(n3862) );
  SDFFX1 DFF_694_Q_reg ( .D(WX4695), .SI(WX4694), .SE(n4533), .CLK(n4993), .Q(
        WX4696), .QN(n3860) );
  SDFFX1 DFF_695_Q_reg ( .D(WX4697), .SI(WX4696), .SE(n4532), .CLK(n4993), .Q(
        WX4698), .QN(n3858) );
  SDFFX1 DFF_696_Q_reg ( .D(WX4699), .SI(WX4698), .SE(n4531), .CLK(n4993), .Q(
        WX4700), .QN(n3856) );
  SDFFX1 DFF_697_Q_reg ( .D(WX4701), .SI(WX4700), .SE(n4531), .CLK(n4994), .Q(
        WX4702), .QN(n3854) );
  SDFFX1 DFF_698_Q_reg ( .D(WX4703), .SI(WX4702), .SE(n4530), .CLK(n4994), .Q(
        WX4704), .QN(n3852) );
  SDFFX1 DFF_699_Q_reg ( .D(WX4705), .SI(WX4704), .SE(n4529), .CLK(n4994), .Q(
        WX4706), .QN(n3850) );
  SDFFX1 DFF_700_Q_reg ( .D(WX4707), .SI(WX4706), .SE(n4529), .CLK(n4995), .Q(
        WX4708), .QN(n3848) );
  SDFFX1 DFF_701_Q_reg ( .D(WX4709), .SI(WX4708), .SE(n4528), .CLK(n4995), .Q(
        WX4710), .QN(n3846) );
  SDFFX1 DFF_702_Q_reg ( .D(WX4711), .SI(WX4710), .SE(n4527), .CLK(n4995), .Q(
        WX4712), .QN(n3844) );
  SDFFX1 DFF_703_Q_reg ( .D(WX4713), .SI(WX4712), .SE(n4527), .CLK(n4996), .Q(
        WX4714) );
  SDFFX1 DFF_704_Q_reg ( .D(WX4715), .SI(WX4714), .SE(n4526), .CLK(n4996), .Q(
        WX4716), .QN(n4101) );
  SDFFX1 DFF_705_Q_reg ( .D(WX4717), .SI(WX4716), .SE(n4526), .CLK(n4996), .Q(
        WX4718), .QN(n4102) );
  SDFFX1 DFF_706_Q_reg ( .D(WX4719), .SI(WX4718), .SE(n4526), .CLK(n4996), .Q(
        WX4720), .QN(n4103) );
  SDFFX1 DFF_707_Q_reg ( .D(WX4721), .SI(WX4720), .SE(n4526), .CLK(n4996), .Q(
        test_so40) );
  SDFFX1 DFF_708_Q_reg ( .D(WX4723), .SI(test_si41), .SE(n4545), .CLK(n4987), 
        .Q(WX4724), .QN(n4104) );
  SDFFX1 DFF_709_Q_reg ( .D(WX4725), .SI(WX4724), .SE(n4544), .CLK(n4987), .Q(
        WX4726), .QN(n4105) );
  SDFFX1 DFF_710_Q_reg ( .D(WX4727), .SI(WX4726), .SE(n4543), .CLK(n4987), .Q(
        WX4728), .QN(n4106) );
  SDFFX1 DFF_711_Q_reg ( .D(WX4729), .SI(WX4728), .SE(n4542), .CLK(n4988), .Q(
        WX4730), .QN(n4107) );
  SDFFX1 DFF_712_Q_reg ( .D(WX4731), .SI(WX4730), .SE(n4542), .CLK(n4988), .Q(
        WX4732), .QN(n4108) );
  SDFFX1 DFF_713_Q_reg ( .D(WX4733), .SI(WX4732), .SE(n4541), .CLK(n4989), .Q(
        WX4734), .QN(n4109) );
  SDFFX1 DFF_714_Q_reg ( .D(WX4735), .SI(WX4734), .SE(n4541), .CLK(n4989), .Q(
        WX4736), .QN(n4110) );
  SDFFX1 DFF_715_Q_reg ( .D(WX4737), .SI(WX4736), .SE(n4540), .CLK(n4989), .Q(
        WX4738), .QN(n4111) );
  SDFFX1 DFF_716_Q_reg ( .D(WX4739), .SI(WX4738), .SE(n4539), .CLK(n4989), .Q(
        WX4740), .QN(n4112) );
  SDFFX1 DFF_717_Q_reg ( .D(WX4741), .SI(WX4740), .SE(n4538), .CLK(n4990), .Q(
        WX4742), .QN(n4113) );
  SDFFX1 DFF_718_Q_reg ( .D(WX4743), .SI(WX4742), .SE(n4538), .CLK(n4990), .Q(
        WX4744), .QN(n4114) );
  SDFFX1 DFF_719_Q_reg ( .D(WX4745), .SI(WX4744), .SE(n4537), .CLK(n4990), .Q(
        WX4746), .QN(n3952) );
  SDFFX1 DFF_720_Q_reg ( .D(WX4747), .SI(WX4746), .SE(n4537), .CLK(n4991), .Q(
        WX4748), .QN(n4115) );
  SDFFX1 DFF_721_Q_reg ( .D(WX4749), .SI(WX4748), .SE(n4536), .CLK(n4991), .Q(
        WX4750), .QN(n4116) );
  SDFFX1 DFF_722_Q_reg ( .D(WX4751), .SI(WX4750), .SE(n4535), .CLK(n4991), .Q(
        WX4752), .QN(n4117) );
  SDFFX1 DFF_723_Q_reg ( .D(WX4753), .SI(WX4752), .SE(n4535), .CLK(n4992), .Q(
        WX4754), .QN(n4118) );
  SDFFX1 DFF_724_Q_reg ( .D(WX4755), .SI(WX4754), .SE(n4534), .CLK(n4992), .Q(
        test_so41) );
  SDFFX1 DFF_725_Q_reg ( .D(WX4757), .SI(test_si42), .SE(n4533), .CLK(n4992), 
        .Q(WX4758), .QN(n4119) );
  SDFFX1 DFF_726_Q_reg ( .D(WX4759), .SI(WX4758), .SE(n4533), .CLK(n4993), .Q(
        WX4760), .QN(n4120) );
  SDFFX1 DFF_727_Q_reg ( .D(WX4761), .SI(WX4760), .SE(n4532), .CLK(n4993), .Q(
        WX4762), .QN(n4121) );
  SDFFX1 DFF_728_Q_reg ( .D(WX4763), .SI(WX4762), .SE(n4531), .CLK(n4993), .Q(
        WX4764), .QN(n4122) );
  SDFFX1 DFF_729_Q_reg ( .D(WX4765), .SI(WX4764), .SE(n4531), .CLK(n4994), .Q(
        WX4766), .QN(n4123) );
  SDFFX1 DFF_730_Q_reg ( .D(WX4767), .SI(WX4766), .SE(n4530), .CLK(n4994), .Q(
        WX4768), .QN(n4124) );
  SDFFX1 DFF_731_Q_reg ( .D(WX4769), .SI(WX4768), .SE(n4529), .CLK(n4994), .Q(
        WX4770), .QN(n3953) );
  SDFFX1 DFF_732_Q_reg ( .D(WX4771), .SI(WX4770), .SE(n4529), .CLK(n4995), .Q(
        WX4772), .QN(n4125) );
  SDFFX1 DFF_733_Q_reg ( .D(WX4773), .SI(WX4772), .SE(n4528), .CLK(n4995), .Q(
        WX4774), .QN(n4126) );
  SDFFX1 DFF_734_Q_reg ( .D(WX4775), .SI(WX4774), .SE(n4527), .CLK(n4995), .Q(
        WX4776), .QN(n4127) );
  SDFFX1 DFF_735_Q_reg ( .D(WX4777), .SI(WX4776), .SE(n4527), .CLK(n4996), .Q(
        WX4778), .QN(n3965) );
  SDFFX1 DFF_736_Q_reg ( .D(WX5143), .SI(WX4778), .SE(n4366), .CLK(n5077), .Q(
        CRC_OUT_6_0), .QN(DFF_736_n1) );
  SDFFX1 DFF_737_Q_reg ( .D(WX5145), .SI(CRC_OUT_6_0), .SE(n4366), .CLK(n5077), 
        .Q(CRC_OUT_6_1), .QN(DFF_737_n1) );
  SDFFX1 DFF_738_Q_reg ( .D(WX5147), .SI(CRC_OUT_6_1), .SE(n4366), .CLK(n5077), 
        .Q(CRC_OUT_6_2), .QN(DFF_738_n1) );
  SDFFX1 DFF_739_Q_reg ( .D(WX5149), .SI(CRC_OUT_6_2), .SE(n4366), .CLK(n5077), 
        .Q(CRC_OUT_6_3), .QN(DFF_739_n1) );
  SDFFX1 DFF_740_Q_reg ( .D(WX5151), .SI(CRC_OUT_6_3), .SE(n4366), .CLK(n5077), 
        .Q(CRC_OUT_6_4), .QN(DFF_740_n1) );
  SDFFX1 DFF_741_Q_reg ( .D(WX5153), .SI(CRC_OUT_6_4), .SE(n4366), .CLK(n5077), 
        .Q(test_so42) );
  SDFFX1 DFF_742_Q_reg ( .D(WX5155), .SI(test_si43), .SE(n4365), .CLK(n5077), 
        .Q(CRC_OUT_6_6), .QN(DFF_742_n1) );
  SDFFX1 DFF_743_Q_reg ( .D(WX5157), .SI(CRC_OUT_6_6), .SE(n4365), .CLK(n5077), 
        .Q(CRC_OUT_6_7), .QN(DFF_743_n1) );
  SDFFX1 DFF_744_Q_reg ( .D(WX5159), .SI(CRC_OUT_6_7), .SE(n4365), .CLK(n5077), 
        .Q(CRC_OUT_6_8), .QN(DFF_744_n1) );
  SDFFX1 DFF_745_Q_reg ( .D(WX5161), .SI(CRC_OUT_6_8), .SE(n4365), .CLK(n5077), 
        .Q(CRC_OUT_6_9), .QN(DFF_745_n1) );
  SDFFX1 DFF_746_Q_reg ( .D(WX5163), .SI(CRC_OUT_6_9), .SE(n4365), .CLK(n5077), 
        .Q(CRC_OUT_6_10), .QN(DFF_746_n1) );
  SDFFX1 DFF_747_Q_reg ( .D(WX5165), .SI(CRC_OUT_6_10), .SE(n4365), .CLK(n5077), .Q(CRC_OUT_6_11), .QN(DFF_747_n1) );
  SDFFX1 DFF_748_Q_reg ( .D(WX5167), .SI(CRC_OUT_6_11), .SE(n4364), .CLK(n5078), .Q(CRC_OUT_6_12), .QN(DFF_748_n1) );
  SDFFX1 DFF_749_Q_reg ( .D(WX5169), .SI(CRC_OUT_6_12), .SE(n4364), .CLK(n5078), .Q(CRC_OUT_6_13), .QN(DFF_749_n1) );
  SDFFX1 DFF_750_Q_reg ( .D(WX5171), .SI(CRC_OUT_6_13), .SE(n4364), .CLK(n5078), .Q(CRC_OUT_6_14), .QN(DFF_750_n1) );
  SDFFX1 DFF_751_Q_reg ( .D(WX5173), .SI(CRC_OUT_6_14), .SE(n4364), .CLK(n5078), .Q(CRC_OUT_6_15), .QN(DFF_751_n1) );
  SDFFX1 DFF_752_Q_reg ( .D(WX5175), .SI(CRC_OUT_6_15), .SE(n4364), .CLK(n5078), .Q(CRC_OUT_6_16), .QN(DFF_752_n1) );
  SDFFX1 DFF_753_Q_reg ( .D(WX5177), .SI(CRC_OUT_6_16), .SE(n4364), .CLK(n5078), .Q(CRC_OUT_6_17), .QN(DFF_753_n1) );
  SDFFX1 DFF_754_Q_reg ( .D(WX5179), .SI(CRC_OUT_6_17), .SE(n4363), .CLK(n5078), .Q(CRC_OUT_6_18), .QN(DFF_754_n1) );
  SDFFX1 DFF_755_Q_reg ( .D(WX5181), .SI(CRC_OUT_6_18), .SE(n4363), .CLK(n5078), .Q(CRC_OUT_6_19), .QN(DFF_755_n1) );
  SDFFX1 DFF_756_Q_reg ( .D(WX5183), .SI(CRC_OUT_6_19), .SE(n4363), .CLK(n5078), .Q(CRC_OUT_6_20), .QN(DFF_756_n1) );
  SDFFX1 DFF_757_Q_reg ( .D(WX5185), .SI(CRC_OUT_6_20), .SE(n4363), .CLK(n5078), .Q(CRC_OUT_6_21), .QN(DFF_757_n1) );
  SDFFX1 DFF_758_Q_reg ( .D(WX5187), .SI(CRC_OUT_6_21), .SE(n4363), .CLK(n5078), .Q(test_so43) );
  SDFFX1 DFF_759_Q_reg ( .D(WX5189), .SI(test_si44), .SE(n4363), .CLK(n5078), 
        .Q(CRC_OUT_6_23), .QN(DFF_759_n1) );
  SDFFX1 DFF_760_Q_reg ( .D(WX5191), .SI(CRC_OUT_6_23), .SE(n4362), .CLK(n5079), .Q(CRC_OUT_6_24), .QN(DFF_760_n1) );
  SDFFX1 DFF_761_Q_reg ( .D(WX5193), .SI(CRC_OUT_6_24), .SE(n4362), .CLK(n5079), .Q(CRC_OUT_6_25), .QN(DFF_761_n1) );
  SDFFX1 DFF_762_Q_reg ( .D(WX5195), .SI(CRC_OUT_6_25), .SE(n4362), .CLK(n5079), .Q(CRC_OUT_6_26), .QN(DFF_762_n1) );
  SDFFX1 DFF_763_Q_reg ( .D(WX5197), .SI(CRC_OUT_6_26), .SE(n4362), .CLK(n5079), .Q(CRC_OUT_6_27), .QN(DFF_763_n1) );
  SDFFX1 DFF_764_Q_reg ( .D(WX5199), .SI(CRC_OUT_6_27), .SE(n4362), .CLK(n5079), .Q(CRC_OUT_6_28), .QN(DFF_764_n1) );
  SDFFX1 DFF_765_Q_reg ( .D(WX5201), .SI(CRC_OUT_6_28), .SE(n4362), .CLK(n5079), .Q(CRC_OUT_6_29), .QN(DFF_765_n1) );
  SDFFX1 DFF_766_Q_reg ( .D(WX5203), .SI(CRC_OUT_6_29), .SE(n4525), .CLK(n4996), .Q(CRC_OUT_6_30), .QN(DFF_766_n1) );
  SDFFX1 DFF_767_Q_reg ( .D(WX5205), .SI(CRC_OUT_6_30), .SE(n4525), .CLK(n4996), .Q(CRC_OUT_6_31), .QN(DFF_767_n1) );
  SDFFX1 DFF_768_Q_reg ( .D(n95), .SI(CRC_OUT_6_31), .SE(n4525), .CLK(n4997), 
        .Q(WX5657), .QN(n3935) );
  SDFFX1 DFF_769_Q_reg ( .D(n96), .SI(WX5657), .SE(n4520), .CLK(n4999), .Q(
        n8528) );
  SDFFX1 DFF_770_Q_reg ( .D(n97), .SI(n8528), .SE(n4520), .CLK(n4999), .Q(
        n8527) );
  SDFFX1 DFF_771_Q_reg ( .D(n98), .SI(n8527), .SE(n4520), .CLK(n4999), .Q(
        n8526) );
  SDFFX1 DFF_772_Q_reg ( .D(n99), .SI(n8526), .SE(n4520), .CLK(n4999), .Q(
        n8525) );
  SDFFX1 DFF_773_Q_reg ( .D(n100), .SI(n8525), .SE(n4521), .CLK(n4999), .Q(
        n8524) );
  SDFFX1 DFF_774_Q_reg ( .D(n101), .SI(n8524), .SE(n4521), .CLK(n4999), .Q(
        n8523) );
  SDFFX1 DFF_775_Q_reg ( .D(n102), .SI(n8523), .SE(n4521), .CLK(n4999), .Q(
        test_so44) );
  SDFFX1 DFF_776_Q_reg ( .D(n103), .SI(test_si45), .SE(n4521), .CLK(n4999), 
        .Q(n8520) );
  SDFFX1 DFF_777_Q_reg ( .D(n104), .SI(n8520), .SE(n4521), .CLK(n4998), .Q(
        n8519) );
  SDFFX1 DFF_778_Q_reg ( .D(n105), .SI(n8519), .SE(n4521), .CLK(n4998), .Q(
        n8518) );
  SDFFX1 DFF_779_Q_reg ( .D(n106), .SI(n8518), .SE(n4522), .CLK(n4998), .Q(
        n8517) );
  SDFFX1 DFF_780_Q_reg ( .D(n107), .SI(n8517), .SE(n4522), .CLK(n4998), .Q(
        n8516) );
  SDFFX1 DFF_781_Q_reg ( .D(n108), .SI(n8516), .SE(n4522), .CLK(n4998), .Q(
        n8515) );
  SDFFX1 DFF_782_Q_reg ( .D(n109), .SI(n8515), .SE(n4522), .CLK(n4998), .Q(
        n8514) );
  SDFFX1 DFF_783_Q_reg ( .D(n110), .SI(n8514), .SE(n4522), .CLK(n4998), .Q(
        n8513) );
  SDFFX1 DFF_784_Q_reg ( .D(n111), .SI(n8513), .SE(n4522), .CLK(n4998), .Q(
        n8512) );
  SDFFX1 DFF_785_Q_reg ( .D(n112), .SI(n8512), .SE(n4523), .CLK(n4998), .Q(
        n8511) );
  SDFFX1 DFF_786_Q_reg ( .D(n113), .SI(n8511), .SE(n4523), .CLK(n4998), .Q(
        n8510) );
  SDFFX1 DFF_787_Q_reg ( .D(n114), .SI(n8510), .SE(n4523), .CLK(n4998), .Q(
        n8509) );
  SDFFX1 DFF_788_Q_reg ( .D(n115), .SI(n8509), .SE(n4523), .CLK(n4998), .Q(
        n8508) );
  SDFFX1 DFF_789_Q_reg ( .D(n116), .SI(n8508), .SE(n4523), .CLK(n4997), .Q(
        n8507) );
  SDFFX1 DFF_790_Q_reg ( .D(n117), .SI(n8507), .SE(n4523), .CLK(n4997), .Q(
        n8506) );
  SDFFX1 DFF_791_Q_reg ( .D(n118), .SI(n8506), .SE(n4524), .CLK(n4997), .Q(
        n8505) );
  SDFFX1 DFF_792_Q_reg ( .D(n119), .SI(n8505), .SE(n4524), .CLK(n4997), .Q(
        test_so45) );
  SDFFX1 DFF_793_Q_reg ( .D(n120), .SI(test_si46), .SE(n4524), .CLK(n4997), 
        .Q(n8502) );
  SDFFX1 DFF_794_Q_reg ( .D(n121), .SI(n8502), .SE(n4524), .CLK(n4997), .Q(
        n8501) );
  SDFFX1 DFF_795_Q_reg ( .D(n122), .SI(n8501), .SE(n4524), .CLK(n4997), .Q(
        n8500) );
  SDFFX1 DFF_796_Q_reg ( .D(n123), .SI(n8500), .SE(n4524), .CLK(n4997), .Q(
        n8499) );
  SDFFX1 DFF_797_Q_reg ( .D(n124), .SI(n8499), .SE(n4525), .CLK(n4997), .Q(
        n8498) );
  SDFFX1 DFF_798_Q_reg ( .D(n125), .SI(n8498), .SE(n4525), .CLK(n4997), .Q(
        n8497) );
  SDFFX1 DFF_799_Q_reg ( .D(WX5718), .SI(n8497), .SE(n4525), .CLK(n4997), .Q(
        n8496) );
  SDFFX1 DFF_800_Q_reg ( .D(WX5816), .SI(n8496), .SE(n4520), .CLK(n4999), .Q(
        n8495), .QN(n8944) );
  SDFFX1 DFF_801_Q_reg ( .D(WX5818), .SI(n8495), .SE(n4519), .CLK(n4999), .Q(
        n8494), .QN(n8943) );
  SDFFX1 DFF_802_Q_reg ( .D(WX5820), .SI(n8494), .SE(n4519), .CLK(n5000), .Q(
        n8493), .QN(n8942) );
  SDFFX1 DFF_803_Q_reg ( .D(WX5822), .SI(n8493), .SE(n4519), .CLK(n5000), .Q(
        n8492), .QN(n8941) );
  SDFFX1 DFF_804_Q_reg ( .D(WX5824), .SI(n8492), .SE(n4518), .CLK(n5000), .Q(
        n8491), .QN(n8940) );
  SDFFX1 DFF_805_Q_reg ( .D(WX5826), .SI(n8491), .SE(n4518), .CLK(n5000), .Q(
        n8490), .QN(n8939) );
  SDFFX1 DFF_806_Q_reg ( .D(WX5828), .SI(n8490), .SE(n4518), .CLK(n5000), .Q(
        n8489), .QN(n8938) );
  SDFFX1 DFF_807_Q_reg ( .D(WX5830), .SI(n8489), .SE(n4517), .CLK(n5000), .Q(
        n8488), .QN(n8937) );
  SDFFX1 DFF_808_Q_reg ( .D(WX5832), .SI(n8488), .SE(n4517), .CLK(n5001), .Q(
        n8487), .QN(n8936) );
  SDFFX1 DFF_809_Q_reg ( .D(WX5834), .SI(n8487), .SE(n4367), .CLK(n5076), .Q(
        test_so46) );
  SDFFX1 DFF_810_Q_reg ( .D(WX5836), .SI(test_si47), .SE(n4516), .CLK(n5001), 
        .Q(n8484), .QN(n8935) );
  SDFFX1 DFF_811_Q_reg ( .D(WX5838), .SI(n8484), .SE(n4516), .CLK(n5001), .Q(
        n8483), .QN(n8932) );
  SDFFX1 DFF_812_Q_reg ( .D(WX5840), .SI(n8483), .SE(n4367), .CLK(n5076), .Q(
        n8482), .QN(n8931) );
  SDFFX1 DFF_813_Q_reg ( .D(WX5842), .SI(n8482), .SE(n4515), .CLK(n5001), .Q(
        n8481), .QN(n8928) );
  SDFFX1 DFF_814_Q_reg ( .D(WX5844), .SI(n8481), .SE(n4515), .CLK(n5002), .Q(
        n8480), .QN(n8927) );
  SDFFX1 DFF_815_Q_reg ( .D(WX5846), .SI(n8480), .SE(n4515), .CLK(n5002), .Q(
        n8479), .QN(n8926) );
  SDFFX1 DFF_816_Q_reg ( .D(WX5848), .SI(n8479), .SE(n4514), .CLK(n5002), .Q(
        WX5849) );
  SDFFX1 DFF_817_Q_reg ( .D(WX5850), .SI(WX5849), .SE(n4513), .CLK(n5002), .Q(
        WX5851) );
  SDFFX1 DFF_818_Q_reg ( .D(WX5852), .SI(WX5851), .SE(n4513), .CLK(n5003), .Q(
        WX5853) );
  SDFFX1 DFF_819_Q_reg ( .D(WX5854), .SI(WX5853), .SE(n4512), .CLK(n5003), .Q(
        WX5855) );
  SDFFX1 DFF_820_Q_reg ( .D(WX5856), .SI(WX5855), .SE(n4511), .CLK(n5003), .Q(
        WX5857) );
  SDFFX1 DFF_821_Q_reg ( .D(WX5858), .SI(WX5857), .SE(n4511), .CLK(n5004), .Q(
        WX5859) );
  SDFFX1 DFF_822_Q_reg ( .D(WX5860), .SI(WX5859), .SE(n4510), .CLK(n5004), .Q(
        WX5861) );
  SDFFX1 DFF_823_Q_reg ( .D(WX5862), .SI(WX5861), .SE(n4509), .CLK(n5004), .Q(
        WX5863) );
  SDFFX1 DFF_824_Q_reg ( .D(WX5864), .SI(WX5863), .SE(n4509), .CLK(n5005), .Q(
        WX5865) );
  SDFFX1 DFF_825_Q_reg ( .D(WX5866), .SI(WX5865), .SE(n4508), .CLK(n5005), .Q(
        WX5867) );
  SDFFX1 DFF_826_Q_reg ( .D(WX5868), .SI(WX5867), .SE(n4507), .CLK(n5005), .Q(
        test_so47) );
  SDFFX1 DFF_827_Q_reg ( .D(WX5870), .SI(test_si48), .SE(n4506), .CLK(n5006), 
        .Q(WX5871) );
  SDFFX1 DFF_828_Q_reg ( .D(WX5872), .SI(WX5871), .SE(n4506), .CLK(n5006), .Q(
        WX5873) );
  SDFFX1 DFF_829_Q_reg ( .D(WX5874), .SI(WX5873), .SE(n4505), .CLK(n5006), .Q(
        WX5875) );
  SDFFX1 DFF_830_Q_reg ( .D(WX5876), .SI(WX5875), .SE(n4505), .CLK(n5007), .Q(
        WX5877) );
  SDFFX1 DFF_831_Q_reg ( .D(WX5878), .SI(WX5877), .SE(n4504), .CLK(n5007), .Q(
        WX5879) );
  SDFFX1 DFF_832_Q_reg ( .D(WX5880), .SI(WX5879), .SE(n4520), .CLK(n4999), .Q(
        WX5881), .QN(n3586) );
  SDFFX1 DFF_833_Q_reg ( .D(WX5882), .SI(WX5881), .SE(n4519), .CLK(n4999), .Q(
        WX5883), .QN(n3654) );
  SDFFX1 DFF_834_Q_reg ( .D(WX5884), .SI(WX5883), .SE(n4519), .CLK(n5000), .Q(
        WX5885), .QN(n3653) );
  SDFFX1 DFF_835_Q_reg ( .D(WX5886), .SI(WX5885), .SE(n4519), .CLK(n5000), .Q(
        WX5887), .QN(n3652) );
  SDFFX1 DFF_836_Q_reg ( .D(WX5888), .SI(WX5887), .SE(n4518), .CLK(n5000), .Q(
        WX5889), .QN(n3651) );
  SDFFX1 DFF_837_Q_reg ( .D(WX5890), .SI(WX5889), .SE(n4518), .CLK(n5000), .Q(
        WX5891), .QN(n3650) );
  SDFFX1 DFF_838_Q_reg ( .D(WX5892), .SI(WX5891), .SE(n4518), .CLK(n5000), .Q(
        WX5893), .QN(n3649) );
  SDFFX1 DFF_839_Q_reg ( .D(WX5894), .SI(WX5893), .SE(n4517), .CLK(n5000), .Q(
        WX5895), .QN(n3648) );
  SDFFX1 DFF_840_Q_reg ( .D(WX5896), .SI(WX5895), .SE(n4517), .CLK(n5001), .Q(
        WX5897), .QN(n3647) );
  SDFFX1 DFF_841_Q_reg ( .D(WX5898), .SI(WX5897), .SE(n4517), .CLK(n5001), .Q(
        WX5899) );
  SDFFX1 DFF_842_Q_reg ( .D(WX5900), .SI(WX5899), .SE(n4517), .CLK(n5001), .Q(
        WX5901), .QN(n3645) );
  SDFFX1 DFF_843_Q_reg ( .D(WX5902), .SI(WX5901), .SE(n4516), .CLK(n5001), .Q(
        test_so48), .QN(n8933) );
  SDFFX1 DFF_844_Q_reg ( .D(WX5904), .SI(test_si49), .SE(n4367), .CLK(n5076), 
        .Q(WX5905), .QN(n3644) );
  SDFFX1 DFF_845_Q_reg ( .D(WX5906), .SI(WX5905), .SE(n4515), .CLK(n5001), .Q(
        WX5907), .QN(n8930) );
  SDFFX1 DFF_846_Q_reg ( .D(WX5908), .SI(WX5907), .SE(n4515), .CLK(n5002), .Q(
        WX5909), .QN(n3643) );
  SDFFX1 DFF_847_Q_reg ( .D(WX5910), .SI(WX5909), .SE(n4514), .CLK(n5002), .Q(
        WX5911) );
  SDFFX1 DFF_848_Q_reg ( .D(WX5912), .SI(WX5911), .SE(n4514), .CLK(n5002), .Q(
        WX5913), .QN(n8925) );
  SDFFX1 DFF_849_Q_reg ( .D(WX5914), .SI(WX5913), .SE(n4513), .CLK(n5002), .Q(
        WX5915), .QN(n8924) );
  SDFFX1 DFF_850_Q_reg ( .D(WX5916), .SI(WX5915), .SE(n4513), .CLK(n5003), .Q(
        WX5917), .QN(n8923) );
  SDFFX1 DFF_851_Q_reg ( .D(WX5918), .SI(WX5917), .SE(n4512), .CLK(n5003), .Q(
        WX5919), .QN(n8922) );
  SDFFX1 DFF_852_Q_reg ( .D(WX5920), .SI(WX5919), .SE(n4511), .CLK(n5003), .Q(
        WX5921), .QN(n8921) );
  SDFFX1 DFF_853_Q_reg ( .D(WX5922), .SI(WX5921), .SE(n4511), .CLK(n5004), .Q(
        WX5923), .QN(n8920) );
  SDFFX1 DFF_854_Q_reg ( .D(WX5924), .SI(WX5923), .SE(n4510), .CLK(n5004), .Q(
        WX5925), .QN(n8919) );
  SDFFX1 DFF_855_Q_reg ( .D(WX5926), .SI(WX5925), .SE(n4509), .CLK(n5004), .Q(
        WX5927), .QN(n8918) );
  SDFFX1 DFF_856_Q_reg ( .D(WX5928), .SI(WX5927), .SE(n4509), .CLK(n5005), .Q(
        WX5929), .QN(n8917) );
  SDFFX1 DFF_857_Q_reg ( .D(WX5930), .SI(WX5929), .SE(n4508), .CLK(n5005), .Q(
        WX5931), .QN(n8916) );
  SDFFX1 DFF_858_Q_reg ( .D(WX5932), .SI(WX5931), .SE(n4507), .CLK(n5005), .Q(
        WX5933), .QN(n8915) );
  SDFFX1 DFF_859_Q_reg ( .D(WX5934), .SI(WX5933), .SE(n4507), .CLK(n5006), .Q(
        WX5935), .QN(n8914) );
  SDFFX1 DFF_860_Q_reg ( .D(WX5936), .SI(WX5935), .SE(n4506), .CLK(n5006), .Q(
        test_so49) );
  SDFFX1 DFF_861_Q_reg ( .D(WX5938), .SI(test_si50), .SE(n4505), .CLK(n5006), 
        .Q(WX5939), .QN(n8912) );
  SDFFX1 DFF_862_Q_reg ( .D(WX5940), .SI(WX5939), .SE(n4505), .CLK(n5007), .Q(
        WX5941), .QN(n8911) );
  SDFFX1 DFF_863_Q_reg ( .D(WX5942), .SI(WX5941), .SE(n4504), .CLK(n5007), .Q(
        WX5943), .QN(n8910) );
  SDFFX1 DFF_864_Q_reg ( .D(WX5944), .SI(WX5943), .SE(n4503), .CLK(n5007), .Q(
        WX5945) );
  SDFFX1 DFF_865_Q_reg ( .D(WX5946), .SI(WX5945), .SE(n4503), .CLK(n5008), .Q(
        WX5947) );
  SDFFX1 DFF_866_Q_reg ( .D(WX5948), .SI(WX5947), .SE(n4503), .CLK(n5008), .Q(
        WX5949) );
  SDFFX1 DFF_867_Q_reg ( .D(WX5950), .SI(WX5949), .SE(n4502), .CLK(n5008), .Q(
        WX5951) );
  SDFFX1 DFF_868_Q_reg ( .D(WX5952), .SI(WX5951), .SE(n4502), .CLK(n5008), .Q(
        WX5953) );
  SDFFX1 DFF_869_Q_reg ( .D(WX5954), .SI(WX5953), .SE(n4502), .CLK(n5008), .Q(
        WX5955) );
  SDFFX1 DFF_870_Q_reg ( .D(WX5956), .SI(WX5955), .SE(n4501), .CLK(n5008), .Q(
        WX5957) );
  SDFFX1 DFF_871_Q_reg ( .D(WX5958), .SI(WX5957), .SE(n4501), .CLK(n5009), .Q(
        WX5959) );
  SDFFX1 DFF_872_Q_reg ( .D(WX5960), .SI(WX5959), .SE(n4501), .CLK(n5009), .Q(
        WX5961) );
  SDFFX1 DFF_873_Q_reg ( .D(WX5962), .SI(WX5961), .SE(n4500), .CLK(n5009), .Q(
        WX5963), .QN(n3646) );
  SDFFX1 DFF_874_Q_reg ( .D(WX5964), .SI(WX5963), .SE(n4500), .CLK(n5009), .Q(
        WX5965) );
  SDFFX1 DFF_875_Q_reg ( .D(WX5966), .SI(WX5965), .SE(n4516), .CLK(n5001), .Q(
        WX5967), .QN(n8934) );
  SDFFX1 DFF_876_Q_reg ( .D(WX5968), .SI(WX5967), .SE(n4516), .CLK(n5001), .Q(
        WX5969) );
  SDFFX1 DFF_877_Q_reg ( .D(WX5970), .SI(WX5969), .SE(n4516), .CLK(n5001), .Q(
        test_so50), .QN(n8929) );
  SDFFX1 DFF_878_Q_reg ( .D(WX5972), .SI(test_si51), .SE(n4515), .CLK(n5002), 
        .Q(WX5973) );
  SDFFX1 DFF_879_Q_reg ( .D(WX5974), .SI(WX5973), .SE(n4514), .CLK(n5002), .Q(
        WX5975), .QN(n3642) );
  SDFFX1 DFF_880_Q_reg ( .D(WX5976), .SI(WX5975), .SE(n4514), .CLK(n5002), .Q(
        WX5977), .QN(n3841) );
  SDFFX1 DFF_881_Q_reg ( .D(WX5978), .SI(WX5977), .SE(n4513), .CLK(n5003), .Q(
        WX5979), .QN(n3839) );
  SDFFX1 DFF_882_Q_reg ( .D(WX5980), .SI(WX5979), .SE(n4512), .CLK(n5003), .Q(
        WX5981), .QN(n3837) );
  SDFFX1 DFF_883_Q_reg ( .D(WX5982), .SI(WX5981), .SE(n4512), .CLK(n5003), .Q(
        WX5983), .QN(n3835) );
  SDFFX1 DFF_884_Q_reg ( .D(WX5984), .SI(WX5983), .SE(n4511), .CLK(n5004), .Q(
        WX5985), .QN(n3833) );
  SDFFX1 DFF_885_Q_reg ( .D(WX5986), .SI(WX5985), .SE(n4510), .CLK(n5004), .Q(
        WX5987), .QN(n3831) );
  SDFFX1 DFF_886_Q_reg ( .D(WX5988), .SI(WX5987), .SE(n4510), .CLK(n5004), .Q(
        WX5989), .QN(n3829) );
  SDFFX1 DFF_887_Q_reg ( .D(WX5990), .SI(WX5989), .SE(n4509), .CLK(n5005), .Q(
        WX5991), .QN(n3827) );
  SDFFX1 DFF_888_Q_reg ( .D(WX5992), .SI(WX5991), .SE(n4508), .CLK(n5005), .Q(
        WX5993), .QN(n3825) );
  SDFFX1 DFF_889_Q_reg ( .D(WX5994), .SI(WX5993), .SE(n4508), .CLK(n5005), .Q(
        WX5995), .QN(n3823) );
  SDFFX1 DFF_890_Q_reg ( .D(WX5996), .SI(WX5995), .SE(n4507), .CLK(n5006), .Q(
        WX5997) );
  SDFFX1 DFF_891_Q_reg ( .D(WX5998), .SI(WX5997), .SE(n4507), .CLK(n5006), .Q(
        WX5999), .QN(n3820) );
  SDFFX1 DFF_892_Q_reg ( .D(WX6000), .SI(WX5999), .SE(n4506), .CLK(n5006), .Q(
        WX6001), .QN(n8913) );
  SDFFX1 DFF_893_Q_reg ( .D(WX6002), .SI(WX6001), .SE(n4505), .CLK(n5007), .Q(
        WX6003), .QN(n3817) );
  SDFFX1 DFF_894_Q_reg ( .D(WX6004), .SI(WX6003), .SE(n4504), .CLK(n5007), .Q(
        test_so51) );
  SDFFX1 DFF_895_Q_reg ( .D(WX6006), .SI(test_si52), .SE(n4504), .CLK(n5007), 
        .Q(WX6007), .QN(n3814) );
  SDFFX1 DFF_896_Q_reg ( .D(WX6008), .SI(WX6007), .SE(n4503), .CLK(n5007), .Q(
        WX6009), .QN(n4073) );
  SDFFX1 DFF_897_Q_reg ( .D(WX6010), .SI(WX6009), .SE(n4503), .CLK(n5008), .Q(
        WX6011), .QN(n4074) );
  SDFFX1 DFF_898_Q_reg ( .D(WX6012), .SI(WX6011), .SE(n4503), .CLK(n5008), .Q(
        WX6013), .QN(n4075) );
  SDFFX1 DFF_899_Q_reg ( .D(WX6014), .SI(WX6013), .SE(n4502), .CLK(n5008), .Q(
        WX6015), .QN(n4076) );
  SDFFX1 DFF_900_Q_reg ( .D(WX6016), .SI(WX6015), .SE(n4502), .CLK(n5008), .Q(
        WX6017), .QN(n4077) );
  SDFFX1 DFF_901_Q_reg ( .D(WX6018), .SI(WX6017), .SE(n4502), .CLK(n5008), .Q(
        WX6019), .QN(n4078) );
  SDFFX1 DFF_902_Q_reg ( .D(WX6020), .SI(WX6019), .SE(n4501), .CLK(n5008), .Q(
        WX6021), .QN(n4079) );
  SDFFX1 DFF_903_Q_reg ( .D(WX6022), .SI(WX6021), .SE(n4501), .CLK(n5009), .Q(
        WX6023), .QN(n4080) );
  SDFFX1 DFF_904_Q_reg ( .D(WX6024), .SI(WX6023), .SE(n4501), .CLK(n5009), .Q(
        WX6025), .QN(n4081) );
  SDFFX1 DFF_905_Q_reg ( .D(WX6026), .SI(WX6025), .SE(n4500), .CLK(n5009), .Q(
        WX6027), .QN(n4082) );
  SDFFX1 DFF_906_Q_reg ( .D(WX6028), .SI(WX6027), .SE(n4500), .CLK(n5009), .Q(
        WX6029), .QN(n4083) );
  SDFFX1 DFF_907_Q_reg ( .D(WX6030), .SI(WX6029), .SE(n4500), .CLK(n5009), .Q(
        WX6031), .QN(n4084) );
  SDFFX1 DFF_908_Q_reg ( .D(WX6032), .SI(WX6031), .SE(n4500), .CLK(n5009), .Q(
        WX6033), .QN(n4085) );
  SDFFX1 DFF_909_Q_reg ( .D(WX6034), .SI(WX6033), .SE(n4499), .CLK(n5009), .Q(
        WX6035), .QN(n4086) );
  SDFFX1 DFF_910_Q_reg ( .D(WX6036), .SI(WX6035), .SE(n4499), .CLK(n5009), .Q(
        WX6037), .QN(n4087) );
  SDFFX1 DFF_911_Q_reg ( .D(WX6038), .SI(WX6037), .SE(n4499), .CLK(n5010), .Q(
        test_so52) );
  SDFFX1 DFF_912_Q_reg ( .D(WX6040), .SI(test_si53), .SE(n4514), .CLK(n5002), 
        .Q(WX6041), .QN(n4088) );
  SDFFX1 DFF_913_Q_reg ( .D(WX6042), .SI(WX6041), .SE(n4513), .CLK(n5003), .Q(
        WX6043), .QN(n4089) );
  SDFFX1 DFF_914_Q_reg ( .D(WX6044), .SI(WX6043), .SE(n4512), .CLK(n5003), .Q(
        WX6045), .QN(n4090) );
  SDFFX1 DFF_915_Q_reg ( .D(WX6046), .SI(WX6045), .SE(n4512), .CLK(n5003), .Q(
        WX6047), .QN(n4091) );
  SDFFX1 DFF_916_Q_reg ( .D(WX6048), .SI(WX6047), .SE(n4511), .CLK(n5004), .Q(
        WX6049), .QN(n3950) );
  SDFFX1 DFF_917_Q_reg ( .D(WX6050), .SI(WX6049), .SE(n4510), .CLK(n5004), .Q(
        WX6051), .QN(n4092) );
  SDFFX1 DFF_918_Q_reg ( .D(WX6052), .SI(WX6051), .SE(n4510), .CLK(n5004), .Q(
        WX6053), .QN(n4093) );
  SDFFX1 DFF_919_Q_reg ( .D(WX6054), .SI(WX6053), .SE(n4509), .CLK(n5005), .Q(
        WX6055), .QN(n4094) );
  SDFFX1 DFF_920_Q_reg ( .D(WX6056), .SI(WX6055), .SE(n4508), .CLK(n5005), .Q(
        WX6057), .QN(n4095) );
  SDFFX1 DFF_921_Q_reg ( .D(WX6058), .SI(WX6057), .SE(n4508), .CLK(n5005), .Q(
        WX6059), .QN(n4096) );
  SDFFX1 DFF_922_Q_reg ( .D(WX6060), .SI(WX6059), .SE(n4507), .CLK(n5006), .Q(
        WX6061), .QN(n4097) );
  SDFFX1 DFF_923_Q_reg ( .D(WX6062), .SI(WX6061), .SE(n4506), .CLK(n5006), .Q(
        WX6063), .QN(n3951) );
  SDFFX1 DFF_924_Q_reg ( .D(WX6064), .SI(WX6063), .SE(n4506), .CLK(n5006), .Q(
        WX6065), .QN(n4098) );
  SDFFX1 DFF_925_Q_reg ( .D(WX6066), .SI(WX6065), .SE(n4505), .CLK(n5007), .Q(
        WX6067), .QN(n4099) );
  SDFFX1 DFF_926_Q_reg ( .D(WX6068), .SI(WX6067), .SE(n4504), .CLK(n5007), .Q(
        WX6069), .QN(n4100) );
  SDFFX1 DFF_927_Q_reg ( .D(WX6070), .SI(WX6069), .SE(n4504), .CLK(n5007), .Q(
        WX6071), .QN(n3964) );
  SDFFX1 DFF_928_Q_reg ( .D(WX6436), .SI(WX6071), .SE(n4492), .CLK(n5013), .Q(
        test_so53) );
  SDFFX1 DFF_929_Q_reg ( .D(WX6438), .SI(test_si54), .SE(n4492), .CLK(n5013), 
        .Q(CRC_OUT_5_1), .QN(DFF_929_n1) );
  SDFFX1 DFF_930_Q_reg ( .D(WX6440), .SI(CRC_OUT_5_1), .SE(n4491), .CLK(n5013), 
        .Q(CRC_OUT_5_2), .QN(DFF_930_n1) );
  SDFFX1 DFF_931_Q_reg ( .D(WX6442), .SI(CRC_OUT_5_2), .SE(n4491), .CLK(n5013), 
        .Q(CRC_OUT_5_3), .QN(DFF_931_n1) );
  SDFFX1 DFF_932_Q_reg ( .D(WX6444), .SI(CRC_OUT_5_3), .SE(n4491), .CLK(n5014), 
        .Q(CRC_OUT_5_4), .QN(DFF_932_n1) );
  SDFFX1 DFF_933_Q_reg ( .D(WX6446), .SI(CRC_OUT_5_4), .SE(n4491), .CLK(n5014), 
        .Q(CRC_OUT_5_5), .QN(DFF_933_n1) );
  SDFFX1 DFF_934_Q_reg ( .D(WX6448), .SI(CRC_OUT_5_5), .SE(n4491), .CLK(n5014), 
        .Q(CRC_OUT_5_6), .QN(DFF_934_n1) );
  SDFFX1 DFF_935_Q_reg ( .D(WX6450), .SI(CRC_OUT_5_6), .SE(n4491), .CLK(n5014), 
        .Q(CRC_OUT_5_7), .QN(DFF_935_n1) );
  SDFFX1 DFF_936_Q_reg ( .D(WX6452), .SI(CRC_OUT_5_7), .SE(n4490), .CLK(n5014), 
        .Q(CRC_OUT_5_8), .QN(DFF_936_n1) );
  SDFFX1 DFF_937_Q_reg ( .D(WX6454), .SI(CRC_OUT_5_8), .SE(n4490), .CLK(n5014), 
        .Q(CRC_OUT_5_9), .QN(DFF_937_n1) );
  SDFFX1 DFF_938_Q_reg ( .D(WX6456), .SI(CRC_OUT_5_9), .SE(n4490), .CLK(n5014), 
        .Q(CRC_OUT_5_10), .QN(DFF_938_n1) );
  SDFFX1 DFF_939_Q_reg ( .D(WX6458), .SI(CRC_OUT_5_10), .SE(n4490), .CLK(n5014), .Q(CRC_OUT_5_11), .QN(DFF_939_n1) );
  SDFFX1 DFF_940_Q_reg ( .D(WX6460), .SI(CRC_OUT_5_11), .SE(n4490), .CLK(n5014), .Q(CRC_OUT_5_12), .QN(DFF_940_n1) );
  SDFFX1 DFF_941_Q_reg ( .D(WX6462), .SI(CRC_OUT_5_12), .SE(n4490), .CLK(n5014), .Q(CRC_OUT_5_13), .QN(DFF_941_n1) );
  SDFFX1 DFF_942_Q_reg ( .D(WX6464), .SI(CRC_OUT_5_13), .SE(n4489), .CLK(n5014), .Q(CRC_OUT_5_14), .QN(DFF_942_n1) );
  SDFFX1 DFF_943_Q_reg ( .D(WX6466), .SI(CRC_OUT_5_14), .SE(n4489), .CLK(n5014), .Q(CRC_OUT_5_15), .QN(DFF_943_n1) );
  SDFFX1 DFF_944_Q_reg ( .D(WX6468), .SI(CRC_OUT_5_15), .SE(n4489), .CLK(n5015), .Q(CRC_OUT_5_16), .QN(DFF_944_n1) );
  SDFFX1 DFF_945_Q_reg ( .D(WX6470), .SI(CRC_OUT_5_16), .SE(n4489), .CLK(n5015), .Q(test_so54) );
  SDFFX1 DFF_946_Q_reg ( .D(WX6472), .SI(test_si55), .SE(n4489), .CLK(n5015), 
        .Q(CRC_OUT_5_18), .QN(DFF_946_n1) );
  SDFFX1 DFF_947_Q_reg ( .D(WX6474), .SI(CRC_OUT_5_18), .SE(n4489), .CLK(n5015), .Q(CRC_OUT_5_19), .QN(DFF_947_n1) );
  SDFFX1 DFF_948_Q_reg ( .D(WX6476), .SI(CRC_OUT_5_19), .SE(n4367), .CLK(n5076), .Q(CRC_OUT_5_20), .QN(DFF_948_n1) );
  SDFFX1 DFF_949_Q_reg ( .D(WX6478), .SI(CRC_OUT_5_20), .SE(n4499), .CLK(n5010), .Q(CRC_OUT_5_21), .QN(DFF_949_n1) );
  SDFFX1 DFF_950_Q_reg ( .D(WX6480), .SI(CRC_OUT_5_21), .SE(n4499), .CLK(n5010), .Q(CRC_OUT_5_22), .QN(DFF_950_n1) );
  SDFFX1 DFF_951_Q_reg ( .D(WX6482), .SI(CRC_OUT_5_22), .SE(n4499), .CLK(n5010), .Q(CRC_OUT_5_23), .QN(DFF_951_n1) );
  SDFFX1 DFF_952_Q_reg ( .D(WX6484), .SI(CRC_OUT_5_23), .SE(n4498), .CLK(n5010), .Q(CRC_OUT_5_24), .QN(DFF_952_n1) );
  SDFFX1 DFF_953_Q_reg ( .D(WX6486), .SI(CRC_OUT_5_24), .SE(n4498), .CLK(n5010), .Q(CRC_OUT_5_25), .QN(DFF_953_n1) );
  SDFFX1 DFF_954_Q_reg ( .D(WX6488), .SI(CRC_OUT_5_25), .SE(n4498), .CLK(n5010), .Q(CRC_OUT_5_26), .QN(DFF_954_n1) );
  SDFFX1 DFF_955_Q_reg ( .D(WX6490), .SI(CRC_OUT_5_26), .SE(n4498), .CLK(n5010), .Q(CRC_OUT_5_27), .QN(DFF_955_n1) );
  SDFFX1 DFF_956_Q_reg ( .D(WX6492), .SI(CRC_OUT_5_27), .SE(n4498), .CLK(n5010), .Q(CRC_OUT_5_28), .QN(DFF_956_n1) );
  SDFFX1 DFF_957_Q_reg ( .D(WX6494), .SI(CRC_OUT_5_28), .SE(n4498), .CLK(n5010), .Q(CRC_OUT_5_29), .QN(DFF_957_n1) );
  SDFFX1 DFF_958_Q_reg ( .D(WX6496), .SI(CRC_OUT_5_29), .SE(n4497), .CLK(n5010), .Q(CRC_OUT_5_30), .QN(DFF_958_n1) );
  SDFFX1 DFF_959_Q_reg ( .D(WX6498), .SI(CRC_OUT_5_30), .SE(n4497), .CLK(n5010), .Q(CRC_OUT_5_31), .QN(DFF_959_n1) );
  SDFFX1 DFF_960_Q_reg ( .D(n126), .SI(CRC_OUT_5_31), .SE(n4497), .CLK(n5011), 
        .Q(WX6950), .QN(n3934) );
  SDFFX1 DFF_961_Q_reg ( .D(n127), .SI(WX6950), .SE(n4492), .CLK(n5013), .Q(
        n8470) );
  SDFFX1 DFF_962_Q_reg ( .D(n128), .SI(n8470), .SE(n4492), .CLK(n5013), .Q(
        test_so55) );
  SDFFX1 DFF_963_Q_reg ( .D(n129), .SI(test_si56), .SE(n4492), .CLK(n5013), 
        .Q(n8467) );
  SDFFX1 DFF_964_Q_reg ( .D(n130), .SI(n8467), .SE(n4492), .CLK(n5013), .Q(
        n8466) );
  SDFFX1 DFF_965_Q_reg ( .D(n131), .SI(n8466), .SE(n4493), .CLK(n5013), .Q(
        n8465) );
  SDFFX1 DFF_966_Q_reg ( .D(n132), .SI(n8465), .SE(n4493), .CLK(n5013), .Q(
        n8464) );
  SDFFX1 DFF_967_Q_reg ( .D(n133), .SI(n8464), .SE(n4493), .CLK(n5013), .Q(
        n8463) );
  SDFFX1 DFF_968_Q_reg ( .D(n134), .SI(n8463), .SE(n4493), .CLK(n5013), .Q(
        n8462) );
  SDFFX1 DFF_969_Q_reg ( .D(n135), .SI(n8462), .SE(n4493), .CLK(n5012), .Q(
        n8461) );
  SDFFX1 DFF_970_Q_reg ( .D(n136), .SI(n8461), .SE(n4493), .CLK(n5012), .Q(
        n8460) );
  SDFFX1 DFF_971_Q_reg ( .D(n137), .SI(n8460), .SE(n4494), .CLK(n5012), .Q(
        n8459) );
  SDFFX1 DFF_972_Q_reg ( .D(n138), .SI(n8459), .SE(n4494), .CLK(n5012), .Q(
        n8458) );
  SDFFX1 DFF_973_Q_reg ( .D(n139), .SI(n8458), .SE(n4494), .CLK(n5012), .Q(
        n8457) );
  SDFFX1 DFF_974_Q_reg ( .D(n140), .SI(n8457), .SE(n4494), .CLK(n5012), .Q(
        n8456) );
  SDFFX1 DFF_975_Q_reg ( .D(n141), .SI(n8456), .SE(n4494), .CLK(n5012), .Q(
        n8455) );
  SDFFX1 DFF_976_Q_reg ( .D(n142), .SI(n8455), .SE(n4494), .CLK(n5012), .Q(
        n8454) );
  SDFFX1 DFF_977_Q_reg ( .D(n143), .SI(n8454), .SE(n4495), .CLK(n5012), .Q(
        n8453) );
  SDFFX1 DFF_978_Q_reg ( .D(n144), .SI(n8453), .SE(n4495), .CLK(n5012), .Q(
        n8452) );
  SDFFX1 DFF_979_Q_reg ( .D(n145), .SI(n8452), .SE(n4495), .CLK(n5012), .Q(
        test_so56) );
  SDFFX1 DFF_980_Q_reg ( .D(n146), .SI(test_si57), .SE(n4495), .CLK(n5012), 
        .Q(n8449) );
  SDFFX1 DFF_981_Q_reg ( .D(n147), .SI(n8449), .SE(n4495), .CLK(n5011), .Q(
        n8448) );
  SDFFX1 DFF_982_Q_reg ( .D(n148), .SI(n8448), .SE(n4495), .CLK(n5011), .Q(
        n8447) );
  SDFFX1 DFF_983_Q_reg ( .D(n149), .SI(n8447), .SE(n4496), .CLK(n5011), .Q(
        n8446) );
  SDFFX1 DFF_984_Q_reg ( .D(n150), .SI(n8446), .SE(n4496), .CLK(n5011), .Q(
        n8445) );
  SDFFX1 DFF_985_Q_reg ( .D(n151), .SI(n8445), .SE(n4496), .CLK(n5011), .Q(
        n8444) );
  SDFFX1 DFF_986_Q_reg ( .D(n152), .SI(n8444), .SE(n4496), .CLK(n5011), .Q(
        n8443) );
  SDFFX1 DFF_987_Q_reg ( .D(n153), .SI(n8443), .SE(n4496), .CLK(n5011), .Q(
        n8442) );
  SDFFX1 DFF_988_Q_reg ( .D(n154), .SI(n8442), .SE(n4496), .CLK(n5011), .Q(
        n8441) );
  SDFFX1 DFF_989_Q_reg ( .D(n155), .SI(n8441), .SE(n4497), .CLK(n5011), .Q(
        n8440) );
  SDFFX1 DFF_990_Q_reg ( .D(n156), .SI(n8440), .SE(n4497), .CLK(n5011), .Q(
        n8439) );
  SDFFX1 DFF_991_Q_reg ( .D(WX7011), .SI(n8439), .SE(n4497), .CLK(n5011), .Q(
        n8438) );
  SDFFX1 DFF_992_Q_reg ( .D(WX7109), .SI(n8438), .SE(n4367), .CLK(n5076), .Q(
        n8437), .QN(n8909) );
  SDFFX1 DFF_993_Q_reg ( .D(WX7111), .SI(n8437), .SE(n4486), .CLK(n5016), .Q(
        n8436), .QN(n8908) );
  SDFFX1 DFF_994_Q_reg ( .D(WX7113), .SI(n8436), .SE(n4485), .CLK(n5017), .Q(
        n8435), .QN(n8907) );
  SDFFX1 DFF_995_Q_reg ( .D(WX7115), .SI(n8435), .SE(n4485), .CLK(n5017), .Q(
        n8434), .QN(n8906) );
  SDFFX1 DFF_996_Q_reg ( .D(WX7117), .SI(n8434), .SE(n4367), .CLK(n5076), .Q(
        test_so57) );
  SDFFX1 DFF_997_Q_reg ( .D(WX7119), .SI(test_si58), .SE(n4484), .CLK(n5017), 
        .Q(n8431), .QN(n8905) );
  SDFFX1 DFF_998_Q_reg ( .D(WX7121), .SI(n8431), .SE(n4484), .CLK(n5017), .Q(
        n8430), .QN(n8902) );
  SDFFX1 DFF_999_Q_reg ( .D(WX7123), .SI(n8430), .SE(n4368), .CLK(n5076), .Q(
        n8429), .QN(n8901) );
  SDFFX1 DFF_1000_Q_reg ( .D(WX7125), .SI(n8429), .SE(n4483), .CLK(n5018), .Q(
        n8428), .QN(n8898) );
  SDFFX1 DFF_1001_Q_reg ( .D(WX7127), .SI(n8428), .SE(n4483), .CLK(n5018), .Q(
        n8427), .QN(n8897) );
  SDFFX1 DFF_1002_Q_reg ( .D(WX7129), .SI(n8427), .SE(n4482), .CLK(n5018), .Q(
        n8426), .QN(n8896) );
  SDFFX1 DFF_1003_Q_reg ( .D(WX7131), .SI(n8426), .SE(n4481), .CLK(n5018), .Q(
        n8425), .QN(n8895) );
  SDFFX1 DFF_1004_Q_reg ( .D(WX7133), .SI(n8425), .SE(n4481), .CLK(n5019), .Q(
        n8424), .QN(n8894) );
  SDFFX1 DFF_1005_Q_reg ( .D(WX7135), .SI(n8424), .SE(n4480), .CLK(n5019), .Q(
        n8423), .QN(n8893) );
  SDFFX1 DFF_1006_Q_reg ( .D(WX7137), .SI(n8423), .SE(n4480), .CLK(n5019), .Q(
        n8422), .QN(n8892) );
  SDFFX1 DFF_1007_Q_reg ( .D(WX7139), .SI(n8422), .SE(n4479), .CLK(n5020), .Q(
        n8421), .QN(n8891) );
  SDFFX1 DFF_1008_Q_reg ( .D(WX7141), .SI(n8421), .SE(n4479), .CLK(n5020), .Q(
        WX7142) );
  SDFFX1 DFF_1009_Q_reg ( .D(WX7143), .SI(WX7142), .SE(n4478), .CLK(n5020), 
        .Q(WX7144) );
  SDFFX1 DFF_1010_Q_reg ( .D(WX7145), .SI(WX7144), .SE(n4477), .CLK(n5021), 
        .Q(WX7146) );
  SDFFX1 DFF_1011_Q_reg ( .D(WX7147), .SI(WX7146), .SE(n4477), .CLK(n5021), 
        .Q(WX7148) );
  SDFFX1 DFF_1012_Q_reg ( .D(WX7149), .SI(WX7148), .SE(n4476), .CLK(n5021), 
        .Q(WX7150) );
  SDFFX1 DFF_1013_Q_reg ( .D(WX7151), .SI(WX7150), .SE(n4475), .CLK(n5022), 
        .Q(test_so58) );
  SDFFX1 DFF_1014_Q_reg ( .D(WX7153), .SI(test_si59), .SE(n4474), .CLK(n5022), 
        .Q(WX7154) );
  SDFFX1 DFF_1015_Q_reg ( .D(WX7155), .SI(WX7154), .SE(n4474), .CLK(n5022), 
        .Q(WX7156) );
  SDFFX1 DFF_1016_Q_reg ( .D(WX7157), .SI(WX7156), .SE(n4473), .CLK(n5023), 
        .Q(WX7158) );
  SDFFX1 DFF_1017_Q_reg ( .D(WX7159), .SI(WX7158), .SE(n4473), .CLK(n5023), 
        .Q(WX7160) );
  SDFFX1 DFF_1018_Q_reg ( .D(WX7161), .SI(WX7160), .SE(n4472), .CLK(n5023), 
        .Q(WX7162) );
  SDFFX1 DFF_1019_Q_reg ( .D(WX7163), .SI(WX7162), .SE(n4471), .CLK(n5024), 
        .Q(WX7164) );
  SDFFX1 DFF_1020_Q_reg ( .D(WX7165), .SI(WX7164), .SE(n4471), .CLK(n5024), 
        .Q(WX7166) );
  SDFFX1 DFF_1021_Q_reg ( .D(WX7167), .SI(WX7166), .SE(n4470), .CLK(n5024), 
        .Q(WX7168) );
  SDFFX1 DFF_1022_Q_reg ( .D(WX7169), .SI(WX7168), .SE(n4469), .CLK(n5025), 
        .Q(WX7170) );
  SDFFX1 DFF_1023_Q_reg ( .D(WX7171), .SI(WX7170), .SE(n4469), .CLK(n5025), 
        .Q(WX7172) );
  SDFFX1 DFF_1024_Q_reg ( .D(WX7173), .SI(WX7172), .SE(n4468), .CLK(n5025), 
        .Q(WX7174), .QN(n3585) );
  SDFFX1 DFF_1025_Q_reg ( .D(WX7175), .SI(WX7174), .SE(n4485), .CLK(n5016), 
        .Q(WX7176), .QN(n3641) );
  SDFFX1 DFF_1026_Q_reg ( .D(WX7177), .SI(WX7176), .SE(n4485), .CLK(n5017), 
        .Q(WX7178), .QN(n3640) );
  SDFFX1 DFF_1027_Q_reg ( .D(WX7179), .SI(WX7178), .SE(n4485), .CLK(n5017), 
        .Q(WX7180), .QN(n3639) );
  SDFFX1 DFF_1028_Q_reg ( .D(WX7181), .SI(WX7180), .SE(n4485), .CLK(n5017), 
        .Q(WX7182) );
  SDFFX1 DFF_1029_Q_reg ( .D(WX7183), .SI(WX7182), .SE(n4484), .CLK(n5017), 
        .Q(WX7184), .QN(n3637) );
  SDFFX1 DFF_1030_Q_reg ( .D(WX7185), .SI(WX7184), .SE(n4484), .CLK(n5017), 
        .Q(test_so59), .QN(n8903) );
  SDFFX1 DFF_1031_Q_reg ( .D(WX7187), .SI(test_si60), .SE(n4368), .CLK(n5076), 
        .Q(WX7188), .QN(n3636) );
  SDFFX1 DFF_1032_Q_reg ( .D(WX7189), .SI(WX7188), .SE(n4483), .CLK(n5018), 
        .Q(WX7190), .QN(n8900) );
  SDFFX1 DFF_1033_Q_reg ( .D(WX7191), .SI(WX7190), .SE(n4483), .CLK(n5018), 
        .Q(WX7192), .QN(n3635) );
  SDFFX1 DFF_1034_Q_reg ( .D(WX7193), .SI(WX7192), .SE(n4482), .CLK(n5018), 
        .Q(WX7194) );
  SDFFX1 DFF_1035_Q_reg ( .D(WX7195), .SI(WX7194), .SE(n4482), .CLK(n5018), 
        .Q(WX7196), .QN(n3633) );
  SDFFX1 DFF_1036_Q_reg ( .D(WX7197), .SI(WX7196), .SE(n4481), .CLK(n5019), 
        .Q(WX7198), .QN(n3632) );
  SDFFX1 DFF_1037_Q_reg ( .D(WX7199), .SI(WX7198), .SE(n4481), .CLK(n5019), 
        .Q(WX7200), .QN(n3631) );
  SDFFX1 DFF_1038_Q_reg ( .D(WX7201), .SI(WX7200), .SE(n4480), .CLK(n5019), 
        .Q(WX7202), .QN(n3630) );
  SDFFX1 DFF_1039_Q_reg ( .D(WX7203), .SI(WX7202), .SE(n4479), .CLK(n5020), 
        .Q(WX7204), .QN(n3629) );
  SDFFX1 DFF_1040_Q_reg ( .D(WX7205), .SI(WX7204), .SE(n4478), .CLK(n5020), 
        .Q(WX7206), .QN(n8890) );
  SDFFX1 DFF_1041_Q_reg ( .D(WX7207), .SI(WX7206), .SE(n4478), .CLK(n5020), 
        .Q(WX7208), .QN(n8889) );
  SDFFX1 DFF_1042_Q_reg ( .D(WX7209), .SI(WX7208), .SE(n4477), .CLK(n5021), 
        .Q(WX7210), .QN(n8888) );
  SDFFX1 DFF_1043_Q_reg ( .D(WX7211), .SI(WX7210), .SE(n4476), .CLK(n5021), 
        .Q(WX7212), .QN(n8887) );
  SDFFX1 DFF_1044_Q_reg ( .D(WX7213), .SI(WX7212), .SE(n4476), .CLK(n5021), 
        .Q(WX7214), .QN(n8886) );
  SDFFX1 DFF_1045_Q_reg ( .D(WX7215), .SI(WX7214), .SE(n4475), .CLK(n5022), 
        .Q(WX7216), .QN(n8885) );
  SDFFX1 DFF_1046_Q_reg ( .D(WX7217), .SI(WX7216), .SE(n4475), .CLK(n5022), 
        .Q(WX7218), .QN(n8884) );
  SDFFX1 DFF_1047_Q_reg ( .D(WX7219), .SI(WX7218), .SE(n4474), .CLK(n5022), 
        .Q(test_so60) );
  SDFFX1 DFF_1048_Q_reg ( .D(WX7221), .SI(test_si61), .SE(n4473), .CLK(n5023), 
        .Q(WX7222), .QN(n8882) );
  SDFFX1 DFF_1049_Q_reg ( .D(WX7223), .SI(WX7222), .SE(n4472), .CLK(n5023), 
        .Q(WX7224), .QN(n8881) );
  SDFFX1 DFF_1050_Q_reg ( .D(WX7225), .SI(WX7224), .SE(n4472), .CLK(n5023), 
        .Q(WX7226), .QN(n8880) );
  SDFFX1 DFF_1051_Q_reg ( .D(WX7227), .SI(WX7226), .SE(n4471), .CLK(n5024), 
        .Q(WX7228), .QN(n8879) );
  SDFFX1 DFF_1052_Q_reg ( .D(WX7229), .SI(WX7228), .SE(n4470), .CLK(n5024), 
        .Q(WX7230), .QN(n8878) );
  SDFFX1 DFF_1053_Q_reg ( .D(WX7231), .SI(WX7230), .SE(n4470), .CLK(n5024), 
        .Q(WX7232), .QN(n8877) );
  SDFFX1 DFF_1054_Q_reg ( .D(WX7233), .SI(WX7232), .SE(n4469), .CLK(n5025), 
        .Q(WX7234), .QN(n8876) );
  SDFFX1 DFF_1055_Q_reg ( .D(WX7235), .SI(WX7234), .SE(n4468), .CLK(n5025), 
        .Q(WX7236), .QN(n8875) );
  SDFFX1 DFF_1056_Q_reg ( .D(WX7237), .SI(WX7236), .SE(n4468), .CLK(n5025), 
        .Q(WX7238) );
  SDFFX1 DFF_1057_Q_reg ( .D(WX7239), .SI(WX7238), .SE(n4467), .CLK(n5025), 
        .Q(WX7240) );
  SDFFX1 DFF_1058_Q_reg ( .D(WX7241), .SI(WX7240), .SE(n4467), .CLK(n5026), 
        .Q(WX7242) );
  SDFFX1 DFF_1059_Q_reg ( .D(WX7243), .SI(WX7242), .SE(n4467), .CLK(n5026), 
        .Q(WX7244) );
  SDFFX1 DFF_1060_Q_reg ( .D(WX7245), .SI(WX7244), .SE(n4466), .CLK(n5026), 
        .Q(WX7246), .QN(n3638) );
  SDFFX1 DFF_1061_Q_reg ( .D(WX7247), .SI(WX7246), .SE(n4466), .CLK(n5026), 
        .Q(WX7248) );
  SDFFX1 DFF_1062_Q_reg ( .D(WX7249), .SI(WX7248), .SE(n4484), .CLK(n5017), 
        .Q(WX7250), .QN(n8904) );
  SDFFX1 DFF_1063_Q_reg ( .D(WX7251), .SI(WX7250), .SE(n4484), .CLK(n5017), 
        .Q(WX7252) );
  SDFFX1 DFF_1064_Q_reg ( .D(WX7253), .SI(WX7252), .SE(n4483), .CLK(n5017), 
        .Q(test_so61), .QN(n8899) );
  SDFFX1 DFF_1065_Q_reg ( .D(WX7255), .SI(test_si62), .SE(n4483), .CLK(n5018), 
        .Q(WX7256) );
  SDFFX1 DFF_1066_Q_reg ( .D(WX7257), .SI(WX7256), .SE(n4482), .CLK(n5018), 
        .Q(WX7258), .QN(n3634) );
  SDFFX1 DFF_1067_Q_reg ( .D(WX7259), .SI(WX7258), .SE(n4482), .CLK(n5018), 
        .Q(WX7260) );
  SDFFX1 DFF_1068_Q_reg ( .D(WX7261), .SI(WX7260), .SE(n4481), .CLK(n5019), 
        .Q(WX7262) );
  SDFFX1 DFF_1069_Q_reg ( .D(WX7263), .SI(WX7262), .SE(n4480), .CLK(n5019), 
        .Q(WX7264) );
  SDFFX1 DFF_1070_Q_reg ( .D(WX7265), .SI(WX7264), .SE(n4480), .CLK(n5019), 
        .Q(WX7266) );
  SDFFX1 DFF_1071_Q_reg ( .D(WX7267), .SI(WX7266), .SE(n4479), .CLK(n5020), 
        .Q(WX7268) );
  SDFFX1 DFF_1072_Q_reg ( .D(WX7269), .SI(WX7268), .SE(n4478), .CLK(n5020), 
        .Q(WX7270), .QN(n3812) );
  SDFFX1 DFF_1073_Q_reg ( .D(WX7271), .SI(WX7270), .SE(n4478), .CLK(n5020), 
        .Q(WX7272), .QN(n3810) );
  SDFFX1 DFF_1074_Q_reg ( .D(WX7273), .SI(WX7272), .SE(n4477), .CLK(n5021), 
        .Q(WX7274), .QN(n3808) );
  SDFFX1 DFF_1075_Q_reg ( .D(WX7275), .SI(WX7274), .SE(n4476), .CLK(n5021), 
        .Q(WX7276), .QN(n3806) );
  SDFFX1 DFF_1076_Q_reg ( .D(WX7277), .SI(WX7276), .SE(n4476), .CLK(n5021), 
        .Q(WX7278), .QN(n3804) );
  SDFFX1 DFF_1077_Q_reg ( .D(WX7279), .SI(WX7278), .SE(n4475), .CLK(n5022), 
        .Q(WX7280) );
  SDFFX1 DFF_1078_Q_reg ( .D(WX7281), .SI(WX7280), .SE(n4474), .CLK(n5022), 
        .Q(WX7282), .QN(n3801) );
  SDFFX1 DFF_1079_Q_reg ( .D(WX7283), .SI(WX7282), .SE(n4474), .CLK(n5022), 
        .Q(WX7284), .QN(n8883) );
  SDFFX1 DFF_1080_Q_reg ( .D(WX7285), .SI(WX7284), .SE(n4473), .CLK(n5023), 
        .Q(WX7286), .QN(n3798) );
  SDFFX1 DFF_1081_Q_reg ( .D(WX7287), .SI(WX7286), .SE(n4472), .CLK(n5023), 
        .Q(test_so62) );
  SDFFX1 DFF_1082_Q_reg ( .D(WX7289), .SI(test_si63), .SE(n4472), .CLK(n5023), 
        .Q(WX7290), .QN(n3795) );
  SDFFX1 DFF_1083_Q_reg ( .D(WX7291), .SI(WX7290), .SE(n4471), .CLK(n5024), 
        .Q(WX7292), .QN(n3793) );
  SDFFX1 DFF_1084_Q_reg ( .D(WX7293), .SI(WX7292), .SE(n4470), .CLK(n5024), 
        .Q(WX7294), .QN(n3791) );
  SDFFX1 DFF_1085_Q_reg ( .D(WX7295), .SI(WX7294), .SE(n4470), .CLK(n5024), 
        .Q(WX7296), .QN(n3789) );
  SDFFX1 DFF_1086_Q_reg ( .D(WX7297), .SI(WX7296), .SE(n4469), .CLK(n5025), 
        .Q(WX7298), .QN(n3787) );
  SDFFX1 DFF_1087_Q_reg ( .D(WX7299), .SI(WX7298), .SE(n4468), .CLK(n5025), 
        .Q(WX7300), .QN(n3785) );
  SDFFX1 DFF_1088_Q_reg ( .D(WX7301), .SI(WX7300), .SE(n4468), .CLK(n5025), 
        .Q(WX7302), .QN(n4046) );
  SDFFX1 DFF_1089_Q_reg ( .D(WX7303), .SI(WX7302), .SE(n4467), .CLK(n5026), 
        .Q(WX7304), .QN(n4047) );
  SDFFX1 DFF_1090_Q_reg ( .D(WX7305), .SI(WX7304), .SE(n4467), .CLK(n5026), 
        .Q(WX7306), .QN(n4048) );
  SDFFX1 DFF_1091_Q_reg ( .D(WX7307), .SI(WX7306), .SE(n4467), .CLK(n5026), 
        .Q(WX7308), .QN(n4049) );
  SDFFX1 DFF_1092_Q_reg ( .D(WX7309), .SI(WX7308), .SE(n4466), .CLK(n5026), 
        .Q(WX7310), .QN(n4050) );
  SDFFX1 DFF_1093_Q_reg ( .D(WX7311), .SI(WX7310), .SE(n4466), .CLK(n5026), 
        .Q(WX7312), .QN(n4051) );
  SDFFX1 DFF_1094_Q_reg ( .D(WX7313), .SI(WX7312), .SE(n4466), .CLK(n5026), 
        .Q(WX7314), .QN(n4052) );
  SDFFX1 DFF_1095_Q_reg ( .D(WX7315), .SI(WX7314), .SE(n4466), .CLK(n5026), 
        .Q(WX7316), .QN(n4053) );
  SDFFX1 DFF_1096_Q_reg ( .D(WX7317), .SI(WX7316), .SE(n4465), .CLK(n5026), 
        .Q(WX7318), .QN(n4054) );
  SDFFX1 DFF_1097_Q_reg ( .D(WX7319), .SI(WX7318), .SE(n4465), .CLK(n5027), 
        .Q(WX7320), .QN(n4055) );
  SDFFX1 DFF_1098_Q_reg ( .D(WX7321), .SI(WX7320), .SE(n4465), .CLK(n5027), 
        .Q(test_so63) );
  SDFFX1 DFF_1099_Q_reg ( .D(WX7323), .SI(test_si64), .SE(n4482), .CLK(n5018), 
        .Q(WX7324), .QN(n4056) );
  SDFFX1 DFF_1100_Q_reg ( .D(WX7325), .SI(WX7324), .SE(n4481), .CLK(n5019), 
        .Q(WX7326), .QN(n4057) );
  SDFFX1 DFF_1101_Q_reg ( .D(WX7327), .SI(WX7326), .SE(n4480), .CLK(n5019), 
        .Q(WX7328), .QN(n4058) );
  SDFFX1 DFF_1102_Q_reg ( .D(WX7329), .SI(WX7328), .SE(n4479), .CLK(n5019), 
        .Q(WX7330), .QN(n4059) );
  SDFFX1 DFF_1103_Q_reg ( .D(WX7331), .SI(WX7330), .SE(n4479), .CLK(n5020), 
        .Q(WX7332), .QN(n3948) );
  SDFFX1 DFF_1104_Q_reg ( .D(WX7333), .SI(WX7332), .SE(n4478), .CLK(n5020), 
        .Q(WX7334), .QN(n4060) );
  SDFFX1 DFF_1105_Q_reg ( .D(WX7335), .SI(WX7334), .SE(n4477), .CLK(n5020), 
        .Q(WX7336), .QN(n4061) );
  SDFFX1 DFF_1106_Q_reg ( .D(WX7337), .SI(WX7336), .SE(n4477), .CLK(n5021), 
        .Q(WX7338), .QN(n4062) );
  SDFFX1 DFF_1107_Q_reg ( .D(WX7339), .SI(WX7338), .SE(n4476), .CLK(n5021), 
        .Q(WX7340), .QN(n4063) );
  SDFFX1 DFF_1108_Q_reg ( .D(WX7341), .SI(WX7340), .SE(n4475), .CLK(n5021), 
        .Q(WX7342), .QN(n3949) );
  SDFFX1 DFF_1109_Q_reg ( .D(WX7343), .SI(WX7342), .SE(n4475), .CLK(n5022), 
        .Q(WX7344), .QN(n4064) );
  SDFFX1 DFF_1110_Q_reg ( .D(WX7345), .SI(WX7344), .SE(n4474), .CLK(n5022), 
        .Q(WX7346), .QN(n4065) );
  SDFFX1 DFF_1111_Q_reg ( .D(WX7347), .SI(WX7346), .SE(n4473), .CLK(n5022), 
        .Q(WX7348), .QN(n4066) );
  SDFFX1 DFF_1112_Q_reg ( .D(WX7349), .SI(WX7348), .SE(n4473), .CLK(n5023), 
        .Q(WX7350), .QN(n4067) );
  SDFFX1 DFF_1113_Q_reg ( .D(WX7351), .SI(WX7350), .SE(n4472), .CLK(n5023), 
        .Q(WX7352), .QN(n4068) );
  SDFFX1 DFF_1114_Q_reg ( .D(WX7353), .SI(WX7352), .SE(n4471), .CLK(n5023), 
        .Q(WX7354), .QN(n4069) );
  SDFFX1 DFF_1115_Q_reg ( .D(WX7355), .SI(WX7354), .SE(n4471), .CLK(n5024), 
        .Q(test_so64) );
  SDFFX1 DFF_1116_Q_reg ( .D(WX7357), .SI(test_si65), .SE(n4470), .CLK(n5024), 
        .Q(WX7358), .QN(n4070) );
  SDFFX1 DFF_1117_Q_reg ( .D(WX7359), .SI(WX7358), .SE(n4469), .CLK(n5024), 
        .Q(WX7360), .QN(n4071) );
  SDFFX1 DFF_1118_Q_reg ( .D(WX7361), .SI(WX7360), .SE(n4469), .CLK(n5025), 
        .Q(WX7362), .QN(n4072) );
  SDFFX1 DFF_1119_Q_reg ( .D(WX7363), .SI(WX7362), .SE(n4468), .CLK(n5025), 
        .Q(WX7364), .QN(n3963) );
  SDFFX1 DFF_1120_Q_reg ( .D(WX7729), .SI(WX7364), .SE(n4372), .CLK(n5074), 
        .Q(CRC_OUT_4_0), .QN(DFF_1120_n1) );
  SDFFX1 DFF_1121_Q_reg ( .D(WX7731), .SI(CRC_OUT_4_0), .SE(n4372), .CLK(n5074), .Q(CRC_OUT_4_1), .QN(DFF_1121_n1) );
  SDFFX1 DFF_1122_Q_reg ( .D(WX7733), .SI(CRC_OUT_4_1), .SE(n4372), .CLK(n5074), .Q(CRC_OUT_4_2), .QN(DFF_1122_n1) );
  SDFFX1 DFF_1123_Q_reg ( .D(WX7735), .SI(CRC_OUT_4_2), .SE(n4372), .CLK(n5074), .Q(CRC_OUT_4_3), .QN(DFF_1123_n1) );
  SDFFX1 DFF_1124_Q_reg ( .D(WX7737), .SI(CRC_OUT_4_3), .SE(n4371), .CLK(n5074), .Q(CRC_OUT_4_4), .QN(DFF_1124_n1) );
  SDFFX1 DFF_1125_Q_reg ( .D(WX7739), .SI(CRC_OUT_4_4), .SE(n4371), .CLK(n5074), .Q(CRC_OUT_4_5), .QN(DFF_1125_n1) );
  SDFFX1 DFF_1126_Q_reg ( .D(WX7741), .SI(CRC_OUT_4_5), .SE(n4371), .CLK(n5074), .Q(CRC_OUT_4_6), .QN(DFF_1126_n1) );
  SDFFX1 DFF_1127_Q_reg ( .D(WX7743), .SI(CRC_OUT_4_6), .SE(n4371), .CLK(n5074), .Q(CRC_OUT_4_7), .QN(DFF_1127_n1) );
  SDFFX1 DFF_1128_Q_reg ( .D(WX7745), .SI(CRC_OUT_4_7), .SE(n4371), .CLK(n5074), .Q(CRC_OUT_4_8), .QN(DFF_1128_n1) );
  SDFFX1 DFF_1129_Q_reg ( .D(WX7747), .SI(CRC_OUT_4_8), .SE(n4371), .CLK(n5074), .Q(CRC_OUT_4_9), .QN(DFF_1129_n1) );
  SDFFX1 DFF_1130_Q_reg ( .D(WX7749), .SI(CRC_OUT_4_9), .SE(n4370), .CLK(n5075), .Q(CRC_OUT_4_10), .QN(DFF_1130_n1) );
  SDFFX1 DFF_1131_Q_reg ( .D(WX7751), .SI(CRC_OUT_4_10), .SE(n4370), .CLK(
        n5075), .Q(CRC_OUT_4_11), .QN(DFF_1131_n1) );
  SDFFX1 DFF_1132_Q_reg ( .D(WX7753), .SI(CRC_OUT_4_11), .SE(n4370), .CLK(
        n5075), .Q(test_so65) );
  SDFFX1 DFF_1133_Q_reg ( .D(WX7755), .SI(test_si66), .SE(n4370), .CLK(n5075), 
        .Q(CRC_OUT_4_13), .QN(DFF_1133_n1) );
  SDFFX1 DFF_1134_Q_reg ( .D(WX7757), .SI(CRC_OUT_4_13), .SE(n4370), .CLK(
        n5075), .Q(CRC_OUT_4_14), .QN(DFF_1134_n1) );
  SDFFX1 DFF_1135_Q_reg ( .D(WX7759), .SI(CRC_OUT_4_14), .SE(n4370), .CLK(
        n5075), .Q(CRC_OUT_4_15), .QN(DFF_1135_n1) );
  SDFFX1 DFF_1136_Q_reg ( .D(WX7761), .SI(CRC_OUT_4_15), .SE(n4369), .CLK(
        n5075), .Q(CRC_OUT_4_16), .QN(DFF_1136_n1) );
  SDFFX1 DFF_1137_Q_reg ( .D(WX7763), .SI(CRC_OUT_4_16), .SE(n4369), .CLK(
        n5075), .Q(CRC_OUT_4_17), .QN(DFF_1137_n1) );
  SDFFX1 DFF_1138_Q_reg ( .D(WX7765), .SI(CRC_OUT_4_17), .SE(n4369), .CLK(
        n5075), .Q(CRC_OUT_4_18), .QN(DFF_1138_n1) );
  SDFFX1 DFF_1139_Q_reg ( .D(WX7767), .SI(CRC_OUT_4_18), .SE(n4369), .CLK(
        n5075), .Q(CRC_OUT_4_19), .QN(DFF_1139_n1) );
  SDFFX1 DFF_1140_Q_reg ( .D(WX7769), .SI(CRC_OUT_4_19), .SE(n4369), .CLK(
        n5075), .Q(CRC_OUT_4_20), .QN(DFF_1140_n1) );
  SDFFX1 DFF_1141_Q_reg ( .D(WX7771), .SI(CRC_OUT_4_20), .SE(n4369), .CLK(
        n5075), .Q(CRC_OUT_4_21), .QN(DFF_1141_n1) );
  SDFFX1 DFF_1142_Q_reg ( .D(WX7773), .SI(CRC_OUT_4_21), .SE(n4368), .CLK(
        n5076), .Q(CRC_OUT_4_22), .QN(DFF_1142_n1) );
  SDFFX1 DFF_1143_Q_reg ( .D(WX7775), .SI(CRC_OUT_4_22), .SE(n4368), .CLK(
        n5076), .Q(CRC_OUT_4_23), .QN(DFF_1143_n1) );
  SDFFX1 DFF_1144_Q_reg ( .D(WX7777), .SI(CRC_OUT_4_23), .SE(n4368), .CLK(
        n5076), .Q(CRC_OUT_4_24), .QN(DFF_1144_n1) );
  SDFFX1 DFF_1145_Q_reg ( .D(WX7779), .SI(CRC_OUT_4_24), .SE(n4368), .CLK(
        n5076), .Q(CRC_OUT_4_25), .QN(DFF_1145_n1) );
  SDFFX1 DFF_1146_Q_reg ( .D(WX7781), .SI(CRC_OUT_4_25), .SE(n4465), .CLK(
        n5027), .Q(CRC_OUT_4_26), .QN(DFF_1146_n1) );
  SDFFX1 DFF_1147_Q_reg ( .D(WX7783), .SI(CRC_OUT_4_26), .SE(n4465), .CLK(
        n5027), .Q(CRC_OUT_4_27), .QN(DFF_1147_n1) );
  SDFFX1 DFF_1148_Q_reg ( .D(WX7785), .SI(CRC_OUT_4_27), .SE(n4465), .CLK(
        n5027), .Q(CRC_OUT_4_28), .QN(DFF_1148_n1) );
  SDFFX1 DFF_1149_Q_reg ( .D(WX7787), .SI(CRC_OUT_4_28), .SE(n4464), .CLK(
        n5027), .Q(test_so66) );
  SDFFX1 DFF_1150_Q_reg ( .D(WX7789), .SI(test_si67), .SE(n4464), .CLK(n5027), 
        .Q(CRC_OUT_4_30), .QN(DFF_1150_n1) );
  SDFFX1 DFF_1151_Q_reg ( .D(WX7791), .SI(CRC_OUT_4_30), .SE(n4464), .CLK(
        n5027), .Q(CRC_OUT_4_31), .QN(DFF_1151_n1) );
  SDFFX1 DFF_1152_Q_reg ( .D(n157), .SI(CRC_OUT_4_31), .SE(n4464), .CLK(n5027), 
        .Q(WX8243), .QN(n3933) );
  SDFFX1 DFF_1153_Q_reg ( .D(n158), .SI(WX8243), .SE(n4372), .CLK(n5074), .Q(
        n8411) );
  SDFFX1 DFF_1154_Q_reg ( .D(n159), .SI(n8411), .SE(n4459), .CLK(n5030), .Q(
        n8410) );
  SDFFX1 DFF_1155_Q_reg ( .D(n160), .SI(n8410), .SE(n4459), .CLK(n5030), .Q(
        n8409) );
  SDFFX1 DFF_1156_Q_reg ( .D(n161), .SI(n8409), .SE(n4459), .CLK(n5030), .Q(
        n8408) );
  SDFFX1 DFF_1157_Q_reg ( .D(n162), .SI(n8408), .SE(n4459), .CLK(n5029), .Q(
        n8407) );
  SDFFX1 DFF_1158_Q_reg ( .D(n163), .SI(n8407), .SE(n4460), .CLK(n5029), .Q(
        n8406) );
  SDFFX1 DFF_1159_Q_reg ( .D(n164), .SI(n8406), .SE(n4460), .CLK(n5029), .Q(
        n8405) );
  SDFFX1 DFF_1160_Q_reg ( .D(n165), .SI(n8405), .SE(n4460), .CLK(n5029), .Q(
        n8404) );
  SDFFX1 DFF_1161_Q_reg ( .D(n166), .SI(n8404), .SE(n4460), .CLK(n5029), .Q(
        n8403) );
  SDFFX1 DFF_1162_Q_reg ( .D(n167), .SI(n8403), .SE(n4460), .CLK(n5029), .Q(
        n8402) );
  SDFFX1 DFF_1163_Q_reg ( .D(n168), .SI(n8402), .SE(n4460), .CLK(n5029), .Q(
        n8401) );
  SDFFX1 DFF_1164_Q_reg ( .D(n169), .SI(n8401), .SE(n4461), .CLK(n5029), .Q(
        n8400) );
  SDFFX1 DFF_1165_Q_reg ( .D(n170), .SI(n8400), .SE(n4461), .CLK(n5029), .Q(
        n8399) );
  SDFFX1 DFF_1166_Q_reg ( .D(n171), .SI(n8399), .SE(n4461), .CLK(n5029), .Q(
        test_so67) );
  SDFFX1 DFF_1167_Q_reg ( .D(n172), .SI(test_si68), .SE(n4461), .CLK(n5029), 
        .Q(n8396) );
  SDFFX1 DFF_1168_Q_reg ( .D(n173), .SI(n8396), .SE(n4461), .CLK(n5029), .Q(
        n8395) );
  SDFFX1 DFF_1169_Q_reg ( .D(n174), .SI(n8395), .SE(n4461), .CLK(n5028), .Q(
        n8394) );
  SDFFX1 DFF_1170_Q_reg ( .D(n175), .SI(n8394), .SE(n4462), .CLK(n5028), .Q(
        n8393) );
  SDFFX1 DFF_1171_Q_reg ( .D(n176), .SI(n8393), .SE(n4462), .CLK(n5028), .Q(
        n8392) );
  SDFFX1 DFF_1172_Q_reg ( .D(n177), .SI(n8392), .SE(n4462), .CLK(n5028), .Q(
        n8391) );
  SDFFX1 DFF_1173_Q_reg ( .D(n178), .SI(n8391), .SE(n4462), .CLK(n5028), .Q(
        n8390) );
  SDFFX1 DFF_1174_Q_reg ( .D(n179), .SI(n8390), .SE(n4462), .CLK(n5028), .Q(
        n8389) );
  SDFFX1 DFF_1175_Q_reg ( .D(n180), .SI(n8389), .SE(n4462), .CLK(n5028), .Q(
        n8388) );
  SDFFX1 DFF_1176_Q_reg ( .D(n181), .SI(n8388), .SE(n4463), .CLK(n5028), .Q(
        n8387) );
  SDFFX1 DFF_1177_Q_reg ( .D(n182), .SI(n8387), .SE(n4463), .CLK(n5028), .Q(
        n8386) );
  SDFFX1 DFF_1178_Q_reg ( .D(n183), .SI(n8386), .SE(n4463), .CLK(n5028), .Q(
        n8385) );
  SDFFX1 DFF_1179_Q_reg ( .D(n184), .SI(n8385), .SE(n4463), .CLK(n5028), .Q(
        n8384) );
  SDFFX1 DFF_1180_Q_reg ( .D(n185), .SI(n8384), .SE(n4463), .CLK(n5028), .Q(
        n8383) );
  SDFFX1 DFF_1181_Q_reg ( .D(n186), .SI(n8383), .SE(n4463), .CLK(n5027), .Q(
        n8382) );
  SDFFX1 DFF_1182_Q_reg ( .D(n187), .SI(n8382), .SE(n4464), .CLK(n5027), .Q(
        n8381) );
  SDFFX1 DFF_1183_Q_reg ( .D(WX8304), .SI(n8381), .SE(n4464), .CLK(n5027), .Q(
        test_so68) );
  SDFFX1 DFF_1184_Q_reg ( .D(WX8402), .SI(test_si69), .SE(n4486), .CLK(n5016), 
        .Q(n8378), .QN(n8874) );
  SDFFX1 DFF_1185_Q_reg ( .D(WX8404), .SI(n8378), .SE(n4486), .CLK(n5016), .Q(
        n8377), .QN(n8871) );
  SDFFX1 DFF_1186_Q_reg ( .D(WX8406), .SI(n8377), .SE(n4459), .CLK(n5030), .Q(
        n8376), .QN(n8870) );
  SDFFX1 DFF_1187_Q_reg ( .D(WX8408), .SI(n8376), .SE(n4458), .CLK(n5030), .Q(
        n8375), .QN(n8867) );
  SDFFX1 DFF_1188_Q_reg ( .D(WX8410), .SI(n8375), .SE(n4458), .CLK(n5030), .Q(
        n8374), .QN(n8866) );
  SDFFX1 DFF_1189_Q_reg ( .D(WX8412), .SI(n8374), .SE(n4373), .CLK(n5073), .Q(
        n8373), .QN(n8865) );
  SDFFX1 DFF_1190_Q_reg ( .D(WX8414), .SI(n8373), .SE(n4457), .CLK(n5031), .Q(
        n8372), .QN(n8864) );
  SDFFX1 DFF_1191_Q_reg ( .D(WX8416), .SI(n8372), .SE(n4457), .CLK(n5031), .Q(
        n8371), .QN(n8863) );
  SDFFX1 DFF_1192_Q_reg ( .D(WX8418), .SI(n8371), .SE(n4455), .CLK(n5031), .Q(
        n8370), .QN(n8862) );
  SDFFX1 DFF_1193_Q_reg ( .D(WX8420), .SI(n8370), .SE(n4455), .CLK(n5032), .Q(
        n8369), .QN(n8861) );
  SDFFX1 DFF_1194_Q_reg ( .D(WX8422), .SI(n8369), .SE(n4454), .CLK(n5032), .Q(
        n8368), .QN(n8860) );
  SDFFX1 DFF_1195_Q_reg ( .D(WX8424), .SI(n8368), .SE(n4454), .CLK(n5032), .Q(
        n8367), .QN(n8859) );
  SDFFX1 DFF_1196_Q_reg ( .D(WX8426), .SI(n8367), .SE(n4453), .CLK(n5033), .Q(
        n8366), .QN(n8858) );
  SDFFX1 DFF_1197_Q_reg ( .D(WX8428), .SI(n8366), .SE(n4453), .CLK(n5033), .Q(
        n8365), .QN(n8857) );
  SDFFX1 DFF_1198_Q_reg ( .D(WX8430), .SI(n8365), .SE(n4451), .CLK(n5033), .Q(
        n8364), .QN(n8856) );
  SDFFX1 DFF_1199_Q_reg ( .D(WX8432), .SI(n8364), .SE(n4451), .CLK(n5034), .Q(
        n8363), .QN(n8855) );
  SDFFX1 DFF_1200_Q_reg ( .D(WX8434), .SI(n8363), .SE(n4372), .CLK(n5074), .Q(
        test_so69) );
  SDFFX1 DFF_1201_Q_reg ( .D(WX8436), .SI(test_si70), .SE(n4450), .CLK(n5034), 
        .Q(WX8437) );
  SDFFX1 DFF_1202_Q_reg ( .D(WX8438), .SI(WX8437), .SE(n4449), .CLK(n5034), 
        .Q(WX8439) );
  SDFFX1 DFF_1203_Q_reg ( .D(WX8440), .SI(WX8439), .SE(n4449), .CLK(n5035), 
        .Q(WX8441) );
  SDFFX1 DFF_1204_Q_reg ( .D(WX8442), .SI(WX8441), .SE(n4448), .CLK(n5035), 
        .Q(WX8443) );
  SDFFX1 DFF_1205_Q_reg ( .D(WX8444), .SI(WX8443), .SE(n4447), .CLK(n5035), 
        .Q(WX8445) );
  SDFFX1 DFF_1206_Q_reg ( .D(WX8446), .SI(WX8445), .SE(n4447), .CLK(n5036), 
        .Q(WX8447) );
  SDFFX1 DFF_1207_Q_reg ( .D(WX8448), .SI(WX8447), .SE(n4446), .CLK(n5036), 
        .Q(WX8449) );
  SDFFX1 DFF_1208_Q_reg ( .D(WX8450), .SI(WX8449), .SE(n4445), .CLK(n5036), 
        .Q(WX8451) );
  SDFFX1 DFF_1209_Q_reg ( .D(WX8452), .SI(WX8451), .SE(n4445), .CLK(n5037), 
        .Q(WX8453) );
  SDFFX1 DFF_1210_Q_reg ( .D(WX8454), .SI(WX8453), .SE(n4444), .CLK(n5037), 
        .Q(WX8455) );
  SDFFX1 DFF_1211_Q_reg ( .D(WX8456), .SI(WX8455), .SE(n4443), .CLK(n5037), 
        .Q(WX8457) );
  SDFFX1 DFF_1212_Q_reg ( .D(WX8458), .SI(WX8457), .SE(n4487), .CLK(n5016), 
        .Q(WX8459) );
  SDFFX1 DFF_1213_Q_reg ( .D(WX8460), .SI(WX8459), .SE(n4487), .CLK(n5016), 
        .Q(WX8461) );
  SDFFX1 DFF_1214_Q_reg ( .D(WX8462), .SI(WX8461), .SE(n4487), .CLK(n5016), 
        .Q(WX8463) );
  SDFFX1 DFF_1215_Q_reg ( .D(WX8464), .SI(WX8463), .SE(n4486), .CLK(n5016), 
        .Q(WX8465) );
  SDFFX1 DFF_1216_Q_reg ( .D(WX8466), .SI(WX8465), .SE(n4486), .CLK(n5016), 
        .Q(WX8467), .QN(n3584) );
  SDFFX1 DFF_1217_Q_reg ( .D(WX8468), .SI(WX8467), .SE(n4486), .CLK(n5016), 
        .Q(test_so70), .QN(n8872) );
  SDFFX1 DFF_1218_Q_reg ( .D(WX8470), .SI(test_si71), .SE(n4459), .CLK(n5030), 
        .Q(WX8471), .QN(n3628) );
  SDFFX1 DFF_1219_Q_reg ( .D(WX8472), .SI(WX8471), .SE(n4458), .CLK(n5030), 
        .Q(WX8473), .QN(n8869) );
  SDFFX1 DFF_1220_Q_reg ( .D(WX8474), .SI(WX8473), .SE(n4458), .CLK(n5030), 
        .Q(WX8475), .QN(n3627) );
  SDFFX1 DFF_1221_Q_reg ( .D(WX8476), .SI(WX8475), .SE(n4458), .CLK(n5030), 
        .Q(WX8477) );
  SDFFX1 DFF_1222_Q_reg ( .D(WX8478), .SI(WX8477), .SE(n4457), .CLK(n5031), 
        .Q(WX8479), .QN(n3625) );
  SDFFX1 DFF_1223_Q_reg ( .D(WX8480), .SI(WX8479), .SE(n4456), .CLK(n5031), 
        .Q(WX8481), .QN(n3624) );
  SDFFX1 DFF_1224_Q_reg ( .D(WX8482), .SI(WX8481), .SE(n4456), .CLK(n5031), 
        .Q(WX8483), .QN(n3623) );
  SDFFX1 DFF_1225_Q_reg ( .D(WX8484), .SI(WX8483), .SE(n4455), .CLK(n5032), 
        .Q(WX8485), .QN(n3622) );
  SDFFX1 DFF_1226_Q_reg ( .D(WX8486), .SI(WX8485), .SE(n4455), .CLK(n5032), 
        .Q(WX8487), .QN(n3621) );
  SDFFX1 DFF_1227_Q_reg ( .D(WX8488), .SI(WX8487), .SE(n4454), .CLK(n5032), 
        .Q(WX8489), .QN(n3620) );
  SDFFX1 DFF_1228_Q_reg ( .D(WX8490), .SI(WX8489), .SE(n4453), .CLK(n5033), 
        .Q(WX8491), .QN(n3619) );
  SDFFX1 DFF_1229_Q_reg ( .D(WX8492), .SI(WX8491), .SE(n4452), .CLK(n5033), 
        .Q(WX8493), .QN(n3618) );
  SDFFX1 DFF_1230_Q_reg ( .D(WX8494), .SI(WX8493), .SE(n4452), .CLK(n5033), 
        .Q(WX8495), .QN(n3617) );
  SDFFX1 DFF_1231_Q_reg ( .D(WX8496), .SI(WX8495), .SE(n4451), .CLK(n5034), 
        .Q(WX8497), .QN(n3616) );
  SDFFX1 DFF_1232_Q_reg ( .D(WX8498), .SI(WX8497), .SE(n4451), .CLK(n5034), 
        .Q(WX8499), .QN(n8854) );
  SDFFX1 DFF_1233_Q_reg ( .D(WX8500), .SI(WX8499), .SE(n4450), .CLK(n5034), 
        .Q(WX8501), .QN(n8853) );
  SDFFX1 DFF_1234_Q_reg ( .D(WX8502), .SI(WX8501), .SE(n4449), .CLK(n5035), 
        .Q(test_so71) );
  SDFFX1 DFF_1235_Q_reg ( .D(WX8504), .SI(test_si72), .SE(n4449), .CLK(n5035), 
        .Q(WX8505), .QN(n8851) );
  SDFFX1 DFF_1236_Q_reg ( .D(WX8506), .SI(WX8505), .SE(n4448), .CLK(n5035), 
        .Q(WX8507), .QN(n8850) );
  SDFFX1 DFF_1237_Q_reg ( .D(WX8508), .SI(WX8507), .SE(n4447), .CLK(n5036), 
        .Q(WX8509), .QN(n8849) );
  SDFFX1 DFF_1238_Q_reg ( .D(WX8510), .SI(WX8509), .SE(n4447), .CLK(n5036), 
        .Q(WX8511), .QN(n8848) );
  SDFFX1 DFF_1239_Q_reg ( .D(WX8512), .SI(WX8511), .SE(n4446), .CLK(n5036), 
        .Q(WX8513), .QN(n8847) );
  SDFFX1 DFF_1240_Q_reg ( .D(WX8514), .SI(WX8513), .SE(n4445), .CLK(n5037), 
        .Q(WX8515), .QN(n8846) );
  SDFFX1 DFF_1241_Q_reg ( .D(WX8516), .SI(WX8515), .SE(n4445), .CLK(n5037), 
        .Q(WX8517), .QN(n8845) );
  SDFFX1 DFF_1242_Q_reg ( .D(WX8518), .SI(WX8517), .SE(n4444), .CLK(n5037), 
        .Q(WX8519), .QN(n8844) );
  SDFFX1 DFF_1243_Q_reg ( .D(WX8520), .SI(WX8519), .SE(n4443), .CLK(n5038), 
        .Q(WX8521), .QN(n8843) );
  SDFFX1 DFF_1244_Q_reg ( .D(WX8522), .SI(WX8521), .SE(n4443), .CLK(n5038), 
        .Q(WX8523), .QN(n8842) );
  SDFFX1 DFF_1245_Q_reg ( .D(WX8524), .SI(WX8523), .SE(n4442), .CLK(n5038), 
        .Q(WX8525), .QN(n8841) );
  SDFFX1 DFF_1246_Q_reg ( .D(WX8526), .SI(WX8525), .SE(n4442), .CLK(n5038), 
        .Q(WX8527), .QN(n8840) );
  SDFFX1 DFF_1247_Q_reg ( .D(WX8528), .SI(WX8527), .SE(n4441), .CLK(n5039), 
        .Q(WX8529), .QN(n8839) );
  SDFFX1 DFF_1248_Q_reg ( .D(WX8530), .SI(WX8529), .SE(n4441), .CLK(n5039), 
        .Q(WX8531) );
  SDFFX1 DFF_1249_Q_reg ( .D(WX8532), .SI(WX8531), .SE(n4440), .CLK(n5039), 
        .Q(WX8533), .QN(n8873) );
  SDFFX1 DFF_1250_Q_reg ( .D(WX8534), .SI(WX8533), .SE(n4440), .CLK(n5039), 
        .Q(WX8535) );
  SDFFX1 DFF_1251_Q_reg ( .D(WX8536), .SI(WX8535), .SE(n4440), .CLK(n5039), 
        .Q(test_so72), .QN(n8868) );
  SDFFX1 DFF_1252_Q_reg ( .D(WX8538), .SI(test_si73), .SE(n4458), .CLK(n5030), 
        .Q(WX8539) );
  SDFFX1 DFF_1253_Q_reg ( .D(WX8540), .SI(WX8539), .SE(n4457), .CLK(n5030), 
        .Q(WX8541), .QN(n3626) );
  SDFFX1 DFF_1254_Q_reg ( .D(WX8542), .SI(WX8541), .SE(n4457), .CLK(n5031), 
        .Q(WX8543) );
  SDFFX1 DFF_1255_Q_reg ( .D(WX8544), .SI(WX8543), .SE(n4456), .CLK(n5031), 
        .Q(WX8545) );
  SDFFX1 DFF_1256_Q_reg ( .D(WX8546), .SI(WX8545), .SE(n4456), .CLK(n5031), 
        .Q(WX8547) );
  SDFFX1 DFF_1257_Q_reg ( .D(WX8548), .SI(WX8547), .SE(n4455), .CLK(n5032), 
        .Q(WX8549) );
  SDFFX1 DFF_1258_Q_reg ( .D(WX8550), .SI(WX8549), .SE(n4454), .CLK(n5032), 
        .Q(WX8551) );
  SDFFX1 DFF_1259_Q_reg ( .D(WX8552), .SI(WX8551), .SE(n4454), .CLK(n5032), 
        .Q(WX8553) );
  SDFFX1 DFF_1260_Q_reg ( .D(WX8554), .SI(WX8553), .SE(n4453), .CLK(n5033), 
        .Q(WX8555) );
  SDFFX1 DFF_1261_Q_reg ( .D(WX8556), .SI(WX8555), .SE(n4452), .CLK(n5033), 
        .Q(WX8557) );
  SDFFX1 DFF_1262_Q_reg ( .D(WX8558), .SI(WX8557), .SE(n4452), .CLK(n5033), 
        .Q(WX8559) );
  SDFFX1 DFF_1263_Q_reg ( .D(WX8560), .SI(WX8559), .SE(n4451), .CLK(n5034), 
        .Q(WX8561) );
  SDFFX1 DFF_1264_Q_reg ( .D(WX8562), .SI(WX8561), .SE(n4450), .CLK(n5034), 
        .Q(WX8563) );
  SDFFX1 DFF_1265_Q_reg ( .D(WX8564), .SI(WX8563), .SE(n4450), .CLK(n5034), 
        .Q(WX8565), .QN(n3782) );
  SDFFX1 DFF_1266_Q_reg ( .D(WX8566), .SI(WX8565), .SE(n4449), .CLK(n5035), 
        .Q(WX8567), .QN(n8852) );
  SDFFX1 DFF_1267_Q_reg ( .D(WX8568), .SI(WX8567), .SE(n4448), .CLK(n5035), 
        .Q(WX8569), .QN(n3779) );
  SDFFX1 DFF_1268_Q_reg ( .D(WX8570), .SI(WX8569), .SE(n4448), .CLK(n5035), 
        .Q(test_so73) );
  SDFFX1 DFF_1269_Q_reg ( .D(WX8572), .SI(test_si74), .SE(n4447), .CLK(n5036), 
        .Q(WX8573), .QN(n3776) );
  SDFFX1 DFF_1270_Q_reg ( .D(WX8574), .SI(WX8573), .SE(n4446), .CLK(n5036), 
        .Q(WX8575), .QN(n3774) );
  SDFFX1 DFF_1271_Q_reg ( .D(WX8576), .SI(WX8575), .SE(n4446), .CLK(n5036), 
        .Q(WX8577), .QN(n3772) );
  SDFFX1 DFF_1272_Q_reg ( .D(WX8578), .SI(WX8577), .SE(n4445), .CLK(n5037), 
        .Q(WX8579), .QN(n3770) );
  SDFFX1 DFF_1273_Q_reg ( .D(WX8580), .SI(WX8579), .SE(n4444), .CLK(n5037), 
        .Q(WX8581), .QN(n3768) );
  SDFFX1 DFF_1274_Q_reg ( .D(WX8582), .SI(WX8581), .SE(n4444), .CLK(n5037), 
        .Q(WX8583), .QN(n3766) );
  SDFFX1 DFF_1275_Q_reg ( .D(WX8584), .SI(WX8583), .SE(n4443), .CLK(n5038), 
        .Q(WX8585), .QN(n3764) );
  SDFFX1 DFF_1276_Q_reg ( .D(WX8586), .SI(WX8585), .SE(n4443), .CLK(n5038), 
        .Q(WX8587), .QN(n3762) );
  SDFFX1 DFF_1277_Q_reg ( .D(WX8588), .SI(WX8587), .SE(n4442), .CLK(n5038), 
        .Q(WX8589), .QN(n3760) );
  SDFFX1 DFF_1278_Q_reg ( .D(WX8590), .SI(WX8589), .SE(n4442), .CLK(n5038), 
        .Q(WX8591), .QN(n3758) );
  SDFFX1 DFF_1279_Q_reg ( .D(WX8592), .SI(WX8591), .SE(n4441), .CLK(n5039), 
        .Q(WX8593), .QN(n3756) );
  SDFFX1 DFF_1280_Q_reg ( .D(WX8594), .SI(WX8593), .SE(n4441), .CLK(n5039), 
        .Q(WX8595), .QN(n4020) );
  SDFFX1 DFF_1281_Q_reg ( .D(WX8596), .SI(WX8595), .SE(n4440), .CLK(n5039), 
        .Q(WX8597), .QN(n4021) );
  SDFFX1 DFF_1282_Q_reg ( .D(WX8598), .SI(WX8597), .SE(n4440), .CLK(n5039), 
        .Q(WX8599), .QN(n4022) );
  SDFFX1 DFF_1283_Q_reg ( .D(WX8600), .SI(WX8599), .SE(n4440), .CLK(n5039), 
        .Q(WX8601), .QN(n4023) );
  SDFFX1 DFF_1284_Q_reg ( .D(WX8602), .SI(WX8601), .SE(n4439), .CLK(n5039), 
        .Q(WX8603), .QN(n4024) );
  SDFFX1 DFF_1285_Q_reg ( .D(WX8604), .SI(WX8603), .SE(n4439), .CLK(n5040), 
        .Q(test_so74) );
  SDFFX1 DFF_1286_Q_reg ( .D(WX8606), .SI(test_si75), .SE(n4457), .CLK(n5031), 
        .Q(WX8607), .QN(n4025) );
  SDFFX1 DFF_1287_Q_reg ( .D(WX8608), .SI(WX8607), .SE(n4456), .CLK(n5031), 
        .Q(WX8609), .QN(n4026) );
  SDFFX1 DFF_1288_Q_reg ( .D(WX8610), .SI(WX8609), .SE(n4456), .CLK(n5031), 
        .Q(WX8611), .QN(n4027) );
  SDFFX1 DFF_1289_Q_reg ( .D(WX8612), .SI(WX8611), .SE(n4455), .CLK(n5032), 
        .Q(WX8613), .QN(n4028) );
  SDFFX1 DFF_1290_Q_reg ( .D(WX8614), .SI(WX8613), .SE(n4454), .CLK(n5032), 
        .Q(WX8615), .QN(n4029) );
  SDFFX1 DFF_1291_Q_reg ( .D(WX8616), .SI(WX8615), .SE(n4453), .CLK(n5032), 
        .Q(WX8617), .QN(n4030) );
  SDFFX1 DFF_1292_Q_reg ( .D(WX8618), .SI(WX8617), .SE(n4453), .CLK(n5033), 
        .Q(WX8619), .QN(n4031) );
  SDFFX1 DFF_1293_Q_reg ( .D(WX8620), .SI(WX8619), .SE(n4452), .CLK(n5033), 
        .Q(WX8621), .QN(n4032) );
  SDFFX1 DFF_1294_Q_reg ( .D(WX8622), .SI(WX8621), .SE(n4452), .CLK(n5033), 
        .Q(WX8623), .QN(n4033) );
  SDFFX1 DFF_1295_Q_reg ( .D(WX8624), .SI(WX8623), .SE(n4451), .CLK(n5034), 
        .Q(WX8625), .QN(n3945) );
  SDFFX1 DFF_1296_Q_reg ( .D(WX8626), .SI(WX8625), .SE(n4450), .CLK(n5034), 
        .Q(WX8627), .QN(n4034) );
  SDFFX1 DFF_1297_Q_reg ( .D(WX8628), .SI(WX8627), .SE(n4450), .CLK(n5034), 
        .Q(WX8629), .QN(n4035) );
  SDFFX1 DFF_1298_Q_reg ( .D(WX8630), .SI(WX8629), .SE(n4449), .CLK(n5035), 
        .Q(WX8631), .QN(n4036) );
  SDFFX1 DFF_1299_Q_reg ( .D(WX8632), .SI(WX8631), .SE(n4448), .CLK(n5035), 
        .Q(WX8633), .QN(n4037) );
  SDFFX1 DFF_1300_Q_reg ( .D(WX8634), .SI(WX8633), .SE(n4448), .CLK(n5035), 
        .Q(WX8635), .QN(n3946) );
  SDFFX1 DFF_1301_Q_reg ( .D(WX8636), .SI(WX8635), .SE(n4447), .CLK(n5036), 
        .Q(WX8637), .QN(n4038) );
  SDFFX1 DFF_1302_Q_reg ( .D(WX8638), .SI(WX8637), .SE(n4446), .CLK(n5036), 
        .Q(test_so75) );
  SDFFX1 DFF_1303_Q_reg ( .D(WX8640), .SI(test_si76), .SE(n4446), .CLK(n5036), 
        .Q(WX8641), .QN(n4039) );
  SDFFX1 DFF_1304_Q_reg ( .D(WX8642), .SI(WX8641), .SE(n4445), .CLK(n5037), 
        .Q(WX8643), .QN(n4040) );
  SDFFX1 DFF_1305_Q_reg ( .D(WX8644), .SI(WX8643), .SE(n4444), .CLK(n5037), 
        .Q(WX8645), .QN(n4041) );
  SDFFX1 DFF_1306_Q_reg ( .D(WX8646), .SI(WX8645), .SE(n4444), .CLK(n5037), 
        .Q(WX8647), .QN(n4042) );
  SDFFX1 DFF_1307_Q_reg ( .D(WX8648), .SI(WX8647), .SE(n4443), .CLK(n5038), 
        .Q(WX8649), .QN(n3947) );
  SDFFX1 DFF_1308_Q_reg ( .D(WX8650), .SI(WX8649), .SE(n4442), .CLK(n5038), 
        .Q(WX8651), .QN(n4043) );
  SDFFX1 DFF_1309_Q_reg ( .D(WX8652), .SI(WX8651), .SE(n4442), .CLK(n5038), 
        .Q(WX8653), .QN(n4044) );
  SDFFX1 DFF_1310_Q_reg ( .D(WX8654), .SI(WX8653), .SE(n4441), .CLK(n5038), 
        .Q(WX8655), .QN(n4045) );
  SDFFX1 DFF_1311_Q_reg ( .D(WX8656), .SI(WX8655), .SE(n4441), .CLK(n5039), 
        .Q(WX8657), .QN(n3962) );
  SDFFX1 DFF_1312_Q_reg ( .D(WX9022), .SI(WX8657), .SE(n4377), .CLK(n5071), 
        .Q(CRC_OUT_3_0), .QN(DFF_1312_n1) );
  SDFFX1 DFF_1313_Q_reg ( .D(WX9024), .SI(CRC_OUT_3_0), .SE(n4377), .CLK(n5071), .Q(CRC_OUT_3_1), .QN(DFF_1313_n1) );
  SDFFX1 DFF_1314_Q_reg ( .D(WX9026), .SI(CRC_OUT_3_1), .SE(n4377), .CLK(n5071), .Q(CRC_OUT_3_2), .QN(DFF_1314_n1) );
  SDFFX1 DFF_1315_Q_reg ( .D(WX9028), .SI(CRC_OUT_3_2), .SE(n4377), .CLK(n5071), .Q(CRC_OUT_3_3), .QN(DFF_1315_n1) );
  SDFFX1 DFF_1316_Q_reg ( .D(WX9030), .SI(CRC_OUT_3_3), .SE(n4377), .CLK(n5071), .Q(CRC_OUT_3_4), .QN(DFF_1316_n1) );
  SDFFX1 DFF_1317_Q_reg ( .D(WX9032), .SI(CRC_OUT_3_4), .SE(n4376), .CLK(n5072), .Q(CRC_OUT_3_5), .QN(DFF_1317_n1) );
  SDFFX1 DFF_1318_Q_reg ( .D(WX9034), .SI(CRC_OUT_3_5), .SE(n4376), .CLK(n5072), .Q(CRC_OUT_3_6), .QN(DFF_1318_n1) );
  SDFFX1 DFF_1319_Q_reg ( .D(WX9036), .SI(CRC_OUT_3_6), .SE(n4376), .CLK(n5072), .Q(test_so76) );
  SDFFX1 DFF_1320_Q_reg ( .D(WX9038), .SI(test_si77), .SE(n4376), .CLK(n5072), 
        .Q(CRC_OUT_3_8), .QN(DFF_1320_n1) );
  SDFFX1 DFF_1321_Q_reg ( .D(WX9040), .SI(CRC_OUT_3_8), .SE(n4376), .CLK(n5072), .Q(CRC_OUT_3_9), .QN(DFF_1321_n1) );
  SDFFX1 DFF_1322_Q_reg ( .D(WX9042), .SI(CRC_OUT_3_9), .SE(n4376), .CLK(n5072), .Q(CRC_OUT_3_10), .QN(DFF_1322_n1) );
  SDFFX1 DFF_1323_Q_reg ( .D(WX9044), .SI(CRC_OUT_3_10), .SE(n4375), .CLK(
        n5072), .Q(CRC_OUT_3_11), .QN(DFF_1323_n1) );
  SDFFX1 DFF_1324_Q_reg ( .D(WX9046), .SI(CRC_OUT_3_11), .SE(n4375), .CLK(
        n5072), .Q(CRC_OUT_3_12), .QN(DFF_1324_n1) );
  SDFFX1 DFF_1325_Q_reg ( .D(WX9048), .SI(CRC_OUT_3_12), .SE(n4375), .CLK(
        n5072), .Q(CRC_OUT_3_13), .QN(DFF_1325_n1) );
  SDFFX1 DFF_1326_Q_reg ( .D(WX9050), .SI(CRC_OUT_3_13), .SE(n4375), .CLK(
        n5072), .Q(CRC_OUT_3_14), .QN(DFF_1326_n1) );
  SDFFX1 DFF_1327_Q_reg ( .D(WX9052), .SI(CRC_OUT_3_14), .SE(n4375), .CLK(
        n5072), .Q(CRC_OUT_3_15), .QN(DFF_1327_n1) );
  SDFFX1 DFF_1328_Q_reg ( .D(WX9054), .SI(CRC_OUT_3_15), .SE(n4375), .CLK(
        n5072), .Q(CRC_OUT_3_16), .QN(DFF_1328_n1) );
  SDFFX1 DFF_1329_Q_reg ( .D(WX9056), .SI(CRC_OUT_3_16), .SE(n4374), .CLK(
        n5073), .Q(CRC_OUT_3_17), .QN(DFF_1329_n1) );
  SDFFX1 DFF_1330_Q_reg ( .D(WX9058), .SI(CRC_OUT_3_17), .SE(n4374), .CLK(
        n5073), .Q(CRC_OUT_3_18), .QN(DFF_1330_n1) );
  SDFFX1 DFF_1331_Q_reg ( .D(WX9060), .SI(CRC_OUT_3_18), .SE(n4374), .CLK(
        n5073), .Q(CRC_OUT_3_19), .QN(DFF_1331_n1) );
  SDFFX1 DFF_1332_Q_reg ( .D(WX9062), .SI(CRC_OUT_3_19), .SE(n4374), .CLK(
        n5073), .Q(CRC_OUT_3_20), .QN(DFF_1332_n1) );
  SDFFX1 DFF_1333_Q_reg ( .D(WX9064), .SI(CRC_OUT_3_20), .SE(n4374), .CLK(
        n5073), .Q(CRC_OUT_3_21), .QN(DFF_1333_n1) );
  SDFFX1 DFF_1334_Q_reg ( .D(WX9066), .SI(CRC_OUT_3_21), .SE(n4374), .CLK(
        n5073), .Q(CRC_OUT_3_22), .QN(DFF_1334_n1) );
  SDFFX1 DFF_1335_Q_reg ( .D(WX9068), .SI(CRC_OUT_3_22), .SE(n4373), .CLK(
        n5073), .Q(CRC_OUT_3_23), .QN(DFF_1335_n1) );
  SDFFX1 DFF_1336_Q_reg ( .D(WX9070), .SI(CRC_OUT_3_23), .SE(n4373), .CLK(
        n5073), .Q(test_so77) );
  SDFFX1 DFF_1337_Q_reg ( .D(WX9072), .SI(test_si78), .SE(n4373), .CLK(n5073), 
        .Q(CRC_OUT_3_25), .QN(DFF_1337_n1) );
  SDFFX1 DFF_1338_Q_reg ( .D(WX9074), .SI(CRC_OUT_3_25), .SE(n4373), .CLK(
        n5073), .Q(CRC_OUT_3_26), .QN(DFF_1338_n1) );
  SDFFX1 DFF_1339_Q_reg ( .D(WX9076), .SI(CRC_OUT_3_26), .SE(n4373), .CLK(
        n5073), .Q(CRC_OUT_3_27), .QN(DFF_1339_n1) );
  SDFFX1 DFF_1340_Q_reg ( .D(WX9078), .SI(CRC_OUT_3_27), .SE(n4439), .CLK(
        n5040), .Q(CRC_OUT_3_28), .QN(DFF_1340_n1) );
  SDFFX1 DFF_1341_Q_reg ( .D(WX9080), .SI(CRC_OUT_3_28), .SE(n4439), .CLK(
        n5040), .Q(CRC_OUT_3_29), .QN(DFF_1341_n1) );
  SDFFX1 DFF_1342_Q_reg ( .D(WX9082), .SI(CRC_OUT_3_29), .SE(n4439), .CLK(
        n5040), .Q(CRC_OUT_3_30), .QN(DFF_1342_n1) );
  SDFFX1 DFF_1343_Q_reg ( .D(WX9084), .SI(CRC_OUT_3_30), .SE(n4439), .CLK(
        n5040), .Q(CRC_OUT_3_31), .QN(DFF_1343_n1) );
  SDFFX1 DFF_1344_Q_reg ( .D(n188), .SI(CRC_OUT_3_31), .SE(n4438), .CLK(n5040), 
        .Q(WX9536), .QN(n3932) );
  SDFFX1 DFF_1345_Q_reg ( .D(n189), .SI(WX9536), .SE(n4433), .CLK(n5043), .Q(
        n8353) );
  SDFFX1 DFF_1346_Q_reg ( .D(n190), .SI(n8353), .SE(n4433), .CLK(n5042), .Q(
        n8352) );
  SDFFX1 DFF_1347_Q_reg ( .D(n191), .SI(n8352), .SE(n4434), .CLK(n5042), .Q(
        n8351) );
  SDFFX1 DFF_1348_Q_reg ( .D(n192), .SI(n8351), .SE(n4434), .CLK(n5042), .Q(
        n8350) );
  SDFFX1 DFF_1349_Q_reg ( .D(n193), .SI(n8350), .SE(n4434), .CLK(n5042), .Q(
        n8349) );
  SDFFX1 DFF_1350_Q_reg ( .D(n194), .SI(n8349), .SE(n4434), .CLK(n5042), .Q(
        n8348) );
  SDFFX1 DFF_1351_Q_reg ( .D(n195), .SI(n8348), .SE(n4434), .CLK(n5042), .Q(
        n8347) );
  SDFFX1 DFF_1352_Q_reg ( .D(n196), .SI(n8347), .SE(n4434), .CLK(n5042), .Q(
        n8346) );
  SDFFX1 DFF_1353_Q_reg ( .D(n197), .SI(n8346), .SE(n4435), .CLK(n5042), .Q(
        test_so78) );
  SDFFX1 DFF_1354_Q_reg ( .D(n198), .SI(test_si79), .SE(n4435), .CLK(n5042), 
        .Q(n8343) );
  SDFFX1 DFF_1355_Q_reg ( .D(n199), .SI(n8343), .SE(n4435), .CLK(n5042), .Q(
        n8342) );
  SDFFX1 DFF_1356_Q_reg ( .D(n200), .SI(n8342), .SE(n4435), .CLK(n5042), .Q(
        n8341) );
  SDFFX1 DFF_1357_Q_reg ( .D(n201), .SI(n8341), .SE(n4435), .CLK(n5042), .Q(
        n8340) );
  SDFFX1 DFF_1358_Q_reg ( .D(n202), .SI(n8340), .SE(n4435), .CLK(n5041), .Q(
        n8339) );
  SDFFX1 DFF_1359_Q_reg ( .D(n203), .SI(n8339), .SE(n4436), .CLK(n5041), .Q(
        n8338) );
  SDFFX1 DFF_1360_Q_reg ( .D(n204), .SI(n8338), .SE(n4436), .CLK(n5041), .Q(
        n8337) );
  SDFFX1 DFF_1361_Q_reg ( .D(n205), .SI(n8337), .SE(n4436), .CLK(n5041), .Q(
        n8336) );
  SDFFX1 DFF_1362_Q_reg ( .D(n206), .SI(n8336), .SE(n4436), .CLK(n5041), .Q(
        n8335) );
  SDFFX1 DFF_1363_Q_reg ( .D(n207), .SI(n8335), .SE(n4436), .CLK(n5041), .Q(
        n8334) );
  SDFFX1 DFF_1364_Q_reg ( .D(n208), .SI(n8334), .SE(n4436), .CLK(n5041), .Q(
        n8333) );
  SDFFX1 DFF_1365_Q_reg ( .D(n209), .SI(n8333), .SE(n4437), .CLK(n5041), .Q(
        n8332) );
  SDFFX1 DFF_1366_Q_reg ( .D(n210), .SI(n8332), .SE(n4437), .CLK(n5041), .Q(
        n8331) );
  SDFFX1 DFF_1367_Q_reg ( .D(n211), .SI(n8331), .SE(n4437), .CLK(n5041), .Q(
        n8330) );
  SDFFX1 DFF_1368_Q_reg ( .D(n212), .SI(n8330), .SE(n4437), .CLK(n5041), .Q(
        n8329) );
  SDFFX1 DFF_1369_Q_reg ( .D(n213), .SI(n8329), .SE(n4437), .CLK(n5041), .Q(
        n8328) );
  SDFFX1 DFF_1370_Q_reg ( .D(n214), .SI(n8328), .SE(n4437), .CLK(n5040), .Q(
        test_so79) );
  SDFFX1 DFF_1371_Q_reg ( .D(n215), .SI(test_si80), .SE(n4438), .CLK(n5040), 
        .Q(n8325) );
  SDFFX1 DFF_1372_Q_reg ( .D(n216), .SI(n8325), .SE(n4438), .CLK(n5040), .Q(
        n8324) );
  SDFFX1 DFF_1373_Q_reg ( .D(n217), .SI(n8324), .SE(n4438), .CLK(n5040), .Q(
        n8323) );
  SDFFX1 DFF_1374_Q_reg ( .D(n218), .SI(n8323), .SE(n4438), .CLK(n5040), .Q(
        n8322) );
  SDFFX1 DFF_1375_Q_reg ( .D(WX9597), .SI(n8322), .SE(n4438), .CLK(n5040), .Q(
        n8321) );
  SDFFX1 DFF_1376_Q_reg ( .D(WX9695), .SI(n8321), .SE(n4433), .CLK(n5043), .Q(
        n8320), .QN(n8838) );
  SDFFX1 DFF_1377_Q_reg ( .D(WX9697), .SI(n8320), .SE(n4433), .CLK(n5043), .Q(
        n8319), .QN(n8837) );
  SDFFX1 DFF_1378_Q_reg ( .D(WX9699), .SI(n8319), .SE(n4432), .CLK(n5043), .Q(
        n8318), .QN(n8836) );
  SDFFX1 DFF_1379_Q_reg ( .D(WX9701), .SI(n8318), .SE(n4432), .CLK(n5043), .Q(
        n8317), .QN(n8835) );
  SDFFX1 DFF_1380_Q_reg ( .D(WX9703), .SI(n8317), .SE(n4432), .CLK(n5043), .Q(
        n8316), .QN(n8834) );
  SDFFX1 DFF_1381_Q_reg ( .D(WX9705), .SI(n8316), .SE(n4431), .CLK(n5044), .Q(
        n8315), .QN(n8833) );
  SDFFX1 DFF_1382_Q_reg ( .D(WX9707), .SI(n8315), .SE(n4431), .CLK(n5044), .Q(
        n8314), .QN(n8832) );
  SDFFX1 DFF_1383_Q_reg ( .D(WX9709), .SI(n8314), .SE(n4431), .CLK(n5044), .Q(
        n8313), .QN(n8831) );
  SDFFX1 DFF_1384_Q_reg ( .D(WX9711), .SI(n8313), .SE(n4430), .CLK(n5044), .Q(
        n8312), .QN(n8830) );
  SDFFX1 DFF_1385_Q_reg ( .D(WX9713), .SI(n8312), .SE(n4430), .CLK(n5044), .Q(
        n8311), .QN(n8829) );
  SDFFX1 DFF_1386_Q_reg ( .D(WX9715), .SI(n8311), .SE(n4430), .CLK(n5044), .Q(
        n8310), .QN(n8828) );
  SDFFX1 DFF_1387_Q_reg ( .D(WX9717), .SI(n8310), .SE(n4377), .CLK(n5071), .Q(
        test_so80) );
  SDFFX1 DFF_1388_Q_reg ( .D(WX9719), .SI(test_si81), .SE(n4429), .CLK(n5045), 
        .Q(n8307), .QN(n8827) );
  SDFFX1 DFF_1389_Q_reg ( .D(WX9721), .SI(n8307), .SE(n4429), .CLK(n5045), .Q(
        n8306), .QN(n8824) );
  SDFFX1 DFF_1390_Q_reg ( .D(WX9723), .SI(n8306), .SE(n4378), .CLK(n5071), .Q(
        n8305), .QN(n8823) );
  SDFFX1 DFF_1391_Q_reg ( .D(WX9725), .SI(n8305), .SE(n4428), .CLK(n5045), .Q(
        n8304), .QN(n8820) );
  SDFFX1 DFF_1392_Q_reg ( .D(WX9727), .SI(n8304), .SE(n4427), .CLK(n5045), .Q(
        WX9728) );
  SDFFX1 DFF_1393_Q_reg ( .D(WX9729), .SI(WX9728), .SE(n4427), .CLK(n5046), 
        .Q(WX9730) );
  SDFFX1 DFF_1394_Q_reg ( .D(WX9731), .SI(WX9730), .SE(n4427), .CLK(n5046), 
        .Q(WX9732) );
  SDFFX1 DFF_1395_Q_reg ( .D(WX9733), .SI(WX9732), .SE(n4426), .CLK(n5046), 
        .Q(WX9734) );
  SDFFX1 DFF_1396_Q_reg ( .D(WX9735), .SI(WX9734), .SE(n4488), .CLK(n5015), 
        .Q(WX9736) );
  SDFFX1 DFF_1397_Q_reg ( .D(WX9737), .SI(WX9736), .SE(n4488), .CLK(n5015), 
        .Q(WX9738) );
  SDFFX1 DFF_1398_Q_reg ( .D(WX9739), .SI(WX9738), .SE(n4488), .CLK(n5015), 
        .Q(WX9740) );
  SDFFX1 DFF_1399_Q_reg ( .D(WX9741), .SI(WX9740), .SE(n4488), .CLK(n5015), 
        .Q(WX9742) );
  SDFFX1 DFF_1400_Q_reg ( .D(WX9743), .SI(WX9742), .SE(n4488), .CLK(n5015), 
        .Q(WX9744) );
  SDFFX1 DFF_1401_Q_reg ( .D(WX9745), .SI(WX9744), .SE(n4488), .CLK(n5015), 
        .Q(WX9746) );
  SDFFX1 DFF_1402_Q_reg ( .D(WX9747), .SI(WX9746), .SE(n4487), .CLK(n5015), 
        .Q(WX9748) );
  SDFFX1 DFF_1403_Q_reg ( .D(WX9749), .SI(WX9748), .SE(n4487), .CLK(n5016), 
        .Q(WX9750) );
  SDFFX1 DFF_1404_Q_reg ( .D(WX9751), .SI(WX9750), .SE(n4487), .CLK(n5016), 
        .Q(test_so81) );
  SDFFX1 DFF_1405_Q_reg ( .D(WX9753), .SI(test_si82), .SE(n4420), .CLK(n5049), 
        .Q(WX9754) );
  SDFFX1 DFF_1406_Q_reg ( .D(WX9755), .SI(WX9754), .SE(n4420), .CLK(n5049), 
        .Q(WX9756) );
  SDFFX1 DFF_1407_Q_reg ( .D(WX9757), .SI(WX9756), .SE(n4420), .CLK(n5049), 
        .Q(WX9758) );
  SDFFX1 DFF_1408_Q_reg ( .D(WX9759), .SI(WX9758), .SE(n4433), .CLK(n5043), 
        .Q(WX9760) );
  SDFFX1 DFF_1409_Q_reg ( .D(WX9761), .SI(WX9760), .SE(n4433), .CLK(n5043), 
        .Q(WX9762), .QN(n3615) );
  SDFFX1 DFF_1410_Q_reg ( .D(WX9763), .SI(WX9762), .SE(n4432), .CLK(n5043), 
        .Q(WX9764), .QN(n3614) );
  SDFFX1 DFF_1411_Q_reg ( .D(WX9765), .SI(WX9764), .SE(n4432), .CLK(n5043), 
        .Q(WX9766), .QN(n3613) );
  SDFFX1 DFF_1412_Q_reg ( .D(WX9767), .SI(WX9766), .SE(n4432), .CLK(n5043), 
        .Q(WX9768), .QN(n3612) );
  SDFFX1 DFF_1413_Q_reg ( .D(WX9769), .SI(WX9768), .SE(n4431), .CLK(n5043), 
        .Q(WX9770), .QN(n3611) );
  SDFFX1 DFF_1414_Q_reg ( .D(WX9771), .SI(WX9770), .SE(n4431), .CLK(n5044), 
        .Q(WX9772), .QN(n3610) );
  SDFFX1 DFF_1415_Q_reg ( .D(WX9773), .SI(WX9772), .SE(n4431), .CLK(n5044), 
        .Q(WX9774), .QN(n3609) );
  SDFFX1 DFF_1416_Q_reg ( .D(WX9775), .SI(WX9774), .SE(n4430), .CLK(n5044), 
        .Q(WX9776), .QN(n3608) );
  SDFFX1 DFF_1417_Q_reg ( .D(WX9777), .SI(WX9776), .SE(n4430), .CLK(n5044), 
        .Q(WX9778), .QN(n3607) );
  SDFFX1 DFF_1418_Q_reg ( .D(WX9779), .SI(WX9778), .SE(n4430), .CLK(n5044), 
        .Q(WX9780), .QN(n3606) );
  SDFFX1 DFF_1419_Q_reg ( .D(WX9781), .SI(WX9780), .SE(n4429), .CLK(n5044), 
        .Q(WX9782) );
  SDFFX1 DFF_1420_Q_reg ( .D(WX9783), .SI(WX9782), .SE(n4429), .CLK(n5045), 
        .Q(WX9784), .QN(n3604) );
  SDFFX1 DFF_1421_Q_reg ( .D(WX9785), .SI(WX9784), .SE(n4429), .CLK(n5045), 
        .Q(test_so82), .QN(n8825) );
  SDFFX1 DFF_1422_Q_reg ( .D(WX9787), .SI(test_si83), .SE(n4378), .CLK(n5071), 
        .Q(WX9788), .QN(n3603) );
  SDFFX1 DFF_1423_Q_reg ( .D(WX9789), .SI(WX9788), .SE(n4428), .CLK(n5045), 
        .Q(WX9790), .QN(n8822) );
  SDFFX1 DFF_1424_Q_reg ( .D(WX9791), .SI(WX9790), .SE(n4428), .CLK(n5045), 
        .Q(WX9792), .QN(n8819) );
  SDFFX1 DFF_1425_Q_reg ( .D(WX9793), .SI(WX9792), .SE(n4427), .CLK(n5046), 
        .Q(WX9794), .QN(n8818) );
  SDFFX1 DFF_1426_Q_reg ( .D(WX9795), .SI(WX9794), .SE(n4427), .CLK(n5046), 
        .Q(WX9796), .QN(n8817) );
  SDFFX1 DFF_1427_Q_reg ( .D(WX9797), .SI(WX9796), .SE(n4426), .CLK(n5046), 
        .Q(WX9798), .QN(n8816) );
  SDFFX1 DFF_1428_Q_reg ( .D(WX9799), .SI(WX9798), .SE(n4425), .CLK(n5046), 
        .Q(WX9800), .QN(n8815) );
  SDFFX1 DFF_1429_Q_reg ( .D(WX9801), .SI(WX9800), .SE(n4425), .CLK(n5047), 
        .Q(WX9802), .QN(n8814) );
  SDFFX1 DFF_1430_Q_reg ( .D(WX9803), .SI(WX9802), .SE(n4424), .CLK(n5047), 
        .Q(WX9804), .QN(n8813) );
  SDFFX1 DFF_1431_Q_reg ( .D(WX9805), .SI(WX9804), .SE(n4424), .CLK(n5047), 
        .Q(WX9806), .QN(n8812) );
  SDFFX1 DFF_1432_Q_reg ( .D(WX9807), .SI(WX9806), .SE(n4423), .CLK(n5047), 
        .Q(WX9808), .QN(n8811) );
  SDFFX1 DFF_1433_Q_reg ( .D(WX9809), .SI(WX9808), .SE(n4423), .CLK(n5048), 
        .Q(WX9810), .QN(n8810) );
  SDFFX1 DFF_1434_Q_reg ( .D(WX9811), .SI(WX9810), .SE(n4422), .CLK(n5048), 
        .Q(WX9812), .QN(n8809) );
  SDFFX1 DFF_1435_Q_reg ( .D(WX9813), .SI(WX9812), .SE(n4422), .CLK(n5048), 
        .Q(WX9814), .QN(n8808) );
  SDFFX1 DFF_1436_Q_reg ( .D(WX9815), .SI(WX9814), .SE(n4421), .CLK(n5048), 
        .Q(WX9816), .QN(n8807) );
  SDFFX1 DFF_1437_Q_reg ( .D(WX9817), .SI(WX9816), .SE(n4421), .CLK(n5049), 
        .Q(WX9818), .QN(n8806) );
  SDFFX1 DFF_1438_Q_reg ( .D(WX9819), .SI(WX9818), .SE(n4420), .CLK(n5049), 
        .Q(test_so83) );
  SDFFX1 DFF_1439_Q_reg ( .D(WX9821), .SI(test_si84), .SE(n4419), .CLK(n5049), 
        .Q(WX9822), .QN(n8804) );
  SDFFX1 DFF_1440_Q_reg ( .D(WX9823), .SI(WX9822), .SE(n4419), .CLK(n5050), 
        .Q(WX9824), .QN(n3583) );
  SDFFX1 DFF_1441_Q_reg ( .D(WX9825), .SI(WX9824), .SE(n4419), .CLK(n5050), 
        .Q(WX9826) );
  SDFFX1 DFF_1442_Q_reg ( .D(WX9827), .SI(WX9826), .SE(n4418), .CLK(n5050), 
        .Q(WX9828) );
  SDFFX1 DFF_1443_Q_reg ( .D(WX9829), .SI(WX9828), .SE(n4418), .CLK(n5050), 
        .Q(WX9830) );
  SDFFX1 DFF_1444_Q_reg ( .D(WX9831), .SI(WX9830), .SE(n4418), .CLK(n5050), 
        .Q(WX9832) );
  SDFFX1 DFF_1445_Q_reg ( .D(WX9833), .SI(WX9832), .SE(n4417), .CLK(n5051), 
        .Q(WX9834) );
  SDFFX1 DFF_1446_Q_reg ( .D(WX9835), .SI(WX9834), .SE(n4417), .CLK(n5051), 
        .Q(WX9836) );
  SDFFX1 DFF_1447_Q_reg ( .D(WX9837), .SI(WX9836), .SE(n4417), .CLK(n5051), 
        .Q(WX9838) );
  SDFFX1 DFF_1448_Q_reg ( .D(WX9839), .SI(WX9838), .SE(n4416), .CLK(n5051), 
        .Q(WX9840) );
  SDFFX1 DFF_1449_Q_reg ( .D(WX9841), .SI(WX9840), .SE(n4416), .CLK(n5051), 
        .Q(WX9842) );
  SDFFX1 DFF_1450_Q_reg ( .D(WX9843), .SI(WX9842), .SE(n4416), .CLK(n5051), 
        .Q(WX9844) );
  SDFFX1 DFF_1451_Q_reg ( .D(WX9845), .SI(WX9844), .SE(n4415), .CLK(n5052), 
        .Q(WX9846), .QN(n3605) );
  SDFFX1 DFF_1452_Q_reg ( .D(WX9847), .SI(WX9846), .SE(n4415), .CLK(n5052), 
        .Q(WX9848) );
  SDFFX1 DFF_1453_Q_reg ( .D(WX9849), .SI(WX9848), .SE(n4429), .CLK(n5045), 
        .Q(WX9850), .QN(n8826) );
  SDFFX1 DFF_1454_Q_reg ( .D(WX9851), .SI(WX9850), .SE(n4428), .CLK(n5045), 
        .Q(WX9852) );
  SDFFX1 DFF_1455_Q_reg ( .D(WX9853), .SI(WX9852), .SE(n4428), .CLK(n5045), 
        .Q(test_so84), .QN(n8821) );
  SDFFX1 DFF_1456_Q_reg ( .D(WX9855), .SI(test_si85), .SE(n4428), .CLK(n5045), 
        .Q(WX9856), .QN(n3754) );
  SDFFX1 DFF_1457_Q_reg ( .D(WX9857), .SI(WX9856), .SE(n4427), .CLK(n5046), 
        .Q(WX9858), .QN(n3752) );
  SDFFX1 DFF_1458_Q_reg ( .D(WX9859), .SI(WX9858), .SE(n4426), .CLK(n5046), 
        .Q(WX9860), .QN(n3750) );
  SDFFX1 DFF_1459_Q_reg ( .D(WX9861), .SI(WX9860), .SE(n4426), .CLK(n5046), 
        .Q(WX9862), .QN(n3748) );
  SDFFX1 DFF_1460_Q_reg ( .D(WX9863), .SI(WX9862), .SE(n4425), .CLK(n5047), 
        .Q(WX9864), .QN(n3746) );
  SDFFX1 DFF_1461_Q_reg ( .D(WX9865), .SI(WX9864), .SE(n4425), .CLK(n5047), 
        .Q(WX9866), .QN(n3744) );
  SDFFX1 DFF_1462_Q_reg ( .D(WX9867), .SI(WX9866), .SE(n4424), .CLK(n5047), 
        .Q(WX9868), .QN(n3742) );
  SDFFX1 DFF_1463_Q_reg ( .D(WX9869), .SI(WX9868), .SE(n4424), .CLK(n5047), 
        .Q(WX9870), .QN(n3740) );
  SDFFX1 DFF_1464_Q_reg ( .D(WX9871), .SI(WX9870), .SE(n4423), .CLK(n5048), 
        .Q(WX9872), .QN(n3738) );
  SDFFX1 DFF_1465_Q_reg ( .D(WX9873), .SI(WX9872), .SE(n4423), .CLK(n5048), 
        .Q(WX9874), .QN(n3736) );
  SDFFX1 DFF_1466_Q_reg ( .D(WX9875), .SI(WX9874), .SE(n4422), .CLK(n5048), 
        .Q(WX9876), .QN(n3734) );
  SDFFX1 DFF_1467_Q_reg ( .D(WX9877), .SI(WX9876), .SE(n4422), .CLK(n5048), 
        .Q(WX9878), .QN(n3732) );
  SDFFX1 DFF_1468_Q_reg ( .D(WX9879), .SI(WX9878), .SE(n4421), .CLK(n5049), 
        .Q(WX9880) );
  SDFFX1 DFF_1469_Q_reg ( .D(WX9881), .SI(WX9880), .SE(n4421), .CLK(n5049), 
        .Q(WX9882), .QN(n3729) );
  SDFFX1 DFF_1470_Q_reg ( .D(WX9883), .SI(WX9882), .SE(n4420), .CLK(n5049), 
        .Q(WX9884), .QN(n8805) );
  SDFFX1 DFF_1471_Q_reg ( .D(WX9885), .SI(WX9884), .SE(n4419), .CLK(n5050), 
        .Q(WX9886), .QN(n3726) );
  SDFFX1 DFF_1472_Q_reg ( .D(WX9887), .SI(WX9886), .SE(n4419), .CLK(n5050), 
        .Q(test_so85) );
  SDFFX1 DFF_1473_Q_reg ( .D(WX9889), .SI(test_si86), .SE(n4418), .CLK(n5050), 
        .Q(WX9890), .QN(n3994) );
  SDFFX1 DFF_1474_Q_reg ( .D(WX9891), .SI(WX9890), .SE(n4418), .CLK(n5050), 
        .Q(WX9892), .QN(n3995) );
  SDFFX1 DFF_1475_Q_reg ( .D(WX9893), .SI(WX9892), .SE(n4418), .CLK(n5050), 
        .Q(WX9894), .QN(n3996) );
  SDFFX1 DFF_1476_Q_reg ( .D(WX9895), .SI(WX9894), .SE(n4417), .CLK(n5050), 
        .Q(WX9896), .QN(n3997) );
  SDFFX1 DFF_1477_Q_reg ( .D(WX9897), .SI(WX9896), .SE(n4417), .CLK(n5051), 
        .Q(WX9898), .QN(n3998) );
  SDFFX1 DFF_1478_Q_reg ( .D(WX9899), .SI(WX9898), .SE(n4417), .CLK(n5051), 
        .Q(WX9900), .QN(n3999) );
  SDFFX1 DFF_1479_Q_reg ( .D(WX9901), .SI(WX9900), .SE(n4416), .CLK(n5051), 
        .Q(WX9902), .QN(n4000) );
  SDFFX1 DFF_1480_Q_reg ( .D(WX9903), .SI(WX9902), .SE(n4416), .CLK(n5051), 
        .Q(WX9904), .QN(n4001) );
  SDFFX1 DFF_1481_Q_reg ( .D(WX9905), .SI(WX9904), .SE(n4416), .CLK(n5051), 
        .Q(WX9906), .QN(n4002) );
  SDFFX1 DFF_1482_Q_reg ( .D(WX9907), .SI(WX9906), .SE(n4415), .CLK(n5051), 
        .Q(WX9908), .QN(n4003) );
  SDFFX1 DFF_1483_Q_reg ( .D(WX9909), .SI(WX9908), .SE(n4415), .CLK(n5052), 
        .Q(WX9910), .QN(n4004) );
  SDFFX1 DFF_1484_Q_reg ( .D(WX9911), .SI(WX9910), .SE(n4415), .CLK(n5052), 
        .Q(WX9912), .QN(n4005) );
  SDFFX1 DFF_1485_Q_reg ( .D(WX9913), .SI(WX9912), .SE(n4415), .CLK(n5052), 
        .Q(WX9914), .QN(n4006) );
  SDFFX1 DFF_1486_Q_reg ( .D(WX9915), .SI(WX9914), .SE(n4414), .CLK(n5052), 
        .Q(WX9916), .QN(n4007) );
  SDFFX1 DFF_1487_Q_reg ( .D(WX9917), .SI(WX9916), .SE(n4414), .CLK(n5052), 
        .Q(WX9918), .QN(n3942) );
  SDFFX1 DFF_1488_Q_reg ( .D(WX9919), .SI(WX9918), .SE(n4414), .CLK(n5052), 
        .Q(WX9920), .QN(n4008) );
  SDFFX1 DFF_1489_Q_reg ( .D(WX9921), .SI(WX9920), .SE(n4414), .CLK(n5052), 
        .Q(test_so86) );
  SDFFX1 DFF_1490_Q_reg ( .D(WX9923), .SI(test_si87), .SE(n4426), .CLK(n5046), 
        .Q(WX9924), .QN(n4009) );
  SDFFX1 DFF_1491_Q_reg ( .D(WX9925), .SI(WX9924), .SE(n4426), .CLK(n5046), 
        .Q(WX9926), .QN(n4010) );
  SDFFX1 DFF_1492_Q_reg ( .D(WX9927), .SI(WX9926), .SE(n4425), .CLK(n5047), 
        .Q(WX9928), .QN(n3943) );
  SDFFX1 DFF_1493_Q_reg ( .D(WX9929), .SI(WX9928), .SE(n4425), .CLK(n5047), 
        .Q(WX9930), .QN(n4011) );
  SDFFX1 DFF_1494_Q_reg ( .D(WX9931), .SI(WX9930), .SE(n4424), .CLK(n5047), 
        .Q(WX9932), .QN(n4012) );
  SDFFX1 DFF_1495_Q_reg ( .D(WX9933), .SI(WX9932), .SE(n4424), .CLK(n5047), 
        .Q(WX9934), .QN(n4013) );
  SDFFX1 DFF_1496_Q_reg ( .D(WX9935), .SI(WX9934), .SE(n4423), .CLK(n5048), 
        .Q(WX9936), .QN(n4014) );
  SDFFX1 DFF_1497_Q_reg ( .D(WX9937), .SI(WX9936), .SE(n4423), .CLK(n5048), 
        .Q(WX9938), .QN(n4015) );
  SDFFX1 DFF_1498_Q_reg ( .D(WX9939), .SI(WX9938), .SE(n4422), .CLK(n5048), 
        .Q(WX9940), .QN(n4016) );
  SDFFX1 DFF_1499_Q_reg ( .D(WX9941), .SI(WX9940), .SE(n4422), .CLK(n5048), 
        .Q(WX9942), .QN(n3944) );
  SDFFX1 DFF_1500_Q_reg ( .D(WX9943), .SI(WX9942), .SE(n4421), .CLK(n5049), 
        .Q(WX9944), .QN(n4017) );
  SDFFX1 DFF_1501_Q_reg ( .D(WX9945), .SI(WX9944), .SE(n4421), .CLK(n5049), 
        .Q(WX9946), .QN(n4018) );
  SDFFX1 DFF_1502_Q_reg ( .D(WX9947), .SI(WX9946), .SE(n4420), .CLK(n5049), 
        .Q(WX9948), .QN(n4019) );
  SDFFX1 DFF_1503_Q_reg ( .D(WX9949), .SI(WX9948), .SE(n4419), .CLK(n5050), 
        .Q(WX9950), .QN(n3961) );
  SDFFX1 DFF_1504_Q_reg ( .D(WX10315), .SI(WX9950), .SE(n4381), .CLK(n5069), 
        .Q(CRC_OUT_2_0), .QN(DFF_1504_n1) );
  SDFFX1 DFF_1505_Q_reg ( .D(WX10317), .SI(CRC_OUT_2_0), .SE(n4381), .CLK(
        n5069), .Q(CRC_OUT_2_1), .QN(DFF_1505_n1) );
  SDFFX1 DFF_1506_Q_reg ( .D(WX10319), .SI(CRC_OUT_2_1), .SE(n4381), .CLK(
        n5069), .Q(test_so87) );
  SDFFX1 DFF_1507_Q_reg ( .D(WX10321), .SI(test_si88), .SE(n4380), .CLK(n5070), 
        .Q(CRC_OUT_2_3), .QN(DFF_1507_n1) );
  SDFFX1 DFF_1508_Q_reg ( .D(WX10323), .SI(CRC_OUT_2_3), .SE(n4380), .CLK(
        n5070), .Q(CRC_OUT_2_4), .QN(DFF_1508_n1) );
  SDFFX1 DFF_1509_Q_reg ( .D(WX10325), .SI(CRC_OUT_2_4), .SE(n4380), .CLK(
        n5070), .Q(CRC_OUT_2_5), .QN(DFF_1509_n1) );
  SDFFX1 DFF_1510_Q_reg ( .D(WX10327), .SI(CRC_OUT_2_5), .SE(n4380), .CLK(
        n5070), .Q(CRC_OUT_2_6), .QN(DFF_1510_n1) );
  SDFFX1 DFF_1511_Q_reg ( .D(WX10329), .SI(CRC_OUT_2_6), .SE(n4380), .CLK(
        n5070), .Q(CRC_OUT_2_7), .QN(DFF_1511_n1) );
  SDFFX1 DFF_1512_Q_reg ( .D(WX10331), .SI(CRC_OUT_2_7), .SE(n4380), .CLK(
        n5070), .Q(CRC_OUT_2_8), .QN(DFF_1512_n1) );
  SDFFX1 DFF_1513_Q_reg ( .D(WX10333), .SI(CRC_OUT_2_8), .SE(n4379), .CLK(
        n5070), .Q(CRC_OUT_2_9), .QN(DFF_1513_n1) );
  SDFFX1 DFF_1514_Q_reg ( .D(WX10335), .SI(CRC_OUT_2_9), .SE(n4379), .CLK(
        n5070), .Q(CRC_OUT_2_10), .QN(DFF_1514_n1) );
  SDFFX1 DFF_1515_Q_reg ( .D(WX10337), .SI(CRC_OUT_2_10), .SE(n4379), .CLK(
        n5070), .Q(CRC_OUT_2_11), .QN(DFF_1515_n1) );
  SDFFX1 DFF_1516_Q_reg ( .D(WX10339), .SI(CRC_OUT_2_11), .SE(n4379), .CLK(
        n5070), .Q(CRC_OUT_2_12), .QN(DFF_1516_n1) );
  SDFFX1 DFF_1517_Q_reg ( .D(WX10341), .SI(CRC_OUT_2_12), .SE(n4379), .CLK(
        n5070), .Q(CRC_OUT_2_13), .QN(DFF_1517_n1) );
  SDFFX1 DFF_1518_Q_reg ( .D(WX10343), .SI(CRC_OUT_2_13), .SE(n4379), .CLK(
        n5070), .Q(CRC_OUT_2_14), .QN(DFF_1518_n1) );
  SDFFX1 DFF_1519_Q_reg ( .D(WX10345), .SI(CRC_OUT_2_14), .SE(n4378), .CLK(
        n5071), .Q(CRC_OUT_2_15), .QN(DFF_1519_n1) );
  SDFFX1 DFF_1520_Q_reg ( .D(WX10347), .SI(CRC_OUT_2_15), .SE(n4378), .CLK(
        n5071), .Q(CRC_OUT_2_16), .QN(DFF_1520_n1) );
  SDFFX1 DFF_1521_Q_reg ( .D(WX10349), .SI(CRC_OUT_2_16), .SE(n4378), .CLK(
        n5071), .Q(CRC_OUT_2_17), .QN(DFF_1521_n1) );
  SDFFX1 DFF_1522_Q_reg ( .D(WX10351), .SI(CRC_OUT_2_17), .SE(n4378), .CLK(
        n5071), .Q(CRC_OUT_2_18), .QN(DFF_1522_n1) );
  SDFFX1 DFF_1523_Q_reg ( .D(WX10353), .SI(CRC_OUT_2_18), .SE(n4414), .CLK(
        n5052), .Q(test_so88) );
  SDFFX1 DFF_1524_Q_reg ( .D(WX10355), .SI(test_si89), .SE(n4414), .CLK(n5052), 
        .Q(CRC_OUT_2_20), .QN(DFF_1524_n1) );
  SDFFX1 DFF_1525_Q_reg ( .D(WX10357), .SI(CRC_OUT_2_20), .SE(n4413), .CLK(
        n5052), .Q(CRC_OUT_2_21), .QN(DFF_1525_n1) );
  SDFFX1 DFF_1526_Q_reg ( .D(WX10359), .SI(CRC_OUT_2_21), .SE(n4413), .CLK(
        n5053), .Q(CRC_OUT_2_22), .QN(DFF_1526_n1) );
  SDFFX1 DFF_1527_Q_reg ( .D(WX10361), .SI(CRC_OUT_2_22), .SE(n4413), .CLK(
        n5053), .Q(CRC_OUT_2_23), .QN(DFF_1527_n1) );
  SDFFX1 DFF_1528_Q_reg ( .D(WX10363), .SI(CRC_OUT_2_23), .SE(n4413), .CLK(
        n5053), .Q(CRC_OUT_2_24), .QN(DFF_1528_n1) );
  SDFFX1 DFF_1529_Q_reg ( .D(WX10365), .SI(CRC_OUT_2_24), .SE(n4413), .CLK(
        n5053), .Q(CRC_OUT_2_25), .QN(DFF_1529_n1) );
  SDFFX1 DFF_1530_Q_reg ( .D(WX10367), .SI(CRC_OUT_2_25), .SE(n4413), .CLK(
        n5053), .Q(CRC_OUT_2_26), .QN(DFF_1530_n1) );
  SDFFX1 DFF_1531_Q_reg ( .D(WX10369), .SI(CRC_OUT_2_26), .SE(n4412), .CLK(
        n5053), .Q(CRC_OUT_2_27), .QN(DFF_1531_n1) );
  SDFFX1 DFF_1532_Q_reg ( .D(WX10371), .SI(CRC_OUT_2_27), .SE(n4412), .CLK(
        n5053), .Q(CRC_OUT_2_28), .QN(DFF_1532_n1) );
  SDFFX1 DFF_1533_Q_reg ( .D(WX10373), .SI(CRC_OUT_2_28), .SE(n4412), .CLK(
        n5053), .Q(CRC_OUT_2_29), .QN(DFF_1533_n1) );
  SDFFX1 DFF_1534_Q_reg ( .D(WX10375), .SI(CRC_OUT_2_29), .SE(n4412), .CLK(
        n5053), .Q(CRC_OUT_2_30), .QN(DFF_1534_n1) );
  SDFFX1 DFF_1535_Q_reg ( .D(WX10377), .SI(CRC_OUT_2_30), .SE(n4412), .CLK(
        n5053), .Q(CRC_OUT_2_31), .QN(DFF_1535_n1) );
  SDFFX1 DFF_1536_Q_reg ( .D(WX10828), .SI(CRC_OUT_2_31), .SE(n4412), .CLK(
        n5053), .Q(WX10829), .QN(n3931) );
  SDFFX1 DFF_1537_Q_reg ( .D(WX10830), .SI(WX10829), .SE(n4406), .CLK(n5056), 
        .Q(n8295) );
  SDFFX1 DFF_1538_Q_reg ( .D(WX10832), .SI(n8295), .SE(n4407), .CLK(n5056), 
        .Q(n8294) );
  SDFFX1 DFF_1539_Q_reg ( .D(WX10834), .SI(n8294), .SE(n4407), .CLK(n5056), 
        .Q(n8293) );
  SDFFX1 DFF_1540_Q_reg ( .D(WX10836), .SI(n8293), .SE(n4407), .CLK(n5056), 
        .Q(test_so89) );
  SDFFX1 DFF_1541_Q_reg ( .D(WX10838), .SI(test_si90), .SE(n4407), .CLK(n5056), 
        .Q(n8290) );
  SDFFX1 DFF_1542_Q_reg ( .D(WX10840), .SI(n8290), .SE(n4407), .CLK(n5056), 
        .Q(n8289) );
  SDFFX1 DFF_1543_Q_reg ( .D(WX10842), .SI(n8289), .SE(n4407), .CLK(n5055), 
        .Q(n8288) );
  SDFFX1 DFF_1544_Q_reg ( .D(WX10844), .SI(n8288), .SE(n4408), .CLK(n5055), 
        .Q(n8287) );
  SDFFX1 DFF_1545_Q_reg ( .D(WX10846), .SI(n8287), .SE(n4408), .CLK(n5055), 
        .Q(n8286) );
  SDFFX1 DFF_1546_Q_reg ( .D(WX10848), .SI(n8286), .SE(n4408), .CLK(n5055), 
        .Q(n8285) );
  SDFFX1 DFF_1547_Q_reg ( .D(WX10850), .SI(n8285), .SE(n4408), .CLK(n5055), 
        .Q(n8284) );
  SDFFX1 DFF_1548_Q_reg ( .D(WX10852), .SI(n8284), .SE(n4408), .CLK(n5055), 
        .Q(n8283) );
  SDFFX1 DFF_1549_Q_reg ( .D(WX10854), .SI(n8283), .SE(n4408), .CLK(n5055), 
        .Q(n8282) );
  SDFFX1 DFF_1550_Q_reg ( .D(WX10856), .SI(n8282), .SE(n4409), .CLK(n5055), 
        .Q(n8281) );
  SDFFX1 DFF_1551_Q_reg ( .D(WX10858), .SI(n8281), .SE(n4409), .CLK(n5055), 
        .Q(n8280) );
  SDFFX1 DFF_1552_Q_reg ( .D(WX10860), .SI(n8280), .SE(n4409), .CLK(n5055), 
        .Q(n8279) );
  SDFFX1 DFF_1553_Q_reg ( .D(WX10862), .SI(n8279), .SE(n4409), .CLK(n5055), 
        .Q(n8278) );
  SDFFX1 DFF_1554_Q_reg ( .D(WX10864), .SI(n8278), .SE(n4409), .CLK(n5055), 
        .Q(n8277) );
  SDFFX1 DFF_1555_Q_reg ( .D(WX10866), .SI(n8277), .SE(n4409), .CLK(n5054), 
        .Q(n8276) );
  SDFFX1 DFF_1556_Q_reg ( .D(WX10868), .SI(n8276), .SE(n4410), .CLK(n5054), 
        .Q(n8275) );
  SDFFX1 DFF_1557_Q_reg ( .D(WX10870), .SI(n8275), .SE(n4410), .CLK(n5054), 
        .Q(test_so90) );
  SDFFX1 DFF_1558_Q_reg ( .D(WX10872), .SI(test_si91), .SE(n4410), .CLK(n5054), 
        .Q(n8272) );
  SDFFX1 DFF_1559_Q_reg ( .D(WX10874), .SI(n8272), .SE(n4410), .CLK(n5054), 
        .Q(n8271) );
  SDFFX1 DFF_1560_Q_reg ( .D(WX10876), .SI(n8271), .SE(n4410), .CLK(n5054), 
        .Q(n8270) );
  SDFFX1 DFF_1561_Q_reg ( .D(WX10878), .SI(n8270), .SE(n4410), .CLK(n5054), 
        .Q(n8269) );
  SDFFX1 DFF_1562_Q_reg ( .D(WX10880), .SI(n8269), .SE(n4411), .CLK(n5054), 
        .Q(n8268) );
  SDFFX1 DFF_1563_Q_reg ( .D(WX10882), .SI(n8268), .SE(n4411), .CLK(n5054), 
        .Q(n8267) );
  SDFFX1 DFF_1564_Q_reg ( .D(WX10884), .SI(n8267), .SE(n4411), .CLK(n5054), 
        .Q(n8266) );
  SDFFX1 DFF_1565_Q_reg ( .D(WX10886), .SI(n8266), .SE(n4411), .CLK(n5054), 
        .Q(n8265) );
  SDFFX1 DFF_1566_Q_reg ( .D(WX10888), .SI(n8265), .SE(n4411), .CLK(n5054), 
        .Q(n8264) );
  SDFFX1 DFF_1567_Q_reg ( .D(WX10890), .SI(n8264), .SE(n4411), .CLK(n5053), 
        .Q(n8263) );
  SDFFX1 DFF_1568_Q_reg ( .D(WX10988), .SI(n8263), .SE(n4406), .CLK(n5056), 
        .Q(n8262), .QN(n9080) );
  SDFFX1 DFF_1569_Q_reg ( .D(WX10990), .SI(n8262), .SE(n4406), .CLK(n5056), 
        .Q(n8261), .QN(n9079) );
  SDFFX1 DFF_1570_Q_reg ( .D(WX10992), .SI(n8261), .SE(n4406), .CLK(n5056), 
        .Q(n8260), .QN(n9078) );
  SDFFX1 DFF_1571_Q_reg ( .D(WX10994), .SI(n8260), .SE(n4405), .CLK(n5057), 
        .Q(n8259), .QN(n9077) );
  SDFFX1 DFF_1572_Q_reg ( .D(WX10996), .SI(n8259), .SE(n4405), .CLK(n5057), 
        .Q(n8258), .QN(n9076) );
  SDFFX1 DFF_1573_Q_reg ( .D(WX10998), .SI(n8258), .SE(n4404), .CLK(n5057), 
        .Q(n8257), .QN(n9075) );
  SDFFX1 DFF_1574_Q_reg ( .D(WX11000), .SI(n8257), .SE(n4404), .CLK(n5057), 
        .Q(test_so91) );
  SDFFX1 DFF_1575_Q_reg ( .D(WX11002), .SI(test_si92), .SE(n4404), .CLK(n5057), 
        .Q(n8254), .QN(n9074) );
  SDFFX1 DFF_1576_Q_reg ( .D(WX11004), .SI(n8254), .SE(n4404), .CLK(n5057), 
        .Q(n8253), .QN(n9071) );
  SDFFX1 DFF_1577_Q_reg ( .D(WX11006), .SI(n8253), .SE(n4381), .CLK(n5069), 
        .Q(n8252), .QN(n9070) );
  SDFFX1 DFF_1578_Q_reg ( .D(WX11008), .SI(n8252), .SE(n4403), .CLK(n5058), 
        .Q(n8251), .QN(n9067) );
  SDFFX1 DFF_1579_Q_reg ( .D(WX11010), .SI(n8251), .SE(n4402), .CLK(n5058), 
        .Q(n8250), .QN(n9066) );
  SDFFX1 DFF_1580_Q_reg ( .D(WX11012), .SI(n8250), .SE(n4402), .CLK(n5058), 
        .Q(n8249), .QN(n9065) );
  SDFFX1 DFF_1581_Q_reg ( .D(WX11014), .SI(n8249), .SE(n4401), .CLK(n5059), 
        .Q(n8248), .QN(n9064) );
  SDFFX1 DFF_1582_Q_reg ( .D(WX11016), .SI(n8248), .SE(n4401), .CLK(n5059), 
        .Q(n8247), .QN(n9063) );
  SDFFX1 DFF_1583_Q_reg ( .D(WX11018), .SI(n8247), .SE(n4400), .CLK(n5059), 
        .Q(n8246), .QN(n9062) );
  SDFFX1 DFF_1584_Q_reg ( .D(WX11020), .SI(n8246), .SE(n4399), .CLK(n5059), 
        .Q(WX11021) );
  SDFFX1 DFF_1585_Q_reg ( .D(WX11022), .SI(WX11021), .SE(n4399), .CLK(n5060), 
        .Q(WX11023) );
  SDFFX1 DFF_1586_Q_reg ( .D(WX11024), .SI(WX11023), .SE(n4398), .CLK(n5060), 
        .Q(WX11025) );
  SDFFX1 DFF_1587_Q_reg ( .D(WX11026), .SI(WX11025), .SE(n4397), .CLK(n5060), 
        .Q(WX11027) );
  SDFFX1 DFF_1588_Q_reg ( .D(WX11028), .SI(WX11027), .SE(n4397), .CLK(n5061), 
        .Q(WX11029) );
  SDFFX1 DFF_1589_Q_reg ( .D(WX11030), .SI(WX11029), .SE(n4396), .CLK(n5061), 
        .Q(WX11031) );
  SDFFX1 DFF_1590_Q_reg ( .D(WX11032), .SI(WX11031), .SE(n4396), .CLK(n5061), 
        .Q(WX11033) );
  SDFFX1 DFF_1591_Q_reg ( .D(WX11034), .SI(WX11033), .SE(n4395), .CLK(n5062), 
        .Q(test_so92) );
  SDFFX1 DFF_1592_Q_reg ( .D(WX11036), .SI(test_si93), .SE(n4394), .CLK(n5062), 
        .Q(WX11037) );
  SDFFX1 DFF_1593_Q_reg ( .D(WX11038), .SI(WX11037), .SE(n4394), .CLK(n5062), 
        .Q(WX11039) );
  SDFFX1 DFF_1594_Q_reg ( .D(WX11040), .SI(WX11039), .SE(n4394), .CLK(n5063), 
        .Q(WX11041) );
  SDFFX1 DFF_1595_Q_reg ( .D(WX11042), .SI(WX11041), .SE(n4393), .CLK(n5063), 
        .Q(WX11043) );
  SDFFX1 DFF_1596_Q_reg ( .D(WX11044), .SI(WX11043), .SE(n4393), .CLK(n5063), 
        .Q(WX11045) );
  SDFFX1 DFF_1597_Q_reg ( .D(WX11046), .SI(WX11045), .SE(n4392), .CLK(n5064), 
        .Q(WX11047) );
  SDFFX1 DFF_1598_Q_reg ( .D(WX11048), .SI(WX11047), .SE(n4391), .CLK(n5064), 
        .Q(WX11049) );
  SDFFX1 DFF_1599_Q_reg ( .D(WX11050), .SI(WX11049), .SE(n4391), .CLK(n5064), 
        .Q(WX11051) );
  SDFFX1 DFF_1600_Q_reg ( .D(WX11052), .SI(WX11051), .SE(n4406), .CLK(n5056), 
        .Q(WX11053), .QN(n3582) );
  SDFFX1 DFF_1601_Q_reg ( .D(WX11054), .SI(WX11053), .SE(n4406), .CLK(n5056), 
        .Q(WX11055), .QN(n3602) );
  SDFFX1 DFF_1602_Q_reg ( .D(WX11056), .SI(WX11055), .SE(n4405), .CLK(n5056), 
        .Q(WX11057), .QN(n3601) );
  SDFFX1 DFF_1603_Q_reg ( .D(WX11058), .SI(WX11057), .SE(n4405), .CLK(n5057), 
        .Q(WX11059), .QN(n3600) );
  SDFFX1 DFF_1604_Q_reg ( .D(WX11060), .SI(WX11059), .SE(n4405), .CLK(n5057), 
        .Q(WX11061), .QN(n3599) );
  SDFFX1 DFF_1605_Q_reg ( .D(WX11062), .SI(WX11061), .SE(n4405), .CLK(n5057), 
        .Q(WX11063), .QN(n3598) );
  SDFFX1 DFF_1606_Q_reg ( .D(WX11064), .SI(WX11063), .SE(n4404), .CLK(n5057), 
        .Q(WX11065) );
  SDFFX1 DFF_1607_Q_reg ( .D(WX11066), .SI(WX11065), .SE(n4404), .CLK(n5057), 
        .Q(WX11067), .QN(n3596) );
  SDFFX1 DFF_1608_Q_reg ( .D(WX11068), .SI(WX11067), .SE(n4403), .CLK(n5057), 
        .Q(test_so93), .QN(n9072) );
  SDFFX1 DFF_1609_Q_reg ( .D(WX11070), .SI(test_si94), .SE(n4381), .CLK(n5069), 
        .Q(WX11071), .QN(n3595) );
  SDFFX1 DFF_1610_Q_reg ( .D(WX11072), .SI(WX11071), .SE(n4403), .CLK(n5058), 
        .Q(WX11073), .QN(n9069) );
  SDFFX1 DFF_1611_Q_reg ( .D(WX11074), .SI(WX11073), .SE(n4402), .CLK(n5058), 
        .Q(WX11075), .QN(n3594) );
  SDFFX1 DFF_1612_Q_reg ( .D(WX11076), .SI(WX11075), .SE(n4402), .CLK(n5058), 
        .Q(WX11077) );
  SDFFX1 DFF_1613_Q_reg ( .D(WX11078), .SI(WX11077), .SE(n4401), .CLK(n5058), 
        .Q(WX11079), .QN(n3592) );
  SDFFX1 DFF_1614_Q_reg ( .D(WX11080), .SI(WX11079), .SE(n4401), .CLK(n5059), 
        .Q(WX11081), .QN(n3591) );
  SDFFX1 DFF_1615_Q_reg ( .D(WX11082), .SI(WX11081), .SE(n4400), .CLK(n5059), 
        .Q(WX11083), .QN(n3590) );
  SDFFX1 DFF_1616_Q_reg ( .D(WX11084), .SI(WX11083), .SE(n4399), .CLK(n5060), 
        .Q(WX11085), .QN(n9061) );
  SDFFX1 DFF_1617_Q_reg ( .D(WX11086), .SI(WX11085), .SE(n4399), .CLK(n5060), 
        .Q(WX11087), .QN(n9060) );
  SDFFX1 DFF_1618_Q_reg ( .D(WX11088), .SI(WX11087), .SE(n4398), .CLK(n5060), 
        .Q(WX11089), .QN(n9059) );
  SDFFX1 DFF_1619_Q_reg ( .D(WX11090), .SI(WX11089), .SE(n4397), .CLK(n5061), 
        .Q(WX11091), .QN(n9058) );
  SDFFX1 DFF_1620_Q_reg ( .D(WX11092), .SI(WX11091), .SE(n4396), .CLK(n5061), 
        .Q(WX11093), .QN(n9057) );
  SDFFX1 DFF_1621_Q_reg ( .D(WX11094), .SI(WX11093), .SE(n4396), .CLK(n5061), 
        .Q(WX11095), .QN(n9056) );
  SDFFX1 DFF_1622_Q_reg ( .D(WX11096), .SI(WX11095), .SE(n4396), .CLK(n5061), 
        .Q(WX11097), .QN(n9055) );
  SDFFX1 DFF_1623_Q_reg ( .D(WX11098), .SI(WX11097), .SE(n4395), .CLK(n5062), 
        .Q(WX11099), .QN(n9054) );
  SDFFX1 DFF_1624_Q_reg ( .D(WX11100), .SI(WX11099), .SE(n4395), .CLK(n5062), 
        .Q(WX11101), .QN(n9053) );
  SDFFX1 DFF_1625_Q_reg ( .D(WX11102), .SI(WX11101), .SE(n4394), .CLK(n5062), 
        .Q(test_so94) );
  SDFFX1 DFF_1626_Q_reg ( .D(WX11104), .SI(test_si95), .SE(n4394), .CLK(n5063), 
        .Q(WX11105), .QN(n9051) );
  SDFFX1 DFF_1627_Q_reg ( .D(WX11106), .SI(WX11105), .SE(n4393), .CLK(n5063), 
        .Q(WX11107), .QN(n9050) );
  SDFFX1 DFF_1628_Q_reg ( .D(WX11108), .SI(WX11107), .SE(n4393), .CLK(n5063), 
        .Q(WX11109), .QN(n9049) );
  SDFFX1 DFF_1629_Q_reg ( .D(WX11110), .SI(WX11109), .SE(n4392), .CLK(n5064), 
        .Q(WX11111), .QN(n9048) );
  SDFFX1 DFF_1630_Q_reg ( .D(WX11112), .SI(WX11111), .SE(n4391), .CLK(n5064), 
        .Q(WX11113), .QN(n9047) );
  SDFFX1 DFF_1631_Q_reg ( .D(WX11114), .SI(WX11113), .SE(n4391), .CLK(n5064), 
        .Q(WX11115), .QN(n9046) );
  SDFFX1 DFF_1632_Q_reg ( .D(WX11116), .SI(WX11115), .SE(n4390), .CLK(n5065), 
        .Q(WX11117) );
  SDFFX1 DFF_1633_Q_reg ( .D(WX11118), .SI(WX11117), .SE(n4390), .CLK(n5065), 
        .Q(WX11119) );
  SDFFX1 DFF_1634_Q_reg ( .D(WX11120), .SI(WX11119), .SE(n4389), .CLK(n5065), 
        .Q(WX11121) );
  SDFFX1 DFF_1635_Q_reg ( .D(WX11122), .SI(WX11121), .SE(n4389), .CLK(n5065), 
        .Q(WX11123) );
  SDFFX1 DFF_1636_Q_reg ( .D(WX11124), .SI(WX11123), .SE(n4389), .CLK(n5065), 
        .Q(WX11125) );
  SDFFX1 DFF_1637_Q_reg ( .D(WX11126), .SI(WX11125), .SE(n4388), .CLK(n5066), 
        .Q(WX11127) );
  SDFFX1 DFF_1638_Q_reg ( .D(WX11128), .SI(WX11127), .SE(n4388), .CLK(n5066), 
        .Q(WX11129), .QN(n3597) );
  SDFFX1 DFF_1639_Q_reg ( .D(WX11130), .SI(WX11129), .SE(n4388), .CLK(n5066), 
        .Q(WX11131) );
  SDFFX1 DFF_1640_Q_reg ( .D(WX11132), .SI(WX11131), .SE(n4403), .CLK(n5058), 
        .Q(WX11133), .QN(n9073) );
  SDFFX1 DFF_1641_Q_reg ( .D(WX11134), .SI(WX11133), .SE(n4403), .CLK(n5058), 
        .Q(WX11135) );
  SDFFX1 DFF_1642_Q_reg ( .D(WX11136), .SI(WX11135), .SE(n4403), .CLK(n5058), 
        .Q(test_so95), .QN(n9068) );
  SDFFX1 DFF_1643_Q_reg ( .D(WX11138), .SI(test_si96), .SE(n4402), .CLK(n5058), 
        .Q(WX11139) );
  SDFFX1 DFF_1644_Q_reg ( .D(WX11140), .SI(WX11139), .SE(n4402), .CLK(n5058), 
        .Q(WX11141), .QN(n3593) );
  SDFFX1 DFF_1645_Q_reg ( .D(WX11142), .SI(WX11141), .SE(n4401), .CLK(n5059), 
        .Q(WX11143) );
  SDFFX1 DFF_1646_Q_reg ( .D(WX11144), .SI(WX11143), .SE(n4400), .CLK(n5059), 
        .Q(WX11145) );
  SDFFX1 DFF_1647_Q_reg ( .D(WX11146), .SI(WX11145), .SE(n4400), .CLK(n5059), 
        .Q(WX11147) );
  SDFFX1 DFF_1648_Q_reg ( .D(WX11148), .SI(WX11147), .SE(n4399), .CLK(n5060), 
        .Q(WX11149), .QN(n3724) );
  SDFFX1 DFF_1649_Q_reg ( .D(WX11150), .SI(WX11149), .SE(n4398), .CLK(n5060), 
        .Q(WX11151), .QN(n3722) );
  SDFFX1 DFF_1650_Q_reg ( .D(WX11152), .SI(WX11151), .SE(n4398), .CLK(n5060), 
        .Q(WX11153), .QN(n3720) );
  SDFFX1 DFF_1651_Q_reg ( .D(WX11154), .SI(WX11153), .SE(n4397), .CLK(n5061), 
        .Q(WX11155), .QN(n3718) );
  SDFFX1 DFF_1652_Q_reg ( .D(WX11156), .SI(WX11155_Tj_Payload), .SE(
        test_se_Trojan), .CLK(n5015), .Q(WX11157), .QN(n3716) );
  SDFFX1 DFF_1653_Q_reg ( .D(WX11158), .SI(WX11157), .SE(test_se_Trojan), 
        .CLK(n5061), .Q(WX11159), .QN(n3714) );
  SDFFX1 DFF_1654_Q_reg ( .D(WX11160), .SI(WX11159), .SE(test_se_Trojan), 
        .CLK(n5062), .Q(WX11161), .QN(n3712) );
  SDFFX1 DFF_1655_Q_reg ( .D(WX11162), .SI(WX11161), .SE(test_se_Trojan), 
        .CLK(n5062), .Q(WX11163) );
  SDFFX1 DFF_1656_Q_reg ( .D(WX11164), .SI(WX11163), .SE(test_se_Trojan), 
        .CLK(n5062), .Q(WX11165), .QN(n3709) );
  SDFFX1 DFF_1657_Q_reg ( .D(WX11166), .SI(WX11165), .SE(test_se_Trojan), 
        .CLK(n5063), .Q(WX11167), .QN(n9052) );
  SDFFX1 DFF_1658_Q_reg ( .D(WX11168), .SI(WX11167), .SE(test_se_Trojan), 
        .CLK(n5063), .Q(WX11169), .QN(n3706) );
  SDFFX1 DFF_1659_Q_reg ( .D(WX11170), .SI(WX11169), .SE(test_se_Trojan), 
        .CLK(n5063), .Q(test_so96) );
  SDFFX1 DFF_1660_Q_reg ( .D(WX11172), .SI(test_si97), .SE(n4392), .CLK(n5064), 
        .Q(WX11173), .QN(n3703) );
  SDFFX1 DFF_1661_Q_reg ( .D(WX11174), .SI(WX11173), .SE(n4392), .CLK(n5064), 
        .Q(WX11175), .QN(n3701) );
  SDFFX1 DFF_1662_Q_reg ( .D(WX11176), .SI(WX11175), .SE(n4391), .CLK(n5064), 
        .Q(WX11177), .QN(n3699) );
  SDFFX1 DFF_1663_Q_reg ( .D(WX11178), .SI(WX11177), .SE(n4390), .CLK(n5065), 
        .Q(WX11179), .QN(n3697) );
  SDFFX1 DFF_1664_Q_reg ( .D(WX11180), .SI(WX11179), .SE(n4390), .CLK(n5065), 
        .Q(WX11181), .QN(n3968) );
  SDFFX1 DFF_1665_Q_reg ( .D(WX11182), .SI(WX11181), .SE(n4390), .CLK(n5065), 
        .Q(WX11183), .QN(n3969) );
  SDFFX1 DFF_1666_Q_reg ( .D(WX11184), .SI(WX11183), .SE(n4389), .CLK(n5065), 
        .Q(WX11185), .QN(n3970) );
  SDFFX1 DFF_1667_Q_reg ( .D(WX11186), .SI(WX11185), .SE(n4389), .CLK(n5065), 
        .Q(WX11187), .QN(n3971) );
  SDFFX1 DFF_1668_Q_reg ( .D(WX11188), .SI(WX11187), .SE(n4389), .CLK(n5065), 
        .Q(WX11189), .QN(n3972) );
  SDFFX1 DFF_1669_Q_reg ( .D(WX11190), .SI(WX11189), .SE(n4388), .CLK(n5066), 
        .Q(WX11191), .QN(n3973) );
  SDFFX1 DFF_1670_Q_reg ( .D(WX11192), .SI(WX11191), .SE(n4388), .CLK(n5066), 
        .Q(WX11193), .QN(n3974) );
  SDFFX1 DFF_1671_Q_reg ( .D(WX11194), .SI(WX11193), .SE(n4388), .CLK(n5066), 
        .Q(WX11195), .QN(n3975) );
  SDFFX1 DFF_1672_Q_reg ( .D(WX11196), .SI(WX11195), .SE(n4387), .CLK(n5066), 
        .Q(WX11197), .QN(n3976) );
  SDFFX1 DFF_1673_Q_reg ( .D(WX11198), .SI(WX11197), .SE(n4387), .CLK(n5066), 
        .Q(WX11199), .QN(n3977) );
  SDFFX1 DFF_1674_Q_reg ( .D(WX11200), .SI(WX11199), .SE(n4387), .CLK(n5066), 
        .Q(WX11201), .QN(n3978) );
  SDFFX1 DFF_1675_Q_reg ( .D(WX11202), .SI(WX11201), .SE(n4387), .CLK(n5066), 
        .Q(WX11203), .QN(n3979) );
  SDFFX1 DFF_1676_Q_reg ( .D(WX11204), .SI(WX11203), .SE(n4387), .CLK(n5066), 
        .Q(test_so97) );
  SDFFX1 DFF_1677_Q_reg ( .D(WX11206), .SI(test_si98), .SE(n4401), .CLK(n5059), 
        .Q(WX11207), .QN(n3980) );
  SDFFX1 DFF_1678_Q_reg ( .D(WX11208), .SI(WX11207), .SE(n4400), .CLK(n5059), 
        .Q(WX11209), .QN(n3981) );
  SDFFX1 DFF_1679_Q_reg ( .D(WX11210), .SI(WX11209), .SE(n4400), .CLK(n5059), 
        .Q(WX11211), .QN(n3939) );
  SDFFX1 DFF_1680_Q_reg ( .D(WX11212), .SI(WX11211), .SE(n4399), .CLK(n5060), 
        .Q(WX11213), .QN(n3982) );
  SDFFX1 DFF_1681_Q_reg ( .D(WX11214), .SI(WX11213), .SE(n4398), .CLK(n5060), 
        .Q(WX11215), .QN(n3983) );
  SDFFX1 DFF_1682_Q_reg ( .D(WX11216), .SI(WX11215), .SE(n4398), .CLK(n5060), 
        .Q(WX11217), .QN(n3984) );
  SDFFX1 DFF_1683_Q_reg ( .D(WX11218), .SI(WX11217), .SE(n4397), .CLK(n5061), 
        .Q(WX11219), .QN(n3985) );
  SDFFX1 DFF_1684_Q_reg ( .D(WX11220), .SI(WX11219), .SE(n4397), .CLK(n5061), 
        .Q(WX11221), .QN(n3940) );
  SDFFX1 DFF_1685_Q_reg ( .D(WX11222), .SI(WX11221), .SE(n4396), .CLK(n5061), 
        .Q(WX11223), .QN(n3986) );
  SDFFX1 DFF_1686_Q_reg ( .D(WX11224), .SI(WX11223), .SE(n4395), .CLK(n5062), 
        .Q(WX11225), .QN(n3987) );
  SDFFX1 DFF_1687_Q_reg ( .D(WX11226), .SI(WX11225), .SE(n4395), .CLK(n5062), 
        .Q(WX11227), .QN(n3988) );
  SDFFX1 DFF_1688_Q_reg ( .D(WX11228), .SI(WX11227), .SE(n4395), .CLK(n5062), 
        .Q(WX11229), .QN(n3989) );
  SDFFX1 DFF_1689_Q_reg ( .D(WX11230), .SI(WX11229), .SE(n4394), .CLK(n5063), 
        .Q(WX11231), .QN(n3990) );
  SDFFX1 DFF_1690_Q_reg ( .D(WX11232), .SI(WX11231), .SE(n4393), .CLK(n5063), 
        .Q(WX11233), .QN(n3991) );
  SDFFX1 DFF_1691_Q_reg ( .D(WX11234), .SI(WX11233), .SE(n4393), .CLK(n5063), 
        .Q(WX11235), .QN(n3941) );
  SDFFX1 DFF_1692_Q_reg ( .D(WX11236), .SI(WX11235), .SE(n4392), .CLK(n5064), 
        .Q(WX11237), .QN(n3992) );
  SDFFX1 DFF_1693_Q_reg ( .D(WX11238), .SI(WX11237), .SE(n4392), .CLK(n5064), 
        .Q(test_so98) );
  SDFFX1 DFF_1694_Q_reg ( .D(WX11240), .SI(test_si99), .SE(n4391), .CLK(n5064), 
        .Q(WX11241), .QN(n3993) );
  SDFFX1 DFF_1695_Q_reg ( .D(WX11242), .SI(WX11241), .SE(n4390), .CLK(n5065), 
        .Q(WX11243), .QN(n3960) );
  SDFFX1 DFF_1696_Q_reg ( .D(WX11608), .SI(WX11243), .SE(n4385), .CLK(n5067), 
        .Q(CRC_OUT_1_0), .QN(DFF_1696_n1) );
  SDFFX1 DFF_1697_Q_reg ( .D(WX11610), .SI(CRC_OUT_1_0), .SE(n4385), .CLK(
        n5067), .Q(CRC_OUT_1_1), .QN(DFF_1697_n1) );
  SDFFX1 DFF_1698_Q_reg ( .D(WX11612), .SI(CRC_OUT_1_1), .SE(n4385), .CLK(
        n5067), .Q(CRC_OUT_1_2), .QN(DFF_1698_n1) );
  SDFFX1 DFF_1699_Q_reg ( .D(WX11614), .SI(CRC_OUT_1_2), .SE(n4385), .CLK(
        n5067), .Q(CRC_OUT_1_3), .QN(DFF_1699_n1) );
  SDFFX1 DFF_1700_Q_reg ( .D(WX11616), .SI(CRC_OUT_1_3), .SE(n4385), .CLK(
        n5067), .Q(CRC_OUT_1_4), .QN(DFF_1700_n1) );
  SDFFX1 DFF_1701_Q_reg ( .D(WX11618), .SI(CRC_OUT_1_4), .SE(n4384), .CLK(
        n5068), .Q(CRC_OUT_1_5), .QN(DFF_1701_n1) );
  SDFFX1 DFF_1702_Q_reg ( .D(WX11620), .SI(CRC_OUT_1_5), .SE(n4384), .CLK(
        n5068), .Q(CRC_OUT_1_6), .QN(DFF_1702_n1) );
  SDFFX1 DFF_1703_Q_reg ( .D(WX11622), .SI(CRC_OUT_1_6), .SE(n4384), .CLK(
        n5068), .Q(CRC_OUT_1_7), .QN(DFF_1703_n1) );
  SDFFX1 DFF_1704_Q_reg ( .D(WX11624), .SI(CRC_OUT_1_7), .SE(n4384), .CLK(
        n5068), .Q(CRC_OUT_1_8), .QN(DFF_1704_n1) );
  SDFFX1 DFF_1705_Q_reg ( .D(WX11626), .SI(CRC_OUT_1_8), .SE(n4384), .CLK(
        n5068), .Q(CRC_OUT_1_9), .QN(DFF_1705_n1) );
  SDFFX1 DFF_1706_Q_reg ( .D(WX11628), .SI(CRC_OUT_1_9), .SE(n4384), .CLK(
        n5068), .Q(CRC_OUT_1_10), .QN(DFF_1706_n1) );
  SDFFX1 DFF_1707_Q_reg ( .D(WX11630), .SI(CRC_OUT_1_10), .SE(n4383), .CLK(
        n5068), .Q(CRC_OUT_1_11), .QN(DFF_1707_n1) );
  SDFFX1 DFF_1708_Q_reg ( .D(WX11632), .SI(CRC_OUT_1_11), .SE(n4383), .CLK(
        n5068), .Q(CRC_OUT_1_12), .QN(DFF_1708_n1) );
  SDFFX1 DFF_1709_Q_reg ( .D(WX11634), .SI(CRC_OUT_1_12), .SE(n4383), .CLK(
        n5068), .Q(CRC_OUT_1_13), .QN(DFF_1709_n1) );
  SDFFX1 DFF_1710_Q_reg ( .D(WX11636), .SI(CRC_OUT_1_13), .SE(n4383), .CLK(
        n5068), .Q(test_so99) );
  SDFFX1 DFF_1711_Q_reg ( .D(WX11638), .SI(test_si100), .SE(n4383), .CLK(n5068), .Q(CRC_OUT_1_15), .QN(DFF_1711_n1) );
  SDFFX1 DFF_1712_Q_reg ( .D(WX11640), .SI(CRC_OUT_1_15), .SE(n4383), .CLK(
        n5068), .Q(CRC_OUT_1_16), .QN(DFF_1712_n1) );
  SDFFX1 DFF_1713_Q_reg ( .D(WX11642), .SI(CRC_OUT_1_16), .SE(n4382), .CLK(
        n5069), .Q(CRC_OUT_1_17), .QN(DFF_1713_n1) );
  SDFFX1 DFF_1714_Q_reg ( .D(WX11644), .SI(CRC_OUT_1_17), .SE(n4382), .CLK(
        n5069), .Q(CRC_OUT_1_18), .QN(DFF_1714_n1) );
  SDFFX1 DFF_1715_Q_reg ( .D(WX11646), .SI(CRC_OUT_1_18), .SE(n4382), .CLK(
        n5069), .Q(CRC_OUT_1_19), .QN(DFF_1715_n1) );
  SDFFX1 DFF_1716_Q_reg ( .D(WX11648), .SI(CRC_OUT_1_19), .SE(n4382), .CLK(
        n5069), .Q(CRC_OUT_1_20), .QN(DFF_1716_n1) );
  SDFFX1 DFF_1717_Q_reg ( .D(WX11650), .SI(CRC_OUT_1_20), .SE(n4382), .CLK(
        n5069), .Q(CRC_OUT_1_21), .QN(DFF_1717_n1) );
  SDFFX1 DFF_1718_Q_reg ( .D(WX11652), .SI(CRC_OUT_1_21), .SE(n4382), .CLK(
        n5069), .Q(CRC_OUT_1_22), .QN(DFF_1718_n1) );
  SDFFX1 DFF_1719_Q_reg ( .D(WX11654), .SI(CRC_OUT_1_22), .SE(n4381), .CLK(
        n5069), .Q(CRC_OUT_1_23), .QN(DFF_1719_n1) );
  SDFFX1 DFF_1720_Q_reg ( .D(WX11656), .SI(CRC_OUT_1_23), .SE(n4387), .CLK(
        n5066), .Q(CRC_OUT_1_24), .QN(DFF_1720_n1) );
  SDFFX1 DFF_1721_Q_reg ( .D(WX11658), .SI(CRC_OUT_1_24), .SE(n4386), .CLK(
        n5067), .Q(CRC_OUT_1_25), .QN(DFF_1721_n1) );
  SDFFX1 DFF_1722_Q_reg ( .D(WX11660), .SI(CRC_OUT_1_25), .SE(n4386), .CLK(
        n5067), .Q(CRC_OUT_1_26), .QN(DFF_1722_n1) );
  SDFFX1 DFF_1723_Q_reg ( .D(WX11662), .SI(CRC_OUT_1_26), .SE(n4386), .CLK(
        n5067), .Q(CRC_OUT_1_27), .QN(DFF_1723_n1) );
  SDFFX1 DFF_1724_Q_reg ( .D(WX11664), .SI(CRC_OUT_1_27), .SE(n4386), .CLK(
        n5067), .Q(CRC_OUT_1_28), .QN(DFF_1724_n1) );
  SDFFX1 DFF_1725_Q_reg ( .D(WX11666), .SI(CRC_OUT_1_28), .SE(n4386), .CLK(
        n5067), .Q(CRC_OUT_1_29), .QN(DFF_1725_n1) );
  SDFFX1 DFF_1726_Q_reg ( .D(WX11668), .SI(CRC_OUT_1_29), .SE(n4386), .CLK(
        n5067), .Q(CRC_OUT_1_30), .QN(DFF_1726_n1) );
  SDFFX1 DFF_1727_Q_reg ( .D(WX11670), .SI(CRC_OUT_1_30), .SE(n4385), .CLK(
        n5067), .Q(test_so100), .QN(n4245) );
  AND2X1 Trojan1 ( .IN1(WX742), .IN2(WX7249), .Q(Tj_OUT1) );
  AND2X1 Trojan2 ( .IN1(WX5922), .IN2(WX5960), .Q(Tj_OUT2) );
  AND2X1 Trojan3 ( .IN1(WX4697), .IN2(WX9032), .Q(Tj_OUT3) );
  AND2X1 Trojan4 ( .IN1(n185), .IN2(WX10846), .Q(Tj_OUT4) );
  NOR4X0 Trojan1234_NOT ( .IN1(Tj_OUT1), .IN2(Tj_OUT2), .IN3(Tj_OUT3), .IN4(
        Tj_OUT4), .QN(Tj_OUT1234) );
  AND2X1 Trojan5 ( .IN1(WX3340), .IN2(WX6476), .Q(Tj_OUT5) );
  AND2X1 Trojan6 ( .IN1(WX9819), .IN2(n20), .Q(Tj_OUT6) );
  AND2X1 Trojan7 ( .IN1(n122), .IN2(WX3458), .Q(Tj_OUT7) );
  AND2X1 Trojan8 ( .IN1(WX9060), .IN2(WX7749), .Q(Tj_OUT8) );
  NOR4X0 Trojan5678_NOT ( .IN1(Tj_OUT5), .IN2(Tj_OUT6), .IN3(Tj_OUT7), .IN4(
        Tj_OUT8), .QN(Tj_OUT5678) );
  INVX0 TrojanINV_test_se ( .INP(n4627), .ZN(test_se_NOT) );
  AND3X1 Trojan_Trigger ( .IN1(Tj_OUT1234), .IN2(Tj_OUT5678), .IN3(test_se_NOT), .Q(Tj_Trigger) );
  DFFX2 TrojanScanEnable ( .D(1'b1), .CLK(Tj_Trigger), .Q(Trojan_SE) );
  MUX21X1 Trojan_Payload1 ( .IN1(n4627), .IN2(1'b1), .S(Trojan_SE), .Q(
        test_se_Trojan) );
  MUX21X1 Trojan_Payload2 ( .IN1(WX11155), .IN2(WX3442), .S(Trojan_SE), .Q(
        WX11155_Tj_Payload) );
  NBUFFX2 U4327 ( .INP(n5118), .Z(n4949) );
  NBUFFX2 U4328 ( .INP(n5118), .Z(n4947) );
  NBUFFX2 U4329 ( .INP(n5118), .Z(n4948) );
  NBUFFX2 U4330 ( .INP(n5118), .Z(n4946) );
  NBUFFX2 U4331 ( .INP(n5094), .Z(n5068) );
  NBUFFX2 U4332 ( .INP(n5094), .Z(n5067) );
  NBUFFX2 U4333 ( .INP(n5094), .Z(n5066) );
  NBUFFX2 U4334 ( .INP(n5094), .Z(n5065) );
  NBUFFX2 U4335 ( .INP(n5095), .Z(n5064) );
  NBUFFX2 U4336 ( .INP(n5095), .Z(n5063) );
  NBUFFX2 U4337 ( .INP(n5095), .Z(n5062) );
  NBUFFX2 U4338 ( .INP(n5095), .Z(n5061) );
  NBUFFX2 U4339 ( .INP(n5095), .Z(n5060) );
  NBUFFX2 U4340 ( .INP(n5096), .Z(n5059) );
  NBUFFX2 U4341 ( .INP(n5096), .Z(n5058) );
  NBUFFX2 U4342 ( .INP(n5096), .Z(n5057) );
  NBUFFX2 U4343 ( .INP(n5097), .Z(n5054) );
  NBUFFX2 U4344 ( .INP(n5096), .Z(n5055) );
  NBUFFX2 U4345 ( .INP(n5096), .Z(n5056) );
  NBUFFX2 U4346 ( .INP(n5097), .Z(n5053) );
  NBUFFX2 U4347 ( .INP(n5093), .Z(n5070) );
  NBUFFX2 U4348 ( .INP(n5094), .Z(n5069) );
  NBUFFX2 U4349 ( .INP(n5097), .Z(n5052) );
  NBUFFX2 U4350 ( .INP(n5097), .Z(n5051) );
  NBUFFX2 U4351 ( .INP(n5097), .Z(n5050) );
  NBUFFX2 U4352 ( .INP(n5098), .Z(n5048) );
  NBUFFX2 U4353 ( .INP(n5098), .Z(n5047) );
  NBUFFX2 U4354 ( .INP(n5098), .Z(n5049) );
  NBUFFX2 U4355 ( .INP(n5098), .Z(n5046) );
  NBUFFX2 U4356 ( .INP(n5098), .Z(n5045) );
  NBUFFX2 U4357 ( .INP(n5099), .Z(n5044) );
  NBUFFX2 U4358 ( .INP(n5099), .Z(n5041) );
  NBUFFX2 U4359 ( .INP(n5099), .Z(n5042) );
  NBUFFX2 U4360 ( .INP(n5099), .Z(n5043) );
  NBUFFX2 U4361 ( .INP(n5093), .Z(n5072) );
  NBUFFX2 U4362 ( .INP(n5093), .Z(n5071) );
  NBUFFX2 U4363 ( .INP(n5099), .Z(n5040) );
  NBUFFX2 U4364 ( .INP(n5100), .Z(n5039) );
  NBUFFX2 U4365 ( .INP(n5100), .Z(n5038) );
  NBUFFX2 U4366 ( .INP(n5100), .Z(n5037) );
  NBUFFX2 U4367 ( .INP(n5100), .Z(n5036) );
  NBUFFX2 U4368 ( .INP(n5100), .Z(n5035) );
  NBUFFX2 U4369 ( .INP(n5101), .Z(n5034) );
  NBUFFX2 U4370 ( .INP(n5101), .Z(n5033) );
  NBUFFX2 U4371 ( .INP(n5101), .Z(n5032) );
  NBUFFX2 U4372 ( .INP(n5101), .Z(n5031) );
  NBUFFX2 U4373 ( .INP(n5093), .Z(n5073) );
  NBUFFX2 U4374 ( .INP(n5102), .Z(n5028) );
  NBUFFX2 U4375 ( .INP(n5102), .Z(n5029) );
  NBUFFX2 U4376 ( .INP(n5101), .Z(n5030) );
  NBUFFX2 U4377 ( .INP(n5092), .Z(n5075) );
  NBUFFX2 U4378 ( .INP(n5093), .Z(n5074) );
  NBUFFX2 U4379 ( .INP(n5102), .Z(n5027) );
  NBUFFX2 U4380 ( .INP(n5102), .Z(n5026) );
  NBUFFX2 U4381 ( .INP(n5102), .Z(n5025) );
  NBUFFX2 U4382 ( .INP(n5103), .Z(n5024) );
  NBUFFX2 U4383 ( .INP(n5103), .Z(n5023) );
  NBUFFX2 U4384 ( .INP(n5103), .Z(n5022) );
  NBUFFX2 U4385 ( .INP(n5103), .Z(n5021) );
  NBUFFX2 U4386 ( .INP(n5103), .Z(n5020) );
  NBUFFX2 U4387 ( .INP(n5104), .Z(n5019) );
  NBUFFX2 U4388 ( .INP(n5104), .Z(n5018) );
  NBUFFX2 U4389 ( .INP(n5104), .Z(n5017) );
  NBUFFX2 U4390 ( .INP(n5104), .Z(n5016) );
  NBUFFX2 U4391 ( .INP(n5105), .Z(n5012) );
  NBUFFX2 U4392 ( .INP(n5105), .Z(n5011) );
  NBUFFX2 U4393 ( .INP(n5104), .Z(n5015) );
  NBUFFX2 U4394 ( .INP(n5105), .Z(n5014) );
  NBUFFX2 U4395 ( .INP(n5105), .Z(n5013) );
  NBUFFX2 U4396 ( .INP(n5105), .Z(n5010) );
  NBUFFX2 U4397 ( .INP(n5106), .Z(n5009) );
  NBUFFX2 U4398 ( .INP(n5106), .Z(n5008) );
  NBUFFX2 U4399 ( .INP(n5106), .Z(n5007) );
  NBUFFX2 U4400 ( .INP(n5106), .Z(n5006) );
  NBUFFX2 U4401 ( .INP(n5106), .Z(n5005) );
  NBUFFX2 U4402 ( .INP(n5107), .Z(n5004) );
  NBUFFX2 U4403 ( .INP(n5107), .Z(n5003) );
  NBUFFX2 U4404 ( .INP(n5107), .Z(n5002) );
  NBUFFX2 U4405 ( .INP(n5092), .Z(n5076) );
  NBUFFX2 U4406 ( .INP(n5107), .Z(n5001) );
  NBUFFX2 U4407 ( .INP(n5107), .Z(n5000) );
  NBUFFX2 U4408 ( .INP(n5108), .Z(n4998) );
  NBUFFX2 U4409 ( .INP(n5108), .Z(n4999) );
  NBUFFX2 U4410 ( .INP(n5108), .Z(n4997) );
  NBUFFX2 U4411 ( .INP(n5092), .Z(n5078) );
  NBUFFX2 U4412 ( .INP(n5092), .Z(n5077) );
  NBUFFX2 U4413 ( .INP(n5108), .Z(n4996) );
  NBUFFX2 U4414 ( .INP(n5108), .Z(n4995) );
  NBUFFX2 U4415 ( .INP(n5109), .Z(n4994) );
  NBUFFX2 U4416 ( .INP(n5109), .Z(n4993) );
  NBUFFX2 U4417 ( .INP(n5109), .Z(n4992) );
  NBUFFX2 U4418 ( .INP(n5109), .Z(n4991) );
  NBUFFX2 U4419 ( .INP(n5109), .Z(n4990) );
  NBUFFX2 U4420 ( .INP(n5110), .Z(n4989) );
  NBUFFX2 U4421 ( .INP(n5110), .Z(n4988) );
  NBUFFX2 U4422 ( .INP(n5110), .Z(n4987) );
  NBUFFX2 U4423 ( .INP(n5111), .Z(n4984) );
  NBUFFX2 U4424 ( .INP(n5110), .Z(n4985) );
  NBUFFX2 U4425 ( .INP(n5110), .Z(n4986) );
  NBUFFX2 U4426 ( .INP(n5091), .Z(n5080) );
  NBUFFX2 U4427 ( .INP(n5092), .Z(n5079) );
  NBUFFX2 U4428 ( .INP(n5111), .Z(n4983) );
  NBUFFX2 U4429 ( .INP(n5111), .Z(n4982) );
  NBUFFX2 U4430 ( .INP(n5111), .Z(n4981) );
  NBUFFX2 U4431 ( .INP(n5111), .Z(n4980) );
  NBUFFX2 U4432 ( .INP(n5112), .Z(n4979) );
  NBUFFX2 U4433 ( .INP(n5112), .Z(n4978) );
  NBUFFX2 U4434 ( .INP(n5112), .Z(n4977) );
  NBUFFX2 U4435 ( .INP(n5112), .Z(n4976) );
  NBUFFX2 U4436 ( .INP(n5112), .Z(n4975) );
  NBUFFX2 U4437 ( .INP(n5113), .Z(n4974) );
  NBUFFX2 U4438 ( .INP(n5113), .Z(n4973) );
  NBUFFX2 U4439 ( .INP(n5113), .Z(n4970) );
  NBUFFX2 U4440 ( .INP(n5113), .Z(n4971) );
  NBUFFX2 U4441 ( .INP(n5113), .Z(n4972) );
  NBUFFX2 U4442 ( .INP(n5091), .Z(n5083) );
  NBUFFX2 U4443 ( .INP(n5091), .Z(n5082) );
  NBUFFX2 U4444 ( .INP(n5091), .Z(n5081) );
  NBUFFX2 U4445 ( .INP(n5090), .Z(n5087) );
  NBUFFX2 U4446 ( .INP(n5090), .Z(n5086) );
  NBUFFX2 U4447 ( .INP(n5090), .Z(n5085) );
  NBUFFX2 U4448 ( .INP(n5114), .Z(n4969) );
  NBUFFX2 U4449 ( .INP(n5114), .Z(n4968) );
  NBUFFX2 U4450 ( .INP(n5114), .Z(n4967) );
  NBUFFX2 U4451 ( .INP(n5114), .Z(n4966) );
  NBUFFX2 U4452 ( .INP(n5114), .Z(n4965) );
  NBUFFX2 U4453 ( .INP(n5115), .Z(n4964) );
  NBUFFX2 U4454 ( .INP(n5091), .Z(n5084) );
  NBUFFX2 U4455 ( .INP(n5115), .Z(n4963) );
  NBUFFX2 U4456 ( .INP(n5115), .Z(n4961) );
  NBUFFX2 U4457 ( .INP(n5115), .Z(n4962) );
  NBUFFX2 U4458 ( .INP(n5115), .Z(n4960) );
  NBUFFX2 U4459 ( .INP(n5090), .Z(n5088) );
  NBUFFX2 U4460 ( .INP(n5116), .Z(n4959) );
  NBUFFX2 U4461 ( .INP(n5116), .Z(n4958) );
  NBUFFX2 U4462 ( .INP(n5116), .Z(n4957) );
  NBUFFX2 U4463 ( .INP(n5116), .Z(n4956) );
  NBUFFX2 U4464 ( .INP(n5116), .Z(n4955) );
  NBUFFX2 U4465 ( .INP(n5117), .Z(n4954) );
  NBUFFX2 U4466 ( .INP(n5090), .Z(n5089) );
  NBUFFX2 U4467 ( .INP(n5117), .Z(n4953) );
  NBUFFX2 U4468 ( .INP(n5117), .Z(n4952) );
  NBUFFX2 U4469 ( .INP(n5117), .Z(n4951) );
  NBUFFX2 U4470 ( .INP(n5117), .Z(n4950) );
  NBUFFX2 U4471 ( .INP(n4272), .Z(n4280) );
  NBUFFX2 U4472 ( .INP(n4325), .Z(n4338) );
  NBUFFX2 U4473 ( .INP(n4325), .Z(n4339) );
  NBUFFX2 U4474 ( .INP(n4325), .Z(n4337) );
  NBUFFX2 U4475 ( .INP(n4272), .Z(n4277) );
  NBUFFX2 U4476 ( .INP(n4272), .Z(n4276) );
  NBUFFX2 U4477 ( .INP(n4272), .Z(n4279) );
  NBUFFX2 U4478 ( .INP(n4272), .Z(n4278) );
  NBUFFX2 U4479 ( .INP(n4275), .Z(n4295) );
  NBUFFX2 U4480 ( .INP(n4323), .Z(n4326) );
  NBUFFX2 U4481 ( .INP(n4323), .Z(n4328) );
  NBUFFX2 U4482 ( .INP(n4323), .Z(n4329) );
  NBUFFX2 U4483 ( .INP(n4324), .Z(n4331) );
  NBUFFX2 U4484 ( .INP(n4325), .Z(n4336) );
  NBUFFX2 U4485 ( .INP(n4324), .Z(n4334) );
  NBUFFX2 U4486 ( .INP(n4324), .Z(n4335) );
  NBUFFX2 U4487 ( .INP(n4324), .Z(n4333) );
  NBUFFX2 U4488 ( .INP(n4324), .Z(n4332) );
  NBUFFX2 U4489 ( .INP(n4323), .Z(n4327) );
  NBUFFX2 U4490 ( .INP(n4323), .Z(n4330) );
  NBUFFX2 U4491 ( .INP(n4274), .Z(n4286) );
  NBUFFX2 U4492 ( .INP(n4273), .Z(n4285) );
  NBUFFX2 U4493 ( .INP(n4273), .Z(n4284) );
  NBUFFX2 U4494 ( .INP(n4273), .Z(n4282) );
  NBUFFX2 U4495 ( .INP(n4273), .Z(n4281) );
  NBUFFX2 U4496 ( .INP(n4273), .Z(n4283) );
  NBUFFX2 U4497 ( .INP(n4275), .Z(n4294) );
  NBUFFX2 U4498 ( .INP(n4275), .Z(n4293) );
  NBUFFX2 U4499 ( .INP(n4275), .Z(n4292) );
  NBUFFX2 U4500 ( .INP(n4274), .Z(n4290) );
  NBUFFX2 U4501 ( .INP(n4275), .Z(n4291) );
  NBUFFX2 U4502 ( .INP(n4274), .Z(n4289) );
  NBUFFX2 U4503 ( .INP(n4274), .Z(n4288) );
  NBUFFX2 U4504 ( .INP(n4274), .Z(n4287) );
  NBUFFX2 U4505 ( .INP(n4325), .Z(n4340) );
  NBUFFX2 U4506 ( .INP(n4786), .Z(n4772) );
  NBUFFX2 U4507 ( .INP(n4786), .Z(n4773) );
  NBUFFX2 U4508 ( .INP(n4786), .Z(n4771) );
  NBUFFX2 U4509 ( .INP(n4785), .Z(n4774) );
  NBUFFX2 U4510 ( .INP(n4785), .Z(n4775) );
  NBUFFX2 U4511 ( .INP(n4785), .Z(n4776) );
  NBUFFX2 U4512 ( .INP(n4785), .Z(n4777) );
  NBUFFX2 U4513 ( .INP(n4785), .Z(n4778) );
  NBUFFX2 U4514 ( .INP(n4784), .Z(n4779) );
  NBUFFX2 U4515 ( .INP(n4784), .Z(n4782) );
  NBUFFX2 U4516 ( .INP(n4784), .Z(n4781) );
  NBUFFX2 U4517 ( .INP(n4784), .Z(n4780) );
  INVX0 U4518 ( .INP(n5352), .ZN(n4271) );
  INVX0 U4519 ( .INP(n5356), .ZN(n4322) );
  NBUFFX2 U4520 ( .INP(n4784), .Z(n4783) );
  INVX0 U4521 ( .INP(n4262), .ZN(n4246) );
  INVX0 U4522 ( .INP(n4262), .ZN(n4247) );
  INVX0 U4523 ( .INP(n4262), .ZN(n4248) );
  INVX0 U4524 ( .INP(n4262), .ZN(n4249) );
  INVX0 U4525 ( .INP(n4262), .ZN(n4250) );
  INVX0 U4526 ( .INP(n4262), .ZN(n4251) );
  INVX0 U4527 ( .INP(n4262), .ZN(n4252) );
  INVX0 U4528 ( .INP(n4262), .ZN(n4253) );
  INVX0 U4529 ( .INP(n4261), .ZN(n4254) );
  INVX0 U4530 ( .INP(n4261), .ZN(n4255) );
  INVX0 U4531 ( .INP(n4261), .ZN(n4256) );
  INVX0 U4532 ( .INP(n4261), .ZN(n4257) );
  INVX0 U4533 ( .INP(n4261), .ZN(n4258) );
  INVX0 U4534 ( .INP(n4261), .ZN(n4259) );
  INVX0 U4535 ( .INP(n4261), .ZN(n4260) );
  NBUFFX2 U4536 ( .INP(n4271), .Z(n4261) );
  NBUFFX2 U4537 ( .INP(n4271), .Z(n4262) );
  NBUFFX2 U4538 ( .INP(n4271), .Z(n4263) );
  NBUFFX2 U4539 ( .INP(n4271), .Z(n4264) );
  NBUFFX2 U4540 ( .INP(n4271), .Z(n4265) );
  NBUFFX2 U4541 ( .INP(n4261), .Z(n4266) );
  NBUFFX2 U4542 ( .INP(n4262), .Z(n4267) );
  NBUFFX2 U4543 ( .INP(n4265), .Z(n4268) );
  NBUFFX2 U4544 ( .INP(n4263), .Z(n4269) );
  NBUFFX2 U4545 ( .INP(n4264), .Z(n4270) );
  NBUFFX2 U4546 ( .INP(n5355), .Z(n4272) );
  NBUFFX2 U4547 ( .INP(n5355), .Z(n4273) );
  NBUFFX2 U4548 ( .INP(n5355), .Z(n4274) );
  NBUFFX2 U4549 ( .INP(n5355), .Z(n4275) );
  INVX0 U4550 ( .INP(n4315), .ZN(n4296) );
  INVX0 U4551 ( .INP(n4315), .ZN(n4297) );
  INVX0 U4552 ( .INP(n4315), .ZN(n4298) );
  INVX0 U4553 ( .INP(n4315), .ZN(n4299) );
  INVX0 U4554 ( .INP(n4314), .ZN(n4300) );
  INVX0 U4555 ( .INP(n4314), .ZN(n4301) );
  INVX0 U4556 ( .INP(n4314), .ZN(n4302) );
  INVX0 U4557 ( .INP(n4314), .ZN(n4303) );
  INVX0 U4558 ( .INP(n4314), .ZN(n4304) );
  INVX0 U4559 ( .INP(n4314), .ZN(n4305) );
  INVX0 U4560 ( .INP(n4314), .ZN(n4306) );
  INVX0 U4561 ( .INP(n4314), .ZN(n4307) );
  INVX0 U4562 ( .INP(n4313), .ZN(n4308) );
  INVX0 U4563 ( .INP(n4313), .ZN(n4309) );
  INVX0 U4564 ( .INP(n4313), .ZN(n4310) );
  INVX0 U4565 ( .INP(n4313), .ZN(n4311) );
  INVX0 U4566 ( .INP(n4313), .ZN(n4312) );
  NBUFFX2 U4567 ( .INP(n4322), .Z(n4313) );
  NBUFFX2 U4568 ( .INP(n4322), .Z(n4314) );
  NBUFFX2 U4569 ( .INP(n4322), .Z(n4315) );
  NBUFFX2 U4570 ( .INP(n4322), .Z(n4316) );
  NBUFFX2 U4571 ( .INP(n4313), .Z(n4317) );
  NBUFFX2 U4572 ( .INP(n4321), .Z(n4318) );
  NBUFFX2 U4573 ( .INP(n4322), .Z(n4319) );
  NBUFFX2 U4574 ( .INP(n4314), .Z(n4320) );
  NBUFFX2 U4575 ( .INP(n4315), .Z(n4321) );
  NBUFFX2 U4576 ( .INP(n5369), .Z(n4323) );
  NBUFFX2 U4577 ( .INP(n5369), .Z(n4324) );
  NBUFFX2 U4578 ( .INP(n5369), .Z(n4325) );
  NBUFFX2 U4579 ( .INP(n4723), .Z(n4341) );
  NBUFFX2 U4580 ( .INP(n4723), .Z(n4342) );
  NBUFFX2 U4581 ( .INP(n4722), .Z(n4343) );
  NBUFFX2 U4582 ( .INP(n4722), .Z(n4344) );
  NBUFFX2 U4583 ( .INP(n4722), .Z(n4345) );
  NBUFFX2 U4584 ( .INP(n4721), .Z(n4346) );
  NBUFFX2 U4585 ( .INP(n4721), .Z(n4347) );
  NBUFFX2 U4586 ( .INP(n4721), .Z(n4348) );
  NBUFFX2 U4587 ( .INP(n4720), .Z(n4349) );
  NBUFFX2 U4588 ( .INP(n4720), .Z(n4350) );
  NBUFFX2 U4589 ( .INP(n4720), .Z(n4351) );
  NBUFFX2 U4590 ( .INP(n4719), .Z(n4352) );
  NBUFFX2 U4591 ( .INP(n4719), .Z(n4353) );
  NBUFFX2 U4592 ( .INP(n4719), .Z(n4354) );
  NBUFFX2 U4593 ( .INP(n4718), .Z(n4355) );
  NBUFFX2 U4594 ( .INP(n4718), .Z(n4356) );
  NBUFFX2 U4595 ( .INP(n4718), .Z(n4357) );
  NBUFFX2 U4596 ( .INP(n4717), .Z(n4358) );
  NBUFFX2 U4597 ( .INP(n4717), .Z(n4359) );
  NBUFFX2 U4598 ( .INP(n4717), .Z(n4360) );
  NBUFFX2 U4599 ( .INP(n4716), .Z(n4361) );
  NBUFFX2 U4600 ( .INP(n4716), .Z(n4362) );
  NBUFFX2 U4601 ( .INP(n4716), .Z(n4363) );
  NBUFFX2 U4602 ( .INP(n4715), .Z(n4364) );
  NBUFFX2 U4603 ( .INP(n4715), .Z(n4365) );
  NBUFFX2 U4604 ( .INP(n4715), .Z(n4366) );
  NBUFFX2 U4605 ( .INP(n4714), .Z(n4367) );
  NBUFFX2 U4606 ( .INP(n4714), .Z(n4368) );
  NBUFFX2 U4607 ( .INP(n4714), .Z(n4369) );
  NBUFFX2 U4608 ( .INP(n4713), .Z(n4370) );
  NBUFFX2 U4609 ( .INP(n4713), .Z(n4371) );
  NBUFFX2 U4610 ( .INP(n4713), .Z(n4372) );
  NBUFFX2 U4611 ( .INP(n4712), .Z(n4373) );
  NBUFFX2 U4612 ( .INP(n4712), .Z(n4374) );
  NBUFFX2 U4613 ( .INP(n4712), .Z(n4375) );
  NBUFFX2 U4614 ( .INP(n4711), .Z(n4376) );
  NBUFFX2 U4615 ( .INP(n4711), .Z(n4377) );
  NBUFFX2 U4616 ( .INP(n4711), .Z(n4378) );
  NBUFFX2 U4617 ( .INP(n4710), .Z(n4379) );
  NBUFFX2 U4618 ( .INP(n4710), .Z(n4380) );
  NBUFFX2 U4619 ( .INP(n4710), .Z(n4381) );
  NBUFFX2 U4620 ( .INP(n4709), .Z(n4382) );
  NBUFFX2 U4621 ( .INP(n4709), .Z(n4383) );
  NBUFFX2 U4622 ( .INP(n4709), .Z(n4384) );
  NBUFFX2 U4623 ( .INP(n4708), .Z(n4385) );
  NBUFFX2 U4624 ( .INP(n4708), .Z(n4386) );
  NBUFFX2 U4625 ( .INP(n4708), .Z(n4387) );
  NBUFFX2 U4626 ( .INP(n4707), .Z(n4388) );
  NBUFFX2 U4627 ( .INP(n4707), .Z(n4389) );
  NBUFFX2 U4628 ( .INP(n4707), .Z(n4390) );
  NBUFFX2 U4629 ( .INP(n4706), .Z(n4391) );
  NBUFFX2 U4630 ( .INP(n4706), .Z(n4392) );
  NBUFFX2 U4631 ( .INP(n4706), .Z(n4393) );
  NBUFFX2 U4632 ( .INP(n4705), .Z(n4394) );
  NBUFFX2 U4633 ( .INP(n4705), .Z(n4395) );
  NBUFFX2 U4634 ( .INP(n4705), .Z(n4396) );
  NBUFFX2 U4635 ( .INP(n4704), .Z(n4397) );
  NBUFFX2 U4636 ( .INP(n4704), .Z(n4398) );
  NBUFFX2 U4637 ( .INP(n4704), .Z(n4399) );
  NBUFFX2 U4638 ( .INP(n4703), .Z(n4400) );
  NBUFFX2 U4639 ( .INP(n4703), .Z(n4401) );
  NBUFFX2 U4640 ( .INP(n4703), .Z(n4402) );
  NBUFFX2 U4641 ( .INP(n4702), .Z(n4403) );
  NBUFFX2 U4642 ( .INP(n4702), .Z(n4404) );
  NBUFFX2 U4643 ( .INP(n4702), .Z(n4405) );
  NBUFFX2 U4644 ( .INP(n4701), .Z(n4406) );
  NBUFFX2 U4645 ( .INP(n4701), .Z(n4407) );
  NBUFFX2 U4646 ( .INP(n4701), .Z(n4408) );
  NBUFFX2 U4647 ( .INP(n4700), .Z(n4409) );
  NBUFFX2 U4648 ( .INP(n4700), .Z(n4410) );
  NBUFFX2 U4649 ( .INP(n4700), .Z(n4411) );
  NBUFFX2 U4650 ( .INP(n4699), .Z(n4412) );
  NBUFFX2 U4651 ( .INP(n4699), .Z(n4413) );
  NBUFFX2 U4652 ( .INP(n4699), .Z(n4414) );
  NBUFFX2 U4653 ( .INP(n4698), .Z(n4415) );
  NBUFFX2 U4654 ( .INP(n4698), .Z(n4416) );
  NBUFFX2 U4655 ( .INP(n4698), .Z(n4417) );
  NBUFFX2 U4656 ( .INP(n4697), .Z(n4418) );
  NBUFFX2 U4657 ( .INP(n4697), .Z(n4419) );
  NBUFFX2 U4658 ( .INP(n4697), .Z(n4420) );
  NBUFFX2 U4659 ( .INP(n4696), .Z(n4421) );
  NBUFFX2 U4660 ( .INP(n4696), .Z(n4422) );
  NBUFFX2 U4661 ( .INP(n4696), .Z(n4423) );
  NBUFFX2 U4662 ( .INP(n4695), .Z(n4424) );
  NBUFFX2 U4663 ( .INP(n4695), .Z(n4425) );
  NBUFFX2 U4664 ( .INP(n4695), .Z(n4426) );
  NBUFFX2 U4665 ( .INP(n4694), .Z(n4427) );
  NBUFFX2 U4666 ( .INP(n4694), .Z(n4428) );
  NBUFFX2 U4667 ( .INP(n4694), .Z(n4429) );
  NBUFFX2 U4668 ( .INP(n4693), .Z(n4430) );
  NBUFFX2 U4669 ( .INP(n4693), .Z(n4431) );
  NBUFFX2 U4670 ( .INP(n4693), .Z(n4432) );
  NBUFFX2 U4671 ( .INP(n4692), .Z(n4433) );
  NBUFFX2 U4672 ( .INP(n4692), .Z(n4434) );
  NBUFFX2 U4673 ( .INP(n4692), .Z(n4435) );
  NBUFFX2 U4674 ( .INP(n4691), .Z(n4436) );
  NBUFFX2 U4675 ( .INP(n4691), .Z(n4437) );
  NBUFFX2 U4676 ( .INP(n4691), .Z(n4438) );
  NBUFFX2 U4677 ( .INP(n4690), .Z(n4439) );
  NBUFFX2 U4678 ( .INP(n4690), .Z(n4440) );
  NBUFFX2 U4679 ( .INP(n4690), .Z(n4441) );
  NBUFFX2 U4680 ( .INP(n4689), .Z(n4442) );
  NBUFFX2 U4681 ( .INP(n4689), .Z(n4443) );
  NBUFFX2 U4682 ( .INP(n4689), .Z(n4444) );
  NBUFFX2 U4683 ( .INP(n4688), .Z(n4445) );
  NBUFFX2 U4684 ( .INP(n4688), .Z(n4446) );
  NBUFFX2 U4685 ( .INP(n4688), .Z(n4447) );
  NBUFFX2 U4686 ( .INP(n4687), .Z(n4448) );
  NBUFFX2 U4687 ( .INP(n4687), .Z(n4449) );
  NBUFFX2 U4688 ( .INP(n4687), .Z(n4450) );
  NBUFFX2 U4689 ( .INP(n4686), .Z(n4451) );
  NBUFFX2 U4690 ( .INP(n4686), .Z(n4452) );
  NBUFFX2 U4691 ( .INP(n4686), .Z(n4453) );
  NBUFFX2 U4692 ( .INP(n4685), .Z(n4454) );
  NBUFFX2 U4693 ( .INP(n4685), .Z(n4455) );
  NBUFFX2 U4694 ( .INP(n4685), .Z(n4456) );
  NBUFFX2 U4695 ( .INP(n4684), .Z(n4457) );
  NBUFFX2 U4696 ( .INP(n4684), .Z(n4458) );
  NBUFFX2 U4697 ( .INP(n4684), .Z(n4459) );
  NBUFFX2 U4698 ( .INP(n4683), .Z(n4460) );
  NBUFFX2 U4699 ( .INP(n4683), .Z(n4461) );
  NBUFFX2 U4700 ( .INP(n4683), .Z(n4462) );
  NBUFFX2 U4701 ( .INP(n4682), .Z(n4463) );
  NBUFFX2 U4702 ( .INP(n4682), .Z(n4464) );
  NBUFFX2 U4703 ( .INP(n4682), .Z(n4465) );
  NBUFFX2 U4704 ( .INP(n4681), .Z(n4466) );
  NBUFFX2 U4705 ( .INP(n4681), .Z(n4467) );
  NBUFFX2 U4706 ( .INP(n4681), .Z(n4468) );
  NBUFFX2 U4707 ( .INP(n4680), .Z(n4469) );
  NBUFFX2 U4708 ( .INP(n4680), .Z(n4470) );
  NBUFFX2 U4709 ( .INP(n4680), .Z(n4471) );
  NBUFFX2 U4710 ( .INP(n4679), .Z(n4472) );
  NBUFFX2 U4711 ( .INP(n4679), .Z(n4473) );
  NBUFFX2 U4712 ( .INP(n4679), .Z(n4474) );
  NBUFFX2 U4713 ( .INP(n4678), .Z(n4475) );
  NBUFFX2 U4714 ( .INP(n4678), .Z(n4476) );
  NBUFFX2 U4715 ( .INP(n4678), .Z(n4477) );
  NBUFFX2 U4716 ( .INP(n4677), .Z(n4478) );
  NBUFFX2 U4717 ( .INP(n4677), .Z(n4479) );
  NBUFFX2 U4718 ( .INP(n4677), .Z(n4480) );
  NBUFFX2 U4719 ( .INP(n4676), .Z(n4481) );
  NBUFFX2 U4720 ( .INP(n4676), .Z(n4482) );
  NBUFFX2 U4721 ( .INP(n4676), .Z(n4483) );
  NBUFFX2 U4722 ( .INP(n4675), .Z(n4484) );
  NBUFFX2 U4723 ( .INP(n4675), .Z(n4485) );
  NBUFFX2 U4724 ( .INP(n4675), .Z(n4486) );
  NBUFFX2 U4725 ( .INP(n4674), .Z(n4487) );
  NBUFFX2 U4726 ( .INP(n4674), .Z(n4488) );
  NBUFFX2 U4727 ( .INP(n4674), .Z(n4489) );
  NBUFFX2 U4728 ( .INP(n4673), .Z(n4490) );
  NBUFFX2 U4729 ( .INP(n4673), .Z(n4491) );
  NBUFFX2 U4730 ( .INP(n4673), .Z(n4492) );
  NBUFFX2 U4731 ( .INP(n4672), .Z(n4493) );
  NBUFFX2 U4732 ( .INP(n4672), .Z(n4494) );
  NBUFFX2 U4733 ( .INP(n4672), .Z(n4495) );
  NBUFFX2 U4734 ( .INP(n4671), .Z(n4496) );
  NBUFFX2 U4735 ( .INP(n4671), .Z(n4497) );
  NBUFFX2 U4736 ( .INP(n4671), .Z(n4498) );
  NBUFFX2 U4737 ( .INP(n4670), .Z(n4499) );
  NBUFFX2 U4738 ( .INP(n4670), .Z(n4500) );
  NBUFFX2 U4739 ( .INP(n4670), .Z(n4501) );
  NBUFFX2 U4740 ( .INP(n4669), .Z(n4502) );
  NBUFFX2 U4741 ( .INP(n4669), .Z(n4503) );
  NBUFFX2 U4742 ( .INP(n4669), .Z(n4504) );
  NBUFFX2 U4743 ( .INP(n4668), .Z(n4505) );
  NBUFFX2 U4744 ( .INP(n4668), .Z(n4506) );
  NBUFFX2 U4745 ( .INP(n4668), .Z(n4507) );
  NBUFFX2 U4746 ( .INP(n4667), .Z(n4508) );
  NBUFFX2 U4747 ( .INP(n4667), .Z(n4509) );
  NBUFFX2 U4748 ( .INP(n4667), .Z(n4510) );
  NBUFFX2 U4749 ( .INP(n4666), .Z(n4511) );
  NBUFFX2 U4750 ( .INP(n4666), .Z(n4512) );
  NBUFFX2 U4751 ( .INP(n4666), .Z(n4513) );
  NBUFFX2 U4752 ( .INP(n4665), .Z(n4514) );
  NBUFFX2 U4753 ( .INP(n4665), .Z(n4515) );
  NBUFFX2 U4754 ( .INP(n4665), .Z(n4516) );
  NBUFFX2 U4755 ( .INP(n4664), .Z(n4517) );
  NBUFFX2 U4756 ( .INP(n4664), .Z(n4518) );
  NBUFFX2 U4757 ( .INP(n4664), .Z(n4519) );
  NBUFFX2 U4758 ( .INP(n4663), .Z(n4520) );
  NBUFFX2 U4759 ( .INP(n4663), .Z(n4521) );
  NBUFFX2 U4760 ( .INP(n4663), .Z(n4522) );
  NBUFFX2 U4761 ( .INP(n4662), .Z(n4523) );
  NBUFFX2 U4762 ( .INP(n4662), .Z(n4524) );
  NBUFFX2 U4763 ( .INP(n4662), .Z(n4525) );
  NBUFFX2 U4764 ( .INP(n4661), .Z(n4526) );
  NBUFFX2 U4765 ( .INP(n4661), .Z(n4527) );
  NBUFFX2 U4766 ( .INP(n4661), .Z(n4528) );
  NBUFFX2 U4767 ( .INP(n4660), .Z(n4529) );
  NBUFFX2 U4768 ( .INP(n4660), .Z(n4530) );
  NBUFFX2 U4769 ( .INP(n4660), .Z(n4531) );
  NBUFFX2 U4770 ( .INP(n4659), .Z(n4532) );
  NBUFFX2 U4771 ( .INP(n4659), .Z(n4533) );
  NBUFFX2 U4772 ( .INP(n4659), .Z(n4534) );
  NBUFFX2 U4773 ( .INP(n4658), .Z(n4535) );
  NBUFFX2 U4774 ( .INP(n4658), .Z(n4536) );
  NBUFFX2 U4775 ( .INP(n4658), .Z(n4537) );
  NBUFFX2 U4776 ( .INP(n4657), .Z(n4538) );
  NBUFFX2 U4777 ( .INP(n4657), .Z(n4539) );
  NBUFFX2 U4778 ( .INP(n4657), .Z(n4540) );
  NBUFFX2 U4779 ( .INP(n4656), .Z(n4541) );
  NBUFFX2 U4780 ( .INP(n4656), .Z(n4542) );
  NBUFFX2 U4781 ( .INP(n4656), .Z(n4543) );
  NBUFFX2 U4782 ( .INP(n4655), .Z(n4544) );
  NBUFFX2 U4783 ( .INP(n4655), .Z(n4545) );
  NBUFFX2 U4784 ( .INP(n4655), .Z(n4546) );
  NBUFFX2 U4785 ( .INP(n4654), .Z(n4547) );
  NBUFFX2 U4786 ( .INP(n4654), .Z(n4548) );
  NBUFFX2 U4787 ( .INP(n4654), .Z(n4549) );
  NBUFFX2 U4788 ( .INP(n4653), .Z(n4550) );
  NBUFFX2 U4789 ( .INP(n4653), .Z(n4551) );
  NBUFFX2 U4790 ( .INP(n4653), .Z(n4552) );
  NBUFFX2 U4791 ( .INP(n4652), .Z(n4553) );
  NBUFFX2 U4792 ( .INP(n4652), .Z(n4554) );
  NBUFFX2 U4793 ( .INP(n4652), .Z(n4555) );
  NBUFFX2 U4794 ( .INP(n4651), .Z(n4556) );
  NBUFFX2 U4795 ( .INP(n4651), .Z(n4557) );
  NBUFFX2 U4796 ( .INP(n4651), .Z(n4558) );
  NBUFFX2 U4797 ( .INP(n4650), .Z(n4559) );
  NBUFFX2 U4798 ( .INP(n4650), .Z(n4560) );
  NBUFFX2 U4799 ( .INP(n4650), .Z(n4561) );
  NBUFFX2 U4800 ( .INP(n4649), .Z(n4562) );
  NBUFFX2 U4801 ( .INP(n4649), .Z(n4563) );
  NBUFFX2 U4802 ( .INP(n4649), .Z(n4564) );
  NBUFFX2 U4803 ( .INP(n4648), .Z(n4565) );
  NBUFFX2 U4804 ( .INP(n4648), .Z(n4566) );
  NBUFFX2 U4805 ( .INP(n4648), .Z(n4567) );
  NBUFFX2 U4806 ( .INP(n4647), .Z(n4568) );
  NBUFFX2 U4807 ( .INP(n4647), .Z(n4569) );
  NBUFFX2 U4808 ( .INP(n4647), .Z(n4570) );
  NBUFFX2 U4809 ( .INP(n4646), .Z(n4571) );
  NBUFFX2 U4810 ( .INP(n4646), .Z(n4572) );
  NBUFFX2 U4811 ( .INP(n4646), .Z(n4573) );
  NBUFFX2 U4812 ( .INP(n4645), .Z(n4574) );
  NBUFFX2 U4813 ( .INP(n4645), .Z(n4575) );
  NBUFFX2 U4814 ( .INP(n4645), .Z(n4576) );
  NBUFFX2 U4815 ( .INP(n4644), .Z(n4577) );
  NBUFFX2 U4816 ( .INP(n4644), .Z(n4578) );
  NBUFFX2 U4817 ( .INP(n4644), .Z(n4579) );
  NBUFFX2 U4818 ( .INP(n4643), .Z(n4580) );
  NBUFFX2 U4819 ( .INP(n4643), .Z(n4581) );
  NBUFFX2 U4820 ( .INP(n4643), .Z(n4582) );
  NBUFFX2 U4821 ( .INP(n4642), .Z(n4583) );
  NBUFFX2 U4822 ( .INP(n4642), .Z(n4584) );
  NBUFFX2 U4823 ( .INP(n4642), .Z(n4585) );
  NBUFFX2 U4824 ( .INP(n4641), .Z(n4586) );
  NBUFFX2 U4825 ( .INP(n4641), .Z(n4587) );
  NBUFFX2 U4826 ( .INP(n4641), .Z(n4588) );
  NBUFFX2 U4827 ( .INP(n4640), .Z(n4589) );
  NBUFFX2 U4828 ( .INP(n4640), .Z(n4590) );
  NBUFFX2 U4829 ( .INP(n4640), .Z(n4591) );
  NBUFFX2 U4830 ( .INP(n4639), .Z(n4592) );
  NBUFFX2 U4831 ( .INP(n4639), .Z(n4593) );
  NBUFFX2 U4832 ( .INP(n4639), .Z(n4594) );
  NBUFFX2 U4833 ( .INP(n4638), .Z(n4595) );
  NBUFFX2 U4834 ( .INP(n4638), .Z(n4596) );
  NBUFFX2 U4835 ( .INP(n4638), .Z(n4597) );
  NBUFFX2 U4836 ( .INP(n4637), .Z(n4598) );
  NBUFFX2 U4837 ( .INP(n4637), .Z(n4599) );
  NBUFFX2 U4838 ( .INP(n4637), .Z(n4600) );
  NBUFFX2 U4839 ( .INP(n4636), .Z(n4601) );
  NBUFFX2 U4840 ( .INP(n4636), .Z(n4602) );
  NBUFFX2 U4841 ( .INP(n4636), .Z(n4603) );
  NBUFFX2 U4842 ( .INP(n4635), .Z(n4604) );
  NBUFFX2 U4843 ( .INP(n4635), .Z(n4605) );
  NBUFFX2 U4844 ( .INP(n4635), .Z(n4606) );
  NBUFFX2 U4845 ( .INP(n4634), .Z(n4607) );
  NBUFFX2 U4846 ( .INP(n4634), .Z(n4608) );
  NBUFFX2 U4847 ( .INP(n4634), .Z(n4609) );
  NBUFFX2 U4848 ( .INP(n4633), .Z(n4610) );
  NBUFFX2 U4849 ( .INP(n4633), .Z(n4611) );
  NBUFFX2 U4850 ( .INP(n4633), .Z(n4612) );
  NBUFFX2 U4851 ( .INP(n4632), .Z(n4613) );
  NBUFFX2 U4852 ( .INP(n4632), .Z(n4614) );
  NBUFFX2 U4853 ( .INP(n4632), .Z(n4615) );
  NBUFFX2 U4854 ( .INP(n4631), .Z(n4616) );
  NBUFFX2 U4855 ( .INP(n4631), .Z(n4617) );
  NBUFFX2 U4856 ( .INP(n4631), .Z(n4618) );
  NBUFFX2 U4857 ( .INP(n4630), .Z(n4619) );
  NBUFFX2 U4858 ( .INP(n4630), .Z(n4620) );
  NBUFFX2 U4859 ( .INP(n4630), .Z(n4621) );
  NBUFFX2 U4860 ( .INP(n4629), .Z(n4622) );
  NBUFFX2 U4861 ( .INP(n4629), .Z(n4623) );
  NBUFFX2 U4862 ( .INP(n4629), .Z(n4624) );
  NBUFFX2 U4863 ( .INP(n4628), .Z(n4625) );
  NBUFFX2 U4864 ( .INP(n4628), .Z(n4626) );
  NBUFFX2 U4865 ( .INP(n4628), .Z(n4627) );
  NBUFFX2 U4866 ( .INP(n4755), .Z(n4628) );
  NBUFFX2 U4867 ( .INP(n4755), .Z(n4629) );
  NBUFFX2 U4868 ( .INP(n4755), .Z(n4630) );
  NBUFFX2 U4869 ( .INP(n4754), .Z(n4631) );
  NBUFFX2 U4870 ( .INP(n4754), .Z(n4632) );
  NBUFFX2 U4871 ( .INP(n4754), .Z(n4633) );
  NBUFFX2 U4872 ( .INP(n4753), .Z(n4634) );
  NBUFFX2 U4873 ( .INP(n4753), .Z(n4635) );
  NBUFFX2 U4874 ( .INP(n4753), .Z(n4636) );
  NBUFFX2 U4875 ( .INP(n4752), .Z(n4637) );
  NBUFFX2 U4876 ( .INP(n4752), .Z(n4638) );
  NBUFFX2 U4877 ( .INP(n4752), .Z(n4639) );
  NBUFFX2 U4878 ( .INP(n4751), .Z(n4640) );
  NBUFFX2 U4879 ( .INP(n4751), .Z(n4641) );
  NBUFFX2 U4880 ( .INP(n4751), .Z(n4642) );
  NBUFFX2 U4881 ( .INP(n4750), .Z(n4643) );
  NBUFFX2 U4882 ( .INP(n4750), .Z(n4644) );
  NBUFFX2 U4883 ( .INP(n4750), .Z(n4645) );
  NBUFFX2 U4884 ( .INP(n4749), .Z(n4646) );
  NBUFFX2 U4885 ( .INP(n4749), .Z(n4647) );
  NBUFFX2 U4886 ( .INP(n4749), .Z(n4648) );
  NBUFFX2 U4887 ( .INP(n4748), .Z(n4649) );
  NBUFFX2 U4888 ( .INP(n4748), .Z(n4650) );
  NBUFFX2 U4889 ( .INP(n4748), .Z(n4651) );
  NBUFFX2 U4890 ( .INP(n4747), .Z(n4652) );
  NBUFFX2 U4891 ( .INP(n4747), .Z(n4653) );
  NBUFFX2 U4892 ( .INP(n4747), .Z(n4654) );
  NBUFFX2 U4893 ( .INP(n4746), .Z(n4655) );
  NBUFFX2 U4894 ( .INP(n4746), .Z(n4656) );
  NBUFFX2 U4895 ( .INP(n4746), .Z(n4657) );
  NBUFFX2 U4896 ( .INP(n4745), .Z(n4658) );
  NBUFFX2 U4897 ( .INP(n4745), .Z(n4659) );
  NBUFFX2 U4898 ( .INP(n4745), .Z(n4660) );
  NBUFFX2 U4899 ( .INP(n4744), .Z(n4661) );
  NBUFFX2 U4900 ( .INP(n4744), .Z(n4662) );
  NBUFFX2 U4901 ( .INP(n4744), .Z(n4663) );
  NBUFFX2 U4902 ( .INP(n4743), .Z(n4664) );
  NBUFFX2 U4903 ( .INP(n4743), .Z(n4665) );
  NBUFFX2 U4904 ( .INP(n4743), .Z(n4666) );
  NBUFFX2 U4905 ( .INP(n4742), .Z(n4667) );
  NBUFFX2 U4906 ( .INP(n4742), .Z(n4668) );
  NBUFFX2 U4907 ( .INP(n4742), .Z(n4669) );
  NBUFFX2 U4908 ( .INP(n4741), .Z(n4670) );
  NBUFFX2 U4909 ( .INP(n4741), .Z(n4671) );
  NBUFFX2 U4910 ( .INP(n4741), .Z(n4672) );
  NBUFFX2 U4911 ( .INP(n4740), .Z(n4673) );
  NBUFFX2 U4912 ( .INP(n4740), .Z(n4674) );
  NBUFFX2 U4913 ( .INP(n4740), .Z(n4675) );
  NBUFFX2 U4914 ( .INP(n4739), .Z(n4676) );
  NBUFFX2 U4915 ( .INP(n4739), .Z(n4677) );
  NBUFFX2 U4916 ( .INP(n4739), .Z(n4678) );
  NBUFFX2 U4917 ( .INP(n4738), .Z(n4679) );
  NBUFFX2 U4918 ( .INP(n4738), .Z(n4680) );
  NBUFFX2 U4919 ( .INP(n4738), .Z(n4681) );
  NBUFFX2 U4920 ( .INP(n4737), .Z(n4682) );
  NBUFFX2 U4921 ( .INP(n4737), .Z(n4683) );
  NBUFFX2 U4922 ( .INP(n4737), .Z(n4684) );
  NBUFFX2 U4923 ( .INP(n4736), .Z(n4685) );
  NBUFFX2 U4924 ( .INP(n4736), .Z(n4686) );
  NBUFFX2 U4925 ( .INP(n4736), .Z(n4687) );
  NBUFFX2 U4926 ( .INP(n4735), .Z(n4688) );
  NBUFFX2 U4927 ( .INP(n4735), .Z(n4689) );
  NBUFFX2 U4928 ( .INP(n4735), .Z(n4690) );
  NBUFFX2 U4929 ( .INP(n4734), .Z(n4691) );
  NBUFFX2 U4930 ( .INP(n4734), .Z(n4692) );
  NBUFFX2 U4931 ( .INP(n4734), .Z(n4693) );
  NBUFFX2 U4932 ( .INP(n4733), .Z(n4694) );
  NBUFFX2 U4933 ( .INP(n4733), .Z(n4695) );
  NBUFFX2 U4934 ( .INP(n4733), .Z(n4696) );
  NBUFFX2 U4935 ( .INP(n4732), .Z(n4697) );
  NBUFFX2 U4936 ( .INP(n4732), .Z(n4698) );
  NBUFFX2 U4937 ( .INP(n4732), .Z(n4699) );
  NBUFFX2 U4938 ( .INP(n4731), .Z(n4700) );
  NBUFFX2 U4939 ( .INP(n4731), .Z(n4701) );
  NBUFFX2 U4940 ( .INP(n4731), .Z(n4702) );
  NBUFFX2 U4941 ( .INP(n4730), .Z(n4703) );
  NBUFFX2 U4942 ( .INP(n4730), .Z(n4704) );
  NBUFFX2 U4943 ( .INP(n4730), .Z(n4705) );
  NBUFFX2 U4944 ( .INP(n4729), .Z(n4706) );
  NBUFFX2 U4945 ( .INP(n4729), .Z(n4707) );
  NBUFFX2 U4946 ( .INP(n4729), .Z(n4708) );
  NBUFFX2 U4947 ( .INP(n4728), .Z(n4709) );
  NBUFFX2 U4948 ( .INP(n4728), .Z(n4710) );
  NBUFFX2 U4949 ( .INP(n4728), .Z(n4711) );
  NBUFFX2 U4950 ( .INP(n4727), .Z(n4712) );
  NBUFFX2 U4951 ( .INP(n4727), .Z(n4713) );
  NBUFFX2 U4952 ( .INP(n4727), .Z(n4714) );
  NBUFFX2 U4953 ( .INP(n4726), .Z(n4715) );
  NBUFFX2 U4954 ( .INP(n4726), .Z(n4716) );
  NBUFFX2 U4955 ( .INP(n4726), .Z(n4717) );
  NBUFFX2 U4956 ( .INP(n4725), .Z(n4718) );
  NBUFFX2 U4957 ( .INP(n4725), .Z(n4719) );
  NBUFFX2 U4958 ( .INP(n4725), .Z(n4720) );
  NBUFFX2 U4959 ( .INP(n4724), .Z(n4721) );
  NBUFFX2 U4960 ( .INP(n4724), .Z(n4722) );
  NBUFFX2 U4961 ( .INP(n4724), .Z(n4723) );
  NBUFFX2 U4962 ( .INP(n4766), .Z(n4724) );
  NBUFFX2 U4963 ( .INP(n4766), .Z(n4725) );
  NBUFFX2 U4964 ( .INP(n4765), .Z(n4726) );
  NBUFFX2 U4965 ( .INP(n4765), .Z(n4727) );
  NBUFFX2 U4966 ( .INP(n4765), .Z(n4728) );
  NBUFFX2 U4967 ( .INP(n4764), .Z(n4729) );
  NBUFFX2 U4968 ( .INP(n4764), .Z(n4730) );
  NBUFFX2 U4969 ( .INP(n4764), .Z(n4731) );
  NBUFFX2 U4970 ( .INP(n4763), .Z(n4732) );
  NBUFFX2 U4971 ( .INP(n4763), .Z(n4733) );
  NBUFFX2 U4972 ( .INP(n4763), .Z(n4734) );
  NBUFFX2 U4973 ( .INP(n4762), .Z(n4735) );
  NBUFFX2 U4974 ( .INP(n4762), .Z(n4736) );
  NBUFFX2 U4975 ( .INP(n4762), .Z(n4737) );
  NBUFFX2 U4976 ( .INP(n4761), .Z(n4738) );
  NBUFFX2 U4977 ( .INP(n4761), .Z(n4739) );
  NBUFFX2 U4978 ( .INP(n4761), .Z(n4740) );
  NBUFFX2 U4979 ( .INP(n4760), .Z(n4741) );
  NBUFFX2 U4980 ( .INP(n4760), .Z(n4742) );
  NBUFFX2 U4981 ( .INP(n4760), .Z(n4743) );
  NBUFFX2 U4982 ( .INP(n4759), .Z(n4744) );
  NBUFFX2 U4983 ( .INP(n4759), .Z(n4745) );
  NBUFFX2 U4984 ( .INP(n4759), .Z(n4746) );
  NBUFFX2 U4985 ( .INP(n4758), .Z(n4747) );
  NBUFFX2 U4986 ( .INP(n4758), .Z(n4748) );
  NBUFFX2 U4987 ( .INP(n4758), .Z(n4749) );
  NBUFFX2 U4988 ( .INP(n4757), .Z(n4750) );
  NBUFFX2 U4989 ( .INP(n4757), .Z(n4751) );
  NBUFFX2 U4990 ( .INP(n4757), .Z(n4752) );
  NBUFFX2 U4991 ( .INP(n4756), .Z(n4753) );
  NBUFFX2 U4992 ( .INP(n4756), .Z(n4754) );
  NBUFFX2 U4993 ( .INP(n4756), .Z(n4755) );
  NBUFFX2 U4994 ( .INP(n4770), .Z(n4756) );
  NBUFFX2 U4995 ( .INP(n4770), .Z(n4757) );
  NBUFFX2 U4996 ( .INP(n4769), .Z(n4758) );
  NBUFFX2 U4997 ( .INP(n4769), .Z(n4759) );
  NBUFFX2 U4998 ( .INP(n4769), .Z(n4760) );
  NBUFFX2 U4999 ( .INP(n4768), .Z(n4761) );
  NBUFFX2 U5000 ( .INP(n4768), .Z(n4762) );
  NBUFFX2 U5001 ( .INP(n4768), .Z(n4763) );
  NBUFFX2 U5002 ( .INP(n4767), .Z(n4764) );
  NBUFFX2 U5003 ( .INP(n4767), .Z(n4765) );
  NBUFFX2 U5004 ( .INP(n4767), .Z(n4766) );
  NBUFFX2 U5005 ( .INP(test_se), .Z(n4767) );
  NBUFFX2 U5006 ( .INP(test_se), .Z(n4768) );
  NBUFFX2 U5007 ( .INP(test_se), .Z(n4769) );
  NBUFFX2 U5008 ( .INP(test_se), .Z(n4770) );
  NBUFFX2 U5009 ( .INP(TM1), .Z(n4784) );
  NBUFFX2 U5010 ( .INP(TM1), .Z(n4785) );
  NBUFFX2 U5011 ( .INP(TM1), .Z(n4786) );
  NBUFFX2 U5012 ( .INP(n4842), .Z(n4787) );
  NBUFFX2 U5013 ( .INP(n4842), .Z(n4788) );
  NBUFFX2 U5014 ( .INP(n4842), .Z(n4789) );
  NBUFFX2 U5015 ( .INP(n4841), .Z(n4790) );
  NBUFFX2 U5016 ( .INP(n4841), .Z(n4791) );
  NBUFFX2 U5017 ( .INP(n4841), .Z(n4792) );
  NBUFFX2 U5018 ( .INP(n4840), .Z(n4793) );
  NBUFFX2 U5019 ( .INP(n4840), .Z(n4794) );
  NBUFFX2 U5020 ( .INP(n4840), .Z(n4795) );
  NBUFFX2 U5021 ( .INP(n4839), .Z(n4796) );
  NBUFFX2 U5022 ( .INP(n4839), .Z(n4797) );
  NBUFFX2 U5023 ( .INP(n4839), .Z(n4798) );
  NBUFFX2 U5024 ( .INP(n4838), .Z(n4799) );
  NBUFFX2 U5025 ( .INP(n4838), .Z(n4800) );
  NBUFFX2 U5026 ( .INP(n4838), .Z(n4801) );
  NBUFFX2 U5027 ( .INP(n4837), .Z(n4802) );
  NBUFFX2 U5028 ( .INP(n4837), .Z(n4803) );
  NBUFFX2 U5029 ( .INP(n4837), .Z(n4804) );
  NBUFFX2 U5030 ( .INP(n4836), .Z(n4805) );
  NBUFFX2 U5031 ( .INP(n4836), .Z(n4806) );
  NBUFFX2 U5032 ( .INP(n4836), .Z(n4807) );
  NBUFFX2 U5033 ( .INP(n4835), .Z(n4808) );
  NBUFFX2 U5034 ( .INP(n4835), .Z(n4809) );
  NBUFFX2 U5035 ( .INP(n4835), .Z(n4810) );
  NBUFFX2 U5036 ( .INP(n4834), .Z(n4811) );
  NBUFFX2 U5037 ( .INP(n4834), .Z(n4812) );
  NBUFFX2 U5038 ( .INP(n4834), .Z(n4813) );
  NBUFFX2 U5039 ( .INP(n4833), .Z(n4814) );
  NBUFFX2 U5040 ( .INP(n4833), .Z(n4815) );
  NBUFFX2 U5041 ( .INP(n4833), .Z(n4816) );
  NBUFFX2 U5042 ( .INP(n4832), .Z(n4817) );
  NBUFFX2 U5043 ( .INP(n4832), .Z(n4818) );
  NBUFFX2 U5044 ( .INP(n4832), .Z(n4819) );
  NBUFFX2 U5045 ( .INP(n4831), .Z(n4820) );
  NBUFFX2 U5046 ( .INP(n4831), .Z(n4821) );
  NBUFFX2 U5047 ( .INP(n4831), .Z(n4822) );
  NBUFFX2 U5048 ( .INP(n4830), .Z(n4823) );
  NBUFFX2 U5049 ( .INP(n4830), .Z(n4824) );
  NBUFFX2 U5050 ( .INP(n4830), .Z(n4825) );
  NBUFFX2 U5051 ( .INP(n4829), .Z(n4826) );
  NBUFFX2 U5052 ( .INP(n4829), .Z(n4827) );
  NBUFFX2 U5053 ( .INP(n4829), .Z(n4828) );
  NBUFFX2 U5054 ( .INP(n4847), .Z(n4829) );
  NBUFFX2 U5055 ( .INP(n4847), .Z(n4830) );
  NBUFFX2 U5056 ( .INP(n4846), .Z(n4831) );
  NBUFFX2 U5057 ( .INP(n4846), .Z(n4832) );
  NBUFFX2 U5058 ( .INP(n4846), .Z(n4833) );
  NBUFFX2 U5059 ( .INP(n4845), .Z(n4834) );
  NBUFFX2 U5060 ( .INP(n4845), .Z(n4835) );
  NBUFFX2 U5061 ( .INP(n4845), .Z(n4836) );
  NBUFFX2 U5062 ( .INP(n4844), .Z(n4837) );
  NBUFFX2 U5063 ( .INP(n4844), .Z(n4838) );
  NBUFFX2 U5064 ( .INP(n4844), .Z(n4839) );
  NBUFFX2 U5065 ( .INP(n4843), .Z(n4840) );
  NBUFFX2 U5066 ( .INP(n4843), .Z(n4841) );
  NBUFFX2 U5067 ( .INP(n4843), .Z(n4842) );
  NBUFFX2 U5068 ( .INP(RESET), .Z(n4843) );
  NBUFFX2 U5069 ( .INP(RESET), .Z(n4844) );
  NBUFFX2 U5070 ( .INP(RESET), .Z(n4845) );
  NBUFFX2 U5071 ( .INP(RESET), .Z(n4846) );
  NBUFFX2 U5072 ( .INP(RESET), .Z(n4847) );
  INVX0 U5073 ( .INP(n4799), .ZN(n4848) );
  INVX0 U5074 ( .INP(n4799), .ZN(n4849) );
  INVX0 U5075 ( .INP(n4799), .ZN(n4850) );
  INVX0 U5076 ( .INP(n4799), .ZN(n4851) );
  INVX0 U5077 ( .INP(n4799), .ZN(n4852) );
  INVX0 U5078 ( .INP(n4799), .ZN(n4853) );
  INVX0 U5079 ( .INP(n4799), .ZN(n4854) );
  INVX0 U5080 ( .INP(n4798), .ZN(n4855) );
  INVX0 U5081 ( .INP(n4798), .ZN(n4856) );
  INVX0 U5082 ( .INP(n4798), .ZN(n4857) );
  INVX0 U5083 ( .INP(n4798), .ZN(n4858) );
  INVX0 U5084 ( .INP(n4797), .ZN(n4859) );
  INVX0 U5085 ( .INP(n4797), .ZN(n4860) );
  INVX0 U5086 ( .INP(n4797), .ZN(n4861) );
  INVX0 U5087 ( .INP(n4797), .ZN(n4862) );
  INVX0 U5088 ( .INP(n4797), .ZN(n4863) );
  INVX0 U5089 ( .INP(n4797), .ZN(n4864) );
  INVX0 U5090 ( .INP(n4797), .ZN(n4865) );
  INVX0 U5091 ( .INP(n4797), .ZN(n4866) );
  INVX0 U5092 ( .INP(n4796), .ZN(n4867) );
  INVX0 U5093 ( .INP(n4796), .ZN(n4868) );
  INVX0 U5094 ( .INP(n4792), .ZN(n4869) );
  INVX0 U5095 ( .INP(n4792), .ZN(n4870) );
  INVX0 U5096 ( .INP(n4788), .ZN(n4871) );
  INVX0 U5097 ( .INP(n4788), .ZN(n4872) );
  INVX0 U5098 ( .INP(n4794), .ZN(n4873) );
  INVX0 U5099 ( .INP(n4787), .ZN(n4874) );
  INVX0 U5100 ( .INP(n4787), .ZN(n4875) );
  INVX0 U5101 ( .INP(n4787), .ZN(n4876) );
  INVX0 U5102 ( .INP(n4787), .ZN(n4877) );
  INVX0 U5103 ( .INP(n4787), .ZN(n4878) );
  INVX0 U5104 ( .INP(n4787), .ZN(n4879) );
  INVX0 U5105 ( .INP(n4787), .ZN(n4880) );
  INVX0 U5106 ( .INP(n4787), .ZN(n4881) );
  INVX0 U5107 ( .INP(n4788), .ZN(n4882) );
  INVX0 U5108 ( .INP(n4788), .ZN(n4883) );
  INVX0 U5109 ( .INP(n4788), .ZN(n4884) );
  INVX0 U5110 ( .INP(n4788), .ZN(n4885) );
  INVX0 U5111 ( .INP(n4788), .ZN(n4886) );
  INVX0 U5112 ( .INP(n4788), .ZN(n4887) );
  INVX0 U5113 ( .INP(n4789), .ZN(n4888) );
  INVX0 U5114 ( .INP(n4789), .ZN(n4889) );
  INVX0 U5115 ( .INP(n4789), .ZN(n4890) );
  INVX0 U5116 ( .INP(n4789), .ZN(n4891) );
  INVX0 U5117 ( .INP(n4789), .ZN(n4892) );
  INVX0 U5118 ( .INP(n4789), .ZN(n4893) );
  INVX0 U5119 ( .INP(n4789), .ZN(n4894) );
  INVX0 U5120 ( .INP(n4790), .ZN(n4895) );
  INVX0 U5121 ( .INP(n4790), .ZN(n4896) );
  INVX0 U5122 ( .INP(n4790), .ZN(n4897) );
  INVX0 U5123 ( .INP(n4790), .ZN(n4898) );
  INVX0 U5124 ( .INP(n4790), .ZN(n4899) );
  INVX0 U5125 ( .INP(n4790), .ZN(n4900) );
  INVX0 U5126 ( .INP(n4790), .ZN(n4901) );
  INVX0 U5127 ( .INP(n4790), .ZN(n4902) );
  INVX0 U5128 ( .INP(n4791), .ZN(n4903) );
  INVX0 U5129 ( .INP(n4791), .ZN(n4904) );
  INVX0 U5130 ( .INP(n4791), .ZN(n4905) );
  INVX0 U5131 ( .INP(n4791), .ZN(n4906) );
  INVX0 U5132 ( .INP(n4791), .ZN(n4907) );
  INVX0 U5133 ( .INP(n4791), .ZN(n4908) );
  INVX0 U5134 ( .INP(n4791), .ZN(n4909) );
  INVX0 U5135 ( .INP(n4791), .ZN(n4910) );
  INVX0 U5136 ( .INP(n4792), .ZN(n4911) );
  INVX0 U5137 ( .INP(n4792), .ZN(n4912) );
  INVX0 U5138 ( .INP(n4792), .ZN(n4913) );
  INVX0 U5139 ( .INP(n4792), .ZN(n4914) );
  INVX0 U5140 ( .INP(n4792), .ZN(n4915) );
  INVX0 U5141 ( .INP(n4792), .ZN(n4916) );
  INVX0 U5142 ( .INP(n4793), .ZN(n4917) );
  INVX0 U5143 ( .INP(n4793), .ZN(n4918) );
  INVX0 U5144 ( .INP(n4793), .ZN(n4919) );
  INVX0 U5145 ( .INP(n4793), .ZN(n4920) );
  INVX0 U5146 ( .INP(n4793), .ZN(n4921) );
  INVX0 U5147 ( .INP(n4793), .ZN(n4922) );
  INVX0 U5148 ( .INP(n4793), .ZN(n4923) );
  INVX0 U5149 ( .INP(n4793), .ZN(n4924) );
  INVX0 U5150 ( .INP(n4794), .ZN(n4925) );
  INVX0 U5151 ( .INP(n4794), .ZN(n4926) );
  INVX0 U5152 ( .INP(n4794), .ZN(n4927) );
  INVX0 U5153 ( .INP(n4794), .ZN(n4928) );
  INVX0 U5154 ( .INP(n4794), .ZN(n4929) );
  INVX0 U5155 ( .INP(n4794), .ZN(n4930) );
  INVX0 U5156 ( .INP(n4794), .ZN(n4931) );
  INVX0 U5157 ( .INP(n4795), .ZN(n4932) );
  INVX0 U5158 ( .INP(n4795), .ZN(n4933) );
  INVX0 U5159 ( .INP(n4795), .ZN(n4934) );
  INVX0 U5160 ( .INP(n4795), .ZN(n4935) );
  INVX0 U5161 ( .INP(n4795), .ZN(n4936) );
  INVX0 U5162 ( .INP(n4795), .ZN(n4937) );
  INVX0 U5163 ( .INP(n4795), .ZN(n4938) );
  INVX0 U5164 ( .INP(n4795), .ZN(n4939) );
  INVX0 U5165 ( .INP(n4796), .ZN(n4940) );
  INVX0 U5166 ( .INP(n4796), .ZN(n4941) );
  INVX0 U5167 ( .INP(n4796), .ZN(n4942) );
  INVX0 U5168 ( .INP(n4796), .ZN(n4943) );
  INVX0 U5169 ( .INP(n4796), .ZN(n4944) );
  INVX0 U5170 ( .INP(n4796), .ZN(n4945) );
  NBUFFX2 U5171 ( .INP(n5128), .Z(n5090) );
  NBUFFX2 U5172 ( .INP(n5128), .Z(n5091) );
  NBUFFX2 U5173 ( .INP(n5127), .Z(n5092) );
  NBUFFX2 U5174 ( .INP(n5127), .Z(n5093) );
  NBUFFX2 U5175 ( .INP(n5127), .Z(n5094) );
  NBUFFX2 U5176 ( .INP(n5126), .Z(n5095) );
  NBUFFX2 U5177 ( .INP(n5126), .Z(n5096) );
  NBUFFX2 U5178 ( .INP(n5126), .Z(n5097) );
  NBUFFX2 U5179 ( .INP(n5125), .Z(n5098) );
  NBUFFX2 U5180 ( .INP(n5125), .Z(n5099) );
  NBUFFX2 U5181 ( .INP(n5125), .Z(n5100) );
  NBUFFX2 U5182 ( .INP(n5124), .Z(n5101) );
  NBUFFX2 U5183 ( .INP(n5124), .Z(n5102) );
  NBUFFX2 U5184 ( .INP(n5124), .Z(n5103) );
  NBUFFX2 U5185 ( .INP(n5123), .Z(n5104) );
  NBUFFX2 U5186 ( .INP(n5123), .Z(n5105) );
  NBUFFX2 U5187 ( .INP(n5123), .Z(n5106) );
  NBUFFX2 U5188 ( .INP(n5122), .Z(n5107) );
  NBUFFX2 U5189 ( .INP(n5122), .Z(n5108) );
  NBUFFX2 U5190 ( .INP(n5122), .Z(n5109) );
  NBUFFX2 U5191 ( .INP(n5121), .Z(n5110) );
  NBUFFX2 U5192 ( .INP(n5121), .Z(n5111) );
  NBUFFX2 U5193 ( .INP(n5121), .Z(n5112) );
  NBUFFX2 U5194 ( .INP(n5120), .Z(n5113) );
  NBUFFX2 U5195 ( .INP(n5120), .Z(n5114) );
  NBUFFX2 U5196 ( .INP(n5120), .Z(n5115) );
  NBUFFX2 U5197 ( .INP(n5119), .Z(n5116) );
  NBUFFX2 U5198 ( .INP(n5119), .Z(n5117) );
  NBUFFX2 U5199 ( .INP(n5119), .Z(n5118) );
  NBUFFX2 U5200 ( .INP(CK), .Z(n5119) );
  NBUFFX2 U5201 ( .INP(CK), .Z(n5120) );
  NBUFFX2 U5202 ( .INP(n5128), .Z(n5121) );
  NBUFFX2 U5203 ( .INP(CK), .Z(n5122) );
  NBUFFX2 U5204 ( .INP(n5124), .Z(n5123) );
  NBUFFX2 U5205 ( .INP(CK), .Z(n5124) );
  NBUFFX2 U5206 ( .INP(n5119), .Z(n5125) );
  NBUFFX2 U5207 ( .INP(n5120), .Z(n5126) );
  NBUFFX2 U5208 ( .INP(n5122), .Z(n5127) );
  NBUFFX2 U5209 ( .INP(n4959), .Z(n5128) );
  INVX0 U5210 ( .INP(n5129), .ZN(n99) );
  INVX0 U5211 ( .INP(n5130), .ZN(n98) );
  INVX0 U5212 ( .INP(n5131), .ZN(n97) );
  INVX0 U5213 ( .INP(n5132), .ZN(n96) );
  INVX0 U5214 ( .INP(n5133), .ZN(n95) );
  INVX0 U5215 ( .INP(n5134), .ZN(n94) );
  INVX0 U5216 ( .INP(n5135), .ZN(n93) );
  INVX0 U5217 ( .INP(n5136), .ZN(n92) );
  INVX0 U5218 ( .INP(n5137), .ZN(n91) );
  INVX0 U5219 ( .INP(n5138), .ZN(n90) );
  INVX0 U5220 ( .INP(n5139), .ZN(n9) );
  INVX0 U5221 ( .INP(n5140), .ZN(n89) );
  INVX0 U5222 ( .INP(n5141), .ZN(n88) );
  INVX0 U5223 ( .INP(n5142), .ZN(n87) );
  INVX0 U5224 ( .INP(n5143), .ZN(n86) );
  INVX0 U5225 ( .INP(n5144), .ZN(n85) );
  INVX0 U5226 ( .INP(n5145), .ZN(n84) );
  INVX0 U5227 ( .INP(n5146), .ZN(n83) );
  INVX0 U5228 ( .INP(n5147), .ZN(n82) );
  INVX0 U5229 ( .INP(n5148), .ZN(n81) );
  INVX0 U5230 ( .INP(n5149), .ZN(n80) );
  INVX0 U5231 ( .INP(n5150), .ZN(n8) );
  INVX0 U5232 ( .INP(n5151), .ZN(n79) );
  INVX0 U5233 ( .INP(n5152), .ZN(n78) );
  INVX0 U5234 ( .INP(n5153), .ZN(n77) );
  INVX0 U5235 ( .INP(n5154), .ZN(n76) );
  INVX0 U5236 ( .INP(n5155), .ZN(n75) );
  INVX0 U5237 ( .INP(n5156), .ZN(n74) );
  INVX0 U5238 ( .INP(n5157), .ZN(n73) );
  INVX0 U5239 ( .INP(n5158), .ZN(n72) );
  INVX0 U5240 ( .INP(n5159), .ZN(n71) );
  INVX0 U5241 ( .INP(n5160), .ZN(n70) );
  INVX0 U5242 ( .INP(n5161), .ZN(n7) );
  INVX0 U5243 ( .INP(n5162), .ZN(n69) );
  INVX0 U5244 ( .INP(n5163), .ZN(n68) );
  INVX0 U5245 ( .INP(n5164), .ZN(n67) );
  INVX0 U5246 ( .INP(n5165), .ZN(n66) );
  INVX0 U5247 ( .INP(n5166), .ZN(n65) );
  INVX0 U5248 ( .INP(n5167), .ZN(n64) );
  INVX0 U5249 ( .INP(n5168), .ZN(n63) );
  INVX0 U5250 ( .INP(n5169), .ZN(n62) );
  INVX0 U5251 ( .INP(n5170), .ZN(n61) );
  INVX0 U5252 ( .INP(n5171), .ZN(n60) );
  INVX0 U5253 ( .INP(n5172), .ZN(n6) );
  INVX0 U5254 ( .INP(n5173), .ZN(n59) );
  INVX0 U5255 ( .INP(n5174), .ZN(n58) );
  INVX0 U5256 ( .INP(n5175), .ZN(n57) );
  INVX0 U5257 ( .INP(n5176), .ZN(n56) );
  INVX0 U5258 ( .INP(n5177), .ZN(n55) );
  INVX0 U5259 ( .INP(n5178), .ZN(n54) );
  INVX0 U5260 ( .INP(n5179), .ZN(n53) );
  INVX0 U5261 ( .INP(n5180), .ZN(n52) );
  INVX0 U5262 ( .INP(n5181), .ZN(n51) );
  INVX0 U5263 ( .INP(n5182), .ZN(n50) );
  INVX0 U5264 ( .INP(n5183), .ZN(n5) );
  INVX0 U5265 ( .INP(n5184), .ZN(n49) );
  INVX0 U5266 ( .INP(n5185), .ZN(n48) );
  INVX0 U5267 ( .INP(n5186), .ZN(n47) );
  INVX0 U5268 ( .INP(n5187), .ZN(n46) );
  INVX0 U5269 ( .INP(n5188), .ZN(n45) );
  INVX0 U5270 ( .INP(n5189), .ZN(n44) );
  INVX0 U5271 ( .INP(n5190), .ZN(n43) );
  INVX0 U5272 ( .INP(n5191), .ZN(n42) );
  INVX0 U5273 ( .INP(n5192), .ZN(n41) );
  INVX0 U5274 ( .INP(n5193), .ZN(n40) );
  INVX0 U5275 ( .INP(n5194), .ZN(n4) );
  INVX0 U5276 ( .INP(n5195), .ZN(n39) );
  INVX0 U5277 ( .INP(n5196), .ZN(n38) );
  INVX0 U5278 ( .INP(n5197), .ZN(n37) );
  INVX0 U5279 ( .INP(n5198), .ZN(n36) );
  INVX0 U5280 ( .INP(n5199), .ZN(n35) );
  INVX0 U5281 ( .INP(n5200), .ZN(n34) );
  INVX0 U5282 ( .INP(n5201), .ZN(n33) );
  NOR2X0 U5283 ( .IN1(n4783), .IN2(n4848), .QN(n3278) );
  INVX0 U5284 ( .INP(n5202), .ZN(n32) );
  INVX0 U5285 ( .INP(n5203), .ZN(n31) );
  INVX0 U5286 ( .INP(n5204), .ZN(n30) );
  INVX0 U5287 ( .INP(n5205), .ZN(n3) );
  INVX0 U5288 ( .INP(n5206), .ZN(n29) );
  INVX0 U5289 ( .INP(n5207), .ZN(n28) );
  INVX0 U5290 ( .INP(n5208), .ZN(n27) );
  INVX0 U5291 ( .INP(n5209), .ZN(n26) );
  INVX0 U5292 ( .INP(n5210), .ZN(n25) );
  INVX0 U5293 ( .INP(n5211), .ZN(n24) );
  INVX0 U5294 ( .INP(n5212), .ZN(n23) );
  INVX0 U5295 ( .INP(TM0), .ZN(n225) );
  INVX0 U5296 ( .INP(n5213), .ZN(n22) );
  INVX0 U5297 ( .INP(n5214), .ZN(n218) );
  INVX0 U5298 ( .INP(n5215), .ZN(n217) );
  INVX0 U5299 ( .INP(n5216), .ZN(n216) );
  INVX0 U5300 ( .INP(n5217), .ZN(n215) );
  INVX0 U5301 ( .INP(n5218), .ZN(n214) );
  INVX0 U5302 ( .INP(n5219), .ZN(n213) );
  INVX0 U5303 ( .INP(n5220), .ZN(n212) );
  INVX0 U5304 ( .INP(n5221), .ZN(n211) );
  INVX0 U5305 ( .INP(n5222), .ZN(n210) );
  INVX0 U5306 ( .INP(n5223), .ZN(n21) );
  INVX0 U5307 ( .INP(n5224), .ZN(n209) );
  INVX0 U5308 ( .INP(n5225), .ZN(n208) );
  INVX0 U5309 ( .INP(n5226), .ZN(n207) );
  INVX0 U5310 ( .INP(n5227), .ZN(n206) );
  INVX0 U5311 ( .INP(n5228), .ZN(n205) );
  INVX0 U5312 ( .INP(n5229), .ZN(n204) );
  INVX0 U5313 ( .INP(n5230), .ZN(n203) );
  INVX0 U5314 ( .INP(n5231), .ZN(n202) );
  INVX0 U5315 ( .INP(n5232), .ZN(n201) );
  INVX0 U5316 ( .INP(n5233), .ZN(n200) );
  INVX0 U5317 ( .INP(n5234), .ZN(n20) );
  INVX0 U5318 ( .INP(n5235), .ZN(n2) );
  INVX0 U5319 ( .INP(n5236), .ZN(n199) );
  INVX0 U5320 ( .INP(n5237), .ZN(n198) );
  INVX0 U5321 ( .INP(n5238), .ZN(n197) );
  INVX0 U5322 ( .INP(n5239), .ZN(n196) );
  INVX0 U5323 ( .INP(n5240), .ZN(n195) );
  INVX0 U5324 ( .INP(n5241), .ZN(n194) );
  INVX0 U5325 ( .INP(n5242), .ZN(n193) );
  INVX0 U5326 ( .INP(n5243), .ZN(n192) );
  INVX0 U5327 ( .INP(n5244), .ZN(n191) );
  INVX0 U5328 ( .INP(n5245), .ZN(n190) );
  INVX0 U5329 ( .INP(n5246), .ZN(n19) );
  INVX0 U5330 ( .INP(n5247), .ZN(n189) );
  INVX0 U5331 ( .INP(n5248), .ZN(n188) );
  INVX0 U5332 ( .INP(n5249), .ZN(n187) );
  INVX0 U5333 ( .INP(n5250), .ZN(n186) );
  INVX0 U5334 ( .INP(n5251), .ZN(n185) );
  INVX0 U5335 ( .INP(n5252), .ZN(n184) );
  INVX0 U5336 ( .INP(n5253), .ZN(n183) );
  INVX0 U5337 ( .INP(n5254), .ZN(n182) );
  INVX0 U5338 ( .INP(n5255), .ZN(n181) );
  INVX0 U5339 ( .INP(n5256), .ZN(n180) );
  INVX0 U5340 ( .INP(n5257), .ZN(n18) );
  INVX0 U5341 ( .INP(n5258), .ZN(n179) );
  INVX0 U5342 ( .INP(n5259), .ZN(n178) );
  INVX0 U5343 ( .INP(n5260), .ZN(n177) );
  INVX0 U5344 ( .INP(n5261), .ZN(n176) );
  INVX0 U5345 ( .INP(n5262), .ZN(n175) );
  INVX0 U5346 ( .INP(n5263), .ZN(n174) );
  INVX0 U5347 ( .INP(n5264), .ZN(n173) );
  INVX0 U5348 ( .INP(n5265), .ZN(n172) );
  INVX0 U5349 ( .INP(n5266), .ZN(n171) );
  INVX0 U5350 ( .INP(n5267), .ZN(n170) );
  INVX0 U5351 ( .INP(n5268), .ZN(n17) );
  INVX0 U5352 ( .INP(n5269), .ZN(n169) );
  INVX0 U5353 ( .INP(n5270), .ZN(n168) );
  INVX0 U5354 ( .INP(n5271), .ZN(n167) );
  INVX0 U5355 ( .INP(n5272), .ZN(n166) );
  INVX0 U5356 ( .INP(n5273), .ZN(n165) );
  INVX0 U5357 ( .INP(n5274), .ZN(n164) );
  INVX0 U5358 ( .INP(n5275), .ZN(n163) );
  INVX0 U5359 ( .INP(n5276), .ZN(n162) );
  INVX0 U5360 ( .INP(n5277), .ZN(n161) );
  INVX0 U5361 ( .INP(n5278), .ZN(n160) );
  INVX0 U5362 ( .INP(n5279), .ZN(n16) );
  INVX0 U5363 ( .INP(n5280), .ZN(n159) );
  INVX0 U5364 ( .INP(n5281), .ZN(n158) );
  INVX0 U5365 ( .INP(n5282), .ZN(n157) );
  INVX0 U5366 ( .INP(n5283), .ZN(n156) );
  INVX0 U5367 ( .INP(n5284), .ZN(n155) );
  INVX0 U5368 ( .INP(n5285), .ZN(n154) );
  INVX0 U5369 ( .INP(n5286), .ZN(n153) );
  INVX0 U5370 ( .INP(n5287), .ZN(n152) );
  INVX0 U5371 ( .INP(n5288), .ZN(n151) );
  INVX0 U5372 ( .INP(n5289), .ZN(n150) );
  INVX0 U5373 ( .INP(n5290), .ZN(n15) );
  INVX0 U5374 ( .INP(n5291), .ZN(n149) );
  INVX0 U5375 ( .INP(n5292), .ZN(n148) );
  INVX0 U5376 ( .INP(n5293), .ZN(n147) );
  INVX0 U5377 ( .INP(n5294), .ZN(n146) );
  INVX0 U5378 ( .INP(n5295), .ZN(n145) );
  INVX0 U5379 ( .INP(n5296), .ZN(n144) );
  INVX0 U5380 ( .INP(n5297), .ZN(n143) );
  INVX0 U5381 ( .INP(n5298), .ZN(n142) );
  INVX0 U5382 ( .INP(n5299), .ZN(n141) );
  INVX0 U5383 ( .INP(n5300), .ZN(n140) );
  INVX0 U5384 ( .INP(n5301), .ZN(n14) );
  INVX0 U5385 ( .INP(n5302), .ZN(n139) );
  INVX0 U5386 ( .INP(n5303), .ZN(n138) );
  INVX0 U5387 ( .INP(n5304), .ZN(n137) );
  INVX0 U5388 ( .INP(n5305), .ZN(n136) );
  INVX0 U5389 ( .INP(n5306), .ZN(n135) );
  INVX0 U5390 ( .INP(n5307), .ZN(n134) );
  INVX0 U5391 ( .INP(n5308), .ZN(n133) );
  INVX0 U5392 ( .INP(n5309), .ZN(n132) );
  INVX0 U5393 ( .INP(n5310), .ZN(n131) );
  INVX0 U5394 ( .INP(n5311), .ZN(n130) );
  INVX0 U5395 ( .INP(n5312), .ZN(n13) );
  INVX0 U5396 ( .INP(n5313), .ZN(n129) );
  INVX0 U5397 ( .INP(n5314), .ZN(n128) );
  INVX0 U5398 ( .INP(n5315), .ZN(n127) );
  INVX0 U5399 ( .INP(n5316), .ZN(n126) );
  INVX0 U5400 ( .INP(n5317), .ZN(n125) );
  INVX0 U5401 ( .INP(n5318), .ZN(n124) );
  INVX0 U5402 ( .INP(n5319), .ZN(n123) );
  INVX0 U5403 ( .INP(n5320), .ZN(n122) );
  INVX0 U5404 ( .INP(n5321), .ZN(n121) );
  INVX0 U5405 ( .INP(n5322), .ZN(n120) );
  INVX0 U5406 ( .INP(n5323), .ZN(n12) );
  INVX0 U5407 ( .INP(n5324), .ZN(n119) );
  INVX0 U5408 ( .INP(n5325), .ZN(n118) );
  INVX0 U5409 ( .INP(n5326), .ZN(n117) );
  INVX0 U5410 ( .INP(n5327), .ZN(n116) );
  INVX0 U5411 ( .INP(n5328), .ZN(n115) );
  INVX0 U5412 ( .INP(n5329), .ZN(n114) );
  INVX0 U5413 ( .INP(n5330), .ZN(n113) );
  INVX0 U5414 ( .INP(n5331), .ZN(n112) );
  INVX0 U5415 ( .INP(n5332), .ZN(n111) );
  INVX0 U5416 ( .INP(n5333), .ZN(n110) );
  INVX0 U5417 ( .INP(n5334), .ZN(n11) );
  INVX0 U5418 ( .INP(n5335), .ZN(n109) );
  INVX0 U5419 ( .INP(n5336), .ZN(n108) );
  INVX0 U5420 ( .INP(n5337), .ZN(n107) );
  INVX0 U5421 ( .INP(n5338), .ZN(n106) );
  INVX0 U5422 ( .INP(n5339), .ZN(n105) );
  INVX0 U5423 ( .INP(n5340), .ZN(n104) );
  INVX0 U5424 ( .INP(n5341), .ZN(n103) );
  INVX0 U5425 ( .INP(n5342), .ZN(n102) );
  INVX0 U5426 ( .INP(n5343), .ZN(n101) );
  INVX0 U5427 ( .INP(n5344), .ZN(n100) );
  INVX0 U5428 ( .INP(n5345), .ZN(n10) );
  NOR2X0 U5429 ( .IN1(n8820), .IN2(n4848), .QN(WX9789) );
  NOR2X0 U5430 ( .IN1(n8823), .IN2(n4848), .QN(WX9787) );
  NOR2X0 U5431 ( .IN1(n8824), .IN2(n4848), .QN(WX9785) );
  NOR2X0 U5432 ( .IN1(n8827), .IN2(n4848), .QN(WX9783) );
  AND2X1 U5433 ( .IN1(n4800), .IN2(test_so80), .Q(WX9781) );
  NOR2X0 U5434 ( .IN1(n8828), .IN2(n4848), .QN(WX9779) );
  NOR2X0 U5435 ( .IN1(n8829), .IN2(n4848), .QN(WX9777) );
  NOR2X0 U5436 ( .IN1(n8830), .IN2(n4848), .QN(WX9775) );
  NOR2X0 U5437 ( .IN1(n8831), .IN2(n4848), .QN(WX9773) );
  NOR2X0 U5438 ( .IN1(n8832), .IN2(n4848), .QN(WX9771) );
  NOR2X0 U5439 ( .IN1(n8833), .IN2(n4848), .QN(WX9769) );
  NOR2X0 U5440 ( .IN1(n8834), .IN2(n4848), .QN(WX9767) );
  NOR2X0 U5441 ( .IN1(n8835), .IN2(n4849), .QN(WX9765) );
  NOR2X0 U5442 ( .IN1(n8836), .IN2(n4849), .QN(WX9763) );
  NOR2X0 U5443 ( .IN1(n8837), .IN2(n4849), .QN(WX9761) );
  NOR2X0 U5444 ( .IN1(n8838), .IN2(n4849), .QN(WX9759) );
  NAND2X0 U5445 ( .IN1(n5346), .IN2(n5347), .QN(WX9757) );
  NOR2X0 U5446 ( .IN1(n5348), .IN2(n5349), .QN(n5347) );
  AND2X1 U5447 ( .IN1(n5350), .IN2(n2153), .Q(n5349) );
  NOR2X0 U5448 ( .IN1(n5351), .IN2(n4253), .QN(n5348) );
  NOR2X0 U5449 ( .IN1(n5353), .IN2(n5354), .QN(n5346) );
  NOR2X0 U5450 ( .IN1(DFF_1504_n1), .IN2(n4287), .QN(n5354) );
  NOR2X0 U5451 ( .IN1(n5356), .IN2(n5214), .QN(n5353) );
  NAND2X0 U5452 ( .IN1(n4805), .IN2(n8321), .QN(n5214) );
  NAND2X0 U5453 ( .IN1(n5357), .IN2(n5358), .QN(WX9755) );
  NOR2X0 U5454 ( .IN1(n5359), .IN2(n5360), .QN(n5358) );
  AND2X1 U5455 ( .IN1(n5361), .IN2(n2153), .Q(n5360) );
  NOR2X0 U5456 ( .IN1(n4258), .IN2(n5362), .QN(n5359) );
  NOR2X0 U5457 ( .IN1(n5363), .IN2(n5364), .QN(n5357) );
  NOR2X0 U5458 ( .IN1(DFF_1505_n1), .IN2(n4280), .QN(n5364) );
  NOR2X0 U5459 ( .IN1(n4312), .IN2(n5215), .QN(n5363) );
  NAND2X0 U5460 ( .IN1(n4805), .IN2(n8322), .QN(n5215) );
  NAND2X0 U5461 ( .IN1(n5365), .IN2(n5366), .QN(WX9753) );
  NOR2X0 U5462 ( .IN1(n5367), .IN2(n5368), .QN(n5366) );
  NOR2X0 U5463 ( .IN1(n4338), .IN2(n5370), .QN(n5368) );
  NOR2X0 U5464 ( .IN1(n5371), .IN2(n4247), .QN(n5367) );
  NOR2X0 U5465 ( .IN1(n5372), .IN2(n5373), .QN(n5365) );
  AND2X1 U5466 ( .IN1(n2152), .IN2(test_so87), .Q(n5373) );
  NOR2X0 U5467 ( .IN1(n4312), .IN2(n5216), .QN(n5372) );
  NAND2X0 U5468 ( .IN1(n4805), .IN2(n8323), .QN(n5216) );
  NAND2X0 U5469 ( .IN1(n5374), .IN2(n5375), .QN(WX9751) );
  NOR2X0 U5470 ( .IN1(n5376), .IN2(n5377), .QN(n5375) );
  AND2X1 U5471 ( .IN1(n5378), .IN2(n2153), .Q(n5377) );
  NOR2X0 U5472 ( .IN1(n4258), .IN2(n5379), .QN(n5376) );
  NOR2X0 U5473 ( .IN1(n5380), .IN2(n5381), .QN(n5374) );
  NOR2X0 U5474 ( .IN1(DFF_1507_n1), .IN2(n4287), .QN(n5381) );
  NOR2X0 U5475 ( .IN1(n4312), .IN2(n5217), .QN(n5380) );
  NAND2X0 U5476 ( .IN1(n4805), .IN2(n8324), .QN(n5217) );
  NAND2X0 U5477 ( .IN1(n5382), .IN2(n5383), .QN(WX9749) );
  NOR2X0 U5478 ( .IN1(n5384), .IN2(n5385), .QN(n5383) );
  NOR2X0 U5479 ( .IN1(n4340), .IN2(n5386), .QN(n5385) );
  NOR2X0 U5480 ( .IN1(n5387), .IN2(n4247), .QN(n5384) );
  NOR2X0 U5481 ( .IN1(n5388), .IN2(n5389), .QN(n5382) );
  NOR2X0 U5482 ( .IN1(DFF_1508_n1), .IN2(n4287), .QN(n5389) );
  NOR2X0 U5483 ( .IN1(n4312), .IN2(n5218), .QN(n5388) );
  NAND2X0 U5484 ( .IN1(n4805), .IN2(n8325), .QN(n5218) );
  NAND2X0 U5485 ( .IN1(n5390), .IN2(n5391), .QN(WX9747) );
  NOR2X0 U5486 ( .IN1(n5392), .IN2(n5393), .QN(n5391) );
  AND2X1 U5487 ( .IN1(n5394), .IN2(n2153), .Q(n5393) );
  NOR2X0 U5488 ( .IN1(n5395), .IN2(n4247), .QN(n5392) );
  NOR2X0 U5489 ( .IN1(n5396), .IN2(n5397), .QN(n5390) );
  NOR2X0 U5490 ( .IN1(DFF_1509_n1), .IN2(n4287), .QN(n5397) );
  NOR2X0 U5491 ( .IN1(n4312), .IN2(n5219), .QN(n5396) );
  NAND2X0 U5492 ( .IN1(test_so79), .IN2(n4827), .QN(n5219) );
  NAND2X0 U5493 ( .IN1(n5398), .IN2(n5399), .QN(WX9745) );
  NOR2X0 U5494 ( .IN1(n5400), .IN2(n5401), .QN(n5399) );
  NOR2X0 U5495 ( .IN1(n4340), .IN2(n5402), .QN(n5401) );
  NOR2X0 U5496 ( .IN1(n5403), .IN2(n4247), .QN(n5400) );
  NOR2X0 U5497 ( .IN1(n5404), .IN2(n5405), .QN(n5398) );
  NOR2X0 U5498 ( .IN1(DFF_1510_n1), .IN2(n4287), .QN(n5405) );
  NOR2X0 U5499 ( .IN1(n4312), .IN2(n5220), .QN(n5404) );
  NAND2X0 U5500 ( .IN1(n4805), .IN2(n8328), .QN(n5220) );
  NAND2X0 U5501 ( .IN1(n5406), .IN2(n5407), .QN(WX9743) );
  NOR2X0 U5502 ( .IN1(n5408), .IN2(n5409), .QN(n5407) );
  AND2X1 U5503 ( .IN1(n5410), .IN2(n2153), .Q(n5409) );
  NOR2X0 U5504 ( .IN1(n5411), .IN2(n4247), .QN(n5408) );
  NOR2X0 U5505 ( .IN1(n5412), .IN2(n5413), .QN(n5406) );
  NOR2X0 U5506 ( .IN1(DFF_1511_n1), .IN2(n4287), .QN(n5413) );
  NOR2X0 U5507 ( .IN1(n4312), .IN2(n5221), .QN(n5412) );
  NAND2X0 U5508 ( .IN1(n4805), .IN2(n8329), .QN(n5221) );
  NAND2X0 U5509 ( .IN1(n5414), .IN2(n5415), .QN(WX9741) );
  NOR2X0 U5510 ( .IN1(n5416), .IN2(n5417), .QN(n5415) );
  NOR2X0 U5511 ( .IN1(n4340), .IN2(n5418), .QN(n5417) );
  NOR2X0 U5512 ( .IN1(n5419), .IN2(n4248), .QN(n5416) );
  NOR2X0 U5513 ( .IN1(n5420), .IN2(n5421), .QN(n5414) );
  NOR2X0 U5514 ( .IN1(DFF_1512_n1), .IN2(n4286), .QN(n5421) );
  NOR2X0 U5515 ( .IN1(n4312), .IN2(n5222), .QN(n5420) );
  NAND2X0 U5516 ( .IN1(n4805), .IN2(n8330), .QN(n5222) );
  NAND2X0 U5517 ( .IN1(n5422), .IN2(n5423), .QN(WX9739) );
  NOR2X0 U5518 ( .IN1(n5424), .IN2(n5425), .QN(n5423) );
  AND2X1 U5519 ( .IN1(n5426), .IN2(n2153), .Q(n5425) );
  NOR2X0 U5520 ( .IN1(n5427), .IN2(n4247), .QN(n5424) );
  NOR2X0 U5521 ( .IN1(n5428), .IN2(n5429), .QN(n5422) );
  NOR2X0 U5522 ( .IN1(DFF_1513_n1), .IN2(n4286), .QN(n5429) );
  NOR2X0 U5523 ( .IN1(n4312), .IN2(n5224), .QN(n5428) );
  NAND2X0 U5524 ( .IN1(n4806), .IN2(n8331), .QN(n5224) );
  NAND2X0 U5525 ( .IN1(n5430), .IN2(n5431), .QN(WX9737) );
  NOR2X0 U5526 ( .IN1(n5432), .IN2(n5433), .QN(n5431) );
  AND2X1 U5527 ( .IN1(n5434), .IN2(n2153), .Q(n5433) );
  NOR2X0 U5528 ( .IN1(n5435), .IN2(n4247), .QN(n5432) );
  NOR2X0 U5529 ( .IN1(n5436), .IN2(n5437), .QN(n5430) );
  NOR2X0 U5530 ( .IN1(DFF_1514_n1), .IN2(n4286), .QN(n5437) );
  NOR2X0 U5531 ( .IN1(n4312), .IN2(n5225), .QN(n5436) );
  NAND2X0 U5532 ( .IN1(n4806), .IN2(n8332), .QN(n5225) );
  NAND2X0 U5533 ( .IN1(n5438), .IN2(n5439), .QN(WX9735) );
  NOR2X0 U5534 ( .IN1(n5440), .IN2(n5441), .QN(n5439) );
  AND2X1 U5535 ( .IN1(n5442), .IN2(n2153), .Q(n5441) );
  NOR2X0 U5536 ( .IN1(n5443), .IN2(n4247), .QN(n5440) );
  NOR2X0 U5537 ( .IN1(n5444), .IN2(n5445), .QN(n5438) );
  NOR2X0 U5538 ( .IN1(DFF_1515_n1), .IN2(n4286), .QN(n5445) );
  NOR2X0 U5539 ( .IN1(n4312), .IN2(n5226), .QN(n5444) );
  NAND2X0 U5540 ( .IN1(n4806), .IN2(n8333), .QN(n5226) );
  NAND2X0 U5541 ( .IN1(n5446), .IN2(n5447), .QN(WX9733) );
  NOR2X0 U5542 ( .IN1(n5448), .IN2(n5449), .QN(n5447) );
  AND2X1 U5543 ( .IN1(n5450), .IN2(n2153), .Q(n5449) );
  NOR2X0 U5544 ( .IN1(n5451), .IN2(n4248), .QN(n5448) );
  NOR2X0 U5545 ( .IN1(n5452), .IN2(n5453), .QN(n5446) );
  NOR2X0 U5546 ( .IN1(DFF_1516_n1), .IN2(n4286), .QN(n5453) );
  NOR2X0 U5547 ( .IN1(n4312), .IN2(n5227), .QN(n5452) );
  NAND2X0 U5548 ( .IN1(n4806), .IN2(n8334), .QN(n5227) );
  NAND2X0 U5549 ( .IN1(n5454), .IN2(n5455), .QN(WX9731) );
  NOR2X0 U5550 ( .IN1(n5456), .IN2(n5457), .QN(n5455) );
  AND2X1 U5551 ( .IN1(n5458), .IN2(n2153), .Q(n5457) );
  NOR2X0 U5552 ( .IN1(n5459), .IN2(n4247), .QN(n5456) );
  NOR2X0 U5553 ( .IN1(n5460), .IN2(n5461), .QN(n5454) );
  NOR2X0 U5554 ( .IN1(DFF_1517_n1), .IN2(n4286), .QN(n5461) );
  NOR2X0 U5555 ( .IN1(n4311), .IN2(n5228), .QN(n5460) );
  NAND2X0 U5556 ( .IN1(n4806), .IN2(n8335), .QN(n5228) );
  NAND2X0 U5557 ( .IN1(n5462), .IN2(n5463), .QN(WX9729) );
  NOR2X0 U5558 ( .IN1(n5464), .IN2(n5465), .QN(n5463) );
  AND2X1 U5559 ( .IN1(n5466), .IN2(n2153), .Q(n5465) );
  NOR2X0 U5560 ( .IN1(n4258), .IN2(n5467), .QN(n5464) );
  NOR2X0 U5561 ( .IN1(n5468), .IN2(n5469), .QN(n5462) );
  NOR2X0 U5562 ( .IN1(DFF_1518_n1), .IN2(n4286), .QN(n5469) );
  NOR2X0 U5563 ( .IN1(n4311), .IN2(n5229), .QN(n5468) );
  NAND2X0 U5564 ( .IN1(n4806), .IN2(n8336), .QN(n5229) );
  NAND2X0 U5565 ( .IN1(n5470), .IN2(n5471), .QN(WX9727) );
  NOR2X0 U5566 ( .IN1(n5472), .IN2(n5473), .QN(n5471) );
  AND2X1 U5567 ( .IN1(n5474), .IN2(n2153), .Q(n5473) );
  NOR2X0 U5568 ( .IN1(n5475), .IN2(n4247), .QN(n5472) );
  NOR2X0 U5569 ( .IN1(n5476), .IN2(n5477), .QN(n5470) );
  NOR2X0 U5570 ( .IN1(DFF_1519_n1), .IN2(n4286), .QN(n5477) );
  NOR2X0 U5571 ( .IN1(n4311), .IN2(n5230), .QN(n5476) );
  NAND2X0 U5572 ( .IN1(n4806), .IN2(n8337), .QN(n5230) );
  NAND2X0 U5573 ( .IN1(n5478), .IN2(n5479), .QN(WX9725) );
  NOR2X0 U5574 ( .IN1(n5480), .IN2(n5481), .QN(n5479) );
  AND2X1 U5575 ( .IN1(n5482), .IN2(n2153), .Q(n5481) );
  NOR2X0 U5576 ( .IN1(n4258), .IN2(n5483), .QN(n5480) );
  NOR2X0 U5577 ( .IN1(n5484), .IN2(n5485), .QN(n5478) );
  NOR2X0 U5578 ( .IN1(DFF_1520_n1), .IN2(n4286), .QN(n5485) );
  NOR2X0 U5579 ( .IN1(n4311), .IN2(n5231), .QN(n5484) );
  NAND2X0 U5580 ( .IN1(n4806), .IN2(n8338), .QN(n5231) );
  NAND2X0 U5581 ( .IN1(n5486), .IN2(n5487), .QN(WX9723) );
  NOR2X0 U5582 ( .IN1(n5488), .IN2(n5489), .QN(n5487) );
  AND2X1 U5583 ( .IN1(n5490), .IN2(n2153), .Q(n5489) );
  NOR2X0 U5584 ( .IN1(n5491), .IN2(n4248), .QN(n5488) );
  NOR2X0 U5585 ( .IN1(n5492), .IN2(n5493), .QN(n5486) );
  NOR2X0 U5586 ( .IN1(DFF_1521_n1), .IN2(n4286), .QN(n5493) );
  NOR2X0 U5587 ( .IN1(n4311), .IN2(n5232), .QN(n5492) );
  NAND2X0 U5588 ( .IN1(n4806), .IN2(n8339), .QN(n5232) );
  NAND2X0 U5589 ( .IN1(n5494), .IN2(n5495), .QN(WX9721) );
  NOR2X0 U5590 ( .IN1(n5496), .IN2(n5497), .QN(n5495) );
  AND2X1 U5591 ( .IN1(n5498), .IN2(n2153), .Q(n5497) );
  NOR2X0 U5592 ( .IN1(n4258), .IN2(n5499), .QN(n5496) );
  NOR2X0 U5593 ( .IN1(n5500), .IN2(n5501), .QN(n5494) );
  NOR2X0 U5594 ( .IN1(DFF_1522_n1), .IN2(n4286), .QN(n5501) );
  NOR2X0 U5595 ( .IN1(n4311), .IN2(n5233), .QN(n5500) );
  NAND2X0 U5596 ( .IN1(n4807), .IN2(n8340), .QN(n5233) );
  NAND2X0 U5597 ( .IN1(n5502), .IN2(n5503), .QN(WX9719) );
  NOR2X0 U5598 ( .IN1(n5504), .IN2(n5505), .QN(n5503) );
  NOR2X0 U5599 ( .IN1(n4340), .IN2(n5506), .QN(n5505) );
  NOR2X0 U5600 ( .IN1(n5507), .IN2(n4248), .QN(n5504) );
  NOR2X0 U5601 ( .IN1(n5508), .IN2(n5509), .QN(n5502) );
  AND2X1 U5602 ( .IN1(n2152), .IN2(test_so88), .Q(n5509) );
  NOR2X0 U5603 ( .IN1(n4311), .IN2(n5236), .QN(n5508) );
  NAND2X0 U5604 ( .IN1(n4807), .IN2(n8341), .QN(n5236) );
  NAND2X0 U5605 ( .IN1(n5510), .IN2(n5511), .QN(WX9717) );
  NOR2X0 U5606 ( .IN1(n5512), .IN2(n5513), .QN(n5511) );
  AND2X1 U5607 ( .IN1(n5514), .IN2(n2153), .Q(n5513) );
  NOR2X0 U5608 ( .IN1(n4258), .IN2(n5515), .QN(n5512) );
  NOR2X0 U5609 ( .IN1(n5516), .IN2(n5517), .QN(n5510) );
  NOR2X0 U5610 ( .IN1(DFF_1524_n1), .IN2(n4286), .QN(n5517) );
  NOR2X0 U5611 ( .IN1(n4311), .IN2(n5237), .QN(n5516) );
  NAND2X0 U5612 ( .IN1(n4807), .IN2(n8342), .QN(n5237) );
  NAND2X0 U5613 ( .IN1(n5518), .IN2(n5519), .QN(WX9715) );
  NOR2X0 U5614 ( .IN1(n5520), .IN2(n5521), .QN(n5519) );
  NOR2X0 U5615 ( .IN1(n4340), .IN2(n5522), .QN(n5521) );
  NOR2X0 U5616 ( .IN1(n5523), .IN2(n4248), .QN(n5520) );
  NOR2X0 U5617 ( .IN1(n5524), .IN2(n5525), .QN(n5518) );
  NOR2X0 U5618 ( .IN1(DFF_1525_n1), .IN2(n4286), .QN(n5525) );
  NOR2X0 U5619 ( .IN1(n4311), .IN2(n5238), .QN(n5524) );
  NAND2X0 U5620 ( .IN1(n4807), .IN2(n8343), .QN(n5238) );
  NAND2X0 U5621 ( .IN1(n5526), .IN2(n5527), .QN(WX9713) );
  NOR2X0 U5622 ( .IN1(n5528), .IN2(n5529), .QN(n5527) );
  AND2X1 U5623 ( .IN1(n5530), .IN2(n2153), .Q(n5529) );
  NOR2X0 U5624 ( .IN1(n5531), .IN2(n4248), .QN(n5528) );
  NOR2X0 U5625 ( .IN1(n5532), .IN2(n5533), .QN(n5526) );
  NOR2X0 U5626 ( .IN1(DFF_1526_n1), .IN2(n4286), .QN(n5533) );
  NOR2X0 U5627 ( .IN1(n4311), .IN2(n5239), .QN(n5532) );
  NAND2X0 U5628 ( .IN1(test_so78), .IN2(n4828), .QN(n5239) );
  NAND2X0 U5629 ( .IN1(n5534), .IN2(n5535), .QN(WX9711) );
  NOR2X0 U5630 ( .IN1(n5536), .IN2(n5537), .QN(n5535) );
  NOR2X0 U5631 ( .IN1(n4340), .IN2(n5538), .QN(n5537) );
  NOR2X0 U5632 ( .IN1(n5539), .IN2(n4248), .QN(n5536) );
  NOR2X0 U5633 ( .IN1(n5540), .IN2(n5541), .QN(n5534) );
  NOR2X0 U5634 ( .IN1(DFF_1527_n1), .IN2(n4285), .QN(n5541) );
  NOR2X0 U5635 ( .IN1(n4311), .IN2(n5240), .QN(n5540) );
  NAND2X0 U5636 ( .IN1(n4807), .IN2(n8346), .QN(n5240) );
  NAND2X0 U5637 ( .IN1(n5542), .IN2(n5543), .QN(WX9709) );
  NOR2X0 U5638 ( .IN1(n5544), .IN2(n5545), .QN(n5543) );
  AND2X1 U5639 ( .IN1(n5546), .IN2(n2153), .Q(n5545) );
  NOR2X0 U5640 ( .IN1(n5547), .IN2(n4248), .QN(n5544) );
  NOR2X0 U5641 ( .IN1(n5548), .IN2(n5549), .QN(n5542) );
  NOR2X0 U5642 ( .IN1(DFF_1528_n1), .IN2(n4285), .QN(n5549) );
  NOR2X0 U5643 ( .IN1(n4311), .IN2(n5241), .QN(n5548) );
  NAND2X0 U5644 ( .IN1(n4807), .IN2(n8347), .QN(n5241) );
  NAND2X0 U5645 ( .IN1(n5550), .IN2(n5551), .QN(WX9707) );
  NOR2X0 U5646 ( .IN1(n5552), .IN2(n5553), .QN(n5551) );
  NOR2X0 U5647 ( .IN1(n4340), .IN2(n5554), .QN(n5553) );
  NOR2X0 U5648 ( .IN1(n5555), .IN2(n4248), .QN(n5552) );
  NOR2X0 U5649 ( .IN1(n5556), .IN2(n5557), .QN(n5550) );
  NOR2X0 U5650 ( .IN1(DFF_1529_n1), .IN2(n4285), .QN(n5557) );
  NOR2X0 U5651 ( .IN1(n4310), .IN2(n5242), .QN(n5556) );
  NAND2X0 U5652 ( .IN1(n4807), .IN2(n8348), .QN(n5242) );
  NAND2X0 U5653 ( .IN1(n5558), .IN2(n5559), .QN(WX9705) );
  NOR2X0 U5654 ( .IN1(n5560), .IN2(n5561), .QN(n5559) );
  AND2X1 U5655 ( .IN1(n5562), .IN2(n2153), .Q(n5561) );
  NOR2X0 U5656 ( .IN1(n5563), .IN2(n4248), .QN(n5560) );
  NOR2X0 U5657 ( .IN1(n5564), .IN2(n5565), .QN(n5558) );
  NOR2X0 U5658 ( .IN1(DFF_1530_n1), .IN2(n4285), .QN(n5565) );
  NOR2X0 U5659 ( .IN1(n4310), .IN2(n5243), .QN(n5564) );
  NAND2X0 U5660 ( .IN1(n4807), .IN2(n8349), .QN(n5243) );
  NAND2X0 U5661 ( .IN1(n5566), .IN2(n5567), .QN(WX9703) );
  NOR2X0 U5662 ( .IN1(n5568), .IN2(n5569), .QN(n5567) );
  AND2X1 U5663 ( .IN1(n5570), .IN2(n2153), .Q(n5569) );
  NOR2X0 U5664 ( .IN1(n5571), .IN2(n4248), .QN(n5568) );
  NOR2X0 U5665 ( .IN1(n5572), .IN2(n5573), .QN(n5566) );
  NOR2X0 U5666 ( .IN1(DFF_1531_n1), .IN2(n4285), .QN(n5573) );
  NOR2X0 U5667 ( .IN1(n4310), .IN2(n5244), .QN(n5572) );
  NAND2X0 U5668 ( .IN1(n4807), .IN2(n8350), .QN(n5244) );
  NAND2X0 U5669 ( .IN1(n5574), .IN2(n5575), .QN(WX9701) );
  NOR2X0 U5670 ( .IN1(n5576), .IN2(n5577), .QN(n5575) );
  AND2X1 U5671 ( .IN1(n5578), .IN2(n2153), .Q(n5577) );
  NOR2X0 U5672 ( .IN1(n5579), .IN2(n4249), .QN(n5576) );
  NOR2X0 U5673 ( .IN1(n5580), .IN2(n5581), .QN(n5574) );
  NOR2X0 U5674 ( .IN1(DFF_1532_n1), .IN2(n4285), .QN(n5581) );
  NOR2X0 U5675 ( .IN1(n4310), .IN2(n5245), .QN(n5580) );
  NAND2X0 U5676 ( .IN1(n4808), .IN2(n8351), .QN(n5245) );
  NAND2X0 U5677 ( .IN1(n5582), .IN2(n5583), .QN(WX9699) );
  NOR2X0 U5678 ( .IN1(n5584), .IN2(n5585), .QN(n5583) );
  AND2X1 U5679 ( .IN1(n5586), .IN2(n2153), .Q(n5585) );
  NOR2X0 U5680 ( .IN1(n5587), .IN2(n4248), .QN(n5584) );
  NOR2X0 U5681 ( .IN1(n5588), .IN2(n5589), .QN(n5582) );
  NOR2X0 U5682 ( .IN1(DFF_1533_n1), .IN2(n4285), .QN(n5589) );
  NOR2X0 U5683 ( .IN1(n4310), .IN2(n5247), .QN(n5588) );
  NAND2X0 U5684 ( .IN1(n4808), .IN2(n8352), .QN(n5247) );
  NAND2X0 U5685 ( .IN1(n5590), .IN2(n5591), .QN(WX9697) );
  NOR2X0 U5686 ( .IN1(n5592), .IN2(n5593), .QN(n5591) );
  AND2X1 U5687 ( .IN1(n5594), .IN2(n2153), .Q(n5593) );
  NOR2X0 U5688 ( .IN1(n5595), .IN2(n4248), .QN(n5592) );
  NOR2X0 U5689 ( .IN1(n5596), .IN2(n5597), .QN(n5590) );
  NOR2X0 U5690 ( .IN1(DFF_1534_n1), .IN2(n4285), .QN(n5597) );
  NOR2X0 U5691 ( .IN1(n4310), .IN2(n5248), .QN(n5596) );
  NAND2X0 U5692 ( .IN1(n4808), .IN2(n8353), .QN(n5248) );
  NAND2X0 U5693 ( .IN1(n5598), .IN2(n5599), .QN(WX9695) );
  NOR2X0 U5694 ( .IN1(n5600), .IN2(n5601), .QN(n5599) );
  AND2X1 U5695 ( .IN1(n5602), .IN2(n2153), .Q(n5601) );
  NOR2X0 U5696 ( .IN1(n4259), .IN2(n5603), .QN(n5600) );
  NOR2X0 U5697 ( .IN1(n5604), .IN2(n5605), .QN(n5598) );
  NOR2X0 U5698 ( .IN1(n3932), .IN2(n5606), .QN(n5605) );
  NOR2X0 U5699 ( .IN1(DFF_1535_n1), .IN2(n4285), .QN(n5604) );
  AND2X1 U5700 ( .IN1(n4800), .IN2(n3932), .Q(WX9597) );
  NOR2X0 U5701 ( .IN1(n4926), .IN2(n5607), .QN(WX9084) );
  XOR2X1 U5702 ( .IN1(n4020), .IN2(DFF_1342_n1), .Q(n5607) );
  NOR2X0 U5703 ( .IN1(n4940), .IN2(n5608), .QN(WX9082) );
  XOR2X1 U5704 ( .IN1(n4021), .IN2(DFF_1341_n1), .Q(n5608) );
  NOR2X0 U5705 ( .IN1(n4934), .IN2(n5609), .QN(WX9080) );
  XOR2X1 U5706 ( .IN1(n4022), .IN2(DFF_1340_n1), .Q(n5609) );
  NOR2X0 U5707 ( .IN1(n4934), .IN2(n5610), .QN(WX9078) );
  XOR2X1 U5708 ( .IN1(n4023), .IN2(DFF_1339_n1), .Q(n5610) );
  NOR2X0 U5709 ( .IN1(n4934), .IN2(n5611), .QN(WX9076) );
  XOR2X1 U5710 ( .IN1(n4024), .IN2(DFF_1338_n1), .Q(n5611) );
  NOR2X0 U5711 ( .IN1(n4934), .IN2(n5612), .QN(WX9074) );
  XNOR2X1 U5712 ( .IN1(DFF_1337_n1), .IN2(test_so74), .Q(n5612) );
  NOR2X0 U5713 ( .IN1(n4934), .IN2(n5613), .QN(WX9072) );
  XNOR2X1 U5714 ( .IN1(n4025), .IN2(test_so77), .Q(n5613) );
  NOR2X0 U5715 ( .IN1(n4934), .IN2(n5614), .QN(WX9070) );
  XOR2X1 U6483 ( .IN1(n4026), .IN2(DFF_1335_n1), .Q(n5614) );
  NOR2X0 U6484 ( .IN1(n4934), .IN2(n5615), .QN(WX9068) );
  XOR2X1 U6485 ( .IN1(n4027), .IN2(DFF_1334_n1), .Q(n5615) );
  NOR2X0 U6486 ( .IN1(n4934), .IN2(n5616), .QN(WX9066) );
  XOR2X1 U6487 ( .IN1(n4028), .IN2(DFF_1333_n1), .Q(n5616) );
  NOR2X0 U6488 ( .IN1(n4934), .IN2(n5617), .QN(WX9064) );
  XOR2X1 U6489 ( .IN1(n4029), .IN2(DFF_1332_n1), .Q(n5617) );
  NOR2X0 U6490 ( .IN1(n4934), .IN2(n5618), .QN(WX9062) );
  XOR2X1 U6491 ( .IN1(n4030), .IN2(DFF_1331_n1), .Q(n5618) );
  NOR2X0 U6492 ( .IN1(n4934), .IN2(n5619), .QN(WX9060) );
  XOR2X1 U6493 ( .IN1(n4031), .IN2(DFF_1330_n1), .Q(n5619) );
  NOR2X0 U6494 ( .IN1(n4934), .IN2(n5620), .QN(WX9058) );
  XOR2X1 U6495 ( .IN1(n4032), .IN2(DFF_1329_n1), .Q(n5620) );
  NOR2X0 U6496 ( .IN1(n4934), .IN2(n5621), .QN(WX9056) );
  XOR2X1 U6497 ( .IN1(n4033), .IN2(DFF_1328_n1), .Q(n5621) );
  NOR2X0 U6498 ( .IN1(n4935), .IN2(n5622), .QN(WX9054) );
  XNOR2X1 U6499 ( .IN1(DFF_1327_n1), .IN2(n5623), .Q(n5622) );
  XOR2X1 U6500 ( .IN1(n3945), .IN2(DFF_1343_n1), .Q(n5623) );
  NOR2X0 U6501 ( .IN1(n4935), .IN2(n5624), .QN(WX9052) );
  XOR2X1 U6502 ( .IN1(n4034), .IN2(DFF_1326_n1), .Q(n5624) );
  NOR2X0 U6503 ( .IN1(n4935), .IN2(n5625), .QN(WX9050) );
  XOR2X1 U6504 ( .IN1(n4035), .IN2(DFF_1325_n1), .Q(n5625) );
  NOR2X0 U6505 ( .IN1(n4935), .IN2(n5626), .QN(WX9048) );
  XOR2X1 U6506 ( .IN1(n4036), .IN2(DFF_1324_n1), .Q(n5626) );
  NOR2X0 U6507 ( .IN1(n4935), .IN2(n5627), .QN(WX9046) );
  XOR2X1 U6508 ( .IN1(n4037), .IN2(DFF_1323_n1), .Q(n5627) );
  NOR2X0 U6509 ( .IN1(n4935), .IN2(n5628), .QN(WX9044) );
  XNOR2X1 U6510 ( .IN1(DFF_1322_n1), .IN2(n5629), .Q(n5628) );
  XOR2X1 U6511 ( .IN1(n3946), .IN2(DFF_1343_n1), .Q(n5629) );
  NOR2X0 U6512 ( .IN1(n4935), .IN2(n5630), .QN(WX9042) );
  XOR2X1 U6513 ( .IN1(n4038), .IN2(DFF_1321_n1), .Q(n5630) );
  NOR2X0 U6514 ( .IN1(n4935), .IN2(n5631), .QN(WX9040) );
  XNOR2X1 U6515 ( .IN1(DFF_1320_n1), .IN2(test_so75), .Q(n5631) );
  NOR2X0 U6516 ( .IN1(n4935), .IN2(n5632), .QN(WX9038) );
  XNOR2X1 U6517 ( .IN1(n4039), .IN2(test_so76), .Q(n5632) );
  NOR2X0 U6518 ( .IN1(n4935), .IN2(n5633), .QN(WX9036) );
  XOR2X1 U6519 ( .IN1(n4040), .IN2(DFF_1318_n1), .Q(n5633) );
  NOR2X0 U6520 ( .IN1(n4935), .IN2(n5634), .QN(WX9034) );
  XOR2X1 U6521 ( .IN1(n4041), .IN2(DFF_1317_n1), .Q(n5634) );
  NOR2X0 U6522 ( .IN1(n4935), .IN2(n5635), .QN(WX9032) );
  XOR2X1 U6523 ( .IN1(n4042), .IN2(DFF_1316_n1), .Q(n5635) );
  NOR2X0 U6524 ( .IN1(n4935), .IN2(n5636), .QN(WX9030) );
  XNOR2X1 U6525 ( .IN1(DFF_1315_n1), .IN2(n5637), .Q(n5636) );
  XOR2X1 U6526 ( .IN1(n3947), .IN2(DFF_1343_n1), .Q(n5637) );
  NOR2X0 U6527 ( .IN1(n4936), .IN2(n5638), .QN(WX9028) );
  XOR2X1 U6528 ( .IN1(n4043), .IN2(DFF_1314_n1), .Q(n5638) );
  NOR2X0 U6529 ( .IN1(n4936), .IN2(n5639), .QN(WX9026) );
  XOR2X1 U6530 ( .IN1(n4044), .IN2(DFF_1313_n1), .Q(n5639) );
  NOR2X0 U6531 ( .IN1(n4936), .IN2(n5640), .QN(WX9024) );
  XOR2X1 U6532 ( .IN1(n4045), .IN2(DFF_1312_n1), .Q(n5640) );
  NOR2X0 U6533 ( .IN1(n4936), .IN2(n5641), .QN(WX9022) );
  XOR2X1 U6534 ( .IN1(n3962), .IN2(DFF_1343_n1), .Q(n5641) );
  NOR2X0 U6535 ( .IN1(n8855), .IN2(n4849), .QN(WX8496) );
  NOR2X0 U6536 ( .IN1(n8856), .IN2(n4849), .QN(WX8494) );
  NOR2X0 U6537 ( .IN1(n8857), .IN2(n4849), .QN(WX8492) );
  NOR2X0 U6538 ( .IN1(n8858), .IN2(n4849), .QN(WX8490) );
  NOR2X0 U6539 ( .IN1(n8859), .IN2(n4849), .QN(WX8488) );
  NOR2X0 U6540 ( .IN1(n8860), .IN2(n4849), .QN(WX8486) );
  NOR2X0 U6541 ( .IN1(n8861), .IN2(n4849), .QN(WX8484) );
  NOR2X0 U6542 ( .IN1(n8862), .IN2(n4849), .QN(WX8482) );
  NOR2X0 U6543 ( .IN1(n8863), .IN2(n4850), .QN(WX8480) );
  NOR2X0 U6544 ( .IN1(n8864), .IN2(n4850), .QN(WX8478) );
  NOR2X0 U6545 ( .IN1(n8865), .IN2(n4850), .QN(WX8476) );
  NOR2X0 U6546 ( .IN1(n8866), .IN2(n4850), .QN(WX8474) );
  NOR2X0 U6547 ( .IN1(n8867), .IN2(n4850), .QN(WX8472) );
  NOR2X0 U6548 ( .IN1(n8870), .IN2(n4850), .QN(WX8470) );
  NOR2X0 U6549 ( .IN1(n8871), .IN2(n4850), .QN(WX8468) );
  NOR2X0 U6550 ( .IN1(n8874), .IN2(n4850), .QN(WX8466) );
  NAND2X0 U6551 ( .IN1(n5642), .IN2(n5643), .QN(WX8464) );
  NOR2X0 U6552 ( .IN1(n5644), .IN2(n5645), .QN(n5643) );
  NOR2X0 U6553 ( .IN1(n5646), .IN2(n4248), .QN(n5645) );
  NOR2X0 U6554 ( .IN1(n5351), .IN2(n4326), .QN(n5644) );
  XOR2X1 U6555 ( .IN1(n5647), .IN2(n5648), .Q(n5351) );
  XOR2X1 U6556 ( .IN1(n8804), .IN2(n3961), .Q(n5648) );
  XOR2X1 U6557 ( .IN1(WX9758), .IN2(n3726), .Q(n5647) );
  NOR2X0 U6558 ( .IN1(n5649), .IN2(n5650), .QN(n5642) );
  NOR2X0 U6559 ( .IN1(DFF_1312_n1), .IN2(n4285), .QN(n5650) );
  NOR2X0 U6560 ( .IN1(n4310), .IN2(n5249), .QN(n5649) );
  NAND2X0 U6561 ( .IN1(test_so68), .IN2(n4828), .QN(n5249) );
  NAND2X0 U6562 ( .IN1(n5651), .IN2(n5652), .QN(WX8462) );
  NOR2X0 U6563 ( .IN1(n5653), .IN2(n5654), .QN(n5652) );
  NOR2X0 U6564 ( .IN1(n5655), .IN2(n4249), .QN(n5654) );
  NOR2X0 U6565 ( .IN1(n4340), .IN2(n5362), .QN(n5653) );
  XNOR2X1 U6566 ( .IN1(n5656), .IN2(n5657), .Q(n5362) );
  XOR2X1 U6567 ( .IN1(test_so83), .IN2(n8805), .Q(n5657) );
  XOR2X1 U6568 ( .IN1(WX9756), .IN2(n4019), .Q(n5656) );
  NOR2X0 U6569 ( .IN1(n5658), .IN2(n5659), .QN(n5651) );
  NOR2X0 U6570 ( .IN1(DFF_1313_n1), .IN2(n4285), .QN(n5659) );
  NOR2X0 U6571 ( .IN1(n4310), .IN2(n5250), .QN(n5658) );
  NAND2X0 U6572 ( .IN1(n4808), .IN2(n8381), .QN(n5250) );
  NAND2X0 U6573 ( .IN1(n5660), .IN2(n5661), .QN(WX8460) );
  NOR2X0 U6574 ( .IN1(n5662), .IN2(n5663), .QN(n5661) );
  NOR2X0 U6575 ( .IN1(n5664), .IN2(n4249), .QN(n5663) );
  NOR2X0 U6576 ( .IN1(n5371), .IN2(n4327), .QN(n5662) );
  XOR2X1 U6577 ( .IN1(n5665), .IN2(n5666), .Q(n5371) );
  XOR2X1 U6578 ( .IN1(n8806), .IN2(n4018), .Q(n5666) );
  XOR2X1 U6579 ( .IN1(WX9754), .IN2(n3729), .Q(n5665) );
  NOR2X0 U6580 ( .IN1(n5667), .IN2(n5668), .QN(n5660) );
  NOR2X0 U6581 ( .IN1(DFF_1314_n1), .IN2(n4285), .QN(n5668) );
  NOR2X0 U6582 ( .IN1(n4310), .IN2(n5251), .QN(n5667) );
  NAND2X0 U6583 ( .IN1(n4808), .IN2(n8382), .QN(n5251) );
  NAND2X0 U6584 ( .IN1(n5669), .IN2(n5670), .QN(WX8458) );
  NOR2X0 U6585 ( .IN1(n5671), .IN2(n5672), .QN(n5670) );
  NOR2X0 U6586 ( .IN1(n5673), .IN2(n4249), .QN(n5672) );
  NOR2X0 U6587 ( .IN1(n4340), .IN2(n5379), .QN(n5671) );
  XNOR2X1 U6588 ( .IN1(n5674), .IN2(n5675), .Q(n5379) );
  XOR2X1 U6589 ( .IN1(test_so81), .IN2(n8807), .Q(n5675) );
  XOR2X1 U6590 ( .IN1(WX9880), .IN2(n4017), .Q(n5674) );
  NOR2X0 U6591 ( .IN1(n5676), .IN2(n5677), .QN(n5669) );
  NOR2X0 U6592 ( .IN1(DFF_1315_n1), .IN2(n4285), .QN(n5677) );
  NOR2X0 U6593 ( .IN1(n4310), .IN2(n5252), .QN(n5676) );
  NAND2X0 U6594 ( .IN1(n4808), .IN2(n8383), .QN(n5252) );
  NAND2X0 U6595 ( .IN1(n5678), .IN2(n5679), .QN(WX8456) );
  NOR2X0 U6596 ( .IN1(n5680), .IN2(n5681), .QN(n5679) );
  NOR2X0 U6597 ( .IN1(n5682), .IN2(n4249), .QN(n5681) );
  NOR2X0 U6598 ( .IN1(n5387), .IN2(n4326), .QN(n5680) );
  XOR2X1 U6599 ( .IN1(n5683), .IN2(n5684), .Q(n5387) );
  XOR2X1 U6600 ( .IN1(n8808), .IN2(n3944), .Q(n5684) );
  XOR2X1 U6601 ( .IN1(WX9750), .IN2(n3732), .Q(n5683) );
  NOR2X0 U6602 ( .IN1(n5685), .IN2(n5686), .QN(n5678) );
  NOR2X0 U6603 ( .IN1(DFF_1316_n1), .IN2(n4285), .QN(n5686) );
  NOR2X0 U6604 ( .IN1(n4310), .IN2(n5253), .QN(n5685) );
  NAND2X0 U6605 ( .IN1(n4808), .IN2(n8384), .QN(n5253) );
  NAND2X0 U6606 ( .IN1(n5687), .IN2(n5688), .QN(WX8454) );
  NOR2X0 U6607 ( .IN1(n5689), .IN2(n5690), .QN(n5688) );
  NOR2X0 U6608 ( .IN1(n5691), .IN2(n4249), .QN(n5690) );
  NOR2X0 U6609 ( .IN1(n5395), .IN2(n4326), .QN(n5689) );
  XOR2X1 U6610 ( .IN1(n5692), .IN2(n5693), .Q(n5395) );
  XOR2X1 U6611 ( .IN1(n8809), .IN2(n4016), .Q(n5693) );
  XOR2X1 U6612 ( .IN1(WX9748), .IN2(n3734), .Q(n5692) );
  NOR2X0 U6613 ( .IN1(n5694), .IN2(n5695), .QN(n5687) );
  NOR2X0 U6614 ( .IN1(DFF_1317_n1), .IN2(n4284), .QN(n5695) );
  NOR2X0 U6615 ( .IN1(n4310), .IN2(n5254), .QN(n5694) );
  NAND2X0 U6616 ( .IN1(n4808), .IN2(n8385), .QN(n5254) );
  NAND2X0 U6617 ( .IN1(n5696), .IN2(n5697), .QN(WX8452) );
  NOR2X0 U6618 ( .IN1(n5698), .IN2(n5699), .QN(n5697) );
  NOR2X0 U6619 ( .IN1(n5700), .IN2(n4249), .QN(n5699) );
  NOR2X0 U6620 ( .IN1(n5403), .IN2(n4326), .QN(n5698) );
  XOR2X1 U6621 ( .IN1(n5701), .IN2(n5702), .Q(n5403) );
  XOR2X1 U6622 ( .IN1(n8810), .IN2(n4015), .Q(n5702) );
  XOR2X1 U6623 ( .IN1(WX9746), .IN2(n3736), .Q(n5701) );
  NOR2X0 U6624 ( .IN1(n5703), .IN2(n5704), .QN(n5696) );
  NOR2X0 U6625 ( .IN1(DFF_1318_n1), .IN2(n4284), .QN(n5704) );
  NOR2X0 U6626 ( .IN1(n4309), .IN2(n5255), .QN(n5703) );
  NAND2X0 U6627 ( .IN1(n4808), .IN2(n8386), .QN(n5255) );
  NAND2X0 U6628 ( .IN1(n5705), .IN2(n5706), .QN(WX8450) );
  NOR2X0 U6629 ( .IN1(n5707), .IN2(n5708), .QN(n5706) );
  NOR2X0 U6630 ( .IN1(n5709), .IN2(n4249), .QN(n5708) );
  NOR2X0 U6631 ( .IN1(n5411), .IN2(n4327), .QN(n5707) );
  XOR2X1 U6632 ( .IN1(n5710), .IN2(n5711), .Q(n5411) );
  XOR2X1 U6633 ( .IN1(n8811), .IN2(n4014), .Q(n5711) );
  XOR2X1 U6634 ( .IN1(WX9744), .IN2(n3738), .Q(n5710) );
  NOR2X0 U6635 ( .IN1(n5712), .IN2(n5713), .QN(n5705) );
  AND2X1 U6636 ( .IN1(n2152), .IN2(test_so76), .Q(n5713) );
  NOR2X0 U6637 ( .IN1(n4309), .IN2(n5256), .QN(n5712) );
  NAND2X0 U6638 ( .IN1(n4809), .IN2(n8387), .QN(n5256) );
  NAND2X0 U6639 ( .IN1(n5714), .IN2(n5715), .QN(WX8448) );
  NOR2X0 U6640 ( .IN1(n5716), .IN2(n5717), .QN(n5715) );
  NOR2X0 U6641 ( .IN1(n5718), .IN2(n4249), .QN(n5717) );
  NOR2X0 U6642 ( .IN1(n5419), .IN2(n4326), .QN(n5716) );
  XOR2X1 U6643 ( .IN1(n5719), .IN2(n5720), .Q(n5419) );
  XOR2X1 U6644 ( .IN1(n8812), .IN2(n4013), .Q(n5720) );
  XOR2X1 U6645 ( .IN1(WX9742), .IN2(n3740), .Q(n5719) );
  NOR2X0 U6646 ( .IN1(n5721), .IN2(n5722), .QN(n5714) );
  NOR2X0 U6647 ( .IN1(DFF_1320_n1), .IN2(n4284), .QN(n5722) );
  NOR2X0 U6648 ( .IN1(n4309), .IN2(n5258), .QN(n5721) );
  NAND2X0 U6649 ( .IN1(n4809), .IN2(n8388), .QN(n5258) );
  NAND2X0 U6650 ( .IN1(n5723), .IN2(n5724), .QN(WX8446) );
  NOR2X0 U6651 ( .IN1(n5725), .IN2(n5726), .QN(n5724) );
  NOR2X0 U6652 ( .IN1(n4259), .IN2(n5727), .QN(n5726) );
  NOR2X0 U6653 ( .IN1(n5427), .IN2(n4326), .QN(n5725) );
  XOR2X1 U6654 ( .IN1(n5728), .IN2(n5729), .Q(n5427) );
  XOR2X1 U6655 ( .IN1(n8813), .IN2(n4012), .Q(n5729) );
  XOR2X1 U6656 ( .IN1(WX9740), .IN2(n3742), .Q(n5728) );
  NOR2X0 U6657 ( .IN1(n5730), .IN2(n5731), .QN(n5723) );
  NOR2X0 U6658 ( .IN1(DFF_1321_n1), .IN2(n4284), .QN(n5731) );
  NOR2X0 U6659 ( .IN1(n4309), .IN2(n5259), .QN(n5730) );
  NAND2X0 U6660 ( .IN1(n4809), .IN2(n8389), .QN(n5259) );
  NAND2X0 U6661 ( .IN1(n5732), .IN2(n5733), .QN(WX8444) );
  NOR2X0 U6662 ( .IN1(n5734), .IN2(n5735), .QN(n5733) );
  NOR2X0 U6663 ( .IN1(n5736), .IN2(n4250), .QN(n5735) );
  NOR2X0 U6664 ( .IN1(n5435), .IN2(n4327), .QN(n5734) );
  XOR2X1 U6665 ( .IN1(n5737), .IN2(n5738), .Q(n5435) );
  XOR2X1 U6666 ( .IN1(n8814), .IN2(n4011), .Q(n5738) );
  XOR2X1 U6667 ( .IN1(WX9738), .IN2(n3744), .Q(n5737) );
  NOR2X0 U6668 ( .IN1(n5739), .IN2(n5740), .QN(n5732) );
  NOR2X0 U6669 ( .IN1(DFF_1322_n1), .IN2(n4284), .QN(n5740) );
  NOR2X0 U6670 ( .IN1(n4309), .IN2(n5260), .QN(n5739) );
  NAND2X0 U6671 ( .IN1(n4809), .IN2(n8390), .QN(n5260) );
  NAND2X0 U6672 ( .IN1(n5741), .IN2(n5742), .QN(WX8442) );
  NOR2X0 U6673 ( .IN1(n5743), .IN2(n5744), .QN(n5742) );
  NOR2X0 U6674 ( .IN1(n4259), .IN2(n5745), .QN(n5744) );
  NOR2X0 U6675 ( .IN1(n5443), .IN2(n4327), .QN(n5743) );
  XOR2X1 U6676 ( .IN1(n5746), .IN2(n5747), .Q(n5443) );
  XOR2X1 U6677 ( .IN1(n8815), .IN2(n3943), .Q(n5747) );
  XOR2X1 U6678 ( .IN1(WX9736), .IN2(n3746), .Q(n5746) );
  NOR2X0 U6679 ( .IN1(n5748), .IN2(n5749), .QN(n5741) );
  NOR2X0 U6680 ( .IN1(DFF_1323_n1), .IN2(n4284), .QN(n5749) );
  NOR2X0 U6681 ( .IN1(n4309), .IN2(n5261), .QN(n5748) );
  NAND2X0 U6682 ( .IN1(n4809), .IN2(n8391), .QN(n5261) );
  NAND2X0 U6683 ( .IN1(n5750), .IN2(n5751), .QN(WX8440) );
  NOR2X0 U6684 ( .IN1(n5752), .IN2(n5753), .QN(n5751) );
  NOR2X0 U6685 ( .IN1(n5754), .IN2(n4249), .QN(n5753) );
  NOR2X0 U6686 ( .IN1(n5451), .IN2(n4327), .QN(n5752) );
  XOR2X1 U6687 ( .IN1(n5755), .IN2(n5756), .Q(n5451) );
  XOR2X1 U6688 ( .IN1(n8816), .IN2(n4010), .Q(n5756) );
  XOR2X1 U6689 ( .IN1(WX9734), .IN2(n3748), .Q(n5755) );
  NOR2X0 U6690 ( .IN1(n5757), .IN2(n5758), .QN(n5750) );
  NOR2X0 U6691 ( .IN1(DFF_1324_n1), .IN2(n4284), .QN(n5758) );
  NOR2X0 U6692 ( .IN1(n4309), .IN2(n5262), .QN(n5757) );
  NAND2X0 U6693 ( .IN1(n4809), .IN2(n8392), .QN(n5262) );
  NAND2X0 U6694 ( .IN1(n5759), .IN2(n5760), .QN(WX8438) );
  NOR2X0 U6695 ( .IN1(n5761), .IN2(n5762), .QN(n5760) );
  NOR2X0 U6696 ( .IN1(n4259), .IN2(n5763), .QN(n5762) );
  NOR2X0 U6697 ( .IN1(n5459), .IN2(n4327), .QN(n5761) );
  XOR2X1 U6698 ( .IN1(n5764), .IN2(n5765), .Q(n5459) );
  XOR2X1 U6699 ( .IN1(n8817), .IN2(n4009), .Q(n5765) );
  XOR2X1 U6700 ( .IN1(WX9732), .IN2(n3750), .Q(n5764) );
  NOR2X0 U6701 ( .IN1(n5766), .IN2(n5767), .QN(n5759) );
  NOR2X0 U6702 ( .IN1(DFF_1325_n1), .IN2(n4284), .QN(n5767) );
  NOR2X0 U6703 ( .IN1(n4309), .IN2(n5263), .QN(n5766) );
  NAND2X0 U6704 ( .IN1(n4809), .IN2(n8393), .QN(n5263) );
  NAND2X0 U6705 ( .IN1(n5768), .IN2(n5769), .QN(WX8436) );
  NOR2X0 U6706 ( .IN1(n5770), .IN2(n5771), .QN(n5769) );
  NOR2X0 U6707 ( .IN1(n5772), .IN2(n4249), .QN(n5771) );
  NOR2X0 U6708 ( .IN1(n4339), .IN2(n5467), .QN(n5770) );
  XNOR2X1 U6709 ( .IN1(n5773), .IN2(n5774), .Q(n5467) );
  XOR2X1 U6710 ( .IN1(test_so86), .IN2(n8818), .Q(n5774) );
  XOR2X1 U6711 ( .IN1(WX9730), .IN2(n3752), .Q(n5773) );
  NOR2X0 U6712 ( .IN1(n5775), .IN2(n5776), .QN(n5768) );
  NOR2X0 U6713 ( .IN1(DFF_1326_n1), .IN2(n4284), .QN(n5776) );
  NOR2X0 U6714 ( .IN1(n4309), .IN2(n5264), .QN(n5775) );
  NAND2X0 U6715 ( .IN1(n4809), .IN2(n8394), .QN(n5264) );
  NAND2X0 U6716 ( .IN1(n5777), .IN2(n5778), .QN(WX8434) );
  NOR2X0 U6717 ( .IN1(n5779), .IN2(n5780), .QN(n5778) );
  NOR2X0 U6718 ( .IN1(n4259), .IN2(n5781), .QN(n5780) );
  NOR2X0 U6719 ( .IN1(n5475), .IN2(n4327), .QN(n5779) );
  XOR2X1 U6720 ( .IN1(n5782), .IN2(n5783), .Q(n5475) );
  XOR2X1 U6721 ( .IN1(n8819), .IN2(n4008), .Q(n5783) );
  XOR2X1 U6722 ( .IN1(WX9728), .IN2(n3754), .Q(n5782) );
  NOR2X0 U6723 ( .IN1(n5784), .IN2(n5785), .QN(n5777) );
  NOR2X0 U6724 ( .IN1(DFF_1327_n1), .IN2(n4284), .QN(n5785) );
  NOR2X0 U6725 ( .IN1(n4309), .IN2(n5265), .QN(n5784) );
  NAND2X0 U6726 ( .IN1(n4809), .IN2(n8395), .QN(n5265) );
  NAND2X0 U6727 ( .IN1(n5786), .IN2(n5787), .QN(WX8432) );
  NOR2X0 U6728 ( .IN1(n5788), .IN2(n5789), .QN(n5787) );
  NOR2X0 U6729 ( .IN1(n5790), .IN2(n4249), .QN(n5789) );
  NOR2X0 U6730 ( .IN1(n4339), .IN2(n5483), .QN(n5788) );
  XNOR2X1 U6731 ( .IN1(n5791), .IN2(n5792), .Q(n5483) );
  XOR2X1 U6732 ( .IN1(n3942), .IN2(n4771), .Q(n5792) );
  XOR2X1 U6733 ( .IN1(n5793), .IN2(n8822), .Q(n5791) );
  XOR2X1 U6734 ( .IN1(n8821), .IN2(n8820), .Q(n5793) );
  NOR2X0 U6735 ( .IN1(n5794), .IN2(n5795), .QN(n5786) );
  NOR2X0 U6736 ( .IN1(DFF_1328_n1), .IN2(n4284), .QN(n5795) );
  NOR2X0 U6737 ( .IN1(n4309), .IN2(n5266), .QN(n5794) );
  NAND2X0 U6738 ( .IN1(n4810), .IN2(n8396), .QN(n5266) );
  NAND2X0 U6739 ( .IN1(n5796), .IN2(n5797), .QN(WX8430) );
  NOR2X0 U6740 ( .IN1(n5798), .IN2(n5799), .QN(n5797) );
  NOR2X0 U6741 ( .IN1(n5800), .IN2(n4250), .QN(n5799) );
  NOR2X0 U6742 ( .IN1(n5491), .IN2(n4327), .QN(n5798) );
  XOR2X1 U6743 ( .IN1(n5801), .IN2(n5802), .Q(n5491) );
  XOR2X1 U6744 ( .IN1(n3603), .IN2(n4771), .Q(n5802) );
  XOR2X1 U6745 ( .IN1(n5803), .IN2(n4007), .Q(n5801) );
  XOR2X1 U6746 ( .IN1(WX9852), .IN2(n8823), .Q(n5803) );
  NOR2X0 U6747 ( .IN1(n5804), .IN2(n5805), .QN(n5796) );
  NOR2X0 U6748 ( .IN1(DFF_1329_n1), .IN2(n4284), .QN(n5805) );
  NOR2X0 U6749 ( .IN1(n4309), .IN2(n5267), .QN(n5804) );
  NAND2X0 U6750 ( .IN1(test_so67), .IN2(n4828), .QN(n5267) );
  NAND2X0 U6751 ( .IN1(n5806), .IN2(n5807), .QN(WX8428) );
  NOR2X0 U6752 ( .IN1(n5808), .IN2(n5809), .QN(n5807) );
  NOR2X0 U6753 ( .IN1(n5810), .IN2(n4249), .QN(n5809) );
  NOR2X0 U6754 ( .IN1(n4339), .IN2(n5499), .QN(n5808) );
  XNOR2X1 U6755 ( .IN1(n5811), .IN2(n5812), .Q(n5499) );
  XOR2X1 U6756 ( .IN1(n4006), .IN2(n4771), .Q(n5812) );
  XOR2X1 U6757 ( .IN1(n5813), .IN2(n8826), .Q(n5811) );
  XOR2X1 U6758 ( .IN1(n8825), .IN2(n8824), .Q(n5813) );
  NOR2X0 U6759 ( .IN1(n5814), .IN2(n5815), .QN(n5806) );
  NOR2X0 U6760 ( .IN1(DFF_1330_n1), .IN2(n4284), .QN(n5815) );
  NOR2X0 U6761 ( .IN1(n4308), .IN2(n5269), .QN(n5814) );
  NAND2X0 U6762 ( .IN1(n4810), .IN2(n8399), .QN(n5269) );
  NAND2X0 U6763 ( .IN1(n5816), .IN2(n5817), .QN(WX8426) );
  NOR2X0 U6764 ( .IN1(n5818), .IN2(n5819), .QN(n5817) );
  NOR2X0 U6765 ( .IN1(n5820), .IN2(n4249), .QN(n5819) );
  NOR2X0 U6766 ( .IN1(n5507), .IN2(n4327), .QN(n5818) );
  XOR2X1 U6767 ( .IN1(n5821), .IN2(n5822), .Q(n5507) );
  XOR2X1 U6768 ( .IN1(n3604), .IN2(n4771), .Q(n5822) );
  XOR2X1 U6769 ( .IN1(n5823), .IN2(n4005), .Q(n5821) );
  XOR2X1 U6770 ( .IN1(WX9848), .IN2(n8827), .Q(n5823) );
  NOR2X0 U6771 ( .IN1(n5824), .IN2(n5825), .QN(n5816) );
  NOR2X0 U6772 ( .IN1(DFF_1331_n1), .IN2(n4284), .QN(n5825) );
  NOR2X0 U6773 ( .IN1(n4308), .IN2(n5270), .QN(n5824) );
  NAND2X0 U6774 ( .IN1(n4810), .IN2(n8400), .QN(n5270) );
  NAND2X0 U6775 ( .IN1(n5826), .IN2(n5827), .QN(WX8424) );
  NOR2X0 U6776 ( .IN1(n5828), .IN2(n5829), .QN(n5827) );
  NOR2X0 U6777 ( .IN1(n5830), .IN2(n4250), .QN(n5829) );
  NOR2X0 U6778 ( .IN1(n4339), .IN2(n5515), .QN(n5828) );
  XNOR2X1 U6779 ( .IN1(n5831), .IN2(n5832), .Q(n5515) );
  XOR2X1 U6780 ( .IN1(n3605), .IN2(n4771), .Q(n5832) );
  XOR2X1 U6781 ( .IN1(n5833), .IN2(n4004), .Q(n5831) );
  XOR2X1 U6782 ( .IN1(WX9782), .IN2(test_so80), .Q(n5833) );
  NOR2X0 U6783 ( .IN1(n5834), .IN2(n5835), .QN(n5826) );
  NOR2X0 U6784 ( .IN1(DFF_1332_n1), .IN2(n4283), .QN(n5835) );
  NOR2X0 U6785 ( .IN1(n4308), .IN2(n5271), .QN(n5834) );
  NAND2X0 U6786 ( .IN1(n4810), .IN2(n8401), .QN(n5271) );
  NAND2X0 U6787 ( .IN1(n5836), .IN2(n5837), .QN(WX8422) );
  NOR2X0 U6788 ( .IN1(n5838), .IN2(n5839), .QN(n5837) );
  NOR2X0 U6789 ( .IN1(n5840), .IN2(n4250), .QN(n5839) );
  NOR2X0 U6790 ( .IN1(n5523), .IN2(n4327), .QN(n5838) );
  XOR2X1 U6791 ( .IN1(n5841), .IN2(n5842), .Q(n5523) );
  XOR2X1 U6792 ( .IN1(n3606), .IN2(n4771), .Q(n5842) );
  XOR2X1 U6793 ( .IN1(n5843), .IN2(n4003), .Q(n5841) );
  XOR2X1 U6794 ( .IN1(WX9844), .IN2(n8828), .Q(n5843) );
  NOR2X0 U6795 ( .IN1(n5844), .IN2(n5845), .QN(n5836) );
  NOR2X0 U6796 ( .IN1(DFF_1333_n1), .IN2(n4283), .QN(n5845) );
  NOR2X0 U6797 ( .IN1(n4308), .IN2(n5272), .QN(n5844) );
  NAND2X0 U6798 ( .IN1(n4810), .IN2(n8402), .QN(n5272) );
  NAND2X0 U6799 ( .IN1(n5846), .IN2(n5847), .QN(WX8420) );
  NOR2X0 U6800 ( .IN1(n5848), .IN2(n5849), .QN(n5847) );
  NOR2X0 U6801 ( .IN1(n5850), .IN2(n4250), .QN(n5849) );
  NOR2X0 U6802 ( .IN1(n5531), .IN2(n4328), .QN(n5848) );
  XOR2X1 U6803 ( .IN1(n5851), .IN2(n5852), .Q(n5531) );
  XOR2X1 U6804 ( .IN1(n3607), .IN2(n4771), .Q(n5852) );
  XOR2X1 U6805 ( .IN1(n5853), .IN2(n4002), .Q(n5851) );
  XOR2X1 U6806 ( .IN1(WX9842), .IN2(n8829), .Q(n5853) );
  NOR2X0 U6807 ( .IN1(n5854), .IN2(n5855), .QN(n5846) );
  NOR2X0 U6808 ( .IN1(DFF_1334_n1), .IN2(n4283), .QN(n5855) );
  NOR2X0 U6809 ( .IN1(n4308), .IN2(n5273), .QN(n5854) );
  NAND2X0 U6810 ( .IN1(n4810), .IN2(n8403), .QN(n5273) );
  NAND2X0 U6811 ( .IN1(n5856), .IN2(n5857), .QN(WX8418) );
  NOR2X0 U6812 ( .IN1(n5858), .IN2(n5859), .QN(n5857) );
  NOR2X0 U6813 ( .IN1(n5860), .IN2(n4250), .QN(n5859) );
  NOR2X0 U6814 ( .IN1(n5539), .IN2(n4328), .QN(n5858) );
  XOR2X1 U6815 ( .IN1(n5861), .IN2(n5862), .Q(n5539) );
  XOR2X1 U6816 ( .IN1(n3608), .IN2(n4771), .Q(n5862) );
  XOR2X1 U6817 ( .IN1(n5863), .IN2(n4001), .Q(n5861) );
  XOR2X1 U6818 ( .IN1(WX9840), .IN2(n8830), .Q(n5863) );
  NOR2X0 U6819 ( .IN1(n5864), .IN2(n5865), .QN(n5856) );
  NOR2X0 U6820 ( .IN1(DFF_1335_n1), .IN2(n4283), .QN(n5865) );
  NOR2X0 U6821 ( .IN1(n4308), .IN2(n5274), .QN(n5864) );
  NAND2X0 U6822 ( .IN1(n4810), .IN2(n8404), .QN(n5274) );
  NAND2X0 U6823 ( .IN1(n5866), .IN2(n5867), .QN(WX8416) );
  NOR2X0 U6824 ( .IN1(n5868), .IN2(n5869), .QN(n5867) );
  NOR2X0 U6825 ( .IN1(n5870), .IN2(n4250), .QN(n5869) );
  NOR2X0 U6826 ( .IN1(n5547), .IN2(n4329), .QN(n5868) );
  XOR2X1 U6827 ( .IN1(n5871), .IN2(n5872), .Q(n5547) );
  XOR2X1 U6828 ( .IN1(n3609), .IN2(n4771), .Q(n5872) );
  XOR2X1 U6829 ( .IN1(n5873), .IN2(n4000), .Q(n5871) );
  XOR2X1 U6830 ( .IN1(WX9838), .IN2(n8831), .Q(n5873) );
  NOR2X0 U6831 ( .IN1(n5874), .IN2(n5875), .QN(n5866) );
  AND2X1 U6832 ( .IN1(n2152), .IN2(test_so77), .Q(n5875) );
  NOR2X0 U6833 ( .IN1(n4308), .IN2(n5275), .QN(n5874) );
  NAND2X0 U6834 ( .IN1(n4810), .IN2(n8405), .QN(n5275) );
  NAND2X0 U6835 ( .IN1(n5876), .IN2(n5877), .QN(WX8414) );
  NOR2X0 U6836 ( .IN1(n5878), .IN2(n5879), .QN(n5877) );
  NOR2X0 U6837 ( .IN1(n5880), .IN2(n4250), .QN(n5879) );
  NOR2X0 U6838 ( .IN1(n5555), .IN2(n4327), .QN(n5878) );
  XOR2X1 U6839 ( .IN1(n5881), .IN2(n5882), .Q(n5555) );
  XOR2X1 U6840 ( .IN1(n3610), .IN2(n4771), .Q(n5882) );
  XOR2X1 U6841 ( .IN1(n5883), .IN2(n3999), .Q(n5881) );
  XOR2X1 U6842 ( .IN1(WX9836), .IN2(n8832), .Q(n5883) );
  NOR2X0 U6843 ( .IN1(n5884), .IN2(n5885), .QN(n5876) );
  NOR2X0 U6844 ( .IN1(DFF_1337_n1), .IN2(n4283), .QN(n5885) );
  NOR2X0 U6845 ( .IN1(n4308), .IN2(n5276), .QN(n5884) );
  NAND2X0 U6846 ( .IN1(n4810), .IN2(n8406), .QN(n5276) );
  NAND2X0 U6847 ( .IN1(n5886), .IN2(n5887), .QN(WX8412) );
  NOR2X0 U6848 ( .IN1(n5888), .IN2(n5889), .QN(n5887) );
  NOR2X0 U6849 ( .IN1(n4260), .IN2(n5890), .QN(n5889) );
  NOR2X0 U6850 ( .IN1(n5563), .IN2(n4328), .QN(n5888) );
  XOR2X1 U6851 ( .IN1(n5891), .IN2(n5892), .Q(n5563) );
  XOR2X1 U6852 ( .IN1(n3611), .IN2(n4771), .Q(n5892) );
  XOR2X1 U6853 ( .IN1(n5893), .IN2(n3998), .Q(n5891) );
  XOR2X1 U6854 ( .IN1(WX9834), .IN2(n8833), .Q(n5893) );
  NOR2X0 U6855 ( .IN1(n5894), .IN2(n5895), .QN(n5886) );
  NOR2X0 U6856 ( .IN1(DFF_1338_n1), .IN2(n4283), .QN(n5895) );
  NOR2X0 U6857 ( .IN1(n4308), .IN2(n5277), .QN(n5894) );
  NAND2X0 U6858 ( .IN1(n4824), .IN2(n8407), .QN(n5277) );
  NAND2X0 U6859 ( .IN1(n5896), .IN2(n5897), .QN(WX8410) );
  NOR2X0 U6860 ( .IN1(n5898), .IN2(n5899), .QN(n5897) );
  NOR2X0 U6861 ( .IN1(n5900), .IN2(n4250), .QN(n5899) );
  NOR2X0 U6862 ( .IN1(n5571), .IN2(n4327), .QN(n5898) );
  XOR2X1 U6863 ( .IN1(n5901), .IN2(n5902), .Q(n5571) );
  XOR2X1 U6864 ( .IN1(n3612), .IN2(n4772), .Q(n5902) );
  XOR2X1 U6865 ( .IN1(n5903), .IN2(n3997), .Q(n5901) );
  XOR2X1 U6866 ( .IN1(WX9832), .IN2(n8834), .Q(n5903) );
  NOR2X0 U6867 ( .IN1(n5904), .IN2(n5905), .QN(n5896) );
  NOR2X0 U6868 ( .IN1(DFF_1339_n1), .IN2(n4283), .QN(n5905) );
  NOR2X0 U6869 ( .IN1(n4308), .IN2(n5278), .QN(n5904) );
  NAND2X0 U6870 ( .IN1(n4827), .IN2(n8408), .QN(n5278) );
  NAND2X0 U6871 ( .IN1(n5906), .IN2(n5907), .QN(WX8408) );
  NOR2X0 U6872 ( .IN1(n5908), .IN2(n5909), .QN(n5907) );
  NOR2X0 U6873 ( .IN1(n4260), .IN2(n5910), .QN(n5909) );
  NOR2X0 U6874 ( .IN1(n5579), .IN2(n4327), .QN(n5908) );
  XOR2X1 U6875 ( .IN1(n5911), .IN2(n5912), .Q(n5579) );
  XOR2X1 U6876 ( .IN1(n3613), .IN2(n4772), .Q(n5912) );
  XOR2X1 U6877 ( .IN1(n5913), .IN2(n3996), .Q(n5911) );
  XOR2X1 U6878 ( .IN1(WX9830), .IN2(n8835), .Q(n5913) );
  NOR2X0 U6879 ( .IN1(n5914), .IN2(n5915), .QN(n5906) );
  NOR2X0 U6880 ( .IN1(DFF_1340_n1), .IN2(n4283), .QN(n5915) );
  NOR2X0 U6881 ( .IN1(n4308), .IN2(n5280), .QN(n5914) );
  NAND2X0 U6882 ( .IN1(n4827), .IN2(n8409), .QN(n5280) );
  NAND2X0 U6883 ( .IN1(n5916), .IN2(n5917), .QN(WX8406) );
  NOR2X0 U6884 ( .IN1(n5918), .IN2(n5919), .QN(n5917) );
  NOR2X0 U6885 ( .IN1(n5920), .IN2(n4250), .QN(n5919) );
  NOR2X0 U6886 ( .IN1(n5587), .IN2(n4328), .QN(n5918) );
  XOR2X1 U6887 ( .IN1(n5921), .IN2(n5922), .Q(n5587) );
  XOR2X1 U6888 ( .IN1(n3614), .IN2(n4772), .Q(n5922) );
  XOR2X1 U6889 ( .IN1(n5923), .IN2(n3995), .Q(n5921) );
  XOR2X1 U6890 ( .IN1(WX9828), .IN2(n8836), .Q(n5923) );
  NOR2X0 U6891 ( .IN1(n5924), .IN2(n5925), .QN(n5916) );
  NOR2X0 U6892 ( .IN1(DFF_1341_n1), .IN2(n4283), .QN(n5925) );
  NOR2X0 U6893 ( .IN1(n4308), .IN2(n5281), .QN(n5924) );
  NAND2X0 U6894 ( .IN1(n4827), .IN2(n8410), .QN(n5281) );
  NAND2X0 U6895 ( .IN1(n5926), .IN2(n5927), .QN(WX8404) );
  NOR2X0 U6896 ( .IN1(n5928), .IN2(n5929), .QN(n5927) );
  NOR2X0 U6897 ( .IN1(n4260), .IN2(n5930), .QN(n5929) );
  NOR2X0 U6898 ( .IN1(n5595), .IN2(n4328), .QN(n5928) );
  XOR2X1 U6899 ( .IN1(n5931), .IN2(n5932), .Q(n5595) );
  XOR2X1 U6900 ( .IN1(n3615), .IN2(n4772), .Q(n5932) );
  XOR2X1 U6901 ( .IN1(n5933), .IN2(n3994), .Q(n5931) );
  XOR2X1 U6902 ( .IN1(WX9826), .IN2(n8837), .Q(n5933) );
  NOR2X0 U6903 ( .IN1(n5934), .IN2(n5935), .QN(n5926) );
  NOR2X0 U6904 ( .IN1(DFF_1342_n1), .IN2(n4283), .QN(n5935) );
  NOR2X0 U6905 ( .IN1(n5356), .IN2(n5282), .QN(n5934) );
  NAND2X0 U6906 ( .IN1(n4827), .IN2(n8411), .QN(n5282) );
  NAND2X0 U6907 ( .IN1(n5936), .IN2(n5937), .QN(WX8402) );
  NOR2X0 U6908 ( .IN1(n5938), .IN2(n5939), .QN(n5937) );
  NOR2X0 U6909 ( .IN1(n5940), .IN2(n4250), .QN(n5939) );
  NOR2X0 U6910 ( .IN1(n4338), .IN2(n5603), .QN(n5938) );
  XNOR2X1 U6911 ( .IN1(n5941), .IN2(n5942), .Q(n5603) );
  XOR2X1 U6912 ( .IN1(n3583), .IN2(n4772), .Q(n5942) );
  XOR2X1 U6913 ( .IN1(WX9760), .IN2(n5943), .Q(n5941) );
  XOR2X1 U6914 ( .IN1(test_so85), .IN2(n8838), .Q(n5943) );
  NOR2X0 U6915 ( .IN1(n5944), .IN2(n5945), .QN(n5936) );
  NOR2X0 U6916 ( .IN1(n3933), .IN2(n5606), .QN(n5945) );
  NOR2X0 U6917 ( .IN1(DFF_1343_n1), .IN2(n4283), .QN(n5944) );
  AND2X1 U6918 ( .IN1(n4800), .IN2(n3933), .Q(WX8304) );
  NOR2X0 U6919 ( .IN1(n4936), .IN2(n5946), .QN(WX7791) );
  XOR2X1 U6920 ( .IN1(n4046), .IN2(DFF_1150_n1), .Q(n5946) );
  NOR2X0 U6921 ( .IN1(n4936), .IN2(n5947), .QN(WX7789) );
  XNOR2X1 U6922 ( .IN1(n4047), .IN2(test_so66), .Q(n5947) );
  NOR2X0 U6923 ( .IN1(n4936), .IN2(n5948), .QN(WX7787) );
  XOR2X1 U6924 ( .IN1(n4048), .IN2(DFF_1148_n1), .Q(n5948) );
  NOR2X0 U6925 ( .IN1(n4936), .IN2(n5949), .QN(WX7785) );
  XOR2X1 U6926 ( .IN1(n4049), .IN2(DFF_1147_n1), .Q(n5949) );
  NOR2X0 U6927 ( .IN1(n4936), .IN2(n5950), .QN(WX7783) );
  XOR2X1 U6928 ( .IN1(n4050), .IN2(DFF_1146_n1), .Q(n5950) );
  NOR2X0 U6929 ( .IN1(n4936), .IN2(n5951), .QN(WX7781) );
  XOR2X1 U6930 ( .IN1(n4051), .IN2(DFF_1145_n1), .Q(n5951) );
  NOR2X0 U6931 ( .IN1(n4936), .IN2(n5952), .QN(WX7779) );
  XOR2X1 U6932 ( .IN1(n4052), .IN2(DFF_1144_n1), .Q(n5952) );
  NOR2X0 U6933 ( .IN1(n4936), .IN2(n5953), .QN(WX7777) );
  XOR2X1 U6934 ( .IN1(n4053), .IN2(DFF_1143_n1), .Q(n5953) );
  NOR2X0 U6935 ( .IN1(n4936), .IN2(n5954), .QN(WX7775) );
  XOR2X1 U6936 ( .IN1(n4054), .IN2(DFF_1142_n1), .Q(n5954) );
  NOR2X0 U6937 ( .IN1(n4937), .IN2(n5955), .QN(WX7773) );
  XOR2X1 U6938 ( .IN1(n4055), .IN2(DFF_1141_n1), .Q(n5955) );
  NOR2X0 U6939 ( .IN1(n4937), .IN2(n5956), .QN(WX7771) );
  XNOR2X1 U6940 ( .IN1(DFF_1140_n1), .IN2(test_so63), .Q(n5956) );
  NOR2X0 U6941 ( .IN1(n4937), .IN2(n5957), .QN(WX7769) );
  XOR2X1 U6942 ( .IN1(n4056), .IN2(DFF_1139_n1), .Q(n5957) );
  NOR2X0 U6943 ( .IN1(n4937), .IN2(n5958), .QN(WX7767) );
  XOR2X1 U6944 ( .IN1(n4057), .IN2(DFF_1138_n1), .Q(n5958) );
  NOR2X0 U6945 ( .IN1(n4937), .IN2(n5959), .QN(WX7765) );
  XOR2X1 U6946 ( .IN1(n4058), .IN2(DFF_1137_n1), .Q(n5959) );
  NOR2X0 U6947 ( .IN1(n4937), .IN2(n5960), .QN(WX7763) );
  XOR2X1 U6948 ( .IN1(n4059), .IN2(DFF_1136_n1), .Q(n5960) );
  NOR2X0 U6949 ( .IN1(n4937), .IN2(n5961), .QN(WX7761) );
  XNOR2X1 U6950 ( .IN1(DFF_1135_n1), .IN2(n5962), .Q(n5961) );
  XOR2X1 U6951 ( .IN1(n3948), .IN2(DFF_1151_n1), .Q(n5962) );
  NOR2X0 U6952 ( .IN1(n4937), .IN2(n5963), .QN(WX7759) );
  XOR2X1 U6953 ( .IN1(n4060), .IN2(DFF_1134_n1), .Q(n5963) );
  NOR2X0 U6954 ( .IN1(n4937), .IN2(n5964), .QN(WX7757) );
  XOR2X1 U6955 ( .IN1(n4061), .IN2(DFF_1133_n1), .Q(n5964) );
  NOR2X0 U6956 ( .IN1(n4937), .IN2(n5965), .QN(WX7755) );
  XNOR2X1 U6957 ( .IN1(n4062), .IN2(test_so65), .Q(n5965) );
  NOR2X0 U6958 ( .IN1(n4937), .IN2(n5966), .QN(WX7753) );
  XOR2X1 U6959 ( .IN1(n4063), .IN2(DFF_1131_n1), .Q(n5966) );
  NOR2X0 U6960 ( .IN1(n4937), .IN2(n5967), .QN(WX7751) );
  XNOR2X1 U6961 ( .IN1(DFF_1130_n1), .IN2(n5968), .Q(n5967) );
  XOR2X1 U6962 ( .IN1(n3949), .IN2(DFF_1151_n1), .Q(n5968) );
  NOR2X0 U6963 ( .IN1(n4937), .IN2(n5969), .QN(WX7749) );
  XOR2X1 U6964 ( .IN1(n4064), .IN2(DFF_1129_n1), .Q(n5969) );
  NOR2X0 U6965 ( .IN1(n4938), .IN2(n5970), .QN(WX7747) );
  XOR2X1 U6966 ( .IN1(n4065), .IN2(DFF_1128_n1), .Q(n5970) );
  NOR2X0 U6967 ( .IN1(n4938), .IN2(n5971), .QN(WX7745) );
  XOR2X1 U6968 ( .IN1(n4066), .IN2(DFF_1127_n1), .Q(n5971) );
  NOR2X0 U6969 ( .IN1(n4938), .IN2(n5972), .QN(WX7743) );
  XOR2X1 U6970 ( .IN1(n4067), .IN2(DFF_1126_n1), .Q(n5972) );
  NOR2X0 U6971 ( .IN1(n4938), .IN2(n5973), .QN(WX7741) );
  XOR2X1 U6972 ( .IN1(n4068), .IN2(DFF_1125_n1), .Q(n5973) );
  NOR2X0 U6973 ( .IN1(n4938), .IN2(n5974), .QN(WX7739) );
  XOR2X1 U6974 ( .IN1(n4069), .IN2(DFF_1124_n1), .Q(n5974) );
  NOR2X0 U6975 ( .IN1(n4938), .IN2(n5975), .QN(WX7737) );
  XOR2X1 U6976 ( .IN1(DFF_1123_n1), .IN2(n5976), .Q(n5975) );
  XOR2X1 U6977 ( .IN1(test_so64), .IN2(DFF_1151_n1), .Q(n5976) );
  NOR2X0 U6978 ( .IN1(n4938), .IN2(n5977), .QN(WX7735) );
  XOR2X1 U6979 ( .IN1(n4070), .IN2(DFF_1122_n1), .Q(n5977) );
  NOR2X0 U6980 ( .IN1(n4938), .IN2(n5978), .QN(WX7733) );
  XOR2X1 U6981 ( .IN1(n4071), .IN2(DFF_1121_n1), .Q(n5978) );
  NOR2X0 U6982 ( .IN1(n4938), .IN2(n5979), .QN(WX7731) );
  XOR2X1 U6983 ( .IN1(n4072), .IN2(DFF_1120_n1), .Q(n5979) );
  NOR2X0 U6984 ( .IN1(n4938), .IN2(n5980), .QN(WX7729) );
  XOR2X1 U6985 ( .IN1(n3963), .IN2(DFF_1151_n1), .Q(n5980) );
  NOR2X0 U6986 ( .IN1(n8891), .IN2(n4850), .QN(WX7203) );
  NOR2X0 U6987 ( .IN1(n8892), .IN2(n4850), .QN(WX7201) );
  NOR2X0 U6988 ( .IN1(n8893), .IN2(n4850), .QN(WX7199) );
  NOR2X0 U6989 ( .IN1(n8894), .IN2(n4850), .QN(WX7197) );
  NOR2X0 U6990 ( .IN1(n8895), .IN2(n4851), .QN(WX7195) );
  NOR2X0 U6991 ( .IN1(n8896), .IN2(n4851), .QN(WX7193) );
  NOR2X0 U6992 ( .IN1(n8897), .IN2(n4851), .QN(WX7191) );
  NOR2X0 U6993 ( .IN1(n8898), .IN2(n4851), .QN(WX7189) );
  NOR2X0 U6994 ( .IN1(n8901), .IN2(n4851), .QN(WX7187) );
  NOR2X0 U6995 ( .IN1(n8902), .IN2(n4851), .QN(WX7185) );
  NOR2X0 U6996 ( .IN1(n8905), .IN2(n4851), .QN(WX7183) );
  AND2X1 U6997 ( .IN1(n4800), .IN2(test_so57), .Q(WX7181) );
  NOR2X0 U6998 ( .IN1(n8906), .IN2(n4851), .QN(WX7179) );
  NOR2X0 U6999 ( .IN1(n8907), .IN2(n4851), .QN(WX7177) );
  NOR2X0 U7000 ( .IN1(n8908), .IN2(n4851), .QN(WX7175) );
  NOR2X0 U7001 ( .IN1(n8909), .IN2(n4851), .QN(WX7173) );
  NAND2X0 U7002 ( .IN1(n5981), .IN2(n5982), .QN(WX7171) );
  NOR2X0 U7003 ( .IN1(n5983), .IN2(n5984), .QN(n5982) );
  NOR2X0 U7004 ( .IN1(n5985), .IN2(n4251), .QN(n5984) );
  NOR2X0 U7005 ( .IN1(n5646), .IN2(n4328), .QN(n5983) );
  XOR2X1 U7006 ( .IN1(n5986), .IN2(n5987), .Q(n5646) );
  XOR2X1 U7007 ( .IN1(n8839), .IN2(n3962), .Q(n5987) );
  XOR2X1 U7008 ( .IN1(WX8465), .IN2(n3756), .Q(n5986) );
  NOR2X0 U7009 ( .IN1(n5988), .IN2(n5989), .QN(n5981) );
  NOR2X0 U7010 ( .IN1(DFF_1120_n1), .IN2(n4283), .QN(n5989) );
  NOR2X0 U7011 ( .IN1(n5356), .IN2(n5283), .QN(n5988) );
  NAND2X0 U7012 ( .IN1(n4826), .IN2(n8438), .QN(n5283) );
  NAND2X0 U7013 ( .IN1(n5990), .IN2(n5991), .QN(WX7169) );
  NOR2X0 U7014 ( .IN1(n5992), .IN2(n5993), .QN(n5991) );
  NOR2X0 U7015 ( .IN1(n5994), .IN2(n4250), .QN(n5993) );
  NOR2X0 U7016 ( .IN1(n5655), .IN2(n4328), .QN(n5992) );
  XOR2X1 U7017 ( .IN1(n5995), .IN2(n5996), .Q(n5655) );
  XOR2X1 U7018 ( .IN1(n8840), .IN2(n4045), .Q(n5996) );
  XOR2X1 U7019 ( .IN1(WX8463), .IN2(n3758), .Q(n5995) );
  NOR2X0 U7020 ( .IN1(n5997), .IN2(n5998), .QN(n5990) );
  NOR2X0 U7021 ( .IN1(DFF_1121_n1), .IN2(n4283), .QN(n5998) );
  NOR2X0 U7022 ( .IN1(n5356), .IN2(n5284), .QN(n5997) );
  NAND2X0 U7023 ( .IN1(n4824), .IN2(n8439), .QN(n5284) );
  NAND2X0 U7024 ( .IN1(n5999), .IN2(n6000), .QN(WX7167) );
  NOR2X0 U7025 ( .IN1(n6001), .IN2(n6002), .QN(n6000) );
  NOR2X0 U7026 ( .IN1(n6003), .IN2(n4250), .QN(n6002) );
  NOR2X0 U7027 ( .IN1(n5664), .IN2(n4328), .QN(n6001) );
  XOR2X1 U7028 ( .IN1(n6004), .IN2(n6005), .Q(n5664) );
  XOR2X1 U7029 ( .IN1(n8841), .IN2(n4044), .Q(n6005) );
  XOR2X1 U7030 ( .IN1(WX8461), .IN2(n3760), .Q(n6004) );
  NOR2X0 U7031 ( .IN1(n6006), .IN2(n6007), .QN(n5999) );
  NOR2X0 U7032 ( .IN1(DFF_1122_n1), .IN2(n4282), .QN(n6007) );
  NOR2X0 U7033 ( .IN1(n5356), .IN2(n5285), .QN(n6006) );
  NAND2X0 U7034 ( .IN1(n4827), .IN2(n8440), .QN(n5285) );
  NAND2X0 U7035 ( .IN1(n6008), .IN2(n6009), .QN(WX7165) );
  NOR2X0 U7036 ( .IN1(n6010), .IN2(n6011), .QN(n6009) );
  NOR2X0 U7037 ( .IN1(n6012), .IN2(n4250), .QN(n6011) );
  NOR2X0 U7038 ( .IN1(n5673), .IN2(n4328), .QN(n6010) );
  XOR2X1 U7039 ( .IN1(n6013), .IN2(n6014), .Q(n5673) );
  XOR2X1 U7040 ( .IN1(n8842), .IN2(n4043), .Q(n6014) );
  XOR2X1 U7041 ( .IN1(WX8459), .IN2(n3762), .Q(n6013) );
  NOR2X0 U7042 ( .IN1(n6015), .IN2(n6016), .QN(n6008) );
  NOR2X0 U7043 ( .IN1(DFF_1123_n1), .IN2(n4282), .QN(n6016) );
  NOR2X0 U7044 ( .IN1(n5356), .IN2(n5286), .QN(n6015) );
  NAND2X0 U7045 ( .IN1(n4826), .IN2(n8441), .QN(n5286) );
  NAND2X0 U7046 ( .IN1(n6017), .IN2(n6018), .QN(WX7163) );
  NOR2X0 U7047 ( .IN1(n6019), .IN2(n6020), .QN(n6018) );
  NOR2X0 U7048 ( .IN1(n4260), .IN2(n6021), .QN(n6020) );
  NOR2X0 U7049 ( .IN1(n5682), .IN2(n4329), .QN(n6019) );
  XOR2X1 U7050 ( .IN1(n6022), .IN2(n6023), .Q(n5682) );
  XOR2X1 U7051 ( .IN1(n8843), .IN2(n3947), .Q(n6023) );
  XOR2X1 U7052 ( .IN1(WX8457), .IN2(n3764), .Q(n6022) );
  NOR2X0 U7053 ( .IN1(n6024), .IN2(n6025), .QN(n6017) );
  NOR2X0 U7054 ( .IN1(DFF_1124_n1), .IN2(n4282), .QN(n6025) );
  NOR2X0 U7055 ( .IN1(n5356), .IN2(n5287), .QN(n6024) );
  NAND2X0 U7056 ( .IN1(n4826), .IN2(n8442), .QN(n5287) );
  NAND2X0 U7057 ( .IN1(n6026), .IN2(n6027), .QN(WX7161) );
  NOR2X0 U7058 ( .IN1(n6028), .IN2(n6029), .QN(n6027) );
  NOR2X0 U7059 ( .IN1(n6030), .IN2(n4251), .QN(n6029) );
  NOR2X0 U7060 ( .IN1(n5691), .IN2(n4328), .QN(n6028) );
  XOR2X1 U7061 ( .IN1(n6031), .IN2(n6032), .Q(n5691) );
  XOR2X1 U7062 ( .IN1(n8844), .IN2(n4042), .Q(n6032) );
  XOR2X1 U7063 ( .IN1(WX8455), .IN2(n3766), .Q(n6031) );
  NOR2X0 U7064 ( .IN1(n6033), .IN2(n6034), .QN(n6026) );
  NOR2X0 U7065 ( .IN1(DFF_1125_n1), .IN2(n4282), .QN(n6034) );
  NOR2X0 U7066 ( .IN1(n5356), .IN2(n5288), .QN(n6033) );
  NAND2X0 U7067 ( .IN1(n4825), .IN2(n8443), .QN(n5288) );
  NAND2X0 U7068 ( .IN1(n6035), .IN2(n6036), .QN(WX7159) );
  NOR2X0 U7069 ( .IN1(n6037), .IN2(n6038), .QN(n6036) );
  NOR2X0 U7070 ( .IN1(n4260), .IN2(n6039), .QN(n6038) );
  NOR2X0 U7071 ( .IN1(n5700), .IN2(n4328), .QN(n6037) );
  XOR2X1 U7072 ( .IN1(n6040), .IN2(n6041), .Q(n5700) );
  XOR2X1 U7073 ( .IN1(n8845), .IN2(n4041), .Q(n6041) );
  XOR2X1 U7074 ( .IN1(WX8453), .IN2(n3768), .Q(n6040) );
  NOR2X0 U7075 ( .IN1(n6042), .IN2(n6043), .QN(n6035) );
  NOR2X0 U7076 ( .IN1(DFF_1126_n1), .IN2(n4282), .QN(n6043) );
  NOR2X0 U7077 ( .IN1(n5356), .IN2(n5289), .QN(n6042) );
  NAND2X0 U7078 ( .IN1(n4826), .IN2(n8444), .QN(n5289) );
  NAND2X0 U7079 ( .IN1(n6044), .IN2(n6045), .QN(WX7157) );
  NOR2X0 U7080 ( .IN1(n6046), .IN2(n6047), .QN(n6045) );
  NOR2X0 U7081 ( .IN1(n6048), .IN2(n4251), .QN(n6047) );
  NOR2X0 U7082 ( .IN1(n5709), .IN2(n4329), .QN(n6046) );
  XOR2X1 U7083 ( .IN1(n6049), .IN2(n6050), .Q(n5709) );
  XOR2X1 U7084 ( .IN1(n8846), .IN2(n4040), .Q(n6050) );
  XOR2X1 U7085 ( .IN1(WX8451), .IN2(n3770), .Q(n6049) );
  NOR2X0 U7086 ( .IN1(n6051), .IN2(n6052), .QN(n6044) );
  NOR2X0 U7087 ( .IN1(DFF_1127_n1), .IN2(n4282), .QN(n6052) );
  NOR2X0 U7088 ( .IN1(n5356), .IN2(n5291), .QN(n6051) );
  NAND2X0 U7089 ( .IN1(n4825), .IN2(n8445), .QN(n5291) );
  NAND2X0 U7090 ( .IN1(n6053), .IN2(n6054), .QN(WX7155) );
  NOR2X0 U7091 ( .IN1(n6055), .IN2(n6056), .QN(n6054) );
  NOR2X0 U7092 ( .IN1(n4260), .IN2(n6057), .QN(n6056) );
  NOR2X0 U7093 ( .IN1(n5718), .IN2(n4328), .QN(n6055) );
  XOR2X1 U7094 ( .IN1(n6058), .IN2(n6059), .Q(n5718) );
  XOR2X1 U7095 ( .IN1(n8847), .IN2(n4039), .Q(n6059) );
  XOR2X1 U7096 ( .IN1(WX8449), .IN2(n3772), .Q(n6058) );
  NOR2X0 U7097 ( .IN1(n6060), .IN2(n6061), .QN(n6053) );
  NOR2X0 U7098 ( .IN1(DFF_1128_n1), .IN2(n4282), .QN(n6061) );
  NOR2X0 U7099 ( .IN1(n5356), .IN2(n5292), .QN(n6060) );
  NAND2X0 U7100 ( .IN1(n4825), .IN2(n8446), .QN(n5292) );
  NAND2X0 U7101 ( .IN1(n6062), .IN2(n6063), .QN(WX7153) );
  NOR2X0 U7102 ( .IN1(n6064), .IN2(n6065), .QN(n6063) );
  NOR2X0 U7103 ( .IN1(n6066), .IN2(n4251), .QN(n6065) );
  NOR2X0 U7104 ( .IN1(n4337), .IN2(n5727), .QN(n6064) );
  XNOR2X1 U7105 ( .IN1(n6067), .IN2(n6068), .Q(n5727) );
  XOR2X1 U7106 ( .IN1(test_so75), .IN2(n8848), .Q(n6068) );
  XOR2X1 U7107 ( .IN1(WX8447), .IN2(n3774), .Q(n6067) );
  NOR2X0 U7108 ( .IN1(n6069), .IN2(n6070), .QN(n6062) );
  NOR2X0 U7109 ( .IN1(DFF_1129_n1), .IN2(n4282), .QN(n6070) );
  NOR2X0 U7110 ( .IN1(n5356), .IN2(n5293), .QN(n6069) );
  NAND2X0 U7111 ( .IN1(n4826), .IN2(n8447), .QN(n5293) );
  NAND2X0 U7112 ( .IN1(n6071), .IN2(n6072), .QN(WX7151) );
  NOR2X0 U7113 ( .IN1(n6073), .IN2(n6074), .QN(n6072) );
  NOR2X0 U7114 ( .IN1(n4260), .IN2(n6075), .QN(n6074) );
  NOR2X0 U7115 ( .IN1(n5736), .IN2(n4328), .QN(n6073) );
  XOR2X1 U7116 ( .IN1(n6076), .IN2(n6077), .Q(n5736) );
  XOR2X1 U7117 ( .IN1(n8849), .IN2(n4038), .Q(n6077) );
  XOR2X1 U7118 ( .IN1(WX8445), .IN2(n3776), .Q(n6076) );
  NOR2X0 U7119 ( .IN1(n6078), .IN2(n6079), .QN(n6071) );
  NOR2X0 U7120 ( .IN1(DFF_1130_n1), .IN2(n4282), .QN(n6079) );
  NOR2X0 U7121 ( .IN1(n4300), .IN2(n5294), .QN(n6078) );
  NAND2X0 U7122 ( .IN1(n4826), .IN2(n8448), .QN(n5294) );
  NAND2X0 U7123 ( .IN1(n6080), .IN2(n6081), .QN(WX7149) );
  NOR2X0 U7124 ( .IN1(n6082), .IN2(n6083), .QN(n6081) );
  NOR2X0 U7125 ( .IN1(n6084), .IN2(n4251), .QN(n6083) );
  NOR2X0 U7126 ( .IN1(n4337), .IN2(n5745), .QN(n6082) );
  XNOR2X1 U7127 ( .IN1(n6085), .IN2(n6086), .Q(n5745) );
  XOR2X1 U7128 ( .IN1(test_so73), .IN2(n8850), .Q(n6086) );
  XOR2X1 U7129 ( .IN1(WX8443), .IN2(n3946), .Q(n6085) );
  NOR2X0 U7130 ( .IN1(n6087), .IN2(n6088), .QN(n6080) );
  NOR2X0 U7131 ( .IN1(DFF_1131_n1), .IN2(n4282), .QN(n6088) );
  NOR2X0 U7132 ( .IN1(n4307), .IN2(n5295), .QN(n6087) );
  NAND2X0 U7133 ( .IN1(n4825), .IN2(n8449), .QN(n5295) );
  NAND2X0 U7134 ( .IN1(n6089), .IN2(n6090), .QN(WX7147) );
  NOR2X0 U7135 ( .IN1(n6091), .IN2(n6092), .QN(n6090) );
  NOR2X0 U7136 ( .IN1(n6093), .IN2(n4251), .QN(n6092) );
  NOR2X0 U7137 ( .IN1(n5754), .IN2(n4330), .QN(n6091) );
  XOR2X1 U7138 ( .IN1(n6094), .IN2(n6095), .Q(n5754) );
  XOR2X1 U7139 ( .IN1(n8851), .IN2(n4037), .Q(n6095) );
  XOR2X1 U7140 ( .IN1(WX8441), .IN2(n3779), .Q(n6094) );
  NOR2X0 U7141 ( .IN1(n6096), .IN2(n6097), .QN(n6089) );
  AND2X1 U7142 ( .IN1(n2152), .IN2(test_so65), .Q(n6097) );
  NOR2X0 U7143 ( .IN1(n4307), .IN2(n5296), .QN(n6096) );
  NAND2X0 U7144 ( .IN1(test_so56), .IN2(n4827), .QN(n5296) );
  NAND2X0 U7145 ( .IN1(n6098), .IN2(n6099), .QN(WX7145) );
  NOR2X0 U7146 ( .IN1(n6100), .IN2(n6101), .QN(n6099) );
  NOR2X0 U7147 ( .IN1(n6102), .IN2(n4251), .QN(n6101) );
  NOR2X0 U7148 ( .IN1(n4337), .IN2(n5763), .QN(n6100) );
  XNOR2X1 U7149 ( .IN1(n6103), .IN2(n6104), .Q(n5763) );
  XOR2X1 U7150 ( .IN1(test_so71), .IN2(n8852), .Q(n6104) );
  XOR2X1 U7151 ( .IN1(WX8439), .IN2(n4036), .Q(n6103) );
  NOR2X0 U7152 ( .IN1(n6105), .IN2(n6106), .QN(n6098) );
  NOR2X0 U7153 ( .IN1(DFF_1133_n1), .IN2(n4282), .QN(n6106) );
  NOR2X0 U7154 ( .IN1(n4307), .IN2(n5297), .QN(n6105) );
  NAND2X0 U7155 ( .IN1(n4826), .IN2(n8452), .QN(n5297) );
  NAND2X0 U7156 ( .IN1(n6107), .IN2(n6108), .QN(WX7143) );
  NOR2X0 U7157 ( .IN1(n6109), .IN2(n6110), .QN(n6108) );
  NOR2X0 U7158 ( .IN1(n6111), .IN2(n4251), .QN(n6110) );
  NOR2X0 U7159 ( .IN1(n5772), .IN2(n4328), .QN(n6109) );
  XOR2X1 U7160 ( .IN1(n6112), .IN2(n6113), .Q(n5772) );
  XOR2X1 U7161 ( .IN1(n8853), .IN2(n4035), .Q(n6113) );
  XOR2X1 U7162 ( .IN1(WX8437), .IN2(n3782), .Q(n6112) );
  NOR2X0 U7163 ( .IN1(n6114), .IN2(n6115), .QN(n6107) );
  NOR2X0 U7164 ( .IN1(DFF_1134_n1), .IN2(n4282), .QN(n6115) );
  NOR2X0 U7165 ( .IN1(n4307), .IN2(n5298), .QN(n6114) );
  NAND2X0 U7166 ( .IN1(n4826), .IN2(n8453), .QN(n5298) );
  NAND2X0 U7167 ( .IN1(n6116), .IN2(n6117), .QN(WX7141) );
  NOR2X0 U7168 ( .IN1(n6118), .IN2(n6119), .QN(n6117) );
  NOR2X0 U7169 ( .IN1(n6120), .IN2(n4251), .QN(n6119) );
  NOR2X0 U7170 ( .IN1(n4337), .IN2(n5781), .QN(n6118) );
  XNOR2X1 U7171 ( .IN1(n6121), .IN2(n6122), .Q(n5781) );
  XOR2X1 U7172 ( .IN1(test_so69), .IN2(n8854), .Q(n6122) );
  XOR2X1 U7173 ( .IN1(WX8563), .IN2(n4034), .Q(n6121) );
  NOR2X0 U7174 ( .IN1(n6123), .IN2(n6124), .QN(n6116) );
  NOR2X0 U7175 ( .IN1(DFF_1135_n1), .IN2(n4282), .QN(n6124) );
  NOR2X0 U7176 ( .IN1(n4307), .IN2(n5299), .QN(n6123) );
  NAND2X0 U7177 ( .IN1(n4826), .IN2(n8454), .QN(n5299) );
  NAND2X0 U7178 ( .IN1(n6125), .IN2(n6126), .QN(WX7139) );
  NOR2X0 U7179 ( .IN1(n6127), .IN2(n6128), .QN(n6126) );
  NOR2X0 U7180 ( .IN1(n6129), .IN2(n4252), .QN(n6128) );
  NOR2X0 U7181 ( .IN1(n5790), .IN2(n4330), .QN(n6127) );
  XOR2X1 U7182 ( .IN1(n6130), .IN2(n6131), .Q(n5790) );
  XOR2X1 U7183 ( .IN1(n3616), .IN2(n4772), .Q(n6131) );
  XOR2X1 U7184 ( .IN1(n6132), .IN2(n3945), .Q(n6130) );
  XOR2X1 U7185 ( .IN1(WX8561), .IN2(n8855), .Q(n6132) );
  NOR2X0 U7186 ( .IN1(n6133), .IN2(n6134), .QN(n6125) );
  NOR2X0 U7187 ( .IN1(DFF_1136_n1), .IN2(n4282), .QN(n6134) );
  NOR2X0 U7188 ( .IN1(n4307), .IN2(n5300), .QN(n6133) );
  NAND2X0 U7189 ( .IN1(n4824), .IN2(n8455), .QN(n5300) );
  NAND2X0 U7190 ( .IN1(n6135), .IN2(n6136), .QN(WX7137) );
  NOR2X0 U7191 ( .IN1(n6137), .IN2(n6138), .QN(n6136) );
  NOR2X0 U7192 ( .IN1(n6139), .IN2(n4251), .QN(n6138) );
  NOR2X0 U7193 ( .IN1(n5800), .IN2(n4329), .QN(n6137) );
  XOR2X1 U7194 ( .IN1(n6140), .IN2(n6141), .Q(n5800) );
  XOR2X1 U7195 ( .IN1(n3617), .IN2(n4772), .Q(n6141) );
  XOR2X1 U7196 ( .IN1(n6142), .IN2(n4033), .Q(n6140) );
  XOR2X1 U7197 ( .IN1(WX8559), .IN2(n8856), .Q(n6142) );
  NOR2X0 U7198 ( .IN1(n6143), .IN2(n6144), .QN(n6135) );
  NOR2X0 U7199 ( .IN1(DFF_1137_n1), .IN2(n4281), .QN(n6144) );
  NOR2X0 U7200 ( .IN1(n4307), .IN2(n5302), .QN(n6143) );
  NAND2X0 U7201 ( .IN1(n4825), .IN2(n8456), .QN(n5302) );
  NAND2X0 U7202 ( .IN1(n6145), .IN2(n6146), .QN(WX7135) );
  NOR2X0 U7203 ( .IN1(n6147), .IN2(n6148), .QN(n6146) );
  NOR2X0 U7204 ( .IN1(n6149), .IN2(n4251), .QN(n6148) );
  NOR2X0 U7205 ( .IN1(n5810), .IN2(n4329), .QN(n6147) );
  XOR2X1 U7206 ( .IN1(n6150), .IN2(n6151), .Q(n5810) );
  XOR2X1 U7207 ( .IN1(n3618), .IN2(n4772), .Q(n6151) );
  XOR2X1 U7208 ( .IN1(n6152), .IN2(n4032), .Q(n6150) );
  XOR2X1 U7209 ( .IN1(WX8557), .IN2(n8857), .Q(n6152) );
  NOR2X0 U7210 ( .IN1(n6153), .IN2(n6154), .QN(n6145) );
  NOR2X0 U7211 ( .IN1(DFF_1138_n1), .IN2(n4281), .QN(n6154) );
  NOR2X0 U7212 ( .IN1(n4307), .IN2(n5303), .QN(n6153) );
  NAND2X0 U7213 ( .IN1(n4825), .IN2(n8457), .QN(n5303) );
  NAND2X0 U7214 ( .IN1(n6155), .IN2(n6156), .QN(WX7133) );
  NOR2X0 U7215 ( .IN1(n6157), .IN2(n6158), .QN(n6156) );
  NOR2X0 U7216 ( .IN1(n6159), .IN2(n4251), .QN(n6158) );
  NOR2X0 U7217 ( .IN1(n5820), .IN2(n4329), .QN(n6157) );
  XOR2X1 U7218 ( .IN1(n6160), .IN2(n6161), .Q(n5820) );
  XOR2X1 U7219 ( .IN1(n3619), .IN2(n4772), .Q(n6161) );
  XOR2X1 U7220 ( .IN1(n6162), .IN2(n4031), .Q(n6160) );
  XOR2X1 U7221 ( .IN1(WX8555), .IN2(n8858), .Q(n6162) );
  NOR2X0 U7222 ( .IN1(n6163), .IN2(n6164), .QN(n6155) );
  NOR2X0 U7223 ( .IN1(DFF_1139_n1), .IN2(n4281), .QN(n6164) );
  NOR2X0 U7224 ( .IN1(n4307), .IN2(n5304), .QN(n6163) );
  NAND2X0 U7225 ( .IN1(n4824), .IN2(n8458), .QN(n5304) );
  NAND2X0 U7226 ( .IN1(n6165), .IN2(n6166), .QN(WX7131) );
  NOR2X0 U7227 ( .IN1(n6167), .IN2(n6168), .QN(n6166) );
  NOR2X0 U7228 ( .IN1(n6169), .IN2(n4252), .QN(n6168) );
  NOR2X0 U7229 ( .IN1(n5830), .IN2(n4329), .QN(n6167) );
  XOR2X1 U7230 ( .IN1(n6170), .IN2(n6171), .Q(n5830) );
  XOR2X1 U7231 ( .IN1(n3620), .IN2(n4772), .Q(n6171) );
  XOR2X1 U7232 ( .IN1(n6172), .IN2(n4030), .Q(n6170) );
  XOR2X1 U7233 ( .IN1(WX8553), .IN2(n8859), .Q(n6172) );
  NOR2X0 U7234 ( .IN1(n6173), .IN2(n6174), .QN(n6165) );
  NOR2X0 U7235 ( .IN1(DFF_1140_n1), .IN2(n4281), .QN(n6174) );
  NOR2X0 U7236 ( .IN1(n4307), .IN2(n5305), .QN(n6173) );
  NAND2X0 U7237 ( .IN1(n4825), .IN2(n8459), .QN(n5305) );
  NAND2X0 U7238 ( .IN1(n6175), .IN2(n6176), .QN(WX7129) );
  NOR2X0 U7239 ( .IN1(n6177), .IN2(n6178), .QN(n6176) );
  NOR2X0 U7240 ( .IN1(n4260), .IN2(n6179), .QN(n6178) );
  NOR2X0 U7241 ( .IN1(n5840), .IN2(n4329), .QN(n6177) );
  XOR2X1 U7242 ( .IN1(n6180), .IN2(n6181), .Q(n5840) );
  XOR2X1 U7243 ( .IN1(n3621), .IN2(n4772), .Q(n6181) );
  XOR2X1 U7244 ( .IN1(n6182), .IN2(n4029), .Q(n6180) );
  XOR2X1 U7245 ( .IN1(WX8551), .IN2(n8860), .Q(n6182) );
  NOR2X0 U7246 ( .IN1(n6183), .IN2(n6184), .QN(n6175) );
  NOR2X0 U7247 ( .IN1(DFF_1141_n1), .IN2(n4281), .QN(n6184) );
  NOR2X0 U7248 ( .IN1(n4307), .IN2(n5306), .QN(n6183) );
  NAND2X0 U7249 ( .IN1(n4824), .IN2(n8460), .QN(n5306) );
  NAND2X0 U7250 ( .IN1(n6185), .IN2(n6186), .QN(WX7127) );
  NOR2X0 U7251 ( .IN1(n6187), .IN2(n6188), .QN(n6186) );
  NOR2X0 U7252 ( .IN1(n6189), .IN2(n4251), .QN(n6188) );
  NOR2X0 U7253 ( .IN1(n5850), .IN2(n4329), .QN(n6187) );
  XOR2X1 U7254 ( .IN1(n6190), .IN2(n6191), .Q(n5850) );
  XOR2X1 U7255 ( .IN1(n3622), .IN2(n4772), .Q(n6191) );
  XOR2X1 U7256 ( .IN1(n6192), .IN2(n4028), .Q(n6190) );
  XOR2X1 U7257 ( .IN1(WX8549), .IN2(n8861), .Q(n6192) );
  NOR2X0 U7258 ( .IN1(n6193), .IN2(n6194), .QN(n6185) );
  NOR2X0 U7259 ( .IN1(DFF_1142_n1), .IN2(n4281), .QN(n6194) );
  NOR2X0 U7260 ( .IN1(n4307), .IN2(n5307), .QN(n6193) );
  NAND2X0 U7261 ( .IN1(n4825), .IN2(n8461), .QN(n5307) );
  NAND2X0 U7262 ( .IN1(n6195), .IN2(n6196), .QN(WX7125) );
  NOR2X0 U7263 ( .IN1(n6197), .IN2(n6198), .QN(n6196) );
  NOR2X0 U7264 ( .IN1(n4260), .IN2(n6199), .QN(n6198) );
  NOR2X0 U7265 ( .IN1(n5860), .IN2(n4329), .QN(n6197) );
  XOR2X1 U7266 ( .IN1(n6200), .IN2(n6201), .Q(n5860) );
  XOR2X1 U7267 ( .IN1(n3623), .IN2(n4773), .Q(n6201) );
  XOR2X1 U7268 ( .IN1(n6202), .IN2(n4027), .Q(n6200) );
  XOR2X1 U7269 ( .IN1(WX8547), .IN2(n8862), .Q(n6202) );
  NOR2X0 U7270 ( .IN1(n6203), .IN2(n6204), .QN(n6195) );
  NOR2X0 U7271 ( .IN1(DFF_1143_n1), .IN2(n4281), .QN(n6204) );
  NOR2X0 U7272 ( .IN1(n4306), .IN2(n5308), .QN(n6203) );
  NAND2X0 U7273 ( .IN1(n4825), .IN2(n8462), .QN(n5308) );
  NAND2X0 U7274 ( .IN1(n6205), .IN2(n6206), .QN(WX7123) );
  NOR2X0 U7275 ( .IN1(n6207), .IN2(n6208), .QN(n6206) );
  NOR2X0 U7276 ( .IN1(n6209), .IN2(n4251), .QN(n6208) );
  NOR2X0 U7277 ( .IN1(n5870), .IN2(n4329), .QN(n6207) );
  XOR2X1 U7278 ( .IN1(n6210), .IN2(n6211), .Q(n5870) );
  XOR2X1 U7279 ( .IN1(n3624), .IN2(n4773), .Q(n6211) );
  XOR2X1 U7280 ( .IN1(n6212), .IN2(n4026), .Q(n6210) );
  XOR2X1 U7281 ( .IN1(WX8545), .IN2(n8863), .Q(n6212) );
  NOR2X0 U7282 ( .IN1(n6213), .IN2(n6214), .QN(n6205) );
  NOR2X0 U7283 ( .IN1(DFF_1144_n1), .IN2(n4281), .QN(n6214) );
  NOR2X0 U7284 ( .IN1(n4306), .IN2(n5309), .QN(n6213) );
  NAND2X0 U7285 ( .IN1(n4824), .IN2(n8463), .QN(n5309) );
  NAND2X0 U7286 ( .IN1(n6215), .IN2(n6216), .QN(WX7121) );
  NOR2X0 U7287 ( .IN1(n6217), .IN2(n6218), .QN(n6216) );
  NOR2X0 U7288 ( .IN1(n4260), .IN2(n6219), .QN(n6218) );
  NOR2X0 U7289 ( .IN1(n5880), .IN2(n4329), .QN(n6217) );
  XOR2X1 U7290 ( .IN1(n6220), .IN2(n6221), .Q(n5880) );
  XOR2X1 U7291 ( .IN1(n3625), .IN2(n4773), .Q(n6221) );
  XOR2X1 U7292 ( .IN1(n6222), .IN2(n4025), .Q(n6220) );
  XOR2X1 U7293 ( .IN1(WX8543), .IN2(n8864), .Q(n6222) );
  NOR2X0 U7294 ( .IN1(n6223), .IN2(n6224), .QN(n6215) );
  NOR2X0 U7295 ( .IN1(DFF_1145_n1), .IN2(n4281), .QN(n6224) );
  NOR2X0 U7296 ( .IN1(n4306), .IN2(n5310), .QN(n6223) );
  NAND2X0 U7297 ( .IN1(n4824), .IN2(n8464), .QN(n5310) );
  NAND2X0 U7298 ( .IN1(n6225), .IN2(n6226), .QN(WX7119) );
  NOR2X0 U7299 ( .IN1(n6227), .IN2(n6228), .QN(n6226) );
  NOR2X0 U7300 ( .IN1(n6229), .IN2(n4252), .QN(n6228) );
  NOR2X0 U7301 ( .IN1(n4338), .IN2(n5890), .QN(n6227) );
  XNOR2X1 U7302 ( .IN1(n6230), .IN2(n6231), .Q(n5890) );
  XOR2X1 U7303 ( .IN1(n3626), .IN2(n4773), .Q(n6231) );
  XOR2X1 U7304 ( .IN1(WX8477), .IN2(n6232), .Q(n6230) );
  XOR2X1 U7305 ( .IN1(test_so74), .IN2(n8865), .Q(n6232) );
  NOR2X0 U7306 ( .IN1(n6233), .IN2(n6234), .QN(n6225) );
  NOR2X0 U7307 ( .IN1(DFF_1146_n1), .IN2(n4281), .QN(n6234) );
  NOR2X0 U7308 ( .IN1(n4306), .IN2(n5311), .QN(n6233) );
  NAND2X0 U7309 ( .IN1(n4823), .IN2(n8465), .QN(n5311) );
  NAND2X0 U7310 ( .IN1(n6235), .IN2(n6236), .QN(WX7117) );
  NOR2X0 U7311 ( .IN1(n6237), .IN2(n6238), .QN(n6236) );
  NOR2X0 U7312 ( .IN1(n5352), .IN2(n6239), .QN(n6238) );
  NOR2X0 U7313 ( .IN1(n5900), .IN2(n4330), .QN(n6237) );
  XOR2X1 U7314 ( .IN1(n6240), .IN2(n6241), .Q(n5900) );
  XOR2X1 U7315 ( .IN1(n3627), .IN2(n4773), .Q(n6241) );
  XOR2X1 U7316 ( .IN1(n6242), .IN2(n4024), .Q(n6240) );
  XOR2X1 U7317 ( .IN1(WX8539), .IN2(n8866), .Q(n6242) );
  NOR2X0 U7318 ( .IN1(n6243), .IN2(n6244), .QN(n6235) );
  NOR2X0 U7319 ( .IN1(DFF_1147_n1), .IN2(n4281), .QN(n6244) );
  NOR2X0 U7320 ( .IN1(n4306), .IN2(n5313), .QN(n6243) );
  NAND2X0 U7321 ( .IN1(n4823), .IN2(n8466), .QN(n5313) );
  NAND2X0 U7322 ( .IN1(n6245), .IN2(n6246), .QN(WX7115) );
  NOR2X0 U7323 ( .IN1(n6247), .IN2(n6248), .QN(n6246) );
  NOR2X0 U7324 ( .IN1(n6249), .IN2(n4252), .QN(n6248) );
  NOR2X0 U7325 ( .IN1(n4337), .IN2(n5910), .QN(n6247) );
  XNOR2X1 U7326 ( .IN1(n6250), .IN2(n6251), .Q(n5910) );
  XOR2X1 U7327 ( .IN1(n4023), .IN2(n4773), .Q(n6251) );
  XOR2X1 U7328 ( .IN1(n6252), .IN2(n8869), .Q(n6250) );
  XOR2X1 U7329 ( .IN1(n8868), .IN2(n8867), .Q(n6252) );
  NOR2X0 U7330 ( .IN1(n6253), .IN2(n6254), .QN(n6245) );
  NOR2X0 U7331 ( .IN1(DFF_1148_n1), .IN2(n4281), .QN(n6254) );
  NOR2X0 U7332 ( .IN1(n4306), .IN2(n5314), .QN(n6253) );
  NAND2X0 U7333 ( .IN1(n4824), .IN2(n8467), .QN(n5314) );
  NAND2X0 U7334 ( .IN1(n6255), .IN2(n6256), .QN(WX7113) );
  NOR2X0 U7335 ( .IN1(n6257), .IN2(n6258), .QN(n6256) );
  NOR2X0 U7336 ( .IN1(n6259), .IN2(n4252), .QN(n6258) );
  NOR2X0 U7337 ( .IN1(n5920), .IN2(n4329), .QN(n6257) );
  XOR2X1 U7338 ( .IN1(n6260), .IN2(n6261), .Q(n5920) );
  XOR2X1 U7339 ( .IN1(n3628), .IN2(n4773), .Q(n6261) );
  XOR2X1 U7340 ( .IN1(n6262), .IN2(n4022), .Q(n6260) );
  XOR2X1 U7341 ( .IN1(WX8535), .IN2(n8870), .Q(n6262) );
  NOR2X0 U7342 ( .IN1(n6263), .IN2(n6264), .QN(n6255) );
  AND2X1 U7343 ( .IN1(n2152), .IN2(test_so66), .Q(n6264) );
  NOR2X0 U7344 ( .IN1(n4306), .IN2(n5315), .QN(n6263) );
  NAND2X0 U7345 ( .IN1(test_so55), .IN2(n4828), .QN(n5315) );
  NAND2X0 U7346 ( .IN1(n6265), .IN2(n6266), .QN(WX7111) );
  NOR2X0 U7347 ( .IN1(n6267), .IN2(n6268), .QN(n6266) );
  NOR2X0 U7348 ( .IN1(n6269), .IN2(n4252), .QN(n6268) );
  NOR2X0 U7349 ( .IN1(n4338), .IN2(n5930), .QN(n6267) );
  XNOR2X1 U7350 ( .IN1(n6270), .IN2(n6271), .Q(n5930) );
  XOR2X1 U7351 ( .IN1(n4021), .IN2(n4773), .Q(n6271) );
  XOR2X1 U7352 ( .IN1(n6272), .IN2(n8873), .Q(n6270) );
  XOR2X1 U7353 ( .IN1(n8872), .IN2(n8871), .Q(n6272) );
  NOR2X0 U7354 ( .IN1(n6273), .IN2(n6274), .QN(n6265) );
  NOR2X0 U7355 ( .IN1(DFF_1150_n1), .IN2(n4281), .QN(n6274) );
  NOR2X0 U7356 ( .IN1(n4306), .IN2(n5316), .QN(n6273) );
  NAND2X0 U7357 ( .IN1(n4824), .IN2(n8470), .QN(n5316) );
  NAND2X0 U7358 ( .IN1(n6275), .IN2(n6276), .QN(WX7109) );
  NOR2X0 U7359 ( .IN1(n6277), .IN2(n6278), .QN(n6276) );
  NOR2X0 U7360 ( .IN1(n6279), .IN2(n4252), .QN(n6278) );
  NOR2X0 U7361 ( .IN1(n5940), .IN2(n4329), .QN(n6277) );
  XOR2X1 U7362 ( .IN1(n6280), .IN2(n6281), .Q(n5940) );
  XOR2X1 U7363 ( .IN1(n3584), .IN2(n4773), .Q(n6281) );
  XOR2X1 U7364 ( .IN1(n6282), .IN2(n4020), .Q(n6280) );
  XOR2X1 U7365 ( .IN1(WX8531), .IN2(n8874), .Q(n6282) );
  NOR2X0 U7366 ( .IN1(n6283), .IN2(n6284), .QN(n6275) );
  NOR2X0 U7367 ( .IN1(n3934), .IN2(n5606), .QN(n6284) );
  NOR2X0 U7368 ( .IN1(DFF_1151_n1), .IN2(n4281), .QN(n6283) );
  OR2X1 U7369 ( .IN1(n6285), .IN2(n6286), .Q(WX706) );
  NAND2X0 U7370 ( .IN1(n6287), .IN2(n6288), .QN(n6286) );
  NAND2X0 U7371 ( .IN1(n4266), .IN2(n6289), .QN(n6288) );
  OR2X1 U7372 ( .IN1(n4280), .IN2(DFF_160_n1), .Q(n6287) );
  NAND2X0 U7373 ( .IN1(n6290), .IN2(n6291), .QN(n6285) );
  OR2X1 U7374 ( .IN1(n6292), .IN2(n4326), .Q(n6291) );
  NAND2X0 U7375 ( .IN1(WX544), .IN2(n4315), .QN(n6290) );
  OR2X1 U7376 ( .IN1(n6293), .IN2(n6294), .Q(WX704) );
  NAND2X0 U7377 ( .IN1(n6295), .IN2(n6296), .QN(n6294) );
  NAND2X0 U7378 ( .IN1(n4270), .IN2(n6297), .QN(n6296) );
  NAND2X0 U7379 ( .IN1(test_so9), .IN2(n2152), .QN(n6295) );
  NAND2X0 U7380 ( .IN1(n6298), .IN2(n6299), .QN(n6293) );
  NAND2X0 U7381 ( .IN1(n2153), .IN2(n6300), .QN(n6299) );
  NAND2X0 U7382 ( .IN1(WX542), .IN2(n4321), .QN(n6298) );
  OR2X1 U7383 ( .IN1(n6301), .IN2(n6302), .Q(WX702) );
  NAND2X0 U7384 ( .IN1(n6303), .IN2(n6304), .QN(n6302) );
  OR2X1 U7385 ( .IN1(n6305), .IN2(n4246), .Q(n6304) );
  OR2X1 U7386 ( .IN1(n4280), .IN2(DFF_162_n1), .Q(n6303) );
  NAND2X0 U7387 ( .IN1(n6306), .IN2(n6307), .QN(n6301) );
  NAND2X0 U7388 ( .IN1(n2153), .IN2(n6308), .QN(n6307) );
  NAND2X0 U7389 ( .IN1(WX540), .IN2(n4321), .QN(n6306) );
  AND2X1 U7390 ( .IN1(n4800), .IN2(n3934), .Q(WX7011) );
  OR2X1 U7391 ( .IN1(n6309), .IN2(n6310), .Q(WX700) );
  NAND2X0 U7392 ( .IN1(n6311), .IN2(n6312), .QN(n6310) );
  NAND2X0 U7393 ( .IN1(n4270), .IN2(n6313), .QN(n6312) );
  OR2X1 U7394 ( .IN1(n4280), .IN2(DFF_163_n1), .Q(n6311) );
  NAND2X0 U7395 ( .IN1(n6314), .IN2(n6315), .QN(n6309) );
  NAND2X0 U7396 ( .IN1(n2153), .IN2(n6316), .QN(n6315) );
  NAND2X0 U7397 ( .IN1(WX538), .IN2(n4321), .QN(n6314) );
  OR2X1 U7398 ( .IN1(n6317), .IN2(n6318), .Q(WX698) );
  NAND2X0 U7399 ( .IN1(n6319), .IN2(n6320), .QN(n6318) );
  NAND2X0 U7400 ( .IN1(n4270), .IN2(n6321), .QN(n6320) );
  OR2X1 U7401 ( .IN1(n4280), .IN2(DFF_164_n1), .Q(n6319) );
  NAND2X0 U7402 ( .IN1(n6322), .IN2(n6323), .QN(n6317) );
  OR2X1 U7403 ( .IN1(n6324), .IN2(n4326), .Q(n6323) );
  NAND2X0 U7404 ( .IN1(WX536), .IN2(n4321), .QN(n6322) );
  OR2X1 U7405 ( .IN1(n6325), .IN2(n6326), .Q(WX696) );
  NAND2X0 U7406 ( .IN1(n6327), .IN2(n6328), .QN(n6326) );
  NAND2X0 U7407 ( .IN1(n4270), .IN2(n6329), .QN(n6328) );
  OR2X1 U7408 ( .IN1(n4280), .IN2(DFF_165_n1), .Q(n6327) );
  NAND2X0 U7409 ( .IN1(n6330), .IN2(n6331), .QN(n6325) );
  NAND2X0 U7410 ( .IN1(n2153), .IN2(n6332), .QN(n6331) );
  NAND2X0 U7411 ( .IN1(WX534), .IN2(n4321), .QN(n6330) );
  OR2X1 U7412 ( .IN1(n6333), .IN2(n6334), .Q(WX694) );
  NAND2X0 U7413 ( .IN1(n6335), .IN2(n6336), .QN(n6334) );
  OR2X1 U7414 ( .IN1(n6337), .IN2(n4246), .Q(n6336) );
  OR2X1 U7415 ( .IN1(n4280), .IN2(DFF_166_n1), .Q(n6335) );
  NAND2X0 U7416 ( .IN1(n6338), .IN2(n6339), .QN(n6333) );
  NAND2X0 U7417 ( .IN1(n2153), .IN2(n6340), .QN(n6339) );
  NAND2X0 U7418 ( .IN1(WX532), .IN2(n4321), .QN(n6338) );
  OR2X1 U7419 ( .IN1(n6341), .IN2(n6342), .Q(WX692) );
  NAND2X0 U7420 ( .IN1(n6343), .IN2(n6344), .QN(n6342) );
  NAND2X0 U7421 ( .IN1(n4270), .IN2(n6345), .QN(n6344) );
  OR2X1 U7422 ( .IN1(n4280), .IN2(DFF_167_n1), .Q(n6343) );
  NAND2X0 U7423 ( .IN1(n6346), .IN2(n6347), .QN(n6341) );
  NAND2X0 U7424 ( .IN1(n2153), .IN2(n6348), .QN(n6347) );
  NAND2X0 U7425 ( .IN1(WX530), .IN2(n4321), .QN(n6346) );
  OR2X1 U7426 ( .IN1(n6349), .IN2(n6350), .Q(WX690) );
  NAND2X0 U7427 ( .IN1(n6351), .IN2(n6352), .QN(n6350) );
  NAND2X0 U7428 ( .IN1(n4270), .IN2(n6353), .QN(n6352) );
  OR2X1 U7429 ( .IN1(n4280), .IN2(DFF_168_n1), .Q(n6351) );
  NAND2X0 U7430 ( .IN1(n6354), .IN2(n6355), .QN(n6349) );
  NAND2X0 U7431 ( .IN1(n2153), .IN2(n6356), .QN(n6355) );
  NAND2X0 U7432 ( .IN1(WX528), .IN2(n4320), .QN(n6354) );
  OR2X1 U7433 ( .IN1(n6357), .IN2(n6358), .Q(WX688) );
  NAND2X0 U7434 ( .IN1(n6359), .IN2(n6360), .QN(n6358) );
  NAND2X0 U7435 ( .IN1(n4270), .IN2(n6361), .QN(n6360) );
  OR2X1 U7436 ( .IN1(n4280), .IN2(DFF_169_n1), .Q(n6359) );
  NAND2X0 U7437 ( .IN1(n6362), .IN2(n6363), .QN(n6357) );
  NAND2X0 U7438 ( .IN1(n2153), .IN2(n6364), .QN(n6363) );
  NAND2X0 U7439 ( .IN1(WX526), .IN2(n4320), .QN(n6362) );
  OR2X1 U7440 ( .IN1(n6365), .IN2(n6366), .Q(WX686) );
  NAND2X0 U7441 ( .IN1(n6367), .IN2(n6368), .QN(n6366) );
  OR2X1 U7442 ( .IN1(n6369), .IN2(n4246), .Q(n6368) );
  OR2X1 U7443 ( .IN1(n4280), .IN2(DFF_170_n1), .Q(n6367) );
  NAND2X0 U7444 ( .IN1(n6370), .IN2(n6371), .QN(n6365) );
  OR2X1 U7445 ( .IN1(n6372), .IN2(n4326), .Q(n6371) );
  NAND2X0 U7446 ( .IN1(WX524), .IN2(n4320), .QN(n6370) );
  OR2X1 U7447 ( .IN1(n6373), .IN2(n6374), .Q(WX684) );
  NAND2X0 U7448 ( .IN1(n6375), .IN2(n6376), .QN(n6374) );
  NAND2X0 U7449 ( .IN1(n4270), .IN2(n6377), .QN(n6376) );
  OR2X1 U7450 ( .IN1(n4280), .IN2(DFF_171_n1), .Q(n6375) );
  NAND2X0 U7451 ( .IN1(n6378), .IN2(n6379), .QN(n6373) );
  NAND2X0 U7452 ( .IN1(n2153), .IN2(n6380), .QN(n6379) );
  NAND2X0 U7453 ( .IN1(WX522), .IN2(n4320), .QN(n6378) );
  OR2X1 U7454 ( .IN1(n6381), .IN2(n6382), .Q(WX682) );
  NAND2X0 U7455 ( .IN1(n6383), .IN2(n6384), .QN(n6382) );
  NAND2X0 U7456 ( .IN1(n4269), .IN2(n6385), .QN(n6384) );
  OR2X1 U7457 ( .IN1(n4279), .IN2(DFF_172_n1), .Q(n6383) );
  NAND2X0 U7458 ( .IN1(n6386), .IN2(n6387), .QN(n6381) );
  NAND2X0 U7459 ( .IN1(n2153), .IN2(n6388), .QN(n6387) );
  NAND2X0 U7460 ( .IN1(WX520), .IN2(n4320), .QN(n6386) );
  OR2X1 U7461 ( .IN1(n6389), .IN2(n6390), .Q(WX680) );
  NAND2X0 U7462 ( .IN1(n6391), .IN2(n6392), .QN(n6390) );
  NAND2X0 U7463 ( .IN1(n4269), .IN2(n6393), .QN(n6392) );
  OR2X1 U7464 ( .IN1(n4279), .IN2(DFF_173_n1), .Q(n6391) );
  NAND2X0 U7465 ( .IN1(n6394), .IN2(n6395), .QN(n6389) );
  NAND2X0 U7466 ( .IN1(n2153), .IN2(n6396), .QN(n6395) );
  NAND2X0 U7467 ( .IN1(WX518), .IN2(n4320), .QN(n6394) );
  OR2X1 U7468 ( .IN1(n6397), .IN2(n6398), .Q(WX678) );
  NAND2X0 U7469 ( .IN1(n6399), .IN2(n6400), .QN(n6398) );
  NAND2X0 U7470 ( .IN1(n4269), .IN2(n6401), .QN(n6400) );
  OR2X1 U7471 ( .IN1(n4279), .IN2(DFF_174_n1), .Q(n6399) );
  NAND2X0 U7472 ( .IN1(n6402), .IN2(n6403), .QN(n6397) );
  OR2X1 U7473 ( .IN1(n6404), .IN2(n4326), .Q(n6403) );
  NAND2X0 U7474 ( .IN1(WX516), .IN2(n4320), .QN(n6402) );
  OR2X1 U7475 ( .IN1(n6405), .IN2(n6406), .Q(WX676) );
  NAND2X0 U7476 ( .IN1(n6407), .IN2(n6408), .QN(n6406) );
  NAND2X0 U7477 ( .IN1(n4269), .IN2(n6409), .QN(n6408) );
  OR2X1 U7478 ( .IN1(n4279), .IN2(DFF_175_n1), .Q(n6407) );
  NAND2X0 U7479 ( .IN1(n6410), .IN2(n6411), .QN(n6405) );
  NAND2X0 U7480 ( .IN1(n2153), .IN2(n6412), .QN(n6411) );
  NAND2X0 U7481 ( .IN1(WX514), .IN2(n4320), .QN(n6410) );
  OR2X1 U7482 ( .IN1(n6413), .IN2(n6414), .Q(WX674) );
  NAND2X0 U7483 ( .IN1(n6415), .IN2(n6416), .QN(n6414) );
  OR2X1 U7484 ( .IN1(n6417), .IN2(n4247), .Q(n6416) );
  OR2X1 U7485 ( .IN1(n4279), .IN2(DFF_176_n1), .Q(n6415) );
  NAND2X0 U7486 ( .IN1(n6418), .IN2(n6419), .QN(n6413) );
  NAND2X0 U7487 ( .IN1(n2153), .IN2(n6420), .QN(n6419) );
  NAND2X0 U7488 ( .IN1(WX512), .IN2(n4320), .QN(n6418) );
  OR2X1 U7489 ( .IN1(n6421), .IN2(n6422), .Q(WX672) );
  NAND2X0 U7490 ( .IN1(n6423), .IN2(n6424), .QN(n6422) );
  NAND2X0 U7491 ( .IN1(n4269), .IN2(n6425), .QN(n6424) );
  OR2X1 U7492 ( .IN1(n4279), .IN2(DFF_177_n1), .Q(n6423) );
  NAND2X0 U7493 ( .IN1(n6426), .IN2(n6427), .QN(n6421) );
  NAND2X0 U7494 ( .IN1(n2153), .IN2(n6428), .QN(n6427) );
  NAND2X0 U7495 ( .IN1(WX510), .IN2(n4320), .QN(n6426) );
  OR2X1 U7496 ( .IN1(n6429), .IN2(n6430), .Q(WX670) );
  NAND2X0 U7497 ( .IN1(n6431), .IN2(n6432), .QN(n6430) );
  NAND2X0 U7498 ( .IN1(n4269), .IN2(n6433), .QN(n6432) );
  OR2X1 U7499 ( .IN1(n4279), .IN2(DFF_178_n1), .Q(n6431) );
  NAND2X0 U7500 ( .IN1(n6434), .IN2(n6435), .QN(n6429) );
  OR2X1 U7501 ( .IN1(n6436), .IN2(n4326), .Q(n6435) );
  NAND2X0 U7502 ( .IN1(WX508), .IN2(n4319), .QN(n6434) );
  OR2X1 U7503 ( .IN1(n6437), .IN2(n6438), .Q(WX668) );
  NAND2X0 U7504 ( .IN1(n6439), .IN2(n6440), .QN(n6438) );
  NAND2X0 U7505 ( .IN1(n4269), .IN2(n6441), .QN(n6440) );
  NAND2X0 U7506 ( .IN1(test_so10), .IN2(n2152), .QN(n6439) );
  NAND2X0 U7507 ( .IN1(n6442), .IN2(n6443), .QN(n6437) );
  NAND2X0 U7508 ( .IN1(n2153), .IN2(n6444), .QN(n6443) );
  NAND2X0 U7509 ( .IN1(WX506), .IN2(n4319), .QN(n6442) );
  OR2X1 U7510 ( .IN1(n6445), .IN2(n6446), .Q(WX666) );
  NAND2X0 U7511 ( .IN1(n6447), .IN2(n6448), .QN(n6446) );
  OR2X1 U7512 ( .IN1(n6449), .IN2(n4246), .Q(n6448) );
  OR2X1 U7513 ( .IN1(n4279), .IN2(DFF_180_n1), .Q(n6447) );
  NAND2X0 U7514 ( .IN1(n6450), .IN2(n6451), .QN(n6445) );
  NAND2X0 U7515 ( .IN1(n2153), .IN2(n6452), .QN(n6451) );
  NAND2X0 U7516 ( .IN1(WX504), .IN2(n4319), .QN(n6450) );
  OR2X1 U7517 ( .IN1(n6453), .IN2(n6454), .Q(WX664) );
  NAND2X0 U7518 ( .IN1(n6455), .IN2(n6456), .QN(n6454) );
  NAND2X0 U7519 ( .IN1(n4269), .IN2(n6457), .QN(n6456) );
  OR2X1 U7520 ( .IN1(n4279), .IN2(DFF_181_n1), .Q(n6455) );
  NAND2X0 U7521 ( .IN1(n6458), .IN2(n6459), .QN(n6453) );
  NAND2X0 U7522 ( .IN1(n2153), .IN2(n6460), .QN(n6459) );
  NAND2X0 U7523 ( .IN1(WX502), .IN2(n4319), .QN(n6458) );
  OR2X1 U7524 ( .IN1(n6461), .IN2(n6462), .Q(WX662) );
  NAND2X0 U7525 ( .IN1(n6463), .IN2(n6464), .QN(n6462) );
  NAND2X0 U7526 ( .IN1(n4269), .IN2(n6465), .QN(n6464) );
  OR2X1 U7527 ( .IN1(n4279), .IN2(DFF_182_n1), .Q(n6463) );
  NAND2X0 U7528 ( .IN1(n6466), .IN2(n6467), .QN(n6461) );
  OR2X1 U7529 ( .IN1(n6468), .IN2(n4326), .Q(n6467) );
  NAND2X0 U7530 ( .IN1(WX500), .IN2(n4319), .QN(n6466) );
  OR2X1 U7531 ( .IN1(n6469), .IN2(n6470), .Q(WX660) );
  NAND2X0 U7532 ( .IN1(n6471), .IN2(n6472), .QN(n6470) );
  NAND2X0 U7533 ( .IN1(n4268), .IN2(n6473), .QN(n6472) );
  OR2X1 U7534 ( .IN1(n4279), .IN2(DFF_183_n1), .Q(n6471) );
  NAND2X0 U7535 ( .IN1(n6474), .IN2(n6475), .QN(n6469) );
  NAND2X0 U7536 ( .IN1(n2153), .IN2(n6476), .QN(n6475) );
  NAND2X0 U7537 ( .IN1(WX498), .IN2(n4319), .QN(n6474) );
  OR2X1 U7538 ( .IN1(n6477), .IN2(n6478), .Q(WX658) );
  NAND2X0 U7539 ( .IN1(n6479), .IN2(n6480), .QN(n6478) );
  OR2X1 U7540 ( .IN1(n6481), .IN2(n4247), .Q(n6480) );
  OR2X1 U7541 ( .IN1(n4279), .IN2(DFF_184_n1), .Q(n6479) );
  NAND2X0 U7542 ( .IN1(n6482), .IN2(n6483), .QN(n6477) );
  NAND2X0 U7543 ( .IN1(n2153), .IN2(n6484), .QN(n6483) );
  NAND2X0 U7544 ( .IN1(WX496), .IN2(n4319), .QN(n6482) );
  OR2X1 U7545 ( .IN1(n6485), .IN2(n6486), .Q(WX656) );
  NAND2X0 U7546 ( .IN1(n6487), .IN2(n6488), .QN(n6486) );
  NAND2X0 U7547 ( .IN1(n4268), .IN2(n6489), .QN(n6488) );
  OR2X1 U7548 ( .IN1(n4278), .IN2(DFF_185_n1), .Q(n6487) );
  NAND2X0 U7549 ( .IN1(n6490), .IN2(n6491), .QN(n6485) );
  NAND2X0 U7550 ( .IN1(n2153), .IN2(n6492), .QN(n6491) );
  NAND2X0 U7551 ( .IN1(WX494), .IN2(n4319), .QN(n6490) );
  OR2X1 U7552 ( .IN1(n6493), .IN2(n6494), .Q(WX654) );
  NAND2X0 U7553 ( .IN1(n6495), .IN2(n6496), .QN(n6494) );
  NAND2X0 U7554 ( .IN1(n4268), .IN2(n6497), .QN(n6496) );
  OR2X1 U7555 ( .IN1(n4278), .IN2(DFF_186_n1), .Q(n6495) );
  NAND2X0 U7556 ( .IN1(n6498), .IN2(n6499), .QN(n6493) );
  NAND2X0 U7557 ( .IN1(n2153), .IN2(n6500), .QN(n6499) );
  NAND2X0 U7558 ( .IN1(WX492), .IN2(n4319), .QN(n6498) );
  OR2X1 U7559 ( .IN1(n6501), .IN2(n6502), .Q(WX652) );
  NAND2X0 U7560 ( .IN1(n6503), .IN2(n6504), .QN(n6502) );
  NAND2X0 U7561 ( .IN1(n4268), .IN2(n6505), .QN(n6504) );
  OR2X1 U7562 ( .IN1(n4278), .IN2(DFF_187_n1), .Q(n6503) );
  NAND2X0 U7563 ( .IN1(n6506), .IN2(n6507), .QN(n6501) );
  NAND2X0 U7564 ( .IN1(n2153), .IN2(n6508), .QN(n6507) );
  NAND2X0 U7565 ( .IN1(WX490), .IN2(n4319), .QN(n6506) );
  OR2X1 U7566 ( .IN1(n6509), .IN2(n6510), .Q(WX650) );
  NAND2X0 U7567 ( .IN1(n6511), .IN2(n6512), .QN(n6510) );
  OR2X1 U7568 ( .IN1(n6513), .IN2(n4247), .Q(n6512) );
  OR2X1 U7569 ( .IN1(n4278), .IN2(DFF_188_n1), .Q(n6511) );
  NAND2X0 U7570 ( .IN1(n6514), .IN2(n6515), .QN(n6509) );
  OR2X1 U7571 ( .IN1(n6516), .IN2(n4326), .Q(n6515) );
  NAND2X0 U7572 ( .IN1(WX488), .IN2(n4318), .QN(n6514) );
  NOR2X0 U7573 ( .IN1(n4938), .IN2(n6517), .QN(WX6498) );
  XOR2X1 U7574 ( .IN1(n4073), .IN2(DFF_958_n1), .Q(n6517) );
  NOR2X0 U7575 ( .IN1(n4938), .IN2(n6518), .QN(WX6496) );
  XOR2X1 U7576 ( .IN1(n4074), .IN2(DFF_957_n1), .Q(n6518) );
  NOR2X0 U7577 ( .IN1(n4938), .IN2(n6519), .QN(WX6494) );
  XOR2X1 U7578 ( .IN1(n4075), .IN2(DFF_956_n1), .Q(n6519) );
  NOR2X0 U7579 ( .IN1(n4939), .IN2(n6520), .QN(WX6492) );
  XOR2X1 U7580 ( .IN1(n4076), .IN2(DFF_955_n1), .Q(n6520) );
  NOR2X0 U7581 ( .IN1(n4939), .IN2(n6521), .QN(WX6490) );
  XOR2X1 U7582 ( .IN1(n4077), .IN2(DFF_954_n1), .Q(n6521) );
  NOR2X0 U7583 ( .IN1(n4939), .IN2(n6522), .QN(WX6488) );
  XOR2X1 U7584 ( .IN1(n4078), .IN2(DFF_953_n1), .Q(n6522) );
  NOR2X0 U7585 ( .IN1(n4939), .IN2(n6523), .QN(WX6486) );
  XOR2X1 U7586 ( .IN1(n4079), .IN2(DFF_952_n1), .Q(n6523) );
  NOR2X0 U7587 ( .IN1(n4939), .IN2(n6524), .QN(WX6484) );
  XOR2X1 U7588 ( .IN1(n4080), .IN2(DFF_951_n1), .Q(n6524) );
  NOR2X0 U7589 ( .IN1(n4939), .IN2(n6525), .QN(WX6482) );
  XOR2X1 U7590 ( .IN1(n4081), .IN2(DFF_950_n1), .Q(n6525) );
  NOR2X0 U7591 ( .IN1(n4939), .IN2(n6526), .QN(WX6480) );
  XOR2X1 U7592 ( .IN1(n4082), .IN2(DFF_949_n1), .Q(n6526) );
  OR2X1 U7593 ( .IN1(n6527), .IN2(n6528), .Q(WX648) );
  NAND2X0 U7594 ( .IN1(n6529), .IN2(n6530), .QN(n6528) );
  NAND2X0 U7595 ( .IN1(n4268), .IN2(n6531), .QN(n6530) );
  OR2X1 U7596 ( .IN1(n4278), .IN2(DFF_189_n1), .Q(n6529) );
  NAND2X0 U7597 ( .IN1(n6532), .IN2(n6533), .QN(n6527) );
  NAND2X0 U7598 ( .IN1(n2153), .IN2(n6534), .QN(n6533) );
  NAND2X0 U7599 ( .IN1(WX486), .IN2(n4318), .QN(n6532) );
  NOR2X0 U7600 ( .IN1(n4939), .IN2(n6535), .QN(WX6478) );
  XOR2X1 U7601 ( .IN1(n4083), .IN2(DFF_948_n1), .Q(n6535) );
  NOR2X0 U7602 ( .IN1(n4939), .IN2(n6536), .QN(WX6476) );
  XOR2X1 U7603 ( .IN1(n4084), .IN2(DFF_947_n1), .Q(n6536) );
  NOR2X0 U7604 ( .IN1(n4939), .IN2(n6537), .QN(WX6474) );
  XOR2X1 U7605 ( .IN1(n4085), .IN2(DFF_946_n1), .Q(n6537) );
  NOR2X0 U7606 ( .IN1(n4939), .IN2(n6538), .QN(WX6472) );
  XNOR2X1 U7607 ( .IN1(n4086), .IN2(test_so54), .Q(n6538) );
  NOR2X0 U7608 ( .IN1(n4939), .IN2(n6539), .QN(WX6470) );
  XOR2X1 U7609 ( .IN1(n4087), .IN2(DFF_944_n1), .Q(n6539) );
  NOR2X0 U7610 ( .IN1(n4939), .IN2(n6540), .QN(WX6468) );
  XOR2X1 U7611 ( .IN1(DFF_943_n1), .IN2(n6541), .Q(n6540) );
  XOR2X1 U7612 ( .IN1(test_so52), .IN2(DFF_959_n1), .Q(n6541) );
  NOR2X0 U7613 ( .IN1(n4940), .IN2(n6542), .QN(WX6466) );
  XOR2X1 U7614 ( .IN1(n4088), .IN2(DFF_942_n1), .Q(n6542) );
  NOR2X0 U7615 ( .IN1(n4940), .IN2(n6543), .QN(WX6464) );
  XOR2X1 U7616 ( .IN1(n4089), .IN2(DFF_941_n1), .Q(n6543) );
  NOR2X0 U7617 ( .IN1(n4940), .IN2(n6544), .QN(WX6462) );
  XOR2X1 U7618 ( .IN1(n4090), .IN2(DFF_940_n1), .Q(n6544) );
  NOR2X0 U7619 ( .IN1(n4940), .IN2(n6545), .QN(WX6460) );
  XOR2X1 U7620 ( .IN1(n4091), .IN2(DFF_939_n1), .Q(n6545) );
  OR2X1 U7621 ( .IN1(n6546), .IN2(n6547), .Q(WX646) );
  NAND2X0 U7622 ( .IN1(n6548), .IN2(n6549), .QN(n6547) );
  NAND2X0 U7623 ( .IN1(n4268), .IN2(n6550), .QN(n6549) );
  OR2X1 U7624 ( .IN1(n4278), .IN2(DFF_190_n1), .Q(n6548) );
  NAND2X0 U7625 ( .IN1(n6551), .IN2(n6552), .QN(n6546) );
  NAND2X0 U7626 ( .IN1(n2153), .IN2(n6553), .QN(n6552) );
  NAND2X0 U7627 ( .IN1(WX484), .IN2(n4318), .QN(n6551) );
  NOR2X0 U7628 ( .IN1(n4940), .IN2(n6554), .QN(WX6458) );
  XNOR2X1 U7629 ( .IN1(DFF_938_n1), .IN2(n6555), .Q(n6554) );
  XOR2X1 U7630 ( .IN1(n3950), .IN2(DFF_959_n1), .Q(n6555) );
  NOR2X0 U7631 ( .IN1(n4940), .IN2(n6556), .QN(WX6456) );
  XOR2X1 U7632 ( .IN1(n4092), .IN2(DFF_937_n1), .Q(n6556) );
  NOR2X0 U7633 ( .IN1(n4940), .IN2(n6557), .QN(WX6454) );
  XOR2X1 U7634 ( .IN1(n4093), .IN2(DFF_936_n1), .Q(n6557) );
  NOR2X0 U7635 ( .IN1(n4940), .IN2(n6558), .QN(WX6452) );
  XOR2X1 U7636 ( .IN1(n4094), .IN2(DFF_935_n1), .Q(n6558) );
  NOR2X0 U7637 ( .IN1(n4940), .IN2(n6559), .QN(WX6450) );
  XOR2X1 U7638 ( .IN1(n4095), .IN2(DFF_934_n1), .Q(n6559) );
  NOR2X0 U7639 ( .IN1(n4940), .IN2(n6560), .QN(WX6448) );
  XOR2X1 U7640 ( .IN1(n4096), .IN2(DFF_933_n1), .Q(n6560) );
  NOR2X0 U7641 ( .IN1(n4940), .IN2(n6561), .QN(WX6446) );
  XOR2X1 U7642 ( .IN1(n4097), .IN2(DFF_932_n1), .Q(n6561) );
  NOR2X0 U7643 ( .IN1(n4940), .IN2(n6562), .QN(WX6444) );
  XNOR2X1 U7644 ( .IN1(DFF_931_n1), .IN2(n6563), .Q(n6562) );
  XOR2X1 U7645 ( .IN1(n3951), .IN2(DFF_959_n1), .Q(n6563) );
  NOR2X0 U7646 ( .IN1(n4941), .IN2(n6564), .QN(WX6442) );
  XOR2X1 U7647 ( .IN1(n4098), .IN2(DFF_930_n1), .Q(n6564) );
  NOR2X0 U7648 ( .IN1(n4941), .IN2(n6565), .QN(WX6440) );
  XOR2X1 U7649 ( .IN1(n4099), .IN2(DFF_929_n1), .Q(n6565) );
  NAND2X0 U7650 ( .IN1(n6566), .IN2(n6567), .QN(WX644) );
  NOR2X0 U7651 ( .IN1(n6568), .IN2(n6569), .QN(n6567) );
  NOR2X0 U7652 ( .IN1(n6570), .IN2(n4252), .QN(n6569) );
  NOR2X0 U7653 ( .IN1(n6571), .IN2(n4330), .QN(n6568) );
  NOR2X0 U7654 ( .IN1(n6572), .IN2(n6573), .QN(n6566) );
  NOR2X0 U7655 ( .IN1(n3930), .IN2(n5606), .QN(n6573) );
  NOR2X0 U7656 ( .IN1(DFF_191_n1), .IN2(n4280), .QN(n6572) );
  NOR2X0 U7657 ( .IN1(n4941), .IN2(n6574), .QN(WX6438) );
  XNOR2X1 U7658 ( .IN1(n4100), .IN2(test_so53), .Q(n6574) );
  NOR2X0 U7659 ( .IN1(n4941), .IN2(n6575), .QN(WX6436) );
  XOR2X1 U7660 ( .IN1(n3964), .IN2(DFF_959_n1), .Q(n6575) );
  NOR2X0 U7661 ( .IN1(n8926), .IN2(n4851), .QN(WX5910) );
  NOR2X0 U7662 ( .IN1(n8927), .IN2(n4852), .QN(WX5908) );
  NOR2X0 U7663 ( .IN1(n8928), .IN2(n4852), .QN(WX5906) );
  NOR2X0 U7664 ( .IN1(n8931), .IN2(n4852), .QN(WX5904) );
  NOR2X0 U7665 ( .IN1(n8932), .IN2(n4852), .QN(WX5902) );
  NOR2X0 U7666 ( .IN1(n8935), .IN2(n4852), .QN(WX5900) );
  AND2X1 U7667 ( .IN1(n4800), .IN2(test_so46), .Q(WX5898) );
  NOR2X0 U7668 ( .IN1(n8936), .IN2(n4852), .QN(WX5896) );
  NOR2X0 U7669 ( .IN1(n8937), .IN2(n4852), .QN(WX5894) );
  NOR2X0 U7670 ( .IN1(n8938), .IN2(n4852), .QN(WX5892) );
  NOR2X0 U7671 ( .IN1(n8939), .IN2(n4852), .QN(WX5890) );
  NOR2X0 U7672 ( .IN1(n8940), .IN2(n4852), .QN(WX5888) );
  NOR2X0 U7673 ( .IN1(n8941), .IN2(n4852), .QN(WX5886) );
  NOR2X0 U7674 ( .IN1(n8942), .IN2(n4852), .QN(WX5884) );
  NOR2X0 U7675 ( .IN1(n8943), .IN2(n4853), .QN(WX5882) );
  NOR2X0 U7676 ( .IN1(n8944), .IN2(n4923), .QN(WX5880) );
  NAND2X0 U7677 ( .IN1(n6576), .IN2(n6577), .QN(WX5878) );
  NOR2X0 U7678 ( .IN1(n6578), .IN2(n6579), .QN(n6577) );
  NOR2X0 U7679 ( .IN1(n6580), .IN2(n4252), .QN(n6579) );
  NOR2X0 U7680 ( .IN1(n5985), .IN2(n4330), .QN(n6578) );
  XOR2X1 U7681 ( .IN1(n6581), .IN2(n6582), .Q(n5985) );
  XOR2X1 U7682 ( .IN1(n8875), .IN2(n3963), .Q(n6582) );
  XOR2X1 U7683 ( .IN1(WX7172), .IN2(n3785), .Q(n6581) );
  NOR2X0 U7684 ( .IN1(n6583), .IN2(n6584), .QN(n6576) );
  AND2X1 U7685 ( .IN1(n2152), .IN2(test_so53), .Q(n6584) );
  NOR2X0 U7686 ( .IN1(n4306), .IN2(n5317), .QN(n6583) );
  NAND2X0 U7687 ( .IN1(n4823), .IN2(n8496), .QN(n5317) );
  NAND2X0 U7688 ( .IN1(n6585), .IN2(n6586), .QN(WX5876) );
  NOR2X0 U7689 ( .IN1(n6587), .IN2(n6588), .QN(n6586) );
  NOR2X0 U7690 ( .IN1(n5352), .IN2(n6589), .QN(n6588) );
  NOR2X0 U7691 ( .IN1(n5994), .IN2(n4330), .QN(n6587) );
  XOR2X1 U7692 ( .IN1(n6590), .IN2(n6591), .Q(n5994) );
  XOR2X1 U7693 ( .IN1(n8876), .IN2(n4072), .Q(n6591) );
  XOR2X1 U7694 ( .IN1(WX7170), .IN2(n3787), .Q(n6590) );
  NOR2X0 U7695 ( .IN1(n6592), .IN2(n6593), .QN(n6585) );
  NOR2X0 U7696 ( .IN1(DFF_929_n1), .IN2(n4283), .QN(n6593) );
  NOR2X0 U7697 ( .IN1(n4306), .IN2(n5318), .QN(n6592) );
  NAND2X0 U7698 ( .IN1(n4823), .IN2(n8497), .QN(n5318) );
  NAND2X0 U7699 ( .IN1(n6594), .IN2(n6595), .QN(WX5874) );
  NOR2X0 U7700 ( .IN1(n6596), .IN2(n6597), .QN(n6595) );
  NOR2X0 U7701 ( .IN1(n6598), .IN2(n4252), .QN(n6597) );
  NOR2X0 U7702 ( .IN1(n6003), .IN2(n4330), .QN(n6596) );
  XOR2X1 U7703 ( .IN1(n6599), .IN2(n6600), .Q(n6003) );
  XOR2X1 U7704 ( .IN1(n8877), .IN2(n4071), .Q(n6600) );
  XOR2X1 U7705 ( .IN1(WX7168), .IN2(n3789), .Q(n6599) );
  NOR2X0 U7706 ( .IN1(n6601), .IN2(n6602), .QN(n6594) );
  NOR2X0 U7707 ( .IN1(DFF_930_n1), .IN2(n4295), .QN(n6602) );
  NOR2X0 U7708 ( .IN1(n4306), .IN2(n5319), .QN(n6601) );
  NAND2X0 U7709 ( .IN1(n4823), .IN2(n8498), .QN(n5319) );
  NAND2X0 U7710 ( .IN1(n6603), .IN2(n6604), .QN(WX5872) );
  NOR2X0 U7711 ( .IN1(n6605), .IN2(n6606), .QN(n6604) );
  NOR2X0 U7712 ( .IN1(n5352), .IN2(n6607), .QN(n6606) );
  NOR2X0 U7713 ( .IN1(n6012), .IN2(n4330), .QN(n6605) );
  XOR2X1 U7714 ( .IN1(n6608), .IN2(n6609), .Q(n6012) );
  XOR2X1 U7715 ( .IN1(n8878), .IN2(n4070), .Q(n6609) );
  XOR2X1 U7716 ( .IN1(WX7166), .IN2(n3791), .Q(n6608) );
  NOR2X0 U7717 ( .IN1(n6610), .IN2(n6611), .QN(n6603) );
  NOR2X0 U7718 ( .IN1(DFF_931_n1), .IN2(n4295), .QN(n6611) );
  NOR2X0 U7719 ( .IN1(n4306), .IN2(n5320), .QN(n6610) );
  NAND2X0 U7720 ( .IN1(n4823), .IN2(n8499), .QN(n5320) );
  NAND2X0 U7721 ( .IN1(n6612), .IN2(n6613), .QN(WX5870) );
  NOR2X0 U7722 ( .IN1(n6614), .IN2(n6615), .QN(n6613) );
  NOR2X0 U7723 ( .IN1(n6616), .IN2(n4252), .QN(n6615) );
  NOR2X0 U7724 ( .IN1(n4338), .IN2(n6021), .QN(n6614) );
  XNOR2X1 U7725 ( .IN1(n6617), .IN2(n6618), .Q(n6021) );
  XOR2X1 U7726 ( .IN1(test_so64), .IN2(n8879), .Q(n6618) );
  XOR2X1 U7727 ( .IN1(WX7164), .IN2(n3793), .Q(n6617) );
  NOR2X0 U7728 ( .IN1(n6619), .IN2(n6620), .QN(n6612) );
  NOR2X0 U7729 ( .IN1(DFF_932_n1), .IN2(n4295), .QN(n6620) );
  NOR2X0 U7730 ( .IN1(n4305), .IN2(n5321), .QN(n6619) );
  NAND2X0 U7731 ( .IN1(n4823), .IN2(n8500), .QN(n5321) );
  NAND2X0 U7732 ( .IN1(n6621), .IN2(n6622), .QN(WX5868) );
  NOR2X0 U7733 ( .IN1(n6623), .IN2(n6624), .QN(n6622) );
  NOR2X0 U7734 ( .IN1(n5352), .IN2(n6625), .QN(n6624) );
  NOR2X0 U7735 ( .IN1(n6030), .IN2(n4330), .QN(n6623) );
  XOR2X1 U7736 ( .IN1(n6626), .IN2(n6627), .Q(n6030) );
  XOR2X1 U7737 ( .IN1(n8880), .IN2(n4069), .Q(n6627) );
  XOR2X1 U7738 ( .IN1(WX7162), .IN2(n3795), .Q(n6626) );
  NOR2X0 U7739 ( .IN1(n6628), .IN2(n6629), .QN(n6621) );
  NOR2X0 U7740 ( .IN1(DFF_933_n1), .IN2(n4295), .QN(n6629) );
  NOR2X0 U7741 ( .IN1(n4305), .IN2(n5322), .QN(n6628) );
  NAND2X0 U7742 ( .IN1(n4823), .IN2(n8501), .QN(n5322) );
  NAND2X0 U7743 ( .IN1(n6630), .IN2(n6631), .QN(WX5866) );
  NOR2X0 U7744 ( .IN1(n6632), .IN2(n6633), .QN(n6631) );
  NOR2X0 U7745 ( .IN1(n6634), .IN2(n4252), .QN(n6633) );
  NOR2X0 U7746 ( .IN1(n4337), .IN2(n6039), .QN(n6632) );
  XNOR2X1 U7747 ( .IN1(n6635), .IN2(n6636), .Q(n6039) );
  XOR2X1 U7748 ( .IN1(test_so62), .IN2(n8881), .Q(n6636) );
  XOR2X1 U7749 ( .IN1(WX7160), .IN2(n4068), .Q(n6635) );
  NOR2X0 U7750 ( .IN1(n6637), .IN2(n6638), .QN(n6630) );
  NOR2X0 U7751 ( .IN1(DFF_934_n1), .IN2(n4295), .QN(n6638) );
  NOR2X0 U7752 ( .IN1(n4305), .IN2(n5324), .QN(n6637) );
  NAND2X0 U7753 ( .IN1(n4822), .IN2(n8502), .QN(n5324) );
  NAND2X0 U7754 ( .IN1(n6639), .IN2(n6640), .QN(WX5864) );
  NOR2X0 U7755 ( .IN1(n6641), .IN2(n6642), .QN(n6640) );
  NOR2X0 U7756 ( .IN1(n6643), .IN2(n4252), .QN(n6642) );
  NOR2X0 U7757 ( .IN1(n6048), .IN2(n4330), .QN(n6641) );
  XOR2X1 U7758 ( .IN1(n6644), .IN2(n6645), .Q(n6048) );
  XOR2X1 U7759 ( .IN1(n8882), .IN2(n4067), .Q(n6645) );
  XOR2X1 U7760 ( .IN1(WX7158), .IN2(n3798), .Q(n6644) );
  NOR2X0 U7761 ( .IN1(n6646), .IN2(n6647), .QN(n6639) );
  NOR2X0 U7762 ( .IN1(DFF_935_n1), .IN2(n4295), .QN(n6647) );
  NOR2X0 U7763 ( .IN1(n4305), .IN2(n5325), .QN(n6646) );
  NAND2X0 U7764 ( .IN1(test_so45), .IN2(n4828), .QN(n5325) );
  NAND2X0 U7765 ( .IN1(n6648), .IN2(n6649), .QN(WX5862) );
  NOR2X0 U7766 ( .IN1(n6650), .IN2(n6651), .QN(n6649) );
  NOR2X0 U7767 ( .IN1(n6652), .IN2(n4252), .QN(n6651) );
  NOR2X0 U7768 ( .IN1(n4338), .IN2(n6057), .QN(n6650) );
  XNOR2X1 U7769 ( .IN1(n6653), .IN2(n6654), .Q(n6057) );
  XOR2X1 U7770 ( .IN1(test_so60), .IN2(n8883), .Q(n6654) );
  XOR2X1 U7771 ( .IN1(WX7156), .IN2(n4066), .Q(n6653) );
  NOR2X0 U7772 ( .IN1(n6655), .IN2(n6656), .QN(n6648) );
  NOR2X0 U7773 ( .IN1(DFF_936_n1), .IN2(n4295), .QN(n6656) );
  NOR2X0 U7774 ( .IN1(n4305), .IN2(n5326), .QN(n6655) );
  NAND2X0 U7775 ( .IN1(n4823), .IN2(n8505), .QN(n5326) );
  NAND2X0 U7776 ( .IN1(n6657), .IN2(n6658), .QN(WX5860) );
  NOR2X0 U7777 ( .IN1(n6659), .IN2(n6660), .QN(n6658) );
  NOR2X0 U7778 ( .IN1(n6661), .IN2(n4253), .QN(n6660) );
  NOR2X0 U7779 ( .IN1(n6066), .IN2(n4330), .QN(n6659) );
  XOR2X1 U7780 ( .IN1(n6662), .IN2(n6663), .Q(n6066) );
  XOR2X1 U7781 ( .IN1(n8884), .IN2(n4065), .Q(n6663) );
  XOR2X1 U7782 ( .IN1(WX7154), .IN2(n3801), .Q(n6662) );
  NOR2X0 U7783 ( .IN1(n6664), .IN2(n6665), .QN(n6657) );
  NOR2X0 U7784 ( .IN1(DFF_937_n1), .IN2(n4295), .QN(n6665) );
  NOR2X0 U7785 ( .IN1(n4305), .IN2(n5327), .QN(n6664) );
  NAND2X0 U7786 ( .IN1(n4822), .IN2(n8506), .QN(n5327) );
  NAND2X0 U7787 ( .IN1(n6666), .IN2(n6667), .QN(WX5858) );
  NOR2X0 U7788 ( .IN1(n6668), .IN2(n6669), .QN(n6667) );
  NOR2X0 U7789 ( .IN1(n6670), .IN2(n4253), .QN(n6669) );
  NOR2X0 U7790 ( .IN1(n4338), .IN2(n6075), .QN(n6668) );
  XNOR2X1 U7791 ( .IN1(n6671), .IN2(n6672), .Q(n6075) );
  XOR2X1 U7792 ( .IN1(test_so58), .IN2(n8885), .Q(n6672) );
  XOR2X1 U7793 ( .IN1(WX7280), .IN2(n4064), .Q(n6671) );
  NOR2X0 U7794 ( .IN1(n6673), .IN2(n6674), .QN(n6666) );
  NOR2X0 U7795 ( .IN1(DFF_938_n1), .IN2(n4295), .QN(n6674) );
  NOR2X0 U7796 ( .IN1(n4305), .IN2(n5328), .QN(n6673) );
  NAND2X0 U7797 ( .IN1(n4822), .IN2(n8507), .QN(n5328) );
  NAND2X0 U7798 ( .IN1(n6675), .IN2(n6676), .QN(WX5856) );
  NOR2X0 U7799 ( .IN1(n6677), .IN2(n6678), .QN(n6676) );
  NOR2X0 U7800 ( .IN1(n6679), .IN2(n4253), .QN(n6678) );
  NOR2X0 U7801 ( .IN1(n6084), .IN2(n4330), .QN(n6677) );
  XOR2X1 U7802 ( .IN1(n6680), .IN2(n6681), .Q(n6084) );
  XOR2X1 U7803 ( .IN1(n8886), .IN2(n3949), .Q(n6681) );
  XOR2X1 U7804 ( .IN1(WX7150), .IN2(n3804), .Q(n6680) );
  NOR2X0 U7805 ( .IN1(n6682), .IN2(n6683), .QN(n6675) );
  NOR2X0 U7806 ( .IN1(DFF_939_n1), .IN2(n4295), .QN(n6683) );
  NOR2X0 U7807 ( .IN1(n4305), .IN2(n5329), .QN(n6682) );
  NAND2X0 U7808 ( .IN1(n4822), .IN2(n8508), .QN(n5329) );
  NAND2X0 U7809 ( .IN1(n6684), .IN2(n6685), .QN(WX5854) );
  NOR2X0 U7810 ( .IN1(n6686), .IN2(n6687), .QN(n6685) );
  NOR2X0 U7811 ( .IN1(n6688), .IN2(n4253), .QN(n6687) );
  NOR2X0 U7812 ( .IN1(n6093), .IN2(n4330), .QN(n6686) );
  XOR2X1 U7813 ( .IN1(n6689), .IN2(n6690), .Q(n6093) );
  XOR2X1 U7814 ( .IN1(n8887), .IN2(n4063), .Q(n6690) );
  XOR2X1 U7815 ( .IN1(WX7148), .IN2(n3806), .Q(n6689) );
  NOR2X0 U7816 ( .IN1(n6691), .IN2(n6692), .QN(n6684) );
  NOR2X0 U7817 ( .IN1(DFF_940_n1), .IN2(n4294), .QN(n6692) );
  NOR2X0 U7818 ( .IN1(n4305), .IN2(n5330), .QN(n6691) );
  NAND2X0 U7819 ( .IN1(n4822), .IN2(n8509), .QN(n5330) );
  NAND2X0 U7820 ( .IN1(n6693), .IN2(n6694), .QN(WX5852) );
  NOR2X0 U7821 ( .IN1(n6695), .IN2(n6696), .QN(n6694) );
  NOR2X0 U7822 ( .IN1(n6697), .IN2(n4253), .QN(n6696) );
  NOR2X0 U7823 ( .IN1(n6102), .IN2(n4330), .QN(n6695) );
  XOR2X1 U7824 ( .IN1(n6698), .IN2(n6699), .Q(n6102) );
  XOR2X1 U7825 ( .IN1(n8888), .IN2(n4062), .Q(n6699) );
  XOR2X1 U7826 ( .IN1(WX7146), .IN2(n3808), .Q(n6698) );
  NOR2X0 U7827 ( .IN1(n6700), .IN2(n6701), .QN(n6693) );
  NOR2X0 U7828 ( .IN1(DFF_941_n1), .IN2(n4295), .QN(n6701) );
  NOR2X0 U7829 ( .IN1(n4305), .IN2(n5331), .QN(n6700) );
  NAND2X0 U7830 ( .IN1(n4822), .IN2(n8510), .QN(n5331) );
  NAND2X0 U7831 ( .IN1(n6702), .IN2(n6703), .QN(WX5850) );
  NOR2X0 U7832 ( .IN1(n6704), .IN2(n6705), .QN(n6703) );
  NOR2X0 U7833 ( .IN1(n6706), .IN2(n4253), .QN(n6705) );
  NOR2X0 U7834 ( .IN1(n6111), .IN2(n4331), .QN(n6704) );
  XOR2X1 U7835 ( .IN1(n6707), .IN2(n6708), .Q(n6111) );
  XOR2X1 U7836 ( .IN1(n8889), .IN2(n4061), .Q(n6708) );
  XOR2X1 U7837 ( .IN1(WX7144), .IN2(n3810), .Q(n6707) );
  NOR2X0 U7838 ( .IN1(n6709), .IN2(n6710), .QN(n6702) );
  NOR2X0 U7839 ( .IN1(DFF_942_n1), .IN2(n4295), .QN(n6710) );
  NOR2X0 U7840 ( .IN1(n4305), .IN2(n5332), .QN(n6709) );
  NAND2X0 U7841 ( .IN1(n4822), .IN2(n8511), .QN(n5332) );
  NAND2X0 U7842 ( .IN1(n6711), .IN2(n6712), .QN(WX5848) );
  NOR2X0 U7843 ( .IN1(n6713), .IN2(n6714), .QN(n6712) );
  NOR2X0 U7844 ( .IN1(n6715), .IN2(n4253), .QN(n6714) );
  NOR2X0 U7845 ( .IN1(n6120), .IN2(n4331), .QN(n6713) );
  XOR2X1 U7846 ( .IN1(n6716), .IN2(n6717), .Q(n6120) );
  XOR2X1 U7847 ( .IN1(n8890), .IN2(n4060), .Q(n6717) );
  XOR2X1 U7848 ( .IN1(WX7142), .IN2(n3812), .Q(n6716) );
  NOR2X0 U7849 ( .IN1(n6718), .IN2(n6719), .QN(n6711) );
  NOR2X0 U7850 ( .IN1(DFF_943_n1), .IN2(n4295), .QN(n6719) );
  NOR2X0 U7851 ( .IN1(n4305), .IN2(n5333), .QN(n6718) );
  NAND2X0 U7852 ( .IN1(n4822), .IN2(n8512), .QN(n5333) );
  NAND2X0 U7853 ( .IN1(n6720), .IN2(n6721), .QN(WX5846) );
  NOR2X0 U7854 ( .IN1(n6722), .IN2(n6723), .QN(n6721) );
  NOR2X0 U7855 ( .IN1(n4258), .IN2(n6724), .QN(n6723) );
  NOR2X0 U7856 ( .IN1(n6129), .IN2(n4331), .QN(n6722) );
  XOR2X1 U7857 ( .IN1(n6725), .IN2(n6726), .Q(n6129) );
  XOR2X1 U7858 ( .IN1(n3629), .IN2(n4773), .Q(n6726) );
  XOR2X1 U7859 ( .IN1(n6727), .IN2(n3948), .Q(n6725) );
  XOR2X1 U7860 ( .IN1(WX7268), .IN2(n8891), .Q(n6727) );
  NOR2X0 U7861 ( .IN1(n6728), .IN2(n6729), .QN(n6720) );
  NOR2X0 U7862 ( .IN1(DFF_944_n1), .IN2(n4294), .QN(n6729) );
  NOR2X0 U7863 ( .IN1(n4304), .IN2(n5335), .QN(n6728) );
  NAND2X0 U7864 ( .IN1(n4821), .IN2(n8513), .QN(n5335) );
  NAND2X0 U7865 ( .IN1(n6730), .IN2(n6731), .QN(WX5844) );
  NOR2X0 U7866 ( .IN1(n6732), .IN2(n6733), .QN(n6731) );
  NOR2X0 U7867 ( .IN1(n6734), .IN2(n4253), .QN(n6733) );
  NOR2X0 U7868 ( .IN1(n6139), .IN2(n4331), .QN(n6732) );
  XOR2X1 U7869 ( .IN1(n6735), .IN2(n6736), .Q(n6139) );
  XOR2X1 U7870 ( .IN1(n3630), .IN2(n4773), .Q(n6736) );
  XOR2X1 U7871 ( .IN1(n6737), .IN2(n4059), .Q(n6735) );
  XOR2X1 U7872 ( .IN1(WX7266), .IN2(n8892), .Q(n6737) );
  NOR2X0 U7873 ( .IN1(n6738), .IN2(n6739), .QN(n6730) );
  AND2X1 U7874 ( .IN1(n2152), .IN2(test_so54), .Q(n6739) );
  NOR2X0 U7875 ( .IN1(n4304), .IN2(n5336), .QN(n6738) );
  NAND2X0 U7876 ( .IN1(n4822), .IN2(n8514), .QN(n5336) );
  NAND2X0 U7877 ( .IN1(n6740), .IN2(n6741), .QN(WX5842) );
  NOR2X0 U7878 ( .IN1(n6742), .IN2(n6743), .QN(n6741) );
  NOR2X0 U7879 ( .IN1(n5352), .IN2(n6744), .QN(n6743) );
  NOR2X0 U7880 ( .IN1(n6149), .IN2(n4331), .QN(n6742) );
  XOR2X1 U7881 ( .IN1(n6745), .IN2(n6746), .Q(n6149) );
  XOR2X1 U7882 ( .IN1(n3631), .IN2(n4773), .Q(n6746) );
  XOR2X1 U7883 ( .IN1(n6747), .IN2(n4058), .Q(n6745) );
  XOR2X1 U7884 ( .IN1(WX7264), .IN2(n8893), .Q(n6747) );
  NOR2X0 U7885 ( .IN1(n6748), .IN2(n6749), .QN(n6740) );
  NOR2X0 U7886 ( .IN1(DFF_946_n1), .IN2(n4294), .QN(n6749) );
  NOR2X0 U7887 ( .IN1(n4304), .IN2(n5337), .QN(n6748) );
  NAND2X0 U7888 ( .IN1(n4821), .IN2(n8515), .QN(n5337) );
  NAND2X0 U7889 ( .IN1(n6750), .IN2(n6751), .QN(WX5840) );
  NOR2X0 U7890 ( .IN1(n6752), .IN2(n6753), .QN(n6751) );
  NOR2X0 U7891 ( .IN1(n6754), .IN2(n4253), .QN(n6753) );
  NOR2X0 U7892 ( .IN1(n6159), .IN2(n4331), .QN(n6752) );
  XOR2X1 U7893 ( .IN1(n6755), .IN2(n6756), .Q(n6159) );
  XOR2X1 U7894 ( .IN1(n3632), .IN2(n4777), .Q(n6756) );
  XOR2X1 U7895 ( .IN1(n6757), .IN2(n4057), .Q(n6755) );
  XOR2X1 U7896 ( .IN1(WX7262), .IN2(n8894), .Q(n6757) );
  NOR2X0 U7897 ( .IN1(n6758), .IN2(n6759), .QN(n6750) );
  NOR2X0 U7898 ( .IN1(DFF_947_n1), .IN2(n4294), .QN(n6759) );
  NOR2X0 U7899 ( .IN1(n4304), .IN2(n5338), .QN(n6758) );
  NAND2X0 U7900 ( .IN1(n4821), .IN2(n8516), .QN(n5338) );
  NAND2X0 U7901 ( .IN1(n6760), .IN2(n6761), .QN(WX5838) );
  NOR2X0 U7902 ( .IN1(n6762), .IN2(n6763), .QN(n6761) );
  NOR2X0 U7903 ( .IN1(n5352), .IN2(n6764), .QN(n6763) );
  NOR2X0 U7904 ( .IN1(n6169), .IN2(n4331), .QN(n6762) );
  XOR2X1 U7905 ( .IN1(n6765), .IN2(n6766), .Q(n6169) );
  XOR2X1 U7906 ( .IN1(n3633), .IN2(n4774), .Q(n6766) );
  XOR2X1 U7907 ( .IN1(n6767), .IN2(n4056), .Q(n6765) );
  XOR2X1 U7908 ( .IN1(WX7260), .IN2(n8895), .Q(n6767) );
  NOR2X0 U7909 ( .IN1(n6768), .IN2(n6769), .QN(n6760) );
  NOR2X0 U7910 ( .IN1(DFF_948_n1), .IN2(n4294), .QN(n6769) );
  NOR2X0 U7911 ( .IN1(n4304), .IN2(n5339), .QN(n6768) );
  NAND2X0 U7912 ( .IN1(n4821), .IN2(n8517), .QN(n5339) );
  NAND2X0 U7913 ( .IN1(n6770), .IN2(n6771), .QN(WX5836) );
  NOR2X0 U7914 ( .IN1(n6772), .IN2(n6773), .QN(n6771) );
  NOR2X0 U7915 ( .IN1(n6774), .IN2(n4254), .QN(n6773) );
  NOR2X0 U7916 ( .IN1(n4339), .IN2(n6179), .QN(n6772) );
  XNOR2X1 U7917 ( .IN1(n6775), .IN2(n6776), .Q(n6179) );
  XOR2X1 U7918 ( .IN1(n3634), .IN2(n4774), .Q(n6776) );
  XOR2X1 U7919 ( .IN1(WX7194), .IN2(n6777), .Q(n6775) );
  XOR2X1 U7920 ( .IN1(test_so63), .IN2(n8896), .Q(n6777) );
  NOR2X0 U7921 ( .IN1(n6778), .IN2(n6779), .QN(n6770) );
  NOR2X0 U7922 ( .IN1(DFF_949_n1), .IN2(n4294), .QN(n6779) );
  NOR2X0 U7923 ( .IN1(n4304), .IN2(n5340), .QN(n6778) );
  NAND2X0 U7924 ( .IN1(n4821), .IN2(n8518), .QN(n5340) );
  NAND2X0 U7925 ( .IN1(n6780), .IN2(n6781), .QN(WX5834) );
  NOR2X0 U7926 ( .IN1(n6782), .IN2(n6783), .QN(n6781) );
  NOR2X0 U7927 ( .IN1(n5352), .IN2(n6784), .QN(n6783) );
  NOR2X0 U7928 ( .IN1(n6189), .IN2(n4331), .QN(n6782) );
  XOR2X1 U7929 ( .IN1(n6785), .IN2(n6786), .Q(n6189) );
  XOR2X1 U7930 ( .IN1(n3635), .IN2(n4774), .Q(n6786) );
  XOR2X1 U7931 ( .IN1(n6787), .IN2(n4055), .Q(n6785) );
  XOR2X1 U7932 ( .IN1(WX7256), .IN2(n8897), .Q(n6787) );
  NOR2X0 U7933 ( .IN1(n6788), .IN2(n6789), .QN(n6780) );
  NOR2X0 U7934 ( .IN1(DFF_950_n1), .IN2(n4294), .QN(n6789) );
  NOR2X0 U7935 ( .IN1(n4304), .IN2(n5341), .QN(n6788) );
  NAND2X0 U7936 ( .IN1(n4821), .IN2(n8519), .QN(n5341) );
  NAND2X0 U7937 ( .IN1(n6790), .IN2(n6791), .QN(WX5832) );
  NOR2X0 U7938 ( .IN1(n6792), .IN2(n6793), .QN(n6791) );
  NOR2X0 U7939 ( .IN1(n6794), .IN2(n4253), .QN(n6793) );
  NOR2X0 U7940 ( .IN1(n4338), .IN2(n6199), .QN(n6792) );
  XNOR2X1 U7941 ( .IN1(n6795), .IN2(n6796), .Q(n6199) );
  XOR2X1 U7942 ( .IN1(n4054), .IN2(n4774), .Q(n6796) );
  XOR2X1 U7943 ( .IN1(n6797), .IN2(n8900), .Q(n6795) );
  XOR2X1 U7944 ( .IN1(n8899), .IN2(n8898), .Q(n6797) );
  NOR2X0 U7945 ( .IN1(n6798), .IN2(n6799), .QN(n6790) );
  NOR2X0 U7946 ( .IN1(DFF_951_n1), .IN2(n4294), .QN(n6799) );
  NOR2X0 U7947 ( .IN1(n4304), .IN2(n5342), .QN(n6798) );
  NAND2X0 U7948 ( .IN1(n4821), .IN2(n8520), .QN(n5342) );
  NAND2X0 U7949 ( .IN1(n6800), .IN2(n6801), .QN(WX5830) );
  NOR2X0 U7950 ( .IN1(n6802), .IN2(n6803), .QN(n6801) );
  NOR2X0 U7951 ( .IN1(n6804), .IN2(n4254), .QN(n6803) );
  NOR2X0 U7952 ( .IN1(n6209), .IN2(n4331), .QN(n6802) );
  XOR2X1 U7953 ( .IN1(n6805), .IN2(n6806), .Q(n6209) );
  XOR2X1 U7954 ( .IN1(n3636), .IN2(n4774), .Q(n6806) );
  XOR2X1 U7955 ( .IN1(n6807), .IN2(n4053), .Q(n6805) );
  XOR2X1 U7956 ( .IN1(WX7252), .IN2(n8901), .Q(n6807) );
  NOR2X0 U7957 ( .IN1(n6808), .IN2(n6809), .QN(n6800) );
  NOR2X0 U7958 ( .IN1(DFF_952_n1), .IN2(n4294), .QN(n6809) );
  NOR2X0 U7959 ( .IN1(n4304), .IN2(n5343), .QN(n6808) );
  NAND2X0 U7960 ( .IN1(test_so44), .IN2(n4827), .QN(n5343) );
  NAND2X0 U7961 ( .IN1(n6810), .IN2(n6811), .QN(WX5828) );
  NOR2X0 U7962 ( .IN1(n6812), .IN2(n6813), .QN(n6811) );
  NOR2X0 U7963 ( .IN1(n6814), .IN2(n4254), .QN(n6813) );
  NOR2X0 U7964 ( .IN1(n4339), .IN2(n6219), .QN(n6812) );
  XNOR2X1 U7965 ( .IN1(n6815), .IN2(n6816), .Q(n6219) );
  XOR2X1 U7966 ( .IN1(n4052), .IN2(n4774), .Q(n6816) );
  XOR2X1 U7967 ( .IN1(n6817), .IN2(n8904), .Q(n6815) );
  XOR2X1 U7968 ( .IN1(n8903), .IN2(n8902), .Q(n6817) );
  NOR2X0 U7969 ( .IN1(n6818), .IN2(n6819), .QN(n6810) );
  NOR2X0 U7970 ( .IN1(DFF_953_n1), .IN2(n4294), .QN(n6819) );
  NOR2X0 U7971 ( .IN1(n4304), .IN2(n5344), .QN(n6818) );
  NAND2X0 U7972 ( .IN1(n4821), .IN2(n8523), .QN(n5344) );
  NAND2X0 U7973 ( .IN1(n6820), .IN2(n6821), .QN(WX5826) );
  NOR2X0 U7974 ( .IN1(n6822), .IN2(n6823), .QN(n6821) );
  NOR2X0 U7975 ( .IN1(n6824), .IN2(n4253), .QN(n6823) );
  NOR2X0 U7976 ( .IN1(n6229), .IN2(n4331), .QN(n6822) );
  XOR2X1 U7977 ( .IN1(n6825), .IN2(n6826), .Q(n6229) );
  XOR2X1 U7978 ( .IN1(n3637), .IN2(n4774), .Q(n6826) );
  XOR2X1 U7979 ( .IN1(n6827), .IN2(n4051), .Q(n6825) );
  XOR2X1 U7980 ( .IN1(WX7248), .IN2(n8905), .Q(n6827) );
  NOR2X0 U7981 ( .IN1(n6828), .IN2(n6829), .QN(n6820) );
  NOR2X0 U7982 ( .IN1(DFF_954_n1), .IN2(n4294), .QN(n6829) );
  NOR2X0 U7983 ( .IN1(n4304), .IN2(n5129), .QN(n6828) );
  NAND2X0 U7984 ( .IN1(n4821), .IN2(n8524), .QN(n5129) );
  NAND2X0 U7985 ( .IN1(n6830), .IN2(n6831), .QN(WX5824) );
  NOR2X0 U7986 ( .IN1(n6832), .IN2(n6833), .QN(n6831) );
  NOR2X0 U7987 ( .IN1(n6834), .IN2(n4254), .QN(n6833) );
  NOR2X0 U7988 ( .IN1(n4339), .IN2(n6239), .QN(n6832) );
  XNOR2X1 U7989 ( .IN1(n6835), .IN2(n6836), .Q(n6239) );
  XOR2X1 U7990 ( .IN1(n3638), .IN2(n4774), .Q(n6836) );
  XOR2X1 U7991 ( .IN1(n6837), .IN2(n4050), .Q(n6835) );
  XOR2X1 U7992 ( .IN1(WX7182), .IN2(test_so57), .Q(n6837) );
  NOR2X0 U7993 ( .IN1(n6838), .IN2(n6839), .QN(n6830) );
  NOR2X0 U7994 ( .IN1(DFF_955_n1), .IN2(n4294), .QN(n6839) );
  NOR2X0 U7995 ( .IN1(n4304), .IN2(n5130), .QN(n6838) );
  NAND2X0 U7996 ( .IN1(n4820), .IN2(n8525), .QN(n5130) );
  NAND2X0 U7997 ( .IN1(n6840), .IN2(n6841), .QN(WX5822) );
  NOR2X0 U7998 ( .IN1(n6842), .IN2(n6843), .QN(n6841) );
  NOR2X0 U7999 ( .IN1(n6844), .IN2(n4254), .QN(n6843) );
  NOR2X0 U8000 ( .IN1(n6249), .IN2(n4331), .QN(n6842) );
  XOR2X1 U8001 ( .IN1(n6845), .IN2(n6846), .Q(n6249) );
  XOR2X1 U8002 ( .IN1(n3639), .IN2(n4774), .Q(n6846) );
  XOR2X1 U8003 ( .IN1(n6847), .IN2(n4049), .Q(n6845) );
  XOR2X1 U8004 ( .IN1(WX7244), .IN2(n8906), .Q(n6847) );
  NOR2X0 U8005 ( .IN1(n6848), .IN2(n6849), .QN(n6840) );
  NOR2X0 U8006 ( .IN1(DFF_956_n1), .IN2(n4293), .QN(n6849) );
  NOR2X0 U8007 ( .IN1(n4303), .IN2(n5131), .QN(n6848) );
  NAND2X0 U8008 ( .IN1(n4820), .IN2(n8526), .QN(n5131) );
  NAND2X0 U8009 ( .IN1(n6850), .IN2(n6851), .QN(WX5820) );
  NOR2X0 U8010 ( .IN1(n6852), .IN2(n6853), .QN(n6851) );
  NOR2X0 U8011 ( .IN1(n6854), .IN2(n4253), .QN(n6853) );
  NOR2X0 U8012 ( .IN1(n6259), .IN2(n4331), .QN(n6852) );
  XOR2X1 U8013 ( .IN1(n6855), .IN2(n6856), .Q(n6259) );
  XOR2X1 U8014 ( .IN1(n3640), .IN2(n4774), .Q(n6856) );
  XOR2X1 U8015 ( .IN1(n6857), .IN2(n4048), .Q(n6855) );
  XOR2X1 U8016 ( .IN1(WX7242), .IN2(n8907), .Q(n6857) );
  NOR2X0 U8017 ( .IN1(n6858), .IN2(n6859), .QN(n6850) );
  NOR2X0 U8018 ( .IN1(DFF_957_n1), .IN2(n4294), .QN(n6859) );
  NOR2X0 U8019 ( .IN1(n4303), .IN2(n5132), .QN(n6858) );
  NAND2X0 U8020 ( .IN1(n4820), .IN2(n8527), .QN(n5132) );
  NAND2X0 U8021 ( .IN1(n6860), .IN2(n6861), .QN(WX5818) );
  NOR2X0 U8022 ( .IN1(n6862), .IN2(n6863), .QN(n6861) );
  NOR2X0 U8023 ( .IN1(n6864), .IN2(n4254), .QN(n6863) );
  NOR2X0 U8024 ( .IN1(n6269), .IN2(n4331), .QN(n6862) );
  XOR2X1 U8025 ( .IN1(n6865), .IN2(n6866), .Q(n6269) );
  XOR2X1 U8026 ( .IN1(n3641), .IN2(n4774), .Q(n6866) );
  XOR2X1 U8027 ( .IN1(n6867), .IN2(n4047), .Q(n6865) );
  XOR2X1 U8028 ( .IN1(WX7240), .IN2(n8908), .Q(n6867) );
  NOR2X0 U8029 ( .IN1(n6868), .IN2(n6869), .QN(n6860) );
  NOR2X0 U8030 ( .IN1(DFF_958_n1), .IN2(n4294), .QN(n6869) );
  NOR2X0 U8031 ( .IN1(n4303), .IN2(n5133), .QN(n6868) );
  NAND2X0 U8032 ( .IN1(n4820), .IN2(n8528), .QN(n5133) );
  NAND2X0 U8033 ( .IN1(n6870), .IN2(n6871), .QN(WX5816) );
  NOR2X0 U8034 ( .IN1(n6872), .IN2(n6873), .QN(n6871) );
  NOR2X0 U8035 ( .IN1(n6874), .IN2(n4254), .QN(n6873) );
  NOR2X0 U8036 ( .IN1(n6279), .IN2(n4331), .QN(n6872) );
  XOR2X1 U8037 ( .IN1(n6875), .IN2(n6876), .Q(n6279) );
  XOR2X1 U8038 ( .IN1(n3585), .IN2(n4774), .Q(n6876) );
  XOR2X1 U8039 ( .IN1(n6877), .IN2(n4046), .Q(n6875) );
  XOR2X1 U8040 ( .IN1(WX7238), .IN2(n8909), .Q(n6877) );
  NOR2X0 U8041 ( .IN1(n6878), .IN2(n6879), .QN(n6870) );
  NOR2X0 U8042 ( .IN1(n3935), .IN2(n5606), .QN(n6879) );
  NOR2X0 U8043 ( .IN1(DFF_959_n1), .IN2(n4293), .QN(n6878) );
  AND2X1 U8044 ( .IN1(n4800), .IN2(n3935), .Q(WX5718) );
  NOR2X0 U8045 ( .IN1(n4941), .IN2(WX485), .QN(WX546) );
  NOR2X0 U8046 ( .IN1(n4941), .IN2(n6880), .QN(WX5205) );
  XOR2X1 U8047 ( .IN1(n4101), .IN2(DFF_766_n1), .Q(n6880) );
  NOR2X0 U8048 ( .IN1(n4941), .IN2(n6881), .QN(WX5203) );
  XOR2X1 U8049 ( .IN1(n4102), .IN2(DFF_765_n1), .Q(n6881) );
  NOR2X0 U8050 ( .IN1(n4941), .IN2(n6882), .QN(WX5201) );
  XOR2X1 U8051 ( .IN1(n4103), .IN2(DFF_764_n1), .Q(n6882) );
  NOR2X0 U8052 ( .IN1(n4941), .IN2(n6883), .QN(WX5199) );
  XNOR2X1 U8053 ( .IN1(DFF_763_n1), .IN2(test_so40), .Q(n6883) );
  NOR2X0 U8054 ( .IN1(n4941), .IN2(n6884), .QN(WX5197) );
  XOR2X1 U8055 ( .IN1(n4104), .IN2(DFF_762_n1), .Q(n6884) );
  NOR2X0 U8056 ( .IN1(n4941), .IN2(n6885), .QN(WX5195) );
  XOR2X1 U8057 ( .IN1(n4105), .IN2(DFF_761_n1), .Q(n6885) );
  NOR2X0 U8058 ( .IN1(n4941), .IN2(n6886), .QN(WX5193) );
  XOR2X1 U8059 ( .IN1(n4106), .IN2(DFF_760_n1), .Q(n6886) );
  NOR2X0 U8060 ( .IN1(n4941), .IN2(n6887), .QN(WX5191) );
  XOR2X1 U8061 ( .IN1(n4107), .IN2(DFF_759_n1), .Q(n6887) );
  NOR2X0 U8062 ( .IN1(n4942), .IN2(n6888), .QN(WX5189) );
  XNOR2X1 U8063 ( .IN1(n4108), .IN2(test_so43), .Q(n6888) );
  NOR2X0 U8064 ( .IN1(n4942), .IN2(n6889), .QN(WX5187) );
  XOR2X1 U8065 ( .IN1(n4109), .IN2(DFF_757_n1), .Q(n6889) );
  NOR2X0 U8066 ( .IN1(n4942), .IN2(n6890), .QN(WX5185) );
  XOR2X1 U8067 ( .IN1(n4110), .IN2(DFF_756_n1), .Q(n6890) );
  NOR2X0 U8068 ( .IN1(n4942), .IN2(n6891), .QN(WX5183) );
  XOR2X1 U8069 ( .IN1(n4111), .IN2(DFF_755_n1), .Q(n6891) );
  NOR2X0 U8070 ( .IN1(n4942), .IN2(n6892), .QN(WX5181) );
  XOR2X1 U8071 ( .IN1(n4112), .IN2(DFF_754_n1), .Q(n6892) );
  NOR2X0 U8072 ( .IN1(n4942), .IN2(n6893), .QN(WX5179) );
  XOR2X1 U8073 ( .IN1(n4113), .IN2(DFF_753_n1), .Q(n6893) );
  NOR2X0 U8074 ( .IN1(n4942), .IN2(n6894), .QN(WX5177) );
  XOR2X1 U8075 ( .IN1(n4114), .IN2(DFF_752_n1), .Q(n6894) );
  NOR2X0 U8076 ( .IN1(n4942), .IN2(n6895), .QN(WX5175) );
  XNOR2X1 U8077 ( .IN1(DFF_751_n1), .IN2(n6896), .Q(n6895) );
  XOR2X1 U8078 ( .IN1(n3952), .IN2(DFF_767_n1), .Q(n6896) );
  NOR2X0 U8079 ( .IN1(n4942), .IN2(n6897), .QN(WX5173) );
  XOR2X1 U8080 ( .IN1(n4115), .IN2(DFF_750_n1), .Q(n6897) );
  NOR2X0 U8081 ( .IN1(n4942), .IN2(n6898), .QN(WX5171) );
  XOR2X1 U8082 ( .IN1(n4116), .IN2(DFF_749_n1), .Q(n6898) );
  NOR2X0 U8083 ( .IN1(n4942), .IN2(n6899), .QN(WX5169) );
  XOR2X1 U8084 ( .IN1(n4117), .IN2(DFF_748_n1), .Q(n6899) );
  NOR2X0 U8085 ( .IN1(n4942), .IN2(n6900), .QN(WX5167) );
  XOR2X1 U8086 ( .IN1(n4118), .IN2(DFF_747_n1), .Q(n6900) );
  NOR2X0 U8087 ( .IN1(n4942), .IN2(n6901), .QN(WX5165) );
  XOR2X1 U8088 ( .IN1(DFF_746_n1), .IN2(n6902), .Q(n6901) );
  XOR2X1 U8089 ( .IN1(test_so41), .IN2(DFF_767_n1), .Q(n6902) );
  NOR2X0 U8090 ( .IN1(n4943), .IN2(n6903), .QN(WX5163) );
  XOR2X1 U8091 ( .IN1(n4119), .IN2(DFF_745_n1), .Q(n6903) );
  NOR2X0 U8092 ( .IN1(n4943), .IN2(n6904), .QN(WX5161) );
  XOR2X1 U8093 ( .IN1(n4120), .IN2(DFF_744_n1), .Q(n6904) );
  NOR2X0 U8094 ( .IN1(n4943), .IN2(n6905), .QN(WX5159) );
  XOR2X1 U8095 ( .IN1(n4121), .IN2(DFF_743_n1), .Q(n6905) );
  NOR2X0 U8096 ( .IN1(n4943), .IN2(n6906), .QN(WX5157) );
  XOR2X1 U8097 ( .IN1(n4122), .IN2(DFF_742_n1), .Q(n6906) );
  NOR2X0 U8098 ( .IN1(n4943), .IN2(n6907), .QN(WX5155) );
  XNOR2X1 U8099 ( .IN1(n4123), .IN2(test_so42), .Q(n6907) );
  NOR2X0 U8100 ( .IN1(n4943), .IN2(n6908), .QN(WX5153) );
  XOR2X1 U8101 ( .IN1(n4124), .IN2(DFF_740_n1), .Q(n6908) );
  NOR2X0 U8102 ( .IN1(n4943), .IN2(n6909), .QN(WX5151) );
  XNOR2X1 U8103 ( .IN1(DFF_739_n1), .IN2(n6910), .Q(n6909) );
  XOR2X1 U8104 ( .IN1(n3953), .IN2(DFF_767_n1), .Q(n6910) );
  NOR2X0 U8105 ( .IN1(n4943), .IN2(n6911), .QN(WX5149) );
  XOR2X1 U8106 ( .IN1(n4125), .IN2(DFF_738_n1), .Q(n6911) );
  NOR2X0 U8107 ( .IN1(n4943), .IN2(n6912), .QN(WX5147) );
  XOR2X1 U8108 ( .IN1(n4126), .IN2(DFF_737_n1), .Q(n6912) );
  NOR2X0 U8109 ( .IN1(n4943), .IN2(n6913), .QN(WX5145) );
  XOR2X1 U8110 ( .IN1(n4127), .IN2(DFF_736_n1), .Q(n6913) );
  NOR2X0 U8111 ( .IN1(n4943), .IN2(n6914), .QN(WX5143) );
  XOR2X1 U8112 ( .IN1(n3965), .IN2(DFF_767_n1), .Q(n6914) );
  NOR2X0 U8113 ( .IN1(n8961), .IN2(n4922), .QN(WX4617) );
  AND2X1 U8114 ( .IN1(n4800), .IN2(test_so35), .Q(WX4615) );
  NOR2X0 U8115 ( .IN1(n8962), .IN2(n4921), .QN(WX4613) );
  NOR2X0 U8116 ( .IN1(n8963), .IN2(n4857), .QN(WX4611) );
  NOR2X0 U8117 ( .IN1(n8964), .IN2(n4857), .QN(WX4609) );
  NOR2X0 U8118 ( .IN1(n8965), .IN2(n4857), .QN(WX4607) );
  NOR2X0 U8119 ( .IN1(n8966), .IN2(n4857), .QN(WX4605) );
  NOR2X0 U8120 ( .IN1(n8967), .IN2(n4857), .QN(WX4603) );
  NOR2X0 U8121 ( .IN1(n8968), .IN2(n4857), .QN(WX4601) );
  NOR2X0 U8122 ( .IN1(n8969), .IN2(n4857), .QN(WX4599) );
  NOR2X0 U8123 ( .IN1(n8970), .IN2(n4857), .QN(WX4597) );
  NOR2X0 U8124 ( .IN1(n8971), .IN2(n4857), .QN(WX4595) );
  NOR2X0 U8125 ( .IN1(n8972), .IN2(n4857), .QN(WX4593) );
  NOR2X0 U8126 ( .IN1(n8973), .IN2(n4857), .QN(WX4591) );
  NOR2X0 U8127 ( .IN1(n8974), .IN2(n4857), .QN(WX4589) );
  NOR2X0 U8128 ( .IN1(n8977), .IN2(n4856), .QN(WX4587) );
  NAND2X0 U8129 ( .IN1(n6915), .IN2(n6916), .QN(WX4585) );
  NOR2X0 U8130 ( .IN1(n6917), .IN2(n6918), .QN(n6916) );
  NOR2X0 U8131 ( .IN1(n5352), .IN2(n6919), .QN(n6918) );
  NOR2X0 U8132 ( .IN1(n6580), .IN2(n4332), .QN(n6917) );
  XOR2X1 U8133 ( .IN1(n6920), .IN2(n6921), .Q(n6580) );
  XOR2X1 U8134 ( .IN1(n8910), .IN2(n3964), .Q(n6921) );
  XOR2X1 U8135 ( .IN1(WX5879), .IN2(n3814), .Q(n6920) );
  NOR2X0 U8136 ( .IN1(n6922), .IN2(n6923), .QN(n6915) );
  NOR2X0 U8137 ( .IN1(DFF_736_n1), .IN2(n4293), .QN(n6923) );
  NOR2X0 U8138 ( .IN1(n4303), .IN2(n5134), .QN(n6922) );
  NAND2X0 U8139 ( .IN1(n4820), .IN2(n8554), .QN(n5134) );
  NAND2X0 U8140 ( .IN1(n6924), .IN2(n6925), .QN(WX4583) );
  NOR2X0 U8141 ( .IN1(n6926), .IN2(n6927), .QN(n6925) );
  NOR2X0 U8142 ( .IN1(n6928), .IN2(n4254), .QN(n6927) );
  NOR2X0 U8143 ( .IN1(n4339), .IN2(n6589), .QN(n6926) );
  XNOR2X1 U8144 ( .IN1(n6929), .IN2(n6930), .Q(n6589) );
  XOR2X1 U8145 ( .IN1(test_so51), .IN2(n8911), .Q(n6930) );
  XOR2X1 U8146 ( .IN1(WX5877), .IN2(n4100), .Q(n6929) );
  NOR2X0 U8147 ( .IN1(n6931), .IN2(n6932), .QN(n6924) );
  NOR2X0 U8148 ( .IN1(DFF_737_n1), .IN2(n4293), .QN(n6932) );
  NOR2X0 U8149 ( .IN1(n4303), .IN2(n5135), .QN(n6931) );
  NAND2X0 U8150 ( .IN1(n4820), .IN2(n8555), .QN(n5135) );
  NAND2X0 U8151 ( .IN1(n6933), .IN2(n6934), .QN(WX4581) );
  NOR2X0 U8152 ( .IN1(n6935), .IN2(n6936), .QN(n6934) );
  NOR2X0 U8153 ( .IN1(n6937), .IN2(n4254), .QN(n6936) );
  NOR2X0 U8154 ( .IN1(n6598), .IN2(n4332), .QN(n6935) );
  XOR2X1 U8155 ( .IN1(n6938), .IN2(n6939), .Q(n6598) );
  XOR2X1 U8156 ( .IN1(n8912), .IN2(n4099), .Q(n6939) );
  XOR2X1 U8157 ( .IN1(WX5875), .IN2(n3817), .Q(n6938) );
  NOR2X0 U8158 ( .IN1(n6940), .IN2(n6941), .QN(n6933) );
  NOR2X0 U8159 ( .IN1(DFF_738_n1), .IN2(n4293), .QN(n6941) );
  NOR2X0 U8160 ( .IN1(n4303), .IN2(n5136), .QN(n6940) );
  NAND2X0 U8161 ( .IN1(test_so34), .IN2(n4827), .QN(n5136) );
  NAND2X0 U8162 ( .IN1(n6942), .IN2(n6943), .QN(WX4579) );
  NOR2X0 U8163 ( .IN1(n6944), .IN2(n6945), .QN(n6943) );
  NOR2X0 U8164 ( .IN1(n6946), .IN2(n4254), .QN(n6945) );
  NOR2X0 U8165 ( .IN1(n4340), .IN2(n6607), .QN(n6944) );
  XNOR2X1 U8166 ( .IN1(n6947), .IN2(n6948), .Q(n6607) );
  XOR2X1 U8167 ( .IN1(test_so49), .IN2(n8913), .Q(n6948) );
  XOR2X1 U8168 ( .IN1(WX5873), .IN2(n4098), .Q(n6947) );
  NOR2X0 U8169 ( .IN1(n6949), .IN2(n6950), .QN(n6942) );
  NOR2X0 U8170 ( .IN1(DFF_739_n1), .IN2(n4293), .QN(n6950) );
  NOR2X0 U8171 ( .IN1(n4303), .IN2(n5137), .QN(n6949) );
  NAND2X0 U8172 ( .IN1(n4820), .IN2(n8558), .QN(n5137) );
  NAND2X0 U8173 ( .IN1(n6951), .IN2(n6952), .QN(WX4577) );
  NOR2X0 U8174 ( .IN1(n6953), .IN2(n6954), .QN(n6952) );
  NOR2X0 U8175 ( .IN1(n6955), .IN2(n4255), .QN(n6954) );
  NOR2X0 U8176 ( .IN1(n6616), .IN2(n4332), .QN(n6953) );
  XOR2X1 U8177 ( .IN1(n6956), .IN2(n6957), .Q(n6616) );
  XOR2X1 U8178 ( .IN1(n8914), .IN2(n3951), .Q(n6957) );
  XOR2X1 U8179 ( .IN1(WX5871), .IN2(n3820), .Q(n6956) );
  NOR2X0 U8180 ( .IN1(n6958), .IN2(n6959), .QN(n6951) );
  NOR2X0 U8181 ( .IN1(DFF_740_n1), .IN2(n4293), .QN(n6959) );
  NOR2X0 U8182 ( .IN1(n4303), .IN2(n5138), .QN(n6958) );
  NAND2X0 U8183 ( .IN1(n4820), .IN2(n8559), .QN(n5138) );
  NAND2X0 U8184 ( .IN1(n6960), .IN2(n6961), .QN(WX4575) );
  NOR2X0 U8185 ( .IN1(n6962), .IN2(n6963), .QN(n6961) );
  NOR2X0 U8186 ( .IN1(n6964), .IN2(n4254), .QN(n6963) );
  NOR2X0 U8187 ( .IN1(n4340), .IN2(n6625), .QN(n6962) );
  XNOR2X1 U8188 ( .IN1(n6965), .IN2(n6966), .Q(n6625) );
  XOR2X1 U8189 ( .IN1(test_so47), .IN2(n8915), .Q(n6966) );
  XOR2X1 U8190 ( .IN1(WX5997), .IN2(n4097), .Q(n6965) );
  NOR2X0 U8191 ( .IN1(n6967), .IN2(n6968), .QN(n6960) );
  AND2X1 U8192 ( .IN1(n2152), .IN2(test_so42), .Q(n6968) );
  NOR2X0 U8193 ( .IN1(n4303), .IN2(n5140), .QN(n6967) );
  NAND2X0 U8194 ( .IN1(n4820), .IN2(n8560), .QN(n5140) );
  NAND2X0 U8195 ( .IN1(n6969), .IN2(n6970), .QN(WX4573) );
  NOR2X0 U8196 ( .IN1(n6971), .IN2(n6972), .QN(n6970) );
  NOR2X0 U8197 ( .IN1(n6973), .IN2(n4255), .QN(n6972) );
  NOR2X0 U8198 ( .IN1(n6634), .IN2(n4332), .QN(n6971) );
  XOR2X1 U8199 ( .IN1(n6974), .IN2(n6975), .Q(n6634) );
  XOR2X1 U8200 ( .IN1(n8916), .IN2(n4096), .Q(n6975) );
  XOR2X1 U8201 ( .IN1(WX5867), .IN2(n3823), .Q(n6974) );
  NOR2X0 U8202 ( .IN1(n6976), .IN2(n6977), .QN(n6969) );
  NOR2X0 U8203 ( .IN1(DFF_742_n1), .IN2(n4293), .QN(n6977) );
  NOR2X0 U8204 ( .IN1(n4303), .IN2(n5141), .QN(n6976) );
  NAND2X0 U8205 ( .IN1(n4819), .IN2(n8561), .QN(n5141) );
  NAND2X0 U8206 ( .IN1(n6978), .IN2(n6979), .QN(WX4571) );
  NOR2X0 U8207 ( .IN1(n6980), .IN2(n6981), .QN(n6979) );
  NOR2X0 U8208 ( .IN1(n6982), .IN2(n4254), .QN(n6981) );
  NOR2X0 U8209 ( .IN1(n6643), .IN2(n4332), .QN(n6980) );
  XOR2X1 U8210 ( .IN1(n6983), .IN2(n6984), .Q(n6643) );
  XOR2X1 U8211 ( .IN1(n8917), .IN2(n4095), .Q(n6984) );
  XOR2X1 U8212 ( .IN1(WX5865), .IN2(n3825), .Q(n6983) );
  NOR2X0 U8213 ( .IN1(n6985), .IN2(n6986), .QN(n6978) );
  NOR2X0 U8214 ( .IN1(DFF_743_n1), .IN2(n4293), .QN(n6986) );
  NOR2X0 U8215 ( .IN1(n4303), .IN2(n5142), .QN(n6985) );
  NAND2X0 U8216 ( .IN1(n4819), .IN2(n8562), .QN(n5142) );
  NAND2X0 U8217 ( .IN1(n6987), .IN2(n6988), .QN(WX4569) );
  NOR2X0 U8218 ( .IN1(n6989), .IN2(n6990), .QN(n6988) );
  NOR2X0 U8219 ( .IN1(n6991), .IN2(n4254), .QN(n6990) );
  NOR2X0 U8220 ( .IN1(n6652), .IN2(n4335), .QN(n6989) );
  XOR2X1 U8221 ( .IN1(n6992), .IN2(n6993), .Q(n6652) );
  XOR2X1 U8222 ( .IN1(n8918), .IN2(n4094), .Q(n6993) );
  XOR2X1 U8223 ( .IN1(WX5863), .IN2(n3827), .Q(n6992) );
  NOR2X0 U8224 ( .IN1(n6994), .IN2(n6995), .QN(n6987) );
  NOR2X0 U8225 ( .IN1(DFF_744_n1), .IN2(n4293), .QN(n6995) );
  NOR2X0 U8226 ( .IN1(n4303), .IN2(n5143), .QN(n6994) );
  NAND2X0 U8227 ( .IN1(n4819), .IN2(n8563), .QN(n5143) );
  NAND2X0 U8228 ( .IN1(n6996), .IN2(n6997), .QN(WX4567) );
  NOR2X0 U8229 ( .IN1(n6998), .IN2(n6999), .QN(n6997) );
  NOR2X0 U8230 ( .IN1(n7000), .IN2(n4255), .QN(n6999) );
  NOR2X0 U8231 ( .IN1(n6661), .IN2(n4336), .QN(n6998) );
  XOR2X1 U8232 ( .IN1(n7001), .IN2(n7002), .Q(n6661) );
  XOR2X1 U8233 ( .IN1(n8919), .IN2(n4093), .Q(n7002) );
  XOR2X1 U8234 ( .IN1(WX5861), .IN2(n3829), .Q(n7001) );
  NOR2X0 U8235 ( .IN1(n7003), .IN2(n7004), .QN(n6996) );
  NOR2X0 U8236 ( .IN1(DFF_745_n1), .IN2(n4293), .QN(n7004) );
  NOR2X0 U8237 ( .IN1(n4302), .IN2(n5144), .QN(n7003) );
  NAND2X0 U8238 ( .IN1(n4819), .IN2(n8564), .QN(n5144) );
  NAND2X0 U8239 ( .IN1(n7005), .IN2(n7006), .QN(WX4565) );
  NOR2X0 U8240 ( .IN1(n7007), .IN2(n7008), .QN(n7006) );
  NOR2X0 U8241 ( .IN1(n7009), .IN2(n4255), .QN(n7008) );
  NOR2X0 U8242 ( .IN1(n6670), .IN2(n4336), .QN(n7007) );
  XOR2X1 U8243 ( .IN1(n7010), .IN2(n7011), .Q(n6670) );
  XOR2X1 U8244 ( .IN1(n8920), .IN2(n4092), .Q(n7011) );
  XOR2X1 U8245 ( .IN1(WX5859), .IN2(n3831), .Q(n7010) );
  NOR2X0 U8246 ( .IN1(n7012), .IN2(n7013), .QN(n7005) );
  NOR2X0 U8247 ( .IN1(DFF_746_n1), .IN2(n4293), .QN(n7013) );
  NOR2X0 U8248 ( .IN1(n4302), .IN2(n5145), .QN(n7012) );
  NAND2X0 U8249 ( .IN1(n4819), .IN2(n8565), .QN(n5145) );
  NAND2X0 U8250 ( .IN1(n7014), .IN2(n7015), .QN(WX4563) );
  NOR2X0 U8251 ( .IN1(n7016), .IN2(n7017), .QN(n7015) );
  NOR2X0 U8252 ( .IN1(n4260), .IN2(n7018), .QN(n7017) );
  NOR2X0 U8253 ( .IN1(n6679), .IN2(n4337), .QN(n7016) );
  XOR2X1 U8254 ( .IN1(n7019), .IN2(n7020), .Q(n6679) );
  XOR2X1 U8255 ( .IN1(n8921), .IN2(n3950), .Q(n7020) );
  XOR2X1 U8256 ( .IN1(WX5857), .IN2(n3833), .Q(n7019) );
  NOR2X0 U8257 ( .IN1(n7021), .IN2(n7022), .QN(n7014) );
  NOR2X0 U8258 ( .IN1(DFF_747_n1), .IN2(n4293), .QN(n7022) );
  NOR2X0 U8259 ( .IN1(n4302), .IN2(n5146), .QN(n7021) );
  NAND2X0 U8260 ( .IN1(n4819), .IN2(n8566), .QN(n5146) );
  NAND2X0 U8261 ( .IN1(n7023), .IN2(n7024), .QN(WX4561) );
  NOR2X0 U8262 ( .IN1(n7025), .IN2(n7026), .QN(n7024) );
  NOR2X0 U8263 ( .IN1(n7027), .IN2(n4255), .QN(n7026) );
  NOR2X0 U8264 ( .IN1(n6688), .IN2(n4336), .QN(n7025) );
  XOR2X1 U8265 ( .IN1(n7028), .IN2(n7029), .Q(n6688) );
  XOR2X1 U8266 ( .IN1(n8922), .IN2(n4091), .Q(n7029) );
  XOR2X1 U8267 ( .IN1(WX5855), .IN2(n3835), .Q(n7028) );
  NOR2X0 U8268 ( .IN1(n7030), .IN2(n7031), .QN(n7023) );
  NOR2X0 U8269 ( .IN1(DFF_748_n1), .IN2(n4293), .QN(n7031) );
  NOR2X0 U8270 ( .IN1(n4302), .IN2(n5147), .QN(n7030) );
  NAND2X0 U8271 ( .IN1(n4819), .IN2(n8567), .QN(n5147) );
  NAND2X0 U8272 ( .IN1(n7032), .IN2(n7033), .QN(WX4559) );
  NOR2X0 U8273 ( .IN1(n7034), .IN2(n7035), .QN(n7033) );
  NOR2X0 U8274 ( .IN1(n4260), .IN2(n7036), .QN(n7035) );
  NOR2X0 U8275 ( .IN1(n6697), .IN2(n4337), .QN(n7034) );
  XOR2X1 U8276 ( .IN1(n7037), .IN2(n7038), .Q(n6697) );
  XOR2X1 U8277 ( .IN1(n8923), .IN2(n4090), .Q(n7038) );
  XOR2X1 U8278 ( .IN1(WX5853), .IN2(n3837), .Q(n7037) );
  NOR2X0 U8279 ( .IN1(n7039), .IN2(n7040), .QN(n7032) );
  NOR2X0 U8280 ( .IN1(DFF_749_n1), .IN2(n4292), .QN(n7040) );
  NOR2X0 U8281 ( .IN1(n4302), .IN2(n5148), .QN(n7039) );
  NAND2X0 U8282 ( .IN1(n4819), .IN2(n8568), .QN(n5148) );
  NAND2X0 U8283 ( .IN1(n7041), .IN2(n7042), .QN(WX4557) );
  NOR2X0 U8284 ( .IN1(n7043), .IN2(n7044), .QN(n7042) );
  NOR2X0 U8285 ( .IN1(n7045), .IN2(n4256), .QN(n7044) );
  NOR2X0 U8286 ( .IN1(n6706), .IN2(n4336), .QN(n7043) );
  XOR2X1 U8287 ( .IN1(n7046), .IN2(n7047), .Q(n6706) );
  XOR2X1 U8288 ( .IN1(n8924), .IN2(n4089), .Q(n7047) );
  XOR2X1 U8289 ( .IN1(WX5851), .IN2(n3839), .Q(n7046) );
  NOR2X0 U8290 ( .IN1(n7048), .IN2(n7049), .QN(n7041) );
  NOR2X0 U8291 ( .IN1(DFF_750_n1), .IN2(n4292), .QN(n7049) );
  NOR2X0 U8292 ( .IN1(n4302), .IN2(n5149), .QN(n7048) );
  NAND2X0 U8293 ( .IN1(n4818), .IN2(n8569), .QN(n5149) );
  NAND2X0 U8294 ( .IN1(n7050), .IN2(n7051), .QN(WX4555) );
  NOR2X0 U8295 ( .IN1(n7052), .IN2(n7053), .QN(n7051) );
  NOR2X0 U8296 ( .IN1(n4260), .IN2(n7054), .QN(n7053) );
  NOR2X0 U8297 ( .IN1(n6715), .IN2(n4337), .QN(n7052) );
  XOR2X1 U8298 ( .IN1(n7055), .IN2(n7056), .Q(n6715) );
  XOR2X1 U8299 ( .IN1(n8925), .IN2(n4088), .Q(n7056) );
  XOR2X1 U8300 ( .IN1(WX5849), .IN2(n3841), .Q(n7055) );
  NOR2X0 U8301 ( .IN1(n7057), .IN2(n7058), .QN(n7050) );
  NOR2X0 U8302 ( .IN1(DFF_751_n1), .IN2(n4292), .QN(n7058) );
  NOR2X0 U8303 ( .IN1(n4302), .IN2(n5151), .QN(n7057) );
  NAND2X0 U8304 ( .IN1(n4818), .IN2(n8570), .QN(n5151) );
  NAND2X0 U8305 ( .IN1(n7059), .IN2(n7060), .QN(WX4553) );
  NOR2X0 U8306 ( .IN1(n7061), .IN2(n7062), .QN(n7060) );
  NOR2X0 U8307 ( .IN1(n7063), .IN2(n4256), .QN(n7062) );
  NOR2X0 U8308 ( .IN1(n4339), .IN2(n6724), .QN(n7061) );
  XNOR2X1 U8309 ( .IN1(n7064), .IN2(n7065), .Q(n6724) );
  XOR2X1 U8310 ( .IN1(n3642), .IN2(n4775), .Q(n7065) );
  XOR2X1 U8311 ( .IN1(WX5911), .IN2(n7066), .Q(n7064) );
  XOR2X1 U8312 ( .IN1(test_so52), .IN2(n8926), .Q(n7066) );
  NOR2X0 U8313 ( .IN1(n7067), .IN2(n7068), .QN(n7059) );
  NOR2X0 U8314 ( .IN1(DFF_752_n1), .IN2(n4292), .QN(n7068) );
  NOR2X0 U8315 ( .IN1(n4302), .IN2(n5152), .QN(n7067) );
  NAND2X0 U8316 ( .IN1(n4818), .IN2(n8571), .QN(n5152) );
  NAND2X0 U8317 ( .IN1(n7069), .IN2(n7070), .QN(WX4551) );
  NOR2X0 U8318 ( .IN1(n7071), .IN2(n7072), .QN(n7070) );
  NOR2X0 U8319 ( .IN1(n4260), .IN2(n7073), .QN(n7072) );
  NOR2X0 U8320 ( .IN1(n6734), .IN2(n4336), .QN(n7071) );
  XOR2X1 U8321 ( .IN1(n7074), .IN2(n7075), .Q(n6734) );
  XOR2X1 U8322 ( .IN1(n3643), .IN2(n4775), .Q(n7075) );
  XOR2X1 U8323 ( .IN1(n7076), .IN2(n4087), .Q(n7074) );
  XOR2X1 U8324 ( .IN1(WX5973), .IN2(n8927), .Q(n7076) );
  NOR2X0 U8325 ( .IN1(n7077), .IN2(n7078), .QN(n7069) );
  NOR2X0 U8326 ( .IN1(DFF_753_n1), .IN2(n4292), .QN(n7078) );
  NOR2X0 U8327 ( .IN1(n4302), .IN2(n5153), .QN(n7077) );
  NAND2X0 U8328 ( .IN1(n4818), .IN2(n8572), .QN(n5153) );
  NAND2X0 U8329 ( .IN1(n7079), .IN2(n7080), .QN(WX4549) );
  NOR2X0 U8330 ( .IN1(n7081), .IN2(n7082), .QN(n7080) );
  NOR2X0 U8331 ( .IN1(n7083), .IN2(n4256), .QN(n7082) );
  NOR2X0 U8332 ( .IN1(n4339), .IN2(n6744), .QN(n7081) );
  XNOR2X1 U8333 ( .IN1(n7084), .IN2(n7085), .Q(n6744) );
  XOR2X1 U8334 ( .IN1(n4086), .IN2(n4775), .Q(n7085) );
  XOR2X1 U8335 ( .IN1(n7086), .IN2(n8930), .Q(n7084) );
  XOR2X1 U8336 ( .IN1(n8929), .IN2(n8928), .Q(n7086) );
  NOR2X0 U8337 ( .IN1(n7087), .IN2(n7088), .QN(n7079) );
  NOR2X0 U8338 ( .IN1(DFF_754_n1), .IN2(n4292), .QN(n7088) );
  NOR2X0 U8339 ( .IN1(n4302), .IN2(n5154), .QN(n7087) );
  NAND2X0 U8340 ( .IN1(n4818), .IN2(n8573), .QN(n5154) );
  NAND2X0 U8341 ( .IN1(n7089), .IN2(n7090), .QN(WX4547) );
  NOR2X0 U8342 ( .IN1(n7091), .IN2(n7092), .QN(n7090) );
  NOR2X0 U8343 ( .IN1(n7093), .IN2(n4255), .QN(n7092) );
  NOR2X0 U8344 ( .IN1(n6754), .IN2(n4336), .QN(n7091) );
  XOR2X1 U8345 ( .IN1(n7094), .IN2(n7095), .Q(n6754) );
  XOR2X1 U8346 ( .IN1(n3644), .IN2(n4775), .Q(n7095) );
  XOR2X1 U8347 ( .IN1(n7096), .IN2(n4085), .Q(n7094) );
  XOR2X1 U8348 ( .IN1(WX5969), .IN2(n8931), .Q(n7096) );
  NOR2X0 U8349 ( .IN1(n7097), .IN2(n7098), .QN(n7089) );
  NOR2X0 U8350 ( .IN1(DFF_755_n1), .IN2(n4292), .QN(n7098) );
  NOR2X0 U8351 ( .IN1(n4302), .IN2(n5155), .QN(n7097) );
  NAND2X0 U8352 ( .IN1(test_so33), .IN2(n4799), .QN(n5155) );
  NAND2X0 U8353 ( .IN1(n7099), .IN2(n7100), .QN(WX4545) );
  NOR2X0 U8354 ( .IN1(n7101), .IN2(n7102), .QN(n7100) );
  NOR2X0 U8355 ( .IN1(n7103), .IN2(n4256), .QN(n7102) );
  NOR2X0 U8356 ( .IN1(n4338), .IN2(n6764), .QN(n7101) );
  XNOR2X1 U8357 ( .IN1(n7104), .IN2(n7105), .Q(n6764) );
  XOR2X1 U8358 ( .IN1(n4084), .IN2(n4775), .Q(n7105) );
  XOR2X1 U8359 ( .IN1(n7106), .IN2(n8934), .Q(n7104) );
  XOR2X1 U8360 ( .IN1(n8933), .IN2(n8932), .Q(n7106) );
  NOR2X0 U8361 ( .IN1(n7107), .IN2(n7108), .QN(n7099) );
  NOR2X0 U8362 ( .IN1(DFF_756_n1), .IN2(n4292), .QN(n7108) );
  NOR2X0 U8363 ( .IN1(n4302), .IN2(n5156), .QN(n7107) );
  NAND2X0 U8364 ( .IN1(n4818), .IN2(n8576), .QN(n5156) );
  NAND2X0 U8365 ( .IN1(n7109), .IN2(n7110), .QN(WX4543) );
  NOR2X0 U8366 ( .IN1(n7111), .IN2(n7112), .QN(n7110) );
  NOR2X0 U8367 ( .IN1(n7113), .IN2(n4256), .QN(n7112) );
  NOR2X0 U8368 ( .IN1(n6774), .IN2(n4336), .QN(n7111) );
  XOR2X1 U8369 ( .IN1(n7114), .IN2(n7115), .Q(n6774) );
  XOR2X1 U8370 ( .IN1(n3645), .IN2(n4775), .Q(n7115) );
  XOR2X1 U8371 ( .IN1(n7116), .IN2(n4083), .Q(n7114) );
  XOR2X1 U8372 ( .IN1(WX5965), .IN2(n8935), .Q(n7116) );
  NOR2X0 U8373 ( .IN1(n7117), .IN2(n7118), .QN(n7109) );
  NOR2X0 U8374 ( .IN1(DFF_757_n1), .IN2(n4292), .QN(n7118) );
  NOR2X0 U8375 ( .IN1(n4301), .IN2(n5157), .QN(n7117) );
  NAND2X0 U8376 ( .IN1(n4818), .IN2(n8577), .QN(n5157) );
  NAND2X0 U8377 ( .IN1(n7119), .IN2(n7120), .QN(WX4541) );
  NOR2X0 U8378 ( .IN1(n7121), .IN2(n7122), .QN(n7120) );
  NOR2X0 U8379 ( .IN1(n7123), .IN2(n4256), .QN(n7122) );
  NOR2X0 U8380 ( .IN1(n4338), .IN2(n6784), .QN(n7121) );
  XNOR2X1 U8381 ( .IN1(n7124), .IN2(n7125), .Q(n6784) );
  XOR2X1 U8382 ( .IN1(n3646), .IN2(n4775), .Q(n7125) );
  XOR2X1 U8383 ( .IN1(n7126), .IN2(n4082), .Q(n7124) );
  XOR2X1 U8384 ( .IN1(WX5899), .IN2(test_so46), .Q(n7126) );
  NOR2X0 U8385 ( .IN1(n7127), .IN2(n7128), .QN(n7119) );
  AND2X1 U8386 ( .IN1(n2152), .IN2(test_so43), .Q(n7128) );
  NOR2X0 U8387 ( .IN1(n4301), .IN2(n5158), .QN(n7127) );
  NAND2X0 U8388 ( .IN1(n4818), .IN2(n8578), .QN(n5158) );
  NAND2X0 U8389 ( .IN1(n7129), .IN2(n7130), .QN(WX4539) );
  NOR2X0 U8390 ( .IN1(n7131), .IN2(n7132), .QN(n7130) );
  NOR2X0 U8391 ( .IN1(n7133), .IN2(n4255), .QN(n7132) );
  NOR2X0 U8392 ( .IN1(n6794), .IN2(n4336), .QN(n7131) );
  XOR2X1 U8393 ( .IN1(n7134), .IN2(n7135), .Q(n6794) );
  XOR2X1 U8394 ( .IN1(n3647), .IN2(n4775), .Q(n7135) );
  XOR2X1 U8395 ( .IN1(n7136), .IN2(n4081), .Q(n7134) );
  XOR2X1 U8396 ( .IN1(WX5961), .IN2(n8936), .Q(n7136) );
  NOR2X0 U8397 ( .IN1(n7137), .IN2(n7138), .QN(n7129) );
  NOR2X0 U8398 ( .IN1(DFF_759_n1), .IN2(n4292), .QN(n7138) );
  NOR2X0 U8399 ( .IN1(n4301), .IN2(n5159), .QN(n7137) );
  NAND2X0 U8400 ( .IN1(n4818), .IN2(n8579), .QN(n5159) );
  NAND2X0 U8401 ( .IN1(n7139), .IN2(n7140), .QN(WX4537) );
  NOR2X0 U8402 ( .IN1(n7141), .IN2(n7142), .QN(n7140) );
  NOR2X0 U8403 ( .IN1(n7143), .IN2(n4257), .QN(n7142) );
  NOR2X0 U8404 ( .IN1(n6804), .IN2(n4335), .QN(n7141) );
  XOR2X1 U8405 ( .IN1(n7144), .IN2(n7145), .Q(n6804) );
  XOR2X1 U8406 ( .IN1(n3648), .IN2(n4775), .Q(n7145) );
  XOR2X1 U8407 ( .IN1(n7146), .IN2(n4080), .Q(n7144) );
  XOR2X1 U8408 ( .IN1(WX5959), .IN2(n8937), .Q(n7146) );
  NOR2X0 U8409 ( .IN1(n7147), .IN2(n7148), .QN(n7139) );
  NOR2X0 U8410 ( .IN1(DFF_760_n1), .IN2(n4292), .QN(n7148) );
  NOR2X0 U8411 ( .IN1(n4301), .IN2(n5160), .QN(n7147) );
  NAND2X0 U8412 ( .IN1(n4817), .IN2(n8580), .QN(n5160) );
  NAND2X0 U8413 ( .IN1(n7149), .IN2(n7150), .QN(WX4535) );
  NOR2X0 U8414 ( .IN1(n7151), .IN2(n7152), .QN(n7150) );
  NOR2X0 U8415 ( .IN1(n7153), .IN2(n4255), .QN(n7152) );
  NOR2X0 U8416 ( .IN1(n6814), .IN2(n4337), .QN(n7151) );
  XOR2X1 U8417 ( .IN1(n7154), .IN2(n7155), .Q(n6814) );
  XOR2X1 U8418 ( .IN1(n3649), .IN2(n4775), .Q(n7155) );
  XOR2X1 U8419 ( .IN1(n7156), .IN2(n4079), .Q(n7154) );
  XOR2X1 U8420 ( .IN1(WX5957), .IN2(n8938), .Q(n7156) );
  NOR2X0 U8421 ( .IN1(n7157), .IN2(n7158), .QN(n7149) );
  NOR2X0 U8422 ( .IN1(DFF_761_n1), .IN2(n4292), .QN(n7158) );
  NOR2X0 U8423 ( .IN1(n4301), .IN2(n5162), .QN(n7157) );
  NAND2X0 U8424 ( .IN1(n4817), .IN2(n8581), .QN(n5162) );
  NAND2X0 U8425 ( .IN1(n7159), .IN2(n7160), .QN(WX4533) );
  NOR2X0 U8426 ( .IN1(n7161), .IN2(n7162), .QN(n7160) );
  NOR2X0 U8427 ( .IN1(n7163), .IN2(n4257), .QN(n7162) );
  NOR2X0 U8428 ( .IN1(n6824), .IN2(n4336), .QN(n7161) );
  XOR2X1 U8429 ( .IN1(n7164), .IN2(n7165), .Q(n6824) );
  XOR2X1 U8430 ( .IN1(n3650), .IN2(n4775), .Q(n7165) );
  XOR2X1 U8431 ( .IN1(n7166), .IN2(n4078), .Q(n7164) );
  XOR2X1 U8432 ( .IN1(WX5955), .IN2(n8939), .Q(n7166) );
  NOR2X0 U8433 ( .IN1(n7167), .IN2(n7168), .QN(n7159) );
  NOR2X0 U8434 ( .IN1(DFF_762_n1), .IN2(n4292), .QN(n7168) );
  NOR2X0 U8435 ( .IN1(n4301), .IN2(n5163), .QN(n7167) );
  NAND2X0 U8436 ( .IN1(n4817), .IN2(n8582), .QN(n5163) );
  NAND2X0 U8437 ( .IN1(n7169), .IN2(n7170), .QN(WX4531) );
  NOR2X0 U8438 ( .IN1(n7171), .IN2(n7172), .QN(n7170) );
  NOR2X0 U8439 ( .IN1(n7173), .IN2(n4257), .QN(n7172) );
  NOR2X0 U8440 ( .IN1(n6834), .IN2(n4336), .QN(n7171) );
  XOR2X1 U8441 ( .IN1(n7174), .IN2(n7175), .Q(n6834) );
  XOR2X1 U8442 ( .IN1(n3651), .IN2(n4775), .Q(n7175) );
  XOR2X1 U8443 ( .IN1(n7176), .IN2(n4077), .Q(n7174) );
  XOR2X1 U8444 ( .IN1(WX5953), .IN2(n8940), .Q(n7176) );
  NOR2X0 U8445 ( .IN1(n7177), .IN2(n7178), .QN(n7169) );
  NOR2X0 U8446 ( .IN1(DFF_763_n1), .IN2(n4292), .QN(n7178) );
  NOR2X0 U8447 ( .IN1(n4301), .IN2(n5164), .QN(n7177) );
  NAND2X0 U8448 ( .IN1(n4817), .IN2(n8583), .QN(n5164) );
  NAND2X0 U8449 ( .IN1(n7179), .IN2(n7180), .QN(WX4529) );
  NOR2X0 U8450 ( .IN1(n7181), .IN2(n7182), .QN(n7180) );
  NOR2X0 U8451 ( .IN1(n4259), .IN2(n7183), .QN(n7182) );
  NOR2X0 U8452 ( .IN1(n6844), .IN2(n4335), .QN(n7181) );
  XOR2X1 U8453 ( .IN1(n7184), .IN2(n7185), .Q(n6844) );
  XOR2X1 U8454 ( .IN1(n3652), .IN2(n4776), .Q(n7185) );
  XOR2X1 U8455 ( .IN1(n7186), .IN2(n4076), .Q(n7184) );
  XOR2X1 U8456 ( .IN1(WX5951), .IN2(n8941), .Q(n7186) );
  NOR2X0 U8457 ( .IN1(n7187), .IN2(n7188), .QN(n7179) );
  NOR2X0 U8458 ( .IN1(DFF_764_n1), .IN2(n4291), .QN(n7188) );
  NOR2X0 U8459 ( .IN1(n4301), .IN2(n5165), .QN(n7187) );
  NAND2X0 U8460 ( .IN1(n4817), .IN2(n8584), .QN(n5165) );
  NAND2X0 U8461 ( .IN1(n7189), .IN2(n7190), .QN(WX4527) );
  NOR2X0 U8462 ( .IN1(n7191), .IN2(n7192), .QN(n7190) );
  NOR2X0 U8463 ( .IN1(n7193), .IN2(n4257), .QN(n7192) );
  NOR2X0 U8464 ( .IN1(n6854), .IN2(n4336), .QN(n7191) );
  XOR2X1 U8465 ( .IN1(n7194), .IN2(n7195), .Q(n6854) );
  XOR2X1 U8466 ( .IN1(n3653), .IN2(n4776), .Q(n7195) );
  XOR2X1 U8467 ( .IN1(n7196), .IN2(n4075), .Q(n7194) );
  XOR2X1 U8468 ( .IN1(WX5949), .IN2(n8942), .Q(n7196) );
  NOR2X0 U8469 ( .IN1(n7197), .IN2(n7198), .QN(n7189) );
  NOR2X0 U8470 ( .IN1(DFF_765_n1), .IN2(n4291), .QN(n7198) );
  NOR2X0 U8471 ( .IN1(n4301), .IN2(n5166), .QN(n7197) );
  NAND2X0 U8472 ( .IN1(n4817), .IN2(n8585), .QN(n5166) );
  NAND2X0 U8473 ( .IN1(n7199), .IN2(n7200), .QN(WX4525) );
  NOR2X0 U8474 ( .IN1(n7201), .IN2(n7202), .QN(n7200) );
  NOR2X0 U8475 ( .IN1(n4259), .IN2(n7203), .QN(n7202) );
  NOR2X0 U8476 ( .IN1(n6864), .IN2(n4336), .QN(n7201) );
  XOR2X1 U8477 ( .IN1(n7204), .IN2(n7205), .Q(n6864) );
  XOR2X1 U8478 ( .IN1(n3654), .IN2(n4776), .Q(n7205) );
  XOR2X1 U8479 ( .IN1(n7206), .IN2(n4074), .Q(n7204) );
  XOR2X1 U8480 ( .IN1(WX5947), .IN2(n8943), .Q(n7206) );
  NOR2X0 U8481 ( .IN1(n7207), .IN2(n7208), .QN(n7199) );
  NOR2X0 U8482 ( .IN1(DFF_766_n1), .IN2(n4291), .QN(n7208) );
  NOR2X0 U8483 ( .IN1(n4301), .IN2(n5167), .QN(n7207) );
  NAND2X0 U8484 ( .IN1(n4817), .IN2(n8586), .QN(n5167) );
  NAND2X0 U8485 ( .IN1(n7209), .IN2(n7210), .QN(WX4523) );
  NOR2X0 U8486 ( .IN1(n7211), .IN2(n7212), .QN(n7210) );
  NOR2X0 U8487 ( .IN1(n7213), .IN2(n4256), .QN(n7212) );
  NOR2X0 U8488 ( .IN1(n6874), .IN2(n4336), .QN(n7211) );
  XOR2X1 U8489 ( .IN1(n7214), .IN2(n7215), .Q(n6874) );
  XOR2X1 U8490 ( .IN1(n3586), .IN2(n4776), .Q(n7215) );
  XOR2X1 U8491 ( .IN1(n7216), .IN2(n4073), .Q(n7214) );
  XOR2X1 U8492 ( .IN1(WX5945), .IN2(n8944), .Q(n7216) );
  NOR2X0 U8493 ( .IN1(n7217), .IN2(n7218), .QN(n7209) );
  NOR2X0 U8494 ( .IN1(n3936), .IN2(n5606), .QN(n7218) );
  NOR2X0 U8495 ( .IN1(DFF_767_n1), .IN2(n4291), .QN(n7217) );
  AND2X1 U8496 ( .IN1(n4801), .IN2(n3936), .Q(WX4425) );
  NOR2X0 U8497 ( .IN1(n4943), .IN2(n7219), .QN(WX3912) );
  XOR2X1 U8498 ( .IN1(n4128), .IN2(DFF_574_n1), .Q(n7219) );
  NOR2X0 U8499 ( .IN1(n4943), .IN2(n7220), .QN(WX3910) );
  XOR2X1 U8500 ( .IN1(n4129), .IN2(DFF_573_n1), .Q(n7220) );
  NOR2X0 U8501 ( .IN1(n4944), .IN2(n7221), .QN(WX3908) );
  XOR2X1 U8502 ( .IN1(n4130), .IN2(DFF_572_n1), .Q(n7221) );
  NOR2X0 U8503 ( .IN1(n4944), .IN2(n7222), .QN(WX3906) );
  XNOR2X1 U8504 ( .IN1(n4131), .IN2(test_so32), .Q(n7222) );
  NOR2X0 U8505 ( .IN1(n4944), .IN2(n7223), .QN(WX3904) );
  XOR2X1 U8506 ( .IN1(n4132), .IN2(DFF_570_n1), .Q(n7223) );
  NOR2X0 U8507 ( .IN1(n4944), .IN2(n7224), .QN(WX3902) );
  XOR2X1 U8508 ( .IN1(n4133), .IN2(DFF_569_n1), .Q(n7224) );
  NOR2X0 U8509 ( .IN1(n4944), .IN2(n7225), .QN(WX3900) );
  XOR2X1 U8510 ( .IN1(n4134), .IN2(DFF_568_n1), .Q(n7225) );
  NOR2X0 U8511 ( .IN1(n4944), .IN2(n7226), .QN(WX3898) );
  XOR2X1 U8512 ( .IN1(n4135), .IN2(DFF_567_n1), .Q(n7226) );
  NOR2X0 U8513 ( .IN1(n4944), .IN2(n7227), .QN(WX3896) );
  XNOR2X1 U8514 ( .IN1(DFF_566_n1), .IN2(test_so29), .Q(n7227) );
  NOR2X0 U8515 ( .IN1(n4944), .IN2(n7228), .QN(WX3894) );
  XOR2X1 U8516 ( .IN1(n4136), .IN2(DFF_565_n1), .Q(n7228) );
  NOR2X0 U8517 ( .IN1(n4944), .IN2(n7229), .QN(WX3892) );
  XOR2X1 U8518 ( .IN1(n4137), .IN2(DFF_564_n1), .Q(n7229) );
  NOR2X0 U8519 ( .IN1(n4944), .IN2(n7230), .QN(WX3890) );
  XOR2X1 U8520 ( .IN1(n4138), .IN2(DFF_563_n1), .Q(n7230) );
  NOR2X0 U8521 ( .IN1(n4944), .IN2(n7231), .QN(WX3888) );
  XOR2X1 U8522 ( .IN1(n4139), .IN2(DFF_562_n1), .Q(n7231) );
  NOR2X0 U8523 ( .IN1(n4944), .IN2(n7232), .QN(WX3886) );
  XOR2X1 U8524 ( .IN1(n4140), .IN2(DFF_561_n1), .Q(n7232) );
  NOR2X0 U8525 ( .IN1(n4944), .IN2(n7233), .QN(WX3884) );
  XOR2X1 U8526 ( .IN1(n4141), .IN2(DFF_560_n1), .Q(n7233) );
  NOR2X0 U8527 ( .IN1(n4945), .IN2(n7234), .QN(WX3882) );
  XNOR2X1 U8528 ( .IN1(DFF_559_n1), .IN2(n7235), .Q(n7234) );
  XOR2X1 U8529 ( .IN1(n3954), .IN2(DFF_575_n1), .Q(n7235) );
  NOR2X0 U8530 ( .IN1(n4945), .IN2(n7236), .QN(WX3880) );
  XOR2X1 U8531 ( .IN1(n4142), .IN2(DFF_558_n1), .Q(n7236) );
  NOR2X0 U8532 ( .IN1(n4945), .IN2(n7237), .QN(WX3878) );
  XOR2X1 U8533 ( .IN1(n4143), .IN2(DFF_557_n1), .Q(n7237) );
  NOR2X0 U8534 ( .IN1(n4945), .IN2(n7238), .QN(WX3876) );
  XOR2X1 U8535 ( .IN1(n4144), .IN2(DFF_556_n1), .Q(n7238) );
  NOR2X0 U8536 ( .IN1(n4945), .IN2(n7239), .QN(WX3874) );
  XOR2X1 U8537 ( .IN1(n4145), .IN2(DFF_555_n1), .Q(n7239) );
  NOR2X0 U8538 ( .IN1(n4945), .IN2(n7240), .QN(WX3872) );
  XOR2X1 U8539 ( .IN1(DFF_575_n1), .IN2(n7241), .Q(n7240) );
  XOR2X1 U8540 ( .IN1(test_so31), .IN2(n3955), .Q(n7241) );
  NOR2X0 U8541 ( .IN1(n4945), .IN2(n7242), .QN(WX3870) );
  XOR2X1 U8542 ( .IN1(n4146), .IN2(DFF_553_n1), .Q(n7242) );
  NOR2X0 U8543 ( .IN1(n4945), .IN2(n7243), .QN(WX3868) );
  XOR2X1 U8544 ( .IN1(n4147), .IN2(DFF_552_n1), .Q(n7243) );
  NOR2X0 U8545 ( .IN1(n4945), .IN2(n7244), .QN(WX3866) );
  XOR2X1 U8546 ( .IN1(n4148), .IN2(DFF_551_n1), .Q(n7244) );
  NOR2X0 U8547 ( .IN1(n4945), .IN2(n7245), .QN(WX3864) );
  XOR2X1 U8548 ( .IN1(n4149), .IN2(DFF_550_n1), .Q(n7245) );
  NOR2X0 U8549 ( .IN1(n4945), .IN2(n7246), .QN(WX3862) );
  XNOR2X1 U8550 ( .IN1(DFF_549_n1), .IN2(test_so30), .Q(n7246) );
  NOR2X0 U8551 ( .IN1(n4945), .IN2(n7247), .QN(WX3860) );
  XOR2X1 U8552 ( .IN1(n4150), .IN2(DFF_548_n1), .Q(n7247) );
  NOR2X0 U8553 ( .IN1(n4945), .IN2(n7248), .QN(WX3858) );
  XNOR2X1 U8554 ( .IN1(DFF_547_n1), .IN2(n7249), .Q(n7248) );
  XOR2X1 U8555 ( .IN1(n3956), .IN2(DFF_575_n1), .Q(n7249) );
  NOR2X0 U8556 ( .IN1(n4860), .IN2(n7250), .QN(WX3856) );
  XOR2X1 U8557 ( .IN1(n4151), .IN2(DFF_546_n1), .Q(n7250) );
  NOR2X0 U8558 ( .IN1(n4859), .IN2(n7251), .QN(WX3854) );
  XOR2X1 U8559 ( .IN1(n4152), .IN2(DFF_545_n1), .Q(n7251) );
  NOR2X0 U8560 ( .IN1(n4868), .IN2(n7252), .QN(WX3852) );
  XOR2X1 U8561 ( .IN1(n4153), .IN2(DFF_544_n1), .Q(n7252) );
  NOR2X0 U8562 ( .IN1(n4867), .IN2(n7253), .QN(WX3850) );
  XOR2X1 U8563 ( .IN1(n3966), .IN2(DFF_575_n1), .Q(n7253) );
  AND2X1 U8564 ( .IN1(n4801), .IN2(test_so24), .Q(WX3324) );
  NOR2X0 U8565 ( .IN1(n9012), .IN2(n4856), .QN(WX3322) );
  NOR2X0 U8566 ( .IN1(n9016), .IN2(n4856), .QN(WX3320) );
  NOR2X0 U8567 ( .IN1(n9018), .IN2(n4856), .QN(WX3318) );
  NOR2X0 U8568 ( .IN1(n9020), .IN2(n4856), .QN(WX3316) );
  NOR2X0 U8569 ( .IN1(n9022), .IN2(n4856), .QN(WX3314) );
  NOR2X0 U8570 ( .IN1(n9023), .IN2(n4856), .QN(WX3312) );
  NOR2X0 U8571 ( .IN1(n9025), .IN2(n4856), .QN(WX3310) );
  NOR2X0 U8572 ( .IN1(n9027), .IN2(n4856), .QN(WX3308) );
  NOR2X0 U8573 ( .IN1(n9029), .IN2(n4856), .QN(WX3306) );
  NOR2X0 U8574 ( .IN1(n9031), .IN2(n4856), .QN(WX3304) );
  NOR2X0 U8575 ( .IN1(n9035), .IN2(n4856), .QN(WX3302) );
  NOR2X0 U8576 ( .IN1(n9037), .IN2(n4855), .QN(WX3300) );
  NOR2X0 U8577 ( .IN1(n9039), .IN2(n4855), .QN(WX3298) );
  NOR2X0 U8578 ( .IN1(n9041), .IN2(n4855), .QN(WX3296) );
  NOR2X0 U8579 ( .IN1(n9044), .IN2(n4855), .QN(WX3294) );
  NAND2X0 U8580 ( .IN1(n7254), .IN2(n7255), .QN(WX3292) );
  NOR2X0 U8581 ( .IN1(n7256), .IN2(n7257), .QN(n7255) );
  NOR2X0 U8582 ( .IN1(n7258), .IN2(n4257), .QN(n7257) );
  NOR2X0 U8583 ( .IN1(n4337), .IN2(n6919), .QN(n7256) );
  XNOR2X1 U8584 ( .IN1(n7259), .IN2(n7260), .Q(n6919) );
  XOR2X1 U8585 ( .IN1(test_so36), .IN2(n8945), .Q(n7260) );
  XOR2X1 U8586 ( .IN1(WX4714), .IN2(n3965), .Q(n7259) );
  NOR2X0 U8587 ( .IN1(n7261), .IN2(n7262), .QN(n7254) );
  NOR2X0 U8588 ( .IN1(DFF_544_n1), .IN2(n4291), .QN(n7262) );
  NOR2X0 U8589 ( .IN1(n4301), .IN2(n5168), .QN(n7261) );
  NAND2X0 U8590 ( .IN1(n4817), .IN2(n8612), .QN(n5168) );
  NAND2X0 U8591 ( .IN1(n7263), .IN2(n7264), .QN(WX3290) );
  NOR2X0 U8592 ( .IN1(n7265), .IN2(n7266), .QN(n7264) );
  NOR2X0 U8593 ( .IN1(n7267), .IN2(n4257), .QN(n7266) );
  NOR2X0 U8594 ( .IN1(n6928), .IN2(n4336), .QN(n7265) );
  XOR2X1 U8595 ( .IN1(n7268), .IN2(n7269), .Q(n6928) );
  XOR2X1 U8596 ( .IN1(n8946), .IN2(n4127), .Q(n7269) );
  XOR2X1 U8597 ( .IN1(WX4584), .IN2(n3844), .Q(n7268) );
  NOR2X0 U8598 ( .IN1(n7270), .IN2(n7271), .QN(n7263) );
  NOR2X0 U8599 ( .IN1(DFF_545_n1), .IN2(n4291), .QN(n7271) );
  NOR2X0 U8600 ( .IN1(n4301), .IN2(n5169), .QN(n7270) );
  NAND2X0 U8601 ( .IN1(n4817), .IN2(n8613), .QN(n5169) );
  NAND2X0 U8602 ( .IN1(n7272), .IN2(n7273), .QN(WX3288) );
  NOR2X0 U8603 ( .IN1(n7274), .IN2(n7275), .QN(n7273) );
  NOR2X0 U8604 ( .IN1(n7276), .IN2(n4255), .QN(n7275) );
  NOR2X0 U8605 ( .IN1(n6937), .IN2(n4335), .QN(n7274) );
  XOR2X1 U8606 ( .IN1(n7277), .IN2(n7278), .Q(n6937) );
  XOR2X1 U8607 ( .IN1(n8947), .IN2(n4126), .Q(n7278) );
  XOR2X1 U8608 ( .IN1(WX4582), .IN2(n3846), .Q(n7277) );
  NOR2X0 U8609 ( .IN1(n7279), .IN2(n7280), .QN(n7272) );
  NOR2X0 U8610 ( .IN1(DFF_546_n1), .IN2(n4291), .QN(n7280) );
  NOR2X0 U8611 ( .IN1(n4300), .IN2(n5170), .QN(n7279) );
  NAND2X0 U8612 ( .IN1(test_so23), .IN2(n4828), .QN(n5170) );
  NAND2X0 U8613 ( .IN1(n7281), .IN2(n7282), .QN(WX3286) );
  NOR2X0 U8614 ( .IN1(n7283), .IN2(n7284), .QN(n7282) );
  NOR2X0 U8615 ( .IN1(n7285), .IN2(n4256), .QN(n7284) );
  NOR2X0 U8616 ( .IN1(n6946), .IN2(n4335), .QN(n7283) );
  XOR2X1 U8617 ( .IN1(n7286), .IN2(n7287), .Q(n6946) );
  XOR2X1 U8618 ( .IN1(n8948), .IN2(n4125), .Q(n7287) );
  XOR2X1 U8619 ( .IN1(WX4580), .IN2(n3848), .Q(n7286) );
  NOR2X0 U8620 ( .IN1(n7288), .IN2(n7289), .QN(n7281) );
  NOR2X0 U8621 ( .IN1(DFF_547_n1), .IN2(n4291), .QN(n7289) );
  NOR2X0 U8622 ( .IN1(n4300), .IN2(n5171), .QN(n7288) );
  NAND2X0 U8623 ( .IN1(n4816), .IN2(n8616), .QN(n5171) );
  NAND2X0 U8624 ( .IN1(n7290), .IN2(n7291), .QN(WX3284) );
  NOR2X0 U8625 ( .IN1(n7292), .IN2(n7293), .QN(n7291) );
  NOR2X0 U8626 ( .IN1(n7294), .IN2(n4257), .QN(n7293) );
  NOR2X0 U8627 ( .IN1(n6955), .IN2(n4335), .QN(n7292) );
  XOR2X1 U8628 ( .IN1(n7295), .IN2(n7296), .Q(n6955) );
  XOR2X1 U8629 ( .IN1(n8949), .IN2(n3953), .Q(n7296) );
  XOR2X1 U8630 ( .IN1(WX4578), .IN2(n3850), .Q(n7295) );
  NOR2X0 U8631 ( .IN1(n7297), .IN2(n7298), .QN(n7290) );
  NOR2X0 U8632 ( .IN1(DFF_548_n1), .IN2(n4291), .QN(n7298) );
  NOR2X0 U8633 ( .IN1(n4300), .IN2(n5173), .QN(n7297) );
  NAND2X0 U8634 ( .IN1(n4816), .IN2(n8617), .QN(n5173) );
  NAND2X0 U8635 ( .IN1(n7299), .IN2(n7300), .QN(WX3282) );
  NOR2X0 U8636 ( .IN1(n7301), .IN2(n7302), .QN(n7300) );
  NOR2X0 U8637 ( .IN1(n7303), .IN2(n4257), .QN(n7302) );
  NOR2X0 U8638 ( .IN1(n6964), .IN2(n4335), .QN(n7301) );
  XOR2X1 U8639 ( .IN1(n7304), .IN2(n7305), .Q(n6964) );
  XOR2X1 U8640 ( .IN1(n8950), .IN2(n4124), .Q(n7305) );
  XOR2X1 U8641 ( .IN1(WX4576), .IN2(n3852), .Q(n7304) );
  NOR2X0 U8642 ( .IN1(n7306), .IN2(n7307), .QN(n7299) );
  NOR2X0 U8643 ( .IN1(DFF_549_n1), .IN2(n4291), .QN(n7307) );
  NOR2X0 U8644 ( .IN1(n4300), .IN2(n5174), .QN(n7306) );
  NAND2X0 U8645 ( .IN1(n4816), .IN2(n8618), .QN(n5174) );
  NAND2X0 U8646 ( .IN1(n7308), .IN2(n7309), .QN(WX3280) );
  NOR2X0 U8647 ( .IN1(n7310), .IN2(n7311), .QN(n7309) );
  NOR2X0 U8648 ( .IN1(n4259), .IN2(n7312), .QN(n7311) );
  NOR2X0 U8649 ( .IN1(n6973), .IN2(n4335), .QN(n7310) );
  XOR2X1 U8650 ( .IN1(n7313), .IN2(n7314), .Q(n6973) );
  XOR2X1 U8651 ( .IN1(n8951), .IN2(n4123), .Q(n7314) );
  XOR2X1 U8652 ( .IN1(WX4574), .IN2(n3854), .Q(n7313) );
  NOR2X0 U8653 ( .IN1(n7315), .IN2(n7316), .QN(n7308) );
  NOR2X0 U8654 ( .IN1(DFF_550_n1), .IN2(n4291), .QN(n7316) );
  NOR2X0 U8655 ( .IN1(n4300), .IN2(n5175), .QN(n7315) );
  NAND2X0 U8656 ( .IN1(n4816), .IN2(n8619), .QN(n5175) );
  NAND2X0 U8657 ( .IN1(n7317), .IN2(n7318), .QN(WX3278) );
  NOR2X0 U8658 ( .IN1(n7319), .IN2(n7320), .QN(n7318) );
  NOR2X0 U8659 ( .IN1(n7321), .IN2(n4256), .QN(n7320) );
  NOR2X0 U8660 ( .IN1(n6982), .IN2(n4335), .QN(n7319) );
  XOR2X1 U8661 ( .IN1(n7322), .IN2(n7323), .Q(n6982) );
  XOR2X1 U8662 ( .IN1(n8952), .IN2(n4122), .Q(n7323) );
  XOR2X1 U8663 ( .IN1(WX4572), .IN2(n3856), .Q(n7322) );
  NOR2X0 U8664 ( .IN1(n7324), .IN2(n7325), .QN(n7317) );
  NOR2X0 U8665 ( .IN1(DFF_551_n1), .IN2(n4291), .QN(n7325) );
  NOR2X0 U8666 ( .IN1(n4300), .IN2(n5176), .QN(n7324) );
  NAND2X0 U8667 ( .IN1(n4811), .IN2(n8620), .QN(n5176) );
  NAND2X0 U8668 ( .IN1(n7326), .IN2(n7327), .QN(WX3276) );
  NOR2X0 U8669 ( .IN1(n7328), .IN2(n7329), .QN(n7327) );
  NOR2X0 U8670 ( .IN1(n4259), .IN2(n7330), .QN(n7329) );
  NOR2X0 U8671 ( .IN1(n6991), .IN2(n4335), .QN(n7328) );
  XOR2X1 U8672 ( .IN1(n7331), .IN2(n7332), .Q(n6991) );
  XOR2X1 U8673 ( .IN1(n8953), .IN2(n4121), .Q(n7332) );
  XOR2X1 U8674 ( .IN1(WX4570), .IN2(n3858), .Q(n7331) );
  NOR2X0 U8675 ( .IN1(n7333), .IN2(n7334), .QN(n7326) );
  NOR2X0 U8676 ( .IN1(DFF_552_n1), .IN2(n4291), .QN(n7334) );
  NOR2X0 U8677 ( .IN1(n4300), .IN2(n5177), .QN(n7333) );
  NAND2X0 U8678 ( .IN1(n4816), .IN2(n8621), .QN(n5177) );
  NAND2X0 U8679 ( .IN1(n7335), .IN2(n7336), .QN(WX3274) );
  NOR2X0 U8680 ( .IN1(n7337), .IN2(n7338), .QN(n7336) );
  NOR2X0 U8681 ( .IN1(n7339), .IN2(n4257), .QN(n7338) );
  NOR2X0 U8682 ( .IN1(n7000), .IN2(n4335), .QN(n7337) );
  XOR2X1 U8683 ( .IN1(n7340), .IN2(n7341), .Q(n7000) );
  XOR2X1 U8684 ( .IN1(n8954), .IN2(n4120), .Q(n7341) );
  XOR2X1 U8685 ( .IN1(WX4568), .IN2(n3860), .Q(n7340) );
  NOR2X0 U8686 ( .IN1(n7342), .IN2(n7343), .QN(n7335) );
  NOR2X0 U8687 ( .IN1(DFF_553_n1), .IN2(n4290), .QN(n7343) );
  NOR2X0 U8688 ( .IN1(n4300), .IN2(n5178), .QN(n7342) );
  NAND2X0 U8689 ( .IN1(n4816), .IN2(n8622), .QN(n5178) );
  NAND2X0 U8690 ( .IN1(n7344), .IN2(n7345), .QN(WX3272) );
  NOR2X0 U8691 ( .IN1(n7346), .IN2(n7347), .QN(n7345) );
  NOR2X0 U8692 ( .IN1(n7348), .IN2(n4256), .QN(n7347) );
  NOR2X0 U8693 ( .IN1(n7009), .IN2(n4335), .QN(n7346) );
  XOR2X1 U8694 ( .IN1(n7349), .IN2(n7350), .Q(n7009) );
  XOR2X1 U8695 ( .IN1(n8955), .IN2(n4119), .Q(n7350) );
  XOR2X1 U8696 ( .IN1(WX4566), .IN2(n3862), .Q(n7349) );
  NOR2X0 U8697 ( .IN1(n7351), .IN2(n7352), .QN(n7344) );
  AND2X1 U8698 ( .IN1(n2152), .IN2(test_so31), .Q(n7352) );
  NOR2X0 U8699 ( .IN1(n4300), .IN2(n5179), .QN(n7351) );
  NAND2X0 U8700 ( .IN1(n4816), .IN2(n8623), .QN(n5179) );
  NAND2X0 U8701 ( .IN1(n7353), .IN2(n7354), .QN(WX3270) );
  NOR2X0 U8702 ( .IN1(n7355), .IN2(n7356), .QN(n7354) );
  NOR2X0 U8703 ( .IN1(n7357), .IN2(n4257), .QN(n7356) );
  NOR2X0 U8704 ( .IN1(n4338), .IN2(n7018), .QN(n7355) );
  XNOR2X1 U8705 ( .IN1(n7358), .IN2(n7359), .Q(n7018) );
  XOR2X1 U8706 ( .IN1(test_so41), .IN2(n8956), .Q(n7359) );
  XOR2X1 U8707 ( .IN1(WX4564), .IN2(n3864), .Q(n7358) );
  NOR2X0 U8708 ( .IN1(n7360), .IN2(n7361), .QN(n7353) );
  NOR2X0 U8709 ( .IN1(DFF_555_n1), .IN2(n4290), .QN(n7361) );
  NOR2X0 U8710 ( .IN1(n4300), .IN2(n5180), .QN(n7360) );
  NAND2X0 U8711 ( .IN1(n4816), .IN2(n8624), .QN(n5180) );
  NAND2X0 U8712 ( .IN1(n7362), .IN2(n7363), .QN(WX3268) );
  NOR2X0 U8713 ( .IN1(n7364), .IN2(n7365), .QN(n7363) );
  NOR2X0 U8714 ( .IN1(n4259), .IN2(n7366), .QN(n7365) );
  NOR2X0 U8715 ( .IN1(n7027), .IN2(n4335), .QN(n7364) );
  XOR2X1 U8716 ( .IN1(n7367), .IN2(n7368), .Q(n7027) );
  XOR2X1 U8717 ( .IN1(n8957), .IN2(n4118), .Q(n7368) );
  XOR2X1 U8718 ( .IN1(WX4562), .IN2(n3866), .Q(n7367) );
  NOR2X0 U8719 ( .IN1(n7369), .IN2(n7370), .QN(n7362) );
  NOR2X0 U8720 ( .IN1(DFF_556_n1), .IN2(n4290), .QN(n7370) );
  NOR2X0 U8721 ( .IN1(n4300), .IN2(n5181), .QN(n7369) );
  NAND2X0 U8722 ( .IN1(n4816), .IN2(n8625), .QN(n5181) );
  NAND2X0 U8723 ( .IN1(n7371), .IN2(n7372), .QN(WX3266) );
  NOR2X0 U8724 ( .IN1(n7373), .IN2(n7374), .QN(n7372) );
  NOR2X0 U8725 ( .IN1(n7375), .IN2(n4256), .QN(n7374) );
  NOR2X0 U8726 ( .IN1(n4337), .IN2(n7036), .QN(n7373) );
  XNOR2X1 U8727 ( .IN1(n7376), .IN2(n7377), .Q(n7036) );
  XOR2X1 U8728 ( .IN1(test_so39), .IN2(n8958), .Q(n7377) );
  XOR2X1 U8729 ( .IN1(WX4560), .IN2(n4117), .Q(n7376) );
  NOR2X0 U8730 ( .IN1(n7378), .IN2(n7379), .QN(n7371) );
  NOR2X0 U8731 ( .IN1(DFF_557_n1), .IN2(n4290), .QN(n7379) );
  NOR2X0 U8732 ( .IN1(n4300), .IN2(n5182), .QN(n7378) );
  NAND2X0 U8733 ( .IN1(n4815), .IN2(n8626), .QN(n5182) );
  NAND2X0 U8734 ( .IN1(n7380), .IN2(n7381), .QN(WX3264) );
  NOR2X0 U8735 ( .IN1(n7382), .IN2(n7383), .QN(n7381) );
  NOR2X0 U8736 ( .IN1(n7384), .IN2(n4257), .QN(n7383) );
  NOR2X0 U8737 ( .IN1(n7045), .IN2(n4334), .QN(n7382) );
  XOR2X1 U8738 ( .IN1(n7385), .IN2(n7386), .Q(n7045) );
  XOR2X1 U8739 ( .IN1(n8959), .IN2(n4116), .Q(n7386) );
  XOR2X1 U8740 ( .IN1(WX4558), .IN2(n3869), .Q(n7385) );
  NOR2X0 U8741 ( .IN1(n7387), .IN2(n7388), .QN(n7380) );
  NOR2X0 U8742 ( .IN1(DFF_558_n1), .IN2(n4290), .QN(n7388) );
  NOR2X0 U8743 ( .IN1(n4299), .IN2(n5184), .QN(n7387) );
  NAND2X0 U8744 ( .IN1(n4815), .IN2(n8627), .QN(n5184) );
  NAND2X0 U8745 ( .IN1(n7389), .IN2(n7390), .QN(WX3262) );
  NOR2X0 U8746 ( .IN1(n7391), .IN2(n7392), .QN(n7390) );
  NOR2X0 U8747 ( .IN1(n7393), .IN2(n4256), .QN(n7392) );
  NOR2X0 U8748 ( .IN1(n4337), .IN2(n7054), .QN(n7391) );
  XNOR2X1 U8749 ( .IN1(n7394), .IN2(n7395), .Q(n7054) );
  XOR2X1 U8750 ( .IN1(test_so37), .IN2(n8960), .Q(n7395) );
  XOR2X1 U8751 ( .IN1(WX4556), .IN2(n4115), .Q(n7394) );
  NOR2X0 U8752 ( .IN1(n7396), .IN2(n7397), .QN(n7389) );
  NOR2X0 U8753 ( .IN1(DFF_559_n1), .IN2(n4290), .QN(n7397) );
  NOR2X0 U8754 ( .IN1(n4299), .IN2(n5185), .QN(n7396) );
  NAND2X0 U8755 ( .IN1(n4815), .IN2(n8628), .QN(n5185) );
  NAND2X0 U8756 ( .IN1(n7398), .IN2(n7399), .QN(WX3260) );
  NOR2X0 U8757 ( .IN1(n7400), .IN2(n7401), .QN(n7399) );
  NOR2X0 U8758 ( .IN1(n4259), .IN2(n7402), .QN(n7401) );
  NOR2X0 U8759 ( .IN1(n7063), .IN2(n4334), .QN(n7400) );
  XOR2X1 U8760 ( .IN1(n7403), .IN2(n7404), .Q(n7063) );
  XOR2X1 U8761 ( .IN1(n3655), .IN2(n4776), .Q(n7404) );
  XOR2X1 U8762 ( .IN1(n7405), .IN2(n3952), .Q(n7403) );
  XOR2X1 U8763 ( .IN1(WX4682), .IN2(n8961), .Q(n7405) );
  NOR2X0 U8764 ( .IN1(n7406), .IN2(n7407), .QN(n7398) );
  NOR2X0 U8765 ( .IN1(DFF_560_n1), .IN2(n4290), .QN(n7407) );
  NOR2X0 U8766 ( .IN1(n4299), .IN2(n5186), .QN(n7406) );
  NAND2X0 U8767 ( .IN1(n4815), .IN2(n8629), .QN(n5186) );
  NAND2X0 U8768 ( .IN1(n7408), .IN2(n7409), .QN(WX3258) );
  NOR2X0 U8769 ( .IN1(n7410), .IN2(n7411), .QN(n7409) );
  NOR2X0 U8770 ( .IN1(n7412), .IN2(n4257), .QN(n7411) );
  NOR2X0 U8771 ( .IN1(n4337), .IN2(n7073), .QN(n7410) );
  XNOR2X1 U8772 ( .IN1(n7413), .IN2(n7414), .Q(n7073) );
  XOR2X1 U8773 ( .IN1(n3656), .IN2(n4776), .Q(n7414) );
  XOR2X1 U8774 ( .IN1(n7415), .IN2(n4114), .Q(n7413) );
  XOR2X1 U8775 ( .IN1(WX4616), .IN2(test_so35), .Q(n7415) );
  NOR2X0 U8776 ( .IN1(n7416), .IN2(n7417), .QN(n7408) );
  NOR2X0 U8777 ( .IN1(DFF_561_n1), .IN2(n4290), .QN(n7417) );
  NOR2X0 U8778 ( .IN1(n4299), .IN2(n5187), .QN(n7416) );
  NAND2X0 U8779 ( .IN1(n4815), .IN2(n8630), .QN(n5187) );
  NAND2X0 U8780 ( .IN1(n7418), .IN2(n7419), .QN(WX3256) );
  NOR2X0 U8781 ( .IN1(n7420), .IN2(n7421), .QN(n7419) );
  NOR2X0 U8782 ( .IN1(n7422), .IN2(n4257), .QN(n7421) );
  NOR2X0 U8783 ( .IN1(n7083), .IN2(n4334), .QN(n7420) );
  XOR2X1 U8784 ( .IN1(n7423), .IN2(n7424), .Q(n7083) );
  XOR2X1 U8785 ( .IN1(n3657), .IN2(n4776), .Q(n7424) );
  XOR2X1 U8786 ( .IN1(n7425), .IN2(n4113), .Q(n7423) );
  XOR2X1 U8787 ( .IN1(WX4678), .IN2(n8962), .Q(n7425) );
  NOR2X0 U8788 ( .IN1(n7426), .IN2(n7427), .QN(n7418) );
  NOR2X0 U8789 ( .IN1(DFF_562_n1), .IN2(n4290), .QN(n7427) );
  NOR2X0 U8790 ( .IN1(n4299), .IN2(n5188), .QN(n7426) );
  NAND2X0 U8791 ( .IN1(n4815), .IN2(n8631), .QN(n5188) );
  NAND2X0 U8792 ( .IN1(n7428), .IN2(n7429), .QN(WX3254) );
  NOR2X0 U8793 ( .IN1(n7430), .IN2(n7431), .QN(n7429) );
  NOR2X0 U8794 ( .IN1(n7432), .IN2(n4256), .QN(n7431) );
  NOR2X0 U8795 ( .IN1(n7093), .IN2(n4334), .QN(n7430) );
  XOR2X1 U8796 ( .IN1(n7433), .IN2(n7434), .Q(n7093) );
  XOR2X1 U8797 ( .IN1(n3658), .IN2(n4776), .Q(n7434) );
  XOR2X1 U8798 ( .IN1(n7435), .IN2(n4112), .Q(n7433) );
  XOR2X1 U8799 ( .IN1(WX4676), .IN2(n8963), .Q(n7435) );
  NOR2X0 U8800 ( .IN1(n7436), .IN2(n7437), .QN(n7428) );
  NOR2X0 U8801 ( .IN1(DFF_563_n1), .IN2(n4290), .QN(n7437) );
  NOR2X0 U8802 ( .IN1(n4299), .IN2(n5189), .QN(n7436) );
  NAND2X0 U8803 ( .IN1(n4815), .IN2(n8632), .QN(n5189) );
  NAND2X0 U8804 ( .IN1(n7438), .IN2(n7439), .QN(WX3252) );
  NOR2X0 U8805 ( .IN1(n7440), .IN2(n7441), .QN(n7439) );
  NOR2X0 U8806 ( .IN1(n7442), .IN2(n4257), .QN(n7441) );
  NOR2X0 U8807 ( .IN1(n7103), .IN2(n4334), .QN(n7440) );
  XOR2X1 U8808 ( .IN1(n7443), .IN2(n7444), .Q(n7103) );
  XOR2X1 U8809 ( .IN1(n3659), .IN2(n4776), .Q(n7444) );
  XOR2X1 U8810 ( .IN1(n7445), .IN2(n4111), .Q(n7443) );
  XOR2X1 U8811 ( .IN1(WX4674), .IN2(n8964), .Q(n7445) );
  NOR2X0 U8812 ( .IN1(n7446), .IN2(n7447), .QN(n7438) );
  NOR2X0 U8813 ( .IN1(DFF_564_n1), .IN2(n4290), .QN(n7447) );
  NOR2X0 U8814 ( .IN1(n4299), .IN2(n5190), .QN(n7446) );
  NAND2X0 U8815 ( .IN1(test_so22), .IN2(n4827), .QN(n5190) );
  NAND2X0 U8816 ( .IN1(n7448), .IN2(n7449), .QN(WX3250) );
  NOR2X0 U8817 ( .IN1(n7450), .IN2(n7451), .QN(n7449) );
  NOR2X0 U8818 ( .IN1(n7452), .IN2(n4255), .QN(n7451) );
  NOR2X0 U8819 ( .IN1(n7113), .IN2(n4334), .QN(n7450) );
  XOR2X1 U8820 ( .IN1(n7453), .IN2(n7454), .Q(n7113) );
  XOR2X1 U8821 ( .IN1(n3660), .IN2(n4776), .Q(n7454) );
  XOR2X1 U8822 ( .IN1(n7455), .IN2(n4110), .Q(n7453) );
  XOR2X1 U8823 ( .IN1(WX4672), .IN2(n8965), .Q(n7455) );
  NOR2X0 U8824 ( .IN1(n7456), .IN2(n7457), .QN(n7448) );
  NOR2X0 U8825 ( .IN1(DFF_565_n1), .IN2(n4290), .QN(n7457) );
  NOR2X0 U8826 ( .IN1(n4299), .IN2(n5191), .QN(n7456) );
  NAND2X0 U8827 ( .IN1(n4815), .IN2(n8635), .QN(n5191) );
  NAND2X0 U8828 ( .IN1(n7458), .IN2(n7459), .QN(WX3248) );
  NOR2X0 U8829 ( .IN1(n7460), .IN2(n7461), .QN(n7459) );
  NOR2X0 U8830 ( .IN1(n7462), .IN2(n4256), .QN(n7461) );
  NOR2X0 U8831 ( .IN1(n7123), .IN2(n4334), .QN(n7460) );
  XOR2X1 U8832 ( .IN1(n7463), .IN2(n7464), .Q(n7123) );
  XOR2X1 U8833 ( .IN1(n3661), .IN2(n4776), .Q(n7464) );
  XOR2X1 U8834 ( .IN1(n7465), .IN2(n4109), .Q(n7463) );
  XOR2X1 U8835 ( .IN1(WX4670), .IN2(n8966), .Q(n7465) );
  NOR2X0 U8836 ( .IN1(n7466), .IN2(n7467), .QN(n7458) );
  NOR2X0 U8837 ( .IN1(DFF_566_n1), .IN2(n4290), .QN(n7467) );
  NOR2X0 U8838 ( .IN1(n4299), .IN2(n5192), .QN(n7466) );
  NAND2X0 U8839 ( .IN1(n4815), .IN2(n8636), .QN(n5192) );
  NAND2X0 U8840 ( .IN1(n7468), .IN2(n7469), .QN(WX3246) );
  NOR2X0 U8841 ( .IN1(n7470), .IN2(n7471), .QN(n7469) );
  NOR2X0 U8842 ( .IN1(n4258), .IN2(n7472), .QN(n7471) );
  NOR2X0 U8843 ( .IN1(n7133), .IN2(n4334), .QN(n7470) );
  XOR2X1 U8844 ( .IN1(n7473), .IN2(n7474), .Q(n7133) );
  XOR2X1 U8845 ( .IN1(n3662), .IN2(n4776), .Q(n7474) );
  XOR2X1 U8846 ( .IN1(n7475), .IN2(n4108), .Q(n7473) );
  XOR2X1 U8847 ( .IN1(WX4668), .IN2(n8967), .Q(n7475) );
  NOR2X0 U8848 ( .IN1(n7476), .IN2(n7477), .QN(n7468) );
  NOR2X0 U8849 ( .IN1(DFF_567_n1), .IN2(n4290), .QN(n7477) );
  NOR2X0 U8850 ( .IN1(n4299), .IN2(n5193), .QN(n7476) );
  NAND2X0 U8851 ( .IN1(n4814), .IN2(n8637), .QN(n5193) );
  NAND2X0 U8852 ( .IN1(n7478), .IN2(n7479), .QN(WX3244) );
  NOR2X0 U8853 ( .IN1(n7480), .IN2(n7481), .QN(n7479) );
  NOR2X0 U8854 ( .IN1(n7482), .IN2(n4255), .QN(n7481) );
  NOR2X0 U8855 ( .IN1(n7143), .IN2(n4334), .QN(n7480) );
  XOR2X1 U8856 ( .IN1(n7483), .IN2(n7484), .Q(n7143) );
  XOR2X1 U8857 ( .IN1(n3663), .IN2(n4777), .Q(n7484) );
  XOR2X1 U8858 ( .IN1(n7485), .IN2(n4107), .Q(n7483) );
  XOR2X1 U8859 ( .IN1(WX4666), .IN2(n8968), .Q(n7485) );
  NOR2X0 U8860 ( .IN1(n7486), .IN2(n7487), .QN(n7478) );
  NOR2X0 U8861 ( .IN1(DFF_568_n1), .IN2(n4289), .QN(n7487) );
  NOR2X0 U8862 ( .IN1(n4299), .IN2(n5195), .QN(n7486) );
  NAND2X0 U8863 ( .IN1(n4814), .IN2(n8638), .QN(n5195) );
  NAND2X0 U8864 ( .IN1(n7488), .IN2(n7489), .QN(WX3242) );
  NOR2X0 U8865 ( .IN1(n7490), .IN2(n7491), .QN(n7489) );
  NOR2X0 U8866 ( .IN1(n7492), .IN2(n4253), .QN(n7491) );
  NOR2X0 U8867 ( .IN1(n7153), .IN2(n4334), .QN(n7490) );
  XOR2X1 U8868 ( .IN1(n7493), .IN2(n7494), .Q(n7153) );
  XOR2X1 U8869 ( .IN1(n3664), .IN2(n4777), .Q(n7494) );
  XOR2X1 U8870 ( .IN1(n7495), .IN2(n4106), .Q(n7493) );
  XOR2X1 U8871 ( .IN1(WX4664), .IN2(n8969), .Q(n7495) );
  NOR2X0 U8872 ( .IN1(n7496), .IN2(n7497), .QN(n7488) );
  NOR2X0 U8873 ( .IN1(DFF_569_n1), .IN2(n4289), .QN(n7497) );
  NOR2X0 U8874 ( .IN1(n4299), .IN2(n5196), .QN(n7496) );
  NAND2X0 U8875 ( .IN1(n4814), .IN2(n8639), .QN(n5196) );
  NAND2X0 U8876 ( .IN1(n7498), .IN2(n7499), .QN(WX3240) );
  NOR2X0 U8877 ( .IN1(n7500), .IN2(n7501), .QN(n7499) );
  NOR2X0 U8878 ( .IN1(n4258), .IN2(n7502), .QN(n7501) );
  NOR2X0 U8879 ( .IN1(n7163), .IN2(n4334), .QN(n7500) );
  XOR2X1 U8880 ( .IN1(n7503), .IN2(n7504), .Q(n7163) );
  XOR2X1 U8881 ( .IN1(n3665), .IN2(n4777), .Q(n7504) );
  XOR2X1 U8882 ( .IN1(n7505), .IN2(n4105), .Q(n7503) );
  XOR2X1 U8883 ( .IN1(WX4662), .IN2(n8970), .Q(n7505) );
  NOR2X0 U8884 ( .IN1(n7506), .IN2(n7507), .QN(n7498) );
  NOR2X0 U8885 ( .IN1(DFF_570_n1), .IN2(n4289), .QN(n7507) );
  NOR2X0 U8886 ( .IN1(n4298), .IN2(n5197), .QN(n7506) );
  NAND2X0 U8887 ( .IN1(n4814), .IN2(n8640), .QN(n5197) );
  NAND2X0 U8888 ( .IN1(n7508), .IN2(n7509), .QN(WX3238) );
  NOR2X0 U8889 ( .IN1(n7510), .IN2(n7511), .QN(n7509) );
  NOR2X0 U8890 ( .IN1(n7512), .IN2(n4255), .QN(n7511) );
  NOR2X0 U8891 ( .IN1(n7173), .IN2(n4334), .QN(n7510) );
  XOR2X1 U8892 ( .IN1(n7513), .IN2(n7514), .Q(n7173) );
  XOR2X1 U8893 ( .IN1(n3666), .IN2(n4777), .Q(n7514) );
  XOR2X1 U8894 ( .IN1(n7515), .IN2(n4104), .Q(n7513) );
  XOR2X1 U8895 ( .IN1(WX4660), .IN2(n8971), .Q(n7515) );
  NOR2X0 U8896 ( .IN1(n7516), .IN2(n7517), .QN(n7508) );
  AND2X1 U8897 ( .IN1(n2152), .IN2(test_so32), .Q(n7517) );
  NOR2X0 U8898 ( .IN1(n4298), .IN2(n5198), .QN(n7516) );
  NAND2X0 U8899 ( .IN1(n4814), .IN2(n8641), .QN(n5198) );
  NAND2X0 U8900 ( .IN1(n7518), .IN2(n7519), .QN(WX3236) );
  NOR2X0 U8901 ( .IN1(n7520), .IN2(n7521), .QN(n7519) );
  NOR2X0 U8902 ( .IN1(n7522), .IN2(n4255), .QN(n7521) );
  NOR2X0 U8903 ( .IN1(n4339), .IN2(n7183), .QN(n7520) );
  XNOR2X1 U8904 ( .IN1(n7523), .IN2(n7524), .Q(n7183) );
  XOR2X1 U8905 ( .IN1(n3667), .IN2(n4777), .Q(n7524) );
  XOR2X1 U8906 ( .IN1(WX4594), .IN2(n7525), .Q(n7523) );
  XOR2X1 U8907 ( .IN1(test_so40), .IN2(n8972), .Q(n7525) );
  NOR2X0 U8908 ( .IN1(n7526), .IN2(n7527), .QN(n7518) );
  NOR2X0 U8909 ( .IN1(DFF_572_n1), .IN2(n4289), .QN(n7527) );
  NOR2X0 U8910 ( .IN1(n4298), .IN2(n5199), .QN(n7526) );
  NAND2X0 U8911 ( .IN1(n4814), .IN2(n8642), .QN(n5199) );
  NAND2X0 U8912 ( .IN1(n7528), .IN2(n7529), .QN(WX3234) );
  NOR2X0 U8913 ( .IN1(n7530), .IN2(n7531), .QN(n7529) );
  NOR2X0 U8914 ( .IN1(n7532), .IN2(n4255), .QN(n7531) );
  NOR2X0 U8915 ( .IN1(n7193), .IN2(n4334), .QN(n7530) );
  XOR2X1 U8916 ( .IN1(n7533), .IN2(n7534), .Q(n7193) );
  XOR2X1 U8917 ( .IN1(n3668), .IN2(n4777), .Q(n7534) );
  XOR2X1 U8918 ( .IN1(n7535), .IN2(n4103), .Q(n7533) );
  XOR2X1 U8919 ( .IN1(WX4656), .IN2(n8973), .Q(n7535) );
  NOR2X0 U8920 ( .IN1(n7536), .IN2(n7537), .QN(n7528) );
  NOR2X0 U8921 ( .IN1(DFF_573_n1), .IN2(n4289), .QN(n7537) );
  NOR2X0 U8922 ( .IN1(n4298), .IN2(n5200), .QN(n7536) );
  NAND2X0 U8923 ( .IN1(n4814), .IN2(n8643), .QN(n5200) );
  NAND2X0 U8924 ( .IN1(n7538), .IN2(n7539), .QN(WX3232) );
  NOR2X0 U8925 ( .IN1(n7540), .IN2(n7541), .QN(n7539) );
  NOR2X0 U8926 ( .IN1(n4258), .IN2(n7542), .QN(n7541) );
  NOR2X0 U8927 ( .IN1(n4338), .IN2(n7203), .QN(n7540) );
  XNOR2X1 U8928 ( .IN1(n7543), .IN2(n7544), .Q(n7203) );
  XOR2X1 U8929 ( .IN1(n4102), .IN2(n4777), .Q(n7544) );
  XOR2X1 U8930 ( .IN1(n7545), .IN2(n8976), .Q(n7543) );
  XOR2X1 U8931 ( .IN1(n8975), .IN2(n8974), .Q(n7545) );
  NOR2X0 U8932 ( .IN1(n7546), .IN2(n7547), .QN(n7538) );
  NOR2X0 U8933 ( .IN1(DFF_574_n1), .IN2(n4289), .QN(n7547) );
  NOR2X0 U8934 ( .IN1(n4298), .IN2(n5201), .QN(n7546) );
  NAND2X0 U8935 ( .IN1(n4814), .IN2(n8644), .QN(n5201) );
  NAND2X0 U8936 ( .IN1(n7548), .IN2(n7549), .QN(WX3230) );
  NOR2X0 U8937 ( .IN1(n7550), .IN2(n7551), .QN(n7549) );
  NOR2X0 U8938 ( .IN1(n7552), .IN2(n4254), .QN(n7551) );
  NOR2X0 U8939 ( .IN1(n7213), .IN2(n4334), .QN(n7550) );
  XOR2X1 U8940 ( .IN1(n7553), .IN2(n7554), .Q(n7213) );
  XOR2X1 U8941 ( .IN1(n3587), .IN2(n4777), .Q(n7554) );
  XOR2X1 U8942 ( .IN1(n7555), .IN2(n4101), .Q(n7553) );
  XOR2X1 U8943 ( .IN1(WX4652), .IN2(n8977), .Q(n7555) );
  NOR2X0 U8944 ( .IN1(n7556), .IN2(n7557), .QN(n7548) );
  NOR2X0 U8945 ( .IN1(n3937), .IN2(n5606), .QN(n7557) );
  NOR2X0 U8946 ( .IN1(DFF_575_n1), .IN2(n4289), .QN(n7556) );
  AND2X1 U8947 ( .IN1(n4801), .IN2(n3937), .Q(WX3132) );
  NOR2X0 U8948 ( .IN1(n4925), .IN2(n7558), .QN(WX2619) );
  XOR2X1 U8949 ( .IN1(n4154), .IN2(DFF_382_n1), .Q(n7558) );
  NOR2X0 U8950 ( .IN1(n4925), .IN2(n7559), .QN(WX2617) );
  XOR2X1 U8951 ( .IN1(n4155), .IN2(DFF_381_n1), .Q(n7559) );
  NOR2X0 U8952 ( .IN1(n4926), .IN2(n7560), .QN(WX2615) );
  XOR2X1 U8953 ( .IN1(n4156), .IN2(DFF_380_n1), .Q(n7560) );
  NOR2X0 U8954 ( .IN1(n4925), .IN2(n7561), .QN(WX2613) );
  XNOR2X1 U8955 ( .IN1(DFF_379_n1), .IN2(test_so18), .Q(n7561) );
  NOR2X0 U8956 ( .IN1(n4926), .IN2(n7562), .QN(WX2611) );
  XOR2X1 U8957 ( .IN1(n4157), .IN2(DFF_378_n1), .Q(n7562) );
  NOR2X0 U8958 ( .IN1(n4926), .IN2(n7563), .QN(WX2609) );
  XNOR2X1 U8959 ( .IN1(n4158), .IN2(test_so21), .Q(n7563) );
  NOR2X0 U8960 ( .IN1(n4925), .IN2(n7564), .QN(WX2607) );
  XOR2X1 U8961 ( .IN1(n4159), .IN2(DFF_376_n1), .Q(n7564) );
  NOR2X0 U8962 ( .IN1(n4925), .IN2(n7565), .QN(WX2605) );
  XOR2X1 U8963 ( .IN1(n4160), .IN2(DFF_375_n1), .Q(n7565) );
  NOR2X0 U8964 ( .IN1(n4926), .IN2(n7566), .QN(WX2603) );
  XOR2X1 U8965 ( .IN1(n4161), .IN2(DFF_374_n1), .Q(n7566) );
  NOR2X0 U8966 ( .IN1(n4925), .IN2(n7567), .QN(WX2601) );
  XOR2X1 U8967 ( .IN1(n4162), .IN2(DFF_373_n1), .Q(n7567) );
  NOR2X0 U8968 ( .IN1(n4925), .IN2(n7568), .QN(WX2599) );
  XOR2X1 U8969 ( .IN1(n4163), .IN2(DFF_372_n1), .Q(n7568) );
  NOR2X0 U8970 ( .IN1(n4925), .IN2(n7569), .QN(WX2597) );
  XOR2X1 U8971 ( .IN1(n4164), .IN2(DFF_371_n1), .Q(n7569) );
  NOR2X0 U8972 ( .IN1(n4925), .IN2(n7570), .QN(WX2595) );
  XOR2X1 U8973 ( .IN1(n4165), .IN2(DFF_370_n1), .Q(n7570) );
  NOR2X0 U8974 ( .IN1(n4924), .IN2(n7571), .QN(WX2593) );
  XOR2X1 U8975 ( .IN1(n4166), .IN2(DFF_369_n1), .Q(n7571) );
  NOR2X0 U8976 ( .IN1(n4924), .IN2(n7572), .QN(WX2591) );
  XOR2X1 U8977 ( .IN1(n4167), .IN2(DFF_368_n1), .Q(n7572) );
  NOR2X0 U8978 ( .IN1(n4925), .IN2(n7573), .QN(WX2589) );
  XNOR2X1 U8979 ( .IN1(DFF_367_n1), .IN2(n7574), .Q(n7573) );
  XOR2X1 U8980 ( .IN1(n3957), .IN2(DFF_383_n1), .Q(n7574) );
  NOR2X0 U8981 ( .IN1(n4924), .IN2(n7575), .QN(WX2587) );
  XOR2X1 U8982 ( .IN1(n4168), .IN2(DFF_366_n1), .Q(n7575) );
  NOR2X0 U8983 ( .IN1(n4924), .IN2(n7576), .QN(WX2585) );
  XOR2X1 U8984 ( .IN1(n4169), .IN2(DFF_365_n1), .Q(n7576) );
  NOR2X0 U8985 ( .IN1(n4924), .IN2(n7577), .QN(WX2583) );
  XOR2X1 U8986 ( .IN1(n4170), .IN2(DFF_364_n1), .Q(n7577) );
  NOR2X0 U8987 ( .IN1(n4924), .IN2(n7578), .QN(WX2581) );
  XOR2X1 U8988 ( .IN1(n4171), .IN2(DFF_363_n1), .Q(n7578) );
  NOR2X0 U8989 ( .IN1(n4925), .IN2(n7579), .QN(WX2579) );
  XNOR2X1 U8990 ( .IN1(DFF_362_n1), .IN2(n7580), .Q(n7579) );
  XOR2X1 U8991 ( .IN1(n3958), .IN2(DFF_383_n1), .Q(n7580) );
  NOR2X0 U8992 ( .IN1(n4926), .IN2(n7581), .QN(WX2577) );
  XNOR2X1 U8993 ( .IN1(DFF_361_n1), .IN2(test_so19), .Q(n7581) );
  NOR2X0 U8994 ( .IN1(n4924), .IN2(n7582), .QN(WX2575) );
  XOR2X1 U8995 ( .IN1(n4172), .IN2(DFF_360_n1), .Q(n7582) );
  NOR2X0 U8996 ( .IN1(n4925), .IN2(n7583), .QN(WX2573) );
  XNOR2X1 U8997 ( .IN1(n4173), .IN2(test_so20), .Q(n7583) );
  NOR2X0 U8998 ( .IN1(n4924), .IN2(n7584), .QN(WX2571) );
  XOR2X1 U8999 ( .IN1(n4174), .IN2(DFF_358_n1), .Q(n7584) );
  NOR2X0 U9000 ( .IN1(n4924), .IN2(n7585), .QN(WX2569) );
  XOR2X1 U9001 ( .IN1(n4175), .IN2(DFF_357_n1), .Q(n7585) );
  NOR2X0 U9002 ( .IN1(n4925), .IN2(n7586), .QN(WX2567) );
  XOR2X1 U9003 ( .IN1(n4176), .IN2(DFF_356_n1), .Q(n7586) );
  NOR2X0 U9004 ( .IN1(n4924), .IN2(n7587), .QN(WX2565) );
  XNOR2X1 U9005 ( .IN1(DFF_355_n1), .IN2(n7588), .Q(n7587) );
  XOR2X1 U9006 ( .IN1(n3959), .IN2(DFF_383_n1), .Q(n7588) );
  NOR2X0 U9007 ( .IN1(n4924), .IN2(n7589), .QN(WX2563) );
  XOR2X1 U9008 ( .IN1(n4177), .IN2(DFF_354_n1), .Q(n7589) );
  NOR2X0 U9009 ( .IN1(n4926), .IN2(n7590), .QN(WX2561) );
  XOR2X1 U9010 ( .IN1(n4178), .IN2(DFF_353_n1), .Q(n7590) );
  NOR2X0 U9011 ( .IN1(n4924), .IN2(n7591), .QN(WX2559) );
  XOR2X1 U9012 ( .IN1(n4179), .IN2(DFF_352_n1), .Q(n7591) );
  NOR2X0 U9013 ( .IN1(n4927), .IN2(n7592), .QN(WX2557) );
  XOR2X1 U9014 ( .IN1(n3967), .IN2(DFF_383_n1), .Q(n7592) );
  NOR2X0 U9015 ( .IN1(n9010), .IN2(n4855), .QN(WX2031) );
  NOR2X0 U9016 ( .IN1(n9011), .IN2(n4855), .QN(WX2029) );
  NOR2X0 U9017 ( .IN1(n9013), .IN2(n4855), .QN(WX2027) );
  NOR2X0 U9018 ( .IN1(n9017), .IN2(n4855), .QN(WX2025) );
  NOR2X0 U9019 ( .IN1(n9019), .IN2(n4855), .QN(WX2023) );
  NOR2X0 U9020 ( .IN1(n9021), .IN2(n4855), .QN(WX2021) );
  AND2X1 U9021 ( .IN1(n4801), .IN2(test_so13), .Q(WX2019) );
  NOR2X0 U9022 ( .IN1(n9024), .IN2(n4855), .QN(WX2017) );
  NOR2X0 U9023 ( .IN1(n9026), .IN2(n4854), .QN(WX2015) );
  NOR2X0 U9024 ( .IN1(n9028), .IN2(n4854), .QN(WX2013) );
  NOR2X0 U9025 ( .IN1(n9030), .IN2(n4854), .QN(WX2011) );
  NOR2X0 U9026 ( .IN1(n9034), .IN2(n4854), .QN(WX2009) );
  NOR2X0 U9027 ( .IN1(n9036), .IN2(n4854), .QN(WX2007) );
  NOR2X0 U9028 ( .IN1(n9038), .IN2(n4854), .QN(WX2005) );
  NOR2X0 U9029 ( .IN1(n9040), .IN2(n4854), .QN(WX2003) );
  NOR2X0 U9030 ( .IN1(n9045), .IN2(n4854), .QN(WX2001) );
  NAND2X0 U9031 ( .IN1(n7593), .IN2(n7594), .QN(WX1999) );
  NOR2X0 U9032 ( .IN1(n7595), .IN2(n7596), .QN(n7594) );
  NOR2X0 U9033 ( .IN1(n7258), .IN2(n4333), .QN(n7596) );
  XOR2X1 U9034 ( .IN1(n7597), .IN2(n7598), .Q(n7258) );
  XOR2X1 U9035 ( .IN1(n8979), .IN2(n3966), .Q(n7598) );
  XOR2X1 U9036 ( .IN1(WX3293), .IN2(n3872), .Q(n7597) );
  NOR2X0 U9037 ( .IN1(n4258), .IN2(n6292), .QN(n7595) );
  XNOR2X1 U9038 ( .IN1(n7599), .IN2(n7600), .Q(n6292) );
  XOR2X1 U9039 ( .IN1(test_so16), .IN2(n8978), .Q(n7600) );
  XOR2X1 U9040 ( .IN1(WX2000), .IN2(n3967), .Q(n7599) );
  NOR2X0 U9041 ( .IN1(n7601), .IN2(n7602), .QN(n7593) );
  NOR2X0 U9042 ( .IN1(DFF_352_n1), .IN2(n4291), .QN(n7602) );
  NOR2X0 U9043 ( .IN1(n4298), .IN2(n5202), .QN(n7601) );
  NAND2X0 U9044 ( .IN1(n4814), .IN2(n8670), .QN(n5202) );
  NAND2X0 U9045 ( .IN1(n7603), .IN2(n7604), .QN(WX1997) );
  NOR2X0 U9046 ( .IN1(n7605), .IN2(n7606), .QN(n7604) );
  NOR2X0 U9047 ( .IN1(n7267), .IN2(n4333), .QN(n7606) );
  XOR2X1 U9048 ( .IN1(n7607), .IN2(n7608), .Q(n7267) );
  XOR2X1 U9049 ( .IN1(n8981), .IN2(n4153), .Q(n7608) );
  XOR2X1 U9050 ( .IN1(WX3291), .IN2(n3874), .Q(n7607) );
  AND2X1 U9051 ( .IN1(n6300), .IN2(n4263), .Q(n7605) );
  XNOR2X1 U9052 ( .IN1(n7609), .IN2(n7610), .Q(n6300) );
  XOR2X1 U9053 ( .IN1(n8980), .IN2(n4179), .Q(n7610) );
  XOR2X1 U9054 ( .IN1(WX1998), .IN2(n3903), .Q(n7609) );
  NOR2X0 U9055 ( .IN1(n7611), .IN2(n7612), .QN(n7603) );
  NOR2X0 U9056 ( .IN1(DFF_353_n1), .IN2(n4289), .QN(n7612) );
  NOR2X0 U9057 ( .IN1(n4298), .IN2(n5203), .QN(n7611) );
  NAND2X0 U9058 ( .IN1(n4813), .IN2(n8671), .QN(n5203) );
  NAND2X0 U9059 ( .IN1(n7613), .IN2(n7614), .QN(WX1995) );
  NOR2X0 U9060 ( .IN1(n7615), .IN2(n7616), .QN(n7614) );
  NOR2X0 U9061 ( .IN1(n7276), .IN2(n4333), .QN(n7616) );
  XOR2X1 U9062 ( .IN1(n7617), .IN2(n7618), .Q(n7276) );
  XOR2X1 U9063 ( .IN1(n8983), .IN2(n4152), .Q(n7618) );
  XOR2X1 U9064 ( .IN1(WX3289), .IN2(n3876), .Q(n7617) );
  AND2X1 U9065 ( .IN1(n6308), .IN2(n4263), .Q(n7615) );
  XNOR2X1 U9066 ( .IN1(n7619), .IN2(n7620), .Q(n6308) );
  XOR2X1 U9067 ( .IN1(n8982), .IN2(n4178), .Q(n7620) );
  XOR2X1 U9068 ( .IN1(WX1996), .IN2(n3905), .Q(n7619) );
  NOR2X0 U9069 ( .IN1(n7621), .IN2(n7622), .QN(n7613) );
  NOR2X0 U9070 ( .IN1(DFF_354_n1), .IN2(n4289), .QN(n7622) );
  NOR2X0 U9071 ( .IN1(n4298), .IN2(n5204), .QN(n7621) );
  NAND2X0 U9072 ( .IN1(n4813), .IN2(n8672), .QN(n5204) );
  NAND2X0 U9073 ( .IN1(n7623), .IN2(n7624), .QN(WX1993) );
  NOR2X0 U9074 ( .IN1(n7625), .IN2(n7626), .QN(n7624) );
  NOR2X0 U9075 ( .IN1(n7285), .IN2(n4333), .QN(n7626) );
  XOR2X1 U9076 ( .IN1(n7627), .IN2(n7628), .Q(n7285) );
  XOR2X1 U9077 ( .IN1(n8985), .IN2(n4151), .Q(n7628) );
  XOR2X1 U9078 ( .IN1(WX3287), .IN2(n3878), .Q(n7627) );
  AND2X1 U9079 ( .IN1(n6316), .IN2(n4263), .Q(n7625) );
  XNOR2X1 U9080 ( .IN1(n7629), .IN2(n7630), .Q(n6316) );
  XOR2X1 U9081 ( .IN1(n8984), .IN2(n4177), .Q(n7630) );
  XOR2X1 U9082 ( .IN1(WX1994), .IN2(n3907), .Q(n7629) );
  NOR2X0 U9083 ( .IN1(n7631), .IN2(n7632), .QN(n7623) );
  NOR2X0 U9084 ( .IN1(DFF_355_n1), .IN2(n4289), .QN(n7632) );
  NOR2X0 U9085 ( .IN1(n4298), .IN2(n5206), .QN(n7631) );
  NAND2X0 U9086 ( .IN1(n4813), .IN2(n8673), .QN(n5206) );
  NAND2X0 U9087 ( .IN1(n7633), .IN2(n7634), .QN(WX1991) );
  NOR2X0 U9088 ( .IN1(n7635), .IN2(n7636), .QN(n7634) );
  NOR2X0 U9089 ( .IN1(n7294), .IN2(n4333), .QN(n7636) );
  XOR2X1 U9090 ( .IN1(n7637), .IN2(n7638), .Q(n7294) );
  XOR2X1 U9091 ( .IN1(n8987), .IN2(n3956), .Q(n7638) );
  XOR2X1 U9092 ( .IN1(WX3285), .IN2(n3880), .Q(n7637) );
  NOR2X0 U9093 ( .IN1(n4258), .IN2(n6324), .QN(n7635) );
  XNOR2X1 U9094 ( .IN1(n7639), .IN2(n7640), .Q(n6324) );
  XOR2X1 U9095 ( .IN1(test_so14), .IN2(n8986), .Q(n7640) );
  XOR2X1 U9096 ( .IN1(WX2120), .IN2(n3959), .Q(n7639) );
  NOR2X0 U9097 ( .IN1(n7641), .IN2(n7642), .QN(n7633) );
  NOR2X0 U9098 ( .IN1(DFF_356_n1), .IN2(n4289), .QN(n7642) );
  NOR2X0 U9099 ( .IN1(n4298), .IN2(n5207), .QN(n7641) );
  NAND2X0 U9100 ( .IN1(n4813), .IN2(n8674), .QN(n5207) );
  NAND2X0 U9101 ( .IN1(n7643), .IN2(n7644), .QN(WX1989) );
  NOR2X0 U9102 ( .IN1(n7645), .IN2(n7646), .QN(n7644) );
  NOR2X0 U9103 ( .IN1(n7303), .IN2(n4332), .QN(n7646) );
  XOR2X1 U9104 ( .IN1(n7647), .IN2(n7648), .Q(n7303) );
  XOR2X1 U9105 ( .IN1(n8989), .IN2(n4150), .Q(n7648) );
  XOR2X1 U9106 ( .IN1(WX3283), .IN2(n3882), .Q(n7647) );
  AND2X1 U9107 ( .IN1(n6332), .IN2(n4263), .Q(n7645) );
  XNOR2X1 U9108 ( .IN1(n7649), .IN2(n7650), .Q(n6332) );
  XOR2X1 U9109 ( .IN1(n8988), .IN2(n4176), .Q(n7650) );
  XOR2X1 U9110 ( .IN1(WX1990), .IN2(n3910), .Q(n7649) );
  NOR2X0 U9111 ( .IN1(n7651), .IN2(n7652), .QN(n7643) );
  NOR2X0 U9112 ( .IN1(DFF_357_n1), .IN2(n4289), .QN(n7652) );
  NOR2X0 U9113 ( .IN1(n4298), .IN2(n5208), .QN(n7651) );
  NAND2X0 U9114 ( .IN1(n4813), .IN2(n8675), .QN(n5208) );
  NAND2X0 U9115 ( .IN1(n7653), .IN2(n7654), .QN(WX1987) );
  NOR2X0 U9116 ( .IN1(n7655), .IN2(n7656), .QN(n7654) );
  NOR2X0 U9117 ( .IN1(n4338), .IN2(n7312), .QN(n7656) );
  XNOR2X1 U9118 ( .IN1(n7657), .IN2(n7658), .Q(n7312) );
  XOR2X1 U9119 ( .IN1(test_so30), .IN2(n8991), .Q(n7658) );
  XOR2X1 U9120 ( .IN1(WX3281), .IN2(n3884), .Q(n7657) );
  AND2X1 U9121 ( .IN1(n6340), .IN2(n4263), .Q(n7655) );
  XNOR2X1 U9122 ( .IN1(n7659), .IN2(n7660), .Q(n6340) );
  XOR2X1 U9123 ( .IN1(n8990), .IN2(n4175), .Q(n7660) );
  XOR2X1 U9124 ( .IN1(WX1988), .IN2(n3912), .Q(n7659) );
  NOR2X0 U9125 ( .IN1(n7661), .IN2(n7662), .QN(n7653) );
  NOR2X0 U9126 ( .IN1(DFF_358_n1), .IN2(n4289), .QN(n7662) );
  NOR2X0 U9127 ( .IN1(n4298), .IN2(n5209), .QN(n7661) );
  NAND2X0 U9128 ( .IN1(n4813), .IN2(n8676), .QN(n5209) );
  NAND2X0 U9129 ( .IN1(n7663), .IN2(n7664), .QN(WX1985) );
  NOR2X0 U9130 ( .IN1(n7665), .IN2(n7666), .QN(n7664) );
  NOR2X0 U9131 ( .IN1(n7321), .IN2(n4333), .QN(n7666) );
  XOR2X1 U9132 ( .IN1(n7667), .IN2(n7668), .Q(n7321) );
  XOR2X1 U9133 ( .IN1(n8993), .IN2(n4149), .Q(n7668) );
  XOR2X1 U9134 ( .IN1(WX3279), .IN2(n3886), .Q(n7667) );
  AND2X1 U9135 ( .IN1(n6348), .IN2(n4263), .Q(n7665) );
  XNOR2X1 U9136 ( .IN1(n7669), .IN2(n7670), .Q(n6348) );
  XOR2X1 U9137 ( .IN1(n8992), .IN2(n4174), .Q(n7670) );
  XOR2X1 U9138 ( .IN1(WX1986), .IN2(n3914), .Q(n7669) );
  NOR2X0 U9139 ( .IN1(n7671), .IN2(n7672), .QN(n7663) );
  AND2X1 U9140 ( .IN1(n2152), .IN2(test_so20), .Q(n7672) );
  NOR2X0 U9141 ( .IN1(n4297), .IN2(n5210), .QN(n7671) );
  NAND2X0 U9142 ( .IN1(n4813), .IN2(n8677), .QN(n5210) );
  NAND2X0 U9143 ( .IN1(n7673), .IN2(n7674), .QN(WX1983) );
  NOR2X0 U9144 ( .IN1(n7675), .IN2(n7676), .QN(n7674) );
  NOR2X0 U9145 ( .IN1(n4340), .IN2(n7330), .QN(n7676) );
  XNOR2X1 U9146 ( .IN1(n7677), .IN2(n7678), .Q(n7330) );
  XOR2X1 U9147 ( .IN1(test_so28), .IN2(n8995), .Q(n7678) );
  XOR2X1 U9148 ( .IN1(WX3277), .IN2(n4148), .Q(n7677) );
  AND2X1 U9149 ( .IN1(n6356), .IN2(n4263), .Q(n7675) );
  XNOR2X1 U9150 ( .IN1(n7679), .IN2(n7680), .Q(n6356) );
  XOR2X1 U9151 ( .IN1(n8994), .IN2(n4173), .Q(n7680) );
  XOR2X1 U9152 ( .IN1(WX1984), .IN2(n3916), .Q(n7679) );
  NOR2X0 U9153 ( .IN1(n7681), .IN2(n7682), .QN(n7673) );
  NOR2X0 U9154 ( .IN1(DFF_360_n1), .IN2(n4289), .QN(n7682) );
  NOR2X0 U9155 ( .IN1(n4297), .IN2(n5211), .QN(n7681) );
  NAND2X0 U9156 ( .IN1(test_so12), .IN2(n4828), .QN(n5211) );
  NAND2X0 U9157 ( .IN1(n7683), .IN2(n7684), .QN(WX1981) );
  NOR2X0 U9158 ( .IN1(n7685), .IN2(n7686), .QN(n7684) );
  NOR2X0 U9159 ( .IN1(n7339), .IN2(n4333), .QN(n7686) );
  XOR2X1 U9160 ( .IN1(n7687), .IN2(n7688), .Q(n7339) );
  XOR2X1 U9161 ( .IN1(n8997), .IN2(n4147), .Q(n7688) );
  XOR2X1 U9162 ( .IN1(WX3275), .IN2(n3889), .Q(n7687) );
  AND2X1 U9163 ( .IN1(n6364), .IN2(n4263), .Q(n7685) );
  XNOR2X1 U9164 ( .IN1(n7689), .IN2(n7690), .Q(n6364) );
  XOR2X1 U9165 ( .IN1(n8996), .IN2(n4172), .Q(n7690) );
  XOR2X1 U9166 ( .IN1(WX1982), .IN2(n3918), .Q(n7689) );
  NOR2X0 U9167 ( .IN1(n7691), .IN2(n7692), .QN(n7683) );
  NOR2X0 U9168 ( .IN1(DFF_361_n1), .IN2(n4288), .QN(n7692) );
  NOR2X0 U9169 ( .IN1(n4297), .IN2(n5212), .QN(n7691) );
  NAND2X0 U9170 ( .IN1(n4819), .IN2(n8680), .QN(n5212) );
  NAND2X0 U9171 ( .IN1(n7693), .IN2(n7694), .QN(WX1979) );
  NOR2X0 U9172 ( .IN1(n7695), .IN2(n7696), .QN(n7694) );
  NOR2X0 U9173 ( .IN1(n7348), .IN2(n4333), .QN(n7696) );
  XOR2X1 U9174 ( .IN1(n7697), .IN2(n7698), .Q(n7348) );
  XOR2X1 U9175 ( .IN1(n8999), .IN2(n4146), .Q(n7698) );
  XOR2X1 U9176 ( .IN1(WX3273), .IN2(n3891), .Q(n7697) );
  NOR2X0 U9177 ( .IN1(n4259), .IN2(n6372), .QN(n7695) );
  XNOR2X1 U9178 ( .IN1(n7699), .IN2(n7700), .Q(n6372) );
  XOR2X1 U9179 ( .IN1(test_so19), .IN2(n8998), .Q(n7700) );
  XOR2X1 U9180 ( .IN1(WX1980), .IN2(n3920), .Q(n7699) );
  NOR2X0 U9181 ( .IN1(n7701), .IN2(n7702), .QN(n7693) );
  NOR2X0 U9182 ( .IN1(DFF_362_n1), .IN2(n4288), .QN(n7702) );
  NOR2X0 U9183 ( .IN1(n4297), .IN2(n5213), .QN(n7701) );
  NAND2X0 U9184 ( .IN1(n4813), .IN2(n8681), .QN(n5213) );
  NAND2X0 U9185 ( .IN1(n7703), .IN2(n7704), .QN(WX1977) );
  NOR2X0 U9186 ( .IN1(n7705), .IN2(n7706), .QN(n7704) );
  NOR2X0 U9187 ( .IN1(n7357), .IN2(n4333), .QN(n7706) );
  XOR2X1 U9188 ( .IN1(n7707), .IN2(n7708), .Q(n7357) );
  XOR2X1 U9189 ( .IN1(n9001), .IN2(n3955), .Q(n7708) );
  XOR2X1 U9190 ( .IN1(WX3271), .IN2(n3893), .Q(n7707) );
  AND2X1 U9191 ( .IN1(n6380), .IN2(n4263), .Q(n7705) );
  XNOR2X1 U9192 ( .IN1(n7709), .IN2(n7710), .Q(n6380) );
  XOR2X1 U9193 ( .IN1(n9000), .IN2(n3958), .Q(n7710) );
  XOR2X1 U9194 ( .IN1(WX1978), .IN2(n3922), .Q(n7709) );
  NOR2X0 U9195 ( .IN1(n7711), .IN2(n7712), .QN(n7703) );
  NOR2X0 U9196 ( .IN1(DFF_363_n1), .IN2(n4288), .QN(n7712) );
  NOR2X0 U9197 ( .IN1(n4297), .IN2(n5223), .QN(n7711) );
  NAND2X0 U9198 ( .IN1(n4812), .IN2(n8682), .QN(n5223) );
  NAND2X0 U9199 ( .IN1(n7713), .IN2(n7714), .QN(WX1975) );
  NOR2X0 U9200 ( .IN1(n7715), .IN2(n7716), .QN(n7714) );
  NOR2X0 U9201 ( .IN1(n4338), .IN2(n7366), .QN(n7716) );
  XNOR2X1 U9202 ( .IN1(n7717), .IN2(n7718), .Q(n7366) );
  XOR2X1 U9203 ( .IN1(test_so26), .IN2(n9003), .Q(n7718) );
  XOR2X1 U9204 ( .IN1(WX3269), .IN2(n4145), .Q(n7717) );
  AND2X1 U9205 ( .IN1(n6388), .IN2(n4264), .Q(n7715) );
  XNOR2X1 U9206 ( .IN1(n7719), .IN2(n7720), .Q(n6388) );
  XOR2X1 U9207 ( .IN1(n9002), .IN2(n4171), .Q(n7720) );
  XOR2X1 U9208 ( .IN1(WX1976), .IN2(n3924), .Q(n7719) );
  NOR2X0 U9209 ( .IN1(n7721), .IN2(n7722), .QN(n7713) );
  NOR2X0 U9210 ( .IN1(DFF_364_n1), .IN2(n4288), .QN(n7722) );
  NOR2X0 U9211 ( .IN1(n4297), .IN2(n5234), .QN(n7721) );
  NAND2X0 U9212 ( .IN1(n4812), .IN2(n8683), .QN(n5234) );
  NAND2X0 U9213 ( .IN1(n7723), .IN2(n7724), .QN(WX1973) );
  NOR2X0 U9214 ( .IN1(n7725), .IN2(n7726), .QN(n7724) );
  NOR2X0 U9215 ( .IN1(n7375), .IN2(n4335), .QN(n7726) );
  XOR2X1 U9216 ( .IN1(n7727), .IN2(n7728), .Q(n7375) );
  XOR2X1 U9217 ( .IN1(n9005), .IN2(n4144), .Q(n7728) );
  XOR2X1 U9218 ( .IN1(WX3267), .IN2(n3896), .Q(n7727) );
  AND2X1 U9219 ( .IN1(n6396), .IN2(n4264), .Q(n7725) );
  XNOR2X1 U9220 ( .IN1(n7729), .IN2(n7730), .Q(n6396) );
  XOR2X1 U9221 ( .IN1(n9004), .IN2(n4170), .Q(n7730) );
  XOR2X1 U9222 ( .IN1(WX1974), .IN2(n3926), .Q(n7729) );
  NOR2X0 U9223 ( .IN1(n7731), .IN2(n7732), .QN(n7723) );
  NOR2X0 U9224 ( .IN1(DFF_365_n1), .IN2(n4288), .QN(n7732) );
  NOR2X0 U9225 ( .IN1(n4297), .IN2(n5246), .QN(n7731) );
  NAND2X0 U9226 ( .IN1(n4812), .IN2(n8684), .QN(n5246) );
  NAND2X0 U9227 ( .IN1(n7733), .IN2(n7734), .QN(WX1971) );
  NOR2X0 U9228 ( .IN1(n7735), .IN2(n7736), .QN(n7734) );
  NOR2X0 U9229 ( .IN1(n7384), .IN2(n4333), .QN(n7736) );
  XOR2X1 U9230 ( .IN1(n7737), .IN2(n7738), .Q(n7384) );
  XOR2X1 U9231 ( .IN1(n9007), .IN2(n4143), .Q(n7738) );
  XOR2X1 U9232 ( .IN1(WX3265), .IN2(n3898), .Q(n7737) );
  NOR2X0 U9233 ( .IN1(n4258), .IN2(n6404), .QN(n7735) );
  XNOR2X1 U9234 ( .IN1(n7739), .IN2(n7740), .Q(n6404) );
  XOR2X1 U9235 ( .IN1(test_so17), .IN2(n9006), .Q(n7740) );
  XOR2X1 U9236 ( .IN1(WX1972), .IN2(n4169), .Q(n7739) );
  NOR2X0 U9237 ( .IN1(n7741), .IN2(n7742), .QN(n7733) );
  NOR2X0 U9238 ( .IN1(DFF_366_n1), .IN2(n4288), .QN(n7742) );
  NOR2X0 U9239 ( .IN1(n4297), .IN2(n5257), .QN(n7741) );
  NAND2X0 U9240 ( .IN1(n4812), .IN2(n8685), .QN(n5257) );
  NAND2X0 U9241 ( .IN1(n7743), .IN2(n7744), .QN(WX1969) );
  NOR2X0 U9242 ( .IN1(n7745), .IN2(n7746), .QN(n7744) );
  NOR2X0 U9243 ( .IN1(n7393), .IN2(n4333), .QN(n7746) );
  XOR2X1 U9244 ( .IN1(n7747), .IN2(n7748), .Q(n7393) );
  XOR2X1 U9245 ( .IN1(n9009), .IN2(n4142), .Q(n7748) );
  XOR2X1 U9246 ( .IN1(WX3263), .IN2(n3900), .Q(n7747) );
  AND2X1 U9247 ( .IN1(n6412), .IN2(n4264), .Q(n7745) );
  XNOR2X1 U9248 ( .IN1(n7749), .IN2(n7750), .Q(n6412) );
  XOR2X1 U9249 ( .IN1(n9008), .IN2(n4168), .Q(n7750) );
  XOR2X1 U9250 ( .IN1(WX1970), .IN2(n3929), .Q(n7749) );
  NOR2X0 U9251 ( .IN1(n7751), .IN2(n7752), .QN(n7743) );
  NOR2X0 U9252 ( .IN1(DFF_367_n1), .IN2(n4288), .QN(n7752) );
  NOR2X0 U9253 ( .IN1(n4297), .IN2(n5268), .QN(n7751) );
  NAND2X0 U9254 ( .IN1(n4812), .IN2(n8686), .QN(n5268) );
  NAND2X0 U9255 ( .IN1(n7753), .IN2(n7754), .QN(WX1967) );
  NOR2X0 U9256 ( .IN1(n7755), .IN2(n7756), .QN(n7754) );
  NOR2X0 U9257 ( .IN1(n4339), .IN2(n7402), .QN(n7756) );
  XNOR2X1 U9258 ( .IN1(n7757), .IN2(n7758), .Q(n7402) );
  XOR2X1 U9259 ( .IN1(n3669), .IN2(n4777), .Q(n7758) );
  XOR2X1 U9260 ( .IN1(n7759), .IN2(n3954), .Q(n7757) );
  XOR2X1 U9261 ( .IN1(WX3325), .IN2(test_so24), .Q(n7759) );
  AND2X1 U9262 ( .IN1(n6420), .IN2(n4264), .Q(n7755) );
  XNOR2X1 U9263 ( .IN1(n7760), .IN2(n7761), .Q(n6420) );
  XOR2X1 U9264 ( .IN1(n3682), .IN2(n4777), .Q(n7761) );
  XOR2X1 U9265 ( .IN1(n7762), .IN2(n3957), .Q(n7760) );
  XOR2X1 U9266 ( .IN1(WX2096), .IN2(n9010), .Q(n7762) );
  NOR2X0 U9267 ( .IN1(n7763), .IN2(n7764), .QN(n7753) );
  NOR2X0 U9268 ( .IN1(DFF_368_n1), .IN2(n4288), .QN(n7764) );
  NOR2X0 U9269 ( .IN1(n4297), .IN2(n5279), .QN(n7763) );
  NAND2X0 U9270 ( .IN1(n4812), .IN2(n8687), .QN(n5279) );
  NAND2X0 U9271 ( .IN1(n7765), .IN2(n7766), .QN(WX1965) );
  NOR2X0 U9272 ( .IN1(n7767), .IN2(n7768), .QN(n7766) );
  NOR2X0 U9273 ( .IN1(n7412), .IN2(n4333), .QN(n7768) );
  XOR2X1 U9274 ( .IN1(n7769), .IN2(n7770), .Q(n7412) );
  XOR2X1 U9275 ( .IN1(n3670), .IN2(n4777), .Q(n7770) );
  XOR2X1 U9276 ( .IN1(n7771), .IN2(n4141), .Q(n7769) );
  XOR2X1 U9277 ( .IN1(WX3387), .IN2(n9012), .Q(n7771) );
  AND2X1 U9278 ( .IN1(n6428), .IN2(n4264), .Q(n7767) );
  XNOR2X1 U9279 ( .IN1(n7772), .IN2(n7773), .Q(n6428) );
  XOR2X1 U9280 ( .IN1(n3683), .IN2(n4778), .Q(n7773) );
  XOR2X1 U9281 ( .IN1(n7774), .IN2(n4167), .Q(n7772) );
  XOR2X1 U9282 ( .IN1(WX2094), .IN2(n9011), .Q(n7774) );
  NOR2X0 U9283 ( .IN1(n7775), .IN2(n7776), .QN(n7765) );
  NOR2X0 U9284 ( .IN1(DFF_369_n1), .IN2(n4288), .QN(n7776) );
  NOR2X0 U9285 ( .IN1(n4297), .IN2(n5290), .QN(n7775) );
  NAND2X0 U9286 ( .IN1(n4812), .IN2(n8688), .QN(n5290) );
  NAND2X0 U9287 ( .IN1(n7777), .IN2(n7778), .QN(WX1963) );
  NOR2X0 U9288 ( .IN1(n7779), .IN2(n7780), .QN(n7778) );
  NOR2X0 U9289 ( .IN1(n7422), .IN2(n4333), .QN(n7780) );
  XOR2X1 U9290 ( .IN1(n7781), .IN2(n7782), .Q(n7422) );
  XOR2X1 U9291 ( .IN1(n3671), .IN2(n4778), .Q(n7782) );
  XOR2X1 U9292 ( .IN1(n7783), .IN2(n4140), .Q(n7781) );
  XOR2X1 U9293 ( .IN1(WX3385), .IN2(n9016), .Q(n7783) );
  NOR2X0 U9294 ( .IN1(n4258), .IN2(n6436), .QN(n7779) );
  XNOR2X1 U9295 ( .IN1(n7784), .IN2(n7785), .Q(n6436) );
  XOR2X1 U9296 ( .IN1(n4166), .IN2(n4778), .Q(n7785) );
  XOR2X1 U9297 ( .IN1(n7786), .IN2(n9015), .Q(n7784) );
  XOR2X1 U9298 ( .IN1(n9014), .IN2(n9013), .Q(n7786) );
  NOR2X0 U9299 ( .IN1(n7787), .IN2(n7788), .QN(n7777) );
  NOR2X0 U9300 ( .IN1(DFF_370_n1), .IN2(n4288), .QN(n7788) );
  NOR2X0 U9301 ( .IN1(n4297), .IN2(n5301), .QN(n7787) );
  NAND2X0 U9302 ( .IN1(n4812), .IN2(n8689), .QN(n5301) );
  NAND2X0 U9303 ( .IN1(n7789), .IN2(n7790), .QN(WX1961) );
  NOR2X0 U9304 ( .IN1(n7791), .IN2(n7792), .QN(n7790) );
  NOR2X0 U9305 ( .IN1(n7432), .IN2(n4333), .QN(n7792) );
  XOR2X1 U9306 ( .IN1(n7793), .IN2(n7794), .Q(n7432) );
  XOR2X1 U9307 ( .IN1(n3672), .IN2(n4778), .Q(n7794) );
  XOR2X1 U9308 ( .IN1(n7795), .IN2(n4139), .Q(n7793) );
  XOR2X1 U9309 ( .IN1(WX3383), .IN2(n9018), .Q(n7795) );
  AND2X1 U9310 ( .IN1(n6444), .IN2(n4264), .Q(n7791) );
  XNOR2X1 U9311 ( .IN1(n7796), .IN2(n7797), .Q(n6444) );
  XOR2X1 U9312 ( .IN1(n3684), .IN2(n4778), .Q(n7797) );
  XOR2X1 U9313 ( .IN1(n7798), .IN2(n4165), .Q(n7796) );
  XOR2X1 U9314 ( .IN1(WX2090), .IN2(n9017), .Q(n7798) );
  NOR2X0 U9315 ( .IN1(n7799), .IN2(n7800), .QN(n7789) );
  NOR2X0 U9316 ( .IN1(DFF_371_n1), .IN2(n4288), .QN(n7800) );
  NOR2X0 U9317 ( .IN1(n4296), .IN2(n5312), .QN(n7799) );
  NAND2X0 U9318 ( .IN1(n4812), .IN2(n8690), .QN(n5312) );
  NAND2X0 U9319 ( .IN1(n7801), .IN2(n7802), .QN(WX1959) );
  NOR2X0 U9320 ( .IN1(n7803), .IN2(n7804), .QN(n7802) );
  NOR2X0 U9321 ( .IN1(n7442), .IN2(n4332), .QN(n7804) );
  XOR2X1 U9322 ( .IN1(n7805), .IN2(n7806), .Q(n7442) );
  XOR2X1 U9323 ( .IN1(n3673), .IN2(n4778), .Q(n7806) );
  XOR2X1 U9324 ( .IN1(n7807), .IN2(n4138), .Q(n7805) );
  XOR2X1 U9325 ( .IN1(WX3381), .IN2(n9020), .Q(n7807) );
  AND2X1 U9326 ( .IN1(n6452), .IN2(n4264), .Q(n7803) );
  XNOR2X1 U9327 ( .IN1(n7808), .IN2(n7809), .Q(n6452) );
  XOR2X1 U9328 ( .IN1(n3685), .IN2(n4778), .Q(n7809) );
  XOR2X1 U9329 ( .IN1(n7810), .IN2(n4164), .Q(n7808) );
  XOR2X1 U9330 ( .IN1(WX2088), .IN2(n9019), .Q(n7810) );
  NOR2X0 U9331 ( .IN1(n7811), .IN2(n7812), .QN(n7801) );
  NOR2X0 U9332 ( .IN1(DFF_372_n1), .IN2(n4288), .QN(n7812) );
  NOR2X0 U9333 ( .IN1(n4296), .IN2(n5323), .QN(n7811) );
  NAND2X0 U9334 ( .IN1(n4811), .IN2(n8691), .QN(n5323) );
  NAND2X0 U9335 ( .IN1(n7813), .IN2(n7814), .QN(WX1957) );
  NOR2X0 U9336 ( .IN1(n7815), .IN2(n7816), .QN(n7814) );
  NOR2X0 U9337 ( .IN1(n7452), .IN2(n4332), .QN(n7816) );
  XOR2X1 U9338 ( .IN1(n7817), .IN2(n7818), .Q(n7452) );
  XOR2X1 U9339 ( .IN1(n3674), .IN2(n4778), .Q(n7818) );
  XOR2X1 U9340 ( .IN1(n7819), .IN2(n4137), .Q(n7817) );
  XOR2X1 U9341 ( .IN1(WX3379), .IN2(n9022), .Q(n7819) );
  AND2X1 U9342 ( .IN1(n6460), .IN2(n4264), .Q(n7815) );
  XNOR2X1 U9343 ( .IN1(n7820), .IN2(n7821), .Q(n6460) );
  XOR2X1 U9344 ( .IN1(n3686), .IN2(n4778), .Q(n7821) );
  XOR2X1 U9345 ( .IN1(n7822), .IN2(n4163), .Q(n7820) );
  XOR2X1 U9346 ( .IN1(WX2086), .IN2(n9021), .Q(n7822) );
  NOR2X0 U9347 ( .IN1(n7823), .IN2(n7824), .QN(n7813) );
  NOR2X0 U9348 ( .IN1(DFF_373_n1), .IN2(n4288), .QN(n7824) );
  NOR2X0 U9349 ( .IN1(n4296), .IN2(n5334), .QN(n7823) );
  NAND2X0 U9350 ( .IN1(n4811), .IN2(n8692), .QN(n5334) );
  NAND2X0 U9351 ( .IN1(n7825), .IN2(n7826), .QN(WX1955) );
  NOR2X0 U9352 ( .IN1(n7827), .IN2(n7828), .QN(n7826) );
  NOR2X0 U9353 ( .IN1(n7462), .IN2(n4332), .QN(n7828) );
  XOR2X1 U9354 ( .IN1(n7829), .IN2(n7830), .Q(n7462) );
  XOR2X1 U9355 ( .IN1(n3675), .IN2(n4778), .Q(n7830) );
  XOR2X1 U9356 ( .IN1(n7831), .IN2(n4136), .Q(n7829) );
  XOR2X1 U9357 ( .IN1(WX3377), .IN2(n9023), .Q(n7831) );
  NOR2X0 U9358 ( .IN1(n4259), .IN2(n6468), .QN(n7827) );
  XNOR2X1 U9359 ( .IN1(n7832), .IN2(n7833), .Q(n6468) );
  XOR2X1 U9360 ( .IN1(n3687), .IN2(n4778), .Q(n7833) );
  XOR2X1 U9361 ( .IN1(n7834), .IN2(n4162), .Q(n7832) );
  XOR2X1 U9362 ( .IN1(WX2020), .IN2(test_so13), .Q(n7834) );
  NOR2X0 U9363 ( .IN1(n7835), .IN2(n7836), .QN(n7825) );
  NOR2X0 U9364 ( .IN1(DFF_374_n1), .IN2(n4288), .QN(n7836) );
  NOR2X0 U9365 ( .IN1(n4296), .IN2(n5345), .QN(n7835) );
  NAND2X0 U9366 ( .IN1(n4811), .IN2(n8693), .QN(n5345) );
  NAND2X0 U9367 ( .IN1(n7837), .IN2(n7838), .QN(WX1953) );
  NOR2X0 U9368 ( .IN1(n7839), .IN2(n7840), .QN(n7838) );
  NOR2X0 U9369 ( .IN1(n4340), .IN2(n7472), .QN(n7840) );
  XNOR2X1 U9370 ( .IN1(n7841), .IN2(n7842), .Q(n7472) );
  XOR2X1 U9371 ( .IN1(n3676), .IN2(n4778), .Q(n7842) );
  XOR2X1 U9372 ( .IN1(WX3311), .IN2(n7843), .Q(n7841) );
  XOR2X1 U9373 ( .IN1(test_so29), .IN2(n9025), .Q(n7843) );
  AND2X1 U9374 ( .IN1(n6476), .IN2(n4264), .Q(n7839) );
  XNOR2X1 U9375 ( .IN1(n7844), .IN2(n7845), .Q(n6476) );
  XOR2X1 U9376 ( .IN1(n3688), .IN2(n4779), .Q(n7845) );
  XOR2X1 U9377 ( .IN1(n7846), .IN2(n4161), .Q(n7844) );
  XOR2X1 U9378 ( .IN1(WX2082), .IN2(n9024), .Q(n7846) );
  NOR2X0 U9379 ( .IN1(n7847), .IN2(n7848), .QN(n7837) );
  NOR2X0 U9380 ( .IN1(DFF_375_n1), .IN2(n4287), .QN(n7848) );
  NOR2X0 U9381 ( .IN1(n4296), .IN2(n5139), .QN(n7847) );
  NAND2X0 U9382 ( .IN1(n4811), .IN2(n8694), .QN(n5139) );
  NAND2X0 U9383 ( .IN1(n7849), .IN2(n7850), .QN(WX1951) );
  NOR2X0 U9384 ( .IN1(n7851), .IN2(n7852), .QN(n7850) );
  NOR2X0 U9385 ( .IN1(n7482), .IN2(n4332), .QN(n7852) );
  XOR2X1 U9386 ( .IN1(n7853), .IN2(n7854), .Q(n7482) );
  XOR2X1 U9387 ( .IN1(n3677), .IN2(n4779), .Q(n7854) );
  XOR2X1 U9388 ( .IN1(n7855), .IN2(n4135), .Q(n7853) );
  XOR2X1 U9389 ( .IN1(WX3373), .IN2(n9027), .Q(n7855) );
  AND2X1 U9390 ( .IN1(n6484), .IN2(n4265), .Q(n7851) );
  XNOR2X1 U9391 ( .IN1(n7856), .IN2(n7857), .Q(n6484) );
  XOR2X1 U9392 ( .IN1(n3689), .IN2(n4779), .Q(n7857) );
  XOR2X1 U9393 ( .IN1(n7858), .IN2(n4160), .Q(n7856) );
  XOR2X1 U9394 ( .IN1(WX2080), .IN2(n9026), .Q(n7858) );
  NOR2X0 U9395 ( .IN1(n7859), .IN2(n7860), .QN(n7849) );
  NOR2X0 U9396 ( .IN1(DFF_376_n1), .IN2(n4287), .QN(n7860) );
  NOR2X0 U9397 ( .IN1(n4296), .IN2(n5150), .QN(n7859) );
  NAND2X0 U9398 ( .IN1(n4811), .IN2(n8695), .QN(n5150) );
  NAND2X0 U9399 ( .IN1(n7861), .IN2(n7862), .QN(WX1949) );
  NOR2X0 U9400 ( .IN1(n7863), .IN2(n7864), .QN(n7862) );
  NOR2X0 U9401 ( .IN1(n7492), .IN2(n4332), .QN(n7864) );
  XOR2X1 U9402 ( .IN1(n7865), .IN2(n7866), .Q(n7492) );
  XOR2X1 U9403 ( .IN1(n3678), .IN2(n4779), .Q(n7866) );
  XOR2X1 U9404 ( .IN1(n7867), .IN2(n4134), .Q(n7865) );
  XOR2X1 U9405 ( .IN1(WX3371), .IN2(n9029), .Q(n7867) );
  AND2X1 U9406 ( .IN1(n6492), .IN2(n4265), .Q(n7863) );
  XNOR2X1 U9407 ( .IN1(n7868), .IN2(n7869), .Q(n6492) );
  XOR2X1 U9408 ( .IN1(n3690), .IN2(n4779), .Q(n7869) );
  XOR2X1 U9409 ( .IN1(n7870), .IN2(n4159), .Q(n7868) );
  XOR2X1 U9410 ( .IN1(WX2078), .IN2(n9028), .Q(n7870) );
  NOR2X0 U9411 ( .IN1(n7871), .IN2(n7872), .QN(n7861) );
  AND2X1 U9412 ( .IN1(n2152), .IN2(test_so21), .Q(n7872) );
  NOR2X0 U9413 ( .IN1(n4296), .IN2(n5161), .QN(n7871) );
  NAND2X0 U9414 ( .IN1(n4811), .IN2(n8696), .QN(n5161) );
  NAND2X0 U9415 ( .IN1(n7873), .IN2(n7874), .QN(WX1947) );
  NOR2X0 U9416 ( .IN1(n7875), .IN2(n7876), .QN(n7874) );
  NOR2X0 U9417 ( .IN1(n4339), .IN2(n7502), .QN(n7876) );
  XNOR2X1 U9418 ( .IN1(n7877), .IN2(n7878), .Q(n7502) );
  XOR2X1 U9419 ( .IN1(n4133), .IN2(n4779), .Q(n7878) );
  XOR2X1 U9420 ( .IN1(n7879), .IN2(n9033), .Q(n7877) );
  XOR2X1 U9421 ( .IN1(n9032), .IN2(n9031), .Q(n7879) );
  AND2X1 U9422 ( .IN1(n6500), .IN2(n4265), .Q(n7875) );
  XNOR2X1 U9423 ( .IN1(n7880), .IN2(n7881), .Q(n6500) );
  XOR2X1 U9424 ( .IN1(n3691), .IN2(n4779), .Q(n7881) );
  XOR2X1 U9425 ( .IN1(n7882), .IN2(n4158), .Q(n7880) );
  XOR2X1 U9426 ( .IN1(WX2076), .IN2(n9030), .Q(n7882) );
  NOR2X0 U9427 ( .IN1(n7883), .IN2(n7884), .QN(n7873) );
  NOR2X0 U9428 ( .IN1(DFF_378_n1), .IN2(n4287), .QN(n7884) );
  NOR2X0 U9429 ( .IN1(n4296), .IN2(n5172), .QN(n7883) );
  NAND2X0 U9430 ( .IN1(test_so11), .IN2(n4828), .QN(n5172) );
  NAND2X0 U9431 ( .IN1(n7885), .IN2(n7886), .QN(WX1945) );
  NOR2X0 U9432 ( .IN1(n7887), .IN2(n7888), .QN(n7886) );
  NOR2X0 U9433 ( .IN1(n7512), .IN2(n4332), .QN(n7888) );
  XOR2X1 U9434 ( .IN1(n7889), .IN2(n7890), .Q(n7512) );
  XOR2X1 U9435 ( .IN1(n3679), .IN2(n4779), .Q(n7890) );
  XOR2X1 U9436 ( .IN1(n7891), .IN2(n4132), .Q(n7889) );
  XOR2X1 U9437 ( .IN1(WX3367), .IN2(n9035), .Q(n7891) );
  AND2X1 U9438 ( .IN1(n6508), .IN2(n4265), .Q(n7887) );
  XNOR2X1 U9439 ( .IN1(n7892), .IN2(n7893), .Q(n6508) );
  XOR2X1 U9440 ( .IN1(n3692), .IN2(n4779), .Q(n7893) );
  XOR2X1 U9441 ( .IN1(n7894), .IN2(n4157), .Q(n7892) );
  XOR2X1 U9442 ( .IN1(WX2074), .IN2(n9034), .Q(n7894) );
  NOR2X0 U9443 ( .IN1(n7895), .IN2(n7896), .QN(n7885) );
  NOR2X0 U9444 ( .IN1(DFF_379_n1), .IN2(n4287), .QN(n7896) );
  NOR2X0 U9445 ( .IN1(n4296), .IN2(n5183), .QN(n7895) );
  NAND2X0 U9446 ( .IN1(n4811), .IN2(n8699), .QN(n5183) );
  NAND2X0 U9447 ( .IN1(n7897), .IN2(n7898), .QN(WX1943) );
  NOR2X0 U9448 ( .IN1(n7899), .IN2(n7900), .QN(n7898) );
  NOR2X0 U9449 ( .IN1(n7522), .IN2(n4332), .QN(n7900) );
  XOR2X1 U9450 ( .IN1(n7901), .IN2(n7902), .Q(n7522) );
  XOR2X1 U9451 ( .IN1(n3680), .IN2(n4779), .Q(n7902) );
  XOR2X1 U9452 ( .IN1(n7903), .IN2(n4131), .Q(n7901) );
  XOR2X1 U9453 ( .IN1(WX3365), .IN2(n9037), .Q(n7903) );
  NOR2X0 U9454 ( .IN1(n4259), .IN2(n6516), .QN(n7899) );
  XNOR2X1 U9455 ( .IN1(n7904), .IN2(n7905), .Q(n6516) );
  XOR2X1 U9456 ( .IN1(n3693), .IN2(n4779), .Q(n7905) );
  XOR2X1 U9457 ( .IN1(WX2008), .IN2(n7906), .Q(n7904) );
  XOR2X1 U9458 ( .IN1(test_so18), .IN2(n9036), .Q(n7906) );
  NOR2X0 U9459 ( .IN1(n7907), .IN2(n7908), .QN(n7897) );
  NOR2X0 U9460 ( .IN1(DFF_380_n1), .IN2(n4287), .QN(n7908) );
  NOR2X0 U9461 ( .IN1(n4296), .IN2(n5194), .QN(n7907) );
  NAND2X0 U9462 ( .IN1(n4811), .IN2(n8700), .QN(n5194) );
  NAND2X0 U9463 ( .IN1(n7909), .IN2(n7910), .QN(WX1941) );
  NOR2X0 U9464 ( .IN1(n7911), .IN2(n7912), .QN(n7910) );
  NOR2X0 U9465 ( .IN1(n7532), .IN2(n4332), .QN(n7912) );
  XOR2X1 U9466 ( .IN1(n7913), .IN2(n7914), .Q(n7532) );
  XOR2X1 U9467 ( .IN1(n3681), .IN2(n4779), .Q(n7914) );
  XOR2X1 U9468 ( .IN1(n7915), .IN2(n4130), .Q(n7913) );
  XOR2X1 U9469 ( .IN1(WX3363), .IN2(n9039), .Q(n7915) );
  AND2X1 U9470 ( .IN1(n6534), .IN2(n4265), .Q(n7911) );
  XNOR2X1 U9471 ( .IN1(n7916), .IN2(n7917), .Q(n6534) );
  XOR2X1 U9472 ( .IN1(n3694), .IN2(n4780), .Q(n7917) );
  XOR2X1 U9473 ( .IN1(n7918), .IN2(n4156), .Q(n7916) );
  XOR2X1 U9474 ( .IN1(WX2070), .IN2(n9038), .Q(n7918) );
  NOR2X0 U9475 ( .IN1(n7919), .IN2(n7920), .QN(n7909) );
  NOR2X0 U9476 ( .IN1(DFF_381_n1), .IN2(n4287), .QN(n7920) );
  NOR2X0 U9477 ( .IN1(n4296), .IN2(n5205), .QN(n7919) );
  NAND2X0 U9478 ( .IN1(n4813), .IN2(n8701), .QN(n5205) );
  NAND2X0 U9479 ( .IN1(n7921), .IN2(n7922), .QN(WX1939) );
  NOR2X0 U9480 ( .IN1(n7923), .IN2(n7924), .QN(n7922) );
  NOR2X0 U9481 ( .IN1(n4339), .IN2(n7542), .QN(n7924) );
  XNOR2X1 U9482 ( .IN1(n7925), .IN2(n7926), .Q(n7542) );
  XOR2X1 U9483 ( .IN1(n4129), .IN2(n4780), .Q(n7926) );
  XOR2X1 U9484 ( .IN1(n7927), .IN2(n9043), .Q(n7925) );
  XOR2X1 U9485 ( .IN1(n9042), .IN2(n9041), .Q(n7927) );
  AND2X1 U9486 ( .IN1(n6553), .IN2(n4265), .Q(n7923) );
  XNOR2X1 U9487 ( .IN1(n7928), .IN2(n7929), .Q(n6553) );
  XOR2X1 U9488 ( .IN1(n3695), .IN2(n4780), .Q(n7929) );
  XOR2X1 U9489 ( .IN1(n7930), .IN2(n4155), .Q(n7928) );
  XOR2X1 U9490 ( .IN1(WX2068), .IN2(n9040), .Q(n7930) );
  NOR2X0 U9491 ( .IN1(n7931), .IN2(n7932), .QN(n7921) );
  NOR2X0 U9492 ( .IN1(DFF_382_n1), .IN2(n4287), .QN(n7932) );
  NOR2X0 U9493 ( .IN1(n4296), .IN2(n5235), .QN(n7931) );
  NAND2X0 U9494 ( .IN1(n4805), .IN2(n8702), .QN(n5235) );
  NAND2X0 U9495 ( .IN1(n7933), .IN2(n7934), .QN(WX1937) );
  NOR2X0 U9496 ( .IN1(n7935), .IN2(n7936), .QN(n7934) );
  NOR2X0 U9497 ( .IN1(n6571), .IN2(n4247), .QN(n7936) );
  XOR2X1 U9498 ( .IN1(n7937), .IN2(n7938), .Q(n6571) );
  XOR2X1 U9499 ( .IN1(n3589), .IN2(n4780), .Q(n7938) );
  XOR2X1 U9500 ( .IN1(n7939), .IN2(n4154), .Q(n7937) );
  XOR2X1 U9501 ( .IN1(WX2066), .IN2(n9045), .Q(n7939) );
  NOR2X0 U9502 ( .IN1(n7552), .IN2(n4327), .QN(n7935) );
  INVX0 U9503 ( .INP(n2153), .ZN(n5369) );
  XOR2X1 U9504 ( .IN1(n7940), .IN2(n7941), .Q(n7552) );
  XOR2X1 U9505 ( .IN1(n3588), .IN2(n4780), .Q(n7941) );
  XOR2X1 U9506 ( .IN1(n7942), .IN2(n4128), .Q(n7940) );
  XOR2X1 U9507 ( .IN1(WX3359), .IN2(n9044), .Q(n7942) );
  NOR2X0 U9508 ( .IN1(n7943), .IN2(n7944), .QN(n7933) );
  NOR2X0 U9509 ( .IN1(n3938), .IN2(n5606), .QN(n7944) );
  NOR2X0 U9510 ( .IN1(DFF_383_n1), .IN2(n4287), .QN(n7943) );
  AND2X1 U9511 ( .IN1(n4801), .IN2(n3938), .Q(WX1839) );
  NOR2X0 U9512 ( .IN1(n4926), .IN2(n7945), .QN(WX1326) );
  XOR2X1 U9513 ( .IN1(n4215), .IN2(DFF_190_n1), .Q(n7945) );
  NOR2X0 U9514 ( .IN1(n4926), .IN2(n7946), .QN(WX1324) );
  XOR2X1 U9515 ( .IN1(n4181), .IN2(DFF_189_n1), .Q(n7946) );
  NOR2X0 U9516 ( .IN1(n4926), .IN2(n7947), .QN(WX1322) );
  XOR2X1 U9517 ( .IN1(n4184), .IN2(DFF_188_n1), .Q(n7947) );
  NOR2X0 U9518 ( .IN1(n4926), .IN2(n7948), .QN(WX1320) );
  XOR2X1 U9519 ( .IN1(n4188), .IN2(DFF_187_n1), .Q(n7948) );
  NOR2X0 U9520 ( .IN1(n4926), .IN2(n7949), .QN(WX1318) );
  XOR2X1 U9521 ( .IN1(n4191), .IN2(DFF_186_n1), .Q(n7949) );
  NOR2X0 U9522 ( .IN1(n4926), .IN2(n7950), .QN(WX1316) );
  XOR2X1 U9523 ( .IN1(n4192), .IN2(DFF_185_n1), .Q(n7950) );
  NOR2X0 U9524 ( .IN1(n4927), .IN2(n7951), .QN(WX1314) );
  XOR2X1 U9525 ( .IN1(n4196), .IN2(DFF_184_n1), .Q(n7951) );
  NOR2X0 U9526 ( .IN1(n4927), .IN2(n7952), .QN(WX1312) );
  XOR2X1 U9527 ( .IN1(n4199), .IN2(DFF_183_n1), .Q(n7952) );
  NOR2X0 U9528 ( .IN1(n4927), .IN2(n7953), .QN(WX1310) );
  XOR2X1 U9529 ( .IN1(n4201), .IN2(DFF_182_n1), .Q(n7953) );
  NOR2X0 U9530 ( .IN1(n4927), .IN2(n7954), .QN(WX1308) );
  XOR2X1 U9531 ( .IN1(n4207), .IN2(DFF_181_n1), .Q(n7954) );
  NOR2X0 U9532 ( .IN1(n4927), .IN2(n7955), .QN(WX1306) );
  XOR2X1 U9533 ( .IN1(n4211), .IN2(DFF_180_n1), .Q(n7955) );
  NOR2X0 U9534 ( .IN1(n4927), .IN2(n7956), .QN(WX1304) );
  XNOR2X1 U9535 ( .IN1(n4213), .IN2(test_so10), .Q(n7956) );
  NOR2X0 U9536 ( .IN1(n4927), .IN2(n7957), .QN(WX1302) );
  XOR2X1 U9537 ( .IN1(n4183), .IN2(DFF_178_n1), .Q(n7957) );
  NOR2X0 U9538 ( .IN1(n4927), .IN2(n7958), .QN(WX1300) );
  XOR2X1 U9539 ( .IN1(n4190), .IN2(DFF_177_n1), .Q(n7958) );
  NOR2X0 U9540 ( .IN1(n4927), .IN2(n7959), .QN(WX1298) );
  XOR2X1 U9541 ( .IN1(n4195), .IN2(DFF_176_n1), .Q(n7959) );
  NOR2X0 U9542 ( .IN1(n4927), .IN2(n7960), .QN(WX1296) );
  XOR2X1 U9543 ( .IN1(DFF_175_n1), .IN2(n7961), .Q(n7960) );
  XOR2X1 U9544 ( .IN1(test_so8), .IN2(DFF_191_n1), .Q(n7961) );
  NOR2X0 U9545 ( .IN1(n4927), .IN2(n7962), .QN(WX1294) );
  XOR2X1 U9546 ( .IN1(n4209), .IN2(DFF_174_n1), .Q(n7962) );
  NOR2X0 U9547 ( .IN1(n4927), .IN2(n7963), .QN(WX1292) );
  XOR2X1 U9548 ( .IN1(n4216), .IN2(DFF_173_n1), .Q(n7963) );
  NOR2X0 U9549 ( .IN1(n4928), .IN2(n7964), .QN(WX1290) );
  XOR2X1 U9550 ( .IN1(n4185), .IN2(DFF_172_n1), .Q(n7964) );
  NOR2X0 U9551 ( .IN1(n4928), .IN2(n7965), .QN(WX1288) );
  XOR2X1 U9552 ( .IN1(n4197), .IN2(DFF_171_n1), .Q(n7965) );
  NOR2X0 U9553 ( .IN1(n4928), .IN2(n7966), .QN(WX1286) );
  XNOR2X1 U9554 ( .IN1(DFF_170_n1), .IN2(n7967), .Q(n7966) );
  XOR2X1 U9555 ( .IN1(n4220), .IN2(DFF_191_n1), .Q(n7967) );
  NOR2X0 U9556 ( .IN1(n4928), .IN2(n7968), .QN(WX1284) );
  XOR2X1 U9557 ( .IN1(n4193), .IN2(DFF_169_n1), .Q(n7968) );
  NOR2X0 U9558 ( .IN1(n4928), .IN2(n7969), .QN(WX1282) );
  XOR2X1 U9559 ( .IN1(n4198), .IN2(DFF_168_n1), .Q(n7969) );
  NOR2X0 U9560 ( .IN1(n4928), .IN2(n7970), .QN(WX1280) );
  XOR2X1 U9561 ( .IN1(n4203), .IN2(DFF_167_n1), .Q(n7970) );
  NOR2X0 U9562 ( .IN1(n4928), .IN2(n7971), .QN(WX1278) );
  XOR2X1 U9563 ( .IN1(n4219), .IN2(DFF_166_n1), .Q(n7971) );
  NOR2X0 U9564 ( .IN1(n4928), .IN2(n7972), .QN(WX1276) );
  XOR2X1 U9565 ( .IN1(n4212), .IN2(DFF_165_n1), .Q(n7972) );
  NOR2X0 U9566 ( .IN1(n4928), .IN2(n7973), .QN(WX1274) );
  XOR2X1 U9567 ( .IN1(n4204), .IN2(DFF_164_n1), .Q(n7973) );
  NOR2X0 U9568 ( .IN1(n4928), .IN2(n7974), .QN(WX1272) );
  XNOR2X1 U9569 ( .IN1(DFF_163_n1), .IN2(n7975), .Q(n7974) );
  XOR2X1 U9570 ( .IN1(n4205), .IN2(DFF_191_n1), .Q(n7975) );
  NOR2X0 U9571 ( .IN1(n4928), .IN2(n7976), .QN(WX1270) );
  XOR2X1 U9572 ( .IN1(n4182), .IN2(DFF_162_n1), .Q(n7976) );
  NOR2X0 U9573 ( .IN1(n4928), .IN2(n7977), .QN(WX1268) );
  XNOR2X1 U9574 ( .IN1(n4217), .IN2(test_so9), .Q(n7977) );
  NOR2X0 U9575 ( .IN1(n4928), .IN2(n7978), .QN(WX1266) );
  XOR2X1 U9576 ( .IN1(n4186), .IN2(DFF_160_n1), .Q(n7978) );
  NOR2X0 U9577 ( .IN1(n4929), .IN2(n7979), .QN(WX1264) );
  XOR2X1 U9578 ( .IN1(n4222), .IN2(DFF_191_n1), .Q(n7979) );
  NOR2X0 U9579 ( .IN1(n4929), .IN2(n7980), .QN(WX11670) );
  XOR2X1 U9580 ( .IN1(n3968), .IN2(DFF_1726_n1), .Q(n7980) );
  NOR2X0 U9581 ( .IN1(n4929), .IN2(n7981), .QN(WX11668) );
  XOR2X1 U9582 ( .IN1(n3969), .IN2(DFF_1725_n1), .Q(n7981) );
  NOR2X0 U9583 ( .IN1(n4929), .IN2(n7982), .QN(WX11666) );
  XOR2X1 U9584 ( .IN1(n3970), .IN2(DFF_1724_n1), .Q(n7982) );
  NOR2X0 U9585 ( .IN1(n4929), .IN2(n7983), .QN(WX11664) );
  XOR2X1 U9586 ( .IN1(n3971), .IN2(DFF_1723_n1), .Q(n7983) );
  NOR2X0 U9587 ( .IN1(n4929), .IN2(n7984), .QN(WX11662) );
  XOR2X1 U9588 ( .IN1(n3972), .IN2(DFF_1722_n1), .Q(n7984) );
  NOR2X0 U9589 ( .IN1(n4929), .IN2(n7985), .QN(WX11660) );
  XOR2X1 U9590 ( .IN1(n3973), .IN2(DFF_1721_n1), .Q(n7985) );
  NOR2X0 U9591 ( .IN1(n4929), .IN2(n7986), .QN(WX11658) );
  XOR2X1 U9592 ( .IN1(n3974), .IN2(DFF_1720_n1), .Q(n7986) );
  NOR2X0 U9593 ( .IN1(n4929), .IN2(n7987), .QN(WX11656) );
  XOR2X1 U9594 ( .IN1(n3975), .IN2(DFF_1719_n1), .Q(n7987) );
  NOR2X0 U9595 ( .IN1(n4929), .IN2(n7988), .QN(WX11654) );
  XOR2X1 U9596 ( .IN1(n3976), .IN2(DFF_1718_n1), .Q(n7988) );
  NOR2X0 U9597 ( .IN1(n4929), .IN2(n7989), .QN(WX11652) );
  XOR2X1 U9598 ( .IN1(n3977), .IN2(DFF_1717_n1), .Q(n7989) );
  NOR2X0 U9599 ( .IN1(n4929), .IN2(n7990), .QN(WX11650) );
  XOR2X1 U9600 ( .IN1(n3978), .IN2(DFF_1716_n1), .Q(n7990) );
  NOR2X0 U9601 ( .IN1(n4929), .IN2(n7991), .QN(WX11648) );
  XOR2X1 U9602 ( .IN1(n3979), .IN2(DFF_1715_n1), .Q(n7991) );
  NOR2X0 U9603 ( .IN1(n4930), .IN2(n7992), .QN(WX11646) );
  XNOR2X1 U9604 ( .IN1(DFF_1714_n1), .IN2(test_so97), .Q(n7992) );
  NOR2X0 U9605 ( .IN1(n4930), .IN2(n7993), .QN(WX11644) );
  XOR2X1 U9606 ( .IN1(n3980), .IN2(DFF_1713_n1), .Q(n7993) );
  NOR2X0 U9607 ( .IN1(n4930), .IN2(n7994), .QN(WX11642) );
  XOR2X1 U9608 ( .IN1(n3981), .IN2(DFF_1712_n1), .Q(n7994) );
  NOR2X0 U9609 ( .IN1(n4930), .IN2(n7995), .QN(WX11640) );
  XOR2X1 U9610 ( .IN1(DFF_1711_n1), .IN2(n7996), .Q(n7995) );
  XOR2X1 U9611 ( .IN1(test_so100), .IN2(n3939), .Q(n7996) );
  NOR2X0 U9612 ( .IN1(n4930), .IN2(n7997), .QN(WX11638) );
  XNOR2X1 U9613 ( .IN1(n3982), .IN2(test_so99), .Q(n7997) );
  NOR2X0 U9614 ( .IN1(n4930), .IN2(n7998), .QN(WX11636) );
  XOR2X1 U9615 ( .IN1(n3983), .IN2(DFF_1709_n1), .Q(n7998) );
  NOR2X0 U9616 ( .IN1(n4930), .IN2(n7999), .QN(WX11634) );
  XOR2X1 U9617 ( .IN1(n3984), .IN2(DFF_1708_n1), .Q(n7999) );
  NOR2X0 U9618 ( .IN1(n4930), .IN2(n8000), .QN(WX11632) );
  XOR2X1 U9619 ( .IN1(n3985), .IN2(DFF_1707_n1), .Q(n8000) );
  NOR2X0 U9620 ( .IN1(n4930), .IN2(n8001), .QN(WX11630) );
  XOR2X1 U9621 ( .IN1(DFF_1706_n1), .IN2(n8002), .Q(n8001) );
  XOR2X1 U9622 ( .IN1(test_so100), .IN2(n3940), .Q(n8002) );
  NOR2X0 U9623 ( .IN1(n4930), .IN2(n8003), .QN(WX11628) );
  XOR2X1 U9624 ( .IN1(n3986), .IN2(DFF_1705_n1), .Q(n8003) );
  NOR2X0 U9625 ( .IN1(n4930), .IN2(n8004), .QN(WX11626) );
  XOR2X1 U9626 ( .IN1(n3987), .IN2(DFF_1704_n1), .Q(n8004) );
  NOR2X0 U9627 ( .IN1(n4930), .IN2(n8005), .QN(WX11624) );
  XOR2X1 U9628 ( .IN1(n3988), .IN2(DFF_1703_n1), .Q(n8005) );
  NOR2X0 U9629 ( .IN1(n4930), .IN2(n8006), .QN(WX11622) );
  XOR2X1 U9630 ( .IN1(n3989), .IN2(DFF_1702_n1), .Q(n8006) );
  NOR2X0 U9631 ( .IN1(n4931), .IN2(n8007), .QN(WX11620) );
  XOR2X1 U9632 ( .IN1(n3990), .IN2(DFF_1701_n1), .Q(n8007) );
  NOR2X0 U9633 ( .IN1(n4931), .IN2(n8008), .QN(WX11618) );
  XOR2X1 U9634 ( .IN1(n3991), .IN2(DFF_1700_n1), .Q(n8008) );
  NOR2X0 U9635 ( .IN1(n4931), .IN2(n8009), .QN(WX11616) );
  XOR2X1 U9636 ( .IN1(DFF_1699_n1), .IN2(n8010), .Q(n8009) );
  XOR2X1 U9637 ( .IN1(test_so100), .IN2(n3941), .Q(n8010) );
  NOR2X0 U9638 ( .IN1(n4931), .IN2(n8011), .QN(WX11614) );
  XOR2X1 U9639 ( .IN1(n3992), .IN2(DFF_1698_n1), .Q(n8011) );
  NOR2X0 U9640 ( .IN1(n4931), .IN2(n8012), .QN(WX11612) );
  XNOR2X1 U9641 ( .IN1(DFF_1697_n1), .IN2(test_so98), .Q(n8012) );
  NOR2X0 U9642 ( .IN1(n4931), .IN2(n8013), .QN(WX11610) );
  XOR2X1 U9643 ( .IN1(n3993), .IN2(DFF_1696_n1), .Q(n8013) );
  NOR2X0 U9644 ( .IN1(n4931), .IN2(n8014), .QN(WX11608) );
  XOR2X1 U9645 ( .IN1(n3960), .IN2(n4245), .Q(n8014) );
  NOR2X0 U9646 ( .IN1(n9062), .IN2(n4854), .QN(WX11082) );
  NOR2X0 U9647 ( .IN1(n9063), .IN2(n4854), .QN(WX11080) );
  NOR2X0 U9648 ( .IN1(n9064), .IN2(n4854), .QN(WX11078) );
  NOR2X0 U9649 ( .IN1(n9065), .IN2(n4854), .QN(WX11076) );
  NOR2X0 U9650 ( .IN1(n9066), .IN2(n4853), .QN(WX11074) );
  NOR2X0 U9651 ( .IN1(n9067), .IN2(n4853), .QN(WX11072) );
  NOR2X0 U9652 ( .IN1(n9070), .IN2(n4853), .QN(WX11070) );
  NOR2X0 U9653 ( .IN1(n9071), .IN2(n4853), .QN(WX11068) );
  NOR2X0 U9654 ( .IN1(n9074), .IN2(n4853), .QN(WX11066) );
  AND2X1 U9655 ( .IN1(n4801), .IN2(test_so91), .Q(WX11064) );
  NOR2X0 U9656 ( .IN1(n9075), .IN2(n4853), .QN(WX11062) );
  NOR2X0 U9657 ( .IN1(n9076), .IN2(n4853), .QN(WX11060) );
  NOR2X0 U9658 ( .IN1(n9077), .IN2(n4853), .QN(WX11058) );
  NOR2X0 U9659 ( .IN1(n9078), .IN2(n4853), .QN(WX11056) );
  NOR2X0 U9660 ( .IN1(n9079), .IN2(n4853), .QN(WX11054) );
  NOR2X0 U9661 ( .IN1(n9080), .IN2(n4853), .QN(WX11052) );
  OR2X1 U9662 ( .IN1(n8015), .IN2(n8016), .Q(WX11050) );
  NAND2X0 U9663 ( .IN1(n8017), .IN2(n8018), .QN(n8016) );
  NAND2X0 U9664 ( .IN1(DATA_0_0), .IN2(n2153), .QN(n8018) );
  OR2X1 U9665 ( .IN1(n4278), .IN2(DFF_1696_n1), .Q(n8017) );
  NAND2X0 U9666 ( .IN1(n8019), .IN2(n8020), .QN(n8015) );
  NAND2X0 U9667 ( .IN1(n4265), .IN2(n5350), .QN(n8020) );
  XNOR2X1 U9668 ( .IN1(n8021), .IN2(n8022), .Q(n5350) );
  XOR2X1 U9669 ( .IN1(n9046), .IN2(n3960), .Q(n8022) );
  XOR2X1 U9670 ( .IN1(WX11051), .IN2(n3697), .Q(n8021) );
  NAND2X0 U9671 ( .IN1(WX10888), .IN2(n4318), .QN(n8019) );
  OR2X1 U9672 ( .IN1(n8023), .IN2(n8024), .Q(WX11048) );
  NAND2X0 U9673 ( .IN1(n8025), .IN2(n8026), .QN(n8024) );
  NAND2X0 U9674 ( .IN1(DATA_0_1), .IN2(n2153), .QN(n8026) );
  OR2X1 U9675 ( .IN1(n4278), .IN2(DFF_1697_n1), .Q(n8025) );
  NAND2X0 U9676 ( .IN1(n8027), .IN2(n8028), .QN(n8023) );
  NAND2X0 U9677 ( .IN1(n4265), .IN2(n5361), .QN(n8028) );
  XNOR2X1 U9678 ( .IN1(n8029), .IN2(n8030), .Q(n5361) );
  XOR2X1 U9679 ( .IN1(n9047), .IN2(n3993), .Q(n8030) );
  XOR2X1 U9680 ( .IN1(WX11049), .IN2(n3699), .Q(n8029) );
  NAND2X0 U9681 ( .IN1(WX10886), .IN2(n4318), .QN(n8027) );
  OR2X1 U9682 ( .IN1(n8031), .IN2(n8032), .Q(WX11046) );
  NAND2X0 U9683 ( .IN1(n8033), .IN2(n8034), .QN(n8032) );
  NAND2X0 U9684 ( .IN1(DATA_0_2), .IN2(n2153), .QN(n8034) );
  OR2X1 U9685 ( .IN1(n4278), .IN2(DFF_1698_n1), .Q(n8033) );
  NAND2X0 U9686 ( .IN1(n8035), .IN2(n8036), .QN(n8031) );
  OR2X1 U9687 ( .IN1(n5370), .IN2(n4246), .Q(n8036) );
  XNOR2X1 U9688 ( .IN1(n8037), .IN2(n8038), .Q(n5370) );
  XOR2X1 U9689 ( .IN1(test_so98), .IN2(n9048), .Q(n8038) );
  XOR2X1 U9690 ( .IN1(WX11047), .IN2(n3701), .Q(n8037) );
  NAND2X0 U9691 ( .IN1(WX10884), .IN2(n4318), .QN(n8035) );
  OR2X1 U9692 ( .IN1(n8039), .IN2(n8040), .Q(WX11044) );
  NAND2X0 U9693 ( .IN1(n8041), .IN2(n8042), .QN(n8040) );
  NAND2X0 U9694 ( .IN1(DATA_0_3), .IN2(n2153), .QN(n8042) );
  OR2X1 U9695 ( .IN1(n4278), .IN2(DFF_1699_n1), .Q(n8041) );
  NAND2X0 U9696 ( .IN1(n8043), .IN2(n8044), .QN(n8039) );
  NAND2X0 U9697 ( .IN1(n4265), .IN2(n5378), .QN(n8044) );
  XNOR2X1 U9698 ( .IN1(n8045), .IN2(n8046), .Q(n5378) );
  XOR2X1 U9699 ( .IN1(n9049), .IN2(n3992), .Q(n8046) );
  XOR2X1 U9700 ( .IN1(WX11045), .IN2(n3703), .Q(n8045) );
  NAND2X0 U9701 ( .IN1(WX10882), .IN2(n4318), .QN(n8043) );
  OR2X1 U9702 ( .IN1(n8047), .IN2(n8048), .Q(WX11042) );
  NAND2X0 U9703 ( .IN1(n8049), .IN2(n8050), .QN(n8048) );
  NAND2X0 U9704 ( .IN1(DATA_0_4), .IN2(n2153), .QN(n8050) );
  OR2X1 U9705 ( .IN1(n4278), .IN2(DFF_1700_n1), .Q(n8049) );
  NAND2X0 U9706 ( .IN1(n8051), .IN2(n8052), .QN(n8047) );
  OR2X1 U9707 ( .IN1(n5386), .IN2(n4246), .Q(n8052) );
  XNOR2X1 U9708 ( .IN1(n8053), .IN2(n8054), .Q(n5386) );
  XOR2X1 U9709 ( .IN1(test_so96), .IN2(n9050), .Q(n8054) );
  XOR2X1 U9710 ( .IN1(WX11043), .IN2(n3941), .Q(n8053) );
  NAND2X0 U9711 ( .IN1(WX10880), .IN2(n4318), .QN(n8051) );
  OR2X1 U9712 ( .IN1(n8055), .IN2(n8056), .Q(WX11040) );
  NAND2X0 U9713 ( .IN1(n8057), .IN2(n8058), .QN(n8056) );
  NAND2X0 U9714 ( .IN1(DATA_0_5), .IN2(n2153), .QN(n8058) );
  OR2X1 U9715 ( .IN1(n4278), .IN2(DFF_1701_n1), .Q(n8057) );
  NAND2X0 U9716 ( .IN1(n8059), .IN2(n8060), .QN(n8055) );
  NAND2X0 U9717 ( .IN1(n4266), .IN2(n5394), .QN(n8060) );
  XNOR2X1 U9718 ( .IN1(n8061), .IN2(n8062), .Q(n5394) );
  XOR2X1 U9719 ( .IN1(n9051), .IN2(n3991), .Q(n8062) );
  XOR2X1 U9720 ( .IN1(WX11041), .IN2(n3706), .Q(n8061) );
  NAND2X0 U9721 ( .IN1(WX10878), .IN2(n4318), .QN(n8059) );
  OR2X1 U9722 ( .IN1(n8063), .IN2(n8064), .Q(WX11038) );
  NAND2X0 U9723 ( .IN1(n8065), .IN2(n8066), .QN(n8064) );
  NAND2X0 U9724 ( .IN1(DATA_0_6), .IN2(n2153), .QN(n8066) );
  OR2X1 U9725 ( .IN1(n4277), .IN2(DFF_1702_n1), .Q(n8065) );
  NAND2X0 U9726 ( .IN1(n8067), .IN2(n8068), .QN(n8063) );
  OR2X1 U9727 ( .IN1(n5402), .IN2(n4246), .Q(n8068) );
  XNOR2X1 U9728 ( .IN1(n8069), .IN2(n8070), .Q(n5402) );
  XOR2X1 U9729 ( .IN1(test_so94), .IN2(n9052), .Q(n8070) );
  XOR2X1 U9730 ( .IN1(WX11039), .IN2(n3990), .Q(n8069) );
  NAND2X0 U9731 ( .IN1(WX10876), .IN2(n4317), .QN(n8067) );
  OR2X1 U9732 ( .IN1(n8071), .IN2(n8072), .Q(WX11036) );
  NAND2X0 U9733 ( .IN1(n8073), .IN2(n8074), .QN(n8072) );
  NAND2X0 U9734 ( .IN1(DATA_0_7), .IN2(n2153), .QN(n8074) );
  OR2X1 U9735 ( .IN1(n4277), .IN2(DFF_1703_n1), .Q(n8073) );
  NAND2X0 U9736 ( .IN1(n8075), .IN2(n8076), .QN(n8071) );
  NAND2X0 U9737 ( .IN1(n4266), .IN2(n5410), .QN(n8076) );
  XNOR2X1 U9738 ( .IN1(n8077), .IN2(n8078), .Q(n5410) );
  XOR2X1 U9739 ( .IN1(n9053), .IN2(n3989), .Q(n8078) );
  XOR2X1 U9740 ( .IN1(WX11037), .IN2(n3709), .Q(n8077) );
  NAND2X0 U9741 ( .IN1(WX10874), .IN2(n4317), .QN(n8075) );
  OR2X1 U9742 ( .IN1(n8079), .IN2(n8080), .Q(WX11034) );
  NAND2X0 U9743 ( .IN1(n8081), .IN2(n8082), .QN(n8080) );
  NAND2X0 U9744 ( .IN1(DATA_0_8), .IN2(n2153), .QN(n8082) );
  OR2X1 U9745 ( .IN1(n4277), .IN2(DFF_1704_n1), .Q(n8081) );
  NAND2X0 U9746 ( .IN1(n8083), .IN2(n8084), .QN(n8079) );
  OR2X1 U9747 ( .IN1(n5418), .IN2(n4246), .Q(n8084) );
  XNOR2X1 U9748 ( .IN1(n8085), .IN2(n8086), .Q(n5418) );
  XOR2X1 U9749 ( .IN1(test_so92), .IN2(n9054), .Q(n8086) );
  XOR2X1 U9750 ( .IN1(WX11163), .IN2(n3988), .Q(n8085) );
  NAND2X0 U9751 ( .IN1(WX10872), .IN2(n4317), .QN(n8083) );
  OR2X1 U9752 ( .IN1(n8087), .IN2(n8088), .Q(WX11032) );
  NAND2X0 U9753 ( .IN1(n8089), .IN2(n8090), .QN(n8088) );
  NAND2X0 U9754 ( .IN1(DATA_0_9), .IN2(n2153), .QN(n8090) );
  OR2X1 U9755 ( .IN1(n4277), .IN2(DFF_1705_n1), .Q(n8089) );
  NAND2X0 U9756 ( .IN1(n8091), .IN2(n8092), .QN(n8087) );
  NAND2X0 U9757 ( .IN1(n4266), .IN2(n5426), .QN(n8092) );
  XNOR2X1 U9758 ( .IN1(n8093), .IN2(n8094), .Q(n5426) );
  XOR2X1 U9759 ( .IN1(n9055), .IN2(n3987), .Q(n8094) );
  XOR2X1 U9760 ( .IN1(WX11033), .IN2(n3712), .Q(n8093) );
  NAND2X0 U9761 ( .IN1(WX10870), .IN2(n4317), .QN(n8091) );
  OR2X1 U9762 ( .IN1(n8095), .IN2(n8096), .Q(WX11030) );
  NAND2X0 U9763 ( .IN1(n8097), .IN2(n8098), .QN(n8096) );
  NAND2X0 U9764 ( .IN1(DATA_0_10), .IN2(n2153), .QN(n8098) );
  OR2X1 U9765 ( .IN1(n4277), .IN2(DFF_1706_n1), .Q(n8097) );
  NAND2X0 U9766 ( .IN1(n8099), .IN2(n8100), .QN(n8095) );
  NAND2X0 U9767 ( .IN1(n4266), .IN2(n5434), .QN(n8100) );
  XNOR2X1 U9768 ( .IN1(n8101), .IN2(n8102), .Q(n5434) );
  XOR2X1 U9769 ( .IN1(n9056), .IN2(n3986), .Q(n8102) );
  XOR2X1 U9770 ( .IN1(WX11031), .IN2(n3714), .Q(n8101) );
  NAND2X0 U9771 ( .IN1(WX10868), .IN2(n4317), .QN(n8099) );
  OR2X1 U9772 ( .IN1(n8103), .IN2(n8104), .Q(WX11028) );
  NAND2X0 U9773 ( .IN1(n8105), .IN2(n8106), .QN(n8104) );
  NAND2X0 U9774 ( .IN1(DATA_0_11), .IN2(n2153), .QN(n8106) );
  OR2X1 U9775 ( .IN1(n4277), .IN2(DFF_1707_n1), .Q(n8105) );
  NAND2X0 U9776 ( .IN1(n8107), .IN2(n8108), .QN(n8103) );
  NAND2X0 U9777 ( .IN1(n4266), .IN2(n5442), .QN(n8108) );
  XNOR2X1 U9778 ( .IN1(n8109), .IN2(n8110), .Q(n5442) );
  XOR2X1 U9779 ( .IN1(n9057), .IN2(n3940), .Q(n8110) );
  XOR2X1 U9780 ( .IN1(WX11029), .IN2(n3716), .Q(n8109) );
  NAND2X0 U9781 ( .IN1(WX10866), .IN2(n4317), .QN(n8107) );
  OR2X1 U9782 ( .IN1(n8111), .IN2(n8112), .Q(WX11026) );
  NAND2X0 U9783 ( .IN1(n8113), .IN2(n8114), .QN(n8112) );
  NAND2X0 U9784 ( .IN1(DATA_0_12), .IN2(n2153), .QN(n8114) );
  OR2X1 U9785 ( .IN1(n4277), .IN2(DFF_1708_n1), .Q(n8113) );
  NAND2X0 U9786 ( .IN1(n8115), .IN2(n8116), .QN(n8111) );
  NAND2X0 U9787 ( .IN1(n4266), .IN2(n5450), .QN(n8116) );
  XNOR2X1 U9788 ( .IN1(n8117), .IN2(n8118), .Q(n5450) );
  XOR2X1 U9789 ( .IN1(n9058), .IN2(n3985), .Q(n8118) );
  XOR2X1 U9790 ( .IN1(WX11027), .IN2(n3718), .Q(n8117) );
  NAND2X0 U9791 ( .IN1(WX10864), .IN2(n4317), .QN(n8115) );
  OR2X1 U9792 ( .IN1(n8119), .IN2(n8120), .Q(WX11024) );
  NAND2X0 U9793 ( .IN1(n8121), .IN2(n8122), .QN(n8120) );
  NAND2X0 U9794 ( .IN1(DATA_0_13), .IN2(n2153), .QN(n8122) );
  OR2X1 U9795 ( .IN1(n4277), .IN2(DFF_1709_n1), .Q(n8121) );
  NAND2X0 U9796 ( .IN1(n8123), .IN2(n8124), .QN(n8119) );
  NAND2X0 U9797 ( .IN1(n4266), .IN2(n5458), .QN(n8124) );
  XNOR2X1 U9798 ( .IN1(n8125), .IN2(n8126), .Q(n5458) );
  XOR2X1 U9799 ( .IN1(n9059), .IN2(n3984), .Q(n8126) );
  XOR2X1 U9800 ( .IN1(WX11025), .IN2(n3720), .Q(n8125) );
  NAND2X0 U9801 ( .IN1(WX10862), .IN2(n4317), .QN(n8123) );
  OR2X1 U9802 ( .IN1(n8127), .IN2(n8128), .Q(WX11022) );
  NAND2X0 U9803 ( .IN1(n8129), .IN2(n8130), .QN(n8128) );
  NAND2X0 U9804 ( .IN1(DATA_0_14), .IN2(n2153), .QN(n8130) );
  NAND2X0 U9805 ( .IN1(test_so99), .IN2(n2152), .QN(n8129) );
  NAND2X0 U9806 ( .IN1(n8131), .IN2(n8132), .QN(n8127) );
  NAND2X0 U9807 ( .IN1(n4266), .IN2(n5466), .QN(n8132) );
  XNOR2X1 U9808 ( .IN1(n8133), .IN2(n8134), .Q(n5466) );
  XOR2X1 U9809 ( .IN1(n9060), .IN2(n3983), .Q(n8134) );
  XOR2X1 U9810 ( .IN1(WX11023), .IN2(n3722), .Q(n8133) );
  NAND2X0 U9811 ( .IN1(WX10860), .IN2(n4317), .QN(n8131) );
  OR2X1 U9812 ( .IN1(n8135), .IN2(n8136), .Q(WX11020) );
  NAND2X0 U9813 ( .IN1(n8137), .IN2(n8138), .QN(n8136) );
  NAND2X0 U9814 ( .IN1(DATA_0_15), .IN2(n2153), .QN(n8138) );
  OR2X1 U9815 ( .IN1(n4277), .IN2(DFF_1711_n1), .Q(n8137) );
  NAND2X0 U9816 ( .IN1(n8139), .IN2(n8140), .QN(n8135) );
  NAND2X0 U9817 ( .IN1(n4267), .IN2(n5474), .QN(n8140) );
  XNOR2X1 U9818 ( .IN1(n8141), .IN2(n8142), .Q(n5474) );
  XOR2X1 U9819 ( .IN1(n9061), .IN2(n3982), .Q(n8142) );
  XOR2X1 U9820 ( .IN1(WX11021), .IN2(n3724), .Q(n8141) );
  NAND2X0 U9821 ( .IN1(WX10858), .IN2(n4317), .QN(n8139) );
  OR2X1 U9822 ( .IN1(n8143), .IN2(n8144), .Q(WX11018) );
  NAND2X0 U9823 ( .IN1(n8145), .IN2(n8146), .QN(n8144) );
  NAND2X0 U9824 ( .IN1(DATA_0_16), .IN2(n2153), .QN(n8146) );
  OR2X1 U9825 ( .IN1(n4277), .IN2(DFF_1712_n1), .Q(n8145) );
  NAND2X0 U9826 ( .IN1(n8147), .IN2(n8148), .QN(n8143) );
  NAND2X0 U9827 ( .IN1(n4267), .IN2(n5482), .QN(n8148) );
  XNOR2X1 U9828 ( .IN1(n8149), .IN2(n8150), .Q(n5482) );
  XOR2X1 U9829 ( .IN1(n3590), .IN2(n4780), .Q(n8150) );
  XOR2X1 U9830 ( .IN1(n8151), .IN2(n3939), .Q(n8149) );
  XOR2X1 U9831 ( .IN1(WX11147), .IN2(n9062), .Q(n8151) );
  NAND2X0 U9832 ( .IN1(WX10856), .IN2(n4316), .QN(n8147) );
  OR2X1 U9833 ( .IN1(n8152), .IN2(n8153), .Q(WX11016) );
  NAND2X0 U9834 ( .IN1(n8154), .IN2(n8155), .QN(n8153) );
  NAND2X0 U9835 ( .IN1(DATA_0_17), .IN2(n2153), .QN(n8155) );
  OR2X1 U9836 ( .IN1(n4277), .IN2(DFF_1713_n1), .Q(n8154) );
  NAND2X0 U9837 ( .IN1(n8156), .IN2(n8157), .QN(n8152) );
  NAND2X0 U9838 ( .IN1(n4267), .IN2(n5490), .QN(n8157) );
  XNOR2X1 U9839 ( .IN1(n8158), .IN2(n8159), .Q(n5490) );
  XOR2X1 U9840 ( .IN1(n3591), .IN2(n4780), .Q(n8159) );
  XOR2X1 U9841 ( .IN1(n8160), .IN2(n3981), .Q(n8158) );
  XOR2X1 U9842 ( .IN1(WX11145), .IN2(n9063), .Q(n8160) );
  NAND2X0 U9843 ( .IN1(WX10854), .IN2(n4316), .QN(n8156) );
  OR2X1 U9844 ( .IN1(n8161), .IN2(n8162), .Q(WX11014) );
  NAND2X0 U9845 ( .IN1(n8163), .IN2(n8164), .QN(n8162) );
  NAND2X0 U9846 ( .IN1(DATA_0_18), .IN2(n2153), .QN(n8164) );
  OR2X1 U9847 ( .IN1(n4277), .IN2(DFF_1714_n1), .Q(n8163) );
  NAND2X0 U9848 ( .IN1(n8165), .IN2(n8166), .QN(n8161) );
  NAND2X0 U9849 ( .IN1(n4267), .IN2(n5498), .QN(n8166) );
  XNOR2X1 U9850 ( .IN1(n8167), .IN2(n8168), .Q(n5498) );
  XOR2X1 U9851 ( .IN1(n3592), .IN2(n4780), .Q(n8168) );
  XOR2X1 U9852 ( .IN1(n8169), .IN2(n3980), .Q(n8167) );
  XOR2X1 U9853 ( .IN1(WX11143), .IN2(n9064), .Q(n8169) );
  NAND2X0 U9854 ( .IN1(WX10852), .IN2(n4316), .QN(n8165) );
  OR2X1 U9855 ( .IN1(n8170), .IN2(n8171), .Q(WX11012) );
  NAND2X0 U9856 ( .IN1(n8172), .IN2(n8173), .QN(n8171) );
  NAND2X0 U9857 ( .IN1(DATA_0_19), .IN2(n2153), .QN(n8173) );
  OR2X1 U9858 ( .IN1(n4276), .IN2(DFF_1715_n1), .Q(n8172) );
  NAND2X0 U9859 ( .IN1(n8174), .IN2(n8175), .QN(n8170) );
  OR2X1 U9860 ( .IN1(n5506), .IN2(n4246), .Q(n8175) );
  XNOR2X1 U9861 ( .IN1(n8176), .IN2(n8177), .Q(n5506) );
  XOR2X1 U9862 ( .IN1(n3593), .IN2(n4780), .Q(n8177) );
  XOR2X1 U9863 ( .IN1(WX11077), .IN2(n8178), .Q(n8176) );
  XOR2X1 U9864 ( .IN1(test_so97), .IN2(n9065), .Q(n8178) );
  NAND2X0 U9865 ( .IN1(WX10850), .IN2(n4316), .QN(n8174) );
  OR2X1 U9866 ( .IN1(n8179), .IN2(n8180), .Q(WX11010) );
  NAND2X0 U9867 ( .IN1(n8181), .IN2(n8182), .QN(n8180) );
  NAND2X0 U9868 ( .IN1(DATA_0_20), .IN2(n2153), .QN(n8182) );
  OR2X1 U9869 ( .IN1(n4276), .IN2(DFF_1716_n1), .Q(n8181) );
  NAND2X0 U9870 ( .IN1(n8183), .IN2(n8184), .QN(n8179) );
  NAND2X0 U9871 ( .IN1(n4267), .IN2(n5514), .QN(n8184) );
  XNOR2X1 U9872 ( .IN1(n8185), .IN2(n8186), .Q(n5514) );
  XOR2X1 U9873 ( .IN1(n3594), .IN2(n4780), .Q(n8186) );
  XOR2X1 U9874 ( .IN1(n8187), .IN2(n3979), .Q(n8185) );
  XOR2X1 U9875 ( .IN1(WX11139), .IN2(n9066), .Q(n8187) );
  NAND2X0 U9876 ( .IN1(WX10848), .IN2(n4316), .QN(n8183) );
  OR2X1 U9877 ( .IN1(n8188), .IN2(n8189), .Q(WX11008) );
  NAND2X0 U9878 ( .IN1(n8190), .IN2(n8191), .QN(n8189) );
  NAND2X0 U9879 ( .IN1(DATA_0_21), .IN2(n2153), .QN(n8191) );
  OR2X1 U9880 ( .IN1(n4276), .IN2(DFF_1717_n1), .Q(n8190) );
  NAND2X0 U9881 ( .IN1(n8192), .IN2(n8193), .QN(n8188) );
  OR2X1 U9882 ( .IN1(n5522), .IN2(n4246), .Q(n8193) );
  XNOR2X1 U9883 ( .IN1(n8194), .IN2(n8195), .Q(n5522) );
  XOR2X1 U9884 ( .IN1(n3978), .IN2(n4780), .Q(n8195) );
  XOR2X1 U9885 ( .IN1(n8196), .IN2(n9069), .Q(n8194) );
  XOR2X1 U9886 ( .IN1(n9068), .IN2(n9067), .Q(n8196) );
  NAND2X0 U9887 ( .IN1(WX10846), .IN2(n4316), .QN(n8192) );
  OR2X1 U9888 ( .IN1(n8197), .IN2(n8198), .Q(WX11006) );
  NAND2X0 U9889 ( .IN1(n8199), .IN2(n8200), .QN(n8198) );
  NAND2X0 U9890 ( .IN1(DATA_0_22), .IN2(n2153), .QN(n8200) );
  OR2X1 U9891 ( .IN1(n4276), .IN2(DFF_1718_n1), .Q(n8199) );
  NAND2X0 U9892 ( .IN1(n8201), .IN2(n8202), .QN(n8197) );
  NAND2X0 U9893 ( .IN1(n4267), .IN2(n5530), .QN(n8202) );
  XNOR2X1 U9894 ( .IN1(n8203), .IN2(n8204), .Q(n5530) );
  XOR2X1 U9895 ( .IN1(n3595), .IN2(n4781), .Q(n8204) );
  XOR2X1 U9896 ( .IN1(n8205), .IN2(n3977), .Q(n8203) );
  XOR2X1 U9897 ( .IN1(WX11135), .IN2(n9070), .Q(n8205) );
  NAND2X0 U9898 ( .IN1(WX10844), .IN2(n4316), .QN(n8201) );
  OR2X1 U9899 ( .IN1(n8206), .IN2(n8207), .Q(WX11004) );
  NAND2X0 U9900 ( .IN1(n8208), .IN2(n8209), .QN(n8207) );
  NAND2X0 U9901 ( .IN1(DATA_0_23), .IN2(n2153), .QN(n8209) );
  OR2X1 U9902 ( .IN1(n4276), .IN2(DFF_1719_n1), .Q(n8208) );
  NAND2X0 U9903 ( .IN1(n8210), .IN2(n8211), .QN(n8206) );
  OR2X1 U9904 ( .IN1(n5538), .IN2(n4246), .Q(n8211) );
  XNOR2X1 U9905 ( .IN1(n8212), .IN2(n8213), .Q(n5538) );
  XOR2X1 U9906 ( .IN1(n3976), .IN2(n4781), .Q(n8213) );
  XOR2X1 U9907 ( .IN1(n8214), .IN2(n9073), .Q(n8212) );
  XOR2X1 U9908 ( .IN1(n9072), .IN2(n9071), .Q(n8214) );
  NAND2X0 U9909 ( .IN1(WX10842), .IN2(n4316), .QN(n8210) );
  OR2X1 U9910 ( .IN1(n8215), .IN2(n8216), .Q(WX11002) );
  NAND2X0 U9911 ( .IN1(n8217), .IN2(n8218), .QN(n8216) );
  NAND2X0 U9912 ( .IN1(DATA_0_24), .IN2(n2153), .QN(n8218) );
  OR2X1 U9913 ( .IN1(n4276), .IN2(DFF_1720_n1), .Q(n8217) );
  NAND2X0 U9914 ( .IN1(n8219), .IN2(n8220), .QN(n8215) );
  NAND2X0 U9915 ( .IN1(n4267), .IN2(n5546), .QN(n8220) );
  XNOR2X1 U9916 ( .IN1(n8221), .IN2(n8222), .Q(n5546) );
  XOR2X1 U9917 ( .IN1(n3596), .IN2(n4780), .Q(n8222) );
  XOR2X1 U9918 ( .IN1(n8223), .IN2(n3975), .Q(n8221) );
  XOR2X1 U9919 ( .IN1(WX11131), .IN2(n9074), .Q(n8223) );
  NAND2X0 U9920 ( .IN1(WX10840), .IN2(n4316), .QN(n8219) );
  OR2X1 U9921 ( .IN1(n8224), .IN2(n8225), .Q(WX11000) );
  NAND2X0 U9922 ( .IN1(n8226), .IN2(n8227), .QN(n8225) );
  NAND2X0 U9923 ( .IN1(DATA_0_25), .IN2(n2153), .QN(n8227) );
  OR2X1 U9924 ( .IN1(n4276), .IN2(DFF_1721_n1), .Q(n8226) );
  NAND2X0 U9925 ( .IN1(n8228), .IN2(n8229), .QN(n8224) );
  OR2X1 U9926 ( .IN1(n5554), .IN2(n4246), .Q(n8229) );
  XNOR2X1 U9927 ( .IN1(n8230), .IN2(n8231), .Q(n5554) );
  XOR2X1 U9928 ( .IN1(n3597), .IN2(n4781), .Q(n8231) );
  XOR2X1 U9929 ( .IN1(n8232), .IN2(n3974), .Q(n8230) );
  XOR2X1 U9930 ( .IN1(WX11065), .IN2(test_so91), .Q(n8232) );
  NAND2X0 U9931 ( .IN1(WX10838), .IN2(n4316), .QN(n8228) );
  OR2X1 U9932 ( .IN1(n8233), .IN2(n8234), .Q(WX10998) );
  NAND2X0 U9933 ( .IN1(n8235), .IN2(n8236), .QN(n8234) );
  NAND2X0 U9934 ( .IN1(DATA_0_26), .IN2(n2153), .QN(n8236) );
  OR2X1 U9935 ( .IN1(n4276), .IN2(DFF_1722_n1), .Q(n8235) );
  NAND2X0 U9936 ( .IN1(n8237), .IN2(n8238), .QN(n8233) );
  NAND2X0 U9937 ( .IN1(n4267), .IN2(n5562), .QN(n8238) );
  XNOR2X1 U9938 ( .IN1(n8239), .IN2(n8240), .Q(n5562) );
  XOR2X1 U9939 ( .IN1(n3598), .IN2(n4781), .Q(n8240) );
  XOR2X1 U9940 ( .IN1(n8241), .IN2(n3973), .Q(n8239) );
  XOR2X1 U9941 ( .IN1(WX11127), .IN2(n9075), .Q(n8241) );
  NAND2X0 U9942 ( .IN1(WX10836), .IN2(n4315), .QN(n8237) );
  OR2X1 U9943 ( .IN1(n8242), .IN2(n8243), .Q(WX10996) );
  NAND2X0 U9944 ( .IN1(n8244), .IN2(n8245), .QN(n8243) );
  NAND2X0 U9945 ( .IN1(DATA_0_27), .IN2(n2153), .QN(n8245) );
  OR2X1 U9946 ( .IN1(n4276), .IN2(DFF_1723_n1), .Q(n8244) );
  NAND2X0 U9947 ( .IN1(n8255), .IN2(n8256), .QN(n8242) );
  NAND2X0 U9948 ( .IN1(n4267), .IN2(n5570), .QN(n8256) );
  XNOR2X1 U9949 ( .IN1(n8273), .IN2(n8274), .Q(n5570) );
  XOR2X1 U9950 ( .IN1(n3599), .IN2(n4781), .Q(n8274) );
  XOR2X1 U9951 ( .IN1(n8291), .IN2(n3972), .Q(n8273) );
  XOR2X1 U9952 ( .IN1(WX11125), .IN2(n9076), .Q(n8291) );
  NAND2X0 U9953 ( .IN1(WX10834), .IN2(n4315), .QN(n8255) );
  OR2X1 U9954 ( .IN1(n8292), .IN2(n8296), .Q(WX10994) );
  NAND2X0 U9955 ( .IN1(n8297), .IN2(n8298), .QN(n8296) );
  NAND2X0 U9956 ( .IN1(DATA_0_28), .IN2(n2153), .QN(n8298) );
  OR2X1 U9957 ( .IN1(n4276), .IN2(DFF_1724_n1), .Q(n8297) );
  NAND2X0 U9958 ( .IN1(n8299), .IN2(n8300), .QN(n8292) );
  NAND2X0 U9959 ( .IN1(n4268), .IN2(n5578), .QN(n8300) );
  XNOR2X1 U9960 ( .IN1(n8301), .IN2(n8302), .Q(n5578) );
  XOR2X1 U9961 ( .IN1(n3600), .IN2(n4781), .Q(n8302) );
  XOR2X1 U9962 ( .IN1(n8303), .IN2(n3971), .Q(n8301) );
  XOR2X1 U9963 ( .IN1(WX11123), .IN2(n9077), .Q(n8303) );
  NAND2X0 U9964 ( .IN1(WX10832), .IN2(n4315), .QN(n8299) );
  OR2X1 U9965 ( .IN1(n8308), .IN2(n8309), .Q(WX10992) );
  NAND2X0 U9966 ( .IN1(n8326), .IN2(n8327), .QN(n8309) );
  NAND2X0 U9967 ( .IN1(DATA_0_29), .IN2(n2153), .QN(n8327) );
  OR2X1 U9968 ( .IN1(n4276), .IN2(DFF_1725_n1), .Q(n8326) );
  NAND2X0 U9969 ( .IN1(n8344), .IN2(n8345), .QN(n8308) );
  NAND2X0 U9970 ( .IN1(n4268), .IN2(n5586), .QN(n8345) );
  XNOR2X1 U9971 ( .IN1(n8354), .IN2(n8355), .Q(n5586) );
  XOR2X1 U9972 ( .IN1(n3601), .IN2(n4781), .Q(n8355) );
  XOR2X1 U9973 ( .IN1(n8356), .IN2(n3970), .Q(n8354) );
  XOR2X1 U9974 ( .IN1(WX11121), .IN2(n9078), .Q(n8356) );
  NAND2X0 U9975 ( .IN1(WX10830), .IN2(n4315), .QN(n8344) );
  OR2X1 U9976 ( .IN1(n8357), .IN2(n8358), .Q(WX10990) );
  NAND2X0 U9977 ( .IN1(n8359), .IN2(n8360), .QN(n8358) );
  NAND2X0 U9978 ( .IN1(DATA_0_30), .IN2(n2153), .QN(n8360) );
  OR2X1 U9979 ( .IN1(n4276), .IN2(DFF_1726_n1), .Q(n8359) );
  NAND2X0 U9980 ( .IN1(n8361), .IN2(n8362), .QN(n8357) );
  NAND2X0 U9981 ( .IN1(n4268), .IN2(n5594), .QN(n8362) );
  XNOR2X1 U9982 ( .IN1(n8379), .IN2(n8380), .Q(n5594) );
  XOR2X1 U9983 ( .IN1(n3602), .IN2(n4781), .Q(n8380) );
  XOR2X1 U9984 ( .IN1(n8397), .IN2(n3969), .Q(n8379) );
  XOR2X1 U9985 ( .IN1(WX11119), .IN2(n9079), .Q(n8397) );
  NAND2X0 U9986 ( .IN1(WX10828), .IN2(n4318), .QN(n8361) );
  NAND2X0 U9987 ( .IN1(n4783), .IN2(TM0), .QN(n5356) );
  NAND2X0 U9988 ( .IN1(n8398), .IN2(n8412), .QN(WX10988) );
  AND2X1 U9989 ( .IN1(n8413), .IN2(n8414), .Q(n8412) );
  NAND2X0 U9990 ( .IN1(n4270), .IN2(n5602), .QN(n8414) );
  XNOR2X1 U9991 ( .IN1(n8415), .IN2(n8416), .Q(n5602) );
  XOR2X1 U9992 ( .IN1(n3582), .IN2(n4781), .Q(n8416) );
  XOR2X1 U9993 ( .IN1(n8417), .IN2(n3968), .Q(n8415) );
  XOR2X1 U9994 ( .IN1(WX11117), .IN2(n9080), .Q(n8417) );
  NAND2X0 U9995 ( .IN1(n8418), .IN2(n4783), .QN(n5352) );
  NOR2X0 U9996 ( .IN1(TM0), .IN2(n4855), .QN(n8418) );
  NAND2X0 U9997 ( .IN1(DATA_0_31), .IN2(n2153), .QN(n8413) );
  NOR2X0 U9998 ( .IN1(n8419), .IN2(n8420), .QN(n8398) );
  NOR2X0 U9999 ( .IN1(n3931), .IN2(n5606), .QN(n8420) );
  INVX0 U10000 ( .INP(n2245), .ZN(n5606) );
  NOR2X0 U10001 ( .IN1(n4295), .IN2(n4245), .QN(n8419) );
  INVX0 U10002 ( .INP(n2152), .ZN(n5355) );
  AND2X1 U10003 ( .IN1(n4801), .IN2(n3931), .Q(WX10890) );
  AND2X1 U10004 ( .IN1(n4802), .IN2(n8263), .Q(WX10888) );
  AND2X1 U10005 ( .IN1(n4802), .IN2(n8264), .Q(WX10886) );
  AND2X1 U10006 ( .IN1(n4801), .IN2(n8265), .Q(WX10884) );
  AND2X1 U10007 ( .IN1(n4802), .IN2(n8266), .Q(WX10882) );
  AND2X1 U10008 ( .IN1(n4802), .IN2(n8267), .Q(WX10880) );
  AND2X1 U10009 ( .IN1(n4802), .IN2(n8268), .Q(WX10878) );
  AND2X1 U10010 ( .IN1(n4802), .IN2(n8269), .Q(WX10876) );
  AND2X1 U10011 ( .IN1(n4802), .IN2(n8270), .Q(WX10874) );
  AND2X1 U10012 ( .IN1(n4802), .IN2(n8271), .Q(WX10872) );
  AND2X1 U10013 ( .IN1(n4803), .IN2(n8272), .Q(WX10870) );
  AND2X1 U10014 ( .IN1(test_so90), .IN2(n4799), .Q(WX10868) );
  AND2X1 U10015 ( .IN1(n4803), .IN2(n8275), .Q(WX10866) );
  AND2X1 U10016 ( .IN1(n4802), .IN2(n8276), .Q(WX10864) );
  AND2X1 U10017 ( .IN1(n4803), .IN2(n8277), .Q(WX10862) );
  AND2X1 U10018 ( .IN1(n4803), .IN2(n8278), .Q(WX10860) );
  AND2X1 U10019 ( .IN1(n4803), .IN2(n8279), .Q(WX10858) );
  AND2X1 U10020 ( .IN1(n4803), .IN2(n8280), .Q(WX10856) );
  AND2X1 U10021 ( .IN1(n4803), .IN2(n8281), .Q(WX10854) );
  AND2X1 U10022 ( .IN1(n4803), .IN2(n8282), .Q(WX10852) );
  AND2X1 U10023 ( .IN1(n4804), .IN2(n8283), .Q(WX10850) );
  AND2X1 U10024 ( .IN1(n4804), .IN2(n8284), .Q(WX10848) );
  AND2X1 U10025 ( .IN1(n4803), .IN2(n8285), .Q(WX10846) );
  AND2X1 U10026 ( .IN1(n4804), .IN2(n8286), .Q(WX10844) );
  AND2X1 U10027 ( .IN1(n4804), .IN2(n8287), .Q(WX10842) );
  AND2X1 U10028 ( .IN1(n4804), .IN2(n8288), .Q(WX10840) );
  AND2X1 U10029 ( .IN1(n4804), .IN2(n8289), .Q(WX10838) );
  AND2X1 U10030 ( .IN1(n4804), .IN2(n8290), .Q(WX10836) );
  AND2X1 U10031 ( .IN1(test_so89), .IN2(n4800), .Q(WX10834) );
  AND2X1 U10032 ( .IN1(n4804), .IN2(n8293), .Q(WX10832) );
  AND2X1 U10033 ( .IN1(n4804), .IN2(n8294), .Q(WX10830) );
  AND2X1 U10034 ( .IN1(n4801), .IN2(n8295), .Q(WX10828) );
  NOR2X0 U10035 ( .IN1(n4931), .IN2(n8432), .QN(WX10377) );
  XNOR2X1 U10036 ( .IN1(DFF_1534_n1), .IN2(test_so85), .Q(n8432) );
  NOR2X0 U10037 ( .IN1(n4931), .IN2(n8433), .QN(WX10375) );
  XOR2X1 U10038 ( .IN1(n3994), .IN2(DFF_1533_n1), .Q(n8433) );
  NOR2X0 U10039 ( .IN1(n4931), .IN2(n8450), .QN(WX10373) );
  XOR2X1 U10040 ( .IN1(n3995), .IN2(DFF_1532_n1), .Q(n8450) );
  NOR2X0 U10041 ( .IN1(n4931), .IN2(n8451), .QN(WX10371) );
  XOR2X1 U10042 ( .IN1(n3996), .IN2(DFF_1531_n1), .Q(n8451) );
  NOR2X0 U10043 ( .IN1(n4931), .IN2(n8468), .QN(WX10369) );
  XOR2X1 U10044 ( .IN1(n3997), .IN2(DFF_1530_n1), .Q(n8468) );
  NOR2X0 U10045 ( .IN1(n4931), .IN2(n8469), .QN(WX10367) );
  XOR2X1 U10046 ( .IN1(n3998), .IN2(DFF_1529_n1), .Q(n8469) );
  NOR2X0 U10047 ( .IN1(n4932), .IN2(n8471), .QN(WX10365) );
  XOR2X1 U10048 ( .IN1(n3999), .IN2(DFF_1528_n1), .Q(n8471) );
  NOR2X0 U10049 ( .IN1(n4932), .IN2(n8472), .QN(WX10363) );
  XOR2X1 U10050 ( .IN1(n4000), .IN2(DFF_1527_n1), .Q(n8472) );
  NOR2X0 U10051 ( .IN1(n4932), .IN2(n8473), .QN(WX10361) );
  XOR2X1 U10052 ( .IN1(n4001), .IN2(DFF_1526_n1), .Q(n8473) );
  NOR2X0 U10053 ( .IN1(n4932), .IN2(n8474), .QN(WX10359) );
  XOR2X1 U10054 ( .IN1(n4002), .IN2(DFF_1525_n1), .Q(n8474) );
  NOR2X0 U10055 ( .IN1(n4932), .IN2(n8475), .QN(WX10357) );
  XOR2X1 U10056 ( .IN1(n4003), .IN2(DFF_1524_n1), .Q(n8475) );
  NOR2X0 U10057 ( .IN1(n4932), .IN2(n8476), .QN(WX10355) );
  XNOR2X1 U10058 ( .IN1(n4004), .IN2(test_so88), .Q(n8476) );
  NOR2X0 U10059 ( .IN1(n4932), .IN2(n8477), .QN(WX10353) );
  XOR2X1 U10060 ( .IN1(n4005), .IN2(DFF_1522_n1), .Q(n8477) );
  NOR2X0 U10061 ( .IN1(n4932), .IN2(n8478), .QN(WX10351) );
  XOR2X1 U10062 ( .IN1(n4006), .IN2(DFF_1521_n1), .Q(n8478) );
  NOR2X0 U10063 ( .IN1(n4932), .IN2(n8485), .QN(WX10349) );
  XOR2X1 U10064 ( .IN1(n4007), .IN2(DFF_1520_n1), .Q(n8485) );
  NOR2X0 U10065 ( .IN1(n4932), .IN2(n8486), .QN(WX10347) );
  XNOR2X1 U10066 ( .IN1(DFF_1519_n1), .IN2(n8503), .Q(n8486) );
  XOR2X1 U10067 ( .IN1(n3942), .IN2(DFF_1535_n1), .Q(n8503) );
  NOR2X0 U10068 ( .IN1(n4932), .IN2(n8504), .QN(WX10345) );
  XOR2X1 U10069 ( .IN1(n4008), .IN2(DFF_1518_n1), .Q(n8504) );
  NOR2X0 U10070 ( .IN1(n4932), .IN2(n8521), .QN(WX10343) );
  XNOR2X1 U10071 ( .IN1(DFF_1517_n1), .IN2(test_so86), .Q(n8521) );
  NOR2X0 U10072 ( .IN1(n4932), .IN2(n8522), .QN(WX10341) );
  XOR2X1 U10073 ( .IN1(n4009), .IN2(DFF_1516_n1), .Q(n8522) );
  NOR2X0 U10074 ( .IN1(n4933), .IN2(n8529), .QN(WX10339) );
  XOR2X1 U10075 ( .IN1(n4010), .IN2(DFF_1515_n1), .Q(n8529) );
  NOR2X0 U10076 ( .IN1(n4933), .IN2(n8530), .QN(WX10337) );
  XNOR2X1 U10077 ( .IN1(DFF_1514_n1), .IN2(n8531), .Q(n8530) );
  XOR2X1 U10078 ( .IN1(n3943), .IN2(DFF_1535_n1), .Q(n8531) );
  NOR2X0 U10079 ( .IN1(n4933), .IN2(n8532), .QN(WX10335) );
  XOR2X1 U10080 ( .IN1(n4011), .IN2(DFF_1513_n1), .Q(n8532) );
  NOR2X0 U10081 ( .IN1(n4933), .IN2(n8533), .QN(WX10333) );
  XOR2X1 U10082 ( .IN1(n4012), .IN2(DFF_1512_n1), .Q(n8533) );
  NOR2X0 U10083 ( .IN1(n4933), .IN2(n8534), .QN(WX10331) );
  XOR2X1 U10084 ( .IN1(n4013), .IN2(DFF_1511_n1), .Q(n8534) );
  NOR2X0 U10085 ( .IN1(n4933), .IN2(n8535), .QN(WX10329) );
  XOR2X1 U10086 ( .IN1(n4014), .IN2(DFF_1510_n1), .Q(n8535) );
  NOR2X0 U10087 ( .IN1(n4933), .IN2(n8536), .QN(WX10327) );
  XOR2X1 U10088 ( .IN1(n4015), .IN2(DFF_1509_n1), .Q(n8536) );
  NOR2X0 U10089 ( .IN1(n4933), .IN2(n8538), .QN(WX10325) );
  XOR2X1 U10090 ( .IN1(n4016), .IN2(DFF_1508_n1), .Q(n8538) );
  NOR2X0 U10091 ( .IN1(n4933), .IN2(n8539), .QN(WX10323) );
  XNOR2X1 U10092 ( .IN1(DFF_1507_n1), .IN2(n8556), .Q(n8539) );
  XOR2X1 U10093 ( .IN1(n3944), .IN2(DFF_1535_n1), .Q(n8556) );
  NOR2X0 U10094 ( .IN1(n4933), .IN2(n8557), .QN(WX10321) );
  XNOR2X1 U10095 ( .IN1(n4017), .IN2(test_so87), .Q(n8557) );
  NOR2X0 U10096 ( .IN1(n4933), .IN2(n8574), .QN(WX10319) );
  XOR2X1 U10097 ( .IN1(n4018), .IN2(DFF_1505_n1), .Q(n8574) );
  NOR2X0 U10098 ( .IN1(n4933), .IN2(n8575), .QN(WX10317) );
  XOR2X1 U10099 ( .IN1(n4019), .IN2(DFF_1504_n1), .Q(n8575) );
  NOR2X0 U10100 ( .IN1(n4933), .IN2(n8587), .QN(WX10315) );
  XOR2X1 U10101 ( .IN1(n3961), .IN2(DFF_1535_n1), .Q(n8587) );
  XNOR2X1 U10102 ( .IN1(n8588), .IN2(n6361), .Q(DATA_9_9) );
  XNOR2X1 U10103 ( .IN1(n8589), .IN2(n8590), .Q(n6361) );
  XOR2X1 U10104 ( .IN1(n3485), .IN2(TM0), .Q(n8590) );
  XOR2X1 U10105 ( .IN1(n8591), .IN2(n4198), .Q(n8589) );
  XOR2X1 U10106 ( .IN1(WX753), .IN2(n9081), .Q(n8591) );
  NAND2X0 U10107 ( .IN1(TM0), .IN2(WX529), .QN(n8588) );
  XNOR2X1 U10108 ( .IN1(n8592), .IN2(n6353), .Q(DATA_9_8) );
  XNOR2X1 U10109 ( .IN1(n8593), .IN2(n8594), .Q(n6353) );
  XOR2X1 U10110 ( .IN1(n3483), .IN2(TM0), .Q(n8594) );
  XOR2X1 U10111 ( .IN1(n8595), .IN2(n4203), .Q(n8593) );
  XOR2X1 U10112 ( .IN1(WX819), .IN2(n9082), .Q(n8595) );
  NAND2X0 U10113 ( .IN1(TM0), .IN2(WX531), .QN(n8592) );
  XNOR2X1 U10114 ( .IN1(n8596), .IN2(n6345), .Q(DATA_9_7) );
  XNOR2X1 U10115 ( .IN1(n8614), .IN2(n8615), .Q(n6345) );
  XOR2X1 U10116 ( .IN1(n3481), .IN2(TM0), .Q(n8615) );
  XOR2X1 U10117 ( .IN1(n8633), .IN2(n4218), .Q(n8614) );
  XOR2X1 U10118 ( .IN1(WX821), .IN2(n4219), .Q(n8633) );
  NAND2X0 U10119 ( .IN1(TM0), .IN2(WX533), .QN(n8596) );
  XOR2X1 U10120 ( .IN1(n8634), .IN2(n6337), .Q(DATA_9_6) );
  XNOR2X1 U10121 ( .IN1(n8645), .IN2(n8646), .Q(n6337) );
  XOR2X1 U10122 ( .IN1(n3479), .IN2(TM0), .Q(n8646) );
  XOR2X1 U10123 ( .IN1(n8647), .IN2(n4212), .Q(n8645) );
  XOR2X1 U10124 ( .IN1(WX823), .IN2(test_so5), .Q(n8647) );
  NAND2X0 U10125 ( .IN1(TM0), .IN2(WX535), .QN(n8634) );
  XNOR2X1 U10126 ( .IN1(n8648), .IN2(n6329), .Q(DATA_9_5) );
  XNOR2X1 U10127 ( .IN1(n8649), .IN2(n8650), .Q(n6329) );
  XOR2X1 U10128 ( .IN1(n3477), .IN2(TM0), .Q(n8650) );
  XOR2X1 U10129 ( .IN1(n8651), .IN2(n4204), .Q(n8649) );
  XOR2X1 U10130 ( .IN1(WX825), .IN2(n9083), .Q(n8651) );
  NAND2X0 U10131 ( .IN1(TM0), .IN2(WX537), .QN(n8648) );
  XNOR2X1 U10132 ( .IN1(n8652), .IN2(n6321), .Q(DATA_9_4) );
  XNOR2X1 U10133 ( .IN1(n8659), .IN2(n8660), .Q(n6321) );
  XOR2X1 U10134 ( .IN1(n3475), .IN2(TM0), .Q(n8660) );
  XOR2X1 U10135 ( .IN1(n8678), .IN2(n4205), .Q(n8659) );
  XOR2X1 U10136 ( .IN1(WX827), .IN2(n9084), .Q(n8678) );
  NAND2X0 U10137 ( .IN1(TM0), .IN2(WX539), .QN(n8652) );
  XOR2X1 U10138 ( .IN1(n8679), .IN2(n6570), .Q(DATA_9_31) );
  XOR2X1 U10139 ( .IN1(n8697), .IN2(n8698), .Q(n6570) );
  XOR2X1 U10140 ( .IN1(n3529), .IN2(n4781), .Q(n8698) );
  XOR2X1 U10141 ( .IN1(n8703), .IN2(n4215), .Q(n8697) );
  XOR2X1 U10142 ( .IN1(WX709), .IN2(n9085), .Q(n8703) );
  NAND2X0 U10143 ( .IN1(TM0), .IN2(WX485), .QN(n8679) );
  XNOR2X1 U10144 ( .IN1(n8704), .IN2(n6550), .Q(DATA_9_30) );
  XNOR2X1 U10145 ( .IN1(n8705), .IN2(n8706), .Q(n6550) );
  XOR2X1 U10146 ( .IN1(n3527), .IN2(n4782), .Q(n8706) );
  XOR2X1 U10147 ( .IN1(n8707), .IN2(n4180), .Q(n8705) );
  XOR2X1 U10148 ( .IN1(WX775), .IN2(n4181), .Q(n8707) );
  NAND2X0 U10149 ( .IN1(TM0), .IN2(WX487), .QN(n8704) );
  XNOR2X1 U10150 ( .IN1(n8708), .IN2(n6313), .Q(DATA_9_3) );
  XNOR2X1 U10151 ( .IN1(n8709), .IN2(n8710), .Q(n6313) );
  XOR2X1 U10152 ( .IN1(n3473), .IN2(TM0), .Q(n8710) );
  XOR2X1 U10153 ( .IN1(n8711), .IN2(n4182), .Q(n8709) );
  XOR2X1 U10154 ( .IN1(WX829), .IN2(n9086), .Q(n8711) );
  NAND2X0 U10155 ( .IN1(TM0), .IN2(WX541), .QN(n8708) );
  XNOR2X1 U10156 ( .IN1(n8712), .IN2(n6531), .Q(DATA_9_29) );
  XNOR2X1 U10157 ( .IN1(n8713), .IN2(n8714), .Q(n6531) );
  XOR2X1 U10158 ( .IN1(n3525), .IN2(n4781), .Q(n8714) );
  XOR2X1 U10159 ( .IN1(n8715), .IN2(n4184), .Q(n8713) );
  XOR2X1 U10160 ( .IN1(WX777), .IN2(n9087), .Q(n8715) );
  NAND2X0 U10161 ( .IN1(TM0), .IN2(WX489), .QN(n8712) );
  XOR2X1 U10162 ( .IN1(n8716), .IN2(n6513), .Q(DATA_9_28) );
  XNOR2X1 U10163 ( .IN1(n8717), .IN2(n8718), .Q(n6513) );
  XOR2X1 U10164 ( .IN1(n4188), .IN2(n4782), .Q(n8718) );
  XOR2X1 U10165 ( .IN1(n8719), .IN2(n4189), .Q(n8717) );
  XOR2X1 U10166 ( .IN1(WX779), .IN2(test_so2), .Q(n8719) );
  NAND2X0 U10167 ( .IN1(TM0), .IN2(WX491), .QN(n8716) );
  XNOR2X1 U10168 ( .IN1(n8720), .IN2(n6505), .Q(DATA_9_27) );
  XNOR2X1 U10169 ( .IN1(n8721), .IN2(n8722), .Q(n6505) );
  XOR2X1 U10170 ( .IN1(n3521), .IN2(n4782), .Q(n8722) );
  XOR2X1 U10171 ( .IN1(n8723), .IN2(n4191), .Q(n8721) );
  XOR2X1 U10172 ( .IN1(WX781), .IN2(n9088), .Q(n8723) );
  NAND2X0 U10173 ( .IN1(TM0), .IN2(WX493), .QN(n8720) );
  XNOR2X1 U10174 ( .IN1(n8724), .IN2(n6497), .Q(DATA_9_26) );
  XNOR2X1 U10175 ( .IN1(n8725), .IN2(n8726), .Q(n6497) );
  XOR2X1 U10176 ( .IN1(n3519), .IN2(n4782), .Q(n8726) );
  XOR2X1 U10177 ( .IN1(n8727), .IN2(n4192), .Q(n8725) );
  XOR2X1 U10178 ( .IN1(WX783), .IN2(n9089), .Q(n8727) );
  NAND2X0 U10179 ( .IN1(TM0), .IN2(WX495), .QN(n8724) );
  XNOR2X1 U10180 ( .IN1(n8728), .IN2(n6489), .Q(DATA_9_25) );
  XNOR2X1 U10181 ( .IN1(n8729), .IN2(n8730), .Q(n6489) );
  XOR2X1 U10182 ( .IN1(n3517), .IN2(n4782), .Q(n8730) );
  XOR2X1 U10183 ( .IN1(n8731), .IN2(n4196), .Q(n8729) );
  XOR2X1 U10184 ( .IN1(WX785), .IN2(n9090), .Q(n8731) );
  NAND2X0 U10185 ( .IN1(TM0), .IN2(WX497), .QN(n8728) );
  XOR2X1 U10186 ( .IN1(n8732), .IN2(n6481), .Q(DATA_9_24) );
  XNOR2X1 U10187 ( .IN1(n8733), .IN2(n8734), .Q(n6481) );
  XOR2X1 U10188 ( .IN1(n3515), .IN2(n4782), .Q(n8734) );
  XOR2X1 U10189 ( .IN1(n8735), .IN2(n4199), .Q(n8733) );
  XOR2X1 U10190 ( .IN1(WX787), .IN2(test_so4), .Q(n8735) );
  NAND2X0 U10191 ( .IN1(TM0), .IN2(WX499), .QN(n8732) );
  XNOR2X1 U10192 ( .IN1(n8736), .IN2(n6473), .Q(DATA_9_23) );
  XNOR2X1 U10193 ( .IN1(n8737), .IN2(n8738), .Q(n6473) );
  XOR2X1 U10194 ( .IN1(n3513), .IN2(n4782), .Q(n8738) );
  XOR2X1 U10195 ( .IN1(n8739), .IN2(n4201), .Q(n8737) );
  XOR2X1 U10196 ( .IN1(WX789), .IN2(n9091), .Q(n8739) );
  NAND2X0 U10197 ( .IN1(TM0), .IN2(WX501), .QN(n8736) );
  XNOR2X1 U10198 ( .IN1(n8740), .IN2(n6465), .Q(DATA_9_22) );
  XNOR2X1 U10199 ( .IN1(n8741), .IN2(n8742), .Q(n6465) );
  XOR2X1 U10200 ( .IN1(n3511), .IN2(n4782), .Q(n8742) );
  XOR2X1 U10201 ( .IN1(n8743), .IN2(n4206), .Q(n8741) );
  XOR2X1 U10202 ( .IN1(WX791), .IN2(n4207), .Q(n8743) );
  NAND2X0 U10203 ( .IN1(TM0), .IN2(WX503), .QN(n8740) );
  XNOR2X1 U10204 ( .IN1(n8744), .IN2(n6457), .Q(DATA_9_21) );
  XNOR2X1 U10205 ( .IN1(n8745), .IN2(n8746), .Q(n6457) );
  XOR2X1 U10206 ( .IN1(n3509), .IN2(n4782), .Q(n8746) );
  XOR2X1 U10207 ( .IN1(n8747), .IN2(n4210), .Q(n8745) );
  XOR2X1 U10208 ( .IN1(WX793), .IN2(n4211), .Q(n8747) );
  NAND2X0 U10209 ( .IN1(TM0), .IN2(WX505), .QN(n8744) );
  XOR2X1 U10210 ( .IN1(n8748), .IN2(n6449), .Q(DATA_9_20) );
  XNOR2X1 U10211 ( .IN1(n8749), .IN2(n8750), .Q(n6449) );
  XOR2X1 U10212 ( .IN1(n3507), .IN2(n4782), .Q(n8750) );
  XOR2X1 U10213 ( .IN1(n8751), .IN2(n4213), .Q(n8749) );
  XOR2X1 U10214 ( .IN1(WX731), .IN2(test_so6), .Q(n8751) );
  NAND2X0 U10215 ( .IN1(TM0), .IN2(WX507), .QN(n8748) );
  XOR2X1 U10216 ( .IN1(n8752), .IN2(n6305), .Q(DATA_9_2) );
  XNOR2X1 U10217 ( .IN1(n8753), .IN2(n8754), .Q(n6305) );
  XOR2X1 U10218 ( .IN1(n3471), .IN2(TM0), .Q(n8754) );
  XOR2X1 U10219 ( .IN1(n8755), .IN2(n4217), .Q(n8753) );
  XOR2X1 U10220 ( .IN1(WX767), .IN2(test_so7), .Q(n8755) );
  NAND2X0 U10221 ( .IN1(TM0), .IN2(WX543), .QN(n8752) );
  XNOR2X1 U10222 ( .IN1(n8756), .IN2(n6441), .Q(DATA_9_19) );
  XNOR2X1 U10223 ( .IN1(n8757), .IN2(n8758), .Q(n6441) );
  XOR2X1 U10224 ( .IN1(n3505), .IN2(n4782), .Q(n8758) );
  XOR2X1 U10225 ( .IN1(n8759), .IN2(n4183), .Q(n8757) );
  XOR2X1 U10226 ( .IN1(WX797), .IN2(n9092), .Q(n8759) );
  NAND2X0 U10227 ( .IN1(TM0), .IN2(WX509), .QN(n8756) );
  XNOR2X1 U10228 ( .IN1(n8760), .IN2(n6433), .Q(DATA_9_18) );
  XNOR2X1 U10229 ( .IN1(n8761), .IN2(n8762), .Q(n6433) );
  XOR2X1 U10230 ( .IN1(n3503), .IN2(n4782), .Q(n8762) );
  XOR2X1 U10231 ( .IN1(n8763), .IN2(n4190), .Q(n8761) );
  XOR2X1 U10232 ( .IN1(WX799), .IN2(n9093), .Q(n8763) );
  NAND2X0 U10233 ( .IN1(TM0), .IN2(WX511), .QN(n8760) );
  XNOR2X1 U10234 ( .IN1(n8764), .IN2(n6425), .Q(DATA_9_17) );
  XNOR2X1 U10235 ( .IN1(n8765), .IN2(n8766), .Q(n6425) );
  XOR2X1 U10236 ( .IN1(n3501), .IN2(n4781), .Q(n8766) );
  XOR2X1 U10237 ( .IN1(n8767), .IN2(n4195), .Q(n8765) );
  XOR2X1 U10238 ( .IN1(WX801), .IN2(n9094), .Q(n8767) );
  NAND2X0 U10239 ( .IN1(TM0), .IN2(WX513), .QN(n8764) );
  XOR2X1 U10240 ( .IN1(n8768), .IN2(n6417), .Q(DATA_9_16) );
  XNOR2X1 U10241 ( .IN1(n8769), .IN2(n8770), .Q(n6417) );
  XOR2X1 U10242 ( .IN1(n3499), .IN2(n4771), .Q(n8770) );
  XOR2X1 U10243 ( .IN1(n8771), .IN2(n4202), .Q(n8769) );
  XOR2X1 U10244 ( .IN1(WX739), .IN2(test_so8), .Q(n8771) );
  NAND2X0 U10245 ( .IN1(TM0), .IN2(WX515), .QN(n8768) );
  XNOR2X1 U10246 ( .IN1(n8772), .IN2(n6409), .Q(DATA_9_15) );
  XNOR2X1 U10247 ( .IN1(n8773), .IN2(n8774), .Q(n6409) );
  XOR2X1 U10248 ( .IN1(n3497), .IN2(TM0), .Q(n8774) );
  XOR2X1 U10249 ( .IN1(n8775), .IN2(n4208), .Q(n8773) );
  XOR2X1 U10250 ( .IN1(WX805), .IN2(n4209), .Q(n8775) );
  NAND2X0 U10251 ( .IN1(TM0), .IN2(WX517), .QN(n8772) );
  XNOR2X1 U10252 ( .IN1(n8776), .IN2(n6401), .Q(DATA_9_14) );
  XNOR2X1 U10253 ( .IN1(n8777), .IN2(n8778), .Q(n6401) );
  XOR2X1 U10254 ( .IN1(n3495), .IN2(TM0), .Q(n8778) );
  XOR2X1 U10255 ( .IN1(n8779), .IN2(n4216), .Q(n8777) );
  XOR2X1 U10256 ( .IN1(WX807), .IN2(n9095), .Q(n8779) );
  NAND2X0 U10257 ( .IN1(test_so1), .IN2(TM0), .QN(n8776) );
  XNOR2X1 U10258 ( .IN1(n8780), .IN2(n6393), .Q(DATA_9_13) );
  XNOR2X1 U10259 ( .IN1(n8781), .IN2(n8782), .Q(n6393) );
  XOR2X1 U10260 ( .IN1(n3493), .IN2(TM0), .Q(n8782) );
  XOR2X1 U10261 ( .IN1(n8783), .IN2(n4185), .Q(n8781) );
  XOR2X1 U10262 ( .IN1(WX809), .IN2(n9096), .Q(n8783) );
  NAND2X0 U10263 ( .IN1(TM0), .IN2(WX521), .QN(n8780) );
  XNOR2X1 U10264 ( .IN1(n8784), .IN2(n6385), .Q(DATA_9_12) );
  XNOR2X1 U10265 ( .IN1(n8785), .IN2(n8786), .Q(n6385) );
  XOR2X1 U10266 ( .IN1(n3491), .IN2(TM0), .Q(n8786) );
  XOR2X1 U10267 ( .IN1(n8787), .IN2(n4197), .Q(n8785) );
  XOR2X1 U10268 ( .IN1(WX811), .IN2(n9097), .Q(n8787) );
  NAND2X0 U10269 ( .IN1(TM0), .IN2(WX523), .QN(n8784) );
  XNOR2X1 U10270 ( .IN1(n8788), .IN2(n6377), .Q(DATA_9_11) );
  XNOR2X1 U10271 ( .IN1(n8789), .IN2(n8790), .Q(n6377) );
  XOR2X1 U10272 ( .IN1(n3489), .IN2(TM0), .Q(n8790) );
  XOR2X1 U10273 ( .IN1(n8791), .IN2(n4220), .Q(n8789) );
  XOR2X1 U10274 ( .IN1(WX813), .IN2(n9098), .Q(n8791) );
  NAND2X0 U10275 ( .IN1(TM0), .IN2(WX525), .QN(n8788) );
  XOR2X1 U10276 ( .IN1(n8792), .IN2(n6369), .Q(DATA_9_10) );
  XNOR2X1 U10277 ( .IN1(n8793), .IN2(n8794), .Q(n6369) );
  XOR2X1 U10278 ( .IN1(n4193), .IN2(TM0), .Q(n8794) );
  XOR2X1 U10279 ( .IN1(n8795), .IN2(n4194), .Q(n8793) );
  XOR2X1 U10280 ( .IN1(WX815), .IN2(test_so3), .Q(n8795) );
  NAND2X0 U10281 ( .IN1(TM0), .IN2(WX527), .QN(n8792) );
  XNOR2X1 U10282 ( .IN1(n8796), .IN2(n6297), .Q(DATA_9_1) );
  XNOR2X1 U10283 ( .IN1(n8797), .IN2(n8798), .Q(n6297) );
  XOR2X1 U10284 ( .IN1(n3469), .IN2(TM0), .Q(n8798) );
  XOR2X1 U10285 ( .IN1(n8799), .IN2(n4186), .Q(n8797) );
  XOR2X1 U10286 ( .IN1(WX833), .IN2(n9099), .Q(n8799) );
  NAND2X0 U10287 ( .IN1(TM0), .IN2(WX545), .QN(n8796) );
  XNOR2X1 U10288 ( .IN1(n8800), .IN2(n6289), .Q(DATA_9_0) );
  XNOR2X1 U10289 ( .IN1(n8801), .IN2(n8802), .Q(n6289) );
  XOR2X1 U10290 ( .IN1(n3467), .IN2(TM0), .Q(n8802) );
  XOR2X1 U10291 ( .IN1(n8803), .IN2(n4221), .Q(n8801) );
  XOR2X1 U10292 ( .IN1(WX835), .IN2(n4222), .Q(n8803) );
  NAND2X0 U10293 ( .IN1(TM0), .IN2(WX547), .QN(n8800) );
  NOR2X0 U3558_U2 ( .IN1(n4900), .IN2(U3558_n1), .QN(n2245) );
  INVX0 U3558_U1 ( .INP(n4313), .ZN(U3558_n1) );
  INVX0 U3871_U2 ( .INP(n3278), .ZN(U3871_n1) );
  NOR2X1 U3871_U1 ( .IN1(TM0), .IN2(U3871_n1), .QN(n2153) );
  INVX0 U3991_U2 ( .INP(n3278), .ZN(U3991_n1) );
  NOR2X0 U3991_U1 ( .IN1(n225), .IN2(U3991_n1), .QN(n2152) );
  INVX0 U5716_U2 ( .INP(WX547), .ZN(U5716_n1) );
  NOR2X0 U5716_U1 ( .IN1(n4883), .IN2(U5716_n1), .QN(WX544) );
  INVX0 U5717_U2 ( .INP(WX545), .ZN(U5717_n1) );
  NOR2X0 U5717_U1 ( .IN1(n4901), .IN2(U5717_n1), .QN(WX542) );
  INVX0 U5718_U2 ( .INP(WX543), .ZN(U5718_n1) );
  NOR2X0 U5718_U1 ( .IN1(n4901), .IN2(U5718_n1), .QN(WX540) );
  INVX0 U5719_U2 ( .INP(WX541), .ZN(U5719_n1) );
  NOR2X0 U5719_U1 ( .IN1(n4901), .IN2(U5719_n1), .QN(WX538) );
  INVX0 U5720_U2 ( .INP(WX539), .ZN(U5720_n1) );
  NOR2X0 U5720_U1 ( .IN1(n4901), .IN2(U5720_n1), .QN(WX536) );
  INVX0 U5721_U2 ( .INP(WX537), .ZN(U5721_n1) );
  NOR2X0 U5721_U1 ( .IN1(n4901), .IN2(U5721_n1), .QN(WX534) );
  INVX0 U5722_U2 ( .INP(WX535), .ZN(U5722_n1) );
  NOR2X0 U5722_U1 ( .IN1(n4901), .IN2(U5722_n1), .QN(WX532) );
  INVX0 U5723_U2 ( .INP(WX533), .ZN(U5723_n1) );
  NOR2X0 U5723_U1 ( .IN1(n4901), .IN2(U5723_n1), .QN(WX530) );
  INVX0 U5724_U2 ( .INP(WX531), .ZN(U5724_n1) );
  NOR2X0 U5724_U1 ( .IN1(n4901), .IN2(U5724_n1), .QN(WX528) );
  INVX0 U5725_U2 ( .INP(WX529), .ZN(U5725_n1) );
  NOR2X0 U5725_U1 ( .IN1(n4901), .IN2(U5725_n1), .QN(WX526) );
  INVX0 U5726_U2 ( .INP(WX527), .ZN(U5726_n1) );
  NOR2X0 U5726_U1 ( .IN1(n4901), .IN2(U5726_n1), .QN(WX524) );
  INVX0 U5727_U2 ( .INP(WX525), .ZN(U5727_n1) );
  NOR2X0 U5727_U1 ( .IN1(n4900), .IN2(U5727_n1), .QN(WX522) );
  INVX0 U5728_U2 ( .INP(WX523), .ZN(U5728_n1) );
  NOR2X0 U5728_U1 ( .IN1(n4900), .IN2(U5728_n1), .QN(WX520) );
  INVX0 U5729_U2 ( .INP(WX521), .ZN(U5729_n1) );
  NOR2X0 U5729_U1 ( .IN1(n4900), .IN2(U5729_n1), .QN(WX518) );
  INVX0 U5730_U2 ( .INP(test_so1), .ZN(U5730_n1) );
  NOR2X0 U5730_U1 ( .IN1(n4900), .IN2(U5730_n1), .QN(WX516) );
  INVX0 U5731_U2 ( .INP(WX517), .ZN(U5731_n1) );
  NOR2X0 U5731_U1 ( .IN1(n4900), .IN2(U5731_n1), .QN(WX514) );
  INVX0 U5732_U2 ( .INP(WX515), .ZN(U5732_n1) );
  NOR2X0 U5732_U1 ( .IN1(n4900), .IN2(U5732_n1), .QN(WX512) );
  INVX0 U5733_U2 ( .INP(WX513), .ZN(U5733_n1) );
  NOR2X0 U5733_U1 ( .IN1(n4897), .IN2(U5733_n1), .QN(WX510) );
  INVX0 U5734_U2 ( .INP(WX511), .ZN(U5734_n1) );
  NOR2X0 U5734_U1 ( .IN1(n4897), .IN2(U5734_n1), .QN(WX508) );
  INVX0 U5735_U2 ( .INP(WX509), .ZN(U5735_n1) );
  NOR2X0 U5735_U1 ( .IN1(n4897), .IN2(U5735_n1), .QN(WX506) );
  INVX0 U5736_U2 ( .INP(WX507), .ZN(U5736_n1) );
  NOR2X0 U5736_U1 ( .IN1(n4897), .IN2(U5736_n1), .QN(WX504) );
  INVX0 U5737_U2 ( .INP(WX505), .ZN(U5737_n1) );
  NOR2X0 U5737_U1 ( .IN1(n4897), .IN2(U5737_n1), .QN(WX502) );
  INVX0 U5738_U2 ( .INP(WX503), .ZN(U5738_n1) );
  NOR2X0 U5738_U1 ( .IN1(n4897), .IN2(U5738_n1), .QN(WX500) );
  INVX0 U5739_U2 ( .INP(WX501), .ZN(U5739_n1) );
  NOR2X0 U5739_U1 ( .IN1(n4897), .IN2(U5739_n1), .QN(WX498) );
  INVX0 U5740_U2 ( .INP(WX499), .ZN(U5740_n1) );
  NOR2X0 U5740_U1 ( .IN1(n4896), .IN2(U5740_n1), .QN(WX496) );
  INVX0 U5741_U2 ( .INP(WX497), .ZN(U5741_n1) );
  NOR2X0 U5741_U1 ( .IN1(n4896), .IN2(U5741_n1), .QN(WX494) );
  INVX0 U5742_U2 ( .INP(WX495), .ZN(U5742_n1) );
  NOR2X0 U5742_U1 ( .IN1(n4896), .IN2(U5742_n1), .QN(WX492) );
  INVX0 U5743_U2 ( .INP(WX493), .ZN(U5743_n1) );
  NOR2X0 U5743_U1 ( .IN1(n4896), .IN2(U5743_n1), .QN(WX490) );
  INVX0 U5744_U2 ( .INP(WX491), .ZN(U5744_n1) );
  NOR2X0 U5744_U1 ( .IN1(n4896), .IN2(U5744_n1), .QN(WX488) );
  INVX0 U5745_U2 ( .INP(WX489), .ZN(U5745_n1) );
  NOR2X0 U5745_U1 ( .IN1(n4896), .IN2(U5745_n1), .QN(WX486) );
  INVX0 U5746_U2 ( .INP(WX487), .ZN(U5746_n1) );
  NOR2X0 U5746_U1 ( .IN1(n4896), .IN2(U5746_n1), .QN(WX484) );
  INVX0 U5747_U2 ( .INP(WX5939), .ZN(U5747_n1) );
  NOR2X0 U5747_U1 ( .IN1(n4896), .IN2(U5747_n1), .QN(WX6002) );
  INVX0 U5748_U2 ( .INP(test_so49), .ZN(U5748_n1) );
  NOR2X0 U5748_U1 ( .IN1(n4894), .IN2(U5748_n1), .QN(WX6000) );
  INVX0 U5749_U2 ( .INP(WX5935), .ZN(U5749_n1) );
  NOR2X0 U5749_U1 ( .IN1(n4894), .IN2(U5749_n1), .QN(WX5998) );
  INVX0 U5750_U2 ( .INP(WX5933), .ZN(U5750_n1) );
  NOR2X0 U5750_U1 ( .IN1(n4903), .IN2(U5750_n1), .QN(WX5996) );
  INVX0 U5751_U2 ( .INP(WX5931), .ZN(U5751_n1) );
  NOR2X0 U5751_U1 ( .IN1(n4898), .IN2(U5751_n1), .QN(WX5994) );
  INVX0 U5752_U2 ( .INP(WX3269), .ZN(U5752_n1) );
  NOR2X0 U5752_U1 ( .IN1(n4893), .IN2(U5752_n1), .QN(WX3332) );
  INVX0 U5753_U2 ( .INP(WX3265), .ZN(U5753_n1) );
  NOR2X0 U5753_U1 ( .IN1(n4893), .IN2(U5753_n1), .QN(WX3328) );
  INVX0 U5754_U2 ( .INP(WX3263), .ZN(U5754_n1) );
  NOR2X0 U5754_U1 ( .IN1(n4893), .IN2(U5754_n1), .QN(WX3326) );
  INVX0 U5755_U2 ( .INP(WX11179), .ZN(U5755_n1) );
  NOR2X0 U5755_U1 ( .IN1(n4894), .IN2(U5755_n1), .QN(WX11242) );
  INVX0 U5756_U2 ( .INP(WX11177), .ZN(U5756_n1) );
  NOR2X0 U5756_U1 ( .IN1(n4894), .IN2(U5756_n1), .QN(WX11240) );
  INVX0 U5757_U2 ( .INP(WX11175), .ZN(U5757_n1) );
  NOR2X0 U5757_U1 ( .IN1(n4894), .IN2(U5757_n1), .QN(WX11238) );
  INVX0 U5758_U2 ( .INP(WX11173), .ZN(U5758_n1) );
  NOR2X0 U5758_U1 ( .IN1(n4894), .IN2(U5758_n1), .QN(WX11236) );
  INVX0 U5759_U2 ( .INP(test_so96), .ZN(U5759_n1) );
  NOR2X0 U5759_U1 ( .IN1(n4894), .IN2(U5759_n1), .QN(WX11234) );
  INVX0 U5760_U2 ( .INP(WX11169), .ZN(U5760_n1) );
  NOR2X0 U5760_U1 ( .IN1(n4894), .IN2(U5760_n1), .QN(WX11232) );
  INVX0 U5761_U2 ( .INP(WX11167), .ZN(U5761_n1) );
  NOR2X0 U5761_U1 ( .IN1(n4894), .IN2(U5761_n1), .QN(WX11230) );
  INVX0 U5762_U2 ( .INP(WX11165), .ZN(U5762_n1) );
  NOR2X0 U5762_U1 ( .IN1(n4894), .IN2(U5762_n1), .QN(WX11228) );
  INVX0 U5763_U2 ( .INP(WX11163), .ZN(U5763_n1) );
  NOR2X0 U5763_U1 ( .IN1(n4894), .IN2(U5763_n1), .QN(WX11226) );
  INVX0 U5764_U2 ( .INP(WX11161), .ZN(U5764_n1) );
  NOR2X0 U5764_U1 ( .IN1(n4895), .IN2(U5764_n1), .QN(WX11224) );
  INVX0 U5765_U2 ( .INP(WX11159), .ZN(U5765_n1) );
  NOR2X0 U5765_U1 ( .IN1(n4895), .IN2(U5765_n1), .QN(WX11222) );
  INVX0 U5766_U2 ( .INP(WX11157), .ZN(U5766_n1) );
  NOR2X0 U5766_U1 ( .IN1(n4895), .IN2(U5766_n1), .QN(WX11220) );
  INVX0 U5767_U2 ( .INP(WX11155), .ZN(U5767_n1) );
  NOR2X0 U5767_U1 ( .IN1(n4895), .IN2(U5767_n1), .QN(WX11218) );
  INVX0 U5768_U2 ( .INP(WX11153), .ZN(U5768_n1) );
  NOR2X0 U5768_U1 ( .IN1(n4895), .IN2(U5768_n1), .QN(WX11216) );
  INVX0 U5769_U2 ( .INP(WX11151), .ZN(U5769_n1) );
  NOR2X0 U5769_U1 ( .IN1(n4895), .IN2(U5769_n1), .QN(WX11214) );
  INVX0 U5770_U2 ( .INP(WX11149), .ZN(U5770_n1) );
  NOR2X0 U5770_U1 ( .IN1(n4895), .IN2(U5770_n1), .QN(WX11212) );
  INVX0 U5771_U2 ( .INP(WX11147), .ZN(U5771_n1) );
  NOR2X0 U5771_U1 ( .IN1(n4895), .IN2(U5771_n1), .QN(WX11210) );
  INVX0 U5772_U2 ( .INP(WX11145), .ZN(U5772_n1) );
  NOR2X0 U5772_U1 ( .IN1(n4895), .IN2(U5772_n1), .QN(WX11208) );
  INVX0 U5773_U2 ( .INP(WX11143), .ZN(U5773_n1) );
  NOR2X0 U5773_U1 ( .IN1(n4895), .IN2(U5773_n1), .QN(WX11206) );
  INVX0 U5774_U2 ( .INP(WX11141), .ZN(U5774_n1) );
  NOR2X0 U5774_U1 ( .IN1(n4895), .IN2(U5774_n1), .QN(WX11204) );
  INVX0 U5775_U2 ( .INP(WX11139), .ZN(U5775_n1) );
  NOR2X0 U5775_U1 ( .IN1(n4896), .IN2(U5775_n1), .QN(WX11202) );
  INVX0 U5776_U2 ( .INP(test_so95), .ZN(U5776_n1) );
  NOR2X0 U5776_U1 ( .IN1(n4896), .IN2(U5776_n1), .QN(WX11200) );
  INVX0 U5777_U2 ( .INP(WX11135), .ZN(U5777_n1) );
  NOR2X0 U5777_U1 ( .IN1(n4896), .IN2(U5777_n1), .QN(WX11198) );
  INVX0 U5778_U2 ( .INP(WX11133), .ZN(U5778_n1) );
  NOR2X0 U5778_U1 ( .IN1(n4897), .IN2(U5778_n1), .QN(WX11196) );
  INVX0 U5779_U2 ( .INP(WX11131), .ZN(U5779_n1) );
  NOR2X0 U5779_U1 ( .IN1(n4897), .IN2(U5779_n1), .QN(WX11194) );
  INVX0 U5780_U2 ( .INP(WX11129), .ZN(U5780_n1) );
  NOR2X0 U5780_U1 ( .IN1(n4897), .IN2(U5780_n1), .QN(WX11192) );
  INVX0 U5781_U2 ( .INP(WX11127), .ZN(U5781_n1) );
  NOR2X0 U5781_U1 ( .IN1(n4897), .IN2(U5781_n1), .QN(WX11190) );
  INVX0 U5782_U2 ( .INP(WX11125), .ZN(U5782_n1) );
  NOR2X0 U5782_U1 ( .IN1(n4898), .IN2(U5782_n1), .QN(WX11188) );
  INVX0 U5783_U2 ( .INP(WX11123), .ZN(U5783_n1) );
  NOR2X0 U5783_U1 ( .IN1(n4898), .IN2(U5783_n1), .QN(WX11186) );
  INVX0 U5784_U2 ( .INP(WX11121), .ZN(U5784_n1) );
  NOR2X0 U5784_U1 ( .IN1(n4898), .IN2(U5784_n1), .QN(WX11184) );
  INVX0 U5785_U2 ( .INP(WX11119), .ZN(U5785_n1) );
  NOR2X0 U5785_U1 ( .IN1(n4898), .IN2(U5785_n1), .QN(WX11182) );
  INVX0 U5786_U2 ( .INP(WX11117), .ZN(U5786_n1) );
  NOR2X0 U5786_U1 ( .IN1(n4898), .IN2(U5786_n1), .QN(WX11180) );
  INVX0 U5787_U2 ( .INP(WX11115), .ZN(U5787_n1) );
  NOR2X0 U5787_U1 ( .IN1(n4898), .IN2(U5787_n1), .QN(WX11178) );
  INVX0 U5788_U2 ( .INP(WX11113), .ZN(U5788_n1) );
  NOR2X0 U5788_U1 ( .IN1(n4898), .IN2(U5788_n1), .QN(WX11176) );
  INVX0 U5789_U2 ( .INP(WX11111), .ZN(U5789_n1) );
  NOR2X0 U5789_U1 ( .IN1(n4898), .IN2(U5789_n1), .QN(WX11174) );
  INVX0 U5790_U2 ( .INP(WX11109), .ZN(U5790_n1) );
  NOR2X0 U5790_U1 ( .IN1(n4898), .IN2(U5790_n1), .QN(WX11172) );
  INVX0 U5791_U2 ( .INP(WX11107), .ZN(U5791_n1) );
  NOR2X0 U5791_U1 ( .IN1(n4898), .IN2(U5791_n1), .QN(WX11170) );
  INVX0 U5792_U2 ( .INP(WX11105), .ZN(U5792_n1) );
  NOR2X0 U5792_U1 ( .IN1(n4899), .IN2(U5792_n1), .QN(WX11168) );
  INVX0 U5793_U2 ( .INP(test_so94), .ZN(U5793_n1) );
  NOR2X0 U5793_U1 ( .IN1(n4899), .IN2(U5793_n1), .QN(WX11166) );
  INVX0 U5794_U2 ( .INP(WX11101), .ZN(U5794_n1) );
  NOR2X0 U5794_U1 ( .IN1(n4899), .IN2(U5794_n1), .QN(WX11164) );
  INVX0 U5795_U2 ( .INP(WX11099), .ZN(U5795_n1) );
  NOR2X0 U5795_U1 ( .IN1(n4899), .IN2(U5795_n1), .QN(WX11162) );
  INVX0 U5796_U2 ( .INP(WX11097), .ZN(U5796_n1) );
  NOR2X0 U5796_U1 ( .IN1(n4899), .IN2(U5796_n1), .QN(WX11160) );
  INVX0 U5797_U2 ( .INP(WX11095), .ZN(U5797_n1) );
  NOR2X0 U5797_U1 ( .IN1(n4899), .IN2(U5797_n1), .QN(WX11158) );
  INVX0 U5798_U2 ( .INP(WX11093), .ZN(U5798_n1) );
  NOR2X0 U5798_U1 ( .IN1(n4899), .IN2(U5798_n1), .QN(WX11156) );
  INVX0 U5799_U2 ( .INP(WX11091), .ZN(U5799_n1) );
  NOR2X0 U5799_U1 ( .IN1(n4899), .IN2(U5799_n1), .QN(WX11154) );
  INVX0 U5800_U2 ( .INP(WX11089), .ZN(U5800_n1) );
  NOR2X0 U5800_U1 ( .IN1(n4899), .IN2(U5800_n1), .QN(WX11152) );
  INVX0 U5801_U2 ( .INP(WX11087), .ZN(U5801_n1) );
  NOR2X0 U5801_U1 ( .IN1(n4899), .IN2(U5801_n1), .QN(WX11150) );
  INVX0 U5802_U2 ( .INP(WX11085), .ZN(U5802_n1) );
  NOR2X0 U5802_U1 ( .IN1(n4899), .IN2(U5802_n1), .QN(WX11148) );
  INVX0 U5803_U2 ( .INP(WX11083), .ZN(U5803_n1) );
  NOR2X0 U5803_U1 ( .IN1(n4900), .IN2(U5803_n1), .QN(WX11146) );
  INVX0 U5804_U2 ( .INP(WX11081), .ZN(U5804_n1) );
  NOR2X0 U5804_U1 ( .IN1(n4900), .IN2(U5804_n1), .QN(WX11144) );
  INVX0 U5805_U2 ( .INP(WX11079), .ZN(U5805_n1) );
  NOR2X0 U5805_U1 ( .IN1(n4900), .IN2(U5805_n1), .QN(WX11142) );
  INVX0 U5806_U2 ( .INP(WX11077), .ZN(U5806_n1) );
  NOR2X0 U5806_U1 ( .IN1(n4900), .IN2(U5806_n1), .QN(WX11140) );
  INVX0 U5807_U2 ( .INP(WX11075), .ZN(U5807_n1) );
  NOR2X0 U5807_U1 ( .IN1(n4900), .IN2(U5807_n1), .QN(WX11138) );
  INVX0 U5808_U2 ( .INP(WX11073), .ZN(U5808_n1) );
  NOR2X0 U5808_U1 ( .IN1(n4901), .IN2(U5808_n1), .QN(WX11136) );
  INVX0 U5809_U2 ( .INP(WX11071), .ZN(U5809_n1) );
  NOR2X0 U5809_U1 ( .IN1(n4902), .IN2(U5809_n1), .QN(WX11134) );
  INVX0 U5810_U2 ( .INP(test_so93), .ZN(U5810_n1) );
  NOR2X0 U5810_U1 ( .IN1(n4902), .IN2(U5810_n1), .QN(WX11132) );
  INVX0 U5811_U2 ( .INP(WX11067), .ZN(U5811_n1) );
  NOR2X0 U5811_U1 ( .IN1(n4902), .IN2(U5811_n1), .QN(WX11130) );
  INVX0 U5812_U2 ( .INP(WX11065), .ZN(U5812_n1) );
  NOR2X0 U5812_U1 ( .IN1(n4902), .IN2(U5812_n1), .QN(WX11128) );
  INVX0 U5813_U2 ( .INP(WX11063), .ZN(U5813_n1) );
  NOR2X0 U5813_U1 ( .IN1(n4902), .IN2(U5813_n1), .QN(WX11126) );
  INVX0 U5814_U2 ( .INP(WX11061), .ZN(U5814_n1) );
  NOR2X0 U5814_U1 ( .IN1(n4902), .IN2(U5814_n1), .QN(WX11124) );
  INVX0 U5815_U2 ( .INP(WX11059), .ZN(U5815_n1) );
  NOR2X0 U5815_U1 ( .IN1(n4902), .IN2(U5815_n1), .QN(WX11122) );
  INVX0 U5816_U2 ( .INP(WX11057), .ZN(U5816_n1) );
  NOR2X0 U5816_U1 ( .IN1(n4902), .IN2(U5816_n1), .QN(WX11120) );
  INVX0 U5817_U2 ( .INP(WX11055), .ZN(U5817_n1) );
  NOR2X0 U5817_U1 ( .IN1(n4902), .IN2(U5817_n1), .QN(WX11118) );
  INVX0 U5818_U2 ( .INP(WX11053), .ZN(U5818_n1) );
  NOR2X0 U5818_U1 ( .IN1(n4902), .IN2(U5818_n1), .QN(WX11116) );
  INVX0 U5819_U2 ( .INP(WX11051), .ZN(U5819_n1) );
  NOR2X0 U5819_U1 ( .IN1(n4902), .IN2(U5819_n1), .QN(WX11114) );
  INVX0 U5820_U2 ( .INP(WX11049), .ZN(U5820_n1) );
  NOR2X0 U5820_U1 ( .IN1(n4903), .IN2(U5820_n1), .QN(WX11112) );
  INVX0 U5821_U2 ( .INP(WX11047), .ZN(U5821_n1) );
  NOR2X0 U5821_U1 ( .IN1(n4903), .IN2(U5821_n1), .QN(WX11110) );
  INVX0 U5822_U2 ( .INP(WX11045), .ZN(U5822_n1) );
  NOR2X0 U5822_U1 ( .IN1(n4903), .IN2(U5822_n1), .QN(WX11108) );
  INVX0 U5823_U2 ( .INP(WX11043), .ZN(U5823_n1) );
  NOR2X0 U5823_U1 ( .IN1(n4903), .IN2(U5823_n1), .QN(WX11106) );
  INVX0 U5824_U2 ( .INP(WX11041), .ZN(U5824_n1) );
  NOR2X0 U5824_U1 ( .IN1(n4903), .IN2(U5824_n1), .QN(WX11104) );
  INVX0 U5825_U2 ( .INP(WX11039), .ZN(U5825_n1) );
  NOR2X0 U5825_U1 ( .IN1(n4903), .IN2(U5825_n1), .QN(WX11102) );
  INVX0 U5826_U2 ( .INP(WX11037), .ZN(U5826_n1) );
  NOR2X0 U5826_U1 ( .IN1(n4903), .IN2(U5826_n1), .QN(WX11100) );
  INVX0 U5827_U2 ( .INP(test_so92), .ZN(U5827_n1) );
  NOR2X0 U5827_U1 ( .IN1(n4903), .IN2(U5827_n1), .QN(WX11098) );
  INVX0 U5828_U2 ( .INP(WX11033), .ZN(U5828_n1) );
  NOR2X0 U5828_U1 ( .IN1(n4903), .IN2(U5828_n1), .QN(WX11096) );
  INVX0 U5829_U2 ( .INP(WX11031), .ZN(U5829_n1) );
  NOR2X0 U5829_U1 ( .IN1(n4888), .IN2(U5829_n1), .QN(WX11094) );
  INVX0 U5830_U2 ( .INP(WX11029), .ZN(U5830_n1) );
  NOR2X0 U5830_U1 ( .IN1(n4883), .IN2(U5830_n1), .QN(WX11092) );
  INVX0 U5831_U2 ( .INP(WX11027), .ZN(U5831_n1) );
  NOR2X0 U5831_U1 ( .IN1(n4883), .IN2(U5831_n1), .QN(WX11090) );
  INVX0 U5832_U2 ( .INP(WX11025), .ZN(U5832_n1) );
  NOR2X0 U5832_U1 ( .IN1(n4883), .IN2(U5832_n1), .QN(WX11088) );
  INVX0 U5833_U2 ( .INP(WX11023), .ZN(U5833_n1) );
  NOR2X0 U5833_U1 ( .IN1(n4883), .IN2(U5833_n1), .QN(WX11086) );
  INVX0 U5834_U2 ( .INP(WX11021), .ZN(U5834_n1) );
  NOR2X0 U5834_U1 ( .IN1(n4884), .IN2(U5834_n1), .QN(WX11084) );
  INVX0 U5835_U2 ( .INP(WX9886), .ZN(U5835_n1) );
  NOR2X0 U5835_U1 ( .IN1(n4884), .IN2(U5835_n1), .QN(WX9949) );
  INVX0 U5836_U2 ( .INP(WX9884), .ZN(U5836_n1) );
  NOR2X0 U5836_U1 ( .IN1(n4884), .IN2(U5836_n1), .QN(WX9947) );
  INVX0 U5837_U2 ( .INP(WX9882), .ZN(U5837_n1) );
  NOR2X0 U5837_U1 ( .IN1(n4884), .IN2(U5837_n1), .QN(WX9945) );
  INVX0 U5838_U2 ( .INP(WX9880), .ZN(U5838_n1) );
  NOR2X0 U5838_U1 ( .IN1(n4884), .IN2(U5838_n1), .QN(WX9943) );
  INVX0 U5839_U2 ( .INP(WX9878), .ZN(U5839_n1) );
  NOR2X0 U5839_U1 ( .IN1(n4884), .IN2(U5839_n1), .QN(WX9941) );
  INVX0 U5840_U2 ( .INP(WX9876), .ZN(U5840_n1) );
  NOR2X0 U5840_U1 ( .IN1(n4884), .IN2(U5840_n1), .QN(WX9939) );
  INVX0 U5841_U2 ( .INP(WX9874), .ZN(U5841_n1) );
  NOR2X0 U5841_U1 ( .IN1(n4884), .IN2(U5841_n1), .QN(WX9937) );
  INVX0 U5842_U2 ( .INP(WX9872), .ZN(U5842_n1) );
  NOR2X0 U5842_U1 ( .IN1(n4884), .IN2(U5842_n1), .QN(WX9935) );
  INVX0 U5843_U2 ( .INP(WX9870), .ZN(U5843_n1) );
  NOR2X0 U5843_U1 ( .IN1(n4884), .IN2(U5843_n1), .QN(WX9933) );
  INVX0 U5844_U2 ( .INP(WX9868), .ZN(U5844_n1) );
  NOR2X0 U5844_U1 ( .IN1(n4884), .IN2(U5844_n1), .QN(WX9931) );
  INVX0 U5845_U2 ( .INP(WX9866), .ZN(U5845_n1) );
  NOR2X0 U5845_U1 ( .IN1(n4885), .IN2(U5845_n1), .QN(WX9929) );
  INVX0 U5846_U2 ( .INP(WX9864), .ZN(U5846_n1) );
  NOR2X0 U5846_U1 ( .IN1(n4885), .IN2(U5846_n1), .QN(WX9927) );
  INVX0 U5847_U2 ( .INP(WX9862), .ZN(U5847_n1) );
  NOR2X0 U5847_U1 ( .IN1(n4885), .IN2(U5847_n1), .QN(WX9925) );
  INVX0 U5848_U2 ( .INP(WX9860), .ZN(U5848_n1) );
  NOR2X0 U5848_U1 ( .IN1(n4885), .IN2(U5848_n1), .QN(WX9923) );
  INVX0 U5849_U2 ( .INP(WX9858), .ZN(U5849_n1) );
  NOR2X0 U5849_U1 ( .IN1(n4885), .IN2(U5849_n1), .QN(WX9921) );
  INVX0 U5850_U2 ( .INP(WX9856), .ZN(U5850_n1) );
  NOR2X0 U5850_U1 ( .IN1(n4885), .IN2(U5850_n1), .QN(WX9919) );
  INVX0 U5851_U2 ( .INP(test_so84), .ZN(U5851_n1) );
  NOR2X0 U5851_U1 ( .IN1(n4885), .IN2(U5851_n1), .QN(WX9917) );
  INVX0 U5852_U2 ( .INP(WX9852), .ZN(U5852_n1) );
  NOR2X0 U5852_U1 ( .IN1(n4885), .IN2(U5852_n1), .QN(WX9915) );
  INVX0 U5853_U2 ( .INP(WX9850), .ZN(U5853_n1) );
  NOR2X0 U5853_U1 ( .IN1(n4885), .IN2(U5853_n1), .QN(WX9913) );
  INVX0 U5854_U2 ( .INP(WX9848), .ZN(U5854_n1) );
  NOR2X0 U5854_U1 ( .IN1(n4885), .IN2(U5854_n1), .QN(WX9911) );
  INVX0 U5855_U2 ( .INP(WX9846), .ZN(U5855_n1) );
  NOR2X0 U5855_U1 ( .IN1(n4885), .IN2(U5855_n1), .QN(WX9909) );
  INVX0 U5856_U2 ( .INP(WX9844), .ZN(U5856_n1) );
  NOR2X0 U5856_U1 ( .IN1(n4886), .IN2(U5856_n1), .QN(WX9907) );
  INVX0 U5857_U2 ( .INP(WX9842), .ZN(U5857_n1) );
  NOR2X0 U5857_U1 ( .IN1(n4886), .IN2(U5857_n1), .QN(WX9905) );
  INVX0 U5858_U2 ( .INP(WX9840), .ZN(U5858_n1) );
  NOR2X0 U5858_U1 ( .IN1(n4886), .IN2(U5858_n1), .QN(WX9903) );
  INVX0 U5859_U2 ( .INP(WX9838), .ZN(U5859_n1) );
  NOR2X0 U5859_U1 ( .IN1(n4886), .IN2(U5859_n1), .QN(WX9901) );
  INVX0 U5860_U2 ( .INP(WX9836), .ZN(U5860_n1) );
  NOR2X0 U5860_U1 ( .IN1(n4886), .IN2(U5860_n1), .QN(WX9899) );
  INVX0 U5861_U2 ( .INP(WX9834), .ZN(U5861_n1) );
  NOR2X0 U5861_U1 ( .IN1(n4886), .IN2(U5861_n1), .QN(WX9897) );
  INVX0 U5862_U2 ( .INP(WX9832), .ZN(U5862_n1) );
  NOR2X0 U5862_U1 ( .IN1(n4886), .IN2(U5862_n1), .QN(WX9895) );
  INVX0 U5863_U2 ( .INP(WX9830), .ZN(U5863_n1) );
  NOR2X0 U5863_U1 ( .IN1(n4886), .IN2(U5863_n1), .QN(WX9893) );
  INVX0 U5864_U2 ( .INP(WX9828), .ZN(U5864_n1) );
  NOR2X0 U5864_U1 ( .IN1(n4886), .IN2(U5864_n1), .QN(WX9891) );
  INVX0 U5865_U2 ( .INP(WX9826), .ZN(U5865_n1) );
  NOR2X0 U5865_U1 ( .IN1(n4886), .IN2(U5865_n1), .QN(WX9889) );
  INVX0 U5866_U2 ( .INP(WX9824), .ZN(U5866_n1) );
  NOR2X0 U5866_U1 ( .IN1(n4886), .IN2(U5866_n1), .QN(WX9887) );
  INVX0 U5867_U2 ( .INP(WX9822), .ZN(U5867_n1) );
  NOR2X0 U5867_U1 ( .IN1(n4887), .IN2(U5867_n1), .QN(WX9885) );
  INVX0 U5868_U2 ( .INP(test_so83), .ZN(U5868_n1) );
  NOR2X0 U5868_U1 ( .IN1(n4887), .IN2(U5868_n1), .QN(WX9883) );
  INVX0 U5869_U2 ( .INP(WX9818), .ZN(U5869_n1) );
  NOR2X0 U5869_U1 ( .IN1(n4887), .IN2(U5869_n1), .QN(WX9881) );
  INVX0 U5870_U2 ( .INP(WX9816), .ZN(U5870_n1) );
  NOR2X0 U5870_U1 ( .IN1(n4887), .IN2(U5870_n1), .QN(WX9879) );
  INVX0 U5871_U2 ( .INP(WX9814), .ZN(U5871_n1) );
  NOR2X0 U5871_U1 ( .IN1(n4887), .IN2(U5871_n1), .QN(WX9877) );
  INVX0 U5872_U2 ( .INP(WX9812), .ZN(U5872_n1) );
  NOR2X0 U5872_U1 ( .IN1(n4887), .IN2(U5872_n1), .QN(WX9875) );
  INVX0 U5873_U2 ( .INP(WX9810), .ZN(U5873_n1) );
  NOR2X0 U5873_U1 ( .IN1(n4887), .IN2(U5873_n1), .QN(WX9873) );
  INVX0 U5874_U2 ( .INP(WX9808), .ZN(U5874_n1) );
  NOR2X0 U5874_U1 ( .IN1(n4887), .IN2(U5874_n1), .QN(WX9871) );
  INVX0 U5875_U2 ( .INP(WX9806), .ZN(U5875_n1) );
  NOR2X0 U5875_U1 ( .IN1(n4887), .IN2(U5875_n1), .QN(WX9869) );
  INVX0 U5876_U2 ( .INP(WX9804), .ZN(U5876_n1) );
  NOR2X0 U5876_U1 ( .IN1(n4887), .IN2(U5876_n1), .QN(WX9867) );
  INVX0 U5877_U2 ( .INP(WX9802), .ZN(U5877_n1) );
  NOR2X0 U5877_U1 ( .IN1(n4887), .IN2(U5877_n1), .QN(WX9865) );
  INVX0 U5878_U2 ( .INP(WX9800), .ZN(U5878_n1) );
  NOR2X0 U5878_U1 ( .IN1(n4888), .IN2(U5878_n1), .QN(WX9863) );
  INVX0 U5879_U2 ( .INP(WX9798), .ZN(U5879_n1) );
  NOR2X0 U5879_U1 ( .IN1(n4888), .IN2(U5879_n1), .QN(WX9861) );
  INVX0 U5880_U2 ( .INP(WX9796), .ZN(U5880_n1) );
  NOR2X0 U5880_U1 ( .IN1(n4888), .IN2(U5880_n1), .QN(WX9859) );
  INVX0 U5881_U2 ( .INP(WX9794), .ZN(U5881_n1) );
  NOR2X0 U5881_U1 ( .IN1(n4888), .IN2(U5881_n1), .QN(WX9857) );
  INVX0 U5882_U2 ( .INP(WX9792), .ZN(U5882_n1) );
  NOR2X0 U5882_U1 ( .IN1(n4888), .IN2(U5882_n1), .QN(WX9855) );
  INVX0 U5883_U2 ( .INP(WX9790), .ZN(U5883_n1) );
  NOR2X0 U5883_U1 ( .IN1(n4888), .IN2(U5883_n1), .QN(WX9853) );
  INVX0 U5884_U2 ( .INP(WX9788), .ZN(U5884_n1) );
  NOR2X0 U5884_U1 ( .IN1(n4888), .IN2(U5884_n1), .QN(WX9851) );
  INVX0 U5885_U2 ( .INP(test_so82), .ZN(U5885_n1) );
  NOR2X0 U5885_U1 ( .IN1(n4888), .IN2(U5885_n1), .QN(WX9849) );
  INVX0 U5886_U2 ( .INP(WX9784), .ZN(U5886_n1) );
  NOR2X0 U5886_U1 ( .IN1(n4888), .IN2(U5886_n1), .QN(WX9847) );
  INVX0 U5887_U2 ( .INP(WX9782), .ZN(U5887_n1) );
  NOR2X0 U5887_U1 ( .IN1(n4888), .IN2(U5887_n1), .QN(WX9845) );
  INVX0 U5888_U2 ( .INP(WX9780), .ZN(U5888_n1) );
  NOR2X0 U5888_U1 ( .IN1(n4889), .IN2(U5888_n1), .QN(WX9843) );
  INVX0 U5889_U2 ( .INP(WX9778), .ZN(U5889_n1) );
  NOR2X0 U5889_U1 ( .IN1(n4889), .IN2(U5889_n1), .QN(WX9841) );
  INVX0 U5890_U2 ( .INP(WX9776), .ZN(U5890_n1) );
  NOR2X0 U5890_U1 ( .IN1(n4889), .IN2(U5890_n1), .QN(WX9839) );
  INVX0 U5891_U2 ( .INP(WX9774), .ZN(U5891_n1) );
  NOR2X0 U5891_U1 ( .IN1(n4889), .IN2(U5891_n1), .QN(WX9837) );
  INVX0 U5892_U2 ( .INP(WX9772), .ZN(U5892_n1) );
  NOR2X0 U5892_U1 ( .IN1(n4889), .IN2(U5892_n1), .QN(WX9835) );
  INVX0 U5893_U2 ( .INP(WX9770), .ZN(U5893_n1) );
  NOR2X0 U5893_U1 ( .IN1(n4889), .IN2(U5893_n1), .QN(WX9833) );
  INVX0 U5894_U2 ( .INP(WX9768), .ZN(U5894_n1) );
  NOR2X0 U5894_U1 ( .IN1(n4889), .IN2(U5894_n1), .QN(WX9831) );
  INVX0 U5895_U2 ( .INP(WX9766), .ZN(U5895_n1) );
  NOR2X0 U5895_U1 ( .IN1(n4889), .IN2(U5895_n1), .QN(WX9829) );
  INVX0 U5896_U2 ( .INP(WX9764), .ZN(U5896_n1) );
  NOR2X0 U5896_U1 ( .IN1(n4889), .IN2(U5896_n1), .QN(WX9827) );
  INVX0 U5897_U2 ( .INP(WX9762), .ZN(U5897_n1) );
  NOR2X0 U5897_U1 ( .IN1(n4889), .IN2(U5897_n1), .QN(WX9825) );
  INVX0 U5898_U2 ( .INP(WX9760), .ZN(U5898_n1) );
  NOR2X0 U5898_U1 ( .IN1(n4889), .IN2(U5898_n1), .QN(WX9823) );
  INVX0 U5899_U2 ( .INP(WX9758), .ZN(U5899_n1) );
  NOR2X0 U5899_U1 ( .IN1(n4890), .IN2(U5899_n1), .QN(WX9821) );
  INVX0 U5900_U2 ( .INP(WX9756), .ZN(U5900_n1) );
  NOR2X0 U5900_U1 ( .IN1(n4890), .IN2(U5900_n1), .QN(WX9819) );
  INVX0 U5901_U2 ( .INP(WX9754), .ZN(U5901_n1) );
  NOR2X0 U5901_U1 ( .IN1(n4890), .IN2(U5901_n1), .QN(WX9817) );
  INVX0 U5902_U2 ( .INP(test_so81), .ZN(U5902_n1) );
  NOR2X0 U5902_U1 ( .IN1(n4890), .IN2(U5902_n1), .QN(WX9815) );
  INVX0 U5903_U2 ( .INP(WX9750), .ZN(U5903_n1) );
  NOR2X0 U5903_U1 ( .IN1(n4890), .IN2(U5903_n1), .QN(WX9813) );
  INVX0 U5904_U2 ( .INP(WX9748), .ZN(U5904_n1) );
  NOR2X0 U5904_U1 ( .IN1(n4890), .IN2(U5904_n1), .QN(WX9811) );
  INVX0 U5905_U2 ( .INP(WX9746), .ZN(U5905_n1) );
  NOR2X0 U5905_U1 ( .IN1(n4890), .IN2(U5905_n1), .QN(WX9809) );
  INVX0 U5906_U2 ( .INP(WX9744), .ZN(U5906_n1) );
  NOR2X0 U5906_U1 ( .IN1(n4890), .IN2(U5906_n1), .QN(WX9807) );
  INVX0 U5907_U2 ( .INP(WX9742), .ZN(U5907_n1) );
  NOR2X0 U5907_U1 ( .IN1(n4890), .IN2(U5907_n1), .QN(WX9805) );
  INVX0 U5908_U2 ( .INP(WX9740), .ZN(U5908_n1) );
  NOR2X0 U5908_U1 ( .IN1(n4890), .IN2(U5908_n1), .QN(WX9803) );
  INVX0 U5909_U2 ( .INP(WX9738), .ZN(U5909_n1) );
  NOR2X0 U5909_U1 ( .IN1(n4890), .IN2(U5909_n1), .QN(WX9801) );
  INVX0 U5910_U2 ( .INP(WX9736), .ZN(U5910_n1) );
  NOR2X0 U5910_U1 ( .IN1(n4891), .IN2(U5910_n1), .QN(WX9799) );
  INVX0 U5911_U2 ( .INP(WX9734), .ZN(U5911_n1) );
  NOR2X0 U5911_U1 ( .IN1(n4891), .IN2(U5911_n1), .QN(WX9797) );
  INVX0 U5912_U2 ( .INP(WX9732), .ZN(U5912_n1) );
  NOR2X0 U5912_U1 ( .IN1(n4891), .IN2(U5912_n1), .QN(WX9795) );
  INVX0 U5913_U2 ( .INP(WX9730), .ZN(U5913_n1) );
  NOR2X0 U5913_U1 ( .IN1(n4891), .IN2(U5913_n1), .QN(WX9793) );
  INVX0 U5914_U2 ( .INP(WX9728), .ZN(U5914_n1) );
  NOR2X0 U5914_U1 ( .IN1(n4891), .IN2(U5914_n1), .QN(WX9791) );
  INVX0 U5915_U2 ( .INP(WX8593), .ZN(U5915_n1) );
  NOR2X0 U5915_U1 ( .IN1(n4891), .IN2(U5915_n1), .QN(WX8656) );
  INVX0 U5916_U2 ( .INP(WX8591), .ZN(U5916_n1) );
  NOR2X0 U5916_U1 ( .IN1(n4891), .IN2(U5916_n1), .QN(WX8654) );
  INVX0 U5917_U2 ( .INP(WX8589), .ZN(U5917_n1) );
  NOR2X0 U5917_U1 ( .IN1(n4891), .IN2(U5917_n1), .QN(WX8652) );
  INVX0 U5918_U2 ( .INP(WX8587), .ZN(U5918_n1) );
  NOR2X0 U5918_U1 ( .IN1(n4891), .IN2(U5918_n1), .QN(WX8650) );
  INVX0 U5919_U2 ( .INP(WX8585), .ZN(U5919_n1) );
  NOR2X0 U5919_U1 ( .IN1(n4891), .IN2(U5919_n1), .QN(WX8648) );
  INVX0 U5920_U2 ( .INP(WX8583), .ZN(U5920_n1) );
  NOR2X0 U5920_U1 ( .IN1(n4891), .IN2(U5920_n1), .QN(WX8646) );
  INVX0 U5921_U2 ( .INP(WX8581), .ZN(U5921_n1) );
  NOR2X0 U5921_U1 ( .IN1(n4892), .IN2(U5921_n1), .QN(WX8644) );
  INVX0 U5922_U2 ( .INP(WX8579), .ZN(U5922_n1) );
  NOR2X0 U5922_U1 ( .IN1(n4892), .IN2(U5922_n1), .QN(WX8642) );
  INVX0 U5923_U2 ( .INP(WX8577), .ZN(U5923_n1) );
  NOR2X0 U5923_U1 ( .IN1(n4892), .IN2(U5923_n1), .QN(WX8640) );
  INVX0 U5924_U2 ( .INP(WX8575), .ZN(U5924_n1) );
  NOR2X0 U5924_U1 ( .IN1(n4892), .IN2(U5924_n1), .QN(WX8638) );
  INVX0 U5925_U2 ( .INP(WX8573), .ZN(U5925_n1) );
  NOR2X0 U5925_U1 ( .IN1(n4892), .IN2(U5925_n1), .QN(WX8636) );
  INVX0 U5926_U2 ( .INP(test_so73), .ZN(U5926_n1) );
  NOR2X0 U5926_U1 ( .IN1(n4892), .IN2(U5926_n1), .QN(WX8634) );
  INVX0 U5927_U2 ( .INP(WX8569), .ZN(U5927_n1) );
  NOR2X0 U5927_U1 ( .IN1(n4892), .IN2(U5927_n1), .QN(WX8632) );
  INVX0 U5928_U2 ( .INP(WX8567), .ZN(U5928_n1) );
  NOR2X0 U5928_U1 ( .IN1(n4892), .IN2(U5928_n1), .QN(WX8630) );
  INVX0 U5929_U2 ( .INP(WX8565), .ZN(U5929_n1) );
  NOR2X0 U5929_U1 ( .IN1(n4892), .IN2(U5929_n1), .QN(WX8628) );
  INVX0 U5930_U2 ( .INP(WX8563), .ZN(U5930_n1) );
  NOR2X0 U5930_U1 ( .IN1(n4892), .IN2(U5930_n1), .QN(WX8626) );
  INVX0 U5931_U2 ( .INP(WX8561), .ZN(U5931_n1) );
  NOR2X0 U5931_U1 ( .IN1(n4892), .IN2(U5931_n1), .QN(WX8624) );
  INVX0 U5932_U2 ( .INP(WX8559), .ZN(U5932_n1) );
  NOR2X0 U5932_U1 ( .IN1(n4893), .IN2(U5932_n1), .QN(WX8622) );
  INVX0 U5933_U2 ( .INP(WX8557), .ZN(U5933_n1) );
  NOR2X0 U5933_U1 ( .IN1(n4893), .IN2(U5933_n1), .QN(WX8620) );
  INVX0 U5934_U2 ( .INP(WX8555), .ZN(U5934_n1) );
  NOR2X0 U5934_U1 ( .IN1(n4893), .IN2(U5934_n1), .QN(WX8618) );
  INVX0 U5935_U2 ( .INP(WX8553), .ZN(U5935_n1) );
  NOR2X0 U5935_U1 ( .IN1(n4893), .IN2(U5935_n1), .QN(WX8616) );
  INVX0 U5936_U2 ( .INP(WX8551), .ZN(U5936_n1) );
  NOR2X0 U5936_U1 ( .IN1(n4893), .IN2(U5936_n1), .QN(WX8614) );
  INVX0 U5937_U2 ( .INP(WX8549), .ZN(U5937_n1) );
  NOR2X0 U5937_U1 ( .IN1(n4893), .IN2(U5937_n1), .QN(WX8612) );
  INVX0 U5938_U2 ( .INP(WX8547), .ZN(U5938_n1) );
  NOR2X0 U5938_U1 ( .IN1(n4893), .IN2(U5938_n1), .QN(WX8610) );
  INVX0 U5939_U2 ( .INP(WX8545), .ZN(U5939_n1) );
  NOR2X0 U5939_U1 ( .IN1(n4893), .IN2(U5939_n1), .QN(WX8608) );
  INVX0 U5940_U2 ( .INP(WX8543), .ZN(U5940_n1) );
  NOR2X0 U5940_U1 ( .IN1(n4919), .IN2(U5940_n1), .QN(WX8606) );
  INVX0 U5941_U2 ( .INP(WX8541), .ZN(U5941_n1) );
  NOR2X0 U5941_U1 ( .IN1(n4914), .IN2(U5941_n1), .QN(WX8604) );
  INVX0 U5942_U2 ( .INP(WX8539), .ZN(U5942_n1) );
  NOR2X0 U5942_U1 ( .IN1(n4914), .IN2(U5942_n1), .QN(WX8602) );
  INVX0 U5943_U2 ( .INP(test_so72), .ZN(U5943_n1) );
  NOR2X0 U5943_U1 ( .IN1(n4914), .IN2(U5943_n1), .QN(WX8600) );
  INVX0 U5944_U2 ( .INP(WX8535), .ZN(U5944_n1) );
  NOR2X0 U5944_U1 ( .IN1(n4914), .IN2(U5944_n1), .QN(WX8598) );
  INVX0 U5945_U2 ( .INP(WX8533), .ZN(U5945_n1) );
  NOR2X0 U5945_U1 ( .IN1(n4914), .IN2(U5945_n1), .QN(WX8596) );
  INVX0 U5946_U2 ( .INP(WX8531), .ZN(U5946_n1) );
  NOR2X0 U5946_U1 ( .IN1(n4914), .IN2(U5946_n1), .QN(WX8594) );
  INVX0 U5947_U2 ( .INP(WX8529), .ZN(U5947_n1) );
  NOR2X0 U5947_U1 ( .IN1(n4914), .IN2(U5947_n1), .QN(WX8592) );
  INVX0 U5948_U2 ( .INP(WX8527), .ZN(U5948_n1) );
  NOR2X0 U5948_U1 ( .IN1(n4914), .IN2(U5948_n1), .QN(WX8590) );
  INVX0 U5949_U2 ( .INP(WX8525), .ZN(U5949_n1) );
  NOR2X0 U5949_U1 ( .IN1(n4914), .IN2(U5949_n1), .QN(WX8588) );
  INVX0 U5950_U2 ( .INP(WX8523), .ZN(U5950_n1) );
  NOR2X0 U5950_U1 ( .IN1(n4914), .IN2(U5950_n1), .QN(WX8586) );
  INVX0 U5951_U2 ( .INP(WX8521), .ZN(U5951_n1) );
  NOR2X0 U5951_U1 ( .IN1(n4914), .IN2(U5951_n1), .QN(WX8584) );
  INVX0 U5952_U2 ( .INP(WX8519), .ZN(U5952_n1) );
  NOR2X0 U5952_U1 ( .IN1(n4915), .IN2(U5952_n1), .QN(WX8582) );
  INVX0 U5953_U2 ( .INP(WX8517), .ZN(U5953_n1) );
  NOR2X0 U5953_U1 ( .IN1(n4915), .IN2(U5953_n1), .QN(WX8580) );
  INVX0 U5954_U2 ( .INP(WX8515), .ZN(U5954_n1) );
  NOR2X0 U5954_U1 ( .IN1(n4915), .IN2(U5954_n1), .QN(WX8578) );
  INVX0 U5955_U2 ( .INP(WX8513), .ZN(U5955_n1) );
  NOR2X0 U5955_U1 ( .IN1(n4915), .IN2(U5955_n1), .QN(WX8576) );
  INVX0 U5956_U2 ( .INP(WX8511), .ZN(U5956_n1) );
  NOR2X0 U5956_U1 ( .IN1(n4915), .IN2(U5956_n1), .QN(WX8574) );
  INVX0 U5957_U2 ( .INP(WX8509), .ZN(U5957_n1) );
  NOR2X0 U5957_U1 ( .IN1(n4915), .IN2(U5957_n1), .QN(WX8572) );
  INVX0 U5958_U2 ( .INP(WX8507), .ZN(U5958_n1) );
  NOR2X0 U5958_U1 ( .IN1(n4915), .IN2(U5958_n1), .QN(WX8570) );
  INVX0 U5959_U2 ( .INP(WX8505), .ZN(U5959_n1) );
  NOR2X0 U5959_U1 ( .IN1(n4915), .IN2(U5959_n1), .QN(WX8568) );
  INVX0 U5960_U2 ( .INP(test_so71), .ZN(U5960_n1) );
  NOR2X0 U5960_U1 ( .IN1(n4915), .IN2(U5960_n1), .QN(WX8566) );
  INVX0 U5961_U2 ( .INP(WX8501), .ZN(U5961_n1) );
  NOR2X0 U5961_U1 ( .IN1(n4915), .IN2(U5961_n1), .QN(WX8564) );
  INVX0 U5962_U2 ( .INP(WX8499), .ZN(U5962_n1) );
  NOR2X0 U5962_U1 ( .IN1(n4915), .IN2(U5962_n1), .QN(WX8562) );
  INVX0 U5963_U2 ( .INP(WX8497), .ZN(U5963_n1) );
  NOR2X0 U5963_U1 ( .IN1(n4916), .IN2(U5963_n1), .QN(WX8560) );
  INVX0 U5964_U2 ( .INP(WX8495), .ZN(U5964_n1) );
  NOR2X0 U5964_U1 ( .IN1(n4916), .IN2(U5964_n1), .QN(WX8558) );
  INVX0 U5965_U2 ( .INP(WX8493), .ZN(U5965_n1) );
  NOR2X0 U5965_U1 ( .IN1(n4916), .IN2(U5965_n1), .QN(WX8556) );
  INVX0 U5966_U2 ( .INP(WX8491), .ZN(U5966_n1) );
  NOR2X0 U5966_U1 ( .IN1(n4916), .IN2(U5966_n1), .QN(WX8554) );
  INVX0 U5967_U2 ( .INP(WX8489), .ZN(U5967_n1) );
  NOR2X0 U5967_U1 ( .IN1(n4916), .IN2(U5967_n1), .QN(WX8552) );
  INVX0 U5968_U2 ( .INP(WX8487), .ZN(U5968_n1) );
  NOR2X0 U5968_U1 ( .IN1(n4916), .IN2(U5968_n1), .QN(WX8550) );
  INVX0 U5969_U2 ( .INP(WX8485), .ZN(U5969_n1) );
  NOR2X0 U5969_U1 ( .IN1(n4916), .IN2(U5969_n1), .QN(WX8548) );
  INVX0 U5970_U2 ( .INP(WX8483), .ZN(U5970_n1) );
  NOR2X0 U5970_U1 ( .IN1(n4916), .IN2(U5970_n1), .QN(WX8546) );
  INVX0 U5971_U2 ( .INP(WX8481), .ZN(U5971_n1) );
  NOR2X0 U5971_U1 ( .IN1(n4916), .IN2(U5971_n1), .QN(WX8544) );
  INVX0 U5972_U2 ( .INP(WX8479), .ZN(U5972_n1) );
  NOR2X0 U5972_U1 ( .IN1(n4916), .IN2(U5972_n1), .QN(WX8542) );
  INVX0 U5973_U2 ( .INP(WX8477), .ZN(U5973_n1) );
  NOR2X0 U5973_U1 ( .IN1(n4916), .IN2(U5973_n1), .QN(WX8540) );
  INVX0 U5974_U2 ( .INP(WX8475), .ZN(U5974_n1) );
  NOR2X0 U5974_U1 ( .IN1(n4917), .IN2(U5974_n1), .QN(WX8538) );
  INVX0 U5975_U2 ( .INP(WX8473), .ZN(U5975_n1) );
  NOR2X0 U5975_U1 ( .IN1(n4917), .IN2(U5975_n1), .QN(WX8536) );
  INVX0 U5976_U2 ( .INP(WX8471), .ZN(U5976_n1) );
  NOR2X0 U5976_U1 ( .IN1(n4917), .IN2(U5976_n1), .QN(WX8534) );
  INVX0 U5977_U2 ( .INP(test_so70), .ZN(U5977_n1) );
  NOR2X0 U5977_U1 ( .IN1(n4917), .IN2(U5977_n1), .QN(WX8532) );
  INVX0 U5978_U2 ( .INP(WX8467), .ZN(U5978_n1) );
  NOR2X0 U5978_U1 ( .IN1(n4917), .IN2(U5978_n1), .QN(WX8530) );
  INVX0 U5979_U2 ( .INP(WX8465), .ZN(U5979_n1) );
  NOR2X0 U5979_U1 ( .IN1(n4917), .IN2(U5979_n1), .QN(WX8528) );
  INVX0 U5980_U2 ( .INP(WX8463), .ZN(U5980_n1) );
  NOR2X0 U5980_U1 ( .IN1(n4917), .IN2(U5980_n1), .QN(WX8526) );
  INVX0 U5981_U2 ( .INP(WX8461), .ZN(U5981_n1) );
  NOR2X0 U5981_U1 ( .IN1(n4917), .IN2(U5981_n1), .QN(WX8524) );
  INVX0 U5982_U2 ( .INP(WX8459), .ZN(U5982_n1) );
  NOR2X0 U5982_U1 ( .IN1(n4917), .IN2(U5982_n1), .QN(WX8522) );
  INVX0 U5983_U2 ( .INP(WX8457), .ZN(U5983_n1) );
  NOR2X0 U5983_U1 ( .IN1(n4917), .IN2(U5983_n1), .QN(WX8520) );
  INVX0 U5984_U2 ( .INP(WX8455), .ZN(U5984_n1) );
  NOR2X0 U5984_U1 ( .IN1(n4917), .IN2(U5984_n1), .QN(WX8518) );
  INVX0 U5985_U2 ( .INP(WX8453), .ZN(U5985_n1) );
  NOR2X0 U5985_U1 ( .IN1(n4918), .IN2(U5985_n1), .QN(WX8516) );
  INVX0 U5986_U2 ( .INP(WX8451), .ZN(U5986_n1) );
  NOR2X0 U5986_U1 ( .IN1(n4918), .IN2(U5986_n1), .QN(WX8514) );
  INVX0 U5987_U2 ( .INP(WX8449), .ZN(U5987_n1) );
  NOR2X0 U5987_U1 ( .IN1(n4918), .IN2(U5987_n1), .QN(WX8512) );
  INVX0 U5988_U2 ( .INP(WX8447), .ZN(U5988_n1) );
  NOR2X0 U5988_U1 ( .IN1(n4918), .IN2(U5988_n1), .QN(WX8510) );
  INVX0 U5989_U2 ( .INP(WX8445), .ZN(U5989_n1) );
  NOR2X0 U5989_U1 ( .IN1(n4918), .IN2(U5989_n1), .QN(WX8508) );
  INVX0 U5990_U2 ( .INP(WX8443), .ZN(U5990_n1) );
  NOR2X0 U5990_U1 ( .IN1(n4918), .IN2(U5990_n1), .QN(WX8506) );
  INVX0 U5991_U2 ( .INP(WX8441), .ZN(U5991_n1) );
  NOR2X0 U5991_U1 ( .IN1(n4918), .IN2(U5991_n1), .QN(WX8504) );
  INVX0 U5992_U2 ( .INP(WX8439), .ZN(U5992_n1) );
  NOR2X0 U5992_U1 ( .IN1(n4918), .IN2(U5992_n1), .QN(WX8502) );
  INVX0 U5993_U2 ( .INP(WX8437), .ZN(U5993_n1) );
  NOR2X0 U5993_U1 ( .IN1(n4918), .IN2(U5993_n1), .QN(WX8500) );
  INVX0 U5994_U2 ( .INP(test_so69), .ZN(U5994_n1) );
  NOR2X0 U5994_U1 ( .IN1(n4918), .IN2(U5994_n1), .QN(WX8498) );
  INVX0 U5995_U2 ( .INP(WX7300), .ZN(U5995_n1) );
  NOR2X0 U5995_U1 ( .IN1(n4918), .IN2(U5995_n1), .QN(WX7363) );
  INVX0 U5996_U2 ( .INP(WX7298), .ZN(U5996_n1) );
  NOR2X0 U5996_U1 ( .IN1(n4919), .IN2(U5996_n1), .QN(WX7361) );
  INVX0 U5997_U2 ( .INP(WX7296), .ZN(U5997_n1) );
  NOR2X0 U5997_U1 ( .IN1(n4919), .IN2(U5997_n1), .QN(WX7359) );
  INVX0 U5998_U2 ( .INP(WX7294), .ZN(U5998_n1) );
  NOR2X0 U5998_U1 ( .IN1(n4919), .IN2(U5998_n1), .QN(WX7357) );
  INVX0 U5999_U2 ( .INP(WX7292), .ZN(U5999_n1) );
  NOR2X0 U5999_U1 ( .IN1(n4919), .IN2(U5999_n1), .QN(WX7355) );
  INVX0 U6000_U2 ( .INP(WX7290), .ZN(U6000_n1) );
  NOR2X0 U6000_U1 ( .IN1(n4919), .IN2(U6000_n1), .QN(WX7353) );
  INVX0 U6001_U2 ( .INP(test_so62), .ZN(U6001_n1) );
  NOR2X0 U6001_U1 ( .IN1(n4919), .IN2(U6001_n1), .QN(WX7351) );
  INVX0 U6002_U2 ( .INP(WX7286), .ZN(U6002_n1) );
  NOR2X0 U6002_U1 ( .IN1(n4919), .IN2(U6002_n1), .QN(WX7349) );
  INVX0 U6003_U2 ( .INP(WX7284), .ZN(U6003_n1) );
  NOR2X0 U6003_U1 ( .IN1(n4919), .IN2(U6003_n1), .QN(WX7347) );
  INVX0 U6004_U2 ( .INP(WX7282), .ZN(U6004_n1) );
  NOR2X0 U6004_U1 ( .IN1(n4919), .IN2(U6004_n1), .QN(WX7345) );
  INVX0 U6005_U2 ( .INP(WX7280), .ZN(U6005_n1) );
  NOR2X0 U6005_U1 ( .IN1(n4919), .IN2(U6005_n1), .QN(WX7343) );
  INVX0 U6006_U2 ( .INP(WX7278), .ZN(U6006_n1) );
  NOR2X0 U6006_U1 ( .IN1(n4920), .IN2(U6006_n1), .QN(WX7341) );
  INVX0 U6007_U2 ( .INP(WX7276), .ZN(U6007_n1) );
  NOR2X0 U6007_U1 ( .IN1(n4920), .IN2(U6007_n1), .QN(WX7339) );
  INVX0 U6008_U2 ( .INP(WX7274), .ZN(U6008_n1) );
  NOR2X0 U6008_U1 ( .IN1(n4920), .IN2(U6008_n1), .QN(WX7337) );
  INVX0 U6009_U2 ( .INP(WX7272), .ZN(U6009_n1) );
  NOR2X0 U6009_U1 ( .IN1(n4920), .IN2(U6009_n1), .QN(WX7335) );
  INVX0 U6010_U2 ( .INP(WX7270), .ZN(U6010_n1) );
  NOR2X0 U6010_U1 ( .IN1(n4920), .IN2(U6010_n1), .QN(WX7333) );
  INVX0 U6011_U2 ( .INP(WX7268), .ZN(U6011_n1) );
  NOR2X0 U6011_U1 ( .IN1(n4921), .IN2(U6011_n1), .QN(WX7331) );
  INVX0 U6012_U2 ( .INP(WX7266), .ZN(U6012_n1) );
  NOR2X0 U6012_U1 ( .IN1(n4921), .IN2(U6012_n1), .QN(WX7329) );
  INVX0 U6013_U2 ( .INP(WX7264), .ZN(U6013_n1) );
  NOR2X0 U6013_U1 ( .IN1(n4920), .IN2(U6013_n1), .QN(WX7327) );
  INVX0 U6014_U2 ( .INP(WX7262), .ZN(U6014_n1) );
  NOR2X0 U6014_U1 ( .IN1(n4921), .IN2(U6014_n1), .QN(WX7325) );
  INVX0 U6015_U2 ( .INP(WX7260), .ZN(U6015_n1) );
  NOR2X0 U6015_U1 ( .IN1(n4921), .IN2(U6015_n1), .QN(WX7323) );
  INVX0 U6016_U2 ( .INP(WX7258), .ZN(U6016_n1) );
  NOR2X0 U6016_U1 ( .IN1(n4920), .IN2(U6016_n1), .QN(WX7321) );
  INVX0 U6017_U2 ( .INP(WX7256), .ZN(U6017_n1) );
  NOR2X0 U6017_U1 ( .IN1(n4921), .IN2(U6017_n1), .QN(WX7319) );
  INVX0 U6018_U2 ( .INP(test_so61), .ZN(U6018_n1) );
  NOR2X0 U6018_U1 ( .IN1(n4921), .IN2(U6018_n1), .QN(WX7317) );
  INVX0 U6019_U2 ( .INP(WX7252), .ZN(U6019_n1) );
  NOR2X0 U6019_U1 ( .IN1(n4920), .IN2(U6019_n1), .QN(WX7315) );
  INVX0 U6020_U2 ( .INP(WX7250), .ZN(U6020_n1) );
  NOR2X0 U6020_U1 ( .IN1(n4921), .IN2(U6020_n1), .QN(WX7313) );
  INVX0 U6021_U2 ( .INP(WX7248), .ZN(U6021_n1) );
  NOR2X0 U6021_U1 ( .IN1(n4921), .IN2(U6021_n1), .QN(WX7311) );
  INVX0 U6022_U2 ( .INP(WX7246), .ZN(U6022_n1) );
  NOR2X0 U6022_U1 ( .IN1(n4920), .IN2(U6022_n1), .QN(WX7309) );
  INVX0 U6023_U2 ( .INP(WX7244), .ZN(U6023_n1) );
  NOR2X0 U6023_U1 ( .IN1(n4922), .IN2(U6023_n1), .QN(WX7307) );
  INVX0 U6024_U2 ( .INP(WX7242), .ZN(U6024_n1) );
  NOR2X0 U6024_U1 ( .IN1(n4922), .IN2(U6024_n1), .QN(WX7305) );
  INVX0 U6025_U2 ( .INP(WX7240), .ZN(U6025_n1) );
  NOR2X0 U6025_U1 ( .IN1(n4920), .IN2(U6025_n1), .QN(WX7303) );
  INVX0 U6026_U2 ( .INP(WX7238), .ZN(U6026_n1) );
  NOR2X0 U6026_U1 ( .IN1(n4922), .IN2(U6026_n1), .QN(WX7301) );
  INVX0 U6027_U2 ( .INP(WX7236), .ZN(U6027_n1) );
  NOR2X0 U6027_U1 ( .IN1(n4922), .IN2(U6027_n1), .QN(WX7299) );
  INVX0 U6028_U2 ( .INP(WX7234), .ZN(U6028_n1) );
  NOR2X0 U6028_U1 ( .IN1(n4921), .IN2(U6028_n1), .QN(WX7297) );
  INVX0 U6029_U2 ( .INP(WX7232), .ZN(U6029_n1) );
  NOR2X0 U6029_U1 ( .IN1(n4922), .IN2(U6029_n1), .QN(WX7295) );
  INVX0 U6030_U2 ( .INP(WX7230), .ZN(U6030_n1) );
  NOR2X0 U6030_U1 ( .IN1(n4922), .IN2(U6030_n1), .QN(WX7293) );
  INVX0 U6031_U2 ( .INP(WX7228), .ZN(U6031_n1) );
  NOR2X0 U6031_U1 ( .IN1(n4921), .IN2(U6031_n1), .QN(WX7291) );
  INVX0 U6032_U2 ( .INP(WX7226), .ZN(U6032_n1) );
  NOR2X0 U6032_U1 ( .IN1(n4922), .IN2(U6032_n1), .QN(WX7289) );
  INVX0 U6033_U2 ( .INP(WX7224), .ZN(U6033_n1) );
  NOR2X0 U6033_U1 ( .IN1(n4922), .IN2(U6033_n1), .QN(WX7287) );
  INVX0 U6034_U2 ( .INP(WX7222), .ZN(U6034_n1) );
  NOR2X0 U6034_U1 ( .IN1(n4923), .IN2(U6034_n1), .QN(WX7285) );
  INVX0 U6035_U2 ( .INP(test_so60), .ZN(U6035_n1) );
  NOR2X0 U6035_U1 ( .IN1(n4923), .IN2(U6035_n1), .QN(WX7283) );
  INVX0 U6036_U2 ( .INP(WX7218), .ZN(U6036_n1) );
  NOR2X0 U6036_U1 ( .IN1(n4922), .IN2(U6036_n1), .QN(WX7281) );
  INVX0 U6037_U2 ( .INP(WX7216), .ZN(U6037_n1) );
  NOR2X0 U6037_U1 ( .IN1(n4923), .IN2(U6037_n1), .QN(WX7279) );
  INVX0 U6038_U2 ( .INP(WX7214), .ZN(U6038_n1) );
  NOR2X0 U6038_U1 ( .IN1(n4923), .IN2(U6038_n1), .QN(WX7277) );
  INVX0 U6039_U2 ( .INP(WX7212), .ZN(U6039_n1) );
  NOR2X0 U6039_U1 ( .IN1(n4921), .IN2(U6039_n1), .QN(WX7275) );
  INVX0 U6040_U2 ( .INP(WX7210), .ZN(U6040_n1) );
  NOR2X0 U6040_U1 ( .IN1(n4923), .IN2(U6040_n1), .QN(WX7273) );
  INVX0 U6041_U2 ( .INP(WX7208), .ZN(U6041_n1) );
  NOR2X0 U6041_U1 ( .IN1(n4923), .IN2(U6041_n1), .QN(WX7271) );
  INVX0 U6042_U2 ( .INP(WX7206), .ZN(U6042_n1) );
  NOR2X0 U6042_U1 ( .IN1(n4922), .IN2(U6042_n1), .QN(WX7269) );
  INVX0 U6043_U2 ( .INP(WX7204), .ZN(U6043_n1) );
  NOR2X0 U6043_U1 ( .IN1(n4923), .IN2(U6043_n1), .QN(WX7267) );
  INVX0 U6044_U2 ( .INP(WX7202), .ZN(U6044_n1) );
  NOR2X0 U6044_U1 ( .IN1(n4923), .IN2(U6044_n1), .QN(WX7265) );
  INVX0 U6045_U2 ( .INP(WX7200), .ZN(U6045_n1) );
  NOR2X0 U6045_U1 ( .IN1(n4922), .IN2(U6045_n1), .QN(WX7263) );
  INVX0 U6046_U2 ( .INP(WX7198), .ZN(U6046_n1) );
  NOR2X0 U6046_U1 ( .IN1(n4923), .IN2(U6046_n1), .QN(WX7261) );
  INVX0 U6047_U2 ( .INP(WX7196), .ZN(U6047_n1) );
  NOR2X0 U6047_U1 ( .IN1(n4923), .IN2(U6047_n1), .QN(WX7259) );
  INVX0 U6048_U2 ( .INP(WX7194), .ZN(U6048_n1) );
  NOR2X0 U6048_U1 ( .IN1(n4923), .IN2(U6048_n1), .QN(WX7257) );
  INVX0 U6049_U2 ( .INP(WX7192), .ZN(U6049_n1) );
  NOR2X0 U6049_U1 ( .IN1(n4924), .IN2(U6049_n1), .QN(WX7255) );
  INVX0 U6050_U2 ( .INP(WX7190), .ZN(U6050_n1) );
  NOR2X0 U6050_U1 ( .IN1(n4920), .IN2(U6050_n1), .QN(WX7253) );
  INVX0 U6051_U2 ( .INP(WX7188), .ZN(U6051_n1) );
  NOR2X0 U6051_U1 ( .IN1(n4908), .IN2(U6051_n1), .QN(WX7251) );
  INVX0 U6052_U2 ( .INP(test_so59), .ZN(U6052_n1) );
  NOR2X0 U6052_U1 ( .IN1(n4903), .IN2(U6052_n1), .QN(WX7249) );
  INVX0 U6053_U2 ( .INP(WX7184), .ZN(U6053_n1) );
  NOR2X0 U6053_U1 ( .IN1(n4904), .IN2(U6053_n1), .QN(WX7247) );
  INVX0 U6054_U2 ( .INP(WX7182), .ZN(U6054_n1) );
  NOR2X0 U6054_U1 ( .IN1(n4904), .IN2(U6054_n1), .QN(WX7245) );
  INVX0 U6055_U2 ( .INP(WX7180), .ZN(U6055_n1) );
  NOR2X0 U6055_U1 ( .IN1(n4905), .IN2(U6055_n1), .QN(WX7243) );
  INVX0 U6056_U2 ( .INP(WX7178), .ZN(U6056_n1) );
  NOR2X0 U6056_U1 ( .IN1(n4905), .IN2(U6056_n1), .QN(WX7241) );
  INVX0 U6057_U2 ( .INP(WX7176), .ZN(U6057_n1) );
  NOR2X0 U6057_U1 ( .IN1(n4905), .IN2(U6057_n1), .QN(WX7239) );
  INVX0 U6058_U2 ( .INP(WX7174), .ZN(U6058_n1) );
  NOR2X0 U6058_U1 ( .IN1(n4905), .IN2(U6058_n1), .QN(WX7237) );
  INVX0 U6059_U2 ( .INP(WX7172), .ZN(U6059_n1) );
  NOR2X0 U6059_U1 ( .IN1(n4905), .IN2(U6059_n1), .QN(WX7235) );
  INVX0 U6060_U2 ( .INP(WX7170), .ZN(U6060_n1) );
  NOR2X0 U6060_U1 ( .IN1(n4905), .IN2(U6060_n1), .QN(WX7233) );
  INVX0 U6061_U2 ( .INP(WX7168), .ZN(U6061_n1) );
  NOR2X0 U6061_U1 ( .IN1(n4906), .IN2(U6061_n1), .QN(WX7231) );
  INVX0 U6062_U2 ( .INP(WX7166), .ZN(U6062_n1) );
  NOR2X0 U6062_U1 ( .IN1(n4906), .IN2(U6062_n1), .QN(WX7229) );
  INVX0 U6063_U2 ( .INP(WX7164), .ZN(U6063_n1) );
  NOR2X0 U6063_U1 ( .IN1(n4906), .IN2(U6063_n1), .QN(WX7227) );
  INVX0 U6064_U2 ( .INP(WX7162), .ZN(U6064_n1) );
  NOR2X0 U6064_U1 ( .IN1(n4906), .IN2(U6064_n1), .QN(WX7225) );
  INVX0 U6065_U2 ( .INP(WX7160), .ZN(U6065_n1) );
  NOR2X0 U6065_U1 ( .IN1(n4906), .IN2(U6065_n1), .QN(WX7223) );
  INVX0 U6066_U2 ( .INP(WX7158), .ZN(U6066_n1) );
  NOR2X0 U6066_U1 ( .IN1(n4906), .IN2(U6066_n1), .QN(WX7221) );
  INVX0 U6067_U2 ( .INP(WX7156), .ZN(U6067_n1) );
  NOR2X0 U6067_U1 ( .IN1(n4906), .IN2(U6067_n1), .QN(WX7219) );
  INVX0 U6068_U2 ( .INP(WX7154), .ZN(U6068_n1) );
  NOR2X0 U6068_U1 ( .IN1(n4906), .IN2(U6068_n1), .QN(WX7217) );
  INVX0 U6069_U2 ( .INP(test_so58), .ZN(U6069_n1) );
  NOR2X0 U6069_U1 ( .IN1(n4906), .IN2(U6069_n1), .QN(WX7215) );
  INVX0 U6070_U2 ( .INP(WX7150), .ZN(U6070_n1) );
  NOR2X0 U6070_U1 ( .IN1(n4906), .IN2(U6070_n1), .QN(WX7213) );
  INVX0 U6071_U2 ( .INP(WX7148), .ZN(U6071_n1) );
  NOR2X0 U6071_U1 ( .IN1(n4906), .IN2(U6071_n1), .QN(WX7211) );
  INVX0 U6072_U2 ( .INP(WX7146), .ZN(U6072_n1) );
  NOR2X0 U6072_U1 ( .IN1(n4907), .IN2(U6072_n1), .QN(WX7209) );
  INVX0 U6073_U2 ( .INP(WX7144), .ZN(U6073_n1) );
  NOR2X0 U6073_U1 ( .IN1(n4907), .IN2(U6073_n1), .QN(WX7207) );
  INVX0 U6074_U2 ( .INP(WX7142), .ZN(U6074_n1) );
  NOR2X0 U6074_U1 ( .IN1(n4907), .IN2(U6074_n1), .QN(WX7205) );
  INVX0 U6075_U2 ( .INP(WX6007), .ZN(U6075_n1) );
  NOR2X0 U6075_U1 ( .IN1(n4907), .IN2(U6075_n1), .QN(WX6070) );
  INVX0 U6076_U2 ( .INP(test_so51), .ZN(U6076_n1) );
  NOR2X0 U6076_U1 ( .IN1(n4907), .IN2(U6076_n1), .QN(WX6068) );
  INVX0 U6077_U2 ( .INP(WX6003), .ZN(U6077_n1) );
  NOR2X0 U6077_U1 ( .IN1(n4907), .IN2(U6077_n1), .QN(WX6066) );
  INVX0 U6078_U2 ( .INP(WX6001), .ZN(U6078_n1) );
  NOR2X0 U6078_U1 ( .IN1(n4907), .IN2(U6078_n1), .QN(WX6064) );
  INVX0 U6079_U2 ( .INP(WX5999), .ZN(U6079_n1) );
  NOR2X0 U6079_U1 ( .IN1(n4907), .IN2(U6079_n1), .QN(WX6062) );
  INVX0 U6080_U2 ( .INP(WX5997), .ZN(U6080_n1) );
  NOR2X0 U6080_U1 ( .IN1(n4907), .IN2(U6080_n1), .QN(WX6060) );
  INVX0 U6081_U2 ( .INP(WX5995), .ZN(U6081_n1) );
  NOR2X0 U6081_U1 ( .IN1(n4907), .IN2(U6081_n1), .QN(WX6058) );
  INVX0 U6082_U2 ( .INP(WX5993), .ZN(U6082_n1) );
  NOR2X0 U6082_U1 ( .IN1(n4907), .IN2(U6082_n1), .QN(WX6056) );
  INVX0 U6083_U2 ( .INP(WX5991), .ZN(U6083_n1) );
  NOR2X0 U6083_U1 ( .IN1(n4908), .IN2(U6083_n1), .QN(WX6054) );
  INVX0 U6084_U2 ( .INP(WX5989), .ZN(U6084_n1) );
  NOR2X0 U6084_U1 ( .IN1(n4908), .IN2(U6084_n1), .QN(WX6052) );
  INVX0 U6085_U2 ( .INP(WX5987), .ZN(U6085_n1) );
  NOR2X0 U6085_U1 ( .IN1(n4908), .IN2(U6085_n1), .QN(WX6050) );
  INVX0 U6086_U2 ( .INP(WX5985), .ZN(U6086_n1) );
  NOR2X0 U6086_U1 ( .IN1(n4908), .IN2(U6086_n1), .QN(WX6048) );
  INVX0 U6087_U2 ( .INP(WX5983), .ZN(U6087_n1) );
  NOR2X0 U6087_U1 ( .IN1(n4908), .IN2(U6087_n1), .QN(WX6046) );
  INVX0 U6088_U2 ( .INP(WX5981), .ZN(U6088_n1) );
  NOR2X0 U6088_U1 ( .IN1(n4908), .IN2(U6088_n1), .QN(WX6044) );
  INVX0 U6089_U2 ( .INP(WX5979), .ZN(U6089_n1) );
  NOR2X0 U6089_U1 ( .IN1(n4908), .IN2(U6089_n1), .QN(WX6042) );
  INVX0 U6090_U2 ( .INP(WX5977), .ZN(U6090_n1) );
  NOR2X0 U6090_U1 ( .IN1(n4909), .IN2(U6090_n1), .QN(WX6040) );
  INVX0 U6091_U2 ( .INP(WX5975), .ZN(U6091_n1) );
  NOR2X0 U6091_U1 ( .IN1(n4909), .IN2(U6091_n1), .QN(WX6038) );
  INVX0 U6092_U2 ( .INP(WX5973), .ZN(U6092_n1) );
  NOR2X0 U6092_U1 ( .IN1(n4909), .IN2(U6092_n1), .QN(WX6036) );
  INVX0 U6093_U2 ( .INP(test_so50), .ZN(U6093_n1) );
  NOR2X0 U6093_U1 ( .IN1(n4909), .IN2(U6093_n1), .QN(WX6034) );
  INVX0 U6094_U2 ( .INP(WX5969), .ZN(U6094_n1) );
  NOR2X0 U6094_U1 ( .IN1(n4909), .IN2(U6094_n1), .QN(WX6032) );
  INVX0 U6095_U2 ( .INP(WX5967), .ZN(U6095_n1) );
  NOR2X0 U6095_U1 ( .IN1(n4909), .IN2(U6095_n1), .QN(WX6030) );
  INVX0 U6096_U2 ( .INP(WX5965), .ZN(U6096_n1) );
  NOR2X0 U6096_U1 ( .IN1(n4909), .IN2(U6096_n1), .QN(WX6028) );
  INVX0 U6097_U2 ( .INP(WX5963), .ZN(U6097_n1) );
  NOR2X0 U6097_U1 ( .IN1(n4909), .IN2(U6097_n1), .QN(WX6026) );
  INVX0 U6098_U2 ( .INP(WX5961), .ZN(U6098_n1) );
  NOR2X0 U6098_U1 ( .IN1(n4909), .IN2(U6098_n1), .QN(WX6024) );
  INVX0 U6099_U2 ( .INP(WX5959), .ZN(U6099_n1) );
  NOR2X0 U6099_U1 ( .IN1(n4909), .IN2(U6099_n1), .QN(WX6022) );
  INVX0 U6100_U2 ( .INP(WX5957), .ZN(U6100_n1) );
  NOR2X0 U6100_U1 ( .IN1(n4909), .IN2(U6100_n1), .QN(WX6020) );
  INVX0 U6101_U2 ( .INP(WX5955), .ZN(U6101_n1) );
  NOR2X0 U6101_U1 ( .IN1(n4910), .IN2(U6101_n1), .QN(WX6018) );
  INVX0 U6102_U2 ( .INP(WX5953), .ZN(U6102_n1) );
  NOR2X0 U6102_U1 ( .IN1(n4912), .IN2(U6102_n1), .QN(WX6016) );
  INVX0 U6103_U2 ( .INP(WX5951), .ZN(U6103_n1) );
  NOR2X0 U6103_U1 ( .IN1(n4912), .IN2(U6103_n1), .QN(WX6014) );
  INVX0 U6104_U2 ( .INP(WX5949), .ZN(U6104_n1) );
  NOR2X0 U6104_U1 ( .IN1(n4912), .IN2(U6104_n1), .QN(WX6012) );
  INVX0 U6105_U2 ( .INP(WX5947), .ZN(U6105_n1) );
  NOR2X0 U6105_U1 ( .IN1(n4912), .IN2(U6105_n1), .QN(WX6010) );
  INVX0 U6106_U2 ( .INP(WX5945), .ZN(U6106_n1) );
  NOR2X0 U6106_U1 ( .IN1(n4912), .IN2(U6106_n1), .QN(WX6008) );
  INVX0 U6107_U2 ( .INP(WX5943), .ZN(U6107_n1) );
  NOR2X0 U6107_U1 ( .IN1(n4913), .IN2(U6107_n1), .QN(WX6006) );
  INVX0 U6108_U2 ( .INP(WX5941), .ZN(U6108_n1) );
  NOR2X0 U6108_U1 ( .IN1(n4913), .IN2(U6108_n1), .QN(WX6004) );
  INVX0 U6109_U2 ( .INP(WX5929), .ZN(U6109_n1) );
  NOR2X0 U6109_U1 ( .IN1(n4913), .IN2(U6109_n1), .QN(WX5992) );
  INVX0 U6110_U2 ( .INP(WX5927), .ZN(U6110_n1) );
  NOR2X0 U6110_U1 ( .IN1(n4913), .IN2(U6110_n1), .QN(WX5990) );
  INVX0 U6111_U2 ( .INP(WX5925), .ZN(U6111_n1) );
  NOR2X0 U6111_U1 ( .IN1(n4913), .IN2(U6111_n1), .QN(WX5988) );
  INVX0 U6112_U2 ( .INP(WX5923), .ZN(U6112_n1) );
  NOR2X0 U6112_U1 ( .IN1(n4913), .IN2(U6112_n1), .QN(WX5986) );
  INVX0 U6113_U2 ( .INP(WX5921), .ZN(U6113_n1) );
  NOR2X0 U6113_U1 ( .IN1(n4913), .IN2(U6113_n1), .QN(WX5984) );
  INVX0 U6114_U2 ( .INP(WX5919), .ZN(U6114_n1) );
  NOR2X0 U6114_U1 ( .IN1(n4913), .IN2(U6114_n1), .QN(WX5982) );
  INVX0 U6115_U2 ( .INP(WX5917), .ZN(U6115_n1) );
  NOR2X0 U6115_U1 ( .IN1(n4913), .IN2(U6115_n1), .QN(WX5980) );
  INVX0 U6116_U2 ( .INP(WX5915), .ZN(U6116_n1) );
  NOR2X0 U6116_U1 ( .IN1(n4913), .IN2(U6116_n1), .QN(WX5978) );
  INVX0 U6117_U2 ( .INP(WX5913), .ZN(U6117_n1) );
  NOR2X0 U6117_U1 ( .IN1(n4912), .IN2(U6117_n1), .QN(WX5976) );
  INVX0 U6118_U2 ( .INP(WX5911), .ZN(U6118_n1) );
  NOR2X0 U6118_U1 ( .IN1(n4912), .IN2(U6118_n1), .QN(WX5974) );
  INVX0 U6119_U2 ( .INP(WX5909), .ZN(U6119_n1) );
  NOR2X0 U6119_U1 ( .IN1(n4912), .IN2(U6119_n1), .QN(WX5972) );
  INVX0 U6120_U2 ( .INP(WX5907), .ZN(U6120_n1) );
  NOR2X0 U6120_U1 ( .IN1(n4912), .IN2(U6120_n1), .QN(WX5970) );
  INVX0 U6121_U2 ( .INP(WX5905), .ZN(U6121_n1) );
  NOR2X0 U6121_U1 ( .IN1(n4912), .IN2(U6121_n1), .QN(WX5968) );
  INVX0 U6122_U2 ( .INP(test_so48), .ZN(U6122_n1) );
  NOR2X0 U6122_U1 ( .IN1(n4912), .IN2(U6122_n1), .QN(WX5966) );
  INVX0 U6123_U2 ( .INP(WX5901), .ZN(U6123_n1) );
  NOR2X0 U6123_U1 ( .IN1(n4911), .IN2(U6123_n1), .QN(WX5964) );
  INVX0 U6124_U2 ( .INP(WX5899), .ZN(U6124_n1) );
  NOR2X0 U6124_U1 ( .IN1(n4911), .IN2(U6124_n1), .QN(WX5962) );
  INVX0 U6125_U2 ( .INP(WX5897), .ZN(U6125_n1) );
  NOR2X0 U6125_U1 ( .IN1(n4911), .IN2(U6125_n1), .QN(WX5960) );
  INVX0 U6126_U2 ( .INP(WX5895), .ZN(U6126_n1) );
  NOR2X0 U6126_U1 ( .IN1(n4911), .IN2(U6126_n1), .QN(WX5958) );
  INVX0 U6127_U2 ( .INP(WX5893), .ZN(U6127_n1) );
  NOR2X0 U6127_U1 ( .IN1(n4911), .IN2(U6127_n1), .QN(WX5956) );
  INVX0 U6128_U2 ( .INP(WX5891), .ZN(U6128_n1) );
  NOR2X0 U6128_U1 ( .IN1(n4911), .IN2(U6128_n1), .QN(WX5954) );
  INVX0 U6129_U2 ( .INP(WX5889), .ZN(U6129_n1) );
  NOR2X0 U6129_U1 ( .IN1(n4911), .IN2(U6129_n1), .QN(WX5952) );
  INVX0 U6130_U2 ( .INP(WX5887), .ZN(U6130_n1) );
  NOR2X0 U6130_U1 ( .IN1(n4911), .IN2(U6130_n1), .QN(WX5950) );
  INVX0 U6131_U2 ( .INP(WX5885), .ZN(U6131_n1) );
  NOR2X0 U6131_U1 ( .IN1(n4911), .IN2(U6131_n1), .QN(WX5948) );
  INVX0 U6132_U2 ( .INP(WX5883), .ZN(U6132_n1) );
  NOR2X0 U6132_U1 ( .IN1(n4911), .IN2(U6132_n1), .QN(WX5946) );
  INVX0 U6133_U2 ( .INP(WX5881), .ZN(U6133_n1) );
  NOR2X0 U6133_U1 ( .IN1(n4911), .IN2(U6133_n1), .QN(WX5944) );
  INVX0 U6134_U2 ( .INP(WX5879), .ZN(U6134_n1) );
  NOR2X0 U6134_U1 ( .IN1(n4910), .IN2(U6134_n1), .QN(WX5942) );
  INVX0 U6135_U2 ( .INP(WX5877), .ZN(U6135_n1) );
  NOR2X0 U6135_U1 ( .IN1(n4910), .IN2(U6135_n1), .QN(WX5940) );
  INVX0 U6136_U2 ( .INP(WX5875), .ZN(U6136_n1) );
  NOR2X0 U6136_U1 ( .IN1(n4910), .IN2(U6136_n1), .QN(WX5938) );
  INVX0 U6137_U2 ( .INP(WX5873), .ZN(U6137_n1) );
  NOR2X0 U6137_U1 ( .IN1(n4910), .IN2(U6137_n1), .QN(WX5936) );
  INVX0 U6138_U2 ( .INP(WX5871), .ZN(U6138_n1) );
  NOR2X0 U6138_U1 ( .IN1(n4910), .IN2(U6138_n1), .QN(WX5934) );
  INVX0 U6139_U2 ( .INP(test_so47), .ZN(U6139_n1) );
  NOR2X0 U6139_U1 ( .IN1(n4910), .IN2(U6139_n1), .QN(WX5932) );
  INVX0 U6140_U2 ( .INP(WX5867), .ZN(U6140_n1) );
  NOR2X0 U6140_U1 ( .IN1(n4910), .IN2(U6140_n1), .QN(WX5930) );
  INVX0 U6141_U2 ( .INP(WX5865), .ZN(U6141_n1) );
  NOR2X0 U6141_U1 ( .IN1(n4910), .IN2(U6141_n1), .QN(WX5928) );
  INVX0 U6142_U2 ( .INP(WX5863), .ZN(U6142_n1) );
  NOR2X0 U6142_U1 ( .IN1(n4910), .IN2(U6142_n1), .QN(WX5926) );
  INVX0 U6143_U2 ( .INP(WX5861), .ZN(U6143_n1) );
  NOR2X0 U6143_U1 ( .IN1(n4910), .IN2(U6143_n1), .QN(WX5924) );
  INVX0 U6144_U2 ( .INP(WX5859), .ZN(U6144_n1) );
  NOR2X0 U6144_U1 ( .IN1(n4908), .IN2(U6144_n1), .QN(WX5922) );
  INVX0 U6145_U2 ( .INP(WX5857), .ZN(U6145_n1) );
  NOR2X0 U6145_U1 ( .IN1(n4908), .IN2(U6145_n1), .QN(WX5920) );
  INVX0 U6146_U2 ( .INP(WX5855), .ZN(U6146_n1) );
  NOR2X0 U6146_U1 ( .IN1(n4908), .IN2(U6146_n1), .QN(WX5918) );
  INVX0 U6147_U2 ( .INP(WX5853), .ZN(U6147_n1) );
  NOR2X0 U6147_U1 ( .IN1(n4905), .IN2(U6147_n1), .QN(WX5916) );
  INVX0 U6148_U2 ( .INP(WX5851), .ZN(U6148_n1) );
  NOR2X0 U6148_U1 ( .IN1(n4905), .IN2(U6148_n1), .QN(WX5914) );
  INVX0 U6149_U2 ( .INP(WX5849), .ZN(U6149_n1) );
  NOR2X0 U6149_U1 ( .IN1(n4905), .IN2(U6149_n1), .QN(WX5912) );
  INVX0 U6150_U2 ( .INP(WX4714), .ZN(U6150_n1) );
  NOR2X0 U6150_U1 ( .IN1(n4905), .IN2(U6150_n1), .QN(WX4777) );
  INVX0 U6151_U2 ( .INP(WX4712), .ZN(U6151_n1) );
  NOR2X0 U6151_U1 ( .IN1(n4905), .IN2(U6151_n1), .QN(WX4775) );
  INVX0 U6152_U2 ( .INP(WX4710), .ZN(U6152_n1) );
  NOR2X0 U6152_U1 ( .IN1(n4904), .IN2(U6152_n1), .QN(WX4773) );
  INVX0 U6153_U2 ( .INP(WX4708), .ZN(U6153_n1) );
  NOR2X0 U6153_U1 ( .IN1(n4904), .IN2(U6153_n1), .QN(WX4771) );
  INVX0 U6154_U2 ( .INP(WX4706), .ZN(U6154_n1) );
  NOR2X0 U6154_U1 ( .IN1(n4904), .IN2(U6154_n1), .QN(WX4769) );
  INVX0 U6155_U2 ( .INP(WX4704), .ZN(U6155_n1) );
  NOR2X0 U6155_U1 ( .IN1(n4904), .IN2(U6155_n1), .QN(WX4767) );
  INVX0 U6156_U2 ( .INP(WX4702), .ZN(U6156_n1) );
  NOR2X0 U6156_U1 ( .IN1(n4904), .IN2(U6156_n1), .QN(WX4765) );
  INVX0 U6157_U2 ( .INP(WX4700), .ZN(U6157_n1) );
  NOR2X0 U6157_U1 ( .IN1(n4904), .IN2(U6157_n1), .QN(WX4763) );
  INVX0 U6158_U2 ( .INP(WX4698), .ZN(U6158_n1) );
  NOR2X0 U6158_U1 ( .IN1(n4904), .IN2(U6158_n1), .QN(WX4761) );
  INVX0 U6159_U2 ( .INP(WX4696), .ZN(U6159_n1) );
  NOR2X0 U6159_U1 ( .IN1(n4904), .IN2(U6159_n1), .QN(WX4759) );
  INVX0 U6160_U2 ( .INP(WX4694), .ZN(U6160_n1) );
  NOR2X0 U6160_U1 ( .IN1(n4904), .IN2(U6160_n1), .QN(WX4757) );
  INVX0 U6161_U2 ( .INP(WX4692), .ZN(U6161_n1) );
  NOR2X0 U6161_U1 ( .IN1(n4913), .IN2(U6161_n1), .QN(WX4755) );
  INVX0 U6162_U2 ( .INP(WX4690), .ZN(U6162_n1) );
  NOR2X0 U6162_U1 ( .IN1(n4868), .IN2(U6162_n1), .QN(WX4753) );
  INVX0 U6163_U2 ( .INP(test_so39), .ZN(U6163_n1) );
  NOR2X0 U6163_U1 ( .IN1(n4868), .IN2(U6163_n1), .QN(WX4751) );
  INVX0 U6164_U2 ( .INP(WX4686), .ZN(U6164_n1) );
  NOR2X0 U6164_U1 ( .IN1(n4868), .IN2(U6164_n1), .QN(WX4749) );
  INVX0 U6165_U2 ( .INP(WX4684), .ZN(U6165_n1) );
  NOR2X0 U6165_U1 ( .IN1(n4868), .IN2(U6165_n1), .QN(WX4747) );
  INVX0 U6166_U2 ( .INP(WX4682), .ZN(U6166_n1) );
  NOR2X0 U6166_U1 ( .IN1(n4868), .IN2(U6166_n1), .QN(WX4745) );
  INVX0 U6167_U2 ( .INP(WX4680), .ZN(U6167_n1) );
  NOR2X0 U6167_U1 ( .IN1(n4868), .IN2(U6167_n1), .QN(WX4743) );
  INVX0 U6168_U2 ( .INP(WX4678), .ZN(U6168_n1) );
  NOR2X0 U6168_U1 ( .IN1(n4868), .IN2(U6168_n1), .QN(WX4741) );
  INVX0 U6169_U2 ( .INP(WX4676), .ZN(U6169_n1) );
  NOR2X0 U6169_U1 ( .IN1(n4868), .IN2(U6169_n1), .QN(WX4739) );
  INVX0 U6170_U2 ( .INP(WX4674), .ZN(U6170_n1) );
  NOR2X0 U6170_U1 ( .IN1(n4868), .IN2(U6170_n1), .QN(WX4737) );
  INVX0 U6171_U2 ( .INP(WX4672), .ZN(U6171_n1) );
  NOR2X0 U6171_U1 ( .IN1(n4868), .IN2(U6171_n1), .QN(WX4735) );
  INVX0 U6172_U2 ( .INP(WX4670), .ZN(U6172_n1) );
  NOR2X0 U6172_U1 ( .IN1(n4868), .IN2(U6172_n1), .QN(WX4733) );
  INVX0 U6173_U2 ( .INP(WX4668), .ZN(U6173_n1) );
  NOR2X0 U6173_U1 ( .IN1(n4867), .IN2(U6173_n1), .QN(WX4731) );
  INVX0 U6174_U2 ( .INP(WX4666), .ZN(U6174_n1) );
  NOR2X0 U6174_U1 ( .IN1(n4867), .IN2(U6174_n1), .QN(WX4729) );
  INVX0 U6175_U2 ( .INP(WX4664), .ZN(U6175_n1) );
  NOR2X0 U6175_U1 ( .IN1(n4867), .IN2(U6175_n1), .QN(WX4727) );
  INVX0 U6176_U2 ( .INP(WX4662), .ZN(U6176_n1) );
  NOR2X0 U6176_U1 ( .IN1(n4867), .IN2(U6176_n1), .QN(WX4725) );
  INVX0 U6177_U2 ( .INP(WX4660), .ZN(U6177_n1) );
  NOR2X0 U6177_U1 ( .IN1(n4867), .IN2(U6177_n1), .QN(WX4723) );
  INVX0 U6178_U2 ( .INP(WX4658), .ZN(U6178_n1) );
  NOR2X0 U6178_U1 ( .IN1(n4867), .IN2(U6178_n1), .QN(WX4721) );
  INVX0 U6179_U2 ( .INP(WX4656), .ZN(U6179_n1) );
  NOR2X0 U6179_U1 ( .IN1(n4867), .IN2(U6179_n1), .QN(WX4719) );
  INVX0 U6180_U2 ( .INP(test_so38), .ZN(U6180_n1) );
  NOR2X0 U6180_U1 ( .IN1(n4867), .IN2(U6180_n1), .QN(WX4717) );
  INVX0 U6181_U2 ( .INP(WX4652), .ZN(U6181_n1) );
  NOR2X0 U6181_U1 ( .IN1(n4867), .IN2(U6181_n1), .QN(WX4715) );
  INVX0 U6182_U2 ( .INP(WX4650), .ZN(U6182_n1) );
  NOR2X0 U6182_U1 ( .IN1(n4867), .IN2(U6182_n1), .QN(WX4713) );
  INVX0 U6183_U2 ( .INP(WX4648), .ZN(U6183_n1) );
  NOR2X0 U6183_U1 ( .IN1(n4867), .IN2(U6183_n1), .QN(WX4711) );
  INVX0 U6184_U2 ( .INP(WX4646), .ZN(U6184_n1) );
  NOR2X0 U6184_U1 ( .IN1(n4866), .IN2(U6184_n1), .QN(WX4709) );
  INVX0 U6185_U2 ( .INP(WX4644), .ZN(U6185_n1) );
  NOR2X0 U6185_U1 ( .IN1(n4866), .IN2(U6185_n1), .QN(WX4707) );
  INVX0 U6186_U2 ( .INP(WX4642), .ZN(U6186_n1) );
  NOR2X0 U6186_U1 ( .IN1(n4866), .IN2(U6186_n1), .QN(WX4705) );
  INVX0 U6187_U2 ( .INP(WX4640), .ZN(U6187_n1) );
  NOR2X0 U6187_U1 ( .IN1(n4866), .IN2(U6187_n1), .QN(WX4703) );
  INVX0 U6188_U2 ( .INP(WX4638), .ZN(U6188_n1) );
  NOR2X0 U6188_U1 ( .IN1(n4866), .IN2(U6188_n1), .QN(WX4701) );
  INVX0 U6189_U2 ( .INP(WX4636), .ZN(U6189_n1) );
  NOR2X0 U6189_U1 ( .IN1(n4866), .IN2(U6189_n1), .QN(WX4699) );
  INVX0 U6190_U2 ( .INP(WX4634), .ZN(U6190_n1) );
  NOR2X0 U6190_U1 ( .IN1(n4866), .IN2(U6190_n1), .QN(WX4697) );
  INVX0 U6191_U2 ( .INP(WX4632), .ZN(U6191_n1) );
  NOR2X0 U6191_U1 ( .IN1(n4866), .IN2(U6191_n1), .QN(WX4695) );
  INVX0 U6192_U2 ( .INP(WX4630), .ZN(U6192_n1) );
  NOR2X0 U6192_U1 ( .IN1(n4866), .IN2(U6192_n1), .QN(WX4693) );
  INVX0 U6193_U2 ( .INP(WX4628), .ZN(U6193_n1) );
  NOR2X0 U6193_U1 ( .IN1(n4866), .IN2(U6193_n1), .QN(WX4691) );
  INVX0 U6194_U2 ( .INP(WX4626), .ZN(U6194_n1) );
  NOR2X0 U6194_U1 ( .IN1(n4866), .IN2(U6194_n1), .QN(WX4689) );
  INVX0 U6195_U2 ( .INP(WX4624), .ZN(U6195_n1) );
  NOR2X0 U6195_U1 ( .IN1(n4865), .IN2(U6195_n1), .QN(WX4687) );
  INVX0 U6196_U2 ( .INP(WX4622), .ZN(U6196_n1) );
  NOR2X0 U6196_U1 ( .IN1(n4865), .IN2(U6196_n1), .QN(WX4685) );
  INVX0 U6197_U2 ( .INP(test_so37), .ZN(U6197_n1) );
  NOR2X0 U6197_U1 ( .IN1(n4865), .IN2(U6197_n1), .QN(WX4683) );
  INVX0 U6198_U2 ( .INP(WX4618), .ZN(U6198_n1) );
  NOR2X0 U6198_U1 ( .IN1(n4865), .IN2(U6198_n1), .QN(WX4681) );
  INVX0 U6199_U2 ( .INP(WX4616), .ZN(U6199_n1) );
  NOR2X0 U6199_U1 ( .IN1(n4865), .IN2(U6199_n1), .QN(WX4679) );
  INVX0 U6200_U2 ( .INP(WX4614), .ZN(U6200_n1) );
  NOR2X0 U6200_U1 ( .IN1(n4865), .IN2(U6200_n1), .QN(WX4677) );
  INVX0 U6201_U2 ( .INP(WX4612), .ZN(U6201_n1) );
  NOR2X0 U6201_U1 ( .IN1(n4865), .IN2(U6201_n1), .QN(WX4675) );
  INVX0 U6202_U2 ( .INP(WX4610), .ZN(U6202_n1) );
  NOR2X0 U6202_U1 ( .IN1(n4865), .IN2(U6202_n1), .QN(WX4673) );
  INVX0 U6203_U2 ( .INP(WX4608), .ZN(U6203_n1) );
  NOR2X0 U6203_U1 ( .IN1(n4865), .IN2(U6203_n1), .QN(WX4671) );
  INVX0 U6204_U2 ( .INP(WX4606), .ZN(U6204_n1) );
  NOR2X0 U6204_U1 ( .IN1(n4865), .IN2(U6204_n1), .QN(WX4669) );
  INVX0 U6205_U2 ( .INP(WX4604), .ZN(U6205_n1) );
  NOR2X0 U6205_U1 ( .IN1(n4865), .IN2(U6205_n1), .QN(WX4667) );
  INVX0 U6206_U2 ( .INP(WX4602), .ZN(U6206_n1) );
  NOR2X0 U6206_U1 ( .IN1(n4864), .IN2(U6206_n1), .QN(WX4665) );
  INVX0 U6207_U2 ( .INP(WX4600), .ZN(U6207_n1) );
  NOR2X0 U6207_U1 ( .IN1(n4864), .IN2(U6207_n1), .QN(WX4663) );
  INVX0 U6208_U2 ( .INP(WX4598), .ZN(U6208_n1) );
  NOR2X0 U6208_U1 ( .IN1(n4864), .IN2(U6208_n1), .QN(WX4661) );
  INVX0 U6209_U2 ( .INP(WX4596), .ZN(U6209_n1) );
  NOR2X0 U6209_U1 ( .IN1(n4864), .IN2(U6209_n1), .QN(WX4659) );
  INVX0 U6210_U2 ( .INP(WX4594), .ZN(U6210_n1) );
  NOR2X0 U6210_U1 ( .IN1(n4864), .IN2(U6210_n1), .QN(WX4657) );
  INVX0 U6211_U2 ( .INP(WX4592), .ZN(U6211_n1) );
  NOR2X0 U6211_U1 ( .IN1(n4864), .IN2(U6211_n1), .QN(WX4655) );
  INVX0 U6212_U2 ( .INP(WX4590), .ZN(U6212_n1) );
  NOR2X0 U6212_U1 ( .IN1(n4864), .IN2(U6212_n1), .QN(WX4653) );
  INVX0 U6213_U2 ( .INP(WX4588), .ZN(U6213_n1) );
  NOR2X0 U6213_U1 ( .IN1(n4864), .IN2(U6213_n1), .QN(WX4651) );
  INVX0 U6214_U2 ( .INP(test_so36), .ZN(U6214_n1) );
  NOR2X0 U6214_U1 ( .IN1(n4864), .IN2(U6214_n1), .QN(WX4649) );
  INVX0 U6215_U2 ( .INP(WX4584), .ZN(U6215_n1) );
  NOR2X0 U6215_U1 ( .IN1(n4864), .IN2(U6215_n1), .QN(WX4647) );
  INVX0 U6216_U2 ( .INP(WX4582), .ZN(U6216_n1) );
  NOR2X0 U6216_U1 ( .IN1(n4864), .IN2(U6216_n1), .QN(WX4645) );
  INVX0 U6217_U2 ( .INP(WX4580), .ZN(U6217_n1) );
  NOR2X0 U6217_U1 ( .IN1(n4863), .IN2(U6217_n1), .QN(WX4643) );
  INVX0 U6218_U2 ( .INP(WX4578), .ZN(U6218_n1) );
  NOR2X0 U6218_U1 ( .IN1(n4863), .IN2(U6218_n1), .QN(WX4641) );
  INVX0 U6219_U2 ( .INP(WX4576), .ZN(U6219_n1) );
  NOR2X0 U6219_U1 ( .IN1(n4863), .IN2(U6219_n1), .QN(WX4639) );
  INVX0 U6220_U2 ( .INP(WX4574), .ZN(U6220_n1) );
  NOR2X0 U6220_U1 ( .IN1(n4863), .IN2(U6220_n1), .QN(WX4637) );
  INVX0 U6221_U2 ( .INP(WX4572), .ZN(U6221_n1) );
  NOR2X0 U6221_U1 ( .IN1(n4863), .IN2(U6221_n1), .QN(WX4635) );
  INVX0 U6222_U2 ( .INP(WX4570), .ZN(U6222_n1) );
  NOR2X0 U6222_U1 ( .IN1(n4863), .IN2(U6222_n1), .QN(WX4633) );
  INVX0 U6223_U2 ( .INP(WX4568), .ZN(U6223_n1) );
  NOR2X0 U6223_U1 ( .IN1(n4863), .IN2(U6223_n1), .QN(WX4631) );
  INVX0 U6224_U2 ( .INP(WX4566), .ZN(U6224_n1) );
  NOR2X0 U6224_U1 ( .IN1(n4863), .IN2(U6224_n1), .QN(WX4629) );
  INVX0 U6225_U2 ( .INP(WX4564), .ZN(U6225_n1) );
  NOR2X0 U6225_U1 ( .IN1(n4863), .IN2(U6225_n1), .QN(WX4627) );
  INVX0 U6226_U2 ( .INP(WX4562), .ZN(U6226_n1) );
  NOR2X0 U6226_U1 ( .IN1(n4863), .IN2(U6226_n1), .QN(WX4625) );
  INVX0 U6227_U2 ( .INP(WX4560), .ZN(U6227_n1) );
  NOR2X0 U6227_U1 ( .IN1(n4863), .IN2(U6227_n1), .QN(WX4623) );
  INVX0 U6228_U2 ( .INP(WX4558), .ZN(U6228_n1) );
  NOR2X0 U6228_U1 ( .IN1(n4862), .IN2(U6228_n1), .QN(WX4621) );
  INVX0 U6229_U2 ( .INP(WX4556), .ZN(U6229_n1) );
  NOR2X0 U6229_U1 ( .IN1(n4862), .IN2(U6229_n1), .QN(WX4619) );
  INVX0 U6230_U2 ( .INP(WX3421), .ZN(U6230_n1) );
  NOR2X0 U6230_U1 ( .IN1(n4862), .IN2(U6230_n1), .QN(WX3484) );
  INVX0 U6231_U2 ( .INP(WX3419), .ZN(U6231_n1) );
  NOR2X0 U6231_U1 ( .IN1(n4862), .IN2(U6231_n1), .QN(WX3482) );
  INVX0 U6232_U2 ( .INP(WX3417), .ZN(U6232_n1) );
  NOR2X0 U6232_U1 ( .IN1(n4862), .IN2(U6232_n1), .QN(WX3480) );
  INVX0 U6233_U2 ( .INP(WX3415), .ZN(U6233_n1) );
  NOR2X0 U6233_U1 ( .IN1(n4862), .IN2(U6233_n1), .QN(WX3478) );
  INVX0 U6234_U2 ( .INP(WX3413), .ZN(U6234_n1) );
  NOR2X0 U6234_U1 ( .IN1(n4862), .IN2(U6234_n1), .QN(WX3476) );
  INVX0 U6235_U2 ( .INP(WX3411), .ZN(U6235_n1) );
  NOR2X0 U6235_U1 ( .IN1(n4862), .IN2(U6235_n1), .QN(WX3474) );
  INVX0 U6236_U2 ( .INP(WX3409), .ZN(U6236_n1) );
  NOR2X0 U6236_U1 ( .IN1(n4862), .IN2(U6236_n1), .QN(WX3472) );
  INVX0 U6237_U2 ( .INP(WX3407), .ZN(U6237_n1) );
  NOR2X0 U6237_U1 ( .IN1(n4862), .IN2(U6237_n1), .QN(WX3470) );
  INVX0 U6238_U2 ( .INP(test_so28), .ZN(U6238_n1) );
  NOR2X0 U6238_U1 ( .IN1(n4862), .IN2(U6238_n1), .QN(WX3468) );
  INVX0 U6239_U2 ( .INP(WX3403), .ZN(U6239_n1) );
  NOR2X0 U6239_U1 ( .IN1(n4861), .IN2(U6239_n1), .QN(WX3466) );
  INVX0 U6240_U2 ( .INP(WX3401), .ZN(U6240_n1) );
  NOR2X0 U6240_U1 ( .IN1(n4861), .IN2(U6240_n1), .QN(WX3464) );
  INVX0 U6241_U2 ( .INP(WX3399), .ZN(U6241_n1) );
  NOR2X0 U6241_U1 ( .IN1(n4861), .IN2(U6241_n1), .QN(WX3462) );
  INVX0 U6242_U2 ( .INP(WX3397), .ZN(U6242_n1) );
  NOR2X0 U6242_U1 ( .IN1(n4861), .IN2(U6242_n1), .QN(WX3460) );
  INVX0 U6243_U2 ( .INP(WX3395), .ZN(U6243_n1) );
  NOR2X0 U6243_U1 ( .IN1(n4904), .IN2(U6243_n1), .QN(WX3458) );
  INVX0 U6244_U2 ( .INP(WX3393), .ZN(U6244_n1) );
  NOR2X0 U6244_U1 ( .IN1(n4901), .IN2(U6244_n1), .QN(WX3456) );
  INVX0 U6245_U2 ( .INP(WX3391), .ZN(U6245_n1) );
  NOR2X0 U6245_U1 ( .IN1(n4902), .IN2(U6245_n1), .QN(WX3454) );
  INVX0 U6246_U2 ( .INP(WX3389), .ZN(U6246_n1) );
  NOR2X0 U6246_U1 ( .IN1(n4873), .IN2(U6246_n1), .QN(WX3452) );
  INVX0 U6247_U2 ( .INP(WX3387), .ZN(U6247_n1) );
  NOR2X0 U6247_U1 ( .IN1(n4917), .IN2(U6247_n1), .QN(WX3450) );
  INVX0 U6248_U2 ( .INP(WX3385), .ZN(U6248_n1) );
  NOR2X0 U6248_U1 ( .IN1(n4918), .IN2(U6248_n1), .QN(WX3448) );
  INVX0 U6249_U2 ( .INP(WX3383), .ZN(U6249_n1) );
  NOR2X0 U6249_U1 ( .IN1(n4919), .IN2(U6249_n1), .QN(WX3446) );
  INVX0 U6250_U2 ( .INP(WX3381), .ZN(U6250_n1) );
  NOR2X0 U6250_U1 ( .IN1(n4920), .IN2(U6250_n1), .QN(WX3444) );
  INVX0 U6251_U2 ( .INP(WX3379), .ZN(U6251_n1) );
  NOR2X0 U6251_U1 ( .IN1(n4858), .IN2(U6251_n1), .QN(WX3442) );
  INVX0 U6252_U2 ( .INP(WX3377), .ZN(U6252_n1) );
  NOR2X0 U6252_U1 ( .IN1(n4858), .IN2(U6252_n1), .QN(WX3440) );
  INVX0 U6253_U2 ( .INP(WX3375), .ZN(U6253_n1) );
  NOR2X0 U6253_U1 ( .IN1(n4858), .IN2(U6253_n1), .QN(WX3438) );
  INVX0 U6254_U2 ( .INP(WX3373), .ZN(U6254_n1) );
  NOR2X0 U6254_U1 ( .IN1(n4858), .IN2(U6254_n1), .QN(WX3436) );
  INVX0 U6255_U2 ( .INP(WX3371), .ZN(U6255_n1) );
  NOR2X0 U6255_U1 ( .IN1(n4858), .IN2(U6255_n1), .QN(WX3434) );
  INVX0 U6256_U2 ( .INP(test_so27), .ZN(U6256_n1) );
  NOR2X0 U6256_U1 ( .IN1(n4858), .IN2(U6256_n1), .QN(WX3432) );
  INVX0 U6257_U2 ( .INP(WX3367), .ZN(U6257_n1) );
  NOR2X0 U6257_U1 ( .IN1(n4858), .IN2(U6257_n1), .QN(WX3430) );
  INVX0 U6258_U2 ( .INP(WX3365), .ZN(U6258_n1) );
  NOR2X0 U6258_U1 ( .IN1(n4858), .IN2(U6258_n1), .QN(WX3428) );
  INVX0 U6259_U2 ( .INP(WX3363), .ZN(U6259_n1) );
  NOR2X0 U6259_U1 ( .IN1(n4858), .IN2(U6259_n1), .QN(WX3426) );
  INVX0 U6260_U2 ( .INP(WX3361), .ZN(U6260_n1) );
  NOR2X0 U6260_U1 ( .IN1(n4858), .IN2(U6260_n1), .QN(WX3424) );
  INVX0 U6261_U2 ( .INP(WX3359), .ZN(U6261_n1) );
  NOR2X0 U6261_U1 ( .IN1(n4858), .IN2(U6261_n1), .QN(WX3422) );
  INVX0 U6262_U2 ( .INP(WX3357), .ZN(U6262_n1) );
  NOR2X0 U6262_U1 ( .IN1(n4872), .IN2(U6262_n1), .QN(WX3420) );
  INVX0 U6263_U2 ( .INP(WX3355), .ZN(U6263_n1) );
  NOR2X0 U6263_U1 ( .IN1(n4871), .IN2(U6263_n1), .QN(WX3418) );
  INVX0 U6264_U2 ( .INP(WX3353), .ZN(U6264_n1) );
  NOR2X0 U6264_U1 ( .IN1(n4886), .IN2(U6264_n1), .QN(WX3416) );
  INVX0 U6265_U2 ( .INP(WX3351), .ZN(U6265_n1) );
  NOR2X0 U6265_U1 ( .IN1(n4887), .IN2(U6265_n1), .QN(WX3414) );
  INVX0 U6266_U2 ( .INP(WX3349), .ZN(U6266_n1) );
  NOR2X0 U6266_U1 ( .IN1(n4874), .IN2(U6266_n1), .QN(WX3412) );
  INVX0 U6267_U2 ( .INP(WX3347), .ZN(U6267_n1) );
  NOR2X0 U6267_U1 ( .IN1(n4875), .IN2(U6267_n1), .QN(WX3410) );
  INVX0 U6268_U2 ( .INP(WX3345), .ZN(U6268_n1) );
  NOR2X0 U6268_U1 ( .IN1(n4876), .IN2(U6268_n1), .QN(WX3408) );
  INVX0 U6269_U2 ( .INP(WX3343), .ZN(U6269_n1) );
  NOR2X0 U6269_U1 ( .IN1(n4877), .IN2(U6269_n1), .QN(WX3406) );
  INVX0 U6270_U2 ( .INP(WX3341), .ZN(U6270_n1) );
  NOR2X0 U6270_U1 ( .IN1(n4878), .IN2(U6270_n1), .QN(WX3404) );
  INVX0 U6271_U2 ( .INP(WX3339), .ZN(U6271_n1) );
  NOR2X0 U6271_U1 ( .IN1(n4879), .IN2(U6271_n1), .QN(WX3402) );
  INVX0 U6272_U2 ( .INP(WX3337), .ZN(U6272_n1) );
  NOR2X0 U6272_U1 ( .IN1(n4880), .IN2(U6272_n1), .QN(WX3400) );
  INVX0 U6273_U2 ( .INP(WX3335), .ZN(U6273_n1) );
  NOR2X0 U6273_U1 ( .IN1(n4881), .IN2(U6273_n1), .QN(WX3398) );
  INVX0 U6274_U2 ( .INP(test_so26), .ZN(U6274_n1) );
  NOR2X0 U6274_U1 ( .IN1(n4911), .IN2(U6274_n1), .QN(WX3396) );
  INVX0 U6275_U2 ( .INP(WX3331), .ZN(U6275_n1) );
  NOR2X0 U6275_U1 ( .IN1(n4912), .IN2(U6275_n1), .QN(WX3394) );
  INVX0 U6276_U2 ( .INP(WX3329), .ZN(U6276_n1) );
  NOR2X0 U6276_U1 ( .IN1(n4913), .IN2(U6276_n1), .QN(WX3392) );
  INVX0 U6277_U2 ( .INP(WX3327), .ZN(U6277_n1) );
  NOR2X0 U6277_U1 ( .IN1(n4914), .IN2(U6277_n1), .QN(WX3390) );
  INVX0 U6278_U2 ( .INP(WX3325), .ZN(U6278_n1) );
  NOR2X0 U6278_U1 ( .IN1(n4915), .IN2(U6278_n1), .QN(WX3388) );
  INVX0 U6279_U2 ( .INP(WX3323), .ZN(U6279_n1) );
  NOR2X0 U6279_U1 ( .IN1(n4870), .IN2(U6279_n1), .QN(WX3386) );
  INVX0 U6280_U2 ( .INP(WX3321), .ZN(U6280_n1) );
  NOR2X0 U6280_U1 ( .IN1(n4869), .IN2(U6280_n1), .QN(WX3384) );
  INVX0 U6281_U2 ( .INP(WX3319), .ZN(U6281_n1) );
  NOR2X0 U6281_U1 ( .IN1(n4916), .IN2(U6281_n1), .QN(WX3382) );
  INVX0 U6282_U2 ( .INP(WX3317), .ZN(U6282_n1) );
  NOR2X0 U6282_U1 ( .IN1(n4903), .IN2(U6282_n1), .QN(WX3380) );
  INVX0 U6283_U2 ( .INP(WX3315), .ZN(U6283_n1) );
  NOR2X0 U6283_U1 ( .IN1(n4905), .IN2(U6283_n1), .QN(WX3378) );
  INVX0 U6284_U2 ( .INP(WX3313), .ZN(U6284_n1) );
  NOR2X0 U6284_U1 ( .IN1(n4906), .IN2(U6284_n1), .QN(WX3376) );
  INVX0 U6285_U2 ( .INP(WX3311), .ZN(U6285_n1) );
  NOR2X0 U6285_U1 ( .IN1(n4907), .IN2(U6285_n1), .QN(WX3374) );
  INVX0 U6286_U2 ( .INP(WX3309), .ZN(U6286_n1) );
  NOR2X0 U6286_U1 ( .IN1(n4908), .IN2(U6286_n1), .QN(WX3372) );
  INVX0 U6287_U2 ( .INP(WX3307), .ZN(U6287_n1) );
  NOR2X0 U6287_U1 ( .IN1(n4909), .IN2(U6287_n1), .QN(WX3370) );
  INVX0 U6288_U2 ( .INP(WX3305), .ZN(U6288_n1) );
  NOR2X0 U6288_U1 ( .IN1(n4910), .IN2(U6288_n1), .QN(WX3368) );
  INVX0 U6289_U2 ( .INP(WX3303), .ZN(U6289_n1) );
  NOR2X0 U6289_U1 ( .IN1(n4895), .IN2(U6289_n1), .QN(WX3366) );
  INVX0 U6290_U2 ( .INP(WX3301), .ZN(U6290_n1) );
  NOR2X0 U6290_U1 ( .IN1(n4896), .IN2(U6290_n1), .QN(WX3364) );
  INVX0 U6291_U2 ( .INP(WX3299), .ZN(U6291_n1) );
  NOR2X0 U6291_U1 ( .IN1(n4897), .IN2(U6291_n1), .QN(WX3362) );
  INVX0 U6292_U2 ( .INP(test_so25), .ZN(U6292_n1) );
  NOR2X0 U6292_U1 ( .IN1(n4898), .IN2(U6292_n1), .QN(WX3360) );
  INVX0 U6293_U2 ( .INP(WX3295), .ZN(U6293_n1) );
  NOR2X0 U6293_U1 ( .IN1(n4899), .IN2(U6293_n1), .QN(WX3358) );
  INVX0 U6294_U2 ( .INP(WX3293), .ZN(U6294_n1) );
  NOR2X0 U6294_U1 ( .IN1(n4859), .IN2(U6294_n1), .QN(WX3356) );
  INVX0 U6295_U2 ( .INP(WX3291), .ZN(U6295_n1) );
  NOR2X0 U6295_U1 ( .IN1(n4859), .IN2(U6295_n1), .QN(WX3354) );
  INVX0 U6296_U2 ( .INP(WX3289), .ZN(U6296_n1) );
  NOR2X0 U6296_U1 ( .IN1(n4859), .IN2(U6296_n1), .QN(WX3352) );
  INVX0 U6297_U2 ( .INP(WX3287), .ZN(U6297_n1) );
  NOR2X0 U6297_U1 ( .IN1(n4859), .IN2(U6297_n1), .QN(WX3350) );
  INVX0 U6298_U2 ( .INP(WX3285), .ZN(U6298_n1) );
  NOR2X0 U6298_U1 ( .IN1(n4859), .IN2(U6298_n1), .QN(WX3348) );
  INVX0 U6299_U2 ( .INP(WX3283), .ZN(U6299_n1) );
  NOR2X0 U6299_U1 ( .IN1(n4859), .IN2(U6299_n1), .QN(WX3346) );
  INVX0 U6300_U2 ( .INP(WX3281), .ZN(U6300_n1) );
  NOR2X0 U6300_U1 ( .IN1(n4859), .IN2(U6300_n1), .QN(WX3344) );
  INVX0 U6301_U2 ( .INP(WX3279), .ZN(U6301_n1) );
  NOR2X0 U6301_U1 ( .IN1(n4859), .IN2(U6301_n1), .QN(WX3342) );
  INVX0 U6302_U2 ( .INP(WX3277), .ZN(U6302_n1) );
  NOR2X0 U6302_U1 ( .IN1(n4859), .IN2(U6302_n1), .QN(WX3340) );
  INVX0 U6303_U2 ( .INP(WX3275), .ZN(U6303_n1) );
  NOR2X0 U6303_U1 ( .IN1(n4859), .IN2(U6303_n1), .QN(WX3338) );
  INVX0 U6304_U2 ( .INP(WX3273), .ZN(U6304_n1) );
  NOR2X0 U6304_U1 ( .IN1(n4859), .IN2(U6304_n1), .QN(WX3336) );
  INVX0 U6305_U2 ( .INP(WX3271), .ZN(U6305_n1) );
  NOR2X0 U6305_U1 ( .IN1(n4860), .IN2(U6305_n1), .QN(WX3334) );
  INVX0 U6306_U2 ( .INP(WX3267), .ZN(U6306_n1) );
  NOR2X0 U6306_U1 ( .IN1(n4860), .IN2(U6306_n1), .QN(WX3330) );
  INVX0 U6307_U2 ( .INP(WX2128), .ZN(U6307_n1) );
  NOR2X0 U6307_U1 ( .IN1(n4860), .IN2(U6307_n1), .QN(WX2191) );
  INVX0 U6308_U2 ( .INP(WX2126), .ZN(U6308_n1) );
  NOR2X0 U6308_U1 ( .IN1(n4860), .IN2(U6308_n1), .QN(WX2189) );
  INVX0 U6309_U2 ( .INP(WX2124), .ZN(U6309_n1) );
  NOR2X0 U6309_U1 ( .IN1(n4860), .IN2(U6309_n1), .QN(WX2187) );
  INVX0 U6310_U2 ( .INP(WX2122), .ZN(U6310_n1) );
  NOR2X0 U6310_U1 ( .IN1(n4860), .IN2(U6310_n1), .QN(WX2185) );
  INVX0 U6311_U2 ( .INP(WX2120), .ZN(U6311_n1) );
  NOR2X0 U6311_U1 ( .IN1(n4860), .IN2(U6311_n1), .QN(WX2183) );
  INVX0 U6312_U2 ( .INP(WX2118), .ZN(U6312_n1) );
  NOR2X0 U6312_U1 ( .IN1(n4860), .IN2(U6312_n1), .QN(WX2181) );
  INVX0 U6313_U2 ( .INP(WX2116), .ZN(U6313_n1) );
  NOR2X0 U6313_U1 ( .IN1(n4860), .IN2(U6313_n1), .QN(WX2179) );
  INVX0 U6314_U2 ( .INP(WX2114), .ZN(U6314_n1) );
  NOR2X0 U6314_U1 ( .IN1(n4860), .IN2(U6314_n1), .QN(WX2177) );
  INVX0 U6315_U2 ( .INP(WX2112), .ZN(U6315_n1) );
  NOR2X0 U6315_U1 ( .IN1(n4860), .IN2(U6315_n1), .QN(WX2175) );
  INVX0 U6316_U2 ( .INP(WX2110), .ZN(U6316_n1) );
  NOR2X0 U6316_U1 ( .IN1(n4861), .IN2(U6316_n1), .QN(WX2173) );
  INVX0 U6317_U2 ( .INP(WX2108), .ZN(U6317_n1) );
  NOR2X0 U6317_U1 ( .IN1(n4861), .IN2(U6317_n1), .QN(WX2171) );
  INVX0 U6318_U2 ( .INP(WX2106), .ZN(U6318_n1) );
  NOR2X0 U6318_U1 ( .IN1(n4861), .IN2(U6318_n1), .QN(WX2169) );
  INVX0 U6319_U2 ( .INP(WX2104), .ZN(U6319_n1) );
  NOR2X0 U6319_U1 ( .IN1(n4861), .IN2(U6319_n1), .QN(WX2167) );
  INVX0 U6320_U2 ( .INP(WX2102), .ZN(U6320_n1) );
  NOR2X0 U6320_U1 ( .IN1(n4861), .IN2(U6320_n1), .QN(WX2165) );
  INVX0 U6321_U2 ( .INP(test_so17), .ZN(U6321_n1) );
  NOR2X0 U6321_U1 ( .IN1(n4861), .IN2(U6321_n1), .QN(WX2163) );
  INVX0 U6322_U2 ( .INP(WX2098), .ZN(U6322_n1) );
  NOR2X0 U6322_U1 ( .IN1(n4861), .IN2(U6322_n1), .QN(WX2161) );
  INVX0 U6323_U2 ( .INP(WX2096), .ZN(U6323_n1) );
  NOR2X0 U6323_U1 ( .IN1(n4883), .IN2(U6323_n1), .QN(WX2159) );
  INVX0 U6324_U2 ( .INP(WX2094), .ZN(U6324_n1) );
  NOR2X0 U6324_U1 ( .IN1(n4883), .IN2(U6324_n1), .QN(WX2157) );
  INVX0 U6325_U2 ( .INP(WX2092), .ZN(U6325_n1) );
  NOR2X0 U6325_U1 ( .IN1(n4883), .IN2(U6325_n1), .QN(WX2155) );
  INVX0 U6326_U2 ( .INP(WX2090), .ZN(U6326_n1) );
  NOR2X0 U6326_U1 ( .IN1(n4883), .IN2(U6326_n1), .QN(WX2153) );
  INVX0 U6327_U2 ( .INP(WX2088), .ZN(U6327_n1) );
  NOR2X0 U6327_U1 ( .IN1(n4883), .IN2(U6327_n1), .QN(WX2151) );
  INVX0 U6328_U2 ( .INP(WX2086), .ZN(U6328_n1) );
  NOR2X0 U6328_U1 ( .IN1(n4883), .IN2(U6328_n1), .QN(WX2149) );
  INVX0 U6329_U2 ( .INP(WX2084), .ZN(U6329_n1) );
  NOR2X0 U6329_U1 ( .IN1(n4882), .IN2(U6329_n1), .QN(WX2147) );
  INVX0 U6330_U2 ( .INP(WX2082), .ZN(U6330_n1) );
  NOR2X0 U6330_U1 ( .IN1(n4882), .IN2(U6330_n1), .QN(WX2145) );
  INVX0 U6331_U2 ( .INP(WX2080), .ZN(U6331_n1) );
  NOR2X0 U6331_U1 ( .IN1(n4882), .IN2(U6331_n1), .QN(WX2143) );
  INVX0 U6332_U2 ( .INP(WX2078), .ZN(U6332_n1) );
  NOR2X0 U6332_U1 ( .IN1(n4882), .IN2(U6332_n1), .QN(WX2141) );
  INVX0 U6333_U2 ( .INP(WX2076), .ZN(U6333_n1) );
  NOR2X0 U6333_U1 ( .IN1(n4882), .IN2(U6333_n1), .QN(WX2139) );
  INVX0 U6334_U2 ( .INP(WX2074), .ZN(U6334_n1) );
  NOR2X0 U6334_U1 ( .IN1(n4882), .IN2(U6334_n1), .QN(WX2137) );
  INVX0 U6335_U2 ( .INP(WX2072), .ZN(U6335_n1) );
  NOR2X0 U6335_U1 ( .IN1(n4882), .IN2(U6335_n1), .QN(WX2135) );
  INVX0 U6336_U2 ( .INP(WX2070), .ZN(U6336_n1) );
  NOR2X0 U6336_U1 ( .IN1(n4882), .IN2(U6336_n1), .QN(WX2133) );
  INVX0 U6337_U2 ( .INP(WX2068), .ZN(U6337_n1) );
  NOR2X0 U6337_U1 ( .IN1(n4882), .IN2(U6337_n1), .QN(WX2131) );
  INVX0 U6338_U2 ( .INP(WX2066), .ZN(U6338_n1) );
  NOR2X0 U6338_U1 ( .IN1(n4882), .IN2(U6338_n1), .QN(WX2129) );
  INVX0 U6339_U2 ( .INP(test_so16), .ZN(U6339_n1) );
  NOR2X0 U6339_U1 ( .IN1(n4882), .IN2(U6339_n1), .QN(WX2127) );
  INVX0 U6340_U2 ( .INP(WX2062), .ZN(U6340_n1) );
  NOR2X0 U6340_U1 ( .IN1(n4881), .IN2(U6340_n1), .QN(WX2125) );
  INVX0 U6341_U2 ( .INP(WX2060), .ZN(U6341_n1) );
  NOR2X0 U6341_U1 ( .IN1(n4881), .IN2(U6341_n1), .QN(WX2123) );
  INVX0 U6342_U2 ( .INP(WX2058), .ZN(U6342_n1) );
  NOR2X0 U6342_U1 ( .IN1(n4881), .IN2(U6342_n1), .QN(WX2121) );
  INVX0 U6343_U2 ( .INP(WX2056), .ZN(U6343_n1) );
  NOR2X0 U6343_U1 ( .IN1(n4881), .IN2(U6343_n1), .QN(WX2119) );
  INVX0 U6344_U2 ( .INP(WX2054), .ZN(U6344_n1) );
  NOR2X0 U6344_U1 ( .IN1(n4881), .IN2(U6344_n1), .QN(WX2117) );
  INVX0 U6345_U2 ( .INP(WX2052), .ZN(U6345_n1) );
  NOR2X0 U6345_U1 ( .IN1(n4881), .IN2(U6345_n1), .QN(WX2115) );
  INVX0 U6346_U2 ( .INP(WX2050), .ZN(U6346_n1) );
  NOR2X0 U6346_U1 ( .IN1(n4881), .IN2(U6346_n1), .QN(WX2113) );
  INVX0 U6347_U2 ( .INP(WX2048), .ZN(U6347_n1) );
  NOR2X0 U6347_U1 ( .IN1(n4881), .IN2(U6347_n1), .QN(WX2111) );
  INVX0 U6348_U2 ( .INP(WX2046), .ZN(U6348_n1) );
  NOR2X0 U6348_U1 ( .IN1(n4881), .IN2(U6348_n1), .QN(WX2109) );
  INVX0 U6349_U2 ( .INP(WX2044), .ZN(U6349_n1) );
  NOR2X0 U6349_U1 ( .IN1(n4881), .IN2(U6349_n1), .QN(WX2107) );
  INVX0 U6350_U2 ( .INP(WX2042), .ZN(U6350_n1) );
  NOR2X0 U6350_U1 ( .IN1(n4881), .IN2(U6350_n1), .QN(WX2105) );
  INVX0 U6351_U2 ( .INP(WX2040), .ZN(U6351_n1) );
  NOR2X0 U6351_U1 ( .IN1(n4880), .IN2(U6351_n1), .QN(WX2103) );
  INVX0 U6352_U2 ( .INP(WX2038), .ZN(U6352_n1) );
  NOR2X0 U6352_U1 ( .IN1(n4880), .IN2(U6352_n1), .QN(WX2101) );
  INVX0 U6353_U2 ( .INP(WX2036), .ZN(U6353_n1) );
  NOR2X0 U6353_U1 ( .IN1(n4880), .IN2(U6353_n1), .QN(WX2099) );
  INVX0 U6354_U2 ( .INP(WX2034), .ZN(U6354_n1) );
  NOR2X0 U6354_U1 ( .IN1(n4880), .IN2(U6354_n1), .QN(WX2097) );
  INVX0 U6355_U2 ( .INP(WX2032), .ZN(U6355_n1) );
  NOR2X0 U6355_U1 ( .IN1(n4880), .IN2(U6355_n1), .QN(WX2095) );
  INVX0 U6356_U2 ( .INP(WX2030), .ZN(U6356_n1) );
  NOR2X0 U6356_U1 ( .IN1(n4880), .IN2(U6356_n1), .QN(WX2093) );
  INVX0 U6357_U2 ( .INP(test_so15), .ZN(U6357_n1) );
  NOR2X0 U6357_U1 ( .IN1(n4880), .IN2(U6357_n1), .QN(WX2091) );
  INVX0 U6358_U2 ( .INP(WX2026), .ZN(U6358_n1) );
  NOR2X0 U6358_U1 ( .IN1(n4880), .IN2(U6358_n1), .QN(WX2089) );
  INVX0 U6359_U2 ( .INP(WX2024), .ZN(U6359_n1) );
  NOR2X0 U6359_U1 ( .IN1(n4880), .IN2(U6359_n1), .QN(WX2087) );
  INVX0 U6360_U2 ( .INP(WX2022), .ZN(U6360_n1) );
  NOR2X0 U6360_U1 ( .IN1(n4880), .IN2(U6360_n1), .QN(WX2085) );
  INVX0 U6361_U2 ( .INP(WX2020), .ZN(U6361_n1) );
  NOR2X0 U6361_U1 ( .IN1(n4880), .IN2(U6361_n1), .QN(WX2083) );
  INVX0 U6362_U2 ( .INP(WX2018), .ZN(U6362_n1) );
  NOR2X0 U6362_U1 ( .IN1(n4879), .IN2(U6362_n1), .QN(WX2081) );
  INVX0 U6363_U2 ( .INP(WX2016), .ZN(U6363_n1) );
  NOR2X0 U6363_U1 ( .IN1(n4879), .IN2(U6363_n1), .QN(WX2079) );
  INVX0 U6364_U2 ( .INP(WX2014), .ZN(U6364_n1) );
  NOR2X0 U6364_U1 ( .IN1(n4879), .IN2(U6364_n1), .QN(WX2077) );
  INVX0 U6365_U2 ( .INP(WX2012), .ZN(U6365_n1) );
  NOR2X0 U6365_U1 ( .IN1(n4879), .IN2(U6365_n1), .QN(WX2075) );
  INVX0 U6366_U2 ( .INP(WX2010), .ZN(U6366_n1) );
  NOR2X0 U6366_U1 ( .IN1(n4879), .IN2(U6366_n1), .QN(WX2073) );
  INVX0 U6367_U2 ( .INP(WX2008), .ZN(U6367_n1) );
  NOR2X0 U6367_U1 ( .IN1(n4879), .IN2(U6367_n1), .QN(WX2071) );
  INVX0 U6368_U2 ( .INP(WX2006), .ZN(U6368_n1) );
  NOR2X0 U6368_U1 ( .IN1(n4879), .IN2(U6368_n1), .QN(WX2069) );
  INVX0 U6369_U2 ( .INP(WX2004), .ZN(U6369_n1) );
  NOR2X0 U6369_U1 ( .IN1(n4879), .IN2(U6369_n1), .QN(WX2067) );
  INVX0 U6370_U2 ( .INP(WX2002), .ZN(U6370_n1) );
  NOR2X0 U6370_U1 ( .IN1(n4879), .IN2(U6370_n1), .QN(WX2065) );
  INVX0 U6371_U2 ( .INP(WX2000), .ZN(U6371_n1) );
  NOR2X0 U6371_U1 ( .IN1(n4879), .IN2(U6371_n1), .QN(WX2063) );
  INVX0 U6372_U2 ( .INP(WX1998), .ZN(U6372_n1) );
  NOR2X0 U6372_U1 ( .IN1(n4879), .IN2(U6372_n1), .QN(WX2061) );
  INVX0 U6373_U2 ( .INP(WX1996), .ZN(U6373_n1) );
  NOR2X0 U6373_U1 ( .IN1(n4878), .IN2(U6373_n1), .QN(WX2059) );
  INVX0 U6374_U2 ( .INP(WX1994), .ZN(U6374_n1) );
  NOR2X0 U6374_U1 ( .IN1(n4878), .IN2(U6374_n1), .QN(WX2057) );
  INVX0 U6375_U2 ( .INP(test_so14), .ZN(U6375_n1) );
  NOR2X0 U6375_U1 ( .IN1(n4878), .IN2(U6375_n1), .QN(WX2055) );
  INVX0 U6376_U2 ( .INP(WX1990), .ZN(U6376_n1) );
  NOR2X0 U6376_U1 ( .IN1(n4878), .IN2(U6376_n1), .QN(WX2053) );
  INVX0 U6377_U2 ( .INP(WX1988), .ZN(U6377_n1) );
  NOR2X0 U6377_U1 ( .IN1(n4878), .IN2(U6377_n1), .QN(WX2051) );
  INVX0 U6378_U2 ( .INP(WX1986), .ZN(U6378_n1) );
  NOR2X0 U6378_U1 ( .IN1(n4878), .IN2(U6378_n1), .QN(WX2049) );
  INVX0 U6379_U2 ( .INP(WX1984), .ZN(U6379_n1) );
  NOR2X0 U6379_U1 ( .IN1(n4878), .IN2(U6379_n1), .QN(WX2047) );
  INVX0 U6380_U2 ( .INP(WX1982), .ZN(U6380_n1) );
  NOR2X0 U6380_U1 ( .IN1(n4878), .IN2(U6380_n1), .QN(WX2045) );
  INVX0 U6381_U2 ( .INP(WX1980), .ZN(U6381_n1) );
  NOR2X0 U6381_U1 ( .IN1(n4878), .IN2(U6381_n1), .QN(WX2043) );
  INVX0 U6382_U2 ( .INP(WX1978), .ZN(U6382_n1) );
  NOR2X0 U6382_U1 ( .IN1(n4878), .IN2(U6382_n1), .QN(WX2041) );
  INVX0 U6383_U2 ( .INP(WX1976), .ZN(U6383_n1) );
  NOR2X0 U6383_U1 ( .IN1(n4878), .IN2(U6383_n1), .QN(WX2039) );
  INVX0 U6384_U2 ( .INP(WX1974), .ZN(U6384_n1) );
  NOR2X0 U6384_U1 ( .IN1(n4877), .IN2(U6384_n1), .QN(WX2037) );
  INVX0 U6385_U2 ( .INP(WX1972), .ZN(U6385_n1) );
  NOR2X0 U6385_U1 ( .IN1(n4877), .IN2(U6385_n1), .QN(WX2035) );
  INVX0 U6386_U2 ( .INP(WX1970), .ZN(U6386_n1) );
  NOR2X0 U6386_U1 ( .IN1(n4877), .IN2(U6386_n1), .QN(WX2033) );
  INVX0 U6387_U2 ( .INP(WX835), .ZN(U6387_n1) );
  NOR2X0 U6387_U1 ( .IN1(n4877), .IN2(U6387_n1), .QN(WX898) );
  INVX0 U6388_U2 ( .INP(WX833), .ZN(U6388_n1) );
  NOR2X0 U6388_U1 ( .IN1(n4877), .IN2(U6388_n1), .QN(WX896) );
  INVX0 U6389_U2 ( .INP(test_so7), .ZN(U6389_n1) );
  NOR2X0 U6389_U1 ( .IN1(n4877), .IN2(U6389_n1), .QN(WX894) );
  INVX0 U6390_U2 ( .INP(WX829), .ZN(U6390_n1) );
  NOR2X0 U6390_U1 ( .IN1(n4877), .IN2(U6390_n1), .QN(WX892) );
  INVX0 U6391_U2 ( .INP(WX827), .ZN(U6391_n1) );
  NOR2X0 U6391_U1 ( .IN1(n4877), .IN2(U6391_n1), .QN(WX890) );
  INVX0 U6392_U2 ( .INP(WX825), .ZN(U6392_n1) );
  NOR2X0 U6392_U1 ( .IN1(n4877), .IN2(U6392_n1), .QN(WX888) );
  INVX0 U6393_U2 ( .INP(WX823), .ZN(U6393_n1) );
  NOR2X0 U6393_U1 ( .IN1(n4877), .IN2(U6393_n1), .QN(WX886) );
  INVX0 U6394_U2 ( .INP(WX821), .ZN(U6394_n1) );
  NOR2X0 U6394_U1 ( .IN1(n4877), .IN2(U6394_n1), .QN(WX884) );
  INVX0 U6395_U2 ( .INP(WX819), .ZN(U6395_n1) );
  NOR2X0 U6395_U1 ( .IN1(n4876), .IN2(U6395_n1), .QN(WX882) );
  INVX0 U6396_U2 ( .INP(WX817), .ZN(U6396_n1) );
  NOR2X0 U6396_U1 ( .IN1(n4876), .IN2(U6396_n1), .QN(WX880) );
  INVX0 U6397_U2 ( .INP(WX815), .ZN(U6397_n1) );
  NOR2X0 U6397_U1 ( .IN1(n4876), .IN2(U6397_n1), .QN(WX878) );
  INVX0 U6398_U2 ( .INP(WX813), .ZN(U6398_n1) );
  NOR2X0 U6398_U1 ( .IN1(n4876), .IN2(U6398_n1), .QN(WX876) );
  INVX0 U6399_U2 ( .INP(WX811), .ZN(U6399_n1) );
  NOR2X0 U6399_U1 ( .IN1(n4876), .IN2(U6399_n1), .QN(WX874) );
  INVX0 U6400_U2 ( .INP(WX809), .ZN(U6400_n1) );
  NOR2X0 U6400_U1 ( .IN1(n4876), .IN2(U6400_n1), .QN(WX872) );
  INVX0 U6401_U2 ( .INP(WX807), .ZN(U6401_n1) );
  NOR2X0 U6401_U1 ( .IN1(n4876), .IN2(U6401_n1), .QN(WX870) );
  INVX0 U6402_U2 ( .INP(WX805), .ZN(U6402_n1) );
  NOR2X0 U6402_U1 ( .IN1(n4876), .IN2(U6402_n1), .QN(WX868) );
  INVX0 U6403_U2 ( .INP(WX803), .ZN(U6403_n1) );
  NOR2X0 U6403_U1 ( .IN1(n4876), .IN2(U6403_n1), .QN(WX866) );
  INVX0 U6404_U2 ( .INP(WX801), .ZN(U6404_n1) );
  NOR2X0 U6404_U1 ( .IN1(n4876), .IN2(U6404_n1), .QN(WX864) );
  INVX0 U6405_U2 ( .INP(WX799), .ZN(U6405_n1) );
  NOR2X0 U6405_U1 ( .IN1(n4875), .IN2(U6405_n1), .QN(WX862) );
  INVX0 U6406_U2 ( .INP(WX797), .ZN(U6406_n1) );
  NOR2X0 U6406_U1 ( .IN1(n4875), .IN2(U6406_n1), .QN(WX860) );
  INVX0 U6407_U2 ( .INP(test_so6), .ZN(U6407_n1) );
  NOR2X0 U6407_U1 ( .IN1(n4875), .IN2(U6407_n1), .QN(WX858) );
  INVX0 U6408_U2 ( .INP(WX793), .ZN(U6408_n1) );
  NOR2X0 U6408_U1 ( .IN1(n4875), .IN2(U6408_n1), .QN(WX856) );
  INVX0 U6409_U2 ( .INP(WX791), .ZN(U6409_n1) );
  NOR2X0 U6409_U1 ( .IN1(n4875), .IN2(U6409_n1), .QN(WX854) );
  INVX0 U6410_U2 ( .INP(WX789), .ZN(U6410_n1) );
  NOR2X0 U6410_U1 ( .IN1(n4875), .IN2(U6410_n1), .QN(WX852) );
  INVX0 U6411_U2 ( .INP(WX787), .ZN(U6411_n1) );
  NOR2X0 U6411_U1 ( .IN1(n4875), .IN2(U6411_n1), .QN(WX850) );
  INVX0 U6412_U2 ( .INP(WX785), .ZN(U6412_n1) );
  NOR2X0 U6412_U1 ( .IN1(n4875), .IN2(U6412_n1), .QN(WX848) );
  INVX0 U6413_U2 ( .INP(WX783), .ZN(U6413_n1) );
  NOR2X0 U6413_U1 ( .IN1(n4875), .IN2(U6413_n1), .QN(WX846) );
  INVX0 U6414_U2 ( .INP(WX781), .ZN(U6414_n1) );
  NOR2X0 U6414_U1 ( .IN1(n4875), .IN2(U6414_n1), .QN(WX844) );
  INVX0 U6415_U2 ( .INP(WX779), .ZN(U6415_n1) );
  NOR2X0 U6415_U1 ( .IN1(n4875), .IN2(U6415_n1), .QN(WX842) );
  INVX0 U6416_U2 ( .INP(WX777), .ZN(U6416_n1) );
  NOR2X0 U6416_U1 ( .IN1(n4874), .IN2(U6416_n1), .QN(WX840) );
  INVX0 U6417_U2 ( .INP(WX775), .ZN(U6417_n1) );
  NOR2X0 U6417_U1 ( .IN1(n4874), .IN2(U6417_n1), .QN(WX838) );
  INVX0 U6418_U2 ( .INP(WX773), .ZN(U6418_n1) );
  NOR2X0 U6418_U1 ( .IN1(n4874), .IN2(U6418_n1), .QN(WX836) );
  INVX0 U6419_U2 ( .INP(WX771), .ZN(U6419_n1) );
  NOR2X0 U6419_U1 ( .IN1(n4874), .IN2(U6419_n1), .QN(WX834) );
  INVX0 U6420_U2 ( .INP(WX769), .ZN(U6420_n1) );
  NOR2X0 U6420_U1 ( .IN1(n4874), .IN2(U6420_n1), .QN(WX832) );
  INVX0 U6421_U2 ( .INP(WX767), .ZN(U6421_n1) );
  NOR2X0 U6421_U1 ( .IN1(n4874), .IN2(U6421_n1), .QN(WX830) );
  INVX0 U6422_U2 ( .INP(WX765), .ZN(U6422_n1) );
  NOR2X0 U6422_U1 ( .IN1(n4874), .IN2(U6422_n1), .QN(WX828) );
  INVX0 U6423_U2 ( .INP(WX763), .ZN(U6423_n1) );
  NOR2X0 U6423_U1 ( .IN1(n4874), .IN2(U6423_n1), .QN(WX826) );
  INVX0 U6424_U2 ( .INP(WX761), .ZN(U6424_n1) );
  NOR2X0 U6424_U1 ( .IN1(n4874), .IN2(U6424_n1), .QN(WX824) );
  INVX0 U6425_U2 ( .INP(test_so5), .ZN(U6425_n1) );
  NOR2X0 U6425_U1 ( .IN1(n4874), .IN2(U6425_n1), .QN(WX822) );
  INVX0 U6426_U2 ( .INP(WX757), .ZN(U6426_n1) );
  NOR2X0 U6426_U1 ( .IN1(n4874), .IN2(U6426_n1), .QN(WX820) );
  INVX0 U6427_U2 ( .INP(WX755), .ZN(U6427_n1) );
  NOR2X0 U6427_U1 ( .IN1(n4873), .IN2(U6427_n1), .QN(WX818) );
  INVX0 U6428_U2 ( .INP(WX753), .ZN(U6428_n1) );
  NOR2X0 U6428_U1 ( .IN1(n4873), .IN2(U6428_n1), .QN(WX816) );
  INVX0 U6429_U2 ( .INP(WX751), .ZN(U6429_n1) );
  NOR2X0 U6429_U1 ( .IN1(n4873), .IN2(U6429_n1), .QN(WX814) );
  INVX0 U6430_U2 ( .INP(WX749), .ZN(U6430_n1) );
  NOR2X0 U6430_U1 ( .IN1(n4873), .IN2(U6430_n1), .QN(WX812) );
  INVX0 U6431_U2 ( .INP(WX747), .ZN(U6431_n1) );
  NOR2X0 U6431_U1 ( .IN1(n4873), .IN2(U6431_n1), .QN(WX810) );
  INVX0 U6432_U2 ( .INP(WX745), .ZN(U6432_n1) );
  NOR2X0 U6432_U1 ( .IN1(n4873), .IN2(U6432_n1), .QN(WX808) );
  INVX0 U6433_U2 ( .INP(WX743), .ZN(U6433_n1) );
  NOR2X0 U6433_U1 ( .IN1(n4873), .IN2(U6433_n1), .QN(WX806) );
  INVX0 U6434_U2 ( .INP(WX741), .ZN(U6434_n1) );
  NOR2X0 U6434_U1 ( .IN1(n4873), .IN2(U6434_n1), .QN(WX804) );
  INVX0 U6435_U2 ( .INP(WX739), .ZN(U6435_n1) );
  NOR2X0 U6435_U1 ( .IN1(n4873), .IN2(U6435_n1), .QN(WX802) );
  INVX0 U6436_U2 ( .INP(WX737), .ZN(U6436_n1) );
  NOR2X0 U6436_U1 ( .IN1(n4873), .IN2(U6436_n1), .QN(WX800) );
  INVX0 U6437_U2 ( .INP(WX735), .ZN(U6437_n1) );
  NOR2X0 U6437_U1 ( .IN1(n4873), .IN2(U6437_n1), .QN(WX798) );
  INVX0 U6438_U2 ( .INP(WX733), .ZN(U6438_n1) );
  NOR2X0 U6438_U1 ( .IN1(n4872), .IN2(U6438_n1), .QN(WX796) );
  INVX0 U6439_U2 ( .INP(WX731), .ZN(U6439_n1) );
  NOR2X0 U6439_U1 ( .IN1(n4872), .IN2(U6439_n1), .QN(WX794) );
  INVX0 U6440_U2 ( .INP(WX729), .ZN(U6440_n1) );
  NOR2X0 U6440_U1 ( .IN1(n4872), .IN2(U6440_n1), .QN(WX792) );
  INVX0 U6441_U2 ( .INP(WX727), .ZN(U6441_n1) );
  NOR2X0 U6441_U1 ( .IN1(n4872), .IN2(U6441_n1), .QN(WX790) );
  INVX0 U6442_U2 ( .INP(WX725), .ZN(U6442_n1) );
  NOR2X0 U6442_U1 ( .IN1(n4872), .IN2(U6442_n1), .QN(WX788) );
  INVX0 U6443_U2 ( .INP(test_so4), .ZN(U6443_n1) );
  NOR2X0 U6443_U1 ( .IN1(n4872), .IN2(U6443_n1), .QN(WX786) );
  INVX0 U6444_U2 ( .INP(WX721), .ZN(U6444_n1) );
  NOR2X0 U6444_U1 ( .IN1(n4872), .IN2(U6444_n1), .QN(WX784) );
  INVX0 U6445_U2 ( .INP(WX719), .ZN(U6445_n1) );
  NOR2X0 U6445_U1 ( .IN1(n4872), .IN2(U6445_n1), .QN(WX782) );
  INVX0 U6446_U2 ( .INP(WX717), .ZN(U6446_n1) );
  NOR2X0 U6446_U1 ( .IN1(n4872), .IN2(U6446_n1), .QN(WX780) );
  INVX0 U6447_U2 ( .INP(WX715), .ZN(U6447_n1) );
  NOR2X0 U6447_U1 ( .IN1(n4872), .IN2(U6447_n1), .QN(WX778) );
  INVX0 U6448_U2 ( .INP(WX713), .ZN(U6448_n1) );
  NOR2X0 U6448_U1 ( .IN1(n4872), .IN2(U6448_n1), .QN(WX776) );
  INVX0 U6449_U2 ( .INP(WX711), .ZN(U6449_n1) );
  NOR2X0 U6449_U1 ( .IN1(n4871), .IN2(U6449_n1), .QN(WX774) );
  INVX0 U6450_U2 ( .INP(WX709), .ZN(U6450_n1) );
  NOR2X0 U6450_U1 ( .IN1(n4871), .IN2(U6450_n1), .QN(WX772) );
  INVX0 U6451_U2 ( .INP(WX707), .ZN(U6451_n1) );
  NOR2X0 U6451_U1 ( .IN1(n4871), .IN2(U6451_n1), .QN(WX770) );
  INVX0 U6452_U2 ( .INP(WX705), .ZN(U6452_n1) );
  NOR2X0 U6452_U1 ( .IN1(n4871), .IN2(U6452_n1), .QN(WX768) );
  INVX0 U6453_U2 ( .INP(WX703), .ZN(U6453_n1) );
  NOR2X0 U6453_U1 ( .IN1(n4871), .IN2(U6453_n1), .QN(WX766) );
  INVX0 U6454_U2 ( .INP(WX701), .ZN(U6454_n1) );
  NOR2X0 U6454_U1 ( .IN1(n4871), .IN2(U6454_n1), .QN(WX764) );
  INVX0 U6455_U2 ( .INP(WX699), .ZN(U6455_n1) );
  NOR2X0 U6455_U1 ( .IN1(n4871), .IN2(U6455_n1), .QN(WX762) );
  INVX0 U6456_U2 ( .INP(WX697), .ZN(U6456_n1) );
  NOR2X0 U6456_U1 ( .IN1(n4871), .IN2(U6456_n1), .QN(WX760) );
  INVX0 U6457_U2 ( .INP(WX695), .ZN(U6457_n1) );
  NOR2X0 U6457_U1 ( .IN1(n4871), .IN2(U6457_n1), .QN(WX758) );
  INVX0 U6458_U2 ( .INP(WX693), .ZN(U6458_n1) );
  NOR2X0 U6458_U1 ( .IN1(n4871), .IN2(U6458_n1), .QN(WX756) );
  INVX0 U6459_U2 ( .INP(WX691), .ZN(U6459_n1) );
  NOR2X0 U6459_U1 ( .IN1(n4871), .IN2(U6459_n1), .QN(WX754) );
  INVX0 U6460_U2 ( .INP(WX689), .ZN(U6460_n1) );
  NOR2X0 U6460_U1 ( .IN1(n4870), .IN2(U6460_n1), .QN(WX752) );
  INVX0 U6461_U2 ( .INP(test_so3), .ZN(U6461_n1) );
  NOR2X0 U6461_U1 ( .IN1(n4870), .IN2(U6461_n1), .QN(WX750) );
  INVX0 U6462_U2 ( .INP(WX685), .ZN(U6462_n1) );
  NOR2X0 U6462_U1 ( .IN1(n4870), .IN2(U6462_n1), .QN(WX748) );
  INVX0 U6463_U2 ( .INP(WX683), .ZN(U6463_n1) );
  NOR2X0 U6463_U1 ( .IN1(n4870), .IN2(U6463_n1), .QN(WX746) );
  INVX0 U6464_U2 ( .INP(WX681), .ZN(U6464_n1) );
  NOR2X0 U6464_U1 ( .IN1(n4870), .IN2(U6464_n1), .QN(WX744) );
  INVX0 U6465_U2 ( .INP(WX679), .ZN(U6465_n1) );
  NOR2X0 U6465_U1 ( .IN1(n4870), .IN2(U6465_n1), .QN(WX742) );
  INVX0 U6466_U2 ( .INP(WX677), .ZN(U6466_n1) );
  NOR2X0 U6466_U1 ( .IN1(n4870), .IN2(U6466_n1), .QN(WX740) );
  INVX0 U6467_U2 ( .INP(WX675), .ZN(U6467_n1) );
  NOR2X0 U6467_U1 ( .IN1(n4870), .IN2(U6467_n1), .QN(WX738) );
  INVX0 U6468_U2 ( .INP(WX673), .ZN(U6468_n1) );
  NOR2X0 U6468_U1 ( .IN1(n4870), .IN2(U6468_n1), .QN(WX736) );
  INVX0 U6469_U2 ( .INP(WX671), .ZN(U6469_n1) );
  NOR2X0 U6469_U1 ( .IN1(n4870), .IN2(U6469_n1), .QN(WX734) );
  INVX0 U6470_U2 ( .INP(WX669), .ZN(U6470_n1) );
  NOR2X0 U6470_U1 ( .IN1(n4870), .IN2(U6470_n1), .QN(WX732) );
  INVX0 U6471_U2 ( .INP(WX667), .ZN(U6471_n1) );
  NOR2X0 U6471_U1 ( .IN1(n4869), .IN2(U6471_n1), .QN(WX730) );
  INVX0 U6472_U2 ( .INP(WX665), .ZN(U6472_n1) );
  NOR2X0 U6472_U1 ( .IN1(n4869), .IN2(U6472_n1), .QN(WX728) );
  INVX0 U6473_U2 ( .INP(WX663), .ZN(U6473_n1) );
  NOR2X0 U6473_U1 ( .IN1(n4869), .IN2(U6473_n1), .QN(WX726) );
  INVX0 U6474_U2 ( .INP(WX661), .ZN(U6474_n1) );
  NOR2X0 U6474_U1 ( .IN1(n4869), .IN2(U6474_n1), .QN(WX724) );
  INVX0 U6475_U2 ( .INP(WX659), .ZN(U6475_n1) );
  NOR2X0 U6475_U1 ( .IN1(n4869), .IN2(U6475_n1), .QN(WX722) );
  INVX0 U6476_U2 ( .INP(WX657), .ZN(U6476_n1) );
  NOR2X0 U6476_U1 ( .IN1(n4869), .IN2(U6476_n1), .QN(WX720) );
  INVX0 U6477_U2 ( .INP(WX655), .ZN(U6477_n1) );
  NOR2X0 U6477_U1 ( .IN1(n4869), .IN2(U6477_n1), .QN(WX718) );
  INVX0 U6478_U2 ( .INP(WX653), .ZN(U6478_n1) );
  NOR2X0 U6478_U1 ( .IN1(n4869), .IN2(U6478_n1), .QN(WX716) );
  INVX0 U6479_U2 ( .INP(test_so2), .ZN(U6479_n1) );
  NOR2X0 U6479_U1 ( .IN1(n4869), .IN2(U6479_n1), .QN(WX714) );
  INVX0 U6480_U2 ( .INP(WX649), .ZN(U6480_n1) );
  NOR2X0 U6480_U1 ( .IN1(n4869), .IN2(U6480_n1), .QN(WX712) );
  INVX0 U6481_U2 ( .INP(WX647), .ZN(U6481_n1) );
  NOR2X0 U6481_U1 ( .IN1(n4869), .IN2(U6481_n1), .QN(WX710) );
  INVX0 U6482_U2 ( .INP(WX645), .ZN(U6482_n1) );
  NOR2X0 U6482_U1 ( .IN1(n4876), .IN2(U6482_n1), .QN(WX708) );
endmodule

