module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n236_, new_n238_, new_n250_, new_n288_, new_n421_, new_n368_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n186_, new_n365_, new_n339_, new_n197_, new_n386_, new_n246_, new_n170_, new_n266_, new_n367_, new_n173_, new_n220_, new_n419_, new_n214_, new_n424_, new_n114_, new_n188_, new_n240_, new_n413_, new_n442_, new_n211_, new_n123_, new_n127_, new_n342_, new_n317_, new_n344_, new_n287_, new_n234_, new_n418_, new_n292_, new_n215_, new_n152_, new_n157_, new_n153_, new_n133_, new_n257_, new_n212_, new_n364_, new_n272_, new_n282_, new_n201_, new_n192_, new_n414_, new_n110_, new_n315_, new_n124_, new_n326_, new_n164_, new_n230_, new_n281_, new_n430_, new_n248_, new_n117_, new_n167_, new_n385_, new_n297_, new_n361_, new_n150_, new_n108_, new_n137_, new_n183_, new_n303_, new_n351_, new_n325_, new_n180_, new_n318_, new_n321_, new_n443_, new_n158_, new_n262_, new_n271_, new_n274_, new_n218_, new_n305_, new_n420_, new_n205_, new_n141_, new_n206_, new_n254_, new_n355_, new_n353_, new_n432_, new_n256_, new_n452_, new_n381_, new_n388_, new_n194_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n314_, new_n118_, new_n165_, new_n441_, new_n216_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n395_, new_n383_, new_n343_, new_n210_, new_n207_, new_n267_, new_n140_, new_n187_, new_n311_, new_n263_, new_n334_, new_n331_, new_n341_, new_n349_, new_n244_, new_n172_, new_n277_, new_n402_, new_n286_, new_n335_, new_n347_, new_n346_, new_n396_, new_n198_, new_n438_, new_n208_, new_n179_, new_n436_, new_n233_, new_n178_, new_n295_, new_n359_, new_n132_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n155_, new_n384_, new_n410_, new_n113_, new_n371_, new_n202_, new_n296_, new_n308_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n291_, new_n261_, new_n309_, new_n323_, new_n259_, new_n362_, new_n227_, new_n416_, new_n222_, new_n400_, new_n328_, new_n130_, new_n268_, new_n374_, new_n380_, new_n138_, new_n310_, new_n144_, new_n275_, new_n352_, new_n126_, new_n177_, new_n264_, new_n379_, new_n273_, new_n224_, new_n270_, new_n143_, new_n125_, new_n145_, new_n253_, new_n237_, new_n149_, new_n260_, new_n251_, new_n189_, new_n300_, new_n106_, new_n411_, new_n107_, new_n182_, new_n407_, new_n151_, new_n219_, new_n231_, new_n313_, new_n239_, new_n428_, new_n199_, new_n146_, new_n360_, new_n302_, new_n191_, new_n225_, new_n112_, new_n121_, new_n415_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n154_, new_n131_, new_n255_, new_n459_, new_n174_, new_n354_, new_n392_, new_n444_, new_n340_, new_n147_, new_n285_, new_n209_, new_n446_, new_n203_, new_n316_, new_n417_, new_n332_, new_n453_, new_n163_, new_n148_, new_n440_, new_n122_, new_n111_, new_n252_, new_n160_, new_n312_, new_n372_, new_n242_, new_n115_, new_n307_, new_n190_, new_n408_, new_n213_, new_n134_, new_n109_, new_n265_, new_n278_, new_n304_, new_n217_, new_n269_, new_n129_, new_n412_, new_n327_, new_n431_, new_n196_, new_n319_, new_n338_, new_n336_, new_n377_, new_n247_, new_n330_, new_n375_, new_n294_, new_n195_, new_n357_, new_n320_, new_n245_, new_n404_, new_n193_, new_n128_, new_n358_, new_n348_, new_n159_, new_n322_, new_n228_, new_n289_, new_n175_, new_n226_, new_n185_, new_n373_, new_n171_, new_n434_, new_n200_, new_n422_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n168_, new_n279_, new_n455_, new_n120_, new_n406_, new_n356_, new_n229_, new_n204_, new_n181_, new_n135_, new_n405_;

not g000 ( new_n106_, keyIn_0_26 );
not g001 ( new_n107_, N1 );
xor g002 ( new_n108_, N73, N77 );
xnor g003 ( new_n109_, N65, N69 );
xnor g004 ( new_n110_, new_n108_, new_n109_ );
xor g005 ( new_n111_, N89, N93 );
xnor g006 ( new_n112_, N81, N85 );
xnor g007 ( new_n113_, new_n111_, new_n112_ );
xor g008 ( new_n114_, new_n110_, new_n113_ );
nand g009 ( new_n115_, N129, N137 );
xnor g010 ( new_n116_, new_n114_, new_n115_ );
xor g011 ( new_n117_, N33, N49 );
xnor g012 ( new_n118_, N1, N17 );
xnor g013 ( new_n119_, new_n117_, new_n118_ );
xnor g014 ( new_n120_, new_n116_, new_n119_ );
not g015 ( new_n121_, new_n120_ );
not g016 ( new_n122_, keyIn_0_18 );
not g017 ( new_n123_, keyIn_0_14 );
not g018 ( new_n124_, keyIn_0_12 );
not g019 ( new_n125_, keyIn_0_10 );
not g020 ( new_n126_, keyIn_0_7 );
not g021 ( new_n127_, keyIn_0_2 );
xnor g022 ( new_n128_, N33, N37 );
xnor g023 ( new_n129_, new_n128_, new_n127_ );
not g024 ( new_n130_, keyIn_0_3 );
xnor g025 ( new_n131_, N41, N45 );
xnor g026 ( new_n132_, new_n131_, new_n130_ );
nand g027 ( new_n133_, new_n129_, new_n132_ );
xnor g028 ( new_n134_, new_n128_, keyIn_0_2 );
xor g029 ( new_n135_, N41, N45 );
nand g030 ( new_n136_, new_n135_, new_n130_ );
nand g031 ( new_n137_, new_n131_, keyIn_0_3 );
nand g032 ( new_n138_, new_n136_, new_n137_ );
nand g033 ( new_n139_, new_n134_, new_n138_ );
nand g034 ( new_n140_, new_n133_, new_n139_ );
xnor g035 ( new_n141_, new_n140_, new_n126_ );
not g036 ( new_n142_, keyIn_0_6 );
not g037 ( new_n143_, keyIn_0_0 );
xnor g038 ( new_n144_, N1, N5 );
xnor g039 ( new_n145_, new_n144_, new_n143_ );
xnor g040 ( new_n146_, N9, N13 );
xnor g041 ( new_n147_, new_n146_, keyIn_0_1 );
xnor g042 ( new_n148_, new_n145_, new_n147_ );
nand g043 ( new_n149_, new_n148_, new_n142_ );
xnor g044 ( new_n150_, new_n144_, keyIn_0_0 );
xnor g045 ( new_n151_, new_n150_, new_n147_ );
nand g046 ( new_n152_, new_n151_, keyIn_0_6 );
nand g047 ( new_n153_, new_n149_, new_n152_ );
xnor g048 ( new_n154_, new_n153_, new_n141_ );
nand g049 ( new_n155_, new_n154_, new_n125_ );
xnor g050 ( new_n156_, new_n140_, keyIn_0_7 );
xnor g051 ( new_n157_, new_n153_, new_n156_ );
nand g052 ( new_n158_, new_n157_, keyIn_0_10 );
nand g053 ( new_n159_, new_n158_, new_n155_ );
nand g054 ( new_n160_, N135, N137 );
not g055 ( new_n161_, new_n160_ );
nand g056 ( new_n162_, new_n159_, new_n161_ );
xnor g057 ( new_n163_, new_n154_, keyIn_0_10 );
nand g058 ( new_n164_, new_n163_, new_n160_ );
nand g059 ( new_n165_, new_n164_, new_n162_ );
nand g060 ( new_n166_, new_n165_, new_n124_ );
xnor g061 ( new_n167_, new_n159_, new_n160_ );
nand g062 ( new_n168_, new_n167_, keyIn_0_12 );
nand g063 ( new_n169_, new_n168_, new_n166_ );
xnor g064 ( new_n170_, N105, N121 );
xnor g065 ( new_n171_, N73, N89 );
xnor g066 ( new_n172_, new_n170_, new_n171_ );
nand g067 ( new_n173_, new_n169_, new_n172_ );
xnor g068 ( new_n174_, new_n165_, keyIn_0_12 );
not g069 ( new_n175_, new_n172_ );
nand g070 ( new_n176_, new_n174_, new_n175_ );
nand g071 ( new_n177_, new_n176_, new_n173_ );
xnor g072 ( new_n178_, new_n177_, new_n123_ );
not g073 ( new_n179_, keyIn_0_8 );
not g074 ( new_n180_, keyIn_0_4 );
xnor g075 ( new_n181_, N49, N53 );
xnor g076 ( new_n182_, new_n181_, new_n180_ );
not g077 ( new_n183_, keyIn_0_5 );
not g078 ( new_n184_, N61 );
nand g079 ( new_n185_, new_n184_, N57 );
not g080 ( new_n186_, N57 );
nand g081 ( new_n187_, new_n186_, N61 );
nand g082 ( new_n188_, new_n185_, new_n187_ );
nand g083 ( new_n189_, new_n188_, new_n183_ );
xnor g084 ( new_n190_, N57, N61 );
nand g085 ( new_n191_, new_n190_, keyIn_0_5 );
nand g086 ( new_n192_, new_n189_, new_n191_ );
nand g087 ( new_n193_, new_n182_, new_n192_ );
xnor g088 ( new_n194_, new_n181_, keyIn_0_4 );
xnor g089 ( new_n195_, new_n190_, new_n183_ );
nand g090 ( new_n196_, new_n194_, new_n195_ );
nand g091 ( new_n197_, new_n196_, new_n193_ );
xnor g092 ( new_n198_, new_n197_, new_n179_ );
xnor g093 ( new_n199_, N25, N29 );
xnor g094 ( new_n200_, N17, N21 );
xnor g095 ( new_n201_, new_n199_, new_n200_ );
xnor g096 ( new_n202_, new_n198_, new_n201_ );
nand g097 ( new_n203_, N136, N137 );
xnor g098 ( new_n204_, new_n202_, new_n203_ );
xor g099 ( new_n205_, N109, N125 );
xnor g100 ( new_n206_, N77, N93 );
xnor g101 ( new_n207_, new_n205_, new_n206_ );
xnor g102 ( new_n208_, new_n204_, new_n207_ );
not g103 ( new_n209_, new_n208_ );
nor g104 ( new_n210_, new_n178_, new_n209_ );
xor g105 ( new_n211_, N121, N125 );
xnor g106 ( new_n212_, N113, N117 );
xnor g107 ( new_n213_, new_n211_, new_n212_ );
xor g108 ( new_n214_, N105, N109 );
xnor g109 ( new_n215_, N97, N101 );
xnor g110 ( new_n216_, new_n214_, new_n215_ );
xor g111 ( new_n217_, new_n213_, new_n216_ );
nand g112 ( new_n218_, N130, N137 );
xnor g113 ( new_n219_, new_n217_, new_n218_ );
xor g114 ( new_n220_, N37, N53 );
xnor g115 ( new_n221_, N5, N21 );
xnor g116 ( new_n222_, new_n220_, new_n221_ );
xnor g117 ( new_n223_, new_n219_, new_n222_ );
not g118 ( new_n224_, new_n223_ );
nor g119 ( new_n225_, new_n224_, new_n120_ );
xor g120 ( new_n226_, new_n110_, new_n216_ );
nand g121 ( new_n227_, N131, N137 );
xnor g122 ( new_n228_, new_n226_, new_n227_ );
xor g123 ( new_n229_, N41, N57 );
xnor g124 ( new_n230_, N9, N25 );
xnor g125 ( new_n231_, new_n229_, new_n230_ );
xnor g126 ( new_n232_, new_n228_, new_n231_ );
nand g127 ( new_n233_, new_n225_, new_n232_ );
nor g128 ( new_n234_, new_n121_, new_n223_ );
nand g129 ( new_n235_, new_n234_, new_n232_ );
nand g130 ( new_n236_, new_n233_, new_n235_ );
xor g131 ( new_n237_, new_n113_, new_n213_ );
nand g132 ( new_n238_, N132, N137 );
xnor g133 ( new_n239_, new_n237_, new_n238_ );
xor g134 ( new_n240_, N45, N61 );
xnor g135 ( new_n241_, N13, N29 );
xnor g136 ( new_n242_, new_n240_, new_n241_ );
xor g137 ( new_n243_, new_n239_, new_n242_ );
not g138 ( new_n244_, new_n243_ );
nand g139 ( new_n245_, new_n236_, new_n244_ );
xnor g140 ( new_n246_, new_n243_, new_n232_ );
nor g141 ( new_n247_, new_n121_, new_n224_ );
nand g142 ( new_n248_, new_n246_, new_n247_ );
nand g143 ( new_n249_, new_n245_, new_n248_ );
xnor g144 ( new_n250_, new_n249_, keyIn_0_17 );
nand g145 ( new_n251_, new_n210_, new_n250_ );
not g146 ( new_n252_, keyIn_0_11 );
not g147 ( new_n253_, keyIn_0_9 );
nand g148 ( new_n254_, new_n197_, keyIn_0_8 );
xnor g149 ( new_n255_, new_n194_, new_n192_ );
nand g150 ( new_n256_, new_n255_, new_n179_ );
nand g151 ( new_n257_, new_n256_, new_n254_ );
nand g152 ( new_n258_, new_n141_, new_n257_ );
nand g153 ( new_n259_, new_n156_, new_n198_ );
nand g154 ( new_n260_, new_n259_, new_n258_ );
nand g155 ( new_n261_, new_n260_, new_n253_ );
xnor g156 ( new_n262_, new_n156_, new_n257_ );
nand g157 ( new_n263_, new_n262_, keyIn_0_9 );
nand g158 ( new_n264_, new_n263_, new_n261_ );
nand g159 ( new_n265_, N134, N137 );
nand g160 ( new_n266_, new_n264_, new_n265_ );
xnor g161 ( new_n267_, new_n260_, keyIn_0_9 );
not g162 ( new_n268_, new_n265_ );
nand g163 ( new_n269_, new_n267_, new_n268_ );
nand g164 ( new_n270_, new_n269_, new_n266_ );
nand g165 ( new_n271_, new_n270_, new_n252_ );
xnor g166 ( new_n272_, new_n264_, new_n268_ );
nand g167 ( new_n273_, new_n272_, keyIn_0_11 );
nand g168 ( new_n274_, new_n273_, new_n271_ );
xnor g169 ( new_n275_, N101, N117 );
xnor g170 ( new_n276_, N69, N85 );
xnor g171 ( new_n277_, new_n275_, new_n276_ );
nand g172 ( new_n278_, new_n274_, new_n277_ );
xnor g173 ( new_n279_, new_n270_, keyIn_0_11 );
not g174 ( new_n280_, new_n277_ );
nand g175 ( new_n281_, new_n279_, new_n280_ );
nand g176 ( new_n282_, new_n281_, new_n278_ );
xnor g177 ( new_n283_, new_n282_, keyIn_0_13 );
nand g178 ( new_n284_, new_n283_, keyIn_0_15 );
not g179 ( new_n285_, keyIn_0_15 );
not g180 ( new_n286_, keyIn_0_13 );
nand g181 ( new_n287_, new_n282_, new_n286_ );
xnor g182 ( new_n288_, new_n274_, new_n280_ );
nand g183 ( new_n289_, new_n288_, keyIn_0_13 );
nand g184 ( new_n290_, new_n289_, new_n287_ );
nand g185 ( new_n291_, new_n290_, new_n285_ );
nand g186 ( new_n292_, new_n284_, new_n291_ );
xor g187 ( new_n293_, new_n153_, new_n201_ );
nand g188 ( new_n294_, N133, N137 );
xnor g189 ( new_n295_, new_n293_, new_n294_ );
xor g190 ( new_n296_, N97, N113 );
xnor g191 ( new_n297_, N65, N81 );
xnor g192 ( new_n298_, new_n296_, new_n297_ );
xnor g193 ( new_n299_, new_n295_, new_n298_ );
not g194 ( new_n300_, new_n299_ );
nand g195 ( new_n301_, new_n292_, new_n300_ );
nor g196 ( new_n302_, new_n301_, new_n251_ );
nand g197 ( new_n303_, new_n302_, new_n122_ );
xnor g198 ( new_n304_, new_n177_, keyIn_0_14 );
nand g199 ( new_n305_, new_n304_, new_n208_ );
not g200 ( new_n306_, new_n250_ );
nor g201 ( new_n307_, new_n305_, new_n306_ );
xnor g202 ( new_n308_, new_n290_, keyIn_0_15 );
nor g203 ( new_n309_, new_n308_, new_n299_ );
nand g204 ( new_n310_, new_n309_, new_n307_ );
nand g205 ( new_n311_, new_n310_, keyIn_0_18 );
nand g206 ( new_n312_, new_n311_, new_n303_ );
nand g207 ( new_n313_, new_n312_, new_n121_ );
nand g208 ( new_n314_, new_n313_, keyIn_0_20 );
not g209 ( new_n315_, keyIn_0_20 );
xnor g210 ( new_n316_, new_n302_, keyIn_0_18 );
nor g211 ( new_n317_, new_n316_, new_n120_ );
nand g212 ( new_n318_, new_n317_, new_n315_ );
nand g213 ( new_n319_, new_n318_, new_n314_ );
nand g214 ( new_n320_, new_n319_, new_n107_ );
xnor g215 ( new_n321_, new_n313_, new_n315_ );
nand g216 ( new_n322_, new_n321_, N1 );
nand g217 ( new_n323_, new_n322_, new_n320_ );
xnor g218 ( N724, new_n323_, new_n106_ );
not g219 ( new_n325_, keyIn_0_27 );
nand g220 ( new_n326_, new_n312_, new_n224_ );
nand g221 ( new_n327_, new_n326_, keyIn_0_21 );
not g222 ( new_n328_, keyIn_0_21 );
nor g223 ( new_n329_, new_n316_, new_n223_ );
nand g224 ( new_n330_, new_n329_, new_n328_ );
nand g225 ( new_n331_, new_n330_, new_n327_ );
nand g226 ( new_n332_, new_n331_, N5 );
not g227 ( new_n333_, N5 );
xnor g228 ( new_n334_, new_n326_, new_n328_ );
nand g229 ( new_n335_, new_n334_, new_n333_ );
nand g230 ( new_n336_, new_n335_, new_n332_ );
xnor g231 ( N725, new_n336_, new_n325_ );
not g232 ( new_n338_, N9 );
not g233 ( new_n339_, new_n232_ );
nand g234 ( new_n340_, new_n312_, new_n339_ );
nand g235 ( new_n341_, new_n340_, keyIn_0_22 );
not g236 ( new_n342_, keyIn_0_22 );
nor g237 ( new_n343_, new_n316_, new_n232_ );
nand g238 ( new_n344_, new_n343_, new_n342_ );
nand g239 ( new_n345_, new_n344_, new_n341_ );
nand g240 ( new_n346_, new_n345_, new_n338_ );
xnor g241 ( new_n347_, new_n340_, new_n342_ );
nand g242 ( new_n348_, new_n347_, N9 );
nand g243 ( new_n349_, new_n348_, new_n346_ );
xnor g244 ( N726, new_n349_, keyIn_0_28 );
not g245 ( new_n351_, keyIn_0_29 );
not g246 ( new_n352_, N13 );
nand g247 ( new_n353_, new_n312_, new_n243_ );
nand g248 ( new_n354_, new_n353_, keyIn_0_23 );
not g249 ( new_n355_, keyIn_0_23 );
nor g250 ( new_n356_, new_n316_, new_n244_ );
nand g251 ( new_n357_, new_n356_, new_n355_ );
nand g252 ( new_n358_, new_n357_, new_n354_ );
nand g253 ( new_n359_, new_n358_, new_n352_ );
xnor g254 ( new_n360_, new_n353_, new_n355_ );
nand g255 ( new_n361_, new_n360_, N13 );
nand g256 ( new_n362_, new_n361_, new_n359_ );
xnor g257 ( N727, new_n362_, new_n351_ );
nor g258 ( new_n364_, new_n283_, new_n299_ );
nand g259 ( new_n365_, new_n250_, new_n209_ );
nor g260 ( new_n366_, new_n304_, new_n365_ );
nand g261 ( new_n367_, new_n366_, new_n364_ );
xnor g262 ( new_n368_, new_n367_, keyIn_0_19 );
nor g263 ( new_n369_, new_n368_, new_n120_ );
xor g264 ( N728, new_n369_, N17 );
not g265 ( new_n371_, keyIn_0_30 );
not g266 ( new_n372_, keyIn_0_24 );
nor g267 ( new_n373_, new_n368_, new_n223_ );
xnor g268 ( new_n374_, new_n373_, new_n372_ );
xnor g269 ( new_n375_, new_n374_, N21 );
xnor g270 ( N729, new_n375_, new_n371_ );
nor g271 ( new_n377_, new_n368_, new_n232_ );
xor g272 ( N730, new_n377_, N25 );
nor g273 ( new_n379_, new_n368_, new_n244_ );
xnor g274 ( new_n380_, new_n379_, keyIn_0_25 );
xnor g275 ( new_n381_, new_n380_, N29 );
xnor g276 ( N731, new_n381_, keyIn_0_31 );
nor g277 ( new_n383_, new_n290_, new_n300_ );
not g278 ( new_n384_, new_n383_ );
nor g279 ( new_n385_, new_n251_, new_n384_ );
nand g280 ( new_n386_, new_n385_, new_n121_ );
xnor g281 ( N732, new_n386_, N33 );
nand g282 ( new_n388_, new_n385_, new_n224_ );
xnor g283 ( N733, new_n388_, N37 );
nand g284 ( new_n390_, new_n385_, new_n339_ );
xnor g285 ( N734, new_n390_, N41 );
nand g286 ( new_n392_, new_n385_, new_n243_ );
xnor g287 ( N735, new_n392_, N45 );
nand g288 ( new_n394_, new_n383_, new_n178_ );
nor g289 ( new_n395_, new_n394_, new_n365_ );
nand g290 ( new_n396_, new_n395_, new_n121_ );
xnor g291 ( N736, new_n396_, N49 );
nand g292 ( new_n398_, new_n395_, new_n224_ );
xnor g293 ( N737, new_n398_, N53 );
nand g294 ( new_n400_, new_n395_, new_n339_ );
xnor g295 ( N738, new_n400_, N57 );
nand g296 ( new_n402_, new_n395_, new_n243_ );
xnor g297 ( N739, new_n402_, N61 );
not g298 ( new_n404_, keyIn_0_16 );
nand g299 ( new_n405_, new_n178_, new_n404_ );
not g300 ( new_n406_, new_n364_ );
nor g301 ( new_n407_, new_n178_, new_n404_ );
nor g302 ( new_n408_, new_n406_, new_n407_ );
nand g303 ( new_n409_, new_n408_, new_n405_ );
nand g304 ( new_n410_, new_n409_, new_n394_ );
nand g305 ( new_n411_, new_n410_, new_n208_ );
nand g306 ( new_n412_, new_n178_, new_n209_ );
nand g307 ( new_n413_, new_n305_, new_n412_ );
nor g308 ( new_n414_, new_n283_, new_n300_ );
nand g309 ( new_n415_, new_n413_, new_n414_ );
nand g310 ( new_n416_, new_n411_, new_n415_ );
not g311 ( new_n417_, new_n225_ );
nand g312 ( new_n418_, new_n244_, new_n339_ );
nor g313 ( new_n419_, new_n417_, new_n418_ );
nand g314 ( new_n420_, new_n416_, new_n419_ );
not g315 ( new_n421_, new_n420_ );
nand g316 ( new_n422_, new_n421_, new_n300_ );
xnor g317 ( N740, new_n422_, N65 );
nand g318 ( new_n424_, new_n421_, new_n283_ );
xnor g319 ( N741, new_n424_, N69 );
nand g320 ( new_n426_, new_n421_, new_n304_ );
xnor g321 ( N742, new_n426_, N73 );
nand g322 ( new_n428_, new_n421_, new_n209_ );
xnor g323 ( N743, new_n428_, N77 );
nand g324 ( new_n430_, new_n416_, new_n243_ );
nor g325 ( new_n431_, new_n430_, new_n233_ );
nand g326 ( new_n432_, new_n431_, new_n300_ );
xnor g327 ( N744, new_n432_, N81 );
nand g328 ( new_n434_, new_n431_, new_n283_ );
xnor g329 ( N745, new_n434_, N85 );
nand g330 ( new_n436_, new_n431_, new_n304_ );
xnor g331 ( N746, new_n436_, N89 );
nand g332 ( new_n438_, new_n431_, new_n209_ );
xnor g333 ( N747, new_n438_, N93 );
not g334 ( new_n440_, new_n234_ );
nor g335 ( new_n441_, new_n440_, new_n418_ );
nand g336 ( new_n442_, new_n416_, new_n441_ );
not g337 ( new_n443_, new_n442_ );
nand g338 ( new_n444_, new_n443_, new_n300_ );
xnor g339 ( N748, new_n444_, N97 );
nand g340 ( new_n446_, new_n443_, new_n283_ );
xnor g341 ( N749, new_n446_, N101 );
nand g342 ( new_n448_, new_n443_, new_n304_ );
xnor g343 ( N750, new_n448_, N105 );
nand g344 ( new_n450_, new_n443_, new_n209_ );
xnor g345 ( N751, new_n450_, N109 );
nor g346 ( new_n452_, new_n430_, new_n235_ );
nand g347 ( new_n453_, new_n452_, new_n300_ );
xnor g348 ( N752, new_n453_, N113 );
nand g349 ( new_n455_, new_n452_, new_n283_ );
xnor g350 ( N753, new_n455_, N117 );
nand g351 ( new_n457_, new_n452_, new_n304_ );
xnor g352 ( N754, new_n457_, N121 );
nand g353 ( new_n459_, new_n452_, new_n209_ );
xnor g354 ( N755, new_n459_, N125 );
endmodule