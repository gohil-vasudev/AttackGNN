module add_mul_8_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, 
        b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, operation, Result_0_, 
        Result_1_, Result_2_, Result_3_, Result_4_, Result_5_, Result_6_, 
        Result_7_, Result_8_, Result_9_, Result_10_, Result_11_, Result_12_, 
        Result_13_, Result_14_, Result_15_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_,
         b_4_, b_5_, b_6_, b_7_, operation;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_;
  wire   n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935;

  OR2_X1 U478 ( .A1(n462), .A2(n463), .ZN(Result_9_) );
  AND2_X1 U479 ( .A1(n464), .A2(operation), .ZN(n463) );
  XNOR2_X1 U480 ( .A(n465), .B(n466), .ZN(n464) );
  XOR2_X1 U481 ( .A(n467), .B(n468), .Z(n466) );
  AND2_X1 U482 ( .A1(n469), .A2(n470), .ZN(n462) );
  OR3_X1 U483 ( .A1(n471), .A2(n472), .A3(n473), .ZN(n469) );
  INV_X1 U484 ( .A(n474), .ZN(n473) );
  OR2_X1 U485 ( .A1(n475), .A2(n476), .ZN(n474) );
  AND2_X1 U486 ( .A1(n477), .A2(n478), .ZN(n472) );
  XOR2_X1 U487 ( .A(n479), .B(n476), .Z(n477) );
  AND3_X1 U488 ( .A1(n476), .A2(n479), .A3(b_1_), .ZN(n471) );
  OR2_X1 U489 ( .A1(n480), .A2(n481), .ZN(Result_8_) );
  AND2_X1 U490 ( .A1(n482), .A2(operation), .ZN(n481) );
  XNOR2_X1 U491 ( .A(n483), .B(n484), .ZN(n482) );
  XOR2_X1 U492 ( .A(n485), .B(n486), .Z(n484) );
  AND2_X1 U493 ( .A1(n487), .A2(n470), .ZN(n480) );
  XOR2_X1 U494 ( .A(n488), .B(n489), .Z(n487) );
  XOR2_X1 U495 ( .A(n490), .B(b_0_), .Z(n489) );
  OR2_X1 U496 ( .A1(n491), .A2(n492), .ZN(n488) );
  AND2_X1 U497 ( .A1(n479), .A2(n478), .ZN(n492) );
  AND2_X1 U498 ( .A1(n476), .A2(n475), .ZN(n491) );
  OR2_X1 U499 ( .A1(n493), .A2(n494), .ZN(n476) );
  AND2_X1 U500 ( .A1(n495), .A2(n496), .ZN(n493) );
  AND2_X1 U501 ( .A1(operation), .A2(n497), .ZN(Result_7_) );
  XOR2_X1 U502 ( .A(n498), .B(n499), .Z(n497) );
  AND3_X1 U503 ( .A1(n500), .A2(n501), .A3(operation), .ZN(Result_6_) );
  OR2_X1 U504 ( .A1(n502), .A2(n503), .ZN(n500) );
  XOR2_X1 U505 ( .A(n504), .B(n505), .Z(n503) );
  INV_X1 U506 ( .A(n506), .ZN(n502) );
  OR2_X1 U507 ( .A1(n498), .A2(n499), .ZN(n506) );
  AND2_X1 U508 ( .A1(operation), .A2(n507), .ZN(Result_5_) );
  XOR2_X1 U509 ( .A(n508), .B(n509), .Z(n507) );
  AND2_X1 U510 ( .A1(operation), .A2(n510), .ZN(Result_4_) );
  XNOR2_X1 U511 ( .A(n511), .B(n512), .ZN(n510) );
  AND2_X1 U512 ( .A1(n513), .A2(n514), .ZN(n511) );
  AND2_X1 U513 ( .A1(operation), .A2(n515), .ZN(Result_3_) );
  XOR2_X1 U514 ( .A(n516), .B(n517), .Z(n515) );
  AND2_X1 U515 ( .A1(n518), .A2(n519), .ZN(n517) );
  OR2_X1 U516 ( .A1(n520), .A2(n521), .ZN(n519) );
  AND2_X1 U517 ( .A1(n522), .A2(n523), .ZN(n521) );
  INV_X1 U518 ( .A(n524), .ZN(n518) );
  AND2_X1 U519 ( .A1(n525), .A2(operation), .ZN(Result_2_) );
  XOR2_X1 U520 ( .A(n526), .B(n527), .Z(n525) );
  AND2_X1 U521 ( .A1(operation), .A2(n528), .ZN(Result_1_) );
  XOR2_X1 U522 ( .A(n529), .B(n530), .Z(n528) );
  AND2_X1 U523 ( .A1(n531), .A2(n532), .ZN(n530) );
  OR2_X1 U524 ( .A1(n533), .A2(n534), .ZN(n532) );
  AND2_X1 U525 ( .A1(n535), .A2(n536), .ZN(n533) );
  INV_X1 U526 ( .A(n537), .ZN(n531) );
  OR2_X1 U527 ( .A1(n538), .A2(n539), .ZN(Result_15_) );
  AND3_X1 U528 ( .A1(b_7_), .A2(a_7_), .A3(operation), .ZN(n539) );
  AND2_X1 U529 ( .A1(n540), .A2(n470), .ZN(n538) );
  XOR2_X1 U530 ( .A(b_7_), .B(a_7_), .Z(n540) );
  OR2_X1 U531 ( .A1(n541), .A2(n542), .ZN(Result_14_) );
  AND2_X1 U532 ( .A1(n543), .A2(operation), .ZN(n542) );
  XNOR2_X1 U533 ( .A(n544), .B(n545), .ZN(n543) );
  AND2_X1 U534 ( .A1(n546), .A2(n470), .ZN(n541) );
  XOR2_X1 U535 ( .A(n547), .B(n548), .Z(n546) );
  XOR2_X1 U536 ( .A(b_6_), .B(a_6_), .Z(n548) );
  AND2_X1 U537 ( .A1(b_7_), .A2(a_7_), .ZN(n547) );
  OR2_X1 U538 ( .A1(n549), .A2(n550), .ZN(Result_13_) );
  AND2_X1 U539 ( .A1(n551), .A2(operation), .ZN(n550) );
  XNOR2_X1 U540 ( .A(n552), .B(n553), .ZN(n551) );
  XOR2_X1 U541 ( .A(n554), .B(n555), .Z(n553) );
  AND2_X1 U542 ( .A1(n556), .A2(n470), .ZN(n549) );
  OR3_X1 U543 ( .A1(n557), .A2(n558), .A3(n559), .ZN(n556) );
  AND2_X1 U544 ( .A1(n560), .A2(n561), .ZN(n559) );
  INV_X1 U545 ( .A(n562), .ZN(n560) );
  AND2_X1 U546 ( .A1(n563), .A2(n564), .ZN(n558) );
  XOR2_X1 U547 ( .A(n561), .B(a_5_), .Z(n563) );
  AND3_X1 U548 ( .A1(n565), .A2(n566), .A3(b_5_), .ZN(n557) );
  OR2_X1 U549 ( .A1(n567), .A2(n568), .ZN(Result_12_) );
  AND2_X1 U550 ( .A1(n569), .A2(operation), .ZN(n568) );
  XNOR2_X1 U551 ( .A(n570), .B(n571), .ZN(n569) );
  XOR2_X1 U552 ( .A(n572), .B(n573), .Z(n571) );
  AND2_X1 U553 ( .A1(n574), .A2(n470), .ZN(n567) );
  XNOR2_X1 U554 ( .A(n575), .B(n576), .ZN(n574) );
  AND2_X1 U555 ( .A1(n577), .A2(n578), .ZN(n576) );
  OR2_X1 U556 ( .A1(n579), .A2(n580), .ZN(Result_11_) );
  AND2_X1 U557 ( .A1(n581), .A2(operation), .ZN(n580) );
  XNOR2_X1 U558 ( .A(n582), .B(n583), .ZN(n581) );
  XOR2_X1 U559 ( .A(n584), .B(n585), .Z(n583) );
  AND2_X1 U560 ( .A1(n586), .A2(n470), .ZN(n579) );
  OR3_X1 U561 ( .A1(n587), .A2(n588), .A3(n589), .ZN(n586) );
  INV_X1 U562 ( .A(n590), .ZN(n589) );
  OR2_X1 U563 ( .A1(n591), .A2(n592), .ZN(n590) );
  AND2_X1 U564 ( .A1(n593), .A2(n594), .ZN(n588) );
  XOR2_X1 U565 ( .A(n595), .B(n591), .Z(n593) );
  AND3_X1 U566 ( .A1(n591), .A2(n595), .A3(b_3_), .ZN(n587) );
  OR2_X1 U567 ( .A1(n596), .A2(n597), .ZN(Result_10_) );
  AND2_X1 U568 ( .A1(n598), .A2(operation), .ZN(n597) );
  XNOR2_X1 U569 ( .A(n599), .B(n600), .ZN(n598) );
  XOR2_X1 U570 ( .A(n601), .B(n602), .Z(n600) );
  AND2_X1 U571 ( .A1(n603), .A2(n470), .ZN(n596) );
  INV_X1 U572 ( .A(operation), .ZN(n470) );
  XOR2_X1 U573 ( .A(n495), .B(n604), .Z(n603) );
  OR2_X1 U574 ( .A1(n494), .A2(n605), .ZN(n604) );
  AND2_X1 U575 ( .A1(n606), .A2(n607), .ZN(n494) );
  OR2_X1 U576 ( .A1(n608), .A2(n609), .ZN(n495) );
  AND2_X1 U577 ( .A1(n595), .A2(n594), .ZN(n609) );
  AND2_X1 U578 ( .A1(n591), .A2(n592), .ZN(n608) );
  OR2_X1 U579 ( .A1(n610), .A2(n611), .ZN(n591) );
  INV_X1 U580 ( .A(n578), .ZN(n611) );
  OR2_X1 U581 ( .A1(a_4_), .A2(b_4_), .ZN(n578) );
  AND2_X1 U582 ( .A1(n575), .A2(n577), .ZN(n610) );
  OR2_X1 U583 ( .A1(n612), .A2(n613), .ZN(n575) );
  AND2_X1 U584 ( .A1(n566), .A2(n564), .ZN(n613) );
  AND2_X1 U585 ( .A1(n565), .A2(n562), .ZN(n612) );
  INV_X1 U586 ( .A(n561), .ZN(n565) );
  OR3_X1 U587 ( .A1(n614), .A2(n615), .A3(n616), .ZN(n561) );
  AND2_X1 U588 ( .A1(b_6_), .A2(a_6_), .ZN(n616) );
  AND2_X1 U589 ( .A1(n617), .A2(a_7_), .ZN(n615) );
  INV_X1 U590 ( .A(n544), .ZN(n617) );
  AND2_X1 U591 ( .A1(b_7_), .A2(n545), .ZN(n614) );
  AND2_X1 U592 ( .A1(operation), .A2(n618), .ZN(Result_0_) );
  OR3_X1 U593 ( .A1(n537), .A2(n619), .A3(n620), .ZN(n618) );
  AND2_X1 U594 ( .A1(n621), .A2(a_0_), .ZN(n620) );
  AND2_X1 U595 ( .A1(n529), .A2(n534), .ZN(n619) );
  AND2_X1 U596 ( .A1(n526), .A2(n527), .ZN(n529) );
  XOR2_X1 U597 ( .A(n536), .B(n535), .Z(n527) );
  OR2_X1 U598 ( .A1(n622), .A2(n623), .ZN(n526) );
  INV_X1 U599 ( .A(n624), .ZN(n623) );
  OR2_X1 U600 ( .A1(n625), .A2(n524), .ZN(n622) );
  AND3_X1 U601 ( .A1(n523), .A2(n522), .A3(n520), .ZN(n524) );
  AND2_X1 U602 ( .A1(n516), .A2(n520), .ZN(n625) );
  AND2_X1 U603 ( .A1(n626), .A2(n624), .ZN(n520) );
  OR2_X1 U604 ( .A1(n627), .A2(n628), .ZN(n624) );
  INV_X1 U605 ( .A(n629), .ZN(n626) );
  AND2_X1 U606 ( .A1(n627), .A2(n628), .ZN(n629) );
  OR2_X1 U607 ( .A1(n630), .A2(n631), .ZN(n628) );
  AND2_X1 U608 ( .A1(n632), .A2(n633), .ZN(n631) );
  AND2_X1 U609 ( .A1(n634), .A2(n635), .ZN(n630) );
  OR2_X1 U610 ( .A1(n633), .A2(n632), .ZN(n635) );
  XOR2_X1 U611 ( .A(n636), .B(n637), .Z(n627) );
  XOR2_X1 U612 ( .A(n638), .B(n639), .Z(n637) );
  AND2_X1 U613 ( .A1(n640), .A2(n512), .ZN(n516) );
  XOR2_X1 U614 ( .A(n523), .B(n522), .Z(n512) );
  INV_X1 U615 ( .A(n641), .ZN(n522) );
  OR2_X1 U616 ( .A1(n642), .A2(n643), .ZN(n641) );
  AND2_X1 U617 ( .A1(n644), .A2(n645), .ZN(n643) );
  AND2_X1 U618 ( .A1(n646), .A2(n647), .ZN(n642) );
  OR2_X1 U619 ( .A1(n645), .A2(n644), .ZN(n647) );
  XOR2_X1 U620 ( .A(n648), .B(n634), .Z(n523) );
  XOR2_X1 U621 ( .A(n649), .B(n650), .Z(n634) );
  XOR2_X1 U622 ( .A(n651), .B(n652), .Z(n650) );
  XNOR2_X1 U623 ( .A(n633), .B(n632), .ZN(n648) );
  OR2_X1 U624 ( .A1(n653), .A2(n654), .ZN(n632) );
  AND2_X1 U625 ( .A1(n655), .A2(n656), .ZN(n654) );
  AND2_X1 U626 ( .A1(n657), .A2(n658), .ZN(n653) );
  OR2_X1 U627 ( .A1(n656), .A2(n655), .ZN(n658) );
  OR2_X1 U628 ( .A1(n594), .A2(n490), .ZN(n633) );
  OR2_X1 U629 ( .A1(n659), .A2(n660), .ZN(n640) );
  INV_X1 U630 ( .A(n513), .ZN(n660) );
  OR2_X1 U631 ( .A1(n508), .A2(n509), .ZN(n513) );
  OR2_X1 U632 ( .A1(n661), .A2(n659), .ZN(n509) );
  AND2_X1 U633 ( .A1(n662), .A2(n663), .ZN(n661) );
  AND2_X1 U634 ( .A1(n501), .A2(n664), .ZN(n508) );
  OR4_X1 U635 ( .A1(n499), .A2(n498), .A3(n665), .A4(n666), .ZN(n501) );
  AND2_X1 U636 ( .A1(n504), .A2(n505), .ZN(n666) );
  INV_X1 U637 ( .A(n664), .ZN(n665) );
  OR2_X1 U638 ( .A1(n504), .A2(n505), .ZN(n664) );
  OR2_X1 U639 ( .A1(n667), .A2(n668), .ZN(n505) );
  AND2_X1 U640 ( .A1(n669), .A2(n670), .ZN(n668) );
  AND2_X1 U641 ( .A1(n671), .A2(n672), .ZN(n667) );
  OR2_X1 U642 ( .A1(n670), .A2(n669), .ZN(n672) );
  XOR2_X1 U643 ( .A(n673), .B(n674), .Z(n504) );
  XOR2_X1 U644 ( .A(n675), .B(n676), .Z(n674) );
  OR2_X1 U645 ( .A1(n677), .A2(n678), .ZN(n498) );
  AND2_X1 U646 ( .A1(n486), .A2(n485), .ZN(n678) );
  AND2_X1 U647 ( .A1(n483), .A2(n679), .ZN(n677) );
  OR2_X1 U648 ( .A1(n485), .A2(n486), .ZN(n679) );
  OR2_X1 U649 ( .A1(n680), .A2(n490), .ZN(n486) );
  OR2_X1 U650 ( .A1(n681), .A2(n682), .ZN(n485) );
  AND2_X1 U651 ( .A1(n468), .A2(n467), .ZN(n682) );
  AND2_X1 U652 ( .A1(n465), .A2(n683), .ZN(n681) );
  OR2_X1 U653 ( .A1(n467), .A2(n468), .ZN(n683) );
  OR2_X1 U654 ( .A1(n680), .A2(n479), .ZN(n468) );
  OR2_X1 U655 ( .A1(n684), .A2(n685), .ZN(n467) );
  AND2_X1 U656 ( .A1(n602), .A2(n601), .ZN(n685) );
  AND2_X1 U657 ( .A1(n599), .A2(n686), .ZN(n684) );
  OR2_X1 U658 ( .A1(n602), .A2(n601), .ZN(n686) );
  OR2_X1 U659 ( .A1(n687), .A2(n688), .ZN(n601) );
  AND2_X1 U660 ( .A1(n585), .A2(n584), .ZN(n688) );
  AND2_X1 U661 ( .A1(n582), .A2(n689), .ZN(n687) );
  OR2_X1 U662 ( .A1(n585), .A2(n584), .ZN(n689) );
  OR2_X1 U663 ( .A1(n690), .A2(n691), .ZN(n584) );
  AND2_X1 U664 ( .A1(n573), .A2(n572), .ZN(n691) );
  AND2_X1 U665 ( .A1(n570), .A2(n692), .ZN(n690) );
  OR2_X1 U666 ( .A1(n573), .A2(n572), .ZN(n692) );
  OR2_X1 U667 ( .A1(n693), .A2(n694), .ZN(n572) );
  AND2_X1 U668 ( .A1(n555), .A2(n554), .ZN(n694) );
  AND2_X1 U669 ( .A1(n552), .A2(n695), .ZN(n693) );
  OR2_X1 U670 ( .A1(n555), .A2(n554), .ZN(n695) );
  OR2_X1 U671 ( .A1(n696), .A2(n544), .ZN(n554) );
  OR2_X1 U672 ( .A1(n697), .A2(n680), .ZN(n544) );
  OR2_X1 U673 ( .A1(n566), .A2(n680), .ZN(n555) );
  XNOR2_X1 U674 ( .A(n698), .B(n699), .ZN(n552) );
  OR2_X1 U675 ( .A1(n697), .A2(n700), .ZN(n698) );
  OR2_X1 U676 ( .A1(n701), .A2(n680), .ZN(n573) );
  XOR2_X1 U677 ( .A(n702), .B(n703), .Z(n570) );
  XOR2_X1 U678 ( .A(n704), .B(n705), .Z(n703) );
  OR2_X1 U679 ( .A1(n595), .A2(n680), .ZN(n585) );
  XOR2_X1 U680 ( .A(n706), .B(n707), .Z(n582) );
  XOR2_X1 U681 ( .A(n708), .B(n709), .Z(n707) );
  OR2_X1 U682 ( .A1(n606), .A2(n680), .ZN(n602) );
  INV_X1 U683 ( .A(b_7_), .ZN(n680) );
  XOR2_X1 U684 ( .A(n710), .B(n711), .Z(n599) );
  XOR2_X1 U685 ( .A(n712), .B(n713), .Z(n711) );
  XOR2_X1 U686 ( .A(n714), .B(n715), .Z(n465) );
  XOR2_X1 U687 ( .A(n716), .B(n717), .Z(n715) );
  XOR2_X1 U688 ( .A(n718), .B(n719), .Z(n483) );
  XOR2_X1 U689 ( .A(n720), .B(n721), .Z(n719) );
  XOR2_X1 U690 ( .A(n671), .B(n722), .Z(n499) );
  XOR2_X1 U691 ( .A(n670), .B(n669), .Z(n722) );
  OR2_X1 U692 ( .A1(n700), .A2(n490), .ZN(n669) );
  OR2_X1 U693 ( .A1(n723), .A2(n724), .ZN(n670) );
  AND2_X1 U694 ( .A1(n721), .A2(n720), .ZN(n724) );
  AND2_X1 U695 ( .A1(n718), .A2(n725), .ZN(n723) );
  OR2_X1 U696 ( .A1(n720), .A2(n721), .ZN(n725) );
  OR2_X1 U697 ( .A1(n700), .A2(n479), .ZN(n721) );
  OR2_X1 U698 ( .A1(n726), .A2(n727), .ZN(n720) );
  AND2_X1 U699 ( .A1(n717), .A2(n716), .ZN(n727) );
  AND2_X1 U700 ( .A1(n714), .A2(n728), .ZN(n726) );
  OR2_X1 U701 ( .A1(n716), .A2(n717), .ZN(n728) );
  OR2_X1 U702 ( .A1(n700), .A2(n606), .ZN(n717) );
  OR2_X1 U703 ( .A1(n729), .A2(n730), .ZN(n716) );
  AND2_X1 U704 ( .A1(n713), .A2(n712), .ZN(n730) );
  AND2_X1 U705 ( .A1(n710), .A2(n731), .ZN(n729) );
  OR2_X1 U706 ( .A1(n713), .A2(n712), .ZN(n731) );
  OR2_X1 U707 ( .A1(n732), .A2(n733), .ZN(n712) );
  AND2_X1 U708 ( .A1(n709), .A2(n708), .ZN(n733) );
  AND2_X1 U709 ( .A1(n706), .A2(n734), .ZN(n732) );
  OR2_X1 U710 ( .A1(n709), .A2(n708), .ZN(n734) );
  OR2_X1 U711 ( .A1(n735), .A2(n736), .ZN(n708) );
  AND2_X1 U712 ( .A1(n705), .A2(n704), .ZN(n736) );
  AND2_X1 U713 ( .A1(n702), .A2(n737), .ZN(n735) );
  OR2_X1 U714 ( .A1(n705), .A2(n704), .ZN(n737) );
  OR2_X1 U715 ( .A1(n696), .A2(n738), .ZN(n704) );
  INV_X1 U716 ( .A(n545), .ZN(n696) );
  AND2_X1 U717 ( .A1(a_7_), .A2(b_6_), .ZN(n545) );
  OR2_X1 U718 ( .A1(n566), .A2(n700), .ZN(n705) );
  XNOR2_X1 U719 ( .A(n739), .B(n738), .ZN(n702) );
  OR2_X1 U720 ( .A1(n697), .A2(n564), .ZN(n738) );
  OR2_X1 U721 ( .A1(n740), .A2(n741), .ZN(n739) );
  OR2_X1 U722 ( .A1(n701), .A2(n700), .ZN(n709) );
  XOR2_X1 U723 ( .A(n742), .B(n743), .Z(n706) );
  XOR2_X1 U724 ( .A(n744), .B(n562), .Z(n743) );
  OR2_X1 U725 ( .A1(n595), .A2(n700), .ZN(n713) );
  INV_X1 U726 ( .A(b_6_), .ZN(n700) );
  XOR2_X1 U727 ( .A(n745), .B(n746), .Z(n710) );
  XOR2_X1 U728 ( .A(n747), .B(n748), .Z(n746) );
  XOR2_X1 U729 ( .A(n749), .B(n750), .Z(n714) );
  XOR2_X1 U730 ( .A(n751), .B(n752), .Z(n750) );
  XOR2_X1 U731 ( .A(n753), .B(n754), .Z(n718) );
  XOR2_X1 U732 ( .A(n755), .B(n756), .Z(n754) );
  XOR2_X1 U733 ( .A(n757), .B(n758), .Z(n671) );
  XOR2_X1 U734 ( .A(n759), .B(n760), .Z(n758) );
  INV_X1 U735 ( .A(n514), .ZN(n659) );
  OR2_X1 U736 ( .A1(n662), .A2(n663), .ZN(n514) );
  OR2_X1 U737 ( .A1(n761), .A2(n762), .ZN(n663) );
  AND2_X1 U738 ( .A1(n673), .A2(n676), .ZN(n762) );
  AND2_X1 U739 ( .A1(n763), .A2(n675), .ZN(n761) );
  OR2_X1 U740 ( .A1(n764), .A2(n765), .ZN(n675) );
  AND2_X1 U741 ( .A1(n760), .A2(n759), .ZN(n765) );
  AND2_X1 U742 ( .A1(n757), .A2(n766), .ZN(n764) );
  OR2_X1 U743 ( .A1(n759), .A2(n760), .ZN(n766) );
  OR2_X1 U744 ( .A1(n564), .A2(n479), .ZN(n760) );
  OR2_X1 U745 ( .A1(n767), .A2(n768), .ZN(n759) );
  AND2_X1 U746 ( .A1(n756), .A2(n755), .ZN(n768) );
  AND2_X1 U747 ( .A1(n753), .A2(n769), .ZN(n767) );
  OR2_X1 U748 ( .A1(n755), .A2(n756), .ZN(n769) );
  OR2_X1 U749 ( .A1(n564), .A2(n606), .ZN(n756) );
  OR2_X1 U750 ( .A1(n770), .A2(n771), .ZN(n755) );
  AND2_X1 U751 ( .A1(n752), .A2(n751), .ZN(n771) );
  AND2_X1 U752 ( .A1(n749), .A2(n772), .ZN(n770) );
  OR2_X1 U753 ( .A1(n751), .A2(n752), .ZN(n772) );
  OR2_X1 U754 ( .A1(n564), .A2(n595), .ZN(n752) );
  OR2_X1 U755 ( .A1(n773), .A2(n774), .ZN(n751) );
  AND2_X1 U756 ( .A1(n748), .A2(n747), .ZN(n774) );
  AND2_X1 U757 ( .A1(n745), .A2(n775), .ZN(n773) );
  OR2_X1 U758 ( .A1(n748), .A2(n747), .ZN(n775) );
  OR2_X1 U759 ( .A1(n776), .A2(n777), .ZN(n747) );
  AND2_X1 U760 ( .A1(n562), .A2(n744), .ZN(n777) );
  AND2_X1 U761 ( .A1(n778), .A2(n742), .ZN(n776) );
  OR2_X1 U762 ( .A1(n779), .A2(n780), .ZN(n742) );
  AND2_X1 U763 ( .A1(n781), .A2(n782), .ZN(n779) );
  OR2_X1 U764 ( .A1(n562), .A2(n744), .ZN(n778) );
  OR2_X1 U765 ( .A1(n781), .A2(n699), .ZN(n744) );
  OR2_X1 U766 ( .A1(n740), .A2(n564), .ZN(n699) );
  OR2_X1 U767 ( .A1(n566), .A2(n564), .ZN(n562) );
  OR2_X1 U768 ( .A1(n701), .A2(n564), .ZN(n748) );
  XNOR2_X1 U769 ( .A(n783), .B(n784), .ZN(n745) );
  XOR2_X1 U770 ( .A(n785), .B(n780), .Z(n783) );
  INV_X1 U771 ( .A(n786), .ZN(n780) );
  XNOR2_X1 U772 ( .A(n787), .B(n788), .ZN(n749) );
  XNOR2_X1 U773 ( .A(n577), .B(n789), .ZN(n787) );
  XOR2_X1 U774 ( .A(n790), .B(n791), .Z(n753) );
  XOR2_X1 U775 ( .A(n792), .B(n793), .Z(n791) );
  XOR2_X1 U776 ( .A(n794), .B(n795), .Z(n757) );
  XOR2_X1 U777 ( .A(n796), .B(n797), .Z(n795) );
  OR2_X1 U778 ( .A1(n676), .A2(n673), .ZN(n763) );
  XOR2_X1 U779 ( .A(n798), .B(n799), .Z(n673) );
  XOR2_X1 U780 ( .A(n800), .B(n801), .Z(n799) );
  OR2_X1 U781 ( .A1(n564), .A2(n490), .ZN(n676) );
  INV_X1 U782 ( .A(b_5_), .ZN(n564) );
  XOR2_X1 U783 ( .A(n646), .B(n802), .Z(n662) );
  XOR2_X1 U784 ( .A(n645), .B(n644), .Z(n802) );
  OR2_X1 U785 ( .A1(n741), .A2(n490), .ZN(n644) );
  OR2_X1 U786 ( .A1(n803), .A2(n804), .ZN(n645) );
  AND2_X1 U787 ( .A1(n798), .A2(n801), .ZN(n804) );
  AND2_X1 U788 ( .A1(n805), .A2(n800), .ZN(n803) );
  OR2_X1 U789 ( .A1(n806), .A2(n807), .ZN(n800) );
  AND2_X1 U790 ( .A1(n797), .A2(n796), .ZN(n807) );
  AND2_X1 U791 ( .A1(n794), .A2(n808), .ZN(n806) );
  OR2_X1 U792 ( .A1(n796), .A2(n797), .ZN(n808) );
  OR2_X1 U793 ( .A1(n741), .A2(n606), .ZN(n797) );
  OR2_X1 U794 ( .A1(n809), .A2(n810), .ZN(n796) );
  AND2_X1 U795 ( .A1(n793), .A2(n792), .ZN(n810) );
  AND2_X1 U796 ( .A1(n790), .A2(n811), .ZN(n809) );
  OR2_X1 U797 ( .A1(n792), .A2(n793), .ZN(n811) );
  OR2_X1 U798 ( .A1(n741), .A2(n595), .ZN(n793) );
  OR2_X1 U799 ( .A1(n812), .A2(n813), .ZN(n792) );
  AND2_X1 U800 ( .A1(n789), .A2(n577), .ZN(n813) );
  AND2_X1 U801 ( .A1(n788), .A2(n814), .ZN(n812) );
  OR2_X1 U802 ( .A1(n577), .A2(n789), .ZN(n814) );
  OR2_X1 U803 ( .A1(n815), .A2(n816), .ZN(n789) );
  AND2_X1 U804 ( .A1(n784), .A2(n786), .ZN(n816) );
  AND2_X1 U805 ( .A1(n817), .A2(n785), .ZN(n815) );
  OR2_X1 U806 ( .A1(n818), .A2(n819), .ZN(n785) );
  INV_X1 U807 ( .A(n820), .ZN(n819) );
  AND2_X1 U808 ( .A1(n821), .A2(n822), .ZN(n818) );
  OR2_X1 U809 ( .A1(n607), .A2(n740), .ZN(n822) );
  OR2_X1 U810 ( .A1(n697), .A2(n594), .ZN(n821) );
  OR2_X1 U811 ( .A1(n784), .A2(n786), .ZN(n817) );
  OR2_X1 U812 ( .A1(n782), .A2(n781), .ZN(n786) );
  OR2_X1 U813 ( .A1(n697), .A2(n741), .ZN(n781) );
  OR2_X1 U814 ( .A1(n566), .A2(n741), .ZN(n784) );
  OR2_X1 U815 ( .A1(n701), .A2(n741), .ZN(n577) );
  XNOR2_X1 U816 ( .A(n823), .B(n820), .ZN(n788) );
  XNOR2_X1 U817 ( .A(n824), .B(n825), .ZN(n823) );
  XNOR2_X1 U818 ( .A(n826), .B(n827), .ZN(n790) );
  XNOR2_X1 U819 ( .A(n828), .B(n829), .ZN(n826) );
  XNOR2_X1 U820 ( .A(n830), .B(n831), .ZN(n794) );
  XNOR2_X1 U821 ( .A(n592), .B(n832), .ZN(n830) );
  OR2_X1 U822 ( .A1(n801), .A2(n798), .ZN(n805) );
  XNOR2_X1 U823 ( .A(n833), .B(n834), .ZN(n798) );
  XNOR2_X1 U824 ( .A(n835), .B(n836), .ZN(n833) );
  OR2_X1 U825 ( .A1(n741), .A2(n479), .ZN(n801) );
  INV_X1 U826 ( .A(b_4_), .ZN(n741) );
  XNOR2_X1 U827 ( .A(n837), .B(n657), .ZN(n646) );
  XNOR2_X1 U828 ( .A(n838), .B(n839), .ZN(n657) );
  XOR2_X1 U829 ( .A(n605), .B(n840), .Z(n838) );
  INV_X1 U830 ( .A(n496), .ZN(n605) );
  XNOR2_X1 U831 ( .A(n656), .B(n655), .ZN(n837) );
  OR2_X1 U832 ( .A1(n841), .A2(n842), .ZN(n655) );
  AND2_X1 U833 ( .A1(n836), .A2(n835), .ZN(n842) );
  AND2_X1 U834 ( .A1(n834), .A2(n843), .ZN(n841) );
  OR2_X1 U835 ( .A1(n835), .A2(n836), .ZN(n843) );
  OR2_X1 U836 ( .A1(n844), .A2(n845), .ZN(n836) );
  AND2_X1 U837 ( .A1(n832), .A2(n592), .ZN(n845) );
  AND2_X1 U838 ( .A1(n831), .A2(n846), .ZN(n844) );
  OR2_X1 U839 ( .A1(n592), .A2(n832), .ZN(n846) );
  OR2_X1 U840 ( .A1(n847), .A2(n848), .ZN(n832) );
  AND2_X1 U841 ( .A1(n829), .A2(n828), .ZN(n848) );
  AND2_X1 U842 ( .A1(n827), .A2(n849), .ZN(n847) );
  OR2_X1 U843 ( .A1(n828), .A2(n829), .ZN(n849) );
  OR2_X1 U844 ( .A1(n850), .A2(n851), .ZN(n829) );
  AND2_X1 U845 ( .A1(n820), .A2(n825), .ZN(n851) );
  AND2_X1 U846 ( .A1(n852), .A2(n824), .ZN(n850) );
  OR2_X1 U847 ( .A1(n853), .A2(n854), .ZN(n824) );
  AND2_X1 U848 ( .A1(n855), .A2(n856), .ZN(n853) );
  OR2_X1 U849 ( .A1(n825), .A2(n820), .ZN(n852) );
  OR2_X1 U850 ( .A1(n782), .A2(n856), .ZN(n820) );
  OR2_X1 U851 ( .A1(n740), .A2(n594), .ZN(n782) );
  OR2_X1 U852 ( .A1(n594), .A2(n566), .ZN(n825) );
  OR2_X1 U853 ( .A1(n594), .A2(n701), .ZN(n828) );
  XNOR2_X1 U854 ( .A(n857), .B(n858), .ZN(n827) );
  XOR2_X1 U855 ( .A(n859), .B(n854), .Z(n857) );
  INV_X1 U856 ( .A(n860), .ZN(n854) );
  OR2_X1 U857 ( .A1(n594), .A2(n595), .ZN(n592) );
  XNOR2_X1 U858 ( .A(n861), .B(n862), .ZN(n831) );
  XNOR2_X1 U859 ( .A(n863), .B(n864), .ZN(n861) );
  OR2_X1 U860 ( .A1(n594), .A2(n606), .ZN(n835) );
  XNOR2_X1 U861 ( .A(n865), .B(n866), .ZN(n834) );
  XNOR2_X1 U862 ( .A(n867), .B(n868), .ZN(n865) );
  OR2_X1 U863 ( .A1(n594), .A2(n479), .ZN(n656) );
  INV_X1 U864 ( .A(b_3_), .ZN(n594) );
  AND3_X1 U865 ( .A1(n536), .A2(n534), .A3(n535), .ZN(n537) );
  INV_X1 U866 ( .A(n869), .ZN(n535) );
  OR2_X1 U867 ( .A1(n870), .A2(n871), .ZN(n869) );
  AND2_X1 U868 ( .A1(n639), .A2(n638), .ZN(n871) );
  AND2_X1 U869 ( .A1(n636), .A2(n872), .ZN(n870) );
  OR2_X1 U870 ( .A1(n638), .A2(n639), .ZN(n872) );
  OR2_X1 U871 ( .A1(n607), .A2(n490), .ZN(n639) );
  OR2_X1 U872 ( .A1(n873), .A2(n874), .ZN(n638) );
  AND2_X1 U873 ( .A1(n652), .A2(n651), .ZN(n874) );
  AND2_X1 U874 ( .A1(n649), .A2(n875), .ZN(n873) );
  OR2_X1 U875 ( .A1(n651), .A2(n652), .ZN(n875) );
  OR2_X1 U876 ( .A1(n607), .A2(n479), .ZN(n652) );
  OR2_X1 U877 ( .A1(n876), .A2(n877), .ZN(n651) );
  AND2_X1 U878 ( .A1(n840), .A2(n496), .ZN(n877) );
  AND2_X1 U879 ( .A1(n839), .A2(n878), .ZN(n876) );
  OR2_X1 U880 ( .A1(n496), .A2(n840), .ZN(n878) );
  OR2_X1 U881 ( .A1(n879), .A2(n880), .ZN(n840) );
  AND2_X1 U882 ( .A1(n867), .A2(n868), .ZN(n880) );
  AND2_X1 U883 ( .A1(n866), .A2(n881), .ZN(n879) );
  OR2_X1 U884 ( .A1(n868), .A2(n867), .ZN(n881) );
  OR2_X1 U885 ( .A1(n882), .A2(n883), .ZN(n867) );
  AND2_X1 U886 ( .A1(n864), .A2(n863), .ZN(n883) );
  AND2_X1 U887 ( .A1(n862), .A2(n884), .ZN(n882) );
  OR2_X1 U888 ( .A1(n863), .A2(n864), .ZN(n884) );
  OR2_X1 U889 ( .A1(n607), .A2(n701), .ZN(n864) );
  OR2_X1 U890 ( .A1(n885), .A2(n886), .ZN(n863) );
  AND2_X1 U891 ( .A1(n858), .A2(n860), .ZN(n886) );
  AND2_X1 U892 ( .A1(n887), .A2(n859), .ZN(n885) );
  OR2_X1 U893 ( .A1(n888), .A2(n889), .ZN(n859) );
  AND2_X1 U894 ( .A1(n890), .A2(n891), .ZN(n888) );
  OR2_X1 U895 ( .A1(n740), .A2(n892), .ZN(n890) );
  OR2_X1 U896 ( .A1(n860), .A2(n858), .ZN(n887) );
  OR2_X1 U897 ( .A1(n607), .A2(n566), .ZN(n858) );
  OR2_X1 U898 ( .A1(n856), .A2(n855), .ZN(n860) );
  OR2_X1 U899 ( .A1(n740), .A2(n478), .ZN(n855) );
  OR2_X1 U900 ( .A1(n697), .A2(n607), .ZN(n856) );
  XOR2_X1 U901 ( .A(n893), .B(n889), .Z(n862) );
  INV_X1 U902 ( .A(n894), .ZN(n889) );
  OR2_X1 U903 ( .A1(n895), .A2(n896), .ZN(n893) );
  INV_X1 U904 ( .A(n897), .ZN(n896) );
  AND2_X1 U905 ( .A1(n898), .A2(n899), .ZN(n895) );
  OR2_X1 U906 ( .A1(n697), .A2(n892), .ZN(n898) );
  OR2_X1 U907 ( .A1(n607), .A2(n595), .ZN(n868) );
  XOR2_X1 U908 ( .A(n900), .B(n901), .Z(n866) );
  XOR2_X1 U909 ( .A(n902), .B(n903), .Z(n900) );
  OR2_X1 U910 ( .A1(n607), .A2(n606), .ZN(n496) );
  INV_X1 U911 ( .A(b_2_), .ZN(n607) );
  XOR2_X1 U912 ( .A(n904), .B(n905), .Z(n839) );
  XOR2_X1 U913 ( .A(n906), .B(n907), .Z(n905) );
  XOR2_X1 U914 ( .A(n908), .B(n909), .Z(n649) );
  XOR2_X1 U915 ( .A(n910), .B(n911), .Z(n909) );
  XNOR2_X1 U916 ( .A(n912), .B(n913), .ZN(n636) );
  XNOR2_X1 U917 ( .A(n475), .B(n914), .ZN(n912) );
  XNOR2_X1 U918 ( .A(n915), .B(n621), .ZN(n534) );
  INV_X1 U919 ( .A(n916), .ZN(n621) );
  OR2_X1 U920 ( .A1(n917), .A2(n918), .ZN(n916) );
  AND2_X1 U921 ( .A1(n919), .A2(n920), .ZN(n918) );
  AND2_X1 U922 ( .A1(n921), .A2(n922), .ZN(n917) );
  OR2_X1 U923 ( .A1(n920), .A2(n919), .ZN(n921) );
  OR2_X1 U924 ( .A1(n892), .A2(n490), .ZN(n915) );
  XNOR2_X1 U925 ( .A(n919), .B(n923), .ZN(n536) );
  XOR2_X1 U926 ( .A(n920), .B(n922), .Z(n923) );
  OR2_X1 U927 ( .A1(n478), .A2(n490), .ZN(n922) );
  INV_X1 U928 ( .A(a_0_), .ZN(n490) );
  OR2_X1 U929 ( .A1(n924), .A2(n925), .ZN(n920) );
  AND2_X1 U930 ( .A1(n913), .A2(n914), .ZN(n925) );
  AND2_X1 U931 ( .A1(n926), .A2(n475), .ZN(n924) );
  OR2_X1 U932 ( .A1(n478), .A2(n479), .ZN(n475) );
  OR2_X1 U933 ( .A1(n914), .A2(n913), .ZN(n926) );
  OR2_X1 U934 ( .A1(n606), .A2(n892), .ZN(n913) );
  OR2_X1 U935 ( .A1(n927), .A2(n928), .ZN(n914) );
  AND2_X1 U936 ( .A1(n908), .A2(n910), .ZN(n928) );
  AND2_X1 U937 ( .A1(n929), .A2(n911), .ZN(n927) );
  OR2_X1 U938 ( .A1(n595), .A2(n892), .ZN(n911) );
  OR2_X1 U939 ( .A1(n910), .A2(n908), .ZN(n929) );
  OR2_X1 U940 ( .A1(n478), .A2(n606), .ZN(n908) );
  INV_X1 U941 ( .A(a_2_), .ZN(n606) );
  OR2_X1 U942 ( .A1(n930), .A2(n931), .ZN(n910) );
  AND2_X1 U943 ( .A1(n904), .A2(n906), .ZN(n931) );
  AND2_X1 U944 ( .A1(n932), .A2(n907), .ZN(n930) );
  OR2_X1 U945 ( .A1(n478), .A2(n595), .ZN(n907) );
  INV_X1 U946 ( .A(a_3_), .ZN(n595) );
  OR2_X1 U947 ( .A1(n906), .A2(n904), .ZN(n932) );
  OR2_X1 U948 ( .A1(n701), .A2(n892), .ZN(n904) );
  OR2_X1 U949 ( .A1(n933), .A2(n934), .ZN(n906) );
  AND2_X1 U950 ( .A1(n901), .A2(n903), .ZN(n934) );
  AND2_X1 U951 ( .A1(n902), .A2(n935), .ZN(n933) );
  OR2_X1 U952 ( .A1(n903), .A2(n901), .ZN(n935) );
  OR2_X1 U953 ( .A1(n566), .A2(n892), .ZN(n901) );
  OR2_X1 U954 ( .A1(n478), .A2(n701), .ZN(n903) );
  INV_X1 U955 ( .A(a_4_), .ZN(n701) );
  AND2_X1 U956 ( .A1(n897), .A2(n894), .ZN(n902) );
  OR3_X1 U957 ( .A1(n740), .A2(n892), .A3(n891), .ZN(n894) );
  OR2_X1 U958 ( .A1(n697), .A2(n478), .ZN(n891) );
  INV_X1 U959 ( .A(a_7_), .ZN(n740) );
  OR3_X1 U960 ( .A1(n697), .A2(n892), .A3(n899), .ZN(n897) );
  OR2_X1 U961 ( .A1(n478), .A2(n566), .ZN(n899) );
  INV_X1 U962 ( .A(a_5_), .ZN(n566) );
  INV_X1 U963 ( .A(b_1_), .ZN(n478) );
  INV_X1 U964 ( .A(a_6_), .ZN(n697) );
  OR2_X1 U965 ( .A1(n479), .A2(n892), .ZN(n919) );
  INV_X1 U966 ( .A(b_0_), .ZN(n892) );
  INV_X1 U967 ( .A(a_1_), .ZN(n479) );
endmodule

