module s38584 ( CK, g100, g10122, g10306, g10500, g10527, g113, g11349, g11388, 
        g114, g11418, g11447, g115, g116, g11678, g11770, g120, g12184, g12238, 
        g12300, g12350, g12368, g124, g12422, g12470, g125, g126, g127, g12832, 
        g12833, g12919, g12923, g13039, g13049, g13068, g13085, g13099, g13259, 
        g13272, g134, g135, g13865, g13881, g13895, g13906, g13926, g13966, 
        g14096, g14125, g14147, g14167, g14189, g14201, g14217, g14421, g14451, 
        g14518, g14597, g14635, g14662, g14673, g14694, g14705, g14738, g14749, 
        g14779, g14828, g16603, g16624, g16627, g16656, g16659, g16686, g16693, 
        g16718, g16722, g16744, g16748, g16775, g16874, g16924, g16955, g17291, 
        g17316, g17320, g17400, g17404, g17423, g17519, g17577, g17580, g17604, 
        g17607, g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711, 
        g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787, g17813, 
        g17819, g17845, g17871, g18092, g18094, g18095, g18096, g18097, g18098, 
        g18099, g18100, g18101, g18881, g19334, g19357, g20049, g20557, g20652, 
        g20654, g20763, g20899, g20901, g21176, g21245, g21270, g21292, g21698, 
        g21727, g23002, g23190, g23612, g23652, g23683, g23759, g24151, g24161, 
        g24162, g24163, g24164, g24165, g24166, g24167, g24168, g24169, g24170, 
        g24171, g24172, g24173, g24174, g24175, g24176, g24177, g24178, g24179, 
        g24180, g24181, g24182, g24183, g24184, g24185, g25114, g25167, g25219, 
        g25259, g25582, g25583, g25584, g25585, g25586, g25587, g25588, g25589, 
        g25590, g26801, g26875, g26876, g26877, g27831, g28030, g28041, g28042, 
        g28753, g29210, g29211, g29212, g29213, g29214, g29215, g29216, g29217, 
        g29218, g29219, g29220, g29221, g30327, g30329, g30330, g30331, g30332, 
        g31521, g31656, g31665, g31793, g31860, g31861, g31862, g31863, g32185, 
        g32429, g32454, g32975, g33079, g33435, g33533, g33636, g33659, g33874, 
        g33894, g33935, g33945, g33946, g33947, g33948, g33949, g33950, g33959, 
        g34201, g34221, g34232, g34233, g34234, g34235, g34236, g34237, g34238, 
        g34239, g34240, g34383, g34425, g34435, g34436, g34437, g34597, g34788, 
        g34839, g34913, g34915, g34917, g34919, g34921, g34923, g34925, g34927, 
        g34956, g34972, g35, g36, g44, g5, g53, g54, g56, g57, g64, g6744, 
        g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6752, g6753, g72, 
        g7243, g7245, g7257, g7260, g73, g7540, g7916, g7946, g8132, g8178, 
        g8215, g8235, g8277, g8279, g8283, g8291, g8342, g8344, g8353, g8358, 
        g8398, g84, g8403, g8416, g8475, g8719, g8783, g8784, g8785, g8786, 
        g8787, g8788, g8789, g8839, g8870, g8915, g8916, g8917, g8918, g8919, 
        g8920, g90, g9019, g9048, g91, g92, g9251, g9497, g9553, g9555, g9615, 
        g9617, g9680, g9682, g9741, g9743, g9817, g99, test_se, test_si1, 
        test_so1, test_si2, test_so2, test_si3, test_so3, test_si4, test_so4, 
        test_si5, test_so5, test_si6, test_so6, test_si7, test_so7, test_si8, 
        test_so8, test_si9, test_so9, test_si10, test_so10, test_si11, 
        test_so11, test_si12, test_so12, test_si13, test_so13, test_si14, 
        test_so14, test_si15, test_so15, test_si16, test_so16, test_si17, 
        test_so17, test_si18, test_so18, test_si19, test_so19, test_si20, 
        test_so20, test_si21, test_so21, test_si22, test_so22, test_si23, 
        test_so23, test_si24, test_so24, test_si25, test_so25, test_si26, 
        test_so26, test_si27, test_so27, test_si28, test_so28, test_si29, 
        test_so29, test_si30, test_so30, test_si31, test_so31, test_si32, 
        test_so32, test_si33, test_so33, test_si34, test_so34, test_si35, 
        test_so35, test_si36, test_so36, test_si37, test_so37, test_si38, 
        test_so38, test_si39, test_so39, test_si40, test_so40, test_si41, 
        test_so41, test_si42, test_so42, test_si43, test_so43, test_si44, 
        test_so44, test_si45, test_so45, test_si46, test_so46, test_si47, 
        test_so47, test_si48, test_so48, test_si49, test_so49, test_si50, 
        test_so50, test_si51, test_so51, test_si52, test_so52, test_si53, 
        test_so53, test_si54, test_so54, test_si55, test_so55, test_si56, 
        test_so56, test_si57, test_so57, test_si58, test_so58, test_si59, 
        test_so59, test_si60, test_so60, test_si61, test_so61, test_si62, 
        test_so62, test_si63, test_so63, test_si64, test_so64, test_si65, 
        test_so65, test_si66, test_so66, test_si67, test_so67, test_si68, 
        test_so68, test_si69, test_so69, test_si70, test_so70, test_si71, 
        test_so71, test_si72, test_so72, test_si73, test_so73, test_si74, 
        test_so74, test_si75, test_so75, test_si76, test_so76, test_si77, 
        test_so77, test_si78, test_so78, test_si79, test_so79, test_si80, 
        test_so80, test_si81, test_so81, test_si82, test_so82, test_si83, 
        test_so83, test_si84, test_so84, test_si85, test_so85, test_si86, 
        test_so86, test_si87, test_so87, test_si88, test_so88, test_si89, 
        test_so89, test_si90, test_so90, test_si91, test_so91, test_si92, 
        test_so92, test_si93, test_so93, test_si94, test_so94, test_si95, 
        test_so95, test_si96, test_so96, test_si97, test_so97, test_si98, 
        test_so98, test_si99, test_so99, test_si100, test_so100 );
  input CK, g100, g113, g114, g115, g116, g120, g124, g125, g126, g127, g134,
         g135, g35, g36, g44, g5, g53, g54, g56, g57, g64, g6744, g6745, g6746,
         g6747, g6748, g6749, g6750, g6751, g6752, g6753, g72, g73, g84, g90,
         g91, g92, g99, test_se, test_si1, test_si2, test_si3, test_si4,
         test_si5, test_si6, test_si7, test_si8, test_si9, test_si10,
         test_si11, test_si12, test_si13, test_si14, test_si15, test_si16,
         test_si17, test_si18, test_si19, test_si20, test_si21, test_si22,
         test_si23, test_si24, test_si25, test_si26, test_si27, test_si28,
         test_si29, test_si30, test_si31, test_si32, test_si33, test_si34,
         test_si35, test_si36, test_si37, test_si38, test_si39, test_si40,
         test_si41, test_si42, test_si43, test_si44, test_si45, test_si46,
         test_si47, test_si48, test_si49, test_si50, test_si51, test_si52,
         test_si53, test_si54, test_si55, test_si56, test_si57, test_si58,
         test_si59, test_si60, test_si61, test_si62, test_si63, test_si64,
         test_si65, test_si66, test_si67, test_si68, test_si69, test_si70,
         test_si71, test_si72, test_si73, test_si74, test_si75, test_si76,
         test_si77, test_si78, test_si79, test_si80, test_si81, test_si82,
         test_si83, test_si84, test_si85, test_si86, test_si87, test_si88,
         test_si89, test_si90, test_si91, test_si92, test_si93, test_si94,
         test_si95, test_si96, test_si97, test_si98, test_si99, test_si100;
  output g10122, g10306, g10500, g10527, g11349, g11388, g11418, g11447,
         g11678, g11770, g12184, g12238, g12300, g12350, g12368, g12422,
         g12470, g12832, g12833, g12919, g12923, g13039, g13049, g13068,
         g13085, g13099, g13259, g13272, g13865, g13881, g13895, g13906,
         g13926, g13966, g14096, g14125, g14147, g14167, g14189, g14201,
         g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673,
         g14694, g14705, g14738, g14749, g14779, g14828, g16603, g16624,
         g16627, g16656, g16659, g16686, g16693, g16718, g16722, g16744,
         g16748, g16775, g16874, g16924, g16955, g17291, g17316, g17320,
         g17400, g17404, g17423, g17519, g17577, g17580, g17604, g17607,
         g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711,
         g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787,
         g17813, g17819, g17845, g17871, g18092, g18094, g18095, g18096,
         g18097, g18098, g18099, g18100, g18101, g18881, g19334, g19357,
         g20049, g20557, g20652, g20654, g20763, g20899, g20901, g21176,
         g21245, g21270, g21292, g21698, g21727, g23002, g23190, g23612,
         g23652, g23683, g23759, g24151, g24161, g24162, g24163, g24164,
         g24165, g24166, g24167, g24168, g24169, g24170, g24171, g24172,
         g24173, g24174, g24175, g24176, g24177, g24178, g24179, g24180,
         g24181, g24182, g24183, g24184, g24185, g25114, g25167, g25219,
         g25259, g25582, g25583, g25584, g25585, g25586, g25587, g25588,
         g25589, g25590, g26801, g26875, g26876, g26877, g27831, g28030,
         g28041, g28042, g28753, g29210, g29211, g29212, g29213, g29214,
         g29215, g29216, g29217, g29218, g29219, g29220, g29221, g30327,
         g30329, g30330, g30331, g30332, g31521, g31656, g31665, g31793,
         g31860, g31861, g31862, g31863, g32185, g32429, g32454, g32975,
         g33079, g33435, g33533, g33636, g33659, g33874, g33894, g33935,
         g33945, g33946, g33947, g33948, g33949, g33950, g33959, g34201,
         g34221, g34232, g34233, g34234, g34235, g34236, g34237, g34238,
         g34239, g34240, g34383, g34425, g34435, g34436, g34437, g34597,
         g34788, g34839, g34913, g34915, g34917, g34919, g34921, g34923,
         g34925, g34927, g34956, g34972, g7243, g7245, g7257, g7260, g7540,
         g7916, g7946, g8132, g8178, g8215, g8235, g8277, g8279, g8283, g8291,
         g8342, g8344, g8353, g8358, g8398, g8403, g8416, g8475, g8719, g8783,
         g8784, g8785, g8786, g8787, g8788, g8789, g8839, g8870, g8915, g8916,
         g8917, g8918, g8919, g8920, g9019, g9048, g9251, g9497, g9553, g9555,
         g9615, g9617, g9680, g9682, g9741, g9743, g9817, test_so1, test_so2,
         test_so3, test_so4, test_so5, test_so6, test_so7, test_so8, test_so9,
         test_so10, test_so11, test_so12, test_so13, test_so14, test_so15,
         test_so16, test_so17, test_so18, test_so19, test_so20, test_so21,
         test_so22, test_so23, test_so24, test_so25, test_so26, test_so27,
         test_so28, test_so29, test_so30, test_so31, test_so32, test_so33,
         test_so34, test_so35, test_so36, test_so37, test_so38, test_so39,
         test_so40, test_so41, test_so42, test_so43, test_so44, test_so45,
         test_so46, test_so47, test_so48, test_so49, test_so50, test_so51,
         test_so52, test_so53, test_so54, test_so55, test_so56, test_so57,
         test_so58, test_so59, test_so60, test_so61, test_so62, test_so63,
         test_so64, test_so65, test_so66, test_so67, test_so68, test_so69,
         test_so70, test_so71, test_so72, test_so73, test_so74, test_so75,
         test_so76, test_so77, test_so78, test_so79, test_so80, test_so81,
         test_so82, test_so83, test_so84, test_so85, test_so86, test_so87,
         test_so88, test_so89, test_so90, test_so91, test_so92, test_so93,
         test_so94, test_so95, test_so96, test_so97, test_so98, test_so99,
         test_so100;
  wire   g100, g113, g114, g115, g116, g120, g124, g125, g126, g127, g134,
         g135, g18881, g23612, g23652, g73, g29211, g29212, g29213, g29214,
         g29215, g29216, g29217, g29219, g29220, g29221, g30327, g30331,
         g30332, g31656, g31665, g33533, g34435, g34788, g34839, g36, g44, g53,
         g54, g56, g57, g64, g6744, g6745, g6746, g6747, g6748, g6749, g6750,
         g6751, g6753, g84, g90, g91, g92, g99, test_so10, test_so26,
         test_so35, test_so39, test_so42, test_so44, test_so46, test_so80,
         test_so86, test_so92, test_so100, g34783, n2730, n4836, n4896, n4895,
         n4837, n4921, n4920, n2787, n4411, n5045, g559, n4959, g33046, g5057,
         n5615, g34441, g2771, n5544, g33982, g1882, g34007, g2299, g24276,
         g4040, n5530, g30381, g2547, n5782, g30405, g3243, g25604, g452,
         g30416, g3542, g30466, g5232, g25736, g5813, g34617, g33974, g1744,
         n5795, g30505, g5909, g33554, g1802, n5536, g30432, g3554, g33064,
         g6219, n5385, g34881, g807, n5479, g6031, g24216, g847, n5709, g24232,
         n9367, DFF_24_n1, g34733, g4172, g34882, g4372, g33026, g3512, g31867,
         n5471, g25668, g3490, n5454, g24344, n5432, g4235, g33966, g1600,
         n5811, g33550, g1714, n5460, g30393, g3155, n5366, g29248, g2236,
         g4571, g4555, g24274, g3698, g33973, g1736, n5817, g30360, g1968,
         n5664, g34460, g30494, g5607, g30384, g2657, n5316, g24340, n5439,
         g29223, g490, n5708, g26881, g311, n5317, g34252, g772, n5334, g30489,
         g5587, g29301, g6177, n5874, g6377, g33022, g3167, n5652, g30496,
         g5615, g33043, g4567, g29263, g30533, g6287, g24256, n5302, g34015,
         g2563, n5816, g34031, g4776, n5707, g34452, g4593, n5303, g34646,
         g6199, n5644, g34001, g2295, n5815, g25633, g1384, g24259, g1339,
         n5381, g33049, g5180, n5384, g34609, g2844, g31869, g1024, g30490,
         g30427, g3598, g21894, g4264, n5823, g33965, g767, n5333, g34645,
         g5853, n5499, n5580, g33571, g2089, g34267, g4933, n5878, g26971,
         g4521, n5752, g34644, g5507, n5643, g30534, g6291, g33535, g294,
         n5680, g30498, g25728, n5722, g25743, g25684, g3813, g25613, g562,
         g34438, g608, n5475, g24244, g1205, n5547, g30439, g3909, g30541,
         g6259, g30519, g5905, g25621, g921, g34807, g2955, g25599, g203,
         g24235, g34036, g4878, n5283, g30476, g5204, g30429, g3606, g32997,
         g1926, n5510, g33063, g6215, n5651, g30424, g3586, g32977, g291,
         n5679, g34026, g4674, n5440, g30420, g3570, g33560, g29226, g676,
         n5751, g25619, g843, g34455, g4332, n5540, g30457, g4153, g33625,
         g6336, n5592, g34790, g622, n5672, g30414, g3506, n5576, g26966,
         g4558, g25656, g3111, g30390, g25688, g34727, g939, n5415, g25594,
         g278, n5627, g26963, g4492, g34034, g4864, n5318, g33541, g1036,
         g28093, g24236, g1178, g30404, g3239, g28051, g718, g29303, g6195,
         g26917, g1135, n5328, g33624, g6395, n5396, g24337, g34911, g554,
         g33963, g496, g34627, g3853, n5641, g29282, g5134, n5807, g25676,
         n5721, g33013, g2485, n5509, g32981, g925, n5725, g34976, n9357,
         g30483, g5555, g32994, g1798, n5833, g28070, g34806, g2941, g30453,
         g3905, g33539, g763, n5332, g30526, g6255, g26951, g4375, g34035,
         g4871, n5443, g34636, g4722, n5345, g32978, g590, n5472, g30348,
         g1632, n5836, g24336, n5438, g3100, g24250, g29236, g1437, n5696,
         g29298, g6154, n5747, g1579, g30499, g5567, g33976, g1752, n5797,
         g32996, g1917, g30335, g744, n5470, g34637, g4737, n5867, g25694,
         g30528, g6267, g24251, g1442, g30521, g26960, g4477, n5849, g24239,
         g34259, g4643, n5382, g30474, g5264, n5703, g33016, g2610, g34643,
         g5160, n5498, g30510, g5933, g29239, g1454, n5866, g26897, g753,
         g34729, g1296, g34625, g3151, n5495, g34800, g24353, g6727, n5531,
         g33029, g3530, n5569, g33615, g4104, g24253, g1532, g24281, g33997,
         n9352, g34971, n9351, g34263, g4754, n5877, g24237, g1189, n5642,
         g33584, g2287, n5353, g24280, g4273, n5764, g26920, g1389, g33548,
         g29296, g5835, n5663, g30338, g1171, n5363, g21895, g4269, n5763,
         g33588, g2399, n5762, g34041, g4983, n5367, g30495, g5611, g29279,
         g4572, g25655, g3143, n5882, g34795, g2898, g24269, g3343, g30403,
         g3235, g33042, g30419, g3566, g34023, n9348, DFF_228_n1, g28090,
         g4961, n5770, g34642, g4927, n5879, g30370, g2259, n5419, g34448,
         g2819, n5609, g26946, g5802, g34610, g2852, g24209, g417, n5358,
         g28047, g681, g24206, g437, g26891, g30504, g5901, g34798, g2886,
         g25669, g3494, n5889, g30480, g5511, n5575, g33027, g3518, n5645,
         g33972, g1604, g25697, g5092, g28099, g4831, g26947, g4382, n5714,
         g24350, g6386, g24210, g479, g30455, g3965, g28084, g33993, g2008,
         g736, g30444, g3933, g33537, g222, g25650, g3050, g25625, g1052,
         g30366, g2122, n5784, g33593, g2465, n5523, g30502, g5889, g33036,
         g4495, g25595, g34462, g33024, g3179, n5390, g33552, g1728, n5352,
         g34014, g2433, g29273, g3835, n5662, g25748, g6187, n5453, g34638,
         g4917, n5408, g30341, g1070, g26899, g822, n5422, g30336, g914, n5560,
         g5339, g26940, g4164, g25622, g34447, g2807, n5379, g33613, g4054,
         n5395, g25749, g6191, n5888, g25704, g5077, n5455, g33053, g5523,
         n5647, g3680, g30555, g6637, g25601, g174, n5402, g33971, g1682,
         g26892, g355, g1087, g26915, g1105, n5478, g33008, g30538, g6307,
         g3802, g25750, g6159, g30369, g2255, n5414, g34446, g2815, n5404,
         g29230, g911, n5559, g43, g33975, g1748, g30497, g5551, g30418, g3558,
         g25721, g5499, n5885, g34622, g30438, g3901, g34266, g4888, n5863,
         g30540, g6251, g32986, g1373, g25648, n5723, g33960, g157, n5678,
         g34442, g2783, n5403, g4281, g30421, g3574, g33573, g2112, n5848,
         g34730, g1283, n5635, g24205, g10122_Tj, g4297, n5698, g32979, g758,
         n5331, g4639, n5727, g25763, g6537, n5884, g30481, g5543, g30517,
         g5961, g30539, g6243, g34880, n9340, g24242, n5654, g30436, g29265,
         g3476, n5786, g32990, g1664, n5407, g24245, g1246, n5756, g30553,
         g6629, g26907, g246, n6008, g24278, g4049, g26955, g24282, g2932,
         g29276, g4575, g31894, g4098, n5350, g33037, g4498, g26894, g528,
         n5327, g34977, n5477, g25654, g3139, n5447, g33962, g34451, g4584,
         n5539, g34250, g142, n5724, g29295, g5831, g26905, g239, g25629,
         g1216, n5442, g34792, g2848, g25703, g5022, g32983, g1030, g30402,
         g3231, g25757, g1430, n9336, g33999, g2241, g24262, g1564, g25729,
         g6148, g30558, g6649, g34781, g110, g26901, g225, n5597, g26961,
         g33039, g4504, g33059, g5873, n5388, g31899, g5037, n5611, g33007,
         g2319, n5375, g25720, g5495, n5446, g21891, g30462, g5208, g30487,
         g5579, g33058, g5869, n5649, g24261, g1589, n5755, g25730, g5752,
         g30531, g6279, g30506, g34804, g2975, n5750, g25747, g6167, n5430,
         n5701, g33601, g2599, n5524, g26922, g1448, n5343, g29250, g2370,
         g30459, g5164, n5570, g1333, n5616, g33534, g153, n5677, g30543,
         g6549, n5571, g29275, g4087, n5480, g34030, g34980, g2984, n5842,
         g30451, g3961, g25627, g962, n5630, g34657, g101, g30552, g6625,
         g34979, n9332, g30337, g1018, g24254, g24277, g4045, g29237, g1467,
         n5693, g30378, g2461, n5840, g33019, n5300, g33623, g5990, n5589,
         g29235, g1256, n5558, g31902, g5029, n5601, g29306, g6519, n5806,
         g25689, g4169, n5729, g33978, g1816, g26970, g4369, g29278, g4578,
         g34253, g4459, n5765, g29272, g3831, n5872, g33595, g2514, g33610,
         g3288, n5400, g33589, g34605, g2145, n5307, g30350, g1700, n5417,
         g25611, g513, n5548, g2841, n5963, g33619, g5297, n5588, g34022,
         g2763, g34033, g4793, n5368, g34726, g952, g31870, g1263, n5674,
         g33985, g1950, g29283, g5138, n5871, g34003, g2307, g25677, g34463,
         g4664, g33006, g2223, n5406, g29292, g5808, n5749, g30557, g6645,
         g33989, g2016, g33033, g3873, n5387, n5699, g34005, g2315, n5802,
         g26932, g2811, g30516, g5957, g33575, g2047, n5831, g33032, g30486,
         g5575, g34974, n9327, g25678, g3752, g30440, g3917, DFF_480_n1, g1585,
         n5757, g26949, g4388, g30530, g6275, g30542, g6311, g25624, g1041,
         g30383, g33597, g2537, n5411, g34598, g26957, g4430, g26967, n9325,
         g28102, g4826, g30524, g6239, g26903, g232, g30475, g5268, g34647,
         g6545, n5497, g30377, n9324, g33553, g1772, n5504, g31903, g5052,
         n5607, g25715, g33984, g1890, n5799, g33602, g2629, n5521, g28045,
         g572, n5337, g34603, g2130, n5487, g33035, g4108, g4308, g24208, g475,
         g990, n5622, g31, n5469, g34970, n9322, g24213, g33614, g3990, n5594,
         g33060, g30362, g1992, n5890, g33023, g3171, n5603, g26898, g812,
         n5733, g25618, g832, g30518, g5897, g4570, n5702, g26959, g4455,
         g34801, g2902, g26884, g333, g25600, g168, g26933, g28066, g3684,
         n5881, g33612, g3639, n5591, n5579, g24268, g3338, n5527, g25716,
         g5406, g26906, g269, g24203, g401, g24346, g6040, g24207, g441,
         g25701, n5690, g29269, g3808, n5745, g9, n5468, g34255, g30450, g3957,
         g30456, g4093, n5340, g32991, g1760, n5602, g24348, n5437, g34249,
         g160, n5843, g30371, g2279, n5778, g29268, g3498, g29224, g586, n5336,
         g33017, g2619, n5508, g30339, g1183, n5599, g33967, g1608, n5792,
         g33559, g1779, n5830, g29255, g2652, g30368, g2193, n5839, g30375,
         g2393, n5421, g28052, g661, g28089, g4950, n5772, g33055, g5535,
         n5566, g30392, g2834, g30343, g1361, g30523, g6235, g24233, g1146,
         n5851, g33018, g32976, g150, n5676, g30349, g1696, n5628, g33067,
         g6555, g26900, g33034, g3881, n5564, g30551, g6621, g25667, g3470,
         n5424, g30452, g3897, g34719, g518, g538, n5491, g33607, g2606, n5311,
         g26923, g1472, n5290, g24211, g33050, g5188, n5567, g24341, g5689,
         n5529, g24201, g405, g30463, g5216, g6494, g34464, g4669, g24243,
         g996, g24335, g4531, g34611, g2860, g34262, g4743, n5876, g30546,
         g6593, g25591, g4411, g30347, g1413, g30556, g6641, g6, g33562, g1936,
         n5534, g55, g25610, g504, n5519, g33015, g2587, n5372, g31896, g4480,
         g34004, n9314, g30428, g30485, g5571, g30422, g3578, g25714, g29294,
         g5827, n5809, g30423, g3582, g30529, g6271, g34028, g4688, n5656,
         g33587, g2380, g30460, g5196, g30401, g3227, g33990, n9312, g29309,
         g6541, g30411, g3203, g33546, g1668, n5598, g28085, g4760, n5775,
         g26904, g262, g33556, g1840, n5451, g25722, g5467, g25605, g460,
         g33062, g6209, g26893, n5704, g28050, g655, g34626, g33583, g2204,
         n5620, g30472, g5256, g34454, g4608, n5274, g34850, g794, n5291,
         n5583, g4423, g24272, g3689, n5532, g5685, g24214, g703, n5821,
         g26909, g862, n5682, g30406, g3247, g33569, g2040, n5505, g34628,
         g4146, n5981, g34458, g4633, n5844, g24240, n5304, g34634, g4732,
         n5296, g25700, n5689, g29293, g5817, g33009, g2351, n5511, g33603,
         g2648, g24355, g6736, g34268, g4944, n5875, g25691, g4072, g26890,
         g29264, g3466, g28072, g4116, g31900, g5041, n5605, g26956, g4434,
         g29271, g3827, n5808, g29304, g6500, n5748, g29261, g3133, n5661,
         g28063, g3333, g979, n5320, g34027, g4681, g33961, g298, n5675,
         g33604, g32995, g1894, n5374, g34624, g2988, g30415, g3538, g33536,
         g301, g26888, n9306, g28055, g827, n5728, g24238, g33600, g2555,
         n5351, g28105, g5011, g34721, g199, g29307, g6523, n5870, g30345,
         g34453, g4601, n5365, g32980, g854, g29238, g1484, n5865, g34639,
         g4922, n5346, g25695, g5080, n5893, g33057, g5863, g26969, g4581,
         n5670, g29253, g2518, g34021, g2567, g26895, g568, n5335, g30413,
         g3263, g30549, g6613, g24347, g25758, g6444, g34808, g2965, g30501,
         g5857, n5573, g33969, n9303, g34440, g890, n5305, g30433, g3562,
         g21900, g26921, g1404, g29270, g3817, n9302, n6010, g33038, g4501,
         g31865, g26926, g2724, n5301, g28083, g4704, n5771, g34797, g22,
         g2878, g30478, g5220, g34724, g617, n5339, g24212, g26883, g316,
         g32985, g1277, g25761, g6513, n5426, g26886, g336, n5824, g34796,
         g2882, g32982, g33561, g1906, n5503, g26880, g305, n5282, g34975, g8,
         g26931, g2799, g34641, g4912, n5297, g34629, g4157, n5983, g33598,
         g2541, n5461, g33576, g2153, n5356, g34720, g550, g26902, g255,
         g29244, g30468, g5240, g26924, g1478, n5289, g33031, g3863, g29245,
         g1959, g29266, g3480, n5868, g30559, g6653, g34794, g2864, n5489,
         g28087, g4894, n5774, g30435, g3857, n5572, g25609, g28057, g1002,
         g34439, g776, n5330, g28, n5324, g1236, g34260, g4646, n5712, g33012,
         g2476, g32989, g1657, n5525, g34006, g2375, g63, g358, g26910, g896,
         n5431, g28043, g33021, g3161, g29251, g2384, n5700, g34456, g4616,
         n5608, g26968, g4561, g33991, g2024, n5801, g3451, g26930, g2795,
         g34599, g613, n5474, g28082, g4527, g33557, g1844, n5847, g30511,
         g5937, g33045, g30379, g2523, n5281, g24267, n5436, g34020, g2643,
         g24249, g1489, n5850, g25592, g30382, n9295, g29285, g5156, n5526,
         n9294, g25662, n5717, g21896, g33563, g1955, g33622, g33582, g2273,
         n5458, n5584, g28086, g4771, n5769, g25744, g6098, g29262, g3147,
         g24270, g3347, g33581, g2269, n5410, g191, g24266, g2712, g34849,
         g626, n5288, g33618, g2729, g5357, n5393, g34038, g34032, g4709,
         n5518, g34803, g2927, g34459, g4340, n5653, g30509, g5929, g34640,
         g4907, n5295, g28069, g4035, g21899, g2946, g31868, g918, n5673,
         g26938, g4082, g25756, n5719, g30363, g30334, g577, n5294, g33970,
         g1620, n5791, g30391, g2831, g25615, g667, g33540, g930, n5731,
         g30445, g3937, g25617, g817, n5822, g24247, g1249, g24215, g837,
         n5562, g33964, g599, n5550, g25719, g5475, n5425, g29228, g30514,
         g5949, g33627, g6682, n5590, g24231, g904, g34615, g2873, n5488,
         g30356, g1854, n5785, g25696, g5084, n5681, g30493, g5603, n5726,
         g33594, g2495, n5522, g34009, g2437, n5789, g30365, g2102, n5666,
         g33004, g2208, g34018, g25685, g4064, n5416, g34040, g4899, n5517,
         g25639, g2719, n5465, g34029, g4785, n5361, g30488, g5583, g34600,
         g781, n5551, g29300, g6173, n5810, g34802, g2917, g25614, g686,
         g28058, g1252, n5554, g29225, g671, g33580, g30532, g6283, n5586,
         DFF_909_n1, g33054, g5527, n5389, g26962, g4489, g33564, g1974, n5450,
         g32984, g1270, n5716, g34039, g4966, n5706, g33065, g6227, n5568,
         g30443, g3929, g29291, g5503, g24279, g30508, g5925, g29232, g1124,
         n5692, g34269, g4955, n5614, g30464, g5224, g33988, g2012, n5790,
         g30522, g6203, n5574, g25708, g5120, g30374, g2389, n5631, g26953,
         g4438, g34008, g2429, n5814, g34444, g2787, n5610, g34731, g33606,
         g2675, n5457, g24334, n5541, g34265, g4836, n5713, g30340, g1199,
         g24257, n5401, g30482, g5547, g34604, g2138, n5275, g33591, g2338,
         n5310, g30525, g6247, g26929, g2791, g30448, g34602, g1291, n2549,
         g30513, g5945, g30469, g5244, g33608, g2759, g33626, g6741, n5398,
         g34725, g785, n5293, g30342, g1259, n5553, g29267, g3484, n5668,
         g25593, g209, g30548, g6609, g33052, g5517, g34012, g2449, n5798,
         g34017, n9281, g24263, g2715, n5299, g26912, g936, n5557, g30364,
         g2098, n5280, g34254, g4462, n5671, g34251, g604, n5473, g30560,
         g6589, g33983, n9280, g24204, g429, g33980, g1870, n5813, g34631,
         g29243, g1825, g25623, g1008, n5321, g26950, g4392, n5710, g30431,
         g3546, g30467, g5236, g30353, g1768, n5834, g34467, g4854, g30442,
         g3925, g29305, g6509, g25616, g732, n5732, g29252, g2504, g4519,
         g4520, g33003, g2185, n5376, g34613, g37, g4031, g33570, g2070, n5535,
         g34734, g4176, n5494, g24275, n5435, g4405, g872, g29302, g6181,
         n5667, g24349, g34264, g4765, n5613, g30484, g5563, g25634, g1395,
         g33567, g1913, n5828, g33585, g2331, n5513, g30527, g6263, g34978,
         n9276, g30447, g3945, g347, n5860, g34256, g4473, g25630, g1266,
         g29290, g5489, n5660, g29227, g31872, g2748, n5516, g29287, g5471,
         g31897, g4540, g6723, g30562, g6605, g34011, n9274, g33996, g2173,
         g21898, g33014, g2491, n5405, g34465, g4849, g33995, g2169, n5788,
         g30372, n9273, g30545, g30389, g33590, g2407, n5459, g34616, g2868,
         g26927, g2767, g32992, g1783, n5596, g25631, g1312, n5466, g30477,
         g5212, g34632, g4245, g28046, g645, g4291, g26896, g25602, g26916,
         g1129, n5329, g33578, g2227, n5538, g33579, g2246, g30354, g1830,
         n5413, g30425, g3590, g24200, g392, g33544, g1592, n5362, g25764,
         g6505, g24246, g1221, g30507, g5921, g26889, g30333, g218, g32998,
         g1932, n5829, g32987, g1624, n5370, g25702, g5062, g29286, g5462,
         n5744, g34606, g2689, n5347, g33070, g6573, n5563, g29240, g1677,
         g32999, g2028, n5371, g33605, g2671, n5278, g24255, g26945, g33558,
         g1848, n5464, g25699, n5669, g29289, g5485, n5869, g30388, g2741,
         n5349, n5482, g29254, g2638, g28074, g4122, g34450, g4322, n5506,
         g30512, g5941, g33572, g2108, n5452, g25, g33551, g33538, g595, n5476,
         g33005, g2217, n5512, g24248, n9267, DFF_1092_n1, g33002, g2066,
         n5832, g24234, g1152, n5618, g30471, g5252, g34000, g2165, g34016,
         g2571, n5787, g33048, g5176, n5650, n5581, g25628, g26934, g2827,
         g34468, g4859, g24202, g424, g33542, g1274, n5730, n9265, g34445,
         g2803, n5545, g33555, g1821, g34013, g2509, g28091, g5073, g26919,
         n5556, g30554, g6633, g29281, g5124, g30537, g6303, g28092, g5069,
         g34732, g2994, n5634, g28049, g650, g33545, g1636, n5549, g30441,
         g3921, g29247, g24354, g6732, g25636, g1306, n5796, g26914, g1061,
         g25670, g3462, g33998, g2181, n5803, g25626, g956, n5341, g33977,
         g1756, n5804, g29297, g5849, g28071, g4112, g30387, n9262, g33577,
         g2197, n5514, g33592, g26913, g1046, g28044, g482, n5820, g26948,
         g4401, g30344, g1514, n5364, g26885, g329, n5766, g33069, g6565,
         n5386, g34621, g2950, g28059, g1345, g25762, g6533, n5445, g34633,
         g4727, n5312, g24352, g26925, g1536, g30446, g3941, g25597, g370,
         g24342, g5694, g30357, g1858, n5892, g26908, g446, g30399, g3219,
         g29242, g1811, g30547, g6601, g34010, g2441, g33986, g1874, g34257,
         g30544, g6581, g30561, g6597, g5008, n5637, g30430, g3610, g34799,
         g2890, g33565, g1978, n5845, g33968, g1612, g34843, g112, g34793,
         g2856, g33566, g1982, n5462, g30465, g28073, g4119, g24351, g6390,
         g30346, g1542, g21893, g4258, g4818, g31904, g5033, g34635, g4717,
         n5344, g25637, g1554, n5768, g29274, g3849, g30396, g3199, g25735,
         g34037, g4975, n5360, g34791, g790, n5292, g30520, g5913, g30358,
         g1902, n5837, g29299, g6163, g25690, g4125, g28096, g4821, g28088,
         g4939, g24241, n5392, g30397, g3207, g4483, g30409, g29284, g5142,
         n5658, g30470, g5248, g30367, g2126, n5891, g24273, g3694, g29288,
         g5481, n5805, g30359, g1964, n5315, g25698, g5097, n5753, g30398,
         g3215, n9255, g26952, g4427, g26928, g2779, n5694, g26954, g30351,
         g1720, n5780, g31871, g1367, g5112, g19, g26939, g4145, g33994, g2161,
         n5812, g25596, g376, n5633, g33586, g2361, n5537, g21901, DFF_1234_n1,
         g31866, g582, n5552, g33000, g2051, g26918, g1193, g30373, g2327,
         n5841, g28056, g907, n5555, g34601, g947, n5286, g30355, g1834, n5665,
         g30426, g3594, g34805, g2999, g34002, g2303, n5794, g28053, g29229,
         g723, n5826, g33620, g5703, n5397, g34722, g546, n5492, g33599, g2472,
         n5619, g30515, g5953, g25649, g33979, g1740, g30417, g3550, g25683,
         g3845, n5886, g33574, g2116, n5463, n5582, g30410, g30454, g3913,
         g34024, g33547, g1687, g30386, g2681, n5777, g33596, g2533, n5761,
         g26887, g324, n5827, g34607, g2697, n5308, g31895, g4417, g33068,
         g6561, n5646, g29233, g1141, n5691, g24258, n5655, g30376, g33549,
         g1710, n5412, g29308, g6527, n5659, g30408, g3255, g29241, g1691,
         g34620, g2936, g33621, g5644, n5593, g25707, g5152, n5883, g24339,
         g5352, g34443, g2775, n5378, g34619, g2922, g29234, g30503, g5893,
         g30550, g6617, g33001, g2060, n5507, g33040, g4512, g30492, g5599,
         g25664, g3401, g26944, g4366, g34614, g29260, g3129, g33047, g5170,
         g24298, g25733, g5821, n5429, g30536, g6299, g29246, g2079, g34261,
         g4698, n5862, g33611, g3703, n5399, g25638, g1559, n5441, g34728,
         n9247, g29222, g411, n5629, g25742, n5718, g30449, g3953, g34608,
         g2704, n5377, g24345, g6035, n5528, n9245, g25635, g1300, g25686,
         g4057, n5711, g30461, g5200, g34466, g4843, g31901, g5046, n5578,
         g29249, g2250, g26882, n5456, g33041, g33011, g2453, n5373, g25734,
         g5841, n5449, n5705, g34618, g2912, g33010, g2357, n5276, g31864,
         g164, n5561, g34630, g4253, n5484, g31898, g5016, n5369, g25653,
         g3119, n5423, g25632, g1351, n5322, g32988, g33616, g29280, g5115,
         n5743, g33609, g3352, n5604, g30563, g6657, g33044, g4552, g30437,
         g3893, g30412, g3211, g30491, g5595, g30434, g3614, g34612, g29259,
         g3125, n5781, g25681, g3821, n5428, g25687, g4141, n5612, g33617,
         g30479, g5272, g29256, g2735, n5600, g28054, g728, g30535, g6295,
         g30385, g2661, n5418, g30361, g1988, n5783, g25705, g24260, g1548,
         n5546, g29257, g3106, n5742, g34461, g4659, g34258, g4358, n5348,
         g32993, g1792, n5359, g33992, g2084, g30394, g3187, g34449, g4311,
         n5323, g34019, g2583, n5800, g18597, n9240, DFF_1381_n1, g29231,
         g1094, n5697, g25682, g21897, g4284, g30395, g3191, g21892, g4239,
         g4180, n5380, g28048, g691, n5520, g34723, g534, n5490, g25598, g385,
         n5632, g33987, g2004, n5818, g30380, g2527, n5420, g5456, g26965,
         n6007, g25706, g30458, g4507, n5846, g24338, g5348, g30400, g3223,
         g34623, g2970, g24343, g5698, g30473, g5260, g24252, g1521, n5577,
         g33028, g3522, n5383, g29258, g3115, g30407, g3251, g26958, g34457,
         g33568, g1996, n5355, g25663, g26964, g4515, g34735, g4300, n5639,
         g30352, n9236, g33543, g1379, g24271, n5433, g33981, g1878, n5793,
         g30500, g5619, g34649, g71, g29277, g25612, n5287, g28060, n2505,
         n2499, n2461, n2396, n2668, n3160, n3141, g72, n5960, n4689, n5961,
         n4708, n3589, n3595, n3570, n3576, n3513, n3519, n3624, n3630, n3551,
         n3557, n3642, n3648, n3532, n3538, n3611, n3607, n3613, n3006, n3765,
         n3505, n3525, n3635, n4888, n3550, n2595, n2527, n3524, n3005, n3623,
         n3549, n3003, n3007, n3569, n3606, n3588, n3165, n3799, n3033, n3622,
         n3587, n3586, n3605, n3604, n3568, n3567, n3548, n3512, n3511, n3531,
         n3530, n3641, n3640, n3131, n3111, n3907, n3773, n3807, n3950, n3841,
         n3983, n3874, n4014, n4537, n4201, n3745, n3684, n3274, n2982, n2706,
         n2649, n2556, n2509, n2487, n2427, n2423, n2421, n4172, n4173, n4190,
         n4191, n4388, n4210, n3479, n3951, n3404, n3774, n3424, n3842, n3414,
         n3808, n3444, n3908, n3489, n3984, n3434, n3875, n3500, n4015, n3446,
         n3914, n3406, n3780, n3481, n3957, n3426, n3848, n3491, n3990, n3416,
         n3814, n3436, n3881, n3502, n4022, n3501, n4027, n3407, n3785, n3482,
         n3962, n3427, n3853, n3437, n3886, n3417, n3819, n3492, n3995, n3447,
         n3919, n3682, n3272, n2980, n2704, n2647, n2554, n2507, n2485, n2425,
         n2419, n3743, n2405, n2760, n2552, n4946, n4198, n2404, n4962, n4948,
         n2726, n2727, n3195, n2774, n3116, n4945, n4525, n3281, n3277, n3276,
         n2989, n2991, n2710, n2707, n3174, n3362, n3676, n2644, n3146, n3115,
         n3833, n3023, n3933, n3729, n4723, n2601, n3664, n3662, n3673, n3671,
         n2607, n3506, n2790, n4490, n4178, n4514, n4196, n3736, n3741, n2598,
         n4814, n4519, n2594, n3084, n2590, n4722, n3125, n3105, n3145, n3164,
         n3910, n3776, n3877, n3810, n3953, n3986, n3844, n3770, n3904, n3804,
         n3947, n3838, n3871, n3980, n4020, n3945, n3836, n3768, n3869, n3978,
         n3802, n3902, n2422, n5121, n4037, n4034, n4039, n3972, n3969, n3929,
         n3926, n3863, n3860, n4003, n4002, n4032, n4035, n3797, n3792, n3790,
         n3795, n3891, n3893, n3827, n3826, n3896, n4007, n3931, n3793, n3924,
         n3831, n3829, n3927, n3974, n3898, n3970, n4000, n3865, n3861, n3824,
         n3894, n3967, n3858, n4005, n3395, n4956, n5026, n3941, n3733, n3660,
         n4798, n4805, n4175, n3734, n4193, n3739, n3738, n3669, n4721, n4523,
         n4524, n4526, n2573, n2577, n2563, n2567, n4938, n4940, n4913, n4915,
         n4714, n4516, n4517, n5111, n4819, n3730, n3121, n3180, n4305, n4283,
         n2608, n4447, n4448, n4402, n4403, n4425, n4426, n4436, n4437, n4391,
         n4392, n4379, n4380, n4414, n4415, n4458, n4459, n5016, n5014, n3064,
         n3065, n4535, n5112, n3675, counter_31, counter_30, counter_29,
         counter_28, counter_27, counter_26, counter_25, counter_24,
         counter_23, counter_22, counter_21, counter_20, counter_19,
         counter_18, counter_17, counter_16, counter_15, counter_14,
         counter_13, counter_12, counter_11, counter_10, counter_9, counter_8,
         counter_7, counter_6, counter_5, counter_4, counter_3, counter_2,
         counter_1, counter_0, carry_31, carry_30, carry_29, carry_28,
         carry_27, carry_26, carry_25, carry_24, carry_23, carry_22, carry_21,
         carry_20, carry_19, carry_18, carry_17, carry_16, carry_15, carry_14,
         carry_13, carry_12, carry_11, carry_10, carry_9, carry_8, carry_7,
         carry_6, carry_5, carry_4, carry_3, carry_2, N31, N5, N6, N7, N8, N9,
         N10, N11, N12, N13, N14, N15, N23, N24, N25, N26, N2, N3, N4, N16,
         N17, N18, N19, N20, N21, N22, N27, N28, N29, N30, N1, N32, n37, n87,
         n73, n86, n85, n84, n83, n82, n81, n80, n79, n78, n77, n76, n75, n74,
         n58, n59, n60, n61, n62, n63, n64, Trigger_out, n65, n66, n67, n68,
         n69, n70, n71, n72, n3, n8, n36, n39, n42, g33959, n195, n291, n333,
         n364, n365, n380, n401, n408, n475, n490, n549, g25114, n572, n780,
         n783, n787, n870, n1019, n1030, n1282, n1289, n9568, n9569, n9570,
         n9571, n9572, n9573, n9575, n9576, n9577, n9578, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9613, n9614, n9615, n9616, n9617, n9618,
         n9621, n9622, n9623, n9624, n9626, n9627, n9629, n9630, n9633, n9638,
         n9639, n9644, n9645, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9663, n9664, n9665, n9668, n9669, n9671,
         n9673, n9675, n9676, n9677, n9678, n9679, n9685, n9686, n9687, n9688,
         n9689, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9703, n9704,
         n9705, n9706, n9708, n9709, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9774,
         n9775, n9776, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9855, n9856, n9858,
         n9859, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9913, n9914, n9915, n9916, n9918, n9919, n9921, n9922,
         n9924, n9925, n9927, n9928, n9930, n9931, n9933, n9934, n9936, n9937,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9970, n9971,
         n9972, n9973, n9975, n9976, n9977, n9978, n9980, n9981, n9982, n9983,
         n9985, n9986, n9987, n9989, n9990, n9991, n9992, n9994, n9995, n9996,
         n9997, n9999, n10000, n10001, n10002, n10004, n10005, n10006, n10007,
         n10009, n10011, n10013, n10015, n10017, n10021, n10023, n10025,
         n10027, n10028, n10029, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10071,
         n10072, n10073, n10074, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10104, n10105,
         n10106, n10107, n10108, g32975, n10110, n10111, n10112, n10113,
         n10114, n10115, g31862, n10117, g31863, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, U5353_n1, U5355_n1, U5961_n1, U5962_n1,
         U5963_n1, U5964_n1, U5965_n1, U5966_n1, U5967_n1, U5968_n1, U6100_n1,
         U6211_n1, U6212_n1, U6213_n1, U6214_n1, U6215_n1, U6216_n1, U6217_n1,
         U6218_n1, U6279_n1, U6280_n1, U6281_n1, U6282_n1, U6283_n1, U6284_n1,
         U6285_n1, U6286_n1, U6287_n1, U6288_n1, U6289_n1, U6290_n1, U6291_n1,
         U6292_n1, U6338_n1, U6341_n1, U6342_n1, U6343_n1, U6344_n1, U6345_n1,
         U6346_n1, U6347_n1, U6348_n1, U6349_n1, U6350_n1, U6351_n1, U6352_n1,
         U6353_n1, U6354_n1, U6355_n1, U6356_n1, U6357_n1, U6358_n1, U6359_n1,
         U6360_n1, U6361_n1, U6362_n1, U6363_n1, U6364_n1, U6365_n1, U6366_n1,
         U6367_n1, U6368_n1, U6369_n1, U6370_n1, U6371_n1, U6372_n1, U6373_n1,
         U6374_n1, U6375_n1, U6417_n1, U6446_n1, U6465_n1, U6497_n1, U6523_n1,
         U6542_n1, U6552_n1, U6553_n1, U6554_n1, U6555_n1, U6556_n1, U6559_n1,
         U6560_n1, U6561_n1, U6570_n1, U6911_n1, U6912_n1, U6917_n1, U6926_n1,
         U6927_n1, U6929_n1, U6931_n1, U6932_n1, U6933_n1, U6934_n1, U6935_n1,
         U6936_n1, U6937_n1, U6938_n1, U6939_n1, U6940_n1, U6941_n1, U6944_n1,
         U6950_n1, U6954_n1, U6955_n1, U6956_n1, U6957_n1, U7174_n1, U7248_n1,
         U7249_n1, U7402_n1, U7405_n1, U7413_n1, U7416_n1, U7427_n1, U7438_n1,
         U7449_n1, U7455_n1, U7464_n1, U7467_n1, U7482_n1, U7492_n1, U7513_n1,
         U7516_n1, U7549_n1, U7561_n1, U7574_n1, U7577_n1, U7585_n1, U7595_n1,
         U7614_n1, U7621_n1, U7629_n1, U7636_n1, U7639_n1, U7649_n1, U7652_n1,
         U7668_n1, U7673_n1, U7690_n1, U7707_n1, U7712_n1, U7792_n1, U7794_n1,
         U7895_n1, U7897_n1, U7977_n1, U8034_n1, U8036_n1, U8050_n1, U8055_n1,
         U8060_n1, U8070_n1, U8074_n1, U8088_n1, U8112_n1, U8113_n1, U8147_n1,
         U8165_n1, U8185_n1, U8192_n1, U8210_n1, U8223_n1, U8224_n1, U8281_n1,
         U8307_n1, U8974_n1, U8975_n1, U9065_n1, U9070_n1, U9075_n1, U9076_n1,
         U9080_n1, U9084_n1, U9085_n1, U9086_n1, U9090_n1, U9098_n1, U9099_n1,
         U9101_n1, U9107_n1, U9111_n1, U9116_n1, U9120_n1, U9124_n1, U9128_n1,
         U9132_n1, U9136_n1, U9315_n1, U9453_n1, U9825_n1, U9886_n1, U9927_n1,
         U9953_n1, U9957_n1, U9958_n1, U9968_n1, U9972_n1, U9992_n1, U10314_n1,
         U10318_n1;
  assign g34240 = 1'b1;
  assign g34239 = 1'b1;
  assign g34238 = 1'b1;
  assign g34237 = 1'b1;
  assign g34236 = 1'b1;
  assign g34235 = 1'b1;
  assign g34234 = 1'b1;
  assign g34233 = 1'b1;
  assign g34232 = 1'b1;
  assign g33950 = 1'b1;
  assign g33949 = 1'b1;
  assign g33948 = 1'b1;
  assign g33947 = 1'b1;
  assign g33946 = 1'b1;
  assign g33945 = 1'b1;
  assign g32454 = 1'b1;
  assign g32429 = 1'b1;
  assign g25590 = 1'b1;
  assign g25589 = 1'b1;
  assign g25588 = 1'b1;
  assign g25587 = 1'b1;
  assign g25586 = 1'b1;
  assign g25585 = 1'b1;
  assign g25584 = 1'b1;
  assign g25583 = 1'b1;
  assign g25582 = 1'b1;
  assign g24151 = 1'b1;
  assign g34597 = 1'b0;
  assign g24173 = g100;
  assign g24174 = g113;
  assign g24175 = g114;
  assign g24176 = g115;
  assign g24177 = g116;
  assign g24178 = g120;
  assign g24179 = g124;
  assign g24180 = g125;
  assign g24181 = g126;
  assign g24182 = g127;
  assign g24183 = g134;
  assign g24184 = g135;
  assign g29218 = g18881;
  assign g30329 = g23612;
  assign g30330 = g23652;
  assign g24167 = g73;
  assign g20763 = g29211;
  assign g20899 = g29212;
  assign g20557 = g29213;
  assign g20652 = g29214;
  assign g20901 = g29215;
  assign g21176 = g29216;
  assign g21270 = g29217;
  assign g20654 = g29219;
  assign g21245 = g29220;
  assign g21292 = g29221;
  assign g23002 = g30327;
  assign g23759 = g30331;
  assign g23683 = g30332;
  assign g34436 = g31656;
  assign g34437 = g31665;
  assign g27831 = g33533;
  assign g31521 = g34435;
  assign g33894 = g34788;
  assign g34956 = g34839;
  assign g21698 = g36;
  assign g24185 = g44;
  assign g24161 = g53;
  assign g24162 = g54;
  assign g24163 = g56;
  assign g24164 = g57;
  assign g24165 = g64;
  assign g18098 = g6744;
  assign g18099 = g6745;
  assign g18101 = g6746;
  assign g18097 = g6747;
  assign g18094 = g6748;
  assign g18095 = g6749;
  assign g18096 = g6750;
  assign g18100 = g6751;
  assign g18092 = g6753;
  assign g24168 = g84;
  assign g24169 = g90;
  assign g24170 = g91;
  assign g24171 = g92;
  assign g24172 = g99;
  assign g31861 = test_so10;
  assign g25219 = test_so10;
  assign g13881 = test_so26;
  assign g9615 = test_so35;
  assign g8785 = test_so39;
  assign g8291 = test_so42;
  assign g17316 = test_so44;
  assign g8178 = test_so46;
  assign g12470 = test_so80;
  assign g11447 = test_so86;
  assign g9682 = test_so92;
  assign g29210 = test_so100;
  assign g20049 = test_so100;
  assign g24166 = g72;
  assign g28753 = g33959;
  assign g31860 = g25114;
  assign g26801 = g32975;
  assign g25259 = g31862;
  assign g25167 = g31863;

  SDFFX1 DFF_0_Q_reg ( .D(g33046), .SI(test_si1), .SE(n10165), .CLK(n10517), 
        .Q(g5057), .QN(n5615) );
  SDFFX1 DFF_1_Q_reg ( .D(g34441), .SI(g5057), .SE(n10267), .CLK(n10619), .Q(
        g2771), .QN(n5544) );
  SDFFX1 DFF_2_Q_reg ( .D(g33982), .SI(g2771), .SE(n10203), .CLK(n10555), .Q(
        g1882) );
  SDFFX1 DFF_4_Q_reg ( .D(g34007), .SI(g1882), .SE(n10263), .CLK(n10615), .Q(
        g2299), .QN(n9644) );
  SDFFX1 DFF_5_Q_reg ( .D(g24276), .SI(g2299), .SE(n10200), .CLK(n10552), .Q(
        g4040), .QN(n5530) );
  SDFFX1 DFF_6_Q_reg ( .D(g30381), .SI(g4040), .SE(n10207), .CLK(n10559), .Q(
        g2547), .QN(n5782) );
  SDFFX1 DFF_7_Q_reg ( .D(g9048), .SI(g2547), .SE(n10223), .CLK(n10575), .Q(
        g559) );
  SDFFX1 DFF_9_Q_reg ( .D(g30405), .SI(g559), .SE(n10232), .CLK(n10584), .Q(
        g3243), .QN(n9843) );
  SDFFX1 DFF_10_Q_reg ( .D(g25604), .SI(g3243), .SE(n10184), .CLK(n10536), .Q(
        g452), .QN(n9914) );
  SDFFX1 DFF_12_Q_reg ( .D(g30416), .SI(g452), .SE(n10184), .CLK(n10536), .Q(
        g3542), .QN(n9805) );
  SDFFX1 DFF_13_Q_reg ( .D(g30466), .SI(g3542), .SE(n10216), .CLK(n10568), .Q(
        g5232), .QN(n9921) );
  SDFFX1 DFF_14_Q_reg ( .D(g25736), .SI(g5232), .SE(n10245), .CLK(n10597), .Q(
        g5813) );
  SDFFX1 DFF_15_Q_reg ( .D(g34617), .SI(g5813), .SE(n10198), .CLK(n10550), .Q(
        test_so1), .QN(n10146) );
  SDFFX1 DFF_16_Q_reg ( .D(g33974), .SI(test_si2), .SE(n10254), .CLK(n10606), 
        .Q(g1744), .QN(n5795) );
  SDFFX1 DFF_17_Q_reg ( .D(g30505), .SI(g1744), .SE(n10187), .CLK(n10539), .Q(
        g5909), .QN(n9925) );
  SDFFX1 DFF_18_Q_reg ( .D(g33554), .SI(g5909), .SE(n10254), .CLK(n10606), .Q(
        g1802), .QN(n5536) );
  SDFFX1 DFF_19_Q_reg ( .D(g30432), .SI(g1802), .SE(n10184), .CLK(n10536), .Q(
        g3554), .QN(n10001) );
  SDFFX1 DFF_20_Q_reg ( .D(g33064), .SI(g3554), .SE(n10242), .CLK(n10594), .Q(
        g6219), .QN(n5385) );
  SDFFX1 DFF_21_Q_reg ( .D(g34881), .SI(g6219), .SE(n10259), .CLK(n10611), .Q(
        g807), .QN(n5479) );
  SDFFX1 DFF_22_Q_reg ( .D(g17715), .SI(g807), .SE(n10260), .CLK(n10612), .Q(
        g6031) );
  SDFFX1 DFF_23_Q_reg ( .D(g24216), .SI(g6031), .SE(n10171), .CLK(n10523), .Q(
        g847), .QN(n5709) );
  SDFFX1 DFF_24_Q_reg ( .D(g24232), .SI(g847), .SE(n10232), .CLK(n10584), .Q(
        n9367), .QN(DFF_24_n1) );
  SDFFX1 DFF_25_Q_reg ( .D(g34733), .SI(n9367), .SE(n10232), .CLK(n10584), .Q(
        g4172) );
  SDFFX1 DFF_26_Q_reg ( .D(g34882), .SI(g4172), .SE(n10173), .CLK(n10525), .Q(
        g4372) );
  SDFFX1 DFF_27_Q_reg ( .D(g33026), .SI(g4372), .SE(n10173), .CLK(n10525), .Q(
        g3512), .QN(n10058) );
  SDFFX1 DFF_28_Q_reg ( .D(g31867), .SI(g3512), .SE(n10191), .CLK(n10543), .Q(
        test_so2), .QN(n5471) );
  SDFFX1 DFF_29_Q_reg ( .D(g25668), .SI(test_si3), .SE(n10173), .CLK(n10525), 
        .Q(g3490), .QN(n5454) );
  SDFFX1 DFF_30_Q_reg ( .D(g24344), .SI(g3490), .SE(n10185), .CLK(n10537), .Q(
        g12350), .QN(n5432) );
  SDFFX1 DFF_31_Q_reg ( .D(g8920), .SI(g12350), .SE(n10219), .CLK(n10571), .Q(
        g4235), .QN(n9834) );
  SDFFX1 DFF_32_Q_reg ( .D(g33966), .SI(g4235), .SE(n10219), .CLK(n10571), .Q(
        g1600), .QN(n5811) );
  SDFFX1 DFF_33_Q_reg ( .D(g33550), .SI(g1600), .SE(n10221), .CLK(n10573), .Q(
        g1714), .QN(n5460) );
  SDFFX1 DFF_34_Q_reg ( .D(g16656), .SI(g1714), .SE(n10221), .CLK(n10573), .Q(
        g14451), .QN(n10028) );
  SDFFX1 DFF_35_Q_reg ( .D(g30393), .SI(g14451), .SE(n10246), .CLK(n10598), 
        .Q(g3155), .QN(n5366) );
  SDFFX1 DFF_37_Q_reg ( .D(g29248), .SI(g3155), .SE(n10209), .CLK(n10561), .Q(
        g2236), .QN(n9822) );
  SDFFX1 DFF_38_Q_reg ( .D(g4571), .SI(g2236), .SE(n10244), .CLK(n10596), .Q(
        g4555) );
  SDFFX1 DFF_39_Q_reg ( .D(g24274), .SI(g4555), .SE(n10168), .CLK(n10520), .Q(
        g3698), .QN(n9901) );
  SDFFX1 DFF_41_Q_reg ( .D(g33973), .SI(g3698), .SE(n10254), .CLK(n10606), .Q(
        g1736), .QN(n5817) );
  SDFFX1 DFF_42_Q_reg ( .D(g30360), .SI(g1736), .SE(n10169), .CLK(n10521), .Q(
        g1968), .QN(n5664) );
  SDFFX1 DFF_43_Q_reg ( .D(g34460), .SI(g1968), .SE(n10224), .CLK(n10576), .Q(
        test_so3), .QN(n10138) );
  SDFFX1 DFF_44_Q_reg ( .D(g30494), .SI(test_si4), .SE(n10271), .CLK(n10623), 
        .Q(g5607), .QN(n9873) );
  SDFFX1 DFF_45_Q_reg ( .D(g30384), .SI(g5607), .SE(n10177), .CLK(n10529), .Q(
        g2657), .QN(n5316) );
  SDFFX1 DFF_46_Q_reg ( .D(g24340), .SI(g2657), .SE(n10182), .CLK(n10534), .Q(
        g12300), .QN(n5439) );
  SDFFX1 DFF_47_Q_reg ( .D(g29223), .SI(g12300), .SE(n10238), .CLK(n10590), 
        .Q(g490), .QN(n5708) );
  SDFFX1 DFF_48_Q_reg ( .D(g26881), .SI(g490), .SE(n10238), .CLK(n10590), .Q(
        g311), .QN(n5317) );
  SDFFX1 DFF_50_Q_reg ( .D(g34252), .SI(g311), .SE(n10238), .CLK(n10590), .Q(
        g772), .QN(n5334) );
  SDFFX1 DFF_51_Q_reg ( .D(g30489), .SI(g772), .SE(n10180), .CLK(n10532), .Q(
        g5587), .QN(n9945) );
  SDFFX1 DFF_52_Q_reg ( .D(g29301), .SI(g5587), .SE(n10179), .CLK(n10531), .Q(
        g6177), .QN(n5874) );
  SDFFX1 DFF_53_Q_reg ( .D(g17743), .SI(g6177), .SE(n10235), .CLK(n10587), .Q(
        g6377) );
  SDFFX1 DFF_54_Q_reg ( .D(g33022), .SI(g6377), .SE(n10235), .CLK(n10587), .Q(
        g3167), .QN(n5652) );
  SDFFX1 DFF_55_Q_reg ( .D(g30496), .SI(g3167), .SE(n10174), .CLK(n10526), .Q(
        g5615), .QN(n9851) );
  SDFFX1 DFF_56_Q_reg ( .D(g33043), .SI(g5615), .SE(n10243), .CLK(n10595), .Q(
        g4567) );
  SDFFX1 DFF_58_Q_reg ( .D(g29263), .SI(g4567), .SE(n10173), .CLK(n10525), .Q(
        test_so4), .QN(n10144) );
  SDFFX1 DFF_59_Q_reg ( .D(g30533), .SI(test_si5), .SE(n10227), .CLK(n10579), 
        .Q(g6287), .QN(n10002) );
  SDFFX1 DFF_60_Q_reg ( .D(g24256), .SI(g6287), .SE(n10227), .CLK(n10579), .Q(
        g7946), .QN(n5302) );
  SDFFX1 DFF_61_Q_reg ( .D(g34015), .SI(g7946), .SE(n10249), .CLK(n10601), .Q(
        g2563), .QN(n5816) );
  SDFFX1 DFF_62_Q_reg ( .D(g34031), .SI(g2563), .SE(n10259), .CLK(n10611), .Q(
        g4776), .QN(n5707) );
  SDFFX1 DFF_63_Q_reg ( .D(g34452), .SI(g4776), .SE(n10259), .CLK(n10611), .Q(
        g4593), .QN(n5303) );
  SDFFX1 DFF_64_Q_reg ( .D(g34646), .SI(g4593), .SE(n10259), .CLK(n10611), .Q(
        g6199), .QN(n5644) );
  SDFFX1 DFF_65_Q_reg ( .D(g34001), .SI(g6199), .SE(n10263), .CLK(n10615), .Q(
        g2295), .QN(n5815) );
  SDFFX1 DFF_66_Q_reg ( .D(g25633), .SI(g2295), .SE(n10201), .CLK(n10553), .Q(
        g1384), .QN(n9592) );
  SDFFX1 DFF_67_Q_reg ( .D(g24259), .SI(g1384), .SE(n10229), .CLK(n10581), .Q(
        g1339), .QN(n5381) );
  SDFFX1 DFF_68_Q_reg ( .D(g33049), .SI(g1339), .SE(n10250), .CLK(n10602), .Q(
        g5180), .QN(n5384) );
  SDFFX1 DFF_69_Q_reg ( .D(g34609), .SI(g5180), .SE(n10250), .CLK(n10602), .Q(
        g2844), .QN(n10078) );
  SDFFX1 DFF_70_Q_reg ( .D(g31869), .SI(g2844), .SE(n10250), .CLK(n10602), .Q(
        g1024), .QN(n9728) );
  SDFFX1 DFF_71_Q_reg ( .D(g30490), .SI(g1024), .SE(n10271), .CLK(n10623), .Q(
        test_so5), .QN(n10147) );
  SDFFX1 DFF_72_Q_reg ( .D(g30427), .SI(test_si6), .SE(n10242), .CLK(n10594), 
        .Q(g3598), .QN(n9803) );
  SDFFX1 DFF_73_Q_reg ( .D(g21894), .SI(g3598), .SE(n10242), .CLK(n10594), .Q(
        g4264), .QN(n5823) );
  SDFFX1 DFF_74_Q_reg ( .D(g33965), .SI(g4264), .SE(n10191), .CLK(n10543), .Q(
        g767), .QN(n5333) );
  SDFFX1 DFF_75_Q_reg ( .D(g34645), .SI(g767), .SE(n10191), .CLK(n10543), .Q(
        g5853), .QN(n5499) );
  SDFFX1 DFF_76_Q_reg ( .D(g16874), .SI(g5853), .SE(n10200), .CLK(n10552), .Q(
        g13865), .QN(n5580) );
  SDFFX1 DFF_77_Q_reg ( .D(g33571), .SI(g13865), .SE(n10213), .CLK(n10565), 
        .Q(g2089), .QN(n9655) );
  SDFFX1 DFF_78_Q_reg ( .D(g34267), .SI(g2089), .SE(n10205), .CLK(n10557), .Q(
        g4933), .QN(n5878) );
  SDFFX1 DFF_79_Q_reg ( .D(g26971), .SI(g4933), .SE(n10205), .CLK(n10557), .Q(
        g4521), .QN(n5752) );
  SDFFX1 DFF_80_Q_reg ( .D(g34644), .SI(g4521), .SE(n10205), .CLK(n10557), .Q(
        g5507), .QN(n5643) );
  SDFFX1 DFF_81_Q_reg ( .D(g16627), .SI(g5507), .SE(n10222), .CLK(n10574), .Q(
        g16656), .QN(n10000) );
  SDFFX1 DFF_82_Q_reg ( .D(g30534), .SI(g16656), .SE(n10226), .CLK(n10578), 
        .Q(g6291), .QN(n9864) );
  SDFFX1 DFF_83_Q_reg ( .D(g33535), .SI(g6291), .SE(n10263), .CLK(n10615), .Q(
        g294), .QN(n5680) );
  SDFFX1 DFF_84_Q_reg ( .D(g30498), .SI(g294), .SE(n10271), .CLK(n10623), .Q(
        test_so6) );
  SDFFX1 DFF_85_Q_reg ( .D(g25728), .SI(test_si7), .SE(n10244), .CLK(n10596), 
        .Q(g9617), .QN(n5722) );
  SDFFX1 DFF_86_Q_reg ( .D(g25743), .SI(g9617), .SE(n10220), .CLK(n10572), .Q(
        g9741) );
  SDFFX1 DFF_87_Q_reg ( .D(g25684), .SI(g9741), .SE(n10220), .CLK(n10572), .Q(
        g3813) );
  SDFFX1 DFF_88_Q_reg ( .D(g25613), .SI(g3813), .SE(n10220), .CLK(n10572), .Q(
        g562), .QN(n9584) );
  SDFFX1 DFF_89_Q_reg ( .D(g34438), .SI(g562), .SE(n10222), .CLK(n10574), .Q(
        g608), .QN(n5475) );
  SDFFX1 DFF_90_Q_reg ( .D(g24244), .SI(g608), .SE(n10240), .CLK(n10592), .Q(
        g1205), .QN(n5547) );
  SDFFX1 DFF_91_Q_reg ( .D(g30439), .SI(g1205), .SE(n10183), .CLK(n10535), .Q(
        g3909), .QN(n9931) );
  SDFFX1 DFF_92_Q_reg ( .D(g30541), .SI(g3909), .SE(n10225), .CLK(n10577), .Q(
        g6259), .QN(n10031) );
  SDFFX1 DFF_93_Q_reg ( .D(g30519), .SI(g6259), .SE(n10187), .CLK(n10539), .Q(
        g5905), .QN(n9982) );
  SDFFX1 DFF_94_Q_reg ( .D(g25621), .SI(g5905), .SE(n10196), .CLK(n10548), .Q(
        g921), .QN(n9740) );
  SDFFX1 DFF_95_Q_reg ( .D(g34807), .SI(g921), .SE(n10165), .CLK(n10517), .Q(
        g2955), .QN(n9733) );
  SDFFX1 DFF_96_Q_reg ( .D(g25599), .SI(g2955), .SE(n10255), .CLK(n10607), .Q(
        g203) );
  SDFFX1 DFF_98_Q_reg ( .D(g24235), .SI(g203), .SE(n10255), .CLK(n10607), .Q(
        test_so7) );
  SDFFX1 DFF_99_Q_reg ( .D(g34036), .SI(test_si8), .SE(n10225), .CLK(n10577), 
        .Q(g4878), .QN(n5283) );
  SDFFX1 DFF_100_Q_reg ( .D(g30476), .SI(g4878), .SE(n10253), .CLK(n10605), 
        .Q(g5204), .QN(n9952) );
  SDFFX1 DFF_101_Q_reg ( .D(g17580), .SI(g5204), .SE(n10233), .CLK(n10585), 
        .Q(g17604), .QN(n9986) );
  SDFFX1 DFF_102_Q_reg ( .D(g30429), .SI(g17604), .SE(n10184), .CLK(n10536), 
        .Q(g3606), .QN(n9999) );
  SDFFX1 DFF_103_Q_reg ( .D(g32997), .SI(g3606), .SE(n10228), .CLK(n10580), 
        .Q(g1926), .QN(n5510) );
  SDFFX1 DFF_104_Q_reg ( .D(g33063), .SI(g1926), .SE(n10228), .CLK(n10580), 
        .Q(g6215), .QN(n5651) );
  SDFFX1 DFF_105_Q_reg ( .D(g30424), .SI(g6215), .SE(n10184), .CLK(n10536), 
        .Q(g3586), .QN(n9893) );
  SDFFX1 DFF_106_Q_reg ( .D(g32977), .SI(g3586), .SE(n10260), .CLK(n10612), 
        .Q(g291), .QN(n5679) );
  SDFFX1 DFF_107_Q_reg ( .D(g34026), .SI(g291), .SE(n10260), .CLK(n10612), .Q(
        g4674), .QN(n5440) );
  SDFFX1 DFF_108_Q_reg ( .D(g30420), .SI(g4674), .SE(n10184), .CLK(n10536), 
        .Q(g3570), .QN(n9841) );
  SDFFX1 DFF_109_Q_reg ( .D(g12368), .SI(g3570), .SE(n10223), .CLK(n10575), 
        .Q(g9048), .QN(n9570) );
  SDFFX1 DFF_110_Q_reg ( .D(g17739), .SI(g9048), .SE(n10223), .CLK(n10575), 
        .Q(g17607), .QN(n9870) );
  SDFFX1 DFF_111_Q_reg ( .D(g33560), .SI(g17607), .SE(n10268), .CLK(n10620), 
        .Q(test_so8), .QN(n10137) );
  SDFFX1 DFF_112_Q_reg ( .D(g29226), .SI(test_si9), .SE(n10199), .CLK(n10551), 
        .Q(g676), .QN(n5751) );
  SDFFX1 DFF_113_Q_reg ( .D(g25619), .SI(g676), .SE(n10199), .CLK(n10551), .Q(
        g843), .QN(n9713) );
  SDFFX1 DFF_115_Q_reg ( .D(g34455), .SI(g843), .SE(n10199), .CLK(n10551), .Q(
        g4332), .QN(n5540) );
  SDFFX1 DFF_116_Q_reg ( .D(g30457), .SI(g4332), .SE(n10233), .CLK(n10585), 
        .Q(g4153), .QN(n10094) );
  SDFFX1 DFF_117_Q_reg ( .D(g14694), .SI(g4153), .SE(n10233), .CLK(n10585), 
        .Q(g17711), .QN(n9887) );
  SDFFX1 DFF_118_Q_reg ( .D(g33625), .SI(g17711), .SE(n10179), .CLK(n10531), 
        .Q(g6336), .QN(n5592) );
  SDFFX1 DFF_119_Q_reg ( .D(g34790), .SI(g6336), .SE(n10223), .CLK(n10575), 
        .Q(g622), .QN(n5672) );
  SDFFX1 DFF_120_Q_reg ( .D(g30414), .SI(g622), .SE(n10241), .CLK(n10593), .Q(
        g3506), .QN(n5576) );
  SDFFX1 DFF_121_Q_reg ( .D(g26966), .SI(g3506), .SE(n10244), .CLK(n10596), 
        .Q(g4558) );
  SDFFX1 DFF_123_Q_reg ( .D(g17649), .SI(g4558), .SE(n10244), .CLK(n10596), 
        .Q(g17685), .QN(n10005) );
  SDFFX1 DFF_124_Q_reg ( .D(g25656), .SI(g17685), .SE(n10256), .CLK(n10608), 
        .Q(g3111) );
  SDFFX1 DFF_125_Q_reg ( .D(g30390), .SI(g3111), .SE(n10256), .CLK(n10608), 
        .Q(g29217) );
  SDFFX1 DFF_126_Q_reg ( .D(g25688), .SI(g29217), .SE(n10256), .CLK(n10608), 
        .Q(test_so9), .QN(n18470) );
  SDFFX1 DFF_127_Q_reg ( .D(g34727), .SI(test_si10), .SE(n10197), .CLK(n10549), 
        .Q(g939), .QN(n5415) );
  SDFFX1 DFF_128_Q_reg ( .D(g25594), .SI(g939), .SE(n10248), .CLK(n10600), .Q(
        g278), .QN(n5627) );
  SDFFX1 DFF_129_Q_reg ( .D(g26963), .SI(g278), .SE(n10248), .CLK(n10600), .Q(
        g4492), .QN(n10061) );
  SDFFX1 DFF_130_Q_reg ( .D(g34034), .SI(g4492), .SE(n10224), .CLK(n10576), 
        .Q(g4864), .QN(n5318) );
  SDFFX1 DFF_131_Q_reg ( .D(g33541), .SI(g4864), .SE(n10191), .CLK(n10543), 
        .Q(g1036), .QN(n9686) );
  SDFFX1 DFF_132_Q_reg ( .D(g28093), .SI(g1036), .SE(n10217), .CLK(n10569), 
        .Q(g29220) );
  SDFFX1 DFF_133_Q_reg ( .D(g24236), .SI(g29220), .SE(n10217), .CLK(n10569), 
        .Q(g1178), .QN(n9756) );
  SDFFX1 DFF_134_Q_reg ( .D(g30404), .SI(g1178), .SE(n10231), .CLK(n10583), 
        .Q(g3239), .QN(n9968) );
  SDFFX1 DFF_135_Q_reg ( .D(g28051), .SI(g3239), .SE(n10237), .CLK(n10589), 
        .Q(g718), .QN(n9819) );
  SDFFX1 DFF_136_Q_reg ( .D(g29303), .SI(g718), .SE(n10242), .CLK(n10594), .Q(
        g6195) );
  SDFFX1 DFF_137_Q_reg ( .D(g26917), .SI(g6195), .SE(n10166), .CLK(n10518), 
        .Q(g1135), .QN(n5328) );
  SDFFX1 DFF_139_Q_reg ( .D(g33624), .SI(g1135), .SE(n10261), .CLK(n10613), 
        .Q(g6395), .QN(n5396) );
  SDFFX1 DFF_141_Q_reg ( .D(g24337), .SI(g6395), .SE(n10207), .CLK(n10559), 
        .Q(test_so10), .QN(n10129) );
  SDFFX1 DFF_142_Q_reg ( .D(g34911), .SI(test_si11), .SE(n10261), .CLK(n10613), 
        .Q(g554), .QN(n9708) );
  SDFFX1 DFF_143_Q_reg ( .D(g33963), .SI(g554), .SE(n10190), .CLK(n10542), .Q(
        g496) );
  SDFFX1 DFF_144_Q_reg ( .D(g34627), .SI(g496), .SE(n10190), .CLK(n10542), .Q(
        g3853), .QN(n5641) );
  SDFFX1 DFF_145_Q_reg ( .D(g29282), .SI(g3853), .SE(n10262), .CLK(n10614), 
        .Q(g5134), .QN(n5807) );
  SDFFX1 DFF_146_Q_reg ( .D(g17320), .SI(g5134), .SE(n10262), .CLK(n10614), 
        .Q(g17404), .QN(n9736) );
  SDFFX1 DFF_147_Q_reg ( .D(g25676), .SI(g17404), .SE(n10262), .CLK(n10614), 
        .Q(g8344), .QN(n5721) );
  SDFFX1 DFF_148_Q_reg ( .D(g33013), .SI(g8344), .SE(n10268), .CLK(n10620), 
        .Q(g2485), .QN(n5509) );
  SDFFX1 DFF_149_Q_reg ( .D(g32981), .SI(g2485), .SE(n10197), .CLK(n10549), 
        .Q(g925), .QN(n5725) );
  SDFFX1 DFF_150_Q_reg ( .D(g34976), .SI(g925), .SE(n10175), .CLK(n10527), .Q(
        n9357) );
  SDFFX1 DFF_151_Q_reg ( .D(g30483), .SI(n9357), .SE(n10175), .CLK(n10527), 
        .Q(g5555), .QN(n10017) );
  SDFFX1 DFF_152_Q_reg ( .D(g14217), .SI(g5555), .SE(n10247), .CLK(n10599), 
        .Q(g14096), .QN(n9594) );
  SDFFX1 DFF_153_Q_reg ( .D(g32994), .SI(g14096), .SE(n10208), .CLK(n10560), 
        .Q(g1798), .QN(n5833) );
  SDFFX1 DFF_154_Q_reg ( .D(g28070), .SI(g1798), .SE(n10239), .CLK(n10591), 
        .Q(test_so11) );
  SDFFX1 DFF_155_Q_reg ( .D(g34806), .SI(test_si12), .SE(n10183), .CLK(n10535), 
        .Q(g2941), .QN(n10084) );
  SDFFX1 DFF_156_Q_reg ( .D(g30453), .SI(g2941), .SE(n10183), .CLK(n10535), 
        .Q(g3905), .QN(n9991) );
  SDFFX1 DFF_157_Q_reg ( .D(g33539), .SI(g3905), .SE(n10191), .CLK(n10543), 
        .Q(g763), .QN(n5332) );
  SDFFX1 DFF_158_Q_reg ( .D(g30526), .SI(g763), .SE(n10225), .CLK(n10577), .Q(
        g6255), .QN(n9940) );
  SDFFX1 DFF_159_Q_reg ( .D(g26951), .SI(g6255), .SE(n10172), .CLK(n10524), 
        .Q(g4375), .QN(n9578) );
  SDFFX1 DFF_160_Q_reg ( .D(g34035), .SI(g4375), .SE(n10225), .CLK(n10577), 
        .Q(g4871), .QN(n5443) );
  SDFFX1 DFF_161_Q_reg ( .D(g34636), .SI(g4871), .SE(n10234), .CLK(n10586), 
        .Q(g4722), .QN(n5345) );
  SDFFX1 DFF_162_Q_reg ( .D(g32978), .SI(g4722), .SE(n10222), .CLK(n10574), 
        .Q(g590), .QN(n5472) );
  SDFFX1 DFF_163_Q_reg ( .D(g17722), .SI(g590), .SE(n10264), .CLK(n10616), .Q(
        g13099) );
  SDFFX1 DFF_164_Q_reg ( .D(g30348), .SI(g13099), .SE(n10219), .CLK(n10571), 
        .Q(g1632), .QN(n5836) );
  SDFFX1 DFF_165_Q_reg ( .D(g24336), .SI(g1632), .SE(n10207), .CLK(n10559), 
        .Q(g12238), .QN(n5438) );
  SDFFX1 DFF_166_Q_reg ( .D(g8215), .SI(g12238), .SE(n10207), .CLK(n10559), 
        .Q(g3100) );
  SDFFX1 DFF_167_Q_reg ( .D(g24250), .SI(g3100), .SE(n10236), .CLK(n10588), 
        .Q(test_so12) );
  SDFFX1 DFF_169_Q_reg ( .D(g29236), .SI(test_si13), .SE(n10236), .CLK(n10588), 
        .Q(g1437), .QN(n5696) );
  SDFFX1 DFF_170_Q_reg ( .D(g29298), .SI(g1437), .SE(n10179), .CLK(n10531), 
        .Q(g6154), .QN(n5747) );
  SDFFX1 DFF_171_Q_reg ( .D(g10527), .SI(g6154), .SE(n10212), .CLK(n10564), 
        .Q(g1579), .QN(n9722) );
  SDFFX1 DFF_172_Q_reg ( .D(g30499), .SI(g1579), .SE(n10175), .CLK(n10527), 
        .Q(g5567), .QN(n10015) );
  SDFFX1 DFF_173_Q_reg ( .D(g33976), .SI(g5567), .SE(n10228), .CLK(n10580), 
        .Q(g1752), .QN(n5797) );
  SDFFX1 DFF_174_Q_reg ( .D(g32996), .SI(g1752), .SE(n10228), .CLK(n10580), 
        .Q(g1917), .QN(n10044) );
  SDFFX1 DFF_175_Q_reg ( .D(g30335), .SI(g1917), .SE(n10228), .CLK(n10580), 
        .Q(g744), .QN(n5470) );
  SDFFX1 DFF_177_Q_reg ( .D(g34637), .SI(g744), .SE(n10234), .CLK(n10586), .Q(
        g4737), .QN(n5867) );
  SDFFX1 DFF_178_Q_reg ( .D(g25694), .SI(g4737), .SE(n10234), .CLK(n10586), 
        .Q(g8132), .QN(n18466) );
  SDFFX1 DFF_179_Q_reg ( .D(g30528), .SI(g8132), .SE(n10226), .CLK(n10578), 
        .Q(g6267), .QN(n9842) );
  SDFFX1 DFF_181_Q_reg ( .D(g16775), .SI(g6267), .SE(n10236), .CLK(n10588), 
        .Q(g16659), .QN(n9874) );
  SDFFX1 DFF_182_Q_reg ( .D(g24251), .SI(g16659), .SE(n10236), .CLK(n10588), 
        .Q(g1442), .QN(n10049) );
  SDFFX1 DFF_183_Q_reg ( .D(g30521), .SI(g1442), .SE(n10187), .CLK(n10539), 
        .Q(test_so13) );
  SDFFX1 DFF_184_Q_reg ( .D(g26960), .SI(test_si14), .SE(n10195), .CLK(n10547), 
        .Q(g4477), .QN(n5849) );
  SDFFX1 DFF_185_Q_reg ( .D(g24239), .SI(g4477), .SE(n10224), .CLK(n10576), 
        .Q(g10500) );
  SDFFX1 DFF_186_Q_reg ( .D(g34259), .SI(g10500), .SE(n10224), .CLK(n10576), 
        .Q(g4643), .QN(n5382) );
  SDFFX1 DFF_187_Q_reg ( .D(g30474), .SI(g4643), .SE(n10216), .CLK(n10568), 
        .Q(g5264), .QN(n9975) );
  SDFFX1 DFF_188_Q_reg ( .D(g12422), .SI(g5264), .SE(n10220), .CLK(n10572), 
        .Q(g14779), .QN(n5703) );
  SDFFX1 DFF_189_Q_reg ( .D(g33016), .SI(g14779), .SE(n10269), .CLK(n10621), 
        .Q(g2610), .QN(n10042) );
  SDFFX1 DFF_190_Q_reg ( .D(g34643), .SI(g2610), .SE(n10269), .CLK(n10621), 
        .Q(g5160), .QN(n5498) );
  SDFFX1 DFF_192_Q_reg ( .D(g30510), .SI(g5160), .SE(n10269), .CLK(n10621), 
        .Q(g5933), .QN(n9944) );
  SDFFX1 DFF_193_Q_reg ( .D(g29239), .SI(g5933), .SE(n10176), .CLK(n10528), 
        .Q(g1454), .QN(n5866) );
  SDFFX1 DFF_194_Q_reg ( .D(g26897), .SI(g1454), .SE(n10255), .CLK(n10607), 
        .Q(g753), .QN(n9678) );
  SDFFX1 DFF_195_Q_reg ( .D(g34729), .SI(g753), .SE(n10255), .CLK(n10607), .Q(
        g1296), .QN(n9576) );
  SDFFX1 DFF_196_Q_reg ( .D(g34625), .SI(g1296), .SE(n10255), .CLK(n10607), 
        .Q(g3151), .QN(n5495) );
  SDFFX1 DFF_197_Q_reg ( .D(g34800), .SI(g3151), .SE(n10197), .CLK(n10549), 
        .Q(test_so14) );
  SDFFX1 DFF_198_Q_reg ( .D(g24353), .SI(test_si15), .SE(n10196), .CLK(n10548), 
        .Q(g6727), .QN(n5531) );
  SDFFX1 DFF_199_Q_reg ( .D(g33029), .SI(g6727), .SE(n10241), .CLK(n10593), 
        .Q(g3530), .QN(n5569) );
  SDFFX1 DFF_201_Q_reg ( .D(g33615), .SI(g3530), .SE(n10240), .CLK(n10592), 
        .Q(g4104), .QN(n9913) );
  SDFFX1 DFF_202_Q_reg ( .D(g24253), .SI(g4104), .SE(n10229), .CLK(n10581), 
        .Q(g1532), .QN(n9907) );
  SDFFX1 DFF_203_Q_reg ( .D(g24281), .SI(g1532), .SE(n10229), .CLK(n10581), 
        .Q(g9251) );
  SDFFX1 DFF_204_Q_reg ( .D(g33997), .SI(g9251), .SE(n10229), .CLK(n10581), 
        .Q(n9352), .QN(n18471) );
  SDFFX1 DFF_206_Q_reg ( .D(g34971), .SI(n9352), .SE(n10270), .CLK(n10622), 
        .Q(n9351) );
  SDFFX1 DFF_207_Q_reg ( .D(g34263), .SI(n9351), .SE(n10185), .CLK(n10537), 
        .Q(g4754), .QN(n5877) );
  SDFFX1 DFF_208_Q_reg ( .D(g24237), .SI(g4754), .SE(n10185), .CLK(n10537), 
        .Q(g1189), .QN(n5642) );
  SDFFX1 DFF_209_Q_reg ( .D(g33584), .SI(g1189), .SE(n10262), .CLK(n10614), 
        .Q(g2287), .QN(n5353) );
  SDFFX1 DFF_210_Q_reg ( .D(g24280), .SI(g2287), .SE(n10227), .CLK(n10579), 
        .Q(g4273), .QN(n5764) );
  SDFFX1 DFF_211_Q_reg ( .D(g26920), .SI(g4273), .SE(n10201), .CLK(n10553), 
        .Q(g1389), .QN(n9758) );
  SDFFX1 DFF_212_Q_reg ( .D(g33548), .SI(g1389), .SE(n10221), .CLK(n10573), 
        .Q(test_so15), .QN(n10158) );
  SDFFX1 DFF_213_Q_reg ( .D(g29296), .SI(test_si16), .SE(n10181), .CLK(n10533), 
        .Q(g5835), .QN(n5663) );
  SDFFX1 DFF_214_Q_reg ( .D(g30338), .SI(g5835), .SE(n10217), .CLK(n10569), 
        .Q(g1171), .QN(n5363) );
  SDFFX1 DFF_215_Q_reg ( .D(g21895), .SI(g1171), .SE(n10227), .CLK(n10579), 
        .Q(g4269), .QN(n5763) );
  SDFFX1 DFF_216_Q_reg ( .D(g33588), .SI(g4269), .SE(n10176), .CLK(n10528), 
        .Q(g2399), .QN(n5762) );
  SDFFX1 DFF_218_Q_reg ( .D(g34041), .SI(g2399), .SE(n10225), .CLK(n10577), 
        .Q(g4983), .QN(n5367) );
  SDFFX1 DFF_219_Q_reg ( .D(g30495), .SI(g4983), .SE(n10175), .CLK(n10527), 
        .Q(g5611), .QN(n9985) );
  SDFFX1 DFF_220_Q_reg ( .D(g16744), .SI(g5611), .SE(n10222), .CLK(n10574), 
        .Q(g16627), .QN(n9878) );
  SDFFX1 DFF_221_Q_reg ( .D(g29279), .SI(g16627), .SE(n10194), .CLK(n10546), 
        .Q(g4572), .QN(n9677) );
  SDFFX1 DFF_222_Q_reg ( .D(g25655), .SI(g4572), .SE(n10270), .CLK(n10622), 
        .Q(g3143), .QN(n5882) );
  SDFFX1 DFF_223_Q_reg ( .D(g34795), .SI(g3143), .SE(n10166), .CLK(n10518), 
        .Q(g2898), .QN(n10088) );
  SDFFX1 DFF_224_Q_reg ( .D(g24269), .SI(g2898), .SE(n10256), .CLK(n10608), 
        .Q(g3343), .QN(n9897) );
  SDFFX1 DFF_225_Q_reg ( .D(g30403), .SI(g3343), .SE(n10231), .CLK(n10583), 
        .Q(g3235), .QN(n9882) );
  SDFFX1 DFF_226_Q_reg ( .D(g33042), .SI(g3235), .SE(n10242), .CLK(n10594), 
        .Q(test_so16) );
  SDFFX1 DFF_227_Q_reg ( .D(g30419), .SI(test_si17), .SE(n10241), .CLK(n10593), 
        .Q(g3566), .QN(n9804) );
  SDFFX1 DFF_228_Q_reg ( .D(g34023), .SI(g3566), .SE(n10263), .CLK(n10615), 
        .Q(n9348), .QN(DFF_228_n1) );
  SDFFX1 DFF_229_Q_reg ( .D(g28090), .SI(n9348), .SE(n10270), .CLK(n10622), 
        .Q(g4961), .QN(n5770) );
  SDFFX1 DFF_231_Q_reg ( .D(g34642), .SI(g4961), .SE(n10270), .CLK(n10622), 
        .Q(g4927), .QN(n5879) );
  SDFFX1 DFF_232_Q_reg ( .D(g30370), .SI(g4927), .SE(n10193), .CLK(n10545), 
        .Q(g2259), .QN(n5419) );
  SDFFX1 DFF_233_Q_reg ( .D(g34448), .SI(g2259), .SE(n10213), .CLK(n10565), 
        .Q(g2819), .QN(n5609) );
  SDFFX1 DFF_234_Q_reg ( .D(g26946), .SI(g2819), .SE(n10252), .CLK(n10604), 
        .Q(g7257) );
  SDFFX1 DFF_235_Q_reg ( .D(g9617), .SI(g7257), .SE(n10252), .CLK(n10604), .Q(
        g5802) );
  SDFFX1 DFF_236_Q_reg ( .D(g34610), .SI(g5802), .SE(n10253), .CLK(n10605), 
        .Q(g2852), .QN(n10077) );
  SDFFX1 DFF_237_Q_reg ( .D(g24209), .SI(g2852), .SE(n10237), .CLK(n10589), 
        .Q(g417), .QN(n5358) );
  SDFFX1 DFF_238_Q_reg ( .D(g28047), .SI(g417), .SE(n10237), .CLK(n10589), .Q(
        g681), .QN(n9734) );
  SDFFX1 DFF_239_Q_reg ( .D(g24206), .SI(g681), .SE(n10237), .CLK(n10589), .Q(
        g437), .QN(n9747) );
  SDFFX1 DFF_240_Q_reg ( .D(g26891), .SI(g437), .SE(n10239), .CLK(n10591), .Q(
        test_so17), .QN(n10124) );
  SDFFX1 DFF_241_Q_reg ( .D(g30504), .SI(test_si18), .SE(n10187), .CLK(n10539), 
        .Q(g5901), .QN(n10013) );
  SDFFX1 DFF_242_Q_reg ( .D(g34798), .SI(g5901), .SE(n10265), .CLK(n10617), 
        .Q(g2886), .QN(n10086) );
  SDFFX1 DFF_243_Q_reg ( .D(g25669), .SI(g2886), .SE(n10174), .CLK(n10526), 
        .Q(g3494), .QN(n5889) );
  SDFFX1 DFF_244_Q_reg ( .D(g30480), .SI(g3494), .SE(n10174), .CLK(n10526), 
        .Q(g5511), .QN(n5575) );
  SDFFX1 DFF_245_Q_reg ( .D(g33027), .SI(g5511), .SE(n10241), .CLK(n10593), 
        .Q(g3518), .QN(n5645) );
  SDFFX1 DFF_246_Q_reg ( .D(g33972), .SI(g3518), .SE(n10192), .CLK(n10544), 
        .Q(g1604), .QN(n9623) );
  SDFFX1 DFF_248_Q_reg ( .D(g25697), .SI(g1604), .SE(n10165), .CLK(n10517), 
        .Q(g5092) );
  SDFFX1 DFF_249_Q_reg ( .D(g28099), .SI(g5092), .SE(n10188), .CLK(n10540), 
        .Q(g4831), .QN(n9668) );
  SDFFX1 DFF_250_Q_reg ( .D(g26947), .SI(g4831), .SE(n10188), .CLK(n10540), 
        .Q(g4382), .QN(n5714) );
  SDFFX1 DFF_251_Q_reg ( .D(g24350), .SI(g4382), .SE(n10265), .CLK(n10617), 
        .Q(g6386), .QN(n9899) );
  SDFFX1 DFF_252_Q_reg ( .D(g24210), .SI(g6386), .SE(n10265), .CLK(n10617), 
        .Q(g479) );
  SDFFX1 DFF_253_Q_reg ( .D(g30455), .SI(g479), .SE(n10265), .CLK(n10617), .Q(
        g3965), .QN(n9816) );
  SDFFX1 DFF_254_Q_reg ( .D(g28084), .SI(g3965), .SE(n10182), .CLK(n10534), 
        .Q(test_so18) );
  SDFFX1 DFF_255_Q_reg ( .D(g33993), .SI(test_si19), .SE(n10213), .CLK(n10565), 
        .Q(g2008), .QN(n9714) );
  SDFFX1 DFF_256_Q_reg ( .D(g11678), .SI(g2008), .SE(n10213), .CLK(n10565), 
        .Q(g736) );
  SDFFX1 DFF_257_Q_reg ( .D(g30444), .SI(g736), .SE(n10214), .CLK(n10566), .Q(
        g3933), .QN(n9946) );
  SDFFX1 DFF_258_Q_reg ( .D(g33537), .SI(g3933), .SE(n10210), .CLK(n10562), 
        .Q(g222), .QN(n10099) );
  SDFFX1 DFF_259_Q_reg ( .D(g25650), .SI(g222), .SE(n10170), .CLK(n10522), .Q(
        g3050) );
  SDFFX1 DFF_261_Q_reg ( .D(g25625), .SI(g3050), .SE(n10265), .CLK(n10617), 
        .Q(g1052), .QN(n9967) );
  SDFFX1 DFF_263_Q_reg ( .D(g17711), .SI(g1052), .SE(n10233), .CLK(n10585), 
        .Q(g17580), .QN(n9872) );
  SDFFX1 DFF_264_Q_reg ( .D(g30366), .SI(g17580), .SE(n10167), .CLK(n10519), 
        .Q(g2122), .QN(n5784) );
  SDFFX1 DFF_265_Q_reg ( .D(g33593), .SI(g2122), .SE(n10211), .CLK(n10563), 
        .Q(g2465), .QN(n5523) );
  SDFFX1 DFF_267_Q_reg ( .D(g30502), .SI(g2465), .SE(n10244), .CLK(n10596), 
        .Q(g5889), .QN(n9956) );
  SDFFX1 DFF_268_Q_reg ( .D(g33036), .SI(g5889), .SE(n10244), .CLK(n10596), 
        .Q(g4495) );
  SDFFX1 DFF_269_Q_reg ( .D(g25595), .SI(g4495), .SE(n10245), .CLK(n10597), 
        .Q(g8719), .QN(n9786) );
  SDFFX1 DFF_270_Q_reg ( .D(g34462), .SI(g8719), .SE(n10260), .CLK(n10612), 
        .Q(test_so19), .QN(n10133) );
  SDFFX1 DFF_271_Q_reg ( .D(g33024), .SI(test_si20), .SE(n10169), .CLK(n10521), 
        .Q(g3179), .QN(n5390) );
  SDFFX1 DFF_272_Q_reg ( .D(g33552), .SI(g3179), .SE(n10254), .CLK(n10606), 
        .Q(g1728), .QN(n5352) );
  SDFFX1 DFF_273_Q_reg ( .D(g34014), .SI(g1728), .SE(n10206), .CLK(n10558), 
        .Q(g2433), .QN(n9624) );
  SDFFX1 DFF_274_Q_reg ( .D(g29273), .SI(g2433), .SE(n10167), .CLK(n10519), 
        .Q(g3835), .QN(n5662) );
  SDFFX1 DFF_275_Q_reg ( .D(g25748), .SI(g3835), .SE(n10179), .CLK(n10531), 
        .Q(g6187), .QN(n5453) );
  SDFFX1 DFF_276_Q_reg ( .D(g34638), .SI(g6187), .SE(n10180), .CLK(n10532), 
        .Q(g4917), .QN(n5408) );
  SDFFX1 DFF_277_Q_reg ( .D(g30341), .SI(g4917), .SE(n10186), .CLK(n10538), 
        .Q(g1070), .QN(n9571) );
  SDFFX1 DFF_278_Q_reg ( .D(g26899), .SI(g1070), .SE(n10186), .CLK(n10538), 
        .Q(g822), .QN(n5422) );
  SDFFX1 DFF_279_Q_reg ( .D(g14673), .SI(g822), .SE(n10251), .CLK(n10603), .Q(
        g17715) );
  SDFFX1 DFF_280_Q_reg ( .D(g30336), .SI(g17715), .SE(n10197), .CLK(n10549), 
        .Q(g914), .QN(n5560) );
  SDFFX1 DFF_281_Q_reg ( .D(g17639), .SI(g914), .SE(n10216), .CLK(n10568), .Q(
        g5339) );
  SDFFX1 DFF_282_Q_reg ( .D(g26940), .SI(g5339), .SE(n10216), .CLK(n10568), 
        .Q(g4164), .QN(n10073) );
  SDFFX1 DFF_283_Q_reg ( .D(g25622), .SI(g4164), .SE(n10191), .CLK(n10543), 
        .Q(test_so20), .QN(n10152) );
  SDFFX1 DFF_284_Q_reg ( .D(g34447), .SI(test_si21), .SE(n10219), .CLK(n10571), 
        .Q(g2807), .QN(n5379) );
  SDFFX1 DFF_286_Q_reg ( .D(g33613), .SI(g2807), .SE(n10261), .CLK(n10613), 
        .Q(g4054), .QN(n5395) );
  SDFFX1 DFF_287_Q_reg ( .D(g25749), .SI(g4054), .SE(n10180), .CLK(n10532), 
        .Q(g6191), .QN(n5888) );
  SDFFX1 DFF_288_Q_reg ( .D(g25704), .SI(g6191), .SE(n10180), .CLK(n10532), 
        .Q(g5077), .QN(n5455) );
  SDFFX1 DFF_289_Q_reg ( .D(g33053), .SI(g5077), .SE(n10180), .CLK(n10532), 
        .Q(g5523), .QN(n5647) );
  SDFFX1 DFF_290_Q_reg ( .D(g16722), .SI(g5523), .SE(n10250), .CLK(n10602), 
        .Q(g3680) );
  SDFFX1 DFF_291_Q_reg ( .D(g30555), .SI(g3680), .SE(n10194), .CLK(n10546), 
        .Q(g6637), .QN(n9858) );
  SDFFX1 DFF_292_Q_reg ( .D(g25601), .SI(g6637), .SE(n10254), .CLK(n10606), 
        .Q(g174), .QN(n5402) );
  SDFFX1 DFF_293_Q_reg ( .D(g33971), .SI(g174), .SE(n10166), .CLK(n10518), .Q(
        g1682), .QN(n9697) );
  SDFFX1 DFF_294_Q_reg ( .D(g26892), .SI(g1682), .SE(n10239), .CLK(n10591), 
        .Q(g355) );
  SDFFX1 DFF_295_Q_reg ( .D(g17400), .SI(g355), .SE(n10240), .CLK(n10592), .Q(
        g1087), .QN(n10069) );
  SDFFX1 DFF_296_Q_reg ( .D(g26915), .SI(g1087), .SE(n10198), .CLK(n10550), 
        .Q(g1105), .QN(n5478) );
  SDFFX1 DFF_297_Q_reg ( .D(g33008), .SI(g1105), .SE(n10208), .CLK(n10560), 
        .Q(test_so21), .QN(n10126) );
  SDFFX1 DFF_298_Q_reg ( .D(g30538), .SI(test_si22), .SE(n10226), .CLK(n10578), 
        .Q(g6307), .QN(n9863) );
  SDFFX1 DFF_299_Q_reg ( .D(g8344), .SI(g6307), .SE(n10262), .CLK(n10614), .Q(
        g3802) );
  SDFFX1 DFF_300_Q_reg ( .D(g25750), .SI(g3802), .SE(n10262), .CLK(n10614), 
        .Q(g6159) );
  SDFFX1 DFF_301_Q_reg ( .D(g30369), .SI(g6159), .SE(n10192), .CLK(n10544), 
        .Q(g2255), .QN(n5414) );
  SDFFX1 DFF_302_Q_reg ( .D(g34446), .SI(g2255), .SE(n10215), .CLK(n10567), 
        .Q(g2815), .QN(n5404) );
  SDFFX1 DFF_303_Q_reg ( .D(g29230), .SI(g2815), .SE(n10197), .CLK(n10549), 
        .Q(g911), .QN(n5559) );
  SDFFX1 DFF_304_Q_reg ( .D(n10105), .SI(g911), .SE(n10235), .CLK(n10587), .Q(
        g43) );
  SDFFX1 DFF_305_Q_reg ( .D(g13966), .SI(g43), .SE(n10235), .CLK(n10587), .Q(
        g16775), .QN(n9888) );
  SDFFX1 DFF_306_Q_reg ( .D(g33975), .SI(g16775), .SE(n10266), .CLK(n10618), 
        .Q(g1748) );
  SDFFX1 DFF_307_Q_reg ( .D(g30497), .SI(g1748), .SE(n10180), .CLK(n10532), 
        .Q(g5551), .QN(n9957) );
  SDFFX1 DFF_309_Q_reg ( .D(g30418), .SI(g5551), .SE(n10270), .CLK(n10622), 
        .Q(g3558), .QN(n9937) );
  SDFFX1 DFF_310_Q_reg ( .D(g25721), .SI(g3558), .SE(n10182), .CLK(n10534), 
        .Q(g5499), .QN(n5885) );
  SDFFX1 DFF_311_Q_reg ( .D(g34622), .SI(g5499), .SE(n10182), .CLK(n10534), 
        .Q(test_so22) );
  SDFFX1 DFF_312_Q_reg ( .D(g30438), .SI(test_si23), .SE(n10183), .CLK(n10535), 
        .Q(g3901), .QN(n10021) );
  SDFFX1 DFF_313_Q_reg ( .D(g34266), .SI(g3901), .SE(n10196), .CLK(n10548), 
        .Q(g4888), .QN(n5863) );
  SDFFX1 DFF_314_Q_reg ( .D(g30540), .SI(g4888), .SE(n10226), .CLK(n10578), 
        .Q(g6251), .QN(n10006) );
  SDFFX1 DFF_315_Q_reg ( .D(g17760), .SI(g6251), .SE(n10226), .CLK(n10578), 
        .Q(g17649), .QN(n9879) );
  SDFFX1 DFF_316_Q_reg ( .D(g32986), .SI(g17649), .SE(n10270), .CLK(n10622), 
        .Q(g1373), .QN(n9762) );
  SDFFX1 DFF_317_Q_reg ( .D(g25648), .SI(g1373), .SE(n10170), .CLK(n10522), 
        .Q(g8215), .QN(n5723) );
  SDFFX1 DFF_318_Q_reg ( .D(g33960), .SI(g8215), .SE(n10210), .CLK(n10562), 
        .Q(g157), .QN(n5678) );
  SDFFX1 DFF_319_Q_reg ( .D(g34442), .SI(g157), .SE(n10257), .CLK(n10609), .Q(
        g2783), .QN(n5403) );
  SDFFX1 DFF_320_Q_reg ( .D(g8839), .SI(g2783), .SE(n10230), .CLK(n10582), .Q(
        g4281), .QN(n10102) );
  SDFFX1 DFF_321_Q_reg ( .D(g30421), .SI(g4281), .SE(n10184), .CLK(n10536), 
        .Q(g3574), .QN(n9936) );
  SDFFX1 DFF_322_Q_reg ( .D(g33573), .SI(g3574), .SE(n10269), .CLK(n10621), 
        .Q(g2112), .QN(n5848) );
  SDFFX1 DFF_323_Q_reg ( .D(g34730), .SI(g2112), .SE(n10269), .CLK(n10621), 
        .Q(g1283), .QN(n5635) );
  SDFFX1 DFF_324_Q_reg ( .D(g24205), .SI(g1283), .SE(n10203), .CLK(n10555), 
        .Q(test_so23) );
  SDFFX1 DFF_325_Q_reg ( .D(g10122_Tj), .SI(test_si24), .SE(n10185), .CLK(
        n10537), .Q(g4297) );
  SDFFX1 DFF_326_Q_reg ( .D(g12350), .SI(g4297), .SE(n10185), .CLK(n10537), 
        .Q(g14738), .QN(n5698) );
  SDFFX1 DFF_327_Q_reg ( .D(g19357), .SI(g14738), .SE(n10212), .CLK(n10564), 
        .Q(g13272), .QN(n9745) );
  SDFFX1 DFF_328_Q_reg ( .D(g32979), .SI(g13272), .SE(n10191), .CLK(n10543), 
        .Q(g758), .QN(n5331) );
  SDFFX1 DFF_331_Q_reg ( .D(n291), .SI(g758), .SE(n10224), .CLK(n10576), .Q(
        g4639), .QN(n5727) );
  SDFFX1 DFF_332_Q_reg ( .D(g25763), .SI(g4639), .SE(n10270), .CLK(n10622), 
        .Q(g6537), .QN(n5884) );
  SDFFX1 DFF_333_Q_reg ( .D(g30481), .SI(g6537), .SE(n10180), .CLK(n10532), 
        .Q(g5543), .QN(n9958) );
  SDFFX1 DFF_334_Q_reg ( .D(g7946), .SI(g5543), .SE(n10227), .CLK(n10579), .Q(
        g8475), .QN(n9651) );
  SDFFX1 DFF_336_Q_reg ( .D(g30517), .SI(g8475), .SE(n10187), .CLK(n10539), 
        .Q(g5961), .QN(n9848) );
  SDFFX1 DFF_337_Q_reg ( .D(g30539), .SI(g5961), .SE(n10266), .CLK(n10618), 
        .Q(g6243), .QN(n9964) );
  SDFFX1 DFF_338_Q_reg ( .D(g34880), .SI(g6243), .SE(n10223), .CLK(n10575), 
        .Q(n9340), .QN(n18472) );
  SDFFX1 DFF_339_Q_reg ( .D(g24242), .SI(n9340), .SE(n10223), .CLK(n10575), 
        .Q(g12919), .QN(n5654) );
  SDFFX1 DFF_340_Q_reg ( .D(g30436), .SI(g12919), .SE(n10214), .CLK(n10566), 
        .Q(test_so24) );
  SDFFX1 DFF_341_Q_reg ( .D(g29265), .SI(test_si25), .SE(n10173), .CLK(n10525), 
        .Q(g3476), .QN(n5786) );
  SDFFX1 DFF_342_Q_reg ( .D(g32990), .SI(g3476), .SE(n10202), .CLK(n10554), 
        .Q(g1664), .QN(n5407) );
  SDFFX1 DFF_343_Q_reg ( .D(g24245), .SI(g1664), .SE(n10224), .CLK(n10576), 
        .Q(g1246), .QN(n5756) );
  SDFFX1 DFF_345_Q_reg ( .D(g30553), .SI(g1246), .SE(n10193), .CLK(n10545), 
        .Q(g6629), .QN(n9891) );
  SDFFX1 DFF_346_Q_reg ( .D(g26907), .SI(g6629), .SE(n10171), .CLK(n10523), 
        .Q(g246), .QN(n6008) );
  SDFFX1 DFF_347_Q_reg ( .D(g24278), .SI(g246), .SE(n10200), .CLK(n10552), .Q(
        g4049), .QN(n9905) );
  SDFFX1 DFF_348_Q_reg ( .D(g26955), .SI(g4049), .SE(n10188), .CLK(n10540), 
        .Q(g7260) );
  SDFFX1 DFF_349_Q_reg ( .D(g24282), .SI(g7260), .SE(n10188), .CLK(n10540), 
        .Q(g2932), .QN(n10091) );
  SDFFX1 DFF_350_Q_reg ( .D(g29276), .SI(g2932), .SE(n10188), .CLK(n10540), 
        .Q(g4575) );
  SDFFX1 DFF_351_Q_reg ( .D(g31894), .SI(g4575), .SE(n10240), .CLK(n10592), 
        .Q(g4098), .QN(n5350) );
  SDFFX1 DFF_352_Q_reg ( .D(g33037), .SI(g4098), .SE(n10244), .CLK(n10596), 
        .Q(g4498) );
  SDFFX1 DFF_353_Q_reg ( .D(g26894), .SI(g4498), .SE(n10245), .CLK(n10597), 
        .Q(g528), .QN(n5327) );
  SDFFX1 DFF_355_Q_reg ( .D(g34977), .SI(g528), .SE(n10175), .CLK(n10527), .Q(
        test_so25), .QN(n5477) );
  SDFFX1 DFF_356_Q_reg ( .D(g25654), .SI(test_si26), .SE(n10190), .CLK(n10542), 
        .Q(g3139), .QN(n5447) );
  SDFFX1 DFF_357_Q_reg ( .D(g33962), .SI(g3139), .SE(n10190), .CLK(n10542), 
        .Q(g29215) );
  SDFFX1 DFF_358_Q_reg ( .D(g34451), .SI(g29215), .SE(n10264), .CLK(n10616), 
        .Q(g4584), .QN(n5539) );
  SDFFX1 DFF_359_Q_reg ( .D(g34250), .SI(g4584), .SE(n10264), .CLK(n10616), 
        .Q(g142), .QN(n5724) );
  SDFFX1 DFF_360_Q_reg ( .D(g14597), .SI(g142), .SE(n10216), .CLK(n10568), .Q(
        g17639) );
  SDFFX1 DFF_361_Q_reg ( .D(g29295), .SI(g17639), .SE(n10181), .CLK(n10533), 
        .Q(g5831) );
  SDFFX1 DFF_362_Q_reg ( .D(g26905), .SI(g5831), .SE(n10248), .CLK(n10600), 
        .Q(g239), .QN(n9909) );
  SDFFX1 DFF_363_Q_reg ( .D(g25629), .SI(g239), .SE(n10228), .CLK(n10580), .Q(
        g1216), .QN(n5442) );
  SDFFX1 DFF_364_Q_reg ( .D(g34792), .SI(g1216), .SE(n10166), .CLK(n10518), 
        .Q(g2848), .QN(n9709) );
  SDFFX1 DFF_366_Q_reg ( .D(g25703), .SI(g2848), .SE(n10202), .CLK(n10554), 
        .Q(g5022), .QN(n9784) );
  SDFFX1 DFF_367_Q_reg ( .D(g14518), .SI(g5022), .SE(n10241), .CLK(n10593), 
        .Q(g16955) );
  SDFFX1 DFF_368_Q_reg ( .D(g32983), .SI(g16955), .SE(n10250), .CLK(n10602), 
        .Q(g1030), .QN(n9764) );
  SDFFX1 DFF_369_Q_reg ( .D(g16924), .SI(g1030), .SE(n10250), .CLK(n10602), 
        .Q(test_so26) );
  SDFFX1 DFF_370_Q_reg ( .D(g30402), .SI(test_si27), .SE(n10257), .CLK(n10609), 
        .Q(g3231), .QN(n9942) );
  SDFFX1 DFF_371_Q_reg ( .D(g25757), .SI(g3231), .SE(n10257), .CLK(n10609), 
        .Q(g9817) );
  SDFFX1 DFF_372_Q_reg ( .D(g17423), .SI(g9817), .SE(n10257), .CLK(n10609), 
        .Q(g1430), .QN(n10067) );
  SDFFX1 DFF_373_Q_reg ( .D(g7245), .SI(g1430), .SE(n10257), .CLK(n10609), .Q(
        n9336), .QN(n18479) );
  SDFFX1 DFF_374_Q_reg ( .D(g33999), .SI(n9336), .SE(n10192), .CLK(n10544), 
        .Q(g2241), .QN(n9696) );
  SDFFX1 DFF_375_Q_reg ( .D(g24262), .SI(g2241), .SE(n10258), .CLK(n10610), 
        .Q(g1564), .QN(n10066) );
  SDFFX1 DFF_376_Q_reg ( .D(g25729), .SI(g1564), .SE(n10266), .CLK(n10618), 
        .Q(g9680) );
  SDFFX1 DFF_377_Q_reg ( .D(test_so92), .SI(g9680), .SE(n10267), .CLK(n10619), 
        .Q(g6148) );
  SDFFX1 DFF_378_Q_reg ( .D(g30558), .SI(g6148), .SE(n10194), .CLK(n10546), 
        .Q(g6649), .QN(n9994) );
  SDFFX1 DFF_379_Q_reg ( .D(g34781), .SI(g6649), .SE(n10208), .CLK(n10560), 
        .Q(g110), .QN(n9568) );
  SDFFX1 DFF_380_Q_reg ( .D(g14125), .SI(g110), .SE(n10247), .CLK(n10599), .Q(
        g14147), .QN(n9597) );
  SDFFX1 DFF_382_Q_reg ( .D(g26901), .SI(g14147), .SE(n10247), .CLK(n10599), 
        .Q(g225), .QN(n5597) );
  SDFFX1 DFF_383_Q_reg ( .D(g26961), .SI(g225), .SE(n10248), .CLK(n10600), .Q(
        test_so27) );
  SDFFX1 DFF_384_Q_reg ( .D(g33039), .SI(test_si28), .SE(n10244), .CLK(n10596), 
        .Q(g4504) );
  SDFFX1 DFF_385_Q_reg ( .D(g33059), .SI(g4504), .SE(n10245), .CLK(n10597), 
        .Q(g5873), .QN(n5388) );
  SDFFX1 DFF_386_Q_reg ( .D(g31899), .SI(g5873), .SE(n10208), .CLK(n10560), 
        .Q(g5037), .QN(n5611) );
  SDFFX1 DFF_387_Q_reg ( .D(g33007), .SI(g5037), .SE(n10208), .CLK(n10560), 
        .Q(g2319), .QN(n5375) );
  SDFFX1 DFF_388_Q_reg ( .D(g25720), .SI(g2319), .SE(n10182), .CLK(n10534), 
        .Q(g5495), .QN(n5446) );
  SDFFX1 DFF_389_Q_reg ( .D(g21891), .SI(g5495), .SE(n10216), .CLK(n10568), 
        .Q(g11770) );
  SDFFX1 DFF_390_Q_reg ( .D(g30462), .SI(g11770), .SE(n10216), .CLK(n10568), 
        .Q(g5208), .QN(n9916) );
  SDFFX1 DFF_392_Q_reg ( .D(g30487), .SI(g5208), .SE(n10175), .CLK(n10527), 
        .Q(g5579), .QN(n9927) );
  SDFFX1 DFF_393_Q_reg ( .D(g33058), .SI(g5579), .SE(n10244), .CLK(n10596), 
        .Q(g5869), .QN(n5649) );
  SDFFX1 DFF_395_Q_reg ( .D(g24261), .SI(g5869), .SE(n10266), .CLK(n10618), 
        .Q(g1589), .QN(n5755) );
  SDFFX1 DFF_396_Q_reg ( .D(g25730), .SI(g1589), .SE(n10266), .CLK(n10618), 
        .Q(g5752) );
  SDFFX1 DFF_397_Q_reg ( .D(g30531), .SI(g5752), .SE(n10266), .CLK(n10618), 
        .Q(g6279), .QN(n9949) );
  SDFFX1 DFF_398_Q_reg ( .D(g30506), .SI(g6279), .SE(n10266), .CLK(n10618), 
        .Q(test_so28) );
  SDFFX1 DFF_399_Q_reg ( .D(g34804), .SI(test_si29), .SE(n10165), .CLK(n10517), 
        .Q(g2975), .QN(n5750) );
  SDFFX1 DFF_400_Q_reg ( .D(g25747), .SI(g2975), .SE(n10179), .CLK(n10531), 
        .Q(g6167), .QN(n5430) );
  SDFFX1 DFF_401_Q_reg ( .D(g11418), .SI(g6167), .SE(n10255), .CLK(n10607), 
        .Q(g13966), .QN(n5701) );
  SDFFX1 DFF_402_Q_reg ( .D(g33601), .SI(g13966), .SE(n10212), .CLK(n10564), 
        .Q(g2599), .QN(n5524) );
  SDFFX1 DFF_403_Q_reg ( .D(g26922), .SI(g2599), .SE(n10176), .CLK(n10528), 
        .Q(g1448), .QN(n5343) );
  SDFFX1 DFF_404_Q_reg ( .D(g14096), .SI(g1448), .SE(n10247), .CLK(n10599), 
        .Q(g14125), .QN(n9596) );
  SDFFX1 DFF_406_Q_reg ( .D(g29250), .SI(g14125), .SE(n10195), .CLK(n10547), 
        .Q(g2370), .QN(n9826) );
  SDFFX1 DFF_407_Q_reg ( .D(g30459), .SI(g2370), .SE(n10250), .CLK(n10602), 
        .Q(g5164), .QN(n5570) );
  SDFFX1 DFF_408_Q_reg ( .D(g8475), .SI(g5164), .SE(n10250), .CLK(n10602), .Q(
        g1333), .QN(n5616) );
  SDFFX1 DFF_409_Q_reg ( .D(g33534), .SI(g1333), .SE(n10209), .CLK(n10561), 
        .Q(g153), .QN(n5677) );
  SDFFX1 DFF_410_Q_reg ( .D(g30543), .SI(g153), .SE(n10238), .CLK(n10590), .Q(
        g6549), .QN(n5571) );
  SDFFX1 DFF_411_Q_reg ( .D(g29275), .SI(g6549), .SE(n10238), .CLK(n10590), 
        .Q(g4087), .QN(n5480) );
  SDFFX1 DFF_412_Q_reg ( .D(g34030), .SI(g4087), .SE(n10259), .CLK(n10611), 
        .Q(test_so29), .QN(n10125) );
  SDFFX1 DFF_413_Q_reg ( .D(g34980), .SI(test_si30), .SE(n10198), .CLK(n10550), 
        .Q(g2984), .QN(n5842) );
  SDFFX1 DFF_414_Q_reg ( .D(g30451), .SI(g2984), .SE(n10241), .CLK(n10593), 
        .Q(g3961) );
  SDFFX1 DFF_416_Q_reg ( .D(g25627), .SI(g3961), .SE(n10268), .CLK(n10620), 
        .Q(g962), .QN(n5630) );
  SDFFX1 DFF_417_Q_reg ( .D(g34657), .SI(g962), .SE(n10179), .CLK(n10531), .Q(
        g101), .QN(n18465) );
  SDFFX1 DFF_418_Q_reg ( .D(g8870), .SI(g101), .SE(n10179), .CLK(n10531), .Q(
        g8918) );
  SDFFX1 DFF_419_Q_reg ( .D(g30552), .SI(g8918), .SE(n10249), .CLK(n10601), 
        .Q(g6625), .QN(n9947) );
  SDFFX1 DFF_420_Q_reg ( .D(g34979), .SI(g6625), .SE(n10191), .CLK(n10543), 
        .Q(n9332) );
  SDFFX1 DFF_421_Q_reg ( .D(g30337), .SI(n9332), .SE(n10191), .CLK(n10543), 
        .Q(g1018), .QN(n9763) );
  SDFFX1 DFF_422_Q_reg ( .D(g24254), .SI(g1018), .SE(n10192), .CLK(n10544), 
        .Q(g17320), .QN(n9737) );
  SDFFX1 DFF_423_Q_reg ( .D(g24277), .SI(g17320), .SE(n10200), .CLK(n10552), 
        .Q(g4045), .QN(n9906) );
  SDFFX1 DFF_424_Q_reg ( .D(g29237), .SI(g4045), .SE(n10200), .CLK(n10552), 
        .Q(g1467), .QN(n5693) );
  SDFFX1 DFF_425_Q_reg ( .D(g30378), .SI(g1467), .SE(n10215), .CLK(n10567), 
        .Q(g2461), .QN(n5840) );
  SDFFX1 DFF_428_Q_reg ( .D(g33019), .SI(g2461), .SE(n10257), .CLK(n10609), 
        .Q(test_so30), .QN(n5300) );
  SDFFX1 DFF_429_Q_reg ( .D(g33623), .SI(test_si31), .SE(n10181), .CLK(n10533), 
        .Q(g5990), .QN(n5589) );
  SDFFX1 DFF_431_Q_reg ( .D(g29235), .SI(g5990), .SE(n10211), .CLK(n10563), 
        .Q(g1256), .QN(n5558) );
  SDFFX1 DFF_432_Q_reg ( .D(g31902), .SI(g1256), .SE(n10202), .CLK(n10554), 
        .Q(g5029), .QN(n5601) );
  SDFFX1 DFF_433_Q_reg ( .D(g29306), .SI(g5029), .SE(n10189), .CLK(n10541), 
        .Q(g6519), .QN(n5806) );
  SDFFX1 DFF_434_Q_reg ( .D(g25689), .SI(g6519), .SE(n10189), .CLK(n10541), 
        .Q(g4169), .QN(n5729) );
  SDFFX1 DFF_435_Q_reg ( .D(g33978), .SI(g4169), .SE(n10267), .CLK(n10619), 
        .Q(g1816), .QN(n9615) );
  SDFFX1 DFF_436_Q_reg ( .D(g26970), .SI(g1816), .SE(n10267), .CLK(n10619), 
        .Q(g4369), .QN(n9911) );
  SDFFX1 DFF_439_Q_reg ( .D(g29278), .SI(g4369), .SE(n10194), .CLK(n10546), 
        .Q(g4578) );
  SDFFX1 DFF_440_Q_reg ( .D(g34253), .SI(g4578), .SE(n10195), .CLK(n10547), 
        .Q(g4459), .QN(n5765) );
  SDFFX1 DFF_441_Q_reg ( .D(g29272), .SI(g4459), .SE(n10167), .CLK(n10519), 
        .Q(g3831), .QN(n5872) );
  SDFFX1 DFF_442_Q_reg ( .D(g33595), .SI(g3831), .SE(n10269), .CLK(n10621), 
        .Q(g2514), .QN(n9657) );
  SDFFX1 DFF_443_Q_reg ( .D(g33610), .SI(g2514), .SE(n10205), .CLK(n10557), 
        .Q(g3288), .QN(n5400) );
  SDFFX1 DFF_444_Q_reg ( .D(g33589), .SI(g3288), .SE(n10176), .CLK(n10528), 
        .Q(test_so31), .QN(n10153) );
  SDFFX1 DFF_445_Q_reg ( .D(g34605), .SI(test_si32), .SE(n10221), .CLK(n10573), 
        .Q(g2145), .QN(n5307) );
  SDFFX1 DFF_446_Q_reg ( .D(g30350), .SI(g2145), .SE(n10221), .CLK(n10573), 
        .Q(g1700), .QN(n5417) );
  SDFFX1 DFF_447_Q_reg ( .D(g25611), .SI(g1700), .SE(n10245), .CLK(n10597), 
        .Q(g513), .QN(n5548) );
  SDFFX1 DFF_448_Q_reg ( .D(test_so9), .SI(g513), .SE(n10256), .CLK(n10608), 
        .Q(g2841), .QN(n5963) );
  SDFFX1 DFF_449_Q_reg ( .D(g33619), .SI(g2841), .SE(n10262), .CLK(n10614), 
        .Q(g5297), .QN(n5588) );
  SDFFX1 DFF_451_Q_reg ( .D(g34022), .SI(g5297), .SE(n10259), .CLK(n10611), 
        .Q(g2763), .QN(n9587) );
  SDFFX1 DFF_452_Q_reg ( .D(g34033), .SI(g2763), .SE(n10259), .CLK(n10611), 
        .Q(g4793), .QN(n5368) );
  SDFFX1 DFF_453_Q_reg ( .D(g34726), .SI(g4793), .SE(n10268), .CLK(n10620), 
        .Q(g952), .QN(n9577) );
  SDFFX1 DFF_454_Q_reg ( .D(g31870), .SI(g952), .SE(n10211), .CLK(n10563), .Q(
        g1263), .QN(n5674) );
  SDFFX1 DFF_455_Q_reg ( .D(g33985), .SI(g1263), .SE(n10198), .CLK(n10550), 
        .Q(g1950), .QN(n9695) );
  SDFFX1 DFF_456_Q_reg ( .D(g29283), .SI(g1950), .SE(n10178), .CLK(n10530), 
        .Q(g5138), .QN(n5871) );
  SDFFX1 DFF_457_Q_reg ( .D(g34003), .SI(g5138), .SE(n10263), .CLK(n10615), 
        .Q(g2307) );
  SDFFX1 DFF_458_Q_reg ( .D(g9497), .SI(g2307), .SE(n10263), .CLK(n10615), .Q(
        test_so32) );
  SDFFX1 DFF_460_Q_reg ( .D(g25677), .SI(test_si33), .SE(n10181), .CLK(n10533), 
        .Q(g8398) );
  SDFFX1 DFF_461_Q_reg ( .D(g34463), .SI(g8398), .SE(n10181), .CLK(n10533), 
        .Q(g4664) );
  SDFFX1 DFF_462_Q_reg ( .D(g33006), .SI(g4664), .SE(n10209), .CLK(n10561), 
        .Q(g2223), .QN(n5406) );
  SDFFX1 DFF_463_Q_reg ( .D(g29292), .SI(g2223), .SE(n10181), .CLK(n10533), 
        .Q(g5808), .QN(n5749) );
  SDFFX1 DFF_464_Q_reg ( .D(g30557), .SI(g5808), .SE(n10193), .CLK(n10545), 
        .Q(g6645), .QN(n9877) );
  SDFFX1 DFF_465_Q_reg ( .D(g33989), .SI(g6645), .SE(n10214), .CLK(n10566), 
        .Q(g2016) );
  SDFFX1 DFF_467_Q_reg ( .D(g33033), .SI(g2016), .SE(n10214), .CLK(n10566), 
        .Q(g3873), .QN(n5387) );
  SDFFX1 DFF_468_Q_reg ( .D(g11388), .SI(g3873), .SE(n10221), .CLK(n10573), 
        .Q(g13926), .QN(n5699) );
  SDFFX1 DFF_469_Q_reg ( .D(g34005), .SI(g13926), .SE(n10263), .CLK(n10615), 
        .Q(g2315), .QN(n5802) );
  SDFFX1 DFF_470_Q_reg ( .D(g26932), .SI(g2315), .SE(n10219), .CLK(n10571), 
        .Q(g2811), .QN(n9608) );
  SDFFX1 DFF_471_Q_reg ( .D(g30516), .SI(g2811), .SE(n10187), .CLK(n10539), 
        .Q(g5957), .QN(n9980) );
  SDFFX1 DFF_472_Q_reg ( .D(g33575), .SI(g5957), .SE(n10217), .CLK(n10569), 
        .Q(g2047), .QN(n5831) );
  SDFFX1 DFF_473_Q_reg ( .D(g33032), .SI(g2047), .SE(n10240), .CLK(n10592), 
        .Q(test_so33) );
  SDFFX1 DFF_474_Q_reg ( .D(g14779), .SI(test_si34), .SE(n10220), .CLK(n10572), 
        .Q(g17760), .QN(n9894) );
  SDFFX1 DFF_476_Q_reg ( .D(g30486), .SI(g17760), .SE(n10180), .CLK(n10532), 
        .Q(g5575), .QN(n9838) );
  SDFFX1 DFF_477_Q_reg ( .D(g34974), .SI(g5575), .SE(n10180), .CLK(n10532), 
        .Q(n9327) );
  SDFFX1 DFF_478_Q_reg ( .D(g25678), .SI(n9327), .SE(n10181), .CLK(n10533), 
        .Q(g3752) );
  SDFFX1 DFF_479_Q_reg ( .D(g30440), .SI(g3752), .SE(n10214), .CLK(n10566), 
        .Q(g3917), .QN(n9817) );
  SDFFX1 DFF_480_Q_reg ( .D(test_so86), .SI(g3917), .SE(n10206), .CLK(n10558), 
        .Q(g8783), .QN(DFF_480_n1) );
  SDFFX1 DFF_481_Q_reg ( .D(g12923), .SI(g8783), .SE(n10206), .CLK(n10558), 
        .Q(g1585), .QN(n5757) );
  SDFFX1 DFF_482_Q_reg ( .D(g26949), .SI(g1585), .SE(n10255), .CLK(n10607), 
        .Q(g4388), .QN(n9676) );
  SDFFX1 DFF_483_Q_reg ( .D(g30530), .SI(g4388), .SE(n10225), .CLK(n10577), 
        .Q(g6275), .QN(n9865) );
  SDFFX1 DFF_484_Q_reg ( .D(g30542), .SI(g6275), .SE(n10226), .CLK(n10578), 
        .Q(g6311), .QN(n9806) );
  SDFFX1 DFF_485_Q_reg ( .D(g8915), .SI(g6311), .SE(n10226), .CLK(n10578), .Q(
        g8916), .QN(n18469) );
  SDFFX1 DFF_486_Q_reg ( .D(g25624), .SI(g8916), .SE(n10253), .CLK(n10605), 
        .Q(g1041), .QN(n9591) );
  SDFFX1 DFF_487_Q_reg ( .D(g30383), .SI(g1041), .SE(n10213), .CLK(n10565), 
        .Q(test_so34) );
  SDFFX1 DFF_488_Q_reg ( .D(g33597), .SI(test_si35), .SE(n10207), .CLK(n10559), 
        .Q(g2537), .QN(n5411) );
  SDFFX1 DFF_489_Q_reg ( .D(g34598), .SI(g2537), .SE(n10172), .CLK(n10524), 
        .Q(g29221), .QN(g23612) );
  SDFFX1 DFF_490_Q_reg ( .D(g26957), .SI(g29221), .SE(n10172), .CLK(n10524), 
        .Q(g4430), .QN(n9679) );
  SDFFX1 DFF_491_Q_reg ( .D(g26967), .SI(g4430), .SE(n10263), .CLK(n10615), 
        .Q(n9325), .QN(n18467) );
  SDFFX1 DFF_493_Q_reg ( .D(g28102), .SI(n9325), .SE(n10226), .CLK(n10578), 
        .Q(g4826) );
  SDFFX1 DFF_494_Q_reg ( .D(g30524), .SI(g4826), .SE(n10226), .CLK(n10578), 
        .Q(g6239), .QN(n9809) );
  SDFFX1 DFF_496_Q_reg ( .D(g26903), .SI(g6239), .SE(n10248), .CLK(n10600), 
        .Q(g232), .QN(n9908) );
  SDFFX1 DFF_497_Q_reg ( .D(g30475), .SI(g232), .SE(n10217), .CLK(n10569), .Q(
        g5268), .QN(n9845) );
  SDFFX1 DFF_498_Q_reg ( .D(g34647), .SI(g5268), .SE(n10217), .CLK(n10569), 
        .Q(g6545), .QN(n5497) );
  SDFFX1 DFF_499_Q_reg ( .D(g30377), .SI(g6545), .SE(n10177), .CLK(n10529), 
        .Q(n9324), .QN(n18483) );
  SDFFX1 DFF_500_Q_reg ( .D(g33553), .SI(n9324), .SE(n10177), .CLK(n10529), 
        .Q(g1772), .QN(n5504) );
  SDFFX1 DFF_502_Q_reg ( .D(g31903), .SI(g1772), .SE(n10202), .CLK(n10554), 
        .Q(g5052), .QN(n5607) );
  SDFFX1 DFF_503_Q_reg ( .D(g25715), .SI(g5052), .SE(n10203), .CLK(n10555), 
        .Q(test_so35) );
  SDFFX1 DFF_504_Q_reg ( .D(g33984), .SI(test_si36), .SE(n10203), .CLK(n10555), 
        .Q(g1890), .QN(n5799) );
  SDFFX1 DFF_505_Q_reg ( .D(g33602), .SI(g1890), .SE(n10249), .CLK(n10601), 
        .Q(g2629), .QN(n5521) );
  SDFFX1 DFF_506_Q_reg ( .D(g28045), .SI(g2629), .SE(n10221), .CLK(n10573), 
        .Q(g572), .QN(n5337) );
  SDFFX1 DFF_507_Q_reg ( .D(g34603), .SI(g572), .SE(n10221), .CLK(n10573), .Q(
        g2130), .QN(n5487) );
  SDFFX1 DFF_508_Q_reg ( .D(g33035), .SI(g2130), .SE(n10240), .CLK(n10592), 
        .Q(g4108) );
  SDFFX1 DFF_509_Q_reg ( .D(g9251), .SI(g4108), .SE(n10240), .CLK(n10592), .Q(
        g4308) );
  SDFFX1 DFF_510_Q_reg ( .D(g24208), .SI(g4308), .SE(n10171), .CLK(n10523), 
        .Q(g475), .QN(n9611) );
  SDFFX1 DFF_511_Q_reg ( .D(g8416), .SI(g475), .SE(n10234), .CLK(n10586), .Q(
        g990), .QN(n5622) );
  SDFFX1 DFF_512_Q_reg ( .D(g34971), .SI(g990), .SE(n10197), .CLK(n10549), .Q(
        g31), .QN(n5469) );
  SDFFX1 DFF_514_Q_reg ( .D(g34970), .SI(g31), .SE(n10190), .CLK(n10542), .Q(
        n9322) );
  SDFFX1 DFF_515_Q_reg ( .D(g24213), .SI(n9322), .SE(n10191), .CLK(n10543), 
        .Q(g12184) );
  SDFFX1 DFF_517_Q_reg ( .D(g33614), .SI(g12184), .SE(n10168), .CLK(n10520), 
        .Q(g3990), .QN(n5594) );
  SDFFX1 DFF_519_Q_reg ( .D(g33060), .SI(g3990), .SE(n10244), .CLK(n10596), 
        .Q(test_so36), .QN(n10139) );
  SDFFX1 DFF_520_Q_reg ( .D(g30362), .SI(test_si37), .SE(n10169), .CLK(n10521), 
        .Q(g1992), .QN(n5890) );
  SDFFX1 DFF_522_Q_reg ( .D(g33023), .SI(g1992), .SE(n10169), .CLK(n10521), 
        .Q(g3171), .QN(n5603) );
  SDFFX1 DFF_524_Q_reg ( .D(g26898), .SI(g3171), .SE(n10186), .CLK(n10538), 
        .Q(g812), .QN(n5733) );
  SDFFX1 DFF_525_Q_reg ( .D(g25618), .SI(g812), .SE(n10186), .CLK(n10538), .Q(
        g832), .QN(n10065) );
  SDFFX1 DFF_526_Q_reg ( .D(g30518), .SI(g832), .SE(n10186), .CLK(n10538), .Q(
        g5897), .QN(n9955) );
  SDFFX1 DFF_527_Q_reg ( .D(g25688), .SI(g5897), .SE(n10186), .CLK(n10538), 
        .Q(g25689), .QN(n9621) );
  SDFFX1 DFF_528_Q_reg ( .D(g4570), .SI(g25689), .SE(n10243), .CLK(n10595), 
        .Q(g4571) );
  SDFFX1 DFF_529_Q_reg ( .D(g11349), .SI(g4571), .SE(n10243), .CLK(n10595), 
        .Q(g13895), .QN(n5702) );
  SDFFX1 DFF_530_Q_reg ( .D(g26959), .SI(g13895), .SE(n10252), .CLK(n10604), 
        .Q(g4455) );
  SDFFX1 DFF_531_Q_reg ( .D(g34801), .SI(g4455), .SE(n10182), .CLK(n10534), 
        .Q(g2902), .QN(n9731) );
  SDFFX1 DFF_532_Q_reg ( .D(g26884), .SI(g2902), .SE(n10209), .CLK(n10561), 
        .Q(g333) );
  SDFFX1 DFF_533_Q_reg ( .D(g25600), .SI(g333), .SE(n10254), .CLK(n10606), .Q(
        g168) );
  SDFFX1 DFF_534_Q_reg ( .D(g26933), .SI(g168), .SE(n10215), .CLK(n10567), .Q(
        test_so37), .QN(n10149) );
  SDFFX1 DFF_535_Q_reg ( .D(g28066), .SI(test_si38), .SE(n10251), .CLK(n10603), 
        .Q(g3684), .QN(n5881) );
  SDFFX1 DFF_536_Q_reg ( .D(g33612), .SI(g3684), .SE(n10216), .CLK(n10568), 
        .Q(g3639), .QN(n5591) );
  SDFFX1 DFF_537_Q_reg ( .D(g17787), .SI(g3639), .SE(n10216), .CLK(n10568), 
        .Q(g14597), .QN(n5579) );
  SDFFX1 DFF_538_Q_reg ( .D(g24268), .SI(g14597), .SE(n10243), .CLK(n10595), 
        .Q(g3338), .QN(n5527) );
  SDFFX1 DFF_539_Q_reg ( .D(g25716), .SI(g3338), .SE(n10203), .CLK(n10555), 
        .Q(g5406) );
  SDFFX1 DFF_541_Q_reg ( .D(g26906), .SI(g5406), .SE(n10203), .CLK(n10555), 
        .Q(g269), .QN(n9783) );
  SDFFX1 DFF_542_Q_reg ( .D(g24203), .SI(g269), .SE(n10270), .CLK(n10622), .Q(
        g401), .QN(n9726) );
  SDFFX1 DFF_543_Q_reg ( .D(g24346), .SI(g401), .SE(n10185), .CLK(n10537), .Q(
        g6040), .QN(n9900) );
  SDFFX1 DFF_544_Q_reg ( .D(g24207), .SI(g6040), .SE(n10171), .CLK(n10523), 
        .Q(g441) );
  SDFFX1 DFF_545_Q_reg ( .D(g25701), .SI(g441), .SE(n10207), .CLK(n10559), .Q(
        g9553), .QN(n5690) );
  SDFFX1 DFF_546_Q_reg ( .D(g29269), .SI(g9553), .SE(n10167), .CLK(n10519), 
        .Q(g3808), .QN(n5745) );
  SDFFX1 DFF_547_Q_reg ( .D(g34976), .SI(g3808), .SE(n10175), .CLK(n10527), 
        .Q(g9), .QN(n5468) );
  SDFFX1 DFF_549_Q_reg ( .D(g34255), .SI(g9), .SE(n10195), .CLK(n10547), .Q(
        test_so38), .QN(n10142) );
  SDFFX1 DFF_550_Q_reg ( .D(g30450), .SI(test_si39), .SE(n10183), .CLK(n10535), 
        .Q(g3957), .QN(n9989) );
  SDFFX1 DFF_551_Q_reg ( .D(g30456), .SI(g3957), .SE(n10239), .CLK(n10591), 
        .Q(g4093), .QN(n5340) );
  SDFFX1 DFF_552_Q_reg ( .D(g32991), .SI(g4093), .SE(n10220), .CLK(n10572), 
        .Q(g1760), .QN(n5602) );
  SDFFX1 DFF_554_Q_reg ( .D(g24348), .SI(g1760), .SE(n10220), .CLK(n10572), 
        .Q(g12422), .QN(n5437) );
  SDFFX1 DFF_555_Q_reg ( .D(g34249), .SI(g12422), .SE(n10210), .CLK(n10562), 
        .Q(g160), .QN(n5843) );
  SDFFX1 DFF_558_Q_reg ( .D(g30371), .SI(g160), .SE(n10193), .CLK(n10545), .Q(
        g2279), .QN(n5778) );
  SDFFX1 DFF_559_Q_reg ( .D(g29268), .SI(g2279), .SE(n10241), .CLK(n10593), 
        .Q(g3498) );
  SDFFX1 DFF_560_Q_reg ( .D(g29224), .SI(g3498), .SE(n10222), .CLK(n10574), 
        .Q(g586), .QN(n5336) );
  SDFFX1 DFF_561_Q_reg ( .D(g14189), .SI(g586), .SE(n10247), .CLK(n10599), .Q(
        g14201), .QN(n9593) );
  SDFFX1 DFF_562_Q_reg ( .D(g33017), .SI(g14201), .SE(n10213), .CLK(n10565), 
        .Q(g2619), .QN(n5508) );
  SDFFX1 DFF_563_Q_reg ( .D(g30339), .SI(g2619), .SE(n10213), .CLK(n10565), 
        .Q(g1183), .QN(n5599) );
  SDFFX1 DFF_564_Q_reg ( .D(g33967), .SI(g1183), .SE(n10219), .CLK(n10571), 
        .Q(g1608), .QN(n5792) );
  SDFFX1 DFF_565_Q_reg ( .D(g8784), .SI(g1608), .SE(n10235), .CLK(n10587), .Q(
        test_so39), .QN(n9765) );
  SDFFX1 DFF_566_Q_reg ( .D(g17519), .SI(test_si40), .SE(n10235), .CLK(n10587), 
        .Q(g17577), .QN(n9976) );
  SDFFX1 DFF_567_Q_reg ( .D(g33559), .SI(g17577), .SE(n10177), .CLK(n10529), 
        .Q(g1779), .QN(n5830) );
  SDFFX1 DFF_568_Q_reg ( .D(g29255), .SI(g1779), .SE(n10177), .CLK(n10529), 
        .Q(g2652), .QN(n9833) );
  SDFFX1 DFF_570_Q_reg ( .D(g30368), .SI(g2652), .SE(n10218), .CLK(n10570), 
        .Q(g2193), .QN(n5839) );
  SDFFX1 DFF_571_Q_reg ( .D(g30375), .SI(g2193), .SE(n10176), .CLK(n10528), 
        .Q(g2393), .QN(n5421) );
  SDFFX1 DFF_573_Q_reg ( .D(g28052), .SI(g2393), .SE(n10254), .CLK(n10606), 
        .Q(g661), .QN(n9789) );
  SDFFX1 DFF_574_Q_reg ( .D(g28089), .SI(g661), .SE(n10168), .CLK(n10520), .Q(
        g4950), .QN(n5772) );
  SDFFX1 DFF_575_Q_reg ( .D(g33055), .SI(g4950), .SE(n10246), .CLK(n10598), 
        .Q(g5535), .QN(n5566) );
  SDFFX1 DFF_576_Q_reg ( .D(g30392), .SI(g5535), .SE(n10201), .CLK(n10553), 
        .Q(g2834), .QN(g23652) );
  SDFFX1 DFF_577_Q_reg ( .D(g30343), .SI(g2834), .SE(n10201), .CLK(n10553), 
        .Q(g1361), .QN(n9761) );
  SDFFX1 DFF_579_Q_reg ( .D(g30523), .SI(g1361), .SE(n10229), .CLK(n10581), 
        .Q(g6235), .QN(n9965) );
  SDFFX1 DFF_580_Q_reg ( .D(g24233), .SI(g6235), .SE(n10229), .CLK(n10581), 
        .Q(g1146), .QN(n5851) );
  SDFFX1 DFF_581_Q_reg ( .D(g33018), .SI(g1146), .SE(n10213), .CLK(n10565), 
        .Q(test_so40), .QN(n10140) );
  SDFFX1 DFF_582_Q_reg ( .D(g32976), .SI(test_si41), .SE(n10209), .CLK(n10561), 
        .Q(g150), .QN(n5676) );
  SDFFX1 DFF_583_Q_reg ( .D(g30349), .SI(g150), .SE(n10166), .CLK(n10518), .Q(
        g1696), .QN(n5628) );
  SDFFX1 DFF_584_Q_reg ( .D(g33067), .SI(g1696), .SE(n10246), .CLK(n10598), 
        .Q(g6555), .QN(n10053) );
  SDFFX1 DFF_585_Q_reg ( .D(g26900), .SI(g6555), .SE(n10247), .CLK(n10599), 
        .Q(g14189), .QN(n9599) );
  SDFFX1 DFF_587_Q_reg ( .D(g33034), .SI(g14189), .SE(n10214), .CLK(n10566), 
        .Q(g3881), .QN(n5564) );
  SDFFX1 DFF_588_Q_reg ( .D(g30551), .SI(g3881), .SE(n10194), .CLK(n10546), 
        .Q(g6621), .QN(n9859) );
  SDFFX1 DFF_589_Q_reg ( .D(g25667), .SI(g6621), .SE(n10173), .CLK(n10525), 
        .Q(g3470), .QN(n5424) );
  SDFFX1 DFF_590_Q_reg ( .D(g30452), .SI(g3470), .SE(n10214), .CLK(n10566), 
        .Q(g3897) );
  SDFFX1 DFF_593_Q_reg ( .D(g34719), .SI(g518), .SE(n10210), .CLK(n10562), .Q(
        g538), .QN(n5491) );
  SDFFX1 DFF_594_Q_reg ( .D(g33607), .SI(g538), .SE(n10212), .CLK(n10564), .Q(
        g2606), .QN(n5311) );
  SDFFX1 DFF_595_Q_reg ( .D(g26923), .SI(g2606), .SE(n10200), .CLK(n10552), 
        .Q(g1472), .QN(n5290) );
  SDFFX1 DFF_597_Q_reg ( .D(g24211), .SI(g1472), .SE(n10172), .CLK(n10524), 
        .Q(test_so41) );
  SDFFX1 DFF_598_Q_reg ( .D(g33050), .SI(test_si42), .SE(n10253), .CLK(n10605), 
        .Q(g5188), .QN(n5567) );
  SDFFX1 DFF_599_Q_reg ( .D(g24341), .SI(g5188), .SE(n10233), .CLK(n10585), 
        .Q(g5689), .QN(n5529) );
  SDFFX1 DFF_600_Q_reg ( .D(g19334), .SI(g5689), .SE(n10233), .CLK(n10585), 
        .Q(g13259), .QN(n9744) );
  SDFFX1 DFF_601_Q_reg ( .D(g24201), .SI(g13259), .SE(n10237), .CLK(n10589), 
        .Q(g405), .QN(n9748) );
  SDFFX1 DFF_602_Q_reg ( .D(g30463), .SI(g405), .SE(n10217), .CLK(n10569), .Q(
        g5216), .QN(n9922) );
  SDFFX1 DFF_603_Q_reg ( .D(g9743), .SI(g5216), .SE(n10248), .CLK(n10600), .Q(
        g6494) );
  SDFFX1 DFF_604_Q_reg ( .D(g34464), .SI(g6494), .SE(n10181), .CLK(n10533), 
        .Q(g4669), .QN(n9590) );
  SDFFX1 DFF_606_Q_reg ( .D(g24243), .SI(g4669), .SE(n10252), .CLK(n10604), 
        .Q(g996), .QN(n9757) );
  SDFFX1 DFF_607_Q_reg ( .D(g24335), .SI(g996), .SE(n10199), .CLK(n10551), .Q(
        g4531) );
  SDFFX1 DFF_608_Q_reg ( .D(g34611), .SI(g4531), .SE(n10199), .CLK(n10551), 
        .Q(g2860), .QN(n10076) );
  SDFFX1 DFF_609_Q_reg ( .D(g34262), .SI(g2860), .SE(n10182), .CLK(n10534), 
        .Q(g4743), .QN(n5876) );
  SDFFX1 DFF_610_Q_reg ( .D(g30546), .SI(g4743), .SE(n10193), .CLK(n10545), 
        .Q(g6593), .QN(n10025) );
  SDFFX1 DFF_612_Q_reg ( .D(g25591), .SI(g6593), .SE(n10210), .CLK(n10562), 
        .Q(test_so42) );
  SDFFX1 DFF_613_Q_reg ( .D(g7257), .SI(test_si43), .SE(n10252), .CLK(n10604), 
        .Q(g4411) );
  SDFFX1 DFF_614_Q_reg ( .D(g30347), .SI(g4411), .SE(n10227), .CLK(n10579), 
        .Q(g1413), .QN(n9572) );
  SDFFX1 DFF_615_Q_reg ( .D(test_so38), .SI(g1413), .SE(n10195), .CLK(n10547), 
        .Q(g26960), .QN(n9788) );
  SDFFX1 DFF_616_Q_reg ( .D(g17577), .SI(g26960), .SE(n10235), .CLK(n10587), 
        .Q(g13039), .QN(n9953) );
  SDFFX1 DFF_617_Q_reg ( .D(g30556), .SI(g13039), .SE(n10249), .CLK(n10601), 
        .Q(g6641), .QN(n9800) );
  SDFFX1 DFF_619_Q_reg ( .D(g34970), .SI(g6641), .SE(n10249), .CLK(n10601), 
        .Q(g6) );
  SDFFX1 DFF_620_Q_reg ( .D(g33562), .SI(g6), .SE(n10218), .CLK(n10570), .Q(
        g1936), .QN(n5534) );
  SDFFX1 DFF_621_Q_reg ( .D(n10104), .SI(g1936), .SE(n10218), .CLK(n10570), 
        .Q(g55) );
  SDFFX1 DFF_622_Q_reg ( .D(g25610), .SI(g55), .SE(n10218), .CLK(n10570), .Q(
        g504), .QN(n5519) );
  SDFFX1 DFF_623_Q_reg ( .D(g33015), .SI(g504), .SE(n10269), .CLK(n10621), .Q(
        g2587), .QN(n5372) );
  SDFFX1 DFF_624_Q_reg ( .D(g31896), .SI(g2587), .SE(n10195), .CLK(n10547), 
        .Q(g4480) );
  SDFFX1 DFF_625_Q_reg ( .D(g34004), .SI(g4480), .SE(n10195), .CLK(n10547), 
        .Q(n9314), .QN(n18473) );
  SDFFX1 DFF_626_Q_reg ( .D(g30428), .SI(n9314), .SE(n10184), .CLK(n10536), 
        .Q(test_so43) );
  SDFFX1 DFF_627_Q_reg ( .D(g30485), .SI(test_si44), .SE(n10180), .CLK(n10532), 
        .Q(g5571), .QN(n9797) );
  SDFFX1 DFF_628_Q_reg ( .D(g30422), .SI(g5571), .SE(n10173), .CLK(n10525), 
        .Q(g3578), .QN(n9862) );
  SDFFX1 DFF_630_Q_reg ( .D(g25714), .SI(g3578), .SE(n10246), .CLK(n10598), 
        .Q(g9555), .QN(n18468) );
  SDFFX1 DFF_632_Q_reg ( .D(g29294), .SI(g9555), .SE(n10181), .CLK(n10533), 
        .Q(g5827), .QN(n5809) );
  SDFFX1 DFF_633_Q_reg ( .D(g30423), .SI(g5827), .SE(n10242), .CLK(n10594), 
        .Q(g3582), .QN(n9948) );
  SDFFX1 DFF_634_Q_reg ( .D(g30529), .SI(g3582), .SE(n10227), .CLK(n10579), 
        .Q(g6271), .QN(n9939) );
  SDFFX1 DFF_635_Q_reg ( .D(g34028), .SI(g6271), .SE(n10260), .CLK(n10612), 
        .Q(g4688), .QN(n5656) );
  SDFFX1 DFF_637_Q_reg ( .D(g33587), .SI(g4688), .SE(n10176), .CLK(n10528), 
        .Q(g2380), .QN(n9656) );
  SDFFX1 DFF_638_Q_reg ( .D(g30460), .SI(g2380), .SE(n10253), .CLK(n10605), 
        .Q(g5196), .QN(n9954) );
  SDFFX1 DFF_640_Q_reg ( .D(g30401), .SI(g5196), .SE(n10232), .CLK(n10584), 
        .Q(g3227), .QN(n9844) );
  SDFFX1 DFF_641_Q_reg ( .D(g33990), .SI(g3227), .SE(n10214), .CLK(n10566), 
        .Q(n9312), .QN(n18474) );
  SDFFX1 DFF_642_Q_reg ( .D(g16693), .SI(n9312), .SE(n10240), .CLK(n10592), 
        .Q(g14518) );
  SDFFX1 DFF_643_Q_reg ( .D(g17291), .SI(g14518), .SE(n10240), .CLK(n10592), 
        .Q(test_so44) );
  SDFFX1 DFF_644_Q_reg ( .D(g29309), .SI(test_si45), .SE(n10228), .CLK(n10580), 
        .Q(g6541) );
  SDFFX1 DFF_645_Q_reg ( .D(g30411), .SI(g6541), .SE(n10231), .CLK(n10583), 
        .Q(g3203), .QN(n9972) );
  SDFFX1 DFF_646_Q_reg ( .D(g33546), .SI(g3203), .SE(n10254), .CLK(n10606), 
        .Q(g1668), .QN(n5598) );
  SDFFX1 DFF_647_Q_reg ( .D(g28085), .SI(g1668), .SE(n10185), .CLK(n10537), 
        .Q(g4760), .QN(n5775) );
  SDFFX1 DFF_648_Q_reg ( .D(g26904), .SI(g4760), .SE(n10248), .CLK(n10600), 
        .Q(g262), .QN(n9782) );
  SDFFX1 DFF_649_Q_reg ( .D(g33556), .SI(g262), .SE(n10170), .CLK(n10522), .Q(
        g1840), .QN(n5451) );
  SDFFX1 DFF_651_Q_reg ( .D(g25722), .SI(g1840), .SE(n10184), .CLK(n10536), 
        .Q(g5467) );
  SDFFX1 DFF_652_Q_reg ( .D(g25605), .SI(g5467), .SE(n10184), .CLK(n10536), 
        .Q(g460), .QN(n9661) );
  SDFFX1 DFF_653_Q_reg ( .D(g33062), .SI(g460), .SE(n10242), .CLK(n10594), .Q(
        g6209), .QN(n10056) );
  SDFFX1 DFF_654_Q_reg ( .D(g26893), .SI(g6209), .SE(n10209), .CLK(n10561), 
        .Q(g29211) );
  SDFFX1 DFF_655_Q_reg ( .D(g12238), .SI(g29211), .SE(n10209), .CLK(n10561), 
        .Q(g14662), .QN(n5704) );
  SDFFX1 DFF_656_Q_reg ( .D(g28050), .SI(g14662), .SE(n10237), .CLK(n10589), 
        .Q(g655), .QN(n9820) );
  SDFFX1 DFF_657_Q_reg ( .D(g34626), .SI(g655), .SE(n10237), .CLK(n10589), .Q(
        test_so45) );
  SDFFX1 DFF_658_Q_reg ( .D(g33583), .SI(test_si46), .SE(n10178), .CLK(n10530), 
        .Q(g2204), .QN(n5620) );
  SDFFX1 DFF_659_Q_reg ( .D(g30472), .SI(g2204), .SE(n10178), .CLK(n10530), 
        .Q(g5256), .QN(n9811) );
  SDFFX1 DFF_660_Q_reg ( .D(g34454), .SI(g5256), .SE(n10259), .CLK(n10611), 
        .Q(g4608), .QN(n5274) );
  SDFFX1 DFF_661_Q_reg ( .D(g34850), .SI(g4608), .SE(n10259), .CLK(n10611), 
        .Q(g794), .QN(n5291) );
  SDFFX1 DFF_662_Q_reg ( .D(g16955), .SI(g794), .SE(n10259), .CLK(n10611), .Q(
        g13906), .QN(n5583) );
  SDFFX1 DFF_663_Q_reg ( .D(g10306), .SI(g13906), .SE(n10188), .CLK(n10540), 
        .Q(g4423), .QN(n9687) );
  SDFFX1 DFF_664_Q_reg ( .D(g24272), .SI(g4423), .SE(n10251), .CLK(n10603), 
        .Q(g3689), .QN(n5532) );
  SDFFX1 DFF_666_Q_reg ( .D(g17678), .SI(g3689), .SE(n10233), .CLK(n10585), 
        .Q(g5685) );
  SDFFX1 DFF_667_Q_reg ( .D(g24214), .SI(g5685), .SE(n10171), .CLK(n10523), 
        .Q(g703), .QN(n5821) );
  SDFFX1 DFF_669_Q_reg ( .D(g26909), .SI(g703), .SE(n10245), .CLK(n10597), .Q(
        g862), .QN(n5682) );
  SDFFX1 DFF_670_Q_reg ( .D(g30406), .SI(g862), .SE(n10265), .CLK(n10617), .Q(
        g3247), .QN(n9792) );
  SDFFX1 DFF_671_Q_reg ( .D(g33569), .SI(g3247), .SE(n10217), .CLK(n10569), 
        .Q(g2040), .QN(n5505) );
  SDFFX1 DFF_672_Q_reg ( .D(g25694), .SI(g2040), .SE(n10218), .CLK(n10570), 
        .Q(test_so46) );
  SDFFX1 DFF_673_Q_reg ( .D(g34628), .SI(test_si47), .SE(n10232), .CLK(n10584), 
        .Q(g4146), .QN(n5981) );
  SDFFX1 DFF_674_Q_reg ( .D(g34458), .SI(g4146), .SE(n10224), .CLK(n10576), 
        .Q(g4633), .QN(n5844) );
  SDFFX1 DFF_675_Q_reg ( .D(g24240), .SI(g4633), .SE(n10233), .CLK(n10585), 
        .Q(g7916), .QN(n5304) );
  SDFFX1 DFF_677_Q_reg ( .D(g34634), .SI(g7916), .SE(n10234), .CLK(n10586), 
        .Q(g4732), .QN(n5296) );
  SDFFX1 DFF_678_Q_reg ( .D(g25700), .SI(g4732), .SE(n10253), .CLK(n10605), 
        .Q(g9497), .QN(n5689) );
  SDFFX1 DFF_679_Q_reg ( .D(g29293), .SI(g9497), .SE(n10181), .CLK(n10533), 
        .Q(g5817), .QN(n9618) );
  SDFFX1 DFF_681_Q_reg ( .D(g33009), .SI(g5817), .SE(n10267), .CLK(n10619), 
        .Q(g2351), .QN(n5511) );
  SDFFX1 DFF_682_Q_reg ( .D(g33603), .SI(g2351), .SE(n10201), .CLK(n10553), 
        .Q(g2648), .QN(n9660) );
  SDFFX1 DFF_683_Q_reg ( .D(g24355), .SI(g2648), .SE(n10196), .CLK(n10548), 
        .Q(g6736), .QN(n10036) );
  SDFFX1 DFF_684_Q_reg ( .D(g34268), .SI(g6736), .SE(n10168), .CLK(n10520), 
        .Q(g4944), .QN(n5875) );
  SDFFX1 DFF_685_Q_reg ( .D(g25691), .SI(g4944), .SE(n10239), .CLK(n10591), 
        .Q(g4072), .QN(n10093) );
  SDFFX1 DFF_686_Q_reg ( .D(g26890), .SI(g4072), .SE(n10239), .CLK(n10591), 
        .Q(g7540), .QN(n9613) );
  SDFFX1 DFF_687_Q_reg ( .D(g7260), .SI(g7540), .SE(n10239), .CLK(n10591), .Q(
        test_so47) );
  SDFFX1 DFF_688_Q_reg ( .D(g29264), .SI(test_si48), .SE(n10173), .CLK(n10525), 
        .Q(g3466), .QN(n9639) );
  SDFFX1 DFF_689_Q_reg ( .D(g28072), .SI(g3466), .SE(n10246), .CLK(n10598), 
        .Q(g4116), .QN(n9589) );
  SDFFX1 DFF_690_Q_reg ( .D(g31900), .SI(g4116), .SE(n10202), .CLK(n10554), 
        .Q(g5041), .QN(n5605) );
  SDFFX1 DFF_692_Q_reg ( .D(g26956), .SI(g5041), .SE(n10258), .CLK(n10610), 
        .Q(g4434), .QN(n9675) );
  SDFFX1 DFF_693_Q_reg ( .D(g29271), .SI(g4434), .SE(n10167), .CLK(n10519), 
        .Q(g3827), .QN(n5808) );
  SDFFX1 DFF_694_Q_reg ( .D(g29304), .SI(g3827), .SE(n10189), .CLK(n10541), 
        .Q(g6500), .QN(n5748) );
  SDFFX1 DFF_695_Q_reg ( .D(g13049), .SI(g6500), .SE(n10233), .CLK(n10585), 
        .Q(g17813) );
  SDFFX1 DFF_696_Q_reg ( .D(g29261), .SI(g17813), .SE(n10190), .CLK(n10542), 
        .Q(g3133), .QN(n5661) );
  SDFFX1 DFF_697_Q_reg ( .D(g28063), .SI(g3133), .SE(n10232), .CLK(n10584), 
        .Q(g3333) );
  SDFFX1 DFF_698_Q_reg ( .D(g13259), .SI(g3333), .SE(n10232), .CLK(n10584), 
        .Q(g979), .QN(n5320) );
  SDFFX1 DFF_699_Q_reg ( .D(g34027), .SI(g979), .SE(n10260), .CLK(n10612), .Q(
        g4681), .QN(n10040) );
  SDFFX1 DFF_700_Q_reg ( .D(g33961), .SI(g4681), .SE(n10263), .CLK(n10615), 
        .Q(g298), .QN(n5675) );
  SDFFX1 DFF_702_Q_reg ( .D(g33604), .SI(g298), .SE(n10177), .CLK(n10529), .Q(
        test_so48), .QN(n10156) );
  SDFFX1 DFF_704_Q_reg ( .D(g8788), .SI(test_si49), .SE(n10206), .CLK(n10558), 
        .Q(g8789), .QN(n9767) );
  SDFFX1 DFF_705_Q_reg ( .D(g32995), .SI(g8789), .SE(n10266), .CLK(n10618), 
        .Q(g1894), .QN(n5374) );
  SDFFX1 DFF_706_Q_reg ( .D(g34624), .SI(g1894), .SE(n10188), .CLK(n10540), 
        .Q(g2988), .QN(n10074) );
  SDFFX1 DFF_707_Q_reg ( .D(g30415), .SI(g2988), .SE(n10241), .CLK(n10593), 
        .Q(g3538), .QN(n9963) );
  SDFFX1 DFF_708_Q_reg ( .D(g33536), .SI(g3538), .SE(n10210), .CLK(n10562), 
        .Q(g301), .QN(n10096) );
  SDFFX1 DFF_709_Q_reg ( .D(g26888), .SI(g301), .SE(n10249), .CLK(n10601), .Q(
        n9306) );
  SDFFX1 DFF_710_Q_reg ( .D(g28055), .SI(n9306), .SE(n10186), .CLK(n10538), 
        .Q(g827), .QN(n5728) );
  SDFFX1 DFF_711_Q_reg ( .D(g24238), .SI(g827), .SE(n10192), .CLK(n10544), .Q(
        g17291), .QN(n9715) );
  SDFFX1 DFF_713_Q_reg ( .D(g33600), .SI(g17291), .SE(n10249), .CLK(n10601), 
        .Q(g2555), .QN(n5351) );
  SDFFX1 DFF_714_Q_reg ( .D(g28105), .SI(g2555), .SE(n10194), .CLK(n10546), 
        .Q(g5011), .QN(n9669) );
  SDFFX1 DFF_715_Q_reg ( .D(g34721), .SI(g5011), .SE(n10210), .CLK(n10562), 
        .Q(g199), .QN(n10098) );
  SDFFX1 DFF_716_Q_reg ( .D(g29307), .SI(g199), .SE(n10189), .CLK(n10541), .Q(
        g6523), .QN(n5870) );
  SDFFX1 DFF_717_Q_reg ( .D(g30345), .SI(g6523), .SE(n10236), .CLK(n10588), 
        .Q(test_so49), .QN(n10127) );
  SDFFX1 DFF_718_Q_reg ( .D(g34453), .SI(test_si50), .SE(n10259), .CLK(n10611), 
        .Q(g4601), .QN(n5365) );
  SDFFX1 DFF_719_Q_reg ( .D(g32980), .SI(g4601), .SE(n10171), .CLK(n10523), 
        .Q(g854) );
  SDFFX1 DFF_720_Q_reg ( .D(g29238), .SI(g854), .SE(n10200), .CLK(n10552), .Q(
        g1484), .QN(n5865) );
  SDFFX1 DFF_721_Q_reg ( .D(g34639), .SI(g1484), .SE(n10200), .CLK(n10552), 
        .Q(g4922), .QN(n5346) );
  SDFFX1 DFF_722_Q_reg ( .D(g25695), .SI(g4922), .SE(n10165), .CLK(n10517), 
        .Q(g5080), .QN(n5893) );
  SDFFX1 DFF_723_Q_reg ( .D(g33057), .SI(g5080), .SE(n10242), .CLK(n10594), 
        .Q(g5863), .QN(n10055) );
  SDFFX1 DFF_724_Q_reg ( .D(g26969), .SI(g5863), .SE(n10242), .CLK(n10594), 
        .Q(g4581), .QN(n5670) );
  SDFFX1 DFF_726_Q_reg ( .D(g29253), .SI(g4581), .SE(n10206), .CLK(n10558), 
        .Q(g2518), .QN(n9831) );
  SDFFX1 DFF_727_Q_reg ( .D(g34021), .SI(g2518), .SE(n10201), .CLK(n10553), 
        .Q(g2567), .QN(n9622) );
  SDFFX1 DFF_728_Q_reg ( .D(g26895), .SI(g2567), .SE(n10223), .CLK(n10575), 
        .Q(g568), .QN(n5335) );
  SDFFX1 DFF_729_Q_reg ( .D(g30413), .SI(g568), .SE(n10232), .CLK(n10584), .Q(
        g3263), .QN(n9791) );
  SDFFX1 DFF_730_Q_reg ( .D(g30549), .SI(g3263), .SE(n10193), .CLK(n10545), 
        .Q(g6613), .QN(n9840) );
  SDFFX1 DFF_731_Q_reg ( .D(g24347), .SI(g6613), .SE(n10185), .CLK(n10537), 
        .Q(test_so50), .QN(n10161) );
  SDFFX1 DFF_732_Q_reg ( .D(g25758), .SI(test_si51), .SE(n10257), .CLK(n10609), 
        .Q(g6444) );
  SDFFX1 DFF_733_Q_reg ( .D(g34808), .SI(g6444), .SE(n10165), .CLK(n10517), 
        .Q(g2965), .QN(n9732) );
  SDFFX1 DFF_734_Q_reg ( .D(g30501), .SI(g2965), .SE(n10244), .CLK(n10596), 
        .Q(g5857), .QN(n5573) );
  SDFFX1 DFF_735_Q_reg ( .D(g33969), .SI(g5857), .SE(n10219), .CLK(n10571), 
        .Q(n9303), .QN(n18475) );
  SDFFX1 DFF_736_Q_reg ( .D(g34440), .SI(n9303), .SE(n10171), .CLK(n10523), 
        .Q(g890), .QN(n5305) );
  SDFFX1 DFF_737_Q_reg ( .D(g17607), .SI(g890), .SE(n10223), .CLK(n10575), .Q(
        g17646), .QN(n9981) );
  SDFFX1 DFF_738_Q_reg ( .D(g30433), .SI(g17646), .SE(n10185), .CLK(n10537), 
        .Q(g3562), .QN(n10027) );
  SDFFX1 DFF_739_Q_reg ( .D(g21900), .SI(g3562), .SE(n10185), .CLK(n10537), 
        .Q(g10122_Tj) );
  SDFFX1 DFF_740_Q_reg ( .D(g26921), .SI(g10122_Tj), .SE(n10212), .CLK(n10564), 
        .Q(g1404), .QN(n9753) );
  SDFFX1 DFF_742_Q_reg ( .D(g29270), .SI(g1404), .SE(n10167), .CLK(n10519), 
        .Q(g3817), .QN(n9617) );
  SDFFX1 DFF_743_Q_reg ( .D(n10110), .SI(g3817), .SE(n10168), .CLK(n10520), 
        .Q(n9302), .QN(n6010) );
  SDFFX1 DFF_744_Q_reg ( .D(g33038), .SI(n9302), .SE(n10244), .CLK(n10596), 
        .Q(g4501) );
  SDFFX1 DFF_745_Q_reg ( .D(g31865), .SI(g4501), .SE(n10260), .CLK(n10612), 
        .Q(test_so51), .QN(n10155) );
  SDFFX1 DFF_746_Q_reg ( .D(g26926), .SI(test_si52), .SE(n10256), .CLK(n10608), 
        .Q(g2724), .QN(n5301) );
  SDFFX1 DFF_747_Q_reg ( .D(g28083), .SI(g2724), .SE(n10178), .CLK(n10530), 
        .Q(g4704), .QN(n5771) );
  SDFFX1 DFF_749_Q_reg ( .D(g34797), .SI(g22), .SE(n10166), .CLK(n10518), .Q(
        g2878), .QN(n10085) );
  SDFFX1 DFF_750_Q_reg ( .D(g30478), .SI(g2878), .SE(n10217), .CLK(n10569), 
        .Q(g5220), .QN(n9915) );
  SDFFX1 DFF_751_Q_reg ( .D(g34724), .SI(g5220), .SE(n10223), .CLK(n10575), 
        .Q(g617), .QN(n5339) );
  SDFFX1 DFF_752_Q_reg ( .D(g24212), .SI(g617), .SE(n10223), .CLK(n10575), .Q(
        g12368) );
  SDFFX1 DFF_753_Q_reg ( .D(g26883), .SI(g12368), .SE(n10249), .CLK(n10601), 
        .Q(g316), .QN(n9663) );
  SDFFX1 DFF_754_Q_reg ( .D(g32985), .SI(g316), .SE(n10269), .CLK(n10621), .Q(
        g1277), .QN(n10095) );
  SDFFX1 DFF_755_Q_reg ( .D(g25761), .SI(g1277), .SE(n10189), .CLK(n10541), 
        .Q(g6513), .QN(n5426) );
  SDFFX1 DFF_756_Q_reg ( .D(g26886), .SI(g6513), .SE(n10238), .CLK(n10590), 
        .Q(g336), .QN(n5824) );
  SDFFX1 DFF_757_Q_reg ( .D(g34796), .SI(g336), .SE(n10166), .CLK(n10518), .Q(
        g2882), .QN(n9575) );
  SDFFX1 DFF_758_Q_reg ( .D(g32982), .SI(g2882), .SE(n10197), .CLK(n10549), 
        .Q(test_so52), .QN(n10100) );
  SDFFX1 DFF_759_Q_reg ( .D(g33561), .SI(test_si53), .SE(n10218), .CLK(n10570), 
        .Q(g1906), .QN(n5503) );
  SDFFX1 DFF_760_Q_reg ( .D(g26880), .SI(g1906), .SE(n10218), .CLK(n10570), 
        .Q(g305), .QN(n5282) );
  SDFFX1 DFF_761_Q_reg ( .D(g34975), .SI(g305), .SE(n10191), .CLK(n10543), .Q(
        g8), .QN(n9673) );
  SDFFX1 DFF_763_Q_reg ( .D(g26931), .SI(g8), .SE(n10219), .CLK(n10571), .Q(
        g2799), .QN(n9605) );
  SDFFX1 DFF_764_Q_reg ( .D(g14147), .SI(g2799), .SE(n10247), .CLK(n10599), 
        .Q(g14167), .QN(n9600) );
  SDFFX1 DFF_765_Q_reg ( .D(g13039), .SI(g14167), .SE(n10247), .CLK(n10599), 
        .Q(g17787) );
  SDFFX1 DFF_766_Q_reg ( .D(g34641), .SI(g17787), .SE(n10247), .CLK(n10599), 
        .Q(g4912), .QN(n5297) );
  SDFFX1 DFF_767_Q_reg ( .D(g34629), .SI(g4912), .SE(n10247), .CLK(n10599), 
        .Q(g4157), .QN(n5983) );
  SDFFX1 DFF_768_Q_reg ( .D(g33598), .SI(g4157), .SE(n10207), .CLK(n10559), 
        .Q(g2541), .QN(n5461) );
  SDFFX1 DFF_769_Q_reg ( .D(g33576), .SI(g2541), .SE(n10218), .CLK(n10570), 
        .Q(g2153), .QN(n5356) );
  SDFFX1 DFF_770_Q_reg ( .D(g34720), .SI(g2153), .SE(n10172), .CLK(n10524), 
        .Q(g550), .QN(n10097) );
  SDFFX1 DFF_771_Q_reg ( .D(g26902), .SI(g550), .SE(n10248), .CLK(n10600), .Q(
        g255), .QN(n9781) );
  SDFFX1 DFF_772_Q_reg ( .D(g29244), .SI(g255), .SE(n10198), .CLK(n10550), .Q(
        test_so53), .QN(n10151) );
  SDFFX1 DFF_773_Q_reg ( .D(g30468), .SI(test_si54), .SE(n10253), .CLK(n10605), 
        .Q(g5240), .QN(n9943) );
  SDFFX1 DFF_774_Q_reg ( .D(g26924), .SI(g5240), .SE(n10236), .CLK(n10588), 
        .Q(g1478), .QN(n5289) );
  SDFFX1 DFF_776_Q_reg ( .D(g33031), .SI(g1478), .SE(n10241), .CLK(n10593), 
        .Q(g3863), .QN(n10054) );
  SDFFX1 DFF_777_Q_reg ( .D(g29245), .SI(g3863), .SE(n10266), .CLK(n10618), 
        .Q(g1959), .QN(n9830) );
  SDFFX1 DFF_778_Q_reg ( .D(g29266), .SI(g1959), .SE(n10173), .CLK(n10525), 
        .Q(g3480), .QN(n5868) );
  SDFFX1 DFF_779_Q_reg ( .D(g30559), .SI(g3480), .SE(n10194), .CLK(n10546), 
        .Q(g6653) );
  SDFFX1 DFF_780_Q_reg ( .D(g14749), .SI(g6653), .SE(n10264), .CLK(n10616), 
        .Q(g17764) );
  SDFFX1 DFF_781_Q_reg ( .D(g34794), .SI(g17764), .SE(n10166), .CLK(n10518), 
        .Q(g2864), .QN(n5489) );
  SDFFX1 DFF_782_Q_reg ( .D(g28087), .SI(g2864), .SE(n10196), .CLK(n10548), 
        .Q(g4894), .QN(n5774) );
  SDFFX1 DFF_783_Q_reg ( .D(g14635), .SI(g4894), .SE(n10233), .CLK(n10585), 
        .Q(g17678) );
  SDFFX1 DFF_784_Q_reg ( .D(g30435), .SI(g17678), .SE(n10240), .CLK(n10592), 
        .Q(g3857), .QN(n5572) );
  SDFFX1 DFF_785_Q_reg ( .D(g16659), .SI(g3857), .SE(n10240), .CLK(n10592), 
        .Q(g16693), .QN(n9990) );
  SDFFX1 DFF_786_Q_reg ( .D(g25609), .SI(g16693), .SE(n10254), .CLK(n10606), 
        .Q(test_so54), .QN(n10135) );
  SDFFX1 DFF_788_Q_reg ( .D(g28057), .SI(test_si55), .SE(n10252), .CLK(n10604), 
        .Q(g1002), .QN(n9751) );
  SDFFX1 DFF_789_Q_reg ( .D(g34439), .SI(g1002), .SE(n10252), .CLK(n10604), 
        .Q(g776), .QN(n5330) );
  SDFFX1 DFF_790_Q_reg ( .D(g34979), .SI(g776), .SE(n10252), .CLK(n10604), .Q(
        g28), .QN(n5324) );
  SDFFX1 DFF_791_Q_reg ( .D(g10500), .SI(g28), .SE(n10252), .CLK(n10604), .Q(
        g1236), .QN(n9721) );
  SDFFX1 DFF_792_Q_reg ( .D(g34260), .SI(g1236), .SE(n10261), .CLK(n10613), 
        .Q(g4646), .QN(n5712) );
  SDFFX1 DFF_793_Q_reg ( .D(g33012), .SI(g4646), .SE(n10268), .CLK(n10620), 
        .Q(g2476), .QN(n10043) );
  SDFFX1 DFF_794_Q_reg ( .D(g32989), .SI(g2476), .SE(n10202), .CLK(n10554), 
        .Q(g1657), .QN(n5525) );
  SDFFX1 DFF_795_Q_reg ( .D(g34006), .SI(g1657), .SE(n10176), .CLK(n10528), 
        .Q(g2375), .QN(n9694) );
  SDFFX1 DFF_796_Q_reg ( .D(g34783), .SI(g2375), .SE(n10205), .CLK(n10557), 
        .Q(g63), .QN(n9738) );
  SDFFX1 DFF_797_Q_reg ( .D(g14738), .SI(g63), .SE(n10205), .CLK(n10557), .Q(
        g17739), .QN(n9885) );
  SDFFX1 DFF_798_Q_reg ( .D(g8719), .SI(g17739), .SE(n10245), .CLK(n10597), 
        .Q(g358), .QN(n9785) );
  SDFFX1 DFF_799_Q_reg ( .D(g26910), .SI(g358), .SE(n10245), .CLK(n10597), .Q(
        g896), .QN(n5431) );
  SDFFX1 DFF_802_Q_reg ( .D(g28043), .SI(g896), .SE(n10260), .CLK(n10612), .Q(
        test_so55), .QN(n10154) );
  SDFFX1 DFF_803_Q_reg ( .D(g33021), .SI(test_si56), .SE(n10246), .CLK(n10598), 
        .Q(g3161), .QN(n10062) );
  SDFFX1 DFF_804_Q_reg ( .D(g29251), .SI(g3161), .SE(n10195), .CLK(n10547), 
        .Q(g2384), .QN(n9825) );
  SDFFX1 DFF_806_Q_reg ( .D(test_so80), .SI(g2384), .SE(n10195), .CLK(n10547), 
        .Q(g14828), .QN(n5700) );
  SDFFX1 DFF_807_Q_reg ( .D(g34456), .SI(g14828), .SE(n10263), .CLK(n10615), 
        .Q(g4616), .QN(n5608) );
  SDFFX1 DFF_808_Q_reg ( .D(g26968), .SI(g4616), .SE(n10263), .CLK(n10615), 
        .Q(g4561) );
  SDFFX1 DFF_809_Q_reg ( .D(g33991), .SI(g4561), .SE(n10214), .CLK(n10566), 
        .Q(g2024), .QN(n5801) );
  SDFFX1 DFF_810_Q_reg ( .D(g8279), .SI(g2024), .SE(n10242), .CLK(n10594), .Q(
        g3451) );
  SDFFX1 DFF_811_Q_reg ( .D(g26930), .SI(g3451), .SE(n10204), .CLK(n10556), 
        .Q(g2795), .QN(n9606) );
  SDFFX1 DFF_812_Q_reg ( .D(g34599), .SI(g2795), .SE(n10222), .CLK(n10574), 
        .Q(g613), .QN(n5474) );
  SDFFX1 DFF_813_Q_reg ( .D(g28082), .SI(g613), .SE(n10205), .CLK(n10557), .Q(
        g4527), .QN(n10071) );
  SDFFX1 DFF_814_Q_reg ( .D(g33557), .SI(g4527), .SE(n10170), .CLK(n10522), 
        .Q(g1844), .QN(n5847) );
  SDFFX1 DFF_815_Q_reg ( .D(g30511), .SI(g1844), .SE(n10186), .CLK(n10538), 
        .Q(g5937), .QN(n9886) );
  SDFFX1 DFF_816_Q_reg ( .D(g33045), .SI(g5937), .SE(n10243), .CLK(n10595), 
        .Q(test_so56) );
  SDFFX1 DFF_818_Q_reg ( .D(g30379), .SI(test_si57), .SE(n10206), .CLK(n10558), 
        .Q(g2523), .QN(n5281) );
  SDFFX1 DFF_819_Q_reg ( .D(g24267), .SI(g2523), .SE(n10243), .CLK(n10595), 
        .Q(g11349), .QN(n5436) );
  SDFFX1 DFF_820_Q_reg ( .D(g34020), .SI(g11349), .SE(n10201), .CLK(n10553), 
        .Q(g2643), .QN(n9693) );
  SDFFX1 DFF_822_Q_reg ( .D(g24249), .SI(g2643), .SE(n10236), .CLK(n10588), 
        .Q(g1489), .QN(n5850) );
  SDFFX1 DFF_824_Q_reg ( .D(g25592), .SI(g1489), .SE(n10210), .CLK(n10562), 
        .Q(g8358), .QN(n9759) );
  SDFFX1 DFF_825_Q_reg ( .D(g30382), .SI(g8358), .SE(n10207), .CLK(n10559), 
        .Q(n9295), .QN(n18481) );
  SDFFX1 DFF_826_Q_reg ( .D(g29285), .SI(n9295), .SE(n10207), .CLK(n10559), 
        .Q(g5156) );
  SDFFX1 DFF_828_Q_reg ( .D(g12919), .SI(g5156), .SE(n10223), .CLK(n10575), 
        .Q(g30332), .QN(n5526) );
  SDFFX1 DFF_829_Q_reg ( .D(g34975), .SI(g30332), .SE(n10224), .CLK(n10576), 
        .Q(n9294) );
  SDFFX1 DFF_830_Q_reg ( .D(g25662), .SI(n9294), .SE(n10242), .CLK(n10594), 
        .Q(g8279), .QN(n5717) );
  SDFFX1 DFF_831_Q_reg ( .D(g21896), .SI(g8279), .SE(n10230), .CLK(n10582), 
        .Q(g8839) );
  SDFFX1 DFF_832_Q_reg ( .D(g33563), .SI(g8839), .SE(n10198), .CLK(n10550), 
        .Q(g1955), .QN(n9653) );
  SDFFX1 DFF_833_Q_reg ( .D(g33622), .SI(g1955), .SE(n10261), .CLK(n10613), 
        .Q(test_so57), .QN(n10122) );
  SDFFX1 DFF_835_Q_reg ( .D(g33582), .SI(test_si58), .SE(n10193), .CLK(n10545), 
        .Q(g2273), .QN(n5458) );
  SDFFX1 DFF_836_Q_reg ( .D(g17871), .SI(g2273), .SE(n10264), .CLK(n10616), 
        .Q(g14749), .QN(n5584) );
  SDFFX1 DFF_837_Q_reg ( .D(g28086), .SI(g14749), .SE(n10220), .CLK(n10572), 
        .Q(g4771), .QN(n5769) );
  SDFFX1 DFF_838_Q_reg ( .D(g25744), .SI(g4771), .SE(n10220), .CLK(n10572), 
        .Q(g6098) );
  SDFFX1 DFF_839_Q_reg ( .D(g29262), .SI(g6098), .SE(n10255), .CLK(n10607), 
        .Q(g3147) );
  SDFFX1 DFF_840_Q_reg ( .D(g24270), .SI(g3147), .SE(n10255), .CLK(n10607), 
        .Q(g3347), .QN(n9896) );
  SDFFX1 DFF_841_Q_reg ( .D(g33581), .SI(g3347), .SE(n10193), .CLK(n10545), 
        .Q(g2269), .QN(n5410) );
  SDFFX1 DFF_842_Q_reg ( .D(g8358), .SI(g2269), .SE(n10210), .CLK(n10562), .Q(
        g191), .QN(n9760) );
  SDFFX1 DFF_843_Q_reg ( .D(g24266), .SI(g191), .SE(n10256), .CLK(n10608), .Q(
        g2712), .QN(n9630) );
  SDFFX1 DFF_844_Q_reg ( .D(g34849), .SI(g2712), .SE(n10223), .CLK(n10575), 
        .Q(g626), .QN(n5288) );
  SDFFX1 DFF_846_Q_reg ( .D(g33618), .SI(g2729), .SE(n10262), .CLK(n10614), 
        .Q(g5357), .QN(n5393) );
  SDFFX1 DFF_847_Q_reg ( .D(g34038), .SI(g5357), .SE(n10225), .CLK(n10577), 
        .Q(test_so58), .QN(n10123) );
  SDFFX1 DFF_848_Q_reg ( .D(g13068), .SI(test_si59), .SE(n10204), .CLK(n10556), 
        .Q(g17819) );
  SDFFX1 DFF_849_Q_reg ( .D(g34032), .SI(g17819), .SE(n10205), .CLK(n10557), 
        .Q(g4709), .QN(n5518) );
  SDFFX1 DFF_852_Q_reg ( .D(g34803), .SI(g4709), .SE(n10183), .CLK(n10535), 
        .Q(g2927), .QN(n9729) );
  SDFFX1 DFF_853_Q_reg ( .D(g34459), .SI(g2927), .SE(n10173), .CLK(n10525), 
        .Q(g4340), .QN(n5653) );
  SDFFX1 DFF_854_Q_reg ( .D(g30509), .SI(g4340), .SE(n10187), .CLK(n10539), 
        .Q(g5929), .QN(n9850) );
  SDFFX1 DFF_855_Q_reg ( .D(g34640), .SI(g5929), .SE(n10200), .CLK(n10552), 
        .Q(g4907), .QN(n5295) );
  SDFFX1 DFF_856_Q_reg ( .D(g14421), .SI(g4907), .SE(n10200), .CLK(n10552), 
        .Q(g16874) );
  SDFFX1 DFF_857_Q_reg ( .D(g28069), .SI(g16874), .SE(n10265), .CLK(n10617), 
        .Q(g4035), .QN(n9671) );
  SDFFX1 DFF_858_Q_reg ( .D(g21899), .SI(g4035), .SE(n10265), .CLK(n10617), 
        .Q(g2946), .QN(n10087) );
  SDFFX1 DFF_859_Q_reg ( .D(g31868), .SI(g2946), .SE(n10197), .CLK(n10549), 
        .Q(g918), .QN(n5673) );
  SDFFX1 DFF_860_Q_reg ( .D(g26938), .SI(g918), .SE(n10239), .CLK(n10591), .Q(
        g4082), .QN(n9739) );
  SDFFX1 DFF_861_Q_reg ( .D(g25756), .SI(g4082), .SE(n10248), .CLK(n10600), 
        .Q(g9743), .QN(n5719) );
  SDFFX1 DFF_862_Q_reg ( .D(g30363), .SI(g9743), .SE(n10268), .CLK(n10620), 
        .Q(test_so59) );
  SDFFX1 DFF_863_Q_reg ( .D(g30334), .SI(test_si60), .SE(n10222), .CLK(n10574), 
        .Q(g577), .QN(n5294) );
  SDFFX1 DFF_864_Q_reg ( .D(g33970), .SI(g577), .SE(n10219), .CLK(n10571), .Q(
        g1620), .QN(n5791) );
  SDFFX1 DFF_865_Q_reg ( .D(g30391), .SI(g1620), .SE(n10199), .CLK(n10551), 
        .Q(g2831), .QN(g30331) );
  SDFFX1 DFF_866_Q_reg ( .D(g25615), .SI(g2831), .SE(n10199), .CLK(n10551), 
        .Q(g667) );
  SDFFX1 DFF_867_Q_reg ( .D(g33540), .SI(g667), .SE(n10197), .CLK(n10549), .Q(
        g930), .QN(n5731) );
  SDFFX1 DFF_868_Q_reg ( .D(g30445), .SI(g930), .SE(n10215), .CLK(n10567), .Q(
        g3937), .QN(n9889) );
  SDFFX1 DFF_870_Q_reg ( .D(g25617), .SI(g3937), .SE(n10186), .CLK(n10538), 
        .Q(g817), .QN(n5822) );
  SDFFX1 DFF_871_Q_reg ( .D(g24247), .SI(g817), .SE(n10229), .CLK(n10581), .Q(
        g1249), .QN(n9742) );
  SDFFX1 DFF_872_Q_reg ( .D(g24215), .SI(g1249), .SE(n10186), .CLK(n10538), 
        .Q(g837), .QN(n5562) );
  SDFFX1 DFF_873_Q_reg ( .D(g14451), .SI(g837), .SE(n10221), .CLK(n10573), .Q(
        g16924) );
  SDFFX1 DFF_874_Q_reg ( .D(g33964), .SI(g16924), .SE(n10222), .CLK(n10574), 
        .Q(g599), .QN(n5550) );
  SDFFX1 DFF_875_Q_reg ( .D(g25719), .SI(g599), .SE(n10169), .CLK(n10521), .Q(
        g5475), .QN(n5425) );
  SDFFX1 DFF_876_Q_reg ( .D(g29228), .SI(g5475), .SE(n10213), .CLK(n10565), 
        .Q(test_so60) );
  SDFFX1 DFF_877_Q_reg ( .D(g30514), .SI(test_si61), .SE(n10269), .CLK(n10621), 
        .Q(g5949), .QN(n9814) );
  SDFFX1 DFF_878_Q_reg ( .D(g33627), .SI(g5949), .SE(n10196), .CLK(n10548), 
        .Q(g6682), .QN(n5590) );
  SDFFX1 DFF_880_Q_reg ( .D(g24231), .SI(g6682), .SE(n10196), .CLK(n10548), 
        .Q(g904), .QN(n9741) );
  SDFFX1 DFF_881_Q_reg ( .D(g34615), .SI(g904), .SE(n10196), .CLK(n10548), .Q(
        g2873), .QN(n5488) );
  SDFFX1 DFF_882_Q_reg ( .D(g30356), .SI(g2873), .SE(n10170), .CLK(n10522), 
        .Q(g1854), .QN(n5785) );
  SDFFX1 DFF_883_Q_reg ( .D(g25696), .SI(g1854), .SE(n10165), .CLK(n10517), 
        .Q(g5084), .QN(n5681) );
  SDFFX1 DFF_884_Q_reg ( .D(g30493), .SI(g5084), .SE(n10180), .CLK(n10532), 
        .Q(g5603), .QN(n9796) );
  SDFFX1 DFF_885_Q_reg ( .D(g8917), .SI(g5603), .SE(n10175), .CLK(n10527), .Q(
        g8870), .QN(n5726) );
  SDFFX1 DFF_886_Q_reg ( .D(g33594), .SI(g8870), .SE(n10211), .CLK(n10563), 
        .Q(g2495), .QN(n5522) );
  SDFFX1 DFF_887_Q_reg ( .D(g34009), .SI(g2495), .SE(n10268), .CLK(n10620), 
        .Q(g2437), .QN(n5789) );
  SDFFX1 DFF_888_Q_reg ( .D(g30365), .SI(g2437), .SE(n10204), .CLK(n10556), 
        .Q(g2102), .QN(n5666) );
  SDFFX1 DFF_889_Q_reg ( .D(g33004), .SI(g2102), .SE(n10264), .CLK(n10616), 
        .Q(g2208), .QN(n10045) );
  SDFFX1 DFF_890_Q_reg ( .D(g34018), .SI(g2208), .SE(n10212), .CLK(n10564), 
        .Q(test_so61) );
  SDFFX1 DFF_891_Q_reg ( .D(g25685), .SI(test_si62), .SE(n10239), .CLK(n10591), 
        .Q(g4064), .QN(n5416) );
  SDFFX1 DFF_892_Q_reg ( .D(g34040), .SI(g4064), .SE(n10205), .CLK(n10557), 
        .Q(g4899), .QN(n5517) );
  SDFFX1 DFF_893_Q_reg ( .D(g25639), .SI(g4899), .SE(n10256), .CLK(n10608), 
        .Q(g2719), .QN(n5465) );
  SDFFX1 DFF_894_Q_reg ( .D(g34029), .SI(g2719), .SE(n10264), .CLK(n10616), 
        .Q(g4785), .QN(n5361) );
  SDFFX1 DFF_895_Q_reg ( .D(g30488), .SI(g4785), .SE(n10174), .CLK(n10526), 
        .Q(g5583), .QN(n9853) );
  SDFFX1 DFF_896_Q_reg ( .D(g34600), .SI(g5583), .SE(n10253), .CLK(n10605), 
        .Q(g781), .QN(n5551) );
  SDFFX1 DFF_897_Q_reg ( .D(g29300), .SI(g781), .SE(n10179), .CLK(n10531), .Q(
        g6173), .QN(n5810) );
  SDFFX1 DFF_898_Q_reg ( .D(g14705), .SI(g6173), .SE(n10235), .CLK(n10587), 
        .Q(g17743) );
  SDFFX1 DFF_899_Q_reg ( .D(g34802), .SI(g17743), .SE(n10183), .CLK(n10535), 
        .Q(g2917), .QN(n9730) );
  SDFFX1 DFF_900_Q_reg ( .D(g25614), .SI(g2917), .SE(n10238), .CLK(n10590), 
        .Q(g686), .QN(n9629) );
  SDFFX1 DFF_901_Q_reg ( .D(g28058), .SI(g686), .SE(n10211), .CLK(n10563), .Q(
        g1252), .QN(n5554) );
  SDFFX1 DFF_902_Q_reg ( .D(g29225), .SI(g1252), .SE(n10199), .CLK(n10551), 
        .Q(g671), .QN(n9626) );
  SDFFX1 DFF_903_Q_reg ( .D(g33580), .SI(g671), .SE(n10193), .CLK(n10545), .Q(
        test_so62), .QN(n10157) );
  SDFFX1 DFF_904_Q_reg ( .D(g30532), .SI(test_si63), .SE(n10226), .CLK(n10578), 
        .Q(g6283), .QN(n9895) );
  SDFFX1 DFF_905_Q_reg ( .D(g17845), .SI(g6283), .SE(n10235), .CLK(n10587), 
        .Q(g14705), .QN(n5586) );
  SDFFX1 DFF_906_Q_reg ( .D(g17674), .SI(g14705), .SE(n10235), .CLK(n10587), 
        .Q(g17519), .QN(n9868) );
  SDFFX1 DFF_909_Q_reg ( .D(g8783), .SI(g17519), .SE(n10235), .CLK(n10587), 
        .Q(g8784), .QN(DFF_909_n1) );
  SDFFX1 DFF_910_Q_reg ( .D(g33054), .SI(g8784), .SE(n10246), .CLK(n10598), 
        .Q(g5527), .QN(n5389) );
  SDFFX1 DFF_911_Q_reg ( .D(g26962), .SI(g5527), .SE(n10248), .CLK(n10600), 
        .Q(g4489), .QN(n10060) );
  SDFFX1 DFF_912_Q_reg ( .D(g33564), .SI(g4489), .SE(n10169), .CLK(n10521), 
        .Q(g1974), .QN(n5450) );
  SDFFX1 DFF_913_Q_reg ( .D(g32984), .SI(g1974), .SE(n10211), .CLK(n10563), 
        .Q(g1270), .QN(n5716) );
  SDFFX1 DFF_914_Q_reg ( .D(g34039), .SI(g1270), .SE(n10225), .CLK(n10577), 
        .Q(g4966), .QN(n5706) );
  SDFFX1 DFF_916_Q_reg ( .D(g33065), .SI(g4966), .SE(n10225), .CLK(n10577), 
        .Q(g6227), .QN(n5568) );
  SDFFX1 DFF_917_Q_reg ( .D(g30443), .SI(g6227), .SE(n10183), .CLK(n10535), 
        .Q(g3929), .QN(n9856) );
  SDFFX1 DFF_918_Q_reg ( .D(g29291), .SI(g3929), .SE(n10183), .CLK(n10535), 
        .Q(g5503) );
  SDFFX1 DFF_919_Q_reg ( .D(g24279), .SI(g5503), .SE(n10175), .CLK(n10527), 
        .Q(test_so63), .QN(n10089) );
  SDFFX1 DFF_920_Q_reg ( .D(g30508), .SI(test_si64), .SE(n10187), .CLK(n10539), 
        .Q(g5925), .QN(n9924) );
  SDFFX1 DFF_921_Q_reg ( .D(g29232), .SI(g5925), .SE(n10198), .CLK(n10550), 
        .Q(g1124), .QN(n5692) );
  SDFFX1 DFF_922_Q_reg ( .D(g34269), .SI(g1124), .SE(n10168), .CLK(n10520), 
        .Q(g4955), .QN(n5614) );
  SDFFX1 DFF_923_Q_reg ( .D(g30464), .SI(g4955), .SE(n10253), .CLK(n10605), 
        .Q(g5224), .QN(n9812) );
  SDFFX1 DFF_924_Q_reg ( .D(g33988), .SI(g5224), .SE(n10214), .CLK(n10566), 
        .Q(g2012), .QN(n5790) );
  SDFFX1 DFF_925_Q_reg ( .D(g30522), .SI(g2012), .SE(n10242), .CLK(n10594), 
        .Q(g6203), .QN(n5574) );
  SDFFX1 DFF_926_Q_reg ( .D(g25708), .SI(g6203), .SE(n10207), .CLK(n10559), 
        .Q(g5120) );
  SDFFX1 DFF_927_Q_reg ( .D(g14662), .SI(g5120), .SE(n10207), .CLK(n10559), 
        .Q(g17674), .QN(n9883) );
  SDFFX1 DFF_928_Q_reg ( .D(g30374), .SI(g17674), .SE(n10176), .CLK(n10528), 
        .Q(g2389), .QN(n5631) );
  SDFFX1 DFF_929_Q_reg ( .D(g26953), .SI(g2389), .SE(n10188), .CLK(n10540), 
        .Q(g4438), .QN(n10051) );
  SDFFX1 DFF_930_Q_reg ( .D(g34008), .SI(g4438), .SE(n10268), .CLK(n10620), 
        .Q(g2429), .QN(n5814) );
  SDFFX1 DFF_931_Q_reg ( .D(g34444), .SI(g2429), .SE(n10204), .CLK(n10556), 
        .Q(g2787), .QN(n5610) );
  SDFFX1 DFF_932_Q_reg ( .D(g34731), .SI(g2787), .SE(n10269), .CLK(n10621), 
        .Q(test_so64) );
  SDFFX1 DFF_933_Q_reg ( .D(g33606), .SI(test_si65), .SE(n10177), .CLK(n10529), 
        .Q(g2675), .QN(n5457) );
  SDFFX1 DFF_934_Q_reg ( .D(g24334), .SI(g2675), .SE(n10224), .CLK(n10576), 
        .Q(g18881), .QN(n5541) );
  SDFFX1 DFF_935_Q_reg ( .D(g34265), .SI(g18881), .SE(n10224), .CLK(n10576), 
        .Q(g4836), .QN(n5713) );
  SDFFX1 DFF_936_Q_reg ( .D(g30340), .SI(g4836), .SE(n10185), .CLK(n10537), 
        .Q(g1199), .QN(n9776) );
  SDFFX1 DFF_937_Q_reg ( .D(g24257), .SI(g1199), .SE(n10212), .CLK(n10564), 
        .Q(g19357), .QN(n5401) );
  SDFFX1 DFF_938_Q_reg ( .D(g30482), .SI(g19357), .SE(n10180), .CLK(n10532), 
        .Q(g5547), .QN(n9798) );
  SDFFX1 DFF_941_Q_reg ( .D(g34604), .SI(g5547), .SE(n10221), .CLK(n10573), 
        .Q(g2138), .QN(n5275) );
  SDFFX1 DFF_942_Q_reg ( .D(g13926), .SI(g2138), .SE(n10222), .CLK(n10574), 
        .Q(g16744), .QN(n9892) );
  SDFFX1 DFF_943_Q_reg ( .D(g33591), .SI(g16744), .SE(n10262), .CLK(n10614), 
        .Q(g2338), .QN(n5310) );
  SDFFX1 DFF_944_Q_reg ( .D(g8918), .SI(g2338), .SE(n10262), .CLK(n10614), .Q(
        g8919) );
  SDFFX1 DFF_945_Q_reg ( .D(g30525), .SI(g8919), .SE(n10226), .CLK(n10578), 
        .Q(g6247), .QN(n10033) );
  SDFFX1 DFF_946_Q_reg ( .D(g26929), .SI(g6247), .SE(n10203), .CLK(n10555), 
        .Q(g2791), .QN(n9607) );
  SDFFX1 DFF_947_Q_reg ( .D(g30448), .SI(g2791), .SE(n10214), .CLK(n10566), 
        .Q(test_so65) );
  SDFFX1 DFF_948_Q_reg ( .D(g34602), .SI(test_si66), .SE(n10165), .CLK(n10517), 
        .Q(g1291), .QN(n2549) );
  SDFFX1 DFF_949_Q_reg ( .D(g30513), .SI(g1291), .SE(n10187), .CLK(n10539), 
        .Q(g5945), .QN(n9849) );
  SDFFX1 DFF_950_Q_reg ( .D(g30469), .SI(g5945), .SE(n10258), .CLK(n10610), 
        .Q(g5244), .QN(n9884) );
  SDFFX1 DFF_951_Q_reg ( .D(g33608), .SI(g5244), .SE(n10258), .CLK(n10610), 
        .Q(g2759), .QN(n9582) );
  SDFFX1 DFF_952_Q_reg ( .D(g33626), .SI(g2759), .SE(n10261), .CLK(n10613), 
        .Q(g6741), .QN(n5398) );
  SDFFX1 DFF_953_Q_reg ( .D(g34725), .SI(g6741), .SE(n10261), .CLK(n10613), 
        .Q(g785), .QN(n5293) );
  SDFFX1 DFF_954_Q_reg ( .D(g30342), .SI(g785), .SE(n10211), .CLK(n10563), .Q(
        g1259), .QN(n5553) );
  SDFFX1 DFF_955_Q_reg ( .D(g29267), .SI(g1259), .SE(n10173), .CLK(n10525), 
        .Q(g3484), .QN(n5668) );
  SDFFX1 DFF_956_Q_reg ( .D(g25593), .SI(g3484), .SE(n10210), .CLK(n10562), 
        .Q(g209) );
  SDFFX1 DFF_957_Q_reg ( .D(g30548), .SI(g209), .SE(n10249), .CLK(n10601), .Q(
        g6609), .QN(n9801) );
  SDFFX1 DFF_958_Q_reg ( .D(g33052), .SI(g6609), .SE(n10174), .CLK(n10526), 
        .Q(g5517), .QN(n10057) );
  SDFFX1 DFF_959_Q_reg ( .D(g34012), .SI(g5517), .SE(n10268), .CLK(n10620), 
        .Q(g2449), .QN(n5798) );
  SDFFX1 DFF_960_Q_reg ( .D(g34017), .SI(g2449), .SE(n10212), .CLK(n10564), 
        .Q(test_so66) );
  SDFFX1 DFF_961_Q_reg ( .D(g18881), .SI(test_si67), .SE(n10224), .CLK(n10576), 
        .Q(n9281) );
  SDFFX1 DFF_962_Q_reg ( .D(g24263), .SI(n9281), .SE(n10256), .CLK(n10608), 
        .Q(g2715), .QN(n5299) );
  SDFFX1 DFF_963_Q_reg ( .D(g26912), .SI(g2715), .SE(n10196), .CLK(n10548), 
        .Q(g936), .QN(n5557) );
  SDFFX1 DFF_964_Q_reg ( .D(g30364), .SI(g936), .SE(n10204), .CLK(n10556), .Q(
        g2098), .QN(n5280) );
  SDFFX1 DFF_965_Q_reg ( .D(g34254), .SI(g2098), .SE(n10195), .CLK(n10547), 
        .Q(g4462), .QN(n5671) );
  SDFFX1 DFF_966_Q_reg ( .D(g34251), .SI(g4462), .SE(n10222), .CLK(n10574), 
        .Q(g604), .QN(n5473) );
  SDFFX1 DFF_967_Q_reg ( .D(g30560), .SI(g604), .SE(n10249), .CLK(n10601), .Q(
        g6589), .QN(n9960) );
  SDFFX1 DFF_968_Q_reg ( .D(g33983), .SI(g6589), .SE(n10203), .CLK(n10555), 
        .Q(n9280), .QN(n18476) );
  SDFFX1 DFF_970_Q_reg ( .D(g13085), .SI(n9280), .SE(n10234), .CLK(n10586), 
        .Q(g17845) );
  SDFFX1 DFF_971_Q_reg ( .D(g13099), .SI(g17845), .SE(n10264), .CLK(n10616), 
        .Q(g17871) );
  SDFFX1 DFF_972_Q_reg ( .D(g24204), .SI(g17871), .SE(n10203), .CLK(n10555), 
        .Q(g429) );
  SDFFX1 DFF_973_Q_reg ( .D(g33980), .SI(g429), .SE(n10203), .CLK(n10555), .Q(
        g1870), .QN(n5813) );
  SDFFX1 DFF_974_Q_reg ( .D(g34631), .SI(g1870), .SE(n10230), .CLK(n10582), 
        .Q(test_so67) );
  SDFFX1 DFF_977_Q_reg ( .D(g29243), .SI(test_si68), .SE(n10170), .CLK(n10522), 
        .Q(g1825), .QN(n9823) );
  SDFFX1 DFF_979_Q_reg ( .D(g25623), .SI(g1825), .SE(n10251), .CLK(n10603), 
        .Q(g1008), .QN(n5321) );
  SDFFX1 DFF_980_Q_reg ( .D(g26950), .SI(g1008), .SE(n10251), .CLK(n10603), 
        .Q(g4392), .QN(n5710) );
  SDFFX1 DFF_981_Q_reg ( .D(test_so46), .SI(g4392), .SE(n10251), .CLK(n10603), 
        .Q(g8283), .QN(n9716) );
  SDFFX1 DFF_982_Q_reg ( .D(g30431), .SI(g8283), .SE(n10252), .CLK(n10604), 
        .Q(g3546), .QN(n9962) );
  SDFFX1 DFF_983_Q_reg ( .D(g30467), .SI(g3546), .SE(n10217), .CLK(n10569), 
        .Q(g5236), .QN(n9847) );
  SDFFX1 DFF_984_Q_reg ( .D(g30353), .SI(g5236), .SE(n10208), .CLK(n10560), 
        .Q(g1768), .QN(n5834) );
  SDFFX1 DFF_985_Q_reg ( .D(g34467), .SI(g1768), .SE(n10225), .CLK(n10577), 
        .Q(g4854) );
  SDFFX1 DFF_986_Q_reg ( .D(g30442), .SI(g4854), .SE(n10183), .CLK(n10535), 
        .Q(g3925), .QN(n9930) );
  SDFFX1 DFF_987_Q_reg ( .D(g29305), .SI(g3925), .SE(n10189), .CLK(n10541), 
        .Q(g6509), .QN(n9665) );
  SDFFX1 DFF_988_Q_reg ( .D(g25616), .SI(g6509), .SE(n10255), .CLK(n10607), 
        .Q(g732), .QN(n5732) );
  SDFFX1 DFF_989_Q_reg ( .D(g29252), .SI(g732), .SE(n10206), .CLK(n10558), .Q(
        g2504), .QN(n9941) );
  SDFFX1 DFF_990_Q_reg ( .D(g13272), .SI(g2504), .SE(n10212), .CLK(n10564), 
        .Q(test_so68), .QN(n10128) );
  SDFFX1 DFF_991_Q_reg ( .D(g4519), .SI(test_si69), .SE(n10174), .CLK(n10526), 
        .Q(g4520) );
  SDFFX1 DFF_992_Q_reg ( .D(g8916), .SI(g4520), .SE(n10174), .CLK(n10526), .Q(
        g8917) );
  SDFFX1 DFF_993_Q_reg ( .D(g33003), .SI(g8917), .SE(n10264), .CLK(n10616), 
        .Q(g2185), .QN(n5376) );
  SDFFX1 DFF_994_Q_reg ( .D(g34613), .SI(g2185), .SE(n10199), .CLK(n10551), 
        .Q(g37), .QN(g30327) );
  SDFFX1 DFF_995_Q_reg ( .D(g16748), .SI(g37), .SE(n10199), .CLK(n10551), .Q(
        g4031) );
  SDFFX1 DFF_996_Q_reg ( .D(g33570), .SI(g4031), .SE(n10218), .CLK(n10570), 
        .Q(g2070), .QN(n5535) );
  SDFFX1 DFF_997_Q_reg ( .D(g8132), .SI(g2070), .SE(n10234), .CLK(n10586), .Q(
        g8235), .QN(n9718) );
  SDFFX1 DFF_1000_Q_reg ( .D(g34734), .SI(g8235), .SE(n10232), .CLK(n10584), 
        .Q(g4176), .QN(n5494) );
  SDFFX1 DFF_1001_Q_reg ( .D(g24275), .SI(g4176), .SE(n10236), .CLK(n10588), 
        .Q(g11418), .QN(n5435) );
  SDFFX1 DFF_1002_Q_reg ( .D(g7243), .SI(g11418), .SE(n10236), .CLK(n10588), 
        .Q(g4405), .QN(n9569) );
  SDFFX1 DFF_1003_Q_reg ( .D(g14167), .SI(g4405), .SE(n10247), .CLK(n10599), 
        .Q(g872), .QN(n9598) );
  SDFFX1 DFF_1004_Q_reg ( .D(g29302), .SI(g872), .SE(n10179), .CLK(n10531), 
        .Q(g6181), .QN(n5667) );
  SDFFX1 DFF_1005_Q_reg ( .D(g24349), .SI(g6181), .SE(n10265), .CLK(n10617), 
        .Q(test_so69), .QN(n10130) );
  SDFFX1 DFF_1006_Q_reg ( .D(g34264), .SI(test_si70), .SE(n10179), .CLK(n10531), .Q(g4765), .QN(n5613) );
  SDFFX1 DFF_1007_Q_reg ( .D(g30484), .SI(g4765), .SE(n10175), .CLK(n10527), 
        .Q(g5563), .QN(n9928) );
  SDFFX1 DFF_1008_Q_reg ( .D(g25634), .SI(g5563), .SE(n10176), .CLK(n10528), 
        .Q(g1395), .QN(n9966) );
  SDFFX1 DFF_1009_Q_reg ( .D(g33567), .SI(g1395), .SE(n10218), .CLK(n10570), 
        .Q(g1913), .QN(n5828) );
  SDFFX1 DFF_1010_Q_reg ( .D(g33585), .SI(g1913), .SE(n10262), .CLK(n10614), 
        .Q(g2331), .QN(n5513) );
  SDFFX1 DFF_1011_Q_reg ( .D(g30527), .SI(g2331), .SE(n10266), .CLK(n10618), 
        .Q(g6263), .QN(n9808) );
  SDFFX1 DFF_1012_Q_reg ( .D(g34978), .SI(g6263), .SE(n10167), .CLK(n10519), 
        .Q(n9276) );
  SDFFX1 DFF_1013_Q_reg ( .D(g30447), .SI(n9276), .SE(n10167), .CLK(n10519), 
        .Q(g3945), .QN(n9855) );
  SDFFX1 DFF_1014_Q_reg ( .D(g7540), .SI(g3945), .SE(n10239), .CLK(n10591), 
        .Q(g347), .QN(n5860) );
  SDFFX1 DFF_1016_Q_reg ( .D(g34256), .SI(g347), .SE(n10195), .CLK(n10547), 
        .Q(g4473), .QN(n9703) );
  SDFFX1 DFF_1017_Q_reg ( .D(g25630), .SI(g4473), .SE(n10266), .CLK(n10618), 
        .Q(g1266), .QN(n9743) );
  SDFFX1 DFF_1018_Q_reg ( .D(g29290), .SI(g1266), .SE(n10182), .CLK(n10534), 
        .Q(g5489), .QN(n5660) );
  SDFFX1 DFF_1019_Q_reg ( .D(g29227), .SI(g5489), .SE(n10172), .CLK(n10524), 
        .Q(test_so70) );
  SDFFX1 DFF_1020_Q_reg ( .D(g31872), .SI(test_si71), .SE(n10257), .CLK(n10609), .Q(g2748), .QN(n5516) );
  SDFFX1 DFF_1021_Q_reg ( .D(g29287), .SI(g2748), .SE(n10169), .CLK(n10521), 
        .Q(g5471), .QN(n9627) );
  SDFFX1 DFF_1022_Q_reg ( .D(g31897), .SI(g5471), .SE(n10189), .CLK(n10541), 
        .Q(g4540) );
  SDFFX1 DFF_1023_Q_reg ( .D(g17764), .SI(g4540), .SE(n10189), .CLK(n10541), 
        .Q(g6723) );
  SDFFX1 DFF_1024_Q_reg ( .D(g30562), .SI(g6723), .SE(n10194), .CLK(n10546), 
        .Q(g6605), .QN(n10023) );
  SDFFX1 DFF_1025_Q_reg ( .D(g34011), .SI(g6605), .SE(n10215), .CLK(n10567), 
        .Q(n9274), .QN(n18477) );
  SDFFX1 DFF_1026_Q_reg ( .D(g33996), .SI(n9274), .SE(n10230), .CLK(n10582), 
        .Q(g2173) );
  SDFFX1 DFF_1027_Q_reg ( .D(g21898), .SI(g2173), .SE(n10230), .CLK(n10582), 
        .Q(g9019) );
  SDFFX1 DFF_1028_Q_reg ( .D(g33014), .SI(g9019), .SE(n10215), .CLK(n10567), 
        .Q(g2491), .QN(n5405) );
  SDFFX1 DFF_1029_Q_reg ( .D(g34465), .SI(g2491), .SE(n10215), .CLK(n10567), 
        .Q(g4849), .QN(n10063) );
  SDFFX1 DFF_1030_Q_reg ( .D(g33995), .SI(g4849), .SE(n10255), .CLK(n10607), 
        .Q(g2169), .QN(n5788) );
  SDFFX1 DFF_1031_Q_reg ( .D(g30372), .SI(g2169), .SE(n10193), .CLK(n10545), 
        .Q(n9273), .QN(n18482) );
  SDFFX1 DFF_1032_Q_reg ( .D(g30545), .SI(n9273), .SE(n10193), .CLK(n10545), 
        .Q(test_so71) );
  SDFFX1 DFF_1033_Q_reg ( .D(g30389), .SI(test_si72), .SE(n10199), .CLK(n10551), .Q(g29219), .QN(n9588) );
  SDFFX1 DFF_1034_Q_reg ( .D(g33590), .SI(g29219), .SE(n10176), .CLK(n10528), 
        .Q(g2407), .QN(n5459) );
  SDFFX1 DFF_1035_Q_reg ( .D(g34616), .SI(g2407), .SE(n10188), .CLK(n10540), 
        .Q(g2868) );
  SDFFX1 DFF_1036_Q_reg ( .D(g26927), .SI(g2868), .SE(n10220), .CLK(n10572), 
        .Q(g2767), .QN(n9610) );
  SDFFX1 DFF_1037_Q_reg ( .D(g32992), .SI(g2767), .SE(n10220), .CLK(n10572), 
        .Q(g1783), .QN(n5596) );
  SDFFX1 DFF_1038_Q_reg ( .D(g13895), .SI(g1783), .SE(n10243), .CLK(n10595), 
        .Q(g16718), .QN(n9881) );
  SDFFX1 DFF_1039_Q_reg ( .D(g25631), .SI(g16718), .SE(n10192), .CLK(n10544), 
        .Q(g1312), .QN(n5466) );
  SDFFX1 DFF_1040_Q_reg ( .D(g30477), .SI(g1312), .SE(n10264), .CLK(n10616), 
        .Q(g5212), .QN(n9977) );
  SDFFX1 DFF_1041_Q_reg ( .D(g34632), .SI(g5212), .SE(n10230), .CLK(n10582), 
        .Q(g4245) );
  SDFFX1 DFF_1042_Q_reg ( .D(g28046), .SI(g4245), .SE(n10230), .CLK(n10582), 
        .Q(g645) );
  SDFFX1 DFF_1043_Q_reg ( .D(g9019), .SI(g645), .SE(n10230), .CLK(n10582), .Q(
        g4291), .QN(n10101) );
  SDFFX1 DFF_1044_Q_reg ( .D(g26896), .SI(g4291), .SE(n10230), .CLK(n10582), 
        .Q(g29212) );
  SDFFX1 DFF_1045_Q_reg ( .D(g25602), .SI(g29212), .SE(n10230), .CLK(n10582), 
        .Q(test_so72), .QN(n10136) );
  SDFFX1 DFF_1046_Q_reg ( .D(g26916), .SI(test_si73), .SE(n10198), .CLK(n10550), .Q(g1129), .QN(n5329) );
  SDFFX1 DFF_1047_Q_reg ( .D(g33578), .SI(g1129), .SE(n10218), .CLK(n10570), 
        .Q(g2227), .QN(n5538) );
  SDFFX1 DFF_1049_Q_reg ( .D(g8787), .SI(g2227), .SE(n10206), .CLK(n10558), 
        .Q(g8788), .QN(n9766) );
  SDFFX1 DFF_1050_Q_reg ( .D(g33579), .SI(g8788), .SE(n10192), .CLK(n10544), 
        .Q(g2246), .QN(n9659) );
  SDFFX1 DFF_1051_Q_reg ( .D(g30354), .SI(g2246), .SE(n10170), .CLK(n10522), 
        .Q(g1830), .QN(n5413) );
  SDFFX1 DFF_1052_Q_reg ( .D(g30425), .SI(g1830), .SE(n10184), .CLK(n10536), 
        .Q(g3590), .QN(n9997) );
  SDFFX1 DFF_1053_Q_reg ( .D(g24200), .SI(g3590), .SE(n10171), .CLK(n10523), 
        .Q(g392), .QN(n9778) );
  SDFFX1 DFF_1054_Q_reg ( .D(g33544), .SI(g392), .SE(n10254), .CLK(n10606), 
        .Q(g1592), .QN(n5362) );
  SDFFX1 DFF_1055_Q_reg ( .D(g25764), .SI(g1592), .SE(n10228), .CLK(n10580), 
        .Q(g6505) );
  SDFFX1 DFF_1057_Q_reg ( .D(g24246), .SI(g6505), .SE(n10228), .CLK(n10580), 
        .Q(g1221), .QN(n10068) );
  SDFFX1 DFF_1058_Q_reg ( .D(g30507), .SI(g1221), .SE(n10186), .CLK(n10538), 
        .Q(g5921), .QN(n9837) );
  SDFFX1 DFF_1059_Q_reg ( .D(g26889), .SI(g5921), .SE(n10209), .CLK(n10561), 
        .Q(g29216) );
  SDFFX1 DFF_1060_Q_reg ( .D(g30333), .SI(g29216), .SE(n10209), .CLK(n10561), 
        .Q(test_so73) );
  SDFFX1 DFF_1061_Q_reg ( .D(test_so42), .SI(test_si74), .SE(n10210), .CLK(
        n10562), .Q(g218), .QN(n10050) );
  SDFFX1 DFF_1063_Q_reg ( .D(g32998), .SI(g218), .SE(n10228), .CLK(n10580), 
        .Q(g1932), .QN(n5829) );
  SDFFX1 DFF_1064_Q_reg ( .D(g32987), .SI(g1932), .SE(n10267), .CLK(n10619), 
        .Q(g1624), .QN(n5370) );
  SDFFX1 DFF_1065_Q_reg ( .D(g25702), .SI(g1624), .SE(n10207), .CLK(n10559), 
        .Q(g5062), .QN(n9755) );
  SDFFX1 DFF_1066_Q_reg ( .D(g29286), .SI(g5062), .SE(n10168), .CLK(n10520), 
        .Q(g5462), .QN(n5744) );
  SDFFX1 DFF_1067_Q_reg ( .D(g34606), .SI(g5462), .SE(n10168), .CLK(n10520), 
        .Q(g2689), .QN(n5347) );
  SDFFX1 DFF_1068_Q_reg ( .D(g33070), .SI(g2689), .SE(n10248), .CLK(n10600), 
        .Q(g6573), .QN(n5563) );
  SDFFX1 DFF_1069_Q_reg ( .D(g29240), .SI(g6573), .SE(n10192), .CLK(n10544), 
        .Q(g1677), .QN(n9828) );
  SDFFX1 DFF_1070_Q_reg ( .D(g32999), .SI(g1677), .SE(n10269), .CLK(n10621), 
        .Q(g2028), .QN(n5371) );
  SDFFX1 DFF_1071_Q_reg ( .D(g33605), .SI(g2028), .SE(n10177), .CLK(n10529), 
        .Q(g2671), .QN(n5278) );
  SDFFX1 DFF_1072_Q_reg ( .D(g24255), .SI(g2671), .SE(n10212), .CLK(n10564), 
        .Q(g10527) );
  SDFFX1 DFF_1073_Q_reg ( .D(g26945), .SI(g10527), .SE(n10252), .CLK(n10604), 
        .Q(g7243) );
  SDFFX1 DFF_1074_Q_reg ( .D(n10104), .SI(g7243), .SE(n10197), .CLK(n10549), 
        .Q(test_so74) );
  SDFFX1 DFF_1075_Q_reg ( .D(g33558), .SI(test_si75), .SE(n10170), .CLK(n10522), .Q(g1848), .QN(n5464) );
  SDFFX1 DFF_1078_Q_reg ( .D(g25699), .SI(g1848), .SE(n10165), .CLK(n10517), 
        .Q(g29213), .QN(n5669) );
  SDFFX1 DFF_1079_Q_reg ( .D(g29289), .SI(g29213), .SE(n10165), .CLK(n10517), 
        .Q(g5485), .QN(n5869) );
  SDFFX1 DFF_1080_Q_reg ( .D(g30388), .SI(g5485), .SE(n10257), .CLK(n10609), 
        .Q(g2741), .QN(n5349) );
  SDFFX1 DFF_1081_Q_reg ( .D(g12184), .SI(g2741), .SE(n10191), .CLK(n10543), 
        .Q(g11678), .QN(n5482) );
  SDFFX1 DFF_1082_Q_reg ( .D(g29254), .SI(g11678), .SE(n10201), .CLK(n10553), 
        .Q(g2638), .QN(n9832) );
  SDFFX1 DFF_1083_Q_reg ( .D(g28074), .SI(g2638), .SE(n10246), .CLK(n10598), 
        .Q(g4122) );
  SDFFX1 DFF_1084_Q_reg ( .D(g34450), .SI(g4122), .SE(n10261), .CLK(n10613), 
        .Q(g4322), .QN(n5506) );
  SDFFX1 DFF_1085_Q_reg ( .D(g30512), .SI(g4322), .SE(n10187), .CLK(n10539), 
        .Q(g5941), .QN(n9978) );
  SDFFX1 DFF_1086_Q_reg ( .D(g33572), .SI(g5941), .SE(n10204), .CLK(n10556), 
        .Q(g2108), .QN(n5452) );
  SDFFX1 DFF_1087_Q_reg ( .D(g17646), .SI(g2108), .SE(n10204), .CLK(n10556), 
        .Q(g13068) );
  SDFFX1 DFF_1088_Q_reg ( .D(g25), .SI(g13068), .SE(n10204), .CLK(n10556), .Q(
        g25) );
  SDFFX1 DFF_1089_Q_reg ( .D(g33551), .SI(g25), .SE(n10254), .CLK(n10606), .Q(
        test_so75), .QN(n10134) );
  SDFFX1 DFF_1090_Q_reg ( .D(g33538), .SI(test_si76), .SE(n10222), .CLK(n10574), .Q(g595), .QN(n5476) );
  SDFFX1 DFF_1091_Q_reg ( .D(g33005), .SI(g595), .SE(n10209), .CLK(n10561), 
        .Q(g2217), .QN(n5512) );
  SDFFX1 DFF_1092_Q_reg ( .D(g24248), .SI(g2217), .SE(n10176), .CLK(n10528), 
        .Q(n9267), .QN(DFF_1092_n1) );
  SDFFX1 DFF_1093_Q_reg ( .D(g33002), .SI(n9267), .SE(n10204), .CLK(n10556), 
        .Q(g2066), .QN(n5832) );
  SDFFX1 DFF_1094_Q_reg ( .D(g24234), .SI(g2066), .SE(n10229), .CLK(n10581), 
        .Q(g1152), .QN(n5618) );
  SDFFX1 DFF_1095_Q_reg ( .D(g30471), .SI(g1152), .SE(n10217), .CLK(n10569), 
        .Q(g5252), .QN(n9846) );
  SDFFX1 DFF_1096_Q_reg ( .D(g34000), .SI(g5252), .SE(n10237), .CLK(n10589), 
        .Q(g2165), .QN(n9652) );
  SDFFX1 DFF_1097_Q_reg ( .D(g34016), .SI(g2165), .SE(n10249), .CLK(n10601), 
        .Q(g2571), .QN(n5787) );
  SDFFX1 DFF_1098_Q_reg ( .D(g33048), .SI(g2571), .SE(n10250), .CLK(n10602), 
        .Q(g5176), .QN(n5650) );
  SDFFX1 DFF_1100_Q_reg ( .D(g8283), .SI(g5176), .SE(n10251), .CLK(n10603), 
        .Q(g8403), .QN(n9717) );
  SDFFX1 DFF_1102_Q_reg ( .D(g17819), .SI(g8403), .SE(n10251), .CLK(n10603), 
        .Q(g14673), .QN(n5581) );
  SDFFX1 DFF_1103_Q_reg ( .D(g25628), .SI(g14673), .SE(n10228), .CLK(n10580), 
        .Q(test_so76) );
  SDFFX1 DFF_1104_Q_reg ( .D(g26934), .SI(test_si77), .SE(n10213), .CLK(n10565), .Q(g2827), .QN(n9609) );
  SDFFX1 DFF_1106_Q_reg ( .D(g14201), .SI(g2827), .SE(n10247), .CLK(n10599), 
        .Q(g14217), .QN(n9595) );
  SDFFX1 DFF_1107_Q_reg ( .D(g34468), .SI(g14217), .SE(n10216), .CLK(n10568), 
        .Q(g4859), .QN(n9586) );
  SDFFX1 DFF_1108_Q_reg ( .D(g24202), .SI(g4859), .SE(n10171), .CLK(n10523), 
        .Q(g424), .QN(n9746) );
  SDFFX1 DFF_1109_Q_reg ( .D(g33542), .SI(g424), .SE(n10211), .CLK(n10563), 
        .Q(g1274), .QN(n5730) );
  SDFFX1 DFF_1110_Q_reg ( .D(g17404), .SI(g1274), .SE(n10212), .CLK(n10564), 
        .Q(g17423), .QN(n9735) );
  SDFFX1 DFF_1111_Q_reg ( .D(g33435), .SI(g17423), .SE(n10208), .CLK(n10560), 
        .Q(n9265) );
  SDFFX1 DFF_1112_Q_reg ( .D(g34445), .SI(n9265), .SE(n10208), .CLK(n10560), 
        .Q(g2803), .QN(n5545) );
  SDFFX1 DFF_1114_Q_reg ( .D(g33555), .SI(g2803), .SE(n10267), .CLK(n10619), 
        .Q(g1821), .QN(n9654) );
  SDFFX1 DFF_1115_Q_reg ( .D(g34013), .SI(g1821), .SE(n10211), .CLK(n10563), 
        .Q(g2509), .QN(n9692) );
  SDFFX1 DFF_1116_Q_reg ( .D(g28091), .SI(g2509), .SE(n10211), .CLK(n10563), 
        .Q(g5073), .QN(n9689) );
  SDFFX1 DFF_1117_Q_reg ( .D(g26919), .SI(g5073), .SE(n10211), .CLK(n10563), 
        .Q(test_so77), .QN(n5556) );
  SDFFX1 DFF_1118_Q_reg ( .D(g8235), .SI(test_si78), .SE(n10234), .CLK(n10586), 
        .Q(g8353), .QN(n9719) );
  SDFFX1 DFF_1119_Q_reg ( .D(g17685), .SI(g8353), .SE(n10234), .CLK(n10586), 
        .Q(g13085), .QN(n10032) );
  SDFFX1 DFF_1120_Q_reg ( .D(g30554), .SI(g13085), .SE(n10194), .CLK(n10546), 
        .Q(g6633), .QN(n9992) );
  SDFFX1 DFF_1121_Q_reg ( .D(g29281), .SI(g6633), .SE(n10178), .CLK(n10530), 
        .Q(g5124), .QN(n9616) );
  SDFFX1 DFF_1122_Q_reg ( .D(test_so44), .SI(g5124), .SE(n10240), .CLK(n10592), 
        .Q(g17400), .QN(n9724) );
  SDFFX1 DFF_1123_Q_reg ( .D(g30537), .SI(g17400), .SE(n10225), .CLK(n10577), 
        .Q(g6303), .QN(n10004) );
  SDFFX1 DFF_1124_Q_reg ( .D(g28092), .SI(g6303), .SE(n10165), .CLK(n10517), 
        .Q(g5069), .QN(n9688) );
  SDFFX1 DFF_1125_Q_reg ( .D(g34732), .SI(g5069), .SE(n10188), .CLK(n10540), 
        .Q(g2994), .QN(n5634) );
  SDFFX1 DFF_1126_Q_reg ( .D(g28049), .SI(g2994), .SE(n10237), .CLK(n10589), 
        .Q(g650), .QN(n9774) );
  SDFFX1 DFF_1127_Q_reg ( .D(g33545), .SI(g650), .SE(n10254), .CLK(n10606), 
        .Q(g1636), .QN(n5549) );
  SDFFX1 DFF_1128_Q_reg ( .D(g30441), .SI(g1636), .SE(n10215), .CLK(n10567), 
        .Q(g3921), .QN(n9839) );
  SDFFX1 DFF_1129_Q_reg ( .D(g29247), .SI(g3921), .SE(n10204), .CLK(n10556), 
        .Q(test_so78) );
  SDFFX1 DFF_1130_Q_reg ( .D(g24354), .SI(test_si79), .SE(n10196), .CLK(n10548), .Q(g6732), .QN(n10037) );
  SDFFX1 DFF_1131_Q_reg ( .D(g25636), .SI(g6732), .SE(n10229), .CLK(n10581), 
        .Q(g1306), .QN(n5796) );
  SDFFX1 DFF_1133_Q_reg ( .D(g26914), .SI(g1306), .SE(n10232), .CLK(n10584), 
        .Q(g1061), .QN(n9754) );
  SDFFX1 DFF_1134_Q_reg ( .D(g25670), .SI(g1061), .SE(n10241), .CLK(n10593), 
        .Q(g3462) );
  SDFFX1 DFF_1135_Q_reg ( .D(g33998), .SI(g3462), .SE(n10255), .CLK(n10607), 
        .Q(g2181), .QN(n5803) );
  SDFFX1 DFF_1136_Q_reg ( .D(g25626), .SI(g2181), .SE(n10213), .CLK(n10565), 
        .Q(g956), .QN(n5341) );
  SDFFX1 DFF_1137_Q_reg ( .D(g33977), .SI(g956), .SE(n10228), .CLK(n10580), 
        .Q(g1756), .QN(n5804) );
  SDFFX1 DFF_1138_Q_reg ( .D(g29297), .SI(g1756), .SE(n10245), .CLK(n10597), 
        .Q(g5849) );
  SDFFX1 DFF_1139_Q_reg ( .D(g28071), .SI(g5849), .SE(n10246), .CLK(n10598), 
        .Q(g4112), .QN(n10035) );
  SDFFX1 DFF_1140_Q_reg ( .D(g30387), .SI(g4112), .SE(n10177), .CLK(n10529), 
        .Q(n9262), .QN(n18484) );
  SDFFX1 DFF_1141_Q_reg ( .D(g33577), .SI(n9262), .SE(n10177), .CLK(n10529), 
        .Q(g2197), .QN(n5514) );
  SDFFX1 DFF_1143_Q_reg ( .D(g33592), .SI(g2197), .SE(n10268), .CLK(n10620), 
        .Q(test_so79), .QN(n10131) );
  SDFFX1 DFF_1144_Q_reg ( .D(g26913), .SI(test_si80), .SE(n10253), .CLK(n10605), .Q(g1046), .QN(n9910) );
  SDFFX1 DFF_1145_Q_reg ( .D(g28044), .SI(g1046), .SE(n10238), .CLK(n10590), 
        .Q(g482), .QN(n5820) );
  SDFFX1 DFF_1146_Q_reg ( .D(g26948), .SI(g482), .SE(n10236), .CLK(n10588), 
        .Q(g4401) );
  SDFFX1 DFF_1148_Q_reg ( .D(g30344), .SI(g4401), .SE(n10236), .CLK(n10588), 
        .Q(g1514), .QN(n5364) );
  SDFFX1 DFF_1149_Q_reg ( .D(g26885), .SI(g1514), .SE(n10236), .CLK(n10588), 
        .Q(g329), .QN(n5766) );
  SDFFX1 DFF_1150_Q_reg ( .D(g33069), .SI(g329), .SE(n10248), .CLK(n10600), 
        .Q(g6565), .QN(n5386) );
  SDFFX1 DFF_1151_Q_reg ( .D(g34621), .SI(g6565), .SE(n10192), .CLK(n10544), 
        .Q(g2950), .QN(n10082) );
  SDFFX1 DFF_1153_Q_reg ( .D(g28059), .SI(g2950), .SE(n10192), .CLK(n10544), 
        .Q(g1345), .QN(n9750) );
  SDFFX1 DFF_1154_Q_reg ( .D(g25762), .SI(g1345), .SE(n10189), .CLK(n10541), 
        .Q(g6533), .QN(n5445) );
  SDFFX1 DFF_1155_Q_reg ( .D(g16624), .SI(g6533), .SE(n10189), .CLK(n10541), 
        .Q(g14421) );
  SDFFX1 DFF_1157_Q_reg ( .D(g34633), .SI(g14421), .SE(n10190), .CLK(n10542), 
        .Q(g4727), .QN(n5312) );
  SDFFX1 DFF_1158_Q_reg ( .D(g24352), .SI(g4727), .SE(n10265), .CLK(n10617), 
        .Q(test_so80) );
  SDFFX1 DFF_1159_Q_reg ( .D(g26925), .SI(test_si81), .SE(n10227), .CLK(n10579), .Q(g1536) );
  SDFFX1 DFF_1160_Q_reg ( .D(g30446), .SI(g1536), .SE(n10183), .CLK(n10535), 
        .Q(g3941), .QN(n9987) );
  SDFFX1 DFF_1161_Q_reg ( .D(g25597), .SI(g3941), .SE(n10237), .CLK(n10589), 
        .Q(g370), .QN(n9787) );
  SDFFX1 DFF_1162_Q_reg ( .D(g24342), .SI(g370), .SE(n10265), .CLK(n10617), 
        .Q(g5694), .QN(n9904) );
  SDFFX1 DFF_1163_Q_reg ( .D(g30357), .SI(g5694), .SE(n10171), .CLK(n10523), 
        .Q(g1858), .QN(n5892) );
  SDFFX1 DFF_1164_Q_reg ( .D(g26908), .SI(g1858), .SE(n10171), .CLK(n10523), 
        .Q(g446) );
  SDFFX1 DFF_1166_Q_reg ( .D(g30399), .SI(g446), .SE(n10231), .CLK(n10583), 
        .Q(g3219), .QN(n9836) );
  SDFFX1 DFF_1167_Q_reg ( .D(g29242), .SI(g3219), .SE(n10170), .CLK(n10522), 
        .Q(g1811), .QN(n9824) );
  SDFFX1 DFF_1169_Q_reg ( .D(g30547), .SI(g1811), .SE(n10194), .CLK(n10546), 
        .Q(g6601), .QN(n9934) );
  SDFFX1 DFF_1171_Q_reg ( .D(g34010), .SI(g6601), .SE(n10215), .CLK(n10567), 
        .Q(g2441) );
  SDFFX1 DFF_1172_Q_reg ( .D(g33986), .SI(g2441), .SE(n10198), .CLK(n10550), 
        .Q(g1874), .QN(n9633) );
  SDFFX1 DFF_1173_Q_reg ( .D(g34257), .SI(g1874), .SE(n10224), .CLK(n10576), 
        .Q(test_so81), .QN(n10132) );
  SDFFX1 DFF_1174_Q_reg ( .D(g30544), .SI(test_si82), .SE(n10249), .CLK(n10601), .Q(g6581), .QN(n9961) );
  SDFFX1 DFF_1175_Q_reg ( .D(g30561), .SI(g6581), .SE(n10193), .CLK(n10545), 
        .Q(g6597), .QN(n9996) );
  SDFFX1 DFF_1176_Q_reg ( .D(g8403), .SI(g6597), .SE(n10251), .CLK(n10603), 
        .Q(g5008), .QN(n5637) );
  SDFFX1 DFF_1177_Q_reg ( .D(g30430), .SI(g5008), .SE(n10251), .CLK(n10603), 
        .Q(g3610) );
  SDFFX1 DFF_1178_Q_reg ( .D(g34799), .SI(g3610), .SE(n10251), .CLK(n10603), 
        .Q(g2890), .QN(n10090) );
  SDFFX1 DFF_1179_Q_reg ( .D(g33565), .SI(g2890), .SE(n10169), .CLK(n10521), 
        .Q(g1978), .QN(n5845) );
  SDFFX1 DFF_1180_Q_reg ( .D(g33968), .SI(g1978), .SE(n10219), .CLK(n10571), 
        .Q(g1612) );
  SDFFX1 DFF_1181_Q_reg ( .D(g34843), .SI(g1612), .SE(n10218), .CLK(n10570), 
        .Q(g112), .QN(n9779) );
  SDFFX1 DFF_1182_Q_reg ( .D(g34793), .SI(g112), .SE(n10166), .CLK(n10518), 
        .Q(g2856), .QN(n9585) );
  SDFFX1 DFF_1184_Q_reg ( .D(g33566), .SI(g2856), .SE(n10169), .CLK(n10521), 
        .Q(g1982), .QN(n5462) );
  SDFFX1 DFF_1185_Q_reg ( .D(g17688), .SI(g1982), .SE(n10258), .CLK(n10610), 
        .Q(g17722), .QN(n9995) );
  SDFFX1 DFF_1186_Q_reg ( .D(g30465), .SI(g17722), .SE(n10258), .CLK(n10610), 
        .Q(test_so82) );
  SDFFX1 DFF_1187_Q_reg ( .D(g28073), .SI(test_si83), .SE(n10246), .CLK(n10598), .Q(g4119) );
  SDFFX1 DFF_1188_Q_reg ( .D(g24351), .SI(g4119), .SE(n10220), .CLK(n10572), 
        .Q(g6390), .QN(n9898) );
  SDFFX1 DFF_1189_Q_reg ( .D(g30346), .SI(g6390), .SE(n10227), .CLK(n10579), 
        .Q(g1542), .QN(n9775) );
  SDFFX1 DFF_1190_Q_reg ( .D(g21893), .SI(g1542), .SE(n10227), .CLK(n10579), 
        .Q(g4258), .QN(n9614) );
  SDFFX1 DFF_1191_Q_reg ( .D(g8353), .SI(g4258), .SE(n10234), .CLK(n10586), 
        .Q(g4818) );
  SDFFX1 DFF_1192_Q_reg ( .D(g31904), .SI(g4818), .SE(n10202), .CLK(n10554), 
        .Q(g5033), .QN(n9752) );
  SDFFX1 DFF_1193_Q_reg ( .D(g34635), .SI(g5033), .SE(n10234), .CLK(n10586), 
        .Q(g4717), .QN(n5344) );
  SDFFX1 DFF_1194_Q_reg ( .D(g25637), .SI(g4717), .SE(n10258), .CLK(n10610), 
        .Q(g1554), .QN(n5768) );
  SDFFX1 DFF_1195_Q_reg ( .D(g29274), .SI(g1554), .SE(n10258), .CLK(n10610), 
        .Q(g3849) );
  SDFFX1 DFF_1196_Q_reg ( .D(g14828), .SI(g3849), .SE(n10258), .CLK(n10610), 
        .Q(g17778), .QN(n9890) );
  SDFFX1 DFF_1197_Q_reg ( .D(g30396), .SI(g17778), .SE(n10231), .CLK(n10583), 
        .Q(g3199), .QN(n10009) );
  SDFFX1 DFF_1198_Q_reg ( .D(g25735), .SI(g3199), .SE(n10270), .CLK(n10622), 
        .Q(test_so83) );
  SDFFX1 DFF_1199_Q_reg ( .D(g34037), .SI(test_si84), .SE(n10205), .CLK(n10557), .Q(g4975), .QN(n5360) );
  SDFFX1 DFF_1200_Q_reg ( .D(g34791), .SI(g4975), .SE(n10261), .CLK(n10613), 
        .Q(g790), .QN(n5292) );
  SDFFX1 DFF_1201_Q_reg ( .D(g30520), .SI(g790), .SE(n10187), .CLK(n10539), 
        .Q(g5913), .QN(n10011) );
  SDFFX1 DFF_1202_Q_reg ( .D(g30358), .SI(g5913), .SE(n10203), .CLK(n10555), 
        .Q(g1902), .QN(n5837) );
  SDFFX1 DFF_1203_Q_reg ( .D(g29299), .SI(g1902), .SE(n10179), .CLK(n10531), 
        .Q(g6163), .QN(n9645) );
  SDFFX1 DFF_1204_Q_reg ( .D(g25690), .SI(g6163), .SE(n10189), .CLK(n10541), 
        .Q(g4125), .QN(n10034) );
  SDFFX1 DFF_1205_Q_reg ( .D(g28096), .SI(g4125), .SE(n10174), .CLK(n10526), 
        .Q(g4821) );
  SDFFX1 DFF_1206_Q_reg ( .D(g28088), .SI(g4821), .SE(n10205), .CLK(n10557), 
        .Q(g4939) );
  SDFFX1 DFF_1207_Q_reg ( .D(g24241), .SI(g4939), .SE(n10253), .CLK(n10605), 
        .Q(g19334), .QN(n5392) );
  SDFFX1 DFF_1208_Q_reg ( .D(g30397), .SI(g19334), .SE(n10231), .CLK(n10583), 
        .Q(g3207), .QN(n9919) );
  SDFFX1 DFF_1209_Q_reg ( .D(g4520), .SI(g3207), .SE(n10232), .CLK(n10584), 
        .Q(g4483) );
  SDFFX1 DFF_1210_Q_reg ( .D(g30409), .SI(g4483), .SE(n10232), .CLK(n10584), 
        .Q(test_so84) );
  SDFFX1 DFF_1211_Q_reg ( .D(g29284), .SI(test_si85), .SE(n10178), .CLK(n10530), .Q(g5142), .QN(n5658) );
  SDFFX1 DFF_1212_Q_reg ( .D(g30470), .SI(g5142), .SE(n10216), .CLK(n10568), 
        .Q(g5248), .QN(n9973) );
  SDFFX1 DFF_1213_Q_reg ( .D(g30367), .SI(g5248), .SE(n10168), .CLK(n10520), 
        .Q(g2126), .QN(n5891) );
  SDFFX1 DFF_1214_Q_reg ( .D(g24273), .SI(g2126), .SE(n10168), .CLK(n10520), 
        .Q(g3694), .QN(n9902) );
  SDFFX1 DFF_1215_Q_reg ( .D(g29288), .SI(g3694), .SE(n10169), .CLK(n10521), 
        .Q(g5481), .QN(n5805) );
  SDFFX1 DFF_1216_Q_reg ( .D(g30359), .SI(g5481), .SE(n10169), .CLK(n10521), 
        .Q(g1964), .QN(n5315) );
  SDFFX1 DFF_1217_Q_reg ( .D(g25698), .SI(g1964), .SE(n10165), .CLK(n10517), 
        .Q(g5097), .QN(n5753) );
  SDFFX1 DFF_1218_Q_reg ( .D(g30398), .SI(g5097), .SE(n10257), .CLK(n10609), 
        .Q(g3215), .QN(n9793) );
  SDFFX1 DFF_1219_Q_reg ( .D(g13906), .SI(g3215), .SE(n10259), .CLK(n10611), 
        .Q(g16748) );
  SDFFX1 DFF_1220_Q_reg ( .D(g33079), .SI(g16748), .SE(n10267), .CLK(n10619), 
        .Q(n9255) );
  SDFFX1 DFF_1221_Q_reg ( .D(g26952), .SI(n9255), .SE(n10172), .CLK(n10524), 
        .Q(g4427), .QN(n9769) );
  SDFFX1 DFF_1222_Q_reg ( .D(g34974), .SI(g4427), .SE(n10270), .CLK(n10622), 
        .Q(test_so85) );
  SDFFX1 DFF_1223_Q_reg ( .D(g26928), .SI(test_si86), .SE(n10208), .CLK(n10560), .Q(g2779), .QN(n9604) );
  SDFFX1 DFF_1224_Q_reg ( .D(test_so39), .SI(g2779), .SE(n10235), .CLK(n10587), 
        .Q(g8786), .QN(n5694) );
  SDFFX1 DFF_1225_Q_reg ( .D(g26954), .SI(g8786), .SE(n10257), .CLK(n10609), 
        .Q(g7245) );
  SDFFX1 DFF_1226_Q_reg ( .D(g30351), .SI(g7245), .SE(n10202), .CLK(n10554), 
        .Q(g1720), .QN(n5780) );
  SDFFX1 DFF_1227_Q_reg ( .D(g31871), .SI(g1720), .SE(n10202), .CLK(n10554), 
        .Q(g1367), .QN(n9727) );
  SDFFX1 DFF_1228_Q_reg ( .D(g9553), .SI(g1367), .SE(n10202), .CLK(n10554), 
        .Q(g5112) );
  SDFFX1 DFF_1229_Q_reg ( .D(g34978), .SI(g5112), .SE(n10202), .CLK(n10554), 
        .Q(g19), .QN(n9583) );
  SDFFX1 DFF_1230_Q_reg ( .D(g26939), .SI(g19), .SE(n10246), .CLK(n10598), .Q(
        g4145), .QN(n10072) );
  SDFFX1 DFF_1231_Q_reg ( .D(g33994), .SI(g4145), .SE(n10237), .CLK(n10589), 
        .Q(g2161), .QN(n5812) );
  SDFFX1 DFF_1232_Q_reg ( .D(g25596), .SI(g2161), .SE(n10237), .CLK(n10589), 
        .Q(g376), .QN(n5633) );
  SDFFX1 DFF_1233_Q_reg ( .D(g33586), .SI(g376), .SE(n10262), .CLK(n10614), 
        .Q(g2361), .QN(n5537) );
  SDFFX1 DFF_1234_Q_reg ( .D(g21901), .SI(g2361), .SE(n10206), .CLK(n10558), 
        .Q(test_so86), .QN(DFF_1234_n1) );
  SDFFX1 DFF_1235_Q_reg ( .D(g31866), .SI(test_si87), .SE(n10222), .CLK(n10574), .Q(g582), .QN(n5552) );
  SDFFX1 DFF_1236_Q_reg ( .D(g33000), .SI(g582), .SE(n10269), .CLK(n10621), 
        .Q(g2051), .QN(n10041) );
  SDFFX1 DFF_1237_Q_reg ( .D(g26918), .SI(g2051), .SE(n10185), .CLK(n10537), 
        .Q(g1193) );
  SDFFX1 DFF_1240_Q_reg ( .D(g30373), .SI(g1193), .SE(n10267), .CLK(n10619), 
        .Q(g2327), .QN(n5841) );
  SDFFX1 DFF_1241_Q_reg ( .D(g28056), .SI(g2327), .SE(n10196), .CLK(n10548), 
        .Q(g907), .QN(n5555) );
  SDFFX1 DFF_1242_Q_reg ( .D(g34601), .SI(g907), .SE(n10196), .CLK(n10548), 
        .Q(g947), .QN(n5286) );
  SDFFX1 DFF_1243_Q_reg ( .D(g30355), .SI(g947), .SE(n10170), .CLK(n10522), 
        .Q(g1834), .QN(n5665) );
  SDFFX1 DFF_1244_Q_reg ( .D(g30426), .SI(g1834), .SE(n10241), .CLK(n10593), 
        .Q(g3594), .QN(n9861) );
  SDFFX1 DFF_1245_Q_reg ( .D(g34805), .SI(g3594), .SE(n10188), .CLK(n10540), 
        .Q(g2999), .QN(n10092) );
  SDFFX1 DFF_1247_Q_reg ( .D(g34002), .SI(g2999), .SE(n10263), .CLK(n10615), 
        .Q(g2303), .QN(n5794) );
  SDFFX1 DFF_1248_Q_reg ( .D(g17778), .SI(g2303), .SE(n10258), .CLK(n10610), 
        .Q(g17688), .QN(n9876) );
  SDFFX1 DFF_1250_Q_reg ( .D(g28053), .SI(g17688), .SE(n10172), .CLK(n10524), 
        .Q(test_so87), .QN(n10145) );
  SDFFX1 DFF_1251_Q_reg ( .D(g29229), .SI(test_si88), .SE(n10270), .CLK(n10622), .Q(g723), .QN(n5826) );
  SDFFX1 DFF_1252_Q_reg ( .D(g33620), .SI(g723), .SE(n10182), .CLK(n10534), 
        .Q(g5703), .QN(n5397) );
  SDFFX1 DFF_1253_Q_reg ( .D(g34722), .SI(g5703), .SE(n10210), .CLK(n10562), 
        .Q(g546), .QN(n5492) );
  SDFFX1 DFF_1254_Q_reg ( .D(g33599), .SI(g546), .SE(n10211), .CLK(n10563), 
        .Q(g2472), .QN(n5619) );
  SDFFX1 DFF_1255_Q_reg ( .D(g30515), .SI(g2472), .SE(n10187), .CLK(n10539), 
        .Q(g5953), .QN(n9871) );
  SDFFX1 DFF_1256_Q_reg ( .D(g25649), .SI(g5953), .SE(n10170), .CLK(n10522), 
        .Q(g8277) );
  SDFFX1 DFF_1258_Q_reg ( .D(g33979), .SI(g8277), .SE(n10170), .CLK(n10522), 
        .Q(g1740), .QN(n9704) );
  SDFFX1 DFF_1259_Q_reg ( .D(g30417), .SI(g1740), .SE(n10184), .CLK(n10536), 
        .Q(g3550), .QN(n10029) );
  SDFFX1 DFF_1260_Q_reg ( .D(g25683), .SI(g3550), .SE(n10167), .CLK(n10519), 
        .Q(g3845), .QN(n5886) );
  SDFFX1 DFF_1261_Q_reg ( .D(g33574), .SI(g3845), .SE(n10167), .CLK(n10519), 
        .Q(g2116), .QN(n5463) );
  SDFFX1 DFF_1262_Q_reg ( .D(g17813), .SI(g2116), .SE(n10233), .CLK(n10585), 
        .Q(g14635), .QN(n5582) );
  SDFFX1 DFF_1263_Q_reg ( .D(g30410), .SI(g14635), .SE(n10265), .CLK(n10617), 
        .Q(test_so88) );
  SDFFX1 DFF_1264_Q_reg ( .D(g30454), .SI(test_si89), .SE(n10183), .CLK(n10535), .Q(g3913) );
  SDFFX1 DFF_1265_Q_reg ( .D(g34024), .SI(g3913), .SE(n10188), .CLK(n10540), 
        .Q(g10306) );
  SDFFX1 DFF_1266_Q_reg ( .D(g33547), .SI(g10306), .SE(n10166), .CLK(n10518), 
        .Q(g1687), .QN(n9658) );
  SDFFX1 DFF_1267_Q_reg ( .D(g30386), .SI(g1687), .SE(n10177), .CLK(n10529), 
        .Q(g2681), .QN(n5777) );
  SDFFX1 DFF_1268_Q_reg ( .D(g33596), .SI(g2681), .SE(n10206), .CLK(n10558), 
        .Q(g2533), .QN(n5761) );
  SDFFX1 DFF_1269_Q_reg ( .D(g26887), .SI(g2533), .SE(n10238), .CLK(n10590), 
        .Q(g324), .QN(n5827) );
  SDFFX1 DFF_1270_Q_reg ( .D(g34607), .SI(g324), .SE(n10238), .CLK(n10590), 
        .Q(g2697), .QN(n5308) );
  SDFFX1 DFF_1272_Q_reg ( .D(g31895), .SI(g2697), .SE(n10238), .CLK(n10590), 
        .Q(g4417), .QN(n9573) );
  SDFFX1 DFF_1273_Q_reg ( .D(g33068), .SI(g4417), .SE(n10238), .CLK(n10590), 
        .Q(g6561), .QN(n5646) );
  SDFFX1 DFF_1274_Q_reg ( .D(g29233), .SI(g6561), .SE(n10229), .CLK(n10581), 
        .Q(g1141), .QN(n5691) );
  SDFFX1 DFF_1275_Q_reg ( .D(g24258), .SI(g1141), .SE(n10229), .CLK(n10581), 
        .Q(g12923), .QN(n5655) );
  SDFFX1 DFF_1276_Q_reg ( .D(g30376), .SI(g12923), .SE(n10176), .CLK(n10528), 
        .Q(test_so89), .QN(n10143) );
  SDFFX1 DFF_1277_Q_reg ( .D(g33549), .SI(test_si90), .SE(n10221), .CLK(n10573), .Q(g1710), .QN(n5412) );
  SDFFX1 DFF_1278_Q_reg ( .D(g29308), .SI(g1710), .SE(n10189), .CLK(n10541), 
        .Q(g6527), .QN(n5659) );
  SDFFX1 DFF_1280_Q_reg ( .D(g30408), .SI(g6527), .SE(n10231), .CLK(n10583), 
        .Q(g3255), .QN(n9970) );
  SDFFX1 DFF_1281_Q_reg ( .D(g29241), .SI(g3255), .SE(n10192), .CLK(n10544), 
        .Q(g1691), .QN(n9827) );
  SDFFX1 DFF_1282_Q_reg ( .D(g34620), .SI(g1691), .SE(n10192), .CLK(n10544), 
        .Q(g2936), .QN(n10083) );
  SDFFX1 DFF_1283_Q_reg ( .D(g33621), .SI(g2936), .SE(n10168), .CLK(n10520), 
        .Q(g5644), .QN(n5593) );
  SDFFX1 DFF_1284_Q_reg ( .D(g25707), .SI(g5644), .SE(n10178), .CLK(n10530), 
        .Q(g5152), .QN(n5883) );
  SDFFX1 DFF_1285_Q_reg ( .D(g24339), .SI(g5152), .SE(n10178), .CLK(n10530), 
        .Q(g5352), .QN(n10038) );
  SDFFX1 DFF_1286_Q_reg ( .D(g11770), .SI(g5352), .SE(n10216), .CLK(n10568), 
        .Q(g8915) );
  SDFFX1 DFF_1288_Q_reg ( .D(g34443), .SI(g8915), .SE(n10208), .CLK(n10560), 
        .Q(g2775), .QN(n5378) );
  SDFFX1 DFF_1289_Q_reg ( .D(g34619), .SI(g2775), .SE(n10198), .CLK(n10550), 
        .Q(g2922), .QN(n10081) );
  SDFFX1 DFF_1290_Q_reg ( .D(g29234), .SI(g2922), .SE(n10198), .CLK(n10550), 
        .Q(test_so90), .QN(n10148) );
  SDFFX1 DFF_1291_Q_reg ( .D(g30503), .SI(test_si91), .SE(n10186), .CLK(n10538), .Q(g5893), .QN(n9815) );
  SDFFX1 DFF_1293_Q_reg ( .D(g16718), .SI(g5893), .SE(n10243), .CLK(n10595), 
        .Q(g16603), .QN(n9866) );
  SDFFX1 DFF_1294_Q_reg ( .D(g30550), .SI(g16603), .SE(n10194), .CLK(n10546), 
        .Q(g6617), .QN(n9933) );
  SDFFX1 DFF_1295_Q_reg ( .D(g33001), .SI(g6617), .SE(n10204), .CLK(n10556), 
        .Q(g2060), .QN(n5507) );
  SDFFX1 DFF_1296_Q_reg ( .D(g33040), .SI(g2060), .SE(n10245), .CLK(n10597), 
        .Q(g4512), .QN(n9768) );
  SDFFX1 DFF_1297_Q_reg ( .D(g30492), .SI(g4512), .SE(n10174), .CLK(n10526), 
        .Q(g5599), .QN(n9852) );
  SDFFX1 DFF_1298_Q_reg ( .D(g25664), .SI(g5599), .SE(n10268), .CLK(n10620), 
        .Q(g3401) );
  SDFFX1 DFF_1299_Q_reg ( .D(g26944), .SI(g3401), .SE(n10173), .CLK(n10525), 
        .Q(g4366) );
  SDFFX1 DFF_1300_Q_reg ( .D(test_so26), .SI(g4366), .SE(n10250), .CLK(n10602), 
        .Q(g16722) );
  SDFFX1 DFF_1301_Q_reg ( .D(g34614), .SI(g16722), .SE(n10250), .CLK(n10602), 
        .Q(g29214) );
  SDFFX1 DFF_1302_Q_reg ( .D(g29260), .SI(g29214), .SE(n10190), .CLK(n10542), 
        .Q(g3129) );
  SDFFX1 DFF_1303_Q_reg ( .D(g16686), .SI(g3129), .SE(n10200), .CLK(n10552), 
        .Q(test_so91) );
  SDFFX1 DFF_1304_Q_reg ( .D(g33047), .SI(test_si92), .SE(n10250), .CLK(n10602), .Q(g5170), .QN(n10052) );
  SDFFX1 DFF_1305_Q_reg ( .D(g24298), .SI(g5170), .SE(n10252), .CLK(n10604), 
        .Q(g26959) );
  SDFFX1 DFF_1306_Q_reg ( .D(g25733), .SI(g26959), .SE(n10181), .CLK(n10533), 
        .Q(g5821), .QN(n5429) );
  SDFFX1 DFF_1307_Q_reg ( .D(g30536), .SI(g5821), .SE(n10226), .CLK(n10578), 
        .Q(g6299), .QN(n9880) );
  SDFFX1 DFF_1308_Q_reg ( .D(g7916), .SI(g6299), .SE(n10234), .CLK(n10586), 
        .Q(g8416), .QN(n9638) );
  SDFFX1 DFF_1310_Q_reg ( .D(g29246), .SI(g8416), .SE(n10204), .CLK(n10556), 
        .Q(g2079), .QN(n9829) );
  SDFFX1 DFF_1311_Q_reg ( .D(g34261), .SI(g2079), .SE(n10179), .CLK(n10531), 
        .Q(g4698), .QN(n5862) );
  SDFFX1 DFF_1312_Q_reg ( .D(g33611), .SI(g4698), .SE(n10261), .CLK(n10613), 
        .Q(g3703), .QN(n5399) );
  SDFFX1 DFF_1313_Q_reg ( .D(g25638), .SI(g3703), .SE(n10258), .CLK(n10610), 
        .Q(g1559), .QN(n5441) );
  SDFFX1 DFF_1314_Q_reg ( .D(g34728), .SI(g1559), .SE(n10197), .CLK(n10549), 
        .Q(n9247), .QN(n18478) );
  SDFFX1 DFF_1315_Q_reg ( .D(g29222), .SI(n9247), .SE(n10171), .CLK(n10523), 
        .Q(g411), .QN(n5629) );
  SDFFX1 DFF_1316_Q_reg ( .D(g25742), .SI(g411), .SE(n10267), .CLK(n10619), 
        .Q(test_so92), .QN(n5718) );
  SDFFX1 DFF_1317_Q_reg ( .D(g30449), .SI(test_si93), .SE(n10215), .CLK(n10567), .Q(g3953), .QN(n9875) );
  SDFFX1 DFF_1319_Q_reg ( .D(g34608), .SI(g3953), .SE(n10215), .CLK(n10567), 
        .Q(g2704), .QN(n5377) );
  SDFFX1 DFF_1320_Q_reg ( .D(g24345), .SI(g2704), .SE(n10260), .CLK(n10612), 
        .Q(g6035), .QN(n5528) );
  SDFFX1 DFF_1322_Q_reg ( .D(g34977), .SI(g6035), .SE(n10260), .CLK(n10612), 
        .Q(n9245) );
  SDFFX1 DFF_1323_Q_reg ( .D(g25635), .SI(n9245), .SE(n10201), .CLK(n10553), 
        .Q(g1300) );
  SDFFX1 DFF_1324_Q_reg ( .D(g25686), .SI(g1300), .SE(n10239), .CLK(n10591), 
        .Q(g4057), .QN(n5711) );
  SDFFX1 DFF_1325_Q_reg ( .D(g30461), .SI(g4057), .SE(n10253), .CLK(n10605), 
        .Q(g5200), .QN(n9813) );
  SDFFX1 DFF_1326_Q_reg ( .D(g34466), .SI(g5200), .SE(n10225), .CLK(n10577), 
        .Q(g4843), .QN(n9705) );
  SDFFX1 DFF_1327_Q_reg ( .D(g31901), .SI(g4843), .SE(n10202), .CLK(n10554), 
        .Q(g5046), .QN(n5578) );
  SDFFX1 DFF_1328_Q_reg ( .D(g29249), .SI(g5046), .SE(n10209), .CLK(n10561), 
        .Q(g2250), .QN(n9821) );
  SDFFX1 DFF_1329_Q_reg ( .D(g26882), .SI(g2250), .SE(n10209), .CLK(n10561), 
        .Q(g26885), .QN(n5456) );
  SDFFX1 DFF_1330_Q_reg ( .D(g33041), .SI(g26885), .SE(n10243), .CLK(n10595), 
        .Q(test_so93) );
  SDFFX1 DFF_1331_Q_reg ( .D(g33011), .SI(test_si94), .SE(n10268), .CLK(n10620), .Q(g2453), .QN(n5373) );
  SDFFX1 DFF_1332_Q_reg ( .D(g25734), .SI(g2453), .SE(n10181), .CLK(n10533), 
        .Q(g5841), .QN(n5449) );
  SDFFX1 DFF_1335_Q_reg ( .D(g12300), .SI(g5841), .SE(n10182), .CLK(n10534), 
        .Q(g14694), .QN(n5705) );
  SDFFX1 DFF_1336_Q_reg ( .D(g34618), .SI(g14694), .SE(n10198), .CLK(n10550), 
        .Q(g2912), .QN(n10080) );
  SDFFX1 DFF_1337_Q_reg ( .D(g33010), .SI(g2912), .SE(n10219), .CLK(n10571), 
        .Q(g2357), .QN(n5276) );
  SDFFX1 DFF_1338_Q_reg ( .D(g8919), .SI(g2357), .SE(n10219), .CLK(n10571), 
        .Q(g8920) );
  SDFFX1 DFF_1339_Q_reg ( .D(g31864), .SI(g8920), .SE(n10230), .CLK(n10582), 
        .Q(g164), .QN(n5561) );
  SDFFX1 DFF_1340_Q_reg ( .D(g34630), .SI(g164), .SE(n10230), .CLK(n10582), 
        .Q(g4253), .QN(n5484) );
  SDFFX1 DFF_1341_Q_reg ( .D(g31898), .SI(g4253), .SE(n10208), .CLK(n10560), 
        .Q(g5016), .QN(n5369) );
  SDFFX1 DFF_1342_Q_reg ( .D(g25653), .SI(g5016), .SE(n10190), .CLK(n10542), 
        .Q(g3119), .QN(n5423) );
  SDFFX1 DFF_1343_Q_reg ( .D(g25632), .SI(g3119), .SE(n10201), .CLK(n10553), 
        .Q(g1351), .QN(n5322) );
  SDFFX1 DFF_1344_Q_reg ( .D(g32988), .SI(g1351), .SE(n10201), .CLK(n10553), 
        .Q(test_so94), .QN(n10121) );
  SDFFX1 DFF_1345_Q_reg ( .D(g33616), .SI(test_si95), .SE(n10174), .CLK(n10526), .Q(g4519) );
  SDFFX1 DFF_1346_Q_reg ( .D(g29280), .SI(g4519), .SE(n10178), .CLK(n10530), 
        .Q(g5115), .QN(n5743) );
  SDFFX1 DFF_1347_Q_reg ( .D(g33609), .SI(g5115), .SE(n10261), .CLK(n10613), 
        .Q(g3352), .QN(n5604) );
  SDFFX1 DFF_1348_Q_reg ( .D(g30563), .SI(g3352), .SE(n10194), .CLK(n10546), 
        .Q(g6657), .QN(n9799) );
  SDFFX1 DFF_1349_Q_reg ( .D(g33044), .SI(g6657), .SE(n10243), .CLK(n10595), 
        .Q(g4552) );
  SDFFX1 DFF_1350_Q_reg ( .D(g30437), .SI(g4552), .SE(n10215), .CLK(n10567), 
        .Q(g3893), .QN(n9818) );
  SDFFX1 DFF_1351_Q_reg ( .D(g30412), .SI(g3893), .SE(n10231), .CLK(n10583), 
        .Q(g3211), .QN(n10007) );
  SDFFX1 DFF_1352_Q_reg ( .D(g17604), .SI(g3211), .SE(n10233), .CLK(n10585), 
        .Q(g13049) );
  SDFFX1 DFF_1354_Q_reg ( .D(g16603), .SI(g13049), .SE(n10243), .CLK(n10595), 
        .Q(g16624), .QN(n9971) );
  SDFFX1 DFF_1355_Q_reg ( .D(g30491), .SI(g16624), .SE(n10175), .CLK(n10527), 
        .Q(g5595), .QN(n9983) );
  SDFFX1 DFF_1356_Q_reg ( .D(g30434), .SI(g5595), .SE(n10251), .CLK(n10603), 
        .Q(g3614), .QN(n9802) );
  SDFFX1 DFF_1357_Q_reg ( .D(g34612), .SI(g3614), .SE(n10199), .CLK(n10551), 
        .Q(test_so95) );
  SDFFX1 DFF_1358_Q_reg ( .D(g29259), .SI(test_si96), .SE(n10190), .CLK(n10542), .Q(g3125), .QN(n5781) );
  SDFFX1 DFF_1359_Q_reg ( .D(g13865), .SI(g3125), .SE(n10200), .CLK(n10552), 
        .Q(g16686) );
  SDFFX1 DFF_1360_Q_reg ( .D(g25681), .SI(g16686), .SE(n10167), .CLK(n10519), 
        .Q(g3821), .QN(n5428) );
  SDFFX1 DFF_1361_Q_reg ( .D(g25687), .SI(g3821), .SE(n10239), .CLK(n10591), 
        .Q(g4141), .QN(n5612) );
  SDFFX1 DFF_1362_Q_reg ( .D(g33617), .SI(g4141), .SE(n10243), .CLK(n10595), 
        .Q(g4570) );
  SDFFX1 DFF_1363_Q_reg ( .D(g30479), .SI(g4570), .SE(n10217), .CLK(n10569), 
        .Q(g5272), .QN(n9810) );
  SDFFX1 DFF_1364_Q_reg ( .D(g29256), .SI(g5272), .SE(n10256), .CLK(n10608), 
        .Q(g2735), .QN(n5600) );
  SDFFX1 DFF_1365_Q_reg ( .D(g28054), .SI(g2735), .SE(n10256), .CLK(n10608), 
        .Q(g728), .QN(n9790) );
  SDFFX1 DFF_1366_Q_reg ( .D(g30535), .SI(g728), .SE(n10266), .CLK(n10618), 
        .Q(g6295), .QN(n9807) );
  SDFFX1 DFF_1368_Q_reg ( .D(g30385), .SI(g6295), .SE(n10177), .CLK(n10529), 
        .Q(g2661), .QN(n5418) );
  SDFFX1 DFF_1369_Q_reg ( .D(g30361), .SI(g2661), .SE(n10169), .CLK(n10521), 
        .Q(g1988), .QN(n5783) );
  SDFFX1 DFF_1370_Q_reg ( .D(g25705), .SI(g1988), .SE(n10178), .CLK(n10530), 
        .Q(test_so96), .QN(n10141) );
  SDFFX1 DFF_1371_Q_reg ( .D(g24260), .SI(test_si97), .SE(n10258), .CLK(n10610), .Q(g1548), .QN(n5546) );
  SDFFX1 DFF_1372_Q_reg ( .D(g29257), .SI(g1548), .SE(n10190), .CLK(n10542), 
        .Q(g3106), .QN(n5742) );
  SDFFX1 DFF_1373_Q_reg ( .D(g34461), .SI(g3106), .SE(n10260), .CLK(n10612), 
        .Q(g4659), .QN(n10064) );
  SDFFX1 DFF_1374_Q_reg ( .D(g34258), .SI(g4659), .SE(n10260), .CLK(n10612), 
        .Q(g4358), .QN(n5348) );
  SDFFX1 DFF_1375_Q_reg ( .D(g32993), .SI(g4358), .SE(n10208), .CLK(n10560), 
        .Q(g1792), .QN(n5359) );
  SDFFX1 DFF_1376_Q_reg ( .D(g33992), .SI(g1792), .SE(n10213), .CLK(n10565), 
        .Q(g2084), .QN(n9691) );
  SDFFX1 DFF_1378_Q_reg ( .D(g30394), .SI(g2084), .SE(n10257), .CLK(n10609), 
        .Q(g3187), .QN(n9950) );
  SDFFX1 DFF_1379_Q_reg ( .D(g34449), .SI(g3187), .SE(n10261), .CLK(n10613), 
        .Q(g4311), .QN(n5323) );
  SDFFX1 DFF_1380_Q_reg ( .D(g34019), .SI(g4311), .SE(n10212), .CLK(n10564), 
        .Q(g2583), .QN(n5800) );
  SDFFX1 DFF_1381_Q_reg ( .D(g18597), .SI(g2583), .SE(n10166), .CLK(n10518), 
        .Q(n9240), .QN(DFF_1381_n1) );
  SDFFX1 DFF_1382_Q_reg ( .D(g29231), .SI(n9240), .SE(n10166), .CLK(n10518), 
        .Q(g1094), .QN(n5697) );
  SDFFX1 DFF_1383_Q_reg ( .D(g25682), .SI(g1094), .SE(n10167), .CLK(n10519), 
        .Q(test_so97), .QN(n10160) );
  SDFFX1 DFF_1384_Q_reg ( .D(g21897), .SI(test_si98), .SE(n10231), .CLK(n10583), .Q(g4284), .QN(n9725) );
  SDFFX1 DFF_1386_Q_reg ( .D(g30395), .SI(g4284), .SE(n10231), .CLK(n10583), 
        .Q(g3191), .QN(n9794) );
  SDFFX1 DFF_1387_Q_reg ( .D(g21892), .SI(g3191), .SE(n10227), .CLK(n10579), 
        .Q(g4239), .QN(n9706) );
  SDFFX1 DFF_1389_Q_reg ( .D(g8789), .SI(g4239), .SE(n10227), .CLK(n10579), 
        .Q(g4180), .QN(n5380) );
  SDFFX1 DFF_1390_Q_reg ( .D(g28048), .SI(g4180), .SE(n10172), .CLK(n10524), 
        .Q(g691), .QN(n5520) );
  SDFFX1 DFF_1391_Q_reg ( .D(g34723), .SI(g691), .SE(n10172), .CLK(n10524), 
        .Q(g534), .QN(n5490) );
  SDFFX1 DFF_1393_Q_reg ( .D(g25598), .SI(g534), .SE(n10245), .CLK(n10597), 
        .Q(g385), .QN(n5632) );
  SDFFX1 DFF_1394_Q_reg ( .D(g33987), .SI(g385), .SE(n10214), .CLK(n10566), 
        .Q(g2004), .QN(n5818) );
  SDFFX1 DFF_1395_Q_reg ( .D(g30380), .SI(g2004), .SE(n10206), .CLK(n10558), 
        .Q(g2527), .QN(n5420) );
  SDFFX1 DFF_1396_Q_reg ( .D(g9555), .SI(g2527), .SE(n10246), .CLK(n10598), 
        .Q(g5456) );
  SDFFX1 DFF_1397_Q_reg ( .D(g26965), .SI(g5456), .SE(n10264), .CLK(n10616), 
        .Q(n6007) );
  SDFFX1 DFF_1398_Q_reg ( .D(g25706), .SI(n6007), .SE(n10178), .CLK(n10530), 
        .Q(test_so98), .QN(n10159) );
  SDFFX1 DFF_1399_Q_reg ( .D(g30458), .SI(test_si99), .SE(n10195), .CLK(n10547), .Q(g4507), .QN(n5846) );
  SDFFX1 DFF_1400_Q_reg ( .D(g24338), .SI(g4507), .SE(n10178), .CLK(n10530), 
        .Q(g5348), .QN(n10039) );
  SDFFX1 DFF_1401_Q_reg ( .D(g30400), .SI(g5348), .SE(n10231), .CLK(n10583), 
        .Q(g3223), .QN(n9918) );
  SDFFX1 DFF_1403_Q_reg ( .D(g34623), .SI(g3223), .SE(n10182), .CLK(n10534), 
        .Q(g2970), .QN(n10079) );
  SDFFX1 DFF_1404_Q_reg ( .D(g24343), .SI(g2970), .SE(n10182), .CLK(n10534), 
        .Q(g5698), .QN(n9903) );
  SDFFX1 DFF_1406_Q_reg ( .D(g30473), .SI(g5698), .SE(n10264), .CLK(n10616), 
        .Q(g5260), .QN(n9869) );
  SDFFX1 DFF_1407_Q_reg ( .D(g24252), .SI(g5260), .SE(n10229), .CLK(n10581), 
        .Q(g1521), .QN(n5577) );
  SDFFX1 DFF_1408_Q_reg ( .D(g33028), .SI(g1521), .SE(n10241), .CLK(n10593), 
        .Q(g3522), .QN(n5383) );
  SDFFX1 DFF_1409_Q_reg ( .D(g29258), .SI(g3522), .SE(n10190), .CLK(n10542), 
        .Q(g3115), .QN(n9664) );
  SDFFX1 DFF_1410_Q_reg ( .D(g30407), .SI(g3115), .SE(n10231), .CLK(n10583), 
        .Q(g3251), .QN(n9867) );
  SDFFX1 DFF_1411_Q_reg ( .D(g26958), .SI(g3251), .SE(n10172), .CLK(n10524), 
        .Q(g12832) );
  SDFFX1 DFF_1412_Q_reg ( .D(g34457), .SI(g12832), .SE(n10172), .CLK(n10524), 
        .Q(test_so99) );
  SDFFX1 DFF_1413_Q_reg ( .D(g33568), .SI(test_si100), .SE(n10267), .CLK(
        n10619), .Q(g1996), .QN(n5355) );
  SDFFX1 DFF_1414_Q_reg ( .D(g25663), .SI(g1996), .SE(n10267), .CLK(n10619), 
        .Q(g8342) );
  SDFFX1 DFF_1415_Q_reg ( .D(g26964), .SI(g8342), .SE(n10205), .CLK(n10557), 
        .Q(g4515), .QN(n10046) );
  SDFFX1 DFF_1416_Q_reg ( .D(g8786), .SI(g4515), .SE(n10206), .CLK(n10558), 
        .Q(g8787) );
  SDFFX1 DFF_1417_Q_reg ( .D(g34735), .SI(g8787), .SE(n10175), .CLK(n10527), 
        .Q(g4300), .QN(n5639) );
  SDFFX1 DFF_1418_Q_reg ( .D(g30352), .SI(g4300), .SE(n10270), .CLK(n10622), 
        .Q(n9236), .QN(n18480) );
  SDFFX1 DFF_1419_Q_reg ( .D(g33543), .SI(n9236), .SE(n10201), .CLK(n10553), 
        .Q(g1379), .QN(n9685) );
  SDFFX1 DFF_1420_Q_reg ( .D(g24271), .SI(g1379), .SE(n10221), .CLK(n10573), 
        .Q(g11388), .QN(n5433) );
  SDFFX1 DFF_1422_Q_reg ( .D(g33981), .SI(g11388), .SE(n10203), .CLK(n10555), 
        .Q(g1878), .QN(n5793) );
  SDFFX1 DFF_1423_Q_reg ( .D(g30500), .SI(g1878), .SE(n10174), .CLK(n10526), 
        .Q(g5619), .QN(n9795) );
  SDFFX1 DFF_1424_Q_reg ( .D(g34649), .SI(g5619), .SE(n10168), .CLK(n10520), 
        .Q(g71), .QN(n18464) );
  SDFFX1 DFF_1425_Q_reg ( .D(g29277), .SI(g71), .SE(n10174), .CLK(n10526), .Q(
        test_so100), .QN(n10150) );
  SDFFX1 DFF_748_Q_reg ( .D(n1030), .SI(g4704), .SE(n10197), .CLK(n10549), .Q(
        g22), .QN(n9723) );
  SDFFX1 DFF_591_Q_reg ( .D(g25612), .SI(g3897), .SE(n10245), .CLK(n10597), 
        .Q(g518), .QN(n5287) );
  SDFFX1 DFF_845_Q_reg ( .D(g28060), .SI(g626), .SE(n10256), .CLK(n10608), .Q(
        g2729), .QN(n9780) );
  HADDX1 Trojan_U1_1_30 ( .A0(counter_30), .B0(carry_30), .C1(carry_31), .SO(
        N31) );
  HADDX1 Trojan_U1_1_4 ( .A0(counter_4), .B0(carry_4), .C1(carry_5), .SO(N5)
         );
  HADDX1 Trojan_U1_1_5 ( .A0(counter_5), .B0(carry_5), .C1(carry_6), .SO(N6)
         );
  HADDX1 Trojan_U1_1_6 ( .A0(counter_6), .B0(carry_6), .C1(carry_7), .SO(N7)
         );
  HADDX1 Trojan_U1_1_7 ( .A0(counter_7), .B0(carry_7), .C1(carry_8), .SO(N8)
         );
  HADDX1 Trojan_U1_1_8 ( .A0(counter_8), .B0(carry_8), .C1(carry_9), .SO(N9)
         );
  HADDX1 Trojan_U1_1_9 ( .A0(counter_9), .B0(carry_9), .C1(carry_10), .SO(N10)
         );
  HADDX1 Trojan_U1_1_10 ( .A0(counter_10), .B0(carry_10), .C1(carry_11), .SO(
        N11) );
  HADDX1 Trojan_U1_1_11 ( .A0(counter_11), .B0(carry_11), .C1(carry_12), .SO(
        N12) );
  HADDX1 Trojan_U1_1_12 ( .A0(counter_12), .B0(carry_12), .C1(carry_13), .SO(
        N13) );
  HADDX1 Trojan_U1_1_13 ( .A0(counter_13), .B0(carry_13), .C1(carry_14), .SO(
        N14) );
  HADDX1 Trojan_U1_1_14 ( .A0(counter_14), .B0(carry_14), .C1(carry_15), .SO(
        N15) );
  HADDX1 Trojan_U1_1_22 ( .A0(counter_22), .B0(carry_22), .C1(carry_23), .SO(
        N23) );
  HADDX1 Trojan_U1_1_23 ( .A0(counter_23), .B0(carry_23), .C1(carry_24), .SO(
        N24) );
  HADDX1 Trojan_U1_1_24 ( .A0(counter_24), .B0(carry_24), .C1(carry_25), .SO(
        N25) );
  HADDX1 Trojan_U1_1_25 ( .A0(counter_25), .B0(carry_25), .C1(carry_26), .SO(
        N26) );
  HADDX1 Trojan_U1_1_1 ( .A0(counter_1), .B0(counter_0), .C1(carry_2), .SO(N2)
         );
  HADDX1 Trojan_U1_1_2 ( .A0(counter_2), .B0(carry_2), .C1(carry_3), .SO(N3)
         );
  HADDX1 Trojan_U1_1_3 ( .A0(counter_3), .B0(carry_3), .C1(carry_4), .SO(N4)
         );
  HADDX1 Trojan_U1_1_15 ( .A0(counter_15), .B0(carry_15), .C1(carry_16), .SO(
        N16) );
  HADDX1 Trojan_U1_1_16 ( .A0(counter_16), .B0(carry_16), .C1(carry_17), .SO(
        N17) );
  HADDX1 Trojan_U1_1_17 ( .A0(counter_17), .B0(carry_17), .C1(carry_18), .SO(
        N18) );
  HADDX1 Trojan_U1_1_18 ( .A0(counter_18), .B0(carry_18), .C1(carry_19), .SO(
        N19) );
  HADDX1 Trojan_U1_1_19 ( .A0(counter_19), .B0(carry_19), .C1(carry_20), .SO(
        N20) );
  HADDX1 Trojan_U1_1_20 ( .A0(counter_20), .B0(carry_20), .C1(carry_21), .SO(
        N21) );
  HADDX1 Trojan_U1_1_21 ( .A0(counter_21), .B0(carry_21), .C1(carry_22), .SO(
        N22) );
  HADDX1 Trojan_U1_1_26 ( .A0(counter_26), .B0(carry_26), .C1(carry_27), .SO(
        N27) );
  HADDX1 Trojan_U1_1_27 ( .A0(counter_27), .B0(carry_27), .C1(carry_28), .SO(
        N28) );
  HADDX1 Trojan_U1_1_28 ( .A0(counter_28), .B0(carry_28), .C1(carry_29), .SO(
        N29) );
  HADDX1 Trojan_U1_1_29 ( .A0(counter_29), .B0(carry_29), .C1(carry_30), .SO(
        N30) );
  INVX0 Trojan_U1 ( .INP(counter_0), .ZN(N1) );
  XOR2X1 Trojan_U2 ( .IN1(carry_31), .IN2(counter_31), .Q(N32) );
  DFFARX1 Trojan_counter_reg_31_ ( .D(N32), .CLK(n37), .RSTB(n10164), .Q(
        counter_31), .QN(n73) );
  DFFARX1 Trojan_counter_reg_1_ ( .D(N2), .CLK(n37), .RSTB(n10163), .Q(
        counter_1) );
  DFFARX1 Trojan_counter_reg_2_ ( .D(N3), .CLK(n37), .RSTB(n87), .Q(counter_2)
         );
  DFFARX1 Trojan_counter_reg_3_ ( .D(N4), .CLK(n37), .RSTB(n10164), .Q(
        counter_3), .QN(n86) );
  DFFARX1 Trojan_counter_reg_15_ ( .D(N16), .CLK(n37), .RSTB(n10163), .Q(
        counter_15), .QN(n85) );
  DFFARX1 Trojan_counter_reg_16_ ( .D(N17), .CLK(n37), .RSTB(n87), .Q(
        counter_16), .QN(n84) );
  DFFARX1 Trojan_counter_reg_17_ ( .D(N18), .CLK(n37), .RSTB(n10164), .Q(
        counter_17), .QN(n83) );
  DFFARX1 Trojan_counter_reg_18_ ( .D(N19), .CLK(n37), .RSTB(n10163), .Q(
        counter_18), .QN(n82) );
  DFFARX1 Trojan_counter_reg_19_ ( .D(N20), .CLK(n37), .RSTB(n87), .Q(
        counter_19), .QN(n81) );
  DFFARX1 Trojan_counter_reg_20_ ( .D(N21), .CLK(n37), .RSTB(n10164), .Q(
        counter_20), .QN(n80) );
  DFFARX1 Trojan_counter_reg_21_ ( .D(N22), .CLK(n37), .RSTB(n10163), .Q(
        counter_21), .QN(n79) );
  DFFARX1 Trojan_counter_reg_26_ ( .D(N27), .CLK(n37), .RSTB(n87), .Q(
        counter_26), .QN(n78) );
  DFFARX1 Trojan_counter_reg_27_ ( .D(N28), .CLK(n37), .RSTB(n10164), .Q(
        counter_27), .QN(n77) );
  DFFARX1 Trojan_counter_reg_28_ ( .D(N29), .CLK(n37), .RSTB(n10163), .Q(
        counter_28), .QN(n76) );
  DFFARX1 Trojan_counter_reg_29_ ( .D(N30), .CLK(n37), .RSTB(n87), .Q(
        counter_29), .QN(n75) );
  DFFARX1 Trojan_counter_reg_30_ ( .D(N31), .CLK(n37), .RSTB(n10164), .Q(
        counter_30), .QN(n74) );
  DFFARX1 Trojan_counter_reg_7_ ( .D(N8), .CLK(n37), .RSTB(n10163), .Q(
        counter_7) );
  DFFARX1 Trojan_counter_reg_11_ ( .D(N12), .CLK(n37), .RSTB(n87), .Q(
        counter_11) );
  DFFARX1 Trojan_counter_reg_25_ ( .D(N26), .CLK(n37), .RSTB(n10164), .Q(
        counter_25) );
  DFFARX1 Trojan_counter_reg_6_ ( .D(N7), .CLK(n37), .RSTB(n10163), .Q(
        counter_6) );
  DFFARX1 Trojan_counter_reg_10_ ( .D(N11), .CLK(n37), .RSTB(n87), .Q(
        counter_10) );
  DFFARX1 Trojan_counter_reg_12_ ( .D(N13), .CLK(n37), .RSTB(n10164), .Q(
        counter_12) );
  DFFARX1 Trojan_counter_reg_24_ ( .D(N25), .CLK(n37), .RSTB(n10163), .Q(
        counter_24) );
  DFFARX1 Trojan_counter_reg_4_ ( .D(N5), .CLK(n37), .RSTB(n87), .Q(counter_4)
         );
  DFFARX1 Trojan_counter_reg_5_ ( .D(N6), .CLK(n37), .RSTB(n10164), .Q(
        counter_5) );
  DFFARX1 Trojan_counter_reg_9_ ( .D(N10), .CLK(n37), .RSTB(n10163), .Q(
        counter_9) );
  DFFARX1 Trojan_counter_reg_14_ ( .D(N15), .CLK(n37), .RSTB(n87), .Q(
        counter_14) );
  DFFARX1 Trojan_counter_reg_23_ ( .D(N24), .CLK(n37), .RSTB(n10164), .Q(
        counter_23) );
  DFFARX1 Trojan_counter_reg_8_ ( .D(N9), .CLK(n37), .RSTB(n10163), .Q(
        counter_8) );
  DFFARX1 Trojan_counter_reg_13_ ( .D(N14), .CLK(n37), .RSTB(n87), .Q(
        counter_13) );
  DFFARX1 Trojan_counter_reg_22_ ( .D(N23), .CLK(n37), .RSTB(n10164), .Q(
        counter_22) );
  DFFARX1 Trojan_counter_reg_0_ ( .D(N1), .CLK(n37), .RSTB(n10163), .Q(
        counter_0) );
  NAND4X0 Trojan_U14 ( .IN1(n3180), .IN2(n3121), .IN3(n2461), .IN4(n58), .QN(
        n87) );
  INVX0 Trojan_U15 ( .INP(n59), .ZN(n58) );
  NOR4X0 Trojan_U16 ( .IN1(n3180), .IN2(n3121), .IN3(n2461), .IN4(n59), .QN(
        n37) );
  NAND3X0 Trojan_U17 ( .IN1(n2601), .IN2(n5111), .IN3(n60), .QN(n59) );
  AND3X1 Trojan_U18 ( .IN1(n2396), .IN2(n36), .IN3(n10106), .Q(n60) );
  NOR4X0 Trojan_U19 ( .IN1(n61), .IN2(n62), .IN3(n63), .IN4(n64), .QN(
        Trigger_out) );
  NAND4X0 Trojan_U20 ( .IN1(n78), .IN2(n77), .IN3(n76), .IN4(n75), .QN(n64) );
  NAND4X0 Trojan_U21 ( .IN1(n74), .IN2(n73), .IN3(counter_6), .IN4(counter_5), 
        .QN(n63) );
  NAND4X0 Trojan_U22 ( .IN1(n80), .IN2(n79), .IN3(n81), .IN4(n65), .QN(n62) );
  NOR4X0 Trojan_U23 ( .IN1(counter_25), .IN2(counter_24), .IN3(counter_23), 
        .IN4(counter_22), .QN(n65) );
  NAND4X0 Trojan_U24 ( .IN1(n66), .IN2(n67), .IN3(n68), .IN4(n69), .QN(n61) );
  NOR4X0 Trojan_U25 ( .IN1(n70), .IN2(counter_12), .IN3(counter_14), .IN4(
        counter_13), .QN(n69) );
  NAND4X0 Trojan_U26 ( .IN1(n85), .IN2(n84), .IN3(n83), .IN4(n82), .QN(n70) );
  NOR4X0 Trojan_U27 ( .IN1(counter_11), .IN2(counter_10), .IN3(counter_9), 
        .IN4(counter_8), .QN(n68) );
  MUX21X1 Trojan_U28 ( .IN1(n71), .IN2(n72), .S(n86), .Q(n67) );
  OA21X1 Trojan_U29 ( .IN1(counter_1), .IN2(counter_0), .IN3(counter_2), .Q(
        n72) );
  NAND2X0 Trojan_U30 ( .IN1(counter_2), .IN2(counter_1), .QN(n71) );
  NOR2X0 Trojan_U31 ( .IN1(counter_7), .IN2(counter_4), .QN(n66) );
  MUX21X1 Trojan_Paylod ( .IN1(g10122_Tj), .IN2(g25715), .S(Trigger_out), .Q(
        g10122) );
  INVX0 U10091 ( .INP(n87), .ZN(n10162) );
  INVX0 U10092 ( .INP(n10162), .ZN(n10163) );
  INVX0 U10093 ( .INP(n10162), .ZN(n10164) );
  NBUFFX2 U10094 ( .INP(n10293), .Z(n10166) );
  NBUFFX2 U10095 ( .INP(n10293), .Z(n10165) );
  NBUFFX2 U10096 ( .INP(n10285), .Z(n10204) );
  NBUFFX2 U10097 ( .INP(n10282), .Z(n10218) );
  NBUFFX2 U10098 ( .INP(n10290), .Z(n10178) );
  NBUFFX2 U10099 ( .INP(n10288), .Z(n10189) );
  NBUFFX2 U10100 ( .INP(n10274), .Z(n10258) );
  NBUFFX2 U10101 ( .INP(n10285), .Z(n10202) );
  NBUFFX2 U10102 ( .INP(n10280), .Z(n10230) );
  NBUFFX2 U10103 ( .INP(n10274), .Z(n10257) );
  NBUFFX2 U10104 ( .INP(n10273), .Z(n10266) );
  NBUFFX2 U10105 ( .INP(n10283), .Z(n10215) );
  NBUFFX2 U10106 ( .INP(n10276), .Z(n10251) );
  NBUFFX2 U10107 ( .INP(n10289), .Z(n10186) );
  NBUFFX2 U10108 ( .INP(n10285), .Z(n10206) );
  NBUFFX2 U10109 ( .INP(n10284), .Z(n10211) );
  NBUFFX2 U10110 ( .INP(n10292), .Z(n10167) );
  NBUFFX2 U10111 ( .INP(n10292), .Z(n10170) );
  NBUFFX2 U10112 ( .INP(n10284), .Z(n10210) );
  NBUFFX2 U10113 ( .INP(n10283), .Z(n10214) );
  NBUFFX2 U10114 ( .INP(n10288), .Z(n10188) );
  NBUFFX2 U10115 ( .INP(n10287), .Z(n10192) );
  NBUFFX2 U10116 ( .INP(n10273), .Z(n10265) );
  NBUFFX2 U10117 ( .INP(n10275), .Z(n10252) );
  NBUFFX2 U10118 ( .INP(n10287), .Z(n10193) );
  NBUFFX2 U10119 ( .INP(n10287), .Z(n10194) );
  NBUFFX2 U10120 ( .INP(n10290), .Z(n10181) );
  NBUFFX2 U10121 ( .INP(n10291), .Z(n10176) );
  NBUFFX2 U10122 ( .INP(n10287), .Z(n10195) );
  NBUFFX2 U10123 ( .INP(n10283), .Z(n10212) );
  NBUFFX2 U10124 ( .INP(n10279), .Z(n10236) );
  NBUFFX2 U10125 ( .INP(n10273), .Z(n10264) );
  NBUFFX2 U10126 ( .INP(n10279), .Z(n10234) );
  NBUFFX2 U10127 ( .INP(n10291), .Z(n10172) );
  NBUFFX2 U10128 ( .INP(n10278), .Z(n10239) );
  NBUFFX2 U10129 ( .INP(n10284), .Z(n10208) );
  NBUFFX2 U10130 ( .INP(n10276), .Z(n10247) );
  NBUFFX2 U10131 ( .INP(n10291), .Z(n10175) );
  NBUFFX2 U10132 ( .INP(n10273), .Z(n10262) );
  NBUFFX2 U10133 ( .INP(n10288), .Z(n10190) );
  NBUFFX2 U10134 ( .INP(n10274), .Z(n10261) );
  NBUFFX2 U10135 ( .INP(n10278), .Z(n10237) );
  NBUFFX2 U10136 ( .INP(n10280), .Z(n10231) );
  NBUFFX2 U10137 ( .INP(n10282), .Z(n10217) );
  NBUFFX2 U10138 ( .INP(n10276), .Z(n10248) );
  NBUFFX2 U10139 ( .INP(n10286), .Z(n10197) );
  NBUFFX2 U10140 ( .INP(n10275), .Z(n10256) );
  NBUFFX2 U10141 ( .INP(n10278), .Z(n10241) );
  NBUFFX2 U10142 ( .INP(n10286), .Z(n10199) );
  NBUFFX2 U10143 ( .INP(n10280), .Z(n10228) );
  NBUFFX2 U10144 ( .INP(n10279), .Z(n10233) );
  NBUFFX2 U10145 ( .INP(n10275), .Z(n10253) );
  NBUFFX2 U10146 ( .INP(n10275), .Z(n10255) );
  NBUFFX2 U10147 ( .INP(n10287), .Z(n10196) );
  NBUFFX2 U10148 ( .INP(n10281), .Z(n10225) );
  NBUFFX2 U10149 ( .INP(n10289), .Z(n10183) );
  NBUFFX2 U10150 ( .INP(n10278), .Z(n10240) );
  NBUFFX2 U10151 ( .INP(n10282), .Z(n10220) );
  NBUFFX2 U10152 ( .INP(n10281), .Z(n10226) );
  NBUFFX2 U10153 ( .INP(n10281), .Z(n10222) );
  NBUFFX2 U10154 ( .INP(n10285), .Z(n10205) );
  NBUFFX2 U10155 ( .INP(n10283), .Z(n10213) );
  NBUFFX2 U10156 ( .INP(n10276), .Z(n10250) );
  NBUFFX2 U10157 ( .INP(n10280), .Z(n10229) );
  NBUFFX2 U10158 ( .INP(n10286), .Z(n10201) );
  NBUFFX2 U10159 ( .INP(n10276), .Z(n10249) );
  NBUFFX2 U10160 ( .INP(n10280), .Z(n10227) );
  NBUFFX2 U10161 ( .INP(n10277), .Z(n10243) );
  NBUFFX2 U10162 ( .INP(n10291), .Z(n10174) );
  NBUFFX2 U10163 ( .INP(n10279), .Z(n10235) );
  NBUFFX2 U10164 ( .INP(n10290), .Z(n10179) );
  NBUFFX2 U10165 ( .INP(n10290), .Z(n10180) );
  NBUFFX2 U10166 ( .INP(n10278), .Z(n10238) );
  NBUFFX2 U10167 ( .INP(n10289), .Z(n10182) );
  NBUFFX2 U10168 ( .INP(n10290), .Z(n10177) );
  NBUFFX2 U10169 ( .INP(n10281), .Z(n10224) );
  NBUFFX2 U10170 ( .INP(n10292), .Z(n10169) );
  NBUFFX2 U10171 ( .INP(n10292), .Z(n10168) );
  NBUFFX2 U10172 ( .INP(n10277), .Z(n10244) );
  NBUFFX2 U10173 ( .INP(n10284), .Z(n10209) );
  NBUFFX2 U10174 ( .INP(n10277), .Z(n10246) );
  NBUFFX2 U10175 ( .INP(n10282), .Z(n10221) );
  NBUFFX2 U10176 ( .INP(n10282), .Z(n10219) );
  NBUFFX2 U10177 ( .INP(n10289), .Z(n10185) );
  NBUFFX2 U10178 ( .INP(n10288), .Z(n10191) );
  NBUFFX2 U10179 ( .INP(n10291), .Z(n10173) );
  NBUFFX2 U10180 ( .INP(n10292), .Z(n10171) );
  NBUFFX2 U10181 ( .INP(n10274), .Z(n10260) );
  NBUFFX2 U10182 ( .INP(n10274), .Z(n10259) );
  NBUFFX2 U10183 ( .INP(n10277), .Z(n10242) );
  NBUFFX2 U10184 ( .INP(n10288), .Z(n10187) );
  NBUFFX2 U10185 ( .INP(n10275), .Z(n10254) );
  NBUFFX2 U10186 ( .INP(n10286), .Z(n10198) );
  NBUFFX2 U10187 ( .INP(n10277), .Z(n10245) );
  NBUFFX2 U10188 ( .INP(n10283), .Z(n10216) );
  NBUFFX2 U10189 ( .INP(n10289), .Z(n10184) );
  NBUFFX2 U10190 ( .INP(n10279), .Z(n10232) );
  NBUFFX2 U10191 ( .INP(n10281), .Z(n10223) );
  NBUFFX2 U10192 ( .INP(n10284), .Z(n10207) );
  NBUFFX2 U10193 ( .INP(n10286), .Z(n10200) );
  NBUFFX2 U10194 ( .INP(n10273), .Z(n10263) );
  NBUFFX2 U10195 ( .INP(n10285), .Z(n10203) );
  NBUFFX2 U10196 ( .INP(n10645), .Z(n10518) );
  NBUFFX2 U10197 ( .INP(n10645), .Z(n10517) );
  NBUFFX2 U10198 ( .INP(n10637), .Z(n10556) );
  NBUFFX2 U10199 ( .INP(n10634), .Z(n10570) );
  NBUFFX2 U10200 ( .INP(n10642), .Z(n10530) );
  NBUFFX2 U10201 ( .INP(n10640), .Z(n10541) );
  NBUFFX2 U10202 ( .INP(n10626), .Z(n10610) );
  NBUFFX2 U10203 ( .INP(n10637), .Z(n10554) );
  NBUFFX2 U10204 ( .INP(n10632), .Z(n10582) );
  NBUFFX2 U10205 ( .INP(n10626), .Z(n10609) );
  NBUFFX2 U10206 ( .INP(n10625), .Z(n10618) );
  NBUFFX2 U10207 ( .INP(n10635), .Z(n10567) );
  NBUFFX2 U10208 ( .INP(n10628), .Z(n10603) );
  NBUFFX2 U10209 ( .INP(n10641), .Z(n10538) );
  NBUFFX2 U10210 ( .INP(n10637), .Z(n10558) );
  NBUFFX2 U10211 ( .INP(n10636), .Z(n10563) );
  NBUFFX2 U10212 ( .INP(n10644), .Z(n10519) );
  NBUFFX2 U10213 ( .INP(n10644), .Z(n10522) );
  NBUFFX2 U10214 ( .INP(n10636), .Z(n10562) );
  NBUFFX2 U10215 ( .INP(n10635), .Z(n10566) );
  NBUFFX2 U10216 ( .INP(n10640), .Z(n10540) );
  NBUFFX2 U10217 ( .INP(n10639), .Z(n10544) );
  NBUFFX2 U10218 ( .INP(n10625), .Z(n10617) );
  NBUFFX2 U10219 ( .INP(n10627), .Z(n10604) );
  NBUFFX2 U10220 ( .INP(n10639), .Z(n10545) );
  NBUFFX2 U10221 ( .INP(n10639), .Z(n10546) );
  NBUFFX2 U10222 ( .INP(n10642), .Z(n10533) );
  NBUFFX2 U10223 ( .INP(n10643), .Z(n10528) );
  NBUFFX2 U10224 ( .INP(n10639), .Z(n10547) );
  NBUFFX2 U10225 ( .INP(n10635), .Z(n10564) );
  NBUFFX2 U10226 ( .INP(n10631), .Z(n10588) );
  NBUFFX2 U10227 ( .INP(n10625), .Z(n10616) );
  NBUFFX2 U10228 ( .INP(n10631), .Z(n10586) );
  NBUFFX2 U10229 ( .INP(n10643), .Z(n10524) );
  NBUFFX2 U10230 ( .INP(n10630), .Z(n10591) );
  NBUFFX2 U10231 ( .INP(n10636), .Z(n10560) );
  NBUFFX2 U10232 ( .INP(n10628), .Z(n10599) );
  NBUFFX2 U10233 ( .INP(n10643), .Z(n10527) );
  NBUFFX2 U10234 ( .INP(n10625), .Z(n10614) );
  NBUFFX2 U10235 ( .INP(n10640), .Z(n10542) );
  NBUFFX2 U10236 ( .INP(n10626), .Z(n10613) );
  NBUFFX2 U10237 ( .INP(n10630), .Z(n10589) );
  NBUFFX2 U10238 ( .INP(n10632), .Z(n10583) );
  NBUFFX2 U10239 ( .INP(n10634), .Z(n10569) );
  NBUFFX2 U10240 ( .INP(n10628), .Z(n10600) );
  NBUFFX2 U10241 ( .INP(n10638), .Z(n10549) );
  NBUFFX2 U10242 ( .INP(n10627), .Z(n10608) );
  NBUFFX2 U10243 ( .INP(n10630), .Z(n10593) );
  NBUFFX2 U10244 ( .INP(n10638), .Z(n10551) );
  NBUFFX2 U10245 ( .INP(n10632), .Z(n10580) );
  NBUFFX2 U10246 ( .INP(n10631), .Z(n10585) );
  NBUFFX2 U10247 ( .INP(n10627), .Z(n10605) );
  NBUFFX2 U10248 ( .INP(n10627), .Z(n10607) );
  NBUFFX2 U10249 ( .INP(n10639), .Z(n10548) );
  NBUFFX2 U10250 ( .INP(n10633), .Z(n10577) );
  NBUFFX2 U10251 ( .INP(n10641), .Z(n10535) );
  NBUFFX2 U10252 ( .INP(n10630), .Z(n10592) );
  NBUFFX2 U10253 ( .INP(n10634), .Z(n10572) );
  NBUFFX2 U10254 ( .INP(n10633), .Z(n10578) );
  NBUFFX2 U10255 ( .INP(n10633), .Z(n10574) );
  NBUFFX2 U10256 ( .INP(n10637), .Z(n10557) );
  NBUFFX2 U10257 ( .INP(n10635), .Z(n10565) );
  NBUFFX2 U10258 ( .INP(n10628), .Z(n10602) );
  NBUFFX2 U10259 ( .INP(n10632), .Z(n10581) );
  NBUFFX2 U10260 ( .INP(n10638), .Z(n10553) );
  NBUFFX2 U10261 ( .INP(n10628), .Z(n10601) );
  NBUFFX2 U10262 ( .INP(n10632), .Z(n10579) );
  NBUFFX2 U10263 ( .INP(n10629), .Z(n10595) );
  NBUFFX2 U10264 ( .INP(n10643), .Z(n10526) );
  NBUFFX2 U10265 ( .INP(n10631), .Z(n10587) );
  NBUFFX2 U10266 ( .INP(n10642), .Z(n10531) );
  NBUFFX2 U10267 ( .INP(n10642), .Z(n10532) );
  NBUFFX2 U10268 ( .INP(n10630), .Z(n10590) );
  NBUFFX2 U10269 ( .INP(n10641), .Z(n10534) );
  NBUFFX2 U10270 ( .INP(n10642), .Z(n10529) );
  NBUFFX2 U10271 ( .INP(n10633), .Z(n10576) );
  NBUFFX2 U10272 ( .INP(n10644), .Z(n10521) );
  NBUFFX2 U10273 ( .INP(n10644), .Z(n10520) );
  NBUFFX2 U10274 ( .INP(n10629), .Z(n10596) );
  NBUFFX2 U10275 ( .INP(n10636), .Z(n10561) );
  NBUFFX2 U10276 ( .INP(n10629), .Z(n10598) );
  NBUFFX2 U10277 ( .INP(n10634), .Z(n10573) );
  NBUFFX2 U10278 ( .INP(n10634), .Z(n10571) );
  NBUFFX2 U10279 ( .INP(n10641), .Z(n10537) );
  NBUFFX2 U10280 ( .INP(n10640), .Z(n10543) );
  NBUFFX2 U10281 ( .INP(n10643), .Z(n10525) );
  NBUFFX2 U10282 ( .INP(n10644), .Z(n10523) );
  NBUFFX2 U10283 ( .INP(n10626), .Z(n10612) );
  NBUFFX2 U10284 ( .INP(n10626), .Z(n10611) );
  NBUFFX2 U10285 ( .INP(n10629), .Z(n10594) );
  NBUFFX2 U10286 ( .INP(n10640), .Z(n10539) );
  NBUFFX2 U10287 ( .INP(n10627), .Z(n10606) );
  NBUFFX2 U10288 ( .INP(n10638), .Z(n10550) );
  NBUFFX2 U10289 ( .INP(n10629), .Z(n10597) );
  NBUFFX2 U10290 ( .INP(n10635), .Z(n10568) );
  NBUFFX2 U10291 ( .INP(n10641), .Z(n10536) );
  NBUFFX2 U10292 ( .INP(n10631), .Z(n10584) );
  NBUFFX2 U10293 ( .INP(n10633), .Z(n10575) );
  NBUFFX2 U10294 ( .INP(n10636), .Z(n10559) );
  NBUFFX2 U10295 ( .INP(n10638), .Z(n10552) );
  NBUFFX2 U10296 ( .INP(n10625), .Z(n10615) );
  NBUFFX2 U10297 ( .INP(n10637), .Z(n10555) );
  NBUFFX2 U10298 ( .INP(n10272), .Z(n10270) );
  NBUFFX2 U10299 ( .INP(n10272), .Z(n10269) );
  NBUFFX2 U10300 ( .INP(n10272), .Z(n10268) );
  NBUFFX2 U10301 ( .INP(n10272), .Z(n10267) );
  NBUFFX2 U10302 ( .INP(n10624), .Z(n10622) );
  NBUFFX2 U10303 ( .INP(n10624), .Z(n10621) );
  NBUFFX2 U10304 ( .INP(n10624), .Z(n10620) );
  NBUFFX2 U10305 ( .INP(n10624), .Z(n10619) );
  NBUFFX2 U10306 ( .INP(n10272), .Z(n10271) );
  NBUFFX2 U10307 ( .INP(n10624), .Z(n10623) );
  NBUFFX2 U10308 ( .INP(n10301), .Z(n10272) );
  NBUFFX2 U10309 ( .INP(n10300), .Z(n10273) );
  NBUFFX2 U10310 ( .INP(n10300), .Z(n10274) );
  NBUFFX2 U10311 ( .INP(n10300), .Z(n10275) );
  NBUFFX2 U10312 ( .INP(n10299), .Z(n10276) );
  NBUFFX2 U10313 ( .INP(n10299), .Z(n10277) );
  NBUFFX2 U10315 ( .INP(n10299), .Z(n10278) );
  NBUFFX2 U10316 ( .INP(n10298), .Z(n10279) );
  NBUFFX2 U10317 ( .INP(n10298), .Z(n10280) );
  NBUFFX2 U10319 ( .INP(n10298), .Z(n10281) );
  NBUFFX2 U10320 ( .INP(n10297), .Z(n10282) );
  NBUFFX2 U10321 ( .INP(n10297), .Z(n10283) );
  NBUFFX2 U10322 ( .INP(n10297), .Z(n10284) );
  NBUFFX2 U10323 ( .INP(n10296), .Z(n10285) );
  NBUFFX2 U10324 ( .INP(n10296), .Z(n10286) );
  NBUFFX2 U10325 ( .INP(n10296), .Z(n10287) );
  NBUFFX2 U10326 ( .INP(n10295), .Z(n10288) );
  NBUFFX2 U10327 ( .INP(n10295), .Z(n10289) );
  NBUFFX2 U10328 ( .INP(n10295), .Z(n10290) );
  NBUFFX2 U10329 ( .INP(n10294), .Z(n10291) );
  NBUFFX2 U10330 ( .INP(n10294), .Z(n10292) );
  NBUFFX2 U10331 ( .INP(n10294), .Z(n10293) );
  NBUFFX2 U10332 ( .INP(n10304), .Z(n10294) );
  NBUFFX2 U10333 ( .INP(n10304), .Z(n10295) );
  NBUFFX2 U10334 ( .INP(n10303), .Z(n10296) );
  NBUFFX2 U10335 ( .INP(n10303), .Z(n10297) );
  NBUFFX2 U10336 ( .INP(n10303), .Z(n10298) );
  NBUFFX2 U10337 ( .INP(n10302), .Z(n10299) );
  NBUFFX2 U10338 ( .INP(n10302), .Z(n10300) );
  NBUFFX2 U10339 ( .INP(n10302), .Z(n10301) );
  NBUFFX2 U10340 ( .INP(test_se), .Z(n10302) );
  NBUFFX2 U10341 ( .INP(test_se), .Z(n10303) );
  NBUFFX2 U10342 ( .INP(test_se), .Z(n10304) );
  NBUFFX2 U10343 ( .INP(n10440), .Z(n10305) );
  NBUFFX2 U10344 ( .INP(n10440), .Z(n10306) );
  NBUFFX2 U10345 ( .INP(n10440), .Z(n10307) );
  NBUFFX2 U10346 ( .INP(n10439), .Z(n10308) );
  NBUFFX2 U10347 ( .INP(n10439), .Z(n10309) );
  NBUFFX2 U10348 ( .INP(n10439), .Z(n10310) );
  NBUFFX2 U10349 ( .INP(n10438), .Z(n10311) );
  NBUFFX2 U10350 ( .INP(n10438), .Z(n10312) );
  NBUFFX2 U10351 ( .INP(n10438), .Z(n10313) );
  NBUFFX2 U10352 ( .INP(n10437), .Z(n10314) );
  NBUFFX2 U10353 ( .INP(n10437), .Z(n10315) );
  NBUFFX2 U10354 ( .INP(n10437), .Z(n10316) );
  NBUFFX2 U10355 ( .INP(n10436), .Z(n10317) );
  NBUFFX2 U10356 ( .INP(n10436), .Z(n10318) );
  NBUFFX2 U10357 ( .INP(n10436), .Z(n10319) );
  NBUFFX2 U10358 ( .INP(n10435), .Z(n10320) );
  NBUFFX2 U10359 ( .INP(n10435), .Z(n10321) );
  NBUFFX2 U10360 ( .INP(n10435), .Z(n10322) );
  NBUFFX2 U10361 ( .INP(n10434), .Z(n10323) );
  NBUFFX2 U10362 ( .INP(n10434), .Z(n10324) );
  NBUFFX2 U10363 ( .INP(n10434), .Z(n10325) );
  NBUFFX2 U10364 ( .INP(n10433), .Z(n10326) );
  NBUFFX2 U10365 ( .INP(n10433), .Z(n10327) );
  NBUFFX2 U10366 ( .INP(n10433), .Z(n10328) );
  NBUFFX2 U10367 ( .INP(n10432), .Z(n10329) );
  NBUFFX2 U10368 ( .INP(n10432), .Z(n10330) );
  NBUFFX2 U10369 ( .INP(n10432), .Z(n10331) );
  NBUFFX2 U10370 ( .INP(n10431), .Z(n10332) );
  NBUFFX2 U10371 ( .INP(n10431), .Z(n10333) );
  NBUFFX2 U10372 ( .INP(n10431), .Z(n10334) );
  NBUFFX2 U10373 ( .INP(n10430), .Z(n10335) );
  NBUFFX2 U10374 ( .INP(n10430), .Z(n10336) );
  NBUFFX2 U10375 ( .INP(n10430), .Z(n10337) );
  NBUFFX2 U10376 ( .INP(n10429), .Z(n10338) );
  NBUFFX2 U10377 ( .INP(n10429), .Z(n10339) );
  NBUFFX2 U10378 ( .INP(n10429), .Z(n10340) );
  NBUFFX2 U10379 ( .INP(n10428), .Z(n10341) );
  NBUFFX2 U10380 ( .INP(n10428), .Z(n10342) );
  NBUFFX2 U10381 ( .INP(n10428), .Z(n10343) );
  NBUFFX2 U10382 ( .INP(n10427), .Z(n10344) );
  NBUFFX2 U10383 ( .INP(n10427), .Z(n10345) );
  NBUFFX2 U10384 ( .INP(n10427), .Z(n10346) );
  NBUFFX2 U10385 ( .INP(n10426), .Z(n10347) );
  NBUFFX2 U10386 ( .INP(n10426), .Z(n10348) );
  NBUFFX2 U10387 ( .INP(n10426), .Z(n10349) );
  NBUFFX2 U10388 ( .INP(n10425), .Z(n10350) );
  NBUFFX2 U10389 ( .INP(n10425), .Z(n10351) );
  NBUFFX2 U10390 ( .INP(n10425), .Z(n10352) );
  NBUFFX2 U10391 ( .INP(n10424), .Z(n10353) );
  NBUFFX2 U10392 ( .INP(n10424), .Z(n10354) );
  NBUFFX2 U10393 ( .INP(n10424), .Z(n10355) );
  NBUFFX2 U10394 ( .INP(n10423), .Z(n10356) );
  NBUFFX2 U10395 ( .INP(n10423), .Z(n10357) );
  NBUFFX2 U10396 ( .INP(n10423), .Z(n10358) );
  NBUFFX2 U10397 ( .INP(n10422), .Z(n10359) );
  NBUFFX2 U10398 ( .INP(n10422), .Z(n10360) );
  NBUFFX2 U10399 ( .INP(n10422), .Z(n10361) );
  NBUFFX2 U10400 ( .INP(n10421), .Z(n10362) );
  NBUFFX2 U10401 ( .INP(n10421), .Z(n10363) );
  NBUFFX2 U10402 ( .INP(n10421), .Z(n10364) );
  NBUFFX2 U10403 ( .INP(n10420), .Z(n10365) );
  NBUFFX2 U10404 ( .INP(n10420), .Z(n10366) );
  NBUFFX2 U10405 ( .INP(n10420), .Z(n10367) );
  NBUFFX2 U10406 ( .INP(n10419), .Z(n10368) );
  NBUFFX2 U10407 ( .INP(n10419), .Z(n10369) );
  NBUFFX2 U10408 ( .INP(n10419), .Z(n10370) );
  NBUFFX2 U10409 ( .INP(n10418), .Z(n10371) );
  NBUFFX2 U10410 ( .INP(n10418), .Z(n10372) );
  NBUFFX2 U10411 ( .INP(n10418), .Z(n10373) );
  NBUFFX2 U10412 ( .INP(n10417), .Z(n10374) );
  NBUFFX2 U10413 ( .INP(n10417), .Z(n10375) );
  NBUFFX2 U10414 ( .INP(n10417), .Z(n10376) );
  NBUFFX2 U10415 ( .INP(n10416), .Z(n10377) );
  NBUFFX2 U10416 ( .INP(n10416), .Z(n10378) );
  NBUFFX2 U10417 ( .INP(n10416), .Z(n10379) );
  NBUFFX2 U10418 ( .INP(n10415), .Z(n10380) );
  NBUFFX2 U10419 ( .INP(n10415), .Z(n10381) );
  NBUFFX2 U10420 ( .INP(n10415), .Z(n10382) );
  NBUFFX2 U10421 ( .INP(n10414), .Z(n10383) );
  NBUFFX2 U10422 ( .INP(n10414), .Z(n10384) );
  NBUFFX2 U10423 ( .INP(n10414), .Z(n10385) );
  NBUFFX2 U10424 ( .INP(n10413), .Z(n10386) );
  NBUFFX2 U10425 ( .INP(n10413), .Z(n10387) );
  NBUFFX2 U10426 ( .INP(n10413), .Z(n10388) );
  NBUFFX2 U10427 ( .INP(n10412), .Z(n10389) );
  NBUFFX2 U10428 ( .INP(n10412), .Z(n10390) );
  NBUFFX2 U10429 ( .INP(n10412), .Z(n10391) );
  NBUFFX2 U10430 ( .INP(n10411), .Z(n10392) );
  NBUFFX2 U10431 ( .INP(n10411), .Z(n10393) );
  NBUFFX2 U10432 ( .INP(n10411), .Z(n10394) );
  NBUFFX2 U10433 ( .INP(n10410), .Z(n10395) );
  NBUFFX2 U10434 ( .INP(n10410), .Z(n10396) );
  NBUFFX2 U10435 ( .INP(n10410), .Z(n10397) );
  NBUFFX2 U10436 ( .INP(n10409), .Z(n10398) );
  NBUFFX2 U10437 ( .INP(n10409), .Z(n10399) );
  NBUFFX2 U10438 ( .INP(n10409), .Z(n10400) );
  NBUFFX2 U10439 ( .INP(n10408), .Z(n10401) );
  NBUFFX2 U10440 ( .INP(n10408), .Z(n10402) );
  NBUFFX2 U10441 ( .INP(n10408), .Z(n10403) );
  NBUFFX2 U10442 ( .INP(n10407), .Z(n10404) );
  NBUFFX2 U10443 ( .INP(n10407), .Z(n10405) );
  NBUFFX2 U10444 ( .INP(n10407), .Z(n10406) );
  NBUFFX2 U10445 ( .INP(n10452), .Z(n10407) );
  NBUFFX2 U10446 ( .INP(n10451), .Z(n10408) );
  NBUFFX2 U10447 ( .INP(n10451), .Z(n10409) );
  NBUFFX2 U10448 ( .INP(n10451), .Z(n10410) );
  NBUFFX2 U10449 ( .INP(n10450), .Z(n10411) );
  NBUFFX2 U10450 ( .INP(n10450), .Z(n10412) );
  NBUFFX2 U10451 ( .INP(n10450), .Z(n10413) );
  NBUFFX2 U10452 ( .INP(n10449), .Z(n10414) );
  NBUFFX2 U10453 ( .INP(n10449), .Z(n10415) );
  NBUFFX2 U10454 ( .INP(n10449), .Z(n10416) );
  NBUFFX2 U10455 ( .INP(n10448), .Z(n10417) );
  NBUFFX2 U10456 ( .INP(n10448), .Z(n10418) );
  NBUFFX2 U10457 ( .INP(n10448), .Z(n10419) );
  NBUFFX2 U10458 ( .INP(n10447), .Z(n10420) );
  NBUFFX2 U10459 ( .INP(n10447), .Z(n10421) );
  NBUFFX2 U10460 ( .INP(n10447), .Z(n10422) );
  NBUFFX2 U10461 ( .INP(n10446), .Z(n10423) );
  NBUFFX2 U10462 ( .INP(n10446), .Z(n10424) );
  NBUFFX2 U10463 ( .INP(n10446), .Z(n10425) );
  NBUFFX2 U10464 ( .INP(n10445), .Z(n10426) );
  NBUFFX2 U10465 ( .INP(n10445), .Z(n10427) );
  NBUFFX2 U10466 ( .INP(n10445), .Z(n10428) );
  NBUFFX2 U10467 ( .INP(n10444), .Z(n10429) );
  NBUFFX2 U10468 ( .INP(n10444), .Z(n10430) );
  NBUFFX2 U10469 ( .INP(n10444), .Z(n10431) );
  NBUFFX2 U10470 ( .INP(n10443), .Z(n10432) );
  NBUFFX2 U10471 ( .INP(n10443), .Z(n10433) );
  NBUFFX2 U10472 ( .INP(n10443), .Z(n10434) );
  NBUFFX2 U10473 ( .INP(n10442), .Z(n10435) );
  NBUFFX2 U10474 ( .INP(n10442), .Z(n10436) );
  NBUFFX2 U10475 ( .INP(n10442), .Z(n10437) );
  NBUFFX2 U10476 ( .INP(n10441), .Z(n10438) );
  NBUFFX2 U10477 ( .INP(n10441), .Z(n10439) );
  NBUFFX2 U10478 ( .INP(n10441), .Z(n10440) );
  NBUFFX2 U10479 ( .INP(n10456), .Z(n10441) );
  NBUFFX2 U10480 ( .INP(n10456), .Z(n10442) );
  NBUFFX2 U10481 ( .INP(n10456), .Z(n10443) );
  NBUFFX2 U10482 ( .INP(n10455), .Z(n10444) );
  NBUFFX2 U10483 ( .INP(n10455), .Z(n10445) );
  NBUFFX2 U10484 ( .INP(n10455), .Z(n10446) );
  NBUFFX2 U10485 ( .INP(n10454), .Z(n10447) );
  NBUFFX2 U10486 ( .INP(n10454), .Z(n10448) );
  NBUFFX2 U10487 ( .INP(n10454), .Z(n10449) );
  NBUFFX2 U10488 ( .INP(n10453), .Z(n10450) );
  NBUFFX2 U10489 ( .INP(n10453), .Z(n10451) );
  NBUFFX2 U10490 ( .INP(n10453), .Z(n10452) );
  NBUFFX2 U10491 ( .INP(g35), .Z(n10453) );
  NBUFFX2 U10492 ( .INP(g35), .Z(n10454) );
  NBUFFX2 U10493 ( .INP(g35), .Z(n10455) );
  NBUFFX2 U10494 ( .INP(g35), .Z(n10456) );
  INVX0 U10495 ( .INP(n10359), .ZN(n10457) );
  INVX0 U10496 ( .INP(n10359), .ZN(n10458) );
  INVX0 U10497 ( .INP(n10358), .ZN(n10459) );
  INVX0 U10498 ( .INP(n10359), .ZN(n10460) );
  INVX0 U10499 ( .INP(n10360), .ZN(n10461) );
  INVX0 U10500 ( .INP(n10359), .ZN(n10462) );
  INVX0 U10501 ( .INP(n10360), .ZN(n10463) );
  INVX0 U10502 ( .INP(n10359), .ZN(n10464) );
  INVX0 U10503 ( .INP(n10360), .ZN(n10465) );
  INVX0 U10504 ( .INP(n10359), .ZN(n10466) );
  INVX0 U10505 ( .INP(n10359), .ZN(n10467) );
  INVX0 U10506 ( .INP(n10360), .ZN(n10468) );
  INVX0 U10507 ( .INP(n10360), .ZN(n10469) );
  INVX0 U10508 ( .INP(n10361), .ZN(n10470) );
  INVX0 U10509 ( .INP(n10360), .ZN(n10471) );
  INVX0 U10510 ( .INP(n10361), .ZN(n10472) );
  INVX0 U10511 ( .INP(n10360), .ZN(n10473) );
  INVX0 U10512 ( .INP(n10361), .ZN(n10474) );
  INVX0 U10513 ( .INP(n10360), .ZN(n10475) );
  INVX0 U10514 ( .INP(n10359), .ZN(n10476) );
  INVX0 U10515 ( .INP(n10361), .ZN(n10477) );
  INVX0 U10516 ( .INP(n10362), .ZN(n10478) );
  INVX0 U10517 ( .INP(n10360), .ZN(n10479) );
  INVX0 U10518 ( .INP(n10358), .ZN(n10480) );
  INVX0 U10519 ( .INP(n10362), .ZN(n10481) );
  INVX0 U10520 ( .INP(n10361), .ZN(n10482) );
  INVX0 U10521 ( .INP(n10362), .ZN(n10483) );
  INVX0 U10522 ( .INP(n10359), .ZN(n10484) );
  INVX0 U10523 ( .INP(n10361), .ZN(n10485) );
  INVX0 U10524 ( .INP(n10362), .ZN(n10486) );
  INVX0 U10525 ( .INP(n10362), .ZN(n10487) );
  INVX0 U10526 ( .INP(n10362), .ZN(n10488) );
  INVX0 U10527 ( .INP(n10363), .ZN(n10489) );
  INVX0 U10528 ( .INP(n10362), .ZN(n10490) );
  INVX0 U10529 ( .INP(n10363), .ZN(n10491) );
  INVX0 U10530 ( .INP(n10361), .ZN(n10492) );
  INVX0 U10531 ( .INP(n10363), .ZN(n10493) );
  INVX0 U10532 ( .INP(n10363), .ZN(n10494) );
  INVX0 U10533 ( .INP(n10364), .ZN(n10495) );
  INVX0 U10534 ( .INP(n10363), .ZN(n10496) );
  INVX0 U10535 ( .INP(n10364), .ZN(n10497) );
  INVX0 U10536 ( .INP(n10361), .ZN(n10498) );
  INVX0 U10537 ( .INP(n10364), .ZN(n10499) );
  INVX0 U10538 ( .INP(n10363), .ZN(n10500) );
  INVX0 U10539 ( .INP(n10361), .ZN(n10501) );
  INVX0 U10540 ( .INP(n10363), .ZN(n10502) );
  INVX0 U10541 ( .INP(n10364), .ZN(n10503) );
  INVX0 U10542 ( .INP(n10362), .ZN(n10504) );
  INVX0 U10543 ( .INP(n10364), .ZN(n10505) );
  INVX0 U10544 ( .INP(n10363), .ZN(n10506) );
  INVX0 U10545 ( .INP(n10364), .ZN(n10507) );
  INVX0 U10546 ( .INP(n10363), .ZN(n10508) );
  INVX0 U10547 ( .INP(n10364), .ZN(n10509) );
  INVX0 U10548 ( .INP(n10362), .ZN(n10510) );
  INVX0 U10549 ( .INP(n10365), .ZN(n10511) );
  INVX0 U10550 ( .INP(n10364), .ZN(n10512) );
  INVX0 U10551 ( .INP(n10365), .ZN(n10513) );
  INVX0 U10552 ( .INP(n10364), .ZN(n10514) );
  INVX0 U10553 ( .INP(n10365), .ZN(n10515) );
  INVX0 U10554 ( .INP(n10358), .ZN(n10516) );
  NBUFFX2 U10555 ( .INP(n10653), .Z(n10624) );
  NBUFFX2 U10556 ( .INP(n10652), .Z(n10625) );
  NBUFFX2 U10557 ( .INP(n10652), .Z(n10626) );
  NBUFFX2 U10558 ( .INP(n10652), .Z(n10627) );
  NBUFFX2 U10559 ( .INP(n10651), .Z(n10628) );
  NBUFFX2 U10560 ( .INP(n10651), .Z(n10629) );
  NBUFFX2 U10561 ( .INP(n10651), .Z(n10630) );
  NBUFFX2 U10562 ( .INP(n10650), .Z(n10631) );
  NBUFFX2 U10563 ( .INP(n10650), .Z(n10632) );
  NBUFFX2 U10564 ( .INP(n10650), .Z(n10633) );
  NBUFFX2 U10565 ( .INP(n10649), .Z(n10634) );
  NBUFFX2 U10566 ( .INP(n10649), .Z(n10635) );
  NBUFFX2 U10567 ( .INP(n10649), .Z(n10636) );
  NBUFFX2 U10568 ( .INP(n10648), .Z(n10637) );
  NBUFFX2 U10569 ( .INP(n10648), .Z(n10638) );
  NBUFFX2 U10570 ( .INP(n10648), .Z(n10639) );
  NBUFFX2 U10571 ( .INP(n10647), .Z(n10640) );
  NBUFFX2 U10572 ( .INP(n10647), .Z(n10641) );
  NBUFFX2 U10573 ( .INP(n10647), .Z(n10642) );
  NBUFFX2 U10574 ( .INP(n10646), .Z(n10643) );
  NBUFFX2 U10575 ( .INP(n10646), .Z(n10644) );
  NBUFFX2 U10576 ( .INP(n10646), .Z(n10645) );
  NBUFFX2 U10577 ( .INP(n10656), .Z(n10646) );
  NBUFFX2 U10578 ( .INP(n10656), .Z(n10647) );
  NBUFFX2 U10579 ( .INP(n10655), .Z(n10648) );
  NBUFFX2 U10580 ( .INP(n10655), .Z(n10649) );
  NBUFFX2 U10581 ( .INP(n10655), .Z(n10650) );
  NBUFFX2 U10582 ( .INP(n10654), .Z(n10651) );
  NBUFFX2 U10583 ( .INP(n10654), .Z(n10652) );
  NBUFFX2 U10584 ( .INP(n10654), .Z(n10653) );
  NBUFFX2 U10585 ( .INP(CK), .Z(n10654) );
  NBUFFX2 U10586 ( .INP(CK), .Z(n10655) );
  NBUFFX2 U10587 ( .INP(CK), .Z(n10656) );
  NAND2X0 U10588 ( .IN1(n10657), .IN2(n10658), .QN(n5961) );
  NOR2X0 U10589 ( .IN1(n10659), .IN2(n10660), .QN(n10658) );
  AND2X1 U10590 ( .IN1(n10661), .IN2(n10039), .Q(n10660) );
  NOR2X0 U10591 ( .IN1(n10039), .IN2(n10662), .QN(n10659) );
  NOR2X0 U10592 ( .IN1(n10663), .IN2(n10664), .QN(n10657) );
  AND2X1 U10593 ( .IN1(n10665), .IN2(n10038), .Q(n10664) );
  NOR2X0 U10594 ( .IN1(n10038), .IN2(n10666), .QN(n10663) );
  NAND2X0 U10595 ( .IN1(n10667), .IN2(n10668), .QN(n5960) );
  NOR2X0 U10596 ( .IN1(n10669), .IN2(n10670), .QN(n10668) );
  AND2X1 U10597 ( .IN1(n10671), .IN2(n10037), .Q(n10670) );
  NOR2X0 U10598 ( .IN1(n10037), .IN2(n10672), .QN(n10669) );
  NOR2X0 U10599 ( .IN1(n10673), .IN2(n10674), .QN(n10667) );
  AND2X1 U10600 ( .IN1(n10675), .IN2(n10036), .Q(n10674) );
  NOR2X0 U10601 ( .IN1(n10036), .IN2(n10676), .QN(n10673) );
  INVX0 U10602 ( .INP(n10677), .ZN(n490) );
  NAND2X0 U10603 ( .IN1(n10678), .IN2(g1677), .QN(n4459) );
  NAND2X0 U10604 ( .IN1(n10679), .IN2(g1811), .QN(n4448) );
  NAND2X0 U10605 ( .IN1(test_so53), .IN2(n10680), .QN(n4437) );
  OR2X1 U10606 ( .IN1(n10681), .IN2(n9829), .Q(n4426) );
  NAND2X0 U10607 ( .IN1(n10682), .IN2(g2236), .QN(n4415) );
  NAND2X0 U10608 ( .IN1(n10683), .IN2(g2370), .QN(n4403) );
  NAND2X0 U10609 ( .IN1(n10684), .IN2(g2504), .QN(n4392) );
  NAND2X0 U10610 ( .IN1(n10685), .IN2(g2638), .QN(n4380) );
  NAND2X0 U10611 ( .IN1(n10686), .IN2(n10687), .QN(n4305) );
  NOR2X0 U10612 ( .IN1(n10688), .IN2(n10689), .QN(n10687) );
  NOR2X0 U10613 ( .IN1(n5440), .IN2(g4821), .QN(n10689) );
  NOR2X0 U10614 ( .IN1(n9668), .IN2(n10040), .QN(n10688) );
  NOR2X0 U10615 ( .IN1(n10690), .IN2(n10691), .QN(n10686) );
  NAND2X0 U10616 ( .IN1(n10692), .IN2(n10693), .QN(n10691) );
  NAND2X0 U10617 ( .IN1(n10694), .IN2(n5712), .QN(n10693) );
  NOR2X0 U10618 ( .IN1(n10695), .IN2(n10696), .QN(n10694) );
  NAND2X0 U10619 ( .IN1(n5656), .IN2(n5440), .QN(n10696) );
  NAND2X0 U10620 ( .IN1(n10040), .IN2(n10697), .QN(n10695) );
  NAND2X0 U10621 ( .IN1(n10698), .IN2(n10699), .QN(n10697) );
  NAND2X0 U10622 ( .IN1(n10700), .IN2(n10701), .QN(n10698) );
  NAND2X0 U10623 ( .IN1(n10702), .IN2(g4776), .QN(n10701) );
  NAND2X0 U10624 ( .IN1(n5368), .IN2(n10703), .QN(n10702) );
  XNOR2X1 U10625 ( .IN1(g34657), .IN2(n10704), .Q(n10703) );
  NOR2X0 U10626 ( .IN1(n10705), .IN2(n10706), .QN(n10704) );
  NAND2X0 U10627 ( .IN1(n10707), .IN2(n10708), .QN(n10706) );
  NAND2X0 U10628 ( .IN1(n10709), .IN2(g4727), .QN(n10708) );
  OR2X1 U10629 ( .IN1(n10710), .IN2(n5345), .Q(n10707) );
  NAND2X0 U10630 ( .IN1(n10711), .IN2(n10712), .QN(n10705) );
  OR2X1 U10631 ( .IN1(n10713), .IN2(n5296), .Q(n10712) );
  OR2X1 U10632 ( .IN1(n10714), .IN2(n5344), .Q(n10711) );
  NOR2X0 U10633 ( .IN1(n10715), .IN2(n10716), .QN(n10700) );
  NOR2X0 U10634 ( .IN1(n10717), .IN2(g4793), .QN(n10716) );
  NOR2X0 U10635 ( .IN1(n10718), .IN2(test_so29), .QN(n10717) );
  NOR2X0 U10636 ( .IN1(n10719), .IN2(n10720), .QN(n10718) );
  NAND2X0 U10637 ( .IN1(n5707), .IN2(n10721), .QN(n10720) );
  NAND2X0 U10638 ( .IN1(n5867), .IN2(n10709), .QN(n10721) );
  NAND2X0 U10639 ( .IN1(n10713), .IN2(n10714), .QN(n10719) );
  NOR2X0 U10640 ( .IN1(n5368), .IN2(g34657), .QN(n10715) );
  NAND2X0 U10641 ( .IN1(g4646), .IN2(g29220), .QN(n10692) );
  NOR2X0 U10642 ( .IN1(n5656), .IN2(g4826), .QN(n10690) );
  NAND2X0 U10643 ( .IN1(n10722), .IN2(n10723), .QN(n4283) );
  NOR2X0 U10644 ( .IN1(n10724), .IN2(n10725), .QN(n10723) );
  NOR2X0 U10645 ( .IN1(n5881), .IN2(n5443), .QN(n10725) );
  NOR2X0 U10646 ( .IN1(n5318), .IN2(g3333), .QN(n10724) );
  NOR2X0 U10647 ( .IN1(n10726), .IN2(n10727), .QN(n10722) );
  NAND2X0 U10648 ( .IN1(n10728), .IN2(n10729), .QN(n10727) );
  NAND2X0 U10649 ( .IN1(n9671), .IN2(g4878), .QN(n10729) );
  NAND2X0 U10650 ( .IN1(n10730), .IN2(n5283), .QN(n10728) );
  NOR2X0 U10651 ( .IN1(n10731), .IN2(n10732), .QN(n10730) );
  NOR2X0 U10652 ( .IN1(n10733), .IN2(n10734), .QN(n10731) );
  NOR2X0 U10653 ( .IN1(n10735), .IN2(n10736), .QN(n10734) );
  NAND2X0 U10654 ( .IN1(n10737), .IN2(n10738), .QN(n10736) );
  OR2X1 U10655 ( .IN1(g34649), .IN2(n5367), .Q(n10738) );
  NAND2X0 U10656 ( .IN1(n5367), .IN2(n10739), .QN(n10737) );
  NAND2X0 U10657 ( .IN1(n10123), .IN2(n10740), .QN(n10739) );
  NAND2X0 U10658 ( .IN1(n10741), .IN2(n10742), .QN(n10740) );
  AND2X1 U10659 ( .IN1(n10743), .IN2(n10744), .Q(n10742) );
  NOR2X0 U10660 ( .IN1(n10745), .IN2(g4966), .QN(n10741) );
  NOR2X0 U10661 ( .IN1(n10746), .IN2(g4927), .QN(n10745) );
  NOR2X0 U10662 ( .IN1(n5706), .IN2(n10747), .QN(n10735) );
  NOR2X0 U10663 ( .IN1(n10748), .IN2(g4983), .QN(n10747) );
  XNOR2X1 U10664 ( .IN1(n10749), .IN2(g34649), .Q(n10748) );
  NAND2X0 U10665 ( .IN1(n10750), .IN2(n10751), .QN(n10749) );
  NOR2X0 U10666 ( .IN1(n10752), .IN2(n10753), .QN(n10751) );
  NOR2X0 U10667 ( .IN1(n5408), .IN2(n10746), .QN(n10753) );
  NOR2X0 U10668 ( .IN1(n5297), .IN2(n10754), .QN(n10752) );
  NOR2X0 U10669 ( .IN1(n10755), .IN2(n10756), .QN(n10750) );
  NOR2X0 U10670 ( .IN1(n5295), .IN2(n10743), .QN(n10756) );
  NOR2X0 U10671 ( .IN1(n5346), .IN2(n10744), .QN(n10755) );
  INVX0 U10672 ( .INP(n10757), .ZN(n10733) );
  NOR2X0 U10673 ( .IN1(n9669), .IN2(n5713), .QN(n10726) );
  INVX0 U10674 ( .INP(n10758), .ZN(n4198) );
  NOR2X0 U10675 ( .IN1(g3167), .IN2(n10759), .QN(n4034) );
  NAND2X0 U10676 ( .IN1(n5366), .IN2(n10062), .QN(n10759) );
  NOR2X0 U10677 ( .IN1(g3518), .IN2(n10760), .QN(n4002) );
  NAND2X0 U10678 ( .IN1(n5576), .IN2(n10058), .QN(n10760) );
  NOR2X0 U10679 ( .IN1(g3857), .IN2(n10761), .QN(n3969) );
  OR2X1 U10680 ( .IN1(g3863), .IN2(test_so33), .Q(n10761) );
  NOR2X0 U10681 ( .IN1(n10762), .IN2(n10763), .QN(n3933) );
  NAND2X0 U10682 ( .IN1(n2760), .IN2(g43), .QN(n10762) );
  NOR2X0 U10683 ( .IN1(g5176), .IN2(n10764), .QN(n3926) );
  NAND2X0 U10684 ( .IN1(n5570), .IN2(n10052), .QN(n10764) );
  INVX0 U10685 ( .INP(n10765), .ZN(n39) );
  NOR2X0 U10686 ( .IN1(g5523), .IN2(n10766), .QN(n3893) );
  NAND2X0 U10687 ( .IN1(n5575), .IN2(n10057), .QN(n10766) );
  NOR2X0 U10688 ( .IN1(g5869), .IN2(n10767), .QN(n3860) );
  NAND2X0 U10689 ( .IN1(n5573), .IN2(n10055), .QN(n10767) );
  NOR2X0 U10690 ( .IN1(g6215), .IN2(n10768), .QN(n3826) );
  NAND2X0 U10691 ( .IN1(n5574), .IN2(n10056), .QN(n10768) );
  NOR2X0 U10692 ( .IN1(g6561), .IN2(n10769), .QN(n3792) );
  NAND2X0 U10693 ( .IN1(n5571), .IN2(n10053), .QN(n10769) );
  INVX0 U10694 ( .INP(n10770), .ZN(n3743) );
  NAND2X0 U10695 ( .IN1(n10771), .IN2(n10772), .QN(n3675) );
  NOR2X0 U10696 ( .IN1(n10773), .IN2(n10774), .QN(n10772) );
  NOR2X0 U10697 ( .IN1(n9778), .IN2(n10775), .QN(n10774) );
  NOR2X0 U10698 ( .IN1(g441), .IN2(n10776), .QN(n10775) );
  XOR2X1 U10699 ( .IN1(test_so72), .IN2(n9914), .Q(n10776) );
  NOR2X0 U10700 ( .IN1(n10777), .IN2(g392), .QN(n10773) );
  NOR2X0 U10701 ( .IN1(g411), .IN2(n10778), .QN(n10777) );
  XOR2X1 U10702 ( .IN1(test_so72), .IN2(n5402), .Q(n10778) );
  NOR2X0 U10703 ( .IN1(g691), .IN2(g417), .QN(n10771) );
  NAND2X0 U10704 ( .IN1(n10779), .IN2(n5516), .QN(n3635) );
  NOR2X0 U10705 ( .IN1(test_so30), .IN2(n5349), .QN(n10779) );
  INVX0 U10706 ( .INP(n10780), .ZN(n36) );
  NOR2X0 U10707 ( .IN1(n10781), .IN2(n10782), .QN(n3174) );
  XOR2X1 U10708 ( .IN1(n5820), .IN2(n10783), .Q(n10782) );
  XOR2X1 U10709 ( .IN1(n5708), .IN2(n10784), .Q(n10781) );
  NOR2X0 U10710 ( .IN1(n1289), .IN2(n6010), .QN(n3084) );
  NAND2X0 U10711 ( .IN1(n10785), .IN2(n10786), .QN(n3065) );
  NAND2X0 U10712 ( .IN1(n10787), .IN2(g4108), .QN(n10786) );
  NOR2X0 U10713 ( .IN1(n9913), .IN2(n10463), .QN(n10785) );
  INVX0 U10714 ( .INP(n10788), .ZN(n3) );
  XOR2X1 U10715 ( .IN1(n5323), .IN2(n2607), .Q(n2608) );
  INVX0 U10716 ( .INP(n10789), .ZN(n2601) );
  NAND2X0 U10717 ( .IN1(n10790), .IN2(g34979), .QN(n2461) );
  NOR2X0 U10718 ( .IN1(n10791), .IN2(n10792), .QN(n2396) );
  INVX0 U10719 ( .INP(n10793), .ZN(n195) );
  NOR2X0 U10720 ( .IN1(n10794), .IN2(n10763), .QN(n10105) );
  NAND2X0 U10721 ( .IN1(n10795), .IN2(n10796), .QN(n10763) );
  NAND2X0 U10722 ( .IN1(n10797), .IN2(n10798), .QN(g34980) );
  NAND2X0 U10723 ( .IN1(test_so14), .IN2(n10515), .QN(n10798) );
  NAND2X0 U10724 ( .IN1(n10799), .IN2(n10378), .QN(n10797) );
  NAND2X0 U10725 ( .IN1(n5842), .IN2(n10800), .QN(n10799) );
  NAND2X0 U10726 ( .IN1(n10801), .IN2(n10802), .QN(n10800) );
  NOR2X0 U10727 ( .IN1(g56), .IN2(g54), .QN(n10802) );
  NOR2X0 U10728 ( .IN1(g53), .IN2(n10803), .QN(n10801) );
  NAND2X0 U10729 ( .IN1(n10803), .IN2(g22), .QN(g34972) );
  INVX0 U10730 ( .INP(n10104), .ZN(n10803) );
  XOR2X1 U10731 ( .IN1(n10804), .IN2(n10805), .Q(n10104) );
  XOR2X1 U10732 ( .IN1(g34978), .IN2(g34977), .Q(n10805) );
  XNOR2X1 U10733 ( .IN1(n10806), .IN2(g34970), .Q(n10804) );
  XOR2X1 U10734 ( .IN1(n10807), .IN2(n10808), .Q(n10806) );
  XNOR2X1 U10735 ( .IN1(g34975), .IN2(n10809), .Q(n10808) );
  XOR2X1 U10736 ( .IN1(g34974), .IN2(g34976), .Q(n10809) );
  XOR2X1 U10737 ( .IN1(g34971), .IN2(n10810), .Q(n10807) );
  XOR2X1 U10738 ( .IN1(n10811), .IN2(g34979), .Q(n10810) );
  NAND2X0 U10739 ( .IN1(n10812), .IN2(g55), .QN(n10811) );
  OR2X1 U10740 ( .IN1(g34979), .IN2(n9723), .Q(g34927) );
  NAND2X0 U10741 ( .IN1(n10813), .IN2(n10814), .QN(g34979) );
  NOR2X0 U10742 ( .IN1(n10815), .IN2(n10816), .QN(n10814) );
  OR2X1 U10743 ( .IN1(n10817), .IN2(n10818), .Q(n10816) );
  NOR2X0 U10744 ( .IN1(n5635), .IN2(n10819), .QN(n10818) );
  NOR2X0 U10745 ( .IN1(n10820), .IN2(n10821), .QN(n10817) );
  NOR2X0 U10746 ( .IN1(n10822), .IN2(n10823), .QN(n10820) );
  NAND2X0 U10747 ( .IN1(n10824), .IN2(n10825), .QN(n10823) );
  NOR2X0 U10748 ( .IN1(n10826), .IN2(n10827), .QN(n10825) );
  NAND2X0 U10749 ( .IN1(n10828), .IN2(n10829), .QN(n10827) );
  NAND2X0 U10750 ( .IN1(n10830), .IN2(g568), .QN(n10829) );
  NAND2X0 U10751 ( .IN1(n10831), .IN2(g744), .QN(n10828) );
  NOR2X0 U10752 ( .IN1(n10079), .IN2(n10832), .QN(n10826) );
  NOR2X0 U10753 ( .IN1(n10833), .IN2(n10834), .QN(n10824) );
  NAND2X0 U10754 ( .IN1(n10835), .IN2(n10836), .QN(n10834) );
  NAND2X0 U10755 ( .IN1(n10837), .IN2(g2886), .QN(n10836) );
  OR2X1 U10756 ( .IN1(n10838), .IN2(n5750), .Q(n10835) );
  NOR2X0 U10757 ( .IN1(n5981), .IN2(n10839), .QN(n10833) );
  NAND2X0 U10758 ( .IN1(n10840), .IN2(n10841), .QN(n10822) );
  NOR2X0 U10759 ( .IN1(n10842), .IN2(n10843), .QN(n10841) );
  NAND2X0 U10760 ( .IN1(n10844), .IN2(n10845), .QN(n10843) );
  NAND2X0 U10761 ( .IN1(g92), .IN2(n10846), .QN(n10845) );
  NAND2X0 U10762 ( .IN1(g127), .IN2(n10847), .QN(n10844) );
  AND2X1 U10763 ( .IN1(n10790), .IN2(test_so14), .Q(n10842) );
  NOR2X0 U10764 ( .IN1(n10848), .IN2(n10849), .QN(n10840) );
  NAND2X0 U10765 ( .IN1(n10850), .IN2(n10851), .QN(n10849) );
  NAND2X0 U10766 ( .IN1(n10852), .IN2(g785), .QN(n10851) );
  NAND2X0 U10767 ( .IN1(g29221), .IN2(n10853), .QN(n10850) );
  NOR2X0 U10768 ( .IN1(n5473), .IN2(n10854), .QN(n10848) );
  NAND2X0 U10769 ( .IN1(n10855), .IN2(n10856), .QN(n10815) );
  NAND2X0 U10770 ( .IN1(test_so67), .IN2(n10857), .QN(n10855) );
  NOR2X0 U10771 ( .IN1(n10858), .IN2(n10859), .QN(n10813) );
  NAND2X0 U10772 ( .IN1(n10860), .IN2(n10861), .QN(n10859) );
  NAND2X0 U10773 ( .IN1(n10862), .IN2(g2138), .QN(n10861) );
  NAND2X0 U10774 ( .IN1(n10863), .IN2(g2697), .QN(n10860) );
  NAND2X0 U10775 ( .IN1(n10864), .IN2(n10865), .QN(n10858) );
  NAND2X0 U10776 ( .IN1(n10866), .IN2(g939), .QN(n10865) );
  NAND2X0 U10777 ( .IN1(n10867), .IN2(n9332), .QN(n10864) );
  OR2X1 U10778 ( .IN1(g34978), .IN2(n9723), .Q(g34925) );
  NAND2X0 U10779 ( .IN1(n10868), .IN2(n10869), .QN(g34978) );
  NOR2X0 U10780 ( .IN1(n10870), .IN2(n10871), .QN(n10869) );
  NAND2X0 U10781 ( .IN1(n10872), .IN2(n10873), .QN(n10871) );
  NAND2X0 U10782 ( .IN1(n1030), .IN2(n10874), .QN(n10873) );
  NAND2X0 U10783 ( .IN1(n10875), .IN2(n10876), .QN(n10874) );
  NOR2X0 U10784 ( .IN1(n10877), .IN2(n10878), .QN(n10876) );
  NAND2X0 U10785 ( .IN1(n10879), .IN2(n10880), .QN(n10878) );
  NAND2X0 U10786 ( .IN1(n10830), .IN2(g572), .QN(n10880) );
  NOR2X0 U10787 ( .IN1(n10881), .IN2(n10882), .QN(n10879) );
  NOR2X0 U10788 ( .IN1(n5475), .IN2(n10854), .QN(n10882) );
  NOR2X0 U10789 ( .IN1(n10883), .IN2(g550), .QN(n10881) );
  NAND2X0 U10790 ( .IN1(n10884), .IN2(n10885), .QN(n10877) );
  NAND2X0 U10791 ( .IN1(n10852), .IN2(g790), .QN(n10885) );
  NOR2X0 U10792 ( .IN1(n10886), .IN2(n10887), .QN(n10884) );
  NOR2X0 U10793 ( .IN1(n5488), .IN2(n10888), .QN(n10887) );
  AND2X1 U10794 ( .IN1(g29214), .IN2(n10846), .Q(n10886) );
  NOR2X0 U10795 ( .IN1(n10889), .IN2(n10890), .QN(n10875) );
  NAND2X0 U10796 ( .IN1(n10891), .IN2(n10892), .QN(n10890) );
  OR2X1 U10797 ( .IN1(n10838), .IN2(n9732), .Q(n10892) );
  NAND2X0 U10798 ( .IN1(n10893), .IN2(g4176), .QN(n10891) );
  NAND2X0 U10799 ( .IN1(n10894), .IN2(n10895), .QN(n10889) );
  NAND2X0 U10800 ( .IN1(n10837), .IN2(g2878), .QN(n10895) );
  INVX0 U10801 ( .INP(n10896), .ZN(n10837) );
  NOR2X0 U10802 ( .IN1(n10897), .IN2(n10898), .QN(n10894) );
  AND2X1 U10803 ( .IN1(n10899), .IN2(test_so22), .Q(n10898) );
  AND2X1 U10804 ( .IN1(n10831), .IN2(test_so2), .Q(n10897) );
  NAND2X0 U10805 ( .IN1(n9576), .IN2(n10900), .QN(n10872) );
  NAND2X0 U10806 ( .IN1(n10901), .IN2(n10856), .QN(n10870) );
  NAND2X0 U10807 ( .IN1(n10857), .IN2(g4253), .QN(n10901) );
  NOR2X0 U10808 ( .IN1(n10902), .IN2(n10903), .QN(n10868) );
  NAND2X0 U10809 ( .IN1(n10904), .IN2(n10905), .QN(n10903) );
  NAND2X0 U10810 ( .IN1(n10862), .IN2(g2130), .QN(n10905) );
  NAND2X0 U10811 ( .IN1(n10863), .IN2(g2689), .QN(n10904) );
  NAND2X0 U10812 ( .IN1(n10906), .IN2(n10907), .QN(n10902) );
  NAND2X0 U10813 ( .IN1(n9577), .IN2(n10866), .QN(n10907) );
  NAND2X0 U10814 ( .IN1(n10867), .IN2(n9276), .QN(n10906) );
  OR2X1 U10815 ( .IN1(g34977), .IN2(n9723), .Q(g34923) );
  NAND2X0 U10816 ( .IN1(n10908), .IN2(n10909), .QN(g34977) );
  NOR2X0 U10817 ( .IN1(n10910), .IN2(n10911), .QN(n10909) );
  NAND2X0 U10818 ( .IN1(n10912), .IN2(n10913), .QN(n10911) );
  NAND2X0 U10819 ( .IN1(n1030), .IN2(n10914), .QN(n10913) );
  NAND2X0 U10820 ( .IN1(n10915), .IN2(n10916), .QN(n10914) );
  NOR2X0 U10821 ( .IN1(n10917), .IN2(n10918), .QN(n10916) );
  NAND2X0 U10822 ( .IN1(n10919), .IN2(n10920), .QN(n10918) );
  NAND2X0 U10823 ( .IN1(n10921), .IN2(g613), .QN(n10920) );
  NOR2X0 U10824 ( .IN1(n10922), .IN2(n10923), .QN(n10919) );
  NOR2X0 U10825 ( .IN1(n5490), .IN2(n10883), .QN(n10923) );
  NOR2X0 U10826 ( .IN1(n5291), .IN2(n10924), .QN(n10922) );
  NAND2X0 U10827 ( .IN1(n10925), .IN2(n10926), .QN(n10917) );
  NAND2X0 U10828 ( .IN1(n10847), .IN2(g2868), .QN(n10926) );
  NOR2X0 U10829 ( .IN1(n10927), .IN2(n10928), .QN(n10925) );
  AND2X1 U10830 ( .IN1(g37), .IN2(n10846), .Q(n10928) );
  NOR2X0 U10831 ( .IN1(n10929), .IN2(n10930), .QN(n10915) );
  NAND2X0 U10832 ( .IN1(n10931), .IN2(n10932), .QN(n10930) );
  NAND2X0 U10833 ( .IN1(n10893), .IN2(g4172), .QN(n10932) );
  NOR2X0 U10834 ( .IN1(n10933), .IN2(n10934), .QN(n10931) );
  NOR2X0 U10835 ( .IN1(n9733), .IN2(n10838), .QN(n10934) );
  NOR2X0 U10836 ( .IN1(n9575), .IN2(n10896), .QN(n10933) );
  NAND2X0 U10837 ( .IN1(n10935), .IN2(n10936), .QN(n10929) );
  NAND2X0 U10838 ( .IN1(n10899), .IN2(g2950), .QN(n10936) );
  NOR2X0 U10839 ( .IN1(n10937), .IN2(n10938), .QN(n10935) );
  NOR2X0 U10840 ( .IN1(n5331), .IN2(n10939), .QN(n10938) );
  NOR2X0 U10841 ( .IN1(n5336), .IN2(n10940), .QN(n10937) );
  NAND2X0 U10842 ( .IN1(n10941), .IN2(n5879), .QN(n10912) );
  NAND2X0 U10843 ( .IN1(n10942), .IN2(n10856), .QN(n10910) );
  NAND2X0 U10844 ( .IN1(n10857), .IN2(g4300), .QN(n10942) );
  NOR2X0 U10845 ( .IN1(n10943), .IN2(n10944), .QN(n10908) );
  NAND2X0 U10846 ( .IN1(n10945), .IN2(n10946), .QN(n10944) );
  NAND2X0 U10847 ( .IN1(n10867), .IN2(n9245), .QN(n10946) );
  NAND2X0 U10848 ( .IN1(n10947), .IN2(n5867), .QN(n10945) );
  NAND2X0 U10849 ( .IN1(n10948), .IN2(n10949), .QN(n10943) );
  NAND2X0 U10850 ( .IN1(n10900), .IN2(g1291), .QN(n10949) );
  NAND2X0 U10851 ( .IN1(n10866), .IN2(g947), .QN(n10948) );
  OR2X1 U10852 ( .IN1(g34976), .IN2(n9723), .Q(g34921) );
  NAND2X0 U10853 ( .IN1(n10950), .IN2(n10951), .QN(g34976) );
  NOR2X0 U10854 ( .IN1(n10952), .IN2(n10953), .QN(n10951) );
  NAND2X0 U10855 ( .IN1(n10954), .IN2(n10955), .QN(n10953) );
  NAND2X0 U10856 ( .IN1(n10956), .IN2(n10900), .QN(n10955) );
  NAND2X0 U10857 ( .IN1(n10957), .IN2(n10866), .QN(n10954) );
  NAND2X0 U10858 ( .IN1(n10958), .IN2(n10959), .QN(n10952) );
  NAND2X0 U10859 ( .IN1(n10941), .IN2(g4912), .QN(n10959) );
  NOR2X0 U10860 ( .IN1(n10960), .IN2(n10961), .QN(n10958) );
  NOR2X0 U10861 ( .IN1(n10962), .IN2(n10821), .QN(n10961) );
  NOR2X0 U10862 ( .IN1(n10963), .IN2(n10964), .QN(n10962) );
  NAND2X0 U10863 ( .IN1(n10965), .IN2(n10966), .QN(n10964) );
  NOR2X0 U10864 ( .IN1(n10967), .IN2(n10968), .QN(n10966) );
  NAND2X0 U10865 ( .IN1(n10969), .IN2(n10970), .QN(n10968) );
  NAND2X0 U10866 ( .IN1(n10831), .IN2(g763), .QN(n10970) );
  NAND2X0 U10867 ( .IN1(n10899), .IN2(g2936), .QN(n10969) );
  NOR2X0 U10868 ( .IN1(n10088), .IN2(n10896), .QN(n10967) );
  NOR2X0 U10869 ( .IN1(n10971), .IN2(n10972), .QN(n10965) );
  AND2X1 U10870 ( .IN1(n10893), .IN2(test_so95), .Q(n10972) );
  NOR2X0 U10871 ( .IN1(n10084), .IN2(n10838), .QN(n10971) );
  NAND2X0 U10872 ( .IN1(n10973), .IN2(n10974), .QN(n10963) );
  NOR2X0 U10873 ( .IN1(n10975), .IN2(n10976), .QN(n10974) );
  NAND2X0 U10874 ( .IN1(n10977), .IN2(n10978), .QN(n10976) );
  NAND2X0 U10875 ( .IN1(n10847), .IN2(g2988), .QN(n10977) );
  NOR2X0 U10876 ( .IN1(n5479), .IN2(n10924), .QN(n10975) );
  NOR2X0 U10877 ( .IN1(n10979), .IN2(n10980), .QN(n10973) );
  NAND2X0 U10878 ( .IN1(n10981), .IN2(n10982), .QN(n10980) );
  NAND2X0 U10879 ( .IN1(test_so41), .IN2(n10853), .QN(n10982) );
  INVX0 U10880 ( .INP(n10883), .ZN(n10853) );
  NAND2X0 U10881 ( .IN1(n10921), .IN2(g617), .QN(n10981) );
  INVX0 U10882 ( .INP(n10854), .ZN(n10921) );
  NOR2X0 U10883 ( .IN1(n5294), .IN2(n10940), .QN(n10979) );
  NOR2X0 U10884 ( .IN1(n10983), .IN2(n10984), .QN(n10950) );
  NAND2X0 U10885 ( .IN1(n10985), .IN2(n10986), .QN(n10984) );
  NAND2X0 U10886 ( .IN1(n10947), .IN2(g4722), .QN(n10986) );
  NAND2X0 U10887 ( .IN1(n10863), .IN2(g6545), .QN(n10985) );
  NAND2X0 U10888 ( .IN1(n10987), .IN2(n10988), .QN(n10983) );
  NAND2X0 U10889 ( .IN1(n10867), .IN2(n9357), .QN(n10988) );
  NAND2X0 U10890 ( .IN1(n10862), .IN2(g5160), .QN(n10987) );
  OR2X1 U10891 ( .IN1(g34975), .IN2(n9723), .Q(g34919) );
  NAND2X0 U10892 ( .IN1(n10989), .IN2(n10990), .QN(g34975) );
  NOR2X0 U10893 ( .IN1(n10991), .IN2(n10992), .QN(n10990) );
  NAND2X0 U10894 ( .IN1(n10993), .IN2(n10994), .QN(n10992) );
  NAND2X0 U10895 ( .IN1(n10995), .IN2(n10900), .QN(n10994) );
  NAND2X0 U10896 ( .IN1(n10996), .IN2(n10866), .QN(n10993) );
  NAND2X0 U10897 ( .IN1(n10997), .IN2(n10998), .QN(n10991) );
  NAND2X0 U10898 ( .IN1(n10941), .IN2(g4907), .QN(n10998) );
  NOR2X0 U10899 ( .IN1(n10960), .IN2(n10999), .QN(n10997) );
  NOR2X0 U10900 ( .IN1(n11000), .IN2(n10821), .QN(n10999) );
  NOR2X0 U10901 ( .IN1(n11001), .IN2(n11002), .QN(n11000) );
  NAND2X0 U10902 ( .IN1(n11003), .IN2(n11004), .QN(n11002) );
  NOR2X0 U10903 ( .IN1(n11005), .IN2(n11006), .QN(n11004) );
  NAND2X0 U10904 ( .IN1(n11007), .IN2(n11008), .QN(n11006) );
  NAND2X0 U10905 ( .IN1(n10831), .IN2(g767), .QN(n11008) );
  NAND2X0 U10906 ( .IN1(n10899), .IN2(g2922), .QN(n11007) );
  INVX0 U10907 ( .INP(n10832), .ZN(n10899) );
  NOR2X0 U10908 ( .IN1(n5489), .IN2(n10896), .QN(n11005) );
  NOR2X0 U10909 ( .IN1(n11009), .IN2(n11010), .QN(n11003) );
  NOR2X0 U10910 ( .IN1(n10076), .IN2(n10839), .QN(n11010) );
  NOR2X0 U10911 ( .IN1(n9729), .IN2(n10838), .QN(n11009) );
  NAND2X0 U10912 ( .IN1(n11011), .IN2(n11012), .QN(n11001) );
  NOR2X0 U10913 ( .IN1(n11013), .IN2(n11014), .QN(n11012) );
  NAND2X0 U10914 ( .IN1(n11015), .IN2(n11016), .QN(n11014) );
  NAND2X0 U10915 ( .IN1(n5634), .IN2(n10847), .QN(n11016) );
  NAND2X0 U10916 ( .IN1(n10852), .IN2(g554), .QN(n11015) );
  NOR2X0 U10917 ( .IN1(n5492), .IN2(n10883), .QN(n11013) );
  NOR2X0 U10918 ( .IN1(n11017), .IN2(n11018), .QN(n11011) );
  NOR2X0 U10919 ( .IN1(n5552), .IN2(n10940), .QN(n11018) );
  NOR2X0 U10920 ( .IN1(n5672), .IN2(n10854), .QN(n11017) );
  INVX0 U10921 ( .INP(n10856), .ZN(n10960) );
  NOR2X0 U10922 ( .IN1(n11019), .IN2(n11020), .QN(n10989) );
  NAND2X0 U10923 ( .IN1(n11021), .IN2(n11022), .QN(n11020) );
  NAND2X0 U10924 ( .IN1(n10947), .IN2(g4717), .QN(n11022) );
  NAND2X0 U10925 ( .IN1(n10863), .IN2(g3151), .QN(n11021) );
  NAND2X0 U10926 ( .IN1(n11023), .IN2(n11024), .QN(n11019) );
  NAND2X0 U10927 ( .IN1(n10867), .IN2(n9294), .QN(n11024) );
  NAND2X0 U10928 ( .IN1(n10862), .IN2(g5507), .QN(n11023) );
  OR2X1 U10929 ( .IN1(g34974), .IN2(n9723), .Q(g34917) );
  NAND2X0 U10930 ( .IN1(n11025), .IN2(n11026), .QN(g34974) );
  NOR2X0 U10931 ( .IN1(n11027), .IN2(n11028), .QN(n11026) );
  NAND2X0 U10932 ( .IN1(n11029), .IN2(n11030), .QN(n11028) );
  NAND2X0 U10933 ( .IN1(n11031), .IN2(n10900), .QN(n11030) );
  NAND2X0 U10934 ( .IN1(n11032), .IN2(n10866), .QN(n11029) );
  NAND2X0 U10935 ( .IN1(n11033), .IN2(n11034), .QN(n11027) );
  NAND2X0 U10936 ( .IN1(n10941), .IN2(g4922), .QN(n11034) );
  NOR2X0 U10937 ( .IN1(n11035), .IN2(n11036), .QN(n11033) );
  NOR2X0 U10938 ( .IN1(n11037), .IN2(n10821), .QN(n11036) );
  NOR2X0 U10939 ( .IN1(n11038), .IN2(n11039), .QN(n11037) );
  NAND2X0 U10940 ( .IN1(n11040), .IN2(n11041), .QN(n11039) );
  NOR2X0 U10941 ( .IN1(n11042), .IN2(n11043), .QN(n11041) );
  NOR2X0 U10942 ( .IN1(n9585), .IN2(n10896), .QN(n11043) );
  NOR2X0 U10943 ( .IN1(n10080), .IN2(n10832), .QN(n11042) );
  NOR2X0 U10944 ( .IN1(n11044), .IN2(n11045), .QN(n11040) );
  NOR2X0 U10945 ( .IN1(n10077), .IN2(n10839), .QN(n11045) );
  NOR2X0 U10946 ( .IN1(n9730), .IN2(n10838), .QN(n11044) );
  NAND2X0 U10947 ( .IN1(n11046), .IN2(n11047), .QN(n11038) );
  NOR2X0 U10948 ( .IN1(n11048), .IN2(n11049), .QN(n11047) );
  NOR2X0 U10949 ( .IN1(n5288), .IN2(n10854), .QN(n11049) );
  NOR2X0 U10950 ( .IN1(n10092), .IN2(n10888), .QN(n11048) );
  NOR2X0 U10951 ( .IN1(n11050), .IN2(n11051), .QN(n11046) );
  NOR2X0 U10952 ( .IN1(n5334), .IN2(n10939), .QN(n11051) );
  NOR2X0 U10953 ( .IN1(n5472), .IN2(n10940), .QN(n11050) );
  NOR2X0 U10954 ( .IN1(n11052), .IN2(n11053), .QN(n11025) );
  NAND2X0 U10955 ( .IN1(n11054), .IN2(n11055), .QN(n11053) );
  NAND2X0 U10956 ( .IN1(n10947), .IN2(g4732), .QN(n11055) );
  NAND2X0 U10957 ( .IN1(test_so45), .IN2(n10863), .QN(n11054) );
  NAND2X0 U10958 ( .IN1(n11056), .IN2(n11057), .QN(n11052) );
  NAND2X0 U10959 ( .IN1(n10867), .IN2(n9327), .QN(n11057) );
  NAND2X0 U10960 ( .IN1(n10862), .IN2(g5853), .QN(n11056) );
  NAND2X0 U10961 ( .IN1(n10791), .IN2(g22), .QN(g34915) );
  INVX0 U10962 ( .INP(g34971), .ZN(n10791) );
  NAND2X0 U10963 ( .IN1(n11058), .IN2(n11059), .QN(g34971) );
  NOR2X0 U10964 ( .IN1(n11060), .IN2(n11061), .QN(n11059) );
  NAND2X0 U10965 ( .IN1(n11062), .IN2(n11063), .QN(n11061) );
  NAND2X0 U10966 ( .IN1(n1030), .IN2(n11064), .QN(n11063) );
  NAND2X0 U10967 ( .IN1(n11065), .IN2(n11066), .QN(n11064) );
  NOR2X0 U10968 ( .IN1(n11067), .IN2(n11068), .QN(n11066) );
  NAND2X0 U10969 ( .IN1(n11069), .IN2(n11070), .QN(n11068) );
  NAND2X0 U10970 ( .IN1(n10790), .IN2(g2984), .QN(n11070) );
  INVX0 U10971 ( .INP(n10792), .ZN(n10790) );
  NAND2X0 U10972 ( .IN1(n11071), .IN2(n5324), .QN(n10792) );
  NOR2X0 U10973 ( .IN1(n11072), .IN2(n11073), .QN(n11071) );
  NAND2X0 U10974 ( .IN1(n10852), .IN2(g781), .QN(n11069) );
  NAND2X0 U10975 ( .IN1(n11074), .IN2(n11075), .QN(n11067) );
  NAND2X0 U10976 ( .IN1(n10847), .IN2(g2890), .QN(n11075) );
  INVX0 U10977 ( .INP(n10888), .ZN(n10847) );
  NAND2X0 U10978 ( .IN1(n11076), .IN2(n5468), .QN(n10888) );
  NOR2X0 U10979 ( .IN1(n11072), .IN2(n11077), .QN(n11076) );
  NOR2X0 U10980 ( .IN1(n10927), .IN2(n11078), .QN(n11074) );
  AND2X1 U10981 ( .IN1(g100), .IN2(n10846), .Q(n11078) );
  NOR2X0 U10982 ( .IN1(n11079), .IN2(n11072), .QN(n10846) );
  INVX0 U10983 ( .INP(n10978), .ZN(n10927) );
  NAND2X0 U10984 ( .IN1(n11080), .IN2(n11081), .QN(n10978) );
  NOR2X0 U10985 ( .IN1(n11082), .IN2(n11083), .QN(n11065) );
  NAND2X0 U10986 ( .IN1(n11084), .IN2(n11085), .QN(n11083) );
  NAND2X0 U10987 ( .IN1(n10831), .IN2(test_so60), .QN(n11085) );
  NAND2X0 U10988 ( .IN1(n10893), .IN2(g4157), .QN(n11084) );
  INVX0 U10989 ( .INP(n10839), .ZN(n10893) );
  NAND2X0 U10990 ( .IN1(n11086), .IN2(n11087), .QN(n11082) );
  NAND2X0 U10991 ( .IN1(n10830), .IN2(g562), .QN(n11087) );
  NOR2X0 U10992 ( .IN1(n11088), .IN2(n11089), .QN(n11086) );
  NOR2X0 U10993 ( .IN1(n5550), .IN2(n10854), .QN(n11089) );
  NOR2X0 U10994 ( .IN1(n10098), .IN2(n10883), .QN(n11088) );
  NAND2X0 U10995 ( .IN1(test_so64), .IN2(n10900), .QN(n11062) );
  NAND2X0 U10996 ( .IN1(n11090), .IN2(n10856), .QN(n11060) );
  NAND2X0 U10997 ( .IN1(n11091), .IN2(n1030), .QN(n10856) );
  NOR2X0 U10998 ( .IN1(n10357), .IN2(n11092), .QN(n11091) );
  NOR2X0 U10999 ( .IN1(n10852), .IN2(n11093), .QN(n11092) );
  INVX0 U11000 ( .INP(n10924), .ZN(n10852) );
  NAND2X0 U11001 ( .IN1(n11094), .IN2(n5468), .QN(n10924) );
  NOR2X0 U11002 ( .IN1(n11077), .IN2(n11095), .QN(n11094) );
  NAND2X0 U11003 ( .IN1(n10857), .IN2(g4245), .QN(n11090) );
  AND2X1 U11004 ( .IN1(n11096), .IN2(n11097), .Q(n10857) );
  NOR2X0 U11005 ( .IN1(n11098), .IN2(n11099), .QN(n11058) );
  NAND2X0 U11006 ( .IN1(n11100), .IN2(n11101), .QN(n11099) );
  NAND2X0 U11007 ( .IN1(n10862), .IN2(g2145), .QN(n11101) );
  NAND2X0 U11008 ( .IN1(n10863), .IN2(g2704), .QN(n11100) );
  NAND2X0 U11009 ( .IN1(n11102), .IN2(n11103), .QN(n11098) );
  NAND2X0 U11010 ( .IN1(n10866), .IN2(n9247), .QN(n11103) );
  NAND2X0 U11011 ( .IN1(n10867), .IN2(n9351), .QN(n11102) );
  OR2X1 U11012 ( .IN1(g34970), .IN2(n9723), .Q(g34913) );
  NAND2X0 U11013 ( .IN1(n11104), .IN2(n11105), .QN(g34970) );
  NOR2X0 U11014 ( .IN1(n11106), .IN2(n11107), .QN(n11105) );
  NAND2X0 U11015 ( .IN1(n11108), .IN2(n11109), .QN(n11107) );
  NAND2X0 U11016 ( .IN1(n11110), .IN2(n10900), .QN(n11109) );
  INVX0 U11017 ( .INP(n10819), .ZN(n10900) );
  NAND2X0 U11018 ( .IN1(n11111), .IN2(n11112), .QN(n10819) );
  NOR2X0 U11019 ( .IN1(n11072), .IN2(g9), .QN(n11112) );
  NAND2X0 U11020 ( .IN1(test_so25), .IN2(n9583), .QN(n11072) );
  NAND2X0 U11021 ( .IN1(n11113), .IN2(n10866), .QN(n11108) );
  AND2X1 U11022 ( .IN1(n11114), .IN2(n1030), .Q(n10866) );
  AND2X1 U11023 ( .IN1(n11097), .IN2(n2552), .Q(n11114) );
  INVX0 U11024 ( .INP(n11077), .ZN(n11097) );
  NAND2X0 U11025 ( .IN1(n11115), .IN2(n11116), .QN(n11106) );
  NAND2X0 U11026 ( .IN1(n10941), .IN2(g4917), .QN(n11116) );
  AND2X1 U11027 ( .IN1(n11117), .IN2(n2527), .Q(n10941) );
  NOR2X0 U11028 ( .IN1(n11077), .IN2(n10821), .QN(n11117) );
  NOR2X0 U11029 ( .IN1(n11035), .IN2(n11118), .QN(n11115) );
  NOR2X0 U11030 ( .IN1(n11119), .IN2(n10821), .QN(n11118) );
  NOR2X0 U11031 ( .IN1(n11120), .IN2(n11121), .QN(n11119) );
  NAND2X0 U11032 ( .IN1(n11122), .IN2(n11123), .QN(n11121) );
  NOR2X0 U11033 ( .IN1(n11124), .IN2(n11125), .QN(n11123) );
  NOR2X0 U11034 ( .IN1(n9709), .IN2(n10896), .QN(n11125) );
  NAND2X0 U11035 ( .IN1(n11126), .IN2(n11127), .QN(n10896) );
  NOR2X0 U11036 ( .IN1(n5468), .IN2(n11077), .QN(n11126) );
  NAND2X0 U11037 ( .IN1(n11128), .IN2(g28), .QN(n11077) );
  NOR2X0 U11038 ( .IN1(n10832), .IN2(n10146), .QN(n11124) );
  NAND2X0 U11039 ( .IN1(n11080), .IN2(n11127), .QN(n10832) );
  NOR2X0 U11040 ( .IN1(n5324), .IN2(n11073), .QN(n11080) );
  NOR2X0 U11041 ( .IN1(n11129), .IN2(n11130), .QN(n11122) );
  NOR2X0 U11042 ( .IN1(n10078), .IN2(n10839), .QN(n11130) );
  NAND2X0 U11043 ( .IN1(n11131), .IN2(n11132), .QN(n10839) );
  NOR2X0 U11044 ( .IN1(n5468), .IN2(n11095), .QN(n11131) );
  NOR2X0 U11045 ( .IN1(n9731), .IN2(n10838), .QN(n11129) );
  NAND2X0 U11046 ( .IN1(n11133), .IN2(n11127), .QN(n10838) );
  INVX0 U11047 ( .INP(n11095), .ZN(n11127) );
  NOR2X0 U11048 ( .IN1(n11073), .IN2(g28), .QN(n11133) );
  NAND2X0 U11049 ( .IN1(n11134), .IN2(n11135), .QN(n11073) );
  NOR2X0 U11050 ( .IN1(n9673), .IN2(n5468), .QN(n11135) );
  AND2X1 U11051 ( .IN1(test_so85), .IN2(n3395), .Q(n11134) );
  NAND2X0 U11052 ( .IN1(n11136), .IN2(n11137), .QN(n11120) );
  NOR2X0 U11053 ( .IN1(n11138), .IN2(n11139), .QN(n11137) );
  NOR2X0 U11054 ( .IN1(n18472), .IN2(n10854), .QN(n11139) );
  NOR2X0 U11055 ( .IN1(n5491), .IN2(n10883), .QN(n11138) );
  NAND2X0 U11056 ( .IN1(n11140), .IN2(n11132), .QN(n10883) );
  NOR2X0 U11057 ( .IN1(n11095), .IN2(g9), .QN(n11140) );
  NOR2X0 U11058 ( .IN1(n11141), .IN2(n11142), .QN(n11136) );
  NOR2X0 U11059 ( .IN1(n5330), .IN2(n10939), .QN(n11142) );
  INVX0 U11060 ( .INP(n10831), .ZN(n10939) );
  NOR2X0 U11061 ( .IN1(n5476), .IN2(n10940), .QN(n11141) );
  AND2X1 U11062 ( .IN1(n11143), .IN2(n1030), .Q(n11035) );
  AND2X1 U11063 ( .IN1(n10497), .IN2(n11093), .Q(n11143) );
  NAND2X0 U11064 ( .IN1(n11144), .IN2(n10854), .QN(n11093) );
  NAND2X0 U11065 ( .IN1(n11132), .IN2(n2552), .QN(n10854) );
  NOR2X0 U11066 ( .IN1(n10831), .IN2(n10830), .QN(n11144) );
  INVX0 U11067 ( .INP(n10940), .ZN(n10830) );
  NAND2X0 U11068 ( .IN1(n11145), .IN2(n2552), .QN(n10940) );
  NOR2X0 U11069 ( .IN1(n11079), .IN2(n11095), .QN(n10831) );
  NAND2X0 U11070 ( .IN1(n9583), .IN2(n5477), .QN(n11095) );
  OR2X1 U11071 ( .IN1(n11146), .IN2(n11147), .Q(n11079) );
  NAND2X0 U11072 ( .IN1(g28), .IN2(n5468), .QN(n11146) );
  NOR2X0 U11073 ( .IN1(n11148), .IN2(n11149), .QN(n11104) );
  NAND2X0 U11074 ( .IN1(n11150), .IN2(n11151), .QN(n11149) );
  NAND2X0 U11075 ( .IN1(n10947), .IN2(g4727), .QN(n11151) );
  AND2X1 U11076 ( .IN1(n11111), .IN2(n2527), .Q(n10947) );
  NOR2X0 U11077 ( .IN1(n11152), .IN2(n10821), .QN(n11111) );
  NAND2X0 U11078 ( .IN1(n10863), .IN2(g3853), .QN(n11150) );
  AND2X1 U11079 ( .IN1(n11145), .IN2(n11096), .Q(n10863) );
  NOR2X0 U11080 ( .IN1(g28), .IN2(n11147), .QN(n11145) );
  NAND2X0 U11081 ( .IN1(n11153), .IN2(n11154), .QN(n11147) );
  NOR2X0 U11082 ( .IN1(test_so85), .IN2(n5469), .QN(n11154) );
  NAND2X0 U11083 ( .IN1(n11155), .IN2(n11156), .QN(n11148) );
  NAND2X0 U11084 ( .IN1(n10867), .IN2(n9322), .QN(n11156) );
  NOR2X0 U11085 ( .IN1(n1030), .IN2(g53), .QN(n10867) );
  INVX0 U11086 ( .INP(n10821), .ZN(n1030) );
  NAND2X0 U11087 ( .IN1(n10862), .IN2(g6199), .QN(n11155) );
  AND2X1 U11088 ( .IN1(n11096), .IN2(n11132), .Q(n10862) );
  INVX0 U11089 ( .INP(n11152), .ZN(n11132) );
  NAND2X0 U11090 ( .IN1(n11128), .IN2(n5324), .QN(n11152) );
  AND2X1 U11091 ( .IN1(n11153), .IN2(n11157), .Q(n11128) );
  NOR2X0 U11092 ( .IN1(test_so85), .IN2(g31), .QN(n11157) );
  NOR2X0 U11093 ( .IN1(g6), .IN2(g8), .QN(n11153) );
  AND2X1 U11094 ( .IN1(n11158), .IN2(n11081), .Q(n11096) );
  NOR2X0 U11095 ( .IN1(test_so25), .IN2(n9583), .QN(n11081) );
  NOR2X0 U11096 ( .IN1(n5468), .IN2(n10821), .QN(n11158) );
  NAND2X0 U11097 ( .IN1(n11159), .IN2(n11160), .QN(n10821) );
  NOR2X0 U11098 ( .IN1(test_so74), .IN2(g57), .QN(n11160) );
  NOR2X0 U11099 ( .IN1(g53), .IN2(n10812), .QN(n11159) );
  NAND2X0 U11100 ( .IN1(g54), .IN2(n11161), .QN(n10812) );
  INVX0 U11101 ( .INP(g56), .ZN(n11161) );
  NAND2X0 U11102 ( .IN1(n11162), .IN2(n11163), .QN(g34911) );
  NAND2X0 U11103 ( .IN1(n11164), .IN2(g807), .QN(n11163) );
  NAND2X0 U11104 ( .IN1(n10367), .IN2(n11165), .QN(n11164) );
  NAND2X0 U11105 ( .IN1(n2404), .IN2(g554), .QN(n11162) );
  NAND2X0 U11106 ( .IN1(n11166), .IN2(n11167), .QN(g34882) );
  NAND2X0 U11107 ( .IN1(n10502), .IN2(g4366), .QN(n11167) );
  NAND2X0 U11108 ( .IN1(n11168), .IN2(n10378), .QN(n11166) );
  NAND2X0 U11109 ( .IN1(n11169), .IN2(n11170), .QN(n11168) );
  NAND2X0 U11110 ( .IN1(n11171), .IN2(n11172), .QN(n11170) );
  NOR2X0 U11111 ( .IN1(n11173), .IN2(g4340), .QN(n11171) );
  NOR2X0 U11112 ( .IN1(g4358), .IN2(n11174), .QN(n11173) );
  NOR2X0 U11113 ( .IN1(n11175), .IN2(n11176), .QN(n11169) );
  NOR2X0 U11114 ( .IN1(g4358), .IN2(n11177), .QN(n11176) );
  NAND2X0 U11115 ( .IN1(n11174), .IN2(n10132), .QN(n11177) );
  NAND2X0 U11116 ( .IN1(n11178), .IN2(n11179), .QN(n11174) );
  NOR2X0 U11117 ( .IN1(n11180), .IN2(n11181), .QN(n11179) );
  NOR2X0 U11118 ( .IN1(n5540), .IN2(n11182), .QN(n11181) );
  NAND2X0 U11119 ( .IN1(n5506), .IN2(g4311), .QN(n11182) );
  NOR2X0 U11120 ( .IN1(n11183), .IN2(g4332), .QN(n11180) );
  NOR2X0 U11121 ( .IN1(n11184), .IN2(n11185), .QN(n11183) );
  NAND2X0 U11122 ( .IN1(n11186), .IN2(n11187), .QN(n11185) );
  NAND2X0 U11123 ( .IN1(n10046), .IN2(g4322), .QN(n11187) );
  NAND2X0 U11124 ( .IN1(n11188), .IN2(n5506), .QN(n11186) );
  AND2X1 U11125 ( .IN1(g90), .IN2(n5634), .Q(n11188) );
  NOR2X0 U11126 ( .IN1(test_so81), .IN2(g4340), .QN(n11178) );
  NOR2X0 U11127 ( .IN1(n5348), .IN2(n11189), .QN(n11175) );
  NAND2X0 U11128 ( .IN1(test_so81), .IN2(g4340), .QN(n11189) );
  NAND2X0 U11129 ( .IN1(n11190), .IN2(n11191), .QN(g34881) );
  NAND2X0 U11130 ( .IN1(n10499), .IN2(g794), .QN(n11191) );
  NOR2X0 U11131 ( .IN1(n11192), .IN2(n11193), .QN(n11190) );
  NOR2X0 U11132 ( .IN1(g807), .IN2(n11165), .QN(n11193) );
  NOR2X0 U11133 ( .IN1(n5479), .IN2(n11194), .QN(n11192) );
  NAND2X0 U11134 ( .IN1(n2404), .IN2(n11165), .QN(n11194) );
  INVX0 U11135 ( .INP(n2405), .ZN(n11165) );
  NAND2X0 U11136 ( .IN1(n11195), .IN2(n11196), .QN(g34880) );
  NAND2X0 U11137 ( .IN1(n10499), .IN2(g626), .QN(n11196) );
  NOR2X0 U11138 ( .IN1(n11197), .IN2(n11198), .QN(n11195) );
  AND2X1 U11139 ( .IN1(n18472), .IN2(n2422), .Q(n11198) );
  NOR2X0 U11140 ( .IN1(n18472), .IN2(n11199), .QN(n11197) );
  OR2X1 U11141 ( .IN1(n11200), .IN2(n2422), .Q(n11199) );
  NAND2X0 U11142 ( .IN1(n11201), .IN2(n11202), .QN(g34850) );
  NAND2X0 U11143 ( .IN1(n10499), .IN2(g790), .QN(n11202) );
  NOR2X0 U11144 ( .IN1(n11203), .IN2(n11204), .QN(n11201) );
  NOR2X0 U11145 ( .IN1(g794), .IN2(n11205), .QN(n11204) );
  NOR2X0 U11146 ( .IN1(n5291), .IN2(n11206), .QN(n11203) );
  NAND2X0 U11147 ( .IN1(n2404), .IN2(n11205), .QN(n11206) );
  INVX0 U11148 ( .INP(n2419), .ZN(n11205) );
  NAND2X0 U11149 ( .IN1(n11207), .IN2(n11208), .QN(g34849) );
  NAND2X0 U11150 ( .IN1(n10500), .IN2(g622), .QN(n11208) );
  NOR2X0 U11151 ( .IN1(n11209), .IN2(n11210), .QN(n11207) );
  NOR2X0 U11152 ( .IN1(g626), .IN2(n11211), .QN(n11210) );
  NOR2X0 U11153 ( .IN1(n5288), .IN2(n11212), .QN(n11209) );
  NAND2X0 U11154 ( .IN1(n2421), .IN2(n11211), .QN(n11212) );
  INVX0 U11155 ( .INP(n2423), .ZN(n11211) );
  NOR2X0 U11156 ( .IN1(n9911), .IN2(n11213), .QN(g34839) );
  NOR2X0 U11157 ( .IN1(g4366), .IN2(n11214), .QN(n11213) );
  NAND2X0 U11158 ( .IN1(n11215), .IN2(n11216), .QN(n11214) );
  NAND2X0 U11159 ( .IN1(n11217), .IN2(g4332), .QN(n11216) );
  NAND2X0 U11160 ( .IN1(n11218), .IN2(g73), .QN(n11217) );
  NOR2X0 U11161 ( .IN1(n11219), .IN2(g4311), .QN(n11218) );
  NAND2X0 U11162 ( .IN1(n5540), .IN2(n11220), .QN(n11215) );
  NAND2X0 U11163 ( .IN1(n11221), .IN2(n5323), .QN(n11220) );
  NOR2X0 U11164 ( .IN1(g73), .IN2(n11219), .QN(n11221) );
  INVX0 U11165 ( .INP(n11222), .ZN(n11219) );
  NAND2X0 U11166 ( .IN1(n11223), .IN2(n11224), .QN(g34808) );
  OR2X1 U11167 ( .IN1(n10305), .IN2(n9733), .Q(n11224) );
  NAND2X0 U11168 ( .IN1(n11225), .IN2(n10378), .QN(n11223) );
  NAND2X0 U11169 ( .IN1(n11226), .IN2(n9732), .QN(n11225) );
  AND2X1 U11170 ( .IN1(n11227), .IN2(g91), .Q(n11226) );
  NAND2X0 U11171 ( .IN1(n11228), .IN2(n11229), .QN(g34807) );
  OR2X1 U11172 ( .IN1(n10305), .IN2(n10084), .Q(n11229) );
  NAND2X0 U11173 ( .IN1(n11230), .IN2(n10378), .QN(n11228) );
  NAND2X0 U11174 ( .IN1(n11231), .IN2(n11232), .QN(n11230) );
  NOR2X0 U11175 ( .IN1(n11233), .IN2(n11234), .QN(n11232) );
  OR2X1 U11176 ( .IN1(n11235), .IN2(n11236), .Q(n11234) );
  NAND2X0 U11177 ( .IN1(n11237), .IN2(n11238), .QN(n11233) );
  NOR2X0 U11178 ( .IN1(n11239), .IN2(n11240), .QN(n11231) );
  NAND2X0 U11179 ( .IN1(n9733), .IN2(n9665), .QN(n11240) );
  NAND2X0 U11180 ( .IN1(n10087), .IN2(n11241), .QN(n11239) );
  NAND2X0 U11181 ( .IN1(n11242), .IN2(n11243), .QN(g34806) );
  OR2X1 U11182 ( .IN1(n10305), .IN2(n9729), .Q(n11243) );
  NAND2X0 U11183 ( .IN1(n11244), .IN2(n10379), .QN(n11242) );
  NAND2X0 U11184 ( .IN1(n11245), .IN2(n10094), .QN(n11244) );
  AND2X1 U11185 ( .IN1(n10084), .IN2(n10093), .Q(n11245) );
  NOR2X0 U11186 ( .IN1(n10492), .IN2(n11246), .QN(g34805) );
  AND2X1 U11187 ( .IN1(n10091), .IN2(n10092), .Q(n11246) );
  NAND2X0 U11188 ( .IN1(n11247), .IN2(n11248), .QN(g34804) );
  NAND2X0 U11189 ( .IN1(n10500), .IN2(g2965), .QN(n11248) );
  NAND2X0 U11190 ( .IN1(n11249), .IN2(n10379), .QN(n11247) );
  NAND2X0 U11191 ( .IN1(n11250), .IN2(n5750), .QN(n11249) );
  NOR2X0 U11192 ( .IN1(n5796), .IN2(n5630), .QN(n11250) );
  NAND2X0 U11193 ( .IN1(n11251), .IN2(n11252), .QN(g34803) );
  OR2X1 U11194 ( .IN1(n10305), .IN2(n9730), .Q(n11252) );
  NAND2X0 U11195 ( .IN1(n11253), .IN2(n10381), .QN(n11251) );
  NAND2X0 U11196 ( .IN1(n11254), .IN2(n9729), .QN(n11253) );
  AND2X1 U11197 ( .IN1(n10091), .IN2(g44), .Q(n11254) );
  NAND2X0 U11198 ( .IN1(n11255), .IN2(n11256), .QN(g34802) );
  OR2X1 U11199 ( .IN1(n10305), .IN2(n9731), .Q(n11256) );
  NAND2X0 U11200 ( .IN1(n11257), .IN2(n10381), .QN(n11255) );
  NAND2X0 U11201 ( .IN1(n11258), .IN2(n9730), .QN(n11257) );
  NOR2X0 U11202 ( .IN1(n11259), .IN2(n11260), .QN(n11258) );
  NAND2X0 U11203 ( .IN1(n11261), .IN2(n11262), .QN(g34801) );
  NAND2X0 U11204 ( .IN1(n10500), .IN2(g2970), .QN(n11262) );
  NAND2X0 U11205 ( .IN1(n11263), .IN2(n10383), .QN(n11261) );
  NAND2X0 U11206 ( .IN1(n11264), .IN2(n9731), .QN(n11263) );
  AND2X1 U11207 ( .IN1(n11265), .IN2(n10096), .Q(n11264) );
  NAND2X0 U11208 ( .IN1(n11266), .IN2(n11267), .QN(g34800) );
  NAND2X0 U11209 ( .IN1(n10500), .IN2(g2886), .QN(n11267) );
  NAND2X0 U11210 ( .IN1(n11268), .IN2(n10385), .QN(n11266) );
  OR2X1 U11211 ( .IN1(test_so74), .IN2(test_so14), .Q(n11268) );
  NAND2X0 U11212 ( .IN1(n11269), .IN2(n11270), .QN(g34799) );
  NAND2X0 U11213 ( .IN1(n10500), .IN2(g2873), .QN(n11270) );
  NAND2X0 U11214 ( .IN1(n11271), .IN2(n10385), .QN(n11269) );
  NAND2X0 U11215 ( .IN1(n10090), .IN2(g44), .QN(n11271) );
  NAND2X0 U11216 ( .IN1(n11272), .IN2(n11273), .QN(g34798) );
  NAND2X0 U11217 ( .IN1(n10500), .IN2(g2878), .QN(n11273) );
  NAND2X0 U11218 ( .IN1(n11274), .IN2(n10385), .QN(n11272) );
  NAND2X0 U11219 ( .IN1(n10086), .IN2(n10087), .QN(n11274) );
  NAND2X0 U11220 ( .IN1(n11275), .IN2(n11276), .QN(g34797) );
  OR2X1 U11221 ( .IN1(n10305), .IN2(n9575), .Q(n11276) );
  NAND2X0 U11222 ( .IN1(n11277), .IN2(n10386), .QN(n11275) );
  NAND2X0 U11223 ( .IN1(n10085), .IN2(g91), .QN(n11277) );
  NAND2X0 U11224 ( .IN1(n11278), .IN2(n11279), .QN(g34796) );
  OR2X1 U11225 ( .IN1(n10306), .IN2(n10088), .Q(n11279) );
  NAND2X0 U11226 ( .IN1(n11280), .IN2(n10386), .QN(n11278) );
  NAND2X0 U11227 ( .IN1(n9575), .IN2(n11227), .QN(n11280) );
  NOR2X0 U11228 ( .IN1(n11281), .IN2(n11282), .QN(n11227) );
  NAND2X0 U11229 ( .IN1(n11283), .IN2(n11284), .QN(g34795) );
  NAND2X0 U11230 ( .IN1(n10500), .IN2(g2864), .QN(n11284) );
  NAND2X0 U11231 ( .IN1(n11285), .IN2(n10378), .QN(n11283) );
  NAND2X0 U11232 ( .IN1(n10088), .IN2(n11237), .QN(n11285) );
  AND2X1 U11233 ( .IN1(n11286), .IN2(n11287), .Q(n11237) );
  NOR2X0 U11234 ( .IN1(n11288), .IN2(n11289), .QN(n11287) );
  NOR2X0 U11235 ( .IN1(g3129), .IN2(g3143), .QN(n11286) );
  NAND2X0 U11236 ( .IN1(n11290), .IN2(n11291), .QN(g34794) );
  NOR2X0 U11237 ( .IN1(n11292), .IN2(n11293), .QN(n11290) );
  NOR2X0 U11238 ( .IN1(n10494), .IN2(n11294), .QN(n11293) );
  NOR2X0 U11239 ( .IN1(n11236), .IN2(g2864), .QN(n11294) );
  NAND2X0 U11240 ( .IN1(n11295), .IN2(n11296), .QN(n11236) );
  NOR2X0 U11241 ( .IN1(n11297), .IN2(n11298), .QN(n11296) );
  OR2X1 U11242 ( .IN1(n11299), .IN2(n11300), .Q(n11298) );
  NOR2X0 U11243 ( .IN1(n9585), .IN2(n10313), .QN(n11292) );
  NAND2X0 U11244 ( .IN1(n11301), .IN2(n11302), .QN(g34793) );
  OR2X1 U11245 ( .IN1(n10306), .IN2(n9709), .Q(n11302) );
  NAND2X0 U11246 ( .IN1(n11303), .IN2(n10386), .QN(n11301) );
  NAND2X0 U11247 ( .IN1(n11304), .IN2(n9585), .QN(n11303) );
  NOR2X0 U11248 ( .IN1(n11235), .IN2(n11305), .QN(n11304) );
  NAND2X0 U11249 ( .IN1(n11306), .IN2(n11307), .QN(g34792) );
  NAND2X0 U11250 ( .IN1(n10500), .IN2(g29214), .QN(n11307) );
  NAND2X0 U11251 ( .IN1(n11308), .IN2(n10386), .QN(n11306) );
  NAND2X0 U11252 ( .IN1(n9709), .IN2(n11238), .QN(n11308) );
  NOR2X0 U11253 ( .IN1(n11309), .IN2(n11310), .QN(n11238) );
  NAND2X0 U11254 ( .IN1(n11311), .IN2(n11312), .QN(g34791) );
  NAND2X0 U11255 ( .IN1(n10500), .IN2(g785), .QN(n11312) );
  NOR2X0 U11256 ( .IN1(n11313), .IN2(n11314), .QN(n11311) );
  NOR2X0 U11257 ( .IN1(g790), .IN2(n11315), .QN(n11314) );
  NOR2X0 U11258 ( .IN1(n5292), .IN2(n11316), .QN(n11313) );
  NAND2X0 U11259 ( .IN1(n2404), .IN2(n11315), .QN(n11316) );
  INVX0 U11260 ( .INP(n2425), .ZN(n11315) );
  NAND2X0 U11261 ( .IN1(n11317), .IN2(n11318), .QN(g34790) );
  NAND2X0 U11262 ( .IN1(n10500), .IN2(g617), .QN(n11318) );
  NOR2X0 U11263 ( .IN1(n11319), .IN2(n11320), .QN(n11317) );
  NOR2X0 U11264 ( .IN1(g622), .IN2(n11321), .QN(n11320) );
  NOR2X0 U11265 ( .IN1(n5672), .IN2(n11322), .QN(n11319) );
  NAND2X0 U11266 ( .IN1(n2421), .IN2(n11321), .QN(n11322) );
  INVX0 U11267 ( .INP(n2427), .ZN(n11321) );
  NOR2X0 U11268 ( .IN1(n5305), .IN2(n11323), .QN(g34788) );
  AND2X1 U11269 ( .IN1(g479), .IN2(n3195), .Q(n11323) );
  NAND2X0 U11270 ( .IN1(n11324), .IN2(n11325), .QN(g34783) );
  NAND2X0 U11271 ( .IN1(n11326), .IN2(n11327), .QN(n11325) );
  NOR2X0 U11272 ( .IN1(n11328), .IN2(n11329), .QN(n11326) );
  NAND2X0 U11273 ( .IN1(n11330), .IN2(n11331), .QN(n11324) );
  NOR2X0 U11274 ( .IN1(n11332), .IN2(n11333), .QN(n11330) );
  NAND2X0 U11275 ( .IN1(n11334), .IN2(n11335), .QN(g34735) );
  NAND2X0 U11276 ( .IN1(n10501), .IN2(g4297), .QN(n11335) );
  NAND2X0 U11277 ( .IN1(n11336), .IN2(n10384), .QN(n11334) );
  NAND2X0 U11278 ( .IN1(n5639), .IN2(n10089), .QN(n11336) );
  NAND2X0 U11279 ( .IN1(n11337), .IN2(n11338), .QN(g34734) );
  NAND2X0 U11280 ( .IN1(n10501), .IN2(g4172), .QN(n11338) );
  NAND2X0 U11281 ( .IN1(n11339), .IN2(n10384), .QN(n11337) );
  NAND2X0 U11282 ( .IN1(n5494), .IN2(n10093), .QN(n11339) );
  NOR2X0 U11283 ( .IN1(n10495), .IN2(n11340), .QN(g34733) );
  NOR2X0 U11284 ( .IN1(g4153), .IN2(g4172), .QN(n11340) );
  NAND2X0 U11285 ( .IN1(n11341), .IN2(n11342), .QN(g34732) );
  NAND2X0 U11286 ( .IN1(n10377), .IN2(g2994), .QN(n11342) );
  OR2X1 U11287 ( .IN1(n10306), .IN2(n10092), .Q(n11341) );
  NAND2X0 U11288 ( .IN1(n11343), .IN2(n11344), .QN(g34731) );
  OR2X1 U11289 ( .IN1(n10306), .IN2(n5635), .Q(n11344) );
  NAND2X0 U11290 ( .IN1(n11345), .IN2(n10384), .QN(n11343) );
  OR2X1 U11291 ( .IN1(n11259), .IN2(test_so64), .Q(n11345) );
  NAND2X0 U11292 ( .IN1(n11346), .IN2(n11347), .QN(g34730) );
  OR2X1 U11293 ( .IN1(n10306), .IN2(n9576), .Q(n11347) );
  NAND2X0 U11294 ( .IN1(n11348), .IN2(n10383), .QN(n11346) );
  NAND2X0 U11295 ( .IN1(n5635), .IN2(n10095), .QN(n11348) );
  OR2X1 U11296 ( .IN1(n2499), .IN2(n11349), .Q(g34729) );
  NAND2X0 U11297 ( .IN1(n11350), .IN2(n11351), .QN(n11349) );
  NAND2X0 U11298 ( .IN1(n5796), .IN2(n10381), .QN(n11351) );
  NAND2X0 U11299 ( .IN1(n10501), .IN2(g1291), .QN(n11350) );
  NAND2X0 U11300 ( .IN1(n11352), .IN2(n11353), .QN(g34728) );
  NAND2X0 U11301 ( .IN1(n10501), .IN2(g939), .QN(n11353) );
  NAND2X0 U11302 ( .IN1(n11354), .IN2(n10380), .QN(n11352) );
  NAND2X0 U11303 ( .IN1(n18478), .IN2(n11355), .QN(n11354) );
  NAND2X0 U11304 ( .IN1(n11356), .IN2(n11357), .QN(g34727) );
  OR2X1 U11305 ( .IN1(n10307), .IN2(n9577), .Q(n11357) );
  NAND2X0 U11306 ( .IN1(n11358), .IN2(n10379), .QN(n11356) );
  NAND2X0 U11307 ( .IN1(n5415), .IN2(n10100), .QN(n11358) );
  OR2X1 U11308 ( .IN1(n2505), .IN2(n11359), .Q(g34726) );
  NAND2X0 U11309 ( .IN1(n11360), .IN2(n11361), .QN(n11359) );
  NAND2X0 U11310 ( .IN1(n5630), .IN2(n10382), .QN(n11361) );
  NAND2X0 U11311 ( .IN1(n10501), .IN2(g947), .QN(n11360) );
  NAND2X0 U11312 ( .IN1(n11362), .IN2(n11363), .QN(g34725) );
  NAND2X0 U11313 ( .IN1(n10501), .IN2(g781), .QN(n11363) );
  NOR2X0 U11314 ( .IN1(n11364), .IN2(n11365), .QN(n11362) );
  NOR2X0 U11315 ( .IN1(g785), .IN2(n11366), .QN(n11365) );
  NOR2X0 U11316 ( .IN1(n5293), .IN2(n11367), .QN(n11364) );
  NAND2X0 U11317 ( .IN1(n2404), .IN2(n11366), .QN(n11367) );
  INVX0 U11318 ( .INP(n2485), .ZN(n11366) );
  NAND2X0 U11319 ( .IN1(n11368), .IN2(n11369), .QN(g34724) );
  NAND2X0 U11320 ( .IN1(n10501), .IN2(g613), .QN(n11369) );
  NOR2X0 U11321 ( .IN1(n11370), .IN2(n11371), .QN(n11368) );
  NOR2X0 U11322 ( .IN1(g617), .IN2(n11372), .QN(n11371) );
  NOR2X0 U11323 ( .IN1(n5339), .IN2(n11373), .QN(n11370) );
  NAND2X0 U11324 ( .IN1(n2421), .IN2(n11372), .QN(n11373) );
  INVX0 U11325 ( .INP(n2487), .ZN(n11372) );
  NAND2X0 U11326 ( .IN1(n11374), .IN2(n11375), .QN(g34723) );
  NAND2X0 U11327 ( .IN1(test_so41), .IN2(n10515), .QN(n11375) );
  NAND2X0 U11328 ( .IN1(n11376), .IN2(n10380), .QN(n11374) );
  NAND2X0 U11329 ( .IN1(n5490), .IN2(n10096), .QN(n11376) );
  NAND2X0 U11330 ( .IN1(n11377), .IN2(n11378), .QN(g34722) );
  NAND2X0 U11331 ( .IN1(n10502), .IN2(g538), .QN(n11378) );
  NAND2X0 U11332 ( .IN1(n11379), .IN2(n10381), .QN(n11377) );
  NAND2X0 U11333 ( .IN1(n5492), .IN2(g691), .QN(n11379) );
  NAND2X0 U11334 ( .IN1(n11380), .IN2(n11381), .QN(g34721) );
  NAND2X0 U11335 ( .IN1(g29221), .IN2(n10514), .QN(n11381) );
  NAND2X0 U11336 ( .IN1(n11382), .IN2(n10381), .QN(n11380) );
  NAND2X0 U11337 ( .IN1(n10099), .IN2(n10098), .QN(n11382) );
  NAND2X0 U11338 ( .IN1(n11383), .IN2(n11384), .QN(g34720) );
  OR2X1 U11339 ( .IN1(n10307), .IN2(n5490), .Q(n11384) );
  NAND2X0 U11340 ( .IN1(n11385), .IN2(n10383), .QN(n11383) );
  NAND2X0 U11341 ( .IN1(n10097), .IN2(g29212), .QN(n11385) );
  NOR2X0 U11342 ( .IN1(n10496), .IN2(n11386), .QN(g34719) );
  NOR2X0 U11343 ( .IN1(g209), .IN2(g538), .QN(n11386) );
  NOR2X0 U11344 ( .IN1(n5497), .IN2(n10463), .QN(g34647) );
  NOR2X0 U11345 ( .IN1(n5644), .IN2(n10463), .QN(g34646) );
  NOR2X0 U11346 ( .IN1(n5499), .IN2(n10462), .QN(g34645) );
  NOR2X0 U11347 ( .IN1(n5643), .IN2(n10462), .QN(g34644) );
  NOR2X0 U11348 ( .IN1(n5498), .IN2(n10462), .QN(g34643) );
  NAND2X0 U11349 ( .IN1(n11387), .IN2(n11388), .QN(g34642) );
  NAND2X0 U11350 ( .IN1(n10377), .IN2(g4927), .QN(n11388) );
  NAND2X0 U11351 ( .IN1(n10502), .IN2(g4912), .QN(n11387) );
  NAND2X0 U11352 ( .IN1(n11389), .IN2(n11390), .QN(g34641) );
  NAND2X0 U11353 ( .IN1(n10375), .IN2(g4912), .QN(n11390) );
  NAND2X0 U11354 ( .IN1(n10502), .IN2(g4907), .QN(n11389) );
  NAND2X0 U11355 ( .IN1(n11391), .IN2(n11392), .QN(g34640) );
  NAND2X0 U11356 ( .IN1(n10377), .IN2(g4907), .QN(n11392) );
  NAND2X0 U11357 ( .IN1(n10502), .IN2(g4922), .QN(n11391) );
  NAND2X0 U11358 ( .IN1(n11393), .IN2(n11394), .QN(g34639) );
  NAND2X0 U11359 ( .IN1(n10376), .IN2(g4922), .QN(n11394) );
  NAND2X0 U11360 ( .IN1(n10502), .IN2(g4917), .QN(n11393) );
  NOR2X0 U11361 ( .IN1(n5408), .IN2(n10461), .QN(g34638) );
  NAND2X0 U11362 ( .IN1(n11395), .IN2(n11396), .QN(g34637) );
  OR2X1 U11363 ( .IN1(n10457), .IN2(n5867), .Q(n11396) );
  NAND2X0 U11364 ( .IN1(n10502), .IN2(g4722), .QN(n11395) );
  NAND2X0 U11365 ( .IN1(n11397), .IN2(n11398), .QN(g34636) );
  NAND2X0 U11366 ( .IN1(n10376), .IN2(g4722), .QN(n11398) );
  NAND2X0 U11367 ( .IN1(n10502), .IN2(g4717), .QN(n11397) );
  NAND2X0 U11368 ( .IN1(n11399), .IN2(n11400), .QN(g34635) );
  NAND2X0 U11369 ( .IN1(n10375), .IN2(g4717), .QN(n11400) );
  NAND2X0 U11370 ( .IN1(n10502), .IN2(g4732), .QN(n11399) );
  NAND2X0 U11371 ( .IN1(n11401), .IN2(n11402), .QN(g34634) );
  NAND2X0 U11372 ( .IN1(n10375), .IN2(g4732), .QN(n11402) );
  NAND2X0 U11373 ( .IN1(n10503), .IN2(g4727), .QN(n11401) );
  NOR2X0 U11374 ( .IN1(n5312), .IN2(n10462), .QN(g34633) );
  NAND2X0 U11375 ( .IN1(n11403), .IN2(n11404), .QN(g34632) );
  NAND2X0 U11376 ( .IN1(n10376), .IN2(g4245), .QN(n11404) );
  NAND2X0 U11377 ( .IN1(test_so67), .IN2(n10515), .QN(n11403) );
  NAND2X0 U11378 ( .IN1(n11405), .IN2(n11406), .QN(g34631) );
  NAND2X0 U11379 ( .IN1(test_so67), .IN2(n10385), .QN(n11406) );
  NAND2X0 U11380 ( .IN1(n10503), .IN2(g4253), .QN(n11405) );
  NAND2X0 U11381 ( .IN1(n11407), .IN2(n11408), .QN(g34630) );
  NAND2X0 U11382 ( .IN1(n10376), .IN2(g4253), .QN(n11408) );
  NAND2X0 U11383 ( .IN1(n10503), .IN2(g4300), .QN(n11407) );
  NAND2X0 U11384 ( .IN1(n11409), .IN2(n11410), .QN(g34629) );
  NAND2X0 U11385 ( .IN1(n10375), .IN2(g4157), .QN(n11410) );
  NAND2X0 U11386 ( .IN1(n10503), .IN2(g4146), .QN(n11409) );
  NAND2X0 U11387 ( .IN1(n11411), .IN2(n11412), .QN(g34628) );
  NAND2X0 U11388 ( .IN1(n10375), .IN2(g4146), .QN(n11412) );
  NAND2X0 U11389 ( .IN1(n10503), .IN2(g4176), .QN(n11411) );
  NOR2X0 U11390 ( .IN1(n5641), .IN2(n10461), .QN(g34627) );
  AND2X1 U11391 ( .IN1(n10366), .IN2(test_so45), .Q(g34626) );
  NOR2X0 U11392 ( .IN1(n5495), .IN2(n10461), .QN(g34625) );
  NAND2X0 U11393 ( .IN1(n11413), .IN2(n11414), .QN(g34624) );
  NAND2X0 U11394 ( .IN1(n10374), .IN2(g2988), .QN(n11414) );
  NAND2X0 U11395 ( .IN1(n10503), .IN2(g2994), .QN(n11413) );
  NAND2X0 U11396 ( .IN1(n11415), .IN2(n11416), .QN(g34623) );
  NAND2X0 U11397 ( .IN1(n10374), .IN2(g2970), .QN(n11416) );
  NAND2X0 U11398 ( .IN1(test_so22), .IN2(n10515), .QN(n11415) );
  NAND2X0 U11399 ( .IN1(n11417), .IN2(n11418), .QN(g34622) );
  NAND2X0 U11400 ( .IN1(test_so22), .IN2(n10386), .QN(n11418) );
  NAND2X0 U11401 ( .IN1(n10503), .IN2(g2950), .QN(n11417) );
  NAND2X0 U11402 ( .IN1(n11419), .IN2(n11420), .QN(g34621) );
  NAND2X0 U11403 ( .IN1(n10374), .IN2(g2950), .QN(n11420) );
  NAND2X0 U11404 ( .IN1(n10503), .IN2(g2936), .QN(n11419) );
  NAND2X0 U11405 ( .IN1(n11421), .IN2(n11422), .QN(g34620) );
  NAND2X0 U11406 ( .IN1(n10373), .IN2(g2936), .QN(n11422) );
  NAND2X0 U11407 ( .IN1(n10503), .IN2(g2922), .QN(n11421) );
  NAND2X0 U11408 ( .IN1(n11423), .IN2(n11424), .QN(g34619) );
  NAND2X0 U11409 ( .IN1(n10373), .IN2(g2922), .QN(n11424) );
  NAND2X0 U11410 ( .IN1(n10503), .IN2(g2912), .QN(n11423) );
  NAND2X0 U11411 ( .IN1(n11425), .IN2(n11426), .QN(g34618) );
  NAND2X0 U11412 ( .IN1(n10373), .IN2(g2912), .QN(n11426) );
  NAND2X0 U11413 ( .IN1(test_so1), .IN2(n10516), .QN(n11425) );
  NAND2X0 U11414 ( .IN1(n11427), .IN2(n11428), .QN(g34617) );
  NAND2X0 U11415 ( .IN1(test_so1), .IN2(n10386), .QN(n11428) );
  NAND2X0 U11416 ( .IN1(n10504), .IN2(g2984), .QN(n11427) );
  NAND2X0 U11417 ( .IN1(n11429), .IN2(n11430), .QN(g34616) );
  NAND2X0 U11418 ( .IN1(n10373), .IN2(g2868), .QN(n11430) );
  NAND2X0 U11419 ( .IN1(n10504), .IN2(g2988), .QN(n11429) );
  NAND2X0 U11420 ( .IN1(n11431), .IN2(n11432), .QN(g34615) );
  NAND2X0 U11421 ( .IN1(n10373), .IN2(g2873), .QN(n11432) );
  NAND2X0 U11422 ( .IN1(n10504), .IN2(g2868), .QN(n11431) );
  NAND2X0 U11423 ( .IN1(n11433), .IN2(n11434), .QN(g34614) );
  NAND2X0 U11424 ( .IN1(n10372), .IN2(g29214), .QN(n11434) );
  NAND2X0 U11425 ( .IN1(g37), .IN2(n10516), .QN(n11433) );
  NAND2X0 U11426 ( .IN1(n11435), .IN2(n11436), .QN(g34613) );
  NAND2X0 U11427 ( .IN1(test_so95), .IN2(n10516), .QN(n11436) );
  NAND2X0 U11428 ( .IN1(g37), .IN2(n10386), .QN(n11435) );
  NAND2X0 U11429 ( .IN1(n11437), .IN2(n11438), .QN(g34612) );
  NAND2X0 U11430 ( .IN1(test_so95), .IN2(n10386), .QN(n11438) );
  NAND2X0 U11431 ( .IN1(n10504), .IN2(g2860), .QN(n11437) );
  NAND2X0 U11432 ( .IN1(n11439), .IN2(n11440), .QN(g34611) );
  NAND2X0 U11433 ( .IN1(n10372), .IN2(g2860), .QN(n11440) );
  NAND2X0 U11434 ( .IN1(n10504), .IN2(g2852), .QN(n11439) );
  NAND2X0 U11435 ( .IN1(n11441), .IN2(n11442), .QN(g34610) );
  NAND2X0 U11436 ( .IN1(n10372), .IN2(g2852), .QN(n11442) );
  NAND2X0 U11437 ( .IN1(n10504), .IN2(g2844), .QN(n11441) );
  NAND2X0 U11438 ( .IN1(n11443), .IN2(n11444), .QN(g34609) );
  NAND2X0 U11439 ( .IN1(n10372), .IN2(g2844), .QN(n11444) );
  NAND2X0 U11440 ( .IN1(n10504), .IN2(g2890), .QN(n11443) );
  NAND2X0 U11441 ( .IN1(n11445), .IN2(n11446), .QN(g34608) );
  NAND2X0 U11442 ( .IN1(n10372), .IN2(g2704), .QN(n11446) );
  NAND2X0 U11443 ( .IN1(n10504), .IN2(g2697), .QN(n11445) );
  NAND2X0 U11444 ( .IN1(n11447), .IN2(n11448), .QN(g34607) );
  NAND2X0 U11445 ( .IN1(n10372), .IN2(g2697), .QN(n11448) );
  NAND2X0 U11446 ( .IN1(n10504), .IN2(g2689), .QN(n11447) );
  NOR2X0 U11447 ( .IN1(n5347), .IN2(n10460), .QN(g34606) );
  NAND2X0 U11448 ( .IN1(n11449), .IN2(n11450), .QN(g34605) );
  NAND2X0 U11449 ( .IN1(n10371), .IN2(g2145), .QN(n11450) );
  NAND2X0 U11450 ( .IN1(n10504), .IN2(g2138), .QN(n11449) );
  NAND2X0 U11451 ( .IN1(n11451), .IN2(n11452), .QN(g34604) );
  NAND2X0 U11452 ( .IN1(n10371), .IN2(g2138), .QN(n11452) );
  NAND2X0 U11453 ( .IN1(n10505), .IN2(g2130), .QN(n11451) );
  NOR2X0 U11454 ( .IN1(n5487), .IN2(n10460), .QN(g34603) );
  NOR2X0 U11455 ( .IN1(n2549), .IN2(n10460), .QN(g34602) );
  NOR2X0 U11456 ( .IN1(n5286), .IN2(n10460), .QN(g34601) );
  NAND2X0 U11457 ( .IN1(n11453), .IN2(n11454), .QN(g34600) );
  NAND2X0 U11458 ( .IN1(n10505), .IN2(g776), .QN(n11454) );
  NOR2X0 U11459 ( .IN1(n11455), .IN2(n11456), .QN(n11453) );
  NOR2X0 U11460 ( .IN1(g781), .IN2(n11457), .QN(n11456) );
  NOR2X0 U11461 ( .IN1(n5551), .IN2(n11458), .QN(n11455) );
  NAND2X0 U11462 ( .IN1(n2404), .IN2(n11457), .QN(n11458) );
  INVX0 U11463 ( .INP(n2507), .ZN(n11457) );
  NAND2X0 U11464 ( .IN1(n11459), .IN2(n11460), .QN(g34599) );
  NAND2X0 U11465 ( .IN1(n10505), .IN2(g608), .QN(n11460) );
  NOR2X0 U11466 ( .IN1(n11461), .IN2(n11462), .QN(n11459) );
  NOR2X0 U11467 ( .IN1(g613), .IN2(n11463), .QN(n11462) );
  NOR2X0 U11468 ( .IN1(n5474), .IN2(n11464), .QN(n11461) );
  NAND2X0 U11469 ( .IN1(n2421), .IN2(n11463), .QN(n11464) );
  INVX0 U11470 ( .INP(n2509), .ZN(n11463) );
  NAND2X0 U11471 ( .IN1(n11465), .IN2(n11466), .QN(g34598) );
  NAND2X0 U11472 ( .IN1(n10505), .IN2(g550), .QN(n11466) );
  NAND2X0 U11473 ( .IN1(g29221), .IN2(n10385), .QN(n11465) );
  NAND2X0 U11474 ( .IN1(n11467), .IN2(n11468), .QN(g34468) );
  NAND2X0 U11475 ( .IN1(n11469), .IN2(g4854), .QN(n11468) );
  NAND2X0 U11476 ( .IN1(n11470), .IN2(n10385), .QN(n11469) );
  NAND2X0 U11477 ( .IN1(n11471), .IN2(n11472), .QN(n11470) );
  OR2X1 U11478 ( .IN1(n11473), .IN2(n9586), .Q(n11467) );
  NAND2X0 U11479 ( .IN1(n11474), .IN2(n11475), .QN(g34467) );
  NAND2X0 U11480 ( .IN1(n11476), .IN2(n11477), .QN(n11475) );
  XOR2X1 U11481 ( .IN1(g4854), .IN2(n11472), .Q(n11476) );
  AND2X1 U11482 ( .IN1(n2563), .IN2(g4849), .Q(n11472) );
  NAND2X0 U11483 ( .IN1(n10505), .IN2(g4849), .QN(n11474) );
  NAND2X0 U11484 ( .IN1(n11478), .IN2(n11479), .QN(g34466) );
  NAND2X0 U11485 ( .IN1(n11480), .IN2(g4878), .QN(n11479) );
  NAND2X0 U11486 ( .IN1(n11481), .IN2(n10385), .QN(n11480) );
  NAND2X0 U11487 ( .IN1(n9705), .IN2(n11471), .QN(n11481) );
  NAND2X0 U11488 ( .IN1(n11482), .IN2(n5283), .QN(n11478) );
  NOR2X0 U11489 ( .IN1(n9705), .IN2(n11473), .QN(n11482) );
  NAND2X0 U11490 ( .IN1(n11483), .IN2(n11484), .QN(g34465) );
  NAND2X0 U11491 ( .IN1(n10505), .IN2(g4843), .QN(n11484) );
  NOR2X0 U11492 ( .IN1(n11485), .IN2(n11486), .QN(n11483) );
  AND2X1 U11493 ( .IN1(n2567), .IN2(n11477), .Q(n11486) );
  INVX0 U11494 ( .INP(n11473), .ZN(n11477) );
  NOR2X0 U11495 ( .IN1(g4849), .IN2(n11487), .QN(n11485) );
  NAND2X0 U11496 ( .IN1(n11471), .IN2(n2563), .QN(n11487) );
  NAND2X0 U11497 ( .IN1(n11488), .IN2(n11489), .QN(g34464) );
  NAND2X0 U11498 ( .IN1(n11490), .IN2(g4664), .QN(n11489) );
  NAND2X0 U11499 ( .IN1(n11491), .IN2(n10385), .QN(n11490) );
  NAND2X0 U11500 ( .IN1(n11492), .IN2(n11493), .QN(n11491) );
  NAND2X0 U11501 ( .IN1(n11494), .IN2(g4669), .QN(n11488) );
  NAND2X0 U11502 ( .IN1(n11495), .IN2(n11496), .QN(g34463) );
  NAND2X0 U11503 ( .IN1(n11497), .IN2(n11494), .QN(n11496) );
  XOR2X1 U11504 ( .IN1(g4664), .IN2(n11493), .Q(n11497) );
  AND2X1 U11505 ( .IN1(n2573), .IN2(g4659), .Q(n11493) );
  NAND2X0 U11506 ( .IN1(n10505), .IN2(g4659), .QN(n11495) );
  NAND2X0 U11507 ( .IN1(n11498), .IN2(n11499), .QN(g34462) );
  NAND2X0 U11508 ( .IN1(n11500), .IN2(g4688), .QN(n11499) );
  NAND2X0 U11509 ( .IN1(n11501), .IN2(n10385), .QN(n11500) );
  NAND2X0 U11510 ( .IN1(n11492), .IN2(n10133), .QN(n11501) );
  NAND2X0 U11511 ( .IN1(n11502), .IN2(n5656), .QN(n11498) );
  NOR2X0 U11512 ( .IN1(n10133), .IN2(n11503), .QN(n11502) );
  NAND2X0 U11513 ( .IN1(n11504), .IN2(n11505), .QN(g34461) );
  NAND2X0 U11514 ( .IN1(test_so19), .IN2(n10514), .QN(n11505) );
  NOR2X0 U11515 ( .IN1(n11506), .IN2(n11507), .QN(n11504) );
  AND2X1 U11516 ( .IN1(n2577), .IN2(n11494), .Q(n11507) );
  NOR2X0 U11517 ( .IN1(g4659), .IN2(n11508), .QN(n11506) );
  NAND2X0 U11518 ( .IN1(n11492), .IN2(n2573), .QN(n11508) );
  NAND2X0 U11519 ( .IN1(n11509), .IN2(n11510), .QN(g34460) );
  NAND2X0 U11520 ( .IN1(n11511), .IN2(g4639), .QN(n11510) );
  NAND2X0 U11521 ( .IN1(n11512), .IN2(n10385), .QN(n11511) );
  NAND2X0 U11522 ( .IN1(n11513), .IN2(n10138), .QN(n11512) );
  NAND2X0 U11523 ( .IN1(n291), .IN2(test_so3), .QN(n11509) );
  INVX0 U11524 ( .INP(n11514), .ZN(n291) );
  NAND2X0 U11525 ( .IN1(n11515), .IN2(n11516), .QN(g34459) );
  NAND2X0 U11526 ( .IN1(n10505), .IN2(g4643), .QN(n11516) );
  NAND2X0 U11527 ( .IN1(n11517), .IN2(n10385), .QN(n11515) );
  NAND2X0 U11528 ( .IN1(n11518), .IN2(n11519), .QN(n11517) );
  NAND2X0 U11529 ( .IN1(n11520), .IN2(n11521), .QN(n11519) );
  NAND2X0 U11530 ( .IN1(n5653), .IN2(n11522), .QN(n11520) );
  NAND2X0 U11531 ( .IN1(n11523), .IN2(test_so99), .QN(n11522) );
  NOR2X0 U11532 ( .IN1(g4639), .IN2(n10138), .QN(n11523) );
  NAND2X0 U11533 ( .IN1(n11524), .IN2(n11525), .QN(g34458) );
  NAND2X0 U11534 ( .IN1(n11526), .IN2(g4633), .QN(n11525) );
  NAND2X0 U11535 ( .IN1(n11527), .IN2(n11528), .QN(n11526) );
  NAND2X0 U11536 ( .IN1(n11529), .IN2(n11513), .QN(n11528) );
  NOR2X0 U11537 ( .IN1(test_so99), .IN2(n10460), .QN(n11529) );
  INVX0 U11538 ( .INP(n11530), .ZN(n11527) );
  NAND2X0 U11539 ( .IN1(test_so99), .IN2(n11531), .QN(n11524) );
  NAND2X0 U11540 ( .IN1(n11532), .IN2(n10387), .QN(n11531) );
  NAND2X0 U11541 ( .IN1(n11533), .IN2(n11534), .QN(n11532) );
  NOR2X0 U11542 ( .IN1(n5727), .IN2(n10138), .QN(n11534) );
  NOR2X0 U11543 ( .IN1(n11535), .IN2(g4633), .QN(n11533) );
  NAND2X0 U11544 ( .IN1(n11536), .IN2(n11537), .QN(g34457) );
  NAND2X0 U11545 ( .IN1(test_so3), .IN2(n11538), .QN(n11537) );
  NAND2X0 U11546 ( .IN1(n11539), .IN2(n10384), .QN(n11538) );
  NAND2X0 U11547 ( .IN1(n11540), .IN2(n11513), .QN(n11539) );
  NOR2X0 U11548 ( .IN1(test_so99), .IN2(n5727), .QN(n11540) );
  NAND2X0 U11549 ( .IN1(test_so99), .IN2(n11530), .QN(n11536) );
  NAND2X0 U11550 ( .IN1(n11514), .IN2(n11541), .QN(n11530) );
  NAND2X0 U11551 ( .IN1(n11542), .IN2(n11513), .QN(n11541) );
  INVX0 U11552 ( .INP(n11535), .ZN(n11513) );
  NOR2X0 U11553 ( .IN1(test_so3), .IN2(n10460), .QN(n11542) );
  NAND2X0 U11554 ( .IN1(n11543), .IN2(n5727), .QN(n11514) );
  NOR2X0 U11555 ( .IN1(n11544), .IN2(g4643), .QN(n11543) );
  NAND2X0 U11556 ( .IN1(n11545), .IN2(n11546), .QN(g34456) );
  NAND2X0 U11557 ( .IN1(n11547), .IN2(g4608), .QN(n11546) );
  NAND2X0 U11558 ( .IN1(n11548), .IN2(n10384), .QN(n11547) );
  NAND2X0 U11559 ( .IN1(n11549), .IN2(n2590), .QN(n11548) );
  NAND2X0 U11560 ( .IN1(n11550), .IN2(g4616), .QN(n11545) );
  NAND2X0 U11561 ( .IN1(n11551), .IN2(n11552), .QN(g34455) );
  NAND2X0 U11562 ( .IN1(n11553), .IN2(g4322), .QN(n11552) );
  NAND2X0 U11563 ( .IN1(n11554), .IN2(n10384), .QN(n11553) );
  NAND2X0 U11564 ( .IN1(n11555), .IN2(n2594), .QN(n11554) );
  NOR2X0 U11565 ( .IN1(n11556), .IN2(n11557), .QN(n11555) );
  NAND2X0 U11566 ( .IN1(n2595), .IN2(g4332), .QN(n11551) );
  NAND2X0 U11567 ( .IN1(n11558), .IN2(n11559), .QN(g34454) );
  NAND2X0 U11568 ( .IN1(n11560), .IN2(n11550), .QN(n11559) );
  XOR2X1 U11569 ( .IN1(n2590), .IN2(g4608), .Q(n11560) );
  NAND2X0 U11570 ( .IN1(n10505), .IN2(g4601), .QN(n11558) );
  NAND2X0 U11571 ( .IN1(n11561), .IN2(n11562), .QN(g34453) );
  NAND2X0 U11572 ( .IN1(n10505), .IN2(g4593), .QN(n11562) );
  NOR2X0 U11573 ( .IN1(n11563), .IN2(n11564), .QN(n11561) );
  NOR2X0 U11574 ( .IN1(g4601), .IN2(n11565), .QN(n11564) );
  NAND2X0 U11575 ( .IN1(n11549), .IN2(n2598), .QN(n11565) );
  NOR2X0 U11576 ( .IN1(n11556), .IN2(n11566), .QN(n11549) );
  NOR2X0 U11577 ( .IN1(n5365), .IN2(n11567), .QN(n11563) );
  NAND2X0 U11578 ( .IN1(n11550), .IN2(n11568), .QN(n11567) );
  INVX0 U11579 ( .INP(n2598), .ZN(n11568) );
  NAND2X0 U11580 ( .IN1(n11569), .IN2(n11570), .QN(g34452) );
  NAND2X0 U11581 ( .IN1(n11571), .IN2(n11550), .QN(n11570) );
  XOR2X1 U11582 ( .IN1(n10789), .IN2(n5303), .Q(n11571) );
  NAND2X0 U11583 ( .IN1(n10505), .IN2(g4584), .QN(n11569) );
  NAND2X0 U11584 ( .IN1(n11572), .IN2(n11573), .QN(g34451) );
  NAND2X0 U11585 ( .IN1(n11574), .IN2(n11550), .QN(n11573) );
  NOR2X0 U11586 ( .IN1(n11544), .IN2(n11566), .QN(n11550) );
  NOR2X0 U11587 ( .IN1(n10789), .IN2(n5608), .QN(n11566) );
  NAND2X0 U11588 ( .IN1(n11557), .IN2(g4584), .QN(n10789) );
  XOR2X1 U11589 ( .IN1(g4584), .IN2(n11557), .Q(n11574) );
  NAND2X0 U11590 ( .IN1(n10498), .IN2(g4332), .QN(n11572) );
  NAND2X0 U11591 ( .IN1(n11575), .IN2(n11576), .QN(g34450) );
  NAND2X0 U11592 ( .IN1(n10499), .IN2(g4311), .QN(n11576) );
  NOR2X0 U11593 ( .IN1(n11577), .IN2(n11578), .QN(n11575) );
  NOR2X0 U11594 ( .IN1(g4322), .IN2(n11579), .QN(n11578) );
  NAND2X0 U11595 ( .IN1(n2594), .IN2(n11518), .QN(n11579) );
  NOR2X0 U11596 ( .IN1(n5506), .IN2(n11580), .QN(n11577) );
  NAND2X0 U11597 ( .IN1(n2595), .IN2(n11581), .QN(n11580) );
  INVX0 U11598 ( .INP(n2594), .ZN(n11581) );
  NOR2X0 U11599 ( .IN1(n11544), .IN2(n11557), .QN(n2595) );
  AND2X1 U11600 ( .IN1(n11582), .IN2(n2607), .Q(n11557) );
  NOR2X0 U11601 ( .IN1(n11583), .IN2(n5348), .QN(n2607) );
  NOR2X0 U11602 ( .IN1(n5540), .IN2(n5506), .QN(n11582) );
  NAND2X0 U11603 ( .IN1(n11584), .IN2(n11585), .QN(g34448) );
  NAND2X0 U11604 ( .IN1(n11586), .IN2(n11587), .QN(n11585) );
  INVX0 U11605 ( .INP(n11588), .ZN(n11587) );
  NOR2X0 U11606 ( .IN1(n11589), .IN2(n11590), .QN(n11586) );
  NOR2X0 U11607 ( .IN1(n9609), .IN2(n11591), .QN(n11589) );
  NOR2X0 U11608 ( .IN1(n11592), .IN2(n11593), .QN(n11584) );
  NOR2X0 U11609 ( .IN1(n9609), .IN2(n10337), .QN(n11593) );
  NOR2X0 U11610 ( .IN1(n10485), .IN2(n11594), .QN(n11592) );
  NAND2X0 U11611 ( .IN1(n11588), .IN2(g2819), .QN(n11594) );
  NAND2X0 U11612 ( .IN1(n11595), .IN2(n11596), .QN(g34447) );
  NAND2X0 U11613 ( .IN1(n11597), .IN2(n11598), .QN(n11596) );
  INVX0 U11614 ( .INP(n11599), .ZN(n11598) );
  NOR2X0 U11615 ( .IN1(n11600), .IN2(n11590), .QN(n11597) );
  NOR2X0 U11616 ( .IN1(n9608), .IN2(n11591), .QN(n11600) );
  NOR2X0 U11617 ( .IN1(n11601), .IN2(n11602), .QN(n11595) );
  NOR2X0 U11618 ( .IN1(n5404), .IN2(n10328), .QN(n11602) );
  NOR2X0 U11619 ( .IN1(n10485), .IN2(n11603), .QN(n11601) );
  NAND2X0 U11620 ( .IN1(n11599), .IN2(g2807), .QN(n11603) );
  NAND2X0 U11621 ( .IN1(n11604), .IN2(n11605), .QN(g34446) );
  NAND2X0 U11622 ( .IN1(n11606), .IN2(n11607), .QN(n11605) );
  NOR2X0 U11623 ( .IN1(n11608), .IN2(n11590), .QN(n11606) );
  NOR2X0 U11624 ( .IN1(n11591), .IN2(n10149), .QN(n11608) );
  NOR2X0 U11625 ( .IN1(n11609), .IN2(n11610), .QN(n11604) );
  NOR2X0 U11626 ( .IN1(n5609), .IN2(n10328), .QN(n11610) );
  NOR2X0 U11627 ( .IN1(n10485), .IN2(n11611), .QN(n11609) );
  NAND2X0 U11628 ( .IN1(n11612), .IN2(g2815), .QN(n11611) );
  NAND2X0 U11629 ( .IN1(n11613), .IN2(n11614), .QN(g34445) );
  NAND2X0 U11630 ( .IN1(n11615), .IN2(n11616), .QN(n11614) );
  NOR2X0 U11631 ( .IN1(n11617), .IN2(n11590), .QN(n11615) );
  NAND2X0 U11632 ( .IN1(n11618), .IN2(n10384), .QN(n11590) );
  NAND2X0 U11633 ( .IN1(n2760), .IN2(n9255), .QN(n11618) );
  NOR2X0 U11634 ( .IN1(n9605), .IN2(n11591), .QN(n11617) );
  NOR2X0 U11635 ( .IN1(n11619), .IN2(n11620), .QN(n11613) );
  NOR2X0 U11636 ( .IN1(n5379), .IN2(n10328), .QN(n11620) );
  NOR2X0 U11637 ( .IN1(n10485), .IN2(n11621), .QN(n11619) );
  NAND2X0 U11638 ( .IN1(n11622), .IN2(g2803), .QN(n11621) );
  NAND2X0 U11639 ( .IN1(n11623), .IN2(n11624), .QN(g34444) );
  NAND2X0 U11640 ( .IN1(n11625), .IN2(n11626), .QN(n11624) );
  NOR2X0 U11641 ( .IN1(n11627), .IN2(n11588), .QN(n11625) );
  NOR2X0 U11642 ( .IN1(n9606), .IN2(n11591), .QN(n11627) );
  NOR2X0 U11643 ( .IN1(n11628), .IN2(n11629), .QN(n11623) );
  NOR2X0 U11644 ( .IN1(n9606), .IN2(n10328), .QN(n11629) );
  NOR2X0 U11645 ( .IN1(n10485), .IN2(n11630), .QN(n11628) );
  NAND2X0 U11646 ( .IN1(n11588), .IN2(g2787), .QN(n11630) );
  NAND2X0 U11647 ( .IN1(n11631), .IN2(n11632), .QN(n11588) );
  NOR2X0 U11648 ( .IN1(n9780), .IN2(n5301), .QN(n11631) );
  NAND2X0 U11649 ( .IN1(n11633), .IN2(n11634), .QN(g34443) );
  NAND2X0 U11650 ( .IN1(n11635), .IN2(n11626), .QN(n11634) );
  NOR2X0 U11651 ( .IN1(n11636), .IN2(n11599), .QN(n11635) );
  NOR2X0 U11652 ( .IN1(n9604), .IN2(n11591), .QN(n11636) );
  NOR2X0 U11653 ( .IN1(n11637), .IN2(n11638), .QN(n11633) );
  NOR2X0 U11654 ( .IN1(n5403), .IN2(n10329), .QN(n11638) );
  NOR2X0 U11655 ( .IN1(n10485), .IN2(n11639), .QN(n11637) );
  NAND2X0 U11656 ( .IN1(n11599), .IN2(g2775), .QN(n11639) );
  NAND2X0 U11657 ( .IN1(n11640), .IN2(n11632), .QN(n11599) );
  NOR2X0 U11658 ( .IN1(n5301), .IN2(g2729), .QN(n11640) );
  NAND2X0 U11659 ( .IN1(n11641), .IN2(n11642), .QN(g34442) );
  NAND2X0 U11660 ( .IN1(n11643), .IN2(n11626), .QN(n11642) );
  NOR2X0 U11661 ( .IN1(n11644), .IN2(n11612), .QN(n11643) );
  NOR2X0 U11662 ( .IN1(n9607), .IN2(n11591), .QN(n11644) );
  NOR2X0 U11663 ( .IN1(n11645), .IN2(n11646), .QN(n11641) );
  NOR2X0 U11664 ( .IN1(n5610), .IN2(n10329), .QN(n11646) );
  NOR2X0 U11665 ( .IN1(n10485), .IN2(n11647), .QN(n11645) );
  NAND2X0 U11666 ( .IN1(n11612), .IN2(g2783), .QN(n11647) );
  INVX0 U11667 ( .INP(n11607), .ZN(n11612) );
  NOR2X0 U11668 ( .IN1(n11648), .IN2(n11649), .QN(n11607) );
  NAND2X0 U11669 ( .IN1(n11650), .IN2(n11651), .QN(g34441) );
  NAND2X0 U11670 ( .IN1(n11652), .IN2(n11626), .QN(n11651) );
  AND2X1 U11671 ( .IN1(n11653), .IN2(n10365), .Q(n11626) );
  NAND2X0 U11672 ( .IN1(n2760), .IN2(n9265), .QN(n11653) );
  NOR2X0 U11673 ( .IN1(n11654), .IN2(n11622), .QN(n11652) );
  NOR2X0 U11674 ( .IN1(n9610), .IN2(n11591), .QN(n11654) );
  NOR2X0 U11675 ( .IN1(n11655), .IN2(n11656), .QN(n11650) );
  NOR2X0 U11676 ( .IN1(n5378), .IN2(n10329), .QN(n11656) );
  NOR2X0 U11677 ( .IN1(n10485), .IN2(n11657), .QN(n11655) );
  NAND2X0 U11678 ( .IN1(n11622), .IN2(g2771), .QN(n11657) );
  INVX0 U11679 ( .INP(n11616), .ZN(n11622) );
  NOR2X0 U11680 ( .IN1(n11649), .IN2(n11658), .QN(n11616) );
  NAND2X0 U11681 ( .IN1(n11659), .IN2(n11660), .QN(g34440) );
  NAND2X0 U11682 ( .IN1(n10498), .IN2(g446), .QN(n11660) );
  NAND2X0 U11683 ( .IN1(n11661), .IN2(n10383), .QN(n11659) );
  NAND2X0 U11684 ( .IN1(n11662), .IN2(n11663), .QN(n11661) );
  NAND2X0 U11685 ( .IN1(n11664), .IN2(g862), .QN(n11663) );
  NAND2X0 U11686 ( .IN1(g896), .IN2(n11665), .QN(n11664) );
  NAND2X0 U11687 ( .IN1(n11666), .IN2(n11667), .QN(n11665) );
  NAND2X0 U11688 ( .IN1(n5821), .IN2(n11668), .QN(n11666) );
  NAND2X0 U11689 ( .IN1(g890), .IN2(g896), .QN(n11662) );
  NAND2X0 U11690 ( .IN1(n11669), .IN2(n11670), .QN(g34439) );
  NAND2X0 U11691 ( .IN1(n10499), .IN2(g772), .QN(n11670) );
  NOR2X0 U11692 ( .IN1(n11671), .IN2(n11672), .QN(n11669) );
  NOR2X0 U11693 ( .IN1(g776), .IN2(n11673), .QN(n11672) );
  NOR2X0 U11694 ( .IN1(n5330), .IN2(n11674), .QN(n11671) );
  NAND2X0 U11695 ( .IN1(n2404), .IN2(n11673), .QN(n11674) );
  INVX0 U11696 ( .INP(n2554), .ZN(n11673) );
  NAND2X0 U11697 ( .IN1(n11675), .IN2(n11676), .QN(g34438) );
  NAND2X0 U11698 ( .IN1(n10498), .IN2(g604), .QN(n11676) );
  NOR2X0 U11699 ( .IN1(n11677), .IN2(n11678), .QN(n11675) );
  NOR2X0 U11700 ( .IN1(g608), .IN2(n11679), .QN(n11678) );
  NOR2X0 U11701 ( .IN1(n5475), .IN2(n11680), .QN(n11677) );
  NAND2X0 U11702 ( .IN1(n2421), .IN2(n11679), .QN(n11680) );
  INVX0 U11703 ( .INP(n2556), .ZN(n11679) );
  NOR2X0 U11704 ( .IN1(n11681), .IN2(n11682), .QN(g34435) );
  NAND2X0 U11705 ( .IN1(n5711), .IN2(n5416), .QN(n11682) );
  NAND2X0 U11706 ( .IN1(n10034), .IN2(n11683), .QN(n11681) );
  NAND2X0 U11707 ( .IN1(n11684), .IN2(n9739), .QN(n11683) );
  NOR2X0 U11708 ( .IN1(n11685), .IN2(g4141), .QN(n11684) );
  NOR2X0 U11709 ( .IN1(n11686), .IN2(n11687), .QN(n11685) );
  NAND2X0 U11710 ( .IN1(test_so11), .IN2(n5350), .QN(n11687) );
  NAND2X0 U11711 ( .IN1(n11688), .IN2(g4112), .QN(n11686) );
  NAND2X0 U11712 ( .IN1(n2730), .IN2(n11689), .QN(g34425) );
  INVX0 U11713 ( .INP(n10110), .ZN(n11689) );
  NAND2X0 U11714 ( .IN1(n11690), .IN2(n11691), .QN(n10110) );
  NAND2X0 U11715 ( .IN1(n5348), .IN2(n11692), .QN(n11691) );
  NAND2X0 U11716 ( .IN1(n11693), .IN2(n11694), .QN(n11692) );
  NOR2X0 U11717 ( .IN1(n11695), .IN2(n11696), .QN(n11694) );
  NOR2X0 U11718 ( .IN1(n10676), .IN2(n11697), .QN(n11696) );
  NOR2X0 U11719 ( .IN1(n10666), .IN2(n11698), .QN(n11695) );
  NOR2X0 U11720 ( .IN1(n11699), .IN2(n11700), .QN(n11693) );
  NOR2X0 U11721 ( .IN1(n11701), .IN2(n11702), .QN(n11700) );
  NOR2X0 U11722 ( .IN1(n11703), .IN2(n11704), .QN(n11699) );
  NAND2X0 U11723 ( .IN1(n11705), .IN2(g4358), .QN(n11690) );
  NAND2X0 U11724 ( .IN1(n11706), .IN2(n11707), .QN(n11705) );
  NOR2X0 U11725 ( .IN1(n11708), .IN2(n11709), .QN(n11707) );
  NOR2X0 U11726 ( .IN1(n11710), .IN2(n11697), .QN(n11709) );
  NOR2X0 U11727 ( .IN1(n11711), .IN2(n11698), .QN(n11708) );
  NOR2X0 U11728 ( .IN1(n11712), .IN2(n11713), .QN(n11706) );
  NOR2X0 U11729 ( .IN1(n11714), .IN2(n11701), .QN(n11713) );
  NOR2X0 U11730 ( .IN1(n11715), .IN2(n11703), .QN(n11712) );
  AND2X1 U11731 ( .IN1(n11716), .IN2(n11717), .Q(n2730) );
  NAND2X0 U11732 ( .IN1(n11332), .IN2(n11328), .QN(n11717) );
  NAND2X0 U11733 ( .IN1(n11718), .IN2(n11716), .QN(g34383) );
  NOR2X0 U11734 ( .IN1(g34843), .IN2(n11719), .QN(n11718) );
  NOR2X0 U11735 ( .IN1(n11720), .IN2(n11721), .QN(n11719) );
  NAND2X0 U11736 ( .IN1(n11722), .IN2(n11723), .QN(n11721) );
  NOR2X0 U11737 ( .IN1(n11724), .IN2(n11725), .QN(n11722) );
  NAND2X0 U11738 ( .IN1(n11726), .IN2(n11727), .QN(n11720) );
  NOR2X0 U11739 ( .IN1(n11728), .IN2(n11729), .QN(n11727) );
  NOR2X0 U11740 ( .IN1(n11730), .IN2(n11731), .QN(n11726) );
  NAND2X0 U11741 ( .IN1(n11732), .IN2(n11733), .QN(g34843) );
  NOR2X0 U11742 ( .IN1(n11734), .IN2(n11735), .QN(n11733) );
  NAND2X0 U11743 ( .IN1(n11736), .IN2(n11737), .QN(n11735) );
  NAND2X0 U11744 ( .IN1(n11738), .IN2(n5513), .QN(n11737) );
  NAND2X0 U11745 ( .IN1(n11739), .IN2(n5514), .QN(n11736) );
  NAND2X0 U11746 ( .IN1(n11740), .IN2(n11741), .QN(n11734) );
  NAND2X0 U11747 ( .IN1(n11742), .IN2(n5504), .QN(n11741) );
  NOR2X0 U11748 ( .IN1(n5536), .IN2(n11743), .QN(n11742) );
  NAND2X0 U11749 ( .IN1(n11744), .IN2(n5524), .QN(n11740) );
  NOR2X0 U11750 ( .IN1(n11745), .IN2(n11746), .QN(n11732) );
  NAND2X0 U11751 ( .IN1(n11747), .IN2(n11748), .QN(n11746) );
  NAND2X0 U11752 ( .IN1(n11749), .IN2(n11728), .QN(n11748) );
  NAND2X0 U11753 ( .IN1(g31862), .IN2(n11724), .QN(n11747) );
  NAND2X0 U11754 ( .IN1(n11750), .IN2(n11751), .QN(n11745) );
  NAND2X0 U11755 ( .IN1(n11752), .IN2(n11753), .QN(n11751) );
  OR2X1 U11756 ( .IN1(n11754), .IN2(n2727), .Q(n11750) );
  NAND2X0 U11757 ( .IN1(n11755), .IN2(n11756), .QN(g34269) );
  NAND2X0 U11758 ( .IN1(n11757), .IN2(n11758), .QN(n11756) );
  NOR2X0 U11759 ( .IN1(n5614), .IN2(n11759), .QN(n11757) );
  NOR2X0 U11760 ( .IN1(n11760), .IN2(n11761), .QN(n11755) );
  NOR2X0 U11761 ( .IN1(n5770), .IN2(n11762), .QN(n11761) );
  NOR2X0 U11762 ( .IN1(n10487), .IN2(n11763), .QN(n11762) );
  AND2X1 U11763 ( .IN1(n11764), .IN2(n11759), .Q(n11763) );
  NAND2X0 U11764 ( .IN1(n11765), .IN2(n11766), .QN(g34268) );
  NAND2X0 U11765 ( .IN1(n11767), .IN2(n11758), .QN(n11766) );
  NOR2X0 U11766 ( .IN1(n5875), .IN2(n11768), .QN(n11767) );
  NOR2X0 U11767 ( .IN1(n11760), .IN2(n11769), .QN(n11765) );
  NOR2X0 U11768 ( .IN1(n5772), .IN2(n11770), .QN(n11769) );
  NOR2X0 U11769 ( .IN1(n10488), .IN2(n11771), .QN(n11770) );
  AND2X1 U11770 ( .IN1(n11764), .IN2(n11768), .Q(n11771) );
  NAND2X0 U11771 ( .IN1(n11772), .IN2(n11773), .QN(g34267) );
  NAND2X0 U11772 ( .IN1(n11774), .IN2(g4939), .QN(n11773) );
  NAND2X0 U11773 ( .IN1(n11775), .IN2(n10383), .QN(n11774) );
  NAND2X0 U11774 ( .IN1(n11776), .IN2(n11764), .QN(n11775) );
  NOR2X0 U11775 ( .IN1(n11760), .IN2(n11777), .QN(n11772) );
  NOR2X0 U11776 ( .IN1(n11778), .IN2(n11779), .QN(n11777) );
  OR2X1 U11777 ( .IN1(n11776), .IN2(n5878), .Q(n11779) );
  NAND2X0 U11778 ( .IN1(n11780), .IN2(n11781), .QN(g34266) );
  NAND2X0 U11779 ( .IN1(n11782), .IN2(n11758), .QN(n11781) );
  INVX0 U11780 ( .INP(n11778), .ZN(n11758) );
  NAND2X0 U11781 ( .IN1(n11764), .IN2(n10383), .QN(n11778) );
  NOR2X0 U11782 ( .IN1(n5863), .IN2(n11783), .QN(n11782) );
  NOR2X0 U11783 ( .IN1(n11760), .IN2(n11784), .QN(n11780) );
  NOR2X0 U11784 ( .IN1(n5774), .IN2(n11785), .QN(n11784) );
  NOR2X0 U11785 ( .IN1(n10488), .IN2(n11786), .QN(n11785) );
  NOR2X0 U11786 ( .IN1(n11787), .IN2(n11333), .QN(n11786) );
  INVX0 U11787 ( .INP(n11783), .ZN(n11333) );
  AND2X1 U11788 ( .IN1(n11788), .IN2(n11787), .Q(n11760) );
  INVX0 U11789 ( .INP(n11764), .ZN(n11787) );
  NAND2X0 U11790 ( .IN1(n11789), .IN2(n5637), .QN(n11764) );
  NOR2X0 U11791 ( .IN1(test_so46), .IN2(n11790), .QN(n11789) );
  NOR2X0 U11792 ( .IN1(n18464), .IN2(n10459), .QN(n11788) );
  NOR2X0 U11793 ( .IN1(n10732), .IN2(n11473), .QN(g34265) );
  NAND2X0 U11794 ( .IN1(n11471), .IN2(n10383), .QN(n11473) );
  NOR2X0 U11795 ( .IN1(n11791), .IN2(n11331), .QN(n11471) );
  NAND2X0 U11796 ( .IN1(n11792), .IN2(n5713), .QN(n10732) );
  NOR2X0 U11797 ( .IN1(g4864), .IN2(g4871), .QN(n11792) );
  NAND2X0 U11798 ( .IN1(n11793), .IN2(n11794), .QN(g34264) );
  NAND2X0 U11799 ( .IN1(n11795), .IN2(n11796), .QN(n11794) );
  NOR2X0 U11800 ( .IN1(n5613), .IN2(n11797), .QN(n11795) );
  NOR2X0 U11801 ( .IN1(n11798), .IN2(n11799), .QN(n11793) );
  NOR2X0 U11802 ( .IN1(n5769), .IN2(n11800), .QN(n11799) );
  NOR2X0 U11803 ( .IN1(n10489), .IN2(n11801), .QN(n11800) );
  AND2X1 U11804 ( .IN1(n11802), .IN2(n11797), .Q(n11801) );
  NAND2X0 U11805 ( .IN1(n11803), .IN2(n11804), .QN(g34263) );
  NAND2X0 U11806 ( .IN1(n11805), .IN2(n11796), .QN(n11804) );
  NOR2X0 U11807 ( .IN1(n5877), .IN2(n11806), .QN(n11805) );
  NOR2X0 U11808 ( .IN1(n11798), .IN2(n11807), .QN(n11803) );
  NOR2X0 U11809 ( .IN1(n5775), .IN2(n11808), .QN(n11807) );
  NOR2X0 U11810 ( .IN1(n10490), .IN2(n11809), .QN(n11808) );
  AND2X1 U11811 ( .IN1(n11802), .IN2(n11806), .Q(n11809) );
  NAND2X0 U11812 ( .IN1(n11810), .IN2(n11811), .QN(g34262) );
  NAND2X0 U11813 ( .IN1(test_so18), .IN2(n11812), .QN(n11811) );
  NAND2X0 U11814 ( .IN1(n11813), .IN2(n10383), .QN(n11812) );
  NAND2X0 U11815 ( .IN1(n11814), .IN2(n11802), .QN(n11813) );
  NOR2X0 U11816 ( .IN1(n11798), .IN2(n11815), .QN(n11810) );
  NOR2X0 U11817 ( .IN1(n11816), .IN2(n11817), .QN(n11815) );
  OR2X1 U11818 ( .IN1(n11814), .IN2(n5876), .Q(n11817) );
  NAND2X0 U11819 ( .IN1(n11818), .IN2(n11819), .QN(g34261) );
  NAND2X0 U11820 ( .IN1(n11820), .IN2(n11796), .QN(n11819) );
  INVX0 U11821 ( .INP(n11816), .ZN(n11796) );
  NAND2X0 U11822 ( .IN1(n11802), .IN2(n10382), .QN(n11816) );
  NOR2X0 U11823 ( .IN1(n5862), .IN2(n11821), .QN(n11820) );
  NOR2X0 U11824 ( .IN1(n11798), .IN2(n11822), .QN(n11818) );
  NOR2X0 U11825 ( .IN1(n5771), .IN2(n11823), .QN(n11822) );
  NOR2X0 U11826 ( .IN1(n10491), .IN2(n11824), .QN(n11823) );
  NOR2X0 U11827 ( .IN1(n11825), .IN2(n11329), .QN(n11824) );
  INVX0 U11828 ( .INP(n11821), .ZN(n11329) );
  AND2X1 U11829 ( .IN1(n11826), .IN2(n11825), .Q(n11798) );
  INVX0 U11830 ( .INP(n11802), .ZN(n11825) );
  NAND2X0 U11831 ( .IN1(n11827), .IN2(n18466), .QN(n11802) );
  NOR2X0 U11832 ( .IN1(n11790), .IN2(g4818), .QN(n11827) );
  NOR2X0 U11833 ( .IN1(n18465), .IN2(n10458), .QN(n11826) );
  NOR2X0 U11834 ( .IN1(n11828), .IN2(n11829), .QN(g34260) );
  NAND2X0 U11835 ( .IN1(n11494), .IN2(n5712), .QN(n11829) );
  INVX0 U11836 ( .INP(n11503), .ZN(n11494) );
  NAND2X0 U11837 ( .IN1(n11492), .IN2(n10382), .QN(n11503) );
  NOR2X0 U11838 ( .IN1(n11830), .IN2(n11327), .QN(n11492) );
  NAND2X0 U11839 ( .IN1(n5440), .IN2(n10040), .QN(n11828) );
  NOR2X0 U11840 ( .IN1(n5844), .IN2(n11831), .QN(g34259) );
  NOR2X0 U11841 ( .IN1(n10496), .IN2(n11832), .QN(n11831) );
  NOR2X0 U11842 ( .IN1(n11535), .IN2(n11833), .QN(n11832) );
  NAND2X0 U11843 ( .IN1(test_so3), .IN2(n5727), .QN(n11833) );
  NAND2X0 U11844 ( .IN1(n5382), .IN2(n11518), .QN(n11535) );
  NAND2X0 U11845 ( .IN1(n11834), .IN2(n11835), .QN(g34258) );
  NAND2X0 U11846 ( .IN1(test_so81), .IN2(n10515), .QN(n11835) );
  NOR2X0 U11847 ( .IN1(n11836), .IN2(n11837), .QN(n11834) );
  NOR2X0 U11848 ( .IN1(g4358), .IN2(n11838), .QN(n11837) );
  OR2X1 U11849 ( .IN1(n11583), .IN2(n11556), .Q(n11838) );
  INVX0 U11850 ( .INP(n11518), .ZN(n11556) );
  NOR2X0 U11851 ( .IN1(n5348), .IN2(n11839), .QN(n11836) );
  NAND2X0 U11852 ( .IN1(n11840), .IN2(n11583), .QN(n11839) );
  NAND2X0 U11853 ( .IN1(test_so81), .IN2(n11841), .QN(n11583) );
  NAND2X0 U11854 ( .IN1(n11842), .IN2(n11843), .QN(g34257) );
  NAND2X0 U11855 ( .IN1(n10497), .IN2(g4340), .QN(n11843) );
  NOR2X0 U11856 ( .IN1(n11844), .IN2(n11845), .QN(n11842) );
  NOR2X0 U11857 ( .IN1(n11521), .IN2(n11846), .QN(n11845) );
  NAND2X0 U11858 ( .IN1(n11518), .IN2(n10132), .QN(n11846) );
  NOR2X0 U11859 ( .IN1(n11841), .IN2(n11847), .QN(n11844) );
  NAND2X0 U11860 ( .IN1(test_so81), .IN2(n11840), .QN(n11847) );
  INVX0 U11861 ( .INP(n11544), .ZN(n11840) );
  NAND2X0 U11862 ( .IN1(n11518), .IN2(n10382), .QN(n11544) );
  NAND2X0 U11863 ( .IN1(n9281), .IN2(n11848), .QN(n11518) );
  NAND2X0 U11864 ( .IN1(n11849), .IN2(n1289), .QN(n11848) );
  INVX0 U11865 ( .INP(n11521), .ZN(n11841) );
  NAND2X0 U11866 ( .IN1(test_so99), .IN2(n11850), .QN(n11521) );
  NAND2X0 U11867 ( .IN1(n11851), .IN2(n11852), .QN(g34256) );
  OR2X1 U11868 ( .IN1(n10308), .IN2(n9911), .Q(n11852) );
  NAND2X0 U11869 ( .IN1(n11853), .IN2(n10382), .QN(n11851) );
  NAND2X0 U11870 ( .IN1(n11854), .IN2(n5765), .QN(n11853) );
  NOR2X0 U11871 ( .IN1(n11855), .IN2(n11856), .QN(n11854) );
  NOR2X0 U11872 ( .IN1(n9703), .IN2(g4462), .QN(n11856) );
  NAND2X0 U11873 ( .IN1(n11857), .IN2(n11858), .QN(g34255) );
  NOR2X0 U11874 ( .IN1(n10495), .IN2(n11855), .QN(n11858) );
  NOR2X0 U11875 ( .IN1(n11859), .IN2(g4462), .QN(n11857) );
  NOR2X0 U11876 ( .IN1(n9703), .IN2(n10142), .QN(n11859) );
  NAND2X0 U11877 ( .IN1(n11860), .IN2(n11861), .QN(g34254) );
  NAND2X0 U11878 ( .IN1(n11862), .IN2(g4473), .QN(n11861) );
  NAND2X0 U11879 ( .IN1(n11863), .IN2(n11864), .QN(n11862) );
  NOR2X0 U11880 ( .IN1(test_so38), .IN2(n5671), .QN(n11864) );
  NOR2X0 U11881 ( .IN1(n5382), .IN2(n10458), .QN(n11863) );
  NAND2X0 U11882 ( .IN1(n11855), .IN2(n10382), .QN(n11860) );
  INVX0 U11883 ( .INP(n11865), .ZN(n11855) );
  NOR2X0 U11884 ( .IN1(n10493), .IN2(n11866), .QN(g34253) );
  NOR2X0 U11885 ( .IN1(n10142), .IN2(n11867), .QN(n11866) );
  NAND2X0 U11886 ( .IN1(n11865), .IN2(g4462), .QN(n11867) );
  NAND2X0 U11887 ( .IN1(n11868), .IN2(n5849), .QN(n11865) );
  NOR2X0 U11888 ( .IN1(n9788), .IN2(n11869), .QN(n11868) );
  NOR2X0 U11889 ( .IN1(n11870), .IN2(n11184), .QN(n11869) );
  AND2X1 U11890 ( .IN1(n2668), .IN2(n5846), .Q(n11870) );
  NAND2X0 U11891 ( .IN1(n11871), .IN2(n11872), .QN(g34252) );
  NAND2X0 U11892 ( .IN1(n10498), .IN2(g767), .QN(n11872) );
  NOR2X0 U11893 ( .IN1(n11873), .IN2(n11874), .QN(n11871) );
  NOR2X0 U11894 ( .IN1(g772), .IN2(n11875), .QN(n11874) );
  NOR2X0 U11895 ( .IN1(n5334), .IN2(n11876), .QN(n11873) );
  NAND2X0 U11896 ( .IN1(n2404), .IN2(n11875), .QN(n11876) );
  INVX0 U11897 ( .INP(n2647), .ZN(n11875) );
  NAND2X0 U11898 ( .IN1(n11877), .IN2(n11878), .QN(g34251) );
  NAND2X0 U11899 ( .IN1(n10498), .IN2(g599), .QN(n11878) );
  NOR2X0 U11900 ( .IN1(n11879), .IN2(n11880), .QN(n11877) );
  NOR2X0 U11901 ( .IN1(g604), .IN2(n11881), .QN(n11880) );
  NOR2X0 U11902 ( .IN1(n5473), .IN2(n11882), .QN(n11879) );
  NAND2X0 U11903 ( .IN1(n2421), .IN2(n11881), .QN(n11882) );
  INVX0 U11904 ( .INP(n2649), .ZN(n11881) );
  NAND2X0 U11905 ( .IN1(n11883), .IN2(n11884), .QN(g34250) );
  NAND2X0 U11906 ( .IN1(n10498), .IN2(g298), .QN(n11884) );
  NOR2X0 U11907 ( .IN1(n11885), .IN2(n11886), .QN(n11883) );
  NOR2X0 U11908 ( .IN1(n11887), .IN2(g142), .QN(n11886) );
  NOR2X0 U11909 ( .IN1(n5724), .IN2(n11888), .QN(n11885) );
  NAND2X0 U11910 ( .IN1(n10106), .IN2(n11887), .QN(n11888) );
  NAND2X0 U11911 ( .IN1(n11889), .IN2(n11890), .QN(g34249) );
  NAND2X0 U11912 ( .IN1(n10499), .IN2(g157), .QN(n11890) );
  NOR2X0 U11913 ( .IN1(n11891), .IN2(n11892), .QN(n11889) );
  AND2X1 U11914 ( .IN1(n5843), .IN2(n2710), .Q(n11892) );
  NOR2X0 U11915 ( .IN1(n5843), .IN2(n11893), .QN(n11891) );
  NAND2X0 U11916 ( .IN1(n11894), .IN2(n11895), .QN(n11893) );
  INVX0 U11917 ( .INP(n2710), .ZN(n11895) );
  NAND2X0 U11918 ( .IN1(n11896), .IN2(n11716), .QN(g34201) );
  NOR2X0 U11919 ( .IN1(g34781), .IN2(n11897), .QN(n11896) );
  NOR2X0 U11920 ( .IN1(n11898), .IN2(n11899), .QN(n11897) );
  NAND2X0 U11921 ( .IN1(n11900), .IN2(n11901), .QN(n11899) );
  NOR2X0 U11922 ( .IN1(n11902), .IN2(n11903), .QN(n11901) );
  NOR2X0 U11923 ( .IN1(n11904), .IN2(n11905), .QN(n11900) );
  NAND2X0 U11924 ( .IN1(n11906), .IN2(n11907), .QN(n11898) );
  NOR2X0 U11925 ( .IN1(n3005), .IN2(n11908), .QN(n11907) );
  NOR2X0 U11926 ( .IN1(n11909), .IN2(n11910), .QN(n11906) );
  NAND2X0 U11927 ( .IN1(n11911), .IN2(n11912), .QN(g34781) );
  NOR2X0 U11928 ( .IN1(n11913), .IN2(n11914), .QN(n11912) );
  NAND2X0 U11929 ( .IN1(n11915), .IN2(n11916), .QN(n11914) );
  NAND2X0 U11930 ( .IN1(n11917), .IN2(n5511), .QN(n11916) );
  NOR2X0 U11931 ( .IN1(n3550), .IN2(n10126), .QN(n11917) );
  NAND2X0 U11932 ( .IN1(n11918), .IN2(n5512), .QN(n11915) );
  NOR2X0 U11933 ( .IN1(n10045), .IN2(n3569), .QN(n11918) );
  NAND2X0 U11934 ( .IN1(n11919), .IN2(n11920), .QN(n11913) );
  NAND2X0 U11935 ( .IN1(n11921), .IN2(n5508), .QN(n11920) );
  NOR2X0 U11936 ( .IN1(n10042), .IN2(n3006), .QN(n11921) );
  NAND2X0 U11937 ( .IN1(n11922), .IN2(n5509), .QN(n11919) );
  NOR2X0 U11938 ( .IN1(n10043), .IN2(n3007), .QN(n11922) );
  NOR2X0 U11939 ( .IN1(n11923), .IN2(n11924), .QN(n11911) );
  NAND2X0 U11940 ( .IN1(n11925), .IN2(n11926), .QN(n11924) );
  NAND2X0 U11941 ( .IN1(n11927), .IN2(n5359), .QN(n11926) );
  NOR2X0 U11942 ( .IN1(n5596), .IN2(n1282), .QN(n11927) );
  INVX0 U11943 ( .INP(n3005), .ZN(n1282) );
  NAND2X0 U11944 ( .IN1(g31863), .IN2(n11908), .QN(n11925) );
  NAND2X0 U11945 ( .IN1(n11928), .IN2(n11929), .QN(n11923) );
  NAND2X0 U11946 ( .IN1(n11930), .IN2(n5507), .QN(n11929) );
  NOR2X0 U11947 ( .IN1(n10041), .IN2(n3588), .QN(n11930) );
  NAND2X0 U11948 ( .IN1(n11931), .IN2(n5510), .QN(n11928) );
  NOR2X0 U11949 ( .IN1(n10044), .IN2(n3606), .QN(n11931) );
  NAND2X0 U11950 ( .IN1(n11932), .IN2(n11933), .QN(g34041) );
  NAND2X0 U11951 ( .IN1(n11934), .IN2(n11935), .QN(n11933) );
  XOR2X1 U11952 ( .IN1(n11936), .IN2(n5367), .Q(n11934) );
  OR2X1 U11953 ( .IN1(n10308), .IN2(n5637), .Q(n11932) );
  NAND2X0 U11954 ( .IN1(n11937), .IN2(n11938), .QN(g34040) );
  NAND2X0 U11955 ( .IN1(n10499), .IN2(g4975), .QN(n11938) );
  NOR2X0 U11956 ( .IN1(n11939), .IN2(n11940), .QN(n11937) );
  NOR2X0 U11957 ( .IN1(n5517), .IN2(n11941), .QN(n11940) );
  NOR2X0 U11958 ( .IN1(n11791), .IN2(n11942), .QN(n11939) );
  NOR2X0 U11959 ( .IN1(n11943), .IN2(n11944), .QN(n11942) );
  NOR2X0 U11960 ( .IN1(n10491), .IN2(n10744), .QN(n11944) );
  NOR2X0 U11961 ( .IN1(n10743), .IN2(n11945), .QN(n11943) );
  NAND2X0 U11962 ( .IN1(n11946), .IN2(n11947), .QN(g34039) );
  NAND2X0 U11963 ( .IN1(test_so58), .IN2(n11948), .QN(n11947) );
  NAND2X0 U11964 ( .IN1(n11949), .IN2(n10382), .QN(n11948) );
  NAND2X0 U11965 ( .IN1(n11935), .IN2(g4966), .QN(n11946) );
  NAND2X0 U11966 ( .IN1(n11950), .IN2(n11951), .QN(g34038) );
  NAND2X0 U11967 ( .IN1(n10510), .IN2(g4983), .QN(n11951) );
  NOR2X0 U11968 ( .IN1(n11952), .IN2(n11953), .QN(n11950) );
  NOR2X0 U11969 ( .IN1(n10123), .IN2(n11954), .QN(n11953) );
  NAND2X0 U11970 ( .IN1(n11935), .IN2(n11955), .QN(n11954) );
  INVX0 U11971 ( .INP(n11941), .ZN(n11935) );
  NOR2X0 U11972 ( .IN1(test_so58), .IN2(n11949), .QN(n11952) );
  NAND2X0 U11973 ( .IN1(n11956), .IN2(n11957), .QN(n11949) );
  NOR2X0 U11974 ( .IN1(n11791), .IN2(n11958), .QN(n11956) );
  NAND2X0 U11975 ( .IN1(n11959), .IN2(n11960), .QN(g34037) );
  NAND2X0 U11976 ( .IN1(n10510), .IN2(g4966), .QN(n11960) );
  NOR2X0 U11977 ( .IN1(n11961), .IN2(n11962), .QN(n11959) );
  NOR2X0 U11978 ( .IN1(g4975), .IN2(n11963), .QN(n11962) );
  NAND2X0 U11979 ( .IN1(n11958), .IN2(n11964), .QN(n11963) );
  INVX0 U11980 ( .INP(n11945), .ZN(n11958) );
  NOR2X0 U11981 ( .IN1(n5360), .IN2(n11941), .QN(n11961) );
  NAND2X0 U11982 ( .IN1(n11965), .IN2(n11945), .QN(n11941) );
  NAND2X0 U11983 ( .IN1(n11957), .IN2(g4966), .QN(n11945) );
  INVX0 U11984 ( .INP(n11955), .ZN(n11957) );
  NAND2X0 U11985 ( .IN1(n11331), .IN2(g4983), .QN(n11955) );
  INVX0 U11986 ( .INP(n11936), .ZN(n11331) );
  NAND2X0 U11987 ( .IN1(n11966), .IN2(n11967), .QN(n11936) );
  NOR2X0 U11988 ( .IN1(n9705), .IN2(n9586), .QN(n11967) );
  NOR2X0 U11989 ( .IN1(n5283), .IN2(n10063), .QN(n11966) );
  NOR2X0 U11990 ( .IN1(n10492), .IN2(n11791), .QN(n11965) );
  INVX0 U11991 ( .INP(n11964), .ZN(n11791) );
  NOR2X0 U11992 ( .IN1(n5443), .IN2(n11968), .QN(g34036) );
  NOR2X0 U11993 ( .IN1(n5318), .IN2(n11968), .QN(g34035) );
  NOR2X0 U11994 ( .IN1(n5713), .IN2(n11968), .QN(g34034) );
  NOR2X0 U11995 ( .IN1(n11964), .IN2(n10458), .QN(n11968) );
  NAND2X0 U11996 ( .IN1(n11969), .IN2(n11970), .QN(n11964) );
  NAND2X0 U11997 ( .IN1(n11971), .IN2(n11972), .QN(g34033) );
  NAND2X0 U11998 ( .IN1(n11973), .IN2(n11974), .QN(n11972) );
  XOR2X1 U11999 ( .IN1(n11975), .IN2(n5368), .Q(n11973) );
  NAND2X0 U12000 ( .IN1(n10510), .IN2(g4818), .QN(n11971) );
  NAND2X0 U12001 ( .IN1(n11976), .IN2(n11977), .QN(g34032) );
  NAND2X0 U12002 ( .IN1(n10510), .IN2(g4785), .QN(n11977) );
  NOR2X0 U12003 ( .IN1(n11978), .IN2(n11979), .QN(n11976) );
  NOR2X0 U12004 ( .IN1(n5518), .IN2(n11980), .QN(n11979) );
  NOR2X0 U12005 ( .IN1(n11830), .IN2(n11981), .QN(n11978) );
  NOR2X0 U12006 ( .IN1(n11982), .IN2(n11983), .QN(n11981) );
  NOR2X0 U12007 ( .IN1(n10492), .IN2(n10713), .QN(n11983) );
  NOR2X0 U12008 ( .IN1(n10714), .IN2(n11984), .QN(n11982) );
  NAND2X0 U12009 ( .IN1(n11985), .IN2(n11986), .QN(g34031) );
  NAND2X0 U12010 ( .IN1(test_so29), .IN2(n11987), .QN(n11986) );
  NAND2X0 U12011 ( .IN1(n11988), .IN2(n10382), .QN(n11987) );
  NAND2X0 U12012 ( .IN1(n11974), .IN2(g4776), .QN(n11985) );
  NAND2X0 U12013 ( .IN1(n11989), .IN2(n11990), .QN(g34030) );
  NAND2X0 U12014 ( .IN1(n10511), .IN2(g4793), .QN(n11990) );
  NOR2X0 U12015 ( .IN1(n11991), .IN2(n11992), .QN(n11989) );
  NOR2X0 U12016 ( .IN1(n10125), .IN2(n11993), .QN(n11992) );
  NAND2X0 U12017 ( .IN1(n11974), .IN2(n11994), .QN(n11993) );
  INVX0 U12018 ( .INP(n11980), .ZN(n11974) );
  NOR2X0 U12019 ( .IN1(test_so29), .IN2(n11988), .QN(n11991) );
  NAND2X0 U12020 ( .IN1(n11995), .IN2(n11996), .QN(n11988) );
  NOR2X0 U12021 ( .IN1(n11830), .IN2(n11997), .QN(n11995) );
  NAND2X0 U12022 ( .IN1(n11998), .IN2(n11999), .QN(g34029) );
  NAND2X0 U12023 ( .IN1(n10511), .IN2(g4776), .QN(n11999) );
  NOR2X0 U12024 ( .IN1(n12000), .IN2(n12001), .QN(n11998) );
  NOR2X0 U12025 ( .IN1(g4785), .IN2(n12002), .QN(n12001) );
  NAND2X0 U12026 ( .IN1(n11997), .IN2(n12003), .QN(n12002) );
  INVX0 U12027 ( .INP(n11984), .ZN(n11997) );
  NOR2X0 U12028 ( .IN1(n5361), .IN2(n11980), .QN(n12000) );
  NAND2X0 U12029 ( .IN1(n12004), .IN2(n11984), .QN(n11980) );
  NAND2X0 U12030 ( .IN1(n11996), .IN2(g4776), .QN(n11984) );
  INVX0 U12031 ( .INP(n11994), .ZN(n11996) );
  NAND2X0 U12032 ( .IN1(n11327), .IN2(g4793), .QN(n11994) );
  INVX0 U12033 ( .INP(n11975), .ZN(n11327) );
  NAND2X0 U12034 ( .IN1(n12005), .IN2(n12006), .QN(n11975) );
  NOR2X0 U12035 ( .IN1(n9590), .IN2(n5656), .QN(n12006) );
  NOR2X0 U12036 ( .IN1(n10064), .IN2(n10133), .QN(n12005) );
  NOR2X0 U12037 ( .IN1(n10492), .IN2(n11830), .QN(n12004) );
  INVX0 U12038 ( .INP(n12003), .ZN(n11830) );
  NOR2X0 U12039 ( .IN1(n5440), .IN2(n2774), .QN(g34027) );
  NOR2X0 U12040 ( .IN1(n5712), .IN2(n2774), .QN(g34026) );
  NOR2X0 U12041 ( .IN1(n12003), .IN2(n10457), .QN(n2774) );
  NAND2X0 U12042 ( .IN1(n11969), .IN2(n12007), .QN(n12003) );
  NOR2X0 U12043 ( .IN1(n9738), .IN2(n1289), .QN(n11969) );
  NAND2X0 U12044 ( .IN1(n12008), .IN2(n12009), .QN(g34024) );
  NOR2X0 U12045 ( .IN1(n12010), .IN2(n12011), .QN(n12009) );
  NOR2X0 U12046 ( .IN1(n10492), .IN2(n12012), .QN(n12011) );
  NOR2X0 U12047 ( .IN1(n12013), .IN2(n12014), .QN(n12012) );
  NOR2X0 U12048 ( .IN1(n11184), .IN2(n12015), .QN(n12014) );
  NOR2X0 U12049 ( .IN1(n9768), .IN2(n11849), .QN(n12013) );
  NOR2X0 U12050 ( .IN1(n10061), .IN2(n10329), .QN(n12010) );
  NAND2X0 U12051 ( .IN1(n12016), .IN2(n12008), .QN(g34023) );
  NOR2X0 U12052 ( .IN1(n12017), .IN2(n12018), .QN(n12008) );
  AND2X1 U12053 ( .IN1(n12019), .IN2(n11849), .Q(n12018) );
  NOR2X0 U12054 ( .IN1(n10074), .IN2(n10457), .QN(n12019) );
  NOR2X0 U12055 ( .IN1(n12020), .IN2(n12021), .QN(n12016) );
  NOR2X0 U12056 ( .IN1(n18467), .IN2(n12022), .QN(n12021) );
  NOR2X0 U12057 ( .IN1(n10493), .IN2(n12023), .QN(n12022) );
  NOR2X0 U12058 ( .IN1(n12024), .IN2(n12025), .QN(n12023) );
  NAND2X0 U12059 ( .IN1(n11849), .IN2(g4555), .QN(n12025) );
  NAND2X0 U12060 ( .IN1(g4558), .IN2(g4561), .QN(n12024) );
  NOR2X0 U12061 ( .IN1(n11849), .IN2(n12026), .QN(n12020) );
  NAND2X0 U12062 ( .IN1(n10368), .IN2(g4552), .QN(n12026) );
  NAND2X0 U12063 ( .IN1(n12027), .IN2(n12028), .QN(g34022) );
  NOR2X0 U12064 ( .IN1(n12029), .IN2(n12030), .QN(n12028) );
  NOR2X0 U12065 ( .IN1(n9582), .IN2(n10329), .QN(n12030) );
  NOR2X0 U12066 ( .IN1(n10493), .IN2(n12031), .QN(n12029) );
  NAND2X0 U12067 ( .IN1(n12032), .IN2(g2763), .QN(n12031) );
  NOR2X0 U12068 ( .IN1(n2787), .IN2(n12033), .QN(n12027) );
  NOR2X0 U12069 ( .IN1(g2763), .IN2(n12032), .QN(n12033) );
  OR2X1 U12070 ( .IN1(n12034), .IN2(n9582), .Q(n12032) );
  NAND2X0 U12071 ( .IN1(n12035), .IN2(n12036), .QN(g34021) );
  NAND2X0 U12072 ( .IN1(n10511), .IN2(g2648), .QN(n12036) );
  NOR2X0 U12073 ( .IN1(n12037), .IN2(n12038), .QN(n12035) );
  NOR2X0 U12074 ( .IN1(n9622), .IN2(n12039), .QN(n12038) );
  NOR2X0 U12075 ( .IN1(n12040), .IN2(n12041), .QN(n12037) );
  NAND2X0 U12076 ( .IN1(n12042), .IN2(n12043), .QN(g34020) );
  NAND2X0 U12077 ( .IN1(n12044), .IN2(n12045), .QN(n12043) );
  NOR2X0 U12078 ( .IN1(n9693), .IN2(n12046), .QN(n12044) );
  NOR2X0 U12079 ( .IN1(n12047), .IN2(g2629), .QN(n12046) );
  NOR2X0 U12080 ( .IN1(n12048), .IN2(n12049), .QN(n12042) );
  NOR2X0 U12081 ( .IN1(n10493), .IN2(n12050), .QN(n12049) );
  NOR2X0 U12082 ( .IN1(n12051), .IN2(n12052), .QN(n12050) );
  NOR2X0 U12083 ( .IN1(n9693), .IN2(n12053), .QN(n12052) );
  NOR2X0 U12084 ( .IN1(n12045), .IN2(n12054), .QN(n12051) );
  NOR2X0 U12085 ( .IN1(n12055), .IN2(n12056), .QN(n12054) );
  NOR2X0 U12086 ( .IN1(n12057), .IN2(g2643), .QN(n12055) );
  AND2X1 U12087 ( .IN1(n12058), .IN2(n12059), .Q(n12045) );
  NAND2X0 U12088 ( .IN1(n5755), .IN2(n12060), .QN(n12059) );
  NOR2X0 U12089 ( .IN1(n5521), .IN2(n10329), .QN(n12048) );
  NAND2X0 U12090 ( .IN1(n12061), .IN2(n12062), .QN(g34019) );
  OR2X1 U12091 ( .IN1(n12063), .IN2(n12040), .Q(n12062) );
  NOR2X0 U12092 ( .IN1(n12064), .IN2(n12065), .QN(n12061) );
  NOR2X0 U12093 ( .IN1(n5787), .IN2(n10329), .QN(n12065) );
  NOR2X0 U12094 ( .IN1(n10494), .IN2(n12066), .QN(n12064) );
  NAND2X0 U12095 ( .IN1(n12063), .IN2(g2583), .QN(n12066) );
  NAND2X0 U12096 ( .IN1(n12067), .IN2(g2629), .QN(n12063) );
  NAND2X0 U12097 ( .IN1(n12068), .IN2(n12069), .QN(g34018) );
  OR2X1 U12098 ( .IN1(n12070), .IN2(n12040), .Q(n12069) );
  NOR2X0 U12099 ( .IN1(n12071), .IN2(n12072), .QN(n12068) );
  NOR2X0 U12100 ( .IN1(n5800), .IN2(n10330), .QN(n12072) );
  NOR2X0 U12101 ( .IN1(n10494), .IN2(n12073), .QN(n12071) );
  NAND2X0 U12102 ( .IN1(test_so61), .IN2(n12070), .QN(n12073) );
  NAND2X0 U12103 ( .IN1(n12074), .IN2(n5351), .QN(n12070) );
  NAND2X0 U12104 ( .IN1(n12075), .IN2(n12076), .QN(g34017) );
  OR2X1 U12105 ( .IN1(n12077), .IN2(n12040), .Q(n12076) );
  NOR2X0 U12106 ( .IN1(n12078), .IN2(n12079), .QN(n12075) );
  AND2X1 U12107 ( .IN1(n10496), .IN2(test_so61), .Q(n12079) );
  NOR2X0 U12108 ( .IN1(n10494), .IN2(n12080), .QN(n12078) );
  NAND2X0 U12109 ( .IN1(test_so66), .IN2(n12077), .QN(n12080) );
  NAND2X0 U12110 ( .IN1(n12081), .IN2(n12053), .QN(n12077) );
  NOR2X0 U12111 ( .IN1(n5521), .IN2(n5351), .QN(n12081) );
  NAND2X0 U12112 ( .IN1(n12082), .IN2(n12083), .QN(g34016) );
  OR2X1 U12113 ( .IN1(n12084), .IN2(n12040), .Q(n12083) );
  NOR2X0 U12114 ( .IN1(n12085), .IN2(n12086), .QN(n12082) );
  NOR2X0 U12115 ( .IN1(n5816), .IN2(n10330), .QN(n12086) );
  NOR2X0 U12116 ( .IN1(n10494), .IN2(n12087), .QN(n12085) );
  NAND2X0 U12117 ( .IN1(n12084), .IN2(g2571), .QN(n12087) );
  NAND2X0 U12118 ( .IN1(n12074), .IN2(n5521), .QN(n12084) );
  NAND2X0 U12119 ( .IN1(n12088), .IN2(n12089), .QN(g34015) );
  OR2X1 U12120 ( .IN1(n12090), .IN2(n12040), .Q(n12089) );
  NAND2X0 U12121 ( .IN1(n12091), .IN2(n10381), .QN(n12040) );
  NAND2X0 U12122 ( .IN1(n12092), .IN2(n12058), .QN(n12091) );
  NAND2X0 U12123 ( .IN1(n12093), .IN2(n12094), .QN(n12058) );
  NAND2X0 U12124 ( .IN1(n12095), .IN2(n12096), .QN(n12094) );
  NAND2X0 U12125 ( .IN1(n5757), .IN2(n12060), .QN(n12092) );
  NOR2X0 U12126 ( .IN1(n12097), .IN2(n12098), .QN(n12088) );
  NOR2X0 U12127 ( .IN1(n9622), .IN2(n10330), .QN(n12098) );
  NOR2X0 U12128 ( .IN1(n10494), .IN2(n12099), .QN(n12097) );
  NAND2X0 U12129 ( .IN1(n12090), .IN2(g2563), .QN(n12099) );
  NAND2X0 U12130 ( .IN1(n12067), .IN2(g2555), .QN(n12090) );
  NAND2X0 U12131 ( .IN1(n12100), .IN2(n12101), .QN(g34014) );
  NAND2X0 U12132 ( .IN1(n10511), .IN2(g2514), .QN(n12101) );
  NOR2X0 U12133 ( .IN1(n12102), .IN2(n12103), .QN(n12100) );
  NOR2X0 U12134 ( .IN1(n9624), .IN2(n12104), .QN(n12103) );
  NOR2X0 U12135 ( .IN1(n12105), .IN2(n12106), .QN(n12102) );
  NAND2X0 U12136 ( .IN1(n12107), .IN2(n12108), .QN(g34013) );
  NAND2X0 U12137 ( .IN1(n12109), .IN2(n12110), .QN(n12108) );
  NOR2X0 U12138 ( .IN1(n9692), .IN2(n12111), .QN(n12109) );
  NOR2X0 U12139 ( .IN1(n12112), .IN2(g2495), .QN(n12111) );
  NOR2X0 U12140 ( .IN1(n10494), .IN2(n10131), .QN(n12112) );
  NOR2X0 U12141 ( .IN1(n12113), .IN2(n12114), .QN(n12107) );
  NOR2X0 U12142 ( .IN1(n10494), .IN2(n12115), .QN(n12114) );
  NOR2X0 U12143 ( .IN1(n12116), .IN2(n12117), .QN(n12115) );
  NOR2X0 U12144 ( .IN1(n9692), .IN2(n12118), .QN(n12117) );
  NOR2X0 U12145 ( .IN1(n12110), .IN2(n12119), .QN(n12116) );
  NOR2X0 U12146 ( .IN1(n12120), .IN2(n12121), .QN(n12119) );
  NOR2X0 U12147 ( .IN1(n12122), .IN2(g2509), .QN(n12120) );
  AND2X1 U12148 ( .IN1(n12123), .IN2(n12124), .Q(n12110) );
  NAND2X0 U12149 ( .IN1(n12125), .IN2(g1589), .QN(n12124) );
  NOR2X0 U12150 ( .IN1(n5522), .IN2(n10330), .QN(n12113) );
  NAND2X0 U12151 ( .IN1(n12126), .IN2(n12127), .QN(g34012) );
  NAND2X0 U12152 ( .IN1(n12128), .IN2(n12129), .QN(n12127) );
  NOR2X0 U12153 ( .IN1(n12130), .IN2(n12131), .QN(n12126) );
  NOR2X0 U12154 ( .IN1(n5789), .IN2(n10330), .QN(n12131) );
  NOR2X0 U12155 ( .IN1(n10494), .IN2(n12132), .QN(n12130) );
  OR2X1 U12156 ( .IN1(n12128), .IN2(n5798), .Q(n12132) );
  NOR2X0 U12157 ( .IN1(n11754), .IN2(n12122), .QN(n12128) );
  NAND2X0 U12158 ( .IN1(n12133), .IN2(n12134), .QN(g34011) );
  NAND2X0 U12159 ( .IN1(n12135), .IN2(n12129), .QN(n12134) );
  NOR2X0 U12160 ( .IN1(n12136), .IN2(n12137), .QN(n12133) );
  NOR2X0 U12161 ( .IN1(n5798), .IN2(n10330), .QN(n12137) );
  NOR2X0 U12162 ( .IN1(n10495), .IN2(n12138), .QN(n12136) );
  OR2X1 U12163 ( .IN1(n12135), .IN2(n18477), .Q(n12138) );
  NOR2X0 U12164 ( .IN1(n12139), .IN2(test_so79), .QN(n12135) );
  NAND2X0 U12165 ( .IN1(n12140), .IN2(n12141), .QN(g34010) );
  OR2X1 U12166 ( .IN1(n12142), .IN2(n12105), .Q(n12141) );
  NOR2X0 U12167 ( .IN1(n12143), .IN2(n12144), .QN(n12140) );
  NOR2X0 U12168 ( .IN1(n18477), .IN2(n10330), .QN(n12144) );
  NOR2X0 U12169 ( .IN1(n10495), .IN2(n12145), .QN(n12143) );
  NAND2X0 U12170 ( .IN1(n12142), .IN2(g2441), .QN(n12145) );
  NAND2X0 U12171 ( .IN1(n12146), .IN2(g2495), .QN(n12142) );
  NAND2X0 U12172 ( .IN1(n12147), .IN2(n12148), .QN(g34009) );
  NAND2X0 U12173 ( .IN1(n12149), .IN2(n12129), .QN(n12148) );
  NOR2X0 U12174 ( .IN1(n12150), .IN2(n12151), .QN(n12147) );
  NOR2X0 U12175 ( .IN1(n5814), .IN2(n10331), .QN(n12151) );
  NOR2X0 U12176 ( .IN1(n10495), .IN2(n12152), .QN(n12150) );
  OR2X1 U12177 ( .IN1(n12149), .IN2(n5789), .Q(n12152) );
  NOR2X0 U12178 ( .IN1(n12139), .IN2(g2495), .QN(n12149) );
  NAND2X0 U12179 ( .IN1(n12153), .IN2(n12154), .QN(g34008) );
  NAND2X0 U12180 ( .IN1(n12155), .IN2(n12129), .QN(n12154) );
  INVX0 U12181 ( .INP(n12105), .ZN(n12129) );
  NAND2X0 U12182 ( .IN1(n12156), .IN2(n10380), .QN(n12105) );
  NAND2X0 U12183 ( .IN1(n12157), .IN2(n12123), .QN(n12156) );
  NAND2X0 U12184 ( .IN1(n12158), .IN2(n12159), .QN(n12123) );
  NAND2X0 U12185 ( .IN1(n12095), .IN2(n12160), .QN(n12159) );
  INVX0 U12186 ( .INP(n11031), .ZN(n12160) );
  NAND2X0 U12187 ( .IN1(n12125), .IN2(g1585), .QN(n12157) );
  NOR2X0 U12188 ( .IN1(n12161), .IN2(n12162), .QN(n12153) );
  NOR2X0 U12189 ( .IN1(n9624), .IN2(n10331), .QN(n12162) );
  NOR2X0 U12190 ( .IN1(n10495), .IN2(n12163), .QN(n12161) );
  OR2X1 U12191 ( .IN1(n12155), .IN2(n5814), .Q(n12163) );
  AND2X1 U12192 ( .IN1(n12146), .IN2(n5523), .Q(n12155) );
  NAND2X0 U12193 ( .IN1(n12164), .IN2(n12165), .QN(g34007) );
  NAND2X0 U12194 ( .IN1(n10511), .IN2(g2380), .QN(n12165) );
  NOR2X0 U12195 ( .IN1(n12166), .IN2(n12167), .QN(n12164) );
  NOR2X0 U12196 ( .IN1(n9644), .IN2(n12168), .QN(n12167) );
  NOR2X0 U12197 ( .IN1(n12169), .IN2(n12170), .QN(n12166) );
  NAND2X0 U12198 ( .IN1(n12171), .IN2(n12172), .QN(g34006) );
  NAND2X0 U12199 ( .IN1(n12173), .IN2(n12174), .QN(n12172) );
  NOR2X0 U12200 ( .IN1(n9694), .IN2(n12175), .QN(n12173) );
  NOR2X0 U12201 ( .IN1(n12176), .IN2(g2361), .QN(n12175) );
  NOR2X0 U12202 ( .IN1(n12177), .IN2(n12178), .QN(n12171) );
  NOR2X0 U12203 ( .IN1(n10496), .IN2(n12179), .QN(n12178) );
  NOR2X0 U12204 ( .IN1(n12180), .IN2(n12181), .QN(n12179) );
  AND2X1 U12205 ( .IN1(g2375), .IN2(n12182), .Q(n12181) );
  NOR2X0 U12206 ( .IN1(n12174), .IN2(n12183), .QN(n12180) );
  NOR2X0 U12207 ( .IN1(n12184), .IN2(n12185), .QN(n12183) );
  NOR2X0 U12208 ( .IN1(n12182), .IN2(g2375), .QN(n12184) );
  AND2X1 U12209 ( .IN1(n12186), .IN2(n12187), .Q(n12174) );
  NAND2X0 U12210 ( .IN1(n12188), .IN2(n5755), .QN(n12187) );
  NOR2X0 U12211 ( .IN1(n5537), .IN2(n10331), .QN(n12177) );
  NAND2X0 U12212 ( .IN1(n12189), .IN2(n12190), .QN(g34005) );
  OR2X1 U12213 ( .IN1(n12191), .IN2(n12169), .Q(n12190) );
  NOR2X0 U12214 ( .IN1(n12192), .IN2(n12193), .QN(n12189) );
  NOR2X0 U12215 ( .IN1(n5794), .IN2(n10331), .QN(n12193) );
  NOR2X0 U12216 ( .IN1(n10495), .IN2(n12194), .QN(n12192) );
  NAND2X0 U12217 ( .IN1(n12191), .IN2(g2315), .QN(n12194) );
  NAND2X0 U12218 ( .IN1(n12195), .IN2(n5513), .QN(n12191) );
  NAND2X0 U12219 ( .IN1(n12196), .IN2(n12197), .QN(g34004) );
  OR2X1 U12220 ( .IN1(n12198), .IN2(n12169), .Q(n12197) );
  NOR2X0 U12221 ( .IN1(n12199), .IN2(n12200), .QN(n12196) );
  NOR2X0 U12222 ( .IN1(n5802), .IN2(n10331), .QN(n12200) );
  NOR2X0 U12223 ( .IN1(n10496), .IN2(n12201), .QN(n12199) );
  NAND2X0 U12224 ( .IN1(n12198), .IN2(n9314), .QN(n12201) );
  NAND2X0 U12225 ( .IN1(n12202), .IN2(n5353), .QN(n12198) );
  NAND2X0 U12226 ( .IN1(n12203), .IN2(n12204), .QN(g34003) );
  OR2X1 U12227 ( .IN1(n12205), .IN2(n12169), .Q(n12204) );
  NOR2X0 U12228 ( .IN1(n12206), .IN2(n12207), .QN(n12203) );
  NOR2X0 U12229 ( .IN1(n18473), .IN2(n10331), .QN(n12207) );
  NOR2X0 U12230 ( .IN1(n10496), .IN2(n12208), .QN(n12206) );
  NAND2X0 U12231 ( .IN1(n12205), .IN2(g2307), .QN(n12208) );
  NAND2X0 U12232 ( .IN1(n12195), .IN2(g2287), .QN(n12205) );
  NOR2X0 U12233 ( .IN1(n5537), .IN2(n12182), .QN(n12195) );
  NAND2X0 U12234 ( .IN1(n12209), .IN2(n12210), .QN(g34002) );
  OR2X1 U12235 ( .IN1(n12211), .IN2(n12169), .Q(n12210) );
  NOR2X0 U12236 ( .IN1(n12212), .IN2(n12213), .QN(n12209) );
  NOR2X0 U12237 ( .IN1(n5815), .IN2(n10331), .QN(n12213) );
  NOR2X0 U12238 ( .IN1(n10496), .IN2(n12214), .QN(n12212) );
  NAND2X0 U12239 ( .IN1(n12211), .IN2(g2303), .QN(n12214) );
  NAND2X0 U12240 ( .IN1(n12202), .IN2(n5537), .QN(n12211) );
  NAND2X0 U12241 ( .IN1(n12215), .IN2(n12216), .QN(g34001) );
  OR2X1 U12242 ( .IN1(n12217), .IN2(n12169), .Q(n12216) );
  NAND2X0 U12243 ( .IN1(n12218), .IN2(n10380), .QN(n12169) );
  NAND2X0 U12244 ( .IN1(n12219), .IN2(n12186), .QN(n12218) );
  NAND2X0 U12245 ( .IN1(n12220), .IN2(n12221), .QN(n12186) );
  NAND2X0 U12246 ( .IN1(n12095), .IN2(n12222), .QN(n12221) );
  NAND2X0 U12247 ( .IN1(n12188), .IN2(n5757), .QN(n12219) );
  INVX0 U12248 ( .INP(n12220), .ZN(n12188) );
  NOR2X0 U12249 ( .IN1(n12223), .IN2(n12224), .QN(n12215) );
  NOR2X0 U12250 ( .IN1(n9644), .IN2(n10332), .QN(n12224) );
  NOR2X0 U12251 ( .IN1(n10494), .IN2(n12225), .QN(n12223) );
  NAND2X0 U12252 ( .IN1(n12217), .IN2(g2295), .QN(n12225) );
  NAND2X0 U12253 ( .IN1(n12226), .IN2(n5513), .QN(n12217) );
  NOR2X0 U12254 ( .IN1(n5353), .IN2(n12182), .QN(n12226) );
  NAND2X0 U12255 ( .IN1(n12227), .IN2(n12228), .QN(g34000) );
  NAND2X0 U12256 ( .IN1(n10511), .IN2(g2246), .QN(n12228) );
  NOR2X0 U12257 ( .IN1(n12229), .IN2(n12230), .QN(n12227) );
  NOR2X0 U12258 ( .IN1(n9652), .IN2(n12231), .QN(n12230) );
  NOR2X0 U12259 ( .IN1(n12232), .IN2(n12233), .QN(n12229) );
  NAND2X0 U12260 ( .IN1(n12234), .IN2(n12235), .QN(g33999) );
  NAND2X0 U12261 ( .IN1(n12236), .IN2(n12237), .QN(n12235) );
  NOR2X0 U12262 ( .IN1(n9696), .IN2(n12238), .QN(n12236) );
  NOR2X0 U12263 ( .IN1(n12239), .IN2(g2227), .QN(n12238) );
  NOR2X0 U12264 ( .IN1(n12240), .IN2(n12241), .QN(n12234) );
  NOR2X0 U12265 ( .IN1(n10495), .IN2(n12242), .QN(n12241) );
  NOR2X0 U12266 ( .IN1(n12243), .IN2(n12244), .QN(n12242) );
  AND2X1 U12267 ( .IN1(g2241), .IN2(n12245), .Q(n12244) );
  NOR2X0 U12268 ( .IN1(n12237), .IN2(n12246), .QN(n12243) );
  NOR2X0 U12269 ( .IN1(n12247), .IN2(n12248), .QN(n12246) );
  NOR2X0 U12270 ( .IN1(n12245), .IN2(g2241), .QN(n12247) );
  AND2X1 U12271 ( .IN1(n12249), .IN2(n12250), .Q(n12237) );
  NAND2X0 U12272 ( .IN1(n12251), .IN2(g1589), .QN(n12250) );
  NOR2X0 U12273 ( .IN1(n5538), .IN2(n10332), .QN(n12240) );
  NAND2X0 U12274 ( .IN1(n12252), .IN2(n12253), .QN(g33998) );
  OR2X1 U12275 ( .IN1(n12254), .IN2(n12232), .Q(n12253) );
  NOR2X0 U12276 ( .IN1(n12255), .IN2(n12256), .QN(n12252) );
  NOR2X0 U12277 ( .IN1(n5788), .IN2(n10332), .QN(n12256) );
  NOR2X0 U12278 ( .IN1(n10495), .IN2(n12257), .QN(n12255) );
  NAND2X0 U12279 ( .IN1(n12254), .IN2(g2181), .QN(n12257) );
  NAND2X0 U12280 ( .IN1(n12258), .IN2(n5514), .QN(n12254) );
  NAND2X0 U12281 ( .IN1(n12259), .IN2(n12260), .QN(g33997) );
  OR2X1 U12282 ( .IN1(n12261), .IN2(n12232), .Q(n12260) );
  NOR2X0 U12283 ( .IN1(n12262), .IN2(n12263), .QN(n12259) );
  NOR2X0 U12284 ( .IN1(n5803), .IN2(n10332), .QN(n12263) );
  NOR2X0 U12285 ( .IN1(n10496), .IN2(n12264), .QN(n12262) );
  NAND2X0 U12286 ( .IN1(n12261), .IN2(n9352), .QN(n12264) );
  NAND2X0 U12287 ( .IN1(n12265), .IN2(n5356), .QN(n12261) );
  NAND2X0 U12288 ( .IN1(n12266), .IN2(n12267), .QN(g33996) );
  OR2X1 U12289 ( .IN1(n12268), .IN2(n12232), .Q(n12267) );
  NOR2X0 U12290 ( .IN1(n12269), .IN2(n12270), .QN(n12266) );
  NOR2X0 U12291 ( .IN1(n18471), .IN2(n10332), .QN(n12270) );
  NOR2X0 U12292 ( .IN1(n10495), .IN2(n12271), .QN(n12269) );
  NAND2X0 U12293 ( .IN1(n12268), .IN2(g2173), .QN(n12271) );
  NAND2X0 U12294 ( .IN1(n12258), .IN2(g2153), .QN(n12268) );
  NOR2X0 U12295 ( .IN1(n5538), .IN2(n12245), .QN(n12258) );
  NAND2X0 U12296 ( .IN1(n12272), .IN2(n12273), .QN(g33995) );
  OR2X1 U12297 ( .IN1(n12274), .IN2(n12232), .Q(n12273) );
  NOR2X0 U12298 ( .IN1(n12275), .IN2(n12276), .QN(n12272) );
  NOR2X0 U12299 ( .IN1(n5812), .IN2(n10332), .QN(n12276) );
  NOR2X0 U12300 ( .IN1(n10495), .IN2(n12277), .QN(n12275) );
  NAND2X0 U12301 ( .IN1(n12274), .IN2(g2169), .QN(n12277) );
  NAND2X0 U12302 ( .IN1(n12265), .IN2(n5538), .QN(n12274) );
  NAND2X0 U12303 ( .IN1(n12278), .IN2(n12279), .QN(g33994) );
  OR2X1 U12304 ( .IN1(n12280), .IN2(n12232), .Q(n12279) );
  NAND2X0 U12305 ( .IN1(n12281), .IN2(n10380), .QN(n12232) );
  NAND2X0 U12306 ( .IN1(n12282), .IN2(n12249), .QN(n12281) );
  NAND2X0 U12307 ( .IN1(n12283), .IN2(n12284), .QN(n12249) );
  NAND2X0 U12308 ( .IN1(n12095), .IN2(n12285), .QN(n12284) );
  INVX0 U12309 ( .INP(n10956), .ZN(n12285) );
  NOR2X0 U12310 ( .IN1(n12286), .IN2(n5380), .QN(n12095) );
  NAND2X0 U12311 ( .IN1(n12251), .IN2(g1585), .QN(n12282) );
  INVX0 U12312 ( .INP(n12283), .ZN(n12251) );
  NOR2X0 U12313 ( .IN1(n12287), .IN2(n12288), .QN(n12278) );
  NOR2X0 U12314 ( .IN1(n9652), .IN2(n10332), .QN(n12288) );
  NOR2X0 U12315 ( .IN1(n10495), .IN2(n12289), .QN(n12287) );
  NAND2X0 U12316 ( .IN1(n12280), .IN2(g2161), .QN(n12289) );
  NAND2X0 U12317 ( .IN1(n12290), .IN2(n5514), .QN(n12280) );
  NOR2X0 U12318 ( .IN1(n5356), .IN2(n12245), .QN(n12290) );
  NAND2X0 U12319 ( .IN1(n12291), .IN2(n12292), .QN(g33993) );
  NAND2X0 U12320 ( .IN1(n10511), .IN2(g2089), .QN(n12292) );
  NOR2X0 U12321 ( .IN1(n12293), .IN2(n12294), .QN(n12291) );
  NOR2X0 U12322 ( .IN1(n9714), .IN2(n12295), .QN(n12294) );
  NOR2X0 U12323 ( .IN1(n12296), .IN2(n12297), .QN(n12293) );
  NAND2X0 U12324 ( .IN1(n12298), .IN2(n12299), .QN(g33992) );
  NAND2X0 U12325 ( .IN1(n12300), .IN2(n12301), .QN(n12299) );
  NOR2X0 U12326 ( .IN1(n9691), .IN2(n12302), .QN(n12300) );
  NOR2X0 U12327 ( .IN1(n12303), .IN2(g2070), .QN(n12302) );
  NOR2X0 U12328 ( .IN1(n5355), .IN2(n10460), .QN(n12303) );
  NOR2X0 U12329 ( .IN1(n12304), .IN2(n12305), .QN(n12298) );
  NOR2X0 U12330 ( .IN1(n10491), .IN2(n12306), .QN(n12305) );
  NOR2X0 U12331 ( .IN1(n12307), .IN2(n12308), .QN(n12306) );
  NOR2X0 U12332 ( .IN1(n9691), .IN2(n12309), .QN(n12308) );
  NOR2X0 U12333 ( .IN1(n12301), .IN2(n12310), .QN(n12307) );
  NOR2X0 U12334 ( .IN1(n12311), .IN2(n12312), .QN(n12310) );
  NOR2X0 U12335 ( .IN1(n12313), .IN2(g2084), .QN(n12311) );
  AND2X1 U12336 ( .IN1(n12314), .IN2(n12315), .Q(n12301) );
  NAND2X0 U12337 ( .IN1(n5756), .IN2(n12316), .QN(n12315) );
  NOR2X0 U12338 ( .IN1(n5535), .IN2(n10333), .QN(n12304) );
  NAND2X0 U12339 ( .IN1(n12317), .IN2(n12318), .QN(g33991) );
  NAND2X0 U12340 ( .IN1(n12319), .IN2(n12320), .QN(n12318) );
  NOR2X0 U12341 ( .IN1(n12321), .IN2(n12322), .QN(n12317) );
  NOR2X0 U12342 ( .IN1(n5790), .IN2(n10333), .QN(n12322) );
  NOR2X0 U12343 ( .IN1(n10491), .IN2(n12323), .QN(n12321) );
  OR2X1 U12344 ( .IN1(n12319), .IN2(n5801), .Q(n12323) );
  NOR2X0 U12345 ( .IN1(n12324), .IN2(n12313), .QN(n12319) );
  NAND2X0 U12346 ( .IN1(n12325), .IN2(n12326), .QN(g33990) );
  NAND2X0 U12347 ( .IN1(n12327), .IN2(n12320), .QN(n12326) );
  NOR2X0 U12348 ( .IN1(n12328), .IN2(n12329), .QN(n12325) );
  NOR2X0 U12349 ( .IN1(n5801), .IN2(n10333), .QN(n12329) );
  NOR2X0 U12350 ( .IN1(n10491), .IN2(n12330), .QN(n12328) );
  OR2X1 U12351 ( .IN1(n12327), .IN2(n18474), .Q(n12330) );
  NOR2X0 U12352 ( .IN1(n12331), .IN2(g1996), .QN(n12327) );
  NAND2X0 U12353 ( .IN1(n12332), .IN2(n12333), .QN(g33989) );
  OR2X1 U12354 ( .IN1(n12334), .IN2(n12296), .Q(n12333) );
  NOR2X0 U12355 ( .IN1(n12335), .IN2(n12336), .QN(n12332) );
  NOR2X0 U12356 ( .IN1(n18474), .IN2(n10333), .QN(n12336) );
  NOR2X0 U12357 ( .IN1(n10490), .IN2(n12337), .QN(n12335) );
  NAND2X0 U12358 ( .IN1(n12334), .IN2(g2016), .QN(n12337) );
  NAND2X0 U12359 ( .IN1(n12338), .IN2(g2070), .QN(n12334) );
  NAND2X0 U12360 ( .IN1(n12339), .IN2(n12340), .QN(g33988) );
  NAND2X0 U12361 ( .IN1(n12341), .IN2(n12320), .QN(n12340) );
  NOR2X0 U12362 ( .IN1(n12342), .IN2(n12343), .QN(n12339) );
  NOR2X0 U12363 ( .IN1(n5818), .IN2(n10333), .QN(n12343) );
  NOR2X0 U12364 ( .IN1(n10490), .IN2(n12344), .QN(n12342) );
  OR2X1 U12365 ( .IN1(n12341), .IN2(n5790), .Q(n12344) );
  NOR2X0 U12366 ( .IN1(n12331), .IN2(g2070), .QN(n12341) );
  NAND2X0 U12367 ( .IN1(n12345), .IN2(n12346), .QN(g33987) );
  NAND2X0 U12368 ( .IN1(n12347), .IN2(n12320), .QN(n12346) );
  INVX0 U12369 ( .INP(n12296), .ZN(n12320) );
  NAND2X0 U12370 ( .IN1(n12348), .IN2(n10379), .QN(n12296) );
  NAND2X0 U12371 ( .IN1(n12349), .IN2(n12314), .QN(n12348) );
  NAND2X0 U12372 ( .IN1(n12350), .IN2(n12351), .QN(n12314) );
  NAND2X0 U12373 ( .IN1(n12352), .IN2(n12353), .QN(n12351) );
  NAND2X0 U12374 ( .IN1(n5526), .IN2(n12316), .QN(n12349) );
  NOR2X0 U12375 ( .IN1(n12354), .IN2(n12355), .QN(n12345) );
  NOR2X0 U12376 ( .IN1(n9714), .IN2(n10333), .QN(n12355) );
  NOR2X0 U12377 ( .IN1(n10490), .IN2(n12356), .QN(n12354) );
  OR2X1 U12378 ( .IN1(n12347), .IN2(n5818), .Q(n12356) );
  AND2X1 U12379 ( .IN1(n12338), .IN2(n5505), .Q(n12347) );
  NAND2X0 U12380 ( .IN1(n12357), .IN2(n12358), .QN(g33986) );
  NAND2X0 U12381 ( .IN1(n10512), .IN2(g1955), .QN(n12358) );
  NOR2X0 U12382 ( .IN1(n12359), .IN2(n12360), .QN(n12357) );
  NOR2X0 U12383 ( .IN1(n9633), .IN2(n12361), .QN(n12360) );
  NOR2X0 U12384 ( .IN1(n12362), .IN2(n12363), .QN(n12359) );
  NAND2X0 U12385 ( .IN1(n12364), .IN2(n12365), .QN(g33985) );
  NAND2X0 U12386 ( .IN1(n12366), .IN2(n12367), .QN(n12365) );
  NOR2X0 U12387 ( .IN1(n9695), .IN2(n12368), .QN(n12366) );
  NOR2X0 U12388 ( .IN1(n12369), .IN2(g1936), .QN(n12368) );
  NOR2X0 U12389 ( .IN1(n10489), .IN2(n10137), .QN(n12369) );
  NOR2X0 U12390 ( .IN1(n12370), .IN2(n12371), .QN(n12364) );
  NOR2X0 U12391 ( .IN1(n10489), .IN2(n12372), .QN(n12371) );
  NOR2X0 U12392 ( .IN1(n12373), .IN2(n12374), .QN(n12372) );
  NOR2X0 U12393 ( .IN1(n9695), .IN2(n12375), .QN(n12374) );
  NOR2X0 U12394 ( .IN1(n12367), .IN2(n12376), .QN(n12373) );
  NOR2X0 U12395 ( .IN1(n12377), .IN2(n12378), .QN(n12376) );
  NOR2X0 U12396 ( .IN1(n12379), .IN2(g1950), .QN(n12377) );
  AND2X1 U12397 ( .IN1(n12380), .IN2(n12381), .Q(n12367) );
  NAND2X0 U12398 ( .IN1(n12382), .IN2(g1246), .QN(n12381) );
  NOR2X0 U12399 ( .IN1(n5534), .IN2(n10333), .QN(n12370) );
  NAND2X0 U12400 ( .IN1(n12383), .IN2(n12384), .QN(g33984) );
  NAND2X0 U12401 ( .IN1(n12385), .IN2(n12386), .QN(n12384) );
  NOR2X0 U12402 ( .IN1(n12387), .IN2(n12388), .QN(n12383) );
  NOR2X0 U12403 ( .IN1(n5793), .IN2(n10334), .QN(n12388) );
  NOR2X0 U12404 ( .IN1(n10489), .IN2(n12389), .QN(n12387) );
  OR2X1 U12405 ( .IN1(n12385), .IN2(n5799), .Q(n12389) );
  NOR2X0 U12406 ( .IN1(n12390), .IN2(n12379), .QN(n12385) );
  NAND2X0 U12407 ( .IN1(n12391), .IN2(n12392), .QN(g33983) );
  NAND2X0 U12408 ( .IN1(n12393), .IN2(n12386), .QN(n12392) );
  NOR2X0 U12409 ( .IN1(n12394), .IN2(n12395), .QN(n12391) );
  NOR2X0 U12410 ( .IN1(n5799), .IN2(n10334), .QN(n12395) );
  NOR2X0 U12411 ( .IN1(n10488), .IN2(n12396), .QN(n12394) );
  OR2X1 U12412 ( .IN1(n12393), .IN2(n18476), .Q(n12396) );
  NOR2X0 U12413 ( .IN1(n12397), .IN2(test_so8), .QN(n12393) );
  NAND2X0 U12414 ( .IN1(n12398), .IN2(n12399), .QN(g33982) );
  OR2X1 U12415 ( .IN1(n12400), .IN2(n12362), .Q(n12399) );
  NOR2X0 U12416 ( .IN1(n12401), .IN2(n12402), .QN(n12398) );
  NOR2X0 U12417 ( .IN1(n18476), .IN2(n10334), .QN(n12402) );
  NOR2X0 U12418 ( .IN1(n10488), .IN2(n12403), .QN(n12401) );
  NAND2X0 U12419 ( .IN1(n12400), .IN2(g1882), .QN(n12403) );
  NAND2X0 U12420 ( .IN1(n12404), .IN2(g1936), .QN(n12400) );
  NAND2X0 U12421 ( .IN1(n12405), .IN2(n12406), .QN(g33981) );
  NAND2X0 U12422 ( .IN1(n12407), .IN2(n12386), .QN(n12406) );
  NOR2X0 U12423 ( .IN1(n12408), .IN2(n12409), .QN(n12405) );
  NOR2X0 U12424 ( .IN1(n5813), .IN2(n10334), .QN(n12409) );
  NOR2X0 U12425 ( .IN1(n10488), .IN2(n12410), .QN(n12408) );
  OR2X1 U12426 ( .IN1(n12407), .IN2(n5793), .Q(n12410) );
  NOR2X0 U12427 ( .IN1(n12397), .IN2(g1936), .QN(n12407) );
  NAND2X0 U12428 ( .IN1(n12411), .IN2(n12412), .QN(g33980) );
  NAND2X0 U12429 ( .IN1(n12413), .IN2(n12386), .QN(n12412) );
  INVX0 U12430 ( .INP(n12362), .ZN(n12386) );
  NAND2X0 U12431 ( .IN1(n12414), .IN2(n10379), .QN(n12362) );
  NAND2X0 U12432 ( .IN1(n12415), .IN2(n12380), .QN(n12414) );
  NAND2X0 U12433 ( .IN1(n12416), .IN2(n12417), .QN(n12380) );
  NAND2X0 U12434 ( .IN1(n12352), .IN2(n12418), .QN(n12417) );
  NAND2X0 U12435 ( .IN1(n12382), .IN2(g30332), .QN(n12415) );
  NOR2X0 U12436 ( .IN1(n12419), .IN2(n12420), .QN(n12411) );
  NOR2X0 U12437 ( .IN1(n9633), .IN2(n10334), .QN(n12420) );
  NOR2X0 U12438 ( .IN1(n10487), .IN2(n12421), .QN(n12419) );
  OR2X1 U12439 ( .IN1(n12413), .IN2(n5813), .Q(n12421) );
  AND2X1 U12440 ( .IN1(n12404), .IN2(n5503), .Q(n12413) );
  NAND2X0 U12441 ( .IN1(n12422), .IN2(n12423), .QN(g33979) );
  NAND2X0 U12442 ( .IN1(n10512), .IN2(g1821), .QN(n12423) );
  NOR2X0 U12443 ( .IN1(n12424), .IN2(n12425), .QN(n12422) );
  NOR2X0 U12444 ( .IN1(n9704), .IN2(n12426), .QN(n12425) );
  NOR2X0 U12445 ( .IN1(n12427), .IN2(n12428), .QN(n12424) );
  NAND2X0 U12446 ( .IN1(n12429), .IN2(n12430), .QN(g33978) );
  NAND2X0 U12447 ( .IN1(n12431), .IN2(n12432), .QN(n12430) );
  NOR2X0 U12448 ( .IN1(n9615), .IN2(n12433), .QN(n12431) );
  NOR2X0 U12449 ( .IN1(n12434), .IN2(g1802), .QN(n12433) );
  NOR2X0 U12450 ( .IN1(n12435), .IN2(n12436), .QN(n12429) );
  NOR2X0 U12451 ( .IN1(n10487), .IN2(n12437), .QN(n12436) );
  NOR2X0 U12452 ( .IN1(n12438), .IN2(n12439), .QN(n12437) );
  NOR2X0 U12453 ( .IN1(n9615), .IN2(n12440), .QN(n12439) );
  NOR2X0 U12454 ( .IN1(n12432), .IN2(n12441), .QN(n12438) );
  NOR2X0 U12455 ( .IN1(n12442), .IN2(n12443), .QN(n12441) );
  NOR2X0 U12456 ( .IN1(n12444), .IN2(g1816), .QN(n12442) );
  AND2X1 U12457 ( .IN1(n12445), .IN2(n12446), .Q(n12432) );
  NAND2X0 U12458 ( .IN1(n12447), .IN2(n5756), .QN(n12446) );
  NOR2X0 U12459 ( .IN1(n5536), .IN2(n10334), .QN(n12435) );
  NAND2X0 U12460 ( .IN1(n12448), .IN2(n12449), .QN(g33977) );
  OR2X1 U12461 ( .IN1(n12450), .IN2(n12427), .Q(n12449) );
  NOR2X0 U12462 ( .IN1(n12451), .IN2(n12452), .QN(n12448) );
  NOR2X0 U12463 ( .IN1(n5795), .IN2(n10334), .QN(n12452) );
  NOR2X0 U12464 ( .IN1(n10487), .IN2(n12453), .QN(n12451) );
  NAND2X0 U12465 ( .IN1(n12450), .IN2(g1756), .QN(n12453) );
  NAND2X0 U12466 ( .IN1(n12454), .IN2(n5504), .QN(n12450) );
  NAND2X0 U12467 ( .IN1(n12455), .IN2(n12456), .QN(g33976) );
  OR2X1 U12468 ( .IN1(n12457), .IN2(n12427), .Q(n12456) );
  NOR2X0 U12469 ( .IN1(n12458), .IN2(n12459), .QN(n12455) );
  NOR2X0 U12470 ( .IN1(n5804), .IN2(n10335), .QN(n12459) );
  NOR2X0 U12471 ( .IN1(n10486), .IN2(n12460), .QN(n12458) );
  NAND2X0 U12472 ( .IN1(n12457), .IN2(g1752), .QN(n12460) );
  NAND2X0 U12473 ( .IN1(n12461), .IN2(n5352), .QN(n12457) );
  NAND2X0 U12474 ( .IN1(n12462), .IN2(n12463), .QN(g33975) );
  OR2X1 U12475 ( .IN1(n12464), .IN2(n12427), .Q(n12463) );
  NOR2X0 U12476 ( .IN1(n12465), .IN2(n12466), .QN(n12462) );
  NOR2X0 U12477 ( .IN1(n5797), .IN2(n10335), .QN(n12466) );
  NOR2X0 U12478 ( .IN1(n10486), .IN2(n12467), .QN(n12465) );
  NAND2X0 U12479 ( .IN1(n12464), .IN2(g1748), .QN(n12467) );
  NAND2X0 U12480 ( .IN1(n12454), .IN2(g1728), .QN(n12464) );
  NOR2X0 U12481 ( .IN1(n5536), .IN2(n12444), .QN(n12454) );
  NAND2X0 U12482 ( .IN1(n12468), .IN2(n12469), .QN(g33974) );
  OR2X1 U12483 ( .IN1(n12470), .IN2(n12427), .Q(n12469) );
  NOR2X0 U12484 ( .IN1(n12471), .IN2(n12472), .QN(n12468) );
  NOR2X0 U12485 ( .IN1(n5817), .IN2(n10335), .QN(n12472) );
  NOR2X0 U12486 ( .IN1(n10486), .IN2(n12473), .QN(n12471) );
  NAND2X0 U12487 ( .IN1(n12470), .IN2(g1744), .QN(n12473) );
  NAND2X0 U12488 ( .IN1(n12461), .IN2(n5536), .QN(n12470) );
  NAND2X0 U12489 ( .IN1(n12474), .IN2(n12475), .QN(g33973) );
  OR2X1 U12490 ( .IN1(n12476), .IN2(n12427), .Q(n12475) );
  NAND2X0 U12491 ( .IN1(n12477), .IN2(n10397), .QN(n12427) );
  NAND2X0 U12492 ( .IN1(n12478), .IN2(n12445), .QN(n12477) );
  NAND2X0 U12493 ( .IN1(n12479), .IN2(n12480), .QN(n12445) );
  NAND2X0 U12494 ( .IN1(n12352), .IN2(n12481), .QN(n12480) );
  INVX0 U12495 ( .INP(n10996), .ZN(n12481) );
  NAND2X0 U12496 ( .IN1(n12447), .IN2(n5526), .QN(n12478) );
  NOR2X0 U12497 ( .IN1(n12482), .IN2(n12483), .QN(n12474) );
  NOR2X0 U12498 ( .IN1(n9704), .IN2(n10335), .QN(n12483) );
  NOR2X0 U12499 ( .IN1(n10486), .IN2(n12484), .QN(n12482) );
  NAND2X0 U12500 ( .IN1(n12476), .IN2(g1736), .QN(n12484) );
  NAND2X0 U12501 ( .IN1(n12485), .IN2(n5504), .QN(n12476) );
  NOR2X0 U12502 ( .IN1(n5352), .IN2(n12444), .QN(n12485) );
  NAND2X0 U12503 ( .IN1(n12486), .IN2(n12487), .QN(g33972) );
  NAND2X0 U12504 ( .IN1(n10512), .IN2(g1687), .QN(n12487) );
  NOR2X0 U12505 ( .IN1(n12488), .IN2(n12489), .QN(n12486) );
  NOR2X0 U12506 ( .IN1(n9623), .IN2(n12490), .QN(n12489) );
  NOR2X0 U12507 ( .IN1(n12491), .IN2(n12492), .QN(n12488) );
  NAND2X0 U12508 ( .IN1(n12493), .IN2(n12494), .QN(g33971) );
  NAND2X0 U12509 ( .IN1(n12495), .IN2(n12496), .QN(n12494) );
  NOR2X0 U12510 ( .IN1(n9697), .IN2(n12497), .QN(n12495) );
  NOR2X0 U12511 ( .IN1(n12498), .IN2(g1668), .QN(n12497) );
  NOR2X0 U12512 ( .IN1(n5362), .IN2(n10461), .QN(n12498) );
  NOR2X0 U12513 ( .IN1(n12499), .IN2(n12500), .QN(n12493) );
  NOR2X0 U12514 ( .IN1(n10486), .IN2(n12501), .QN(n12500) );
  NOR2X0 U12515 ( .IN1(n12502), .IN2(n12503), .QN(n12501) );
  NOR2X0 U12516 ( .IN1(n9697), .IN2(n12504), .QN(n12503) );
  NOR2X0 U12517 ( .IN1(n12496), .IN2(n12505), .QN(n12502) );
  NOR2X0 U12518 ( .IN1(n12506), .IN2(n12507), .QN(n12505) );
  NOR2X0 U12519 ( .IN1(n12508), .IN2(g1682), .QN(n12506) );
  AND2X1 U12520 ( .IN1(n12509), .IN2(n12510), .Q(n12496) );
  NAND2X0 U12521 ( .IN1(n12511), .IN2(g1246), .QN(n12510) );
  NOR2X0 U12522 ( .IN1(n5598), .IN2(n10335), .QN(n12499) );
  NAND2X0 U12523 ( .IN1(n12512), .IN2(n12513), .QN(g33970) );
  OR2X1 U12524 ( .IN1(n12514), .IN2(n12491), .Q(n12513) );
  NOR2X0 U12525 ( .IN1(n12515), .IN2(n12516), .QN(n12512) );
  NOR2X0 U12526 ( .IN1(n5792), .IN2(n10335), .QN(n12516) );
  NOR2X0 U12527 ( .IN1(n10486), .IN2(n12517), .QN(n12515) );
  NAND2X0 U12528 ( .IN1(n12514), .IN2(g1620), .QN(n12517) );
  NAND2X0 U12529 ( .IN1(g31862), .IN2(n12504), .QN(n12514) );
  NAND2X0 U12530 ( .IN1(n12518), .IN2(n12519), .QN(g33969) );
  NAND2X0 U12531 ( .IN1(n12520), .IN2(n12521), .QN(n12519) );
  NOR2X0 U12532 ( .IN1(n12522), .IN2(n12523), .QN(n12518) );
  NOR2X0 U12533 ( .IN1(n5791), .IN2(n10335), .QN(n12523) );
  NOR2X0 U12534 ( .IN1(n10486), .IN2(n12524), .QN(n12522) );
  OR2X1 U12535 ( .IN1(n12520), .IN2(n18475), .Q(n12524) );
  NOR2X0 U12536 ( .IN1(n12525), .IN2(g1592), .QN(n12520) );
  NAND2X0 U12537 ( .IN1(n12526), .IN2(n12527), .QN(g33968) );
  OR2X1 U12538 ( .IN1(n12528), .IN2(n12491), .Q(n12527) );
  NOR2X0 U12539 ( .IN1(n12529), .IN2(n12530), .QN(n12526) );
  NOR2X0 U12540 ( .IN1(n18475), .IN2(n10336), .QN(n12530) );
  NOR2X0 U12541 ( .IN1(n10486), .IN2(n12531), .QN(n12529) );
  NAND2X0 U12542 ( .IN1(n12528), .IN2(g1612), .QN(n12531) );
  NAND2X0 U12543 ( .IN1(n12532), .IN2(g1668), .QN(n12528) );
  NAND2X0 U12544 ( .IN1(n12533), .IN2(n12534), .QN(g33967) );
  NAND2X0 U12545 ( .IN1(n12535), .IN2(n12521), .QN(n12534) );
  INVX0 U12546 ( .INP(n12491), .ZN(n12521) );
  NOR2X0 U12547 ( .IN1(n12536), .IN2(n12537), .QN(n12533) );
  NOR2X0 U12548 ( .IN1(n5811), .IN2(n10336), .QN(n12537) );
  NOR2X0 U12549 ( .IN1(n10486), .IN2(n12538), .QN(n12536) );
  OR2X1 U12550 ( .IN1(n12535), .IN2(n5792), .Q(n12538) );
  NOR2X0 U12551 ( .IN1(n12525), .IN2(g1668), .QN(n12535) );
  NAND2X0 U12552 ( .IN1(n12539), .IN2(n12540), .QN(g33966) );
  OR2X1 U12553 ( .IN1(n12541), .IN2(n12491), .Q(n12540) );
  NAND2X0 U12554 ( .IN1(n12542), .IN2(n10397), .QN(n12491) );
  NAND2X0 U12555 ( .IN1(n12543), .IN2(n12509), .QN(n12542) );
  NAND2X0 U12556 ( .IN1(n12544), .IN2(n12545), .QN(n12509) );
  NAND2X0 U12557 ( .IN1(n12352), .IN2(n12546), .QN(n12545) );
  NOR2X0 U12558 ( .IN1(n12547), .IN2(n5380), .QN(n12352) );
  NAND2X0 U12559 ( .IN1(n12511), .IN2(g30332), .QN(n12543) );
  INVX0 U12560 ( .INP(n12544), .ZN(n12511) );
  NOR2X0 U12561 ( .IN1(n12548), .IN2(n12549), .QN(n12539) );
  NOR2X0 U12562 ( .IN1(n9623), .IN2(n10336), .QN(n12549) );
  NOR2X0 U12563 ( .IN1(n10486), .IN2(n12550), .QN(n12548) );
  NAND2X0 U12564 ( .IN1(n12541), .IN2(g1600), .QN(n12550) );
  NAND2X0 U12565 ( .IN1(n12532), .IN2(n5549), .QN(n12541) );
  NAND2X0 U12566 ( .IN1(n12551), .IN2(n12552), .QN(g33965) );
  NAND2X0 U12567 ( .IN1(n10513), .IN2(g763), .QN(n12552) );
  NOR2X0 U12568 ( .IN1(n12553), .IN2(n12554), .QN(n12551) );
  NOR2X0 U12569 ( .IN1(g767), .IN2(n12555), .QN(n12554) );
  NOR2X0 U12570 ( .IN1(n5333), .IN2(n12556), .QN(n12553) );
  NAND2X0 U12571 ( .IN1(n2404), .IN2(n12555), .QN(n12556) );
  INVX0 U12572 ( .INP(n2704), .ZN(n12555) );
  NAND2X0 U12573 ( .IN1(n12557), .IN2(n12558), .QN(g33964) );
  NAND2X0 U12574 ( .IN1(n10513), .IN2(g595), .QN(n12558) );
  NOR2X0 U12575 ( .IN1(n12559), .IN2(n12560), .QN(n12557) );
  NOR2X0 U12576 ( .IN1(g599), .IN2(n12561), .QN(n12560) );
  NOR2X0 U12577 ( .IN1(n5550), .IN2(n12562), .QN(n12559) );
  NAND2X0 U12578 ( .IN1(n2421), .IN2(n12561), .QN(n12562) );
  INVX0 U12579 ( .INP(n2706), .ZN(n12561) );
  NAND2X0 U12580 ( .IN1(n12563), .IN2(n12564), .QN(g33963) );
  NAND2X0 U12581 ( .IN1(n10513), .IN2(g29215), .QN(n12564) );
  NAND2X0 U12582 ( .IN1(n12565), .IN2(n10397), .QN(n12563) );
  NOR2X0 U12583 ( .IN1(n12566), .IN2(n12567), .QN(n12565) );
  NOR2X0 U12584 ( .IN1(n12568), .IN2(n12569), .QN(n12567) );
  NOR2X0 U12585 ( .IN1(n9781), .IN2(g72), .QN(n12568) );
  NOR2X0 U12586 ( .IN1(n12570), .IN2(n12571), .QN(n12566) );
  NAND2X0 U12587 ( .IN1(n12572), .IN2(n10784), .QN(n12571) );
  NAND2X0 U12588 ( .IN1(n12573), .IN2(g269), .QN(n12572) );
  NOR2X0 U12589 ( .IN1(n9782), .IN2(n10783), .QN(n12570) );
  NAND2X0 U12590 ( .IN1(n12574), .IN2(n12575), .QN(g33962) );
  NAND2X0 U12591 ( .IN1(n10513), .IN2(g479), .QN(n12575) );
  NAND2X0 U12592 ( .IN1(n12576), .IN2(n10397), .QN(n12574) );
  NOR2X0 U12593 ( .IN1(n12577), .IN2(n12578), .QN(n12576) );
  NAND2X0 U12594 ( .IN1(n12579), .IN2(n12580), .QN(n12578) );
  NAND2X0 U12595 ( .IN1(n12581), .IN2(g73), .QN(n12580) );
  NOR2X0 U12596 ( .IN1(g225), .IN2(n12573), .QN(n12581) );
  NAND2X0 U12597 ( .IN1(n12582), .IN2(n10783), .QN(n12579) );
  NAND2X0 U12598 ( .IN1(n12583), .IN2(n12584), .QN(n12582) );
  NAND2X0 U12599 ( .IN1(g73), .IN2(n9908), .QN(n12584) );
  NOR2X0 U12600 ( .IN1(g239), .IN2(n12583), .QN(n12577) );
  NAND2X0 U12601 ( .IN1(n10784), .IN2(n12585), .QN(n12583) );
  NAND2X0 U12602 ( .IN1(n12573), .IN2(g246), .QN(n12585) );
  INVX0 U12603 ( .INP(g73), .ZN(n10784) );
  NAND2X0 U12604 ( .IN1(n12586), .IN2(n12587), .QN(g33961) );
  NAND2X0 U12605 ( .IN1(n10513), .IN2(g294), .QN(n12587) );
  NOR2X0 U12606 ( .IN1(n12588), .IN2(n12589), .QN(n12586) );
  NOR2X0 U12607 ( .IN1(g298), .IN2(n12590), .QN(n12589) );
  NOR2X0 U12608 ( .IN1(n5675), .IN2(n12591), .QN(n12588) );
  NAND2X0 U12609 ( .IN1(n10106), .IN2(n12590), .QN(n12591) );
  INVX0 U12610 ( .INP(n2989), .ZN(n12590) );
  NAND2X0 U12611 ( .IN1(n12592), .IN2(n12593), .QN(g33960) );
  NAND2X0 U12612 ( .IN1(n10513), .IN2(g153), .QN(n12593) );
  NOR2X0 U12613 ( .IN1(n12594), .IN2(n12595), .QN(n12592) );
  NOR2X0 U12614 ( .IN1(g157), .IN2(n12596), .QN(n12595) );
  NOR2X0 U12615 ( .IN1(n5678), .IN2(n12597), .QN(n12594) );
  NAND2X0 U12616 ( .IN1(n11894), .IN2(n12596), .QN(n12597) );
  INVX0 U12617 ( .INP(n2991), .ZN(n12596) );
  NAND2X0 U12618 ( .IN1(n12598), .IN2(n12599), .QN(g33935) );
  NOR2X0 U12619 ( .IN1(n9717), .IN2(n9716), .QN(n12599) );
  NOR2X0 U12620 ( .IN1(g34649), .IN2(n11790), .QN(n12598) );
  NAND2X0 U12621 ( .IN1(n12600), .IN2(n12601), .QN(g34649) );
  NOR2X0 U12622 ( .IN1(n12602), .IN2(n12603), .QN(n12601) );
  NOR2X0 U12623 ( .IN1(n12604), .IN2(n12605), .QN(n12600) );
  NAND2X0 U12624 ( .IN1(n12606), .IN2(n5541), .QN(g33874) );
  NOR2X0 U12625 ( .IN1(n5846), .IN2(n11790), .QN(n12606) );
  NAND2X0 U12626 ( .IN1(n12607), .IN2(n12608), .QN(g33659) );
  AND2X1 U12627 ( .IN1(n10796), .IN2(n10795), .Q(n12608) );
  XOR2X1 U12628 ( .IN1(n9913), .IN2(g73), .Q(n10795) );
  XOR2X1 U12629 ( .IN1(g4108), .IN2(n10783), .Q(n10796) );
  INVX0 U12630 ( .INP(g72), .ZN(n10783) );
  AND2X1 U12631 ( .IN1(n11716), .IN2(n10794), .Q(n12607) );
  AND2X1 U12632 ( .IN1(n12609), .IN2(n12610), .Q(n10794) );
  NAND2X0 U12633 ( .IN1(n5350), .IN2(n12611), .QN(n12610) );
  NAND2X0 U12634 ( .IN1(n12612), .IN2(n12613), .QN(n12611) );
  NAND2X0 U12635 ( .IN1(n12614), .IN2(n12615), .QN(n12613) );
  NOR2X0 U12636 ( .IN1(n12616), .IN2(n12617), .QN(n12612) );
  NOR2X0 U12637 ( .IN1(n12618), .IN2(n12619), .QN(n12617) );
  NOR2X0 U12638 ( .IN1(n5340), .IN2(n12620), .QN(n12616) );
  NAND2X0 U12639 ( .IN1(n12621), .IN2(n12622), .QN(n12620) );
  NAND2X0 U12640 ( .IN1(n5480), .IN2(n12623), .QN(n12622) );
  NAND2X0 U12641 ( .IN1(n12624), .IN2(g4087), .QN(n12621) );
  NAND2X0 U12642 ( .IN1(n12625), .IN2(g4098), .QN(n12609) );
  NAND2X0 U12643 ( .IN1(n12626), .IN2(n12627), .QN(n12625) );
  NAND2X0 U12644 ( .IN1(n12615), .IN2(n12628), .QN(n12627) );
  NOR2X0 U12645 ( .IN1(n12629), .IN2(n12630), .QN(n12626) );
  NOR2X0 U12646 ( .IN1(n12618), .IN2(n12631), .QN(n12630) );
  NOR2X0 U12647 ( .IN1(n5340), .IN2(n12632), .QN(n12629) );
  NAND2X0 U12648 ( .IN1(n12633), .IN2(n12634), .QN(n12632) );
  NAND2X0 U12649 ( .IN1(n5480), .IN2(n12635), .QN(n12634) );
  NAND2X0 U12650 ( .IN1(n12636), .IN2(g4087), .QN(n12633) );
  AND2X1 U12651 ( .IN1(g113), .IN2(n2668), .Q(n11716) );
  NAND2X0 U12652 ( .IN1(n12637), .IN2(n12638), .QN(g33636) );
  NOR2X0 U12653 ( .IN1(n9719), .IN2(n9718), .QN(n12638) );
  NOR2X0 U12654 ( .IN1(g34657), .IN2(n11790), .QN(n12637) );
  INVX0 U12655 ( .INP(n2668), .ZN(n11790) );
  NAND2X0 U12656 ( .IN1(n12639), .IN2(n12640), .QN(n2668) );
  NAND2X0 U12657 ( .IN1(g99), .IN2(g37), .QN(n12640) );
  NAND2X0 U12658 ( .IN1(n12641), .IN2(n12642), .QN(g34657) );
  NOR2X0 U12659 ( .IN1(n12643), .IN2(n12644), .QN(n12642) );
  NOR2X0 U12660 ( .IN1(n12645), .IN2(n12646), .QN(n12641) );
  NAND2X0 U12661 ( .IN1(n12647), .IN2(n12648), .QN(g33627) );
  NAND2X0 U12662 ( .IN1(n12649), .IN2(n12650), .QN(n12648) );
  NAND2X0 U12663 ( .IN1(n12651), .IN2(n12652), .QN(n12649) );
  NAND2X0 U12664 ( .IN1(n12653), .IN2(n10398), .QN(n12652) );
  NAND2X0 U12665 ( .IN1(n10672), .IN2(n12654), .QN(n12653) );
  NAND2X0 U12666 ( .IN1(n10113), .IN2(g6682), .QN(n12654) );
  NAND2X0 U12667 ( .IN1(n10675), .IN2(n12655), .QN(n12651) );
  NAND2X0 U12668 ( .IN1(n10513), .IN2(g6741), .QN(n12647) );
  NAND2X0 U12669 ( .IN1(n12656), .IN2(n12657), .QN(g33626) );
  NAND2X0 U12670 ( .IN1(n12658), .IN2(g6741), .QN(n12657) );
  NOR2X0 U12671 ( .IN1(n12659), .IN2(n12660), .QN(n12656) );
  NOR2X0 U12672 ( .IN1(n10036), .IN2(n10336), .QN(n12660) );
  NOR2X0 U12673 ( .IN1(n10485), .IN2(n12661), .QN(n12659) );
  NAND2X0 U12674 ( .IN1(n12662), .IN2(n5398), .QN(n12661) );
  AND2X1 U12675 ( .IN1(n12655), .IN2(n12650), .Q(n12662) );
  NAND2X0 U12676 ( .IN1(n12663), .IN2(n3023), .QN(n12650) );
  NOR2X0 U12677 ( .IN1(n10113), .IN2(n11697), .QN(n12663) );
  NAND2X0 U12678 ( .IN1(n12664), .IN2(n12665), .QN(g33625) );
  NAND2X0 U12679 ( .IN1(n12666), .IN2(n12667), .QN(n12665) );
  NAND2X0 U12680 ( .IN1(n12668), .IN2(n12669), .QN(n12666) );
  NAND2X0 U12681 ( .IN1(n12670), .IN2(n10398), .QN(n12669) );
  NAND2X0 U12682 ( .IN1(n12671), .IN2(n12672), .QN(n12670) );
  NAND2X0 U12683 ( .IN1(n12673), .IN2(g6336), .QN(n12672) );
  NAND2X0 U12684 ( .IN1(n12674), .IN2(n12675), .QN(n12668) );
  NAND2X0 U12685 ( .IN1(n10514), .IN2(g6395), .QN(n12664) );
  NAND2X0 U12686 ( .IN1(n12676), .IN2(n12677), .QN(g33624) );
  NAND2X0 U12687 ( .IN1(n12678), .IN2(g6395), .QN(n12677) );
  NOR2X0 U12688 ( .IN1(n12679), .IN2(n12680), .QN(n12676) );
  NOR2X0 U12689 ( .IN1(n9898), .IN2(n10336), .QN(n12680) );
  NOR2X0 U12690 ( .IN1(n10485), .IN2(n12681), .QN(n12679) );
  NAND2X0 U12691 ( .IN1(n12682), .IN2(n5396), .QN(n12681) );
  AND2X1 U12692 ( .IN1(n12667), .IN2(n12675), .Q(n12682) );
  NAND2X0 U12693 ( .IN1(n12683), .IN2(n3033), .QN(n12667) );
  NOR2X0 U12694 ( .IN1(n11703), .IN2(n12673), .QN(n12683) );
  NAND2X0 U12695 ( .IN1(n12684), .IN2(n12685), .QN(g33623) );
  NAND2X0 U12696 ( .IN1(n12686), .IN2(n12687), .QN(n12685) );
  NAND2X0 U12697 ( .IN1(n12688), .IN2(n12689), .QN(n12686) );
  NAND2X0 U12698 ( .IN1(n12690), .IN2(n10398), .QN(n12689) );
  NAND2X0 U12699 ( .IN1(n12691), .IN2(n12692), .QN(n12690) );
  NAND2X0 U12700 ( .IN1(n12693), .IN2(g5990), .QN(n12692) );
  NAND2X0 U12701 ( .IN1(n12694), .IN2(n12695), .QN(n12688) );
  NAND2X0 U12702 ( .IN1(test_so57), .IN2(n10515), .QN(n12684) );
  NAND2X0 U12703 ( .IN1(n12696), .IN2(n12697), .QN(g33622) );
  NAND2X0 U12704 ( .IN1(test_so50), .IN2(n10514), .QN(n12697) );
  NOR2X0 U12705 ( .IN1(n12698), .IN2(n12699), .QN(n12696) );
  NOR2X0 U12706 ( .IN1(n10122), .IN2(n12700), .QN(n12699) );
  NOR2X0 U12707 ( .IN1(test_so57), .IN2(n12701), .QN(n12698) );
  NAND2X0 U12708 ( .IN1(n12702), .IN2(n12687), .QN(n12701) );
  NAND2X0 U12709 ( .IN1(n12703), .IN2(n12695), .QN(n12687) );
  NOR2X0 U12710 ( .IN1(n11698), .IN2(n12704), .QN(n12703) );
  INVX0 U12711 ( .INP(n12705), .ZN(n12702) );
  NAND2X0 U12712 ( .IN1(n12706), .IN2(n12707), .QN(g33621) );
  NAND2X0 U12713 ( .IN1(n12708), .IN2(n12709), .QN(n12707) );
  NAND2X0 U12714 ( .IN1(n12710), .IN2(n12711), .QN(n12708) );
  NAND2X0 U12715 ( .IN1(n12712), .IN2(n10398), .QN(n12711) );
  NAND2X0 U12716 ( .IN1(n12713), .IN2(n12714), .QN(n12712) );
  NAND2X0 U12717 ( .IN1(n12715), .IN2(g5644), .QN(n12714) );
  NAND2X0 U12718 ( .IN1(n12716), .IN2(n12717), .QN(n12710) );
  NAND2X0 U12719 ( .IN1(n10513), .IN2(g5703), .QN(n12706) );
  NAND2X0 U12720 ( .IN1(n12718), .IN2(n12719), .QN(g33620) );
  NAND2X0 U12721 ( .IN1(n12720), .IN2(g5703), .QN(n12719) );
  NOR2X0 U12722 ( .IN1(n12721), .IN2(n12722), .QN(n12718) );
  NOR2X0 U12723 ( .IN1(n9903), .IN2(n10336), .QN(n12722) );
  NOR2X0 U12724 ( .IN1(n10485), .IN2(n12723), .QN(n12721) );
  NAND2X0 U12725 ( .IN1(n12724), .IN2(n5397), .QN(n12723) );
  AND2X1 U12726 ( .IN1(n12709), .IN2(n12717), .Q(n12724) );
  NAND2X0 U12727 ( .IN1(n12725), .IN2(n12717), .QN(n12709) );
  NOR2X0 U12728 ( .IN1(n11703), .IN2(n12726), .QN(n12725) );
  NAND2X0 U12729 ( .IN1(test_so81), .IN2(n12007), .QN(n11703) );
  NAND2X0 U12730 ( .IN1(n12727), .IN2(n12728), .QN(g33619) );
  NAND2X0 U12731 ( .IN1(n12729), .IN2(n12730), .QN(n12728) );
  NAND2X0 U12732 ( .IN1(n12731), .IN2(n12732), .QN(n12729) );
  NAND2X0 U12733 ( .IN1(n12733), .IN2(n10398), .QN(n12732) );
  NAND2X0 U12734 ( .IN1(n10662), .IN2(n12734), .QN(n12733) );
  NAND2X0 U12735 ( .IN1(n10108), .IN2(g5297), .QN(n12734) );
  NAND2X0 U12736 ( .IN1(n10665), .IN2(g33959), .QN(n12731) );
  NAND2X0 U12737 ( .IN1(n10514), .IN2(g5357), .QN(n12727) );
  NAND2X0 U12738 ( .IN1(n12735), .IN2(n12736), .QN(g33618) );
  NAND2X0 U12739 ( .IN1(n12737), .IN2(g5357), .QN(n12736) );
  NOR2X0 U12740 ( .IN1(n12738), .IN2(n12739), .QN(n12735) );
  NOR2X0 U12741 ( .IN1(n10038), .IN2(n10336), .QN(n12739) );
  NOR2X0 U12742 ( .IN1(n10485), .IN2(n12740), .QN(n12738) );
  NAND2X0 U12743 ( .IN1(n12741), .IN2(n5393), .QN(n12740) );
  AND2X1 U12744 ( .IN1(g33959), .IN2(n12730), .Q(n12741) );
  NAND2X0 U12745 ( .IN1(n12742), .IN2(n3023), .QN(n12730) );
  NOR2X0 U12746 ( .IN1(n10108), .IN2(n11698), .QN(n12742) );
  NAND2X0 U12747 ( .IN1(n12007), .IN2(n10132), .QN(n11698) );
  INVX0 U12748 ( .INP(n11328), .ZN(n12007) );
  NAND2X0 U12749 ( .IN1(n5323), .IN2(n12743), .QN(n11328) );
  NAND2X0 U12750 ( .IN1(n12744), .IN2(n12745), .QN(g33617) );
  NAND2X0 U12751 ( .IN1(n12746), .IN2(g4552), .QN(n12745) );
  NOR2X0 U12752 ( .IN1(n12017), .IN2(n12747), .QN(n12744) );
  NAND2X0 U12753 ( .IN1(n12748), .IN2(n12749), .QN(g33616) );
  NOR2X0 U12754 ( .IN1(n12017), .IN2(n12750), .QN(n12749) );
  NOR2X0 U12755 ( .IN1(n12751), .IN2(n12752), .QN(n12748) );
  NOR2X0 U12756 ( .IN1(n10046), .IN2(n10337), .QN(n12752) );
  NOR2X0 U12757 ( .IN1(n9768), .IN2(n12753), .QN(n12751) );
  NAND2X0 U12758 ( .IN1(n3064), .IN2(n12754), .QN(g33615) );
  NAND2X0 U12759 ( .IN1(n12755), .IN2(g4108), .QN(n12754) );
  NAND2X0 U12760 ( .IN1(n12756), .IN2(n10398), .QN(n12755) );
  NAND2X0 U12761 ( .IN1(n10787), .IN2(n9913), .QN(n12756) );
  NAND2X0 U12762 ( .IN1(n12757), .IN2(n12758), .QN(g33614) );
  NAND2X0 U12763 ( .IN1(n12759), .IN2(n12760), .QN(n12758) );
  NAND2X0 U12764 ( .IN1(n12761), .IN2(n12762), .QN(n12759) );
  NAND2X0 U12765 ( .IN1(n12763), .IN2(n10398), .QN(n12762) );
  NAND2X0 U12766 ( .IN1(n12764), .IN2(n12765), .QN(n12763) );
  NAND2X0 U12767 ( .IN1(n12766), .IN2(g3990), .QN(n12765) );
  NAND2X0 U12768 ( .IN1(n12767), .IN2(n12768), .QN(n12761) );
  NAND2X0 U12769 ( .IN1(n10513), .IN2(g4054), .QN(n12757) );
  NAND2X0 U12770 ( .IN1(n12769), .IN2(n12770), .QN(g33613) );
  NAND2X0 U12771 ( .IN1(n12771), .IN2(g4054), .QN(n12770) );
  NOR2X0 U12772 ( .IN1(n12772), .IN2(n12773), .QN(n12769) );
  NOR2X0 U12773 ( .IN1(n9905), .IN2(n10337), .QN(n12773) );
  NOR2X0 U12774 ( .IN1(n10485), .IN2(n12774), .QN(n12772) );
  NAND2X0 U12775 ( .IN1(n12775), .IN2(n5395), .QN(n12774) );
  AND2X1 U12776 ( .IN1(n12760), .IN2(n12768), .Q(n12775) );
  NAND2X0 U12777 ( .IN1(n12776), .IN2(n12768), .QN(n12760) );
  NOR2X0 U12778 ( .IN1(n11701), .IN2(n12704), .QN(n12776) );
  NAND2X0 U12779 ( .IN1(n12777), .IN2(n12778), .QN(g33612) );
  NAND2X0 U12780 ( .IN1(n12779), .IN2(n12780), .QN(n12778) );
  NAND2X0 U12781 ( .IN1(n12781), .IN2(n12782), .QN(n12779) );
  NAND2X0 U12782 ( .IN1(n12783), .IN2(n10399), .QN(n12782) );
  NAND2X0 U12783 ( .IN1(n12784), .IN2(n12785), .QN(n12783) );
  NAND2X0 U12784 ( .IN1(n12786), .IN2(g3639), .QN(n12785) );
  NAND2X0 U12785 ( .IN1(n12787), .IN2(n12788), .QN(n12781) );
  NAND2X0 U12786 ( .IN1(n10514), .IN2(g3703), .QN(n12777) );
  NAND2X0 U12787 ( .IN1(n12789), .IN2(n12790), .QN(g33611) );
  NAND2X0 U12788 ( .IN1(n12791), .IN2(g3703), .QN(n12790) );
  NOR2X0 U12789 ( .IN1(n12792), .IN2(n12793), .QN(n12789) );
  NOR2X0 U12790 ( .IN1(n9901), .IN2(n10337), .QN(n12793) );
  NOR2X0 U12791 ( .IN1(n10486), .IN2(n12794), .QN(n12792) );
  NAND2X0 U12792 ( .IN1(n12795), .IN2(n5399), .QN(n12794) );
  AND2X1 U12793 ( .IN1(n12780), .IN2(n12788), .Q(n12795) );
  NAND2X0 U12794 ( .IN1(n12796), .IN2(n12788), .QN(n12780) );
  NOR2X0 U12795 ( .IN1(n11697), .IN2(n12704), .QN(n12796) );
  INVX0 U12796 ( .INP(n3033), .ZN(n12704) );
  NAND2X0 U12797 ( .IN1(n11970), .IN2(n10132), .QN(n11697) );
  NAND2X0 U12798 ( .IN1(n12797), .IN2(n12798), .QN(g33610) );
  NAND2X0 U12799 ( .IN1(n10514), .IN2(g3352), .QN(n12798) );
  NAND2X0 U12800 ( .IN1(n12799), .IN2(n10399), .QN(n12797) );
  NOR2X0 U12801 ( .IN1(n12800), .IN2(n12801), .QN(n12799) );
  NOR2X0 U12802 ( .IN1(n12802), .IN2(n12803), .QN(n12801) );
  NAND2X0 U12803 ( .IN1(n12804), .IN2(n12805), .QN(n12803) );
  NAND2X0 U12804 ( .IN1(n12806), .IN2(g3288), .QN(n12805) );
  NAND2X0 U12805 ( .IN1(n12807), .IN2(n12808), .QN(n12804) );
  NAND2X0 U12806 ( .IN1(n12809), .IN2(n12810), .QN(g33609) );
  NAND2X0 U12807 ( .IN1(n12811), .IN2(g3352), .QN(n12810) );
  NOR2X0 U12808 ( .IN1(n12812), .IN2(n12813), .QN(n12809) );
  NOR2X0 U12809 ( .IN1(n9896), .IN2(n10337), .QN(n12813) );
  NOR2X0 U12810 ( .IN1(n10486), .IN2(n12814), .QN(n12812) );
  NAND2X0 U12811 ( .IN1(n12815), .IN2(n5604), .QN(n12814) );
  NOR2X0 U12812 ( .IN1(n12800), .IN2(n12806), .QN(n12815) );
  AND2X1 U12813 ( .IN1(n12816), .IN2(n12808), .Q(n12800) );
  NOR2X0 U12814 ( .IN1(n11701), .IN2(n12726), .QN(n12816) );
  INVX0 U12815 ( .INP(n3023), .ZN(n12726) );
  NAND2X0 U12816 ( .IN1(n11970), .IN2(test_so81), .QN(n11701) );
  INVX0 U12817 ( .INP(n11332), .ZN(n11970) );
  NAND2X0 U12818 ( .IN1(n12743), .IN2(g4311), .QN(n11332) );
  AND2X1 U12819 ( .IN1(n12817), .IN2(n11222), .Q(n12743) );
  XNOR2X1 U12820 ( .IN1(n12573), .IN2(n5506), .Q(n11222) );
  XOR2X1 U12821 ( .IN1(n5540), .IN2(g73), .Q(n12817) );
  NAND2X0 U12822 ( .IN1(n12818), .IN2(n12819), .QN(g33608) );
  NOR2X0 U12823 ( .IN1(n12820), .IN2(n12821), .QN(n12819) );
  AND2X1 U12824 ( .IN1(n10496), .IN2(test_so30), .Q(n12821) );
  NOR2X0 U12825 ( .IN1(n10486), .IN2(n12822), .QN(n12820) );
  NAND2X0 U12826 ( .IN1(n12034), .IN2(g2759), .QN(n12822) );
  NOR2X0 U12827 ( .IN1(n2787), .IN2(n12823), .QN(n12818) );
  NOR2X0 U12828 ( .IN1(g2759), .IN2(n12034), .QN(n12823) );
  NAND2X0 U12829 ( .IN1(n2790), .IN2(test_so30), .QN(n12034) );
  NAND2X0 U12830 ( .IN1(n12824), .IN2(n12825), .QN(g33607) );
  NAND2X0 U12831 ( .IN1(n10510), .IN2(g2555), .QN(n12825) );
  NOR2X0 U12832 ( .IN1(n12826), .IN2(n12827), .QN(n12824) );
  NOR2X0 U12833 ( .IN1(n5311), .IN2(n12828), .QN(n12827) );
  NOR2X0 U12834 ( .IN1(n12829), .IN2(n12830), .QN(n12828) );
  NOR2X0 U12835 ( .IN1(n3105), .IN2(n10463), .QN(n12829) );
  NOR2X0 U12836 ( .IN1(n12831), .IN2(n12832), .QN(n12826) );
  NAND2X0 U12837 ( .IN1(n12833), .IN2(n12834), .QN(n12832) );
  NAND2X0 U12838 ( .IN1(n12835), .IN2(n12836), .QN(n12834) );
  NAND2X0 U12839 ( .IN1(n12837), .IN2(n11744), .QN(n12836) );
  NOR2X0 U12840 ( .IN1(n5521), .IN2(n2726), .QN(n11744) );
  NAND2X0 U12841 ( .IN1(n11731), .IN2(n5519), .QN(n2726) );
  NOR2X0 U12842 ( .IN1(n12838), .IN2(g2599), .QN(n12837) );
  NAND2X0 U12843 ( .IN1(n3111), .IN2(n10399), .QN(n12835) );
  NAND2X0 U12844 ( .IN1(n12839), .IN2(n5524), .QN(n12833) );
  NOR2X0 U12845 ( .IN1(n9779), .IN2(n5521), .QN(n12839) );
  NAND2X0 U12846 ( .IN1(n12840), .IN2(n12841), .QN(g33606) );
  NAND2X0 U12847 ( .IN1(n12842), .IN2(g2675), .QN(n12841) );
  NOR2X0 U12848 ( .IN1(n12843), .IN2(n12844), .QN(n12840) );
  NOR2X0 U12849 ( .IN1(n5278), .IN2(n10337), .QN(n12844) );
  NOR2X0 U12850 ( .IN1(n10486), .IN2(n12845), .QN(n12843) );
  NAND2X0 U12851 ( .IN1(n5457), .IN2(n12056), .QN(n12845) );
  INVX0 U12852 ( .INP(n12041), .ZN(n12056) );
  NAND2X0 U12853 ( .IN1(n12846), .IN2(n12847), .QN(g33605) );
  OR2X1 U12854 ( .IN1(n12039), .IN2(n5278), .Q(n12847) );
  NOR2X0 U12855 ( .IN1(n12848), .IN2(n12849), .QN(n12846) );
  NOR2X0 U12856 ( .IN1(test_so48), .IN2(n12850), .QN(n12849) );
  NAND2X0 U12857 ( .IN1(n12851), .IN2(n5418), .QN(n12850) );
  NOR2X0 U12858 ( .IN1(n10487), .IN2(n12041), .QN(n12851) );
  NOR2X0 U12859 ( .IN1(n12852), .IN2(n10156), .QN(n12848) );
  NOR2X0 U12860 ( .IN1(n10487), .IN2(n12853), .QN(n12852) );
  NOR2X0 U12861 ( .IN1(n5418), .IN2(n12041), .QN(n12853) );
  NAND2X0 U12862 ( .IN1(n12854), .IN2(n12855), .QN(g33604) );
  NAND2X0 U12863 ( .IN1(test_so48), .IN2(n12842), .QN(n12855) );
  NAND2X0 U12864 ( .IN1(n12039), .IN2(g2661), .QN(n12854) );
  NAND2X0 U12865 ( .IN1(n12856), .IN2(n12857), .QN(g33603) );
  NAND2X0 U12866 ( .IN1(n12842), .IN2(g2648), .QN(n12857) );
  INVX0 U12867 ( .INP(n12039), .ZN(n12842) );
  NAND2X0 U12868 ( .IN1(n12039), .IN2(g2643), .QN(n12856) );
  NAND2X0 U12869 ( .IN1(n12041), .IN2(n10399), .QN(n12039) );
  NAND2X0 U12870 ( .IN1(n12858), .IN2(n5521), .QN(n12041) );
  NOR2X0 U12871 ( .IN1(n12057), .IN2(g2555), .QN(n12858) );
  NAND2X0 U12872 ( .IN1(n12859), .IN2(n12860), .QN(g33602) );
  NAND2X0 U12873 ( .IN1(n12074), .IN2(n12861), .QN(n12860) );
  INVX0 U12874 ( .INP(n3111), .ZN(n12861) );
  NOR2X0 U12875 ( .IN1(n5524), .IN2(n12057), .QN(n12074) );
  NOR2X0 U12876 ( .IN1(n12862), .IN2(n12863), .QN(n12859) );
  NOR2X0 U12877 ( .IN1(n10487), .IN2(n12864), .QN(n12863) );
  NAND2X0 U12878 ( .IN1(n12057), .IN2(g2629), .QN(n12864) );
  NOR2X0 U12879 ( .IN1(n5524), .IN2(n10337), .QN(n12862) );
  NAND2X0 U12880 ( .IN1(n12865), .IN2(n12866), .QN(g33601) );
  NAND2X0 U12881 ( .IN1(n12867), .IN2(n12047), .QN(n12866) );
  NOR2X0 U12882 ( .IN1(n3111), .IN2(n12057), .QN(n12867) );
  NOR2X0 U12883 ( .IN1(n12868), .IN2(n12869), .QN(n12865) );
  NOR2X0 U12884 ( .IN1(n5311), .IN2(n10338), .QN(n12869) );
  NOR2X0 U12885 ( .IN1(n10487), .IN2(n12870), .QN(n12868) );
  NAND2X0 U12886 ( .IN1(n12057), .IN2(g2599), .QN(n12870) );
  NAND2X0 U12887 ( .IN1(n12871), .IN2(n12872), .QN(g33600) );
  NAND2X0 U12888 ( .IN1(n12873), .IN2(n12874), .QN(n12872) );
  NOR2X0 U12889 ( .IN1(n3111), .IN2(n10463), .QN(n12874) );
  NOR2X0 U12890 ( .IN1(n12875), .IN2(g2629), .QN(n12873) );
  NOR2X0 U12891 ( .IN1(n12067), .IN2(g2555), .QN(n12875) );
  NOR2X0 U12892 ( .IN1(g2599), .IN2(n12057), .QN(n12067) );
  NAND2X0 U12893 ( .IN1(n12047), .IN2(n12057), .QN(n12871) );
  INVX0 U12894 ( .INP(n12053), .ZN(n12057) );
  NAND2X0 U12895 ( .IN1(n12060), .IN2(n12831), .QN(n12053) );
  INVX0 U12896 ( .INP(n475), .ZN(n12831) );
  NOR2X0 U12897 ( .IN1(n10067), .IN2(n12876), .QN(n475) );
  AND2X1 U12898 ( .IN1(n12877), .IN2(n5364), .Q(n12876) );
  NOR2X0 U12899 ( .IN1(test_so49), .IN2(n12878), .QN(n12877) );
  INVX0 U12900 ( .INP(n12093), .ZN(n12060) );
  NAND2X0 U12901 ( .IN1(n12879), .IN2(n12880), .QN(n12093) );
  NAND2X0 U12902 ( .IN1(n12881), .IN2(g2697), .QN(n12880) );
  NOR2X0 U12903 ( .IN1(n12286), .IN2(n11110), .QN(n12879) );
  INVX0 U12904 ( .INP(n12096), .ZN(n11110) );
  NAND2X0 U12905 ( .IN1(n2549), .IN2(g1300), .QN(n12096) );
  NOR2X0 U12906 ( .IN1(n10487), .IN2(n5351), .QN(n12047) );
  NAND2X0 U12907 ( .IN1(n12882), .IN2(n12883), .QN(g33599) );
  NOR2X0 U12908 ( .IN1(n12884), .IN2(n12885), .QN(n12883) );
  NOR2X0 U12909 ( .IN1(n10487), .IN2(n12886), .QN(n12885) );
  NAND2X0 U12910 ( .IN1(n12887), .IN2(n3131), .QN(n12886) );
  NOR2X0 U12911 ( .IN1(n12888), .IN2(n10677), .QN(n12887) );
  NOR2X0 U12912 ( .IN1(n9779), .IN2(n11754), .QN(n12888) );
  NOR2X0 U12913 ( .IN1(n10358), .IN2(n10131), .QN(n12884) );
  NOR2X0 U12914 ( .IN1(n12889), .IN2(n12890), .QN(n12882) );
  NOR2X0 U12915 ( .IN1(n5619), .IN2(n12891), .QN(n12890) );
  NOR2X0 U12916 ( .IN1(n12892), .IN2(n12830), .QN(n12891) );
  NOR2X0 U12917 ( .IN1(n3125), .IN2(n10463), .QN(n12892) );
  INVX0 U12918 ( .INP(n3121), .ZN(n12889) );
  NAND2X0 U12919 ( .IN1(n12893), .IN2(n12894), .QN(n3121) );
  NOR2X0 U12920 ( .IN1(g112), .IN2(n12895), .QN(n12894) );
  OR2X1 U12921 ( .IN1(n12838), .IN2(n2727), .Q(n12895) );
  NAND2X0 U12922 ( .IN1(n11731), .IN2(g504), .QN(n2727) );
  AND2X1 U12923 ( .IN1(n3116), .IN2(g518), .Q(n11731) );
  NOR2X0 U12924 ( .IN1(n11754), .IN2(n10677), .QN(n12893) );
  NAND2X0 U12925 ( .IN1(n5523), .IN2(g2495), .QN(n11754) );
  NAND2X0 U12926 ( .IN1(n12896), .IN2(n12897), .QN(g33598) );
  NAND2X0 U12927 ( .IN1(n12898), .IN2(g2541), .QN(n12897) );
  NOR2X0 U12928 ( .IN1(n12899), .IN2(n12900), .QN(n12896) );
  NOR2X0 U12929 ( .IN1(n5411), .IN2(n10338), .QN(n12900) );
  NOR2X0 U12930 ( .IN1(n10487), .IN2(n12901), .QN(n12899) );
  NAND2X0 U12931 ( .IN1(n5461), .IN2(n12121), .QN(n12901) );
  INVX0 U12932 ( .INP(n12106), .ZN(n12121) );
  NAND2X0 U12933 ( .IN1(n12902), .IN2(n12903), .QN(g33597) );
  OR2X1 U12934 ( .IN1(n12104), .IN2(n5411), .Q(n12903) );
  NOR2X0 U12935 ( .IN1(n12904), .IN2(n12905), .QN(n12902) );
  NOR2X0 U12936 ( .IN1(g2533), .IN2(n12906), .QN(n12905) );
  NAND2X0 U12937 ( .IN1(n12907), .IN2(n5420), .QN(n12906) );
  NOR2X0 U12938 ( .IN1(n10491), .IN2(n12106), .QN(n12907) );
  NOR2X0 U12939 ( .IN1(n5761), .IN2(n12908), .QN(n12904) );
  NOR2X0 U12940 ( .IN1(n10487), .IN2(n12909), .QN(n12908) );
  NOR2X0 U12941 ( .IN1(n5420), .IN2(n12106), .QN(n12909) );
  NAND2X0 U12942 ( .IN1(n12910), .IN2(n12911), .QN(g33596) );
  NAND2X0 U12943 ( .IN1(n12898), .IN2(g2533), .QN(n12911) );
  NAND2X0 U12944 ( .IN1(n12104), .IN2(g2527), .QN(n12910) );
  NAND2X0 U12945 ( .IN1(n12912), .IN2(n12913), .QN(g33595) );
  NAND2X0 U12946 ( .IN1(n12898), .IN2(g2514), .QN(n12913) );
  INVX0 U12947 ( .INP(n12104), .ZN(n12898) );
  NAND2X0 U12948 ( .IN1(n12104), .IN2(g2509), .QN(n12912) );
  NAND2X0 U12949 ( .IN1(n12106), .IN2(n10399), .QN(n12104) );
  NAND2X0 U12950 ( .IN1(n12914), .IN2(n5522), .QN(n12106) );
  NOR2X0 U12951 ( .IN1(test_so79), .IN2(n12122), .QN(n12914) );
  NAND2X0 U12952 ( .IN1(n12915), .IN2(n12916), .QN(g33594) );
  NAND2X0 U12953 ( .IN1(n10510), .IN2(g2465), .QN(n12916) );
  NOR2X0 U12954 ( .IN1(n12917), .IN2(n12918), .QN(n12915) );
  NOR2X0 U12955 ( .IN1(n3131), .IN2(n12139), .QN(n12918) );
  NAND2X0 U12956 ( .IN1(g2465), .IN2(n12118), .QN(n12139) );
  AND2X1 U12957 ( .IN1(g2495), .IN2(n12919), .Q(n12917) );
  NAND2X0 U12958 ( .IN1(n12920), .IN2(n12921), .QN(g33593) );
  NAND2X0 U12959 ( .IN1(n12919), .IN2(g2465), .QN(n12921) );
  NOR2X0 U12960 ( .IN1(n12922), .IN2(n12923), .QN(n12920) );
  NOR2X0 U12961 ( .IN1(n10487), .IN2(n12924), .QN(n12923) );
  NAND2X0 U12962 ( .IN1(n12146), .IN2(n12925), .QN(n12924) );
  INVX0 U12963 ( .INP(n3131), .ZN(n12925) );
  NOR2X0 U12964 ( .IN1(n10131), .IN2(n12122), .QN(n12146) );
  NOR2X0 U12965 ( .IN1(n5619), .IN2(n10338), .QN(n12922) );
  NAND2X0 U12966 ( .IN1(n12926), .IN2(n12927), .QN(g33592) );
  NAND2X0 U12967 ( .IN1(n12928), .IN2(n12929), .QN(n12927) );
  NOR2X0 U12968 ( .IN1(n3131), .IN2(n10462), .QN(n12929) );
  NOR2X0 U12969 ( .IN1(n12930), .IN2(g2495), .QN(n12928) );
  NOR2X0 U12970 ( .IN1(n12931), .IN2(test_so79), .QN(n12930) );
  NOR2X0 U12971 ( .IN1(n12122), .IN2(g2465), .QN(n12931) );
  INVX0 U12972 ( .INP(n12118), .ZN(n12122) );
  NAND2X0 U12973 ( .IN1(n12919), .IN2(test_so79), .QN(n12926) );
  NOR2X0 U12974 ( .IN1(n12118), .IN2(n10462), .QN(n12919) );
  NAND2X0 U12975 ( .IN1(n12125), .IN2(n10677), .QN(n12118) );
  NAND2X0 U12976 ( .IN1(g17423), .IN2(n12932), .QN(n10677) );
  NAND2X0 U12977 ( .IN1(n12933), .IN2(test_so49), .QN(n12932) );
  NOR2X0 U12978 ( .IN1(n5364), .IN2(n12878), .QN(n12933) );
  INVX0 U12979 ( .INP(n12158), .ZN(n12125) );
  NAND2X0 U12980 ( .IN1(n12934), .IN2(n12935), .QN(n12158) );
  NAND2X0 U12981 ( .IN1(n12936), .IN2(g2697), .QN(n12935) );
  NOR2X0 U12982 ( .IN1(n12286), .IN2(n11031), .QN(n12934) );
  NOR2X0 U12983 ( .IN1(g1291), .IN2(n5290), .QN(n11031) );
  NAND2X0 U12984 ( .IN1(n12937), .IN2(n12938), .QN(g33591) );
  NAND2X0 U12985 ( .IN1(n10509), .IN2(g2287), .QN(n12938) );
  NOR2X0 U12986 ( .IN1(n12939), .IN2(n12940), .QN(n12937) );
  NOR2X0 U12987 ( .IN1(n5310), .IN2(n12941), .QN(n12940) );
  NOR2X0 U12988 ( .IN1(n12942), .IN2(n12830), .QN(n12941) );
  NOR2X0 U12989 ( .IN1(n3145), .IN2(n10462), .QN(n12942) );
  NOR2X0 U12990 ( .IN1(n12943), .IN2(n12944), .QN(n12939) );
  NAND2X0 U12991 ( .IN1(n12945), .IN2(n12946), .QN(n12944) );
  NAND2X0 U12992 ( .IN1(n12947), .IN2(n12948), .QN(n12946) );
  NAND2X0 U12993 ( .IN1(n12949), .IN2(n11738), .QN(n12948) );
  NOR2X0 U12994 ( .IN1(n5537), .IN2(n3146), .QN(n11738) );
  NOR2X0 U12995 ( .IN1(n12838), .IN2(g2331), .QN(n12949) );
  NAND2X0 U12996 ( .IN1(n12950), .IN2(n10400), .QN(n12947) );
  NAND2X0 U12997 ( .IN1(n12951), .IN2(n5513), .QN(n12945) );
  NOR2X0 U12998 ( .IN1(n9779), .IN2(n5537), .QN(n12951) );
  INVX0 U12999 ( .INP(n3141), .ZN(n12943) );
  NAND2X0 U13000 ( .IN1(n12952), .IN2(n12953), .QN(g33590) );
  NAND2X0 U13001 ( .IN1(n12954), .IN2(g2407), .QN(n12953) );
  NOR2X0 U13002 ( .IN1(n12955), .IN2(n12956), .QN(n12952) );
  NOR2X0 U13003 ( .IN1(n10358), .IN2(n10153), .QN(n12956) );
  NOR2X0 U13004 ( .IN1(n10487), .IN2(n12957), .QN(n12955) );
  NAND2X0 U13005 ( .IN1(n5459), .IN2(n12185), .QN(n12957) );
  INVX0 U13006 ( .INP(n12170), .ZN(n12185) );
  NAND2X0 U13007 ( .IN1(n12958), .IN2(n12959), .QN(g33589) );
  NAND2X0 U13008 ( .IN1(test_so31), .IN2(n12954), .QN(n12959) );
  NOR2X0 U13009 ( .IN1(n12960), .IN2(n12961), .QN(n12958) );
  NOR2X0 U13010 ( .IN1(g2399), .IN2(n12962), .QN(n12961) );
  NAND2X0 U13011 ( .IN1(n12963), .IN2(n5421), .QN(n12962) );
  NOR2X0 U13012 ( .IN1(n10488), .IN2(n12170), .QN(n12963) );
  NOR2X0 U13013 ( .IN1(n5762), .IN2(n12964), .QN(n12960) );
  NOR2X0 U13014 ( .IN1(n10488), .IN2(n12965), .QN(n12964) );
  NOR2X0 U13015 ( .IN1(n5421), .IN2(n12170), .QN(n12965) );
  NAND2X0 U13016 ( .IN1(n12966), .IN2(n12967), .QN(g33588) );
  NAND2X0 U13017 ( .IN1(n12954), .IN2(g2399), .QN(n12967) );
  NAND2X0 U13018 ( .IN1(n12168), .IN2(g2393), .QN(n12966) );
  NAND2X0 U13019 ( .IN1(n12968), .IN2(n12969), .QN(g33587) );
  NAND2X0 U13020 ( .IN1(n12954), .IN2(g2380), .QN(n12969) );
  INVX0 U13021 ( .INP(n12168), .ZN(n12954) );
  NAND2X0 U13022 ( .IN1(n12168), .IN2(g2375), .QN(n12968) );
  NAND2X0 U13023 ( .IN1(n12170), .IN2(n10400), .QN(n12168) );
  NAND2X0 U13024 ( .IN1(n12970), .IN2(n5537), .QN(n12170) );
  NOR2X0 U13025 ( .IN1(n12182), .IN2(g2287), .QN(n12970) );
  NAND2X0 U13026 ( .IN1(n12971), .IN2(n12972), .QN(g33586) );
  NAND2X0 U13027 ( .IN1(n12202), .IN2(n12973), .QN(n12972) );
  NOR2X0 U13028 ( .IN1(n5513), .IN2(n12182), .QN(n12202) );
  NOR2X0 U13029 ( .IN1(n12974), .IN2(n12975), .QN(n12971) );
  NOR2X0 U13030 ( .IN1(n10488), .IN2(n12976), .QN(n12975) );
  NAND2X0 U13031 ( .IN1(n12182), .IN2(g2361), .QN(n12976) );
  NOR2X0 U13032 ( .IN1(n5513), .IN2(n10338), .QN(n12974) );
  NAND2X0 U13033 ( .IN1(n12977), .IN2(n12978), .QN(g33585) );
  NAND2X0 U13034 ( .IN1(n12979), .IN2(n12176), .QN(n12978) );
  NOR2X0 U13035 ( .IN1(n12182), .IN2(n12950), .QN(n12979) );
  NOR2X0 U13036 ( .IN1(n12980), .IN2(n12981), .QN(n12977) );
  NOR2X0 U13037 ( .IN1(n5310), .IN2(n10338), .QN(n12981) );
  NOR2X0 U13038 ( .IN1(n10488), .IN2(n12982), .QN(n12980) );
  NAND2X0 U13039 ( .IN1(n12182), .IN2(g2331), .QN(n12982) );
  NAND2X0 U13040 ( .IN1(n12983), .IN2(n12984), .QN(g33584) );
  NAND2X0 U13041 ( .IN1(n12985), .IN2(n12986), .QN(n12984) );
  NOR2X0 U13042 ( .IN1(n10488), .IN2(n12950), .QN(n12986) );
  INVX0 U13043 ( .INP(n12973), .ZN(n12950) );
  NAND2X0 U13044 ( .IN1(n3115), .IN2(n11730), .QN(n12973) );
  INVX0 U13045 ( .INP(n3146), .ZN(n11730) );
  NAND2X0 U13046 ( .IN1(n12987), .IN2(n3116), .QN(n3146) );
  NOR2X0 U13047 ( .IN1(n12988), .IN2(g2361), .QN(n12985) );
  NOR2X0 U13048 ( .IN1(n12989), .IN2(g2287), .QN(n12988) );
  NOR2X0 U13049 ( .IN1(n12182), .IN2(g2331), .QN(n12989) );
  NAND2X0 U13050 ( .IN1(n12176), .IN2(n12182), .QN(n12983) );
  NOR2X0 U13051 ( .IN1(n12220), .IN2(n3141), .QN(n12182) );
  NOR2X0 U13052 ( .IN1(n12990), .IN2(n9736), .QN(n3141) );
  AND2X1 U13053 ( .IN1(n12991), .IN2(n12992), .Q(n12990) );
  NAND2X0 U13054 ( .IN1(n12993), .IN2(n12994), .QN(n12220) );
  NAND2X0 U13055 ( .IN1(n5308), .IN2(n12881), .QN(n12994) );
  NOR2X0 U13056 ( .IN1(n5377), .IN2(n5347), .QN(n12881) );
  NOR2X0 U13057 ( .IN1(n12286), .IN2(n10995), .QN(n12993) );
  INVX0 U13058 ( .INP(n12222), .ZN(n10995) );
  NAND2X0 U13059 ( .IN1(n2549), .IN2(g1448), .QN(n12222) );
  NOR2X0 U13060 ( .IN1(n10488), .IN2(n5353), .QN(n12176) );
  NAND2X0 U13061 ( .IN1(n12995), .IN2(n12996), .QN(g33583) );
  NAND2X0 U13062 ( .IN1(n10509), .IN2(g2153), .QN(n12996) );
  NOR2X0 U13063 ( .IN1(n12997), .IN2(n12998), .QN(n12995) );
  NOR2X0 U13064 ( .IN1(n5620), .IN2(n12999), .QN(n12998) );
  NOR2X0 U13065 ( .IN1(n13000), .IN2(n12830), .QN(n12999) );
  NOR2X0 U13066 ( .IN1(n3164), .IN2(n10460), .QN(n13000) );
  NOR2X0 U13067 ( .IN1(n13001), .IN2(n13002), .QN(n12997) );
  NAND2X0 U13068 ( .IN1(n13003), .IN2(n13004), .QN(n13002) );
  NAND2X0 U13069 ( .IN1(n13005), .IN2(n13006), .QN(n13004) );
  NAND2X0 U13070 ( .IN1(n13007), .IN2(n11739), .QN(n13006) );
  NOR2X0 U13071 ( .IN1(n5538), .IN2(n3165), .QN(n11739) );
  NOR2X0 U13072 ( .IN1(n12838), .IN2(g2197), .QN(n13007) );
  NAND2X0 U13073 ( .IN1(n13008), .IN2(n10400), .QN(n13005) );
  NAND2X0 U13074 ( .IN1(n13009), .IN2(n5514), .QN(n13003) );
  NOR2X0 U13075 ( .IN1(n9779), .IN2(n5538), .QN(n13009) );
  INVX0 U13076 ( .INP(n3160), .ZN(n13001) );
  NAND2X0 U13077 ( .IN1(n13010), .IN2(n13011), .QN(g33582) );
  NAND2X0 U13078 ( .IN1(n13012), .IN2(g2273), .QN(n13011) );
  NOR2X0 U13079 ( .IN1(n13013), .IN2(n13014), .QN(n13010) );
  NOR2X0 U13080 ( .IN1(n5410), .IN2(n10338), .QN(n13014) );
  NOR2X0 U13081 ( .IN1(n10488), .IN2(n13015), .QN(n13013) );
  NAND2X0 U13082 ( .IN1(n5458), .IN2(n12248), .QN(n13015) );
  INVX0 U13083 ( .INP(n12233), .ZN(n12248) );
  NAND2X0 U13084 ( .IN1(n13016), .IN2(n13017), .QN(g33581) );
  OR2X1 U13085 ( .IN1(n12231), .IN2(n5410), .Q(n13017) );
  NOR2X0 U13086 ( .IN1(n13018), .IN2(n13019), .QN(n13016) );
  NOR2X0 U13087 ( .IN1(test_so62), .IN2(n13020), .QN(n13019) );
  NAND2X0 U13088 ( .IN1(n13021), .IN2(n5419), .QN(n13020) );
  NOR2X0 U13089 ( .IN1(n10488), .IN2(n12233), .QN(n13021) );
  NOR2X0 U13090 ( .IN1(n13022), .IN2(n10157), .QN(n13018) );
  NOR2X0 U13091 ( .IN1(n10488), .IN2(n13023), .QN(n13022) );
  NOR2X0 U13092 ( .IN1(n5419), .IN2(n12233), .QN(n13023) );
  NAND2X0 U13093 ( .IN1(n13024), .IN2(n13025), .QN(g33580) );
  NAND2X0 U13094 ( .IN1(test_so62), .IN2(n13012), .QN(n13025) );
  NAND2X0 U13095 ( .IN1(n12231), .IN2(g2259), .QN(n13024) );
  NAND2X0 U13096 ( .IN1(n13026), .IN2(n13027), .QN(g33579) );
  NAND2X0 U13097 ( .IN1(n13012), .IN2(g2246), .QN(n13027) );
  INVX0 U13098 ( .INP(n12231), .ZN(n13012) );
  NAND2X0 U13099 ( .IN1(n12231), .IN2(g2241), .QN(n13026) );
  NAND2X0 U13100 ( .IN1(n12233), .IN2(n10400), .QN(n12231) );
  NAND2X0 U13101 ( .IN1(n13028), .IN2(n5538), .QN(n12233) );
  NOR2X0 U13102 ( .IN1(n12245), .IN2(g2153), .QN(n13028) );
  NAND2X0 U13103 ( .IN1(n13029), .IN2(n13030), .QN(g33578) );
  NAND2X0 U13104 ( .IN1(n12265), .IN2(n13031), .QN(n13030) );
  NOR2X0 U13105 ( .IN1(n5514), .IN2(n12245), .QN(n12265) );
  NOR2X0 U13106 ( .IN1(n13032), .IN2(n13033), .QN(n13029) );
  NOR2X0 U13107 ( .IN1(n10489), .IN2(n13034), .QN(n13033) );
  NAND2X0 U13108 ( .IN1(n12245), .IN2(g2227), .QN(n13034) );
  NOR2X0 U13109 ( .IN1(n5514), .IN2(n10338), .QN(n13032) );
  NAND2X0 U13110 ( .IN1(n13035), .IN2(n13036), .QN(g33577) );
  NAND2X0 U13111 ( .IN1(n13037), .IN2(n12239), .QN(n13036) );
  NOR2X0 U13112 ( .IN1(n12245), .IN2(n13008), .QN(n13037) );
  NOR2X0 U13113 ( .IN1(n13038), .IN2(n13039), .QN(n13035) );
  NOR2X0 U13114 ( .IN1(n5620), .IN2(n10339), .QN(n13039) );
  NOR2X0 U13115 ( .IN1(n10489), .IN2(n13040), .QN(n13038) );
  NAND2X0 U13116 ( .IN1(n12245), .IN2(g2197), .QN(n13040) );
  NAND2X0 U13117 ( .IN1(n13041), .IN2(n13042), .QN(g33576) );
  NAND2X0 U13118 ( .IN1(n13043), .IN2(n13044), .QN(n13042) );
  NOR2X0 U13119 ( .IN1(n10489), .IN2(n13008), .QN(n13044) );
  INVX0 U13120 ( .INP(n13031), .ZN(n13008) );
  NAND2X0 U13121 ( .IN1(n3115), .IN2(n11729), .QN(n13031) );
  INVX0 U13122 ( .INP(n3165), .ZN(n11729) );
  NAND2X0 U13123 ( .IN1(n13045), .IN2(n3116), .QN(n3165) );
  NOR2X0 U13124 ( .IN1(n13046), .IN2(g2227), .QN(n13043) );
  NOR2X0 U13125 ( .IN1(n13047), .IN2(g2153), .QN(n13046) );
  NOR2X0 U13126 ( .IN1(n12245), .IN2(g2197), .QN(n13047) );
  NAND2X0 U13127 ( .IN1(n12239), .IN2(n12245), .QN(n13041) );
  NOR2X0 U13128 ( .IN1(n12283), .IN2(n3160), .QN(n12245) );
  NOR2X0 U13129 ( .IN1(n13048), .IN2(n9737), .QN(n3160) );
  AND2X1 U13130 ( .IN1(n13049), .IN2(n12992), .Q(n13048) );
  INVX0 U13131 ( .INP(n12878), .ZN(n12992) );
  NAND2X0 U13132 ( .IN1(n13050), .IN2(n13051), .QN(n12878) );
  NOR2X0 U13133 ( .IN1(g1564), .IN2(n13052), .QN(n13051) );
  OR2X1 U13134 ( .IN1(n10128), .IN2(n9753), .Q(n13052) );
  NOR2X0 U13135 ( .IN1(g1554), .IN2(n13053), .QN(n13050) );
  NAND2X0 U13136 ( .IN1(n5546), .IN2(n5441), .QN(n13053) );
  NOR2X0 U13137 ( .IN1(test_so49), .IN2(n5364), .QN(n13049) );
  NAND2X0 U13138 ( .IN1(n13054), .IN2(n13055), .QN(n12283) );
  NAND2X0 U13139 ( .IN1(n5308), .IN2(n12936), .QN(n13055) );
  NOR2X0 U13140 ( .IN1(g2704), .IN2(n5347), .QN(n12936) );
  NOR2X0 U13141 ( .IN1(n12286), .IN2(n10956), .QN(n13054) );
  NOR2X0 U13142 ( .IN1(g1291), .IN2(n5289), .QN(n10956) );
  AND2X1 U13143 ( .IN1(n13056), .IN2(n12639), .Q(n12286) );
  NAND2X0 U13144 ( .IN1(n11265), .IN2(n13057), .QN(n13056) );
  NOR2X0 U13145 ( .IN1(n10489), .IN2(n5356), .QN(n12239) );
  NAND2X0 U13146 ( .IN1(n13058), .IN2(n13059), .QN(g33575) );
  NOR2X0 U13147 ( .IN1(n13060), .IN2(n13061), .QN(n13059) );
  NOR2X0 U13148 ( .IN1(n10489), .IN2(n13062), .QN(n13061) );
  NAND2X0 U13149 ( .IN1(n13063), .IN2(n13064), .QN(n13062) );
  NOR2X0 U13150 ( .IN1(n13065), .IN2(n13066), .QN(n13063) );
  NOR2X0 U13151 ( .IN1(n9779), .IN2(n12324), .QN(n13065) );
  NOR2X0 U13152 ( .IN1(n5355), .IN2(n10339), .QN(n13060) );
  NOR2X0 U13153 ( .IN1(n13067), .IN2(n13068), .QN(n13058) );
  NOR2X0 U13154 ( .IN1(n5831), .IN2(n13069), .QN(n13068) );
  NOR2X0 U13155 ( .IN1(n13070), .IN2(n12830), .QN(n13069) );
  NOR2X0 U13156 ( .IN1(n10489), .IN2(n13071), .QN(n13070) );
  INVX0 U13157 ( .INP(n3180), .ZN(n13067) );
  NAND2X0 U13158 ( .IN1(n13072), .IN2(n13073), .QN(n3180) );
  AND2X1 U13159 ( .IN1(n13071), .IN2(n11749), .Q(n13073) );
  INVX0 U13160 ( .INP(n12324), .ZN(n11749) );
  NAND2X0 U13161 ( .IN1(n5505), .IN2(g2070), .QN(n12324) );
  NOR2X0 U13162 ( .IN1(n13074), .IN2(n13066), .QN(n13071) );
  NAND2X0 U13163 ( .IN1(n13075), .IN2(n13076), .QN(g33574) );
  NAND2X0 U13164 ( .IN1(n13077), .IN2(g2116), .QN(n13076) );
  NOR2X0 U13165 ( .IN1(n13078), .IN2(n13079), .QN(n13075) );
  NOR2X0 U13166 ( .IN1(n5848), .IN2(n10339), .QN(n13079) );
  NOR2X0 U13167 ( .IN1(n10489), .IN2(n13080), .QN(n13078) );
  NAND2X0 U13168 ( .IN1(n5463), .IN2(n12312), .QN(n13080) );
  INVX0 U13169 ( .INP(n12297), .ZN(n12312) );
  NAND2X0 U13170 ( .IN1(n13081), .IN2(n13082), .QN(g33573) );
  OR2X1 U13171 ( .IN1(n12295), .IN2(n5848), .Q(n13082) );
  NOR2X0 U13172 ( .IN1(n13083), .IN2(n13084), .QN(n13081) );
  NOR2X0 U13173 ( .IN1(g2108), .IN2(n13085), .QN(n13084) );
  NAND2X0 U13174 ( .IN1(n13086), .IN2(n5666), .QN(n13085) );
  NOR2X0 U13175 ( .IN1(n10489), .IN2(n12297), .QN(n13086) );
  NOR2X0 U13176 ( .IN1(n5452), .IN2(n13087), .QN(n13083) );
  NOR2X0 U13177 ( .IN1(n10489), .IN2(n13088), .QN(n13087) );
  NOR2X0 U13178 ( .IN1(n5666), .IN2(n12297), .QN(n13088) );
  NAND2X0 U13179 ( .IN1(n13089), .IN2(n13090), .QN(g33572) );
  NAND2X0 U13180 ( .IN1(n13077), .IN2(g2108), .QN(n13090) );
  NAND2X0 U13181 ( .IN1(n12295), .IN2(g2102), .QN(n13089) );
  NAND2X0 U13182 ( .IN1(n13091), .IN2(n13092), .QN(g33571) );
  NAND2X0 U13183 ( .IN1(n13077), .IN2(g2089), .QN(n13092) );
  INVX0 U13184 ( .INP(n12295), .ZN(n13077) );
  NAND2X0 U13185 ( .IN1(n12295), .IN2(g2084), .QN(n13091) );
  NAND2X0 U13186 ( .IN1(n12297), .IN2(n10400), .QN(n12295) );
  NAND2X0 U13187 ( .IN1(n13093), .IN2(n5535), .QN(n12297) );
  NOR2X0 U13188 ( .IN1(n12313), .IN2(g1996), .QN(n13093) );
  NAND2X0 U13189 ( .IN1(n13094), .IN2(n13095), .QN(g33570) );
  NAND2X0 U13190 ( .IN1(n10509), .IN2(g2040), .QN(n13095) );
  NOR2X0 U13191 ( .IN1(n13096), .IN2(n13097), .QN(n13094) );
  NOR2X0 U13192 ( .IN1(n13064), .IN2(n12331), .QN(n13097) );
  NAND2X0 U13193 ( .IN1(g2040), .IN2(n12309), .QN(n12331) );
  AND2X1 U13194 ( .IN1(g2070), .IN2(n13098), .Q(n13096) );
  NAND2X0 U13195 ( .IN1(n13099), .IN2(n13100), .QN(g33569) );
  NAND2X0 U13196 ( .IN1(n13098), .IN2(g2040), .QN(n13100) );
  NOR2X0 U13197 ( .IN1(n13101), .IN2(n13102), .QN(n13099) );
  NOR2X0 U13198 ( .IN1(n10489), .IN2(n13103), .QN(n13102) );
  NAND2X0 U13199 ( .IN1(n12338), .IN2(n13104), .QN(n13103) );
  NOR2X0 U13200 ( .IN1(n5355), .IN2(n12313), .QN(n12338) );
  NOR2X0 U13201 ( .IN1(n5831), .IN2(n10339), .QN(n13101) );
  NAND2X0 U13202 ( .IN1(n13105), .IN2(n13106), .QN(g33568) );
  NAND2X0 U13203 ( .IN1(n13107), .IN2(n13108), .QN(n13106) );
  NOR2X0 U13204 ( .IN1(n10490), .IN2(n13064), .QN(n13108) );
  INVX0 U13205 ( .INP(n13104), .ZN(n13064) );
  NAND2X0 U13206 ( .IN1(n3115), .IN2(n11728), .QN(n13104) );
  INVX0 U13207 ( .INP(n13074), .ZN(n11728) );
  NAND2X0 U13208 ( .IN1(n13109), .IN2(n3195), .QN(n13074) );
  NOR2X0 U13209 ( .IN1(n5287), .IN2(g504), .QN(n13109) );
  NOR2X0 U13210 ( .IN1(n13110), .IN2(g2070), .QN(n13107) );
  NOR2X0 U13211 ( .IN1(n13111), .IN2(g1996), .QN(n13110) );
  NOR2X0 U13212 ( .IN1(n12313), .IN2(g2040), .QN(n13111) );
  INVX0 U13213 ( .INP(n12309), .ZN(n12313) );
  NAND2X0 U13214 ( .IN1(n13098), .IN2(g1996), .QN(n13105) );
  NOR2X0 U13215 ( .IN1(n12309), .IN2(n10459), .QN(n13098) );
  NAND2X0 U13216 ( .IN1(n12316), .IN2(n13066), .QN(n12309) );
  NAND2X0 U13217 ( .IN1(g1087), .IN2(n13112), .QN(n13066) );
  NAND2X0 U13218 ( .IN1(n13113), .IN2(n5599), .QN(n13112) );
  NOR2X0 U13219 ( .IN1(n13114), .IN2(g1171), .QN(n13113) );
  INVX0 U13220 ( .INP(n12350), .ZN(n12316) );
  NAND2X0 U13221 ( .IN1(n13115), .IN2(n13116), .QN(n12350) );
  NAND2X0 U13222 ( .IN1(n13117), .IN2(g2138), .QN(n13116) );
  NOR2X0 U13223 ( .IN1(n12547), .IN2(n11113), .QN(n13115) );
  INVX0 U13224 ( .INP(n12353), .ZN(n11113) );
  NAND2X0 U13225 ( .IN1(n5286), .IN2(g956), .QN(n12353) );
  NAND2X0 U13226 ( .IN1(n13118), .IN2(n13119), .QN(g33567) );
  NAND2X0 U13227 ( .IN1(test_so8), .IN2(n10515), .QN(n13119) );
  NOR2X0 U13228 ( .IN1(n13120), .IN2(n13121), .QN(n13118) );
  NOR2X0 U13229 ( .IN1(n5828), .IN2(n13122), .QN(n13121) );
  NOR2X0 U13230 ( .IN1(n13123), .IN2(n12830), .QN(n13122) );
  NOR2X0 U13231 ( .IN1(n10490), .IN2(n13124), .QN(n13123) );
  NOR2X0 U13232 ( .IN1(n11723), .IN2(n13125), .QN(n13124) );
  NOR2X0 U13233 ( .IN1(n13126), .IN2(n13125), .QN(n13120) );
  NOR2X0 U13234 ( .IN1(n13127), .IN2(n13128), .QN(n13126) );
  NOR2X0 U13235 ( .IN1(n13129), .IN2(g112), .QN(n13128) );
  NOR2X0 U13236 ( .IN1(n13130), .IN2(n13131), .QN(n13129) );
  NOR2X0 U13237 ( .IN1(n10490), .IN2(n13132), .QN(n13131) );
  NOR2X0 U13238 ( .IN1(n11723), .IN2(n13133), .QN(n13130) );
  NAND2X0 U13239 ( .IN1(n11753), .IN2(n11591), .QN(n13133) );
  INVX0 U13240 ( .INP(n12390), .ZN(n11753) );
  NOR2X0 U13241 ( .IN1(n13132), .IN2(n13134), .QN(n13127) );
  NAND2X0 U13242 ( .IN1(n12390), .IN2(n10401), .QN(n13134) );
  NAND2X0 U13243 ( .IN1(n5503), .IN2(g1936), .QN(n12390) );
  NAND2X0 U13244 ( .IN1(n13135), .IN2(n13136), .QN(g33566) );
  NAND2X0 U13245 ( .IN1(n13137), .IN2(g1982), .QN(n13136) );
  NOR2X0 U13246 ( .IN1(n13138), .IN2(n13139), .QN(n13135) );
  NOR2X0 U13247 ( .IN1(n5845), .IN2(n10339), .QN(n13139) );
  NOR2X0 U13248 ( .IN1(n10490), .IN2(n13140), .QN(n13138) );
  NAND2X0 U13249 ( .IN1(n5462), .IN2(n12378), .QN(n13140) );
  INVX0 U13250 ( .INP(n12363), .ZN(n12378) );
  NAND2X0 U13251 ( .IN1(n13141), .IN2(n13142), .QN(g33565) );
  OR2X1 U13252 ( .IN1(n12361), .IN2(n5845), .Q(n13142) );
  NOR2X0 U13253 ( .IN1(n13143), .IN2(n13144), .QN(n13141) );
  NOR2X0 U13254 ( .IN1(g1974), .IN2(n13145), .QN(n13144) );
  NAND2X0 U13255 ( .IN1(n13146), .IN2(n5664), .QN(n13145) );
  NOR2X0 U13256 ( .IN1(n10490), .IN2(n12363), .QN(n13146) );
  NOR2X0 U13257 ( .IN1(n5450), .IN2(n13147), .QN(n13143) );
  NOR2X0 U13258 ( .IN1(n10490), .IN2(n13148), .QN(n13147) );
  NOR2X0 U13259 ( .IN1(n5664), .IN2(n12363), .QN(n13148) );
  NAND2X0 U13260 ( .IN1(n13149), .IN2(n13150), .QN(g33564) );
  NAND2X0 U13261 ( .IN1(n13137), .IN2(g1974), .QN(n13150) );
  NAND2X0 U13262 ( .IN1(n12361), .IN2(g1968), .QN(n13149) );
  NAND2X0 U13263 ( .IN1(n13151), .IN2(n13152), .QN(g33563) );
  NAND2X0 U13264 ( .IN1(n13137), .IN2(g1955), .QN(n13152) );
  INVX0 U13265 ( .INP(n12361), .ZN(n13137) );
  NAND2X0 U13266 ( .IN1(n12361), .IN2(g1950), .QN(n13151) );
  NAND2X0 U13267 ( .IN1(n12363), .IN2(n10401), .QN(n12361) );
  NAND2X0 U13268 ( .IN1(n13153), .IN2(n5534), .QN(n12363) );
  NOR2X0 U13269 ( .IN1(test_so8), .IN2(n12379), .QN(n13153) );
  NAND2X0 U13270 ( .IN1(n13154), .IN2(n13155), .QN(g33562) );
  NAND2X0 U13271 ( .IN1(n10509), .IN2(g1906), .QN(n13155) );
  NOR2X0 U13272 ( .IN1(n13156), .IN2(n13157), .QN(n13154) );
  NOR2X0 U13273 ( .IN1(n13158), .IN2(n12397), .QN(n13157) );
  NAND2X0 U13274 ( .IN1(g1906), .IN2(n12375), .QN(n12397) );
  AND2X1 U13275 ( .IN1(g1936), .IN2(n13159), .Q(n13156) );
  NAND2X0 U13276 ( .IN1(n13160), .IN2(n13161), .QN(g33561) );
  NAND2X0 U13277 ( .IN1(n13159), .IN2(g1906), .QN(n13161) );
  NOR2X0 U13278 ( .IN1(n13162), .IN2(n13163), .QN(n13160) );
  NOR2X0 U13279 ( .IN1(n10490), .IN2(n13164), .QN(n13163) );
  NAND2X0 U13280 ( .IN1(n12404), .IN2(n13132), .QN(n13164) );
  NOR2X0 U13281 ( .IN1(n10137), .IN2(n12379), .QN(n12404) );
  NOR2X0 U13282 ( .IN1(n5828), .IN2(n10339), .QN(n13162) );
  NAND2X0 U13283 ( .IN1(n13165), .IN2(n13166), .QN(g33560) );
  NAND2X0 U13284 ( .IN1(n13167), .IN2(n13168), .QN(n13166) );
  NOR2X0 U13285 ( .IN1(n10490), .IN2(n13158), .QN(n13168) );
  INVX0 U13286 ( .INP(n13132), .ZN(n13158) );
  NAND2X0 U13287 ( .IN1(n3115), .IN2(n11752), .QN(n13132) );
  INVX0 U13288 ( .INP(n11723), .ZN(n11752) );
  NAND2X0 U13289 ( .IN1(n13169), .IN2(n3195), .QN(n11723) );
  NOR2X0 U13290 ( .IN1(n5519), .IN2(n5287), .QN(n13169) );
  NOR2X0 U13291 ( .IN1(n13170), .IN2(g1936), .QN(n13167) );
  NOR2X0 U13292 ( .IN1(n13171), .IN2(test_so8), .QN(n13170) );
  NOR2X0 U13293 ( .IN1(n12379), .IN2(g1906), .QN(n13171) );
  INVX0 U13294 ( .INP(n12375), .ZN(n12379) );
  NAND2X0 U13295 ( .IN1(n13159), .IN2(test_so8), .QN(n13165) );
  NOR2X0 U13296 ( .IN1(n12375), .IN2(n10458), .QN(n13159) );
  NAND2X0 U13297 ( .IN1(n12382), .IN2(n13125), .QN(n12375) );
  NAND2X0 U13298 ( .IN1(g17400), .IN2(n13172), .QN(n13125) );
  NAND2X0 U13299 ( .IN1(n13173), .IN2(n13174), .QN(n13172) );
  INVX0 U13300 ( .INP(n12416), .ZN(n12382) );
  NAND2X0 U13301 ( .IN1(n13175), .IN2(n13176), .QN(n12416) );
  NAND2X0 U13302 ( .IN1(n13177), .IN2(g2138), .QN(n13176) );
  NOR2X0 U13303 ( .IN1(n12547), .IN2(n11032), .QN(n13175) );
  INVX0 U13304 ( .INP(n12418), .ZN(n11032) );
  NAND2X0 U13305 ( .IN1(n5286), .IN2(g1129), .QN(n12418) );
  NAND2X0 U13306 ( .IN1(n13178), .IN2(n13179), .QN(g33559) );
  NAND2X0 U13307 ( .IN1(n10509), .IN2(g1728), .QN(n13179) );
  NOR2X0 U13308 ( .IN1(n13180), .IN2(n13181), .QN(n13178) );
  NOR2X0 U13309 ( .IN1(n5830), .IN2(n13182), .QN(n13181) );
  NOR2X0 U13310 ( .IN1(n13183), .IN2(n12830), .QN(n13182) );
  INVX0 U13311 ( .INP(n13184), .ZN(n12830) );
  NOR2X0 U13312 ( .IN1(n10490), .IN2(n13185), .QN(n13183) );
  NOR2X0 U13313 ( .IN1(n11743), .IN2(n13186), .QN(n13185) );
  NOR2X0 U13314 ( .IN1(n13186), .IN2(n13187), .QN(n13180) );
  NAND2X0 U13315 ( .IN1(n13188), .IN2(n13189), .QN(n13187) );
  NAND2X0 U13316 ( .IN1(n13190), .IN2(n13191), .QN(n13189) );
  NAND2X0 U13317 ( .IN1(n13192), .IN2(n13193), .QN(n13191) );
  NOR2X0 U13318 ( .IN1(n5536), .IN2(n12838), .QN(n13193) );
  NOR2X0 U13319 ( .IN1(n11743), .IN2(g1772), .QN(n13192) );
  NAND2X0 U13320 ( .IN1(n13194), .IN2(n10401), .QN(n13190) );
  NAND2X0 U13321 ( .IN1(n13195), .IN2(n5504), .QN(n13188) );
  NOR2X0 U13322 ( .IN1(n9779), .IN2(n5536), .QN(n13195) );
  NAND2X0 U13323 ( .IN1(n13196), .IN2(n13197), .QN(g33558) );
  NAND2X0 U13324 ( .IN1(n13198), .IN2(g1848), .QN(n13197) );
  NOR2X0 U13325 ( .IN1(n13199), .IN2(n13200), .QN(n13196) );
  NOR2X0 U13326 ( .IN1(n5847), .IN2(n10339), .QN(n13200) );
  NOR2X0 U13327 ( .IN1(n10490), .IN2(n13201), .QN(n13199) );
  NAND2X0 U13328 ( .IN1(n5464), .IN2(n12443), .QN(n13201) );
  INVX0 U13329 ( .INP(n12428), .ZN(n12443) );
  NAND2X0 U13330 ( .IN1(n13202), .IN2(n13203), .QN(g33557) );
  OR2X1 U13331 ( .IN1(n12426), .IN2(n5847), .Q(n13203) );
  NOR2X0 U13332 ( .IN1(n13204), .IN2(n13205), .QN(n13202) );
  NOR2X0 U13333 ( .IN1(g1840), .IN2(n13206), .QN(n13205) );
  NAND2X0 U13334 ( .IN1(n13207), .IN2(n5665), .QN(n13206) );
  NOR2X0 U13335 ( .IN1(n10491), .IN2(n12428), .QN(n13207) );
  NOR2X0 U13336 ( .IN1(n5451), .IN2(n13208), .QN(n13204) );
  NOR2X0 U13337 ( .IN1(n10491), .IN2(n13209), .QN(n13208) );
  NOR2X0 U13338 ( .IN1(n5665), .IN2(n12428), .QN(n13209) );
  NAND2X0 U13339 ( .IN1(n13210), .IN2(n13211), .QN(g33556) );
  NAND2X0 U13340 ( .IN1(n13198), .IN2(g1840), .QN(n13211) );
  NAND2X0 U13341 ( .IN1(n12426), .IN2(g1834), .QN(n13210) );
  NAND2X0 U13342 ( .IN1(n13212), .IN2(n13213), .QN(g33555) );
  NAND2X0 U13343 ( .IN1(n13198), .IN2(g1821), .QN(n13213) );
  INVX0 U13344 ( .INP(n12426), .ZN(n13198) );
  NAND2X0 U13345 ( .IN1(n12426), .IN2(g1816), .QN(n13212) );
  NAND2X0 U13346 ( .IN1(n12428), .IN2(n10401), .QN(n12426) );
  NAND2X0 U13347 ( .IN1(n13214), .IN2(n5536), .QN(n12428) );
  NOR2X0 U13348 ( .IN1(n12444), .IN2(g1728), .QN(n13214) );
  NAND2X0 U13349 ( .IN1(n13215), .IN2(n13216), .QN(g33554) );
  NAND2X0 U13350 ( .IN1(n12461), .IN2(n13217), .QN(n13216) );
  NOR2X0 U13351 ( .IN1(n5504), .IN2(n12444), .QN(n12461) );
  NOR2X0 U13352 ( .IN1(n13218), .IN2(n13219), .QN(n13215) );
  NOR2X0 U13353 ( .IN1(n10491), .IN2(n13220), .QN(n13219) );
  NAND2X0 U13354 ( .IN1(n12444), .IN2(g1802), .QN(n13220) );
  NOR2X0 U13355 ( .IN1(n5504), .IN2(n10340), .QN(n13218) );
  NAND2X0 U13356 ( .IN1(n13221), .IN2(n13222), .QN(g33553) );
  NAND2X0 U13357 ( .IN1(n13223), .IN2(n12434), .QN(n13222) );
  NOR2X0 U13358 ( .IN1(n12444), .IN2(n13194), .QN(n13223) );
  NOR2X0 U13359 ( .IN1(n13224), .IN2(n13225), .QN(n13221) );
  NOR2X0 U13360 ( .IN1(n5830), .IN2(n10340), .QN(n13225) );
  NOR2X0 U13361 ( .IN1(n10491), .IN2(n13226), .QN(n13224) );
  NAND2X0 U13362 ( .IN1(n12444), .IN2(g1772), .QN(n13226) );
  NAND2X0 U13363 ( .IN1(n13227), .IN2(n13228), .QN(g33552) );
  NAND2X0 U13364 ( .IN1(n13229), .IN2(n13230), .QN(n13228) );
  NOR2X0 U13365 ( .IN1(n10491), .IN2(n13194), .QN(n13230) );
  INVX0 U13366 ( .INP(n13217), .ZN(n13194) );
  NAND2X0 U13367 ( .IN1(n3115), .IN2(n11725), .QN(n13217) );
  INVX0 U13368 ( .INP(n11743), .ZN(n11725) );
  NAND2X0 U13369 ( .IN1(n12987), .IN2(n3195), .QN(n11743) );
  NOR2X0 U13370 ( .IN1(n5519), .IN2(g518), .QN(n12987) );
  NOR2X0 U13371 ( .IN1(n13231), .IN2(g1802), .QN(n13229) );
  NOR2X0 U13372 ( .IN1(n13232), .IN2(g1728), .QN(n13231) );
  NOR2X0 U13373 ( .IN1(n12444), .IN2(g1772), .QN(n13232) );
  NAND2X0 U13374 ( .IN1(n12434), .IN2(n12444), .QN(n13227) );
  INVX0 U13375 ( .INP(n12440), .ZN(n12444) );
  NAND2X0 U13376 ( .IN1(n12447), .IN2(n13186), .QN(n12440) );
  NAND2X0 U13377 ( .IN1(test_so44), .IN2(n13233), .QN(n13186) );
  NAND2X0 U13378 ( .IN1(n13234), .IN2(n13174), .QN(n13233) );
  INVX0 U13379 ( .INP(n13114), .ZN(n13174) );
  INVX0 U13380 ( .INP(n12479), .ZN(n12447) );
  NAND2X0 U13381 ( .IN1(n13235), .IN2(n13236), .QN(n12479) );
  NAND2X0 U13382 ( .IN1(n5275), .IN2(n13117), .QN(n13236) );
  NOR2X0 U13383 ( .IN1(n5487), .IN2(n5307), .QN(n13117) );
  NOR2X0 U13384 ( .IN1(n12547), .IN2(n10996), .QN(n13235) );
  NOR2X0 U13385 ( .IN1(g947), .IN2(n5478), .QN(n10996) );
  NOR2X0 U13386 ( .IN1(n10491), .IN2(n5352), .QN(n12434) );
  NAND2X0 U13387 ( .IN1(n13237), .IN2(n13238), .QN(g33551) );
  NOR2X0 U13388 ( .IN1(n13239), .IN2(n13240), .QN(n13238) );
  NOR2X0 U13389 ( .IN1(n10491), .IN2(n13241), .QN(n13240) );
  NOR2X0 U13390 ( .IN1(n13242), .IN2(n13243), .QN(n13241) );
  NOR2X0 U13391 ( .IN1(n13244), .IN2(n10134), .QN(n13243) );
  AND2X1 U13392 ( .IN1(n11724), .IN2(g33533), .Q(n13244) );
  NOR2X0 U13393 ( .IN1(n13245), .IN2(n13246), .QN(n13242) );
  NAND2X0 U13394 ( .IN1(g33533), .IN2(n13247), .QN(n13246) );
  NAND2X0 U13395 ( .IN1(g31862), .IN2(g112), .QN(n13247) );
  NOR2X0 U13396 ( .IN1(n5362), .IN2(n10340), .QN(n13239) );
  NOR2X0 U13397 ( .IN1(n13248), .IN2(n13249), .QN(n13237) );
  NOR2X0 U13398 ( .IN1(n13184), .IN2(n10134), .QN(n13249) );
  NOR2X0 U13399 ( .IN1(n13250), .IN2(n13251), .QN(n13248) );
  NAND2X0 U13400 ( .IN1(g33533), .IN2(g31862), .QN(n13251) );
  NAND2X0 U13401 ( .IN1(n13072), .IN2(n11724), .QN(n13250) );
  NOR2X0 U13402 ( .IN1(n12838), .IN2(g112), .QN(n13072) );
  NAND2X0 U13403 ( .IN1(n13252), .IN2(n13253), .QN(g33550) );
  NAND2X0 U13404 ( .IN1(n13254), .IN2(g1714), .QN(n13253) );
  NOR2X0 U13405 ( .IN1(n13255), .IN2(n13256), .QN(n13252) );
  NOR2X0 U13406 ( .IN1(n5412), .IN2(n10340), .QN(n13256) );
  NOR2X0 U13407 ( .IN1(n10491), .IN2(n13257), .QN(n13255) );
  NAND2X0 U13408 ( .IN1(n5460), .IN2(n12507), .QN(n13257) );
  INVX0 U13409 ( .INP(n12492), .ZN(n12507) );
  NAND2X0 U13410 ( .IN1(n13258), .IN2(n13259), .QN(g33549) );
  OR2X1 U13411 ( .IN1(n12490), .IN2(n5412), .Q(n13259) );
  NOR2X0 U13412 ( .IN1(n13260), .IN2(n13261), .QN(n13258) );
  NOR2X0 U13413 ( .IN1(test_so15), .IN2(n13262), .QN(n13261) );
  NAND2X0 U13414 ( .IN1(n13263), .IN2(n5417), .QN(n13262) );
  NOR2X0 U13415 ( .IN1(n10495), .IN2(n12492), .QN(n13263) );
  NOR2X0 U13416 ( .IN1(n13264), .IN2(n10158), .QN(n13260) );
  NOR2X0 U13417 ( .IN1(n10496), .IN2(n13265), .QN(n13264) );
  NOR2X0 U13418 ( .IN1(n5417), .IN2(n12492), .QN(n13265) );
  NAND2X0 U13419 ( .IN1(n13266), .IN2(n13267), .QN(g33548) );
  NAND2X0 U13420 ( .IN1(test_so15), .IN2(n13254), .QN(n13267) );
  NAND2X0 U13421 ( .IN1(n12490), .IN2(g1700), .QN(n13266) );
  NAND2X0 U13422 ( .IN1(n13268), .IN2(n13269), .QN(g33547) );
  NAND2X0 U13423 ( .IN1(n13254), .IN2(g1687), .QN(n13269) );
  INVX0 U13424 ( .INP(n12490), .ZN(n13254) );
  NAND2X0 U13425 ( .IN1(n12490), .IN2(g1682), .QN(n13268) );
  NAND2X0 U13426 ( .IN1(n12492), .IN2(n10402), .QN(n12490) );
  NAND2X0 U13427 ( .IN1(n13270), .IN2(n5598), .QN(n12492) );
  NOR2X0 U13428 ( .IN1(n12508), .IN2(g1592), .QN(n13270) );
  NAND2X0 U13429 ( .IN1(n13271), .IN2(n13272), .QN(g33546) );
  NAND2X0 U13430 ( .IN1(n10508), .IN2(g1636), .QN(n13272) );
  NOR2X0 U13431 ( .IN1(n13273), .IN2(n13274), .QN(n13271) );
  NOR2X0 U13432 ( .IN1(n13275), .IN2(n12525), .QN(n13274) );
  NAND2X0 U13433 ( .IN1(g1636), .IN2(n12504), .QN(n12525) );
  AND2X1 U13434 ( .IN1(g1668), .IN2(n13276), .Q(n13273) );
  NAND2X0 U13435 ( .IN1(n13277), .IN2(n13278), .QN(g33545) );
  NAND2X0 U13436 ( .IN1(n13276), .IN2(g1636), .QN(n13278) );
  NOR2X0 U13437 ( .IN1(n13279), .IN2(n13280), .QN(n13277) );
  NOR2X0 U13438 ( .IN1(n10495), .IN2(n13281), .QN(n13280) );
  NAND2X0 U13439 ( .IN1(n12532), .IN2(n13245), .QN(n13281) );
  NOR2X0 U13440 ( .IN1(n5362), .IN2(n12508), .QN(n12532) );
  NOR2X0 U13441 ( .IN1(n10358), .IN2(n10134), .QN(n13279) );
  NAND2X0 U13442 ( .IN1(n13282), .IN2(n13283), .QN(g33544) );
  NAND2X0 U13443 ( .IN1(n13284), .IN2(n13285), .QN(n13283) );
  NOR2X0 U13444 ( .IN1(n10496), .IN2(n13275), .QN(n13285) );
  INVX0 U13445 ( .INP(n13245), .ZN(n13275) );
  NAND2X0 U13446 ( .IN1(n3115), .IN2(n11724), .QN(n13245) );
  AND2X1 U13447 ( .IN1(n13045), .IN2(n3195), .Q(n11724) );
  NOR2X0 U13448 ( .IN1(g504), .IN2(g518), .QN(n13045) );
  NOR2X0 U13449 ( .IN1(n13286), .IN2(g1668), .QN(n13284) );
  NOR2X0 U13450 ( .IN1(n13287), .IN2(g1592), .QN(n13286) );
  NOR2X0 U13451 ( .IN1(n12508), .IN2(g1636), .QN(n13287) );
  NAND2X0 U13452 ( .IN1(n13276), .IN2(g1592), .QN(n13282) );
  NOR2X0 U13453 ( .IN1(n12504), .IN2(n10458), .QN(n13276) );
  INVX0 U13454 ( .INP(n12508), .ZN(n12504) );
  NOR2X0 U13455 ( .IN1(n12544), .IN2(g33533), .QN(n12508) );
  NAND2X0 U13456 ( .IN1(n13288), .IN2(n13289), .QN(n12544) );
  NAND2X0 U13457 ( .IN1(n5275), .IN2(n13177), .QN(n13289) );
  NOR2X0 U13458 ( .IN1(g2145), .IN2(n5487), .QN(n13177) );
  NOR2X0 U13459 ( .IN1(n12547), .IN2(n10957), .QN(n13288) );
  INVX0 U13460 ( .INP(n12546), .ZN(n10957) );
  NAND2X0 U13461 ( .IN1(n5286), .IN2(g1135), .QN(n12546) );
  AND2X1 U13462 ( .IN1(n13290), .IN2(n12639), .Q(n12547) );
  INVX0 U13463 ( .INP(g134), .ZN(n12639) );
  NAND2X0 U13464 ( .IN1(n11265), .IN2(n11355), .QN(n13290) );
  NOR2X0 U13465 ( .IN1(g209), .IN2(n5520), .QN(n11265) );
  NAND2X0 U13466 ( .IN1(n13291), .IN2(n13292), .QN(g33543) );
  NAND2X0 U13467 ( .IN1(n13293), .IN2(n13294), .QN(n13292) );
  NAND2X0 U13468 ( .IN1(n13295), .IN2(n13296), .QN(n13294) );
  NAND2X0 U13469 ( .IN1(n9762), .IN2(n13297), .QN(n13296) );
  INVX0 U13470 ( .INP(n13298), .ZN(n13295) );
  NOR2X0 U13471 ( .IN1(n9685), .IN2(n10458), .QN(n13293) );
  NAND2X0 U13472 ( .IN1(n13299), .IN2(g1373), .QN(n13291) );
  NAND2X0 U13473 ( .IN1(n13300), .IN2(n10402), .QN(n13299) );
  NAND2X0 U13474 ( .IN1(n13301), .IN2(n9685), .QN(n13300) );
  NOR2X0 U13475 ( .IN1(n13302), .IN2(n13298), .QN(n13301) );
  NAND2X0 U13476 ( .IN1(n13303), .IN2(n13304), .QN(g33542) );
  NAND2X0 U13477 ( .IN1(n10508), .IN2(g1270), .QN(n13304) );
  NOR2X0 U13478 ( .IN1(n13305), .IN2(n13306), .QN(n13303) );
  NOR2X0 U13479 ( .IN1(n13307), .IN2(g1274), .QN(n13306) );
  NOR2X0 U13480 ( .IN1(n5730), .IN2(n13308), .QN(n13305) );
  NAND2X0 U13481 ( .IN1(n13309), .IN2(n13307), .QN(n13308) );
  NAND2X0 U13482 ( .IN1(n13310), .IN2(n13311), .QN(g33541) );
  NAND2X0 U13483 ( .IN1(n13312), .IN2(n13313), .QN(n13311) );
  NAND2X0 U13484 ( .IN1(n13314), .IN2(n13315), .QN(n13313) );
  NAND2X0 U13485 ( .IN1(n9764), .IN2(n13316), .QN(n13315) );
  INVX0 U13486 ( .INP(n13317), .ZN(n13314) );
  NOR2X0 U13487 ( .IN1(n9686), .IN2(n10459), .QN(n13312) );
  NAND2X0 U13488 ( .IN1(n13318), .IN2(g1030), .QN(n13310) );
  NAND2X0 U13489 ( .IN1(n13319), .IN2(n10402), .QN(n13318) );
  NAND2X0 U13490 ( .IN1(n13320), .IN2(n9686), .QN(n13319) );
  NOR2X0 U13491 ( .IN1(n13321), .IN2(n13317), .QN(n13320) );
  NAND2X0 U13492 ( .IN1(n13322), .IN2(n13323), .QN(g33540) );
  NAND2X0 U13493 ( .IN1(n10508), .IN2(g925), .QN(n13323) );
  NOR2X0 U13494 ( .IN1(n13324), .IN2(n13325), .QN(n13322) );
  NOR2X0 U13495 ( .IN1(n13326), .IN2(g930), .QN(n13325) );
  NOR2X0 U13496 ( .IN1(n5731), .IN2(n13327), .QN(n13324) );
  NAND2X0 U13497 ( .IN1(n13328), .IN2(n13326), .QN(n13327) );
  NAND2X0 U13498 ( .IN1(n13329), .IN2(n13330), .QN(g33539) );
  NAND2X0 U13499 ( .IN1(n10508), .IN2(g758), .QN(n13330) );
  NOR2X0 U13500 ( .IN1(n13331), .IN2(n13332), .QN(n13329) );
  NOR2X0 U13501 ( .IN1(g763), .IN2(n13333), .QN(n13332) );
  NOR2X0 U13502 ( .IN1(n5332), .IN2(n13334), .QN(n13331) );
  NAND2X0 U13503 ( .IN1(n2404), .IN2(n13333), .QN(n13334) );
  INVX0 U13504 ( .INP(n2980), .ZN(n13333) );
  NAND2X0 U13505 ( .IN1(n13335), .IN2(n13336), .QN(g33538) );
  NAND2X0 U13506 ( .IN1(n10508), .IN2(g590), .QN(n13336) );
  NOR2X0 U13507 ( .IN1(n13337), .IN2(n13338), .QN(n13335) );
  NOR2X0 U13508 ( .IN1(g595), .IN2(n13339), .QN(n13338) );
  NOR2X0 U13509 ( .IN1(n5476), .IN2(n13340), .QN(n13337) );
  NAND2X0 U13510 ( .IN1(n2421), .IN2(n13339), .QN(n13340) );
  INVX0 U13511 ( .INP(n2982), .ZN(n13339) );
  NAND2X0 U13512 ( .IN1(n13341), .IN2(n13342), .QN(g33537) );
  OR2X1 U13513 ( .IN1(n10310), .IN2(n10096), .Q(n13342) );
  NAND2X0 U13514 ( .IN1(n13343), .IN2(n10402), .QN(n13341) );
  NOR2X0 U13515 ( .IN1(n5724), .IN2(n11887), .QN(n13343) );
  INVX0 U13516 ( .INP(n2707), .ZN(n11887) );
  NOR2X0 U13517 ( .IN1(n5843), .IN2(n13344), .QN(g33536) );
  NOR2X0 U13518 ( .IN1(n2710), .IN2(n10459), .QN(n13344) );
  NAND2X0 U13519 ( .IN1(n13345), .IN2(n13346), .QN(g33535) );
  NAND2X0 U13520 ( .IN1(n10508), .IN2(g291), .QN(n13346) );
  NOR2X0 U13521 ( .IN1(n13347), .IN2(n13348), .QN(n13345) );
  NOR2X0 U13522 ( .IN1(g294), .IN2(n13349), .QN(n13348) );
  NOR2X0 U13523 ( .IN1(n5680), .IN2(n13350), .QN(n13347) );
  NAND2X0 U13524 ( .IN1(n10106), .IN2(n13349), .QN(n13350) );
  INVX0 U13525 ( .INP(n3276), .ZN(n13349) );
  NAND2X0 U13526 ( .IN1(n13351), .IN2(n13352), .QN(g33534) );
  NAND2X0 U13527 ( .IN1(n10508), .IN2(g150), .QN(n13352) );
  NOR2X0 U13528 ( .IN1(n13353), .IN2(n13354), .QN(n13351) );
  NOR2X0 U13529 ( .IN1(g153), .IN2(n13355), .QN(n13354) );
  NOR2X0 U13530 ( .IN1(n5677), .IN2(n13356), .QN(n13353) );
  NAND2X0 U13531 ( .IN1(n11894), .IN2(n13355), .QN(n13356) );
  INVX0 U13532 ( .INP(n3277), .ZN(n13355) );
  NOR2X0 U13533 ( .IN1(n13357), .IN2(n9715), .QN(g33533) );
  AND2X1 U13534 ( .IN1(n13358), .IN2(n5599), .Q(n13357) );
  NOR2X0 U13535 ( .IN1(n5363), .IN2(n13114), .QN(n13358) );
  NAND2X0 U13536 ( .IN1(n13359), .IN2(n13360), .QN(n13114) );
  NOR2X0 U13537 ( .IN1(n5320), .IN2(n13361), .QN(n13360) );
  OR2X1 U13538 ( .IN1(n9754), .IN2(test_so76), .Q(n13361) );
  NOR2X0 U13539 ( .IN1(g1205), .IN2(n13362), .QN(n13359) );
  NAND2X0 U13540 ( .IN1(n5442), .IN2(n10068), .QN(n13362) );
  NOR2X0 U13541 ( .IN1(n13363), .IN2(n13364), .QN(g33435) );
  NAND2X0 U13542 ( .IN1(n13365), .IN2(n13366), .QN(n13364) );
  NAND2X0 U13543 ( .IN1(n13367), .IN2(g2724), .QN(n13366) );
  NOR2X0 U13544 ( .IN1(n13368), .IN2(n13369), .QN(n13367) );
  NOR2X0 U13545 ( .IN1(g2729), .IN2(g2775), .QN(n13369) );
  NOR2X0 U13546 ( .IN1(n9780), .IN2(g2787), .QN(n13368) );
  NAND2X0 U13547 ( .IN1(n13370), .IN2(g2771), .QN(n13365) );
  NOR2X0 U13548 ( .IN1(n5403), .IN2(n11648), .QN(n13363) );
  NOR2X0 U13549 ( .IN1(n13371), .IN2(n13372), .QN(g33079) );
  NAND2X0 U13550 ( .IN1(n13373), .IN2(n13374), .QN(n13372) );
  NAND2X0 U13551 ( .IN1(n13375), .IN2(g2724), .QN(n13374) );
  NOR2X0 U13552 ( .IN1(n13376), .IN2(n13377), .QN(n13375) );
  NOR2X0 U13553 ( .IN1(g2729), .IN2(g2807), .QN(n13377) );
  NOR2X0 U13554 ( .IN1(n9780), .IN2(g2819), .QN(n13376) );
  NAND2X0 U13555 ( .IN1(n13370), .IN2(g2803), .QN(n13373) );
  NOR2X0 U13556 ( .IN1(n5404), .IN2(n11648), .QN(n13371) );
  NAND2X0 U13557 ( .IN1(n5301), .IN2(g2729), .QN(n11648) );
  NAND2X0 U13558 ( .IN1(n13378), .IN2(n13379), .QN(g33070) );
  NAND2X0 U13559 ( .IN1(n13380), .IN2(n13381), .QN(n13379) );
  NAND2X0 U13560 ( .IN1(n13382), .IN2(n13383), .QN(n13380) );
  NAND2X0 U13561 ( .IN1(n10369), .IN2(n13384), .QN(n13383) );
  NOR2X0 U13562 ( .IN1(n13385), .IN2(n13386), .QN(n13382) );
  AND2X1 U13563 ( .IN1(n5646), .IN2(g25756), .Q(n13386) );
  NAND2X0 U13564 ( .IN1(n10508), .IN2(g6565), .QN(n13378) );
  NAND2X0 U13565 ( .IN1(n13387), .IN2(n13388), .QN(g33069) );
  NAND2X0 U13566 ( .IN1(n13389), .IN2(g6561), .QN(n13388) );
  NAND2X0 U13567 ( .IN1(n13390), .IN2(n10402), .QN(n13389) );
  NAND2X0 U13568 ( .IN1(n5386), .IN2(n13381), .QN(n13390) );
  OR2X1 U13569 ( .IN1(n13391), .IN2(n5386), .Q(n13387) );
  NAND2X0 U13570 ( .IN1(n13392), .IN2(n13393), .QN(g33068) );
  NAND2X0 U13571 ( .IN1(n13394), .IN2(n5646), .QN(n13393) );
  NOR2X0 U13572 ( .IN1(n3404), .IN2(n13395), .QN(n13394) );
  NAND2X0 U13573 ( .IN1(n10508), .IN2(g6555), .QN(n13392) );
  NAND2X0 U13574 ( .IN1(n13396), .IN2(n13397), .QN(g33067) );
  NAND2X0 U13575 ( .IN1(n13398), .IN2(n13381), .QN(n13397) );
  NAND2X0 U13576 ( .IN1(n3407), .IN2(n13399), .QN(n13398) );
  NAND2X0 U13577 ( .IN1(n10369), .IN2(n13400), .QN(n13399) );
  NAND2X0 U13578 ( .IN1(n10508), .IN2(g6549), .QN(n13396) );
  NAND2X0 U13579 ( .IN1(n13401), .IN2(n13402), .QN(g33065) );
  NAND2X0 U13580 ( .IN1(n13403), .IN2(n13404), .QN(n13402) );
  NAND2X0 U13581 ( .IN1(n13405), .IN2(n13406), .QN(n13403) );
  NAND2X0 U13582 ( .IN1(n10369), .IN2(n13407), .QN(n13406) );
  NOR2X0 U13583 ( .IN1(n13408), .IN2(n13409), .QN(n13405) );
  AND2X1 U13584 ( .IN1(n5651), .IN2(g25742), .Q(n13409) );
  NAND2X0 U13585 ( .IN1(n10508), .IN2(g6219), .QN(n13401) );
  NAND2X0 U13586 ( .IN1(n13410), .IN2(n13411), .QN(g33064) );
  NAND2X0 U13587 ( .IN1(n13412), .IN2(g6215), .QN(n13411) );
  NAND2X0 U13588 ( .IN1(n13413), .IN2(n10402), .QN(n13412) );
  NAND2X0 U13589 ( .IN1(n5385), .IN2(n13404), .QN(n13413) );
  OR2X1 U13590 ( .IN1(n13414), .IN2(n5385), .Q(n13410) );
  NAND2X0 U13591 ( .IN1(n13415), .IN2(n13416), .QN(g33063) );
  NAND2X0 U13592 ( .IN1(n13417), .IN2(n5651), .QN(n13416) );
  NOR2X0 U13593 ( .IN1(n3414), .IN2(n13418), .QN(n13417) );
  NAND2X0 U13594 ( .IN1(n10508), .IN2(g6209), .QN(n13415) );
  NAND2X0 U13595 ( .IN1(n13419), .IN2(n13420), .QN(g33062) );
  NAND2X0 U13596 ( .IN1(n13421), .IN2(n13404), .QN(n13420) );
  NAND2X0 U13597 ( .IN1(n3417), .IN2(n13422), .QN(n13421) );
  NAND2X0 U13598 ( .IN1(n10369), .IN2(n13423), .QN(n13422) );
  NAND2X0 U13599 ( .IN1(n10510), .IN2(g6203), .QN(n13419) );
  NAND2X0 U13600 ( .IN1(n13424), .IN2(n13425), .QN(g33060) );
  NAND2X0 U13601 ( .IN1(n13426), .IN2(n13427), .QN(n13425) );
  NAND2X0 U13602 ( .IN1(n13428), .IN2(n13429), .QN(n13426) );
  NAND2X0 U13603 ( .IN1(n10369), .IN2(n13430), .QN(n13429) );
  NOR2X0 U13604 ( .IN1(n13431), .IN2(n13432), .QN(n13428) );
  AND2X1 U13605 ( .IN1(n5649), .IN2(g25728), .Q(n13432) );
  NAND2X0 U13606 ( .IN1(n10508), .IN2(g5873), .QN(n13424) );
  NAND2X0 U13607 ( .IN1(n13433), .IN2(n13434), .QN(g33059) );
  NAND2X0 U13608 ( .IN1(n13435), .IN2(g5869), .QN(n13434) );
  NAND2X0 U13609 ( .IN1(n13436), .IN2(n10402), .QN(n13435) );
  NAND2X0 U13610 ( .IN1(n5388), .IN2(n13427), .QN(n13436) );
  OR2X1 U13611 ( .IN1(n13437), .IN2(n5388), .Q(n13433) );
  NAND2X0 U13612 ( .IN1(n13438), .IN2(n13439), .QN(g33058) );
  NAND2X0 U13613 ( .IN1(n13440), .IN2(n5649), .QN(n13439) );
  NOR2X0 U13614 ( .IN1(n3424), .IN2(n13441), .QN(n13440) );
  NAND2X0 U13615 ( .IN1(n10508), .IN2(g5863), .QN(n13438) );
  NAND2X0 U13616 ( .IN1(n13442), .IN2(n13443), .QN(g33057) );
  NAND2X0 U13617 ( .IN1(n13444), .IN2(n13427), .QN(n13443) );
  NAND2X0 U13618 ( .IN1(n3427), .IN2(n13445), .QN(n13444) );
  NAND2X0 U13619 ( .IN1(n10370), .IN2(n13446), .QN(n13445) );
  NAND2X0 U13620 ( .IN1(n10507), .IN2(g5857), .QN(n13442) );
  NAND2X0 U13621 ( .IN1(n13447), .IN2(n13448), .QN(g33055) );
  NAND2X0 U13622 ( .IN1(n13449), .IN2(n13450), .QN(n13448) );
  NAND2X0 U13623 ( .IN1(n13451), .IN2(n13452), .QN(n13449) );
  NAND2X0 U13624 ( .IN1(n10370), .IN2(n13453), .QN(n13452) );
  NOR2X0 U13625 ( .IN1(n13454), .IN2(n13455), .QN(n13451) );
  AND2X1 U13626 ( .IN1(n5647), .IN2(g25714), .Q(n13455) );
  NAND2X0 U13627 ( .IN1(n10507), .IN2(g5527), .QN(n13447) );
  NAND2X0 U13628 ( .IN1(n13456), .IN2(n13457), .QN(g33054) );
  NAND2X0 U13629 ( .IN1(n13458), .IN2(g5523), .QN(n13457) );
  NAND2X0 U13630 ( .IN1(n13459), .IN2(n10402), .QN(n13458) );
  NAND2X0 U13631 ( .IN1(n5389), .IN2(n13450), .QN(n13459) );
  OR2X1 U13632 ( .IN1(n13460), .IN2(n5389), .Q(n13456) );
  NAND2X0 U13633 ( .IN1(n13461), .IN2(n13462), .QN(g33053) );
  NAND2X0 U13634 ( .IN1(n13463), .IN2(n5647), .QN(n13462) );
  NOR2X0 U13635 ( .IN1(n3434), .IN2(n13464), .QN(n13463) );
  NAND2X0 U13636 ( .IN1(n10507), .IN2(g5517), .QN(n13461) );
  NAND2X0 U13637 ( .IN1(n13465), .IN2(n13466), .QN(g33052) );
  NAND2X0 U13638 ( .IN1(n13467), .IN2(n13450), .QN(n13466) );
  NAND2X0 U13639 ( .IN1(n3437), .IN2(n13468), .QN(n13467) );
  NAND2X0 U13640 ( .IN1(n10370), .IN2(n13469), .QN(n13468) );
  NAND2X0 U13641 ( .IN1(n10507), .IN2(g5511), .QN(n13465) );
  NAND2X0 U13642 ( .IN1(n13470), .IN2(n13471), .QN(g33050) );
  NAND2X0 U13643 ( .IN1(n13472), .IN2(n13473), .QN(n13471) );
  NAND2X0 U13644 ( .IN1(n13474), .IN2(n13475), .QN(n13472) );
  NAND2X0 U13645 ( .IN1(n10370), .IN2(n13476), .QN(n13475) );
  NOR2X0 U13646 ( .IN1(n13477), .IN2(n13478), .QN(n13474) );
  AND2X1 U13647 ( .IN1(n5650), .IN2(g25700), .Q(n13478) );
  NAND2X0 U13648 ( .IN1(n10507), .IN2(g5180), .QN(n13470) );
  NAND2X0 U13649 ( .IN1(n13479), .IN2(n13480), .QN(g33049) );
  NAND2X0 U13650 ( .IN1(n13481), .IN2(g5176), .QN(n13480) );
  NAND2X0 U13651 ( .IN1(n13482), .IN2(n10402), .QN(n13481) );
  NAND2X0 U13652 ( .IN1(n5384), .IN2(n13473), .QN(n13482) );
  OR2X1 U13653 ( .IN1(n13483), .IN2(n5384), .Q(n13479) );
  NAND2X0 U13654 ( .IN1(n13484), .IN2(n13485), .QN(g33048) );
  NAND2X0 U13655 ( .IN1(n13486), .IN2(n5650), .QN(n13485) );
  NOR2X0 U13656 ( .IN1(n3444), .IN2(n13487), .QN(n13486) );
  NAND2X0 U13657 ( .IN1(n10507), .IN2(g5170), .QN(n13484) );
  NAND2X0 U13658 ( .IN1(n13488), .IN2(n13489), .QN(g33047) );
  NAND2X0 U13659 ( .IN1(n13490), .IN2(n13473), .QN(n13489) );
  NAND2X0 U13660 ( .IN1(n3447), .IN2(n13491), .QN(n13490) );
  NAND2X0 U13661 ( .IN1(n10370), .IN2(n13492), .QN(n13491) );
  NAND2X0 U13662 ( .IN1(n10507), .IN2(g5164), .QN(n13488) );
  NAND2X0 U13663 ( .IN1(n13493), .IN2(n13494), .QN(g33046) );
  NAND2X0 U13664 ( .IN1(n10507), .IN2(g5052), .QN(n13494) );
  NOR2X0 U13665 ( .IN1(n13495), .IN2(n13496), .QN(n13493) );
  NOR2X0 U13666 ( .IN1(n5615), .IN2(n13497), .QN(n13496) );
  OR2X1 U13667 ( .IN1(n13498), .IN2(n13499), .Q(n13497) );
  NOR2X0 U13668 ( .IN1(n13500), .IN2(g5057), .QN(n13495) );
  NOR2X0 U13669 ( .IN1(n13499), .IN2(n13501), .QN(n13500) );
  NOR2X0 U13670 ( .IN1(n13502), .IN2(n5607), .QN(n13499) );
  NAND2X0 U13671 ( .IN1(n13503), .IN2(n13504), .QN(g33045) );
  NAND2X0 U13672 ( .IN1(n12746), .IN2(g4567), .QN(n13504) );
  NOR2X0 U13673 ( .IN1(n13505), .IN2(n13506), .QN(n13503) );
  NAND2X0 U13674 ( .IN1(n13507), .IN2(n13508), .QN(g33044) );
  NAND2X0 U13675 ( .IN1(test_so93), .IN2(n12746), .QN(n13508) );
  NOR2X0 U13676 ( .IN1(n12017), .IN2(n13506), .QN(n13507) );
  NAND2X0 U13677 ( .IN1(n13509), .IN2(n13510), .QN(g33043) );
  NAND2X0 U13678 ( .IN1(test_so16), .IN2(n12746), .QN(n13510) );
  NOR2X0 U13679 ( .IN1(n13511), .IN2(n12747), .QN(n13509) );
  NAND2X0 U13680 ( .IN1(n13512), .IN2(n13513), .QN(g33042) );
  NAND2X0 U13681 ( .IN1(n12746), .IN2(g4540), .QN(n13513) );
  NOR2X0 U13682 ( .IN1(n13511), .IN2(n13506), .QN(n13512) );
  AND2X1 U13683 ( .IN1(n13514), .IN2(g4578), .Q(n13506) );
  NAND2X0 U13684 ( .IN1(n13515), .IN2(n13516), .QN(g33041) );
  NAND2X0 U13685 ( .IN1(test_so56), .IN2(n12746), .QN(n13516) );
  NOR2X0 U13686 ( .IN1(n13505), .IN2(n12747), .QN(n13515) );
  NAND2X0 U13687 ( .IN1(n13517), .IN2(n13518), .QN(g33040) );
  NAND2X0 U13688 ( .IN1(n12746), .IN2(g4504), .QN(n13518) );
  NOR2X0 U13689 ( .IN1(n12017), .IN2(n13519), .QN(n13517) );
  NOR2X0 U13690 ( .IN1(n12746), .IN2(n11849), .QN(n12017) );
  INVX0 U13691 ( .INP(n11184), .ZN(n11849) );
  NAND2X0 U13692 ( .IN1(n12573), .IN2(n12569), .QN(n11184) );
  NAND2X0 U13693 ( .IN1(n13520), .IN2(n13521), .QN(g33039) );
  NAND2X0 U13694 ( .IN1(n12746), .IN2(g4501), .QN(n13521) );
  NOR2X0 U13695 ( .IN1(n13505), .IN2(n12750), .QN(n13520) );
  NAND2X0 U13696 ( .IN1(n13522), .IN2(n13523), .QN(g33038) );
  NAND2X0 U13697 ( .IN1(n12746), .IN2(g4498), .QN(n13523) );
  NOR2X0 U13698 ( .IN1(n13505), .IN2(n13519), .QN(n13522) );
  AND2X1 U13699 ( .IN1(n13514), .IN2(n13524), .Q(n13505) );
  NAND2X0 U13700 ( .IN1(g72), .IN2(n12569), .QN(n13524) );
  INVX0 U13701 ( .INP(g73), .ZN(n12569) );
  NAND2X0 U13702 ( .IN1(n13525), .IN2(n13526), .QN(g33037) );
  NAND2X0 U13703 ( .IN1(n12746), .IN2(g4495), .QN(n13526) );
  NOR2X0 U13704 ( .IN1(n13511), .IN2(n12750), .QN(n13525) );
  NAND2X0 U13705 ( .IN1(n13527), .IN2(n13528), .QN(g33036) );
  NAND2X0 U13706 ( .IN1(n12746), .IN2(g4480), .QN(n13528) );
  NOR2X0 U13707 ( .IN1(n13511), .IN2(n13519), .QN(n13527) );
  NOR2X0 U13708 ( .IN1(n12746), .IN2(n9677), .QN(n13519) );
  AND2X1 U13709 ( .IN1(n13514), .IN2(n13529), .Q(n13511) );
  NAND2X0 U13710 ( .IN1(g73), .IN2(n12573), .QN(n13529) );
  INVX0 U13711 ( .INP(g72), .ZN(n12573) );
  NAND2X0 U13712 ( .IN1(n13530), .IN2(n13531), .QN(g33035) );
  NOR2X0 U13713 ( .IN1(n13532), .IN2(n13533), .QN(n13531) );
  NOR2X0 U13714 ( .IN1(n5350), .IN2(n10340), .QN(n13533) );
  NOR2X0 U13715 ( .IN1(n10494), .IN2(n13534), .QN(n13532) );
  NAND2X0 U13716 ( .IN1(n13535), .IN2(g4108), .QN(n13534) );
  NOR2X0 U13717 ( .IN1(n10114), .IN2(n13536), .QN(n13530) );
  NOR2X0 U13718 ( .IN1(g4108), .IN2(n13535), .QN(n13536) );
  INVX0 U13719 ( .INP(n10787), .ZN(n13535) );
  NOR2X0 U13720 ( .IN1(n13537), .IN2(n5350), .QN(n10787) );
  NAND2X0 U13721 ( .IN1(n13538), .IN2(n13539), .QN(g33034) );
  NAND2X0 U13722 ( .IN1(n13540), .IN2(n13541), .QN(n13539) );
  NAND2X0 U13723 ( .IN1(n13542), .IN2(n13543), .QN(n13540) );
  NAND2X0 U13724 ( .IN1(n10370), .IN2(n13544), .QN(n13543) );
  NOR2X0 U13725 ( .IN1(n13545), .IN2(n13546), .QN(n13542) );
  NOR2X0 U13726 ( .IN1(test_so33), .IN2(n13547), .QN(n13546) );
  NAND2X0 U13727 ( .IN1(n10507), .IN2(g3873), .QN(n13538) );
  NAND2X0 U13728 ( .IN1(n13548), .IN2(n13549), .QN(g33033) );
  NAND2X0 U13729 ( .IN1(test_so33), .IN2(n13550), .QN(n13549) );
  NAND2X0 U13730 ( .IN1(n13551), .IN2(n10403), .QN(n13550) );
  NAND2X0 U13731 ( .IN1(n5387), .IN2(n13541), .QN(n13551) );
  OR2X1 U13732 ( .IN1(n13552), .IN2(n5387), .Q(n13548) );
  NAND2X0 U13733 ( .IN1(n13553), .IN2(n13554), .QN(g33032) );
  NAND2X0 U13734 ( .IN1(n13555), .IN2(n13541), .QN(n13554) );
  NOR2X0 U13735 ( .IN1(test_so33), .IN2(n3479), .QN(n13555) );
  NAND2X0 U13736 ( .IN1(n10507), .IN2(g3863), .QN(n13553) );
  NAND2X0 U13737 ( .IN1(n13556), .IN2(n13557), .QN(g33031) );
  NAND2X0 U13738 ( .IN1(n13558), .IN2(n13541), .QN(n13557) );
  NAND2X0 U13739 ( .IN1(n3482), .IN2(n13559), .QN(n13558) );
  NAND2X0 U13740 ( .IN1(n10370), .IN2(n13560), .QN(n13559) );
  NAND2X0 U13741 ( .IN1(n10507), .IN2(g3857), .QN(n13556) );
  NAND2X0 U13742 ( .IN1(n13561), .IN2(n13562), .QN(g33029) );
  NAND2X0 U13743 ( .IN1(n13563), .IN2(n13564), .QN(n13562) );
  NAND2X0 U13744 ( .IN1(n13565), .IN2(n13566), .QN(n13563) );
  NAND2X0 U13745 ( .IN1(n10370), .IN2(n13567), .QN(n13566) );
  NOR2X0 U13746 ( .IN1(n13568), .IN2(n13569), .QN(n13565) );
  AND2X1 U13747 ( .IN1(n5645), .IN2(g25662), .Q(n13569) );
  NAND2X0 U13748 ( .IN1(n10507), .IN2(g3522), .QN(n13561) );
  NAND2X0 U13749 ( .IN1(n13570), .IN2(n13571), .QN(g33028) );
  NAND2X0 U13750 ( .IN1(n13572), .IN2(g3518), .QN(n13571) );
  NAND2X0 U13751 ( .IN1(n13573), .IN2(n10403), .QN(n13572) );
  NAND2X0 U13752 ( .IN1(n5383), .IN2(n13564), .QN(n13573) );
  OR2X1 U13753 ( .IN1(n13574), .IN2(n5383), .Q(n13570) );
  NAND2X0 U13754 ( .IN1(n13575), .IN2(n13576), .QN(g33027) );
  NAND2X0 U13755 ( .IN1(n13577), .IN2(n5645), .QN(n13576) );
  NOR2X0 U13756 ( .IN1(n3489), .IN2(n13578), .QN(n13577) );
  NAND2X0 U13757 ( .IN1(n10507), .IN2(g3512), .QN(n13575) );
  NAND2X0 U13758 ( .IN1(n13579), .IN2(n13580), .QN(g33026) );
  NAND2X0 U13759 ( .IN1(n13581), .IN2(n13564), .QN(n13580) );
  NAND2X0 U13760 ( .IN1(n3492), .IN2(n13582), .QN(n13581) );
  NAND2X0 U13761 ( .IN1(n10370), .IN2(n13583), .QN(n13582) );
  NAND2X0 U13762 ( .IN1(n10507), .IN2(g3506), .QN(n13579) );
  NAND2X0 U13763 ( .IN1(n13584), .IN2(n13585), .QN(g33024) );
  NAND2X0 U13764 ( .IN1(n10507), .IN2(g3171), .QN(n13585) );
  NOR2X0 U13765 ( .IN1(n13586), .IN2(n13587), .QN(n13584) );
  AND2X1 U13766 ( .IN1(n13588), .IN2(g25648), .Q(n13587) );
  NOR2X0 U13767 ( .IN1(n13589), .IN2(n13590), .QN(n13586) );
  NOR2X0 U13768 ( .IN1(n13591), .IN2(n13592), .QN(n13589) );
  NAND2X0 U13769 ( .IN1(n13593), .IN2(n13594), .QN(g33023) );
  NAND2X0 U13770 ( .IN1(n13595), .IN2(n13588), .QN(n13594) );
  NOR2X0 U13771 ( .IN1(n5603), .IN2(n10461), .QN(n13595) );
  NAND2X0 U13772 ( .IN1(n13596), .IN2(g3167), .QN(n13593) );
  NAND2X0 U13773 ( .IN1(n13597), .IN2(n10403), .QN(n13596) );
  NAND2X0 U13774 ( .IN1(n5603), .IN2(n13598), .QN(n13597) );
  NAND2X0 U13775 ( .IN1(n13599), .IN2(n13600), .QN(g33022) );
  NAND2X0 U13776 ( .IN1(n13588), .IN2(n13601), .QN(n13600) );
  INVX0 U13777 ( .INP(n13602), .ZN(n13588) );
  NAND2X0 U13778 ( .IN1(n10506), .IN2(g3161), .QN(n13599) );
  NAND2X0 U13779 ( .IN1(n13603), .IN2(n13604), .QN(g33021) );
  NAND2X0 U13780 ( .IN1(n10506), .IN2(g3155), .QN(n13604) );
  NOR2X0 U13781 ( .IN1(n13605), .IN2(n13606), .QN(n13603) );
  NOR2X0 U13782 ( .IN1(n3502), .IN2(n13590), .QN(n13606) );
  NAND2X0 U13783 ( .IN1(n13598), .IN2(n10403), .QN(n13590) );
  AND2X1 U13784 ( .IN1(n13607), .IN2(n13598), .Q(n13605) );
  NAND2X0 U13785 ( .IN1(n13608), .IN2(n13609), .QN(g33019) );
  NOR2X0 U13786 ( .IN1(n13610), .IN2(n13611), .QN(n13608) );
  NOR2X0 U13787 ( .IN1(n10494), .IN2(n13612), .QN(n13611) );
  XNOR2X1 U13788 ( .IN1(n2790), .IN2(test_so30), .Q(n13612) );
  NOR2X0 U13789 ( .IN1(n5516), .IN2(n10340), .QN(n13610) );
  NAND2X0 U13790 ( .IN1(n13613), .IN2(n13614), .QN(g33018) );
  NOR2X0 U13791 ( .IN1(n13615), .IN2(n13616), .QN(n13614) );
  NOR2X0 U13792 ( .IN1(g2610), .IN2(n13617), .QN(n13616) );
  NAND2X0 U13793 ( .IN1(n13618), .IN2(n13619), .QN(n13617) );
  NOR2X0 U13794 ( .IN1(n5508), .IN2(n13620), .QN(n13619) );
  AND2X1 U13795 ( .IN1(n3511), .IN2(n11591), .Q(n13618) );
  NOR2X0 U13796 ( .IN1(n10042), .IN2(n10340), .QN(n13615) );
  NOR2X0 U13797 ( .IN1(n13621), .IN2(n13622), .QN(n13613) );
  NOR2X0 U13798 ( .IN1(n13623), .IN2(n10140), .QN(n13622) );
  NOR2X0 U13799 ( .IN1(n13624), .IN2(n13625), .QN(n13623) );
  NAND2X0 U13800 ( .IN1(n13626), .IN2(n13184), .QN(n13625) );
  NOR2X0 U13801 ( .IN1(n10494), .IN2(n11905), .QN(n13624) );
  NOR2X0 U13802 ( .IN1(n13627), .IN2(n13628), .QN(n13621) );
  NAND2X0 U13803 ( .IN1(n3512), .IN2(n13629), .QN(n13628) );
  INVX0 U13804 ( .INP(n3513), .ZN(n13629) );
  NAND2X0 U13805 ( .IN1(n3524), .IN2(n11905), .QN(n3513) );
  INVX0 U13806 ( .INP(n3006), .ZN(n11905) );
  NAND2X0 U13807 ( .IN1(n3525), .IN2(n3505), .QN(n3006) );
  NAND2X0 U13808 ( .IN1(n13630), .IN2(n10042), .QN(n3512) );
  NOR2X0 U13809 ( .IN1(n9568), .IN2(n5508), .QN(n13630) );
  NAND2X0 U13810 ( .IN1(n13631), .IN2(n13632), .QN(g33017) );
  NOR2X0 U13811 ( .IN1(n3519), .IN2(n13633), .QN(n13632) );
  NOR2X0 U13812 ( .IN1(n5508), .IN2(n13626), .QN(n13633) );
  NOR2X0 U13813 ( .IN1(n13634), .IN2(n13635), .QN(n13631) );
  NOR2X0 U13814 ( .IN1(n10358), .IN2(n10140), .QN(n13635) );
  NOR2X0 U13815 ( .IN1(n10042), .IN2(n13627), .QN(n13634) );
  NAND2X0 U13816 ( .IN1(n13636), .IN2(n13637), .QN(g33016) );
  INVX0 U13817 ( .INP(n3519), .ZN(n13637) );
  NOR2X0 U13818 ( .IN1(n13638), .IN2(n13639), .QN(n13636) );
  NOR2X0 U13819 ( .IN1(n5372), .IN2(n13640), .QN(n13639) );
  NOR2X0 U13820 ( .IN1(n10042), .IN2(n13626), .QN(n13638) );
  NAND2X0 U13821 ( .IN1(n13641), .IN2(n13642), .QN(g33015) );
  NOR2X0 U13822 ( .IN1(n3519), .IN2(n13643), .QN(n13642) );
  NOR2X0 U13823 ( .IN1(n13627), .IN2(n13644), .QN(n13643) );
  NAND2X0 U13824 ( .IN1(n5508), .IN2(n13645), .QN(n13644) );
  NOR2X0 U13825 ( .IN1(n13646), .IN2(n13647), .QN(n13641) );
  AND2X1 U13826 ( .IN1(n10496), .IN2(test_so34), .Q(n13647) );
  NOR2X0 U13827 ( .IN1(n5372), .IN2(n13626), .QN(n13646) );
  NAND2X0 U13828 ( .IN1(n13648), .IN2(n13649), .QN(g33014) );
  NOR2X0 U13829 ( .IN1(n13650), .IN2(n13651), .QN(n13649) );
  NOR2X0 U13830 ( .IN1(g2476), .IN2(n13652), .QN(n13651) );
  NAND2X0 U13831 ( .IN1(n13653), .IN2(n13654), .QN(n13652) );
  NOR2X0 U13832 ( .IN1(n5509), .IN2(n13655), .QN(n13654) );
  AND2X1 U13833 ( .IN1(n3530), .IN2(n11591), .Q(n13653) );
  NOR2X0 U13834 ( .IN1(n10043), .IN2(n10341), .QN(n13650) );
  NOR2X0 U13835 ( .IN1(n13656), .IN2(n13657), .QN(n13648) );
  NOR2X0 U13836 ( .IN1(n5405), .IN2(n13658), .QN(n13657) );
  NOR2X0 U13837 ( .IN1(n13659), .IN2(n13660), .QN(n13658) );
  NAND2X0 U13838 ( .IN1(n13661), .IN2(n13184), .QN(n13660) );
  NOR2X0 U13839 ( .IN1(n10494), .IN2(n11904), .QN(n13659) );
  NOR2X0 U13840 ( .IN1(n13662), .IN2(n13663), .QN(n13656) );
  NAND2X0 U13841 ( .IN1(n3531), .IN2(n13664), .QN(n13663) );
  INVX0 U13842 ( .INP(n3532), .ZN(n13664) );
  NAND2X0 U13843 ( .IN1(n3524), .IN2(n11904), .QN(n3532) );
  INVX0 U13844 ( .INP(n3007), .ZN(n11904) );
  NAND2X0 U13845 ( .IN1(n13665), .IN2(n3525), .QN(n3007) );
  NOR2X0 U13846 ( .IN1(n5516), .IN2(g2741), .QN(n13665) );
  NAND2X0 U13847 ( .IN1(n13666), .IN2(n10043), .QN(n3531) );
  NOR2X0 U13848 ( .IN1(n9568), .IN2(n5509), .QN(n13666) );
  NAND2X0 U13849 ( .IN1(n13667), .IN2(n13668), .QN(g33013) );
  NOR2X0 U13850 ( .IN1(n3538), .IN2(n13669), .QN(n13668) );
  NOR2X0 U13851 ( .IN1(n5509), .IN2(n13661), .QN(n13669) );
  NOR2X0 U13852 ( .IN1(n13670), .IN2(n13671), .QN(n13667) );
  NOR2X0 U13853 ( .IN1(n5405), .IN2(n10341), .QN(n13671) );
  NOR2X0 U13854 ( .IN1(n10043), .IN2(n13662), .QN(n13670) );
  NAND2X0 U13855 ( .IN1(n13672), .IN2(n13673), .QN(g33012) );
  INVX0 U13856 ( .INP(n3538), .ZN(n13673) );
  NOR2X0 U13857 ( .IN1(n13674), .IN2(n13675), .QN(n13672) );
  NOR2X0 U13858 ( .IN1(n5373), .IN2(n13676), .QN(n13675) );
  NOR2X0 U13859 ( .IN1(n10043), .IN2(n13661), .QN(n13674) );
  NAND2X0 U13860 ( .IN1(n13677), .IN2(n13678), .QN(g33011) );
  NOR2X0 U13861 ( .IN1(n3538), .IN2(n13679), .QN(n13678) );
  NOR2X0 U13862 ( .IN1(n13662), .IN2(n13680), .QN(n13679) );
  NAND2X0 U13863 ( .IN1(n5509), .IN2(n13681), .QN(n13680) );
  NOR2X0 U13864 ( .IN1(n13682), .IN2(n13683), .QN(n13677) );
  NOR2X0 U13865 ( .IN1(n5840), .IN2(n10341), .QN(n13683) );
  NOR2X0 U13866 ( .IN1(n5373), .IN2(n13661), .QN(n13682) );
  NAND2X0 U13867 ( .IN1(n13684), .IN2(n13685), .QN(g33010) );
  NOR2X0 U13868 ( .IN1(n13686), .IN2(n13687), .QN(n13685) );
  NOR2X0 U13869 ( .IN1(test_so21), .IN2(n13688), .QN(n13687) );
  NAND2X0 U13870 ( .IN1(n13689), .IN2(n13690), .QN(n13688) );
  NOR2X0 U13871 ( .IN1(n5511), .IN2(n13691), .QN(n13690) );
  AND2X1 U13872 ( .IN1(n3548), .IN2(n11591), .Q(n13689) );
  NOR2X0 U13873 ( .IN1(n10357), .IN2(n10126), .QN(n13686) );
  NOR2X0 U13874 ( .IN1(n13692), .IN2(n13693), .QN(n13684) );
  NOR2X0 U13875 ( .IN1(n5276), .IN2(n13694), .QN(n13693) );
  NOR2X0 U13876 ( .IN1(n13695), .IN2(n13696), .QN(n13694) );
  NAND2X0 U13877 ( .IN1(n13697), .IN2(n13184), .QN(n13696) );
  NOR2X0 U13878 ( .IN1(n10493), .IN2(n11903), .QN(n13695) );
  NOR2X0 U13879 ( .IN1(n13698), .IN2(n13699), .QN(n13692) );
  NAND2X0 U13880 ( .IN1(n3549), .IN2(n13700), .QN(n13699) );
  INVX0 U13881 ( .INP(n3551), .ZN(n13700) );
  NAND2X0 U13882 ( .IN1(n3524), .IN2(n11903), .QN(n3551) );
  INVX0 U13883 ( .INP(n3550), .ZN(n11903) );
  NAND2X0 U13884 ( .IN1(n13701), .IN2(n3525), .QN(n3550) );
  NOR2X0 U13885 ( .IN1(n5349), .IN2(g2748), .QN(n13701) );
  NAND2X0 U13886 ( .IN1(n13702), .IN2(g2351), .QN(n3549) );
  NOR2X0 U13887 ( .IN1(test_so21), .IN2(n9568), .QN(n13702) );
  NAND2X0 U13888 ( .IN1(n13703), .IN2(n13704), .QN(g33009) );
  NOR2X0 U13889 ( .IN1(n3557), .IN2(n13705), .QN(n13704) );
  NOR2X0 U13890 ( .IN1(n5511), .IN2(n13697), .QN(n13705) );
  NOR2X0 U13891 ( .IN1(n13706), .IN2(n13707), .QN(n13703) );
  NOR2X0 U13892 ( .IN1(n5276), .IN2(n10341), .QN(n13707) );
  NOR2X0 U13893 ( .IN1(n10126), .IN2(n13698), .QN(n13706) );
  NAND2X0 U13894 ( .IN1(n13708), .IN2(n13709), .QN(g33008) );
  INVX0 U13895 ( .INP(n3557), .ZN(n13709) );
  NOR2X0 U13896 ( .IN1(n13710), .IN2(n13711), .QN(n13708) );
  NOR2X0 U13897 ( .IN1(n5375), .IN2(n13712), .QN(n13711) );
  NOR2X0 U13898 ( .IN1(n10126), .IN2(n13697), .QN(n13710) );
  NAND2X0 U13899 ( .IN1(n13713), .IN2(n13714), .QN(g33007) );
  NOR2X0 U13900 ( .IN1(n3557), .IN2(n13715), .QN(n13714) );
  NOR2X0 U13901 ( .IN1(n13698), .IN2(n13716), .QN(n13715) );
  NAND2X0 U13902 ( .IN1(n5511), .IN2(n13717), .QN(n13716) );
  NOR2X0 U13903 ( .IN1(n13718), .IN2(n13719), .QN(n13713) );
  NOR2X0 U13904 ( .IN1(n5841), .IN2(n10341), .QN(n13719) );
  NOR2X0 U13905 ( .IN1(n5375), .IN2(n13697), .QN(n13718) );
  NAND2X0 U13906 ( .IN1(n13720), .IN2(n13721), .QN(g33006) );
  NOR2X0 U13907 ( .IN1(n13722), .IN2(n13723), .QN(n13721) );
  NOR2X0 U13908 ( .IN1(g2208), .IN2(n13724), .QN(n13723) );
  NAND2X0 U13909 ( .IN1(n13725), .IN2(n13726), .QN(n13724) );
  NOR2X0 U13910 ( .IN1(n5512), .IN2(n13727), .QN(n13726) );
  AND2X1 U13911 ( .IN1(n3567), .IN2(n11591), .Q(n13725) );
  NOR2X0 U13912 ( .IN1(n10045), .IN2(n10341), .QN(n13722) );
  NOR2X0 U13913 ( .IN1(n13728), .IN2(n13729), .QN(n13720) );
  NOR2X0 U13914 ( .IN1(n5406), .IN2(n13730), .QN(n13729) );
  NOR2X0 U13915 ( .IN1(n13731), .IN2(n13732), .QN(n13730) );
  NAND2X0 U13916 ( .IN1(n13733), .IN2(n13184), .QN(n13732) );
  NOR2X0 U13917 ( .IN1(n10493), .IN2(n11902), .QN(n13731) );
  NOR2X0 U13918 ( .IN1(n13734), .IN2(n13735), .QN(n13728) );
  NAND2X0 U13919 ( .IN1(n3568), .IN2(n13736), .QN(n13735) );
  INVX0 U13920 ( .INP(n3570), .ZN(n13736) );
  NAND2X0 U13921 ( .IN1(n3524), .IN2(n11902), .QN(n3570) );
  INVX0 U13922 ( .INP(n3569), .ZN(n11902) );
  NAND2X0 U13923 ( .IN1(n13737), .IN2(n3525), .QN(n3569) );
  NOR2X0 U13924 ( .IN1(g2741), .IN2(g2748), .QN(n13737) );
  NAND2X0 U13925 ( .IN1(n13738), .IN2(n10045), .QN(n3568) );
  NOR2X0 U13926 ( .IN1(n9568), .IN2(n5512), .QN(n13738) );
  NAND2X0 U13927 ( .IN1(n13739), .IN2(n13740), .QN(g33005) );
  NOR2X0 U13928 ( .IN1(n3576), .IN2(n13741), .QN(n13740) );
  NOR2X0 U13929 ( .IN1(n5512), .IN2(n13733), .QN(n13741) );
  NOR2X0 U13930 ( .IN1(n13742), .IN2(n13743), .QN(n13739) );
  NOR2X0 U13931 ( .IN1(n5406), .IN2(n10341), .QN(n13743) );
  NOR2X0 U13932 ( .IN1(n10045), .IN2(n13734), .QN(n13742) );
  NAND2X0 U13933 ( .IN1(n13744), .IN2(n13745), .QN(g33004) );
  INVX0 U13934 ( .INP(n3576), .ZN(n13745) );
  NOR2X0 U13935 ( .IN1(n13746), .IN2(n13747), .QN(n13744) );
  NOR2X0 U13936 ( .IN1(n5376), .IN2(n13748), .QN(n13747) );
  NOR2X0 U13937 ( .IN1(n10045), .IN2(n13733), .QN(n13746) );
  NAND2X0 U13938 ( .IN1(n13749), .IN2(n13750), .QN(g33003) );
  NOR2X0 U13939 ( .IN1(n3576), .IN2(n13751), .QN(n13750) );
  NOR2X0 U13940 ( .IN1(n13734), .IN2(n13752), .QN(n13751) );
  NAND2X0 U13941 ( .IN1(n5512), .IN2(n13753), .QN(n13752) );
  NOR2X0 U13942 ( .IN1(n13754), .IN2(n13755), .QN(n13749) );
  NOR2X0 U13943 ( .IN1(n5839), .IN2(n10342), .QN(n13755) );
  NOR2X0 U13944 ( .IN1(n5376), .IN2(n13733), .QN(n13754) );
  NAND2X0 U13945 ( .IN1(n13756), .IN2(n13757), .QN(g33002) );
  NOR2X0 U13946 ( .IN1(n13758), .IN2(n13759), .QN(n13757) );
  NOR2X0 U13947 ( .IN1(g2051), .IN2(n13760), .QN(n13759) );
  NAND2X0 U13948 ( .IN1(n13761), .IN2(n13762), .QN(n13760) );
  NOR2X0 U13949 ( .IN1(n5507), .IN2(n13763), .QN(n13762) );
  AND2X1 U13950 ( .IN1(n3586), .IN2(n11591), .Q(n13761) );
  NOR2X0 U13951 ( .IN1(n10041), .IN2(n10342), .QN(n13758) );
  NOR2X0 U13952 ( .IN1(n13764), .IN2(n13765), .QN(n13756) );
  NOR2X0 U13953 ( .IN1(n5832), .IN2(n13766), .QN(n13765) );
  NOR2X0 U13954 ( .IN1(n13767), .IN2(n13768), .QN(n13766) );
  NAND2X0 U13955 ( .IN1(n13769), .IN2(n13184), .QN(n13768) );
  NOR2X0 U13956 ( .IN1(n10493), .IN2(n11910), .QN(n13767) );
  NOR2X0 U13957 ( .IN1(n13770), .IN2(n13771), .QN(n13764) );
  NAND2X0 U13958 ( .IN1(n3587), .IN2(n13772), .QN(n13771) );
  INVX0 U13959 ( .INP(n3589), .ZN(n13772) );
  NAND2X0 U13960 ( .IN1(n3524), .IN2(n11910), .QN(n3589) );
  INVX0 U13961 ( .INP(n3588), .ZN(n11910) );
  NAND2X0 U13962 ( .IN1(n13773), .IN2(n3505), .QN(n3588) );
  NOR2X0 U13963 ( .IN1(test_so30), .IN2(n13774), .QN(n13773) );
  NAND2X0 U13964 ( .IN1(n13775), .IN2(n10041), .QN(n3587) );
  NOR2X0 U13965 ( .IN1(n9568), .IN2(n5507), .QN(n13775) );
  NAND2X0 U13966 ( .IN1(n13776), .IN2(n13777), .QN(g33001) );
  NOR2X0 U13967 ( .IN1(n3595), .IN2(n13778), .QN(n13777) );
  NOR2X0 U13968 ( .IN1(n5507), .IN2(n13769), .QN(n13778) );
  NOR2X0 U13969 ( .IN1(n13779), .IN2(n13780), .QN(n13776) );
  NOR2X0 U13970 ( .IN1(n5832), .IN2(n10342), .QN(n13780) );
  NOR2X0 U13971 ( .IN1(n10041), .IN2(n13770), .QN(n13779) );
  NAND2X0 U13972 ( .IN1(n13781), .IN2(n13782), .QN(g33000) );
  INVX0 U13973 ( .INP(n3595), .ZN(n13782) );
  NOR2X0 U13974 ( .IN1(n13783), .IN2(n13784), .QN(n13781) );
  NOR2X0 U13975 ( .IN1(n5371), .IN2(n13785), .QN(n13784) );
  NOR2X0 U13976 ( .IN1(n10041), .IN2(n13769), .QN(n13783) );
  NAND2X0 U13977 ( .IN1(n13786), .IN2(n13787), .QN(g32999) );
  NOR2X0 U13978 ( .IN1(n3595), .IN2(n13788), .QN(n13787) );
  NOR2X0 U13979 ( .IN1(n13770), .IN2(n13789), .QN(n13788) );
  NAND2X0 U13980 ( .IN1(n5507), .IN2(n13790), .QN(n13789) );
  NOR2X0 U13981 ( .IN1(n13791), .IN2(n13792), .QN(n13786) );
  AND2X1 U13982 ( .IN1(n10496), .IN2(test_so59), .Q(n13792) );
  NOR2X0 U13983 ( .IN1(n5371), .IN2(n13769), .QN(n13791) );
  NAND2X0 U13984 ( .IN1(n13793), .IN2(n13794), .QN(g32998) );
  NOR2X0 U13985 ( .IN1(n13795), .IN2(n13796), .QN(n13794) );
  NOR2X0 U13986 ( .IN1(g1917), .IN2(n13797), .QN(n13796) );
  NAND2X0 U13987 ( .IN1(n13798), .IN2(n13799), .QN(n13797) );
  NOR2X0 U13988 ( .IN1(n5510), .IN2(n13800), .QN(n13799) );
  AND2X1 U13989 ( .IN1(n3604), .IN2(n11591), .Q(n13798) );
  NOR2X0 U13990 ( .IN1(n10044), .IN2(n10342), .QN(n13795) );
  NOR2X0 U13991 ( .IN1(n13801), .IN2(n13802), .QN(n13793) );
  NOR2X0 U13992 ( .IN1(n5829), .IN2(n13803), .QN(n13802) );
  NOR2X0 U13993 ( .IN1(n13804), .IN2(n13805), .QN(n13803) );
  NAND2X0 U13994 ( .IN1(n13806), .IN2(n13184), .QN(n13805) );
  NOR2X0 U13995 ( .IN1(n10493), .IN2(n11909), .QN(n13804) );
  NOR2X0 U13996 ( .IN1(n13807), .IN2(n13808), .QN(n13801) );
  NAND2X0 U13997 ( .IN1(n3605), .IN2(n13809), .QN(n13808) );
  INVX0 U13998 ( .INP(n3607), .ZN(n13809) );
  NAND2X0 U13999 ( .IN1(n3524), .IN2(n11909), .QN(n3607) );
  INVX0 U14000 ( .INP(n3606), .ZN(n11909) );
  NAND2X0 U14001 ( .IN1(n13810), .IN2(n13811), .QN(n3606) );
  NOR2X0 U14002 ( .IN1(test_so30), .IN2(n5516), .QN(n13811) );
  NOR2X0 U14003 ( .IN1(g2741), .IN2(n13774), .QN(n13810) );
  NAND2X0 U14004 ( .IN1(n13812), .IN2(n10044), .QN(n3605) );
  NOR2X0 U14005 ( .IN1(n9568), .IN2(n5510), .QN(n13812) );
  NAND2X0 U14006 ( .IN1(n13813), .IN2(n13814), .QN(g32997) );
  NOR2X0 U14007 ( .IN1(n3613), .IN2(n13815), .QN(n13814) );
  NOR2X0 U14008 ( .IN1(n5510), .IN2(n13806), .QN(n13815) );
  NOR2X0 U14009 ( .IN1(n13816), .IN2(n13817), .QN(n13813) );
  NOR2X0 U14010 ( .IN1(n5829), .IN2(n10342), .QN(n13817) );
  NOR2X0 U14011 ( .IN1(n10044), .IN2(n13807), .QN(n13816) );
  NAND2X0 U14012 ( .IN1(n13818), .IN2(n13819), .QN(g32996) );
  INVX0 U14013 ( .INP(n3613), .ZN(n13819) );
  NOR2X0 U14014 ( .IN1(n13820), .IN2(n13821), .QN(n13818) );
  NOR2X0 U14015 ( .IN1(n5374), .IN2(n13822), .QN(n13821) );
  NOR2X0 U14016 ( .IN1(n10044), .IN2(n13806), .QN(n13820) );
  NAND2X0 U14017 ( .IN1(n13823), .IN2(n13824), .QN(g32995) );
  NOR2X0 U14018 ( .IN1(n3613), .IN2(n13825), .QN(n13824) );
  NOR2X0 U14019 ( .IN1(n13807), .IN2(n13826), .QN(n13825) );
  NAND2X0 U14020 ( .IN1(n5510), .IN2(n13827), .QN(n13826) );
  NOR2X0 U14021 ( .IN1(n13828), .IN2(n13829), .QN(n13823) );
  NOR2X0 U14022 ( .IN1(n5837), .IN2(n10342), .QN(n13829) );
  NOR2X0 U14023 ( .IN1(n5374), .IN2(n13806), .QN(n13828) );
  NAND2X0 U14024 ( .IN1(n13830), .IN2(n13831), .QN(g32994) );
  NOR2X0 U14025 ( .IN1(n13832), .IN2(n13833), .QN(n13831) );
  NOR2X0 U14026 ( .IN1(g1783), .IN2(n13834), .QN(n13833) );
  NAND2X0 U14027 ( .IN1(n13835), .IN2(n13836), .QN(n13834) );
  NOR2X0 U14028 ( .IN1(n5359), .IN2(n13837), .QN(n13836) );
  AND2X1 U14029 ( .IN1(n3622), .IN2(n11591), .Q(n13835) );
  NOR2X0 U14030 ( .IN1(n5596), .IN2(n10342), .QN(n13832) );
  NOR2X0 U14031 ( .IN1(n13838), .IN2(n13839), .QN(n13830) );
  NOR2X0 U14032 ( .IN1(n5833), .IN2(n13840), .QN(n13839) );
  NOR2X0 U14033 ( .IN1(n13841), .IN2(n13842), .QN(n13840) );
  NAND2X0 U14034 ( .IN1(n13843), .IN2(n13184), .QN(n13842) );
  NOR2X0 U14035 ( .IN1(n3005), .IN2(n10461), .QN(n13841) );
  NOR2X0 U14036 ( .IN1(n13844), .IN2(n13845), .QN(n13838) );
  NAND2X0 U14037 ( .IN1(n3623), .IN2(n13846), .QN(n13845) );
  INVX0 U14038 ( .INP(n3624), .ZN(n13846) );
  NAND2X0 U14039 ( .IN1(n3524), .IN2(n3005), .QN(n3624) );
  NAND2X0 U14040 ( .IN1(n13847), .IN2(n5596), .QN(n3623) );
  NOR2X0 U14041 ( .IN1(n9568), .IN2(n5359), .QN(n13847) );
  NAND2X0 U14042 ( .IN1(n13848), .IN2(n13849), .QN(g32993) );
  NOR2X0 U14043 ( .IN1(n3630), .IN2(n13850), .QN(n13849) );
  NOR2X0 U14044 ( .IN1(n5359), .IN2(n13843), .QN(n13850) );
  NOR2X0 U14045 ( .IN1(n13851), .IN2(n13852), .QN(n13848) );
  NOR2X0 U14046 ( .IN1(n5833), .IN2(n10343), .QN(n13852) );
  NOR2X0 U14047 ( .IN1(n5596), .IN2(n13844), .QN(n13851) );
  NAND2X0 U14048 ( .IN1(n13853), .IN2(n13854), .QN(g32992) );
  INVX0 U14049 ( .INP(n3630), .ZN(n13854) );
  NOR2X0 U14050 ( .IN1(n13855), .IN2(n13856), .QN(n13853) );
  NOR2X0 U14051 ( .IN1(n5602), .IN2(n13857), .QN(n13856) );
  NOR2X0 U14052 ( .IN1(n5596), .IN2(n13843), .QN(n13855) );
  NAND2X0 U14053 ( .IN1(n13858), .IN2(n13859), .QN(g32991) );
  NOR2X0 U14054 ( .IN1(n3630), .IN2(n13860), .QN(n13859) );
  NOR2X0 U14055 ( .IN1(n13844), .IN2(n13861), .QN(n13860) );
  NAND2X0 U14056 ( .IN1(n5359), .IN2(n13862), .QN(n13861) );
  NOR2X0 U14057 ( .IN1(n13863), .IN2(n13864), .QN(n13858) );
  NOR2X0 U14058 ( .IN1(n5834), .IN2(n10343), .QN(n13864) );
  NOR2X0 U14059 ( .IN1(n5602), .IN2(n13843), .QN(n13863) );
  NAND2X0 U14060 ( .IN1(n13865), .IN2(n13866), .QN(g32990) );
  NOR2X0 U14061 ( .IN1(n13867), .IN2(n13868), .QN(n13866) );
  NOR2X0 U14062 ( .IN1(test_so94), .IN2(n13869), .QN(n13868) );
  NAND2X0 U14063 ( .IN1(n13870), .IN2(n13871), .QN(n13869) );
  NOR2X0 U14064 ( .IN1(n5525), .IN2(n13872), .QN(n13871) );
  AND2X1 U14065 ( .IN1(n3640), .IN2(n11591), .Q(n13870) );
  INVX0 U14066 ( .INP(n12838), .ZN(n11591) );
  NOR2X0 U14067 ( .IN1(n10358), .IN2(n10121), .QN(n13867) );
  NOR2X0 U14068 ( .IN1(n13873), .IN2(n13874), .QN(n13865) );
  NOR2X0 U14069 ( .IN1(n5407), .IN2(n13875), .QN(n13874) );
  NOR2X0 U14070 ( .IN1(n13876), .IN2(n13877), .QN(n13875) );
  NAND2X0 U14071 ( .IN1(n13878), .IN2(n13184), .QN(n13877) );
  NAND2X0 U14072 ( .IN1(n10371), .IN2(n1289), .QN(n13184) );
  INVX0 U14073 ( .INP(n2760), .ZN(n1289) );
  NOR2X0 U14074 ( .IN1(n10493), .IN2(n11908), .QN(n13876) );
  NOR2X0 U14075 ( .IN1(n13879), .IN2(n13880), .QN(n13873) );
  NAND2X0 U14076 ( .IN1(n3641), .IN2(n13881), .QN(n13880) );
  INVX0 U14077 ( .INP(n3642), .ZN(n13881) );
  NAND2X0 U14078 ( .IN1(n3524), .IN2(n11908), .QN(n3642) );
  INVX0 U14079 ( .INP(n3003), .ZN(n11908) );
  NAND2X0 U14080 ( .IN1(n549), .IN2(n572), .QN(n3003) );
  INVX0 U14081 ( .INP(n13774), .ZN(n572) );
  NAND2X0 U14082 ( .IN1(n13882), .IN2(n13883), .QN(n13774) );
  XOR2X1 U14083 ( .IN1(n9587), .IN2(g73), .Q(n13883) );
  XOR2X1 U14084 ( .IN1(n9582), .IN2(g72), .Q(n13882) );
  INVX0 U14085 ( .INP(n13884), .ZN(n549) );
  NAND2X0 U14086 ( .IN1(n13885), .IN2(g1657), .QN(n3641) );
  NOR2X0 U14087 ( .IN1(test_so94), .IN2(n9568), .QN(n13885) );
  NAND2X0 U14088 ( .IN1(n13886), .IN2(n13887), .QN(g32989) );
  NOR2X0 U14089 ( .IN1(n3648), .IN2(n13888), .QN(n13887) );
  NOR2X0 U14090 ( .IN1(n5525), .IN2(n13878), .QN(n13888) );
  NOR2X0 U14091 ( .IN1(n13889), .IN2(n13890), .QN(n13886) );
  NOR2X0 U14092 ( .IN1(n5407), .IN2(n10343), .QN(n13890) );
  NOR2X0 U14093 ( .IN1(n10121), .IN2(n13879), .QN(n13889) );
  NAND2X0 U14094 ( .IN1(n13891), .IN2(n13892), .QN(g32988) );
  INVX0 U14095 ( .INP(n3648), .ZN(n13892) );
  NOR2X0 U14096 ( .IN1(n13893), .IN2(n13894), .QN(n13891) );
  NOR2X0 U14097 ( .IN1(n5370), .IN2(n13895), .QN(n13894) );
  NOR2X0 U14098 ( .IN1(n10121), .IN2(n13878), .QN(n13893) );
  NAND2X0 U14099 ( .IN1(n13896), .IN2(n13897), .QN(g32987) );
  NOR2X0 U14100 ( .IN1(n3648), .IN2(n13898), .QN(n13897) );
  NOR2X0 U14101 ( .IN1(n13879), .IN2(n13899), .QN(n13898) );
  NAND2X0 U14102 ( .IN1(n5525), .IN2(n13900), .QN(n13899) );
  NOR2X0 U14103 ( .IN1(n13901), .IN2(n13902), .QN(n13896) );
  NOR2X0 U14104 ( .IN1(n5836), .IN2(n10343), .QN(n13902) );
  NOR2X0 U14105 ( .IN1(n5370), .IN2(n13878), .QN(n13901) );
  NAND2X0 U14106 ( .IN1(n13903), .IN2(n13904), .QN(g32986) );
  NAND2X0 U14107 ( .IN1(n13905), .IN2(n13906), .QN(n13904) );
  NOR2X0 U14108 ( .IN1(g1373), .IN2(n13298), .QN(n13905) );
  NOR2X0 U14109 ( .IN1(n13907), .IN2(n13908), .QN(n13903) );
  NOR2X0 U14110 ( .IN1(n9727), .IN2(n10343), .QN(n13908) );
  NOR2X0 U14111 ( .IN1(n10493), .IN2(n13909), .QN(n13907) );
  NAND2X0 U14112 ( .IN1(n13298), .IN2(g1373), .QN(n13909) );
  NAND2X0 U14113 ( .IN1(n3660), .IN2(n13910), .QN(n13298) );
  NAND2X0 U14114 ( .IN1(n9727), .IN2(n13297), .QN(n13910) );
  NOR2X0 U14115 ( .IN1(n5730), .IN2(n13911), .QN(g32985) );
  NOR2X0 U14116 ( .IN1(n10493), .IN2(n13912), .QN(n13911) );
  NOR2X0 U14117 ( .IN1(n13057), .IN2(n13307), .QN(n13912) );
  NAND2X0 U14118 ( .IN1(n3662), .IN2(g1270), .QN(n13307) );
  NAND2X0 U14119 ( .IN1(n13913), .IN2(n13914), .QN(g32984) );
  NAND2X0 U14120 ( .IN1(n10506), .IN2(g1263), .QN(n13914) );
  NOR2X0 U14121 ( .IN1(n13915), .IN2(n13916), .QN(n13913) );
  NOR2X0 U14122 ( .IN1(n13917), .IN2(g1270), .QN(n13916) );
  NOR2X0 U14123 ( .IN1(n5716), .IN2(n13918), .QN(n13915) );
  NAND2X0 U14124 ( .IN1(n13309), .IN2(n13917), .QN(n13918) );
  INVX0 U14125 ( .INP(n3662), .ZN(n13917) );
  NAND2X0 U14126 ( .IN1(n13919), .IN2(n13920), .QN(g32983) );
  NAND2X0 U14127 ( .IN1(n13921), .IN2(n13922), .QN(n13920) );
  NOR2X0 U14128 ( .IN1(g1030), .IN2(n13317), .QN(n13921) );
  NOR2X0 U14129 ( .IN1(n13923), .IN2(n13924), .QN(n13919) );
  NOR2X0 U14130 ( .IN1(n9728), .IN2(n10343), .QN(n13924) );
  NOR2X0 U14131 ( .IN1(n10493), .IN2(n13925), .QN(n13923) );
  NAND2X0 U14132 ( .IN1(n13317), .IN2(g1030), .QN(n13925) );
  NAND2X0 U14133 ( .IN1(n3669), .IN2(n13926), .QN(n13317) );
  NAND2X0 U14134 ( .IN1(n9728), .IN2(n13316), .QN(n13926) );
  NOR2X0 U14135 ( .IN1(n5731), .IN2(n13927), .QN(g32982) );
  NOR2X0 U14136 ( .IN1(n10493), .IN2(n13928), .QN(n13927) );
  NOR2X0 U14137 ( .IN1(n11355), .IN2(n13326), .QN(n13928) );
  NAND2X0 U14138 ( .IN1(n3671), .IN2(g925), .QN(n13326) );
  NAND2X0 U14139 ( .IN1(n13929), .IN2(n13930), .QN(g32981) );
  NAND2X0 U14140 ( .IN1(n10506), .IN2(g918), .QN(n13930) );
  NOR2X0 U14141 ( .IN1(n13931), .IN2(n13932), .QN(n13929) );
  NOR2X0 U14142 ( .IN1(n13933), .IN2(g925), .QN(n13932) );
  NOR2X0 U14143 ( .IN1(n5725), .IN2(n13934), .QN(n13931) );
  NAND2X0 U14144 ( .IN1(n13328), .IN2(n13933), .QN(n13934) );
  INVX0 U14145 ( .INP(n3671), .ZN(n13933) );
  NOR2X0 U14146 ( .IN1(n10493), .IN2(n13935), .QN(g32980) );
  NOR2X0 U14147 ( .IN1(n13936), .IN2(n11668), .QN(n13935) );
  NOR2X0 U14148 ( .IN1(n2644), .IN2(n13937), .QN(n11668) );
  AND2X1 U14149 ( .IN1(g854), .IN2(n13937), .Q(n13936) );
  NAND2X0 U14150 ( .IN1(n13938), .IN2(n13939), .QN(n13937) );
  NOR2X0 U14151 ( .IN1(n9787), .IN2(n9786), .QN(n13939) );
  NOR2X0 U14152 ( .IN1(n5633), .IN2(g385), .QN(n13938) );
  NAND2X0 U14153 ( .IN1(n13940), .IN2(n13941), .QN(g32979) );
  NAND2X0 U14154 ( .IN1(test_so2), .IN2(n10516), .QN(n13941) );
  NOR2X0 U14155 ( .IN1(n13942), .IN2(n13943), .QN(n13940) );
  NOR2X0 U14156 ( .IN1(g758), .IN2(n13944), .QN(n13943) );
  NOR2X0 U14157 ( .IN1(n5331), .IN2(n13945), .QN(n13942) );
  NAND2X0 U14158 ( .IN1(n2404), .IN2(n13944), .QN(n13945) );
  INVX0 U14159 ( .INP(n3272), .ZN(n13944) );
  NAND2X0 U14160 ( .IN1(n13946), .IN2(n13947), .QN(g32978) );
  NAND2X0 U14161 ( .IN1(n10506), .IN2(g582), .QN(n13947) );
  NOR2X0 U14162 ( .IN1(n13948), .IN2(n13949), .QN(n13946) );
  NOR2X0 U14163 ( .IN1(g590), .IN2(n13950), .QN(n13949) );
  NOR2X0 U14164 ( .IN1(n5472), .IN2(n13951), .QN(n13948) );
  NAND2X0 U14165 ( .IN1(n2421), .IN2(n13950), .QN(n13951) );
  INVX0 U14166 ( .INP(n3274), .ZN(n13950) );
  NAND2X0 U14167 ( .IN1(n13952), .IN2(n13953), .QN(g32977) );
  NAND2X0 U14168 ( .IN1(test_so51), .IN2(n10516), .QN(n13953) );
  NOR2X0 U14169 ( .IN1(n13954), .IN2(n13955), .QN(n13952) );
  NOR2X0 U14170 ( .IN1(g291), .IN2(n10780), .QN(n13955) );
  NOR2X0 U14171 ( .IN1(n5679), .IN2(n13956), .QN(n13954) );
  NAND2X0 U14172 ( .IN1(n10106), .IN2(n10780), .QN(n13956) );
  NAND2X0 U14173 ( .IN1(n13957), .IN2(test_so55), .QN(n10780) );
  NOR2X0 U14174 ( .IN1(n13958), .IN2(n10155), .QN(n13957) );
  NAND2X0 U14175 ( .IN1(n13959), .IN2(n13960), .QN(g32976) );
  NAND2X0 U14176 ( .IN1(n10506), .IN2(g164), .QN(n13960) );
  NOR2X0 U14177 ( .IN1(n13961), .IN2(n13962), .QN(n13959) );
  NOR2X0 U14178 ( .IN1(g150), .IN2(n13963), .QN(n13962) );
  NOR2X0 U14179 ( .IN1(n5676), .IN2(n13964), .QN(n13961) );
  NAND2X0 U14180 ( .IN1(n11894), .IN2(n13963), .QN(n13964) );
  INVX0 U14181 ( .INP(n3281), .ZN(n13963) );
  NOR2X0 U14182 ( .IN1(n13965), .IN2(n13966), .QN(g32185) );
  NAND2X0 U14183 ( .IN1(n13967), .IN2(n13968), .QN(n13966) );
  NAND2X0 U14184 ( .IN1(test_so22), .IN2(g2965), .QN(n13968) );
  NOR2X0 U14185 ( .IN1(n13969), .IN2(n13970), .QN(n13967) );
  NOR2X0 U14186 ( .IN1(n9733), .IN2(n10082), .QN(n13970) );
  NOR2X0 U14187 ( .IN1(n5750), .IN2(n10079), .QN(n13969) );
  NAND2X0 U14188 ( .IN1(n13971), .IN2(n13972), .QN(n13965) );
  NOR2X0 U14189 ( .IN1(n13973), .IN2(n13974), .QN(n13972) );
  NOR2X0 U14190 ( .IN1(n9729), .IN2(n10081), .QN(n13974) );
  NOR2X0 U14191 ( .IN1(n9730), .IN2(n10080), .QN(n13973) );
  NOR2X0 U14192 ( .IN1(n13975), .IN2(n13976), .QN(n13971) );
  NOR2X0 U14193 ( .IN1(n9731), .IN2(n10146), .QN(n13976) );
  NOR2X0 U14194 ( .IN1(n10084), .IN2(n10083), .QN(n13975) );
  NAND2X0 U14195 ( .IN1(n13977), .IN2(n13978), .QN(g31904) );
  NOR2X0 U14196 ( .IN1(n13979), .IN2(n13980), .QN(n13978) );
  AND2X1 U14197 ( .IN1(n13981), .IN2(n9752), .Q(n13980) );
  NOR2X0 U14198 ( .IN1(n9752), .IN2(n13982), .QN(n13979) );
  NAND2X0 U14199 ( .IN1(n13983), .IN2(n13984), .QN(n13982) );
  NOR2X0 U14200 ( .IN1(n13981), .IN2(n13985), .QN(n13983) );
  INVX0 U14201 ( .INP(n13986), .ZN(n13981) );
  NOR2X0 U14202 ( .IN1(n13987), .IN2(n13988), .QN(n13977) );
  NOR2X0 U14203 ( .IN1(n5601), .IN2(n10343), .QN(n13987) );
  NAND2X0 U14204 ( .IN1(n13989), .IN2(n13990), .QN(g31903) );
  NOR2X0 U14205 ( .IN1(n13991), .IN2(n13992), .QN(n13990) );
  NOR2X0 U14206 ( .IN1(g5052), .IN2(n13502), .QN(n13992) );
  NOR2X0 U14207 ( .IN1(n5607), .IN2(n13993), .QN(n13991) );
  NAND2X0 U14208 ( .IN1(n13994), .IN2(n13984), .QN(n13993) );
  AND2X1 U14209 ( .IN1(n13995), .IN2(n13502), .Q(n13994) );
  NAND2X0 U14210 ( .IN1(n13996), .IN2(g5046), .QN(n13502) );
  NOR2X0 U14211 ( .IN1(n13501), .IN2(n13997), .QN(n13989) );
  NOR2X0 U14212 ( .IN1(n5578), .IN2(n10344), .QN(n13997) );
  NOR2X0 U14213 ( .IN1(n13998), .IN2(n13995), .QN(n13501) );
  NAND2X0 U14214 ( .IN1(n10372), .IN2(n5607), .QN(n13998) );
  NAND2X0 U14215 ( .IN1(n13999), .IN2(n14000), .QN(g31902) );
  NAND2X0 U14216 ( .IN1(n13985), .IN2(n10404), .QN(n14000) );
  NOR2X0 U14217 ( .IN1(n14001), .IN2(n14002), .QN(n13999) );
  NOR2X0 U14218 ( .IN1(n5369), .IN2(n14003), .QN(n14002) );
  NOR2X0 U14219 ( .IN1(n10492), .IN2(n14004), .QN(n14003) );
  NOR2X0 U14220 ( .IN1(n9755), .IN2(g5029), .QN(n14004) );
  NOR2X0 U14221 ( .IN1(n14005), .IN2(n14006), .QN(n14001) );
  NAND2X0 U14222 ( .IN1(n13984), .IN2(g5029), .QN(n14006) );
  NAND2X0 U14223 ( .IN1(n14007), .IN2(n14008), .QN(n14005) );
  NAND2X0 U14224 ( .IN1(n5369), .IN2(g5022), .QN(n14008) );
  NAND2X0 U14225 ( .IN1(g5016), .IN2(g5062), .QN(n14007) );
  NAND2X0 U14226 ( .IN1(n14009), .IN2(n14010), .QN(g31901) );
  NOR2X0 U14227 ( .IN1(n14011), .IN2(n14012), .QN(n14010) );
  NOR2X0 U14228 ( .IN1(g5046), .IN2(n14013), .QN(n14012) );
  NOR2X0 U14229 ( .IN1(n5578), .IN2(n14014), .QN(n14011) );
  NAND2X0 U14230 ( .IN1(n14015), .IN2(n13984), .QN(n14014) );
  NOR2X0 U14231 ( .IN1(n13996), .IN2(n14016), .QN(n14015) );
  INVX0 U14232 ( .INP(n14013), .ZN(n13996) );
  NAND2X0 U14233 ( .IN1(n14017), .IN2(g5041), .QN(n14013) );
  NOR2X0 U14234 ( .IN1(n14018), .IN2(n14019), .QN(n14009) );
  NOR2X0 U14235 ( .IN1(n10492), .IN2(n13995), .QN(n14019) );
  NAND2X0 U14236 ( .IN1(n14016), .IN2(n5578), .QN(n13995) );
  AND2X1 U14237 ( .IN1(n14020), .IN2(n5611), .Q(n14016) );
  NOR2X0 U14238 ( .IN1(g5041), .IN2(n14021), .QN(n14020) );
  NOR2X0 U14239 ( .IN1(n5605), .IN2(n10344), .QN(n14018) );
  NAND2X0 U14240 ( .IN1(n14022), .IN2(n14023), .QN(g31900) );
  NAND2X0 U14241 ( .IN1(n5605), .IN2(n14024), .QN(n14023) );
  OR2X1 U14242 ( .IN1(n14017), .IN2(n14025), .Q(n14024) );
  NOR2X0 U14243 ( .IN1(n14026), .IN2(n14027), .QN(n14022) );
  NOR2X0 U14244 ( .IN1(n5611), .IN2(n10344), .QN(n14027) );
  NOR2X0 U14245 ( .IN1(n10492), .IN2(n14028), .QN(n14026) );
  NAND2X0 U14246 ( .IN1(n14029), .IN2(n14030), .QN(n14028) );
  NOR2X0 U14247 ( .IN1(n5605), .IN2(n14017), .QN(n14030) );
  NOR2X0 U14248 ( .IN1(n14031), .IN2(n5611), .QN(n14017) );
  NOR2X0 U14249 ( .IN1(n14032), .IN2(n14033), .QN(n14029) );
  NOR2X0 U14250 ( .IN1(n14021), .IN2(g5037), .QN(n14032) );
  NAND2X0 U14251 ( .IN1(n14034), .IN2(n14035), .QN(g31899) );
  NOR2X0 U14252 ( .IN1(n14036), .IN2(n14037), .QN(n14035) );
  NOR2X0 U14253 ( .IN1(n14031), .IN2(g5037), .QN(n14037) );
  NOR2X0 U14254 ( .IN1(n5611), .IN2(n14038), .QN(n14036) );
  NAND2X0 U14255 ( .IN1(n14039), .IN2(n13984), .QN(n14038) );
  AND2X1 U14256 ( .IN1(n14021), .IN2(n14031), .Q(n14039) );
  OR2X1 U14257 ( .IN1(n13986), .IN2(n9752), .Q(n14031) );
  NAND2X0 U14258 ( .IN1(n14040), .IN2(g5016), .QN(n13986) );
  NOR2X0 U14259 ( .IN1(n9755), .IN2(n5601), .QN(n14040) );
  NOR2X0 U14260 ( .IN1(n14025), .IN2(n14041), .QN(n14034) );
  NOR2X0 U14261 ( .IN1(n9752), .IN2(n10344), .QN(n14041) );
  AND2X1 U14262 ( .IN1(n13988), .IN2(n5611), .Q(n14025) );
  NOR2X0 U14263 ( .IN1(n10492), .IN2(n14021), .QN(n13988) );
  NAND2X0 U14264 ( .IN1(n9752), .IN2(n13985), .QN(n14021) );
  AND2X1 U14265 ( .IN1(n14042), .IN2(n5601), .Q(n13985) );
  NOR2X0 U14266 ( .IN1(n9784), .IN2(g5016), .QN(n14042) );
  NAND2X0 U14267 ( .IN1(n14043), .IN2(n14044), .QN(g31898) );
  NAND2X0 U14268 ( .IN1(n14045), .IN2(n5369), .QN(n14044) );
  NOR2X0 U14269 ( .IN1(n14046), .IN2(n13498), .QN(n14045) );
  INVX0 U14270 ( .INP(n13984), .ZN(n13498) );
  NOR2X0 U14271 ( .IN1(n14033), .IN2(n10463), .QN(n13984) );
  NAND2X0 U14272 ( .IN1(n14047), .IN2(n14048), .QN(n14033) );
  NOR2X0 U14273 ( .IN1(n14049), .IN2(n14050), .QN(n14048) );
  NOR2X0 U14274 ( .IN1(n14051), .IN2(n14052), .QN(n14047) );
  NOR2X0 U14275 ( .IN1(n14053), .IN2(n14054), .QN(n14043) );
  NOR2X0 U14276 ( .IN1(n9784), .IN2(n10344), .QN(n14054) );
  NOR2X0 U14277 ( .IN1(n10492), .IN2(n14055), .QN(n14053) );
  NAND2X0 U14278 ( .IN1(n14046), .IN2(g5016), .QN(n14055) );
  NOR2X0 U14279 ( .IN1(g5022), .IN2(g5062), .QN(n14046) );
  NAND2X0 U14280 ( .IN1(n14056), .IN2(n14057), .QN(g31897) );
  NOR2X0 U14281 ( .IN1(n12747), .IN2(n14058), .QN(n14056) );
  NOR2X0 U14282 ( .IN1(n9687), .IN2(n10344), .QN(n14058) );
  AND2X1 U14283 ( .IN1(n13514), .IN2(g4575), .Q(n12747) );
  NAND2X0 U14284 ( .IN1(n14059), .IN2(n14057), .QN(g31896) );
  AND2X1 U14285 ( .IN1(n14060), .IN2(n14061), .Q(n14057) );
  NAND2X0 U14286 ( .IN1(n13514), .IN2(n14062), .QN(n14061) );
  NAND2X0 U14287 ( .IN1(g72), .IN2(g73), .QN(n14062) );
  NAND2X0 U14288 ( .IN1(n14063), .IN2(g4372), .QN(n14060) );
  INVX0 U14289 ( .INP(n12753), .ZN(n14063) );
  NOR2X0 U14290 ( .IN1(n12750), .IN2(n14064), .QN(n14059) );
  NOR2X0 U14291 ( .IN1(n5849), .IN2(n10344), .QN(n14064) );
  NOR2X0 U14292 ( .IN1(n10150), .IN2(n12746), .QN(n12750) );
  INVX0 U14293 ( .INP(n13514), .ZN(n12746) );
  NOR2X0 U14294 ( .IN1(n10492), .IN2(n5670), .QN(n13514) );
  NAND2X0 U14295 ( .IN1(n12838), .IN2(n14065), .QN(g31895) );
  OR2X1 U14296 ( .IN1(n10309), .IN2(n5714), .Q(n14065) );
  NAND2X0 U14297 ( .IN1(n2760), .IN2(n10405), .QN(n12838) );
  NAND2X0 U14298 ( .IN1(n14066), .IN2(n14067), .QN(g31894) );
  NOR2X0 U14299 ( .IN1(n14068), .IN2(n14069), .QN(n14066) );
  NOR2X0 U14300 ( .IN1(n10492), .IN2(n14070), .QN(n14069) );
  XOR2X1 U14301 ( .IN1(g4098), .IN2(n13537), .Q(n14070) );
  OR2X1 U14302 ( .IN1(n3729), .IN2(n5340), .Q(n13537) );
  OR2X1 U14303 ( .IN1(n14071), .IN2(n5480), .Q(n3729) );
  NOR2X0 U14304 ( .IN1(n5340), .IN2(n10345), .QN(n14068) );
  NAND2X0 U14305 ( .IN1(n14072), .IN2(n14073), .QN(g31872) );
  NAND2X0 U14306 ( .IN1(n14074), .IN2(n3730), .QN(n14073) );
  XOR2X1 U14307 ( .IN1(g2748), .IN2(n14075), .Q(n14074) );
  NOR2X0 U14308 ( .IN1(n5349), .IN2(n3506), .QN(n14075) );
  NAND2X0 U14309 ( .IN1(n10506), .IN2(g2741), .QN(n14072) );
  NAND2X0 U14310 ( .IN1(n14076), .IN2(n14077), .QN(g31871) );
  NAND2X0 U14311 ( .IN1(n3733), .IN2(n13906), .QN(n14077) );
  NOR2X0 U14312 ( .IN1(n14078), .IN2(n14079), .QN(n14076) );
  NOR2X0 U14313 ( .IN1(n10492), .IN2(n14080), .QN(n14079) );
  OR2X1 U14314 ( .IN1(n3660), .IN2(n9727), .Q(n14080) );
  AND2X1 U14315 ( .IN1(n3734), .IN2(n14081), .Q(n3660) );
  NAND2X0 U14316 ( .IN1(n9761), .IN2(n13297), .QN(n14081) );
  NOR2X0 U14317 ( .IN1(n9761), .IN2(n10345), .QN(n14078) );
  NAND2X0 U14318 ( .IN1(n14082), .IN2(n14083), .QN(g31870) );
  NAND2X0 U14319 ( .IN1(n10506), .IN2(g1259), .QN(n14083) );
  NOR2X0 U14320 ( .IN1(n14084), .IN2(n14085), .QN(n14082) );
  NOR2X0 U14321 ( .IN1(g1263), .IN2(n14086), .QN(n14085) );
  NOR2X0 U14322 ( .IN1(n5674), .IN2(n14087), .QN(n14084) );
  NAND2X0 U14323 ( .IN1(n13309), .IN2(n14086), .QN(n14087) );
  INVX0 U14324 ( .INP(n3664), .ZN(n14086) );
  NAND2X0 U14325 ( .IN1(n14088), .IN2(n14089), .QN(g31869) );
  NAND2X0 U14326 ( .IN1(n3738), .IN2(n13922), .QN(n14089) );
  NOR2X0 U14327 ( .IN1(n14090), .IN2(n14091), .QN(n14088) );
  NOR2X0 U14328 ( .IN1(n10492), .IN2(n14092), .QN(n14091) );
  OR2X1 U14329 ( .IN1(n3669), .IN2(n9728), .Q(n14092) );
  AND2X1 U14330 ( .IN1(n3739), .IN2(n14093), .Q(n3669) );
  NAND2X0 U14331 ( .IN1(n9763), .IN2(n13316), .QN(n14093) );
  INVX0 U14332 ( .INP(n14094), .ZN(n3739) );
  NOR2X0 U14333 ( .IN1(n9763), .IN2(n10345), .QN(n14090) );
  NAND2X0 U14334 ( .IN1(n14095), .IN2(n14096), .QN(g31868) );
  NAND2X0 U14335 ( .IN1(n10506), .IN2(g914), .QN(n14096) );
  NOR2X0 U14336 ( .IN1(n14097), .IN2(n14098), .QN(n14095) );
  NOR2X0 U14337 ( .IN1(g918), .IN2(n14099), .QN(n14098) );
  NOR2X0 U14338 ( .IN1(n5673), .IN2(n14100), .QN(n14097) );
  NAND2X0 U14339 ( .IN1(n13328), .IN2(n14099), .QN(n14100) );
  INVX0 U14340 ( .INP(n3673), .ZN(n14099) );
  NAND2X0 U14341 ( .IN1(n14101), .IN2(n14102), .QN(g31867) );
  NAND2X0 U14342 ( .IN1(n10506), .IN2(g744), .QN(n14102) );
  NOR2X0 U14343 ( .IN1(n14103), .IN2(n14104), .QN(n14101) );
  NOR2X0 U14344 ( .IN1(test_so2), .IN2(n14105), .QN(n14104) );
  INVX0 U14345 ( .INP(n3682), .ZN(n14105) );
  NOR2X0 U14346 ( .IN1(n3682), .IN2(n14106), .QN(n14103) );
  NAND2X0 U14347 ( .IN1(n2404), .IN2(test_so2), .QN(n14106) );
  NAND2X0 U14348 ( .IN1(n14107), .IN2(n14108), .QN(g31866) );
  NAND2X0 U14349 ( .IN1(n10505), .IN2(g577), .QN(n14108) );
  NOR2X0 U14350 ( .IN1(n14109), .IN2(n14110), .QN(n14107) );
  NOR2X0 U14351 ( .IN1(g582), .IN2(n14111), .QN(n14110) );
  NOR2X0 U14352 ( .IN1(n5552), .IN2(n14112), .QN(n14109) );
  NAND2X0 U14353 ( .IN1(n2421), .IN2(n14111), .QN(n14112) );
  INVX0 U14354 ( .INP(n3684), .ZN(n14111) );
  NAND2X0 U14355 ( .IN1(n14113), .IN2(n14114), .QN(g31865) );
  NAND2X0 U14356 ( .IN1(test_so55), .IN2(n14115), .QN(n14114) );
  NAND2X0 U14357 ( .IN1(n14116), .IN2(n10405), .QN(n14115) );
  OR2X1 U14358 ( .IN1(n13958), .IN2(test_so51), .Q(n14116) );
  NAND2X0 U14359 ( .IN1(n14117), .IN2(n10154), .QN(n14113) );
  AND2X1 U14360 ( .IN1(test_so51), .IN2(n10106), .Q(n14117) );
  NAND2X0 U14361 ( .IN1(n14118), .IN2(n14119), .QN(g31864) );
  NAND2X0 U14362 ( .IN1(test_so73), .IN2(n10515), .QN(n14119) );
  NOR2X0 U14363 ( .IN1(n14120), .IN2(n14121), .QN(n14118) );
  NOR2X0 U14364 ( .IN1(g164), .IN2(n10765), .QN(n14121) );
  NOR2X0 U14365 ( .IN1(n5561), .IN2(n14122), .QN(n14120) );
  NAND2X0 U14366 ( .IN1(n11894), .IN2(n10765), .QN(n14122) );
  NAND2X0 U14367 ( .IN1(n14123), .IN2(test_so73), .QN(n10765) );
  NOR2X0 U14368 ( .IN1(n14124), .IN2(n14125), .QN(n14123) );
  NOR2X0 U14369 ( .IN1(g1636), .IN2(n5598), .QN(g31862) );
  NAND2X0 U14370 ( .IN1(n14126), .IN2(n14127), .QN(g31793) );
  NAND2X0 U14371 ( .IN1(n14128), .IN2(n14129), .QN(n14127) );
  NOR2X0 U14372 ( .IN1(n11300), .IN2(n14130), .QN(n14129) );
  NOR2X0 U14373 ( .IN1(n14131), .IN2(n11297), .QN(n14128) );
  NOR2X0 U14374 ( .IN1(n14132), .IN2(n14133), .QN(n14131) );
  NOR2X0 U14375 ( .IN1(n6007), .IN2(n14134), .QN(n14132) );
  NAND2X0 U14376 ( .IN1(n9769), .IN2(n14135), .QN(n14134) );
  NAND2X0 U14377 ( .IN1(n14136), .IN2(n14137), .QN(n14135) );
  NAND2X0 U14378 ( .IN1(n14138), .IN2(n14139), .QN(n14137) );
  INVX0 U14379 ( .INP(n14140), .ZN(n14139) );
  NAND2X0 U14380 ( .IN1(n14141), .IN2(n14142), .QN(n14138) );
  NAND2X0 U14381 ( .IN1(n9645), .IN2(n14143), .QN(n14142) );
  NAND2X0 U14382 ( .IN1(g5471), .IN2(g5817), .QN(n14143) );
  NAND2X0 U14383 ( .IN1(n9627), .IN2(n9618), .QN(n14141) );
  NAND2X0 U14384 ( .IN1(n11295), .IN2(n14144), .QN(n14126) );
  NOR2X0 U14385 ( .IN1(n14145), .IN2(n11299), .QN(n14144) );
  INVX0 U14386 ( .INP(n14133), .ZN(n11299) );
  NOR2X0 U14387 ( .IN1(n14136), .IN2(n14140), .QN(n14133) );
  AND2X1 U14388 ( .IN1(n14146), .IN2(n10365), .Q(n14136) );
  NAND2X0 U14389 ( .IN1(n14147), .IN2(n9645), .QN(n14146) );
  NOR2X0 U14390 ( .IN1(g5817), .IN2(g5471), .QN(n14147) );
  NOR2X0 U14391 ( .IN1(n14148), .IN2(n14149), .QN(n14145) );
  NOR2X0 U14392 ( .IN1(n11300), .IN2(n11297), .QN(n14149) );
  NOR2X0 U14393 ( .IN1(g6509), .IN2(n14150), .QN(n14148) );
  NAND2X0 U14394 ( .IN1(n14151), .IN2(n14152), .QN(n14150) );
  NAND2X0 U14395 ( .IN1(n14153), .IN2(g3466), .QN(n14152) );
  NAND2X0 U14396 ( .IN1(n11300), .IN2(n11297), .QN(n14151) );
  NAND2X0 U14397 ( .IN1(n14154), .IN2(n14155), .QN(n11297) );
  INVX0 U14398 ( .INP(n14153), .ZN(n14155) );
  NAND2X0 U14399 ( .IN1(n10373), .IN2(g3466), .QN(n14154) );
  NOR2X0 U14400 ( .IN1(g4427), .IN2(n6007), .QN(n11295) );
  NAND2X0 U14401 ( .IN1(g113), .IN2(g2868), .QN(g31665) );
  NAND2X0 U14402 ( .IN1(g113), .IN2(g2873), .QN(g31656) );
  NAND2X0 U14403 ( .IN1(n14156), .IN2(n14157), .QN(g30563) );
  NAND2X0 U14404 ( .IN1(n10505), .IN2(g6653), .QN(n14157) );
  NOR2X0 U14405 ( .IN1(n14158), .IN2(n14159), .QN(n14156) );
  NOR2X0 U14406 ( .IN1(n12631), .IN2(n14160), .QN(n14159) );
  NOR2X0 U14407 ( .IN1(n9799), .IN2(n14161), .QN(n14158) );
  NAND2X0 U14408 ( .IN1(n14162), .IN2(n14163), .QN(g30562) );
  NAND2X0 U14409 ( .IN1(n14164), .IN2(n3765), .QN(n14163) );
  NOR2X0 U14410 ( .IN1(n14165), .IN2(n14166), .QN(n14162) );
  NOR2X0 U14411 ( .IN1(n9994), .IN2(n10345), .QN(n14166) );
  NOR2X0 U14412 ( .IN1(n10474), .IN2(n14167), .QN(n14165) );
  OR2X1 U14413 ( .IN1(n14164), .IN2(n10023), .Q(n14167) );
  NOR2X0 U14414 ( .IN1(n3768), .IN2(n5646), .QN(n14164) );
  NAND2X0 U14415 ( .IN1(n14168), .IN2(n14169), .QN(g30561) );
  NAND2X0 U14416 ( .IN1(n13385), .IN2(n3765), .QN(n14169) );
  NOR2X0 U14417 ( .IN1(n14170), .IN2(n14171), .QN(n14168) );
  NOR2X0 U14418 ( .IN1(n9877), .IN2(n10345), .QN(n14171) );
  NOR2X0 U14419 ( .IN1(n10474), .IN2(n14172), .QN(n14170) );
  OR2X1 U14420 ( .IN1(n13385), .IN2(n9996), .Q(n14172) );
  NOR2X0 U14421 ( .IN1(n3770), .IN2(n5646), .QN(n13385) );
  NAND2X0 U14422 ( .IN1(n14173), .IN2(n14174), .QN(g30560) );
  NAND2X0 U14423 ( .IN1(n14175), .IN2(n3765), .QN(n14174) );
  NOR2X0 U14424 ( .IN1(n14176), .IN2(n14177), .QN(n14173) );
  NOR2X0 U14425 ( .IN1(n9800), .IN2(n10345), .QN(n14177) );
  NOR2X0 U14426 ( .IN1(n10474), .IN2(n14178), .QN(n14176) );
  OR2X1 U14427 ( .IN1(n14175), .IN2(n9960), .Q(n14178) );
  NOR2X0 U14428 ( .IN1(n3773), .IN2(n5646), .QN(n14175) );
  NAND2X0 U14429 ( .IN1(n14179), .IN2(n14180), .QN(g30559) );
  NAND2X0 U14430 ( .IN1(n3774), .IN2(n14181), .QN(n14180) );
  NOR2X0 U14431 ( .IN1(n14182), .IN2(n14183), .QN(n14179) );
  NOR2X0 U14432 ( .IN1(n10474), .IN2(n14184), .QN(n14183) );
  NAND2X0 U14433 ( .IN1(n14185), .IN2(g6653), .QN(n14184) );
  NAND2X0 U14434 ( .IN1(n14186), .IN2(n14181), .QN(n14185) );
  NOR2X0 U14435 ( .IN1(n9858), .IN2(n10345), .QN(n14182) );
  NAND2X0 U14436 ( .IN1(n14187), .IN2(n14188), .QN(g30558) );
  NAND2X0 U14437 ( .IN1(n3774), .IN2(n13384), .QN(n14188) );
  NOR2X0 U14438 ( .IN1(n14189), .IN2(n14190), .QN(n14187) );
  NOR2X0 U14439 ( .IN1(n10474), .IN2(n14191), .QN(n14190) );
  NAND2X0 U14440 ( .IN1(n14192), .IN2(g6649), .QN(n14191) );
  NAND2X0 U14441 ( .IN1(n14186), .IN2(n13384), .QN(n14192) );
  NOR2X0 U14442 ( .IN1(n9992), .IN2(n10346), .QN(n14189) );
  NAND2X0 U14443 ( .IN1(n14193), .IN2(n14194), .QN(g30557) );
  NAND2X0 U14444 ( .IN1(n3774), .IN2(n14195), .QN(n14194) );
  NOR2X0 U14445 ( .IN1(n14196), .IN2(n14197), .QN(n14193) );
  NOR2X0 U14446 ( .IN1(n10474), .IN2(n14198), .QN(n14197) );
  NAND2X0 U14447 ( .IN1(n14199), .IN2(g6645), .QN(n14198) );
  NAND2X0 U14448 ( .IN1(n14186), .IN2(n14195), .QN(n14199) );
  NOR2X0 U14449 ( .IN1(n9891), .IN2(n10346), .QN(n14196) );
  NAND2X0 U14450 ( .IN1(n14200), .IN2(n14201), .QN(g30556) );
  NAND2X0 U14451 ( .IN1(n3774), .IN2(n14202), .QN(n14201) );
  NOR2X0 U14452 ( .IN1(n14203), .IN2(n14204), .QN(n14200) );
  NOR2X0 U14453 ( .IN1(n10474), .IN2(n14205), .QN(n14204) );
  NAND2X0 U14454 ( .IN1(n14206), .IN2(g6641), .QN(n14205) );
  NAND2X0 U14455 ( .IN1(n14186), .IN2(n14202), .QN(n14206) );
  INVX0 U14456 ( .INP(n3404), .ZN(n14186) );
  NAND2X0 U14457 ( .IN1(g6549), .IN2(g6555), .QN(n3404) );
  NOR2X0 U14458 ( .IN1(n9947), .IN2(n10346), .QN(n14203) );
  NAND2X0 U14459 ( .IN1(n14207), .IN2(n14208), .QN(g30555) );
  NAND2X0 U14460 ( .IN1(n3780), .IN2(n14181), .QN(n14208) );
  NOR2X0 U14461 ( .IN1(n14209), .IN2(n14210), .QN(n14207) );
  NOR2X0 U14462 ( .IN1(n10474), .IN2(n14211), .QN(n14210) );
  NAND2X0 U14463 ( .IN1(n14212), .IN2(g6637), .QN(n14211) );
  NAND2X0 U14464 ( .IN1(n13400), .IN2(n14181), .QN(n14212) );
  NOR2X0 U14465 ( .IN1(n9859), .IN2(n10346), .QN(n14209) );
  NAND2X0 U14466 ( .IN1(n14213), .IN2(n14214), .QN(g30554) );
  NAND2X0 U14467 ( .IN1(n3780), .IN2(n13384), .QN(n14214) );
  NOR2X0 U14468 ( .IN1(n14215), .IN2(n14216), .QN(n14213) );
  NOR2X0 U14469 ( .IN1(n10474), .IN2(n14217), .QN(n14216) );
  NAND2X0 U14470 ( .IN1(n14218), .IN2(g6633), .QN(n14217) );
  NAND2X0 U14471 ( .IN1(n13400), .IN2(n13384), .QN(n14218) );
  NOR2X0 U14472 ( .IN1(n9933), .IN2(n10346), .QN(n14215) );
  NAND2X0 U14473 ( .IN1(n14219), .IN2(n14220), .QN(g30553) );
  NAND2X0 U14474 ( .IN1(n3780), .IN2(n14195), .QN(n14220) );
  NOR2X0 U14475 ( .IN1(n14221), .IN2(n14222), .QN(n14219) );
  NOR2X0 U14476 ( .IN1(n10474), .IN2(n14223), .QN(n14222) );
  NAND2X0 U14477 ( .IN1(n14224), .IN2(g6629), .QN(n14223) );
  NAND2X0 U14478 ( .IN1(n13400), .IN2(n14195), .QN(n14224) );
  NOR2X0 U14479 ( .IN1(n9840), .IN2(n10319), .QN(n14221) );
  NAND2X0 U14480 ( .IN1(n14225), .IN2(n14226), .QN(g30552) );
  NAND2X0 U14481 ( .IN1(n3780), .IN2(n14202), .QN(n14226) );
  NOR2X0 U14482 ( .IN1(n14227), .IN2(n14228), .QN(n14225) );
  NOR2X0 U14483 ( .IN1(n10473), .IN2(n14229), .QN(n14228) );
  NAND2X0 U14484 ( .IN1(n14230), .IN2(g6625), .QN(n14229) );
  NAND2X0 U14485 ( .IN1(n13400), .IN2(n14202), .QN(n14230) );
  INVX0 U14486 ( .INP(n3406), .ZN(n13400) );
  NAND2X0 U14487 ( .IN1(n5571), .IN2(g6555), .QN(n3406) );
  NOR2X0 U14488 ( .IN1(n9801), .IN2(n10312), .QN(n14227) );
  NAND2X0 U14489 ( .IN1(n14231), .IN2(n14232), .QN(g30551) );
  NAND2X0 U14490 ( .IN1(n3785), .IN2(n14181), .QN(n14232) );
  NOR2X0 U14491 ( .IN1(n14233), .IN2(n14234), .QN(n14231) );
  NOR2X0 U14492 ( .IN1(n10473), .IN2(n14235), .QN(n14234) );
  NAND2X0 U14493 ( .IN1(n14236), .IN2(g6621), .QN(n14235) );
  NAND2X0 U14494 ( .IN1(n14237), .IN2(n14181), .QN(n14236) );
  NOR2X0 U14495 ( .IN1(n9934), .IN2(n10314), .QN(n14233) );
  NAND2X0 U14496 ( .IN1(n14238), .IN2(n14239), .QN(g30550) );
  NAND2X0 U14497 ( .IN1(n3785), .IN2(n13384), .QN(n14239) );
  NOR2X0 U14498 ( .IN1(n14240), .IN2(n14241), .QN(n14238) );
  NOR2X0 U14499 ( .IN1(n10473), .IN2(n14242), .QN(n14241) );
  NAND2X0 U14500 ( .IN1(n14243), .IN2(g6617), .QN(n14242) );
  NAND2X0 U14501 ( .IN1(n14237), .IN2(n13384), .QN(n14243) );
  INVX0 U14502 ( .INP(n3768), .ZN(n13384) );
  NAND2X0 U14503 ( .IN1(n5386), .IN2(g6573), .QN(n3768) );
  NOR2X0 U14504 ( .IN1(n10025), .IN2(n10312), .QN(n14240) );
  NAND2X0 U14505 ( .IN1(n14244), .IN2(n14245), .QN(g30549) );
  NAND2X0 U14506 ( .IN1(n3785), .IN2(n14195), .QN(n14245) );
  NOR2X0 U14507 ( .IN1(n14246), .IN2(n14247), .QN(n14244) );
  NOR2X0 U14508 ( .IN1(n10473), .IN2(n14248), .QN(n14247) );
  NAND2X0 U14509 ( .IN1(n14249), .IN2(g6613), .QN(n14248) );
  NAND2X0 U14510 ( .IN1(n14237), .IN2(n14195), .QN(n14249) );
  INVX0 U14511 ( .INP(n3770), .ZN(n14195) );
  NAND2X0 U14512 ( .IN1(n5563), .IN2(g6565), .QN(n3770) );
  AND2X1 U14513 ( .IN1(n10497), .IN2(test_so71), .Q(n14246) );
  NAND2X0 U14514 ( .IN1(n14250), .IN2(n14251), .QN(g30548) );
  NAND2X0 U14515 ( .IN1(n3785), .IN2(n14202), .QN(n14251) );
  NOR2X0 U14516 ( .IN1(n14252), .IN2(n14253), .QN(n14250) );
  NOR2X0 U14517 ( .IN1(n10473), .IN2(n14254), .QN(n14253) );
  NAND2X0 U14518 ( .IN1(n14255), .IN2(g6609), .QN(n14254) );
  NAND2X0 U14519 ( .IN1(n14237), .IN2(n14202), .QN(n14255) );
  INVX0 U14520 ( .INP(n3773), .ZN(n14202) );
  NAND2X0 U14521 ( .IN1(n5563), .IN2(n5386), .QN(n3773) );
  INVX0 U14522 ( .INP(n3407), .ZN(n14237) );
  NAND2X0 U14523 ( .IN1(n10053), .IN2(g6549), .QN(n3407) );
  NOR2X0 U14524 ( .IN1(n9961), .IN2(n10312), .QN(n14252) );
  NAND2X0 U14525 ( .IN1(n14256), .IN2(n14257), .QN(g30547) );
  NAND2X0 U14526 ( .IN1(n10506), .IN2(g6605), .QN(n14257) );
  NOR2X0 U14527 ( .IN1(n14258), .IN2(n14259), .QN(n14256) );
  AND2X1 U14528 ( .IN1(n3765), .IN2(n3790), .Q(n14259) );
  NOR2X0 U14529 ( .IN1(n3790), .IN2(n14260), .QN(n14258) );
  NAND2X0 U14530 ( .IN1(n10375), .IN2(g6601), .QN(n14260) );
  NAND2X0 U14531 ( .IN1(n14261), .IN2(n14262), .QN(g30546) );
  OR2X1 U14532 ( .IN1(n10307), .IN2(n9996), .Q(n14262) );
  NOR2X0 U14533 ( .IN1(n14263), .IN2(n14264), .QN(n14261) );
  AND2X1 U14534 ( .IN1(n3765), .IN2(n3793), .Q(n14264) );
  NOR2X0 U14535 ( .IN1(n3793), .IN2(n14265), .QN(n14263) );
  NAND2X0 U14536 ( .IN1(n10375), .IN2(g6593), .QN(n14265) );
  NAND2X0 U14537 ( .IN1(n14266), .IN2(n14267), .QN(g30545) );
  NAND2X0 U14538 ( .IN1(n10506), .IN2(g6589), .QN(n14267) );
  NOR2X0 U14539 ( .IN1(n14268), .IN2(n14269), .QN(n14266) );
  AND2X1 U14540 ( .IN1(n3765), .IN2(n3795), .Q(n14269) );
  NOR2X0 U14541 ( .IN1(n3795), .IN2(n14270), .QN(n14268) );
  NAND2X0 U14542 ( .IN1(test_so71), .IN2(n10406), .QN(n14270) );
  NAND2X0 U14543 ( .IN1(n14271), .IN2(n14272), .QN(g30544) );
  NAND2X0 U14544 ( .IN1(n10506), .IN2(g6573), .QN(n14272) );
  NOR2X0 U14545 ( .IN1(n14273), .IN2(n14274), .QN(n14271) );
  AND2X1 U14546 ( .IN1(n3765), .IN2(n3797), .Q(n14274) );
  NOR2X0 U14547 ( .IN1(n3797), .IN2(n14275), .QN(n14273) );
  NAND2X0 U14548 ( .IN1(n10374), .IN2(g6581), .QN(n14275) );
  NOR2X0 U14549 ( .IN1(g6549), .IN2(n13391), .QN(g30543) );
  NAND2X0 U14550 ( .IN1(n14276), .IN2(n5646), .QN(n13391) );
  NOR2X0 U14551 ( .IN1(n10473), .IN2(n13395), .QN(n14276) );
  INVX0 U14552 ( .INP(n13381), .ZN(n13395) );
  NAND2X0 U14553 ( .IN1(n3799), .IN2(n11688), .QN(n13381) );
  NAND2X0 U14554 ( .IN1(n14277), .IN2(n14278), .QN(g30542) );
  NAND2X0 U14555 ( .IN1(n10506), .IN2(g6307), .QN(n14278) );
  NOR2X0 U14556 ( .IN1(n14279), .IN2(n14280), .QN(n14277) );
  NOR2X0 U14557 ( .IN1(n14160), .IN2(n12624), .QN(n14280) );
  NOR2X0 U14558 ( .IN1(n9806), .IN2(n14281), .QN(n14279) );
  NAND2X0 U14559 ( .IN1(n14282), .IN2(n14283), .QN(g30541) );
  NAND2X0 U14560 ( .IN1(n14284), .IN2(n3765), .QN(n14283) );
  NOR2X0 U14561 ( .IN1(n14285), .IN2(n14286), .QN(n14282) );
  NOR2X0 U14562 ( .IN1(n10004), .IN2(n10312), .QN(n14286) );
  NOR2X0 U14563 ( .IN1(n10473), .IN2(n14287), .QN(n14285) );
  OR2X1 U14564 ( .IN1(n14284), .IN2(n10031), .Q(n14287) );
  NOR2X0 U14565 ( .IN1(n3802), .IN2(n5651), .QN(n14284) );
  NAND2X0 U14566 ( .IN1(n14288), .IN2(n14289), .QN(g30540) );
  NAND2X0 U14567 ( .IN1(n13408), .IN2(n3765), .QN(n14289) );
  NOR2X0 U14568 ( .IN1(n14290), .IN2(n14291), .QN(n14288) );
  NOR2X0 U14569 ( .IN1(n9880), .IN2(n10312), .QN(n14291) );
  NOR2X0 U14570 ( .IN1(n10473), .IN2(n14292), .QN(n14290) );
  OR2X1 U14571 ( .IN1(n13408), .IN2(n10006), .Q(n14292) );
  NOR2X0 U14572 ( .IN1(n3804), .IN2(n5651), .QN(n13408) );
  NAND2X0 U14573 ( .IN1(n14293), .IN2(n14294), .QN(g30539) );
  NAND2X0 U14574 ( .IN1(n14295), .IN2(n3765), .QN(n14294) );
  NOR2X0 U14575 ( .IN1(n14296), .IN2(n14297), .QN(n14293) );
  NOR2X0 U14576 ( .IN1(n9807), .IN2(n10314), .QN(n14297) );
  NOR2X0 U14577 ( .IN1(n10473), .IN2(n14298), .QN(n14296) );
  OR2X1 U14578 ( .IN1(n14295), .IN2(n9964), .Q(n14298) );
  NOR2X0 U14579 ( .IN1(n3807), .IN2(n5651), .QN(n14295) );
  NAND2X0 U14580 ( .IN1(n14299), .IN2(n14300), .QN(g30538) );
  NAND2X0 U14581 ( .IN1(n3808), .IN2(n14301), .QN(n14300) );
  NOR2X0 U14582 ( .IN1(n14302), .IN2(n14303), .QN(n14299) );
  NOR2X0 U14583 ( .IN1(n10473), .IN2(n14304), .QN(n14303) );
  NAND2X0 U14584 ( .IN1(n14305), .IN2(g6307), .QN(n14304) );
  NAND2X0 U14585 ( .IN1(n14306), .IN2(n14301), .QN(n14305) );
  NOR2X0 U14586 ( .IN1(n9864), .IN2(n10316), .QN(n14302) );
  NAND2X0 U14587 ( .IN1(n14307), .IN2(n14308), .QN(g30537) );
  NAND2X0 U14588 ( .IN1(n3808), .IN2(n13407), .QN(n14308) );
  NOR2X0 U14589 ( .IN1(n14309), .IN2(n14310), .QN(n14307) );
  NOR2X0 U14590 ( .IN1(n10473), .IN2(n14311), .QN(n14310) );
  NAND2X0 U14591 ( .IN1(n14312), .IN2(g6303), .QN(n14311) );
  NAND2X0 U14592 ( .IN1(n14306), .IN2(n13407), .QN(n14312) );
  NOR2X0 U14593 ( .IN1(n10002), .IN2(n10312), .QN(n14309) );
  NAND2X0 U14594 ( .IN1(n14313), .IN2(n14314), .QN(g30536) );
  NAND2X0 U14595 ( .IN1(n3808), .IN2(n14315), .QN(n14314) );
  NOR2X0 U14596 ( .IN1(n14316), .IN2(n14317), .QN(n14313) );
  NOR2X0 U14597 ( .IN1(n10473), .IN2(n14318), .QN(n14317) );
  NAND2X0 U14598 ( .IN1(n14319), .IN2(g6299), .QN(n14318) );
  NAND2X0 U14599 ( .IN1(n14306), .IN2(n14315), .QN(n14319) );
  NOR2X0 U14600 ( .IN1(n9895), .IN2(n10312), .QN(n14316) );
  NAND2X0 U14601 ( .IN1(n14320), .IN2(n14321), .QN(g30535) );
  NAND2X0 U14602 ( .IN1(n3808), .IN2(n14322), .QN(n14321) );
  NOR2X0 U14603 ( .IN1(n14323), .IN2(n14324), .QN(n14320) );
  NOR2X0 U14604 ( .IN1(n10473), .IN2(n14325), .QN(n14324) );
  NAND2X0 U14605 ( .IN1(n14326), .IN2(g6295), .QN(n14325) );
  NAND2X0 U14606 ( .IN1(n14306), .IN2(n14322), .QN(n14326) );
  INVX0 U14607 ( .INP(n3414), .ZN(n14306) );
  NAND2X0 U14608 ( .IN1(g6203), .IN2(g6209), .QN(n3414) );
  NOR2X0 U14609 ( .IN1(n9949), .IN2(n10315), .QN(n14323) );
  NAND2X0 U14610 ( .IN1(n14327), .IN2(n14328), .QN(g30534) );
  NAND2X0 U14611 ( .IN1(n3814), .IN2(n14301), .QN(n14328) );
  NOR2X0 U14612 ( .IN1(n14329), .IN2(n14330), .QN(n14327) );
  NOR2X0 U14613 ( .IN1(n10473), .IN2(n14331), .QN(n14330) );
  NAND2X0 U14614 ( .IN1(n14332), .IN2(g6291), .QN(n14331) );
  NAND2X0 U14615 ( .IN1(n13423), .IN2(n14301), .QN(n14332) );
  NOR2X0 U14616 ( .IN1(n9865), .IN2(n10313), .QN(n14329) );
  NAND2X0 U14617 ( .IN1(n14333), .IN2(n14334), .QN(g30533) );
  NAND2X0 U14618 ( .IN1(n3814), .IN2(n13407), .QN(n14334) );
  NOR2X0 U14619 ( .IN1(n14335), .IN2(n14336), .QN(n14333) );
  NOR2X0 U14620 ( .IN1(n10472), .IN2(n14337), .QN(n14336) );
  NAND2X0 U14621 ( .IN1(n14338), .IN2(g6287), .QN(n14337) );
  NAND2X0 U14622 ( .IN1(n13423), .IN2(n13407), .QN(n14338) );
  NOR2X0 U14623 ( .IN1(n9939), .IN2(n10313), .QN(n14335) );
  NAND2X0 U14624 ( .IN1(n14339), .IN2(n14340), .QN(g30532) );
  NAND2X0 U14625 ( .IN1(n3814), .IN2(n14315), .QN(n14340) );
  NOR2X0 U14626 ( .IN1(n14341), .IN2(n14342), .QN(n14339) );
  NOR2X0 U14627 ( .IN1(n10472), .IN2(n14343), .QN(n14342) );
  NAND2X0 U14628 ( .IN1(n14344), .IN2(g6283), .QN(n14343) );
  NAND2X0 U14629 ( .IN1(n13423), .IN2(n14315), .QN(n14344) );
  NOR2X0 U14630 ( .IN1(n9842), .IN2(n10313), .QN(n14341) );
  NAND2X0 U14631 ( .IN1(n14345), .IN2(n14346), .QN(g30531) );
  NAND2X0 U14632 ( .IN1(n3814), .IN2(n14322), .QN(n14346) );
  NOR2X0 U14633 ( .IN1(n14347), .IN2(n14348), .QN(n14345) );
  NOR2X0 U14634 ( .IN1(n10472), .IN2(n14349), .QN(n14348) );
  NAND2X0 U14635 ( .IN1(n14350), .IN2(g6279), .QN(n14349) );
  NAND2X0 U14636 ( .IN1(n13423), .IN2(n14322), .QN(n14350) );
  INVX0 U14637 ( .INP(n3416), .ZN(n13423) );
  NAND2X0 U14638 ( .IN1(n5574), .IN2(g6209), .QN(n3416) );
  NOR2X0 U14639 ( .IN1(n9808), .IN2(n10315), .QN(n14347) );
  NAND2X0 U14640 ( .IN1(n14351), .IN2(n14352), .QN(g30530) );
  NAND2X0 U14641 ( .IN1(n3819), .IN2(n14301), .QN(n14352) );
  NOR2X0 U14642 ( .IN1(n14353), .IN2(n14354), .QN(n14351) );
  NOR2X0 U14643 ( .IN1(n10472), .IN2(n14355), .QN(n14354) );
  NAND2X0 U14644 ( .IN1(n14356), .IN2(g6275), .QN(n14355) );
  NAND2X0 U14645 ( .IN1(n14357), .IN2(n14301), .QN(n14356) );
  NOR2X0 U14646 ( .IN1(n9940), .IN2(n10313), .QN(n14353) );
  NAND2X0 U14647 ( .IN1(n14358), .IN2(n14359), .QN(g30529) );
  NAND2X0 U14648 ( .IN1(n3819), .IN2(n13407), .QN(n14359) );
  NOR2X0 U14649 ( .IN1(n14360), .IN2(n14361), .QN(n14358) );
  NOR2X0 U14650 ( .IN1(n10472), .IN2(n14362), .QN(n14361) );
  NAND2X0 U14651 ( .IN1(n14363), .IN2(g6271), .QN(n14362) );
  NAND2X0 U14652 ( .IN1(n14357), .IN2(n13407), .QN(n14363) );
  INVX0 U14653 ( .INP(n3802), .ZN(n13407) );
  NAND2X0 U14654 ( .IN1(n5385), .IN2(g6227), .QN(n3802) );
  NOR2X0 U14655 ( .IN1(n10033), .IN2(n10313), .QN(n14360) );
  NAND2X0 U14656 ( .IN1(n14364), .IN2(n14365), .QN(g30528) );
  NAND2X0 U14657 ( .IN1(n3819), .IN2(n14315), .QN(n14365) );
  NOR2X0 U14658 ( .IN1(n14366), .IN2(n14367), .QN(n14364) );
  NOR2X0 U14659 ( .IN1(n10472), .IN2(n14368), .QN(n14367) );
  NAND2X0 U14660 ( .IN1(n14369), .IN2(g6267), .QN(n14368) );
  NAND2X0 U14661 ( .IN1(n14357), .IN2(n14315), .QN(n14369) );
  INVX0 U14662 ( .INP(n3804), .ZN(n14315) );
  NAND2X0 U14663 ( .IN1(n5568), .IN2(g6219), .QN(n3804) );
  NOR2X0 U14664 ( .IN1(n9809), .IN2(n10314), .QN(n14366) );
  NAND2X0 U14665 ( .IN1(n14370), .IN2(n14371), .QN(g30527) );
  NAND2X0 U14666 ( .IN1(n3819), .IN2(n14322), .QN(n14371) );
  NOR2X0 U14667 ( .IN1(n14372), .IN2(n14373), .QN(n14370) );
  NOR2X0 U14668 ( .IN1(n10472), .IN2(n14374), .QN(n14373) );
  NAND2X0 U14669 ( .IN1(n14375), .IN2(g6263), .QN(n14374) );
  NAND2X0 U14670 ( .IN1(n14357), .IN2(n14322), .QN(n14375) );
  INVX0 U14671 ( .INP(n3807), .ZN(n14322) );
  NAND2X0 U14672 ( .IN1(n5568), .IN2(n5385), .QN(n3807) );
  INVX0 U14673 ( .INP(n3417), .ZN(n14357) );
  NAND2X0 U14674 ( .IN1(n10056), .IN2(g6203), .QN(n3417) );
  NOR2X0 U14675 ( .IN1(n9965), .IN2(n10313), .QN(n14372) );
  NAND2X0 U14676 ( .IN1(n14376), .IN2(n14377), .QN(g30526) );
  NAND2X0 U14677 ( .IN1(n10506), .IN2(g6259), .QN(n14377) );
  NOR2X0 U14678 ( .IN1(n14378), .IN2(n14379), .QN(n14376) );
  AND2X1 U14679 ( .IN1(n3765), .IN2(n3824), .Q(n14379) );
  NOR2X0 U14680 ( .IN1(n3824), .IN2(n14380), .QN(n14378) );
  NAND2X0 U14681 ( .IN1(n10377), .IN2(g6255), .QN(n14380) );
  NAND2X0 U14682 ( .IN1(n14381), .IN2(n14382), .QN(g30525) );
  NAND2X0 U14683 ( .IN1(n10506), .IN2(g6251), .QN(n14382) );
  NOR2X0 U14684 ( .IN1(n14383), .IN2(n14384), .QN(n14381) );
  AND2X1 U14685 ( .IN1(n3765), .IN2(n3827), .Q(n14384) );
  NOR2X0 U14686 ( .IN1(n3827), .IN2(n14385), .QN(n14383) );
  NAND2X0 U14687 ( .IN1(n10376), .IN2(g6247), .QN(n14385) );
  NAND2X0 U14688 ( .IN1(n14386), .IN2(n14387), .QN(g30524) );
  NAND2X0 U14689 ( .IN1(n10506), .IN2(g6243), .QN(n14387) );
  NOR2X0 U14690 ( .IN1(n14388), .IN2(n14389), .QN(n14386) );
  AND2X1 U14691 ( .IN1(n3765), .IN2(n3829), .Q(n14389) );
  NOR2X0 U14692 ( .IN1(n3829), .IN2(n14390), .QN(n14388) );
  NAND2X0 U14693 ( .IN1(n10377), .IN2(g6239), .QN(n14390) );
  NAND2X0 U14694 ( .IN1(n14391), .IN2(n14392), .QN(g30523) );
  NAND2X0 U14695 ( .IN1(n10506), .IN2(g6227), .QN(n14392) );
  NOR2X0 U14696 ( .IN1(n14393), .IN2(n14394), .QN(n14391) );
  AND2X1 U14697 ( .IN1(n3765), .IN2(n3831), .Q(n14394) );
  NOR2X0 U14698 ( .IN1(n3831), .IN2(n14395), .QN(n14393) );
  NAND2X0 U14699 ( .IN1(n10376), .IN2(g6235), .QN(n14395) );
  NOR2X0 U14700 ( .IN1(g6203), .IN2(n13414), .QN(g30522) );
  NAND2X0 U14701 ( .IN1(n14396), .IN2(n5651), .QN(n13414) );
  NOR2X0 U14702 ( .IN1(n10472), .IN2(n13418), .QN(n14396) );
  INVX0 U14703 ( .INP(n13404), .ZN(n13418) );
  NAND2X0 U14704 ( .IN1(n14397), .IN2(n3833), .QN(n13404) );
  NAND2X0 U14705 ( .IN1(n14398), .IN2(n14399), .QN(g30521) );
  NAND2X0 U14706 ( .IN1(n10506), .IN2(g5961), .QN(n14399) );
  NOR2X0 U14707 ( .IN1(n14400), .IN2(n14401), .QN(n14398) );
  NOR2X0 U14708 ( .IN1(n14160), .IN2(n12623), .QN(n14401) );
  AND2X1 U14709 ( .IN1(n14402), .IN2(test_so13), .Q(n14400) );
  NAND2X0 U14710 ( .IN1(n14403), .IN2(n14404), .QN(g30520) );
  NAND2X0 U14711 ( .IN1(n14405), .IN2(n3765), .QN(n14404) );
  NOR2X0 U14712 ( .IN1(n14406), .IN2(n14407), .QN(n14403) );
  NOR2X0 U14713 ( .IN1(n9980), .IN2(n10316), .QN(n14407) );
  NOR2X0 U14714 ( .IN1(n10472), .IN2(n14408), .QN(n14406) );
  OR2X1 U14715 ( .IN1(n14405), .IN2(n10011), .Q(n14408) );
  NOR2X0 U14716 ( .IN1(n3836), .IN2(n5649), .QN(n14405) );
  NAND2X0 U14717 ( .IN1(n14409), .IN2(n14410), .QN(g30519) );
  NAND2X0 U14718 ( .IN1(n13431), .IN2(n3765), .QN(n14410) );
  NOR2X0 U14719 ( .IN1(n14411), .IN2(n14412), .QN(n14409) );
  NOR2X0 U14720 ( .IN1(n9871), .IN2(n10314), .QN(n14412) );
  NOR2X0 U14721 ( .IN1(n10472), .IN2(n14413), .QN(n14411) );
  OR2X1 U14722 ( .IN1(n13431), .IN2(n9982), .Q(n14413) );
  NOR2X0 U14723 ( .IN1(n3838), .IN2(n5649), .QN(n13431) );
  NAND2X0 U14724 ( .IN1(n14414), .IN2(n14415), .QN(g30518) );
  NAND2X0 U14725 ( .IN1(n14416), .IN2(n3765), .QN(n14415) );
  NOR2X0 U14726 ( .IN1(n14417), .IN2(n14418), .QN(n14414) );
  NOR2X0 U14727 ( .IN1(n9814), .IN2(n10314), .QN(n14418) );
  NOR2X0 U14728 ( .IN1(n10472), .IN2(n14419), .QN(n14417) );
  OR2X1 U14729 ( .IN1(n14416), .IN2(n9955), .Q(n14419) );
  NOR2X0 U14730 ( .IN1(n3841), .IN2(n5649), .QN(n14416) );
  NAND2X0 U14731 ( .IN1(n14420), .IN2(n14421), .QN(g30517) );
  NAND2X0 U14732 ( .IN1(n3842), .IN2(n14422), .QN(n14421) );
  NOR2X0 U14733 ( .IN1(n14423), .IN2(n14424), .QN(n14420) );
  NOR2X0 U14734 ( .IN1(n10472), .IN2(n14425), .QN(n14424) );
  NAND2X0 U14735 ( .IN1(n14426), .IN2(g5961), .QN(n14425) );
  NAND2X0 U14736 ( .IN1(n14427), .IN2(n14422), .QN(n14426) );
  NOR2X0 U14737 ( .IN1(n9849), .IN2(n10314), .QN(n14423) );
  NAND2X0 U14738 ( .IN1(n14428), .IN2(n14429), .QN(g30516) );
  NAND2X0 U14739 ( .IN1(n3842), .IN2(n13430), .QN(n14429) );
  NOR2X0 U14740 ( .IN1(n14430), .IN2(n14431), .QN(n14428) );
  NOR2X0 U14741 ( .IN1(n10472), .IN2(n14432), .QN(n14431) );
  NAND2X0 U14742 ( .IN1(n14433), .IN2(g5957), .QN(n14432) );
  NAND2X0 U14743 ( .IN1(n14427), .IN2(n13430), .QN(n14433) );
  NOR2X0 U14744 ( .IN1(n9978), .IN2(n10315), .QN(n14430) );
  NAND2X0 U14745 ( .IN1(n14434), .IN2(n14435), .QN(g30515) );
  NAND2X0 U14746 ( .IN1(n3842), .IN2(n14436), .QN(n14435) );
  NOR2X0 U14747 ( .IN1(n14437), .IN2(n14438), .QN(n14434) );
  NOR2X0 U14748 ( .IN1(n10472), .IN2(n14439), .QN(n14438) );
  NAND2X0 U14749 ( .IN1(n14440), .IN2(g5953), .QN(n14439) );
  NAND2X0 U14750 ( .IN1(n14427), .IN2(n14436), .QN(n14440) );
  NOR2X0 U14751 ( .IN1(n9886), .IN2(n10316), .QN(n14437) );
  NAND2X0 U14752 ( .IN1(n14441), .IN2(n14442), .QN(g30514) );
  NAND2X0 U14753 ( .IN1(n3842), .IN2(n14443), .QN(n14442) );
  NOR2X0 U14754 ( .IN1(n14444), .IN2(n14445), .QN(n14441) );
  NOR2X0 U14755 ( .IN1(n10471), .IN2(n14446), .QN(n14445) );
  NAND2X0 U14756 ( .IN1(n14447), .IN2(g5949), .QN(n14446) );
  NAND2X0 U14757 ( .IN1(n14427), .IN2(n14443), .QN(n14447) );
  INVX0 U14758 ( .INP(n3424), .ZN(n14427) );
  NAND2X0 U14759 ( .IN1(g5857), .IN2(g5863), .QN(n3424) );
  NOR2X0 U14760 ( .IN1(n9944), .IN2(n10314), .QN(n14444) );
  NAND2X0 U14761 ( .IN1(n14448), .IN2(n14449), .QN(g30513) );
  NAND2X0 U14762 ( .IN1(n3848), .IN2(n14422), .QN(n14449) );
  NOR2X0 U14763 ( .IN1(n14450), .IN2(n14451), .QN(n14448) );
  NOR2X0 U14764 ( .IN1(n10471), .IN2(n14452), .QN(n14451) );
  NAND2X0 U14765 ( .IN1(n14453), .IN2(g5945), .QN(n14452) );
  NAND2X0 U14766 ( .IN1(n13446), .IN2(n14422), .QN(n14453) );
  NOR2X0 U14767 ( .IN1(n9850), .IN2(n10315), .QN(n14450) );
  NAND2X0 U14768 ( .IN1(n14454), .IN2(n14455), .QN(g30512) );
  NAND2X0 U14769 ( .IN1(n3848), .IN2(n13430), .QN(n14455) );
  NOR2X0 U14770 ( .IN1(n14456), .IN2(n14457), .QN(n14454) );
  NOR2X0 U14771 ( .IN1(n10471), .IN2(n14458), .QN(n14457) );
  NAND2X0 U14772 ( .IN1(n14459), .IN2(g5941), .QN(n14458) );
  NAND2X0 U14773 ( .IN1(n13446), .IN2(n13430), .QN(n14459) );
  NOR2X0 U14774 ( .IN1(n9924), .IN2(n10316), .QN(n14456) );
  NAND2X0 U14775 ( .IN1(n14460), .IN2(n14461), .QN(g30511) );
  NAND2X0 U14776 ( .IN1(n3848), .IN2(n14436), .QN(n14461) );
  NOR2X0 U14777 ( .IN1(n14462), .IN2(n14463), .QN(n14460) );
  NOR2X0 U14778 ( .IN1(n10471), .IN2(n14464), .QN(n14463) );
  NAND2X0 U14779 ( .IN1(n14465), .IN2(g5937), .QN(n14464) );
  NAND2X0 U14780 ( .IN1(n13446), .IN2(n14436), .QN(n14465) );
  NOR2X0 U14781 ( .IN1(n9837), .IN2(n10315), .QN(n14462) );
  NAND2X0 U14782 ( .IN1(n14466), .IN2(n14467), .QN(g30510) );
  NAND2X0 U14783 ( .IN1(n3848), .IN2(n14443), .QN(n14467) );
  NOR2X0 U14784 ( .IN1(n14468), .IN2(n14469), .QN(n14466) );
  NOR2X0 U14785 ( .IN1(n10471), .IN2(n14470), .QN(n14469) );
  NAND2X0 U14786 ( .IN1(n14471), .IN2(g5933), .QN(n14470) );
  NAND2X0 U14787 ( .IN1(n13446), .IN2(n14443), .QN(n14471) );
  INVX0 U14788 ( .INP(n3426), .ZN(n13446) );
  NAND2X0 U14789 ( .IN1(n5573), .IN2(g5863), .QN(n3426) );
  AND2X1 U14790 ( .IN1(n10496), .IN2(test_so28), .Q(n14468) );
  NAND2X0 U14791 ( .IN1(n14472), .IN2(n14473), .QN(g30509) );
  NAND2X0 U14792 ( .IN1(n3853), .IN2(n14422), .QN(n14473) );
  NOR2X0 U14793 ( .IN1(n14474), .IN2(n14475), .QN(n14472) );
  NOR2X0 U14794 ( .IN1(n10471), .IN2(n14476), .QN(n14475) );
  NAND2X0 U14795 ( .IN1(n14477), .IN2(g5929), .QN(n14476) );
  NAND2X0 U14796 ( .IN1(n14478), .IN2(n14422), .QN(n14477) );
  NOR2X0 U14797 ( .IN1(n9925), .IN2(n10315), .QN(n14474) );
  NAND2X0 U14798 ( .IN1(n14479), .IN2(n14480), .QN(g30508) );
  NAND2X0 U14799 ( .IN1(n3853), .IN2(n13430), .QN(n14480) );
  NOR2X0 U14800 ( .IN1(n14481), .IN2(n14482), .QN(n14479) );
  NOR2X0 U14801 ( .IN1(n10471), .IN2(n14483), .QN(n14482) );
  NAND2X0 U14802 ( .IN1(n14484), .IN2(g5925), .QN(n14483) );
  NAND2X0 U14803 ( .IN1(n14478), .IN2(n13430), .QN(n14484) );
  INVX0 U14804 ( .INP(n3836), .ZN(n13430) );
  NAND2X0 U14805 ( .IN1(n5388), .IN2(test_so36), .QN(n3836) );
  NOR2X0 U14806 ( .IN1(n10013), .IN2(n10317), .QN(n14481) );
  NAND2X0 U14807 ( .IN1(n14485), .IN2(n14486), .QN(g30507) );
  NAND2X0 U14808 ( .IN1(n3853), .IN2(n14436), .QN(n14486) );
  NOR2X0 U14809 ( .IN1(n14487), .IN2(n14488), .QN(n14485) );
  NOR2X0 U14810 ( .IN1(n10471), .IN2(n14489), .QN(n14488) );
  NAND2X0 U14811 ( .IN1(n14490), .IN2(g5921), .QN(n14489) );
  NAND2X0 U14812 ( .IN1(n14478), .IN2(n14436), .QN(n14490) );
  INVX0 U14813 ( .INP(n3838), .ZN(n14436) );
  NAND2X0 U14814 ( .IN1(n10139), .IN2(g5873), .QN(n3838) );
  NOR2X0 U14815 ( .IN1(n9815), .IN2(n10318), .QN(n14487) );
  NAND2X0 U14816 ( .IN1(n14491), .IN2(n14492), .QN(g30506) );
  NAND2X0 U14817 ( .IN1(n3853), .IN2(n14443), .QN(n14492) );
  NOR2X0 U14818 ( .IN1(n14493), .IN2(n14494), .QN(n14491) );
  NOR2X0 U14819 ( .IN1(n10471), .IN2(n14495), .QN(n14494) );
  NAND2X0 U14820 ( .IN1(test_so28), .IN2(n14496), .QN(n14495) );
  NAND2X0 U14821 ( .IN1(n14478), .IN2(n14443), .QN(n14496) );
  INVX0 U14822 ( .INP(n3841), .ZN(n14443) );
  NAND2X0 U14823 ( .IN1(n5388), .IN2(n10139), .QN(n3841) );
  INVX0 U14824 ( .INP(n3427), .ZN(n14478) );
  NAND2X0 U14825 ( .IN1(n10055), .IN2(g5857), .QN(n3427) );
  NOR2X0 U14826 ( .IN1(n9956), .IN2(n10315), .QN(n14493) );
  NAND2X0 U14827 ( .IN1(n14497), .IN2(n14498), .QN(g30505) );
  NAND2X0 U14828 ( .IN1(n10507), .IN2(g5913), .QN(n14498) );
  NOR2X0 U14829 ( .IN1(n14499), .IN2(n14500), .QN(n14497) );
  AND2X1 U14830 ( .IN1(n3765), .IN2(n3858), .Q(n14500) );
  NOR2X0 U14831 ( .IN1(n3858), .IN2(n14501), .QN(n14499) );
  NAND2X0 U14832 ( .IN1(n10377), .IN2(g5909), .QN(n14501) );
  NAND2X0 U14833 ( .IN1(n14502), .IN2(n14503), .QN(g30504) );
  NAND2X0 U14834 ( .IN1(n10507), .IN2(g5905), .QN(n14503) );
  NOR2X0 U14835 ( .IN1(n14504), .IN2(n14505), .QN(n14502) );
  AND2X1 U14836 ( .IN1(n3765), .IN2(n3861), .Q(n14505) );
  NOR2X0 U14837 ( .IN1(n3861), .IN2(n14506), .QN(n14504) );
  NAND2X0 U14838 ( .IN1(n10377), .IN2(g5901), .QN(n14506) );
  NAND2X0 U14839 ( .IN1(n14507), .IN2(n14508), .QN(g30503) );
  NAND2X0 U14840 ( .IN1(n10507), .IN2(g5897), .QN(n14508) );
  NOR2X0 U14841 ( .IN1(n14509), .IN2(n14510), .QN(n14507) );
  AND2X1 U14842 ( .IN1(n3765), .IN2(n3863), .Q(n14510) );
  NOR2X0 U14843 ( .IN1(n3863), .IN2(n14511), .QN(n14509) );
  NAND2X0 U14844 ( .IN1(n10376), .IN2(g5893), .QN(n14511) );
  NAND2X0 U14845 ( .IN1(n14512), .IN2(n14513), .QN(g30502) );
  NAND2X0 U14846 ( .IN1(test_so36), .IN2(n10515), .QN(n14513) );
  NOR2X0 U14847 ( .IN1(n14514), .IN2(n14515), .QN(n14512) );
  AND2X1 U14848 ( .IN1(n3765), .IN2(n3865), .Q(n14515) );
  NOR2X0 U14849 ( .IN1(n3865), .IN2(n14516), .QN(n14514) );
  NAND2X0 U14850 ( .IN1(n10377), .IN2(g5889), .QN(n14516) );
  NOR2X0 U14851 ( .IN1(g5857), .IN2(n13437), .QN(g30501) );
  NAND2X0 U14852 ( .IN1(n14517), .IN2(n5649), .QN(n13437) );
  NOR2X0 U14853 ( .IN1(n10471), .IN2(n13441), .QN(n14517) );
  INVX0 U14854 ( .INP(n13427), .ZN(n13441) );
  NAND2X0 U14855 ( .IN1(n14518), .IN2(n3833), .QN(n13427) );
  NAND2X0 U14856 ( .IN1(n14519), .IN2(n14520), .QN(g30500) );
  NAND2X0 U14857 ( .IN1(n10507), .IN2(g5615), .QN(n14520) );
  NOR2X0 U14858 ( .IN1(n14521), .IN2(n14522), .QN(n14519) );
  NOR2X0 U14859 ( .IN1(n14523), .IN2(n14160), .QN(n14522) );
  NOR2X0 U14860 ( .IN1(n9795), .IN2(n14524), .QN(n14521) );
  NAND2X0 U14861 ( .IN1(n14525), .IN2(n14526), .QN(g30499) );
  NAND2X0 U14862 ( .IN1(n14527), .IN2(n3765), .QN(n14526) );
  NOR2X0 U14863 ( .IN1(n14528), .IN2(n14529), .QN(n14525) );
  NOR2X0 U14864 ( .IN1(n9985), .IN2(n10316), .QN(n14529) );
  NOR2X0 U14865 ( .IN1(n10471), .IN2(n14530), .QN(n14528) );
  OR2X1 U14866 ( .IN1(n14527), .IN2(n10015), .Q(n14530) );
  NOR2X0 U14867 ( .IN1(n3869), .IN2(n5647), .QN(n14527) );
  NAND2X0 U14868 ( .IN1(n14531), .IN2(n14532), .QN(g30498) );
  NAND2X0 U14869 ( .IN1(n13454), .IN2(n3765), .QN(n14532) );
  INVX0 U14870 ( .INP(n14533), .ZN(n13454) );
  NOR2X0 U14871 ( .IN1(n14534), .IN2(n14535), .QN(n14531) );
  NOR2X0 U14872 ( .IN1(n9873), .IN2(n10317), .QN(n14535) );
  NOR2X0 U14873 ( .IN1(n10471), .IN2(n14536), .QN(n14534) );
  NAND2X0 U14874 ( .IN1(test_so6), .IN2(n14533), .QN(n14536) );
  NAND2X0 U14875 ( .IN1(n14537), .IN2(g5523), .QN(n14533) );
  NAND2X0 U14876 ( .IN1(n14538), .IN2(n14539), .QN(g30497) );
  NAND2X0 U14877 ( .IN1(n14540), .IN2(n3765), .QN(n14539) );
  NOR2X0 U14878 ( .IN1(n14541), .IN2(n14542), .QN(n14538) );
  NOR2X0 U14879 ( .IN1(n9796), .IN2(n10316), .QN(n14542) );
  NOR2X0 U14880 ( .IN1(n10471), .IN2(n14543), .QN(n14541) );
  OR2X1 U14881 ( .IN1(n14540), .IN2(n9957), .Q(n14543) );
  NOR2X0 U14882 ( .IN1(n3874), .IN2(n5647), .QN(n14540) );
  NAND2X0 U14883 ( .IN1(n14544), .IN2(n14545), .QN(g30496) );
  NAND2X0 U14884 ( .IN1(n3875), .IN2(n14546), .QN(n14545) );
  NOR2X0 U14885 ( .IN1(n14547), .IN2(n14548), .QN(n14544) );
  NOR2X0 U14886 ( .IN1(n10471), .IN2(n14549), .QN(n14548) );
  NAND2X0 U14887 ( .IN1(n14550), .IN2(g5615), .QN(n14549) );
  NAND2X0 U14888 ( .IN1(n14551), .IN2(n14546), .QN(n14550) );
  NOR2X0 U14889 ( .IN1(n9852), .IN2(n10317), .QN(n14547) );
  NAND2X0 U14890 ( .IN1(n14552), .IN2(n14553), .QN(g30495) );
  NAND2X0 U14891 ( .IN1(n3875), .IN2(n13453), .QN(n14553) );
  NOR2X0 U14892 ( .IN1(n14554), .IN2(n14555), .QN(n14552) );
  NOR2X0 U14893 ( .IN1(n10470), .IN2(n14556), .QN(n14555) );
  NAND2X0 U14894 ( .IN1(n14557), .IN2(g5611), .QN(n14556) );
  NAND2X0 U14895 ( .IN1(n14551), .IN2(n13453), .QN(n14557) );
  NOR2X0 U14896 ( .IN1(n9983), .IN2(n10316), .QN(n14554) );
  NAND2X0 U14897 ( .IN1(n14558), .IN2(n14559), .QN(g30494) );
  NAND2X0 U14898 ( .IN1(n3875), .IN2(n14537), .QN(n14559) );
  NOR2X0 U14899 ( .IN1(n14560), .IN2(n14561), .QN(n14558) );
  NOR2X0 U14900 ( .IN1(n10470), .IN2(n14562), .QN(n14561) );
  NAND2X0 U14901 ( .IN1(n14563), .IN2(g5607), .QN(n14562) );
  NAND2X0 U14902 ( .IN1(n14551), .IN2(n14537), .QN(n14563) );
  NOR2X0 U14903 ( .IN1(n10357), .IN2(n10147), .QN(n14560) );
  NAND2X0 U14904 ( .IN1(n14564), .IN2(n14565), .QN(g30493) );
  NAND2X0 U14905 ( .IN1(n3875), .IN2(n14566), .QN(n14565) );
  NOR2X0 U14906 ( .IN1(n14567), .IN2(n14568), .QN(n14564) );
  NOR2X0 U14907 ( .IN1(n10470), .IN2(n14569), .QN(n14568) );
  NAND2X0 U14908 ( .IN1(n14570), .IN2(g5603), .QN(n14569) );
  NAND2X0 U14909 ( .IN1(n14551), .IN2(n14566), .QN(n14570) );
  INVX0 U14910 ( .INP(n3434), .ZN(n14551) );
  NAND2X0 U14911 ( .IN1(g5511), .IN2(g5517), .QN(n3434) );
  NOR2X0 U14912 ( .IN1(n9945), .IN2(n10317), .QN(n14567) );
  NAND2X0 U14913 ( .IN1(n14571), .IN2(n14572), .QN(g30492) );
  NAND2X0 U14914 ( .IN1(n3881), .IN2(n14546), .QN(n14572) );
  NOR2X0 U14915 ( .IN1(n14573), .IN2(n14574), .QN(n14571) );
  NOR2X0 U14916 ( .IN1(n10470), .IN2(n14575), .QN(n14574) );
  NAND2X0 U14917 ( .IN1(n14576), .IN2(g5599), .QN(n14575) );
  NAND2X0 U14918 ( .IN1(n13469), .IN2(n14546), .QN(n14576) );
  NOR2X0 U14919 ( .IN1(n9853), .IN2(n10317), .QN(n14573) );
  NAND2X0 U14920 ( .IN1(n14577), .IN2(n14578), .QN(g30491) );
  NAND2X0 U14921 ( .IN1(n3881), .IN2(n13453), .QN(n14578) );
  NOR2X0 U14922 ( .IN1(n14579), .IN2(n14580), .QN(n14577) );
  NOR2X0 U14923 ( .IN1(n10470), .IN2(n14581), .QN(n14580) );
  NAND2X0 U14924 ( .IN1(n14582), .IN2(g5595), .QN(n14581) );
  NAND2X0 U14925 ( .IN1(n13469), .IN2(n13453), .QN(n14582) );
  NOR2X0 U14926 ( .IN1(n9927), .IN2(n10318), .QN(n14579) );
  NAND2X0 U14927 ( .IN1(n14583), .IN2(n14584), .QN(g30490) );
  NAND2X0 U14928 ( .IN1(n3881), .IN2(n14537), .QN(n14584) );
  NOR2X0 U14929 ( .IN1(n14585), .IN2(n14586), .QN(n14583) );
  NOR2X0 U14930 ( .IN1(n10470), .IN2(n14587), .QN(n14586) );
  NAND2X0 U14931 ( .IN1(test_so5), .IN2(n14588), .QN(n14587) );
  NAND2X0 U14932 ( .IN1(n13469), .IN2(n14537), .QN(n14588) );
  NOR2X0 U14933 ( .IN1(n9838), .IN2(n10317), .QN(n14585) );
  NAND2X0 U14934 ( .IN1(n14589), .IN2(n14590), .QN(g30489) );
  NAND2X0 U14935 ( .IN1(n3881), .IN2(n14566), .QN(n14590) );
  NOR2X0 U14936 ( .IN1(n14591), .IN2(n14592), .QN(n14589) );
  NOR2X0 U14937 ( .IN1(n10470), .IN2(n14593), .QN(n14592) );
  NAND2X0 U14938 ( .IN1(n14594), .IN2(g5587), .QN(n14593) );
  NAND2X0 U14939 ( .IN1(n13469), .IN2(n14566), .QN(n14594) );
  INVX0 U14940 ( .INP(n3436), .ZN(n13469) );
  NAND2X0 U14941 ( .IN1(n5575), .IN2(g5517), .QN(n3436) );
  NOR2X0 U14942 ( .IN1(n9797), .IN2(n10318), .QN(n14591) );
  NAND2X0 U14943 ( .IN1(n14595), .IN2(n14596), .QN(g30488) );
  NAND2X0 U14944 ( .IN1(n3886), .IN2(n14546), .QN(n14596) );
  NOR2X0 U14945 ( .IN1(n14597), .IN2(n14598), .QN(n14595) );
  NOR2X0 U14946 ( .IN1(n10470), .IN2(n14599), .QN(n14598) );
  NAND2X0 U14947 ( .IN1(n14600), .IN2(g5583), .QN(n14599) );
  NAND2X0 U14948 ( .IN1(n14601), .IN2(n14546), .QN(n14600) );
  NOR2X0 U14949 ( .IN1(n9928), .IN2(n10317), .QN(n14597) );
  NAND2X0 U14950 ( .IN1(n14602), .IN2(n14603), .QN(g30487) );
  NAND2X0 U14951 ( .IN1(n3886), .IN2(n13453), .QN(n14603) );
  NOR2X0 U14952 ( .IN1(n14604), .IN2(n14605), .QN(n14602) );
  NOR2X0 U14953 ( .IN1(n10470), .IN2(n14606), .QN(n14605) );
  NAND2X0 U14954 ( .IN1(n14607), .IN2(g5579), .QN(n14606) );
  NAND2X0 U14955 ( .IN1(n14601), .IN2(n13453), .QN(n14607) );
  INVX0 U14956 ( .INP(n3869), .ZN(n13453) );
  NAND2X0 U14957 ( .IN1(n5389), .IN2(g5535), .QN(n3869) );
  NOR2X0 U14958 ( .IN1(n10017), .IN2(n10318), .QN(n14604) );
  NAND2X0 U14959 ( .IN1(n14608), .IN2(n14609), .QN(g30486) );
  NAND2X0 U14960 ( .IN1(n3886), .IN2(n14537), .QN(n14609) );
  NOR2X0 U14961 ( .IN1(n14610), .IN2(n14611), .QN(n14608) );
  NOR2X0 U14962 ( .IN1(n10470), .IN2(n14612), .QN(n14611) );
  NAND2X0 U14963 ( .IN1(n14613), .IN2(g5575), .QN(n14612) );
  NAND2X0 U14964 ( .IN1(n14601), .IN2(n14537), .QN(n14613) );
  INVX0 U14965 ( .INP(n3871), .ZN(n14537) );
  NAND2X0 U14966 ( .IN1(n5566), .IN2(g5527), .QN(n3871) );
  NOR2X0 U14967 ( .IN1(n9798), .IN2(n10318), .QN(n14610) );
  NAND2X0 U14968 ( .IN1(n14614), .IN2(n14615), .QN(g30485) );
  NAND2X0 U14969 ( .IN1(n3886), .IN2(n14566), .QN(n14615) );
  NOR2X0 U14970 ( .IN1(n14616), .IN2(n14617), .QN(n14614) );
  NOR2X0 U14971 ( .IN1(n10470), .IN2(n14618), .QN(n14617) );
  NAND2X0 U14972 ( .IN1(n14619), .IN2(g5571), .QN(n14618) );
  NAND2X0 U14973 ( .IN1(n14601), .IN2(n14566), .QN(n14619) );
  INVX0 U14974 ( .INP(n3874), .ZN(n14566) );
  NAND2X0 U14975 ( .IN1(n5566), .IN2(n5389), .QN(n3874) );
  INVX0 U14976 ( .INP(n3437), .ZN(n14601) );
  NAND2X0 U14977 ( .IN1(n10057), .IN2(g5511), .QN(n3437) );
  NOR2X0 U14978 ( .IN1(n9958), .IN2(n10318), .QN(n14616) );
  NAND2X0 U14979 ( .IN1(n14620), .IN2(n14621), .QN(g30484) );
  NAND2X0 U14980 ( .IN1(n10508), .IN2(g5567), .QN(n14621) );
  NOR2X0 U14981 ( .IN1(n14622), .IN2(n14623), .QN(n14620) );
  AND2X1 U14982 ( .IN1(n3765), .IN2(n3891), .Q(n14623) );
  NOR2X0 U14983 ( .IN1(n3891), .IN2(n14624), .QN(n14622) );
  NAND2X0 U14984 ( .IN1(n10374), .IN2(g5563), .QN(n14624) );
  NAND2X0 U14985 ( .IN1(n14625), .IN2(n14626), .QN(g30483) );
  NAND2X0 U14986 ( .IN1(test_so6), .IN2(n10514), .QN(n14626) );
  NOR2X0 U14987 ( .IN1(n14627), .IN2(n14628), .QN(n14625) );
  AND2X1 U14988 ( .IN1(n3765), .IN2(n3894), .Q(n14628) );
  NOR2X0 U14989 ( .IN1(n3894), .IN2(n14629), .QN(n14627) );
  NAND2X0 U14990 ( .IN1(n10374), .IN2(g5555), .QN(n14629) );
  NAND2X0 U14991 ( .IN1(n14630), .IN2(n14631), .QN(g30482) );
  NAND2X0 U14992 ( .IN1(n10508), .IN2(g5551), .QN(n14631) );
  NOR2X0 U14993 ( .IN1(n14632), .IN2(n14633), .QN(n14630) );
  AND2X1 U14994 ( .IN1(n3765), .IN2(n3896), .Q(n14633) );
  NOR2X0 U14995 ( .IN1(n3896), .IN2(n14634), .QN(n14632) );
  NAND2X0 U14996 ( .IN1(n10374), .IN2(g5547), .QN(n14634) );
  NAND2X0 U14997 ( .IN1(n14635), .IN2(n14636), .QN(g30481) );
  NAND2X0 U14998 ( .IN1(n10508), .IN2(g5535), .QN(n14636) );
  NOR2X0 U14999 ( .IN1(n14637), .IN2(n14638), .QN(n14635) );
  AND2X1 U15000 ( .IN1(n3765), .IN2(n3898), .Q(n14638) );
  NOR2X0 U15001 ( .IN1(n3898), .IN2(n14639), .QN(n14637) );
  NAND2X0 U15002 ( .IN1(n10375), .IN2(g5543), .QN(n14639) );
  NOR2X0 U15003 ( .IN1(g5511), .IN2(n13460), .QN(g30480) );
  NAND2X0 U15004 ( .IN1(n14640), .IN2(n5647), .QN(n13460) );
  NOR2X0 U15005 ( .IN1(n10470), .IN2(n13464), .QN(n14640) );
  INVX0 U15006 ( .INP(n13450), .ZN(n13464) );
  NAND2X0 U15007 ( .IN1(n3833), .IN2(n12615), .QN(n13450) );
  NAND2X0 U15008 ( .IN1(n14641), .IN2(n14642), .QN(g30479) );
  NAND2X0 U15009 ( .IN1(n10508), .IN2(g5268), .QN(n14642) );
  NOR2X0 U15010 ( .IN1(n14643), .IN2(n14644), .QN(n14641) );
  NOR2X0 U15011 ( .IN1(n12619), .IN2(n14160), .QN(n14644) );
  NOR2X0 U15012 ( .IN1(n9810), .IN2(n14645), .QN(n14643) );
  NAND2X0 U15013 ( .IN1(n14646), .IN2(n14647), .QN(g30478) );
  NAND2X0 U15014 ( .IN1(n14648), .IN2(n3765), .QN(n14647) );
  NOR2X0 U15015 ( .IN1(n14649), .IN2(n14650), .QN(n14646) );
  NOR2X0 U15016 ( .IN1(n9975), .IN2(n10318), .QN(n14650) );
  NOR2X0 U15017 ( .IN1(n10470), .IN2(n14651), .QN(n14649) );
  OR2X1 U15018 ( .IN1(n14648), .IN2(n9915), .Q(n14651) );
  NOR2X0 U15019 ( .IN1(n3902), .IN2(n5650), .QN(n14648) );
  NAND2X0 U15020 ( .IN1(n14652), .IN2(n14653), .QN(g30477) );
  NAND2X0 U15021 ( .IN1(n13477), .IN2(n3765), .QN(n14653) );
  NOR2X0 U15022 ( .IN1(n14654), .IN2(n14655), .QN(n14652) );
  NOR2X0 U15023 ( .IN1(n9869), .IN2(n10319), .QN(n14655) );
  NOR2X0 U15024 ( .IN1(n10470), .IN2(n14656), .QN(n14654) );
  OR2X1 U15025 ( .IN1(n13477), .IN2(n9977), .Q(n14656) );
  NOR2X0 U15026 ( .IN1(n3904), .IN2(n5650), .QN(n13477) );
  NAND2X0 U15027 ( .IN1(n14657), .IN2(n14658), .QN(g30476) );
  NAND2X0 U15028 ( .IN1(n14659), .IN2(n3765), .QN(n14658) );
  NOR2X0 U15029 ( .IN1(n14660), .IN2(n14661), .QN(n14657) );
  NOR2X0 U15030 ( .IN1(n9811), .IN2(n10319), .QN(n14661) );
  NOR2X0 U15031 ( .IN1(n10469), .IN2(n14662), .QN(n14660) );
  OR2X1 U15032 ( .IN1(n14659), .IN2(n9952), .Q(n14662) );
  NOR2X0 U15033 ( .IN1(n3907), .IN2(n5650), .QN(n14659) );
  NAND2X0 U15034 ( .IN1(n14663), .IN2(n14664), .QN(g30475) );
  NAND2X0 U15035 ( .IN1(n3908), .IN2(n14665), .QN(n14664) );
  NOR2X0 U15036 ( .IN1(n14666), .IN2(n14667), .QN(n14663) );
  NOR2X0 U15037 ( .IN1(n10469), .IN2(n14668), .QN(n14667) );
  NAND2X0 U15038 ( .IN1(n14669), .IN2(g5268), .QN(n14668) );
  NAND2X0 U15039 ( .IN1(n14670), .IN2(n14665), .QN(n14669) );
  NOR2X0 U15040 ( .IN1(n9846), .IN2(n10319), .QN(n14666) );
  NAND2X0 U15041 ( .IN1(n14671), .IN2(n14672), .QN(g30474) );
  NAND2X0 U15042 ( .IN1(n3908), .IN2(n13476), .QN(n14672) );
  NOR2X0 U15043 ( .IN1(n14673), .IN2(n14674), .QN(n14671) );
  NOR2X0 U15044 ( .IN1(n10469), .IN2(n14675), .QN(n14674) );
  NAND2X0 U15045 ( .IN1(n14676), .IN2(g5264), .QN(n14675) );
  NAND2X0 U15046 ( .IN1(n14670), .IN2(n13476), .QN(n14676) );
  NOR2X0 U15047 ( .IN1(n9973), .IN2(n10319), .QN(n14673) );
  NAND2X0 U15048 ( .IN1(n14677), .IN2(n14678), .QN(g30473) );
  NAND2X0 U15049 ( .IN1(n3908), .IN2(n14679), .QN(n14678) );
  NOR2X0 U15050 ( .IN1(n14680), .IN2(n14681), .QN(n14677) );
  NOR2X0 U15051 ( .IN1(n10469), .IN2(n14682), .QN(n14681) );
  NAND2X0 U15052 ( .IN1(n14683), .IN2(g5260), .QN(n14682) );
  NAND2X0 U15053 ( .IN1(n14670), .IN2(n14679), .QN(n14683) );
  NOR2X0 U15054 ( .IN1(n9884), .IN2(n10319), .QN(n14680) );
  NAND2X0 U15055 ( .IN1(n14684), .IN2(n14685), .QN(g30472) );
  NAND2X0 U15056 ( .IN1(n3908), .IN2(n14686), .QN(n14685) );
  NOR2X0 U15057 ( .IN1(n14687), .IN2(n14688), .QN(n14684) );
  NOR2X0 U15058 ( .IN1(n10469), .IN2(n14689), .QN(n14688) );
  NAND2X0 U15059 ( .IN1(n14690), .IN2(g5256), .QN(n14689) );
  NAND2X0 U15060 ( .IN1(n14670), .IN2(n14686), .QN(n14690) );
  INVX0 U15061 ( .INP(n3444), .ZN(n14670) );
  NAND2X0 U15062 ( .IN1(g5164), .IN2(g5170), .QN(n3444) );
  NOR2X0 U15063 ( .IN1(n9943), .IN2(n10319), .QN(n14687) );
  NAND2X0 U15064 ( .IN1(n14691), .IN2(n14692), .QN(g30471) );
  NAND2X0 U15065 ( .IN1(n3914), .IN2(n14665), .QN(n14692) );
  NOR2X0 U15066 ( .IN1(n14693), .IN2(n14694), .QN(n14691) );
  NOR2X0 U15067 ( .IN1(n10469), .IN2(n14695), .QN(n14694) );
  NAND2X0 U15068 ( .IN1(n14696), .IN2(g5252), .QN(n14695) );
  NAND2X0 U15069 ( .IN1(n13492), .IN2(n14665), .QN(n14696) );
  NOR2X0 U15070 ( .IN1(n9847), .IN2(n10320), .QN(n14693) );
  NAND2X0 U15071 ( .IN1(n14697), .IN2(n14698), .QN(g30470) );
  NAND2X0 U15072 ( .IN1(n3914), .IN2(n13476), .QN(n14698) );
  NOR2X0 U15073 ( .IN1(n14699), .IN2(n14700), .QN(n14697) );
  NOR2X0 U15074 ( .IN1(n10469), .IN2(n14701), .QN(n14700) );
  NAND2X0 U15075 ( .IN1(n14702), .IN2(g5248), .QN(n14701) );
  NAND2X0 U15076 ( .IN1(n13492), .IN2(n13476), .QN(n14702) );
  NOR2X0 U15077 ( .IN1(n9921), .IN2(n10320), .QN(n14699) );
  NAND2X0 U15078 ( .IN1(n14703), .IN2(n14704), .QN(g30469) );
  NAND2X0 U15079 ( .IN1(n3914), .IN2(n14679), .QN(n14704) );
  NOR2X0 U15080 ( .IN1(n14705), .IN2(n14706), .QN(n14703) );
  NOR2X0 U15081 ( .IN1(n10469), .IN2(n14707), .QN(n14706) );
  NAND2X0 U15082 ( .IN1(n14708), .IN2(g5244), .QN(n14707) );
  NAND2X0 U15083 ( .IN1(n13492), .IN2(n14679), .QN(n14708) );
  AND2X1 U15084 ( .IN1(n10497), .IN2(test_so82), .Q(n14705) );
  NAND2X0 U15085 ( .IN1(n14709), .IN2(n14710), .QN(g30468) );
  NAND2X0 U15086 ( .IN1(n3914), .IN2(n14686), .QN(n14710) );
  NOR2X0 U15087 ( .IN1(n14711), .IN2(n14712), .QN(n14709) );
  NOR2X0 U15088 ( .IN1(n10469), .IN2(n14713), .QN(n14712) );
  NAND2X0 U15089 ( .IN1(n14714), .IN2(g5240), .QN(n14713) );
  NAND2X0 U15090 ( .IN1(n13492), .IN2(n14686), .QN(n14714) );
  INVX0 U15091 ( .INP(n3446), .ZN(n13492) );
  NAND2X0 U15092 ( .IN1(n5570), .IN2(g5170), .QN(n3446) );
  NOR2X0 U15093 ( .IN1(n9812), .IN2(n10320), .QN(n14711) );
  NAND2X0 U15094 ( .IN1(n14715), .IN2(n14716), .QN(g30467) );
  NAND2X0 U15095 ( .IN1(n3919), .IN2(n14665), .QN(n14716) );
  NOR2X0 U15096 ( .IN1(n14717), .IN2(n14718), .QN(n14715) );
  NOR2X0 U15097 ( .IN1(n10469), .IN2(n14719), .QN(n14718) );
  NAND2X0 U15098 ( .IN1(n14720), .IN2(g5236), .QN(n14719) );
  NAND2X0 U15099 ( .IN1(n14721), .IN2(n14665), .QN(n14720) );
  NOR2X0 U15100 ( .IN1(n9922), .IN2(n10320), .QN(n14717) );
  NAND2X0 U15101 ( .IN1(n14722), .IN2(n14723), .QN(g30466) );
  NAND2X0 U15102 ( .IN1(n3919), .IN2(n13476), .QN(n14723) );
  NOR2X0 U15103 ( .IN1(n14724), .IN2(n14725), .QN(n14722) );
  NOR2X0 U15104 ( .IN1(n10469), .IN2(n14726), .QN(n14725) );
  NAND2X0 U15105 ( .IN1(n14727), .IN2(g5232), .QN(n14726) );
  NAND2X0 U15106 ( .IN1(n14721), .IN2(n13476), .QN(n14727) );
  INVX0 U15107 ( .INP(n3902), .ZN(n13476) );
  NAND2X0 U15108 ( .IN1(n5384), .IN2(g5188), .QN(n3902) );
  NOR2X0 U15109 ( .IN1(n9916), .IN2(n10320), .QN(n14724) );
  NAND2X0 U15110 ( .IN1(n14728), .IN2(n14729), .QN(g30465) );
  NAND2X0 U15111 ( .IN1(n3919), .IN2(n14679), .QN(n14729) );
  NOR2X0 U15112 ( .IN1(n14730), .IN2(n14731), .QN(n14728) );
  NOR2X0 U15113 ( .IN1(n10469), .IN2(n14732), .QN(n14731) );
  NAND2X0 U15114 ( .IN1(test_so82), .IN2(n14733), .QN(n14732) );
  NAND2X0 U15115 ( .IN1(n14721), .IN2(n14679), .QN(n14733) );
  INVX0 U15116 ( .INP(n3904), .ZN(n14679) );
  NAND2X0 U15117 ( .IN1(n5567), .IN2(g5180), .QN(n3904) );
  NOR2X0 U15118 ( .IN1(n9813), .IN2(n10320), .QN(n14730) );
  NAND2X0 U15119 ( .IN1(n14734), .IN2(n14735), .QN(g30464) );
  NAND2X0 U15120 ( .IN1(n3919), .IN2(n14686), .QN(n14735) );
  NOR2X0 U15121 ( .IN1(n14736), .IN2(n14737), .QN(n14734) );
  NOR2X0 U15122 ( .IN1(n10469), .IN2(n14738), .QN(n14737) );
  NAND2X0 U15123 ( .IN1(n14739), .IN2(g5224), .QN(n14738) );
  NAND2X0 U15124 ( .IN1(n14721), .IN2(n14686), .QN(n14739) );
  INVX0 U15125 ( .INP(n3907), .ZN(n14686) );
  NAND2X0 U15126 ( .IN1(n5567), .IN2(n5384), .QN(n3907) );
  INVX0 U15127 ( .INP(n3447), .ZN(n14721) );
  NAND2X0 U15128 ( .IN1(n10052), .IN2(g5164), .QN(n3447) );
  NOR2X0 U15129 ( .IN1(n9954), .IN2(n10320), .QN(n14736) );
  NAND2X0 U15130 ( .IN1(n14740), .IN2(n14741), .QN(g30463) );
  NAND2X0 U15131 ( .IN1(n10508), .IN2(g5220), .QN(n14741) );
  NOR2X0 U15132 ( .IN1(n14742), .IN2(n14743), .QN(n14740) );
  AND2X1 U15133 ( .IN1(n3765), .IN2(n3924), .Q(n14743) );
  NOR2X0 U15134 ( .IN1(n3924), .IN2(n14744), .QN(n14742) );
  NAND2X0 U15135 ( .IN1(n10376), .IN2(g5216), .QN(n14744) );
  NAND2X0 U15136 ( .IN1(n14745), .IN2(n14746), .QN(g30462) );
  OR2X1 U15137 ( .IN1(n10311), .IN2(n9977), .Q(n14746) );
  NOR2X0 U15138 ( .IN1(n14747), .IN2(n14748), .QN(n14745) );
  AND2X1 U15139 ( .IN1(n3765), .IN2(n3927), .Q(n14748) );
  NOR2X0 U15140 ( .IN1(n3927), .IN2(n14749), .QN(n14747) );
  NAND2X0 U15141 ( .IN1(n10376), .IN2(g5208), .QN(n14749) );
  NAND2X0 U15142 ( .IN1(n14750), .IN2(n14751), .QN(g30461) );
  NAND2X0 U15143 ( .IN1(n10509), .IN2(g5204), .QN(n14751) );
  NOR2X0 U15144 ( .IN1(n14752), .IN2(n14753), .QN(n14750) );
  AND2X1 U15145 ( .IN1(n3765), .IN2(n3929), .Q(n14753) );
  NOR2X0 U15146 ( .IN1(n3929), .IN2(n14754), .QN(n14752) );
  NAND2X0 U15147 ( .IN1(n10375), .IN2(g5200), .QN(n14754) );
  NAND2X0 U15148 ( .IN1(n14755), .IN2(n14756), .QN(g30460) );
  NAND2X0 U15149 ( .IN1(n10509), .IN2(g5188), .QN(n14756) );
  NOR2X0 U15150 ( .IN1(n14757), .IN2(n14758), .QN(n14755) );
  AND2X1 U15151 ( .IN1(n3765), .IN2(n3931), .Q(n14758) );
  NOR2X0 U15152 ( .IN1(n3931), .IN2(n14759), .QN(n14757) );
  NAND2X0 U15153 ( .IN1(n10373), .IN2(g5196), .QN(n14759) );
  NOR2X0 U15154 ( .IN1(g5164), .IN2(n13483), .QN(g30459) );
  NAND2X0 U15155 ( .IN1(n14760), .IN2(n5650), .QN(n13483) );
  NOR2X0 U15156 ( .IN1(n10468), .IN2(n13487), .QN(n14760) );
  INVX0 U15157 ( .INP(n13473), .ZN(n13487) );
  NAND2X0 U15158 ( .IN1(n3833), .IN2(n11688), .QN(n13473) );
  INVX0 U15159 ( .INP(n12618), .ZN(n11688) );
  NAND2X0 U15160 ( .IN1(n14761), .IN2(n10389), .QN(g30458) );
  NOR2X0 U15161 ( .IN1(n14762), .IN2(n14763), .QN(n14761) );
  NOR2X0 U15162 ( .IN1(n5846), .IN2(n14764), .QN(n14763) );
  AND2X1 U15163 ( .IN1(g113), .IN2(n14764), .Q(n14762) );
  NOR2X0 U15164 ( .IN1(g4459), .IN2(n9703), .QN(n14764) );
  NAND2X0 U15165 ( .IN1(n14765), .IN2(n14766), .QN(g30457) );
  NAND2X0 U15166 ( .IN1(n10509), .IN2(g4122), .QN(n14766) );
  NAND2X0 U15167 ( .IN1(n14767), .IN2(n10389), .QN(n14765) );
  NAND2X0 U15168 ( .IN1(n14768), .IN2(n14769), .QN(n14767) );
  NAND2X0 U15169 ( .IN1(n14770), .IN2(n5981), .QN(n14769) );
  XNOR2X1 U15170 ( .IN1(g126), .IN2(n14771), .Q(n14770) );
  NAND2X0 U15171 ( .IN1(n14772), .IN2(n5983), .QN(n14768) );
  XNOR2X1 U15172 ( .IN1(g115), .IN2(n14773), .Q(n14772) );
  NAND2X0 U15173 ( .IN1(n14774), .IN2(n14775), .QN(g30456) );
  NAND2X0 U15174 ( .IN1(n10509), .IN2(g4087), .QN(n14775) );
  NOR2X0 U15175 ( .IN1(n14776), .IN2(n14777), .QN(n14774) );
  AND2X1 U15176 ( .IN1(n3941), .IN2(n14778), .Q(n14777) );
  NOR2X0 U15177 ( .IN1(n14779), .IN2(n14780), .QN(n14776) );
  OR2X1 U15178 ( .IN1(n14071), .IN2(n5729), .Q(n14780) );
  NAND2X0 U15179 ( .IN1(n14781), .IN2(n14782), .QN(g30455) );
  NAND2X0 U15180 ( .IN1(n10509), .IN2(g3961), .QN(n14782) );
  NOR2X0 U15181 ( .IN1(n14783), .IN2(n14784), .QN(n14781) );
  NOR2X0 U15182 ( .IN1(n14160), .IN2(n12636), .QN(n14784) );
  NOR2X0 U15183 ( .IN1(n9816), .IN2(n14785), .QN(n14783) );
  NAND2X0 U15184 ( .IN1(n14786), .IN2(n14787), .QN(g30454) );
  OR2X1 U15185 ( .IN1(n14788), .IN2(n14160), .Q(n14787) );
  NOR2X0 U15186 ( .IN1(n14789), .IN2(n14790), .QN(n14786) );
  NOR2X0 U15187 ( .IN1(n9989), .IN2(n10321), .QN(n14790) );
  NOR2X0 U15188 ( .IN1(n10468), .IN2(n14791), .QN(n14789) );
  NAND2X0 U15189 ( .IN1(n14788), .IN2(g3913), .QN(n14791) );
  NAND2X0 U15190 ( .IN1(test_so33), .IN2(n13544), .QN(n14788) );
  NAND2X0 U15191 ( .IN1(n14792), .IN2(n14793), .QN(g30453) );
  NAND2X0 U15192 ( .IN1(n13545), .IN2(n3765), .QN(n14793) );
  INVX0 U15193 ( .INP(n14794), .ZN(n13545) );
  NOR2X0 U15194 ( .IN1(n14795), .IN2(n14796), .QN(n14792) );
  NOR2X0 U15195 ( .IN1(n9875), .IN2(n10321), .QN(n14796) );
  NOR2X0 U15196 ( .IN1(n10468), .IN2(n14797), .QN(n14795) );
  NAND2X0 U15197 ( .IN1(n14794), .IN2(g3905), .QN(n14797) );
  NAND2X0 U15198 ( .IN1(test_so33), .IN2(n14798), .QN(n14794) );
  NAND2X0 U15199 ( .IN1(n14799), .IN2(n14800), .QN(g30452) );
  OR2X1 U15200 ( .IN1(n14801), .IN2(n14160), .Q(n14800) );
  NOR2X0 U15201 ( .IN1(n14802), .IN2(n14803), .QN(n14799) );
  AND2X1 U15202 ( .IN1(n10497), .IN2(test_so65), .Q(n14803) );
  NOR2X0 U15203 ( .IN1(n10468), .IN2(n14804), .QN(n14802) );
  NAND2X0 U15204 ( .IN1(n14801), .IN2(g3897), .QN(n14804) );
  NAND2X0 U15205 ( .IN1(test_so33), .IN2(n14805), .QN(n14801) );
  NAND2X0 U15206 ( .IN1(n14806), .IN2(n14807), .QN(g30451) );
  NAND2X0 U15207 ( .IN1(n3951), .IN2(n14808), .QN(n14807) );
  NOR2X0 U15208 ( .IN1(n14809), .IN2(n14810), .QN(n14806) );
  NOR2X0 U15209 ( .IN1(n10468), .IN2(n14811), .QN(n14810) );
  NAND2X0 U15210 ( .IN1(n14812), .IN2(g3961), .QN(n14811) );
  NAND2X0 U15211 ( .IN1(n14813), .IN2(n14808), .QN(n14812) );
  NOR2X0 U15212 ( .IN1(n9855), .IN2(n10321), .QN(n14809) );
  NAND2X0 U15213 ( .IN1(n14814), .IN2(n14815), .QN(g30450) );
  NAND2X0 U15214 ( .IN1(n3951), .IN2(n13544), .QN(n14815) );
  NOR2X0 U15215 ( .IN1(n14816), .IN2(n14817), .QN(n14814) );
  NOR2X0 U15216 ( .IN1(n10468), .IN2(n14818), .QN(n14817) );
  NAND2X0 U15217 ( .IN1(n14819), .IN2(g3957), .QN(n14818) );
  NAND2X0 U15218 ( .IN1(n14813), .IN2(n13544), .QN(n14819) );
  NOR2X0 U15219 ( .IN1(n9987), .IN2(n10321), .QN(n14816) );
  NAND2X0 U15220 ( .IN1(n14820), .IN2(n14821), .QN(g30449) );
  NAND2X0 U15221 ( .IN1(n3951), .IN2(n14798), .QN(n14821) );
  NOR2X0 U15222 ( .IN1(n14822), .IN2(n14823), .QN(n14820) );
  NOR2X0 U15223 ( .IN1(n10468), .IN2(n14824), .QN(n14823) );
  NAND2X0 U15224 ( .IN1(n14825), .IN2(g3953), .QN(n14824) );
  NAND2X0 U15225 ( .IN1(n14813), .IN2(n14798), .QN(n14825) );
  NOR2X0 U15226 ( .IN1(n9889), .IN2(n10321), .QN(n14822) );
  NAND2X0 U15227 ( .IN1(n14826), .IN2(n14827), .QN(g30448) );
  NAND2X0 U15228 ( .IN1(n3951), .IN2(n14805), .QN(n14827) );
  NOR2X0 U15229 ( .IN1(n14828), .IN2(n14829), .QN(n14826) );
  NOR2X0 U15230 ( .IN1(n10468), .IN2(n14830), .QN(n14829) );
  NAND2X0 U15231 ( .IN1(test_so65), .IN2(n14831), .QN(n14830) );
  NAND2X0 U15232 ( .IN1(n14813), .IN2(n14805), .QN(n14831) );
  INVX0 U15233 ( .INP(n3479), .ZN(n14813) );
  NAND2X0 U15234 ( .IN1(g3857), .IN2(g3863), .QN(n3479) );
  NOR2X0 U15235 ( .IN1(n9946), .IN2(n10321), .QN(n14828) );
  NAND2X0 U15236 ( .IN1(n14832), .IN2(n14833), .QN(g30447) );
  NAND2X0 U15237 ( .IN1(n3957), .IN2(n14808), .QN(n14833) );
  NOR2X0 U15238 ( .IN1(n14834), .IN2(n14835), .QN(n14832) );
  NOR2X0 U15239 ( .IN1(n10467), .IN2(n14836), .QN(n14835) );
  NAND2X0 U15240 ( .IN1(n14837), .IN2(g3945), .QN(n14836) );
  NAND2X0 U15241 ( .IN1(n13560), .IN2(n14808), .QN(n14837) );
  NOR2X0 U15242 ( .IN1(n9856), .IN2(n10321), .QN(n14834) );
  NAND2X0 U15243 ( .IN1(n14838), .IN2(n14839), .QN(g30446) );
  NAND2X0 U15244 ( .IN1(n3957), .IN2(n13544), .QN(n14839) );
  NOR2X0 U15245 ( .IN1(n14840), .IN2(n14841), .QN(n14838) );
  NOR2X0 U15246 ( .IN1(n10467), .IN2(n14842), .QN(n14841) );
  NAND2X0 U15247 ( .IN1(n14843), .IN2(g3941), .QN(n14842) );
  NAND2X0 U15248 ( .IN1(n13560), .IN2(n13544), .QN(n14843) );
  NOR2X0 U15249 ( .IN1(n9930), .IN2(n10322), .QN(n14840) );
  NAND2X0 U15250 ( .IN1(n14844), .IN2(n14845), .QN(g30445) );
  NAND2X0 U15251 ( .IN1(n3957), .IN2(n14798), .QN(n14845) );
  NOR2X0 U15252 ( .IN1(n14846), .IN2(n14847), .QN(n14844) );
  NOR2X0 U15253 ( .IN1(n10467), .IN2(n14848), .QN(n14847) );
  NAND2X0 U15254 ( .IN1(n14849), .IN2(g3937), .QN(n14848) );
  NAND2X0 U15255 ( .IN1(n13560), .IN2(n14798), .QN(n14849) );
  NOR2X0 U15256 ( .IN1(n9839), .IN2(n10322), .QN(n14846) );
  NAND2X0 U15257 ( .IN1(n14850), .IN2(n14851), .QN(g30444) );
  NAND2X0 U15258 ( .IN1(n3957), .IN2(n14805), .QN(n14851) );
  NOR2X0 U15259 ( .IN1(n14852), .IN2(n14853), .QN(n14850) );
  NOR2X0 U15260 ( .IN1(n10467), .IN2(n14854), .QN(n14853) );
  NAND2X0 U15261 ( .IN1(n14855), .IN2(g3933), .QN(n14854) );
  NAND2X0 U15262 ( .IN1(n13560), .IN2(n14805), .QN(n14855) );
  INVX0 U15263 ( .INP(n3481), .ZN(n13560) );
  NAND2X0 U15264 ( .IN1(n5572), .IN2(g3863), .QN(n3481) );
  NOR2X0 U15265 ( .IN1(n9817), .IN2(n10322), .QN(n14852) );
  NAND2X0 U15266 ( .IN1(n14856), .IN2(n14857), .QN(g30443) );
  NAND2X0 U15267 ( .IN1(n3962), .IN2(n14808), .QN(n14857) );
  NOR2X0 U15268 ( .IN1(n14858), .IN2(n14859), .QN(n14856) );
  NOR2X0 U15269 ( .IN1(n10467), .IN2(n14860), .QN(n14859) );
  NAND2X0 U15270 ( .IN1(n14861), .IN2(g3929), .QN(n14860) );
  NAND2X0 U15271 ( .IN1(n14862), .IN2(n14808), .QN(n14861) );
  NOR2X0 U15272 ( .IN1(n9931), .IN2(n10322), .QN(n14858) );
  NAND2X0 U15273 ( .IN1(n14863), .IN2(n14864), .QN(g30442) );
  NAND2X0 U15274 ( .IN1(n3962), .IN2(n13544), .QN(n14864) );
  NOR2X0 U15275 ( .IN1(n14865), .IN2(n14866), .QN(n14863) );
  NOR2X0 U15276 ( .IN1(n10467), .IN2(n14867), .QN(n14866) );
  NAND2X0 U15277 ( .IN1(n14868), .IN2(g3925), .QN(n14867) );
  NAND2X0 U15278 ( .IN1(n14862), .IN2(n13544), .QN(n14868) );
  INVX0 U15279 ( .INP(n3945), .ZN(n13544) );
  NAND2X0 U15280 ( .IN1(n5387), .IN2(g3881), .QN(n3945) );
  NOR2X0 U15281 ( .IN1(n10021), .IN2(n10322), .QN(n14865) );
  NAND2X0 U15282 ( .IN1(n14869), .IN2(n14870), .QN(g30441) );
  NAND2X0 U15283 ( .IN1(n3962), .IN2(n14798), .QN(n14870) );
  NOR2X0 U15284 ( .IN1(n14871), .IN2(n14872), .QN(n14869) );
  NOR2X0 U15285 ( .IN1(n10467), .IN2(n14873), .QN(n14872) );
  NAND2X0 U15286 ( .IN1(n14874), .IN2(g3921), .QN(n14873) );
  NAND2X0 U15287 ( .IN1(n14862), .IN2(n14798), .QN(n14874) );
  INVX0 U15288 ( .INP(n3947), .ZN(n14798) );
  NAND2X0 U15289 ( .IN1(n5564), .IN2(g3873), .QN(n3947) );
  NOR2X0 U15290 ( .IN1(n9818), .IN2(n10322), .QN(n14871) );
  NAND2X0 U15291 ( .IN1(n14875), .IN2(n14876), .QN(g30440) );
  NAND2X0 U15292 ( .IN1(n3962), .IN2(n14805), .QN(n14876) );
  NOR2X0 U15293 ( .IN1(n14877), .IN2(n14878), .QN(n14875) );
  NOR2X0 U15294 ( .IN1(n10466), .IN2(n14879), .QN(n14878) );
  NAND2X0 U15295 ( .IN1(n14880), .IN2(g3917), .QN(n14879) );
  NAND2X0 U15296 ( .IN1(n14862), .IN2(n14805), .QN(n14880) );
  INVX0 U15297 ( .INP(n3950), .ZN(n14805) );
  NAND2X0 U15298 ( .IN1(n5564), .IN2(n5387), .QN(n3950) );
  INVX0 U15299 ( .INP(n3482), .ZN(n14862) );
  NAND2X0 U15300 ( .IN1(n10054), .IN2(g3857), .QN(n3482) );
  AND2X1 U15301 ( .IN1(n10496), .IN2(test_so24), .Q(n14877) );
  NAND2X0 U15302 ( .IN1(n14881), .IN2(n14882), .QN(g30439) );
  NAND2X0 U15303 ( .IN1(n10509), .IN2(g3913), .QN(n14882) );
  NOR2X0 U15304 ( .IN1(n14883), .IN2(n14884), .QN(n14881) );
  AND2X1 U15305 ( .IN1(n3765), .IN2(n3967), .Q(n14884) );
  NOR2X0 U15306 ( .IN1(n3967), .IN2(n14885), .QN(n14883) );
  NAND2X0 U15307 ( .IN1(n10371), .IN2(g3909), .QN(n14885) );
  NAND2X0 U15308 ( .IN1(n14886), .IN2(n14887), .QN(g30438) );
  NAND2X0 U15309 ( .IN1(n10509), .IN2(g3905), .QN(n14887) );
  NOR2X0 U15310 ( .IN1(n14888), .IN2(n14889), .QN(n14886) );
  AND2X1 U15311 ( .IN1(n3765), .IN2(n3970), .Q(n14889) );
  NOR2X0 U15312 ( .IN1(n3970), .IN2(n14890), .QN(n14888) );
  NAND2X0 U15313 ( .IN1(n10371), .IN2(g3901), .QN(n14890) );
  NAND2X0 U15314 ( .IN1(n14891), .IN2(n14892), .QN(g30437) );
  NAND2X0 U15315 ( .IN1(n10509), .IN2(g3897), .QN(n14892) );
  NOR2X0 U15316 ( .IN1(n14893), .IN2(n14894), .QN(n14891) );
  AND2X1 U15317 ( .IN1(n3765), .IN2(n3972), .Q(n14894) );
  NOR2X0 U15318 ( .IN1(n3972), .IN2(n14895), .QN(n14893) );
  NAND2X0 U15319 ( .IN1(n10371), .IN2(g3893), .QN(n14895) );
  NAND2X0 U15320 ( .IN1(n14896), .IN2(n14897), .QN(g30436) );
  NAND2X0 U15321 ( .IN1(n10509), .IN2(g3881), .QN(n14897) );
  NOR2X0 U15322 ( .IN1(n14898), .IN2(n14899), .QN(n14896) );
  AND2X1 U15323 ( .IN1(n3765), .IN2(n3974), .Q(n14899) );
  NOR2X0 U15324 ( .IN1(n3974), .IN2(n14900), .QN(n14898) );
  NAND2X0 U15325 ( .IN1(test_so24), .IN2(n10389), .QN(n14900) );
  NOR2X0 U15326 ( .IN1(g3857), .IN2(n13552), .QN(g30435) );
  NAND2X0 U15327 ( .IN1(n14901), .IN2(n13541), .QN(n13552) );
  NAND2X0 U15328 ( .IN1(n14397), .IN2(n3799), .QN(n13541) );
  NOR2X0 U15329 ( .IN1(n5480), .IN2(n5340), .QN(n14397) );
  NOR2X0 U15330 ( .IN1(test_so33), .IN2(n10460), .QN(n14901) );
  NAND2X0 U15331 ( .IN1(n14902), .IN2(n14903), .QN(g30434) );
  NAND2X0 U15332 ( .IN1(n10509), .IN2(g3610), .QN(n14903) );
  NOR2X0 U15333 ( .IN1(n14904), .IN2(n14905), .QN(n14902) );
  NOR2X0 U15334 ( .IN1(n14160), .IN2(n12635), .QN(n14905) );
  NOR2X0 U15335 ( .IN1(n9802), .IN2(n14906), .QN(n14904) );
  NAND2X0 U15336 ( .IN1(n14907), .IN2(n14908), .QN(g30433) );
  NAND2X0 U15337 ( .IN1(n14909), .IN2(n3765), .QN(n14908) );
  NOR2X0 U15338 ( .IN1(n14910), .IN2(n14911), .QN(n14907) );
  NOR2X0 U15339 ( .IN1(n9999), .IN2(n10322), .QN(n14911) );
  NOR2X0 U15340 ( .IN1(n10466), .IN2(n14912), .QN(n14910) );
  OR2X1 U15341 ( .IN1(n14909), .IN2(n10027), .Q(n14912) );
  NOR2X0 U15342 ( .IN1(n3978), .IN2(n5645), .QN(n14909) );
  NAND2X0 U15343 ( .IN1(n14913), .IN2(n14914), .QN(g30432) );
  NAND2X0 U15344 ( .IN1(n13568), .IN2(n3765), .QN(n14914) );
  NOR2X0 U15345 ( .IN1(n14915), .IN2(n14916), .QN(n14913) );
  AND2X1 U15346 ( .IN1(n10497), .IN2(test_so43), .Q(n14916) );
  NOR2X0 U15347 ( .IN1(n10468), .IN2(n14917), .QN(n14915) );
  OR2X1 U15348 ( .IN1(n13568), .IN2(n10001), .Q(n14917) );
  NOR2X0 U15349 ( .IN1(n3980), .IN2(n5645), .QN(n13568) );
  NAND2X0 U15350 ( .IN1(n14918), .IN2(n14919), .QN(g30431) );
  NAND2X0 U15351 ( .IN1(n14920), .IN2(n3765), .QN(n14919) );
  NOR2X0 U15352 ( .IN1(n14921), .IN2(n14922), .QN(n14918) );
  NOR2X0 U15353 ( .IN1(n9803), .IN2(n10323), .QN(n14922) );
  NOR2X0 U15354 ( .IN1(n10466), .IN2(n14923), .QN(n14921) );
  OR2X1 U15355 ( .IN1(n14920), .IN2(n9962), .Q(n14923) );
  NOR2X0 U15356 ( .IN1(n3983), .IN2(n5645), .QN(n14920) );
  NAND2X0 U15357 ( .IN1(n14924), .IN2(n14925), .QN(g30430) );
  NAND2X0 U15358 ( .IN1(n3984), .IN2(n14926), .QN(n14925) );
  NOR2X0 U15359 ( .IN1(n14927), .IN2(n14928), .QN(n14924) );
  NOR2X0 U15360 ( .IN1(n10467), .IN2(n14929), .QN(n14928) );
  NAND2X0 U15361 ( .IN1(n14930), .IN2(g3610), .QN(n14929) );
  NAND2X0 U15362 ( .IN1(n14931), .IN2(n14926), .QN(n14930) );
  NOR2X0 U15363 ( .IN1(n9861), .IN2(n10323), .QN(n14927) );
  NAND2X0 U15364 ( .IN1(n14932), .IN2(n14933), .QN(g30429) );
  NAND2X0 U15365 ( .IN1(n3984), .IN2(n13567), .QN(n14933) );
  NOR2X0 U15366 ( .IN1(n14934), .IN2(n14935), .QN(n14932) );
  NOR2X0 U15367 ( .IN1(n10466), .IN2(n14936), .QN(n14935) );
  NAND2X0 U15368 ( .IN1(n14937), .IN2(g3606), .QN(n14936) );
  NAND2X0 U15369 ( .IN1(n14931), .IN2(n13567), .QN(n14937) );
  NOR2X0 U15370 ( .IN1(n9997), .IN2(n10323), .QN(n14934) );
  NAND2X0 U15371 ( .IN1(n14938), .IN2(n14939), .QN(g30428) );
  NAND2X0 U15372 ( .IN1(n3984), .IN2(n14940), .QN(n14939) );
  NOR2X0 U15373 ( .IN1(n14941), .IN2(n14942), .QN(n14938) );
  NOR2X0 U15374 ( .IN1(n10466), .IN2(n14943), .QN(n14942) );
  NAND2X0 U15375 ( .IN1(test_so43), .IN2(n14944), .QN(n14943) );
  NAND2X0 U15376 ( .IN1(n14931), .IN2(n14940), .QN(n14944) );
  NOR2X0 U15377 ( .IN1(n9893), .IN2(n10323), .QN(n14941) );
  NAND2X0 U15378 ( .IN1(n14945), .IN2(n14946), .QN(g30427) );
  NAND2X0 U15379 ( .IN1(n3984), .IN2(n14947), .QN(n14946) );
  NOR2X0 U15380 ( .IN1(n14948), .IN2(n14949), .QN(n14945) );
  NOR2X0 U15381 ( .IN1(n10468), .IN2(n14950), .QN(n14949) );
  NAND2X0 U15382 ( .IN1(n14951), .IN2(g3598), .QN(n14950) );
  NAND2X0 U15383 ( .IN1(n14931), .IN2(n14947), .QN(n14951) );
  INVX0 U15384 ( .INP(n3489), .ZN(n14931) );
  NAND2X0 U15385 ( .IN1(g3506), .IN2(g3512), .QN(n3489) );
  NOR2X0 U15386 ( .IN1(n9948), .IN2(n10323), .QN(n14948) );
  NAND2X0 U15387 ( .IN1(n14952), .IN2(n14953), .QN(g30426) );
  NAND2X0 U15388 ( .IN1(n3990), .IN2(n14926), .QN(n14953) );
  NOR2X0 U15389 ( .IN1(n14954), .IN2(n14955), .QN(n14952) );
  NOR2X0 U15390 ( .IN1(n10466), .IN2(n14956), .QN(n14955) );
  NAND2X0 U15391 ( .IN1(n14957), .IN2(g3594), .QN(n14956) );
  NAND2X0 U15392 ( .IN1(n13583), .IN2(n14926), .QN(n14957) );
  NOR2X0 U15393 ( .IN1(n9862), .IN2(n10323), .QN(n14954) );
  NAND2X0 U15394 ( .IN1(n14958), .IN2(n14959), .QN(g30425) );
  NAND2X0 U15395 ( .IN1(n3990), .IN2(n13567), .QN(n14959) );
  NOR2X0 U15396 ( .IN1(n14960), .IN2(n14961), .QN(n14958) );
  NOR2X0 U15397 ( .IN1(n10465), .IN2(n14962), .QN(n14961) );
  NAND2X0 U15398 ( .IN1(n14963), .IN2(g3590), .QN(n14962) );
  NAND2X0 U15399 ( .IN1(n13583), .IN2(n13567), .QN(n14963) );
  NOR2X0 U15400 ( .IN1(n9936), .IN2(n10323), .QN(n14960) );
  NAND2X0 U15401 ( .IN1(n14964), .IN2(n14965), .QN(g30424) );
  NAND2X0 U15402 ( .IN1(n3990), .IN2(n14940), .QN(n14965) );
  NOR2X0 U15403 ( .IN1(n14966), .IN2(n14967), .QN(n14964) );
  NOR2X0 U15404 ( .IN1(n10467), .IN2(n14968), .QN(n14967) );
  NAND2X0 U15405 ( .IN1(n14969), .IN2(g3586), .QN(n14968) );
  NAND2X0 U15406 ( .IN1(n13583), .IN2(n14940), .QN(n14969) );
  NOR2X0 U15407 ( .IN1(n9841), .IN2(n10324), .QN(n14966) );
  NAND2X0 U15408 ( .IN1(n14970), .IN2(n14971), .QN(g30423) );
  NAND2X0 U15409 ( .IN1(n3990), .IN2(n14947), .QN(n14971) );
  NOR2X0 U15410 ( .IN1(n14972), .IN2(n14973), .QN(n14970) );
  NOR2X0 U15411 ( .IN1(n10465), .IN2(n14974), .QN(n14973) );
  NAND2X0 U15412 ( .IN1(n14975), .IN2(g3582), .QN(n14974) );
  NAND2X0 U15413 ( .IN1(n13583), .IN2(n14947), .QN(n14975) );
  INVX0 U15414 ( .INP(n3491), .ZN(n13583) );
  NAND2X0 U15415 ( .IN1(n5576), .IN2(g3512), .QN(n3491) );
  NOR2X0 U15416 ( .IN1(n9804), .IN2(n10324), .QN(n14972) );
  NAND2X0 U15417 ( .IN1(n14976), .IN2(n14977), .QN(g30422) );
  NAND2X0 U15418 ( .IN1(n3995), .IN2(n14926), .QN(n14977) );
  NOR2X0 U15419 ( .IN1(n14978), .IN2(n14979), .QN(n14976) );
  NOR2X0 U15420 ( .IN1(n10467), .IN2(n14980), .QN(n14979) );
  NAND2X0 U15421 ( .IN1(n14981), .IN2(g3578), .QN(n14980) );
  NAND2X0 U15422 ( .IN1(n14982), .IN2(n14926), .QN(n14981) );
  NOR2X0 U15423 ( .IN1(n9937), .IN2(n10324), .QN(n14978) );
  NAND2X0 U15424 ( .IN1(n14983), .IN2(n14984), .QN(g30421) );
  NAND2X0 U15425 ( .IN1(n3995), .IN2(n13567), .QN(n14984) );
  NOR2X0 U15426 ( .IN1(n14985), .IN2(n14986), .QN(n14983) );
  NOR2X0 U15427 ( .IN1(n10465), .IN2(n14987), .QN(n14986) );
  NAND2X0 U15428 ( .IN1(n14988), .IN2(g3574), .QN(n14987) );
  NAND2X0 U15429 ( .IN1(n14982), .IN2(n13567), .QN(n14988) );
  INVX0 U15430 ( .INP(n3978), .ZN(n13567) );
  NAND2X0 U15431 ( .IN1(n5383), .IN2(g3530), .QN(n3978) );
  NOR2X0 U15432 ( .IN1(n10029), .IN2(n10324), .QN(n14985) );
  NAND2X0 U15433 ( .IN1(n14989), .IN2(n14990), .QN(g30420) );
  NAND2X0 U15434 ( .IN1(n3995), .IN2(n14940), .QN(n14990) );
  NOR2X0 U15435 ( .IN1(n14991), .IN2(n14992), .QN(n14989) );
  NOR2X0 U15436 ( .IN1(n10465), .IN2(n14993), .QN(n14992) );
  NAND2X0 U15437 ( .IN1(n14994), .IN2(g3570), .QN(n14993) );
  NAND2X0 U15438 ( .IN1(n14982), .IN2(n14940), .QN(n14994) );
  INVX0 U15439 ( .INP(n3980), .ZN(n14940) );
  NAND2X0 U15440 ( .IN1(n5569), .IN2(g3522), .QN(n3980) );
  NOR2X0 U15441 ( .IN1(n9805), .IN2(n10324), .QN(n14991) );
  NAND2X0 U15442 ( .IN1(n14995), .IN2(n14996), .QN(g30419) );
  NAND2X0 U15443 ( .IN1(n3995), .IN2(n14947), .QN(n14996) );
  NOR2X0 U15444 ( .IN1(n14997), .IN2(n14998), .QN(n14995) );
  NOR2X0 U15445 ( .IN1(n10467), .IN2(n14999), .QN(n14998) );
  NAND2X0 U15446 ( .IN1(n15000), .IN2(g3566), .QN(n14999) );
  NAND2X0 U15447 ( .IN1(n14982), .IN2(n14947), .QN(n15000) );
  INVX0 U15448 ( .INP(n3983), .ZN(n14947) );
  NAND2X0 U15449 ( .IN1(n5569), .IN2(n5383), .QN(n3983) );
  INVX0 U15450 ( .INP(n3492), .ZN(n14982) );
  NAND2X0 U15451 ( .IN1(n10058), .IN2(g3506), .QN(n3492) );
  NOR2X0 U15452 ( .IN1(n9963), .IN2(n10324), .QN(n14997) );
  NAND2X0 U15453 ( .IN1(n15001), .IN2(n15002), .QN(g30418) );
  NAND2X0 U15454 ( .IN1(n10509), .IN2(g3562), .QN(n15002) );
  NOR2X0 U15455 ( .IN1(n15003), .IN2(n15004), .QN(n15001) );
  AND2X1 U15456 ( .IN1(n3765), .IN2(n4000), .Q(n15004) );
  NOR2X0 U15457 ( .IN1(n4000), .IN2(n15005), .QN(n15003) );
  NAND2X0 U15458 ( .IN1(n10369), .IN2(g3558), .QN(n15005) );
  NAND2X0 U15459 ( .IN1(n15006), .IN2(n15007), .QN(g30417) );
  NAND2X0 U15460 ( .IN1(n10509), .IN2(g3554), .QN(n15007) );
  NOR2X0 U15461 ( .IN1(n15008), .IN2(n15009), .QN(n15006) );
  AND2X1 U15462 ( .IN1(n3765), .IN2(n4003), .Q(n15009) );
  NOR2X0 U15463 ( .IN1(n4003), .IN2(n15010), .QN(n15008) );
  NAND2X0 U15464 ( .IN1(n10369), .IN2(g3550), .QN(n15010) );
  NAND2X0 U15465 ( .IN1(n15011), .IN2(n15012), .QN(g30416) );
  NAND2X0 U15466 ( .IN1(n10509), .IN2(g3546), .QN(n15012) );
  NOR2X0 U15467 ( .IN1(n15013), .IN2(n15014), .QN(n15011) );
  AND2X1 U15468 ( .IN1(n3765), .IN2(n4005), .Q(n15014) );
  NOR2X0 U15469 ( .IN1(n4005), .IN2(n15015), .QN(n15013) );
  NAND2X0 U15470 ( .IN1(n10369), .IN2(g3542), .QN(n15015) );
  NAND2X0 U15471 ( .IN1(n15016), .IN2(n15017), .QN(g30415) );
  NAND2X0 U15472 ( .IN1(n10509), .IN2(g3530), .QN(n15017) );
  NOR2X0 U15473 ( .IN1(n15018), .IN2(n15019), .QN(n15016) );
  AND2X1 U15474 ( .IN1(n3765), .IN2(n4007), .Q(n15019) );
  NOR2X0 U15475 ( .IN1(n4007), .IN2(n15020), .QN(n15018) );
  NAND2X0 U15476 ( .IN1(n10368), .IN2(g3538), .QN(n15020) );
  NOR2X0 U15477 ( .IN1(g3506), .IN2(n13574), .QN(g30414) );
  NAND2X0 U15478 ( .IN1(n15021), .IN2(n5645), .QN(n13574) );
  NOR2X0 U15479 ( .IN1(n10463), .IN2(n13578), .QN(n15021) );
  INVX0 U15480 ( .INP(n13564), .ZN(n13578) );
  NAND2X0 U15481 ( .IN1(n14518), .IN2(n3799), .QN(n13564) );
  NOR2X0 U15482 ( .IN1(n5340), .IN2(g4087), .QN(n14518) );
  NAND2X0 U15483 ( .IN1(n15022), .IN2(n15023), .QN(g30413) );
  NAND2X0 U15484 ( .IN1(test_so84), .IN2(n10515), .QN(n15023) );
  NOR2X0 U15485 ( .IN1(n15024), .IN2(n15025), .QN(n15022) );
  NOR2X0 U15486 ( .IN1(n15026), .IN2(n14160), .QN(n15025) );
  NOR2X0 U15487 ( .IN1(n9791), .IN2(n15027), .QN(n15024) );
  NAND2X0 U15488 ( .IN1(n15028), .IN2(n15029), .QN(g30412) );
  NAND2X0 U15489 ( .IN1(n15030), .IN2(n3765), .QN(n15029) );
  NOR2X0 U15490 ( .IN1(n15031), .IN2(n15032), .QN(n15028) );
  NOR2X0 U15491 ( .IN1(n9970), .IN2(n10324), .QN(n15032) );
  NOR2X0 U15492 ( .IN1(n10467), .IN2(n15033), .QN(n15031) );
  OR2X1 U15493 ( .IN1(n15030), .IN2(n10007), .Q(n15033) );
  NOR2X0 U15494 ( .IN1(n364), .IN2(n5652), .QN(n15030) );
  NAND2X0 U15495 ( .IN1(n15034), .IN2(n15035), .QN(g30411) );
  NAND2X0 U15496 ( .IN1(n13591), .IN2(n3765), .QN(n15035) );
  NOR2X0 U15497 ( .IN1(n15036), .IN2(n15037), .QN(n15034) );
  NOR2X0 U15498 ( .IN1(n9867), .IN2(n10325), .QN(n15037) );
  NOR2X0 U15499 ( .IN1(n10465), .IN2(n15038), .QN(n15036) );
  OR2X1 U15500 ( .IN1(n13591), .IN2(n9972), .Q(n15038) );
  NOR2X0 U15501 ( .IN1(n4020), .IN2(n5652), .QN(n13591) );
  NAND2X0 U15502 ( .IN1(n15039), .IN2(n15040), .QN(g30410) );
  OR2X1 U15503 ( .IN1(n15041), .IN2(n14160), .Q(n15040) );
  NOR2X0 U15504 ( .IN1(n15042), .IN2(n15043), .QN(n15039) );
  NOR2X0 U15505 ( .IN1(n9792), .IN2(n10325), .QN(n15043) );
  NOR2X0 U15506 ( .IN1(n10468), .IN2(n15044), .QN(n15042) );
  NAND2X0 U15507 ( .IN1(test_so88), .IN2(n15041), .QN(n15044) );
  NAND2X0 U15508 ( .IN1(n15045), .IN2(g3167), .QN(n15041) );
  NAND2X0 U15509 ( .IN1(n15046), .IN2(n15047), .QN(g30409) );
  NAND2X0 U15510 ( .IN1(n4015), .IN2(n15048), .QN(n15047) );
  NOR2X0 U15511 ( .IN1(n15049), .IN2(n15050), .QN(n15046) );
  NOR2X0 U15512 ( .IN1(n10466), .IN2(n15051), .QN(n15050) );
  NAND2X0 U15513 ( .IN1(test_so84), .IN2(n15052), .QN(n15051) );
  NAND2X0 U15514 ( .IN1(n13601), .IN2(n15048), .QN(n15052) );
  NOR2X0 U15515 ( .IN1(n9843), .IN2(n10325), .QN(n15049) );
  NAND2X0 U15516 ( .IN1(n15053), .IN2(n15054), .QN(g30408) );
  NAND2X0 U15517 ( .IN1(n4015), .IN2(n13592), .QN(n15054) );
  NOR2X0 U15518 ( .IN1(n15055), .IN2(n15056), .QN(n15053) );
  NOR2X0 U15519 ( .IN1(n10466), .IN2(n15057), .QN(n15056) );
  NAND2X0 U15520 ( .IN1(n15058), .IN2(g3255), .QN(n15057) );
  NAND2X0 U15521 ( .IN1(n13601), .IN2(n13592), .QN(n15058) );
  NOR2X0 U15522 ( .IN1(n9968), .IN2(n10325), .QN(n15055) );
  NAND2X0 U15523 ( .IN1(n15059), .IN2(n15060), .QN(g30407) );
  NAND2X0 U15524 ( .IN1(n4015), .IN2(n15061), .QN(n15060) );
  NOR2X0 U15525 ( .IN1(n15062), .IN2(n15063), .QN(n15059) );
  NOR2X0 U15526 ( .IN1(n10466), .IN2(n15064), .QN(n15063) );
  NAND2X0 U15527 ( .IN1(n15065), .IN2(g3251), .QN(n15064) );
  NAND2X0 U15528 ( .IN1(n13601), .IN2(n15061), .QN(n15065) );
  NOR2X0 U15529 ( .IN1(n9882), .IN2(n10325), .QN(n15062) );
  NAND2X0 U15530 ( .IN1(n15066), .IN2(n15067), .QN(g30406) );
  NAND2X0 U15531 ( .IN1(n4015), .IN2(n15045), .QN(n15067) );
  NOR2X0 U15532 ( .IN1(n15068), .IN2(n15069), .QN(n15066) );
  NOR2X0 U15533 ( .IN1(n10468), .IN2(n15070), .QN(n15069) );
  NAND2X0 U15534 ( .IN1(n15071), .IN2(g3247), .QN(n15070) );
  NAND2X0 U15535 ( .IN1(n13601), .IN2(n15045), .QN(n15071) );
  INVX0 U15536 ( .INP(n3500), .ZN(n13601) );
  NAND2X0 U15537 ( .IN1(g3155), .IN2(g3161), .QN(n3500) );
  NOR2X0 U15538 ( .IN1(n9942), .IN2(n10325), .QN(n15068) );
  NAND2X0 U15539 ( .IN1(n15072), .IN2(n15073), .QN(g30405) );
  NAND2X0 U15540 ( .IN1(n4022), .IN2(n15048), .QN(n15073) );
  NOR2X0 U15541 ( .IN1(n15074), .IN2(n15075), .QN(n15072) );
  NOR2X0 U15542 ( .IN1(n10466), .IN2(n15076), .QN(n15075) );
  NAND2X0 U15543 ( .IN1(n15077), .IN2(g3243), .QN(n15076) );
  NAND2X0 U15544 ( .IN1(n15078), .IN2(n15048), .QN(n15077) );
  NOR2X0 U15545 ( .IN1(n9844), .IN2(n10325), .QN(n15074) );
  NAND2X0 U15546 ( .IN1(n15079), .IN2(n15080), .QN(g30404) );
  NAND2X0 U15547 ( .IN1(n4022), .IN2(n13592), .QN(n15080) );
  NOR2X0 U15548 ( .IN1(n15081), .IN2(n15082), .QN(n15079) );
  NOR2X0 U15549 ( .IN1(n10466), .IN2(n15083), .QN(n15082) );
  NAND2X0 U15550 ( .IN1(n15084), .IN2(g3239), .QN(n15083) );
  NAND2X0 U15551 ( .IN1(n15078), .IN2(n13592), .QN(n15084) );
  NOR2X0 U15552 ( .IN1(n9918), .IN2(n10326), .QN(n15081) );
  NAND2X0 U15553 ( .IN1(n15085), .IN2(n15086), .QN(g30403) );
  NAND2X0 U15554 ( .IN1(n4022), .IN2(n15061), .QN(n15086) );
  NOR2X0 U15555 ( .IN1(n15087), .IN2(n15088), .QN(n15085) );
  NOR2X0 U15556 ( .IN1(n10466), .IN2(n15089), .QN(n15088) );
  NAND2X0 U15557 ( .IN1(n15090), .IN2(g3235), .QN(n15089) );
  NAND2X0 U15558 ( .IN1(n15078), .IN2(n15061), .QN(n15090) );
  NOR2X0 U15559 ( .IN1(n9836), .IN2(n10326), .QN(n15087) );
  NAND2X0 U15560 ( .IN1(n15091), .IN2(n15092), .QN(g30402) );
  NAND2X0 U15561 ( .IN1(n4022), .IN2(n15045), .QN(n15092) );
  NOR2X0 U15562 ( .IN1(n15093), .IN2(n15094), .QN(n15091) );
  NOR2X0 U15563 ( .IN1(n10466), .IN2(n15095), .QN(n15094) );
  NAND2X0 U15564 ( .IN1(n15096), .IN2(g3231), .QN(n15095) );
  NAND2X0 U15565 ( .IN1(n15078), .IN2(n15045), .QN(n15096) );
  INVX0 U15566 ( .INP(n3502), .ZN(n15078) );
  NAND2X0 U15567 ( .IN1(n5366), .IN2(g3161), .QN(n3502) );
  NOR2X0 U15568 ( .IN1(n9793), .IN2(n10326), .QN(n15093) );
  NAND2X0 U15569 ( .IN1(n15097), .IN2(n15098), .QN(g30401) );
  NAND2X0 U15570 ( .IN1(n4027), .IN2(n15048), .QN(n15098) );
  NOR2X0 U15571 ( .IN1(n15099), .IN2(n15100), .QN(n15097) );
  NOR2X0 U15572 ( .IN1(n10466), .IN2(n15101), .QN(n15100) );
  NAND2X0 U15573 ( .IN1(n15102), .IN2(g3227), .QN(n15101) );
  NAND2X0 U15574 ( .IN1(n13607), .IN2(n15048), .QN(n15102) );
  NOR2X0 U15575 ( .IN1(n9919), .IN2(n10326), .QN(n15099) );
  NAND2X0 U15576 ( .IN1(n15103), .IN2(n15104), .QN(g30400) );
  NAND2X0 U15577 ( .IN1(n4027), .IN2(n13592), .QN(n15104) );
  NOR2X0 U15578 ( .IN1(n15105), .IN2(n15106), .QN(n15103) );
  NOR2X0 U15579 ( .IN1(n10468), .IN2(n15107), .QN(n15106) );
  NAND2X0 U15580 ( .IN1(n15108), .IN2(g3223), .QN(n15107) );
  NAND2X0 U15581 ( .IN1(n13607), .IN2(n13592), .QN(n15108) );
  INVX0 U15582 ( .INP(n364), .ZN(n13592) );
  NAND2X0 U15583 ( .IN1(n5603), .IN2(g3179), .QN(n364) );
  NOR2X0 U15584 ( .IN1(n10009), .IN2(n10326), .QN(n15105) );
  NAND2X0 U15585 ( .IN1(n15109), .IN2(n15110), .QN(g30399) );
  NAND2X0 U15586 ( .IN1(n4027), .IN2(n15061), .QN(n15110) );
  NOR2X0 U15587 ( .IN1(n15111), .IN2(n15112), .QN(n15109) );
  NOR2X0 U15588 ( .IN1(n10468), .IN2(n15113), .QN(n15112) );
  NAND2X0 U15589 ( .IN1(n15114), .IN2(g3219), .QN(n15113) );
  NAND2X0 U15590 ( .IN1(n13607), .IN2(n15061), .QN(n15114) );
  INVX0 U15591 ( .INP(n4020), .ZN(n15061) );
  NAND2X0 U15592 ( .IN1(n5390), .IN2(g3171), .QN(n4020) );
  NOR2X0 U15593 ( .IN1(n9794), .IN2(n10326), .QN(n15111) );
  NAND2X0 U15594 ( .IN1(n15115), .IN2(n15116), .QN(g30398) );
  NAND2X0 U15595 ( .IN1(n4027), .IN2(n15045), .QN(n15116) );
  NOR2X0 U15596 ( .IN1(n15117), .IN2(n15118), .QN(n15115) );
  NOR2X0 U15597 ( .IN1(n10467), .IN2(n15119), .QN(n15118) );
  NAND2X0 U15598 ( .IN1(n15120), .IN2(g3215), .QN(n15119) );
  NAND2X0 U15599 ( .IN1(n13607), .IN2(n15045), .QN(n15120) );
  INVX0 U15600 ( .INP(n4014), .ZN(n15045) );
  NAND2X0 U15601 ( .IN1(n5603), .IN2(n5390), .QN(n4014) );
  INVX0 U15602 ( .INP(n3501), .ZN(n13607) );
  NAND2X0 U15603 ( .IN1(n10062), .IN2(g3155), .QN(n3501) );
  NOR2X0 U15604 ( .IN1(n9950), .IN2(n10326), .QN(n15117) );
  NAND2X0 U15605 ( .IN1(n15121), .IN2(n15122), .QN(g30397) );
  NAND2X0 U15606 ( .IN1(n10510), .IN2(g3211), .QN(n15122) );
  NOR2X0 U15607 ( .IN1(n15123), .IN2(n15124), .QN(n15121) );
  AND2X1 U15608 ( .IN1(n3765), .IN2(n4032), .Q(n15124) );
  NOR2X0 U15609 ( .IN1(n4032), .IN2(n15125), .QN(n15123) );
  NAND2X0 U15610 ( .IN1(n10368), .IN2(g3207), .QN(n15125) );
  NAND2X0 U15611 ( .IN1(n15126), .IN2(n15127), .QN(g30396) );
  OR2X1 U15612 ( .IN1(n10309), .IN2(n9972), .Q(n15127) );
  NOR2X0 U15613 ( .IN1(n15128), .IN2(n15129), .QN(n15126) );
  AND2X1 U15614 ( .IN1(n3765), .IN2(n4035), .Q(n15129) );
  NOR2X0 U15615 ( .IN1(n4035), .IN2(n15130), .QN(n15128) );
  NAND2X0 U15616 ( .IN1(n10368), .IN2(g3199), .QN(n15130) );
  NAND2X0 U15617 ( .IN1(n15131), .IN2(n15132), .QN(g30395) );
  NAND2X0 U15618 ( .IN1(test_so88), .IN2(n10516), .QN(n15132) );
  NOR2X0 U15619 ( .IN1(n15133), .IN2(n15134), .QN(n15131) );
  AND2X1 U15620 ( .IN1(n3765), .IN2(n4037), .Q(n15134) );
  NOR2X0 U15621 ( .IN1(n4037), .IN2(n15135), .QN(n15133) );
  NAND2X0 U15622 ( .IN1(n10368), .IN2(g3191), .QN(n15135) );
  NAND2X0 U15623 ( .IN1(n15136), .IN2(n15137), .QN(g30394) );
  NAND2X0 U15624 ( .IN1(n10510), .IN2(g3179), .QN(n15137) );
  NOR2X0 U15625 ( .IN1(n15138), .IN2(n15139), .QN(n15136) );
  AND2X1 U15626 ( .IN1(n3765), .IN2(n4039), .Q(n15139) );
  NOR2X0 U15627 ( .IN1(n4039), .IN2(n15140), .QN(n15138) );
  NAND2X0 U15628 ( .IN1(n10367), .IN2(g3187), .QN(n15140) );
  NOR2X0 U15629 ( .IN1(n13602), .IN2(n15141), .QN(g30393) );
  NAND2X0 U15630 ( .IN1(n5366), .IN2(n10390), .QN(n15141) );
  NAND2X0 U15631 ( .IN1(n5652), .IN2(n13598), .QN(n13602) );
  NAND2X0 U15632 ( .IN1(n3799), .IN2(n12615), .QN(n13598) );
  NAND2X0 U15633 ( .IN1(n15142), .IN2(n15143), .QN(g30392) );
  NAND2X0 U15634 ( .IN1(n10510), .IN2(g2803), .QN(n15143) );
  NAND2X0 U15635 ( .IN1(n15144), .IN2(n15145), .QN(g30391) );
  NAND2X0 U15636 ( .IN1(n10510), .IN2(g2771), .QN(n15145) );
  NAND2X0 U15637 ( .IN1(n15142), .IN2(n15146), .QN(g30390) );
  NAND2X0 U15638 ( .IN1(g2834), .IN2(n10516), .QN(n15146) );
  NAND2X0 U15639 ( .IN1(n15147), .IN2(n10390), .QN(n15142) );
  NAND2X0 U15640 ( .IN1(n15148), .IN2(n15149), .QN(n15147) );
  NAND2X0 U15641 ( .IN1(n15150), .IN2(n15151), .QN(n15149) );
  NOR2X0 U15642 ( .IN1(n15152), .IN2(n15153), .QN(n15150) );
  NAND2X0 U15643 ( .IN1(n15154), .IN2(n15155), .QN(n15153) );
  NAND2X0 U15644 ( .IN1(n9941), .IN2(n15156), .QN(n15155) );
  NAND2X0 U15645 ( .IN1(n9826), .IN2(n15157), .QN(n15154) );
  NAND2X0 U15646 ( .IN1(n15158), .IN2(n15159), .QN(n15152) );
  NAND2X0 U15647 ( .IN1(n9822), .IN2(n15160), .QN(n15159) );
  NAND2X0 U15648 ( .IN1(n9832), .IN2(n15161), .QN(n15158) );
  NAND2X0 U15649 ( .IN1(n15162), .IN2(n15163), .QN(n15148) );
  NOR2X0 U15650 ( .IN1(n15164), .IN2(n15165), .QN(n15162) );
  NAND2X0 U15651 ( .IN1(n15166), .IN2(n15167), .QN(n15165) );
  NAND2X0 U15652 ( .IN1(n15156), .IN2(g2815), .QN(n15167) );
  NAND2X0 U15653 ( .IN1(n15157), .IN2(g2807), .QN(n15166) );
  NAND2X0 U15654 ( .IN1(n15168), .IN2(n15169), .QN(n15164) );
  NAND2X0 U15655 ( .IN1(n15160), .IN2(g2803), .QN(n15169) );
  NAND2X0 U15656 ( .IN1(n15161), .IN2(g2819), .QN(n15168) );
  NAND2X0 U15657 ( .IN1(n15144), .IN2(n15170), .QN(g30389) );
  NAND2X0 U15658 ( .IN1(g2831), .IN2(n10515), .QN(n15170) );
  NAND2X0 U15659 ( .IN1(n15171), .IN2(n10390), .QN(n15144) );
  NAND2X0 U15660 ( .IN1(n15172), .IN2(n15173), .QN(n15171) );
  NAND2X0 U15661 ( .IN1(n15174), .IN2(n15151), .QN(n15173) );
  NOR2X0 U15662 ( .IN1(n15175), .IN2(n15176), .QN(n15174) );
  NAND2X0 U15663 ( .IN1(n15177), .IN2(n15178), .QN(n15176) );
  NAND2X0 U15664 ( .IN1(n15156), .IN2(n10151), .QN(n15178) );
  NAND2X0 U15665 ( .IN1(n9824), .IN2(n15157), .QN(n15177) );
  NAND2X0 U15666 ( .IN1(n15179), .IN2(n15180), .QN(n15175) );
  NAND2X0 U15667 ( .IN1(n9828), .IN2(n15160), .QN(n15180) );
  NAND2X0 U15668 ( .IN1(n9829), .IN2(n15161), .QN(n15179) );
  NAND2X0 U15669 ( .IN1(n15181), .IN2(n15163), .QN(n15172) );
  INVX0 U15670 ( .INP(n15151), .ZN(n15163) );
  NAND2X0 U15671 ( .IN1(n15182), .IN2(n5600), .QN(n15151) );
  NOR2X0 U15672 ( .IN1(n11658), .IN2(n13884), .QN(n15182) );
  NAND2X0 U15673 ( .IN1(n15183), .IN2(n5516), .QN(n13884) );
  NOR2X0 U15674 ( .IN1(test_so30), .IN2(g2741), .QN(n15183) );
  NOR2X0 U15675 ( .IN1(n15184), .IN2(n15185), .QN(n15181) );
  NAND2X0 U15676 ( .IN1(n15186), .IN2(n15187), .QN(n15185) );
  NAND2X0 U15677 ( .IN1(n15156), .IN2(g2783), .QN(n15187) );
  NAND2X0 U15678 ( .IN1(n15157), .IN2(g2775), .QN(n15186) );
  INVX0 U15679 ( .INP(n4411), .ZN(n15157) );
  NAND2X0 U15680 ( .IN1(n15188), .IN2(n15189), .QN(n15184) );
  NAND2X0 U15681 ( .IN1(n15160), .IN2(g2771), .QN(n15189) );
  NAND2X0 U15682 ( .IN1(n15161), .IN2(g2787), .QN(n15188) );
  NAND2X0 U15683 ( .IN1(n15190), .IN2(n15191), .QN(g30388) );
  NAND2X0 U15684 ( .IN1(n15192), .IN2(n3730), .QN(n15191) );
  XOR2X1 U15685 ( .IN1(n3506), .IN2(n5349), .Q(n15192) );
  NAND2X0 U15686 ( .IN1(n15193), .IN2(g2735), .QN(n3506) );
  NAND2X0 U15687 ( .IN1(n10510), .IN2(g2735), .QN(n15190) );
  NAND2X0 U15688 ( .IN1(n15194), .IN2(n15195), .QN(g30387) );
  OR2X1 U15689 ( .IN1(n15196), .IN2(n18484), .Q(n15195) );
  NOR2X0 U15690 ( .IN1(n15197), .IN2(n15198), .QN(n15194) );
  NOR2X0 U15691 ( .IN1(g2681), .IN2(n15199), .QN(n15198) );
  NAND2X0 U15692 ( .IN1(n15200), .IN2(n5457), .QN(n15199) );
  NOR2X0 U15693 ( .IN1(n5777), .IN2(n15201), .QN(n15197) );
  NOR2X0 U15694 ( .IN1(n10469), .IN2(n15202), .QN(n15201) );
  NOR2X0 U15695 ( .IN1(n5457), .IN2(n15203), .QN(n15202) );
  NAND2X0 U15696 ( .IN1(n15204), .IN2(n15205), .QN(g30386) );
  OR2X1 U15697 ( .IN1(n15196), .IN2(n5777), .Q(n15205) );
  NAND2X0 U15698 ( .IN1(n15196), .IN2(g2675), .QN(n15204) );
  NAND2X0 U15699 ( .IN1(n15206), .IN2(n15207), .QN(g30385) );
  NAND2X0 U15700 ( .IN1(n10510), .IN2(g2657), .QN(n15207) );
  NOR2X0 U15701 ( .IN1(n15208), .IN2(n15209), .QN(n15206) );
  NOR2X0 U15702 ( .IN1(g2661), .IN2(n15210), .QN(n15209) );
  NOR2X0 U15703 ( .IN1(n5418), .IN2(n15196), .QN(n15208) );
  NAND2X0 U15704 ( .IN1(n15203), .IN2(n10390), .QN(n15196) );
  NAND2X0 U15705 ( .IN1(n15211), .IN2(n15212), .QN(g30384) );
  NAND2X0 U15706 ( .IN1(n10510), .IN2(g2652), .QN(n15212) );
  NOR2X0 U15707 ( .IN1(n15213), .IN2(n15214), .QN(n15211) );
  NOR2X0 U15708 ( .IN1(n5316), .IN2(n15215), .QN(n15214) );
  NOR2X0 U15709 ( .IN1(n15216), .IN2(n13640), .QN(n15215) );
  INVX0 U15710 ( .INP(n13626), .ZN(n13640) );
  NOR2X0 U15711 ( .IN1(n10484), .IN2(n10112), .QN(n15216) );
  NOR2X0 U15712 ( .IN1(n13645), .IN2(n15217), .QN(n15213) );
  NAND2X0 U15713 ( .IN1(n333), .IN2(n15218), .QN(n15217) );
  XOR2X1 U15714 ( .IN1(n9833), .IN2(n9660), .Q(n15218) );
  INVX0 U15715 ( .INP(n13627), .ZN(n333) );
  NAND2X0 U15716 ( .IN1(n15219), .IN2(n15220), .QN(g30383) );
  NAND2X0 U15717 ( .IN1(test_so66), .IN2(n10516), .QN(n15220) );
  NAND2X0 U15718 ( .IN1(n15221), .IN2(n10390), .QN(n15219) );
  NAND2X0 U15719 ( .IN1(n15222), .IN2(n15223), .QN(n15221) );
  NAND2X0 U15720 ( .IN1(test_so34), .IN2(n15224), .QN(n15223) );
  NAND2X0 U15721 ( .IN1(n15225), .IN2(n15226), .QN(n15222) );
  NAND2X0 U15722 ( .IN1(n5351), .IN2(g2599), .QN(n15226) );
  INVX0 U15723 ( .INP(n15224), .ZN(n15225) );
  NAND2X0 U15724 ( .IN1(n15227), .IN2(n5508), .QN(n15224) );
  NOR2X0 U15725 ( .IN1(n10042), .IN2(n13620), .QN(n15227) );
  NAND2X0 U15726 ( .IN1(n15228), .IN2(n15229), .QN(g30382) );
  OR2X1 U15727 ( .IN1(n15230), .IN2(n18481), .Q(n15229) );
  NOR2X0 U15728 ( .IN1(n15231), .IN2(n15232), .QN(n15228) );
  NOR2X0 U15729 ( .IN1(g2547), .IN2(n15233), .QN(n15232) );
  NAND2X0 U15730 ( .IN1(n15234), .IN2(n5461), .QN(n15233) );
  NOR2X0 U15731 ( .IN1(n5782), .IN2(n15235), .QN(n15231) );
  NOR2X0 U15732 ( .IN1(n10484), .IN2(n15236), .QN(n15235) );
  NOR2X0 U15733 ( .IN1(n5461), .IN2(n15237), .QN(n15236) );
  NAND2X0 U15734 ( .IN1(n15238), .IN2(n15239), .QN(g30381) );
  OR2X1 U15735 ( .IN1(n15230), .IN2(n5782), .Q(n15239) );
  NAND2X0 U15736 ( .IN1(n15230), .IN2(g2541), .QN(n15238) );
  NAND2X0 U15737 ( .IN1(n15240), .IN2(n15241), .QN(g30380) );
  NAND2X0 U15738 ( .IN1(n10510), .IN2(g2523), .QN(n15241) );
  NOR2X0 U15739 ( .IN1(n15242), .IN2(n15243), .QN(n15240) );
  NOR2X0 U15740 ( .IN1(g2527), .IN2(n15244), .QN(n15243) );
  NOR2X0 U15741 ( .IN1(n5420), .IN2(n15230), .QN(n15242) );
  NAND2X0 U15742 ( .IN1(n15237), .IN2(n10391), .QN(n15230) );
  NAND2X0 U15743 ( .IN1(n15245), .IN2(n15246), .QN(g30379) );
  NAND2X0 U15744 ( .IN1(n10510), .IN2(g2518), .QN(n15246) );
  NOR2X0 U15745 ( .IN1(n15247), .IN2(n15248), .QN(n15245) );
  NOR2X0 U15746 ( .IN1(n5281), .IN2(n15249), .QN(n15248) );
  NOR2X0 U15747 ( .IN1(n15250), .IN2(n13676), .QN(n15249) );
  INVX0 U15748 ( .INP(n13661), .ZN(n13676) );
  NOR2X0 U15749 ( .IN1(n10484), .IN2(n10117), .QN(n15250) );
  NOR2X0 U15750 ( .IN1(n13681), .IN2(n15251), .QN(n15247) );
  NAND2X0 U15751 ( .IN1(n408), .IN2(n15252), .QN(n15251) );
  XOR2X1 U15752 ( .IN1(n9831), .IN2(n9657), .Q(n15252) );
  INVX0 U15753 ( .INP(n13662), .ZN(n408) );
  NAND2X0 U15754 ( .IN1(n15253), .IN2(n15254), .QN(g30378) );
  NAND2X0 U15755 ( .IN1(n10510), .IN2(g2441), .QN(n15254) );
  NAND2X0 U15756 ( .IN1(n15255), .IN2(n10391), .QN(n15253) );
  NAND2X0 U15757 ( .IN1(n15256), .IN2(n15257), .QN(n15255) );
  NAND2X0 U15758 ( .IN1(n15258), .IN2(g2461), .QN(n15257) );
  NAND2X0 U15759 ( .IN1(n15259), .IN2(n15260), .QN(n15256) );
  NAND2X0 U15760 ( .IN1(g2465), .IN2(n10131), .QN(n15260) );
  INVX0 U15761 ( .INP(n15258), .ZN(n15259) );
  NAND2X0 U15762 ( .IN1(n15261), .IN2(n5509), .QN(n15258) );
  NOR2X0 U15763 ( .IN1(n10043), .IN2(n13655), .QN(n15261) );
  NAND2X0 U15764 ( .IN1(n15262), .IN2(n15263), .QN(g30377) );
  OR2X1 U15765 ( .IN1(n15264), .IN2(n18483), .Q(n15263) );
  NOR2X0 U15766 ( .IN1(n15265), .IN2(n15266), .QN(n15262) );
  NOR2X0 U15767 ( .IN1(test_so89), .IN2(n15267), .QN(n15266) );
  NAND2X0 U15768 ( .IN1(n15268), .IN2(n5459), .QN(n15267) );
  NOR2X0 U15769 ( .IN1(n15269), .IN2(n10143), .QN(n15265) );
  NOR2X0 U15770 ( .IN1(n10484), .IN2(n15270), .QN(n15269) );
  NOR2X0 U15771 ( .IN1(n5459), .IN2(n15271), .QN(n15270) );
  NAND2X0 U15772 ( .IN1(n15272), .IN2(n15273), .QN(g30376) );
  OR2X1 U15773 ( .IN1(n10143), .IN2(n15264), .Q(n15273) );
  NAND2X0 U15774 ( .IN1(n15264), .IN2(g2407), .QN(n15272) );
  NAND2X0 U15775 ( .IN1(n15274), .IN2(n15275), .QN(g30375) );
  NAND2X0 U15776 ( .IN1(n10514), .IN2(g2389), .QN(n15275) );
  NOR2X0 U15777 ( .IN1(n15276), .IN2(n15277), .QN(n15274) );
  NOR2X0 U15778 ( .IN1(g2393), .IN2(n15278), .QN(n15277) );
  NOR2X0 U15779 ( .IN1(n5421), .IN2(n15264), .QN(n15276) );
  NAND2X0 U15780 ( .IN1(n15271), .IN2(n10391), .QN(n15264) );
  NAND2X0 U15781 ( .IN1(n15279), .IN2(n15280), .QN(g30374) );
  NAND2X0 U15782 ( .IN1(n10514), .IN2(g2384), .QN(n15280) );
  NOR2X0 U15783 ( .IN1(n15281), .IN2(n15282), .QN(n15279) );
  NOR2X0 U15784 ( .IN1(n5631), .IN2(n15283), .QN(n15282) );
  NOR2X0 U15785 ( .IN1(n15284), .IN2(n13712), .QN(n15283) );
  INVX0 U15786 ( .INP(n13697), .ZN(n13712) );
  NOR2X0 U15787 ( .IN1(n10484), .IN2(n401), .QN(n15284) );
  NOR2X0 U15788 ( .IN1(n13717), .IN2(n15285), .QN(n15281) );
  NAND2X0 U15789 ( .IN1(n380), .IN2(n15286), .QN(n15285) );
  XOR2X1 U15790 ( .IN1(n9825), .IN2(n9656), .Q(n15286) );
  INVX0 U15791 ( .INP(n13698), .ZN(n380) );
  NAND2X0 U15792 ( .IN1(n15287), .IN2(n15288), .QN(g30373) );
  NAND2X0 U15793 ( .IN1(n10514), .IN2(g2307), .QN(n15288) );
  NAND2X0 U15794 ( .IN1(n15289), .IN2(n10391), .QN(n15287) );
  NAND2X0 U15795 ( .IN1(n15290), .IN2(n15291), .QN(n15289) );
  NAND2X0 U15796 ( .IN1(n15292), .IN2(g2327), .QN(n15291) );
  NAND2X0 U15797 ( .IN1(n15293), .IN2(n15294), .QN(n15290) );
  NAND2X0 U15798 ( .IN1(n5353), .IN2(g2331), .QN(n15294) );
  INVX0 U15799 ( .INP(n15292), .ZN(n15293) );
  NAND2X0 U15800 ( .IN1(n15295), .IN2(n5511), .QN(n15292) );
  NOR2X0 U15801 ( .IN1(n10126), .IN2(n13691), .QN(n15295) );
  NAND2X0 U15802 ( .IN1(n15296), .IN2(n15297), .QN(g30372) );
  OR2X1 U15803 ( .IN1(n15298), .IN2(n18482), .Q(n15297) );
  NOR2X0 U15804 ( .IN1(n15299), .IN2(n15300), .QN(n15296) );
  NOR2X0 U15805 ( .IN1(g2279), .IN2(n15301), .QN(n15300) );
  NAND2X0 U15806 ( .IN1(n15302), .IN2(n5458), .QN(n15301) );
  NOR2X0 U15807 ( .IN1(n5778), .IN2(n15303), .QN(n15299) );
  NOR2X0 U15808 ( .IN1(n10484), .IN2(n15304), .QN(n15303) );
  NOR2X0 U15809 ( .IN1(n5458), .IN2(n15305), .QN(n15304) );
  NAND2X0 U15810 ( .IN1(n15306), .IN2(n15307), .QN(g30371) );
  OR2X1 U15811 ( .IN1(n15298), .IN2(n5778), .Q(n15307) );
  NAND2X0 U15812 ( .IN1(n15298), .IN2(g2273), .QN(n15306) );
  NAND2X0 U15813 ( .IN1(n15308), .IN2(n15309), .QN(g30370) );
  NAND2X0 U15814 ( .IN1(n10514), .IN2(g2255), .QN(n15309) );
  NOR2X0 U15815 ( .IN1(n15310), .IN2(n15311), .QN(n15308) );
  NOR2X0 U15816 ( .IN1(g2259), .IN2(n15312), .QN(n15311) );
  NOR2X0 U15817 ( .IN1(n5419), .IN2(n15298), .QN(n15310) );
  NAND2X0 U15818 ( .IN1(n15305), .IN2(n10391), .QN(n15298) );
  NAND2X0 U15819 ( .IN1(n15313), .IN2(n15314), .QN(g30369) );
  NAND2X0 U15820 ( .IN1(n10514), .IN2(g2250), .QN(n15314) );
  NOR2X0 U15821 ( .IN1(n15315), .IN2(n15316), .QN(n15313) );
  NOR2X0 U15822 ( .IN1(n5414), .IN2(n15317), .QN(n15316) );
  NOR2X0 U15823 ( .IN1(n15318), .IN2(n13748), .QN(n15317) );
  INVX0 U15824 ( .INP(n13733), .ZN(n13748) );
  NOR2X0 U15825 ( .IN1(n10484), .IN2(n10119), .QN(n15318) );
  NOR2X0 U15826 ( .IN1(n13753), .IN2(n15319), .QN(n15315) );
  NAND2X0 U15827 ( .IN1(n780), .IN2(n15320), .QN(n15319) );
  XOR2X1 U15828 ( .IN1(n9821), .IN2(n9659), .Q(n15320) );
  INVX0 U15829 ( .INP(n13734), .ZN(n780) );
  NAND2X0 U15830 ( .IN1(n15321), .IN2(n15322), .QN(g30368) );
  NAND2X0 U15831 ( .IN1(n10513), .IN2(g2173), .QN(n15322) );
  NAND2X0 U15832 ( .IN1(n15323), .IN2(n10391), .QN(n15321) );
  NAND2X0 U15833 ( .IN1(n15324), .IN2(n15325), .QN(n15323) );
  NAND2X0 U15834 ( .IN1(n15326), .IN2(g2193), .QN(n15325) );
  NAND2X0 U15835 ( .IN1(n15327), .IN2(n15328), .QN(n15324) );
  NAND2X0 U15836 ( .IN1(n5356), .IN2(g2197), .QN(n15328) );
  INVX0 U15837 ( .INP(n15326), .ZN(n15327) );
  NAND2X0 U15838 ( .IN1(n15329), .IN2(n5512), .QN(n15326) );
  NOR2X0 U15839 ( .IN1(n10045), .IN2(n13727), .QN(n15329) );
  NAND2X0 U15840 ( .IN1(n15330), .IN2(n15331), .QN(g30367) );
  OR2X1 U15841 ( .IN1(n15332), .IN2(n5891), .Q(n15331) );
  NOR2X0 U15842 ( .IN1(n15333), .IN2(n15334), .QN(n15330) );
  NOR2X0 U15843 ( .IN1(g2122), .IN2(n15335), .QN(n15334) );
  NAND2X0 U15844 ( .IN1(n15336), .IN2(n5463), .QN(n15335) );
  NOR2X0 U15845 ( .IN1(n5784), .IN2(n15337), .QN(n15333) );
  NOR2X0 U15846 ( .IN1(n10484), .IN2(n15338), .QN(n15337) );
  NOR2X0 U15847 ( .IN1(n5463), .IN2(n15339), .QN(n15338) );
  NAND2X0 U15848 ( .IN1(n15340), .IN2(n15341), .QN(g30366) );
  OR2X1 U15849 ( .IN1(n15332), .IN2(n5784), .Q(n15341) );
  NAND2X0 U15850 ( .IN1(n15332), .IN2(g2116), .QN(n15340) );
  NAND2X0 U15851 ( .IN1(n15342), .IN2(n15343), .QN(g30365) );
  NAND2X0 U15852 ( .IN1(n10514), .IN2(g2098), .QN(n15343) );
  NOR2X0 U15853 ( .IN1(n15344), .IN2(n15345), .QN(n15342) );
  NOR2X0 U15854 ( .IN1(g2102), .IN2(n15346), .QN(n15345) );
  NOR2X0 U15855 ( .IN1(n5666), .IN2(n15332), .QN(n15344) );
  NAND2X0 U15856 ( .IN1(n15339), .IN2(n10391), .QN(n15332) );
  NAND2X0 U15857 ( .IN1(n15347), .IN2(n15348), .QN(g30364) );
  NAND2X0 U15858 ( .IN1(test_so78), .IN2(n10515), .QN(n15348) );
  NOR2X0 U15859 ( .IN1(n15349), .IN2(n15350), .QN(n15347) );
  NOR2X0 U15860 ( .IN1(n5280), .IN2(n15351), .QN(n15350) );
  NOR2X0 U15861 ( .IN1(n15352), .IN2(n13785), .QN(n15351) );
  INVX0 U15862 ( .INP(n13769), .ZN(n13785) );
  NOR2X0 U15863 ( .IN1(n10484), .IN2(n10120), .QN(n15352) );
  NOR2X0 U15864 ( .IN1(n15353), .IN2(n15354), .QN(n15349) );
  NAND2X0 U15865 ( .IN1(n10120), .IN2(n787), .QN(n15354) );
  INVX0 U15866 ( .INP(n13770), .ZN(n787) );
  INVX0 U15867 ( .INP(n13790), .ZN(n10120) );
  XOR2X1 U15868 ( .IN1(test_so78), .IN2(n9655), .Q(n15353) );
  NAND2X0 U15869 ( .IN1(n15355), .IN2(n15356), .QN(g30363) );
  NAND2X0 U15870 ( .IN1(n10514), .IN2(g2016), .QN(n15356) );
  NAND2X0 U15871 ( .IN1(n15357), .IN2(n10391), .QN(n15355) );
  NAND2X0 U15872 ( .IN1(n15358), .IN2(n15359), .QN(n15357) );
  NAND2X0 U15873 ( .IN1(test_so59), .IN2(n15360), .QN(n15359) );
  NAND2X0 U15874 ( .IN1(n15361), .IN2(n15362), .QN(n15358) );
  NAND2X0 U15875 ( .IN1(n5355), .IN2(g2040), .QN(n15362) );
  INVX0 U15876 ( .INP(n15360), .ZN(n15361) );
  NAND2X0 U15877 ( .IN1(n15363), .IN2(n5507), .QN(n15360) );
  NOR2X0 U15878 ( .IN1(n10041), .IN2(n13763), .QN(n15363) );
  NAND2X0 U15879 ( .IN1(n15364), .IN2(n15365), .QN(g30362) );
  OR2X1 U15880 ( .IN1(n15366), .IN2(n5890), .Q(n15365) );
  NOR2X0 U15881 ( .IN1(n15367), .IN2(n15368), .QN(n15364) );
  NOR2X0 U15882 ( .IN1(g1988), .IN2(n15369), .QN(n15368) );
  NAND2X0 U15883 ( .IN1(n15370), .IN2(n5462), .QN(n15369) );
  NOR2X0 U15884 ( .IN1(n5783), .IN2(n15371), .QN(n15367) );
  NOR2X0 U15885 ( .IN1(n10484), .IN2(n15372), .QN(n15371) );
  NOR2X0 U15886 ( .IN1(n5462), .IN2(n15373), .QN(n15372) );
  NAND2X0 U15887 ( .IN1(n15374), .IN2(n15375), .QN(g30361) );
  OR2X1 U15888 ( .IN1(n15366), .IN2(n5783), .Q(n15375) );
  NAND2X0 U15889 ( .IN1(n15366), .IN2(g1982), .QN(n15374) );
  NAND2X0 U15890 ( .IN1(n15376), .IN2(n15377), .QN(g30360) );
  NAND2X0 U15891 ( .IN1(n10514), .IN2(g1964), .QN(n15377) );
  NOR2X0 U15892 ( .IN1(n15378), .IN2(n15379), .QN(n15376) );
  NOR2X0 U15893 ( .IN1(g1968), .IN2(n15380), .QN(n15379) );
  NOR2X0 U15894 ( .IN1(n5664), .IN2(n15366), .QN(n15378) );
  NAND2X0 U15895 ( .IN1(n15373), .IN2(n10391), .QN(n15366) );
  NAND2X0 U15896 ( .IN1(n15381), .IN2(n15382), .QN(g30359) );
  NAND2X0 U15897 ( .IN1(n10514), .IN2(g1959), .QN(n15382) );
  NOR2X0 U15898 ( .IN1(n15383), .IN2(n15384), .QN(n15381) );
  NOR2X0 U15899 ( .IN1(n5315), .IN2(n15385), .QN(n15384) );
  NOR2X0 U15900 ( .IN1(n15386), .IN2(n13822), .QN(n15385) );
  INVX0 U15901 ( .INP(n13806), .ZN(n13822) );
  NOR2X0 U15902 ( .IN1(n10484), .IN2(n10111), .QN(n15386) );
  NOR2X0 U15903 ( .IN1(n13827), .IN2(n15387), .QN(n15383) );
  NAND2X0 U15904 ( .IN1(n3611), .IN2(n15388), .QN(n15387) );
  XOR2X1 U15905 ( .IN1(n9830), .IN2(n9653), .Q(n15388) );
  INVX0 U15906 ( .INP(n13807), .ZN(n3611) );
  NAND2X0 U15907 ( .IN1(n15389), .IN2(n15390), .QN(g30358) );
  NAND2X0 U15908 ( .IN1(n10513), .IN2(g1882), .QN(n15390) );
  NAND2X0 U15909 ( .IN1(n15391), .IN2(n10391), .QN(n15389) );
  NAND2X0 U15910 ( .IN1(n15392), .IN2(n15393), .QN(n15391) );
  NAND2X0 U15911 ( .IN1(n15394), .IN2(g1902), .QN(n15393) );
  NAND2X0 U15912 ( .IN1(n15395), .IN2(n15396), .QN(n15392) );
  NAND2X0 U15913 ( .IN1(g1906), .IN2(n10137), .QN(n15396) );
  INVX0 U15914 ( .INP(n15394), .ZN(n15395) );
  NAND2X0 U15915 ( .IN1(n15397), .IN2(n5510), .QN(n15394) );
  NOR2X0 U15916 ( .IN1(n10044), .IN2(n13800), .QN(n15397) );
  NAND2X0 U15917 ( .IN1(n15398), .IN2(n15399), .QN(g30357) );
  OR2X1 U15918 ( .IN1(n15400), .IN2(n5892), .Q(n15399) );
  NOR2X0 U15919 ( .IN1(n15401), .IN2(n15402), .QN(n15398) );
  NOR2X0 U15920 ( .IN1(g1854), .IN2(n15403), .QN(n15402) );
  NAND2X0 U15921 ( .IN1(n15404), .IN2(n5464), .QN(n15403) );
  NOR2X0 U15922 ( .IN1(n5785), .IN2(n15405), .QN(n15401) );
  NOR2X0 U15923 ( .IN1(n10484), .IN2(n15406), .QN(n15405) );
  NOR2X0 U15924 ( .IN1(n5464), .IN2(n15407), .QN(n15406) );
  NAND2X0 U15925 ( .IN1(n15408), .IN2(n15409), .QN(g30356) );
  OR2X1 U15926 ( .IN1(n15400), .IN2(n5785), .Q(n15409) );
  NAND2X0 U15927 ( .IN1(n15400), .IN2(g1848), .QN(n15408) );
  NAND2X0 U15928 ( .IN1(n15410), .IN2(n15411), .QN(g30355) );
  OR2X1 U15929 ( .IN1(n10308), .IN2(n5413), .Q(n15411) );
  NOR2X0 U15930 ( .IN1(n15412), .IN2(n15413), .QN(n15410) );
  NOR2X0 U15931 ( .IN1(g1834), .IN2(n15414), .QN(n15413) );
  NOR2X0 U15932 ( .IN1(n5665), .IN2(n15400), .QN(n15412) );
  NAND2X0 U15933 ( .IN1(n15407), .IN2(n10392), .QN(n15400) );
  NAND2X0 U15934 ( .IN1(n15415), .IN2(n15416), .QN(g30354) );
  NAND2X0 U15935 ( .IN1(n10513), .IN2(g1825), .QN(n15416) );
  NOR2X0 U15936 ( .IN1(n15417), .IN2(n15418), .QN(n15415) );
  NOR2X0 U15937 ( .IN1(n5413), .IN2(n15419), .QN(n15418) );
  NOR2X0 U15938 ( .IN1(n15420), .IN2(n13857), .QN(n15419) );
  INVX0 U15939 ( .INP(n13843), .ZN(n13857) );
  NOR2X0 U15940 ( .IN1(n10484), .IN2(n10115), .QN(n15420) );
  NOR2X0 U15941 ( .IN1(n13862), .IN2(n15421), .QN(n15417) );
  NAND2X0 U15942 ( .IN1(n783), .IN2(n15422), .QN(n15421) );
  XOR2X1 U15943 ( .IN1(n9823), .IN2(n9654), .Q(n15422) );
  INVX0 U15944 ( .INP(n13844), .ZN(n783) );
  NAND2X0 U15945 ( .IN1(n15423), .IN2(n15424), .QN(g30353) );
  NAND2X0 U15946 ( .IN1(n10513), .IN2(g1748), .QN(n15424) );
  NAND2X0 U15947 ( .IN1(n15425), .IN2(n10392), .QN(n15423) );
  NAND2X0 U15948 ( .IN1(n15426), .IN2(n15427), .QN(n15425) );
  NAND2X0 U15949 ( .IN1(n15428), .IN2(g1768), .QN(n15427) );
  NAND2X0 U15950 ( .IN1(n15429), .IN2(n15430), .QN(n15426) );
  NAND2X0 U15951 ( .IN1(n5352), .IN2(g1772), .QN(n15430) );
  INVX0 U15952 ( .INP(n15428), .ZN(n15429) );
  NAND2X0 U15953 ( .IN1(n15431), .IN2(n5359), .QN(n15428) );
  NOR2X0 U15954 ( .IN1(n5596), .IN2(n13837), .QN(n15431) );
  NAND2X0 U15955 ( .IN1(n15432), .IN2(n15433), .QN(g30352) );
  OR2X1 U15956 ( .IN1(n15434), .IN2(n18480), .Q(n15433) );
  NOR2X0 U15957 ( .IN1(n15435), .IN2(n15436), .QN(n15432) );
  NOR2X0 U15958 ( .IN1(g1720), .IN2(n15437), .QN(n15436) );
  NAND2X0 U15959 ( .IN1(n15438), .IN2(n15439), .QN(n15437) );
  NOR2X0 U15960 ( .IN1(n10484), .IN2(g1714), .QN(n15438) );
  NOR2X0 U15961 ( .IN1(n5780), .IN2(n15440), .QN(n15435) );
  NOR2X0 U15962 ( .IN1(n10483), .IN2(n15441), .QN(n15440) );
  NOR2X0 U15963 ( .IN1(n5460), .IN2(n15442), .QN(n15441) );
  NAND2X0 U15964 ( .IN1(n15443), .IN2(n15444), .QN(g30351) );
  NAND2X0 U15965 ( .IN1(n15445), .IN2(g1720), .QN(n15444) );
  NAND2X0 U15966 ( .IN1(n15434), .IN2(g1714), .QN(n15443) );
  NAND2X0 U15967 ( .IN1(n15446), .IN2(n15447), .QN(g30350) );
  NAND2X0 U15968 ( .IN1(n15445), .IN2(g1700), .QN(n15447) );
  INVX0 U15969 ( .INP(n15434), .ZN(n15445) );
  NAND2X0 U15970 ( .IN1(n15442), .IN2(n10392), .QN(n15434) );
  NOR2X0 U15971 ( .IN1(n15448), .IN2(n15449), .QN(n15446) );
  NOR2X0 U15972 ( .IN1(n5628), .IN2(n10327), .QN(n15449) );
  NOR2X0 U15973 ( .IN1(n10483), .IN2(n15450), .QN(n15448) );
  NAND2X0 U15974 ( .IN1(n15439), .IN2(n5417), .QN(n15450) );
  INVX0 U15975 ( .INP(n15442), .ZN(n15439) );
  NAND2X0 U15976 ( .IN1(n15451), .IN2(n15452), .QN(g30349) );
  NAND2X0 U15977 ( .IN1(n10514), .IN2(g1691), .QN(n15452) );
  NOR2X0 U15978 ( .IN1(n15453), .IN2(n15454), .QN(n15451) );
  NOR2X0 U15979 ( .IN1(n5628), .IN2(n15455), .QN(n15454) );
  NOR2X0 U15980 ( .IN1(n15456), .IN2(n13895), .QN(n15455) );
  NOR2X0 U15981 ( .IN1(n10483), .IN2(n1019), .QN(n15456) );
  NOR2X0 U15982 ( .IN1(n13900), .IN2(n15457), .QN(n15453) );
  NAND2X0 U15983 ( .IN1(n8), .IN2(n15458), .QN(n15457) );
  XOR2X1 U15984 ( .IN1(n9827), .IN2(n9658), .Q(n15458) );
  INVX0 U15985 ( .INP(n13879), .ZN(n8) );
  NAND2X0 U15986 ( .IN1(n15459), .IN2(n15460), .QN(g30348) );
  NAND2X0 U15987 ( .IN1(n10513), .IN2(g1612), .QN(n15460) );
  NOR2X0 U15988 ( .IN1(n15461), .IN2(n15462), .QN(n15459) );
  NOR2X0 U15989 ( .IN1(n5836), .IN2(n15463), .QN(n15462) );
  NOR2X0 U15990 ( .IN1(n15464), .IN2(n13895), .QN(n15463) );
  INVX0 U15991 ( .INP(n13878), .ZN(n13895) );
  NOR2X0 U15992 ( .IN1(n10483), .IN2(g31863), .QN(n15464) );
  NOR2X0 U15993 ( .IN1(n13879), .IN2(n15465), .QN(n15461) );
  NAND2X0 U15994 ( .IN1(g31863), .IN2(n15466), .QN(n15465) );
  NAND2X0 U15995 ( .IN1(n5362), .IN2(g1636), .QN(n15466) );
  NAND2X0 U15996 ( .IN1(n15467), .IN2(n15468), .QN(g30347) );
  NAND2X0 U15997 ( .IN1(n15469), .IN2(n15470), .QN(n15468) );
  INVX0 U15998 ( .INP(n15471), .ZN(n15470) );
  NOR2X0 U15999 ( .IN1(n15472), .IN2(n15473), .QN(n15469) );
  NOR2X0 U16000 ( .IN1(n15474), .IN2(n15475), .QN(n15473) );
  NOR2X0 U16001 ( .IN1(n9572), .IN2(n10463), .QN(n15475) );
  NOR2X0 U16002 ( .IN1(n9572), .IN2(n15476), .QN(n15472) );
  OR2X1 U16003 ( .IN1(n10309), .IN2(n9775), .Q(n15467) );
  NAND2X0 U16004 ( .IN1(n15477), .IN2(n15478), .QN(g30346) );
  NAND2X0 U16005 ( .IN1(n10513), .IN2(g1536), .QN(n15478) );
  NAND2X0 U16006 ( .IN1(n15479), .IN2(n10392), .QN(n15477) );
  NOR2X0 U16007 ( .IN1(n15471), .IN2(n15480), .QN(n15479) );
  NAND2X0 U16008 ( .IN1(n15481), .IN2(n15476), .QN(n15480) );
  NAND2X0 U16009 ( .IN1(n9775), .IN2(n15482), .QN(n15481) );
  NAND2X0 U16010 ( .IN1(n15483), .IN2(n15484), .QN(g30345) );
  NAND2X0 U16011 ( .IN1(n15485), .IN2(n10392), .QN(n15484) );
  OR2X1 U16012 ( .IN1(n15471), .IN2(n12991), .Q(n15485) );
  NAND2X0 U16013 ( .IN1(n15486), .IN2(g1514), .QN(n15483) );
  NAND2X0 U16014 ( .IN1(n15487), .IN2(n10392), .QN(n15486) );
  XOR2X1 U16015 ( .IN1(test_so49), .IN2(n5302), .Q(n15487) );
  NOR2X0 U16016 ( .IN1(n10483), .IN2(n15488), .QN(g30344) );
  NOR2X0 U16017 ( .IN1(n15471), .IN2(n15489), .QN(n15488) );
  XOR2X1 U16018 ( .IN1(n5364), .IN2(n5302), .Q(n15489) );
  NAND2X0 U16019 ( .IN1(n15490), .IN2(n15491), .QN(n15471) );
  NAND2X0 U16020 ( .IN1(n4172), .IN2(n12991), .QN(n15491) );
  NOR2X0 U16021 ( .IN1(n15492), .IN2(n15493), .QN(n4172) );
  NAND2X0 U16022 ( .IN1(n9907), .IN2(n4895), .QN(n15493) );
  NAND2X0 U16023 ( .IN1(n15494), .IN2(g7946), .QN(n15492) );
  NOR2X0 U16024 ( .IN1(n5577), .IN2(n5381), .QN(n15494) );
  NAND2X0 U16025 ( .IN1(n15495), .IN2(n15496), .QN(g30343) );
  NAND2X0 U16026 ( .IN1(n4175), .IN2(n13906), .QN(n15496) );
  NOR2X0 U16027 ( .IN1(n15497), .IN2(n15498), .QN(n15495) );
  NOR2X0 U16028 ( .IN1(n10483), .IN2(n15499), .QN(n15498) );
  OR2X1 U16029 ( .IN1(n3734), .IN2(n9761), .Q(n15499) );
  AND2X1 U16030 ( .IN1(n15500), .IN2(n15501), .Q(n3734) );
  NAND2X0 U16031 ( .IN1(n9750), .IN2(n13297), .QN(n15500) );
  INVX0 U16032 ( .INP(n13302), .ZN(n13297) );
  NOR2X0 U16033 ( .IN1(n9750), .IN2(n10327), .QN(n15497) );
  NAND2X0 U16034 ( .IN1(n15502), .IN2(n15503), .QN(g30342) );
  NAND2X0 U16035 ( .IN1(n10513), .IN2(g1256), .QN(n15503) );
  NOR2X0 U16036 ( .IN1(n15504), .IN2(n15505), .QN(n15502) );
  NOR2X0 U16037 ( .IN1(g1259), .IN2(n15506), .QN(n15505) );
  NOR2X0 U16038 ( .IN1(n5553), .IN2(n15507), .QN(n15504) );
  NAND2X0 U16039 ( .IN1(n13309), .IN2(n15506), .QN(n15507) );
  INVX0 U16040 ( .INP(n3736), .ZN(n15506) );
  NAND2X0 U16041 ( .IN1(n15508), .IN2(n15509), .QN(g30341) );
  NAND2X0 U16042 ( .IN1(n15510), .IN2(n15511), .QN(n15509) );
  INVX0 U16043 ( .INP(n15512), .ZN(n15511) );
  NOR2X0 U16044 ( .IN1(n15513), .IN2(n15514), .QN(n15510) );
  NOR2X0 U16045 ( .IN1(n15515), .IN2(n15516), .QN(n15514) );
  NOR2X0 U16046 ( .IN1(n9571), .IN2(n10462), .QN(n15516) );
  NOR2X0 U16047 ( .IN1(n9571), .IN2(n15517), .QN(n15513) );
  OR2X1 U16048 ( .IN1(n10308), .IN2(n9776), .Q(n15508) );
  NAND2X0 U16049 ( .IN1(n15518), .IN2(n15519), .QN(g30340) );
  NAND2X0 U16050 ( .IN1(n10513), .IN2(g1193), .QN(n15519) );
  NAND2X0 U16051 ( .IN1(n15520), .IN2(n10392), .QN(n15518) );
  NOR2X0 U16052 ( .IN1(n15512), .IN2(n15521), .QN(n15520) );
  NAND2X0 U16053 ( .IN1(n15522), .IN2(n15517), .QN(n15521) );
  NAND2X0 U16054 ( .IN1(n9776), .IN2(n15523), .QN(n15522) );
  NAND2X0 U16055 ( .IN1(n15524), .IN2(n15525), .QN(g30339) );
  NAND2X0 U16056 ( .IN1(n15526), .IN2(n10392), .QN(n15525) );
  OR2X1 U16057 ( .IN1(n15512), .IN2(n13234), .Q(n15526) );
  NAND2X0 U16058 ( .IN1(n15527), .IN2(g1171), .QN(n15524) );
  NAND2X0 U16059 ( .IN1(n15528), .IN2(n10393), .QN(n15527) );
  XOR2X1 U16060 ( .IN1(g7916), .IN2(n5599), .Q(n15528) );
  NOR2X0 U16061 ( .IN1(n10483), .IN2(n15529), .QN(g30338) );
  NOR2X0 U16062 ( .IN1(n15512), .IN2(n15530), .QN(n15529) );
  XOR2X1 U16063 ( .IN1(n5363), .IN2(n5304), .Q(n15530) );
  NAND2X0 U16064 ( .IN1(n15531), .IN2(n15532), .QN(n15512) );
  NAND2X0 U16065 ( .IN1(n4190), .IN2(n13234), .QN(n15532) );
  NOR2X0 U16066 ( .IN1(n15533), .IN2(n15534), .QN(n4190) );
  NAND2X0 U16067 ( .IN1(n5642), .IN2(n4920), .QN(n15534) );
  NAND2X0 U16068 ( .IN1(n15535), .IN2(g7916), .QN(n15533) );
  NOR2X0 U16069 ( .IN1(n9757), .IN2(n9756), .QN(n15535) );
  NAND2X0 U16070 ( .IN1(n15536), .IN2(n15537), .QN(g30337) );
  NAND2X0 U16071 ( .IN1(n4193), .IN2(n13922), .QN(n15537) );
  NOR2X0 U16072 ( .IN1(n15538), .IN2(n15539), .QN(n15536) );
  NOR2X0 U16073 ( .IN1(n10483), .IN2(n15540), .QN(n15539) );
  NAND2X0 U16074 ( .IN1(n14094), .IN2(g1018), .QN(n15540) );
  NAND2X0 U16075 ( .IN1(n15541), .IN2(n15542), .QN(n14094) );
  NAND2X0 U16076 ( .IN1(n9751), .IN2(n13316), .QN(n15541) );
  INVX0 U16077 ( .INP(n13321), .ZN(n13316) );
  NOR2X0 U16078 ( .IN1(n9751), .IN2(n10327), .QN(n15538) );
  NAND2X0 U16079 ( .IN1(n15543), .IN2(n15544), .QN(g30336) );
  NAND2X0 U16080 ( .IN1(n10513), .IN2(g911), .QN(n15544) );
  NOR2X0 U16081 ( .IN1(n15545), .IN2(n15546), .QN(n15543) );
  NOR2X0 U16082 ( .IN1(g914), .IN2(n15547), .QN(n15546) );
  NOR2X0 U16083 ( .IN1(n5560), .IN2(n15548), .QN(n15545) );
  NAND2X0 U16084 ( .IN1(n13328), .IN2(n15547), .QN(n15548) );
  INVX0 U16085 ( .INP(n3741), .ZN(n15547) );
  NAND2X0 U16086 ( .IN1(n15549), .IN2(n15550), .QN(g30335) );
  NAND2X0 U16087 ( .IN1(test_so60), .IN2(n10514), .QN(n15550) );
  NOR2X0 U16088 ( .IN1(n15551), .IN2(n15552), .QN(n15549) );
  NOR2X0 U16089 ( .IN1(g744), .IN2(n10770), .QN(n15552) );
  NOR2X0 U16090 ( .IN1(n5470), .IN2(n15553), .QN(n15551) );
  NAND2X0 U16091 ( .IN1(n2404), .IN2(n10770), .QN(n15553) );
  NAND2X0 U16092 ( .IN1(n15554), .IN2(test_so60), .QN(n10770) );
  NOR2X0 U16093 ( .IN1(n10758), .IN2(n15555), .QN(n15554) );
  NOR2X0 U16094 ( .IN1(g736), .IN2(n5482), .QN(n10758) );
  NAND2X0 U16095 ( .IN1(n15556), .IN2(n15557), .QN(g30334) );
  NAND2X0 U16096 ( .IN1(n10513), .IN2(g586), .QN(n15557) );
  NOR2X0 U16097 ( .IN1(n15558), .IN2(n15559), .QN(n15556) );
  NOR2X0 U16098 ( .IN1(g577), .IN2(n15560), .QN(n15559) );
  NOR2X0 U16099 ( .IN1(n5294), .IN2(n15561), .QN(n15558) );
  NAND2X0 U16100 ( .IN1(n2421), .IN2(n15560), .QN(n15561) );
  INVX0 U16101 ( .INP(n3745), .ZN(n15560) );
  NAND2X0 U16102 ( .IN1(n15562), .IN2(n15563), .QN(g30333) );
  NAND2X0 U16103 ( .IN1(n11894), .IN2(n15564), .QN(n15563) );
  XOR2X1 U16104 ( .IN1(test_so73), .IN2(n15565), .Q(n15564) );
  NOR2X0 U16105 ( .IN1(n14125), .IN2(n10462), .QN(n11894) );
  NAND2X0 U16106 ( .IN1(n15566), .IN2(n15567), .QN(n14125) );
  NAND2X0 U16107 ( .IN1(n15565), .IN2(n15568), .QN(n15567) );
  NAND2X0 U16108 ( .IN1(n15569), .IN2(n10136), .QN(n15568) );
  INVX0 U16109 ( .INP(n14124), .ZN(n15565) );
  NAND2X0 U16110 ( .IN1(n10512), .IN2(g142), .QN(n15562) );
  NAND2X0 U16111 ( .IN1(n15570), .IN2(n15571), .QN(g29309) );
  NAND2X0 U16112 ( .IN1(n3765), .IN2(n15572), .QN(n15571) );
  NAND2X0 U16113 ( .IN1(g6541), .IN2(n12631), .QN(n15572) );
  NOR2X0 U16114 ( .IN1(n15573), .IN2(n15574), .QN(n15570) );
  NOR2X0 U16115 ( .IN1(n14161), .IN2(n15575), .QN(n15574) );
  NAND2X0 U16116 ( .IN1(n15576), .IN2(g6541), .QN(n15575) );
  NAND2X0 U16117 ( .IN1(n15577), .IN2(n15578), .QN(g29308) );
  NAND2X0 U16118 ( .IN1(n10512), .IN2(g6523), .QN(n15578) );
  NOR2X0 U16119 ( .IN1(n15579), .IN2(n15580), .QN(n15577) );
  AND2X1 U16120 ( .IN1(n15581), .IN2(n5659), .Q(n15580) );
  NOR2X0 U16121 ( .IN1(n5659), .IN2(n15582), .QN(n15579) );
  NAND2X0 U16122 ( .IN1(n15583), .IN2(n15584), .QN(g29307) );
  NAND2X0 U16123 ( .IN1(n15585), .IN2(g6523), .QN(n15584) );
  NOR2X0 U16124 ( .IN1(n15586), .IN2(n15587), .QN(n15583) );
  NOR2X0 U16125 ( .IN1(g6519), .IN2(n15588), .QN(n15587) );
  NAND2X0 U16126 ( .IN1(n5426), .IN2(n15581), .QN(n15588) );
  NOR2X0 U16127 ( .IN1(n5806), .IN2(n15589), .QN(n15586) );
  NOR2X0 U16128 ( .IN1(n10483), .IN2(n15590), .QN(n15589) );
  NOR2X0 U16129 ( .IN1(n5426), .IN2(n15591), .QN(n15590) );
  NAND2X0 U16130 ( .IN1(n15592), .IN2(n15593), .QN(g29306) );
  NAND2X0 U16131 ( .IN1(n15585), .IN2(g6519), .QN(n15593) );
  INVX0 U16132 ( .INP(n15582), .ZN(n15585) );
  NAND2X0 U16133 ( .IN1(n15582), .IN2(g6513), .QN(n15592) );
  NAND2X0 U16134 ( .IN1(n15591), .IN2(n10393), .QN(n15582) );
  NAND2X0 U16135 ( .IN1(n15594), .IN2(n15595), .QN(g29305) );
  NAND2X0 U16136 ( .IN1(n14130), .IN2(n15591), .QN(n15595) );
  INVX0 U16137 ( .INP(n11291), .ZN(n14130) );
  NAND2X0 U16138 ( .IN1(n10367), .IN2(g6509), .QN(n11291) );
  NOR2X0 U16139 ( .IN1(n15596), .IN2(n15597), .QN(n15594) );
  NOR2X0 U16140 ( .IN1(g6500), .IN2(n15598), .QN(n15597) );
  NAND2X0 U16141 ( .IN1(n15581), .IN2(g6505), .QN(n15598) );
  NOR2X0 U16142 ( .IN1(n15591), .IN2(n10461), .QN(n15581) );
  NOR2X0 U16143 ( .IN1(n5748), .IN2(n15599), .QN(n15596) );
  NOR2X0 U16144 ( .IN1(n10483), .IN2(n15600), .QN(n15599) );
  NOR2X0 U16145 ( .IN1(n15591), .IN2(g6505), .QN(n15600) );
  NAND2X0 U16146 ( .IN1(n15601), .IN2(n12655), .QN(n15591) );
  NAND2X0 U16147 ( .IN1(n15602), .IN2(n15603), .QN(g29304) );
  NAND2X0 U16148 ( .IN1(n10512), .IN2(g6505), .QN(n15603) );
  NAND2X0 U16149 ( .IN1(n15604), .IN2(n10393), .QN(n15602) );
  NAND2X0 U16150 ( .IN1(n15605), .IN2(n15606), .QN(n15604) );
  NAND2X0 U16151 ( .IN1(n10113), .IN2(g6500), .QN(n15606) );
  INVX0 U16152 ( .INP(n12655), .ZN(n10113) );
  NAND2X0 U16153 ( .IN1(n15607), .IN2(n12655), .QN(n15605) );
  XOR2X1 U16154 ( .IN1(n15608), .IN2(n15609), .Q(n15607) );
  NOR2X0 U16155 ( .IN1(n15601), .IN2(n5748), .QN(n15609) );
  AND2X1 U16156 ( .IN1(n15610), .IN2(n15611), .Q(n15601) );
  NOR2X0 U16157 ( .IN1(n9995), .IN2(n5531), .QN(n15610) );
  NAND2X0 U16158 ( .IN1(n15612), .IN2(n15613), .QN(g29303) );
  NAND2X0 U16159 ( .IN1(n3765), .IN2(n15614), .QN(n15613) );
  NAND2X0 U16160 ( .IN1(g6195), .IN2(n12624), .QN(n15614) );
  NOR2X0 U16161 ( .IN1(n15573), .IN2(n15615), .QN(n15612) );
  NOR2X0 U16162 ( .IN1(n14281), .IN2(n15616), .QN(n15615) );
  NAND2X0 U16163 ( .IN1(n15576), .IN2(g6195), .QN(n15616) );
  NAND2X0 U16164 ( .IN1(n15617), .IN2(n15618), .QN(g29302) );
  NAND2X0 U16165 ( .IN1(n10512), .IN2(g6177), .QN(n15618) );
  NOR2X0 U16166 ( .IN1(n15619), .IN2(n15620), .QN(n15617) );
  AND2X1 U16167 ( .IN1(n15621), .IN2(n5667), .Q(n15620) );
  NOR2X0 U16168 ( .IN1(n5667), .IN2(n15622), .QN(n15619) );
  NAND2X0 U16169 ( .IN1(n15623), .IN2(n15624), .QN(g29301) );
  NAND2X0 U16170 ( .IN1(n15625), .IN2(g6177), .QN(n15624) );
  NOR2X0 U16171 ( .IN1(n15626), .IN2(n15627), .QN(n15623) );
  NOR2X0 U16172 ( .IN1(g6173), .IN2(n15628), .QN(n15627) );
  NAND2X0 U16173 ( .IN1(n5430), .IN2(n15621), .QN(n15628) );
  NOR2X0 U16174 ( .IN1(n5810), .IN2(n15629), .QN(n15626) );
  NOR2X0 U16175 ( .IN1(n10483), .IN2(n15630), .QN(n15629) );
  NOR2X0 U16176 ( .IN1(n5430), .IN2(n15631), .QN(n15630) );
  NAND2X0 U16177 ( .IN1(n15632), .IN2(n15633), .QN(g29300) );
  NAND2X0 U16178 ( .IN1(n15625), .IN2(g6173), .QN(n15633) );
  INVX0 U16179 ( .INP(n15622), .ZN(n15625) );
  NAND2X0 U16180 ( .IN1(n15622), .IN2(g6167), .QN(n15632) );
  NAND2X0 U16181 ( .IN1(n15634), .IN2(n15635), .QN(g29299) );
  OR2X1 U16182 ( .IN1(n15622), .IN2(n9645), .Q(n15635) );
  NAND2X0 U16183 ( .IN1(n15631), .IN2(n10393), .QN(n15622) );
  NOR2X0 U16184 ( .IN1(n15636), .IN2(n15637), .QN(n15634) );
  NOR2X0 U16185 ( .IN1(g6154), .IN2(n15638), .QN(n15637) );
  NAND2X0 U16186 ( .IN1(n15621), .IN2(g6159), .QN(n15638) );
  NOR2X0 U16187 ( .IN1(n15631), .IN2(n10461), .QN(n15621) );
  NOR2X0 U16188 ( .IN1(n5747), .IN2(n15639), .QN(n15636) );
  NOR2X0 U16189 ( .IN1(n10483), .IN2(n15640), .QN(n15639) );
  NOR2X0 U16190 ( .IN1(n15631), .IN2(g6159), .QN(n15640) );
  OR2X1 U16191 ( .IN1(n15641), .IN2(n12673), .Q(n15631) );
  NAND2X0 U16192 ( .IN1(n15642), .IN2(n15643), .QN(g29298) );
  NAND2X0 U16193 ( .IN1(n10512), .IN2(g6159), .QN(n15643) );
  NAND2X0 U16194 ( .IN1(n15644), .IN2(n10393), .QN(n15642) );
  NAND2X0 U16195 ( .IN1(n15645), .IN2(n15646), .QN(n15644) );
  NAND2X0 U16196 ( .IN1(n12673), .IN2(g6154), .QN(n15646) );
  NAND2X0 U16197 ( .IN1(n15647), .IN2(n12675), .QN(n15645) );
  XNOR2X1 U16198 ( .IN1(n15648), .IN2(n15649), .Q(n15647) );
  NAND2X0 U16199 ( .IN1(g6154), .IN2(n15641), .QN(n15648) );
  NAND2X0 U16200 ( .IN1(n15650), .IN2(test_so69), .QN(n15641) );
  NOR2X0 U16201 ( .IN1(n10005), .IN2(n11715), .QN(n15650) );
  NAND2X0 U16202 ( .IN1(n15651), .IN2(n15652), .QN(g29297) );
  NAND2X0 U16203 ( .IN1(n3765), .IN2(n15653), .QN(n15652) );
  NAND2X0 U16204 ( .IN1(g5849), .IN2(n12623), .QN(n15653) );
  NOR2X0 U16205 ( .IN1(n15573), .IN2(n15654), .QN(n15651) );
  NOR2X0 U16206 ( .IN1(n15655), .IN2(n15656), .QN(n15654) );
  NAND2X0 U16207 ( .IN1(n15576), .IN2(g5849), .QN(n15656) );
  NAND2X0 U16208 ( .IN1(n15657), .IN2(n15658), .QN(g29296) );
  NAND2X0 U16209 ( .IN1(n10512), .IN2(g5831), .QN(n15658) );
  NOR2X0 U16210 ( .IN1(n15659), .IN2(n15660), .QN(n15657) );
  AND2X1 U16211 ( .IN1(n15661), .IN2(n5663), .Q(n15660) );
  NOR2X0 U16212 ( .IN1(n5663), .IN2(n15662), .QN(n15659) );
  NAND2X0 U16213 ( .IN1(n15663), .IN2(n15664), .QN(g29295) );
  NAND2X0 U16214 ( .IN1(n15665), .IN2(g5831), .QN(n15664) );
  NOR2X0 U16215 ( .IN1(n15666), .IN2(n15667), .QN(n15663) );
  NOR2X0 U16216 ( .IN1(g5827), .IN2(n15668), .QN(n15667) );
  NAND2X0 U16217 ( .IN1(n5429), .IN2(n15661), .QN(n15668) );
  NOR2X0 U16218 ( .IN1(n5809), .IN2(n15669), .QN(n15666) );
  NOR2X0 U16219 ( .IN1(n10483), .IN2(n15670), .QN(n15669) );
  NOR2X0 U16220 ( .IN1(n5429), .IN2(n15671), .QN(n15670) );
  NAND2X0 U16221 ( .IN1(n15672), .IN2(n15673), .QN(g29294) );
  NAND2X0 U16222 ( .IN1(n15665), .IN2(g5827), .QN(n15673) );
  NAND2X0 U16223 ( .IN1(n15662), .IN2(g5821), .QN(n15672) );
  NAND2X0 U16224 ( .IN1(n15674), .IN2(n15675), .QN(g29293) );
  NAND2X0 U16225 ( .IN1(n15665), .IN2(g5817), .QN(n15675) );
  INVX0 U16226 ( .INP(n15662), .ZN(n15665) );
  NAND2X0 U16227 ( .IN1(n15671), .IN2(n10393), .QN(n15662) );
  NOR2X0 U16228 ( .IN1(n15676), .IN2(n15677), .QN(n15674) );
  NOR2X0 U16229 ( .IN1(g5808), .IN2(n15678), .QN(n15677) );
  NAND2X0 U16230 ( .IN1(n15661), .IN2(g5813), .QN(n15678) );
  NOR2X0 U16231 ( .IN1(n15671), .IN2(n10461), .QN(n15661) );
  NOR2X0 U16232 ( .IN1(n5749), .IN2(n15679), .QN(n15676) );
  NOR2X0 U16233 ( .IN1(n10483), .IN2(n15680), .QN(n15679) );
  NOR2X0 U16234 ( .IN1(n15671), .IN2(g5813), .QN(n15680) );
  NAND2X0 U16235 ( .IN1(n15681), .IN2(n12695), .QN(n15671) );
  NAND2X0 U16236 ( .IN1(n15682), .IN2(n15683), .QN(g29292) );
  NAND2X0 U16237 ( .IN1(n10512), .IN2(g5813), .QN(n15683) );
  NOR2X0 U16238 ( .IN1(n15684), .IN2(n15685), .QN(n15682) );
  NOR2X0 U16239 ( .IN1(n5749), .IN2(n12700), .QN(n15685) );
  NOR2X0 U16240 ( .IN1(n12705), .IN2(n15686), .QN(n15684) );
  XOR2X1 U16241 ( .IN1(n15687), .IN2(n15688), .Q(n15686) );
  NOR2X0 U16242 ( .IN1(n15681), .IN2(n5749), .QN(n15688) );
  AND2X1 U16243 ( .IN1(n15689), .IN2(n15690), .Q(n15681) );
  NOR2X0 U16244 ( .IN1(n9981), .IN2(n5528), .QN(n15689) );
  NAND2X0 U16245 ( .IN1(n15691), .IN2(n15692), .QN(g29291) );
  NAND2X0 U16246 ( .IN1(n3765), .IN2(n15693), .QN(n15692) );
  NAND2X0 U16247 ( .IN1(g5503), .IN2(n14523), .QN(n15693) );
  NOR2X0 U16248 ( .IN1(n15573), .IN2(n15694), .QN(n15691) );
  NOR2X0 U16249 ( .IN1(n14524), .IN2(n15695), .QN(n15694) );
  NAND2X0 U16250 ( .IN1(n15576), .IN2(g5503), .QN(n15695) );
  NAND2X0 U16251 ( .IN1(n15696), .IN2(n15697), .QN(g29290) );
  NAND2X0 U16252 ( .IN1(n10512), .IN2(g5485), .QN(n15697) );
  NOR2X0 U16253 ( .IN1(n15698), .IN2(n15699), .QN(n15696) );
  AND2X1 U16254 ( .IN1(n15700), .IN2(n5660), .Q(n15699) );
  NOR2X0 U16255 ( .IN1(n5660), .IN2(n15701), .QN(n15698) );
  NAND2X0 U16256 ( .IN1(n15702), .IN2(n15703), .QN(g29289) );
  NAND2X0 U16257 ( .IN1(n15704), .IN2(g5485), .QN(n15703) );
  NOR2X0 U16258 ( .IN1(n15705), .IN2(n15706), .QN(n15702) );
  NOR2X0 U16259 ( .IN1(g5481), .IN2(n15707), .QN(n15706) );
  NAND2X0 U16260 ( .IN1(n5425), .IN2(n15700), .QN(n15707) );
  NOR2X0 U16261 ( .IN1(n5805), .IN2(n15708), .QN(n15705) );
  NOR2X0 U16262 ( .IN1(n10482), .IN2(n15709), .QN(n15708) );
  NOR2X0 U16263 ( .IN1(n5425), .IN2(n15710), .QN(n15709) );
  NAND2X0 U16264 ( .IN1(n15711), .IN2(n15712), .QN(g29288) );
  NAND2X0 U16265 ( .IN1(n15704), .IN2(g5481), .QN(n15712) );
  NAND2X0 U16266 ( .IN1(n15701), .IN2(g5475), .QN(n15711) );
  NAND2X0 U16267 ( .IN1(n15713), .IN2(n15714), .QN(g29287) );
  NAND2X0 U16268 ( .IN1(n15704), .IN2(g5471), .QN(n15714) );
  INVX0 U16269 ( .INP(n15701), .ZN(n15704) );
  NAND2X0 U16270 ( .IN1(n15710), .IN2(n10393), .QN(n15701) );
  NOR2X0 U16271 ( .IN1(n15715), .IN2(n15716), .QN(n15713) );
  NOR2X0 U16272 ( .IN1(g5462), .IN2(n15717), .QN(n15716) );
  NAND2X0 U16273 ( .IN1(n15700), .IN2(g5467), .QN(n15717) );
  NOR2X0 U16274 ( .IN1(n15710), .IN2(n10461), .QN(n15700) );
  NOR2X0 U16275 ( .IN1(n5744), .IN2(n15718), .QN(n15715) );
  NOR2X0 U16276 ( .IN1(n10482), .IN2(n15719), .QN(n15718) );
  NOR2X0 U16277 ( .IN1(n15710), .IN2(g5467), .QN(n15719) );
  NAND2X0 U16278 ( .IN1(n15720), .IN2(n12717), .QN(n15710) );
  NAND2X0 U16279 ( .IN1(n15721), .IN2(n15722), .QN(g29286) );
  NAND2X0 U16280 ( .IN1(n10512), .IN2(g5467), .QN(n15722) );
  NAND2X0 U16281 ( .IN1(n15723), .IN2(n10393), .QN(n15721) );
  NAND2X0 U16282 ( .IN1(n15724), .IN2(n15725), .QN(n15723) );
  NAND2X0 U16283 ( .IN1(n12715), .IN2(g5462), .QN(n15725) );
  NAND2X0 U16284 ( .IN1(n15726), .IN2(n12717), .QN(n15724) );
  XOR2X1 U16285 ( .IN1(n15727), .IN2(n15728), .Q(n15726) );
  NOR2X0 U16286 ( .IN1(n15720), .IN2(n5744), .QN(n15728) );
  AND2X1 U16287 ( .IN1(n15729), .IN2(n15730), .Q(n15720) );
  NOR2X0 U16288 ( .IN1(n9986), .IN2(n5529), .QN(n15729) );
  NAND2X0 U16289 ( .IN1(n15731), .IN2(n15732), .QN(g29285) );
  NAND2X0 U16290 ( .IN1(n3765), .IN2(n15733), .QN(n15732) );
  NAND2X0 U16291 ( .IN1(g5156), .IN2(n12619), .QN(n15733) );
  NOR2X0 U16292 ( .IN1(n15573), .IN2(n15734), .QN(n15731) );
  NOR2X0 U16293 ( .IN1(n14645), .IN2(n15735), .QN(n15734) );
  NAND2X0 U16294 ( .IN1(n15576), .IN2(g5156), .QN(n15735) );
  NAND2X0 U16295 ( .IN1(n15736), .IN2(n15737), .QN(g29284) );
  NAND2X0 U16296 ( .IN1(n10512), .IN2(g5138), .QN(n15737) );
  NOR2X0 U16297 ( .IN1(n15738), .IN2(n15739), .QN(n15736) );
  AND2X1 U16298 ( .IN1(n15740), .IN2(n5658), .Q(n15739) );
  NOR2X0 U16299 ( .IN1(n5658), .IN2(n15741), .QN(n15738) );
  NAND2X0 U16300 ( .IN1(n15742), .IN2(n15743), .QN(g29283) );
  NAND2X0 U16301 ( .IN1(n15744), .IN2(g5138), .QN(n15743) );
  NOR2X0 U16302 ( .IN1(n15745), .IN2(n15746), .QN(n15742) );
  NOR2X0 U16303 ( .IN1(g5134), .IN2(n15747), .QN(n15746) );
  NAND2X0 U16304 ( .IN1(n15740), .IN2(n10141), .QN(n15747) );
  NOR2X0 U16305 ( .IN1(n5807), .IN2(n15748), .QN(n15745) );
  NOR2X0 U16306 ( .IN1(n10482), .IN2(n15749), .QN(n15748) );
  NOR2X0 U16307 ( .IN1(n15750), .IN2(n10141), .QN(n15749) );
  NAND2X0 U16308 ( .IN1(n15751), .IN2(n15752), .QN(g29282) );
  NAND2X0 U16309 ( .IN1(n15744), .IN2(g5134), .QN(n15752) );
  INVX0 U16310 ( .INP(n15741), .ZN(n15744) );
  NAND2X0 U16311 ( .IN1(test_so96), .IN2(n15741), .QN(n15751) );
  NAND2X0 U16312 ( .IN1(n15750), .IN2(n10393), .QN(n15741) );
  NAND2X0 U16313 ( .IN1(n15753), .IN2(n15754), .QN(g29281) );
  NAND2X0 U16314 ( .IN1(n14140), .IN2(n15750), .QN(n15754) );
  NOR2X0 U16315 ( .IN1(n10482), .IN2(n9616), .QN(n14140) );
  NOR2X0 U16316 ( .IN1(n15755), .IN2(n15756), .QN(n15753) );
  NOR2X0 U16317 ( .IN1(g5115), .IN2(n15757), .QN(n15756) );
  NAND2X0 U16318 ( .IN1(n15740), .IN2(g5120), .QN(n15757) );
  NOR2X0 U16319 ( .IN1(n15750), .IN2(n10461), .QN(n15740) );
  NOR2X0 U16320 ( .IN1(n5743), .IN2(n15758), .QN(n15755) );
  NOR2X0 U16321 ( .IN1(n10482), .IN2(n15759), .QN(n15758) );
  NOR2X0 U16322 ( .IN1(n15750), .IN2(g5120), .QN(n15759) );
  NAND2X0 U16323 ( .IN1(n15760), .IN2(g33959), .QN(n15750) );
  NAND2X0 U16324 ( .IN1(n15761), .IN2(n15762), .QN(g29280) );
  NAND2X0 U16325 ( .IN1(n10512), .IN2(g5120), .QN(n15762) );
  NAND2X0 U16326 ( .IN1(n15763), .IN2(n10393), .QN(n15761) );
  NAND2X0 U16327 ( .IN1(n15764), .IN2(n15765), .QN(n15763) );
  NAND2X0 U16328 ( .IN1(n10108), .IN2(g5115), .QN(n15765) );
  NAND2X0 U16329 ( .IN1(n15766), .IN2(g33959), .QN(n15764) );
  XOR2X1 U16330 ( .IN1(n15767), .IN2(n15768), .Q(n15766) );
  NOR2X0 U16331 ( .IN1(n15760), .IN2(n5743), .QN(n15768) );
  AND2X1 U16332 ( .IN1(n15769), .IN2(test_so10), .Q(n15760) );
  NOR2X0 U16333 ( .IN1(n9976), .IN2(n10666), .QN(n15769) );
  OR2X1 U16334 ( .IN1(n15770), .IN2(g29279), .Q(g29278) );
  NOR2X0 U16335 ( .IN1(n9677), .IN2(n10327), .QN(n15770) );
  OR2X1 U16336 ( .IN1(n15771), .IN2(g29277), .Q(g29276) );
  NOR2X0 U16337 ( .IN1(n10357), .IN2(n10150), .QN(n15771) );
  NAND2X0 U16338 ( .IN1(n15772), .IN2(n15773), .QN(g29275) );
  NAND2X0 U16339 ( .IN1(n15774), .IN2(n14778), .QN(n15773) );
  XOR2X1 U16340 ( .IN1(n14071), .IN2(n5480), .Q(n15774) );
  NAND2X0 U16341 ( .IN1(test_so11), .IN2(n15775), .QN(n14071) );
  NAND2X0 U16342 ( .IN1(test_so11), .IN2(n10514), .QN(n15772) );
  NAND2X0 U16343 ( .IN1(n15776), .IN2(n15777), .QN(g29274) );
  NAND2X0 U16344 ( .IN1(n3765), .IN2(n15778), .QN(n15777) );
  NAND2X0 U16345 ( .IN1(g3849), .IN2(n12636), .QN(n15778) );
  NOR2X0 U16346 ( .IN1(n15573), .IN2(n15779), .QN(n15776) );
  NOR2X0 U16347 ( .IN1(n14785), .IN2(n15780), .QN(n15779) );
  NAND2X0 U16348 ( .IN1(n15576), .IN2(g3849), .QN(n15780) );
  NAND2X0 U16349 ( .IN1(n15781), .IN2(n15782), .QN(g29273) );
  NAND2X0 U16350 ( .IN1(n10512), .IN2(g3831), .QN(n15782) );
  NOR2X0 U16351 ( .IN1(n15783), .IN2(n15784), .QN(n15781) );
  AND2X1 U16352 ( .IN1(n15785), .IN2(n5662), .Q(n15784) );
  NOR2X0 U16353 ( .IN1(n5662), .IN2(n15786), .QN(n15783) );
  NAND2X0 U16354 ( .IN1(n15787), .IN2(n15788), .QN(g29272) );
  NAND2X0 U16355 ( .IN1(n15789), .IN2(g3831), .QN(n15788) );
  NOR2X0 U16356 ( .IN1(n15790), .IN2(n15791), .QN(n15787) );
  NOR2X0 U16357 ( .IN1(g3827), .IN2(n15792), .QN(n15791) );
  NAND2X0 U16358 ( .IN1(n5428), .IN2(n15785), .QN(n15792) );
  NOR2X0 U16359 ( .IN1(n5808), .IN2(n15793), .QN(n15790) );
  NOR2X0 U16360 ( .IN1(n10482), .IN2(n15794), .QN(n15793) );
  NOR2X0 U16361 ( .IN1(n5428), .IN2(n15795), .QN(n15794) );
  NAND2X0 U16362 ( .IN1(n15796), .IN2(n15797), .QN(g29271) );
  NAND2X0 U16363 ( .IN1(n15789), .IN2(g3827), .QN(n15797) );
  INVX0 U16364 ( .INP(n15786), .ZN(n15789) );
  NAND2X0 U16365 ( .IN1(n15786), .IN2(g3821), .QN(n15796) );
  NAND2X0 U16366 ( .IN1(n15795), .IN2(n10394), .QN(n15786) );
  NAND2X0 U16367 ( .IN1(n15798), .IN2(n15799), .QN(g29270) );
  NAND2X0 U16368 ( .IN1(n14153), .IN2(n15795), .QN(n15799) );
  NOR2X0 U16369 ( .IN1(n10482), .IN2(n9617), .QN(n14153) );
  NOR2X0 U16370 ( .IN1(n15800), .IN2(n15801), .QN(n15798) );
  NOR2X0 U16371 ( .IN1(g3808), .IN2(n15802), .QN(n15801) );
  NAND2X0 U16372 ( .IN1(n15785), .IN2(g3813), .QN(n15802) );
  NOR2X0 U16373 ( .IN1(n15795), .IN2(n10460), .QN(n15785) );
  NOR2X0 U16374 ( .IN1(n5745), .IN2(n15803), .QN(n15800) );
  NOR2X0 U16375 ( .IN1(n10482), .IN2(n15804), .QN(n15803) );
  NOR2X0 U16376 ( .IN1(n15795), .IN2(g3813), .QN(n15804) );
  OR2X1 U16377 ( .IN1(n15805), .IN2(n12766), .Q(n15795) );
  NAND2X0 U16378 ( .IN1(n15806), .IN2(n15807), .QN(g29269) );
  NAND2X0 U16379 ( .IN1(n10512), .IN2(g3813), .QN(n15807) );
  NAND2X0 U16380 ( .IN1(n15808), .IN2(n10394), .QN(n15806) );
  NAND2X0 U16381 ( .IN1(n15809), .IN2(n15810), .QN(n15808) );
  NAND2X0 U16382 ( .IN1(n12766), .IN2(g3808), .QN(n15810) );
  NAND2X0 U16383 ( .IN1(n15811), .IN2(n12768), .QN(n15809) );
  XNOR2X1 U16384 ( .IN1(n15812), .IN2(n15813), .Q(n15811) );
  NAND2X0 U16385 ( .IN1(g3808), .IN2(n15805), .QN(n15812) );
  NAND2X0 U16386 ( .IN1(n15814), .IN2(n15815), .QN(n15805) );
  NOR2X0 U16387 ( .IN1(n9990), .IN2(n5530), .QN(n15814) );
  NAND2X0 U16388 ( .IN1(n15816), .IN2(n15817), .QN(g29268) );
  NAND2X0 U16389 ( .IN1(n3765), .IN2(n15818), .QN(n15817) );
  NAND2X0 U16390 ( .IN1(g3498), .IN2(n12635), .QN(n15818) );
  NOR2X0 U16391 ( .IN1(n15573), .IN2(n15819), .QN(n15816) );
  NOR2X0 U16392 ( .IN1(n14906), .IN2(n15820), .QN(n15819) );
  NAND2X0 U16393 ( .IN1(n15576), .IN2(g3498), .QN(n15820) );
  NAND2X0 U16394 ( .IN1(n15821), .IN2(n15822), .QN(g29267) );
  NAND2X0 U16395 ( .IN1(n10512), .IN2(g3480), .QN(n15822) );
  NOR2X0 U16396 ( .IN1(n15823), .IN2(n15824), .QN(n15821) );
  AND2X1 U16397 ( .IN1(n15825), .IN2(n5668), .Q(n15824) );
  NOR2X0 U16398 ( .IN1(n5668), .IN2(n15826), .QN(n15823) );
  NAND2X0 U16399 ( .IN1(n15827), .IN2(n15828), .QN(g29266) );
  NAND2X0 U16400 ( .IN1(n15829), .IN2(g3480), .QN(n15828) );
  NOR2X0 U16401 ( .IN1(n15830), .IN2(n15831), .QN(n15827) );
  NOR2X0 U16402 ( .IN1(g3476), .IN2(n15832), .QN(n15831) );
  NAND2X0 U16403 ( .IN1(n5424), .IN2(n15825), .QN(n15832) );
  NOR2X0 U16404 ( .IN1(n5786), .IN2(n15833), .QN(n15830) );
  NOR2X0 U16405 ( .IN1(n10482), .IN2(n15834), .QN(n15833) );
  NOR2X0 U16406 ( .IN1(n5424), .IN2(n15835), .QN(n15834) );
  NAND2X0 U16407 ( .IN1(n15836), .IN2(n15837), .QN(g29265) );
  NAND2X0 U16408 ( .IN1(n15829), .IN2(g3476), .QN(n15837) );
  NAND2X0 U16409 ( .IN1(n15826), .IN2(g3470), .QN(n15836) );
  NAND2X0 U16410 ( .IN1(n15838), .IN2(n15839), .QN(g29264) );
  NAND2X0 U16411 ( .IN1(n15829), .IN2(g3466), .QN(n15839) );
  INVX0 U16412 ( .INP(n15826), .ZN(n15829) );
  NAND2X0 U16413 ( .IN1(n15835), .IN2(n10394), .QN(n15826) );
  NOR2X0 U16414 ( .IN1(n15840), .IN2(n15841), .QN(n15838) );
  NOR2X0 U16415 ( .IN1(test_so4), .IN2(n15842), .QN(n15841) );
  NAND2X0 U16416 ( .IN1(n15825), .IN2(g3462), .QN(n15842) );
  NOR2X0 U16417 ( .IN1(n15835), .IN2(n10460), .QN(n15825) );
  NOR2X0 U16418 ( .IN1(n15843), .IN2(n10144), .QN(n15840) );
  NOR2X0 U16419 ( .IN1(n10482), .IN2(n15844), .QN(n15843) );
  NOR2X0 U16420 ( .IN1(n15835), .IN2(g3462), .QN(n15844) );
  NAND2X0 U16421 ( .IN1(n15845), .IN2(n12788), .QN(n15835) );
  NAND2X0 U16422 ( .IN1(n15846), .IN2(n15847), .QN(g29263) );
  NAND2X0 U16423 ( .IN1(n10512), .IN2(g3462), .QN(n15847) );
  NAND2X0 U16424 ( .IN1(n15848), .IN2(n10394), .QN(n15846) );
  NAND2X0 U16425 ( .IN1(n15849), .IN2(n15850), .QN(n15848) );
  NAND2X0 U16426 ( .IN1(test_so4), .IN2(n12786), .QN(n15850) );
  NAND2X0 U16427 ( .IN1(n15851), .IN2(n12788), .QN(n15849) );
  XOR2X1 U16428 ( .IN1(n15852), .IN2(n15853), .Q(n15851) );
  NOR2X0 U16429 ( .IN1(n15845), .IN2(n10144), .QN(n15853) );
  AND2X1 U16430 ( .IN1(n15854), .IN2(n15855), .Q(n15845) );
  NOR2X0 U16431 ( .IN1(n5532), .IN2(n10000), .QN(n15854) );
  NAND2X0 U16432 ( .IN1(n15856), .IN2(n15857), .QN(g29262) );
  NAND2X0 U16433 ( .IN1(n3765), .IN2(n15858), .QN(n15857) );
  NAND2X0 U16434 ( .IN1(g3147), .IN2(n15026), .QN(n15858) );
  NOR2X0 U16435 ( .IN1(n15573), .IN2(n15859), .QN(n15856) );
  NOR2X0 U16436 ( .IN1(n15027), .IN2(n15860), .QN(n15859) );
  NAND2X0 U16437 ( .IN1(n15576), .IN2(g3147), .QN(n15860) );
  INVX0 U16438 ( .INP(n4210), .ZN(n15576) );
  NOR2X0 U16439 ( .IN1(n14160), .IN2(n4210), .QN(n15573) );
  NAND2X0 U16440 ( .IN1(n9725), .IN2(g4180), .QN(n4210) );
  INVX0 U16441 ( .INP(n3765), .ZN(n14160) );
  NAND2X0 U16442 ( .IN1(n15861), .IN2(n15862), .QN(g29261) );
  NAND2X0 U16443 ( .IN1(n10512), .IN2(g3129), .QN(n15862) );
  NOR2X0 U16444 ( .IN1(n15863), .IN2(n15864), .QN(n15861) );
  AND2X1 U16445 ( .IN1(n15865), .IN2(n5661), .Q(n15864) );
  NOR2X0 U16446 ( .IN1(n5661), .IN2(n15866), .QN(n15863) );
  NAND2X0 U16447 ( .IN1(n15867), .IN2(n15868), .QN(g29260) );
  NAND2X0 U16448 ( .IN1(n15869), .IN2(g3129), .QN(n15868) );
  NOR2X0 U16449 ( .IN1(n15870), .IN2(n15871), .QN(n15867) );
  NOR2X0 U16450 ( .IN1(g3125), .IN2(n15872), .QN(n15871) );
  NAND2X0 U16451 ( .IN1(n5423), .IN2(n15865), .QN(n15872) );
  NOR2X0 U16452 ( .IN1(n5781), .IN2(n15873), .QN(n15870) );
  NOR2X0 U16453 ( .IN1(n10482), .IN2(n15874), .QN(n15873) );
  NOR2X0 U16454 ( .IN1(n5423), .IN2(n15875), .QN(n15874) );
  NAND2X0 U16455 ( .IN1(n15876), .IN2(n15877), .QN(g29259) );
  NAND2X0 U16456 ( .IN1(n15869), .IN2(g3125), .QN(n15877) );
  INVX0 U16457 ( .INP(n15866), .ZN(n15869) );
  NAND2X0 U16458 ( .IN1(n15866), .IN2(g3119), .QN(n15876) );
  NAND2X0 U16459 ( .IN1(n15875), .IN2(n10394), .QN(n15866) );
  NAND2X0 U16460 ( .IN1(n15878), .IN2(n15879), .QN(g29258) );
  NAND2X0 U16461 ( .IN1(n11300), .IN2(n15875), .QN(n15879) );
  NOR2X0 U16462 ( .IN1(n10482), .IN2(n9664), .QN(n11300) );
  NOR2X0 U16463 ( .IN1(n15880), .IN2(n15881), .QN(n15878) );
  NOR2X0 U16464 ( .IN1(g3106), .IN2(n15882), .QN(n15881) );
  NAND2X0 U16465 ( .IN1(n15865), .IN2(g3111), .QN(n15882) );
  NOR2X0 U16466 ( .IN1(n15875), .IN2(n10460), .QN(n15865) );
  NOR2X0 U16467 ( .IN1(n5742), .IN2(n15883), .QN(n15880) );
  NOR2X0 U16468 ( .IN1(n10482), .IN2(n15884), .QN(n15883) );
  NOR2X0 U16469 ( .IN1(n15875), .IN2(g3111), .QN(n15884) );
  OR2X1 U16470 ( .IN1(n15885), .IN2(n12806), .Q(n15875) );
  NAND2X0 U16471 ( .IN1(n15886), .IN2(n15887), .QN(g29257) );
  NAND2X0 U16472 ( .IN1(n10511), .IN2(g3111), .QN(n15887) );
  NAND2X0 U16473 ( .IN1(n15888), .IN2(n10394), .QN(n15886) );
  NAND2X0 U16474 ( .IN1(n15889), .IN2(n15890), .QN(n15888) );
  NAND2X0 U16475 ( .IN1(n12806), .IN2(g3106), .QN(n15890) );
  NAND2X0 U16476 ( .IN1(n15891), .IN2(n12808), .QN(n15889) );
  XNOR2X1 U16477 ( .IN1(n15892), .IN2(n15893), .Q(n15891) );
  NAND2X0 U16478 ( .IN1(g3106), .IN2(n15885), .QN(n15892) );
  NAND2X0 U16479 ( .IN1(n15894), .IN2(n15895), .QN(n15885) );
  NOR2X0 U16480 ( .IN1(n9971), .IN2(n5527), .QN(n15894) );
  NAND2X0 U16481 ( .IN1(n15896), .IN2(n15897), .QN(g29256) );
  NOR2X0 U16482 ( .IN1(n15898), .IN2(n15899), .QN(n15897) );
  NOR2X0 U16483 ( .IN1(n9780), .IN2(n10327), .QN(n15899) );
  NOR2X0 U16484 ( .IN1(n10482), .IN2(n15900), .QN(n15898) );
  NAND2X0 U16485 ( .IN1(n15901), .IN2(g2735), .QN(n15900) );
  NOR2X0 U16486 ( .IN1(n2787), .IN2(n15902), .QN(n15896) );
  NOR2X0 U16487 ( .IN1(n15901), .IN2(g2735), .QN(n15902) );
  INVX0 U16488 ( .INP(n15193), .ZN(n15901) );
  NOR2X0 U16489 ( .IN1(n15903), .IN2(n9780), .QN(n15193) );
  NAND2X0 U16490 ( .IN1(n15904), .IN2(n15905), .QN(g29255) );
  NAND2X0 U16491 ( .IN1(n15906), .IN2(g2638), .QN(n15905) );
  NAND2X0 U16492 ( .IN1(n15907), .IN2(n10394), .QN(n15906) );
  OR2X1 U16493 ( .IN1(n13620), .IN2(n10685), .Q(n15907) );
  NOR2X0 U16494 ( .IN1(n9833), .IN2(n10112), .QN(n10685) );
  INVX0 U16495 ( .INP(n13645), .ZN(n10112) );
  NAND2X0 U16496 ( .IN1(n15908), .IN2(g2652), .QN(n15904) );
  NAND2X0 U16497 ( .IN1(n13626), .IN2(n15909), .QN(n15908) );
  NAND2X0 U16498 ( .IN1(n4379), .IN2(n10394), .QN(n15909) );
  NAND2X0 U16499 ( .IN1(n15910), .IN2(n15911), .QN(g29254) );
  NOR2X0 U16500 ( .IN1(n15912), .IN2(n15913), .QN(n15911) );
  NOR2X0 U16501 ( .IN1(n15914), .IN2(n13627), .QN(n15913) );
  NAND2X0 U16502 ( .IN1(n15915), .IN2(n10394), .QN(n13627) );
  NOR2X0 U16503 ( .IN1(n15916), .IN2(n15917), .QN(n15914) );
  NAND2X0 U16504 ( .IN1(n15918), .IN2(n15919), .QN(n15917) );
  NAND2X0 U16505 ( .IN1(n10042), .IN2(n15920), .QN(n15919) );
  NAND2X0 U16506 ( .IN1(n15921), .IN2(n15922), .QN(n15920) );
  NAND2X0 U16507 ( .IN1(test_so61), .IN2(g2587), .QN(n15922) );
  OR2X1 U16508 ( .IN1(n5508), .IN2(n5787), .Q(n15921) );
  NAND2X0 U16509 ( .IN1(n5508), .IN2(n15923), .QN(n15918) );
  NAND2X0 U16510 ( .IN1(n15924), .IN2(n15925), .QN(n15923) );
  NAND2X0 U16511 ( .IN1(g2610), .IN2(g2583), .QN(n15925) );
  NAND2X0 U16512 ( .IN1(test_so66), .IN2(n5372), .QN(n15924) );
  NOR2X0 U16513 ( .IN1(n5816), .IN2(n13645), .QN(n15916) );
  NAND2X0 U16514 ( .IN1(n5372), .IN2(g2610), .QN(n13645) );
  NOR2X0 U16515 ( .IN1(n9622), .IN2(n15210), .QN(n15912) );
  INVX0 U16516 ( .INP(n15200), .ZN(n15210) );
  NOR2X0 U16517 ( .IN1(n15203), .IN2(n10459), .QN(n15200) );
  NAND2X0 U16518 ( .IN1(n15926), .IN2(n15915), .QN(n15203) );
  INVX0 U16519 ( .INP(n13620), .ZN(n15915) );
  NOR2X0 U16520 ( .IN1(n5508), .IN2(n5372), .QN(n15926) );
  NOR2X0 U16521 ( .IN1(n15927), .IN2(n15928), .QN(n15910) );
  NOR2X0 U16522 ( .IN1(n5508), .IN2(n10327), .QN(n15928) );
  NOR2X0 U16523 ( .IN1(n9832), .IN2(n13626), .QN(n15927) );
  NAND2X0 U16524 ( .IN1(n13620), .IN2(n10395), .QN(n13626) );
  NAND2X0 U16525 ( .IN1(n15929), .IN2(n15161), .QN(n13620) );
  NOR2X0 U16526 ( .IN1(n15930), .IN2(n15931), .QN(n15929) );
  NOR2X0 U16527 ( .IN1(n5609), .IN2(n11658), .QN(n15931) );
  NAND2X0 U16528 ( .IN1(n15932), .IN2(n15933), .QN(g29253) );
  NAND2X0 U16529 ( .IN1(n15934), .IN2(g2518), .QN(n15933) );
  NAND2X0 U16530 ( .IN1(n13661), .IN2(n15935), .QN(n15934) );
  NAND2X0 U16531 ( .IN1(n4391), .IN2(n10395), .QN(n15935) );
  NAND2X0 U16532 ( .IN1(n15936), .IN2(g2504), .QN(n15932) );
  NAND2X0 U16533 ( .IN1(n15937), .IN2(n10395), .QN(n15936) );
  OR2X1 U16534 ( .IN1(n13655), .IN2(n10684), .Q(n15937) );
  NOR2X0 U16535 ( .IN1(n9831), .IN2(n10117), .QN(n10684) );
  INVX0 U16536 ( .INP(n13681), .ZN(n10117) );
  NAND2X0 U16537 ( .IN1(n15938), .IN2(n15939), .QN(g29252) );
  NOR2X0 U16538 ( .IN1(n15940), .IN2(n15941), .QN(n15939) );
  NOR2X0 U16539 ( .IN1(n15942), .IN2(n13662), .QN(n15941) );
  NAND2X0 U16540 ( .IN1(n15943), .IN2(n10395), .QN(n13662) );
  NOR2X0 U16541 ( .IN1(n15944), .IN2(n15945), .QN(n15942) );
  NAND2X0 U16542 ( .IN1(n15946), .IN2(n15947), .QN(n15945) );
  NAND2X0 U16543 ( .IN1(n10043), .IN2(n15948), .QN(n15947) );
  NAND2X0 U16544 ( .IN1(n15949), .IN2(n15950), .QN(n15948) );
  OR2X1 U16545 ( .IN1(n5373), .IN2(n18477), .Q(n15950) );
  OR2X1 U16546 ( .IN1(n5509), .IN2(n5789), .Q(n15949) );
  NAND2X0 U16547 ( .IN1(n5509), .IN2(n15951), .QN(n15946) );
  NAND2X0 U16548 ( .IN1(n15952), .IN2(n15953), .QN(n15951) );
  OR2X1 U16549 ( .IN1(n10043), .IN2(n5798), .Q(n15953) );
  NAND2X0 U16550 ( .IN1(n5373), .IN2(g2441), .QN(n15952) );
  NOR2X0 U16551 ( .IN1(n5814), .IN2(n13681), .QN(n15944) );
  NAND2X0 U16552 ( .IN1(n5373), .IN2(g2476), .QN(n13681) );
  NOR2X0 U16553 ( .IN1(n9624), .IN2(n15244), .QN(n15940) );
  INVX0 U16554 ( .INP(n15234), .ZN(n15244) );
  NOR2X0 U16555 ( .IN1(n15237), .IN2(n10460), .QN(n15234) );
  NAND2X0 U16556 ( .IN1(n15954), .IN2(n15943), .QN(n15237) );
  INVX0 U16557 ( .INP(n13655), .ZN(n15943) );
  NOR2X0 U16558 ( .IN1(n5509), .IN2(n5373), .QN(n15954) );
  NOR2X0 U16559 ( .IN1(n15955), .IN2(n15956), .QN(n15938) );
  NOR2X0 U16560 ( .IN1(n5509), .IN2(n10327), .QN(n15956) );
  NOR2X0 U16561 ( .IN1(n9941), .IN2(n13661), .QN(n15955) );
  NAND2X0 U16562 ( .IN1(n13655), .IN2(n10395), .QN(n13661) );
  NAND2X0 U16563 ( .IN1(n15957), .IN2(n15156), .QN(n13655) );
  NOR2X0 U16564 ( .IN1(n15930), .IN2(n15958), .QN(n15957) );
  NOR2X0 U16565 ( .IN1(n5404), .IN2(n11658), .QN(n15958) );
  NAND2X0 U16566 ( .IN1(n15959), .IN2(n15960), .QN(g29251) );
  NAND2X0 U16567 ( .IN1(n15961), .IN2(g2384), .QN(n15960) );
  NAND2X0 U16568 ( .IN1(n13697), .IN2(n15962), .QN(n15961) );
  NAND2X0 U16569 ( .IN1(n4402), .IN2(n10395), .QN(n15962) );
  NAND2X0 U16570 ( .IN1(n15963), .IN2(g2370), .QN(n15959) );
  NAND2X0 U16571 ( .IN1(n15964), .IN2(n10395), .QN(n15963) );
  OR2X1 U16572 ( .IN1(n13691), .IN2(n10683), .Q(n15964) );
  NOR2X0 U16573 ( .IN1(n9825), .IN2(n401), .QN(n10683) );
  INVX0 U16574 ( .INP(n13717), .ZN(n401) );
  NAND2X0 U16575 ( .IN1(n15965), .IN2(n15966), .QN(g29250) );
  NOR2X0 U16576 ( .IN1(n15967), .IN2(n15968), .QN(n15966) );
  NOR2X0 U16577 ( .IN1(n15969), .IN2(n13698), .QN(n15968) );
  NAND2X0 U16578 ( .IN1(n15970), .IN2(n10395), .QN(n13698) );
  NOR2X0 U16579 ( .IN1(n15971), .IN2(n15972), .QN(n15969) );
  NAND2X0 U16580 ( .IN1(n15973), .IN2(n15974), .QN(n15972) );
  NAND2X0 U16581 ( .IN1(n5511), .IN2(n15975), .QN(n15974) );
  NAND2X0 U16582 ( .IN1(n15976), .IN2(n15977), .QN(n15975) );
  NAND2X0 U16583 ( .IN1(n5375), .IN2(g2307), .QN(n15977) );
  NAND2X0 U16584 ( .IN1(test_so21), .IN2(g2315), .QN(n15976) );
  NAND2X0 U16585 ( .IN1(n15978), .IN2(n10126), .QN(n15973) );
  NAND2X0 U16586 ( .IN1(n15979), .IN2(n15980), .QN(n15978) );
  OR2X1 U16587 ( .IN1(n5375), .IN2(n18473), .Q(n15980) );
  NAND2X0 U16588 ( .IN1(g2351), .IN2(g2303), .QN(n15979) );
  NOR2X0 U16589 ( .IN1(n5815), .IN2(n13717), .QN(n15971) );
  NAND2X0 U16590 ( .IN1(test_so21), .IN2(n5375), .QN(n13717) );
  NOR2X0 U16591 ( .IN1(n9644), .IN2(n15278), .QN(n15967) );
  INVX0 U16592 ( .INP(n15268), .ZN(n15278) );
  NOR2X0 U16593 ( .IN1(n15271), .IN2(n10459), .QN(n15268) );
  NAND2X0 U16594 ( .IN1(n15981), .IN2(n15970), .QN(n15271) );
  INVX0 U16595 ( .INP(n13691), .ZN(n15970) );
  NOR2X0 U16596 ( .IN1(n5511), .IN2(n5375), .QN(n15981) );
  NOR2X0 U16597 ( .IN1(n15982), .IN2(n15983), .QN(n15965) );
  NOR2X0 U16598 ( .IN1(n5511), .IN2(n10328), .QN(n15983) );
  NOR2X0 U16599 ( .IN1(n9826), .IN2(n13697), .QN(n15982) );
  NAND2X0 U16600 ( .IN1(n13691), .IN2(n10395), .QN(n13697) );
  NAND2X0 U16601 ( .IN1(n15984), .IN2(n15985), .QN(n13691) );
  NAND2X0 U16602 ( .IN1(n13370), .IN2(g2807), .QN(n15985) );
  NAND2X0 U16603 ( .IN1(n15986), .IN2(n15987), .QN(g29249) );
  NAND2X0 U16604 ( .IN1(n15988), .IN2(g2250), .QN(n15987) );
  NAND2X0 U16605 ( .IN1(n13733), .IN2(n15989), .QN(n15988) );
  NAND2X0 U16606 ( .IN1(n4414), .IN2(n10396), .QN(n15989) );
  NAND2X0 U16607 ( .IN1(n15990), .IN2(g2236), .QN(n15986) );
  NAND2X0 U16608 ( .IN1(n15991), .IN2(n10396), .QN(n15990) );
  OR2X1 U16609 ( .IN1(n13727), .IN2(n10682), .Q(n15991) );
  NOR2X0 U16610 ( .IN1(n9821), .IN2(n10119), .QN(n10682) );
  INVX0 U16611 ( .INP(n13753), .ZN(n10119) );
  NAND2X0 U16612 ( .IN1(n15992), .IN2(n15993), .QN(g29248) );
  NOR2X0 U16613 ( .IN1(n15994), .IN2(n15995), .QN(n15993) );
  NOR2X0 U16614 ( .IN1(n15996), .IN2(n13734), .QN(n15995) );
  NAND2X0 U16615 ( .IN1(n15997), .IN2(n10396), .QN(n13734) );
  NOR2X0 U16616 ( .IN1(n15998), .IN2(n15999), .QN(n15996) );
  NAND2X0 U16617 ( .IN1(n16000), .IN2(n16001), .QN(n15999) );
  NAND2X0 U16618 ( .IN1(n10045), .IN2(n16002), .QN(n16001) );
  NAND2X0 U16619 ( .IN1(n16003), .IN2(n16004), .QN(n16002) );
  OR2X1 U16620 ( .IN1(n5376), .IN2(n18471), .Q(n16004) );
  OR2X1 U16621 ( .IN1(n5512), .IN2(n5788), .Q(n16003) );
  NAND2X0 U16622 ( .IN1(n5512), .IN2(n16005), .QN(n16000) );
  NAND2X0 U16623 ( .IN1(n16006), .IN2(n16007), .QN(n16005) );
  NAND2X0 U16624 ( .IN1(g2208), .IN2(g2181), .QN(n16007) );
  NAND2X0 U16625 ( .IN1(n5376), .IN2(g2173), .QN(n16006) );
  NOR2X0 U16626 ( .IN1(n5812), .IN2(n13753), .QN(n15998) );
  NAND2X0 U16627 ( .IN1(n5376), .IN2(g2208), .QN(n13753) );
  NOR2X0 U16628 ( .IN1(n9652), .IN2(n15312), .QN(n15994) );
  INVX0 U16629 ( .INP(n15302), .ZN(n15312) );
  NOR2X0 U16630 ( .IN1(n15305), .IN2(n10459), .QN(n15302) );
  NAND2X0 U16631 ( .IN1(n16008), .IN2(n15997), .QN(n15305) );
  INVX0 U16632 ( .INP(n13727), .ZN(n15997) );
  NOR2X0 U16633 ( .IN1(n5512), .IN2(n5376), .QN(n16008) );
  NOR2X0 U16634 ( .IN1(n16009), .IN2(n16010), .QN(n15992) );
  NOR2X0 U16635 ( .IN1(n5512), .IN2(n10328), .QN(n16010) );
  NOR2X0 U16636 ( .IN1(n9822), .IN2(n13733), .QN(n16009) );
  NAND2X0 U16637 ( .IN1(n13727), .IN2(n10396), .QN(n13733) );
  NAND2X0 U16638 ( .IN1(n16011), .IN2(n15160), .QN(n13727) );
  NOR2X0 U16639 ( .IN1(n15930), .IN2(n16012), .QN(n16011) );
  NOR2X0 U16640 ( .IN1(n5545), .IN2(n11658), .QN(n16012) );
  NAND2X0 U16641 ( .IN1(n16013), .IN2(n16014), .QN(g29247) );
  NAND2X0 U16642 ( .IN1(n16015), .IN2(g2079), .QN(n16014) );
  NAND2X0 U16643 ( .IN1(n16016), .IN2(n10396), .QN(n16015) );
  NAND2X0 U16644 ( .IN1(n16017), .IN2(n10681), .QN(n16016) );
  NAND2X0 U16645 ( .IN1(test_so78), .IN2(n13790), .QN(n10681) );
  NAND2X0 U16646 ( .IN1(test_so78), .IN2(n16018), .QN(n16013) );
  NAND2X0 U16647 ( .IN1(n13769), .IN2(n16019), .QN(n16018) );
  NAND2X0 U16648 ( .IN1(n4425), .IN2(n10396), .QN(n16019) );
  NAND2X0 U16649 ( .IN1(n16020), .IN2(n16021), .QN(g29246) );
  NOR2X0 U16650 ( .IN1(n16022), .IN2(n16023), .QN(n16021) );
  NOR2X0 U16651 ( .IN1(n16024), .IN2(n13770), .QN(n16023) );
  NAND2X0 U16652 ( .IN1(n16017), .IN2(n10396), .QN(n13770) );
  NOR2X0 U16653 ( .IN1(n16025), .IN2(n16026), .QN(n16024) );
  NAND2X0 U16654 ( .IN1(n16027), .IN2(n16028), .QN(n16026) );
  NAND2X0 U16655 ( .IN1(n10041), .IN2(n16029), .QN(n16028) );
  NAND2X0 U16656 ( .IN1(n16030), .IN2(n16031), .QN(n16029) );
  OR2X1 U16657 ( .IN1(n5371), .IN2(n18474), .Q(n16031) );
  OR2X1 U16658 ( .IN1(n5507), .IN2(n5790), .Q(n16030) );
  NAND2X0 U16659 ( .IN1(n5507), .IN2(n16032), .QN(n16027) );
  NAND2X0 U16660 ( .IN1(n16033), .IN2(n16034), .QN(n16032) );
  OR2X1 U16661 ( .IN1(n10041), .IN2(n5801), .Q(n16034) );
  NAND2X0 U16662 ( .IN1(n5371), .IN2(g2016), .QN(n16033) );
  NOR2X0 U16663 ( .IN1(n5818), .IN2(n13790), .QN(n16025) );
  NAND2X0 U16664 ( .IN1(n5371), .IN2(g2051), .QN(n13790) );
  NOR2X0 U16665 ( .IN1(n9714), .IN2(n15346), .QN(n16022) );
  INVX0 U16666 ( .INP(n15336), .ZN(n15346) );
  NOR2X0 U16667 ( .IN1(n15339), .IN2(n10459), .QN(n15336) );
  NAND2X0 U16668 ( .IN1(n16035), .IN2(n16017), .QN(n15339) );
  INVX0 U16669 ( .INP(n13763), .ZN(n16017) );
  NOR2X0 U16670 ( .IN1(n5507), .IN2(n5371), .QN(n16035) );
  NOR2X0 U16671 ( .IN1(n16036), .IN2(n16037), .QN(n16020) );
  NOR2X0 U16672 ( .IN1(n5507), .IN2(n10328), .QN(n16037) );
  NOR2X0 U16673 ( .IN1(n9829), .IN2(n13769), .QN(n16036) );
  NAND2X0 U16674 ( .IN1(n13763), .IN2(n10396), .QN(n13769) );
  NAND2X0 U16675 ( .IN1(n16038), .IN2(n15161), .QN(n13763) );
  NOR2X0 U16676 ( .IN1(n15930), .IN2(n16039), .QN(n16038) );
  NOR2X0 U16677 ( .IN1(n5610), .IN2(n11658), .QN(n16039) );
  NAND2X0 U16678 ( .IN1(n16040), .IN2(n16041), .QN(g29245) );
  NAND2X0 U16679 ( .IN1(n16042), .IN2(g1959), .QN(n16041) );
  NAND2X0 U16680 ( .IN1(n13806), .IN2(n16043), .QN(n16042) );
  NAND2X0 U16681 ( .IN1(n4436), .IN2(n10396), .QN(n16043) );
  NAND2X0 U16682 ( .IN1(test_so53), .IN2(n16044), .QN(n16040) );
  NAND2X0 U16683 ( .IN1(n16045), .IN2(n10396), .QN(n16044) );
  OR2X1 U16684 ( .IN1(n13800), .IN2(n10680), .Q(n16045) );
  NOR2X0 U16685 ( .IN1(n9830), .IN2(n10111), .QN(n10680) );
  INVX0 U16686 ( .INP(n13827), .ZN(n10111) );
  NAND2X0 U16687 ( .IN1(n16046), .IN2(n16047), .QN(g29244) );
  NOR2X0 U16688 ( .IN1(n16048), .IN2(n16049), .QN(n16047) );
  NOR2X0 U16689 ( .IN1(n16050), .IN2(n13807), .QN(n16049) );
  NAND2X0 U16690 ( .IN1(n16051), .IN2(n10386), .QN(n13807) );
  NOR2X0 U16691 ( .IN1(n16052), .IN2(n16053), .QN(n16050) );
  NAND2X0 U16692 ( .IN1(n16054), .IN2(n16055), .QN(n16053) );
  NAND2X0 U16693 ( .IN1(n10044), .IN2(n16056), .QN(n16055) );
  NAND2X0 U16694 ( .IN1(n16057), .IN2(n16058), .QN(n16056) );
  OR2X1 U16695 ( .IN1(n5374), .IN2(n18476), .Q(n16058) );
  OR2X1 U16696 ( .IN1(n5510), .IN2(n5793), .Q(n16057) );
  NAND2X0 U16697 ( .IN1(n5510), .IN2(n16059), .QN(n16054) );
  NAND2X0 U16698 ( .IN1(n16060), .IN2(n16061), .QN(n16059) );
  OR2X1 U16699 ( .IN1(n10044), .IN2(n5799), .Q(n16061) );
  NAND2X0 U16700 ( .IN1(n5374), .IN2(g1882), .QN(n16060) );
  NOR2X0 U16701 ( .IN1(n5813), .IN2(n13827), .QN(n16052) );
  NAND2X0 U16702 ( .IN1(n5374), .IN2(g1917), .QN(n13827) );
  NOR2X0 U16703 ( .IN1(n9633), .IN2(n15380), .QN(n16048) );
  INVX0 U16704 ( .INP(n15370), .ZN(n15380) );
  NOR2X0 U16705 ( .IN1(n15373), .IN2(n10458), .QN(n15370) );
  NAND2X0 U16706 ( .IN1(n16062), .IN2(n16051), .QN(n15373) );
  INVX0 U16707 ( .INP(n13800), .ZN(n16051) );
  NOR2X0 U16708 ( .IN1(n5510), .IN2(n5374), .QN(n16062) );
  NOR2X0 U16709 ( .IN1(n16063), .IN2(n16064), .QN(n16046) );
  NOR2X0 U16710 ( .IN1(n5510), .IN2(n10347), .QN(n16064) );
  NOR2X0 U16711 ( .IN1(n10151), .IN2(n13806), .QN(n16063) );
  NAND2X0 U16712 ( .IN1(n13800), .IN2(n10396), .QN(n13806) );
  NAND2X0 U16713 ( .IN1(n16065), .IN2(n15156), .QN(n13800) );
  NOR2X0 U16714 ( .IN1(n15930), .IN2(n16066), .QN(n16065) );
  NOR2X0 U16715 ( .IN1(n5403), .IN2(n11658), .QN(n16066) );
  NAND2X0 U16716 ( .IN1(n16067), .IN2(n16068), .QN(g29243) );
  NAND2X0 U16717 ( .IN1(n16069), .IN2(g1825), .QN(n16068) );
  NAND2X0 U16718 ( .IN1(n13843), .IN2(n16070), .QN(n16069) );
  NAND2X0 U16719 ( .IN1(n4447), .IN2(n10395), .QN(n16070) );
  NAND2X0 U16720 ( .IN1(n16071), .IN2(g1811), .QN(n16067) );
  NAND2X0 U16721 ( .IN1(n16072), .IN2(n10395), .QN(n16071) );
  OR2X1 U16722 ( .IN1(n13837), .IN2(n10679), .Q(n16072) );
  NOR2X0 U16723 ( .IN1(n9823), .IN2(n10115), .QN(n10679) );
  INVX0 U16724 ( .INP(n13862), .ZN(n10115) );
  NAND2X0 U16725 ( .IN1(n16073), .IN2(n16074), .QN(g29242) );
  NOR2X0 U16726 ( .IN1(n16075), .IN2(n16076), .QN(n16074) );
  NOR2X0 U16727 ( .IN1(n16077), .IN2(n13844), .QN(n16076) );
  NAND2X0 U16728 ( .IN1(n16078), .IN2(n10394), .QN(n13844) );
  NOR2X0 U16729 ( .IN1(n16079), .IN2(n16080), .QN(n16077) );
  NAND2X0 U16730 ( .IN1(n16081), .IN2(n16082), .QN(n16080) );
  NAND2X0 U16731 ( .IN1(n5359), .IN2(n16083), .QN(n16082) );
  NAND2X0 U16732 ( .IN1(n16084), .IN2(n16085), .QN(n16083) );
  NAND2X0 U16733 ( .IN1(g1783), .IN2(g1756), .QN(n16085) );
  NAND2X0 U16734 ( .IN1(n5602), .IN2(g1748), .QN(n16084) );
  NAND2X0 U16735 ( .IN1(n5596), .IN2(n16086), .QN(n16081) );
  NAND2X0 U16736 ( .IN1(n16087), .IN2(n16088), .QN(n16086) );
  OR2X1 U16737 ( .IN1(n5359), .IN2(n5795), .Q(n16088) );
  OR2X1 U16738 ( .IN1(n5602), .IN2(n5797), .Q(n16087) );
  NOR2X0 U16739 ( .IN1(n5817), .IN2(n13862), .QN(n16079) );
  NAND2X0 U16740 ( .IN1(n5602), .IN2(g1783), .QN(n13862) );
  NOR2X0 U16741 ( .IN1(n9704), .IN2(n15414), .QN(n16075) );
  INVX0 U16742 ( .INP(n15404), .ZN(n15414) );
  NOR2X0 U16743 ( .IN1(n15407), .IN2(n10458), .QN(n15404) );
  NAND2X0 U16744 ( .IN1(n16089), .IN2(n16078), .QN(n15407) );
  INVX0 U16745 ( .INP(n13837), .ZN(n16078) );
  NOR2X0 U16746 ( .IN1(n5602), .IN2(n5359), .QN(n16089) );
  NOR2X0 U16747 ( .IN1(n16090), .IN2(n16091), .QN(n16073) );
  NOR2X0 U16748 ( .IN1(n5359), .IN2(n10350), .QN(n16091) );
  NOR2X0 U16749 ( .IN1(n9824), .IN2(n13843), .QN(n16090) );
  NAND2X0 U16750 ( .IN1(n13837), .IN2(n10394), .QN(n13843) );
  NAND2X0 U16751 ( .IN1(n15984), .IN2(n16092), .QN(n13837) );
  NAND2X0 U16752 ( .IN1(n13370), .IN2(g2775), .QN(n16092) );
  INVX0 U16753 ( .INP(n11658), .ZN(n13370) );
  NOR2X0 U16754 ( .IN1(n4411), .IN2(n15930), .QN(n15984) );
  NAND2X0 U16755 ( .IN1(n5465), .IN2(g2715), .QN(n4411) );
  NAND2X0 U16756 ( .IN1(n16093), .IN2(n16094), .QN(g29241) );
  NAND2X0 U16757 ( .IN1(n16095), .IN2(g1691), .QN(n16094) );
  NAND2X0 U16758 ( .IN1(n13878), .IN2(n16096), .QN(n16095) );
  NAND2X0 U16759 ( .IN1(n4458), .IN2(n10393), .QN(n16096) );
  NAND2X0 U16760 ( .IN1(n16097), .IN2(g1677), .QN(n16093) );
  NAND2X0 U16761 ( .IN1(n16098), .IN2(n10392), .QN(n16097) );
  OR2X1 U16762 ( .IN1(n13872), .IN2(n10678), .Q(n16098) );
  NOR2X0 U16763 ( .IN1(n9827), .IN2(n1019), .QN(n10678) );
  NAND2X0 U16764 ( .IN1(n16099), .IN2(n16100), .QN(g29240) );
  NOR2X0 U16765 ( .IN1(n16101), .IN2(n16102), .QN(n16100) );
  NOR2X0 U16766 ( .IN1(n9828), .IN2(n13878), .QN(n16102) );
  NAND2X0 U16767 ( .IN1(n13872), .IN2(n10392), .QN(n13878) );
  NOR2X0 U16768 ( .IN1(n16103), .IN2(n13879), .QN(n16101) );
  NAND2X0 U16769 ( .IN1(n16104), .IN2(n10392), .QN(n13879) );
  NOR2X0 U16770 ( .IN1(n16105), .IN2(n16106), .QN(n16103) );
  NAND2X0 U16771 ( .IN1(n16107), .IN2(n16108), .QN(n16106) );
  NAND2X0 U16772 ( .IN1(n1019), .IN2(g1600), .QN(n16108) );
  INVX0 U16773 ( .INP(n13900), .ZN(n1019) );
  NAND2X0 U16774 ( .IN1(test_so94), .IN2(n5370), .QN(n13900) );
  NAND2X0 U16775 ( .IN1(g31863), .IN2(g1620), .QN(n16107) );
  NOR2X0 U16776 ( .IN1(g1657), .IN2(n10121), .QN(g31863) );
  NAND2X0 U16777 ( .IN1(n16109), .IN2(n16110), .QN(n16105) );
  NAND2X0 U16778 ( .IN1(n16111), .IN2(n5525), .QN(n16110) );
  AND2X1 U16779 ( .IN1(g1612), .IN2(n5370), .Q(n16111) );
  NAND2X0 U16780 ( .IN1(n16112), .IN2(n10121), .QN(n16109) );
  NAND2X0 U16781 ( .IN1(n16113), .IN2(n16114), .QN(n16112) );
  OR2X1 U16782 ( .IN1(n5370), .IN2(n18475), .Q(n16114) );
  OR2X1 U16783 ( .IN1(n5525), .IN2(n5792), .Q(n16113) );
  NOR2X0 U16784 ( .IN1(n16115), .IN2(n16116), .QN(n16099) );
  NOR2X0 U16785 ( .IN1(n5525), .IN2(n10354), .QN(n16116) );
  NOR2X0 U16786 ( .IN1(n9623), .IN2(n15442), .QN(n16115) );
  NAND2X0 U16787 ( .IN1(n16117), .IN2(n16104), .QN(n15442) );
  INVX0 U16788 ( .INP(n13872), .ZN(n16104) );
  NAND2X0 U16789 ( .IN1(n16118), .IN2(n15160), .QN(n13872) );
  NOR2X0 U16790 ( .IN1(g2719), .IN2(g2715), .QN(n15160) );
  NOR2X0 U16791 ( .IN1(n15930), .IN2(n16119), .QN(n16118) );
  NOR2X0 U16792 ( .IN1(n5544), .IN2(n11658), .QN(n16119) );
  NOR2X0 U16793 ( .IN1(n4388), .IN2(n11658), .QN(n15930) );
  NAND2X0 U16794 ( .IN1(n9780), .IN2(n5301), .QN(n11658) );
  NOR2X0 U16795 ( .IN1(n5525), .IN2(n5370), .QN(n16117) );
  NAND2X0 U16796 ( .IN1(n16120), .IN2(n16121), .QN(g29239) );
  NAND2X0 U16797 ( .IN1(n16122), .IN2(n16123), .QN(n16121) );
  INVX0 U16798 ( .INP(n16124), .ZN(n16123) );
  NOR2X0 U16799 ( .IN1(n16125), .IN2(n16126), .QN(n16122) );
  NOR2X0 U16800 ( .IN1(n16127), .IN2(n16128), .QN(n16120) );
  NOR2X0 U16801 ( .IN1(n10481), .IN2(n16129), .QN(n16128) );
  NAND2X0 U16802 ( .IN1(n16130), .IN2(g1454), .QN(n16129) );
  NAND2X0 U16803 ( .IN1(n16131), .IN2(n16126), .QN(n16130) );
  XOR2X1 U16804 ( .IN1(n5343), .IN2(n16132), .Q(n16126) );
  INVX0 U16805 ( .INP(n16125), .ZN(n16131) );
  NOR2X0 U16806 ( .IN1(n5289), .IN2(n10355), .QN(n16127) );
  NAND2X0 U16807 ( .IN1(n16133), .IN2(n16134), .QN(g29238) );
  NAND2X0 U16808 ( .IN1(n16135), .IN2(g1484), .QN(n16134) );
  NOR2X0 U16809 ( .IN1(n16136), .IN2(n16137), .QN(n16133) );
  NOR2X0 U16810 ( .IN1(n10481), .IN2(n16138), .QN(n16137) );
  NAND2X0 U16811 ( .IN1(n16139), .IN2(n16140), .QN(n16138) );
  NAND2X0 U16812 ( .IN1(n5865), .IN2(n16141), .QN(n16140) );
  NAND2X0 U16813 ( .IN1(n16142), .IN2(n16143), .QN(n16141) );
  NOR2X0 U16814 ( .IN1(g1442), .IN2(g1489), .QN(n16142) );
  XOR2X1 U16815 ( .IN1(g1300), .IN2(n16132), .Q(n16139) );
  NOR2X0 U16816 ( .IN1(n5290), .IN2(n10355), .QN(n16136) );
  NAND2X0 U16817 ( .IN1(n16144), .IN2(n16145), .QN(g29237) );
  NAND2X0 U16818 ( .IN1(n16146), .IN2(n16147), .QN(n16145) );
  NOR2X0 U16819 ( .IN1(n10127), .IN2(n16124), .QN(n16147) );
  NOR2X0 U16820 ( .IN1(n16148), .IN2(n16149), .QN(n16146) );
  NOR2X0 U16821 ( .IN1(n16150), .IN2(n16151), .QN(n16144) );
  NOR2X0 U16822 ( .IN1(n10481), .IN2(n16152), .QN(n16151) );
  NAND2X0 U16823 ( .IN1(n16153), .IN2(g1467), .QN(n16152) );
  NAND2X0 U16824 ( .IN1(n16154), .IN2(n16155), .QN(n16153) );
  AND2X1 U16825 ( .IN1(n16149), .IN2(test_so49), .Q(n16154) );
  XOR2X1 U16826 ( .IN1(n5290), .IN2(n16132), .Q(n16149) );
  NOR2X0 U16827 ( .IN1(n5343), .IN2(n10356), .QN(n16150) );
  NAND2X0 U16828 ( .IN1(n16156), .IN2(n16157), .QN(g29236) );
  NAND2X0 U16829 ( .IN1(n16158), .IN2(n16159), .QN(n16157) );
  NOR2X0 U16830 ( .IN1(test_so49), .IN2(n16124), .QN(n16159) );
  NAND2X0 U16831 ( .IN1(n16160), .IN2(n5850), .QN(n16124) );
  NOR2X0 U16832 ( .IN1(n16148), .IN2(n16161), .QN(n16158) );
  NOR2X0 U16833 ( .IN1(n16162), .IN2(n16163), .QN(n16156) );
  NOR2X0 U16834 ( .IN1(n10481), .IN2(n16164), .QN(n16163) );
  NAND2X0 U16835 ( .IN1(n16165), .IN2(g1437), .QN(n16164) );
  NAND2X0 U16836 ( .IN1(n16166), .IN2(n16155), .QN(n16165) );
  INVX0 U16837 ( .INP(n16148), .ZN(n16155) );
  AND2X1 U16838 ( .IN1(n10127), .IN2(n16161), .Q(n16166) );
  XOR2X1 U16839 ( .IN1(n5289), .IN2(n16132), .Q(n16161) );
  AND2X1 U16840 ( .IN1(n13057), .IN2(DFF_1092_n1), .Q(n16132) );
  INVX0 U16841 ( .INP(n11259), .ZN(n13057) );
  NOR2X0 U16842 ( .IN1(n10049), .IN2(n10353), .QN(n16162) );
  NAND2X0 U16843 ( .IN1(n16167), .IN2(n16168), .QN(g29235) );
  NAND2X0 U16844 ( .IN1(n10511), .IN2(g1252), .QN(n16168) );
  NOR2X0 U16845 ( .IN1(n16169), .IN2(n16170), .QN(n16167) );
  NOR2X0 U16846 ( .IN1(g1256), .IN2(n16171), .QN(n16170) );
  NOR2X0 U16847 ( .IN1(n5558), .IN2(n16172), .QN(n16169) );
  NAND2X0 U16848 ( .IN1(n13309), .IN2(n16171), .QN(n16172) );
  INVX0 U16849 ( .INP(n4178), .ZN(n16171) );
  NAND2X0 U16850 ( .IN1(n16173), .IN2(n16174), .QN(g29234) );
  NAND2X0 U16851 ( .IN1(n16175), .IN2(n16176), .QN(n16174) );
  INVX0 U16852 ( .INP(n16177), .ZN(n16176) );
  NOR2X0 U16853 ( .IN1(n16178), .IN2(n16179), .QN(n16175) );
  NOR2X0 U16854 ( .IN1(n16180), .IN2(n16181), .QN(n16173) );
  NOR2X0 U16855 ( .IN1(n10481), .IN2(n16182), .QN(n16181) );
  NAND2X0 U16856 ( .IN1(test_so90), .IN2(n16183), .QN(n16182) );
  NAND2X0 U16857 ( .IN1(n16184), .IN2(n16179), .QN(n16183) );
  XNOR2X1 U16858 ( .IN1(n16185), .IN2(n5478), .Q(n16179) );
  INVX0 U16859 ( .INP(n16178), .ZN(n16184) );
  NOR2X0 U16860 ( .IN1(n5328), .IN2(n10356), .QN(n16180) );
  NAND2X0 U16861 ( .IN1(n16186), .IN2(n16187), .QN(g29233) );
  NAND2X0 U16862 ( .IN1(n16188), .IN2(g1141), .QN(n16187) );
  NOR2X0 U16863 ( .IN1(n16189), .IN2(n16190), .QN(n16186) );
  NOR2X0 U16864 ( .IN1(n10481), .IN2(n16191), .QN(n16190) );
  NAND2X0 U16865 ( .IN1(n16192), .IN2(n16193), .QN(n16191) );
  NAND2X0 U16866 ( .IN1(n5691), .IN2(n16194), .QN(n16193) );
  NAND2X0 U16867 ( .IN1(n16195), .IN2(n16196), .QN(n16194) );
  NOR2X0 U16868 ( .IN1(test_so7), .IN2(g1146), .QN(n16195) );
  XOR2X1 U16869 ( .IN1(n16185), .IN2(n5341), .Q(n16192) );
  NOR2X0 U16870 ( .IN1(n5329), .IN2(n10355), .QN(n16189) );
  NAND2X0 U16871 ( .IN1(n16197), .IN2(n16198), .QN(g29232) );
  NAND2X0 U16872 ( .IN1(n16199), .IN2(n16200), .QN(n16198) );
  NOR2X0 U16873 ( .IN1(n5599), .IN2(n16177), .QN(n16200) );
  NOR2X0 U16874 ( .IN1(n16201), .IN2(n16202), .QN(n16199) );
  NOR2X0 U16875 ( .IN1(n16203), .IN2(n16204), .QN(n16197) );
  NOR2X0 U16876 ( .IN1(n10481), .IN2(n16205), .QN(n16204) );
  NAND2X0 U16877 ( .IN1(n16206), .IN2(g1124), .QN(n16205) );
  NAND2X0 U16878 ( .IN1(n16207), .IN2(n16208), .QN(n16206) );
  AND2X1 U16879 ( .IN1(g1183), .IN2(n16202), .Q(n16207) );
  XNOR2X1 U16880 ( .IN1(n16185), .IN2(n5329), .Q(n16202) );
  NOR2X0 U16881 ( .IN1(n5478), .IN2(n10356), .QN(n16203) );
  NAND2X0 U16882 ( .IN1(n16209), .IN2(n16210), .QN(g29231) );
  NAND2X0 U16883 ( .IN1(n16211), .IN2(n16212), .QN(n16210) );
  NOR2X0 U16884 ( .IN1(g1183), .IN2(n16177), .QN(n16212) );
  NAND2X0 U16885 ( .IN1(n16213), .IN2(n5851), .QN(n16177) );
  NOR2X0 U16886 ( .IN1(n16201), .IN2(n16214), .QN(n16211) );
  NOR2X0 U16887 ( .IN1(n16215), .IN2(n16216), .QN(n16209) );
  NOR2X0 U16888 ( .IN1(n10481), .IN2(n16217), .QN(n16216) );
  NAND2X0 U16889 ( .IN1(n16218), .IN2(g1094), .QN(n16217) );
  NAND2X0 U16890 ( .IN1(n16219), .IN2(n16208), .QN(n16218) );
  INVX0 U16891 ( .INP(n16201), .ZN(n16208) );
  AND2X1 U16892 ( .IN1(n16214), .IN2(n5599), .Q(n16219) );
  XNOR2X1 U16893 ( .IN1(n16185), .IN2(n5328), .Q(n16214) );
  NAND2X0 U16894 ( .IN1(n11355), .IN2(DFF_24_n1), .QN(n16185) );
  AND2X1 U16895 ( .IN1(n10496), .IN2(test_so7), .Q(n16215) );
  NAND2X0 U16896 ( .IN1(n16220), .IN2(n16221), .QN(g29230) );
  NAND2X0 U16897 ( .IN1(n10511), .IN2(g907), .QN(n16221) );
  NOR2X0 U16898 ( .IN1(n16222), .IN2(n16223), .QN(n16220) );
  NOR2X0 U16899 ( .IN1(g911), .IN2(n16224), .QN(n16223) );
  NOR2X0 U16900 ( .IN1(n5559), .IN2(n16225), .QN(n16222) );
  NAND2X0 U16901 ( .IN1(n13328), .IN2(n16224), .QN(n16225) );
  INVX0 U16902 ( .INP(n4196), .ZN(n16224) );
  NAND2X0 U16903 ( .IN1(n16226), .IN2(n16227), .QN(g29229) );
  NAND2X0 U16904 ( .IN1(n10511), .IN2(g827), .QN(n16227) );
  NOR2X0 U16905 ( .IN1(n16228), .IN2(n16229), .QN(n16226) );
  NOR2X0 U16906 ( .IN1(g723), .IN2(n16230), .QN(n16229) );
  NAND2X0 U16907 ( .IN1(n4516), .IN2(n16231), .QN(n16230) );
  AND2X1 U16908 ( .IN1(n4517), .IN2(g723), .Q(n16228) );
  NAND2X0 U16909 ( .IN1(n16232), .IN2(n16233), .QN(g29228) );
  NAND2X0 U16910 ( .IN1(n2404), .IN2(n16234), .QN(n16233) );
  XNOR2X1 U16911 ( .IN1(test_so60), .IN2(n15555), .Q(n16234) );
  NAND2X0 U16912 ( .IN1(n16235), .IN2(n16236), .QN(n15555) );
  NAND2X0 U16913 ( .IN1(n5482), .IN2(g12184), .QN(n16236) );
  NAND2X0 U16914 ( .IN1(n10511), .IN2(g736), .QN(n16232) );
  NAND2X0 U16915 ( .IN1(n16237), .IN2(n16238), .QN(g29227) );
  NAND2X0 U16916 ( .IN1(n10511), .IN2(g676), .QN(n16238) );
  NOR2X0 U16917 ( .IN1(n16239), .IN2(n16240), .QN(n16237) );
  AND2X1 U16918 ( .IN1(n4524), .IN2(test_so70), .Q(n16240) );
  NOR2X0 U16919 ( .IN1(test_so70), .IN2(n16241), .QN(n16239) );
  NAND2X0 U16920 ( .IN1(n4523), .IN2(n16242), .QN(n16241) );
  NAND2X0 U16921 ( .IN1(n16243), .IN2(n16244), .QN(g29226) );
  OR2X1 U16922 ( .IN1(n10309), .IN2(n9626), .Q(n16244) );
  NOR2X0 U16923 ( .IN1(n16245), .IN2(n16246), .QN(n16243) );
  NOR2X0 U16924 ( .IN1(g676), .IN2(n16247), .QN(n16246) );
  NAND2X0 U16925 ( .IN1(n4526), .IN2(n16242), .QN(n16247) );
  NOR2X0 U16926 ( .IN1(n5751), .IN2(n16248), .QN(n16245) );
  NAND2X0 U16927 ( .IN1(n4525), .IN2(n16249), .QN(n16248) );
  INVX0 U16928 ( .INP(n4526), .ZN(n16249) );
  NAND2X0 U16929 ( .IN1(n16250), .IN2(n16251), .QN(g29225) );
  NAND2X0 U16930 ( .IN1(n16252), .IN2(n4525), .QN(n16251) );
  AND2X1 U16931 ( .IN1(n16242), .IN2(n10365), .Q(n4525) );
  AND2X1 U16932 ( .IN1(g703), .IN2(n16253), .Q(n16242) );
  NAND2X0 U16933 ( .IN1(n16254), .IN2(n16255), .QN(n16253) );
  NOR2X0 U16934 ( .IN1(n9734), .IN2(n10107), .QN(n16255) );
  NOR2X0 U16935 ( .IN1(n16256), .IN2(n4535), .QN(n16254) );
  XOR2X1 U16936 ( .IN1(n9819), .IN2(n9820), .Q(n4535) );
  XOR2X1 U16937 ( .IN1(n10107), .IN2(n9626), .Q(n16252) );
  NAND2X0 U16938 ( .IN1(n10511), .IN2(g667), .QN(n16250) );
  NAND2X0 U16939 ( .IN1(n16257), .IN2(n16258), .QN(g29224) );
  NAND2X0 U16940 ( .IN1(n10511), .IN2(g572), .QN(n16258) );
  NOR2X0 U16941 ( .IN1(n16259), .IN2(n16260), .QN(n16257) );
  NOR2X0 U16942 ( .IN1(g586), .IN2(n16261), .QN(n16260) );
  NOR2X0 U16943 ( .IN1(n5336), .IN2(n16262), .QN(n16259) );
  NAND2X0 U16944 ( .IN1(n2421), .IN2(n16261), .QN(n16262) );
  INVX0 U16945 ( .INP(n4201), .ZN(n16261) );
  NAND2X0 U16946 ( .IN1(n16263), .IN2(n16264), .QN(g29223) );
  NAND2X0 U16947 ( .IN1(n16265), .IN2(n5708), .QN(n16264) );
  NOR2X0 U16948 ( .IN1(n16266), .IN2(n16267), .QN(n16263) );
  NOR2X0 U16949 ( .IN1(n10481), .IN2(n16268), .QN(n16267) );
  NOR2X0 U16950 ( .IN1(n16269), .IN2(n4962), .QN(n16268) );
  NOR2X0 U16951 ( .IN1(n5708), .IN2(n16265), .QN(n16269) );
  NOR2X0 U16952 ( .IN1(n16270), .IN2(n5820), .QN(n16265) );
  NOR2X0 U16953 ( .IN1(n5820), .IN2(n10356), .QN(n16266) );
  NAND2X0 U16954 ( .IN1(n16271), .IN2(n16272), .QN(g29222) );
  NAND2X0 U16955 ( .IN1(n16273), .IN2(g411), .QN(n16272) );
  NOR2X0 U16956 ( .IN1(n16274), .IN2(n16275), .QN(n16271) );
  NOR2X0 U16957 ( .IN1(g417), .IN2(n16276), .QN(n16275) );
  NAND2X0 U16958 ( .IN1(n16277), .IN2(n3676), .QN(n16276) );
  NOR2X0 U16959 ( .IN1(n5358), .IN2(n16278), .QN(n16274) );
  NOR2X0 U16960 ( .IN1(n10481), .IN2(n16279), .QN(n16278) );
  NOR2X0 U16961 ( .IN1(n3676), .IN2(n16280), .QN(n16279) );
  XOR2X1 U16962 ( .IN1(g417), .IN2(n16281), .Q(n3676) );
  NOR2X0 U16963 ( .IN1(n16282), .IN2(n16283), .QN(n16281) );
  NOR2X0 U16964 ( .IN1(g392), .IN2(n16284), .QN(n16283) );
  NOR2X0 U16965 ( .IN1(n16285), .IN2(n16286), .QN(n16284) );
  NOR2X0 U16966 ( .IN1(n9746), .IN2(g405), .QN(n16286) );
  NOR2X0 U16967 ( .IN1(n9748), .IN2(n9747), .QN(n16285) );
  NOR2X0 U16968 ( .IN1(n9778), .IN2(n16287), .QN(n16282) );
  NOR2X0 U16969 ( .IN1(n16288), .IN2(n16289), .QN(n16287) );
  NOR2X0 U16970 ( .IN1(n9748), .IN2(n9726), .QN(n16289) );
  NOR2X0 U16971 ( .IN1(n9747), .IN2(g405), .QN(n16288) );
  NAND2X0 U16972 ( .IN1(n16290), .IN2(n16291), .QN(g28105) );
  NAND2X0 U16973 ( .IN1(n12658), .IN2(g5011), .QN(n16291) );
  NOR2X0 U16974 ( .IN1(n16292), .IN2(n16293), .QN(n16290) );
  NOR2X0 U16975 ( .IN1(n10481), .IN2(n16294), .QN(n16293) );
  NAND2X0 U16976 ( .IN1(n12655), .IN2(n15608), .QN(n16294) );
  NAND2X0 U16977 ( .IN1(n16295), .IN2(n16296), .QN(n15608) );
  NOR2X0 U16978 ( .IN1(n16297), .IN2(n16298), .QN(n16296) );
  NOR2X0 U16979 ( .IN1(n5531), .IN2(n16299), .QN(n16298) );
  NOR2X0 U16980 ( .IN1(n16300), .IN2(n16301), .QN(n16299) );
  NAND2X0 U16981 ( .IN1(n16302), .IN2(n16303), .QN(n16301) );
  NAND2X0 U16982 ( .IN1(n10671), .IN2(n16304), .QN(n16303) );
  NAND2X0 U16983 ( .IN1(n16305), .IN2(n16306), .QN(n16304) );
  NAND2X0 U16984 ( .IN1(g6723), .IN2(g6589), .QN(n16306) );
  NAND2X0 U16985 ( .IN1(g13099), .IN2(g6581), .QN(n16305) );
  NAND2X0 U16986 ( .IN1(n10675), .IN2(n16307), .QN(n16302) );
  NAND2X0 U16987 ( .IN1(n16308), .IN2(n16309), .QN(n16307) );
  NAND2X0 U16988 ( .IN1(g6609), .IN2(g17871), .QN(n16309) );
  NAND2X0 U16989 ( .IN1(test_so80), .IN2(test_so71), .QN(n16308) );
  NAND2X0 U16990 ( .IN1(n16310), .IN2(n16311), .QN(n16300) );
  NAND2X0 U16991 ( .IN1(n16312), .IN2(n16313), .QN(n16311) );
  NOR2X0 U16992 ( .IN1(n9947), .IN2(n5584), .QN(n16312) );
  NAND2X0 U16993 ( .IN1(n15611), .IN2(n16314), .QN(n16310) );
  NAND2X0 U16994 ( .IN1(n16315), .IN2(n16316), .QN(n16314) );
  OR2X1 U16995 ( .IN1(n9799), .IN2(n9995), .Q(n16316) );
  NAND2X0 U16996 ( .IN1(g6641), .IN2(g17764), .QN(n16315) );
  NOR2X0 U16997 ( .IN1(n16317), .IN2(g6727), .QN(n16297) );
  NOR2X0 U16998 ( .IN1(n16318), .IN2(n16319), .QN(n16317) );
  NAND2X0 U16999 ( .IN1(n16320), .IN2(n16321), .QN(n16319) );
  NAND2X0 U17000 ( .IN1(n10675), .IN2(n16322), .QN(n16321) );
  NAND2X0 U17001 ( .IN1(n16323), .IN2(n16324), .QN(n16322) );
  NAND2X0 U17002 ( .IN1(g17764), .IN2(g6649), .QN(n16324) );
  OR2X1 U17003 ( .IN1(n9995), .IN2(n9996), .Q(n16323) );
  NAND2X0 U17004 ( .IN1(n16313), .IN2(n16325), .QN(n16320) );
  NAND2X0 U17005 ( .IN1(n16326), .IN2(n16327), .QN(n16325) );
  NAND2X0 U17006 ( .IN1(g6723), .IN2(g6605), .QN(n16327) );
  NAND2X0 U17007 ( .IN1(g13099), .IN2(g6593), .QN(n16326) );
  NAND2X0 U17008 ( .IN1(n16328), .IN2(n16329), .QN(n16318) );
  NAND2X0 U17009 ( .IN1(n16330), .IN2(n10671), .QN(n16329) );
  NOR2X0 U17010 ( .IN1(n9992), .IN2(n5584), .QN(n16330) );
  NAND2X0 U17011 ( .IN1(n15611), .IN2(n16331), .QN(n16328) );
  NAND2X0 U17012 ( .IN1(n16332), .IN2(n16333), .QN(n16331) );
  NAND2X0 U17013 ( .IN1(g17871), .IN2(g6617), .QN(n16333) );
  NAND2X0 U17014 ( .IN1(test_so80), .IN2(g6601), .QN(n16332) );
  NOR2X0 U17015 ( .IN1(n16334), .IN2(n16335), .QN(n16295) );
  NOR2X0 U17016 ( .IN1(n16336), .IN2(n16337), .QN(n16335) );
  NOR2X0 U17017 ( .IN1(n16338), .IN2(n16339), .QN(n16336) );
  NAND2X0 U17018 ( .IN1(n16340), .IN2(n16341), .QN(n16339) );
  NAND2X0 U17019 ( .IN1(n16342), .IN2(n10671), .QN(n16341) );
  INVX0 U17020 ( .INP(n16343), .ZN(n10671) );
  NOR2X0 U17021 ( .IN1(n9859), .IN2(n5700), .QN(n16342) );
  NAND2X0 U17022 ( .IN1(n16344), .IN2(n10675), .QN(n16340) );
  NOR2X0 U17023 ( .IN1(g6682), .IN2(n5398), .QN(n10675) );
  NOR2X0 U17024 ( .IN1(n9890), .IN2(n9858), .QN(n16344) );
  NOR2X0 U17025 ( .IN1(n10672), .IN2(n16345), .QN(n16338) );
  NAND2X0 U17026 ( .IN1(g6653), .IN2(g17688), .QN(n16345) );
  NOR2X0 U17027 ( .IN1(n16346), .IN2(n16347), .QN(n16334) );
  INVX0 U17028 ( .INP(n16337), .ZN(n16347) );
  XOR2X1 U17029 ( .IN1(test_so80), .IN2(n5531), .Q(n16337) );
  NOR2X0 U17030 ( .IN1(n16348), .IN2(n16349), .QN(n16346) );
  NAND2X0 U17031 ( .IN1(n16350), .IN2(n16351), .QN(n16349) );
  NAND2X0 U17032 ( .IN1(n16352), .IN2(n16313), .QN(n16351) );
  INVX0 U17033 ( .INP(n10672), .ZN(n16313) );
  NAND2X0 U17034 ( .IN1(n5398), .IN2(g6682), .QN(n10672) );
  NOR2X0 U17035 ( .IN1(n9840), .IN2(n5700), .QN(n16352) );
  NAND2X0 U17036 ( .IN1(n16353), .IN2(n15611), .QN(n16350) );
  INVX0 U17037 ( .INP(n10676), .ZN(n15611) );
  NAND2X0 U17038 ( .IN1(g6682), .IN2(g6741), .QN(n10676) );
  NOR2X0 U17039 ( .IN1(n9891), .IN2(n9890), .QN(n16353) );
  NOR2X0 U17040 ( .IN1(n16343), .IN2(n16354), .QN(n16348) );
  NAND2X0 U17041 ( .IN1(g17688), .IN2(g6645), .QN(n16354) );
  NAND2X0 U17042 ( .IN1(n5590), .IN2(n5398), .QN(n16343) );
  NOR2X0 U17043 ( .IN1(n9799), .IN2(n10354), .QN(n16292) );
  NAND2X0 U17044 ( .IN1(n16355), .IN2(n16356), .QN(g28102) );
  NAND2X0 U17045 ( .IN1(n12678), .IN2(g4826), .QN(n16356) );
  NOR2X0 U17046 ( .IN1(n16357), .IN2(n16358), .QN(n16355) );
  NOR2X0 U17047 ( .IN1(n10481), .IN2(n16359), .QN(n16358) );
  NAND2X0 U17048 ( .IN1(n12675), .IN2(n15649), .QN(n16359) );
  NAND2X0 U17049 ( .IN1(n16360), .IN2(n16361), .QN(n15649) );
  NOR2X0 U17050 ( .IN1(n16362), .IN2(n16363), .QN(n16361) );
  NOR2X0 U17051 ( .IN1(test_so69), .IN2(n16364), .QN(n16363) );
  NOR2X0 U17052 ( .IN1(n16365), .IN2(n16366), .QN(n16364) );
  NAND2X0 U17053 ( .IN1(n16367), .IN2(n16368), .QN(n16366) );
  NAND2X0 U17054 ( .IN1(n16369), .IN2(n16370), .QN(n16368) );
  NAND2X0 U17055 ( .IN1(n16371), .IN2(n16372), .QN(n16370) );
  NAND2X0 U17056 ( .IN1(g6377), .IN2(g6259), .QN(n16372) );
  NAND2X0 U17057 ( .IN1(g13085), .IN2(g6247), .QN(n16371) );
  NAND2X0 U17058 ( .IN1(n16373), .IN2(n16374), .QN(n16367) );
  NAND2X0 U17059 ( .IN1(n16375), .IN2(n16376), .QN(n16374) );
  NAND2X0 U17060 ( .IN1(g12422), .IN2(g6255), .QN(n16376) );
  NAND2X0 U17061 ( .IN1(g17845), .IN2(g6271), .QN(n16375) );
  NAND2X0 U17062 ( .IN1(n16377), .IN2(n16378), .QN(n16365) );
  NAND2X0 U17063 ( .IN1(n16379), .IN2(n16380), .QN(n16378) );
  NOR2X0 U17064 ( .IN1(n5586), .IN2(n10002), .QN(n16379) );
  NAND2X0 U17065 ( .IN1(n12674), .IN2(n16381), .QN(n16377) );
  NAND2X0 U17066 ( .IN1(n16382), .IN2(n16383), .QN(n16381) );
  NAND2X0 U17067 ( .IN1(g17743), .IN2(g6303), .QN(n16383) );
  NAND2X0 U17068 ( .IN1(g17685), .IN2(g6251), .QN(n16382) );
  NOR2X0 U17069 ( .IN1(n16384), .IN2(n10130), .QN(n16362) );
  NOR2X0 U17070 ( .IN1(n16385), .IN2(n16386), .QN(n16384) );
  NAND2X0 U17071 ( .IN1(n16387), .IN2(n16388), .QN(n16386) );
  NAND2X0 U17072 ( .IN1(n16373), .IN2(n16389), .QN(n16388) );
  NAND2X0 U17073 ( .IN1(n16390), .IN2(n16391), .QN(n16389) );
  NAND2X0 U17074 ( .IN1(g17743), .IN2(g6295), .QN(n16391) );
  OR2X1 U17075 ( .IN1(n10005), .IN2(n9806), .Q(n16390) );
  NAND2X0 U17076 ( .IN1(n16380), .IN2(n16392), .QN(n16387) );
  NAND2X0 U17077 ( .IN1(n16393), .IN2(n16394), .QN(n16392) );
  NAND2X0 U17078 ( .IN1(g6377), .IN2(g6243), .QN(n16394) );
  NAND2X0 U17079 ( .IN1(g13085), .IN2(g6235), .QN(n16393) );
  NAND2X0 U17080 ( .IN1(n16395), .IN2(n16396), .QN(n16385) );
  NAND2X0 U17081 ( .IN1(n16397), .IN2(n16369), .QN(n16396) );
  NOR2X0 U17082 ( .IN1(n9949), .IN2(n5586), .QN(n16397) );
  NAND2X0 U17083 ( .IN1(n12674), .IN2(n16398), .QN(n16395) );
  NAND2X0 U17084 ( .IN1(n16399), .IN2(n16400), .QN(n16398) );
  NAND2X0 U17085 ( .IN1(g12422), .IN2(g6239), .QN(n16400) );
  NAND2X0 U17086 ( .IN1(g6263), .IN2(g17845), .QN(n16399) );
  NOR2X0 U17087 ( .IN1(n16401), .IN2(n16402), .QN(n16360) );
  NOR2X0 U17088 ( .IN1(n16403), .IN2(n16404), .QN(n16402) );
  NOR2X0 U17089 ( .IN1(n16405), .IN2(n16406), .QN(n16403) );
  NAND2X0 U17090 ( .IN1(n16407), .IN2(n16408), .QN(n16406) );
  NAND2X0 U17091 ( .IN1(n16409), .IN2(n16369), .QN(n16408) );
  NOR2X0 U17092 ( .IN1(n9879), .IN2(n9863), .QN(n16409) );
  NAND2X0 U17093 ( .IN1(n16410), .IN2(n12674), .QN(n16407) );
  NOR2X0 U17094 ( .IN1(n9894), .IN2(n9864), .QN(n16410) );
  NOR2X0 U17095 ( .IN1(n16411), .IN2(n16412), .QN(n16405) );
  NAND2X0 U17096 ( .IN1(g14779), .IN2(g6275), .QN(n16412) );
  NOR2X0 U17097 ( .IN1(n16413), .IN2(n16414), .QN(n16401) );
  INVX0 U17098 ( .INP(n16404), .ZN(n16414) );
  XNOR2X1 U17099 ( .IN1(g12422), .IN2(test_so69), .Q(n16404) );
  NOR2X0 U17100 ( .IN1(n16415), .IN2(n16416), .QN(n16413) );
  NAND2X0 U17101 ( .IN1(n16417), .IN2(n16418), .QN(n16416) );
  NAND2X0 U17102 ( .IN1(n16419), .IN2(n16369), .QN(n16418) );
  INVX0 U17103 ( .INP(n12671), .ZN(n16369) );
  NOR2X0 U17104 ( .IN1(n9842), .IN2(n5703), .QN(n16419) );
  NAND2X0 U17105 ( .IN1(n16420), .IN2(n16380), .QN(n16417) );
  NOR2X0 U17106 ( .IN1(n9880), .IN2(n9879), .QN(n16420) );
  NOR2X0 U17107 ( .IN1(n11715), .IN2(n16421), .QN(n16415) );
  OR2X1 U17108 ( .IN1(n9894), .IN2(n9895), .Q(n16421) );
  NOR2X0 U17109 ( .IN1(n9806), .IN2(n10354), .QN(n16357) );
  NAND2X0 U17110 ( .IN1(n16422), .IN2(n16423), .QN(g28099) );
  NAND2X0 U17111 ( .IN1(test_so13), .IN2(n10515), .QN(n16423) );
  NOR2X0 U17112 ( .IN1(n16424), .IN2(n16425), .QN(n16422) );
  NOR2X0 U17113 ( .IN1(n9668), .IN2(n12700), .QN(n16425) );
  NOR2X0 U17114 ( .IN1(n15687), .IN2(n12705), .QN(n16424) );
  NAND2X0 U17115 ( .IN1(n12695), .IN2(n10390), .QN(n12705) );
  AND2X1 U17116 ( .IN1(n16426), .IN2(n16427), .Q(n15687) );
  NOR2X0 U17117 ( .IN1(n16428), .IN2(n16429), .QN(n16427) );
  NOR2X0 U17118 ( .IN1(n5528), .IN2(n16430), .QN(n16429) );
  NOR2X0 U17119 ( .IN1(n16431), .IN2(n16432), .QN(n16430) );
  NAND2X0 U17120 ( .IN1(n16433), .IN2(n16434), .QN(n16432) );
  NAND2X0 U17121 ( .IN1(n15690), .IN2(n16435), .QN(n16434) );
  NAND2X0 U17122 ( .IN1(n16436), .IN2(n16437), .QN(n16435) );
  NAND2X0 U17123 ( .IN1(g5949), .IN2(g17715), .QN(n16437) );
  NAND2X0 U17124 ( .IN1(test_so13), .IN2(g17646), .QN(n16436) );
  NAND2X0 U17125 ( .IN1(n16438), .IN2(n16439), .QN(n16433) );
  NAND2X0 U17126 ( .IN1(n16440), .IN2(n16441), .QN(n16439) );
  NAND2X0 U17127 ( .IN1(g6031), .IN2(g5897), .QN(n16441) );
  NAND2X0 U17128 ( .IN1(g13068), .IN2(g5889), .QN(n16440) );
  NAND2X0 U17129 ( .IN1(n16442), .IN2(n16443), .QN(n16431) );
  NAND2X0 U17130 ( .IN1(n16444), .IN2(n16445), .QN(n16443) );
  NOR2X0 U17131 ( .IN1(n9944), .IN2(n5581), .QN(n16444) );
  NAND2X0 U17132 ( .IN1(n12694), .IN2(n16446), .QN(n16442) );
  NAND2X0 U17133 ( .IN1(n16447), .IN2(n16448), .QN(n16446) );
  NAND2X0 U17134 ( .IN1(g12350), .IN2(g5893), .QN(n16448) );
  NAND2X0 U17135 ( .IN1(test_so28), .IN2(g17819), .QN(n16447) );
  NOR2X0 U17136 ( .IN1(n16449), .IN2(g6035), .QN(n16428) );
  NOR2X0 U17137 ( .IN1(n16450), .IN2(n16451), .QN(n16449) );
  NAND2X0 U17138 ( .IN1(n16452), .IN2(n16453), .QN(n16451) );
  NAND2X0 U17139 ( .IN1(n16445), .IN2(n16454), .QN(n16453) );
  NAND2X0 U17140 ( .IN1(n16455), .IN2(n16456), .QN(n16454) );
  NAND2X0 U17141 ( .IN1(g6031), .IN2(g5913), .QN(n16456) );
  NAND2X0 U17142 ( .IN1(g13068), .IN2(g5901), .QN(n16455) );
  NAND2X0 U17143 ( .IN1(n15690), .IN2(n16457), .QN(n16452) );
  NAND2X0 U17144 ( .IN1(n16458), .IN2(n16459), .QN(n16457) );
  NAND2X0 U17145 ( .IN1(g12350), .IN2(g5909), .QN(n16459) );
  NAND2X0 U17146 ( .IN1(g17819), .IN2(g5925), .QN(n16458) );
  NAND2X0 U17147 ( .IN1(n16460), .IN2(n16461), .QN(n16450) );
  NAND2X0 U17148 ( .IN1(n16462), .IN2(n16438), .QN(n16461) );
  NOR2X0 U17149 ( .IN1(n9978), .IN2(n5581), .QN(n16462) );
  NAND2X0 U17150 ( .IN1(n12694), .IN2(n16463), .QN(n16460) );
  NAND2X0 U17151 ( .IN1(n16464), .IN2(n16465), .QN(n16463) );
  NAND2X0 U17152 ( .IN1(g17715), .IN2(g5957), .QN(n16465) );
  NAND2X0 U17153 ( .IN1(g17646), .IN2(g5905), .QN(n16464) );
  NOR2X0 U17154 ( .IN1(n16466), .IN2(n16467), .QN(n16426) );
  NOR2X0 U17155 ( .IN1(n16468), .IN2(n16469), .QN(n16467) );
  NOR2X0 U17156 ( .IN1(n16470), .IN2(n16471), .QN(n16468) );
  NAND2X0 U17157 ( .IN1(n16472), .IN2(n16473), .QN(n16471) );
  NAND2X0 U17158 ( .IN1(n16474), .IN2(n16445), .QN(n16473) );
  NOR2X0 U17159 ( .IN1(n9837), .IN2(n5698), .QN(n16474) );
  NAND2X0 U17160 ( .IN1(n16475), .IN2(n16438), .QN(n16472) );
  NOR2X0 U17161 ( .IN1(n9871), .IN2(n9870), .QN(n16475) );
  NOR2X0 U17162 ( .IN1(n11711), .IN2(n16476), .QN(n16470) );
  OR2X1 U17163 ( .IN1(n9885), .IN2(n9886), .Q(n16476) );
  NOR2X0 U17164 ( .IN1(n16477), .IN2(n16478), .QN(n16466) );
  INVX0 U17165 ( .INP(n16469), .ZN(n16478) );
  XNOR2X1 U17166 ( .IN1(g12350), .IN2(n5528), .Q(n16469) );
  NOR2X0 U17167 ( .IN1(n16479), .IN2(n16480), .QN(n16477) );
  NAND2X0 U17168 ( .IN1(n16481), .IN2(n16482), .QN(n16480) );
  NAND2X0 U17169 ( .IN1(n16483), .IN2(n16445), .QN(n16482) );
  INVX0 U17170 ( .INP(n12691), .ZN(n16445) );
  NOR2X0 U17171 ( .IN1(n9870), .IN2(n9848), .QN(n16483) );
  NAND2X0 U17172 ( .IN1(n16484), .IN2(n12694), .QN(n16481) );
  NOR2X0 U17173 ( .IN1(n9885), .IN2(n9849), .QN(n16484) );
  NOR2X0 U17174 ( .IN1(n16485), .IN2(n16486), .QN(n16479) );
  NAND2X0 U17175 ( .IN1(g14738), .IN2(g5929), .QN(n16486) );
  NAND2X0 U17176 ( .IN1(n16487), .IN2(n16488), .QN(g28096) );
  NAND2X0 U17177 ( .IN1(n12720), .IN2(g4821), .QN(n16488) );
  NOR2X0 U17178 ( .IN1(n16489), .IN2(n16490), .QN(n16487) );
  NOR2X0 U17179 ( .IN1(n10481), .IN2(n16491), .QN(n16490) );
  NAND2X0 U17180 ( .IN1(n12717), .IN2(n15727), .QN(n16491) );
  NAND2X0 U17181 ( .IN1(n16492), .IN2(n16493), .QN(n15727) );
  NOR2X0 U17182 ( .IN1(n16494), .IN2(n16495), .QN(n16493) );
  NOR2X0 U17183 ( .IN1(n5529), .IN2(n16496), .QN(n16495) );
  NOR2X0 U17184 ( .IN1(n16497), .IN2(n16498), .QN(n16496) );
  NAND2X0 U17185 ( .IN1(n16499), .IN2(n16500), .QN(n16498) );
  NAND2X0 U17186 ( .IN1(n15730), .IN2(n16501), .QN(n16500) );
  NAND2X0 U17187 ( .IN1(n16502), .IN2(n16503), .QN(n16501) );
  OR2X1 U17188 ( .IN1(n9795), .IN2(n9986), .Q(n16503) );
  NAND2X0 U17189 ( .IN1(g5603), .IN2(g17678), .QN(n16502) );
  NAND2X0 U17190 ( .IN1(n16504), .IN2(n16505), .QN(n16499) );
  NAND2X0 U17191 ( .IN1(n16506), .IN2(n16507), .QN(n16505) );
  NAND2X0 U17192 ( .IN1(g5685), .IN2(g5551), .QN(n16507) );
  NAND2X0 U17193 ( .IN1(g13049), .IN2(g5543), .QN(n16506) );
  NAND2X0 U17194 ( .IN1(n16508), .IN2(n16509), .QN(n16497) );
  NAND2X0 U17195 ( .IN1(n16510), .IN2(n16511), .QN(n16509) );
  NOR2X0 U17196 ( .IN1(n9945), .IN2(n5582), .QN(n16510) );
  NAND2X0 U17197 ( .IN1(n12716), .IN2(n16512), .QN(n16508) );
  NAND2X0 U17198 ( .IN1(n16513), .IN2(n16514), .QN(n16512) );
  NAND2X0 U17199 ( .IN1(g12300), .IN2(g5547), .QN(n16514) );
  NAND2X0 U17200 ( .IN1(g5571), .IN2(g17813), .QN(n16513) );
  NOR2X0 U17201 ( .IN1(n16515), .IN2(g5689), .QN(n16494) );
  NOR2X0 U17202 ( .IN1(n16516), .IN2(n16517), .QN(n16515) );
  NAND2X0 U17203 ( .IN1(n16518), .IN2(n16519), .QN(n16517) );
  NAND2X0 U17204 ( .IN1(n16511), .IN2(n16520), .QN(n16519) );
  NAND2X0 U17205 ( .IN1(n16521), .IN2(n16522), .QN(n16520) );
  NAND2X0 U17206 ( .IN1(g5685), .IN2(g5567), .QN(n16522) );
  NAND2X0 U17207 ( .IN1(g13049), .IN2(g5555), .QN(n16521) );
  NAND2X0 U17208 ( .IN1(n15730), .IN2(n16523), .QN(n16518) );
  NAND2X0 U17209 ( .IN1(n16524), .IN2(n16525), .QN(n16523) );
  NAND2X0 U17210 ( .IN1(g12300), .IN2(g5563), .QN(n16525) );
  NAND2X0 U17211 ( .IN1(g17813), .IN2(g5579), .QN(n16524) );
  NAND2X0 U17212 ( .IN1(n16526), .IN2(n16527), .QN(n16516) );
  NAND2X0 U17213 ( .IN1(n16528), .IN2(n16504), .QN(n16527) );
  NOR2X0 U17214 ( .IN1(n9983), .IN2(n5582), .QN(n16528) );
  NAND2X0 U17215 ( .IN1(n12716), .IN2(n16529), .QN(n16526) );
  NAND2X0 U17216 ( .IN1(n16530), .IN2(n16531), .QN(n16529) );
  NAND2X0 U17217 ( .IN1(g17678), .IN2(g5611), .QN(n16531) );
  NAND2X0 U17218 ( .IN1(test_so6), .IN2(g17604), .QN(n16530) );
  NOR2X0 U17219 ( .IN1(n16532), .IN2(n16533), .QN(n16492) );
  NOR2X0 U17220 ( .IN1(n16534), .IN2(n16535), .QN(n16533) );
  NOR2X0 U17221 ( .IN1(n16536), .IN2(n16537), .QN(n16534) );
  NAND2X0 U17222 ( .IN1(n16538), .IN2(n16539), .QN(n16537) );
  NAND2X0 U17223 ( .IN1(n16540), .IN2(n16511), .QN(n16539) );
  NOR2X0 U17224 ( .IN1(n9838), .IN2(n5705), .QN(n16540) );
  NAND2X0 U17225 ( .IN1(n16541), .IN2(n16504), .QN(n16538) );
  NOR2X0 U17226 ( .IN1(n9873), .IN2(n9872), .QN(n16541) );
  NOR2X0 U17227 ( .IN1(n10147), .IN2(n16542), .QN(n16536) );
  OR2X1 U17228 ( .IN1(n11704), .IN2(n9887), .Q(n16542) );
  NOR2X0 U17229 ( .IN1(n16543), .IN2(n16544), .QN(n16532) );
  INVX0 U17230 ( .INP(n16535), .ZN(n16544) );
  XNOR2X1 U17231 ( .IN1(g12300), .IN2(n5529), .Q(n16535) );
  NOR2X0 U17232 ( .IN1(n16545), .IN2(n16546), .QN(n16543) );
  NAND2X0 U17233 ( .IN1(n16547), .IN2(n16548), .QN(n16546) );
  NAND2X0 U17234 ( .IN1(n16549), .IN2(n16511), .QN(n16548) );
  INVX0 U17235 ( .INP(n12713), .ZN(n16511) );
  NOR2X0 U17236 ( .IN1(n9872), .IN2(n9851), .QN(n16549) );
  NAND2X0 U17237 ( .IN1(n16550), .IN2(n12716), .QN(n16547) );
  NOR2X0 U17238 ( .IN1(n9887), .IN2(n9852), .QN(n16550) );
  NOR2X0 U17239 ( .IN1(n16551), .IN2(n16552), .QN(n16545) );
  NAND2X0 U17240 ( .IN1(g14694), .IN2(g5583), .QN(n16552) );
  NOR2X0 U17241 ( .IN1(n9795), .IN2(n10353), .QN(n16489) );
  NAND2X0 U17242 ( .IN1(n16553), .IN2(n16554), .QN(g28093) );
  NAND2X0 U17243 ( .IN1(n12737), .IN2(g29220), .QN(n16554) );
  NOR2X0 U17244 ( .IN1(n16555), .IN2(n16556), .QN(n16553) );
  NOR2X0 U17245 ( .IN1(n10481), .IN2(n16557), .QN(n16556) );
  NAND2X0 U17246 ( .IN1(g33959), .IN2(n15767), .QN(n16557) );
  NAND2X0 U17247 ( .IN1(n16558), .IN2(n16559), .QN(n15767) );
  NOR2X0 U17248 ( .IN1(n16560), .IN2(n16561), .QN(n16559) );
  NOR2X0 U17249 ( .IN1(test_so10), .IN2(n16562), .QN(n16561) );
  NOR2X0 U17250 ( .IN1(n16563), .IN2(n16564), .QN(n16562) );
  NAND2X0 U17251 ( .IN1(n16565), .IN2(n16566), .QN(n16564) );
  NAND2X0 U17252 ( .IN1(n16567), .IN2(n16568), .QN(n16566) );
  NAND2X0 U17253 ( .IN1(n16569), .IN2(n16570), .QN(n16568) );
  NAND2X0 U17254 ( .IN1(g5220), .IN2(g5339), .QN(n16570) );
  NAND2X0 U17255 ( .IN1(g5208), .IN2(g13039), .QN(n16569) );
  NAND2X0 U17256 ( .IN1(n10665), .IN2(n16571), .QN(n16565) );
  NAND2X0 U17257 ( .IN1(n16572), .IN2(n16573), .QN(n16571) );
  NAND2X0 U17258 ( .IN1(g17639), .IN2(g5264), .QN(n16573) );
  OR2X1 U17259 ( .IN1(n9976), .IN2(n9977), .Q(n16572) );
  NAND2X0 U17260 ( .IN1(n16574), .IN2(n16575), .QN(n16563) );
  NAND2X0 U17261 ( .IN1(n16576), .IN2(n10661), .QN(n16575) );
  NOR2X0 U17262 ( .IN1(n9973), .IN2(n5579), .QN(n16576) );
  NAND2X0 U17263 ( .IN1(g25114), .IN2(n16577), .QN(n16574) );
  NAND2X0 U17264 ( .IN1(n16578), .IN2(n16579), .QN(n16577) );
  NAND2X0 U17265 ( .IN1(g12238), .IN2(g5216), .QN(n16579) );
  NAND2X0 U17266 ( .IN1(g17787), .IN2(g5232), .QN(n16578) );
  NOR2X0 U17267 ( .IN1(n16580), .IN2(n10129), .QN(n16560) );
  NOR2X0 U17268 ( .IN1(n16581), .IN2(n16582), .QN(n16580) );
  NAND2X0 U17269 ( .IN1(n16583), .IN2(n16584), .QN(n16582) );
  NAND2X0 U17270 ( .IN1(n10665), .IN2(n16585), .QN(n16584) );
  NAND2X0 U17271 ( .IN1(n16586), .IN2(n16587), .QN(n16585) );
  NAND2X0 U17272 ( .IN1(g12238), .IN2(g5200), .QN(n16587) );
  NAND2X0 U17273 ( .IN1(g5224), .IN2(g17787), .QN(n16586) );
  NAND2X0 U17274 ( .IN1(n10661), .IN2(n16588), .QN(n16583) );
  NAND2X0 U17275 ( .IN1(n16589), .IN2(n16590), .QN(n16588) );
  NAND2X0 U17276 ( .IN1(g5339), .IN2(g5204), .QN(n16590) );
  NAND2X0 U17277 ( .IN1(g13039), .IN2(g5196), .QN(n16589) );
  INVX0 U17278 ( .INP(n16591), .ZN(n10661) );
  NAND2X0 U17279 ( .IN1(n16592), .IN2(n16593), .QN(n16581) );
  NAND2X0 U17280 ( .IN1(n16594), .IN2(n16567), .QN(n16593) );
  NOR2X0 U17281 ( .IN1(n9943), .IN2(n5579), .QN(n16594) );
  NAND2X0 U17282 ( .IN1(g25114), .IN2(n16595), .QN(n16592) );
  NAND2X0 U17283 ( .IN1(n16596), .IN2(n16597), .QN(n16595) );
  OR2X1 U17284 ( .IN1(n9810), .IN2(n9976), .Q(n16597) );
  NAND2X0 U17285 ( .IN1(g5256), .IN2(g17639), .QN(n16596) );
  NOR2X0 U17286 ( .IN1(n16598), .IN2(n16599), .QN(n16558) );
  NOR2X0 U17287 ( .IN1(n16600), .IN2(n16601), .QN(n16599) );
  NOR2X0 U17288 ( .IN1(n16602), .IN2(n16603), .QN(n16600) );
  NAND2X0 U17289 ( .IN1(n16604), .IN2(n16605), .QN(n16603) );
  NAND2X0 U17290 ( .IN1(n16606), .IN2(n16567), .QN(n16605) );
  INVX0 U17291 ( .INP(n10662), .ZN(n16567) );
  NOR2X0 U17292 ( .IN1(n9868), .IN2(n9845), .QN(n16606) );
  NAND2X0 U17293 ( .IN1(n16607), .IN2(n10665), .QN(n16604) );
  NOR2X0 U17294 ( .IN1(g5297), .IN2(n5393), .QN(n10665) );
  NOR2X0 U17295 ( .IN1(n9883), .IN2(n9846), .QN(n16607) );
  NOR2X0 U17296 ( .IN1(n16591), .IN2(n16608), .QN(n16602) );
  NAND2X0 U17297 ( .IN1(g14662), .IN2(g5236), .QN(n16608) );
  NOR2X0 U17298 ( .IN1(n16609), .IN2(n16610), .QN(n16598) );
  INVX0 U17299 ( .INP(n16601), .ZN(n16610) );
  XNOR2X1 U17300 ( .IN1(g12238), .IN2(test_so10), .Q(n16601) );
  NOR2X0 U17301 ( .IN1(n16611), .IN2(n16612), .QN(n16609) );
  NAND2X0 U17302 ( .IN1(n16613), .IN2(n16614), .QN(n16612) );
  NAND2X0 U17303 ( .IN1(n16615), .IN2(test_so82), .QN(n16614) );
  NOR2X0 U17304 ( .IN1(n5704), .IN2(n10662), .QN(n16615) );
  NAND2X0 U17305 ( .IN1(n5393), .IN2(g5297), .QN(n10662) );
  NAND2X0 U17306 ( .IN1(n16616), .IN2(g25114), .QN(n16613) );
  NOR2X0 U17307 ( .IN1(n9884), .IN2(n9883), .QN(n16616) );
  NOR2X0 U17308 ( .IN1(n16591), .IN2(n16617), .QN(n16611) );
  NAND2X0 U17309 ( .IN1(g17519), .IN2(g5260), .QN(n16617) );
  NAND2X0 U17310 ( .IN1(n5588), .IN2(n5393), .QN(n16591) );
  NOR2X0 U17311 ( .IN1(n9810), .IN2(n10355), .QN(n16555) );
  NAND2X0 U17312 ( .IN1(n16618), .IN2(n16619), .QN(g28092) );
  NAND2X0 U17313 ( .IN1(n10511), .IN2(g5057), .QN(n16619) );
  NAND2X0 U17314 ( .IN1(n16620), .IN2(n10390), .QN(n16618) );
  NOR2X0 U17315 ( .IN1(n14050), .IN2(n14052), .QN(n16620) );
  AND2X1 U17316 ( .IN1(n16621), .IN2(n16622), .Q(n14052) );
  NOR2X0 U17317 ( .IN1(g5046), .IN2(n16623), .QN(n16622) );
  NOR2X0 U17318 ( .IN1(n16624), .IN2(g5041), .QN(n16621) );
  AND2X1 U17319 ( .IN1(n16625), .IN2(n16626), .Q(n14050) );
  NOR2X0 U17320 ( .IN1(g84), .IN2(n16623), .QN(n16626) );
  NAND2X0 U17321 ( .IN1(g5057), .IN2(g5022), .QN(n16623) );
  NOR2X0 U17322 ( .IN1(g5046), .IN2(g5052), .QN(n16625) );
  NAND2X0 U17323 ( .IN1(n16627), .IN2(n16628), .QN(g28091) );
  NAND2X0 U17324 ( .IN1(n10511), .IN2(g5069), .QN(n16628) );
  NAND2X0 U17325 ( .IN1(n16629), .IN2(n10390), .QN(n16627) );
  NOR2X0 U17326 ( .IN1(n14049), .IN2(n14051), .QN(n16629) );
  AND2X1 U17327 ( .IN1(n16630), .IN2(n16631), .Q(n14051) );
  NOR2X0 U17328 ( .IN1(n5578), .IN2(n16632), .QN(n16631) );
  NAND2X0 U17329 ( .IN1(g5041), .IN2(g5062), .QN(n16632) );
  NOR2X0 U17330 ( .IN1(g5057), .IN2(n16624), .QN(n16630) );
  INVX0 U17331 ( .INP(g84), .ZN(n16624) );
  AND2X1 U17332 ( .IN1(n16633), .IN2(n16634), .Q(n14049) );
  NOR2X0 U17333 ( .IN1(n5578), .IN2(n16635), .QN(n16634) );
  NAND2X0 U17334 ( .IN1(g5052), .IN2(g5062), .QN(n16635) );
  NOR2X0 U17335 ( .IN1(g84), .IN2(g5057), .QN(n16633) );
  NAND2X0 U17336 ( .IN1(n16636), .IN2(n16637), .QN(g28090) );
  NAND2X0 U17337 ( .IN1(n16638), .IN2(n11759), .QN(n16637) );
  NOR2X0 U17338 ( .IN1(n10757), .IN2(n10744), .QN(n11759) );
  NOR2X0 U17339 ( .IN1(n10480), .IN2(n16639), .QN(n16638) );
  NOR2X0 U17340 ( .IN1(n16640), .IN2(g4961), .QN(n16639) );
  NOR2X0 U17341 ( .IN1(n16641), .IN2(n12766), .QN(n16640) );
  NOR2X0 U17342 ( .IN1(n16642), .IN2(n16643), .QN(n16641) );
  NAND2X0 U17343 ( .IN1(n16644), .IN2(n16645), .QN(n16643) );
  NAND2X0 U17344 ( .IN1(n15815), .IN2(g4049), .QN(n16645) );
  NAND2X0 U17345 ( .IN1(n9905), .IN2(n12767), .QN(n16644) );
  NAND2X0 U17346 ( .IN1(n16646), .IN2(n16647), .QN(n16642) );
  OR2X1 U17347 ( .IN1(n12764), .IN2(n9906), .Q(n16647) );
  NAND2X0 U17348 ( .IN1(n9906), .IN2(n16648), .QN(n16646) );
  NAND2X0 U17349 ( .IN1(n12771), .IN2(g4961), .QN(n16636) );
  NAND2X0 U17350 ( .IN1(n16649), .IN2(n16650), .QN(g28089) );
  NAND2X0 U17351 ( .IN1(n16651), .IN2(n11768), .QN(n16650) );
  NOR2X0 U17352 ( .IN1(n10757), .IN2(n10743), .QN(n11768) );
  NOR2X0 U17353 ( .IN1(n10485), .IN2(n16652), .QN(n16651) );
  NOR2X0 U17354 ( .IN1(n16653), .IN2(g4950), .QN(n16652) );
  NOR2X0 U17355 ( .IN1(n16654), .IN2(n12786), .QN(n16653) );
  NOR2X0 U17356 ( .IN1(n16655), .IN2(n16656), .QN(n16654) );
  NAND2X0 U17357 ( .IN1(n16657), .IN2(n16658), .QN(n16656) );
  NAND2X0 U17358 ( .IN1(n15855), .IN2(g3698), .QN(n16658) );
  NAND2X0 U17359 ( .IN1(n9901), .IN2(n12787), .QN(n16657) );
  NAND2X0 U17360 ( .IN1(n16659), .IN2(n16660), .QN(n16655) );
  OR2X1 U17361 ( .IN1(n12784), .IN2(n9902), .Q(n16660) );
  NAND2X0 U17362 ( .IN1(n9902), .IN2(n16661), .QN(n16659) );
  NAND2X0 U17363 ( .IN1(n12791), .IN2(g4950), .QN(n16649) );
  NAND2X0 U17364 ( .IN1(n16662), .IN2(n16663), .QN(g28088) );
  NAND2X0 U17365 ( .IN1(n16664), .IN2(n11776), .QN(n16663) );
  NOR2X0 U17366 ( .IN1(n10757), .IN2(n10754), .QN(n11776) );
  NOR2X0 U17367 ( .IN1(n10480), .IN2(n16665), .QN(n16664) );
  NOR2X0 U17368 ( .IN1(n16666), .IN2(g4939), .QN(n16665) );
  NOR2X0 U17369 ( .IN1(n16667), .IN2(n12806), .QN(n16666) );
  NOR2X0 U17370 ( .IN1(n16668), .IN2(n16669), .QN(n16667) );
  NAND2X0 U17371 ( .IN1(n16670), .IN2(n16671), .QN(n16669) );
  NAND2X0 U17372 ( .IN1(n15895), .IN2(g3347), .QN(n16671) );
  NAND2X0 U17373 ( .IN1(n9896), .IN2(n12807), .QN(n16670) );
  NAND2X0 U17374 ( .IN1(n16672), .IN2(n16673), .QN(n16668) );
  OR2X1 U17375 ( .IN1(n16674), .IN2(n9897), .Q(n16673) );
  NAND2X0 U17376 ( .IN1(n9897), .IN2(n16675), .QN(n16672) );
  NAND2X0 U17377 ( .IN1(n12811), .IN2(g4939), .QN(n16662) );
  NAND2X0 U17378 ( .IN1(n16676), .IN2(n16677), .QN(g28087) );
  NAND2X0 U17379 ( .IN1(n16678), .IN2(n11783), .QN(n16677) );
  NOR2X0 U17380 ( .IN1(n10757), .IN2(n10746), .QN(n11783) );
  NAND2X0 U17381 ( .IN1(n16679), .IN2(g4983), .QN(n10757) );
  NOR2X0 U17382 ( .IN1(test_so58), .IN2(n5706), .QN(n16679) );
  NOR2X0 U17383 ( .IN1(n10480), .IN2(n16680), .QN(n16678) );
  NOR2X0 U17384 ( .IN1(n4689), .IN2(g4894), .QN(n16680) );
  NAND2X0 U17385 ( .IN1(n12658), .IN2(g4894), .QN(n16676) );
  NOR2X0 U17386 ( .IN1(n12655), .IN2(n10461), .QN(n12658) );
  NOR2X0 U17387 ( .IN1(n5713), .IN2(n16681), .QN(n12655) );
  AND2X1 U17388 ( .IN1(n12602), .IN2(n16682), .Q(n16681) );
  NOR2X0 U17389 ( .IN1(n5863), .IN2(n10754), .QN(n12602) );
  NAND2X0 U17390 ( .IN1(n5517), .IN2(n5360), .QN(n10754) );
  NAND2X0 U17391 ( .IN1(n16683), .IN2(n16684), .QN(g28086) );
  NAND2X0 U17392 ( .IN1(n16685), .IN2(n11797), .QN(n16684) );
  NOR2X0 U17393 ( .IN1(n10699), .IN2(n10713), .QN(n11797) );
  NOR2X0 U17394 ( .IN1(n10480), .IN2(n16686), .QN(n16685) );
  NOR2X0 U17395 ( .IN1(n16687), .IN2(g4771), .QN(n16686) );
  NOR2X0 U17396 ( .IN1(n16688), .IN2(n12673), .QN(n16687) );
  NOR2X0 U17397 ( .IN1(n16689), .IN2(n16690), .QN(n16688) );
  NAND2X0 U17398 ( .IN1(n16691), .IN2(n16692), .QN(n16690) );
  NAND2X0 U17399 ( .IN1(n16373), .IN2(g6390), .QN(n16692) );
  INVX0 U17400 ( .INP(n11715), .ZN(n16373) );
  NAND2X0 U17401 ( .IN1(g6336), .IN2(g6395), .QN(n11715) );
  NAND2X0 U17402 ( .IN1(n9898), .IN2(n12674), .QN(n16691) );
  NOR2X0 U17403 ( .IN1(g6336), .IN2(n5396), .QN(n12674) );
  NAND2X0 U17404 ( .IN1(n16693), .IN2(n16694), .QN(n16689) );
  OR2X1 U17405 ( .IN1(n12671), .IN2(n9899), .Q(n16694) );
  NAND2X0 U17406 ( .IN1(n5396), .IN2(g6336), .QN(n12671) );
  NAND2X0 U17407 ( .IN1(n9899), .IN2(n16380), .QN(n16693) );
  INVX0 U17408 ( .INP(n16411), .ZN(n16380) );
  NAND2X0 U17409 ( .IN1(n5592), .IN2(n5396), .QN(n16411) );
  NAND2X0 U17410 ( .IN1(n12678), .IN2(g4771), .QN(n16683) );
  NOR2X0 U17411 ( .IN1(n12675), .IN2(n10457), .QN(n12678) );
  INVX0 U17412 ( .INP(n12673), .ZN(n12675) );
  NAND2X0 U17413 ( .IN1(g4688), .IN2(n16695), .QN(n12673) );
  NAND2X0 U17414 ( .IN1(n12645), .IN2(n16696), .QN(n16695) );
  NOR2X0 U17415 ( .IN1(n5613), .IN2(n16697), .QN(n12645) );
  NAND2X0 U17416 ( .IN1(n16698), .IN2(n16699), .QN(g28085) );
  NAND2X0 U17417 ( .IN1(n16700), .IN2(n11806), .QN(n16699) );
  NOR2X0 U17418 ( .IN1(n10699), .IN2(n10714), .QN(n11806) );
  NOR2X0 U17419 ( .IN1(n10480), .IN2(n16701), .QN(n16700) );
  NOR2X0 U17420 ( .IN1(n16702), .IN2(g4760), .QN(n16701) );
  NOR2X0 U17421 ( .IN1(n16703), .IN2(n12693), .QN(n16702) );
  NOR2X0 U17422 ( .IN1(n16704), .IN2(n16705), .QN(n16703) );
  NAND2X0 U17423 ( .IN1(n16706), .IN2(n16707), .QN(n16705) );
  NAND2X0 U17424 ( .IN1(n12694), .IN2(n10161), .QN(n16707) );
  NOR2X0 U17425 ( .IN1(g5990), .IN2(n10122), .QN(n12694) );
  NAND2X0 U17426 ( .IN1(test_so50), .IN2(n15690), .QN(n16706) );
  INVX0 U17427 ( .INP(n11711), .ZN(n15690) );
  NAND2X0 U17428 ( .IN1(test_so57), .IN2(g5990), .QN(n11711) );
  NAND2X0 U17429 ( .IN1(n16708), .IN2(n16709), .QN(n16704) );
  OR2X1 U17430 ( .IN1(n12691), .IN2(n9900), .Q(n16709) );
  NAND2X0 U17431 ( .IN1(n10122), .IN2(g5990), .QN(n12691) );
  NAND2X0 U17432 ( .IN1(n9900), .IN2(n16438), .QN(n16708) );
  INVX0 U17433 ( .INP(n16485), .ZN(n16438) );
  NAND2X0 U17434 ( .IN1(n5589), .IN2(n10122), .QN(n16485) );
  OR2X1 U17435 ( .IN1(n12700), .IN2(n5775), .Q(n16698) );
  NAND2X0 U17436 ( .IN1(n12693), .IN2(n10390), .QN(n12700) );
  INVX0 U17437 ( .INP(n12695), .ZN(n12693) );
  NOR2X0 U17438 ( .IN1(n10040), .IN2(n16710), .QN(n12695) );
  AND2X1 U17439 ( .IN1(n12643), .IN2(n16696), .Q(n16710) );
  NOR2X0 U17440 ( .IN1(n5877), .IN2(n10713), .QN(n12643) );
  OR2X1 U17441 ( .IN1(g4785), .IN2(n5518), .Q(n10713) );
  NAND2X0 U17442 ( .IN1(n16711), .IN2(n16712), .QN(g28084) );
  NAND2X0 U17443 ( .IN1(n16713), .IN2(n11814), .QN(n16712) );
  NOR2X0 U17444 ( .IN1(n10699), .IN2(n10710), .QN(n11814) );
  NOR2X0 U17445 ( .IN1(n10480), .IN2(n16714), .QN(n16713) );
  NOR2X0 U17446 ( .IN1(n16715), .IN2(test_so18), .QN(n16714) );
  NOR2X0 U17447 ( .IN1(n16716), .IN2(n12715), .QN(n16715) );
  INVX0 U17448 ( .INP(n12717), .ZN(n12715) );
  NOR2X0 U17449 ( .IN1(n16717), .IN2(n16718), .QN(n16716) );
  NAND2X0 U17450 ( .IN1(n16719), .IN2(n16720), .QN(n16718) );
  NAND2X0 U17451 ( .IN1(n15730), .IN2(g5698), .QN(n16720) );
  INVX0 U17452 ( .INP(n11704), .ZN(n15730) );
  NAND2X0 U17453 ( .IN1(g5644), .IN2(g5703), .QN(n11704) );
  NAND2X0 U17454 ( .IN1(n9903), .IN2(n12716), .QN(n16719) );
  NOR2X0 U17455 ( .IN1(g5644), .IN2(n5397), .QN(n12716) );
  NAND2X0 U17456 ( .IN1(n16721), .IN2(n16722), .QN(n16717) );
  OR2X1 U17457 ( .IN1(n12713), .IN2(n9904), .Q(n16722) );
  NAND2X0 U17458 ( .IN1(n5397), .IN2(g5644), .QN(n12713) );
  NAND2X0 U17459 ( .IN1(n9904), .IN2(n16504), .QN(n16721) );
  INVX0 U17460 ( .INP(n16551), .ZN(n16504) );
  NAND2X0 U17461 ( .IN1(n5593), .IN2(n5397), .QN(n16551) );
  NAND2X0 U17462 ( .IN1(n12720), .IN2(test_so18), .QN(n16711) );
  NOR2X0 U17463 ( .IN1(n12717), .IN2(n10458), .QN(n12720) );
  NOR2X0 U17464 ( .IN1(n5440), .IN2(n16723), .QN(n12717) );
  AND2X1 U17465 ( .IN1(n12644), .IN2(n16696), .Q(n16723) );
  NOR2X0 U17466 ( .IN1(n5876), .IN2(n10714), .QN(n12644) );
  NAND2X0 U17467 ( .IN1(n5518), .IN2(g4785), .QN(n10714) );
  NAND2X0 U17468 ( .IN1(n16724), .IN2(n16725), .QN(g28083) );
  NAND2X0 U17469 ( .IN1(n16726), .IN2(n11821), .QN(n16725) );
  NOR2X0 U17470 ( .IN1(n10699), .IN2(n16697), .QN(n11821) );
  INVX0 U17471 ( .INP(n10709), .ZN(n16697) );
  NOR2X0 U17472 ( .IN1(n5518), .IN2(n5361), .QN(n10709) );
  NAND2X0 U17473 ( .IN1(n16727), .IN2(g4793), .QN(n10699) );
  NOR2X0 U17474 ( .IN1(test_so29), .IN2(n5707), .QN(n16727) );
  NOR2X0 U17475 ( .IN1(n10480), .IN2(n16728), .QN(n16726) );
  NOR2X0 U17476 ( .IN1(n4708), .IN2(g4704), .QN(n16728) );
  NAND2X0 U17477 ( .IN1(n12737), .IN2(g4704), .QN(n16724) );
  NOR2X0 U17478 ( .IN1(g33959), .IN2(n10458), .QN(n12737) );
  INVX0 U17479 ( .INP(n10108), .ZN(g33959) );
  NAND2X0 U17480 ( .IN1(g4646), .IN2(n16729), .QN(n10108) );
  NAND2X0 U17481 ( .IN1(n12646), .IN2(n16696), .QN(n16729) );
  AND2X1 U17482 ( .IN1(n16730), .IN2(n16731), .Q(n16696) );
  NOR2X0 U17483 ( .IN1(n5707), .IN2(n16732), .QN(n16731) );
  NAND2X0 U17484 ( .IN1(g4669), .IN2(n10125), .QN(n16732) );
  NOR2X0 U17485 ( .IN1(n10133), .IN2(n16733), .QN(n16730) );
  NAND2X0 U17486 ( .IN1(n5368), .IN2(g4659), .QN(n16733) );
  NOR2X0 U17487 ( .IN1(n5862), .IN2(n10710), .QN(n12646) );
  NAND2X0 U17488 ( .IN1(n5518), .IN2(n5361), .QN(n10710) );
  NAND2X0 U17489 ( .IN1(n16734), .IN2(n16735), .QN(g28082) );
  NAND2X0 U17490 ( .IN1(n16736), .IN2(g4521), .QN(n16735) );
  NAND2X0 U17491 ( .IN1(n16737), .IN2(n10390), .QN(n16736) );
  NAND2X0 U17492 ( .IN1(n16738), .IN2(n5752), .QN(n16734) );
  AND2X1 U17493 ( .IN1(n10367), .IN2(n11172), .Q(n16738) );
  NAND2X0 U17494 ( .IN1(n16739), .IN2(n16740), .QN(g28074) );
  NAND2X0 U17495 ( .IN1(n10511), .IN2(g4119), .QN(n16740) );
  NOR2X0 U17496 ( .IN1(n16741), .IN2(n16742), .QN(n16739) );
  AND2X1 U17497 ( .IN1(n4721), .IN2(n4714), .Q(n16742) );
  NOR2X0 U17498 ( .IN1(n4714), .IN2(n16743), .QN(n16741) );
  NAND2X0 U17499 ( .IN1(n10370), .IN2(g4122), .QN(n16743) );
  NAND2X0 U17500 ( .IN1(n16744), .IN2(n16745), .QN(g28073) );
  NAND2X0 U17501 ( .IN1(n16746), .IN2(n4721), .QN(n16745) );
  INVX0 U17502 ( .INP(n16747), .ZN(n16746) );
  NOR2X0 U17503 ( .IN1(n16748), .IN2(n16749), .QN(n16744) );
  NOR2X0 U17504 ( .IN1(n9589), .IN2(n10354), .QN(n16749) );
  NOR2X0 U17505 ( .IN1(n10480), .IN2(n16750), .QN(n16748) );
  NAND2X0 U17506 ( .IN1(n16747), .IN2(g4119), .QN(n16750) );
  NAND2X0 U17507 ( .IN1(n16751), .IN2(g4057), .QN(n16747) );
  NAND2X0 U17508 ( .IN1(n16752), .IN2(n16753), .QN(g28072) );
  NAND2X0 U17509 ( .IN1(n16754), .IN2(n4721), .QN(n16753) );
  NOR2X0 U17510 ( .IN1(n16755), .IN2(n16756), .QN(n16752) );
  NOR2X0 U17511 ( .IN1(n10035), .IN2(n10352), .QN(n16756) );
  NOR2X0 U17512 ( .IN1(n10480), .IN2(n16757), .QN(n16755) );
  OR2X1 U17513 ( .IN1(n16754), .IN2(n9589), .Q(n16757) );
  AND2X1 U17514 ( .IN1(n16758), .IN2(n4722), .Q(n16754) );
  NOR2X0 U17515 ( .IN1(n5416), .IN2(g4057), .QN(n16758) );
  NAND2X0 U17516 ( .IN1(n16759), .IN2(n16760), .QN(g28071) );
  NAND2X0 U17517 ( .IN1(n16761), .IN2(g4112), .QN(n16760) );
  OR2X1 U17518 ( .IN1(n16761), .IN2(n10072), .Q(n16759) );
  AND2X1 U17519 ( .IN1(n16762), .IN2(n10365), .Q(n16761) );
  NAND2X0 U17520 ( .IN1(n16751), .IN2(n5711), .QN(n16762) );
  AND2X1 U17521 ( .IN1(n4722), .IN2(n5416), .Q(n16751) );
  AND2X1 U17522 ( .IN1(n16763), .IN2(n16764), .Q(n4722) );
  NOR2X0 U17523 ( .IN1(g4098), .IN2(n16765), .QN(n16764) );
  OR2X1 U17524 ( .IN1(n12618), .IN2(test_so11), .Q(n16765) );
  NAND2X0 U17525 ( .IN1(n5480), .IN2(n5340), .QN(n12618) );
  AND2X1 U17526 ( .IN1(n5612), .IN2(n9739), .Q(n16763) );
  NAND2X0 U17527 ( .IN1(n16766), .IN2(n16767), .QN(g28070) );
  NOR2X0 U17528 ( .IN1(n16768), .IN2(n16769), .QN(n16767) );
  NOR2X0 U17529 ( .IN1(n9739), .IN2(n10354), .QN(n16769) );
  NOR2X0 U17530 ( .IN1(n10480), .IN2(n16770), .QN(n16768) );
  NAND2X0 U17531 ( .IN1(test_so11), .IN2(n16771), .QN(n16770) );
  NOR2X0 U17532 ( .IN1(n10114), .IN2(n16772), .QN(n16766) );
  NOR2X0 U17533 ( .IN1(test_so11), .IN2(n16771), .QN(n16772) );
  INVX0 U17534 ( .INP(n15775), .ZN(n16771) );
  NOR2X0 U17535 ( .IN1(n16773), .IN2(n9739), .QN(n15775) );
  NAND2X0 U17536 ( .IN1(n16774), .IN2(n16775), .QN(g28069) );
  NAND2X0 U17537 ( .IN1(n12771), .IN2(g4035), .QN(n16775) );
  NOR2X0 U17538 ( .IN1(n12768), .IN2(n10457), .QN(n12771) );
  NOR2X0 U17539 ( .IN1(n16776), .IN2(n16777), .QN(n16774) );
  NOR2X0 U17540 ( .IN1(n10480), .IN2(n16778), .QN(n16777) );
  NAND2X0 U17541 ( .IN1(n12768), .IN2(n15813), .QN(n16778) );
  NAND2X0 U17542 ( .IN1(n16779), .IN2(n16780), .QN(n15813) );
  NOR2X0 U17543 ( .IN1(n16781), .IN2(n16782), .QN(n16780) );
  NOR2X0 U17544 ( .IN1(n5530), .IN2(n16783), .QN(n16782) );
  NOR2X0 U17545 ( .IN1(n16784), .IN2(n16785), .QN(n16783) );
  NAND2X0 U17546 ( .IN1(n16786), .IN2(n16787), .QN(n16785) );
  NAND2X0 U17547 ( .IN1(n16648), .IN2(n16788), .QN(n16787) );
  NAND2X0 U17548 ( .IN1(n16789), .IN2(n16790), .QN(n16788) );
  NAND2X0 U17549 ( .IN1(g4031), .IN2(g3897), .QN(n16790) );
  NAND2X0 U17550 ( .IN1(test_so24), .IN2(g14518), .QN(n16789) );
  NAND2X0 U17551 ( .IN1(n12767), .IN2(n16791), .QN(n16786) );
  NAND2X0 U17552 ( .IN1(n16792), .IN2(n16793), .QN(n16791) );
  NAND2X0 U17553 ( .IN1(g11418), .IN2(g3893), .QN(n16793) );
  NAND2X0 U17554 ( .IN1(g3917), .IN2(g16955), .QN(n16792) );
  NAND2X0 U17555 ( .IN1(n16794), .IN2(n16795), .QN(n16784) );
  NAND2X0 U17556 ( .IN1(n16796), .IN2(n16797), .QN(n16795) );
  NOR2X0 U17557 ( .IN1(n9946), .IN2(n5583), .QN(n16796) );
  NAND2X0 U17558 ( .IN1(n15815), .IN2(n16798), .QN(n16794) );
  NAND2X0 U17559 ( .IN1(n16799), .IN2(n16800), .QN(n16798) );
  OR2X1 U17560 ( .IN1(n9816), .IN2(n9990), .Q(n16800) );
  NAND2X0 U17561 ( .IN1(test_so65), .IN2(g16748), .QN(n16799) );
  NOR2X0 U17562 ( .IN1(n16801), .IN2(g4040), .QN(n16781) );
  NOR2X0 U17563 ( .IN1(n16802), .IN2(n16803), .QN(n16801) );
  NAND2X0 U17564 ( .IN1(n16804), .IN2(n16805), .QN(n16803) );
  NAND2X0 U17565 ( .IN1(n12767), .IN2(n16806), .QN(n16805) );
  NAND2X0 U17566 ( .IN1(n16807), .IN2(n16808), .QN(n16806) );
  NAND2X0 U17567 ( .IN1(g16748), .IN2(g3957), .QN(n16808) );
  OR2X1 U17568 ( .IN1(n9990), .IN2(n9991), .Q(n16807) );
  NAND2X0 U17569 ( .IN1(n16797), .IN2(n16809), .QN(n16804) );
  NAND2X0 U17570 ( .IN1(n16810), .IN2(n16811), .QN(n16809) );
  NAND2X0 U17571 ( .IN1(g4031), .IN2(g3913), .QN(n16811) );
  NAND2X0 U17572 ( .IN1(g14518), .IN2(g3901), .QN(n16810) );
  NAND2X0 U17573 ( .IN1(n16812), .IN2(n16813), .QN(n16802) );
  NAND2X0 U17574 ( .IN1(n16814), .IN2(n16648), .QN(n16813) );
  NOR2X0 U17575 ( .IN1(n9987), .IN2(n5583), .QN(n16814) );
  NAND2X0 U17576 ( .IN1(n15815), .IN2(n16815), .QN(n16812) );
  NAND2X0 U17577 ( .IN1(n16816), .IN2(n16817), .QN(n16815) );
  NAND2X0 U17578 ( .IN1(g11418), .IN2(g3909), .QN(n16817) );
  NAND2X0 U17579 ( .IN1(g16955), .IN2(g3925), .QN(n16816) );
  NOR2X0 U17580 ( .IN1(n16818), .IN2(n16819), .QN(n16779) );
  NOR2X0 U17581 ( .IN1(n16820), .IN2(n16821), .QN(n16819) );
  NOR2X0 U17582 ( .IN1(n16822), .IN2(n16823), .QN(n16820) );
  NAND2X0 U17583 ( .IN1(n16824), .IN2(n16825), .QN(n16823) );
  NAND2X0 U17584 ( .IN1(n16826), .IN2(n16797), .QN(n16825) );
  INVX0 U17585 ( .INP(n12764), .ZN(n16797) );
  NOR2X0 U17586 ( .IN1(n9839), .IN2(n5701), .QN(n16826) );
  NAND2X0 U17587 ( .IN1(n16827), .IN2(n15815), .QN(n16824) );
  INVX0 U17588 ( .INP(n11714), .ZN(n15815) );
  NAND2X0 U17589 ( .IN1(g3990), .IN2(g4054), .QN(n11714) );
  NOR2X0 U17590 ( .IN1(n9889), .IN2(n9888), .QN(n16827) );
  NOR2X0 U17591 ( .IN1(n16828), .IN2(n16829), .QN(n16822) );
  NAND2X0 U17592 ( .IN1(g16659), .IN2(g3953), .QN(n16829) );
  NOR2X0 U17593 ( .IN1(n16830), .IN2(n16831), .QN(n16818) );
  INVX0 U17594 ( .INP(n16821), .ZN(n16831) );
  XNOR2X1 U17595 ( .IN1(g11418), .IN2(n5530), .Q(n16821) );
  NOR2X0 U17596 ( .IN1(n16832), .IN2(n16833), .QN(n16830) );
  NAND2X0 U17597 ( .IN1(n16834), .IN2(n16835), .QN(n16833) );
  NAND2X0 U17598 ( .IN1(n16836), .IN2(n16648), .QN(n16835) );
  INVX0 U17599 ( .INP(n16828), .ZN(n16648) );
  NAND2X0 U17600 ( .IN1(n5594), .IN2(n5395), .QN(n16828) );
  NOR2X0 U17601 ( .IN1(n9856), .IN2(n5701), .QN(n16836) );
  NAND2X0 U17602 ( .IN1(n16837), .IN2(n12767), .QN(n16834) );
  NOR2X0 U17603 ( .IN1(g3990), .IN2(n5395), .QN(n12767) );
  NOR2X0 U17604 ( .IN1(n9888), .IN2(n9855), .QN(n16837) );
  NOR2X0 U17605 ( .IN1(n12764), .IN2(n16838), .QN(n16832) );
  NAND2X0 U17606 ( .IN1(g3961), .IN2(g16659), .QN(n16838) );
  NAND2X0 U17607 ( .IN1(n5395), .IN2(g3990), .QN(n12764) );
  INVX0 U17608 ( .INP(n12766), .ZN(n12768) );
  NAND2X0 U17609 ( .IN1(g4878), .IN2(n16839), .QN(n12766) );
  NAND2X0 U17610 ( .IN1(n12603), .IN2(n16682), .QN(n16839) );
  NOR2X0 U17611 ( .IN1(n5614), .IN2(n10746), .QN(n12603) );
  NAND2X0 U17612 ( .IN1(g4899), .IN2(g4975), .QN(n10746) );
  NOR2X0 U17613 ( .IN1(n9816), .IN2(n10353), .QN(n16776) );
  NAND2X0 U17614 ( .IN1(n16840), .IN2(n16841), .QN(g28066) );
  NAND2X0 U17615 ( .IN1(n12791), .IN2(g3684), .QN(n16841) );
  NOR2X0 U17616 ( .IN1(n12788), .IN2(n10457), .QN(n12791) );
  NOR2X0 U17617 ( .IN1(n16842), .IN2(n16843), .QN(n16840) );
  NOR2X0 U17618 ( .IN1(n10480), .IN2(n16844), .QN(n16843) );
  NAND2X0 U17619 ( .IN1(n12788), .IN2(n15852), .QN(n16844) );
  NAND2X0 U17620 ( .IN1(n16845), .IN2(n16846), .QN(n15852) );
  NOR2X0 U17621 ( .IN1(n16847), .IN2(n16848), .QN(n16846) );
  NOR2X0 U17622 ( .IN1(n5532), .IN2(n16849), .QN(n16848) );
  NOR2X0 U17623 ( .IN1(n16850), .IN2(n16851), .QN(n16849) );
  NAND2X0 U17624 ( .IN1(n16852), .IN2(n16853), .QN(n16851) );
  NAND2X0 U17625 ( .IN1(n16661), .IN2(n16854), .QN(n16853) );
  NAND2X0 U17626 ( .IN1(n16855), .IN2(n16856), .QN(n16854) );
  NAND2X0 U17627 ( .IN1(g3680), .IN2(g3546), .QN(n16856) );
  NAND2X0 U17628 ( .IN1(g14451), .IN2(g3538), .QN(n16855) );
  NAND2X0 U17629 ( .IN1(n12787), .IN2(n16857), .QN(n16852) );
  NAND2X0 U17630 ( .IN1(n16858), .IN2(n16859), .QN(n16857) );
  NAND2X0 U17631 ( .IN1(g11388), .IN2(g3542), .QN(n16859) );
  NAND2X0 U17632 ( .IN1(g3566), .IN2(g16924), .QN(n16858) );
  NAND2X0 U17633 ( .IN1(n16860), .IN2(n16861), .QN(n16850) );
  NAND2X0 U17634 ( .IN1(n16862), .IN2(test_so26), .QN(n16861) );
  NOR2X0 U17635 ( .IN1(n9948), .IN2(n12784), .QN(n16862) );
  NAND2X0 U17636 ( .IN1(n15855), .IN2(n16863), .QN(n16860) );
  NAND2X0 U17637 ( .IN1(n16864), .IN2(n16865), .QN(n16863) );
  OR2X1 U17638 ( .IN1(n10000), .IN2(n9802), .Q(n16865) );
  NAND2X0 U17639 ( .IN1(g3598), .IN2(g16722), .QN(n16864) );
  NOR2X0 U17640 ( .IN1(n16866), .IN2(g3689), .QN(n16847) );
  NOR2X0 U17641 ( .IN1(n16867), .IN2(n16868), .QN(n16866) );
  NAND2X0 U17642 ( .IN1(n16869), .IN2(n16870), .QN(n16868) );
  NAND2X0 U17643 ( .IN1(n12787), .IN2(n16871), .QN(n16870) );
  NAND2X0 U17644 ( .IN1(n16872), .IN2(n16873), .QN(n16871) );
  NAND2X0 U17645 ( .IN1(g16656), .IN2(g3554), .QN(n16873) );
  NAND2X0 U17646 ( .IN1(g16722), .IN2(g3606), .QN(n16872) );
  NAND2X0 U17647 ( .IN1(n16874), .IN2(n16875), .QN(n16869) );
  NAND2X0 U17648 ( .IN1(n16876), .IN2(n16877), .QN(n16875) );
  NAND2X0 U17649 ( .IN1(g3680), .IN2(g3562), .QN(n16877) );
  NAND2X0 U17650 ( .IN1(g14451), .IN2(g3550), .QN(n16876) );
  NAND2X0 U17651 ( .IN1(n16878), .IN2(n16879), .QN(n16867) );
  NAND2X0 U17652 ( .IN1(n16880), .IN2(n16661), .QN(n16879) );
  AND2X1 U17653 ( .IN1(g3590), .IN2(test_so26), .Q(n16880) );
  NAND2X0 U17654 ( .IN1(n15855), .IN2(n16881), .QN(n16878) );
  NAND2X0 U17655 ( .IN1(n16882), .IN2(n16883), .QN(n16881) );
  NAND2X0 U17656 ( .IN1(g11388), .IN2(g3558), .QN(n16883) );
  NAND2X0 U17657 ( .IN1(g16924), .IN2(g3574), .QN(n16882) );
  NOR2X0 U17658 ( .IN1(n16884), .IN2(n16885), .QN(n16845) );
  NOR2X0 U17659 ( .IN1(n16886), .IN2(n16887), .QN(n16885) );
  NOR2X0 U17660 ( .IN1(n16888), .IN2(n16889), .QN(n16886) );
  NAND2X0 U17661 ( .IN1(n16890), .IN2(n16891), .QN(n16889) );
  NAND2X0 U17662 ( .IN1(n16892), .IN2(n16874), .QN(n16891) );
  INVX0 U17663 ( .INP(n12784), .ZN(n16874) );
  NOR2X0 U17664 ( .IN1(n9841), .IN2(n5699), .QN(n16892) );
  NAND2X0 U17665 ( .IN1(n16893), .IN2(n15855), .QN(n16890) );
  INVX0 U17666 ( .INP(n11710), .ZN(n15855) );
  NAND2X0 U17667 ( .IN1(g3639), .IN2(g3703), .QN(n11710) );
  NOR2X0 U17668 ( .IN1(n9893), .IN2(n9892), .QN(n16893) );
  NOR2X0 U17669 ( .IN1(n16894), .IN2(n16895), .QN(n16888) );
  NAND2X0 U17670 ( .IN1(test_so43), .IN2(g16627), .QN(n16895) );
  NOR2X0 U17671 ( .IN1(n16896), .IN2(n16897), .QN(n16884) );
  INVX0 U17672 ( .INP(n16887), .ZN(n16897) );
  XNOR2X1 U17673 ( .IN1(g11388), .IN2(n5532), .Q(n16887) );
  NOR2X0 U17674 ( .IN1(n16898), .IN2(n16899), .QN(n16896) );
  NAND2X0 U17675 ( .IN1(n16900), .IN2(n16901), .QN(n16899) );
  NAND2X0 U17676 ( .IN1(n16902), .IN2(n16661), .QN(n16901) );
  INVX0 U17677 ( .INP(n16894), .ZN(n16661) );
  NAND2X0 U17678 ( .IN1(n5591), .IN2(n5399), .QN(n16894) );
  NOR2X0 U17679 ( .IN1(n9862), .IN2(n5699), .QN(n16902) );
  NAND2X0 U17680 ( .IN1(n16903), .IN2(n12787), .QN(n16900) );
  NOR2X0 U17681 ( .IN1(g3639), .IN2(n5399), .QN(n12787) );
  NOR2X0 U17682 ( .IN1(n9892), .IN2(n9861), .QN(n16903) );
  NOR2X0 U17683 ( .IN1(n12784), .IN2(n16904), .QN(n16898) );
  NAND2X0 U17684 ( .IN1(g3610), .IN2(g16627), .QN(n16904) );
  NAND2X0 U17685 ( .IN1(n5399), .IN2(g3639), .QN(n12784) );
  INVX0 U17686 ( .INP(n12786), .ZN(n12788) );
  NAND2X0 U17687 ( .IN1(g4871), .IN2(n16905), .QN(n12786) );
  NAND2X0 U17688 ( .IN1(n12604), .IN2(n16682), .QN(n16905) );
  NOR2X0 U17689 ( .IN1(n5875), .IN2(n10744), .QN(n12604) );
  NAND2X0 U17690 ( .IN1(n5360), .IN2(g4899), .QN(n10744) );
  NOR2X0 U17691 ( .IN1(n9802), .IN2(n10352), .QN(n16842) );
  NAND2X0 U17692 ( .IN1(n16906), .IN2(n16907), .QN(g28063) );
  NAND2X0 U17693 ( .IN1(n12811), .IN2(g3333), .QN(n16907) );
  NOR2X0 U17694 ( .IN1(n12808), .IN2(n10457), .QN(n12811) );
  NOR2X0 U17695 ( .IN1(n16908), .IN2(n16909), .QN(n16906) );
  NOR2X0 U17696 ( .IN1(n10480), .IN2(n16910), .QN(n16909) );
  NAND2X0 U17697 ( .IN1(n12808), .IN2(n15893), .QN(n16910) );
  NAND2X0 U17698 ( .IN1(n16911), .IN2(n16912), .QN(n15893) );
  NOR2X0 U17699 ( .IN1(n16913), .IN2(n16914), .QN(n16912) );
  NOR2X0 U17700 ( .IN1(n5527), .IN2(n16915), .QN(n16914) );
  NOR2X0 U17701 ( .IN1(n16916), .IN2(n16917), .QN(n16915) );
  NAND2X0 U17702 ( .IN1(n16918), .IN2(n16919), .QN(n16917) );
  NAND2X0 U17703 ( .IN1(n16675), .IN2(n16920), .QN(n16919) );
  NAND2X0 U17704 ( .IN1(n16921), .IN2(n16922), .QN(n16920) );
  NAND2X0 U17705 ( .IN1(g14421), .IN2(g3187), .QN(n16922) );
  NAND2X0 U17706 ( .IN1(test_so91), .IN2(test_so88), .QN(n16921) );
  NAND2X0 U17707 ( .IN1(n12807), .IN2(n16923), .QN(n16918) );
  NAND2X0 U17708 ( .IN1(n16924), .IN2(n16925), .QN(n16923) );
  NAND2X0 U17709 ( .IN1(g11349), .IN2(g3191), .QN(n16925) );
  NAND2X0 U17710 ( .IN1(g3215), .IN2(g16874), .QN(n16924) );
  NAND2X0 U17711 ( .IN1(n16926), .IN2(n16927), .QN(n16916) );
  NAND2X0 U17712 ( .IN1(n16928), .IN2(n12802), .QN(n16927) );
  NOR2X0 U17713 ( .IN1(n9942), .IN2(n5580), .QN(n16928) );
  NAND2X0 U17714 ( .IN1(n15895), .IN2(n16929), .QN(n16926) );
  NAND2X0 U17715 ( .IN1(n16930), .IN2(n16931), .QN(n16929) );
  OR2X1 U17716 ( .IN1(n9791), .IN2(n9971), .Q(n16931) );
  NAND2X0 U17717 ( .IN1(g3247), .IN2(g16686), .QN(n16930) );
  NOR2X0 U17718 ( .IN1(n16932), .IN2(g3338), .QN(n16913) );
  NOR2X0 U17719 ( .IN1(n16933), .IN2(n16934), .QN(n16932) );
  NAND2X0 U17720 ( .IN1(n16935), .IN2(n16936), .QN(n16934) );
  NAND2X0 U17721 ( .IN1(n12807), .IN2(n16937), .QN(n16936) );
  NAND2X0 U17722 ( .IN1(n16938), .IN2(n16939), .QN(n16937) );
  NAND2X0 U17723 ( .IN1(g16686), .IN2(g3255), .QN(n16939) );
  OR2X1 U17724 ( .IN1(n9971), .IN2(n9972), .Q(n16938) );
  NAND2X0 U17725 ( .IN1(n12802), .IN2(n16940), .QN(n16935) );
  NAND2X0 U17726 ( .IN1(n16941), .IN2(n16942), .QN(n16940) );
  NAND2X0 U17727 ( .IN1(test_so91), .IN2(g3211), .QN(n16942) );
  NAND2X0 U17728 ( .IN1(g14421), .IN2(g3199), .QN(n16941) );
  NAND2X0 U17729 ( .IN1(n16943), .IN2(n16944), .QN(n16933) );
  NAND2X0 U17730 ( .IN1(n16945), .IN2(n16675), .QN(n16944) );
  NOR2X0 U17731 ( .IN1(n9968), .IN2(n5580), .QN(n16945) );
  NAND2X0 U17732 ( .IN1(n15895), .IN2(n16946), .QN(n16943) );
  NAND2X0 U17733 ( .IN1(n16947), .IN2(n16948), .QN(n16946) );
  NAND2X0 U17734 ( .IN1(g11349), .IN2(g3207), .QN(n16948) );
  NAND2X0 U17735 ( .IN1(g16874), .IN2(g3223), .QN(n16947) );
  NOR2X0 U17736 ( .IN1(n16949), .IN2(n16950), .QN(n16911) );
  NOR2X0 U17737 ( .IN1(n16951), .IN2(n16952), .QN(n16950) );
  NOR2X0 U17738 ( .IN1(n16953), .IN2(n16954), .QN(n16951) );
  NAND2X0 U17739 ( .IN1(n16955), .IN2(n16956), .QN(n16954) );
  NAND2X0 U17740 ( .IN1(n16957), .IN2(n12802), .QN(n16956) );
  INVX0 U17741 ( .INP(n16674), .ZN(n12802) );
  NOR2X0 U17742 ( .IN1(n9836), .IN2(n5702), .QN(n16957) );
  NAND2X0 U17743 ( .IN1(n16958), .IN2(n15895), .QN(n16955) );
  INVX0 U17744 ( .INP(n11702), .ZN(n15895) );
  NAND2X0 U17745 ( .IN1(g3352), .IN2(g3288), .QN(n11702) );
  NOR2X0 U17746 ( .IN1(n9882), .IN2(n9881), .QN(n16958) );
  NOR2X0 U17747 ( .IN1(n16959), .IN2(n16960), .QN(n16953) );
  NAND2X0 U17748 ( .IN1(g16603), .IN2(g3251), .QN(n16960) );
  NOR2X0 U17749 ( .IN1(n16961), .IN2(n16962), .QN(n16949) );
  INVX0 U17750 ( .INP(n16952), .ZN(n16962) );
  XNOR2X1 U17751 ( .IN1(g11349), .IN2(n5527), .Q(n16952) );
  NOR2X0 U17752 ( .IN1(n16963), .IN2(n16964), .QN(n16961) );
  NAND2X0 U17753 ( .IN1(n16965), .IN2(n16966), .QN(n16964) );
  NAND2X0 U17754 ( .IN1(n16967), .IN2(n16675), .QN(n16966) );
  INVX0 U17755 ( .INP(n16959), .ZN(n16675) );
  NAND2X0 U17756 ( .IN1(n5400), .IN2(n5604), .QN(n16959) );
  NOR2X0 U17757 ( .IN1(n9844), .IN2(n5702), .QN(n16967) );
  NAND2X0 U17758 ( .IN1(n16968), .IN2(n12807), .QN(n16965) );
  NOR2X0 U17759 ( .IN1(g3288), .IN2(n5604), .QN(n12807) );
  NOR2X0 U17760 ( .IN1(n9881), .IN2(n9843), .QN(n16968) );
  NOR2X0 U17761 ( .IN1(n16674), .IN2(n16969), .QN(n16963) );
  NAND2X0 U17762 ( .IN1(test_so84), .IN2(g16603), .QN(n16969) );
  NAND2X0 U17763 ( .IN1(n5604), .IN2(g3288), .QN(n16674) );
  INVX0 U17764 ( .INP(n12806), .ZN(n12808) );
  NAND2X0 U17765 ( .IN1(g4864), .IN2(n16970), .QN(n12806) );
  NAND2X0 U17766 ( .IN1(n12605), .IN2(n16682), .QN(n16970) );
  AND2X1 U17767 ( .IN1(n16971), .IN2(n16972), .Q(n16682) );
  NOR2X0 U17768 ( .IN1(n9586), .IN2(n16973), .QN(n16972) );
  NAND2X0 U17769 ( .IN1(g4843), .IN2(n10123), .QN(n16973) );
  NOR2X0 U17770 ( .IN1(g4983), .IN2(n16974), .QN(n16971) );
  NAND2X0 U17771 ( .IN1(g4849), .IN2(g4966), .QN(n16974) );
  NOR2X0 U17772 ( .IN1(n5878), .IN2(n10743), .QN(n12605) );
  NAND2X0 U17773 ( .IN1(n5517), .IN2(g4975), .QN(n10743) );
  NOR2X0 U17774 ( .IN1(n9791), .IN2(n10350), .QN(n16908) );
  NAND2X0 U17775 ( .IN1(n16975), .IN2(n16976), .QN(g28060) );
  NOR2X0 U17776 ( .IN1(n16977), .IN2(n16978), .QN(n16976) );
  NOR2X0 U17777 ( .IN1(n5301), .IN2(n10353), .QN(n16978) );
  NOR2X0 U17778 ( .IN1(n10480), .IN2(n16979), .QN(n16977) );
  NAND2X0 U17779 ( .IN1(n15903), .IN2(g2729), .QN(n16979) );
  NOR2X0 U17780 ( .IN1(n2787), .IN2(n16980), .QN(n16975) );
  NOR2X0 U17781 ( .IN1(g2729), .IN2(n15903), .QN(n16980) );
  NAND2X0 U17782 ( .IN1(n15161), .IN2(g2724), .QN(n15903) );
  INVX0 U17783 ( .INP(n13609), .ZN(n2787) );
  OR2X1 U17784 ( .IN1(n16981), .IN2(n16982), .Q(g28059) );
  NAND2X0 U17785 ( .IN1(n16983), .IN2(n16984), .QN(n16982) );
  NAND2X0 U17786 ( .IN1(n16985), .IN2(n15501), .QN(n16984) );
  AND2X1 U17787 ( .IN1(n9750), .IN2(n13906), .Q(n16985) );
  NOR2X0 U17788 ( .IN1(n13302), .IN2(n10458), .QN(n13906) );
  NAND2X0 U17789 ( .IN1(n16986), .IN2(n16987), .QN(n13302) );
  NOR2X0 U17790 ( .IN1(n16988), .IN2(n16989), .QN(n16987) );
  NOR2X0 U17791 ( .IN1(n16990), .IN2(n16991), .QN(n16989) );
  NAND2X0 U17792 ( .IN1(n16992), .IN2(g1351), .QN(n16991) );
  NOR2X0 U17793 ( .IN1(g1351), .IN2(n16993), .QN(n16988) );
  NOR2X0 U17794 ( .IN1(n16994), .IN2(g1312), .QN(n16986) );
  NAND2X0 U17795 ( .IN1(n4798), .IN2(n16995), .QN(n16983) );
  NOR2X0 U17796 ( .IN1(n5322), .IN2(n10351), .QN(n16981) );
  NAND2X0 U17797 ( .IN1(n16996), .IN2(n16997), .QN(g28058) );
  NAND2X0 U17798 ( .IN1(test_so77), .IN2(n10516), .QN(n16997) );
  NOR2X0 U17799 ( .IN1(n16998), .IN2(n16999), .QN(n16996) );
  NOR2X0 U17800 ( .IN1(g1252), .IN2(n17000), .QN(n16999) );
  NOR2X0 U17801 ( .IN1(n5554), .IN2(n17001), .QN(n16998) );
  NAND2X0 U17802 ( .IN1(n13309), .IN2(n17000), .QN(n17001) );
  INVX0 U17803 ( .INP(n4490), .ZN(n17000) );
  OR2X1 U17804 ( .IN1(n17002), .IN2(n17003), .Q(g28057) );
  NAND2X0 U17805 ( .IN1(n17004), .IN2(n17005), .QN(n17003) );
  NAND2X0 U17806 ( .IN1(n17006), .IN2(n15542), .QN(n17005) );
  AND2X1 U17807 ( .IN1(n9751), .IN2(n13922), .Q(n17006) );
  NOR2X0 U17808 ( .IN1(n13321), .IN2(n10459), .QN(n13922) );
  NAND2X0 U17809 ( .IN1(n17007), .IN2(n17008), .QN(n13321) );
  NOR2X0 U17810 ( .IN1(n17009), .IN2(n17010), .QN(n17008) );
  NOR2X0 U17811 ( .IN1(n17011), .IN2(g1008), .QN(n17010) );
  NOR2X0 U17812 ( .IN1(n17012), .IN2(n17013), .QN(n17009) );
  NOR2X0 U17813 ( .IN1(test_so20), .IN2(n17014), .QN(n17007) );
  NAND2X0 U17814 ( .IN1(n4805), .IN2(n17015), .QN(n17004) );
  NOR2X0 U17815 ( .IN1(n5321), .IN2(n10353), .QN(n17002) );
  NAND2X0 U17816 ( .IN1(n17016), .IN2(n17017), .QN(g28056) );
  NAND2X0 U17817 ( .IN1(n10510), .IN2(g936), .QN(n17017) );
  NOR2X0 U17818 ( .IN1(n17018), .IN2(n17019), .QN(n17016) );
  NOR2X0 U17819 ( .IN1(g907), .IN2(n17020), .QN(n17019) );
  NOR2X0 U17820 ( .IN1(n5555), .IN2(n17021), .QN(n17018) );
  NAND2X0 U17821 ( .IN1(n13328), .IN2(n17020), .QN(n17021) );
  INVX0 U17822 ( .INP(n4514), .ZN(n17020) );
  NAND2X0 U17823 ( .IN1(n17022), .IN2(n17023), .QN(g28055) );
  OR2X1 U17824 ( .IN1(n10309), .IN2(n5422), .Q(n17023) );
  NOR2X0 U17825 ( .IN1(n17024), .IN2(n17025), .QN(n17022) );
  NOR2X0 U17826 ( .IN1(g827), .IN2(n17026), .QN(n17025) );
  NAND2X0 U17827 ( .IN1(n4519), .IN2(n16231), .QN(n17026) );
  NOR2X0 U17828 ( .IN1(n5728), .IN2(n17027), .QN(n17024) );
  NAND2X0 U17829 ( .IN1(n42), .IN2(n17028), .QN(n17027) );
  INVX0 U17830 ( .INP(n4519), .ZN(n17028) );
  NAND2X0 U17831 ( .IN1(n17029), .IN2(n17030), .QN(g28054) );
  OR2X1 U17832 ( .IN1(n17031), .IN2(n9790), .Q(n17030) );
  NAND2X0 U17833 ( .IN1(n17031), .IN2(g661), .QN(n17029) );
  NAND2X0 U17834 ( .IN1(n17032), .IN2(n17033), .QN(g28053) );
  NAND2X0 U17835 ( .IN1(n10510), .IN2(g681), .QN(n17033) );
  NOR2X0 U17836 ( .IN1(n17034), .IN2(n17035), .QN(n17032) );
  NOR2X0 U17837 ( .IN1(n10145), .IN2(n17036), .QN(n17035) );
  NAND2X0 U17838 ( .IN1(n17037), .IN2(n17038), .QN(g28052) );
  NAND2X0 U17839 ( .IN1(n17039), .IN2(g661), .QN(n17038) );
  NAND2X0 U17840 ( .IN1(n17031), .IN2(g718), .QN(n17037) );
  NAND2X0 U17841 ( .IN1(n17040), .IN2(n17041), .QN(g28051) );
  NAND2X0 U17842 ( .IN1(n17039), .IN2(g718), .QN(n17041) );
  NAND2X0 U17843 ( .IN1(n17031), .IN2(g655), .QN(n17040) );
  NAND2X0 U17844 ( .IN1(n17042), .IN2(n17043), .QN(g28050) );
  NAND2X0 U17845 ( .IN1(n17039), .IN2(g655), .QN(n17043) );
  NAND2X0 U17846 ( .IN1(n17031), .IN2(g650), .QN(n17042) );
  NAND2X0 U17847 ( .IN1(n17044), .IN2(n17045), .QN(g28049) );
  NAND2X0 U17848 ( .IN1(test_so87), .IN2(n10515), .QN(n17045) );
  NOR2X0 U17849 ( .IN1(n17046), .IN2(n17047), .QN(n17044) );
  NOR2X0 U17850 ( .IN1(n9774), .IN2(n17031), .QN(n17047) );
  AND2X1 U17851 ( .IN1(g681), .IN2(n17034), .Q(n17046) );
  NAND2X0 U17852 ( .IN1(n17048), .IN2(n17049), .QN(g28048) );
  NAND2X0 U17853 ( .IN1(n10499), .IN2(g29212), .QN(n17049) );
  NOR2X0 U17854 ( .IN1(n17050), .IN2(n17051), .QN(n17048) );
  NOR2X0 U17855 ( .IN1(n4819), .IN2(n17052), .QN(n17051) );
  NAND2X0 U17856 ( .IN1(n17053), .IN2(n17054), .QN(n4819) );
  NOR2X0 U17857 ( .IN1(n5821), .IN2(n16256), .QN(n17054) );
  NAND2X0 U17858 ( .IN1(n17055), .IN2(n17056), .QN(n16256) );
  NOR2X0 U17859 ( .IN1(g645), .IN2(g650), .QN(n17056) );
  NOR2X0 U17860 ( .IN1(n10145), .IN2(n17057), .QN(n17055) );
  XOR2X1 U17861 ( .IN1(n9790), .IN2(n9789), .Q(n17057) );
  AND2X1 U17862 ( .IN1(n5520), .IN2(n5112), .Q(n17053) );
  NOR2X0 U17863 ( .IN1(n5520), .IN2(n17058), .QN(n17050) );
  NOR2X0 U17864 ( .IN1(n17059), .IN2(n17060), .QN(n17058) );
  NOR2X0 U17865 ( .IN1(n10479), .IN2(n17061), .QN(n17059) );
  OR2X1 U17866 ( .IN1(n5821), .IN2(test_so70), .Q(n17061) );
  NAND2X0 U17867 ( .IN1(n17062), .IN2(n17063), .QN(g28047) );
  NAND2X0 U17868 ( .IN1(n17039), .IN2(g681), .QN(n17063) );
  NAND2X0 U17869 ( .IN1(n17031), .IN2(g645), .QN(n17062) );
  NAND2X0 U17870 ( .IN1(n17064), .IN2(n17065), .QN(g28046) );
  NAND2X0 U17871 ( .IN1(n17034), .IN2(g446), .QN(n17065) );
  NOR2X0 U17872 ( .IN1(n17066), .IN2(n10458), .QN(n17034) );
  NAND2X0 U17873 ( .IN1(n17039), .IN2(g645), .QN(n17064) );
  INVX0 U17874 ( .INP(n17031), .ZN(n17039) );
  NAND2X0 U17875 ( .IN1(n17066), .IN2(n10390), .QN(n17031) );
  NAND2X0 U17876 ( .IN1(n17067), .IN2(n17068), .QN(n17066) );
  NOR2X0 U17877 ( .IN1(n17069), .IN2(n17070), .QN(n17068) );
  NOR2X0 U17878 ( .IN1(n17071), .IN2(g691), .QN(n17070) );
  NOR2X0 U17879 ( .IN1(g424), .IN2(n17072), .QN(n17071) );
  NAND2X0 U17880 ( .IN1(n5629), .IN2(g417), .QN(n17072) );
  AND2X1 U17881 ( .IN1(g691), .IN2(n17073), .Q(n17069) );
  NOR2X0 U17882 ( .IN1(n5121), .IN2(g370), .QN(n17067) );
  NAND2X0 U17883 ( .IN1(n17074), .IN2(n17075), .QN(g28045) );
  NAND2X0 U17884 ( .IN1(n10499), .IN2(g568), .QN(n17075) );
  NOR2X0 U17885 ( .IN1(n17076), .IN2(n17077), .QN(n17074) );
  NOR2X0 U17886 ( .IN1(g572), .IN2(n17078), .QN(n17077) );
  NOR2X0 U17887 ( .IN1(n5337), .IN2(n17079), .QN(n17076) );
  NAND2X0 U17888 ( .IN1(n2421), .IN2(n17078), .QN(n17079) );
  INVX0 U17889 ( .INP(n4537), .ZN(n17078) );
  NAND2X0 U17890 ( .IN1(n17080), .IN2(n17081), .QN(g28044) );
  NAND2X0 U17891 ( .IN1(n10499), .IN2(g528), .QN(n17081) );
  NAND2X0 U17892 ( .IN1(n17082), .IN2(n10389), .QN(n17080) );
  NAND2X0 U17893 ( .IN1(n17083), .IN2(n17084), .QN(n17082) );
  XNOR2X1 U17894 ( .IN1(n5820), .IN2(n16270), .Q(n17083) );
  NAND2X0 U17895 ( .IN1(n17085), .IN2(n17086), .QN(n16270) );
  NOR2X0 U17896 ( .IN1(n17087), .IN2(n17088), .QN(n17085) );
  AND2X1 U17897 ( .IN1(n17089), .IN2(n5327), .Q(n17087) );
  NAND2X0 U17898 ( .IN1(n17090), .IN2(n17091), .QN(g28043) );
  NAND2X0 U17899 ( .IN1(n10106), .IN2(n10154), .QN(n17091) );
  NOR2X0 U17900 ( .IN1(n13958), .IN2(n10458), .QN(n10106) );
  NAND2X0 U17901 ( .IN1(n17092), .IN2(n15566), .QN(n13958) );
  NOR2X0 U17902 ( .IN1(n16235), .IN2(n5520), .QN(n15566) );
  AND2X1 U17903 ( .IN1(n17093), .IN2(n17094), .Q(n16235) );
  NOR2X0 U17904 ( .IN1(n17095), .IN2(n17096), .QN(n17094) );
  NOR2X0 U17905 ( .IN1(g655), .IN2(n17097), .QN(n17096) );
  NAND2X0 U17906 ( .IN1(n9678), .IN2(n9819), .QN(n17097) );
  NOR2X0 U17907 ( .IN1(n9820), .IN2(n17098), .QN(n17095) );
  NAND2X0 U17908 ( .IN1(g753), .IN2(g718), .QN(n17098) );
  NOR2X0 U17909 ( .IN1(n17099), .IN2(n17100), .QN(n17093) );
  NOR2X0 U17910 ( .IN1(n9708), .IN2(n5479), .QN(n17099) );
  NOR2X0 U17911 ( .IN1(n17101), .IN2(n17102), .QN(n17092) );
  AND2X1 U17912 ( .IN1(g278), .IN2(n17103), .Q(n17102) );
  NAND2X0 U17913 ( .IN1(n10498), .IN2(g278), .QN(n17090) );
  NAND2X0 U17914 ( .IN1(n17104), .IN2(n5630), .QN(g28042) );
  NOR2X0 U17915 ( .IN1(n10479), .IN2(g1306), .QN(n17104) );
  NAND2X0 U17916 ( .IN1(n17105), .IN2(n11259), .QN(g28041) );
  NAND2X0 U17917 ( .IN1(g1536), .IN2(n4836), .QN(n11259) );
  NOR2X0 U17918 ( .IN1(n10479), .IN2(n11355), .QN(n17105) );
  INVX0 U17919 ( .INP(n11260), .ZN(n11355) );
  NAND2X0 U17920 ( .IN1(g1193), .IN2(n4837), .QN(n11260) );
  NAND2X0 U17921 ( .IN1(n17106), .IN2(n17107), .QN(g28030) );
  NAND2X0 U17922 ( .IN1(n17108), .IN2(n5882), .QN(n17107) );
  NOR2X0 U17923 ( .IN1(n17109), .IN2(g3129), .QN(n17108) );
  NOR2X0 U17924 ( .IN1(n17110), .IN2(n17111), .QN(n17109) );
  NOR2X0 U17925 ( .IN1(n17112), .IN2(n11288), .QN(n17111) );
  INVX0 U17926 ( .INP(n17113), .ZN(n11288) );
  NOR2X0 U17927 ( .IN1(n17114), .IN2(n17115), .QN(n17112) );
  NOR2X0 U17928 ( .IN1(n17116), .IN2(n17117), .QN(n17115) );
  NOR2X0 U17929 ( .IN1(n17118), .IN2(n17119), .QN(n17116) );
  NOR2X0 U17930 ( .IN1(n17120), .IN2(n17121), .QN(n17118) );
  NOR2X0 U17931 ( .IN1(n17122), .IN2(n17123), .QN(n17121) );
  NOR2X0 U17932 ( .IN1(n17124), .IN2(n17125), .QN(n17122) );
  NAND2X0 U17933 ( .IN1(n17126), .IN2(n17127), .QN(n17124) );
  NAND2X0 U17934 ( .IN1(n17128), .IN2(n17129), .QN(n17127) );
  OR2X1 U17935 ( .IN1(g5831), .IN2(test_so83), .Q(n17129) );
  NAND2X0 U17936 ( .IN1(n5888), .IN2(n5874), .QN(n17128) );
  NAND2X0 U17937 ( .IN1(n17130), .IN2(n17131), .QN(n17126) );
  INVX0 U17938 ( .INP(n17132), .ZN(n17120) );
  NAND2X0 U17939 ( .IN1(n17110), .IN2(n17113), .QN(n17106) );
  NAND2X0 U17940 ( .IN1(n17133), .IN2(n10389), .QN(n17113) );
  NAND2X0 U17941 ( .IN1(n5889), .IN2(n5868), .QN(n17133) );
  INVX0 U17942 ( .INP(n11289), .ZN(n17110) );
  NAND2X0 U17943 ( .IN1(n17114), .IN2(n17134), .QN(n11289) );
  NAND2X0 U17944 ( .IN1(n17117), .IN2(n10389), .QN(n17134) );
  NAND2X0 U17945 ( .IN1(n5886), .IN2(n5872), .QN(n17117) );
  AND2X1 U17946 ( .IN1(n17119), .IN2(n17132), .Q(n17114) );
  NAND2X0 U17947 ( .IN1(n17135), .IN2(n10389), .QN(n17132) );
  NAND2X0 U17948 ( .IN1(n5883), .IN2(n5871), .QN(n17135) );
  AND2X1 U17949 ( .IN1(n17123), .IN2(n17136), .Q(n17119) );
  NAND2X0 U17950 ( .IN1(n17125), .IN2(n10389), .QN(n17136) );
  NAND2X0 U17951 ( .IN1(n5885), .IN2(n5869), .QN(n17125) );
  NOR2X0 U17952 ( .IN1(n17130), .IN2(n17131), .QN(n17123) );
  AND2X1 U17953 ( .IN1(n17137), .IN2(n10365), .Q(n17131) );
  NAND2X0 U17954 ( .IN1(n17138), .IN2(n17139), .QN(n17137) );
  NOR2X0 U17955 ( .IN1(test_so83), .IN2(g5831), .QN(n17139) );
  NOR2X0 U17956 ( .IN1(g6177), .IN2(g6191), .QN(n17138) );
  AND2X1 U17957 ( .IN1(n17140), .IN2(n10365), .Q(n17130) );
  NAND2X0 U17958 ( .IN1(n5884), .IN2(n5870), .QN(n17140) );
  NAND2X0 U17959 ( .IN1(n17141), .IN2(n12753), .QN(g26971) );
  NAND2X0 U17960 ( .IN1(n5670), .IN2(n10389), .QN(n12753) );
  NOR2X0 U17961 ( .IN1(n17142), .IN2(n17143), .QN(n17141) );
  NOR2X0 U17962 ( .IN1(n9768), .IN2(n10348), .QN(n17143) );
  NOR2X0 U17963 ( .IN1(n10479), .IN2(g4531), .QN(n17142) );
  NAND2X0 U17964 ( .IN1(n17144), .IN2(n17145), .QN(g26970) );
  NAND2X0 U17965 ( .IN1(n10373), .IN2(g4473), .QN(n17145) );
  NAND2X0 U17966 ( .IN1(n10497), .IN2(g4459), .QN(n17144) );
  NAND2X0 U17967 ( .IN1(n17146), .IN2(n17147), .QN(g26969) );
  NAND2X0 U17968 ( .IN1(n10498), .IN2(g4462), .QN(n17147) );
  NAND2X0 U17969 ( .IN1(n17148), .IN2(n10389), .QN(n17146) );
  NOR2X0 U17970 ( .IN1(test_so38), .IN2(g4473), .QN(n17148) );
  NAND2X0 U17971 ( .IN1(n17149), .IN2(n17150), .QN(g26968) );
  NAND2X0 U17972 ( .IN1(n10497), .IN2(g4558), .QN(n17149) );
  NAND2X0 U17973 ( .IN1(n17151), .IN2(n17152), .QN(g26967) );
  NAND2X0 U17974 ( .IN1(n10497), .IN2(g4561), .QN(n17151) );
  NAND2X0 U17975 ( .IN1(n17153), .IN2(n17154), .QN(g26966) );
  NAND2X0 U17976 ( .IN1(n10497), .IN2(g4555), .QN(n17153) );
  XOR2X1 U17977 ( .IN1(DFF_228_n1), .IN2(n17155), .Q(g26965) );
  NAND2X0 U17978 ( .IN1(n10374), .IN2(g10306), .QN(n17155) );
  NAND2X0 U17979 ( .IN1(n17156), .IN2(n17157), .QN(g26964) );
  OR2X1 U17980 ( .IN1(n10310), .IN2(n10071), .Q(n17157) );
  NAND2X0 U17981 ( .IN1(n17158), .IN2(n10389), .QN(n17156) );
  NAND2X0 U17982 ( .IN1(n17159), .IN2(n17160), .QN(n17158) );
  OR2X1 U17983 ( .IN1(n10046), .IN2(n5752), .Q(n17160) );
  OR2X1 U17984 ( .IN1(g4521), .IN2(n16737), .Q(n17159) );
  XNOR2X1 U17985 ( .IN1(n12015), .IN2(n10071), .Q(n16737) );
  NAND2X0 U17986 ( .IN1(n17161), .IN2(n17162), .QN(n12015) );
  NOR2X0 U17987 ( .IN1(n10061), .IN2(n10060), .QN(n17162) );
  AND2X1 U17988 ( .IN1(g4483), .IN2(test_so27), .Q(n17161) );
  NAND2X0 U17989 ( .IN1(n17163), .IN2(n17152), .QN(g26963) );
  NAND2X0 U17990 ( .IN1(g6750), .IN2(n10388), .QN(n17152) );
  OR2X1 U17991 ( .IN1(n10310), .IN2(n10060), .Q(n17163) );
  NAND2X0 U17992 ( .IN1(n17150), .IN2(n17164), .QN(g26962) );
  NAND2X0 U17993 ( .IN1(test_so27), .IN2(n10515), .QN(n17164) );
  NAND2X0 U17994 ( .IN1(g6749), .IN2(n10388), .QN(n17150) );
  NAND2X0 U17995 ( .IN1(n17165), .IN2(n17154), .QN(g26961) );
  NAND2X0 U17996 ( .IN1(g6748), .IN2(n10388), .QN(n17154) );
  NAND2X0 U17997 ( .IN1(n10497), .IN2(g4483), .QN(n17165) );
  NAND2X0 U17998 ( .IN1(n17166), .IN2(n17167), .QN(g26958) );
  NAND2X0 U17999 ( .IN1(n10498), .IN2(g4455), .QN(n17167) );
  NAND2X0 U18000 ( .IN1(n17168), .IN2(n17169), .QN(g26957) );
  NAND2X0 U18001 ( .IN1(n17170), .IN2(g4434), .QN(n17169) );
  NAND2X0 U18002 ( .IN1(n17171), .IN2(n10388), .QN(n17170) );
  NAND2X0 U18003 ( .IN1(n17172), .IN2(g4392), .QN(n17171) );
  NAND2X0 U18004 ( .IN1(test_so47), .IN2(n10388), .QN(n17168) );
  NAND2X0 U18005 ( .IN1(n18479), .IN2(n17173), .QN(g26956) );
  NAND2X0 U18006 ( .IN1(n17174), .IN2(n17175), .QN(n17173) );
  NOR2X0 U18007 ( .IN1(n9679), .IN2(n17176), .QN(n17174) );
  NAND2X0 U18008 ( .IN1(n17177), .IN2(n17178), .QN(g26955) );
  NAND2X0 U18009 ( .IN1(n17179), .IN2(n17172), .QN(n17178) );
  INVX0 U18010 ( .INP(n17176), .ZN(n17172) );
  NAND2X0 U18011 ( .IN1(n17180), .IN2(g4438), .QN(n17177) );
  NAND2X0 U18012 ( .IN1(n17181), .IN2(n17182), .QN(g26954) );
  NAND2X0 U18013 ( .IN1(test_so47), .IN2(n10515), .QN(n17182) );
  NOR2X0 U18014 ( .IN1(n17183), .IN2(n17184), .QN(n17181) );
  NOR2X0 U18015 ( .IN1(n10051), .IN2(n17180), .QN(n17184) );
  NOR2X0 U18016 ( .IN1(n17176), .IN2(n17185), .QN(n17183) );
  NAND2X0 U18017 ( .IN1(n17186), .IN2(n17187), .QN(n17176) );
  NOR2X0 U18018 ( .IN1(n9336), .IN2(n17188), .QN(n17187) );
  OR2X1 U18019 ( .IN1(g4438), .IN2(test_so47), .Q(n17188) );
  NOR2X0 U18020 ( .IN1(g7245), .IN2(g7260), .QN(n17186) );
  NAND2X0 U18021 ( .IN1(n17189), .IN2(n17190), .QN(g26952) );
  NAND2X0 U18022 ( .IN1(n17191), .IN2(g4430), .QN(n17190) );
  NAND2X0 U18023 ( .IN1(n10376), .IN2(g4388), .QN(n17191) );
  NAND2X0 U18024 ( .IN1(n17192), .IN2(n10388), .QN(n17189) );
  NAND2X0 U18025 ( .IN1(n17193), .IN2(n17194), .QN(n17192) );
  NAND2X0 U18026 ( .IN1(n9679), .IN2(g4388), .QN(n17194) );
  XOR2X1 U18027 ( .IN1(g4401), .IN2(n9675), .Q(n17193) );
  OR2X1 U18028 ( .IN1(n17195), .IN2(g26953), .Q(g26951) );
  NOR2X0 U18029 ( .IN1(n9769), .IN2(n10349), .QN(n17195) );
  NAND2X0 U18030 ( .IN1(n17166), .IN2(n17196), .QN(g26950) );
  OR2X1 U18031 ( .IN1(n10311), .IN2(n9573), .Q(n17196) );
  NAND2X0 U18032 ( .IN1(n17197), .IN2(n10388), .QN(n17166) );
  NAND2X0 U18033 ( .IN1(n17198), .IN2(n17199), .QN(n17197) );
  NAND2X0 U18034 ( .IN1(n17200), .IN2(g4392), .QN(n17199) );
  NAND2X0 U18035 ( .IN1(n17201), .IN2(n17202), .QN(g26949) );
  NAND2X0 U18036 ( .IN1(n17203), .IN2(g4401), .QN(n17202) );
  NAND2X0 U18037 ( .IN1(n17204), .IN2(n10388), .QN(n17203) );
  NAND2X0 U18038 ( .IN1(n17205), .IN2(g4392), .QN(n17204) );
  NAND2X0 U18039 ( .IN1(n10377), .IN2(g4411), .QN(n17201) );
  NAND2X0 U18040 ( .IN1(n9569), .IN2(n17206), .QN(g26948) );
  NAND2X0 U18041 ( .IN1(n17207), .IN2(n17175), .QN(n17206) );
  INVX0 U18042 ( .INP(n17185), .ZN(n17175) );
  NOR2X0 U18043 ( .IN1(n9676), .IN2(n17200), .QN(n17207) );
  NAND2X0 U18044 ( .IN1(n17208), .IN2(n17209), .QN(g26947) );
  NAND2X0 U18045 ( .IN1(n10497), .IN2(g4388), .QN(n17209) );
  NAND2X0 U18046 ( .IN1(n17210), .IN2(n10388), .QN(n17208) );
  NAND2X0 U18047 ( .IN1(n17198), .IN2(n17211), .QN(n17210) );
  NAND2X0 U18048 ( .IN1(n17212), .IN2(n17200), .QN(n17211) );
  XOR2X1 U18049 ( .IN1(n9578), .IN2(n5714), .Q(n17212) );
  NAND2X0 U18050 ( .IN1(n17213), .IN2(n9573), .QN(n17198) );
  NOR2X0 U18051 ( .IN1(n17200), .IN2(g4392), .QN(n17213) );
  NAND2X0 U18052 ( .IN1(n17214), .IN2(n17215), .QN(g26946) );
  NAND2X0 U18053 ( .IN1(n17179), .IN2(n17205), .QN(n17215) );
  INVX0 U18054 ( .INP(n17200), .ZN(n17205) );
  NOR2X0 U18055 ( .IN1(n5710), .IN2(n10458), .QN(n17179) );
  NAND2X0 U18056 ( .IN1(n17180), .IN2(g4375), .QN(n17214) );
  NAND2X0 U18057 ( .IN1(n17216), .IN2(n17217), .QN(g26945) );
  NAND2X0 U18058 ( .IN1(n10497), .IN2(g4411), .QN(n17217) );
  NOR2X0 U18059 ( .IN1(n17218), .IN2(n17219), .QN(n17216) );
  NOR2X0 U18060 ( .IN1(n9578), .IN2(n17180), .QN(n17219) );
  NAND2X0 U18061 ( .IN1(n5714), .IN2(n10388), .QN(n17180) );
  NOR2X0 U18062 ( .IN1(n17200), .IN2(n17185), .QN(n17218) );
  NAND2X0 U18063 ( .IN1(n5710), .IN2(n10388), .QN(n17185) );
  NAND2X0 U18064 ( .IN1(n17220), .IN2(n17221), .QN(n17200) );
  NOR2X0 U18065 ( .IN1(g4411), .IN2(n17222), .QN(n17221) );
  NAND2X0 U18066 ( .IN1(n9578), .IN2(n9569), .QN(n17222) );
  NOR2X0 U18067 ( .IN1(g7257), .IN2(g7243), .QN(n17220) );
  NOR2X0 U18068 ( .IN1(n10479), .IN2(n17223), .QN(g26944) );
  NOR2X0 U18069 ( .IN1(n17224), .IN2(n17225), .QN(n17223) );
  NAND2X0 U18070 ( .IN1(n11172), .IN2(test_so81), .QN(n17225) );
  NOR2X0 U18071 ( .IN1(g135), .IN2(n17226), .QN(n11172) );
  NOR2X0 U18072 ( .IN1(n17227), .IN2(n17228), .QN(n17226) );
  NAND2X0 U18073 ( .IN1(n17229), .IN2(n17230), .QN(n17228) );
  NAND2X0 U18074 ( .IN1(n17231), .IN2(g4584), .QN(n17230) );
  NOR2X0 U18075 ( .IN1(g4608), .IN2(n17232), .QN(n17231) );
  NAND2X0 U18076 ( .IN1(n5365), .IN2(g4593), .QN(n17232) );
  NAND2X0 U18077 ( .IN1(n17233), .IN2(n5539), .QN(n17229) );
  NOR2X0 U18078 ( .IN1(n5274), .IN2(g4593), .QN(n17233) );
  NOR2X0 U18079 ( .IN1(n17234), .IN2(n17235), .QN(n17227) );
  NAND2X0 U18080 ( .IN1(n17236), .IN2(n5608), .QN(n17235) );
  XOR2X1 U18081 ( .IN1(g4593), .IN2(n5365), .Q(n17236) );
  XOR2X1 U18082 ( .IN1(n5539), .IN2(n5274), .Q(n17234) );
  NAND2X0 U18083 ( .IN1(n17237), .IN2(n11850), .QN(n17224) );
  NOR2X0 U18084 ( .IN1(n5844), .IN2(n5348), .QN(n17237) );
  NAND2X0 U18085 ( .IN1(n17238), .IN2(n17239), .QN(g26940) );
  NAND2X0 U18086 ( .IN1(n10497), .IN2(g4153), .QN(n17239) );
  NAND2X0 U18087 ( .IN1(n14773), .IN2(n10387), .QN(n17238) );
  NAND2X0 U18088 ( .IN1(n17240), .IN2(n17241), .QN(n14773) );
  NAND2X0 U18089 ( .IN1(g116), .IN2(g4157), .QN(n17241) );
  NAND2X0 U18090 ( .IN1(g114), .IN2(n5983), .QN(n17240) );
  NAND2X0 U18091 ( .IN1(n17242), .IN2(n17243), .QN(g26939) );
  OR2X1 U18092 ( .IN1(n10311), .IN2(n9913), .Q(n17243) );
  NAND2X0 U18093 ( .IN1(n14771), .IN2(n10387), .QN(n17242) );
  NAND2X0 U18094 ( .IN1(n17244), .IN2(n17245), .QN(n14771) );
  NAND2X0 U18095 ( .IN1(g124), .IN2(g4146), .QN(n17245) );
  NAND2X0 U18096 ( .IN1(g120), .IN2(n5981), .QN(n17244) );
  NAND2X0 U18097 ( .IN1(n17246), .IN2(n14067), .QN(g26938) );
  NOR2X0 U18098 ( .IN1(n17247), .IN2(n17248), .QN(n17246) );
  NOR2X0 U18099 ( .IN1(n10479), .IN2(n17249), .QN(n17248) );
  XNOR2X1 U18100 ( .IN1(n9739), .IN2(n16773), .Q(n17249) );
  NAND2X0 U18101 ( .IN1(n17250), .IN2(g4141), .QN(n16773) );
  NOR2X0 U18102 ( .IN1(n5612), .IN2(n10347), .QN(n17247) );
  NAND2X0 U18103 ( .IN1(n17251), .IN2(n17252), .QN(g26934) );
  NAND2X0 U18104 ( .IN1(n4888), .IN2(g2827), .QN(n17252) );
  NOR2X0 U18105 ( .IN1(n17253), .IN2(n17254), .QN(n17251) );
  NOR2X0 U18106 ( .IN1(n10357), .IN2(n10149), .QN(n17254) );
  NOR2X0 U18107 ( .IN1(test_so34), .IN2(n17255), .QN(n17253) );
  NAND2X0 U18108 ( .IN1(n17256), .IN2(n17257), .QN(g26933) );
  NAND2X0 U18109 ( .IN1(n4888), .IN2(test_so37), .QN(n17257) );
  NOR2X0 U18110 ( .IN1(n17258), .IN2(n17259), .QN(n17256) );
  NOR2X0 U18111 ( .IN1(n9608), .IN2(n10346), .QN(n17259) );
  NOR2X0 U18112 ( .IN1(n17255), .IN2(g2461), .QN(n17258) );
  NAND2X0 U18113 ( .IN1(n17260), .IN2(n17261), .QN(g26932) );
  NAND2X0 U18114 ( .IN1(n4888), .IN2(g2811), .QN(n17261) );
  NOR2X0 U18115 ( .IN1(n17262), .IN2(n17263), .QN(n17260) );
  NOR2X0 U18116 ( .IN1(n9605), .IN2(n10352), .QN(n17263) );
  NOR2X0 U18117 ( .IN1(n17255), .IN2(g2327), .QN(n17262) );
  NAND2X0 U18118 ( .IN1(n17264), .IN2(n17265), .QN(g26931) );
  NAND2X0 U18119 ( .IN1(n4888), .IN2(g2799), .QN(n17265) );
  NOR2X0 U18120 ( .IN1(n17266), .IN2(n17267), .QN(n17264) );
  NOR2X0 U18121 ( .IN1(n9588), .IN2(n10347), .QN(n17267) );
  NOR2X0 U18122 ( .IN1(n17255), .IN2(g2193), .QN(n17266) );
  NAND2X0 U18123 ( .IN1(n17268), .IN2(n17269), .QN(g26930) );
  NAND2X0 U18124 ( .IN1(n4888), .IN2(g2795), .QN(n17269) );
  NOR2X0 U18125 ( .IN1(n17270), .IN2(n17271), .QN(n17268) );
  NOR2X0 U18126 ( .IN1(n9607), .IN2(n10347), .QN(n17271) );
  NOR2X0 U18127 ( .IN1(test_so59), .IN2(n17255), .QN(n17270) );
  NAND2X0 U18128 ( .IN1(n17272), .IN2(n17273), .QN(g26929) );
  NAND2X0 U18129 ( .IN1(n4888), .IN2(g2791), .QN(n17273) );
  NOR2X0 U18130 ( .IN1(n17274), .IN2(n17275), .QN(n17272) );
  NOR2X0 U18131 ( .IN1(n9604), .IN2(n10347), .QN(n17275) );
  NOR2X0 U18132 ( .IN1(n17255), .IN2(g1902), .QN(n17274) );
  NAND2X0 U18133 ( .IN1(n17276), .IN2(n17277), .QN(g26928) );
  NAND2X0 U18134 ( .IN1(n4888), .IN2(g2779), .QN(n17277) );
  NOR2X0 U18135 ( .IN1(n17278), .IN2(n17279), .QN(n17276) );
  NOR2X0 U18136 ( .IN1(n9610), .IN2(n10347), .QN(n17279) );
  NOR2X0 U18137 ( .IN1(n17255), .IN2(g1768), .QN(n17278) );
  NAND2X0 U18138 ( .IN1(n17280), .IN2(n17281), .QN(g26927) );
  NAND2X0 U18139 ( .IN1(n4888), .IN2(g2767), .QN(n17281) );
  NOR2X0 U18140 ( .IN1(n17282), .IN2(n17283), .QN(n17280) );
  NOR2X0 U18141 ( .IN1(n9587), .IN2(n10348), .QN(n17283) );
  NOR2X0 U18142 ( .IN1(n17255), .IN2(g1632), .QN(n17282) );
  NAND2X0 U18143 ( .IN1(n17284), .IN2(n4888), .QN(n17255) );
  NOR2X0 U18144 ( .IN1(n11632), .IN2(n17285), .QN(n17284) );
  NOR2X0 U18145 ( .IN1(test_so30), .IN2(g2748), .QN(n17285) );
  INVX0 U18146 ( .INP(n11649), .ZN(n11632) );
  NAND2X0 U18147 ( .IN1(n17286), .IN2(test_so30), .QN(n11649) );
  AND2X1 U18148 ( .IN1(g2735), .IN2(n3505), .Q(n17286) );
  NOR2X0 U18149 ( .IN1(n5349), .IN2(n5516), .QN(n3505) );
  NAND2X0 U18150 ( .IN1(n17287), .IN2(n17288), .QN(g26926) );
  NAND2X0 U18151 ( .IN1(n17289), .IN2(n3730), .QN(n17288) );
  XOR2X1 U18152 ( .IN1(g2724), .IN2(n15161), .Q(n17289) );
  NOR2X0 U18153 ( .IN1(n5465), .IN2(n5299), .QN(n15161) );
  NAND2X0 U18154 ( .IN1(n10498), .IN2(g2719), .QN(n17287) );
  NAND2X0 U18155 ( .IN1(n17290), .IN2(n17291), .QN(g26925) );
  NAND2X0 U18156 ( .IN1(n10498), .IN2(g1532), .QN(n17291) );
  NAND2X0 U18157 ( .IN1(n17292), .IN2(n10387), .QN(n17290) );
  NAND2X0 U18158 ( .IN1(n15490), .IN2(n17293), .QN(n17292) );
  NAND2X0 U18159 ( .IN1(n17294), .IN2(g1536), .QN(n17293) );
  OR2X1 U18160 ( .IN1(n15476), .IN2(n9572), .Q(n17294) );
  INVX0 U18161 ( .INP(n15474), .ZN(n15476) );
  NOR2X0 U18162 ( .IN1(n15482), .IN2(n9775), .QN(n15474) );
  NAND2X0 U18163 ( .IN1(n17295), .IN2(n12991), .QN(n15482) );
  NOR2X0 U18164 ( .IN1(n5302), .IN2(n17296), .QN(n17295) );
  NOR2X0 U18165 ( .IN1(g1532), .IN2(n17297), .QN(n17296) );
  NAND2X0 U18166 ( .IN1(g1339), .IN2(g1521), .QN(n17297) );
  INVX0 U18167 ( .INP(n4173), .ZN(n15490) );
  NAND2X0 U18168 ( .IN1(n17298), .IN2(n17299), .QN(g26924) );
  NAND2X0 U18169 ( .IN1(n17300), .IN2(n5289), .QN(n17299) );
  NOR2X0 U18170 ( .IN1(n17301), .IN2(n17302), .QN(n17298) );
  NOR2X0 U18171 ( .IN1(n5696), .IN2(n10348), .QN(n17302) );
  NOR2X0 U18172 ( .IN1(n10479), .IN2(n17303), .QN(n17301) );
  OR2X1 U18173 ( .IN1(n17300), .IN2(n5289), .Q(n17303) );
  AND2X1 U18174 ( .IN1(n17304), .IN2(n17305), .Q(n17300) );
  NOR2X0 U18175 ( .IN1(test_so49), .IN2(n5696), .QN(n17305) );
  NAND2X0 U18176 ( .IN1(n17306), .IN2(n17307), .QN(g26923) );
  NAND2X0 U18177 ( .IN1(n17308), .IN2(n5290), .QN(n17307) );
  NOR2X0 U18178 ( .IN1(n17309), .IN2(n17310), .QN(n17306) );
  NOR2X0 U18179 ( .IN1(n5693), .IN2(n10347), .QN(n17310) );
  NOR2X0 U18180 ( .IN1(n10479), .IN2(n17311), .QN(n17309) );
  OR2X1 U18181 ( .IN1(n17308), .IN2(n5290), .Q(n17311) );
  AND2X1 U18182 ( .IN1(n17304), .IN2(n17312), .Q(n17308) );
  NOR2X0 U18183 ( .IN1(n5693), .IN2(n10127), .QN(n17312) );
  NOR2X0 U18184 ( .IN1(n16148), .IN2(n17313), .QN(n17304) );
  INVX0 U18185 ( .INP(n17314), .ZN(n17313) );
  NAND2X0 U18186 ( .IN1(g13272), .IN2(g1514), .QN(n16148) );
  NAND2X0 U18187 ( .IN1(n17315), .IN2(n17316), .QN(g26922) );
  OR2X1 U18188 ( .IN1(n17317), .IN2(g1448), .Q(n17316) );
  NOR2X0 U18189 ( .IN1(n17318), .IN2(n17319), .QN(n17315) );
  NOR2X0 U18190 ( .IN1(n5866), .IN2(n10348), .QN(n17319) );
  NOR2X0 U18191 ( .IN1(n10479), .IN2(n17320), .QN(n17318) );
  NAND2X0 U18192 ( .IN1(n17317), .IN2(g1448), .QN(n17320) );
  NAND2X0 U18193 ( .IN1(n17321), .IN2(n17314), .QN(n17317) );
  NOR2X0 U18194 ( .IN1(n5866), .IN2(n16125), .QN(n17321) );
  NAND2X0 U18195 ( .IN1(n12991), .IN2(g13272), .QN(n16125) );
  NOR2X0 U18196 ( .IN1(g1514), .IN2(n10127), .QN(n12991) );
  NAND2X0 U18197 ( .IN1(n17322), .IN2(n17323), .QN(g26921) );
  OR2X1 U18198 ( .IN1(n10311), .IN2(n9966), .Q(n17323) );
  NAND2X0 U18199 ( .IN1(n17324), .IN2(n10387), .QN(n17322) );
  NOR2X0 U18200 ( .IN1(test_so68), .IN2(n17325), .QN(n17324) );
  XNOR2X1 U18201 ( .IN1(n9753), .IN2(n17326), .Q(n17325) );
  NAND2X0 U18202 ( .IN1(n17327), .IN2(n17328), .QN(g26920) );
  NAND2X0 U18203 ( .IN1(n10497), .IN2(g1384), .QN(n17328) );
  NAND2X0 U18204 ( .IN1(n17329), .IN2(n10387), .QN(n17327) );
  NAND2X0 U18205 ( .IN1(n17330), .IN2(n17331), .QN(n17329) );
  OR2X1 U18206 ( .IN1(n4915), .IN2(n9758), .Q(n17331) );
  AND2X1 U18207 ( .IN1(n17332), .IN2(n17333), .Q(n4915) );
  NAND2X0 U18208 ( .IN1(n9592), .IN2(g1351), .QN(n17333) );
  NAND2X0 U18209 ( .IN1(n4913), .IN2(g1351), .QN(n17330) );
  NAND2X0 U18210 ( .IN1(n17334), .IN2(n17335), .QN(g26919) );
  NAND2X0 U18211 ( .IN1(n10497), .IN2(g1266), .QN(n17335) );
  NOR2X0 U18212 ( .IN1(n17336), .IN2(n17337), .QN(n17334) );
  NOR2X0 U18213 ( .IN1(test_so77), .IN2(n17338), .QN(n17337) );
  NOR2X0 U18214 ( .IN1(n870), .IN2(n17339), .QN(n17336) );
  NAND2X0 U18215 ( .IN1(test_so77), .IN2(n13309), .QN(n17339) );
  INVX0 U18216 ( .INP(n17338), .ZN(n870) );
  NAND2X0 U18217 ( .IN1(n17340), .IN2(g12923), .QN(n17338) );
  NOR2X0 U18218 ( .IN1(n9743), .IN2(n9742), .QN(n17340) );
  NAND2X0 U18219 ( .IN1(n17341), .IN2(n17342), .QN(g26918) );
  NAND2X0 U18220 ( .IN1(n10497), .IN2(g1189), .QN(n17342) );
  NAND2X0 U18221 ( .IN1(n17343), .IN2(n10387), .QN(n17341) );
  NAND2X0 U18222 ( .IN1(n15531), .IN2(n17344), .QN(n17343) );
  NAND2X0 U18223 ( .IN1(n17345), .IN2(g1193), .QN(n17344) );
  OR2X1 U18224 ( .IN1(n15517), .IN2(n9571), .Q(n17345) );
  INVX0 U18225 ( .INP(n15515), .ZN(n15517) );
  NOR2X0 U18226 ( .IN1(n15523), .IN2(n9776), .QN(n15515) );
  NAND2X0 U18227 ( .IN1(n17346), .IN2(n13234), .QN(n15523) );
  NOR2X0 U18228 ( .IN1(n5304), .IN2(n17347), .QN(n17346) );
  NOR2X0 U18229 ( .IN1(g1189), .IN2(n17348), .QN(n17347) );
  NAND2X0 U18230 ( .IN1(g1178), .IN2(g996), .QN(n17348) );
  INVX0 U18231 ( .INP(n4191), .ZN(n15531) );
  NAND2X0 U18232 ( .IN1(n17349), .IN2(n17350), .QN(g26917) );
  OR2X1 U18233 ( .IN1(n17351), .IN2(g1135), .Q(n17350) );
  NOR2X0 U18234 ( .IN1(n17352), .IN2(n17353), .QN(n17349) );
  NOR2X0 U18235 ( .IN1(n5697), .IN2(n10348), .QN(n17353) );
  NOR2X0 U18236 ( .IN1(n10479), .IN2(n17354), .QN(n17352) );
  NAND2X0 U18237 ( .IN1(n17351), .IN2(g1135), .QN(n17354) );
  NAND2X0 U18238 ( .IN1(n17355), .IN2(n17356), .QN(n17351) );
  NOR2X0 U18239 ( .IN1(n5697), .IN2(g1183), .QN(n17356) );
  NAND2X0 U18240 ( .IN1(n17357), .IN2(n17358), .QN(g26916) );
  OR2X1 U18241 ( .IN1(n17359), .IN2(g1129), .Q(n17358) );
  NOR2X0 U18242 ( .IN1(n17360), .IN2(n17361), .QN(n17357) );
  NOR2X0 U18243 ( .IN1(n5692), .IN2(n10348), .QN(n17361) );
  NOR2X0 U18244 ( .IN1(n10479), .IN2(n17362), .QN(n17360) );
  NAND2X0 U18245 ( .IN1(n17359), .IN2(g1129), .QN(n17362) );
  NAND2X0 U18246 ( .IN1(n17355), .IN2(n17363), .QN(n17359) );
  NOR2X0 U18247 ( .IN1(n5692), .IN2(n5599), .QN(n17363) );
  NOR2X0 U18248 ( .IN1(n16201), .IN2(n17364), .QN(n17355) );
  NAND2X0 U18249 ( .IN1(g13259), .IN2(g1171), .QN(n16201) );
  NAND2X0 U18250 ( .IN1(n17365), .IN2(n17366), .QN(g26915) );
  NAND2X0 U18251 ( .IN1(n17367), .IN2(n5478), .QN(n17366) );
  NOR2X0 U18252 ( .IN1(n17368), .IN2(n17369), .QN(n17365) );
  NOR2X0 U18253 ( .IN1(n10357), .IN2(n10148), .QN(n17369) );
  NOR2X0 U18254 ( .IN1(n10479), .IN2(n17370), .QN(n17368) );
  OR2X1 U18255 ( .IN1(n17367), .IN2(n5478), .Q(n17370) );
  AND2X1 U18256 ( .IN1(n17371), .IN2(n17372), .Q(n17367) );
  NOR2X0 U18257 ( .IN1(n16178), .IN2(n10148), .QN(n17371) );
  NAND2X0 U18258 ( .IN1(n13234), .IN2(g13259), .QN(n16178) );
  NOR2X0 U18259 ( .IN1(g1171), .IN2(n5599), .QN(n13234) );
  NAND2X0 U18260 ( .IN1(n17373), .IN2(n17374), .QN(g26914) );
  NAND2X0 U18261 ( .IN1(n10497), .IN2(g1052), .QN(n17374) );
  NAND2X0 U18262 ( .IN1(n17375), .IN2(n10387), .QN(n17373) );
  NOR2X0 U18263 ( .IN1(n17376), .IN2(g979), .QN(n17375) );
  XNOR2X1 U18264 ( .IN1(n9754), .IN2(n17377), .Q(n17376) );
  NAND2X0 U18265 ( .IN1(n17378), .IN2(n17379), .QN(g26913) );
  NAND2X0 U18266 ( .IN1(n4938), .IN2(n17380), .QN(n17379) );
  NOR2X0 U18267 ( .IN1(n17381), .IN2(n17382), .QN(n17378) );
  NOR2X0 U18268 ( .IN1(n10479), .IN2(n17383), .QN(n17382) );
  OR2X1 U18269 ( .IN1(n4940), .IN2(n9910), .Q(n17383) );
  AND2X1 U18270 ( .IN1(n17384), .IN2(n17385), .Q(n4940) );
  NAND2X0 U18271 ( .IN1(n9591), .IN2(g1008), .QN(n17385) );
  NOR2X0 U18272 ( .IN1(n9591), .IN2(n10348), .QN(n17381) );
  NAND2X0 U18273 ( .IN1(n17386), .IN2(n17387), .QN(g26912) );
  NAND2X0 U18274 ( .IN1(n10498), .IN2(g921), .QN(n17387) );
  NOR2X0 U18275 ( .IN1(n17388), .IN2(n17389), .QN(n17386) );
  NOR2X0 U18276 ( .IN1(g936), .IN2(n10793), .QN(n17389) );
  NOR2X0 U18277 ( .IN1(n5557), .IN2(n17390), .QN(n17388) );
  NAND2X0 U18278 ( .IN1(n13328), .IN2(n10793), .QN(n17390) );
  NAND2X0 U18279 ( .IN1(n17391), .IN2(g12919), .QN(n10793) );
  NOR2X0 U18280 ( .IN1(n9741), .IN2(n9740), .QN(n17391) );
  XOR2X1 U18281 ( .IN1(n17392), .IN2(n5682), .Q(g26910) );
  NAND2X0 U18282 ( .IN1(n5305), .IN2(n10387), .QN(n17392) );
  NAND2X0 U18283 ( .IN1(n17393), .IN2(n17394), .QN(g26909) );
  NAND2X0 U18284 ( .IN1(n10498), .IN2(g890), .QN(n17394) );
  NAND2X0 U18285 ( .IN1(n17395), .IN2(n10387), .QN(n17393) );
  NAND2X0 U18286 ( .IN1(n17396), .IN2(n17397), .QN(n17395) );
  NAND2X0 U18287 ( .IN1(n5431), .IN2(g862), .QN(n17397) );
  NAND2X0 U18288 ( .IN1(n5305), .IN2(g896), .QN(n17396) );
  NAND2X0 U18289 ( .IN1(n17398), .IN2(n17399), .QN(g26908) );
  NAND2X0 U18290 ( .IN1(n4945), .IN2(g446), .QN(n17399) );
  NOR2X0 U18291 ( .IN1(n17400), .IN2(n17401), .QN(n17398) );
  NOR2X0 U18292 ( .IN1(n6008), .IN2(n10349), .QN(n17401) );
  NOR2X0 U18293 ( .IN1(n9598), .IN2(n17402), .QN(n17400) );
  NAND2X0 U18294 ( .IN1(n17403), .IN2(n17404), .QN(g26907) );
  NAND2X0 U18295 ( .IN1(n4945), .IN2(g246), .QN(n17404) );
  NOR2X0 U18296 ( .IN1(n17405), .IN2(n17406), .QN(n17403) );
  NOR2X0 U18297 ( .IN1(n9783), .IN2(n10349), .QN(n17406) );
  NOR2X0 U18298 ( .IN1(n9600), .IN2(n17402), .QN(n17405) );
  NAND2X0 U18299 ( .IN1(n17407), .IN2(n17408), .QN(g26906) );
  NAND2X0 U18300 ( .IN1(n4945), .IN2(g269), .QN(n17408) );
  NOR2X0 U18301 ( .IN1(n17409), .IN2(n17410), .QN(n17407) );
  NOR2X0 U18302 ( .IN1(n9909), .IN2(n10349), .QN(n17410) );
  NOR2X0 U18303 ( .IN1(n9597), .IN2(n17402), .QN(n17409) );
  NAND2X0 U18304 ( .IN1(n17411), .IN2(n17412), .QN(g26905) );
  NAND2X0 U18305 ( .IN1(n4945), .IN2(g239), .QN(n17412) );
  NOR2X0 U18306 ( .IN1(n17413), .IN2(n17414), .QN(n17411) );
  NOR2X0 U18307 ( .IN1(n9782), .IN2(n10349), .QN(n17414) );
  NOR2X0 U18308 ( .IN1(n9596), .IN2(n17402), .QN(n17413) );
  NAND2X0 U18309 ( .IN1(n17415), .IN2(n17416), .QN(g26904) );
  NAND2X0 U18310 ( .IN1(n4945), .IN2(g262), .QN(n17416) );
  NOR2X0 U18311 ( .IN1(n17417), .IN2(n17418), .QN(n17415) );
  NOR2X0 U18312 ( .IN1(n9908), .IN2(n10349), .QN(n17418) );
  NOR2X0 U18313 ( .IN1(n9594), .IN2(n17402), .QN(n17417) );
  NAND2X0 U18314 ( .IN1(n17419), .IN2(n17420), .QN(g26903) );
  NAND2X0 U18315 ( .IN1(n4945), .IN2(g232), .QN(n17420) );
  NOR2X0 U18316 ( .IN1(n17421), .IN2(n17422), .QN(n17419) );
  NOR2X0 U18317 ( .IN1(n9781), .IN2(n10349), .QN(n17422) );
  NOR2X0 U18318 ( .IN1(n9595), .IN2(n17402), .QN(n17421) );
  NAND2X0 U18319 ( .IN1(n17423), .IN2(n17424), .QN(g26902) );
  NAND2X0 U18320 ( .IN1(n4945), .IN2(g255), .QN(n17424) );
  NOR2X0 U18321 ( .IN1(n17425), .IN2(n17426), .QN(n17423) );
  NOR2X0 U18322 ( .IN1(n5597), .IN2(n10350), .QN(n17426) );
  NOR2X0 U18323 ( .IN1(n9593), .IN2(n17402), .QN(n17425) );
  NAND2X0 U18324 ( .IN1(n17427), .IN2(n17428), .QN(g26901) );
  NAND2X0 U18325 ( .IN1(n4945), .IN2(g225), .QN(n17428) );
  NOR2X0 U18326 ( .IN1(n17429), .IN2(n17430), .QN(n17427) );
  NOR2X0 U18327 ( .IN1(n9598), .IN2(n10350), .QN(n17430) );
  NOR2X0 U18328 ( .IN1(n9599), .IN2(n17402), .QN(n17429) );
  OR2X1 U18329 ( .IN1(n10457), .IN2(n4946), .Q(n17402) );
  NAND2X0 U18330 ( .IN1(n17431), .IN2(n5682), .QN(n4946) );
  NOR2X0 U18331 ( .IN1(n5305), .IN2(g896), .QN(n17431) );
  NAND2X0 U18332 ( .IN1(n17432), .IN2(n17433), .QN(g26899) );
  NAND2X0 U18333 ( .IN1(n17434), .IN2(n42), .QN(n17433) );
  XNOR2X1 U18334 ( .IN1(n4814), .IN2(n5422), .Q(n17434) );
  AND2X1 U18335 ( .IN1(n17435), .IN2(n4948), .Q(n4814) );
  NOR2X0 U18336 ( .IN1(n5822), .IN2(n10065), .QN(n17435) );
  NAND2X0 U18337 ( .IN1(n10497), .IN2(g832), .QN(n17432) );
  NAND2X0 U18338 ( .IN1(n17436), .IN2(n17437), .QN(g26898) );
  NAND2X0 U18339 ( .IN1(n17438), .IN2(n17439), .QN(n17437) );
  NAND2X0 U18340 ( .IN1(n17440), .IN2(n17441), .QN(n17439) );
  NAND2X0 U18341 ( .IN1(n9713), .IN2(n10387), .QN(n17441) );
  NAND2X0 U18342 ( .IN1(n17442), .IN2(g843), .QN(n17436) );
  NAND2X0 U18343 ( .IN1(n17443), .IN2(n10391), .QN(n17442) );
  NAND2X0 U18344 ( .IN1(n17444), .IN2(n17445), .QN(n17443) );
  NOR2X0 U18345 ( .IN1(n5562), .IN2(g812), .QN(n17444) );
  NAND2X0 U18346 ( .IN1(n17446), .IN2(n17447), .QN(g26897) );
  NAND2X0 U18347 ( .IN1(n17448), .IN2(g753), .QN(n17447) );
  OR2X1 U18348 ( .IN1(n17448), .IN2(n5732), .Q(n17446) );
  NOR2X0 U18349 ( .IN1(n17449), .IN2(n10459), .QN(n17448) );
  NAND2X0 U18350 ( .IN1(n17450), .IN2(n17451), .QN(g26896) );
  NAND2X0 U18351 ( .IN1(n4956), .IN2(n17452), .QN(n17451) );
  NOR2X0 U18352 ( .IN1(n17453), .IN2(n17454), .QN(n17450) );
  NOR2X0 U18353 ( .IN1(n9790), .IN2(n17455), .QN(n17454) );
  AND2X1 U18354 ( .IN1(g29212), .IN2(n17455), .Q(n17453) );
  NOR2X0 U18355 ( .IN1(n17452), .IN2(n10459), .QN(n17455) );
  INVX0 U18356 ( .INP(n10107), .ZN(n17452) );
  NAND2X0 U18357 ( .IN1(n17456), .IN2(n17457), .QN(n10107) );
  NOR2X0 U18358 ( .IN1(n16280), .IN2(n17089), .QN(n17457) );
  NOR2X0 U18359 ( .IN1(g504), .IN2(n10135), .QN(n17456) );
  NAND2X0 U18360 ( .IN1(n17458), .IN2(n17459), .QN(g26895) );
  NAND2X0 U18361 ( .IN1(n10498), .IN2(g562), .QN(n17459) );
  NOR2X0 U18362 ( .IN1(n17460), .IN2(n17461), .QN(n17458) );
  NOR2X0 U18363 ( .IN1(g568), .IN2(n10788), .QN(n17461) );
  NOR2X0 U18364 ( .IN1(n5335), .IN2(n17462), .QN(n17460) );
  NAND2X0 U18365 ( .IN1(n2421), .IN2(n10788), .QN(n17462) );
  NAND2X0 U18366 ( .IN1(n17463), .IN2(n4959), .QN(n10788) );
  NOR2X0 U18367 ( .IN1(n9584), .IN2(n17464), .QN(n17463) );
  NAND2X0 U18368 ( .IN1(n17465), .IN2(n17466), .QN(g26894) );
  NAND2X0 U18369 ( .IN1(n17467), .IN2(n17084), .QN(n17466) );
  NOR2X0 U18370 ( .IN1(n17468), .IN2(n17469), .QN(n17467) );
  NOR2X0 U18371 ( .IN1(n5327), .IN2(n17470), .QN(n17469) );
  NAND2X0 U18372 ( .IN1(n17471), .IN2(n17472), .QN(n17470) );
  NAND2X0 U18373 ( .IN1(n17088), .IN2(n10406), .QN(n17471) );
  NOR2X0 U18374 ( .IN1(n17473), .IN2(g528), .QN(n17468) );
  NOR2X0 U18375 ( .IN1(n17474), .IN2(n17475), .QN(n17473) );
  NAND2X0 U18376 ( .IN1(n17476), .IN2(n17089), .QN(n17475) );
  NAND2X0 U18377 ( .IN1(n17477), .IN2(n5327), .QN(n17089) );
  NOR2X0 U18378 ( .IN1(n5820), .IN2(n5708), .QN(n17477) );
  NAND2X0 U18379 ( .IN1(n10498), .IN2(g518), .QN(n17465) );
  NAND2X0 U18380 ( .IN1(n17478), .IN2(n17479), .QN(g26893) );
  NAND2X0 U18381 ( .IN1(n10498), .IN2(g355), .QN(n17479) );
  NAND2X0 U18382 ( .IN1(n17480), .IN2(n10406), .QN(n17478) );
  NAND2X0 U18383 ( .IN1(n17481), .IN2(n17482), .QN(n17480) );
  NAND2X0 U18384 ( .IN1(g29211), .IN2(n10124), .QN(n17482) );
  OR2X1 U18385 ( .IN1(n10124), .IN2(n17483), .Q(n17481) );
  NAND2X0 U18386 ( .IN1(n17484), .IN2(n17485), .QN(g26892) );
  NAND2X0 U18387 ( .IN1(n17486), .IN2(n10124), .QN(n17485) );
  NOR2X0 U18388 ( .IN1(n17483), .IN2(n10459), .QN(n17486) );
  NOR2X0 U18389 ( .IN1(g355), .IN2(g333), .QN(n17483) );
  NAND2X0 U18390 ( .IN1(test_so17), .IN2(n10515), .QN(n17484) );
  NAND2X0 U18391 ( .IN1(n17487), .IN2(n17488), .QN(g26891) );
  OR2X1 U18392 ( .IN1(n10308), .IN2(n5860), .Q(n17488) );
  NAND2X0 U18393 ( .IN1(n17489), .IN2(n5860), .QN(n17487) );
  NOR2X0 U18394 ( .IN1(n9613), .IN2(n10459), .QN(n17489) );
  NAND2X0 U18395 ( .IN1(n17490), .IN2(n17491), .QN(g26890) );
  NAND2X0 U18396 ( .IN1(n5860), .IN2(n10406), .QN(n17491) );
  NAND2X0 U18397 ( .IN1(n10498), .IN2(g333), .QN(n17490) );
  NAND2X0 U18398 ( .IN1(n17492), .IN2(n17493), .QN(g26889) );
  NAND2X0 U18399 ( .IN1(n10498), .IN2(g29211), .QN(n17493) );
  NAND2X0 U18400 ( .IN1(n17494), .IN2(n10406), .QN(n17492) );
  NOR2X0 U18401 ( .IN1(n9306), .IN2(n17495), .QN(n17494) );
  NAND2X0 U18402 ( .IN1(n17496), .IN2(g329), .QN(n17495) );
  NAND2X0 U18403 ( .IN1(n17497), .IN2(n17498), .QN(g26888) );
  OR2X1 U18404 ( .IN1(n10457), .IN2(n9663), .Q(n17498) );
  NAND2X0 U18405 ( .IN1(n10499), .IN2(g29216), .QN(n17497) );
  NAND2X0 U18406 ( .IN1(n17499), .IN2(n17500), .QN(g26887) );
  NOR2X0 U18407 ( .IN1(n17501), .IN2(n17502), .QN(n17499) );
  NOR2X0 U18408 ( .IN1(n10478), .IN2(n17503), .QN(n17502) );
  NAND2X0 U18409 ( .IN1(n5317), .IN2(g324), .QN(n17503) );
  NOR2X0 U18410 ( .IN1(n5824), .IN2(n10350), .QN(n17501) );
  NAND2X0 U18411 ( .IN1(n17504), .IN2(n17505), .QN(g26886) );
  OR2X1 U18412 ( .IN1(n17500), .IN2(n17496), .Q(n17505) );
  NOR2X0 U18413 ( .IN1(n17506), .IN2(n17507), .QN(n17504) );
  NOR2X0 U18414 ( .IN1(n5317), .IN2(n10350), .QN(n17507) );
  NOR2X0 U18415 ( .IN1(n10478), .IN2(n17508), .QN(n17506) );
  NAND2X0 U18416 ( .IN1(n17496), .IN2(g336), .QN(n17508) );
  INVX0 U18417 ( .INP(n17509), .ZN(n17496) );
  NAND2X0 U18418 ( .IN1(n17510), .IN2(n17511), .QN(g26884) );
  NAND2X0 U18419 ( .IN1(n10499), .IN2(g329), .QN(n17511) );
  NAND2X0 U18420 ( .IN1(n17512), .IN2(n10406), .QN(n17510) );
  NAND2X0 U18421 ( .IN1(n17513), .IN2(n17514), .QN(n17512) );
  NAND2X0 U18422 ( .IN1(n17515), .IN2(n17516), .QN(n17514) );
  NOR2X0 U18423 ( .IN1(g311), .IN2(g305), .QN(n17516) );
  AND2X1 U18424 ( .IN1(n5456), .IN2(n5766), .Q(n17515) );
  NAND2X0 U18425 ( .IN1(n17509), .IN2(n17517), .QN(n17513) );
  NAND2X0 U18426 ( .IN1(n17518), .IN2(n5456), .QN(n17517) );
  NOR2X0 U18427 ( .IN1(n17519), .IN2(n17520), .QN(n17518) );
  NOR2X0 U18428 ( .IN1(n5824), .IN2(n5282), .QN(n17520) );
  NOR2X0 U18429 ( .IN1(n5317), .IN2(g336), .QN(n17519) );
  NAND2X0 U18430 ( .IN1(n17521), .IN2(n17522), .QN(g26883) );
  NAND2X0 U18431 ( .IN1(n10499), .IN2(g324), .QN(n17522) );
  NAND2X0 U18432 ( .IN1(n17509), .IN2(n10406), .QN(n17521) );
  NAND2X0 U18433 ( .IN1(n17523), .IN2(n17524), .QN(n17509) );
  NAND2X0 U18434 ( .IN1(n5827), .IN2(g311), .QN(n17524) );
  NAND2X0 U18435 ( .IN1(g305), .IN2(g324), .QN(n17523) );
  NAND2X0 U18436 ( .IN1(n17525), .IN2(n17500), .QN(g26882) );
  NAND2X0 U18437 ( .IN1(n10375), .IN2(g305), .QN(n17500) );
  NOR2X0 U18438 ( .IN1(n17526), .IN2(n17527), .QN(n17525) );
  NOR2X0 U18439 ( .IN1(n9663), .IN2(n10350), .QN(n17527) );
  NOR2X0 U18440 ( .IN1(n5317), .IN2(n10459), .QN(n17526) );
  NAND2X0 U18441 ( .IN1(n17528), .IN2(n17529), .QN(g26881) );
  NAND2X0 U18442 ( .IN1(g6744), .IN2(n10406), .QN(n17529) );
  NAND2X0 U18443 ( .IN1(n10499), .IN2(g305), .QN(n17528) );
  NAND2X0 U18444 ( .IN1(n17530), .IN2(n11282), .QN(g26877) );
  NAND2X0 U18445 ( .IN1(n17531), .IN2(n17532), .QN(n11282) );
  NOR2X0 U18446 ( .IN1(n17533), .IN2(n17534), .QN(n17532) );
  NAND2X0 U18447 ( .IN1(n5311), .IN2(n5310), .QN(n17534) );
  NAND2X0 U18448 ( .IN1(n5276), .IN2(n10140), .QN(n17533) );
  NOR2X0 U18449 ( .IN1(n17535), .IN2(n17536), .QN(n17531) );
  NAND2X0 U18450 ( .IN1(n5620), .IN2(n5619), .QN(n17536) );
  NAND2X0 U18451 ( .IN1(n5406), .IN2(n5405), .QN(n17535) );
  AND2X1 U18452 ( .IN1(n10366), .IN2(n11281), .Q(n17530) );
  NAND2X0 U18453 ( .IN1(n17537), .IN2(n17538), .QN(n11281) );
  NOR2X0 U18454 ( .IN1(n17539), .IN2(n17540), .QN(n17538) );
  NAND2X0 U18455 ( .IN1(n5829), .IN2(n5828), .QN(n17540) );
  NAND2X0 U18456 ( .IN1(n5407), .IN2(n10134), .QN(n17539) );
  NOR2X0 U18457 ( .IN1(n17541), .IN2(n17542), .QN(n17537) );
  NAND2X0 U18458 ( .IN1(n5833), .IN2(n5832), .QN(n17542) );
  NAND2X0 U18459 ( .IN1(n5831), .IN2(n5830), .QN(n17541) );
  NAND2X0 U18460 ( .IN1(n17543), .IN2(n11235), .QN(g26876) );
  NAND2X0 U18461 ( .IN1(n17544), .IN2(n17545), .QN(n11235) );
  NOR2X0 U18462 ( .IN1(n17546), .IN2(n17547), .QN(n17545) );
  NAND2X0 U18463 ( .IN1(n5848), .IN2(n5847), .QN(n17547) );
  NAND2X0 U18464 ( .IN1(n5845), .IN2(n5412), .QN(n17546) );
  NOR2X0 U18465 ( .IN1(n17548), .IN2(n17549), .QN(n17544) );
  NAND2X0 U18466 ( .IN1(n18480), .IN2(n5892), .QN(n17549) );
  NAND2X0 U18467 ( .IN1(n5891), .IN2(n5890), .QN(n17548) );
  NOR2X0 U18468 ( .IN1(n10478), .IN2(n11241), .QN(n17543) );
  INVX0 U18469 ( .INP(n11305), .ZN(n11241) );
  NAND2X0 U18470 ( .IN1(n17550), .IN2(n17551), .QN(n11305) );
  NOR2X0 U18471 ( .IN1(n17552), .IN2(n17553), .QN(n17551) );
  NAND2X0 U18472 ( .IN1(n5411), .IN2(n5410), .QN(n17553) );
  NAND2X0 U18473 ( .IN1(n5278), .IN2(n10153), .QN(n17552) );
  NOR2X0 U18474 ( .IN1(n17554), .IN2(n17555), .QN(n17550) );
  NAND2X0 U18475 ( .IN1(n18481), .IN2(n18482), .QN(n17555) );
  NAND2X0 U18476 ( .IN1(n18483), .IN2(n18484), .QN(n17554) );
  NAND2X0 U18477 ( .IN1(n17556), .IN2(n11310), .QN(g26875) );
  NAND2X0 U18478 ( .IN1(n17557), .IN2(n17558), .QN(n11310) );
  NOR2X0 U18479 ( .IN1(g2523), .IN2(g2657), .QN(n17558) );
  NOR2X0 U18480 ( .IN1(g2255), .IN2(g2389), .QN(n17557) );
  AND2X1 U18481 ( .IN1(n10366), .IN2(n11309), .Q(n17556) );
  NAND2X0 U18482 ( .IN1(n17559), .IN2(n17560), .QN(n11309) );
  NOR2X0 U18483 ( .IN1(g2098), .IN2(g1964), .QN(n17560) );
  AND2X1 U18484 ( .IN1(n5413), .IN2(n5628), .Q(n17559) );
  NAND2X0 U18485 ( .IN1(n17561), .IN2(n17562), .QN(g25764) );
  NAND2X0 U18486 ( .IN1(n17563), .IN2(g6505), .QN(n17562) );
  NAND2X0 U18487 ( .IN1(n14161), .IN2(g6541), .QN(n17561) );
  NAND2X0 U18488 ( .IN1(n17564), .IN2(n17565), .QN(g25763) );
  OR2X1 U18489 ( .IN1(n14161), .IN2(n5884), .Q(n17565) );
  NOR2X0 U18490 ( .IN1(n17566), .IN2(n17567), .QN(n17564) );
  NOR2X0 U18491 ( .IN1(g6533), .IN2(n17568), .QN(n17567) );
  NAND2X0 U18492 ( .IN1(n17569), .IN2(n5659), .QN(n17568) );
  NOR2X0 U18493 ( .IN1(n10478), .IN2(n12631), .QN(n17569) );
  NOR2X0 U18494 ( .IN1(n5445), .IN2(n17570), .QN(n17566) );
  NOR2X0 U18495 ( .IN1(n10478), .IN2(n17571), .QN(n17570) );
  NOR2X0 U18496 ( .IN1(n5659), .IN2(n12631), .QN(n17571) );
  NAND2X0 U18497 ( .IN1(n17572), .IN2(n17573), .QN(g25762) );
  NAND2X0 U18498 ( .IN1(n17563), .IN2(g6533), .QN(n17573) );
  OR2X1 U18499 ( .IN1(n17563), .IN2(n5659), .Q(n17572) );
  NAND2X0 U18500 ( .IN1(n17574), .IN2(n17575), .QN(g25761) );
  NAND2X0 U18501 ( .IN1(n17563), .IN2(g6513), .QN(n17575) );
  INVX0 U18502 ( .INP(n14161), .ZN(n17563) );
  NAND2X0 U18503 ( .IN1(n12631), .IN2(n10406), .QN(n14161) );
  NOR2X0 U18504 ( .IN1(n17576), .IN2(n17577), .QN(n17574) );
  NOR2X0 U18505 ( .IN1(n9665), .IN2(n10351), .QN(n17577) );
  NOR2X0 U18506 ( .IN1(n10478), .IN2(n17578), .QN(n17576) );
  OR2X1 U18507 ( .IN1(g6513), .IN2(n12631), .Q(n17578) );
  NAND2X0 U18508 ( .IN1(n14181), .IN2(g6561), .QN(n12631) );
  INVX0 U18509 ( .INP(n3776), .ZN(n14181) );
  NAND2X0 U18510 ( .IN1(g6573), .IN2(g6565), .QN(n3776) );
  NAND2X0 U18511 ( .IN1(n17579), .IN2(n17580), .QN(g25758) );
  NAND2X0 U18512 ( .IN1(n10505), .IN2(g6494), .QN(n17580) );
  NAND2X0 U18513 ( .IN1(n17581), .IN2(n10406), .QN(n17579) );
  NOR2X0 U18514 ( .IN1(n17582), .IN2(g9817), .QN(n17581) );
  NOR2X0 U18515 ( .IN1(n17583), .IN2(g6444), .QN(n17582) );
  NOR2X0 U18516 ( .IN1(n5719), .IN2(g6494), .QN(n17583) );
  NAND2X0 U18517 ( .IN1(n17584), .IN2(n17585), .QN(g25757) );
  NAND2X0 U18518 ( .IN1(n10374), .IN2(g6727), .QN(n17585) );
  NAND2X0 U18519 ( .IN1(n10505), .IN2(g6444), .QN(n17584) );
  NOR2X0 U18520 ( .IN1(n10478), .IN2(n5563), .QN(g25756) );
  NAND2X0 U18521 ( .IN1(n17586), .IN2(n17587), .QN(g25750) );
  NAND2X0 U18522 ( .IN1(n17588), .IN2(g6159), .QN(n17587) );
  NAND2X0 U18523 ( .IN1(n14281), .IN2(g6195), .QN(n17586) );
  NAND2X0 U18524 ( .IN1(n17589), .IN2(n17590), .QN(g25749) );
  NAND2X0 U18525 ( .IN1(n17588), .IN2(g6191), .QN(n17590) );
  NOR2X0 U18526 ( .IN1(n17591), .IN2(n17592), .QN(n17589) );
  NOR2X0 U18527 ( .IN1(g6187), .IN2(n17593), .QN(n17592) );
  NAND2X0 U18528 ( .IN1(n17594), .IN2(n5667), .QN(n17593) );
  NOR2X0 U18529 ( .IN1(n10478), .IN2(n12624), .QN(n17594) );
  NOR2X0 U18530 ( .IN1(n5453), .IN2(n17595), .QN(n17591) );
  NOR2X0 U18531 ( .IN1(n10478), .IN2(n17596), .QN(n17595) );
  NOR2X0 U18532 ( .IN1(n5667), .IN2(n12624), .QN(n17596) );
  NAND2X0 U18533 ( .IN1(n17597), .IN2(n17598), .QN(g25748) );
  NAND2X0 U18534 ( .IN1(n17588), .IN2(g6187), .QN(n17598) );
  OR2X1 U18535 ( .IN1(n17588), .IN2(n5667), .Q(n17597) );
  NAND2X0 U18536 ( .IN1(n17599), .IN2(n17600), .QN(g25747) );
  NAND2X0 U18537 ( .IN1(n17588), .IN2(g6167), .QN(n17600) );
  INVX0 U18538 ( .INP(n14281), .ZN(n17588) );
  NAND2X0 U18539 ( .IN1(n12624), .IN2(n10405), .QN(n14281) );
  NOR2X0 U18540 ( .IN1(n17601), .IN2(n17602), .QN(n17599) );
  NOR2X0 U18541 ( .IN1(n9645), .IN2(n10351), .QN(n17602) );
  NOR2X0 U18542 ( .IN1(n10478), .IN2(n17603), .QN(n17601) );
  OR2X1 U18543 ( .IN1(g6167), .IN2(n12624), .Q(n17603) );
  NAND2X0 U18544 ( .IN1(n14301), .IN2(g6215), .QN(n12624) );
  INVX0 U18545 ( .INP(n3810), .ZN(n14301) );
  NAND2X0 U18546 ( .IN1(g6227), .IN2(g6219), .QN(n3810) );
  NAND2X0 U18547 ( .IN1(n17604), .IN2(n17605), .QN(g25744) );
  NAND2X0 U18548 ( .IN1(n10505), .IN2(g6148), .QN(n17605) );
  NAND2X0 U18549 ( .IN1(n17606), .IN2(n10405), .QN(n17604) );
  NOR2X0 U18550 ( .IN1(n17607), .IN2(g9741), .QN(n17606) );
  NOR2X0 U18551 ( .IN1(n17608), .IN2(g6098), .QN(n17607) );
  NOR2X0 U18552 ( .IN1(g6148), .IN2(n5718), .QN(n17608) );
  NAND2X0 U18553 ( .IN1(n17609), .IN2(n17610), .QN(g25743) );
  NAND2X0 U18554 ( .IN1(test_so69), .IN2(n10405), .QN(n17610) );
  NAND2X0 U18555 ( .IN1(n10505), .IN2(g6098), .QN(n17609) );
  NOR2X0 U18556 ( .IN1(n10478), .IN2(n5568), .QN(g25742) );
  NAND2X0 U18557 ( .IN1(n17611), .IN2(n17612), .QN(g25736) );
  NAND2X0 U18558 ( .IN1(n14402), .IN2(g5813), .QN(n17612) );
  NAND2X0 U18559 ( .IN1(n15655), .IN2(g5849), .QN(n17611) );
  NAND2X0 U18560 ( .IN1(n17613), .IN2(n17614), .QN(g25735) );
  NAND2X0 U18561 ( .IN1(test_so83), .IN2(n14402), .QN(n17614) );
  NOR2X0 U18562 ( .IN1(n17615), .IN2(n17616), .QN(n17613) );
  NOR2X0 U18563 ( .IN1(g5841), .IN2(n17617), .QN(n17616) );
  NAND2X0 U18564 ( .IN1(n17618), .IN2(n5663), .QN(n17617) );
  NOR2X0 U18565 ( .IN1(n10478), .IN2(n12623), .QN(n17618) );
  NOR2X0 U18566 ( .IN1(n5449), .IN2(n17619), .QN(n17615) );
  NOR2X0 U18567 ( .IN1(n10478), .IN2(n17620), .QN(n17619) );
  NOR2X0 U18568 ( .IN1(n5663), .IN2(n12623), .QN(n17620) );
  NAND2X0 U18569 ( .IN1(n17621), .IN2(n17622), .QN(g25734) );
  NAND2X0 U18570 ( .IN1(n14402), .IN2(g5841), .QN(n17622) );
  OR2X1 U18571 ( .IN1(n14402), .IN2(n5663), .Q(n17621) );
  NAND2X0 U18572 ( .IN1(n17623), .IN2(n17624), .QN(g25733) );
  NAND2X0 U18573 ( .IN1(n14402), .IN2(g5821), .QN(n17624) );
  INVX0 U18574 ( .INP(n15655), .ZN(n14402) );
  NAND2X0 U18575 ( .IN1(n12623), .IN2(n10405), .QN(n15655) );
  NOR2X0 U18576 ( .IN1(n17625), .IN2(n17626), .QN(n17623) );
  NOR2X0 U18577 ( .IN1(n9618), .IN2(n10351), .QN(n17626) );
  NOR2X0 U18578 ( .IN1(n10478), .IN2(n17627), .QN(n17625) );
  OR2X1 U18579 ( .IN1(g5821), .IN2(n12623), .Q(n17627) );
  NAND2X0 U18580 ( .IN1(n14422), .IN2(g5869), .QN(n12623) );
  INVX0 U18581 ( .INP(n3844), .ZN(n14422) );
  NAND2X0 U18582 ( .IN1(test_so36), .IN2(g5873), .QN(n3844) );
  NAND2X0 U18583 ( .IN1(n17628), .IN2(n17629), .QN(g25730) );
  NAND2X0 U18584 ( .IN1(n10505), .IN2(g5802), .QN(n17629) );
  NAND2X0 U18585 ( .IN1(n17630), .IN2(n10405), .QN(n17628) );
  NOR2X0 U18586 ( .IN1(n17631), .IN2(g9680), .QN(n17630) );
  NOR2X0 U18587 ( .IN1(n17632), .IN2(g5752), .QN(n17631) );
  NOR2X0 U18588 ( .IN1(n5722), .IN2(g5802), .QN(n17632) );
  NAND2X0 U18589 ( .IN1(n17633), .IN2(n17634), .QN(g25729) );
  NAND2X0 U18590 ( .IN1(n10373), .IN2(g6035), .QN(n17634) );
  NAND2X0 U18591 ( .IN1(n10505), .IN2(g5752), .QN(n17633) );
  NOR2X0 U18592 ( .IN1(n10139), .IN2(n10460), .QN(g25728) );
  NAND2X0 U18593 ( .IN1(n17635), .IN2(n17636), .QN(g25722) );
  NAND2X0 U18594 ( .IN1(n17637), .IN2(g5467), .QN(n17636) );
  NAND2X0 U18595 ( .IN1(n14524), .IN2(g5503), .QN(n17635) );
  NAND2X0 U18596 ( .IN1(n17638), .IN2(n17639), .QN(g25721) );
  OR2X1 U18597 ( .IN1(n14524), .IN2(n5885), .Q(n17639) );
  NOR2X0 U18598 ( .IN1(n17640), .IN2(n17641), .QN(n17638) );
  NOR2X0 U18599 ( .IN1(g5495), .IN2(n17642), .QN(n17641) );
  NAND2X0 U18600 ( .IN1(n17643), .IN2(n5660), .QN(n17642) );
  NOR2X0 U18601 ( .IN1(n10477), .IN2(n14523), .QN(n17643) );
  NOR2X0 U18602 ( .IN1(n5446), .IN2(n17644), .QN(n17640) );
  NOR2X0 U18603 ( .IN1(n10477), .IN2(n17645), .QN(n17644) );
  NOR2X0 U18604 ( .IN1(n5660), .IN2(n14523), .QN(n17645) );
  NAND2X0 U18605 ( .IN1(n17646), .IN2(n17647), .QN(g25720) );
  NAND2X0 U18606 ( .IN1(n17637), .IN2(g5495), .QN(n17647) );
  OR2X1 U18607 ( .IN1(n17637), .IN2(n5660), .Q(n17646) );
  NAND2X0 U18608 ( .IN1(n17648), .IN2(n17649), .QN(g25719) );
  NAND2X0 U18609 ( .IN1(n17637), .IN2(g5475), .QN(n17649) );
  INVX0 U18610 ( .INP(n14524), .ZN(n17637) );
  NAND2X0 U18611 ( .IN1(n14523), .IN2(n10405), .QN(n14524) );
  NOR2X0 U18612 ( .IN1(n17650), .IN2(n17651), .QN(n17648) );
  NOR2X0 U18613 ( .IN1(n9627), .IN2(n10351), .QN(n17651) );
  NOR2X0 U18614 ( .IN1(n10477), .IN2(n17652), .QN(n17650) );
  NAND2X0 U18615 ( .IN1(n5425), .IN2(n12614), .QN(n17652) );
  INVX0 U18616 ( .INP(n14523), .ZN(n12614) );
  NAND2X0 U18617 ( .IN1(n14546), .IN2(g5523), .QN(n14523) );
  INVX0 U18618 ( .INP(n3877), .ZN(n14546) );
  NAND2X0 U18619 ( .IN1(g5535), .IN2(g5527), .QN(n3877) );
  NAND2X0 U18620 ( .IN1(n17653), .IN2(n17654), .QN(g25716) );
  NAND2X0 U18621 ( .IN1(n10504), .IN2(g5456), .QN(n17654) );
  NAND2X0 U18622 ( .IN1(n17655), .IN2(n10405), .QN(n17653) );
  NOR2X0 U18623 ( .IN1(test_so35), .IN2(n17656), .QN(n17655) );
  NOR2X0 U18624 ( .IN1(n17657), .IN2(g5406), .QN(n17656) );
  NOR2X0 U18625 ( .IN1(n18468), .IN2(g5456), .QN(n17657) );
  NAND2X0 U18626 ( .IN1(n17658), .IN2(n17659), .QN(g25715) );
  NAND2X0 U18627 ( .IN1(n10373), .IN2(g5689), .QN(n17659) );
  NAND2X0 U18628 ( .IN1(n10504), .IN2(g5406), .QN(n17658) );
  NOR2X0 U18629 ( .IN1(n10477), .IN2(n5566), .QN(g25714) );
  NAND2X0 U18630 ( .IN1(n17660), .IN2(n17661), .QN(g25708) );
  NAND2X0 U18631 ( .IN1(n17662), .IN2(g5120), .QN(n17661) );
  NAND2X0 U18632 ( .IN1(n14645), .IN2(g5156), .QN(n17660) );
  NAND2X0 U18633 ( .IN1(n17663), .IN2(n17664), .QN(g25707) );
  OR2X1 U18634 ( .IN1(n14645), .IN2(n5883), .Q(n17664) );
  NOR2X0 U18635 ( .IN1(n17665), .IN2(n17666), .QN(n17663) );
  NOR2X0 U18636 ( .IN1(test_so98), .IN2(n17667), .QN(n17666) );
  NAND2X0 U18637 ( .IN1(n17668), .IN2(n5658), .QN(n17667) );
  NOR2X0 U18638 ( .IN1(n10477), .IN2(n12619), .QN(n17668) );
  NOR2X0 U18639 ( .IN1(n17669), .IN2(n10159), .QN(n17665) );
  NOR2X0 U18640 ( .IN1(n10477), .IN2(n17670), .QN(n17669) );
  NOR2X0 U18641 ( .IN1(n5658), .IN2(n12619), .QN(n17670) );
  NAND2X0 U18642 ( .IN1(n17671), .IN2(n17672), .QN(g25706) );
  NAND2X0 U18643 ( .IN1(test_so98), .IN2(n17662), .QN(n17672) );
  OR2X1 U18644 ( .IN1(n17662), .IN2(n5658), .Q(n17671) );
  NAND2X0 U18645 ( .IN1(n17673), .IN2(n17674), .QN(g25705) );
  NAND2X0 U18646 ( .IN1(test_so96), .IN2(n17662), .QN(n17674) );
  INVX0 U18647 ( .INP(n14645), .ZN(n17662) );
  NAND2X0 U18648 ( .IN1(n12619), .IN2(n10405), .QN(n14645) );
  NOR2X0 U18649 ( .IN1(n17675), .IN2(n17676), .QN(n17673) );
  NOR2X0 U18650 ( .IN1(n9616), .IN2(n10351), .QN(n17676) );
  NOR2X0 U18651 ( .IN1(n10477), .IN2(n17677), .QN(n17675) );
  NAND2X0 U18652 ( .IN1(g32975), .IN2(n10141), .QN(n17677) );
  INVX0 U18653 ( .INP(n12619), .ZN(g32975) );
  NAND2X0 U18654 ( .IN1(n14665), .IN2(g5176), .QN(n12619) );
  INVX0 U18655 ( .INP(n3910), .ZN(n14665) );
  NAND2X0 U18656 ( .IN1(g5188), .IN2(g5180), .QN(n3910) );
  NOR2X0 U18657 ( .IN1(n9689), .IN2(n17678), .QN(g25704) );
  NOR2X0 U18658 ( .IN1(n10477), .IN2(g5069), .QN(n17678) );
  NAND2X0 U18659 ( .IN1(n17679), .IN2(n17680), .QN(g25703) );
  NAND2X0 U18660 ( .IN1(n10504), .IN2(g5112), .QN(n17680) );
  NAND2X0 U18661 ( .IN1(n17681), .IN2(n10405), .QN(n17679) );
  NOR2X0 U18662 ( .IN1(n17682), .IN2(g9497), .QN(n17681) );
  NOR2X0 U18663 ( .IN1(n17683), .IN2(g5022), .QN(n17682) );
  NOR2X0 U18664 ( .IN1(n5690), .IN2(g5112), .QN(n17683) );
  NAND2X0 U18665 ( .IN1(n17684), .IN2(n17685), .QN(g25702) );
  NAND2X0 U18666 ( .IN1(test_so32), .IN2(n10516), .QN(n17685) );
  NAND2X0 U18667 ( .IN1(n17686), .IN2(n10404), .QN(n17684) );
  NOR2X0 U18668 ( .IN1(n17687), .IN2(g9553), .QN(n17686) );
  NOR2X0 U18669 ( .IN1(n17688), .IN2(g5062), .QN(n17687) );
  NOR2X0 U18670 ( .IN1(test_so32), .IN2(n5689), .QN(n17688) );
  NAND2X0 U18671 ( .IN1(n17689), .IN2(n17690), .QN(g25701) );
  NAND2X0 U18672 ( .IN1(test_so10), .IN2(n10404), .QN(n17690) );
  NAND2X0 U18673 ( .IN1(n10504), .IN2(g5062), .QN(n17689) );
  NOR2X0 U18674 ( .IN1(n10477), .IN2(n5567), .QN(g25700) );
  NAND2X0 U18675 ( .IN1(n17691), .IN2(n17692), .QN(g25699) );
  NAND2X0 U18676 ( .IN1(n10504), .IN2(g5097), .QN(n17692) );
  NOR2X0 U18677 ( .IN1(n17693), .IN2(n17694), .QN(n17691) );
  AND2X1 U18678 ( .IN1(n5669), .IN2(n5014), .Q(n17694) );
  NOR2X0 U18679 ( .IN1(n5669), .IN2(n17695), .QN(n17693) );
  OR2X1 U18680 ( .IN1(n10457), .IN2(n5014), .Q(n17695) );
  NAND2X0 U18681 ( .IN1(n17696), .IN2(n17697), .QN(g25698) );
  NAND2X0 U18682 ( .IN1(n10504), .IN2(g5092), .QN(n17697) );
  NOR2X0 U18683 ( .IN1(n17698), .IN2(n17699), .QN(n17696) );
  NOR2X0 U18684 ( .IN1(g5097), .IN2(n17700), .QN(n17699) );
  NOR2X0 U18685 ( .IN1(n5753), .IN2(n17701), .QN(n17698) );
  NAND2X0 U18686 ( .IN1(n10372), .IN2(n17700), .QN(n17701) );
  INVX0 U18687 ( .INP(n5016), .ZN(n17700) );
  XOR2X1 U18688 ( .IN1(n17702), .IN2(n5681), .Q(g25697) );
  NAND2X0 U18689 ( .IN1(n10372), .IN2(g5092), .QN(n17702) );
  NAND2X0 U18690 ( .IN1(n17703), .IN2(n17704), .QN(g25696) );
  NAND2X0 U18691 ( .IN1(n17705), .IN2(n9689), .QN(n17704) );
  NOR2X0 U18692 ( .IN1(n5455), .IN2(n10461), .QN(n17705) );
  NOR2X0 U18693 ( .IN1(n17706), .IN2(n17707), .QN(n17703) );
  NOR2X0 U18694 ( .IN1(g5080), .IN2(n17708), .QN(n17707) );
  NAND2X0 U18695 ( .IN1(n17709), .IN2(n17710), .QN(n17708) );
  OR2X1 U18696 ( .IN1(g5069), .IN2(n5455), .Q(n17710) );
  NOR2X0 U18697 ( .IN1(n5893), .IN2(n17709), .QN(n17706) );
  NOR2X0 U18698 ( .IN1(g5084), .IN2(n10461), .QN(n17709) );
  NOR2X0 U18699 ( .IN1(n5455), .IN2(n17711), .QN(g25695) );
  NOR2X0 U18700 ( .IN1(n10477), .IN2(n17712), .QN(n17711) );
  NAND2X0 U18701 ( .IN1(n17713), .IN2(n17714), .QN(n17712) );
  NAND2X0 U18702 ( .IN1(n9688), .IN2(g5084), .QN(n17714) );
  NAND2X0 U18703 ( .IN1(n9689), .IN2(n5681), .QN(n17713) );
  NAND2X0 U18704 ( .IN1(n17715), .IN2(n17716), .QN(g25691) );
  NAND2X0 U18705 ( .IN1(n10114), .IN2(n17717), .QN(n17716) );
  NAND2X0 U18706 ( .IN1(n17718), .IN2(n17719), .QN(n17717) );
  NOR2X0 U18707 ( .IN1(n17720), .IN2(n17721), .QN(n17719) );
  NAND2X0 U18708 ( .IN1(test_so11), .IN2(n9739), .QN(n17721) );
  NAND2X0 U18709 ( .IN1(n5612), .IN2(g4098), .QN(n17720) );
  NOR2X0 U18710 ( .IN1(g4057), .IN2(n17722), .QN(n17718) );
  NAND2X0 U18711 ( .IN1(n5416), .IN2(n12615), .QN(n17722) );
  INVX0 U18712 ( .INP(n14779), .ZN(n12615) );
  NAND2X0 U18713 ( .IN1(n5340), .IN2(g4087), .QN(n14779) );
  INVX0 U18714 ( .INP(n14067), .ZN(n10114) );
  NAND2X0 U18715 ( .IN1(n10504), .IN2(g4125), .QN(n17715) );
  NAND2X0 U18716 ( .IN1(n17723), .IN2(n17724), .QN(g25690) );
  NAND2X0 U18717 ( .IN1(n10504), .IN2(g4169), .QN(n17724) );
  NAND2X0 U18718 ( .IN1(n17725), .IN2(n10404), .QN(n17723) );
  NOR2X0 U18719 ( .IN1(n9621), .IN2(g4125), .QN(n17725) );
  NAND2X0 U18720 ( .IN1(n17726), .IN2(n17727), .QN(g25687) );
  NAND2X0 U18721 ( .IN1(n10504), .IN2(g4057), .QN(n17727) );
  NOR2X0 U18722 ( .IN1(n17728), .IN2(n17729), .QN(n17726) );
  AND2X1 U18723 ( .IN1(n5026), .IN2(n14778), .Q(n17729) );
  NOR2X0 U18724 ( .IN1(g4141), .IN2(n17730), .QN(n17728) );
  NAND2X0 U18725 ( .IN1(n17250), .IN2(g4169), .QN(n17730) );
  INVX0 U18726 ( .INP(n4723), .ZN(n17250) );
  NAND2X0 U18727 ( .IN1(g4057), .IN2(g4064), .QN(n4723) );
  NAND2X0 U18728 ( .IN1(n17731), .IN2(n17732), .QN(g25686) );
  NAND2X0 U18729 ( .IN1(n17733), .IN2(g4064), .QN(n17732) );
  NAND2X0 U18730 ( .IN1(n17734), .IN2(n10404), .QN(n17733) );
  NAND2X0 U18731 ( .IN1(n5711), .IN2(g4169), .QN(n17734) );
  NAND2X0 U18732 ( .IN1(n17735), .IN2(n5416), .QN(n17731) );
  AND2X1 U18733 ( .IN1(g4057), .IN2(n14778), .Q(n17735) );
  NOR2X0 U18734 ( .IN1(n10477), .IN2(n5729), .QN(n14778) );
  NAND2X0 U18735 ( .IN1(n17736), .IN2(n14067), .QN(g25685) );
  NAND2X0 U18736 ( .IN1(n5729), .IN2(n10404), .QN(n14067) );
  NOR2X0 U18737 ( .IN1(n17737), .IN2(n17738), .QN(n17736) );
  NOR2X0 U18738 ( .IN1(n10093), .IN2(n10352), .QN(n17738) );
  NOR2X0 U18739 ( .IN1(n10477), .IN2(g4064), .QN(n17737) );
  NAND2X0 U18740 ( .IN1(n17739), .IN2(n17740), .QN(g25684) );
  NAND2X0 U18741 ( .IN1(n17741), .IN2(g3813), .QN(n17740) );
  NAND2X0 U18742 ( .IN1(n14785), .IN2(g3849), .QN(n17739) );
  NAND2X0 U18743 ( .IN1(n17742), .IN2(n17743), .QN(g25683) );
  OR2X1 U18744 ( .IN1(n14785), .IN2(n5886), .Q(n17743) );
  NOR2X0 U18745 ( .IN1(n17744), .IN2(n17745), .QN(n17742) );
  NOR2X0 U18746 ( .IN1(test_so97), .IN2(n17746), .QN(n17745) );
  NAND2X0 U18747 ( .IN1(n17747), .IN2(n5662), .QN(n17746) );
  NOR2X0 U18748 ( .IN1(n10477), .IN2(n12636), .QN(n17747) );
  NOR2X0 U18749 ( .IN1(n17748), .IN2(n10160), .QN(n17744) );
  NOR2X0 U18750 ( .IN1(n10477), .IN2(n17749), .QN(n17748) );
  NOR2X0 U18751 ( .IN1(n5662), .IN2(n12636), .QN(n17749) );
  NAND2X0 U18752 ( .IN1(n17750), .IN2(n17751), .QN(g25682) );
  NAND2X0 U18753 ( .IN1(test_so97), .IN2(n17741), .QN(n17751) );
  OR2X1 U18754 ( .IN1(n17741), .IN2(n5662), .Q(n17750) );
  NAND2X0 U18755 ( .IN1(n17752), .IN2(n17753), .QN(g25681) );
  NAND2X0 U18756 ( .IN1(n17741), .IN2(g3821), .QN(n17753) );
  INVX0 U18757 ( .INP(n14785), .ZN(n17741) );
  NAND2X0 U18758 ( .IN1(n12636), .IN2(n10404), .QN(n14785) );
  NOR2X0 U18759 ( .IN1(n17754), .IN2(n17755), .QN(n17752) );
  NOR2X0 U18760 ( .IN1(n9617), .IN2(n10352), .QN(n17755) );
  NOR2X0 U18761 ( .IN1(n10476), .IN2(n17756), .QN(n17754) );
  OR2X1 U18762 ( .IN1(g3821), .IN2(n12636), .Q(n17756) );
  NAND2X0 U18763 ( .IN1(test_so33), .IN2(n14808), .QN(n12636) );
  INVX0 U18764 ( .INP(n3953), .ZN(n14808) );
  NAND2X0 U18765 ( .IN1(g3881), .IN2(g3873), .QN(n3953) );
  NAND2X0 U18766 ( .IN1(n17757), .IN2(n17758), .QN(g25678) );
  NAND2X0 U18767 ( .IN1(n10503), .IN2(g3802), .QN(n17758) );
  NAND2X0 U18768 ( .IN1(n17759), .IN2(n10404), .QN(n17757) );
  NOR2X0 U18769 ( .IN1(n17760), .IN2(g8398), .QN(n17759) );
  NOR2X0 U18770 ( .IN1(n17761), .IN2(g3752), .QN(n17760) );
  NOR2X0 U18771 ( .IN1(n5721), .IN2(g3802), .QN(n17761) );
  NAND2X0 U18772 ( .IN1(n17762), .IN2(n17763), .QN(g25677) );
  NAND2X0 U18773 ( .IN1(n10371), .IN2(g4040), .QN(n17763) );
  NAND2X0 U18774 ( .IN1(n10503), .IN2(g3752), .QN(n17762) );
  INVX0 U18775 ( .INP(n13547), .ZN(g25676) );
  NAND2X0 U18776 ( .IN1(n10371), .IN2(g3881), .QN(n13547) );
  NAND2X0 U18777 ( .IN1(n17764), .IN2(n17765), .QN(g25670) );
  NAND2X0 U18778 ( .IN1(n17766), .IN2(g3462), .QN(n17765) );
  NAND2X0 U18779 ( .IN1(n14906), .IN2(g3498), .QN(n17764) );
  NAND2X0 U18780 ( .IN1(n17767), .IN2(n17768), .QN(g25669) );
  OR2X1 U18781 ( .IN1(n14906), .IN2(n5889), .Q(n17768) );
  NOR2X0 U18782 ( .IN1(n17769), .IN2(n17770), .QN(n17767) );
  NOR2X0 U18783 ( .IN1(g3490), .IN2(n17771), .QN(n17770) );
  NAND2X0 U18784 ( .IN1(n17772), .IN2(n5668), .QN(n17771) );
  NOR2X0 U18785 ( .IN1(n10476), .IN2(n12635), .QN(n17772) );
  NOR2X0 U18786 ( .IN1(n5454), .IN2(n17773), .QN(n17769) );
  NOR2X0 U18787 ( .IN1(n10476), .IN2(n17774), .QN(n17773) );
  NOR2X0 U18788 ( .IN1(n5668), .IN2(n12635), .QN(n17774) );
  NAND2X0 U18789 ( .IN1(n17775), .IN2(n17776), .QN(g25668) );
  NAND2X0 U18790 ( .IN1(n17766), .IN2(g3490), .QN(n17776) );
  OR2X1 U18791 ( .IN1(n17766), .IN2(n5668), .Q(n17775) );
  NAND2X0 U18792 ( .IN1(n17777), .IN2(n17778), .QN(g25667) );
  NAND2X0 U18793 ( .IN1(n17766), .IN2(g3470), .QN(n17778) );
  INVX0 U18794 ( .INP(n14906), .ZN(n17766) );
  NAND2X0 U18795 ( .IN1(n12635), .IN2(n10404), .QN(n14906) );
  NOR2X0 U18796 ( .IN1(n17779), .IN2(n17780), .QN(n17777) );
  NOR2X0 U18797 ( .IN1(n9639), .IN2(n10351), .QN(n17780) );
  NOR2X0 U18798 ( .IN1(n10476), .IN2(n17781), .QN(n17779) );
  OR2X1 U18799 ( .IN1(g3470), .IN2(n12635), .Q(n17781) );
  NAND2X0 U18800 ( .IN1(n14926), .IN2(g3518), .QN(n12635) );
  INVX0 U18801 ( .INP(n3986), .ZN(n14926) );
  NAND2X0 U18802 ( .IN1(g3530), .IN2(g3522), .QN(n3986) );
  NAND2X0 U18803 ( .IN1(n17782), .IN2(n17783), .QN(g25664) );
  NAND2X0 U18804 ( .IN1(n10503), .IN2(g3451), .QN(n17783) );
  NAND2X0 U18805 ( .IN1(n17784), .IN2(n10404), .QN(n17782) );
  NOR2X0 U18806 ( .IN1(n17785), .IN2(g8342), .QN(n17784) );
  NOR2X0 U18807 ( .IN1(n17786), .IN2(g3401), .QN(n17785) );
  NOR2X0 U18808 ( .IN1(n5717), .IN2(g3451), .QN(n17786) );
  NAND2X0 U18809 ( .IN1(n17787), .IN2(n17788), .QN(g25663) );
  NAND2X0 U18810 ( .IN1(n10371), .IN2(g3689), .QN(n17788) );
  NAND2X0 U18811 ( .IN1(n10503), .IN2(g3401), .QN(n17787) );
  NOR2X0 U18812 ( .IN1(n10476), .IN2(n5569), .QN(g25662) );
  NAND2X0 U18813 ( .IN1(n17789), .IN2(n17790), .QN(g25656) );
  NAND2X0 U18814 ( .IN1(n17791), .IN2(g3111), .QN(n17790) );
  NAND2X0 U18815 ( .IN1(n15027), .IN2(g3147), .QN(n17789) );
  NAND2X0 U18816 ( .IN1(n17792), .IN2(n17793), .QN(g25655) );
  NAND2X0 U18817 ( .IN1(n17791), .IN2(g3143), .QN(n17793) );
  NOR2X0 U18818 ( .IN1(n17794), .IN2(n17795), .QN(n17792) );
  NOR2X0 U18819 ( .IN1(g3139), .IN2(n17796), .QN(n17795) );
  NAND2X0 U18820 ( .IN1(n17797), .IN2(n5661), .QN(n17796) );
  NOR2X0 U18821 ( .IN1(n10476), .IN2(n15026), .QN(n17797) );
  NOR2X0 U18822 ( .IN1(n5447), .IN2(n17798), .QN(n17794) );
  NOR2X0 U18823 ( .IN1(n10476), .IN2(n17799), .QN(n17798) );
  NOR2X0 U18824 ( .IN1(n5661), .IN2(n15026), .QN(n17799) );
  NAND2X0 U18825 ( .IN1(n17800), .IN2(n17801), .QN(g25654) );
  NAND2X0 U18826 ( .IN1(n17791), .IN2(g3139), .QN(n17801) );
  OR2X1 U18827 ( .IN1(n17791), .IN2(n5661), .Q(n17800) );
  NAND2X0 U18828 ( .IN1(n17802), .IN2(n17803), .QN(g25653) );
  NAND2X0 U18829 ( .IN1(n17791), .IN2(g3119), .QN(n17803) );
  INVX0 U18830 ( .INP(n15027), .ZN(n17791) );
  NAND2X0 U18831 ( .IN1(n15026), .IN2(n10404), .QN(n15027) );
  NOR2X0 U18832 ( .IN1(n17804), .IN2(n17805), .QN(n17802) );
  NOR2X0 U18833 ( .IN1(n9664), .IN2(n10352), .QN(n17805) );
  NOR2X0 U18834 ( .IN1(n10476), .IN2(n17806), .QN(n17804) );
  NAND2X0 U18835 ( .IN1(n5423), .IN2(n12628), .QN(n17806) );
  INVX0 U18836 ( .INP(n15026), .ZN(n12628) );
  NAND2X0 U18837 ( .IN1(n15048), .IN2(g3167), .QN(n15026) );
  INVX0 U18838 ( .INP(n365), .ZN(n15048) );
  NAND2X0 U18839 ( .IN1(g3179), .IN2(g3171), .QN(n365) );
  NAND2X0 U18840 ( .IN1(n17807), .IN2(n17808), .QN(g25650) );
  NAND2X0 U18841 ( .IN1(n10503), .IN2(g3100), .QN(n17808) );
  NAND2X0 U18842 ( .IN1(n17809), .IN2(n10403), .QN(n17807) );
  NOR2X0 U18843 ( .IN1(n17810), .IN2(g8277), .QN(n17809) );
  NOR2X0 U18844 ( .IN1(n17811), .IN2(g3050), .QN(n17810) );
  NOR2X0 U18845 ( .IN1(n5723), .IN2(g3100), .QN(n17811) );
  NAND2X0 U18846 ( .IN1(n17812), .IN2(n17813), .QN(g25649) );
  NAND2X0 U18847 ( .IN1(n10371), .IN2(g3338), .QN(n17813) );
  NAND2X0 U18848 ( .IN1(n10503), .IN2(g3050), .QN(n17812) );
  NOR2X0 U18849 ( .IN1(n10476), .IN2(n5390), .QN(g25648) );
  OR2X1 U18850 ( .IN1(n5045), .IN2(n17814), .Q(g25639) );
  NAND2X0 U18851 ( .IN1(n17815), .IN2(n17816), .QN(n17814) );
  NAND2X0 U18852 ( .IN1(n10503), .IN2(g2715), .QN(n17816) );
  NAND2X0 U18853 ( .IN1(n15156), .IN2(n10403), .QN(n17815) );
  NOR2X0 U18854 ( .IN1(g2715), .IN2(n5465), .QN(n15156) );
  NAND2X0 U18855 ( .IN1(n17817), .IN2(n17818), .QN(g25638) );
  NAND2X0 U18856 ( .IN1(n10503), .IN2(g1564), .QN(n17818) );
  NAND2X0 U18857 ( .IN1(n17819), .IN2(n10403), .QN(n17817) );
  NAND2X0 U18858 ( .IN1(n17820), .IN2(n17821), .QN(n17819) );
  NAND2X0 U18859 ( .IN1(n17822), .IN2(g1559), .QN(n17821) );
  NAND2X0 U18860 ( .IN1(n17823), .IN2(n5441), .QN(n17820) );
  NOR2X0 U18861 ( .IN1(g1554), .IN2(n17822), .QN(n17823) );
  NAND2X0 U18862 ( .IN1(n17824), .IN2(n17825), .QN(g25637) );
  NAND2X0 U18863 ( .IN1(n17826), .IN2(n17822), .QN(n17825) );
  NOR2X0 U18864 ( .IN1(n5768), .IN2(n10462), .QN(n17826) );
  NAND2X0 U18865 ( .IN1(n17827), .IN2(g1559), .QN(n17824) );
  NAND2X0 U18866 ( .IN1(n17828), .IN2(n10403), .QN(n17827) );
  OR2X1 U18867 ( .IN1(n17822), .IN2(g1554), .Q(n17828) );
  NAND2X0 U18868 ( .IN1(n17829), .IN2(n17830), .QN(g25636) );
  NAND2X0 U18869 ( .IN1(n10503), .IN2(g1521), .QN(n17830) );
  NAND2X0 U18870 ( .IN1(n17831), .IN2(n10403), .QN(n17829) );
  NAND2X0 U18871 ( .IN1(n17832), .IN2(n17833), .QN(n17831) );
  OR2X1 U18872 ( .IN1(n17834), .IN2(n5381), .Q(n17833) );
  NAND2X0 U18873 ( .IN1(n17834), .IN2(g1306), .QN(n17832) );
  NAND2X0 U18874 ( .IN1(n17835), .IN2(test_so49), .QN(n17834) );
  NOR2X0 U18875 ( .IN1(n5364), .IN2(n5302), .QN(n17835) );
  NAND2X0 U18876 ( .IN1(n17836), .IN2(n17837), .QN(g25635) );
  NAND2X0 U18877 ( .IN1(n17838), .IN2(g1484), .QN(n17837) );
  NAND2X0 U18878 ( .IN1(n17839), .IN2(n10403), .QN(n17838) );
  NAND2X0 U18879 ( .IN1(n17840), .IN2(n17314), .QN(n17839) );
  NOR2X0 U18880 ( .IN1(n17841), .IN2(g1300), .QN(n17840) );
  NAND2X0 U18881 ( .IN1(n17842), .IN2(g1300), .QN(n17836) );
  NAND2X0 U18882 ( .IN1(n17843), .IN2(n17844), .QN(n17842) );
  NAND2X0 U18883 ( .IN1(n17845), .IN2(n10403), .QN(n17844) );
  NAND2X0 U18884 ( .IN1(n17314), .IN2(g1484), .QN(n17845) );
  NOR2X0 U18885 ( .IN1(n10049), .IN2(test_so12), .QN(n17314) );
  NOR2X0 U18886 ( .IN1(n17846), .IN2(n17847), .QN(g25634) );
  NAND2X0 U18887 ( .IN1(n17326), .IN2(n10128), .QN(n17847) );
  NAND2X0 U18888 ( .IN1(n17848), .IN2(n17849), .QN(n17326) );
  NOR2X0 U18889 ( .IN1(n9966), .IN2(n5655), .QN(n17848) );
  NOR2X0 U18890 ( .IN1(n17850), .IN2(n17851), .QN(n17846) );
  NOR2X0 U18891 ( .IN1(n9966), .IN2(n10462), .QN(n17851) );
  NOR2X0 U18892 ( .IN1(n17852), .IN2(n17853), .QN(n17850) );
  NAND2X0 U18893 ( .IN1(n17854), .IN2(n17855), .QN(g25633) );
  OR2X1 U18894 ( .IN1(n10311), .IN2(n9685), .Q(n17855) );
  NAND2X0 U18895 ( .IN1(n17856), .IN2(n10402), .QN(n17854) );
  NAND2X0 U18896 ( .IN1(n17857), .IN2(n17858), .QN(n17856) );
  NAND2X0 U18897 ( .IN1(n17859), .IN2(g1384), .QN(n17858) );
  NAND2X0 U18898 ( .IN1(n17860), .IN2(n9592), .QN(n17857) );
  NOR2X0 U18899 ( .IN1(n5322), .IN2(n17859), .QN(n17860) );
  NAND2X0 U18900 ( .IN1(n17861), .IN2(n17862), .QN(g25632) );
  NAND2X0 U18901 ( .IN1(n17863), .IN2(g1312), .QN(n17862) );
  NAND2X0 U18902 ( .IN1(n17859), .IN2(n10402), .QN(n17863) );
  NAND2X0 U18903 ( .IN1(n17864), .IN2(n17865), .QN(n17861) );
  NOR2X0 U18904 ( .IN1(n5322), .IN2(n10462), .QN(n17865) );
  NOR2X0 U18905 ( .IN1(n17866), .IN2(n17867), .QN(n17864) );
  NOR2X0 U18906 ( .IN1(n9758), .IN2(n17859), .QN(n17867) );
  AND2X1 U18907 ( .IN1(n15501), .IN2(n16992), .Q(n17866) );
  NOR2X0 U18908 ( .IN1(n10476), .IN2(n17868), .QN(g25631) );
  NOR2X0 U18909 ( .IN1(n17869), .IN2(n17870), .QN(n17868) );
  NOR2X0 U18910 ( .IN1(n5466), .IN2(n17332), .QN(n17870) );
  INVX0 U18911 ( .INP(n17859), .ZN(n17332) );
  NOR2X0 U18912 ( .IN1(n16995), .IN2(n17871), .QN(n17869) );
  NAND2X0 U18913 ( .IN1(n17872), .IN2(n17873), .QN(n17871) );
  NAND2X0 U18914 ( .IN1(n5322), .IN2(n4896), .QN(n17873) );
  NAND2X0 U18915 ( .IN1(n17874), .IN2(n17875), .QN(n4896) );
  NOR2X0 U18916 ( .IN1(n9750), .IN2(n9727), .QN(n17875) );
  NOR2X0 U18917 ( .IN1(n9685), .IN2(n16990), .QN(n17874) );
  NAND2X0 U18918 ( .IN1(n17876), .IN2(g1351), .QN(n17872) );
  NAND2X0 U18919 ( .IN1(n16992), .IN2(n17877), .QN(n17876) );
  INVX0 U18920 ( .INP(n16994), .ZN(n17877) );
  NOR2X0 U18921 ( .IN1(n16993), .IN2(n9758), .QN(n16994) );
  NOR2X0 U18922 ( .IN1(n9761), .IN2(n9762), .QN(n16992) );
  INVX0 U18923 ( .INP(n15501), .ZN(n16995) );
  NAND2X0 U18924 ( .IN1(n17878), .IN2(n17879), .QN(g25630) );
  NAND2X0 U18925 ( .IN1(n17880), .IN2(g1249), .QN(n17879) );
  NAND2X0 U18926 ( .IN1(n17881), .IN2(n10401), .QN(n17880) );
  NAND2X0 U18927 ( .IN1(n9743), .IN2(g12923), .QN(n17881) );
  NAND2X0 U18928 ( .IN1(g24247), .IN2(g1266), .QN(n17878) );
  NAND2X0 U18929 ( .IN1(n17882), .IN2(n17883), .QN(g25629) );
  NAND2X0 U18930 ( .IN1(n10502), .IN2(g1221), .QN(n17883) );
  NAND2X0 U18931 ( .IN1(n17884), .IN2(n10401), .QN(n17882) );
  NAND2X0 U18932 ( .IN1(n17885), .IN2(n17886), .QN(n17884) );
  NAND2X0 U18933 ( .IN1(n17887), .IN2(g1216), .QN(n17886) );
  NAND2X0 U18934 ( .IN1(n17888), .IN2(n5442), .QN(n17885) );
  NOR2X0 U18935 ( .IN1(test_so76), .IN2(n17887), .QN(n17888) );
  NAND2X0 U18936 ( .IN1(n17889), .IN2(n17890), .QN(g25628) );
  NAND2X0 U18937 ( .IN1(n17891), .IN2(test_so76), .QN(n17890) );
  AND2X1 U18938 ( .IN1(n10366), .IN2(n17887), .Q(n17891) );
  NAND2X0 U18939 ( .IN1(n17892), .IN2(g1216), .QN(n17889) );
  NAND2X0 U18940 ( .IN1(n17893), .IN2(n10401), .QN(n17892) );
  OR2X1 U18941 ( .IN1(n17887), .IN2(test_so76), .Q(n17893) );
  NAND2X0 U18942 ( .IN1(n17894), .IN2(n17895), .QN(g25627) );
  NAND2X0 U18943 ( .IN1(n10502), .IN2(g1178), .QN(n17895) );
  NAND2X0 U18944 ( .IN1(n17896), .IN2(n10401), .QN(n17894) );
  NAND2X0 U18945 ( .IN1(n17897), .IN2(n17898), .QN(n17896) );
  OR2X1 U18946 ( .IN1(n17899), .IN2(n9757), .Q(n17898) );
  NAND2X0 U18947 ( .IN1(n17899), .IN2(g962), .QN(n17897) );
  NAND2X0 U18948 ( .IN1(n13173), .IN2(g7916), .QN(n17899) );
  NOR2X0 U18949 ( .IN1(n5599), .IN2(n5363), .QN(n13173) );
  NAND2X0 U18950 ( .IN1(n17900), .IN2(n17901), .QN(g25626) );
  NAND2X0 U18951 ( .IN1(n17902), .IN2(g1141), .QN(n17901) );
  NAND2X0 U18952 ( .IN1(n17903), .IN2(n10401), .QN(n17902) );
  NAND2X0 U18953 ( .IN1(n17904), .IN2(n17372), .QN(n17903) );
  NOR2X0 U18954 ( .IN1(n17905), .IN2(g956), .QN(n17904) );
  NAND2X0 U18955 ( .IN1(n17906), .IN2(g956), .QN(n17900) );
  NAND2X0 U18956 ( .IN1(n17907), .IN2(n17908), .QN(n17906) );
  NAND2X0 U18957 ( .IN1(n17909), .IN2(n10401), .QN(n17908) );
  NAND2X0 U18958 ( .IN1(n17372), .IN2(g1141), .QN(n17909) );
  INVX0 U18959 ( .INP(n17364), .ZN(n17372) );
  NAND2X0 U18960 ( .IN1(n5618), .IN2(test_so7), .QN(n17364) );
  NOR2X0 U18961 ( .IN1(g979), .IN2(n17910), .QN(g25625) );
  NAND2X0 U18962 ( .IN1(n17911), .IN2(n17377), .QN(n17910) );
  NAND2X0 U18963 ( .IN1(n17912), .IN2(n17913), .QN(n17377) );
  NOR2X0 U18964 ( .IN1(n9967), .IN2(n5654), .QN(n17912) );
  NAND2X0 U18965 ( .IN1(n17914), .IN2(n17915), .QN(n17911) );
  NAND2X0 U18966 ( .IN1(n13328), .IN2(n17913), .QN(n17915) );
  NAND2X0 U18967 ( .IN1(n10369), .IN2(g1052), .QN(n17914) );
  NAND2X0 U18968 ( .IN1(n17916), .IN2(n17917), .QN(g25624) );
  NAND2X0 U18969 ( .IN1(n17918), .IN2(n17380), .QN(n17917) );
  NOR2X0 U18970 ( .IN1(g1041), .IN2(n17919), .QN(n17918) );
  NOR2X0 U18971 ( .IN1(n17920), .IN2(n17921), .QN(n17916) );
  NOR2X0 U18972 ( .IN1(n9686), .IN2(n10355), .QN(n17921) );
  NOR2X0 U18973 ( .IN1(n10476), .IN2(n17922), .QN(n17920) );
  NAND2X0 U18974 ( .IN1(n17919), .IN2(g1041), .QN(n17922) );
  NAND2X0 U18975 ( .IN1(n17923), .IN2(n17924), .QN(g25623) );
  NAND2X0 U18976 ( .IN1(test_so20), .IN2(n17925), .QN(n17924) );
  NAND2X0 U18977 ( .IN1(n17919), .IN2(n10400), .QN(n17925) );
  NAND2X0 U18978 ( .IN1(n17380), .IN2(n17926), .QN(n17923) );
  NAND2X0 U18979 ( .IN1(n15542), .IN2(n17927), .QN(n17926) );
  NAND2X0 U18980 ( .IN1(n17928), .IN2(n17929), .QN(n17927) );
  INVX0 U18981 ( .INP(n17014), .ZN(n17929) );
  NAND2X0 U18982 ( .IN1(g1030), .IN2(g1018), .QN(n17928) );
  NOR2X0 U18983 ( .IN1(n10476), .IN2(n5321), .QN(n17380) );
  NOR2X0 U18984 ( .IN1(n10476), .IN2(n17930), .QN(g25622) );
  NOR2X0 U18985 ( .IN1(n17931), .IN2(n17932), .QN(n17930) );
  NOR2X0 U18986 ( .IN1(n17384), .IN2(n10152), .QN(n17932) );
  NOR2X0 U18987 ( .IN1(n17015), .IN2(n17933), .QN(n17931) );
  NOR2X0 U18988 ( .IN1(n17934), .IN2(n17935), .QN(n17933) );
  NOR2X0 U18989 ( .IN1(n4921), .IN2(g1008), .QN(n17935) );
  NAND2X0 U18990 ( .IN1(n17936), .IN2(n17937), .QN(n4921) );
  NOR2X0 U18991 ( .IN1(n9751), .IN2(n9728), .QN(n17937) );
  NOR2X0 U18992 ( .IN1(n9686), .IN2(n17013), .QN(n17936) );
  NOR2X0 U18993 ( .IN1(n17014), .IN2(n17012), .QN(n17934) );
  NAND2X0 U18994 ( .IN1(n17938), .IN2(g1008), .QN(n17012) );
  NOR2X0 U18995 ( .IN1(n9764), .IN2(n9763), .QN(n17938) );
  NOR2X0 U18996 ( .IN1(n17011), .IN2(n9910), .QN(n17014) );
  INVX0 U18997 ( .INP(n17013), .ZN(n17011) );
  INVX0 U18998 ( .INP(n15542), .ZN(n17015) );
  NAND2X0 U18999 ( .IN1(n17939), .IN2(n17940), .QN(g25621) );
  NAND2X0 U19000 ( .IN1(n17941), .IN2(g904), .QN(n17940) );
  NAND2X0 U19001 ( .IN1(n17942), .IN2(n10400), .QN(n17941) );
  NAND2X0 U19002 ( .IN1(n9740), .IN2(g12919), .QN(n17942) );
  NAND2X0 U19003 ( .IN1(g24231), .IN2(g921), .QN(n17939) );
  NOR2X0 U19004 ( .IN1(n5562), .IN2(n17943), .QN(g25619) );
  NOR2X0 U19005 ( .IN1(n10476), .IN2(n17944), .QN(n17943) );
  XOR2X1 U19006 ( .IN1(n17445), .IN2(g843), .Q(n17944) );
  NAND2X0 U19007 ( .IN1(n17945), .IN2(n17946), .QN(g25618) );
  NAND2X0 U19008 ( .IN1(n17947), .IN2(g832), .QN(n17946) );
  NAND2X0 U19009 ( .IN1(n17948), .IN2(n17949), .QN(n17947) );
  NAND2X0 U19010 ( .IN1(n16273), .IN2(n16231), .QN(n17949) );
  NAND2X0 U19011 ( .IN1(n5822), .IN2(n42), .QN(n17948) );
  NOR2X0 U19012 ( .IN1(n17950), .IN2(n10463), .QN(n42) );
  NAND2X0 U19013 ( .IN1(n17951), .IN2(g817), .QN(n17945) );
  NAND2X0 U19014 ( .IN1(n17952), .IN2(n10400), .QN(n17951) );
  NAND2X0 U19015 ( .IN1(n17953), .IN2(n10065), .QN(n17952) );
  NOR2X0 U19016 ( .IN1(n17950), .IN2(n16280), .QN(n17953) );
  INVX0 U19017 ( .INP(n16231), .ZN(n17950) );
  NAND2X0 U19018 ( .IN1(n17954), .IN2(n17955), .QN(g25617) );
  NAND2X0 U19019 ( .IN1(n17956), .IN2(n16231), .QN(n17955) );
  NAND2X0 U19020 ( .IN1(g847), .IN2(n17957), .QN(n16231) );
  NAND2X0 U19021 ( .IN1(n5733), .IN2(g837), .QN(n17957) );
  NOR2X0 U19022 ( .IN1(n17958), .IN2(n17959), .QN(n17956) );
  NOR2X0 U19023 ( .IN1(n5822), .IN2(n16273), .QN(n17959) );
  NOR2X0 U19024 ( .IN1(n16277), .IN2(g817), .QN(n17958) );
  NAND2X0 U19025 ( .IN1(n10502), .IN2(g812), .QN(n17954) );
  NOR2X0 U19026 ( .IN1(n10475), .IN2(n17960), .QN(g25616) );
  NOR2X0 U19027 ( .IN1(n17961), .IN2(n17962), .QN(n17960) );
  NAND2X0 U19028 ( .IN1(n17963), .IN2(n17964), .QN(n17962) );
  NAND2X0 U19029 ( .IN1(n17965), .IN2(g732), .QN(n17964) );
  NOR2X0 U19030 ( .IN1(n17449), .IN2(n17966), .QN(n17965) );
  NAND2X0 U19031 ( .IN1(n17966), .IN2(n5732), .QN(n17963) );
  AND2X1 U19032 ( .IN1(n17449), .IN2(n17966), .Q(n17961) );
  XOR2X1 U19033 ( .IN1(n17967), .IN2(n17968), .Q(n17966) );
  XOR2X1 U19034 ( .IN1(n17969), .IN2(n17970), .Q(n17968) );
  XOR2X1 U19035 ( .IN1(n9783), .IN2(n9782), .Q(n17970) );
  XOR2X1 U19036 ( .IN1(n9909), .IN2(n9908), .Q(n17969) );
  XOR2X1 U19037 ( .IN1(g225), .IN2(n17971), .Q(n17967) );
  XOR2X1 U19038 ( .IN1(n9781), .IN2(n6008), .Q(n17971) );
  INVX0 U19039 ( .INP(n17100), .ZN(n17449) );
  NAND2X0 U19040 ( .IN1(n17972), .IN2(n17973), .QN(n17100) );
  NOR2X0 U19041 ( .IN1(n17073), .IN2(n17974), .QN(n17973) );
  NAND2X0 U19042 ( .IN1(n5327), .IN2(n17975), .QN(n17974) );
  NAND2X0 U19043 ( .IN1(n5287), .IN2(n10135), .QN(n17073) );
  NOR2X0 U19044 ( .IN1(g370), .IN2(n17976), .QN(n17972) );
  NAND2X0 U19045 ( .IN1(n5820), .IN2(n5708), .QN(n17976) );
  NAND2X0 U19046 ( .IN1(n17977), .IN2(n17978), .QN(g25615) );
  NAND2X0 U19047 ( .IN1(n17060), .IN2(g667), .QN(n17978) );
  OR2X1 U19048 ( .IN1(n17060), .IN2(n9629), .Q(n17977) );
  NAND2X0 U19049 ( .IN1(n17979), .IN2(n17980), .QN(g25614) );
  NAND2X0 U19050 ( .IN1(n10502), .IN2(g691), .QN(n17980) );
  NOR2X0 U19051 ( .IN1(n17981), .IN2(n17982), .QN(n17979) );
  AND2X1 U19052 ( .IN1(n5111), .IN2(n17086), .Q(n17982) );
  NOR2X0 U19053 ( .IN1(n9629), .IN2(n17472), .QN(n17981) );
  NAND2X0 U19054 ( .IN1(n17983), .IN2(n17984), .QN(g25613) );
  NAND2X0 U19055 ( .IN1(n10502), .IN2(g559), .QN(n17984) );
  NAND2X0 U19056 ( .IN1(n17985), .IN2(n17986), .QN(n17983) );
  XOR2X1 U19057 ( .IN1(n9584), .IN2(n17464), .Q(n17986) );
  NAND2X0 U19058 ( .IN1(g29211), .IN2(n17987), .QN(n17464) );
  NAND2X0 U19059 ( .IN1(n9570), .IN2(g12368), .QN(n17987) );
  NOR2X0 U19060 ( .IN1(n17988), .IN2(n11200), .QN(n17985) );
  INVX0 U19061 ( .INP(n2421), .ZN(n11200) );
  NOR2X0 U19062 ( .IN1(n18472), .IN2(n5288), .QN(n17988) );
  NAND2X0 U19063 ( .IN1(n17989), .IN2(n17990), .QN(g25612) );
  NAND2X0 U19064 ( .IN1(n17991), .IN2(g513), .QN(n17990) );
  NAND2X0 U19065 ( .IN1(n17060), .IN2(g518), .QN(n17989) );
  NAND2X0 U19066 ( .IN1(n17992), .IN2(n17993), .QN(g25611) );
  NAND2X0 U19067 ( .IN1(n17991), .IN2(g504), .QN(n17993) );
  NAND2X0 U19068 ( .IN1(n17994), .IN2(n10400), .QN(n17991) );
  NAND2X0 U19069 ( .IN1(n17086), .IN2(n17084), .QN(n17994) );
  INVX0 U19070 ( .INP(n4962), .ZN(n17084) );
  NAND2X0 U19071 ( .IN1(n17060), .IN2(g513), .QN(n17992) );
  NAND2X0 U19072 ( .IN1(n17995), .IN2(n17996), .QN(g25610) );
  NOR2X0 U19073 ( .IN1(n17997), .IN2(n17998), .QN(n17995) );
  NOR2X0 U19074 ( .IN1(n17060), .IN2(n10135), .QN(n17998) );
  NOR2X0 U19075 ( .IN1(n5519), .IN2(n17472), .QN(n17997) );
  NAND2X0 U19076 ( .IN1(n17999), .IN2(n18000), .QN(g25609) );
  NAND2X0 U19077 ( .IN1(n18001), .IN2(n5287), .QN(n18000) );
  NOR2X0 U19078 ( .IN1(n18002), .IN2(n18003), .QN(n17999) );
  NOR2X0 U19079 ( .IN1(n18004), .IN2(n10135), .QN(n18003) );
  NOR2X0 U19080 ( .IN1(n18005), .IN2(n17060), .QN(n18004) );
  INVX0 U19081 ( .INP(n17472), .ZN(n17060) );
  NAND2X0 U19082 ( .IN1(n17474), .IN2(n10400), .QN(n17472) );
  NOR2X0 U19083 ( .IN1(n10475), .IN2(g513), .QN(n18005) );
  INVX0 U19084 ( .INP(n17996), .ZN(n18002) );
  NAND2X0 U19085 ( .IN1(n4962), .IN2(n18001), .QN(n17996) );
  INVX0 U19086 ( .INP(n17052), .ZN(n18001) );
  NAND2X0 U19087 ( .IN1(n17086), .IN2(n10400), .QN(n17052) );
  INVX0 U19088 ( .INP(n17474), .ZN(n17086) );
  NAND2X0 U19089 ( .IN1(n18006), .IN2(n5633), .QN(n17474) );
  NOR2X0 U19090 ( .IN1(n9785), .IN2(n5632), .QN(n18006) );
  NAND2X0 U19091 ( .IN1(n18007), .IN2(n18008), .QN(g25605) );
  NAND2X0 U19092 ( .IN1(n10502), .IN2(g168), .QN(n18008) );
  NOR2X0 U19093 ( .IN1(n18009), .IN2(n18010), .QN(n18007) );
  NOR2X0 U19094 ( .IN1(n9661), .IN2(n18011), .QN(n18010) );
  NOR2X0 U19095 ( .IN1(n18012), .IN2(n18013), .QN(n18009) );
  NAND2X0 U19096 ( .IN1(n17975), .IN2(g246), .QN(n18013) );
  NAND2X0 U19097 ( .IN1(n18014), .IN2(n18015), .QN(g25604) );
  OR2X1 U19098 ( .IN1(n18011), .IN2(n9914), .Q(n18015) );
  OR2X1 U19099 ( .IN1(n18016), .IN2(n9661), .Q(n18014) );
  NAND2X0 U19100 ( .IN1(n18017), .IN2(n18018), .QN(g25602) );
  NAND2X0 U19101 ( .IN1(n10502), .IN2(g405), .QN(n18018) );
  NOR2X0 U19102 ( .IN1(n18019), .IN2(n18020), .QN(n18017) );
  NOR2X0 U19103 ( .IN1(n10136), .IN2(n18011), .QN(n18020) );
  NOR2X0 U19104 ( .IN1(n18012), .IN2(n18021), .QN(n18019) );
  NAND2X0 U19105 ( .IN1(n17975), .IN2(g446), .QN(n18021) );
  NAND2X0 U19106 ( .IN1(n18022), .IN2(n18023), .QN(g25601) );
  NAND2X0 U19107 ( .IN1(n18016), .IN2(g174), .QN(n18023) );
  NAND2X0 U19108 ( .IN1(test_so72), .IN2(n18011), .QN(n18022) );
  NAND2X0 U19109 ( .IN1(n18024), .IN2(n18025), .QN(g25600) );
  NAND2X0 U19110 ( .IN1(n18016), .IN2(g168), .QN(n18025) );
  INVX0 U19111 ( .INP(n18011), .ZN(n18016) );
  NAND2X0 U19112 ( .IN1(n18011), .IN2(g174), .QN(n18024) );
  NAND2X0 U19113 ( .IN1(n18026), .IN2(n10399), .QN(n18011) );
  NAND2X0 U19114 ( .IN1(n9787), .IN2(n17975), .QN(n18026) );
  NAND2X0 U19115 ( .IN1(n11667), .IN2(n18027), .QN(g25599) );
  NAND2X0 U19116 ( .IN1(n10502), .IN2(g385), .QN(n18027) );
  NAND2X0 U19117 ( .IN1(n18028), .IN2(n18029), .QN(g25598) );
  NAND2X0 U19118 ( .IN1(n18030), .IN2(n5121), .QN(n18029) );
  NOR2X0 U19119 ( .IN1(n5632), .IN2(n10463), .QN(n18030) );
  NAND2X0 U19120 ( .IN1(n18031), .IN2(g376), .QN(n18028) );
  NAND2X0 U19121 ( .IN1(n18032), .IN2(n10399), .QN(n18031) );
  OR2X1 U19122 ( .IN1(n17975), .IN2(n9785), .Q(n18032) );
  INVX0 U19123 ( .INP(n5121), .ZN(n17975) );
  NAND2X0 U19124 ( .IN1(n18033), .IN2(g385), .QN(n5121) );
  NOR2X0 U19125 ( .IN1(n9785), .IN2(n5633), .QN(n18033) );
  NAND2X0 U19126 ( .IN1(n18034), .IN2(n18035), .QN(g25597) );
  OR2X1 U19127 ( .IN1(n11667), .IN2(n18012), .Q(n18035) );
  NAND2X0 U19128 ( .IN1(n9787), .IN2(n10399), .QN(n18012) );
  NOR2X0 U19129 ( .IN1(n18036), .IN2(n18037), .QN(n18034) );
  NOR2X0 U19130 ( .IN1(n9785), .IN2(n10356), .QN(n18037) );
  NOR2X0 U19131 ( .IN1(n10475), .IN2(n18038), .QN(n18036) );
  NAND2X0 U19132 ( .IN1(n11667), .IN2(g370), .QN(n18038) );
  NAND2X0 U19133 ( .IN1(n18039), .IN2(g385), .QN(n11667) );
  NOR2X0 U19134 ( .IN1(n9786), .IN2(n5633), .QN(n18039) );
  NAND2X0 U19135 ( .IN1(n18040), .IN2(n18041), .QN(g25596) );
  NAND2X0 U19136 ( .IN1(n10502), .IN2(g370), .QN(n18041) );
  NAND2X0 U19137 ( .IN1(n18042), .IN2(n10399), .QN(n18040) );
  XOR2X1 U19138 ( .IN1(n9785), .IN2(n5633), .Q(n18042) );
  NOR2X0 U19139 ( .IN1(g8719), .IN2(n18043), .QN(g25595) );
  NAND2X0 U19140 ( .IN1(n9785), .IN2(n10399), .QN(n18043) );
  NOR2X0 U19141 ( .IN1(n17101), .IN2(n18044), .QN(g25594) );
  NAND2X0 U19142 ( .IN1(n17103), .IN2(n10399), .QN(n18044) );
  NAND2X0 U19143 ( .IN1(n18045), .IN2(n18046), .QN(n17103) );
  NOR2X0 U19144 ( .IN1(n18047), .IN2(n18048), .QN(n18046) );
  NAND2X0 U19145 ( .IN1(g225), .IN2(g246), .QN(n18048) );
  NAND2X0 U19146 ( .IN1(g232), .IN2(g239), .QN(n18047) );
  NOR2X0 U19147 ( .IN1(g269), .IN2(n18049), .QN(n18045) );
  NAND2X0 U19148 ( .IN1(n9782), .IN2(n9781), .QN(n18049) );
  AND2X1 U19149 ( .IN1(n5627), .IN2(n18050), .Q(n17101) );
  NAND2X0 U19150 ( .IN1(n18051), .IN2(n18052), .QN(n18050) );
  NOR2X0 U19151 ( .IN1(n18053), .IN2(n18054), .QN(n18052) );
  NAND2X0 U19152 ( .IN1(n5597), .IN2(g255), .QN(n18054) );
  NAND2X0 U19153 ( .IN1(g262), .IN2(g269), .QN(n18053) );
  NOR2X0 U19154 ( .IN1(g239), .IN2(n18055), .QN(n18051) );
  NAND2X0 U19155 ( .IN1(n9908), .IN2(n6008), .QN(n18055) );
  NAND2X0 U19156 ( .IN1(n18056), .IN2(n18057), .QN(g25593) );
  OR2X1 U19157 ( .IN1(n10310), .IN2(n9760), .Q(n18057) );
  NAND2X0 U19158 ( .IN1(n18058), .IN2(n10398), .QN(n18056) );
  NAND2X0 U19159 ( .IN1(n18059), .IN2(n18060), .QN(n18058) );
  NAND2X0 U19160 ( .IN1(n18061), .IN2(g209), .QN(n18060) );
  NAND2X0 U19161 ( .IN1(n18062), .IN2(n18063), .QN(n18059) );
  INVX0 U19162 ( .INP(n18061), .ZN(n18063) );
  NAND2X0 U19163 ( .IN1(n18064), .IN2(n18065), .QN(g25592) );
  OR2X1 U19164 ( .IN1(n10310), .IN2(n10099), .Q(n18065) );
  NAND2X0 U19165 ( .IN1(n18066), .IN2(n10398), .QN(n18064) );
  XNOR2X1 U19166 ( .IN1(n9759), .IN2(n18067), .Q(n18066) );
  NOR2X0 U19167 ( .IN1(n18061), .IN2(n18062), .QN(n18067) );
  XOR2X1 U19168 ( .IN1(n9759), .IN2(n9760), .Q(n18062) );
  NAND2X0 U19169 ( .IN1(test_so42), .IN2(g218), .QN(n18061) );
  NAND2X0 U19170 ( .IN1(n18068), .IN2(n18069), .QN(g25591) );
  NAND2X0 U19171 ( .IN1(n10050), .IN2(n10398), .QN(n18069) );
  NAND2X0 U19172 ( .IN1(n10502), .IN2(g209), .QN(n18068) );
  INVX0 U19173 ( .INP(n10666), .ZN(g25114) );
  NAND2X0 U19174 ( .IN1(g5297), .IN2(g5357), .QN(n10666) );
  NOR2X0 U19175 ( .IN1(n10037), .IN2(n18070), .QN(g24355) );
  AND2X1 U19176 ( .IN1(n10366), .IN2(n18071), .Q(n18070) );
  NAND2X0 U19177 ( .IN1(n18072), .IN2(n18073), .QN(g24354) );
  NAND2X0 U19178 ( .IN1(n10501), .IN2(g6727), .QN(n18073) );
  NAND2X0 U19179 ( .IN1(n18074), .IN2(n10398), .QN(n18072) );
  NOR2X0 U19180 ( .IN1(n18071), .IN2(g6736), .QN(n18074) );
  NOR2X0 U19181 ( .IN1(n18075), .IN2(n5531), .QN(n18071) );
  NAND2X0 U19182 ( .IN1(n18076), .IN2(n18077), .QN(g24353) );
  NAND2X0 U19183 ( .IN1(n10501), .IN2(g6723), .QN(n18077) );
  NAND2X0 U19184 ( .IN1(n18078), .IN2(n10397), .QN(n18076) );
  XOR2X1 U19185 ( .IN1(n18075), .IN2(n5531), .Q(n18078) );
  NAND2X0 U19186 ( .IN1(n18079), .IN2(n18080), .QN(n18075) );
  NOR2X0 U19187 ( .IN1(n9890), .IN2(n9876), .QN(n18080) );
  AND2X1 U19188 ( .IN1(g14828), .IN2(test_so80), .Q(n18079) );
  NOR2X0 U19189 ( .IN1(n18081), .IN2(n18082), .QN(g24352) );
  NAND2X0 U19190 ( .IN1(n18083), .IN2(n9995), .QN(n18082) );
  NOR2X0 U19191 ( .IN1(n18084), .IN2(n18085), .QN(n18083) );
  NOR2X0 U19192 ( .IN1(test_so80), .IN2(n5700), .QN(n18085) );
  NOR2X0 U19193 ( .IN1(n9890), .IN2(g14828), .QN(n18084) );
  NAND2X0 U19194 ( .IN1(n18086), .IN2(n9876), .QN(n18081) );
  NOR2X0 U19195 ( .IN1(n10475), .IN2(g13099), .QN(n18086) );
  NOR2X0 U19196 ( .IN1(n9899), .IN2(n18087), .QN(g24351) );
  AND2X1 U19197 ( .IN1(n10366), .IN2(n18088), .Q(n18087) );
  NAND2X0 U19198 ( .IN1(n18089), .IN2(n18090), .QN(g24350) );
  NAND2X0 U19199 ( .IN1(test_so69), .IN2(n10515), .QN(n18090) );
  NAND2X0 U19200 ( .IN1(n18091), .IN2(n10397), .QN(n18089) );
  NOR2X0 U19201 ( .IN1(n18088), .IN2(g6390), .QN(n18091) );
  NOR2X0 U19202 ( .IN1(n18092), .IN2(n10130), .QN(n18088) );
  NAND2X0 U19203 ( .IN1(n18093), .IN2(n18094), .QN(g24349) );
  NAND2X0 U19204 ( .IN1(n10501), .IN2(g6377), .QN(n18094) );
  NAND2X0 U19205 ( .IN1(n18095), .IN2(n10397), .QN(n18093) );
  XOR2X1 U19206 ( .IN1(n10130), .IN2(n18092), .Q(n18095) );
  NAND2X0 U19207 ( .IN1(n18096), .IN2(n18097), .QN(n18092) );
  NOR2X0 U19208 ( .IN1(n9894), .IN2(n9879), .QN(n18097) );
  NOR2X0 U19209 ( .IN1(n5703), .IN2(n5437), .QN(n18096) );
  NOR2X0 U19210 ( .IN1(n18098), .IN2(n18099), .QN(g24348) );
  NAND2X0 U19211 ( .IN1(n18100), .IN2(n9879), .QN(n18099) );
  NOR2X0 U19212 ( .IN1(n18101), .IN2(n18102), .QN(n18100) );
  NOR2X0 U19213 ( .IN1(n5703), .IN2(g12422), .QN(n18102) );
  NOR2X0 U19214 ( .IN1(n9894), .IN2(g14779), .QN(n18101) );
  NAND2X0 U19215 ( .IN1(n18103), .IN2(n10032), .QN(n18098) );
  NOR2X0 U19216 ( .IN1(n10475), .IN2(g17685), .QN(n18103) );
  NOR2X0 U19217 ( .IN1(n9900), .IN2(n18104), .QN(g24347) );
  AND2X1 U19218 ( .IN1(n10366), .IN2(n18105), .Q(n18104) );
  NAND2X0 U19219 ( .IN1(n18106), .IN2(n18107), .QN(g24346) );
  NAND2X0 U19220 ( .IN1(n10501), .IN2(g6035), .QN(n18107) );
  NAND2X0 U19221 ( .IN1(n18108), .IN2(n10397), .QN(n18106) );
  NOR2X0 U19222 ( .IN1(test_so50), .IN2(n18105), .QN(n18108) );
  NOR2X0 U19223 ( .IN1(n18109), .IN2(n5528), .QN(n18105) );
  NAND2X0 U19224 ( .IN1(n18110), .IN2(n18111), .QN(g24345) );
  NAND2X0 U19225 ( .IN1(n10501), .IN2(g6031), .QN(n18111) );
  NAND2X0 U19226 ( .IN1(n18112), .IN2(n10397), .QN(n18110) );
  XOR2X1 U19227 ( .IN1(n18109), .IN2(n5528), .Q(n18112) );
  NAND2X0 U19228 ( .IN1(n18113), .IN2(n18114), .QN(n18109) );
  NOR2X0 U19229 ( .IN1(n9885), .IN2(n9870), .QN(n18114) );
  NOR2X0 U19230 ( .IN1(n5698), .IN2(n5432), .QN(n18113) );
  NOR2X0 U19231 ( .IN1(n18115), .IN2(n18116), .QN(g24344) );
  NAND2X0 U19232 ( .IN1(n18117), .IN2(n9981), .QN(n18116) );
  NOR2X0 U19233 ( .IN1(n18118), .IN2(n18119), .QN(n18117) );
  NOR2X0 U19234 ( .IN1(n5698), .IN2(g12350), .QN(n18119) );
  NOR2X0 U19235 ( .IN1(n9885), .IN2(g14738), .QN(n18118) );
  NAND2X0 U19236 ( .IN1(n18120), .IN2(n9870), .QN(n18115) );
  NOR2X0 U19237 ( .IN1(n10475), .IN2(g13068), .QN(n18120) );
  NOR2X0 U19238 ( .IN1(n9904), .IN2(n18121), .QN(g24343) );
  AND2X1 U19239 ( .IN1(n10367), .IN2(n18122), .Q(n18121) );
  NAND2X0 U19240 ( .IN1(n18123), .IN2(n18124), .QN(g24342) );
  NAND2X0 U19241 ( .IN1(n10501), .IN2(g5689), .QN(n18124) );
  NAND2X0 U19242 ( .IN1(n18125), .IN2(n10397), .QN(n18123) );
  NOR2X0 U19243 ( .IN1(n18122), .IN2(g5698), .QN(n18125) );
  NOR2X0 U19244 ( .IN1(n18126), .IN2(n5529), .QN(n18122) );
  NAND2X0 U19245 ( .IN1(n18127), .IN2(n18128), .QN(g24341) );
  NAND2X0 U19246 ( .IN1(n10501), .IN2(g5685), .QN(n18128) );
  NAND2X0 U19247 ( .IN1(n18129), .IN2(n10397), .QN(n18127) );
  XOR2X1 U19248 ( .IN1(n18126), .IN2(n5529), .Q(n18129) );
  NAND2X0 U19249 ( .IN1(n18130), .IN2(n18131), .QN(n18126) );
  NOR2X0 U19250 ( .IN1(n9887), .IN2(n9872), .QN(n18131) );
  NOR2X0 U19251 ( .IN1(n5705), .IN2(n5439), .QN(n18130) );
  NOR2X0 U19252 ( .IN1(n18132), .IN2(n18133), .QN(g24340) );
  NAND2X0 U19253 ( .IN1(n18134), .IN2(n9986), .QN(n18133) );
  NOR2X0 U19254 ( .IN1(n18135), .IN2(n18136), .QN(n18134) );
  NOR2X0 U19255 ( .IN1(n5705), .IN2(g12300), .QN(n18136) );
  NOR2X0 U19256 ( .IN1(n9887), .IN2(g14694), .QN(n18135) );
  NAND2X0 U19257 ( .IN1(n18137), .IN2(n9872), .QN(n18132) );
  NOR2X0 U19258 ( .IN1(n10475), .IN2(g13049), .QN(n18137) );
  NOR2X0 U19259 ( .IN1(n10039), .IN2(n18138), .QN(g24339) );
  AND2X1 U19260 ( .IN1(n10367), .IN2(n18139), .Q(n18138) );
  NAND2X0 U19261 ( .IN1(n18140), .IN2(n18141), .QN(g24338) );
  NAND2X0 U19262 ( .IN1(test_so10), .IN2(n10515), .QN(n18141) );
  NAND2X0 U19263 ( .IN1(n18142), .IN2(n10401), .QN(n18140) );
  NOR2X0 U19264 ( .IN1(n18139), .IN2(g5352), .QN(n18142) );
  NOR2X0 U19265 ( .IN1(n18143), .IN2(n10129), .QN(n18139) );
  NAND2X0 U19266 ( .IN1(n18144), .IN2(n18145), .QN(g24337) );
  NAND2X0 U19267 ( .IN1(n10501), .IN2(g5339), .QN(n18145) );
  NAND2X0 U19268 ( .IN1(n18146), .IN2(n10378), .QN(n18144) );
  XOR2X1 U19269 ( .IN1(n10129), .IN2(n18143), .Q(n18146) );
  NAND2X0 U19270 ( .IN1(n18147), .IN2(n18148), .QN(n18143) );
  NOR2X0 U19271 ( .IN1(n9883), .IN2(n9868), .QN(n18148) );
  NOR2X0 U19272 ( .IN1(n5704), .IN2(n5438), .QN(n18147) );
  NOR2X0 U19273 ( .IN1(n18149), .IN2(n18150), .QN(g24336) );
  NAND2X0 U19274 ( .IN1(n18151), .IN2(n9976), .QN(n18150) );
  NOR2X0 U19275 ( .IN1(n18152), .IN2(n18153), .QN(n18151) );
  NOR2X0 U19276 ( .IN1(n5704), .IN2(g12238), .QN(n18153) );
  NOR2X0 U19277 ( .IN1(n9883), .IN2(g14662), .QN(n18152) );
  NAND2X0 U19278 ( .IN1(n18154), .IN2(n9953), .QN(n18149) );
  NOR2X0 U19279 ( .IN1(n10475), .IN2(g17519), .QN(n18154) );
  NAND2X0 U19280 ( .IN1(n18155), .IN2(n18156), .QN(g24335) );
  NAND2X0 U19281 ( .IN1(n18157), .IN2(n18158), .QN(n18156) );
  NOR2X0 U19282 ( .IN1(n5382), .IN2(g4340), .QN(n18157) );
  OR2X1 U19283 ( .IN1(n10311), .IN2(n5541), .Q(n18155) );
  NAND2X0 U19284 ( .IN1(n18159), .IN2(n18160), .QN(g24334) );
  NAND2X0 U19285 ( .IN1(n18161), .IN2(n18162), .QN(n18160) );
  NOR2X0 U19286 ( .IN1(n18163), .IN2(n18164), .QN(n18162) );
  NAND2X0 U19287 ( .IN1(n5303), .IN2(n5365), .QN(n18164) );
  NAND2X0 U19288 ( .IN1(n11850), .IN2(g4633), .QN(n18163) );
  AND2X1 U19289 ( .IN1(n18165), .IN2(test_so3), .Q(n11850) );
  NOR2X0 U19290 ( .IN1(n5653), .IN2(g4639), .QN(n18165) );
  NOR2X0 U19291 ( .IN1(n18166), .IN2(n18167), .QN(n18161) );
  NAND2X0 U19292 ( .IN1(n18158), .IN2(n5608), .QN(n18167) );
  AND2X1 U19293 ( .IN1(n18168), .IN2(n18169), .Q(n18158) );
  NOR2X0 U19294 ( .IN1(g4322), .IN2(n18170), .QN(n18169) );
  NAND2X0 U19295 ( .IN1(n10367), .IN2(n10132), .QN(n18170) );
  NOR2X0 U19296 ( .IN1(g4358), .IN2(n18171), .QN(n18168) );
  NAND2X0 U19297 ( .IN1(n5323), .IN2(n5540), .QN(n18171) );
  NAND2X0 U19298 ( .IN1(n5274), .IN2(n5539), .QN(n18166) );
  NAND2X0 U19299 ( .IN1(n10501), .IN2(g4358), .QN(n18159) );
  NOR2X0 U19300 ( .IN1(n5710), .IN2(n10353), .QN(g24298) );
  NAND2X0 U19301 ( .IN1(n18172), .IN2(n18173), .QN(g24282) );
  NAND2X0 U19302 ( .IN1(n18174), .IN2(g4308), .QN(n18173) );
  NAND2X0 U19303 ( .IN1(n10367), .IN2(g9251), .QN(n18174) );
  NAND2X0 U19304 ( .IN1(g24281), .IN2(g9251), .QN(n18172) );
  NOR2X0 U19305 ( .IN1(g4308), .IN2(n10462), .QN(g24281) );
  NAND2X0 U19306 ( .IN1(n18175), .IN2(n18176), .QN(g24280) );
  NAND2X0 U19307 ( .IN1(n18177), .IN2(g4269), .QN(n18176) );
  NAND2X0 U19308 ( .IN1(n18178), .IN2(n10380), .QN(n18177) );
  NAND2X0 U19309 ( .IN1(n18179), .IN2(n5764), .QN(n18178) );
  NOR2X0 U19310 ( .IN1(n9614), .IN2(n5823), .QN(n18179) );
  NAND2X0 U19311 ( .IN1(n18180), .IN2(g4273), .QN(n18175) );
  NAND2X0 U19312 ( .IN1(n18181), .IN2(n18182), .QN(n18180) );
  NAND2X0 U19313 ( .IN1(n5763), .IN2(n10378), .QN(n18182) );
  NAND2X0 U19314 ( .IN1(n18183), .IN2(n18184), .QN(g24279) );
  NAND2X0 U19315 ( .IN1(n18185), .IN2(n18186), .QN(n18184) );
  NOR2X0 U19316 ( .IN1(n18187), .IN2(n18188), .QN(n18183) );
  NOR2X0 U19317 ( .IN1(n10475), .IN2(n18189), .QN(n18188) );
  NOR2X0 U19318 ( .IN1(n18190), .IN2(n18191), .QN(n18189) );
  AND2X1 U19319 ( .IN1(n18186), .IN2(n18192), .Q(n18191) );
  NOR2X0 U19320 ( .IN1(n18192), .IN2(n18193), .QN(n18190) );
  OR2X1 U19321 ( .IN1(n18186), .IN2(n18185), .Q(n18193) );
  NOR2X0 U19322 ( .IN1(n9834), .IN2(n5726), .QN(n18185) );
  AND2X1 U19323 ( .IN1(n18194), .IN2(n9834), .Q(n18192) );
  NOR2X0 U19324 ( .IN1(n18195), .IN2(g8870), .QN(n18194) );
  NOR2X0 U19325 ( .IN1(n18196), .IN2(n18197), .QN(n18195) );
  NAND2X0 U19326 ( .IN1(n18198), .IN2(n18469), .QN(n18197) );
  NOR2X0 U19327 ( .IN1(g8919), .IN2(g11770), .QN(n18198) );
  NAND2X0 U19328 ( .IN1(n18199), .IN2(n18200), .QN(n18196) );
  NOR2X0 U19329 ( .IN1(g8915), .IN2(g8918), .QN(n18200) );
  NOR2X0 U19330 ( .IN1(g8917), .IN2(g8920), .QN(n18199) );
  NOR2X0 U19331 ( .IN1(n9834), .IN2(n10353), .QN(n18187) );
  NOR2X0 U19332 ( .IN1(n9906), .IN2(n18201), .QN(g24278) );
  AND2X1 U19333 ( .IN1(n10366), .IN2(n18202), .Q(n18201) );
  NAND2X0 U19334 ( .IN1(n18203), .IN2(n18204), .QN(g24277) );
  NAND2X0 U19335 ( .IN1(n10501), .IN2(g4040), .QN(n18204) );
  NAND2X0 U19336 ( .IN1(n18205), .IN2(n10379), .QN(n18203) );
  NOR2X0 U19337 ( .IN1(n18202), .IN2(g4049), .QN(n18205) );
  NOR2X0 U19338 ( .IN1(n18206), .IN2(n5530), .QN(n18202) );
  NAND2X0 U19339 ( .IN1(n18207), .IN2(n18208), .QN(g24276) );
  NAND2X0 U19340 ( .IN1(n10501), .IN2(g4031), .QN(n18208) );
  NAND2X0 U19341 ( .IN1(n18209), .IN2(n10379), .QN(n18207) );
  XOR2X1 U19342 ( .IN1(n18206), .IN2(n5530), .Q(n18209) );
  NAND2X0 U19343 ( .IN1(n18210), .IN2(n18211), .QN(n18206) );
  NOR2X0 U19344 ( .IN1(n9888), .IN2(n9874), .QN(n18211) );
  NOR2X0 U19345 ( .IN1(n5701), .IN2(n5435), .QN(n18210) );
  NOR2X0 U19346 ( .IN1(n18212), .IN2(n18213), .QN(g24275) );
  NAND2X0 U19347 ( .IN1(n18214), .IN2(n9990), .QN(n18213) );
  NOR2X0 U19348 ( .IN1(n18215), .IN2(n18216), .QN(n18214) );
  NOR2X0 U19349 ( .IN1(n5701), .IN2(g11418), .QN(n18216) );
  NOR2X0 U19350 ( .IN1(n9888), .IN2(g13966), .QN(n18215) );
  NAND2X0 U19351 ( .IN1(n18217), .IN2(n9874), .QN(n18212) );
  NOR2X0 U19352 ( .IN1(n10475), .IN2(g14518), .QN(n18217) );
  NOR2X0 U19353 ( .IN1(n9902), .IN2(n18218), .QN(g24274) );
  AND2X1 U19354 ( .IN1(n10367), .IN2(n18219), .Q(n18218) );
  NAND2X0 U19355 ( .IN1(n18220), .IN2(n18221), .QN(g24273) );
  NAND2X0 U19356 ( .IN1(n10501), .IN2(g3689), .QN(n18221) );
  NAND2X0 U19357 ( .IN1(n18222), .IN2(n10378), .QN(n18220) );
  NOR2X0 U19358 ( .IN1(n18219), .IN2(g3698), .QN(n18222) );
  NOR2X0 U19359 ( .IN1(n18223), .IN2(n5532), .QN(n18219) );
  NAND2X0 U19360 ( .IN1(n18224), .IN2(n18225), .QN(g24272) );
  NAND2X0 U19361 ( .IN1(n10500), .IN2(g3680), .QN(n18225) );
  NAND2X0 U19362 ( .IN1(n18226), .IN2(n10378), .QN(n18224) );
  XOR2X1 U19363 ( .IN1(n18223), .IN2(n5532), .Q(n18226) );
  NAND2X0 U19364 ( .IN1(n18227), .IN2(n18228), .QN(n18223) );
  NOR2X0 U19365 ( .IN1(n9892), .IN2(n9878), .QN(n18228) );
  NOR2X0 U19366 ( .IN1(n5699), .IN2(n5433), .QN(n18227) );
  NOR2X0 U19367 ( .IN1(n18229), .IN2(n18230), .QN(g24271) );
  NAND2X0 U19368 ( .IN1(n18231), .IN2(n9878), .QN(n18230) );
  NOR2X0 U19369 ( .IN1(n18232), .IN2(n18233), .QN(n18231) );
  NOR2X0 U19370 ( .IN1(n5699), .IN2(g11388), .QN(n18233) );
  NOR2X0 U19371 ( .IN1(n9892), .IN2(g13926), .QN(n18232) );
  NAND2X0 U19372 ( .IN1(n18234), .IN2(n10028), .QN(n18229) );
  NOR2X0 U19373 ( .IN1(n10475), .IN2(g16656), .QN(n18234) );
  NOR2X0 U19374 ( .IN1(n9897), .IN2(n18235), .QN(g24270) );
  AND2X1 U19375 ( .IN1(n10367), .IN2(n18236), .Q(n18235) );
  NAND2X0 U19376 ( .IN1(n18237), .IN2(n18238), .QN(g24269) );
  NAND2X0 U19377 ( .IN1(n10500), .IN2(g3338), .QN(n18238) );
  NAND2X0 U19378 ( .IN1(n18239), .IN2(n10379), .QN(n18237) );
  NOR2X0 U19379 ( .IN1(n18236), .IN2(g3347), .QN(n18239) );
  NOR2X0 U19380 ( .IN1(n18240), .IN2(n5527), .QN(n18236) );
  NAND2X0 U19381 ( .IN1(n18241), .IN2(n18242), .QN(g24268) );
  NAND2X0 U19382 ( .IN1(test_so91), .IN2(n10515), .QN(n18242) );
  NAND2X0 U19383 ( .IN1(n18243), .IN2(n10379), .QN(n18241) );
  XOR2X1 U19384 ( .IN1(n18240), .IN2(n5527), .Q(n18243) );
  NAND2X0 U19385 ( .IN1(n18244), .IN2(n18245), .QN(n18240) );
  NOR2X0 U19386 ( .IN1(n9881), .IN2(n9866), .QN(n18245) );
  NOR2X0 U19387 ( .IN1(n5702), .IN2(n5436), .QN(n18244) );
  NOR2X0 U19388 ( .IN1(n18246), .IN2(n18247), .QN(g24267) );
  NAND2X0 U19389 ( .IN1(n18248), .IN2(n9971), .QN(n18247) );
  NOR2X0 U19390 ( .IN1(n18249), .IN2(n18250), .QN(n18248) );
  NOR2X0 U19391 ( .IN1(n5702), .IN2(g11349), .QN(n18250) );
  NOR2X0 U19392 ( .IN1(n9881), .IN2(g13895), .QN(n18249) );
  NAND2X0 U19393 ( .IN1(n18251), .IN2(n9866), .QN(n18246) );
  NOR2X0 U19394 ( .IN1(n10475), .IN2(g14421), .QN(n18251) );
  NAND2X0 U19395 ( .IN1(n18252), .IN2(n18253), .QN(g24266) );
  OR2X1 U19396 ( .IN1(n10309), .IN2(n5963), .Q(n18253) );
  NAND2X0 U19397 ( .IN1(n18254), .IN2(n10379), .QN(n18252) );
  NOR2X0 U19398 ( .IN1(g2712), .IN2(n18470), .QN(n18254) );
  NAND2X0 U19399 ( .IN1(n18255), .IN2(n13609), .QN(g24263) );
  NAND2X0 U19400 ( .IN1(n5963), .IN2(n10379), .QN(n13609) );
  NOR2X0 U19401 ( .IN1(n18256), .IN2(n18257), .QN(n18255) );
  NOR2X0 U19402 ( .IN1(n9630), .IN2(n10356), .QN(n18257) );
  NOR2X0 U19403 ( .IN1(n10475), .IN2(g2715), .QN(n18256) );
  NAND2X0 U19404 ( .IN1(n18258), .IN2(n18259), .QN(g24262) );
  NAND2X0 U19405 ( .IN1(n18260), .IN2(n10066), .QN(n18259) );
  NOR2X0 U19406 ( .IN1(n18261), .IN2(n18262), .QN(n18258) );
  NOR2X0 U19407 ( .IN1(n5546), .IN2(n10356), .QN(n18262) );
  NOR2X0 U19408 ( .IN1(n10475), .IN2(n18263), .QN(n18261) );
  OR2X1 U19409 ( .IN1(n18260), .IN2(n10066), .Q(n18263) );
  NAND2X0 U19410 ( .IN1(n17853), .IN2(n18264), .QN(g24261) );
  NAND2X0 U19411 ( .IN1(n10500), .IN2(g1585), .QN(n18264) );
  XOR2X1 U19412 ( .IN1(n18265), .IN2(n10067), .Q(g24260) );
  OR2X1 U19413 ( .IN1(n10457), .IN2(n5546), .Q(n18265) );
  NAND2X0 U19414 ( .IN1(n17853), .IN2(n18266), .QN(g24259) );
  OR2X1 U19415 ( .IN1(n10310), .IN2(n9722), .Q(n18266) );
  NAND2X0 U19416 ( .IN1(n18267), .IN2(n18268), .QN(g24258) );
  NAND2X0 U19417 ( .IN1(n10368), .IN2(g496), .QN(n18268) );
  NAND2X0 U19418 ( .IN1(n10500), .IN2(g1554), .QN(n18267) );
  XOR2X1 U19419 ( .IN1(n18269), .IN2(n5616), .Q(g24257) );
  NAND2X0 U19420 ( .IN1(n18270), .IN2(n10380), .QN(n18269) );
  NAND2X0 U19421 ( .IN1(n18271), .IN2(n18272), .QN(g24256) );
  NAND2X0 U19422 ( .IN1(n10500), .IN2(g1339), .QN(n18272) );
  NAND2X0 U19423 ( .IN1(n18273), .IN2(n10380), .QN(n18271) );
  XOR2X1 U19424 ( .IN1(n18270), .IN2(n18274), .Q(n18273) );
  NOR2X0 U19425 ( .IN1(g13272), .IN2(n18275), .QN(n18274) );
  NAND2X0 U19426 ( .IN1(n9651), .IN2(n17852), .QN(n18275) );
  INVX0 U19427 ( .INP(n17849), .ZN(n17852) );
  NAND2X0 U19428 ( .IN1(n18276), .IN2(n5401), .QN(n17849) );
  NOR2X0 U19429 ( .IN1(g1333), .IN2(g7946), .QN(n18276) );
  AND2X1 U19430 ( .IN1(n18277), .IN2(n18278), .Q(n18270) );
  XOR2X1 U19431 ( .IN1(n9722), .IN2(n10128), .Q(n18278) );
  NOR2X0 U19432 ( .IN1(n4836), .IN2(n17859), .QN(n18277) );
  NAND2X0 U19433 ( .IN1(n18279), .IN2(n18280), .QN(g24255) );
  NAND2X0 U19434 ( .IN1(n13309), .IN2(g17423), .QN(n18280) );
  INVX0 U19435 ( .INP(n17853), .ZN(n13309) );
  NOR2X0 U19436 ( .IN1(n18281), .IN2(n18282), .QN(n18279) );
  NOR2X0 U19437 ( .IN1(n5755), .IN2(n10355), .QN(n18282) );
  NOR2X0 U19438 ( .IN1(n10474), .IN2(n18283), .QN(n18281) );
  NAND2X0 U19439 ( .IN1(n9735), .IN2(g10527), .QN(n18283) );
  NOR2X0 U19440 ( .IN1(n18284), .IN2(n18285), .QN(g24254) );
  NAND2X0 U19441 ( .IN1(n9737), .IN2(n9736), .QN(n18285) );
  NAND2X0 U19442 ( .IN1(n18286), .IN2(n9735), .QN(n18284) );
  NOR2X0 U19443 ( .IN1(n10474), .IN2(n18287), .QN(n18286) );
  NOR2X0 U19444 ( .IN1(n17822), .IN2(n18288), .QN(n18287) );
  NAND2X0 U19445 ( .IN1(n18289), .IN2(g1554), .QN(n18288) );
  OR2X1 U19446 ( .IN1(n17859), .IN2(n4836), .Q(n18289) );
  NAND2X0 U19447 ( .IN1(n5466), .IN2(n5322), .QN(n4836) );
  NAND2X0 U19448 ( .IN1(n16990), .IN2(n15501), .QN(n17859) );
  NAND2X0 U19449 ( .IN1(n5616), .IN2(n10128), .QN(n15501) );
  INVX0 U19450 ( .INP(n16993), .ZN(n16990) );
  XNOR2X1 U19451 ( .IN1(g1339), .IN2(test_so68), .Q(n16993) );
  NAND2X0 U19452 ( .IN1(n18260), .IN2(g1564), .QN(n17822) );
  NOR2X0 U19453 ( .IN1(n5546), .IN2(n10067), .QN(n18260) );
  NAND2X0 U19454 ( .IN1(n18290), .IN2(n18291), .QN(g24253) );
  NAND2X0 U19455 ( .IN1(n10500), .IN2(g1306), .QN(n18291) );
  NAND2X0 U19456 ( .IN1(n18292), .IN2(n10380), .QN(n18290) );
  NAND2X0 U19457 ( .IN1(n18293), .IN2(n18294), .QN(n18292) );
  NAND2X0 U19458 ( .IN1(n5302), .IN2(g1532), .QN(n18294) );
  NAND2X0 U19459 ( .IN1(g7946), .IN2(g1521), .QN(n18293) );
  NAND2X0 U19460 ( .IN1(n18295), .IN2(n18296), .QN(g24252) );
  NAND2X0 U19461 ( .IN1(test_so49), .IN2(n10515), .QN(n18296) );
  NAND2X0 U19462 ( .IN1(n18297), .IN2(n10380), .QN(n18295) );
  NAND2X0 U19463 ( .IN1(n18298), .IN2(n18299), .QN(n18297) );
  NAND2X0 U19464 ( .IN1(n5302), .IN2(g1521), .QN(n18299) );
  NAND2X0 U19465 ( .IN1(g7946), .IN2(g1339), .QN(n18298) );
  NAND2X0 U19466 ( .IN1(n18300), .IN2(n18301), .QN(g24251) );
  NAND2X0 U19467 ( .IN1(n16135), .IN2(g1442), .QN(n18301) );
  NAND2X0 U19468 ( .IN1(test_so12), .IN2(n17843), .QN(n18300) );
  NAND2X0 U19469 ( .IN1(n18302), .IN2(n18303), .QN(g24250) );
  NAND2X0 U19470 ( .IN1(test_so12), .IN2(n16135), .QN(n18303) );
  INVX0 U19471 ( .INP(n17843), .ZN(n16135) );
  NAND2X0 U19472 ( .IN1(n17843), .IN2(g1489), .QN(n18302) );
  NAND2X0 U19473 ( .IN1(n18304), .IN2(n18305), .QN(g24249) );
  NAND2X0 U19474 ( .IN1(n16160), .IN2(n16143), .QN(n18305) );
  INVX0 U19475 ( .INP(n17841), .ZN(n16143) );
  NOR2X0 U19476 ( .IN1(n10474), .IN2(g1442), .QN(n16160) );
  NAND2X0 U19477 ( .IN1(n18306), .IN2(g1489), .QN(n18304) );
  NAND2X0 U19478 ( .IN1(n17843), .IN2(n18307), .QN(n18306) );
  OR2X1 U19479 ( .IN1(n10457), .IN2(test_so12), .Q(n18307) );
  NAND2X0 U19480 ( .IN1(n17841), .IN2(n10380), .QN(n17843) );
  NAND2X0 U19481 ( .IN1(n18308), .IN2(n5364), .QN(n17841) );
  NOR2X0 U19482 ( .IN1(test_so49), .IN2(n9745), .QN(n18308) );
  NAND2X0 U19483 ( .IN1(n18309), .IN2(n18310), .QN(g24248) );
  XNOR2X1 U19484 ( .IN1(n9753), .IN2(n18311), .Q(n18310) );
  NAND2X0 U19485 ( .IN1(n5655), .IN2(n10381), .QN(n18311) );
  NOR2X0 U19486 ( .IN1(n18312), .IN2(n18313), .QN(n18309) );
  AND2X1 U19487 ( .IN1(n10366), .IN2(n5401), .Q(n18313) );
  NOR2X0 U19488 ( .IN1(n9966), .IN2(n17853), .QN(n18312) );
  NOR2X0 U19489 ( .IN1(g1249), .IN2(n17853), .QN(g24247) );
  NAND2X0 U19490 ( .IN1(n10368), .IN2(g12923), .QN(n17853) );
  NAND2X0 U19491 ( .IN1(n18314), .IN2(n18315), .QN(g24246) );
  NAND2X0 U19492 ( .IN1(n18316), .IN2(n10068), .QN(n18315) );
  NOR2X0 U19493 ( .IN1(n18317), .IN2(n18318), .QN(n18314) );
  NOR2X0 U19494 ( .IN1(n5547), .IN2(n10355), .QN(n18318) );
  NOR2X0 U19495 ( .IN1(n10474), .IN2(n18319), .QN(n18317) );
  OR2X1 U19496 ( .IN1(n18316), .IN2(n10068), .Q(n18319) );
  NAND2X0 U19497 ( .IN1(n18320), .IN2(n18321), .QN(g24245) );
  NAND2X0 U19498 ( .IN1(n10500), .IN2(g30332), .QN(n18321) );
  XOR2X1 U19499 ( .IN1(n18322), .IN2(n10069), .Q(g24244) );
  NAND2X0 U19500 ( .IN1(n10368), .IN2(g1205), .QN(n18322) );
  NAND2X0 U19501 ( .IN1(n18320), .IN2(n18323), .QN(g24243) );
  OR2X1 U19502 ( .IN1(n10308), .IN2(n9721), .Q(n18323) );
  NAND2X0 U19503 ( .IN1(n18324), .IN2(n18325), .QN(g24242) );
  NAND2X0 U19504 ( .IN1(n10368), .IN2(g29215), .QN(n18325) );
  NAND2X0 U19505 ( .IN1(test_so76), .IN2(n10516), .QN(n18324) );
  XOR2X1 U19506 ( .IN1(n18326), .IN2(n5622), .Q(g24241) );
  NAND2X0 U19507 ( .IN1(n18327), .IN2(n10381), .QN(n18326) );
  NAND2X0 U19508 ( .IN1(n18328), .IN2(n18329), .QN(g24240) );
  NAND2X0 U19509 ( .IN1(n10500), .IN2(g996), .QN(n18329) );
  NAND2X0 U19510 ( .IN1(n18330), .IN2(n10381), .QN(n18328) );
  XOR2X1 U19511 ( .IN1(n18327), .IN2(n18331), .Q(n18330) );
  NOR2X0 U19512 ( .IN1(g13259), .IN2(n18332), .QN(n18331) );
  NAND2X0 U19513 ( .IN1(n9638), .IN2(n18333), .QN(n18332) );
  INVX0 U19514 ( .INP(n17913), .ZN(n18333) );
  NAND2X0 U19515 ( .IN1(n18334), .IN2(n5392), .QN(n17913) );
  NOR2X0 U19516 ( .IN1(g990), .IN2(g7916), .QN(n18334) );
  AND2X1 U19517 ( .IN1(n18335), .IN2(n17384), .Q(n18327) );
  INVX0 U19518 ( .INP(n17919), .ZN(n17384) );
  NOR2X0 U19519 ( .IN1(n4837), .IN2(n18336), .QN(n18335) );
  XOR2X1 U19520 ( .IN1(n9721), .IN2(g979), .Q(n18336) );
  NAND2X0 U19521 ( .IN1(n18337), .IN2(n18338), .QN(g24239) );
  NAND2X0 U19522 ( .IN1(n13328), .IN2(g17400), .QN(n18338) );
  INVX0 U19523 ( .INP(n18320), .ZN(n13328) );
  NOR2X0 U19524 ( .IN1(n18339), .IN2(n18340), .QN(n18337) );
  NOR2X0 U19525 ( .IN1(n5756), .IN2(n10354), .QN(n18340) );
  NOR2X0 U19526 ( .IN1(n10479), .IN2(n18341), .QN(n18339) );
  NAND2X0 U19527 ( .IN1(n9724), .IN2(g10500), .QN(n18341) );
  NOR2X0 U19528 ( .IN1(n18342), .IN2(n18343), .QN(g24238) );
  NAND2X0 U19529 ( .IN1(n9715), .IN2(n9724), .QN(n18343) );
  NAND2X0 U19530 ( .IN1(n18344), .IN2(n18345), .QN(n18342) );
  NAND2X0 U19531 ( .IN1(n18346), .IN2(test_so76), .QN(n18345) );
  NOR2X0 U19532 ( .IN1(n18347), .IN2(n17887), .QN(n18346) );
  NAND2X0 U19533 ( .IN1(n18316), .IN2(g1221), .QN(n17887) );
  NOR2X0 U19534 ( .IN1(n5547), .IN2(n10069), .QN(n18316) );
  NOR2X0 U19535 ( .IN1(n4837), .IN2(n17919), .QN(n18347) );
  NAND2X0 U19536 ( .IN1(n17013), .IN2(n15542), .QN(n17919) );
  NAND2X0 U19537 ( .IN1(n5622), .IN2(n5320), .QN(n15542) );
  XNOR2X1 U19538 ( .IN1(g979), .IN2(n9757), .Q(n17013) );
  NAND2X0 U19539 ( .IN1(n5321), .IN2(n10152), .QN(n4837) );
  NOR2X0 U19540 ( .IN1(test_so44), .IN2(n10463), .QN(n18344) );
  NAND2X0 U19541 ( .IN1(n18348), .IN2(n18349), .QN(g24237) );
  NAND2X0 U19542 ( .IN1(n10500), .IN2(g962), .QN(n18349) );
  NAND2X0 U19543 ( .IN1(n18350), .IN2(n10382), .QN(n18348) );
  NAND2X0 U19544 ( .IN1(n18351), .IN2(n18352), .QN(n18350) );
  NAND2X0 U19545 ( .IN1(n5304), .IN2(g1189), .QN(n18352) );
  NAND2X0 U19546 ( .IN1(g7916), .IN2(g1178), .QN(n18351) );
  NAND2X0 U19547 ( .IN1(n18353), .IN2(n18354), .QN(g24236) );
  NAND2X0 U19548 ( .IN1(n10499), .IN2(g1183), .QN(n18354) );
  NAND2X0 U19549 ( .IN1(n18355), .IN2(n10382), .QN(n18353) );
  NAND2X0 U19550 ( .IN1(n18356), .IN2(n18357), .QN(n18355) );
  NAND2X0 U19551 ( .IN1(n5304), .IN2(g1178), .QN(n18357) );
  NAND2X0 U19552 ( .IN1(g7916), .IN2(g996), .QN(n18356) );
  NAND2X0 U19553 ( .IN1(n18358), .IN2(n18359), .QN(g24235) );
  NAND2X0 U19554 ( .IN1(test_so7), .IN2(n16188), .QN(n18359) );
  NAND2X0 U19555 ( .IN1(n17907), .IN2(g1152), .QN(n18358) );
  NAND2X0 U19556 ( .IN1(n18360), .IN2(n18361), .QN(g24234) );
  NAND2X0 U19557 ( .IN1(n16188), .IN2(g1152), .QN(n18361) );
  INVX0 U19558 ( .INP(n17907), .ZN(n16188) );
  NAND2X0 U19559 ( .IN1(n17907), .IN2(g1146), .QN(n18360) );
  NAND2X0 U19560 ( .IN1(n18362), .IN2(n18363), .QN(g24233) );
  NAND2X0 U19561 ( .IN1(n16213), .IN2(n16196), .QN(n18363) );
  INVX0 U19562 ( .INP(n17905), .ZN(n16196) );
  NOR2X0 U19563 ( .IN1(test_so7), .IN2(n10462), .QN(n16213) );
  NAND2X0 U19564 ( .IN1(n18364), .IN2(g1146), .QN(n18362) );
  NAND2X0 U19565 ( .IN1(n17907), .IN2(n18365), .QN(n18364) );
  NAND2X0 U19566 ( .IN1(n5618), .IN2(n10382), .QN(n18365) );
  NAND2X0 U19567 ( .IN1(n17905), .IN2(n10383), .QN(n17907) );
  NAND2X0 U19568 ( .IN1(n18366), .IN2(n5599), .QN(n17905) );
  NOR2X0 U19569 ( .IN1(n9744), .IN2(g1171), .QN(n18366) );
  NAND2X0 U19570 ( .IN1(n18367), .IN2(n18368), .QN(g24232) );
  XNOR2X1 U19571 ( .IN1(n9754), .IN2(n18369), .Q(n18368) );
  NAND2X0 U19572 ( .IN1(n5654), .IN2(n10383), .QN(n18369) );
  NOR2X0 U19573 ( .IN1(n18370), .IN2(n18371), .QN(n18367) );
  AND2X1 U19574 ( .IN1(n10366), .IN2(n5392), .Q(n18371) );
  NOR2X0 U19575 ( .IN1(n9967), .IN2(n18320), .QN(n18370) );
  NOR2X0 U19576 ( .IN1(g904), .IN2(n18320), .QN(g24231) );
  NAND2X0 U19577 ( .IN1(n10369), .IN2(g12919), .QN(n18320) );
  NAND2X0 U19578 ( .IN1(n18372), .IN2(n18373), .QN(g24216) );
  NAND2X0 U19579 ( .IN1(n16273), .IN2(g847), .QN(n18373) );
  NAND2X0 U19580 ( .IN1(n17036), .IN2(g854), .QN(n18372) );
  NAND2X0 U19581 ( .IN1(n18374), .IN2(n18375), .QN(g24215) );
  NAND2X0 U19582 ( .IN1(n18376), .IN2(g837), .QN(n18375) );
  NAND2X0 U19583 ( .IN1(n17036), .IN2(n18377), .QN(n18376) );
  NAND2X0 U19584 ( .IN1(n18378), .IN2(n18379), .QN(n18377) );
  NAND2X0 U19585 ( .IN1(g847), .IN2(g812), .QN(n18379) );
  NOR2X0 U19586 ( .IN1(n10467), .IN2(n18380), .QN(n18378) );
  NOR2X0 U19587 ( .IN1(n5728), .IN2(n10065), .QN(n18380) );
  NAND2X0 U19588 ( .IN1(n18381), .IN2(g703), .QN(n18374) );
  NAND2X0 U19589 ( .IN1(n18382), .IN2(n10384), .QN(n18381) );
  NAND2X0 U19590 ( .IN1(n5562), .IN2(n17445), .QN(n18382) );
  NOR2X0 U19591 ( .IN1(n16280), .IN2(n5709), .QN(n17445) );
  NAND2X0 U19592 ( .IN1(n18383), .IN2(n18384), .QN(g24214) );
  NAND2X0 U19593 ( .IN1(n18385), .IN2(g703), .QN(n18384) );
  NAND2X0 U19594 ( .IN1(n17440), .IN2(n18386), .QN(n18385) );
  OR2X1 U19595 ( .IN1(n17438), .IN2(n10457), .Q(n18386) );
  NOR2X0 U19596 ( .IN1(n5733), .IN2(n5562), .QN(n17438) );
  AND2X1 U19597 ( .IN1(n17036), .IN2(n18387), .Q(n17440) );
  NAND2X0 U19598 ( .IN1(n5709), .IN2(n10384), .QN(n18387) );
  NOR2X0 U19599 ( .IN1(n18388), .IN2(n18389), .QN(n18383) );
  NOR2X0 U19600 ( .IN1(g847), .IN2(n18390), .QN(n18389) );
  NAND2X0 U19601 ( .IN1(n18391), .IN2(n18392), .QN(n18390) );
  NOR2X0 U19602 ( .IN1(n5826), .IN2(n5822), .QN(n18392) );
  NOR2X0 U19603 ( .IN1(n5422), .IN2(n18393), .QN(n18391) );
  NOR2X0 U19604 ( .IN1(n5709), .IN2(n10354), .QN(n18388) );
  OR2X1 U19605 ( .IN1(n18394), .IN2(g24212), .Q(g24213) );
  NOR2X0 U19606 ( .IN1(n9678), .IN2(n10352), .QN(n18394) );
  NAND2X0 U19607 ( .IN1(n18395), .IN2(n18396), .QN(g24211) );
  NAND2X0 U19608 ( .IN1(n2404), .IN2(n18397), .QN(n18396) );
  OR2X1 U19609 ( .IN1(test_so41), .IN2(n5520), .Q(n18397) );
  OR2X1 U19610 ( .IN1(n10307), .IN2(n5492), .Q(n18395) );
  NOR2X0 U19611 ( .IN1(n14124), .IN2(n18398), .QN(g24210) );
  NAND2X0 U19612 ( .IN1(n18399), .IN2(n10381), .QN(n18398) );
  NAND2X0 U19613 ( .IN1(n18400), .IN2(n18401), .QN(n18399) );
  OR2X1 U19614 ( .IN1(n10136), .IN2(n15569), .Q(n18401) );
  NOR2X0 U19615 ( .IN1(g168), .IN2(g174), .QN(n15569) );
  NAND2X0 U19616 ( .IN1(g174), .IN2(g168), .QN(n18400) );
  NAND2X0 U19617 ( .IN1(n17476), .IN2(g203), .QN(n14124) );
  INVX0 U19618 ( .INP(n17088), .ZN(n17476) );
  NAND2X0 U19619 ( .IN1(n5548), .IN2(g518), .QN(n17088) );
  NAND2X0 U19620 ( .IN1(n18402), .IN2(n18403), .QN(g24209) );
  NAND2X0 U19621 ( .IN1(n16273), .IN2(g417), .QN(n18403) );
  NAND2X0 U19622 ( .IN1(n16277), .IN2(g446), .QN(n18402) );
  INVX0 U19623 ( .INP(n18393), .ZN(n16277) );
  NAND2X0 U19624 ( .IN1(n18404), .IN2(n18405), .QN(g24208) );
  NAND2X0 U19625 ( .IN1(n10499), .IN2(g424), .QN(n18405) );
  NOR2X0 U19626 ( .IN1(n18406), .IN2(n18407), .QN(n18404) );
  NOR2X0 U19627 ( .IN1(n6008), .IN2(n18393), .QN(n18407) );
  NOR2X0 U19628 ( .IN1(n9611), .IN2(n17036), .QN(n18406) );
  NAND2X0 U19629 ( .IN1(n18408), .IN2(n18409), .QN(g24207) );
  NAND2X0 U19630 ( .IN1(n16273), .IN2(g441), .QN(n18409) );
  OR2X1 U19631 ( .IN1(n16273), .IN2(n9611), .Q(n18408) );
  NAND2X0 U19632 ( .IN1(n18410), .IN2(n18411), .QN(g24206) );
  NAND2X0 U19633 ( .IN1(n16273), .IN2(g437), .QN(n18411) );
  NAND2X0 U19634 ( .IN1(n17036), .IN2(g441), .QN(n18410) );
  NAND2X0 U19635 ( .IN1(n18412), .IN2(n18413), .QN(g24205) );
  NAND2X0 U19636 ( .IN1(n10499), .IN2(g437), .QN(n18413) );
  NOR2X0 U19637 ( .IN1(n18414), .IN2(n18415), .QN(n18412) );
  NOR2X0 U19638 ( .IN1(n9783), .IN2(n18393), .QN(n18415) );
  AND2X1 U19639 ( .IN1(n16273), .IN2(test_so23), .Q(n18414) );
  NAND2X0 U19640 ( .IN1(n18416), .IN2(n18417), .QN(g24204) );
  NAND2X0 U19641 ( .IN1(n16273), .IN2(g429), .QN(n18417) );
  NAND2X0 U19642 ( .IN1(test_so23), .IN2(n17036), .QN(n18416) );
  NAND2X0 U19643 ( .IN1(n18418), .IN2(n18419), .QN(g24203) );
  NAND2X0 U19644 ( .IN1(n16273), .IN2(g401), .QN(n18419) );
  NAND2X0 U19645 ( .IN1(n17036), .IN2(g429), .QN(n18418) );
  NAND2X0 U19646 ( .IN1(n18420), .IN2(n18421), .QN(g24202) );
  NAND2X0 U19647 ( .IN1(n16273), .IN2(g424), .QN(n18421) );
  NAND2X0 U19648 ( .IN1(n17036), .IN2(g411), .QN(n18420) );
  NAND2X0 U19649 ( .IN1(n18422), .IN2(n18423), .QN(g24201) );
  NAND2X0 U19650 ( .IN1(n16273), .IN2(g405), .QN(n18423) );
  INVX0 U19651 ( .INP(n17036), .ZN(n16273) );
  NAND2X0 U19652 ( .IN1(n17036), .IN2(g392), .QN(n18422) );
  NAND2X0 U19653 ( .IN1(n18424), .IN2(n18425), .QN(g24200) );
  NAND2X0 U19654 ( .IN1(n10499), .IN2(g401), .QN(n18425) );
  NOR2X0 U19655 ( .IN1(n18426), .IN2(n18427), .QN(n18424) );
  NOR2X0 U19656 ( .IN1(n9778), .IN2(n17036), .QN(n18427) );
  NAND2X0 U19657 ( .IN1(n10377), .IN2(n16280), .QN(n17036) );
  INVX0 U19658 ( .INP(n4948), .ZN(n16280) );
  NOR2X0 U19659 ( .IN1(n18393), .IN2(n18428), .QN(n18426) );
  NAND2X0 U19660 ( .IN1(n5821), .IN2(g854), .QN(n18428) );
  NAND2X0 U19661 ( .IN1(n4948), .IN2(n10383), .QN(n18393) );
  NOR2X0 U19662 ( .IN1(g22), .IN2(g25), .QN(g23190) );
  NAND2X0 U19663 ( .IN1(n18429), .IN2(n18430), .QN(g21901) );
  OR2X1 U19664 ( .IN1(n10307), .IN2(n10087), .Q(n18430) );
  NAND2X0 U19665 ( .IN1(n18431), .IN2(n10384), .QN(n18429) );
  NAND2X0 U19666 ( .IN1(n18432), .IN2(n18433), .QN(n18431) );
  NAND2X0 U19667 ( .IN1(n5694), .IN2(g4180), .QN(n18433) );
  NAND2X0 U19668 ( .IN1(n5380), .IN2(n18434), .QN(n18432) );
  NAND2X0 U19669 ( .IN1(n5694), .IN2(n18435), .QN(n18434) );
  NAND2X0 U19670 ( .IN1(n18436), .IN2(n18437), .QN(n18435) );
  NOR2X0 U19671 ( .IN1(n18438), .IN2(n18439), .QN(n18437) );
  NAND2X0 U19672 ( .IN1(DFF_480_n1), .IN2(DFF_909_n1), .QN(n18439) );
  NAND2X0 U19673 ( .IN1(n9765), .IN2(DFF_1234_n1), .QN(n18438) );
  NOR2X0 U19674 ( .IN1(g8787), .IN2(n18440), .QN(n18436) );
  NAND2X0 U19675 ( .IN1(n9767), .IN2(n9766), .QN(n18440) );
  NAND2X0 U19676 ( .IN1(n18441), .IN2(n18442), .QN(g21900) );
  OR2X1 U19677 ( .IN1(n10307), .IN2(n9706), .Q(n18442) );
  NAND2X0 U19678 ( .IN1(n18443), .IN2(n10384), .QN(n18441) );
  NOR2X0 U19679 ( .IN1(g10122_Tj), .IN2(g4297), .QN(n18443) );
  XOR2X1 U19680 ( .IN1(n18444), .IN2(n10101), .Q(g21899) );
  NAND2X0 U19681 ( .IN1(n10374), .IN2(g9019), .QN(n18444) );
  NAND2X0 U19682 ( .IN1(n18445), .IN2(n18446), .QN(g21898) );
  NAND2X0 U19683 ( .IN1(n10101), .IN2(n10386), .QN(n18446) );
  OR2X1 U19684 ( .IN1(n10306), .IN2(n9725), .Q(n18445) );
  XOR2X1 U19685 ( .IN1(n18447), .IN2(n10102), .Q(g21897) );
  NAND2X0 U19686 ( .IN1(n10372), .IN2(g8839), .QN(n18447) );
  NAND2X0 U19687 ( .IN1(n18448), .IN2(n18449), .QN(g21896) );
  NAND2X0 U19688 ( .IN1(n10102), .IN2(n10386), .QN(n18449) );
  NAND2X0 U19689 ( .IN1(n10499), .IN2(g4245), .QN(n18448) );
  NAND2X0 U19690 ( .IN1(n18450), .IN2(n18451), .QN(g21895) );
  NAND2X0 U19691 ( .IN1(n18452), .IN2(g4264), .QN(n18451) );
  NAND2X0 U19692 ( .IN1(n18453), .IN2(n10381), .QN(n18452) );
  NAND2X0 U19693 ( .IN1(n5763), .IN2(g4258), .QN(n18453) );
  OR2X1 U19694 ( .IN1(n18181), .IN2(n5763), .Q(n18450) );
  NOR2X0 U19695 ( .IN1(g21893), .IN2(n18454), .QN(n18181) );
  NOR2X0 U19696 ( .IN1(g4264), .IN2(n10463), .QN(n18454) );
  NAND2X0 U19697 ( .IN1(n18455), .IN2(n18456), .QN(g21894) );
  NAND2X0 U19698 ( .IN1(n18457), .IN2(g4258), .QN(n18456) );
  NAND2X0 U19699 ( .IN1(n10368), .IN2(g4264), .QN(n18457) );
  NAND2X0 U19700 ( .IN1(g21893), .IN2(g4264), .QN(n18455) );
  NOR2X0 U19701 ( .IN1(g4258), .IN2(n10463), .QN(g21893) );
  NAND2X0 U19702 ( .IN1(n18458), .IN2(n18459), .QN(g21892) );
  NAND2X0 U19703 ( .IN1(n9706), .IN2(n10378), .QN(n18459) );
  NAND2X0 U19704 ( .IN1(n10498), .IN2(g4273), .QN(n18458) );
  NAND2X0 U19705 ( .IN1(n18460), .IN2(n18461), .QN(g21891) );
  NAND2X0 U19706 ( .IN1(n10511), .IN2(g4180), .QN(n18461) );
  NAND2X0 U19707 ( .IN1(n18186), .IN2(n10378), .QN(n18460) );
  NAND2X0 U19708 ( .IN1(n18462), .IN2(n18463), .QN(n18186) );
  NAND2X0 U19709 ( .IN1(n10073), .IN2(g4253), .QN(n18463) );
  NAND2X0 U19710 ( .IN1(n5484), .IN2(n10072), .QN(n18462) );
  NOR2X0 U19711 ( .IN1(n10357), .IN2(DFF_1381_n1), .QN(g21727) );
  NOR2X0 U19712 ( .IN1(n5750), .IN2(n10346), .QN(g18597) );
  INVX0 U19713 ( .INP(g5), .ZN(g12833) );
  OR2X1 U5116_U1 ( .IN1(g34783), .IN2(n2730), .Q(g34221) );
  OR2X1 U5126_U1 ( .IN1(n4836), .IN2(n4896), .Q(n4895) );
  OR2X1 U5127_U1 ( .IN1(n4837), .IN2(n4921), .Q(n4920) );
  OR2X1 U5128_U1 ( .IN1(n2787), .IN2(n4411), .Q(n5045) );
  OR2X1 U5129_U1 ( .IN1(g559), .IN2(g9048), .Q(n4959) );
  INVX0 U5353_U2 ( .INP(n5960), .ZN(U5353_n1) );
  NOR2X0 U5353_U1 ( .IN1(n10113), .IN2(U5353_n1), .QN(n4689) );
  INVX0 U5355_U2 ( .INP(n5961), .ZN(U5355_n1) );
  NOR2X0 U5355_U1 ( .IN1(n10108), .IN2(U5355_n1), .QN(n4708) );
  INVX0 U5961_U2 ( .INP(n787), .ZN(U5961_n1) );
  NOR2X0 U5961_U1 ( .IN1(n3589), .IN2(U5961_n1), .QN(n3595) );
  INVX0 U5962_U2 ( .INP(n780), .ZN(U5962_n1) );
  NOR2X0 U5962_U1 ( .IN1(n3570), .IN2(U5962_n1), .QN(n3576) );
  INVX0 U5963_U2 ( .INP(n333), .ZN(U5963_n1) );
  NOR2X0 U5963_U1 ( .IN1(n3513), .IN2(U5963_n1), .QN(n3519) );
  INVX0 U5964_U2 ( .INP(n783), .ZN(U5964_n1) );
  NOR2X0 U5964_U1 ( .IN1(n3624), .IN2(U5964_n1), .QN(n3630) );
  INVX0 U5965_U2 ( .INP(n380), .ZN(U5965_n1) );
  NOR2X0 U5965_U1 ( .IN1(n3551), .IN2(U5965_n1), .QN(n3557) );
  INVX0 U5966_U2 ( .INP(n8), .ZN(U5966_n1) );
  NOR2X0 U5966_U1 ( .IN1(n3642), .IN2(U5966_n1), .QN(n3648) );
  INVX0 U5967_U2 ( .INP(n408), .ZN(U5967_n1) );
  NOR2X0 U5967_U1 ( .IN1(n3532), .IN2(U5967_n1), .QN(n3538) );
  INVX0 U5968_U2 ( .INP(n3611), .ZN(U5968_n1) );
  NOR2X0 U5968_U1 ( .IN1(n3607), .IN2(U5968_n1), .QN(n3613) );
  INVX0 U6100_U2 ( .INP(n3635), .ZN(U6100_n1) );
  NOR2X0 U6100_U1 ( .IN1(n10464), .IN2(U6100_n1), .QN(n4888) );
  INVX0 U6211_U2 ( .INP(n3623), .ZN(U6211_n1) );
  NOR2X0 U6211_U1 ( .IN1(n1282), .IN2(U6211_n1), .QN(n3622) );
  INVX0 U6212_U2 ( .INP(n3587), .ZN(U6212_n1) );
  NOR2X0 U6212_U1 ( .IN1(n3588), .IN2(U6212_n1), .QN(n3586) );
  INVX0 U6213_U2 ( .INP(n3605), .ZN(U6213_n1) );
  NOR2X0 U6213_U1 ( .IN1(n3606), .IN2(U6213_n1), .QN(n3604) );
  INVX0 U6214_U2 ( .INP(n3568), .ZN(U6214_n1) );
  NOR2X0 U6214_U1 ( .IN1(n3569), .IN2(U6214_n1), .QN(n3567) );
  INVX0 U6215_U2 ( .INP(n3549), .ZN(U6215_n1) );
  NOR2X0 U6215_U1 ( .IN1(n3550), .IN2(U6215_n1), .QN(n3548) );
  INVX0 U6216_U2 ( .INP(n3512), .ZN(U6216_n1) );
  NOR2X0 U6216_U1 ( .IN1(n3006), .IN2(U6216_n1), .QN(n3511) );
  INVX0 U6217_U2 ( .INP(n3531), .ZN(U6217_n1) );
  NOR2X0 U6217_U1 ( .IN1(n3007), .IN2(U6217_n1), .QN(n3530) );
  INVX0 U6218_U2 ( .INP(n3641), .ZN(U6218_n1) );
  NOR2X0 U6218_U1 ( .IN1(n3003), .IN2(U6218_n1), .QN(n3640) );
  INVX0 U6279_U2 ( .INP(n4537), .ZN(U6279_n1) );
  NOR2X0 U6279_U1 ( .IN1(n5337), .IN2(U6279_n1), .QN(n4201) );
  INVX0 U6280_U2 ( .INP(n4201), .ZN(U6280_n1) );
  NOR2X0 U6280_U1 ( .IN1(n5336), .IN2(U6280_n1), .QN(n3745) );
  INVX0 U6281_U2 ( .INP(n3745), .ZN(U6281_n1) );
  NOR2X0 U6281_U1 ( .IN1(n5294), .IN2(U6281_n1), .QN(n3684) );
  INVX0 U6282_U2 ( .INP(n3684), .ZN(U6282_n1) );
  NOR2X0 U6282_U1 ( .IN1(n5552), .IN2(U6282_n1), .QN(n3274) );
  INVX0 U6283_U2 ( .INP(n3274), .ZN(U6283_n1) );
  NOR2X0 U6283_U1 ( .IN1(n5472), .IN2(U6283_n1), .QN(n2982) );
  INVX0 U6284_U2 ( .INP(n2982), .ZN(U6284_n1) );
  NOR2X0 U6284_U1 ( .IN1(n5476), .IN2(U6284_n1), .QN(n2706) );
  INVX0 U6285_U2 ( .INP(n2706), .ZN(U6285_n1) );
  NOR2X0 U6285_U1 ( .IN1(n5550), .IN2(U6285_n1), .QN(n2649) );
  INVX0 U6286_U2 ( .INP(n2649), .ZN(U6286_n1) );
  NOR2X0 U6286_U1 ( .IN1(n5473), .IN2(U6286_n1), .QN(n2556) );
  INVX0 U6287_U2 ( .INP(n2556), .ZN(U6287_n1) );
  NOR2X0 U6287_U1 ( .IN1(n5475), .IN2(U6287_n1), .QN(n2509) );
  INVX0 U6288_U2 ( .INP(n2509), .ZN(U6288_n1) );
  NOR2X0 U6288_U1 ( .IN1(n5474), .IN2(U6288_n1), .QN(n2487) );
  INVX0 U6289_U2 ( .INP(n2487), .ZN(U6289_n1) );
  NOR2X0 U6289_U1 ( .IN1(n5339), .IN2(U6289_n1), .QN(n2427) );
  INVX0 U6290_U2 ( .INP(n2427), .ZN(U6290_n1) );
  NOR2X0 U6290_U1 ( .IN1(n5672), .IN2(U6290_n1), .QN(n2423) );
  INVX0 U6291_U2 ( .INP(n3), .ZN(U6291_n1) );
  NOR2X0 U6291_U1 ( .IN1(n5335), .IN2(U6291_n1), .QN(n4537) );
  INVX0 U6292_U2 ( .INP(n4959), .ZN(U6292_n1) );
  NOR2X0 U6292_U1 ( .IN1(n10465), .IN2(U6292_n1), .QN(n2421) );
  INVX0 U6338_U2 ( .INP(n4210), .ZN(U6338_n1) );
  NOR2X1 U6338_U1 ( .IN1(n10464), .IN2(U6338_n1), .QN(n3765) );
  INVX0 U6341_U2 ( .INP(n3765), .ZN(U6341_n1) );
  NOR2X0 U6341_U1 ( .IN1(n3479), .IN2(U6341_n1), .QN(n3951) );
  INVX0 U6342_U2 ( .INP(n3765), .ZN(U6342_n1) );
  NOR2X0 U6342_U1 ( .IN1(n3404), .IN2(U6342_n1), .QN(n3774) );
  INVX0 U6343_U2 ( .INP(n3765), .ZN(U6343_n1) );
  NOR2X0 U6343_U1 ( .IN1(n3424), .IN2(U6343_n1), .QN(n3842) );
  INVX0 U6344_U2 ( .INP(n3765), .ZN(U6344_n1) );
  NOR2X0 U6344_U1 ( .IN1(n3414), .IN2(U6344_n1), .QN(n3808) );
  INVX0 U6345_U2 ( .INP(n3765), .ZN(U6345_n1) );
  NOR2X0 U6345_U1 ( .IN1(n3444), .IN2(U6345_n1), .QN(n3908) );
  INVX0 U6346_U2 ( .INP(n3765), .ZN(U6346_n1) );
  NOR2X0 U6346_U1 ( .IN1(n3489), .IN2(U6346_n1), .QN(n3984) );
  INVX0 U6347_U2 ( .INP(n3765), .ZN(U6347_n1) );
  NOR2X0 U6347_U1 ( .IN1(n3434), .IN2(U6347_n1), .QN(n3875) );
  INVX0 U6348_U2 ( .INP(n3765), .ZN(U6348_n1) );
  NOR2X0 U6348_U1 ( .IN1(n3500), .IN2(U6348_n1), .QN(n4015) );
  INVX0 U6349_U2 ( .INP(n3765), .ZN(U6349_n1) );
  NOR2X0 U6349_U1 ( .IN1(n3446), .IN2(U6349_n1), .QN(n3914) );
  INVX0 U6350_U2 ( .INP(n3765), .ZN(U6350_n1) );
  NOR2X0 U6350_U1 ( .IN1(n3406), .IN2(U6350_n1), .QN(n3780) );
  INVX0 U6351_U2 ( .INP(n3765), .ZN(U6351_n1) );
  NOR2X0 U6351_U1 ( .IN1(n3481), .IN2(U6351_n1), .QN(n3957) );
  INVX0 U6352_U2 ( .INP(n3765), .ZN(U6352_n1) );
  NOR2X0 U6352_U1 ( .IN1(n3426), .IN2(U6352_n1), .QN(n3848) );
  INVX0 U6353_U2 ( .INP(n3765), .ZN(U6353_n1) );
  NOR2X0 U6353_U1 ( .IN1(n3491), .IN2(U6353_n1), .QN(n3990) );
  INVX0 U6354_U2 ( .INP(n3765), .ZN(U6354_n1) );
  NOR2X0 U6354_U1 ( .IN1(n3416), .IN2(U6354_n1), .QN(n3814) );
  INVX0 U6355_U2 ( .INP(n3765), .ZN(U6355_n1) );
  NOR2X0 U6355_U1 ( .IN1(n3436), .IN2(U6355_n1), .QN(n3881) );
  INVX0 U6356_U2 ( .INP(n3765), .ZN(U6356_n1) );
  NOR2X0 U6356_U1 ( .IN1(n3502), .IN2(U6356_n1), .QN(n4022) );
  INVX0 U6357_U2 ( .INP(n3765), .ZN(U6357_n1) );
  NOR2X0 U6357_U1 ( .IN1(n3501), .IN2(U6357_n1), .QN(n4027) );
  INVX0 U6358_U2 ( .INP(n3765), .ZN(U6358_n1) );
  NOR2X0 U6358_U1 ( .IN1(n3407), .IN2(U6358_n1), .QN(n3785) );
  INVX0 U6359_U2 ( .INP(n3765), .ZN(U6359_n1) );
  NOR2X0 U6359_U1 ( .IN1(n3482), .IN2(U6359_n1), .QN(n3962) );
  INVX0 U6360_U2 ( .INP(n3765), .ZN(U6360_n1) );
  NOR2X0 U6360_U1 ( .IN1(n3427), .IN2(U6360_n1), .QN(n3853) );
  INVX0 U6361_U2 ( .INP(n3765), .ZN(U6361_n1) );
  NOR2X0 U6361_U1 ( .IN1(n3437), .IN2(U6361_n1), .QN(n3886) );
  INVX0 U6362_U2 ( .INP(n3765), .ZN(U6362_n1) );
  NOR2X0 U6362_U1 ( .IN1(n3417), .IN2(U6362_n1), .QN(n3819) );
  INVX0 U6363_U2 ( .INP(n3765), .ZN(U6363_n1) );
  NOR2X0 U6363_U1 ( .IN1(n3492), .IN2(U6363_n1), .QN(n3995) );
  INVX0 U6364_U2 ( .INP(n3765), .ZN(U6364_n1) );
  NOR2X0 U6364_U1 ( .IN1(n3447), .IN2(U6364_n1), .QN(n3919) );
  INVX0 U6365_U2 ( .INP(n3682), .ZN(U6365_n1) );
  NOR2X0 U6365_U1 ( .IN1(n5471), .IN2(U6365_n1), .QN(n3272) );
  INVX0 U6366_U2 ( .INP(n3272), .ZN(U6366_n1) );
  NOR2X0 U6366_U1 ( .IN1(n5331), .IN2(U6366_n1), .QN(n2980) );
  INVX0 U6367_U2 ( .INP(n2980), .ZN(U6367_n1) );
  NOR2X0 U6367_U1 ( .IN1(n5332), .IN2(U6367_n1), .QN(n2704) );
  INVX0 U6368_U2 ( .INP(n2704), .ZN(U6368_n1) );
  NOR2X0 U6368_U1 ( .IN1(n5333), .IN2(U6368_n1), .QN(n2647) );
  INVX0 U6369_U2 ( .INP(n2647), .ZN(U6369_n1) );
  NOR2X0 U6369_U1 ( .IN1(n5334), .IN2(U6369_n1), .QN(n2554) );
  INVX0 U6370_U2 ( .INP(n2554), .ZN(U6370_n1) );
  NOR2X0 U6370_U1 ( .IN1(n5330), .IN2(U6370_n1), .QN(n2507) );
  INVX0 U6371_U2 ( .INP(n2507), .ZN(U6371_n1) );
  NOR2X0 U6371_U1 ( .IN1(n5551), .IN2(U6371_n1), .QN(n2485) );
  INVX0 U6372_U2 ( .INP(n2485), .ZN(U6372_n1) );
  NOR2X0 U6372_U1 ( .IN1(n5293), .IN2(U6372_n1), .QN(n2425) );
  INVX0 U6373_U2 ( .INP(n2425), .ZN(U6373_n1) );
  NOR2X0 U6373_U1 ( .IN1(n5292), .IN2(U6373_n1), .QN(n2419) );
  INVX0 U6374_U2 ( .INP(n3743), .ZN(U6374_n1) );
  NOR2X0 U6374_U1 ( .IN1(n5470), .IN2(U6374_n1), .QN(n3682) );
  INVX0 U6375_U2 ( .INP(n2419), .ZN(U6375_n1) );
  NOR2X0 U6375_U1 ( .IN1(n5291), .IN2(U6375_n1), .QN(n2405) );
  INVX0 U6417_U2 ( .INP(n4198), .ZN(U6417_n1) );
  NOR2X0 U6417_U1 ( .IN1(n10465), .IN2(U6417_n1), .QN(n2404) );
  INVX0 U6446_U2 ( .INP(g110), .ZN(U6446_n1) );
  NOR2X0 U6446_U1 ( .IN1(n1289), .IN2(U6446_n1), .QN(n3524) );
  INVX0 U6465_U2 ( .INP(n549), .ZN(U6465_n1) );
  NOR2X0 U6465_U1 ( .IN1(n5600), .IN2(U6465_n1), .QN(n4388) );
  INVX0 U6497_U2 ( .INP(n572), .ZN(U6497_n1) );
  NOR2X0 U6497_U1 ( .IN1(n3635), .IN2(U6497_n1), .QN(n3005) );
  INVX0 U6523_U2 ( .INP(n4946), .ZN(U6523_n1) );
  NOR2X0 U6523_U1 ( .IN1(n10465), .IN2(U6523_n1), .QN(n4945) );
  INVX0 U6542_U2 ( .INP(n572), .ZN(U6542_n1) );
  NOR2X0 U6542_U1 ( .IN1(n5300), .IN2(U6542_n1), .QN(n3525) );
  INVX0 U6552_U2 ( .INP(n3281), .ZN(U6552_n1) );
  NOR2X0 U6552_U1 ( .IN1(n5676), .IN2(U6552_n1), .QN(n3277) );
  INVX0 U6553_U2 ( .INP(n3276), .ZN(U6553_n1) );
  NOR2X0 U6553_U1 ( .IN1(n5680), .IN2(U6553_n1), .QN(n2989) );
  INVX0 U6554_U2 ( .INP(n3277), .ZN(U6554_n1) );
  NOR2X0 U6554_U1 ( .IN1(n5677), .IN2(U6554_n1), .QN(n2991) );
  INVX0 U6555_U2 ( .INP(n39), .ZN(U6555_n1) );
  NOR2X0 U6555_U1 ( .IN1(n5561), .IN2(U6555_n1), .QN(n3281) );
  INVX0 U6556_U2 ( .INP(n36), .ZN(U6556_n1) );
  NOR2X0 U6556_U1 ( .IN1(n5679), .IN2(U6556_n1), .QN(n3276) );
  INVX0 U6559_U2 ( .INP(n2991), .ZN(U6559_n1) );
  NOR2X0 U6559_U1 ( .IN1(n5678), .IN2(U6559_n1), .QN(n2710) );
  INVX0 U6560_U2 ( .INP(n2989), .ZN(U6560_n1) );
  NOR2X0 U6560_U1 ( .IN1(n5675), .IN2(U6560_n1), .QN(n2707) );
  INVX0 U6561_U2 ( .INP(n3174), .ZN(U6561_n1) );
  NOR2X0 U6561_U1 ( .IN1(n5327), .IN2(U6561_n1), .QN(n3116) );
  INVX0 U6570_U2 ( .INP(n3362), .ZN(U6570_n1) );
  NOR2X0 U6570_U1 ( .IN1(n5477), .IN2(U6570_n1), .QN(n2527) );
  INVX0 U6911_U2 ( .INP(n3115), .ZN(U6911_n1) );
  NOR2X0 U6911_U1 ( .IN1(n2726), .IN2(U6911_n1), .QN(n3111) );
  INVX0 U6912_U2 ( .INP(n3115), .ZN(U6912_n1) );
  NOR2X0 U6912_U1 ( .IN1(n2727), .IN2(U6912_n1), .QN(n3131) );
  INVX0 U6917_U2 ( .INP(n3933), .ZN(U6917_n1) );
  NOR2X0 U6917_U1 ( .IN1(n5350), .IN2(U6917_n1), .QN(n3799) );
  INVX0 U6926_U2 ( .INP(n3664), .ZN(U6926_n1) );
  NOR2X0 U6926_U1 ( .IN1(n5674), .IN2(U6926_n1), .QN(n3662) );
  INVX0 U6927_U2 ( .INP(n3673), .ZN(U6927_n1) );
  NOR2X0 U6927_U1 ( .IN1(n5673), .IN2(U6927_n1), .QN(n3671) );
  INVX0 U6929_U2 ( .INP(n3505), .ZN(U6929_n1) );
  NOR2X0 U6929_U1 ( .IN1(n3506), .IN2(U6929_n1), .QN(n2790) );
  INVX0 U6931_U2 ( .INP(n4490), .ZN(U6931_n1) );
  NOR2X0 U6931_U1 ( .IN1(n5554), .IN2(U6931_n1), .QN(n4178) );
  INVX0 U6932_U2 ( .INP(n4514), .ZN(U6932_n1) );
  NOR2X0 U6932_U1 ( .IN1(n5555), .IN2(U6932_n1), .QN(n4196) );
  INVX0 U6933_U2 ( .INP(n4178), .ZN(U6933_n1) );
  NOR2X0 U6933_U1 ( .IN1(n5558), .IN2(U6933_n1), .QN(n3736) );
  INVX0 U6934_U2 ( .INP(n4196), .ZN(U6934_n1) );
  NOR2X0 U6934_U1 ( .IN1(n5559), .IN2(U6934_n1), .QN(n3741) );
  INVX0 U6935_U2 ( .INP(n3736), .ZN(U6935_n1) );
  NOR2X0 U6935_U1 ( .IN1(n5553), .IN2(U6935_n1), .QN(n3664) );
  INVX0 U6936_U2 ( .INP(n3741), .ZN(U6936_n1) );
  NOR2X0 U6936_U1 ( .IN1(n5560), .IN2(U6936_n1), .QN(n3673) );
  INVX0 U6937_U2 ( .INP(n2601), .ZN(U6937_n1) );
  NOR2X0 U6937_U1 ( .IN1(n5303), .IN2(U6937_n1), .QN(n2598) );
  INVX0 U6938_U2 ( .INP(n870), .ZN(U6938_n1) );
  NOR2X0 U6938_U1 ( .IN1(n5556), .IN2(U6938_n1), .QN(n4490) );
  INVX0 U6939_U2 ( .INP(n195), .ZN(U6939_n1) );
  NOR2X0 U6939_U1 ( .IN1(n5557), .IN2(U6939_n1), .QN(n4514) );
  INVX0 U6940_U2 ( .INP(n4814), .ZN(U6940_n1) );
  NOR2X0 U6940_U1 ( .IN1(n5422), .IN2(U6940_n1), .QN(n4519) );
  INVX0 U6941_U2 ( .INP(n2607), .ZN(U6941_n1) );
  NOR2X0 U6941_U1 ( .IN1(n5323), .IN2(U6941_n1), .QN(n2594) );
  INVX0 U6944_U2 ( .INP(n3084), .ZN(U6944_n1) );
  NOR2X0 U6944_U1 ( .IN1(n5348), .IN2(U6944_n1), .QN(n3033) );
  INVX0 U6950_U2 ( .INP(n2598), .ZN(U6950_n1) );
  NOR2X0 U6950_U1 ( .IN1(n5365), .IN2(U6950_n1), .QN(n2590) );
  INVX0 U6954_U2 ( .INP(n490), .ZN(U6954_n1) );
  NOR2X0 U6954_U1 ( .IN1(n2727), .IN2(U6954_n1), .QN(n3125) );
  INVX0 U6955_U2 ( .INP(n475), .ZN(U6955_n1) );
  NOR2X0 U6955_U1 ( .IN1(n2726), .IN2(U6955_n1), .QN(n3105) );
  INVX0 U6956_U2 ( .INP(n3141), .ZN(U6956_n1) );
  NOR2X0 U6956_U1 ( .IN1(n3146), .IN2(U6956_n1), .QN(n3145) );
  INVX0 U6957_U2 ( .INP(n3160), .ZN(U6957_n1) );
  NOR2X0 U6957_U1 ( .IN1(n3165), .IN2(U6957_n1), .QN(n3164) );
  INVX0 U7174_U2 ( .INP(n2423), .ZN(U7174_n1) );
  NOR2X0 U7174_U1 ( .IN1(n5288), .IN2(U7174_n1), .QN(n2422) );
  INVX0 U7248_U2 ( .INP(n4172), .ZN(U7248_n1) );
  NOR2X0 U7248_U1 ( .IN1(g1536), .IN2(U7248_n1), .QN(n4173) );
  INVX0 U7249_U2 ( .INP(n4190), .ZN(U7249_n1) );
  NOR2X0 U7249_U1 ( .IN1(g1193), .IN2(U7249_n1), .QN(n4191) );
  INVX0 U7402_U2 ( .INP(n4034), .ZN(U7402_n1) );
  NOR2X0 U7402_U1 ( .IN1(n4020), .IN2(U7402_n1), .QN(n4037) );
  INVX0 U7405_U2 ( .INP(n4034), .ZN(U7405_n1) );
  NOR2X0 U7405_U1 ( .IN1(n4014), .IN2(U7405_n1), .QN(n4039) );
  INVX0 U7413_U2 ( .INP(n3969), .ZN(U7413_n1) );
  NOR2X0 U7413_U1 ( .IN1(n3947), .IN2(U7413_n1), .QN(n3972) );
  INVX0 U7416_U2 ( .INP(n3926), .ZN(U7416_n1) );
  NOR2X0 U7416_U1 ( .IN1(n3904), .IN2(U7416_n1), .QN(n3929) );
  INVX0 U7427_U2 ( .INP(n3860), .ZN(U7427_n1) );
  NOR2X0 U7427_U1 ( .IN1(n3838), .IN2(U7427_n1), .QN(n3863) );
  INVX0 U7438_U2 ( .INP(n4002), .ZN(U7438_n1) );
  NOR2X0 U7438_U1 ( .IN1(n3978), .IN2(U7438_n1), .QN(n4003) );
  INVX0 U7449_U2 ( .INP(n4034), .ZN(U7449_n1) );
  NOR2X0 U7449_U1 ( .IN1(n365), .IN2(U7449_n1), .QN(n4032) );
  INVX0 U7455_U2 ( .INP(n4034), .ZN(U7455_n1) );
  NOR2X0 U7455_U1 ( .IN1(n364), .IN2(U7455_n1), .QN(n4035) );
  INVX0 U7464_U2 ( .INP(n3792), .ZN(U7464_n1) );
  NOR2X0 U7464_U1 ( .IN1(n3773), .IN2(U7464_n1), .QN(n3797) );
  INVX0 U7467_U2 ( .INP(n3792), .ZN(U7467_n1) );
  NOR2X0 U7467_U1 ( .IN1(n3776), .IN2(U7467_n1), .QN(n3790) );
  INVX0 U7482_U2 ( .INP(n3792), .ZN(U7482_n1) );
  NOR2X0 U7482_U1 ( .IN1(n3770), .IN2(U7482_n1), .QN(n3795) );
  INVX0 U7492_U2 ( .INP(n3893), .ZN(U7492_n1) );
  NOR2X0 U7492_U1 ( .IN1(n3877), .IN2(U7492_n1), .QN(n3891) );
  INVX0 U7513_U2 ( .INP(n3826), .ZN(U7513_n1) );
  NOR2X0 U7513_U1 ( .IN1(n3802), .IN2(U7513_n1), .QN(n3827) );
  INVX0 U7516_U2 ( .INP(n3893), .ZN(U7516_n1) );
  NOR2X0 U7516_U1 ( .IN1(n3871), .IN2(U7516_n1), .QN(n3896) );
  INVX0 U7549_U2 ( .INP(n4002), .ZN(U7549_n1) );
  NOR2X0 U7549_U1 ( .IN1(n3983), .IN2(U7549_n1), .QN(n4007) );
  INVX0 U7561_U2 ( .INP(n3926), .ZN(U7561_n1) );
  NOR2X0 U7561_U1 ( .IN1(n3907), .IN2(U7561_n1), .QN(n3931) );
  INVX0 U7574_U2 ( .INP(n3792), .ZN(U7574_n1) );
  NOR2X0 U7574_U1 ( .IN1(n3768), .IN2(U7574_n1), .QN(n3793) );
  INVX0 U7577_U2 ( .INP(n3926), .ZN(U7577_n1) );
  NOR2X0 U7577_U1 ( .IN1(n3910), .IN2(U7577_n1), .QN(n3924) );
  INVX0 U7585_U2 ( .INP(n3826), .ZN(U7585_n1) );
  NOR2X0 U7585_U1 ( .IN1(n3807), .IN2(U7585_n1), .QN(n3831) );
  INVX0 U7595_U2 ( .INP(n3826), .ZN(U7595_n1) );
  NOR2X0 U7595_U1 ( .IN1(n3804), .IN2(U7595_n1), .QN(n3829) );
  INVX0 U7614_U2 ( .INP(n3926), .ZN(U7614_n1) );
  NOR2X0 U7614_U1 ( .IN1(n3902), .IN2(U7614_n1), .QN(n3927) );
  INVX0 U7621_U2 ( .INP(n3969), .ZN(U7621_n1) );
  NOR2X0 U7621_U1 ( .IN1(n3950), .IN2(U7621_n1), .QN(n3974) );
  INVX0 U7629_U2 ( .INP(n3893), .ZN(U7629_n1) );
  NOR2X0 U7629_U1 ( .IN1(n3874), .IN2(U7629_n1), .QN(n3898) );
  INVX0 U7636_U2 ( .INP(n3969), .ZN(U7636_n1) );
  NOR2X0 U7636_U1 ( .IN1(n3945), .IN2(U7636_n1), .QN(n3970) );
  INVX0 U7639_U2 ( .INP(n4002), .ZN(U7639_n1) );
  NOR2X0 U7639_U1 ( .IN1(n3986), .IN2(U7639_n1), .QN(n4000) );
  INVX0 U7649_U2 ( .INP(n3860), .ZN(U7649_n1) );
  NOR2X0 U7649_U1 ( .IN1(n3841), .IN2(U7649_n1), .QN(n3865) );
  INVX0 U7652_U2 ( .INP(n3860), .ZN(U7652_n1) );
  NOR2X0 U7652_U1 ( .IN1(n3836), .IN2(U7652_n1), .QN(n3861) );
  INVX0 U7668_U2 ( .INP(n3826), .ZN(U7668_n1) );
  NOR2X0 U7668_U1 ( .IN1(n3810), .IN2(U7668_n1), .QN(n3824) );
  INVX0 U7673_U2 ( .INP(n3893), .ZN(U7673_n1) );
  NOR2X0 U7673_U1 ( .IN1(n3869), .IN2(U7673_n1), .QN(n3894) );
  INVX0 U7690_U2 ( .INP(n3969), .ZN(U7690_n1) );
  NOR2X0 U7690_U1 ( .IN1(n3953), .IN2(U7690_n1), .QN(n3967) );
  INVX0 U7707_U2 ( .INP(n3860), .ZN(U7707_n1) );
  NOR2X0 U7707_U1 ( .IN1(n3844), .IN2(U7707_n1), .QN(n3858) );
  INVX0 U7712_U2 ( .INP(n4002), .ZN(U7712_n1) );
  NOR2X0 U7712_U1 ( .IN1(n3980), .IN2(U7712_n1), .QN(n4005) );
  INVX0 U7792_U2 ( .INP(g952), .ZN(U7792_n1) );
  NOR2X0 U7792_U1 ( .IN1(n10464), .IN2(U7792_n1), .QN(n2505) );
  INVX0 U7794_U2 ( .INP(g1296), .ZN(U7794_n1) );
  NOR2X0 U7794_U1 ( .IN1(n10464), .IN2(U7794_n1), .QN(n2499) );
  INVX0 U7895_U2 ( .INP(n2668), .ZN(U7895_n1) );
  NOR2X0 U7895_U1 ( .IN1(g113), .IN2(U7895_n1), .QN(n2760) );
  INVX0 U7897_U2 ( .INP(g6), .ZN(U7897_n1) );
  NOR2X0 U7897_U1 ( .IN1(g31), .IN2(U7897_n1), .QN(n3395) );
  INVX0 U7977_U2 ( .INP(g661), .ZN(U7977_n1) );
  NOR2X0 U7977_U1 ( .IN1(n10464), .IN2(U7977_n1), .QN(n4956) );
  INVX0 U8034_U2 ( .INP(n4723), .ZN(U8034_n1) );
  NOR2X0 U8034_U1 ( .IN1(n5612), .IN2(U8034_n1), .QN(n5026) );
  INVX0 U8036_U2 ( .INP(n3729), .ZN(U8036_n1) );
  NOR2X0 U8036_U1 ( .IN1(n5340), .IN2(U8036_n1), .QN(n3941) );
  INVX0 U8050_U2 ( .INP(n3660), .ZN(U8050_n1) );
  NOR2X0 U8050_U1 ( .IN1(g1367), .IN2(U8050_n1), .QN(n3733) );
  INVX0 U8055_U2 ( .INP(g1345), .ZN(U8055_n1) );
  NOR2X0 U8055_U1 ( .IN1(n10465), .IN2(U8055_n1), .QN(n4798) );
  INVX0 U8060_U2 ( .INP(g1002), .ZN(U8060_n1) );
  NOR2X0 U8060_U1 ( .IN1(n10464), .IN2(U8060_n1), .QN(n4805) );
  INVX0 U8070_U2 ( .INP(n3734), .ZN(U8070_n1) );
  NOR2X0 U8070_U1 ( .IN1(g1361), .IN2(U8070_n1), .QN(n4175) );
  INVX0 U8074_U2 ( .INP(n3739), .ZN(U8074_n1) );
  NOR2X0 U8074_U1 ( .IN1(g1018), .IN2(U8074_n1), .QN(n4193) );
  INVX0 U8088_U2 ( .INP(n3669), .ZN(U8088_n1) );
  NOR2X0 U8088_U1 ( .IN1(g1024), .IN2(U8088_n1), .QN(n3738) );
  INVX0 U8112_U2 ( .INP(n4525), .ZN(U8112_n1) );
  NOR2X0 U8112_U1 ( .IN1(n4523), .IN2(U8112_n1), .QN(n4524) );
  INVX0 U8113_U2 ( .INP(n4526), .ZN(U8113_n1) );
  NOR2X0 U8113_U1 ( .IN1(n5751), .IN2(U8113_n1), .QN(n4523) );
  INVX0 U8147_U2 ( .INP(g4659), .ZN(U8147_n1) );
  NOR2X0 U8147_U1 ( .IN1(n2573), .IN2(U8147_n1), .QN(n2577) );
  INVX0 U8165_U2 ( .INP(g4849), .ZN(U8165_n1) );
  NOR2X0 U8165_U1 ( .IN1(n2563), .IN2(U8165_n1), .QN(n2567) );
  INVX0 U8185_U2 ( .INP(n4940), .ZN(U8185_n1) );
  NOR2X0 U8185_U1 ( .IN1(g1046), .IN2(U8185_n1), .QN(n4938) );
  INVX0 U8192_U2 ( .INP(n4915), .ZN(U8192_n1) );
  NOR2X0 U8192_U1 ( .IN1(g1389), .IN2(U8192_n1), .QN(n4913) );
  INVX0 U8210_U2 ( .INP(n4722), .ZN(U8210_n1) );
  NOR2X0 U8210_U1 ( .IN1(n4723), .IN2(U8210_n1), .QN(n4714) );
  INVX0 U8223_U2 ( .INP(n42), .ZN(U8223_n1) );
  NOR2X0 U8223_U1 ( .IN1(n4516), .IN2(U8223_n1), .QN(n4517) );
  INVX0 U8224_U2 ( .INP(n4519), .ZN(U8224_n1) );
  NOR2X0 U8224_U1 ( .IN1(n5728), .IN2(U8224_n1), .QN(n4516) );
  INVX0 U8281_U2 ( .INP(n4819), .ZN(U8281_n1) );
  NOR2X0 U8281_U1 ( .IN1(n10465), .IN2(U8281_n1), .QN(n5111) );
  INVX0 U8307_U2 ( .INP(g29216), .ZN(U8307_n1) );
  NOR2X0 U8307_U1 ( .IN1(n10464), .IN2(U8307_n1), .QN(g26900) );
  INVX0 U8974_U2 ( .INP(n3362), .ZN(U8974_n1) );
  NOR2X0 U8974_U1 ( .IN1(test_so25), .IN2(U8974_n1), .QN(n2552) );
  INVX0 U8975_U2 ( .INP(n3174), .ZN(U8975_n1) );
  NOR2X0 U8975_U1 ( .IN1(g528), .IN2(U8975_n1), .QN(n3195) );
  INVX0 U9065_U2 ( .INP(g4145), .ZN(U9065_n1) );
  NOR2X0 U9065_U1 ( .IN1(n10465), .IN2(U9065_n1), .QN(n4721) );
  INVX0 U9070_U2 ( .INP(g2841), .ZN(U9070_n1) );
  NOR2X0 U9070_U1 ( .IN1(n10465), .IN2(U9070_n1), .QN(n3730) );
  INVX0 U9075_U2 ( .INP(g19), .ZN(U9075_n1) );
  NOR2X0 U9075_U1 ( .IN1(g9), .IN2(U9075_n1), .QN(n3362) );
  INVX0 U9076_U2 ( .INP(g113), .ZN(U9076_n1) );
  NOR2X0 U9076_U1 ( .IN1(n10464), .IN2(U9076_n1), .QN(g25694) );
  INVX0 U9080_U2 ( .INP(n4305), .ZN(U9080_n1) );
  NOR2X0 U9080_U1 ( .IN1(n10465), .IN2(U9080_n1), .QN(g29277) );
  INVX0 U9084_U2 ( .INP(g4423), .ZN(U9084_n1) );
  NOR2X0 U9084_U1 ( .IN1(n10464), .IN2(U9084_n1), .QN(g26953) );
  INVX0 U9085_U2 ( .INP(g64), .ZN(U9085_n1) );
  NOR2X0 U9085_U1 ( .IN1(n10464), .IN2(U9085_n1), .QN(g24212) );
  INVX0 U9086_U2 ( .INP(n4283), .ZN(U9086_n1) );
  NOR2X0 U9086_U1 ( .IN1(n10465), .IN2(U9086_n1), .QN(g29279) );
  INVX0 U9090_U2 ( .INP(g125), .ZN(U9090_n1) );
  NOR2X0 U9090_U1 ( .IN1(n10464), .IN2(U9090_n1), .QN(g25688) );
  INVX0 U9098_U2 ( .INP(g4681), .ZN(U9098_n1) );
  NOR2X0 U9098_U1 ( .IN1(n2774), .IN2(U9098_n1), .QN(g34028) );
  INVX0 U9099_U2 ( .INP(n2595), .ZN(U9099_n1) );
  NOR2X0 U9099_U1 ( .IN1(n2608), .IN2(U9099_n1), .QN(g34449) );
  INVX0 U9101_U2 ( .INP(g6745), .ZN(U9101_n1) );
  NOR2X0 U9101_U1 ( .IN1(n10464), .IN2(U9101_n1), .QN(g26880) );
  INVX0 U9107_U2 ( .INP(n4448), .ZN(U9107_n1) );
  NOR2X0 U9107_U1 ( .IN1(n10115), .IN2(U9107_n1), .QN(n4447) );
  INVX0 U9111_U2 ( .INP(n4403), .ZN(U9111_n1) );
  NOR2X0 U9111_U1 ( .IN1(n401), .IN2(U9111_n1), .QN(n4402) );
  INVX0 U9116_U2 ( .INP(n4426), .ZN(U9116_n1) );
  NOR2X0 U9116_U1 ( .IN1(n10120), .IN2(U9116_n1), .QN(n4425) );
  INVX0 U9120_U2 ( .INP(n4437), .ZN(U9120_n1) );
  NOR2X0 U9120_U1 ( .IN1(n10111), .IN2(U9120_n1), .QN(n4436) );
  INVX0 U9124_U2 ( .INP(n4392), .ZN(U9124_n1) );
  NOR2X0 U9124_U1 ( .IN1(n10117), .IN2(U9124_n1), .QN(n4391) );
  INVX0 U9128_U2 ( .INP(n4380), .ZN(U9128_n1) );
  NOR2X0 U9128_U1 ( .IN1(n10112), .IN2(U9128_n1), .QN(n4379) );
  INVX0 U9132_U2 ( .INP(n4415), .ZN(U9132_n1) );
  NOR2X0 U9132_U1 ( .IN1(n10119), .IN2(U9132_n1), .QN(n4414) );
  INVX0 U9136_U2 ( .INP(n4459), .ZN(U9136_n1) );
  NOR2X0 U9136_U1 ( .IN1(n1019), .IN2(U9136_n1), .QN(n4458) );
  INVX0 U9315_U2 ( .INP(n5016), .ZN(U9315_n1) );
  NOR2X0 U9315_U1 ( .IN1(n5753), .IN2(U9315_n1), .QN(n5014) );
  INVX0 U9453_U2 ( .INP(n3065), .ZN(U9453_n1) );
  NOR2X0 U9453_U1 ( .IN1(n10114), .IN2(U9453_n1), .QN(n3064) );
  INVX0 U9825_U2 ( .INP(g112), .ZN(U9825_n1) );
  NOR2X0 U9825_U1 ( .IN1(n1289), .IN2(U9825_n1), .QN(n3115) );
  INVX0 U9886_U2 ( .INP(g370), .ZN(U9886_n1) );
  NOR2X0 U9886_U1 ( .IN1(n5121), .IN2(U9886_n1), .QN(n4948) );
  INVX0 U9927_U2 ( .INP(n3933), .ZN(U9927_n1) );
  NOR2X0 U9927_U1 ( .IN1(g4098), .IN2(U9927_n1), .QN(n3833) );
  INVX0 U9953_U2 ( .INP(g671), .ZN(U9953_n1) );
  NOR2X0 U9953_U1 ( .IN1(n10107), .IN2(U9953_n1), .QN(n4526) );
  INVX0 U9957_U2 ( .INP(g4843), .ZN(U9957_n1) );
  NOR2X0 U9957_U1 ( .IN1(n5283), .IN2(U9957_n1), .QN(n2563) );
  INVX0 U9958_U2 ( .INP(test_so19), .ZN(U9958_n1) );
  NOR2X0 U9958_U1 ( .IN1(n5656), .IN2(U9958_n1), .QN(n2573) );
  INVX0 U9968_U2 ( .INP(n3084), .ZN(U9968_n1) );
  NOR2X0 U9968_U1 ( .IN1(g4358), .IN2(U9968_n1), .QN(n3023) );
  INVX0 U9972_U2 ( .INP(g681), .ZN(U9972_n1) );
  NOR2X0 U9972_U1 ( .IN1(n4535), .IN2(U9972_n1), .QN(n5112) );
  INVX0 U9992_U2 ( .INP(n3675), .ZN(U9992_n1) );
  NOR2X0 U9992_U1 ( .IN1(n3676), .IN2(U9992_n1), .QN(n2644) );
  INVX0 U10314_U2 ( .INP(g667), .ZN(U10314_n1) );
  NOR2X0 U10314_U1 ( .IN1(g686), .IN2(U10314_n1), .QN(n4962) );
  INVX0 U10318_U2 ( .INP(g5092), .ZN(U10318_n1) );
  NOR2X0 U10318_U1 ( .IN1(n5681), .IN2(U10318_n1), .QN(n5016) );
endmodule

