module add_mul_comp_16_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, 
        b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, 
        b_14_, b_15_, Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, 
        Result_5_, Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, 
        Result_11_, Result_12_, Result_13_, Result_14_, Result_15_, Result_16_, 
        Result_17_, Result_18_, Result_19_, Result_20_, Result_21_, Result_22_, 
        Result_23_, Result_24_, Result_25_, Result_26_, Result_27_, Result_28_, 
        Result_29_, Result_30_, Result_31_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_,
         b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_;
  wire   n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303;

  NOR2_X2 U2174 ( .A1(n4172), .A2(n2194), .ZN(n2450) );
  INV_X2 U2175 ( .A(n2195), .ZN(n2142) );
  NOR2_X1 U2176 ( .A1(n2142), .A2(n2143), .ZN(Result_9_) );
  XOR2_X1 U2177 ( .A(n2144), .B(n2145), .Z(n2143) );
  NOR2_X1 U2178 ( .A1(n2146), .A2(n2147), .ZN(n2145) );
  NAND2_X1 U2179 ( .A1(n2148), .A2(n2149), .ZN(n2144) );
  NAND2_X1 U2180 ( .A1(n2150), .A2(n2151), .ZN(n2148) );
  NAND2_X1 U2181 ( .A1(n2152), .A2(n2153), .ZN(n2151) );
  NOR2_X1 U2182 ( .A1(n2142), .A2(n2154), .ZN(Result_8_) );
  XNOR2_X1 U2183 ( .A(n2155), .B(n2156), .ZN(n2154) );
  NOR2_X1 U2184 ( .A1(n2142), .A2(n2157), .ZN(Result_7_) );
  XOR2_X1 U2185 ( .A(n2158), .B(n2159), .Z(n2157) );
  NOR2_X1 U2186 ( .A1(n2155), .A2(n2156), .ZN(n2159) );
  NAND2_X1 U2187 ( .A1(n2160), .A2(n2161), .ZN(n2158) );
  NAND2_X1 U2188 ( .A1(n2162), .A2(n2163), .ZN(n2160) );
  NAND2_X1 U2189 ( .A1(n2164), .A2(n2165), .ZN(n2163) );
  NOR2_X1 U2190 ( .A1(n2142), .A2(n2166), .ZN(Result_6_) );
  XNOR2_X1 U2191 ( .A(n2167), .B(n2168), .ZN(n2166) );
  NOR2_X1 U2192 ( .A1(n2142), .A2(n2169), .ZN(Result_5_) );
  XOR2_X1 U2193 ( .A(n2170), .B(n2171), .Z(n2169) );
  NOR2_X1 U2194 ( .A1(n2172), .A2(n2173), .ZN(n2171) );
  NOR2_X1 U2195 ( .A1(n2174), .A2(n2175), .ZN(n2173) );
  NOR2_X1 U2196 ( .A1(n2176), .A2(n2177), .ZN(n2174) );
  NAND2_X1 U2197 ( .A1(n2168), .A2(n2167), .ZN(n2170) );
  NOR2_X1 U2198 ( .A1(n2142), .A2(n2178), .ZN(Result_4_) );
  XNOR2_X1 U2199 ( .A(n2179), .B(n2180), .ZN(n2178) );
  NOR2_X1 U2200 ( .A1(n2142), .A2(n2181), .ZN(Result_3_) );
  XOR2_X1 U2201 ( .A(n2182), .B(n2183), .Z(n2181) );
  NOR2_X1 U2202 ( .A1(n2184), .A2(n2185), .ZN(n2183) );
  NOR2_X1 U2203 ( .A1(n2186), .A2(n2187), .ZN(n2185) );
  NOR2_X1 U2204 ( .A1(n2188), .A2(n2189), .ZN(n2186) );
  NAND2_X1 U2205 ( .A1(n2180), .A2(n2179), .ZN(n2182) );
  NAND2_X1 U2206 ( .A1(n2190), .A2(n2191), .ZN(Result_31_) );
  NAND3_X1 U2207 ( .A1(n2142), .A2(a_15_), .A3(n2192), .ZN(n2191) );
  NAND2_X1 U2208 ( .A1(n2193), .A2(b_15_), .ZN(n2190) );
  XOR2_X1 U2209 ( .A(n2194), .B(n2195), .Z(n2193) );
  NAND2_X1 U2210 ( .A1(n2196), .A2(n2197), .ZN(Result_30_) );
  NAND2_X1 U2211 ( .A1(n2198), .A2(n2195), .ZN(n2197) );
  NAND2_X1 U2212 ( .A1(n2199), .A2(n2200), .ZN(n2198) );
  NAND2_X1 U2213 ( .A1(b_14_), .A2(n2201), .ZN(n2200) );
  NAND2_X1 U2214 ( .A1(n2202), .A2(n2203), .ZN(n2201) );
  NAND2_X1 U2215 ( .A1(b_15_), .A2(n2204), .ZN(n2199) );
  NAND2_X1 U2216 ( .A1(n2205), .A2(n2206), .ZN(n2204) );
  NAND2_X1 U2217 ( .A1(a_14_), .A2(n2207), .ZN(n2206) );
  NAND2_X1 U2218 ( .A1(n2208), .A2(n2142), .ZN(n2196) );
  XOR2_X1 U2219 ( .A(n2209), .B(n2210), .Z(n2208) );
  XOR2_X1 U2220 ( .A(b_14_), .B(a_14_), .Z(n2210) );
  NOR2_X1 U2221 ( .A1(n2192), .A2(n2194), .ZN(n2209) );
  NOR2_X1 U2222 ( .A1(n2142), .A2(n2211), .ZN(Result_2_) );
  XNOR2_X1 U2223 ( .A(n2212), .B(n2213), .ZN(n2211) );
  NAND2_X1 U2224 ( .A1(n2214), .A2(n2215), .ZN(Result_29_) );
  NAND2_X1 U2225 ( .A1(n2142), .A2(n2216), .ZN(n2215) );
  NAND3_X1 U2226 ( .A1(n2217), .A2(n2218), .A3(n2219), .ZN(n2216) );
  NAND2_X1 U2227 ( .A1(n2220), .A2(n2221), .ZN(n2219) );
  NAND3_X1 U2228 ( .A1(n2222), .A2(n2223), .A3(b_13_), .ZN(n2218) );
  NAND2_X1 U2229 ( .A1(n2224), .A2(n2225), .ZN(n2217) );
  XOR2_X1 U2230 ( .A(n2223), .B(n2222), .Z(n2224) );
  INV_X1 U2231 ( .A(n2221), .ZN(n2222) );
  NAND2_X1 U2232 ( .A1(n2226), .A2(n2195), .ZN(n2214) );
  XOR2_X1 U2233 ( .A(n2227), .B(n2228), .Z(n2226) );
  XOR2_X1 U2234 ( .A(n2229), .B(n2230), .Z(n2228) );
  NAND2_X1 U2235 ( .A1(n2231), .A2(n2232), .ZN(Result_28_) );
  NAND2_X1 U2236 ( .A1(n2233), .A2(n2195), .ZN(n2232) );
  XNOR2_X1 U2237 ( .A(n2234), .B(n2235), .ZN(n2233) );
  XNOR2_X1 U2238 ( .A(n2236), .B(n2237), .ZN(n2235) );
  NOR2_X1 U2239 ( .A1(n2192), .A2(n2238), .ZN(n2237) );
  NAND2_X1 U2240 ( .A1(n2239), .A2(n2142), .ZN(n2231) );
  XNOR2_X1 U2241 ( .A(n2240), .B(n2241), .ZN(n2239) );
  NAND2_X1 U2242 ( .A1(n2242), .A2(n2243), .ZN(n2240) );
  NAND2_X1 U2243 ( .A1(n2244), .A2(n2245), .ZN(Result_27_) );
  NAND2_X1 U2244 ( .A1(n2142), .A2(n2246), .ZN(n2245) );
  NAND3_X1 U2245 ( .A1(n2247), .A2(n2248), .A3(n2249), .ZN(n2246) );
  NAND2_X1 U2246 ( .A1(n2250), .A2(n2251), .ZN(n2249) );
  INV_X1 U2247 ( .A(n2252), .ZN(n2250) );
  NAND3_X1 U2248 ( .A1(n2253), .A2(n2254), .A3(b_11_), .ZN(n2248) );
  INV_X1 U2249 ( .A(n2251), .ZN(n2253) );
  NAND2_X1 U2250 ( .A1(n2255), .A2(n2256), .ZN(n2247) );
  XOR2_X1 U2251 ( .A(n2251), .B(a_11_), .Z(n2255) );
  NAND2_X1 U2252 ( .A1(n2257), .A2(n2195), .ZN(n2244) );
  XNOR2_X1 U2253 ( .A(n2258), .B(n2259), .ZN(n2257) );
  XNOR2_X1 U2254 ( .A(n2260), .B(n2261), .ZN(n2258) );
  NAND2_X1 U2255 ( .A1(n2262), .A2(n2263), .ZN(Result_26_) );
  NAND2_X1 U2256 ( .A1(n2264), .A2(n2195), .ZN(n2263) );
  XNOR2_X1 U2257 ( .A(n2265), .B(n2266), .ZN(n2264) );
  XOR2_X1 U2258 ( .A(n2267), .B(n2268), .Z(n2266) );
  NAND2_X1 U2259 ( .A1(n2269), .A2(n2142), .ZN(n2262) );
  XNOR2_X1 U2260 ( .A(n2270), .B(n2271), .ZN(n2269) );
  NAND2_X1 U2261 ( .A1(n2272), .A2(n2273), .ZN(n2271) );
  NAND2_X1 U2262 ( .A1(n2274), .A2(n2275), .ZN(Result_25_) );
  NAND2_X1 U2263 ( .A1(n2142), .A2(n2276), .ZN(n2275) );
  NAND3_X1 U2264 ( .A1(n2277), .A2(n2278), .A3(n2279), .ZN(n2276) );
  NAND2_X1 U2265 ( .A1(n2280), .A2(n2281), .ZN(n2279) );
  NAND3_X1 U2266 ( .A1(n2282), .A2(n2283), .A3(b_9_), .ZN(n2278) );
  NAND2_X1 U2267 ( .A1(n2284), .A2(n2285), .ZN(n2277) );
  XOR2_X1 U2268 ( .A(n2281), .B(a_9_), .Z(n2284) );
  NAND2_X1 U2269 ( .A1(n2286), .A2(n2195), .ZN(n2274) );
  XNOR2_X1 U2270 ( .A(n2287), .B(n2288), .ZN(n2286) );
  XNOR2_X1 U2271 ( .A(n2289), .B(n2290), .ZN(n2287) );
  NAND2_X1 U2272 ( .A1(n2291), .A2(n2292), .ZN(Result_24_) );
  NAND2_X1 U2273 ( .A1(n2293), .A2(n2195), .ZN(n2292) );
  XOR2_X1 U2274 ( .A(n2294), .B(n2295), .Z(n2293) );
  XNOR2_X1 U2275 ( .A(n2296), .B(n2297), .ZN(n2294) );
  NAND2_X1 U2276 ( .A1(n2298), .A2(n2142), .ZN(n2291) );
  XNOR2_X1 U2277 ( .A(n2299), .B(n2300), .ZN(n2298) );
  NOR2_X1 U2278 ( .A1(n2301), .A2(n2302), .ZN(n2300) );
  NAND2_X1 U2279 ( .A1(n2303), .A2(n2304), .ZN(Result_23_) );
  NAND2_X1 U2280 ( .A1(n2142), .A2(n2305), .ZN(n2304) );
  NAND3_X1 U2281 ( .A1(n2306), .A2(n2307), .A3(n2308), .ZN(n2305) );
  NAND2_X1 U2282 ( .A1(n2309), .A2(n2310), .ZN(n2308) );
  NAND3_X1 U2283 ( .A1(n2311), .A2(n2312), .A3(b_7_), .ZN(n2307) );
  NAND2_X1 U2284 ( .A1(n2313), .A2(n2314), .ZN(n2306) );
  XOR2_X1 U2285 ( .A(n2310), .B(a_7_), .Z(n2313) );
  NAND2_X1 U2286 ( .A1(n2315), .A2(n2195), .ZN(n2303) );
  XNOR2_X1 U2287 ( .A(n2316), .B(n2317), .ZN(n2315) );
  NAND2_X1 U2288 ( .A1(n2318), .A2(n2319), .ZN(n2316) );
  NAND2_X1 U2289 ( .A1(n2320), .A2(n2321), .ZN(Result_22_) );
  NAND2_X1 U2290 ( .A1(n2322), .A2(n2195), .ZN(n2321) );
  XNOR2_X1 U2291 ( .A(n2323), .B(n2324), .ZN(n2322) );
  XOR2_X1 U2292 ( .A(n2325), .B(n2326), .Z(n2324) );
  NAND2_X1 U2293 ( .A1(n2327), .A2(n2142), .ZN(n2320) );
  XNOR2_X1 U2294 ( .A(n2328), .B(n2329), .ZN(n2327) );
  NAND2_X1 U2295 ( .A1(n2330), .A2(n2331), .ZN(n2329) );
  NAND2_X1 U2296 ( .A1(n2332), .A2(n2333), .ZN(Result_21_) );
  NAND2_X1 U2297 ( .A1(n2142), .A2(n2334), .ZN(n2333) );
  NAND3_X1 U2298 ( .A1(n2335), .A2(n2336), .A3(n2337), .ZN(n2334) );
  NAND2_X1 U2299 ( .A1(n2338), .A2(n2339), .ZN(n2337) );
  NAND3_X1 U2300 ( .A1(n2340), .A2(n2341), .A3(b_5_), .ZN(n2336) );
  NAND2_X1 U2301 ( .A1(n2342), .A2(n2343), .ZN(n2335) );
  XOR2_X1 U2302 ( .A(n2340), .B(n2341), .Z(n2342) );
  INV_X1 U2303 ( .A(n2339), .ZN(n2340) );
  NAND2_X1 U2304 ( .A1(n2344), .A2(n2195), .ZN(n2332) );
  XNOR2_X1 U2305 ( .A(n2345), .B(n2346), .ZN(n2344) );
  NAND2_X1 U2306 ( .A1(n2347), .A2(n2348), .ZN(n2345) );
  NAND2_X1 U2307 ( .A1(n2349), .A2(n2350), .ZN(Result_20_) );
  NAND2_X1 U2308 ( .A1(n2351), .A2(n2195), .ZN(n2350) );
  XOR2_X1 U2309 ( .A(n2352), .B(n2353), .Z(n2351) );
  XOR2_X1 U2310 ( .A(n2354), .B(n2355), .Z(n2353) );
  NAND2_X1 U2311 ( .A1(n2356), .A2(n2142), .ZN(n2349) );
  XNOR2_X1 U2312 ( .A(n2357), .B(n2358), .ZN(n2356) );
  NAND2_X1 U2313 ( .A1(n2359), .A2(n2360), .ZN(n2358) );
  NOR2_X1 U2314 ( .A1(n2142), .A2(n2361), .ZN(Result_1_) );
  XOR2_X1 U2315 ( .A(n2362), .B(n2363), .Z(n2361) );
  NOR2_X1 U2316 ( .A1(n2364), .A2(n2365), .ZN(n2363) );
  NAND2_X1 U2317 ( .A1(n2366), .A2(n2367), .ZN(Result_19_) );
  NAND2_X1 U2318 ( .A1(n2142), .A2(n2368), .ZN(n2367) );
  NAND3_X1 U2319 ( .A1(n2369), .A2(n2370), .A3(n2371), .ZN(n2368) );
  NAND2_X1 U2320 ( .A1(n2372), .A2(n2373), .ZN(n2371) );
  INV_X1 U2321 ( .A(n2374), .ZN(n2372) );
  NAND3_X1 U2322 ( .A1(n2375), .A2(n2376), .A3(b_3_), .ZN(n2370) );
  INV_X1 U2323 ( .A(n2373), .ZN(n2375) );
  NAND2_X1 U2324 ( .A1(n2377), .A2(n2378), .ZN(n2369) );
  XOR2_X1 U2325 ( .A(n2373), .B(a_3_), .Z(n2377) );
  NAND2_X1 U2326 ( .A1(n2379), .A2(n2195), .ZN(n2366) );
  XOR2_X1 U2327 ( .A(n2380), .B(n2381), .Z(n2379) );
  XOR2_X1 U2328 ( .A(n2382), .B(n2383), .Z(n2380) );
  NAND2_X1 U2329 ( .A1(n2384), .A2(n2385), .ZN(Result_18_) );
  NAND2_X1 U2330 ( .A1(n2386), .A2(n2195), .ZN(n2385) );
  XNOR2_X1 U2331 ( .A(n2387), .B(n2388), .ZN(n2386) );
  XOR2_X1 U2332 ( .A(n2389), .B(n2390), .Z(n2388) );
  NAND2_X1 U2333 ( .A1(a_2_), .A2(b_15_), .ZN(n2390) );
  NAND2_X1 U2334 ( .A1(n2391), .A2(n2142), .ZN(n2384) );
  XNOR2_X1 U2335 ( .A(n2392), .B(n2393), .ZN(n2391) );
  NAND2_X1 U2336 ( .A1(n2394), .A2(n2395), .ZN(n2393) );
  NAND2_X1 U2337 ( .A1(n2396), .A2(n2397), .ZN(Result_17_) );
  NAND2_X1 U2338 ( .A1(n2398), .A2(n2195), .ZN(n2397) );
  XOR2_X1 U2339 ( .A(n2399), .B(n2400), .Z(n2398) );
  XNOR2_X1 U2340 ( .A(n2401), .B(n2402), .ZN(n2400) );
  NAND2_X1 U2341 ( .A1(b_15_), .A2(a_1_), .ZN(n2402) );
  NAND2_X1 U2342 ( .A1(n2403), .A2(n2142), .ZN(n2396) );
  NAND2_X1 U2343 ( .A1(n2404), .A2(n2405), .ZN(n2403) );
  NAND2_X1 U2344 ( .A1(n2406), .A2(n2407), .ZN(n2405) );
  INV_X1 U2345 ( .A(n2408), .ZN(n2406) );
  NOR2_X1 U2346 ( .A1(n2409), .A2(n2410), .ZN(n2408) );
  NAND2_X1 U2347 ( .A1(n2411), .A2(n2412), .ZN(n2404) );
  INV_X1 U2348 ( .A(n2407), .ZN(n2412) );
  XOR2_X1 U2349 ( .A(b_1_), .B(a_1_), .Z(n2411) );
  NAND2_X1 U2350 ( .A1(n2413), .A2(n2414), .ZN(Result_16_) );
  NAND2_X1 U2351 ( .A1(n2415), .A2(n2195), .ZN(n2414) );
  XOR2_X1 U2352 ( .A(n2416), .B(n2417), .Z(n2415) );
  XOR2_X1 U2353 ( .A(n2418), .B(n2419), .Z(n2416) );
  NOR2_X1 U2354 ( .A1(n2192), .A2(n2420), .ZN(n2419) );
  NAND2_X1 U2355 ( .A1(n2421), .A2(n2142), .ZN(n2413) );
  XNOR2_X1 U2356 ( .A(n2422), .B(n2423), .ZN(n2421) );
  NOR2_X1 U2357 ( .A1(n2410), .A2(n2424), .ZN(n2422) );
  NOR2_X1 U2358 ( .A1(n2409), .A2(n2407), .ZN(n2424) );
  NAND2_X1 U2359 ( .A1(n2395), .A2(n2425), .ZN(n2407) );
  NAND2_X1 U2360 ( .A1(n2394), .A2(n2392), .ZN(n2425) );
  NAND2_X1 U2361 ( .A1(n2374), .A2(n2426), .ZN(n2392) );
  NAND2_X1 U2362 ( .A1(n2427), .A2(n2373), .ZN(n2426) );
  NAND2_X1 U2363 ( .A1(n2360), .A2(n2428), .ZN(n2373) );
  NAND2_X1 U2364 ( .A1(n2359), .A2(n2357), .ZN(n2428) );
  NAND2_X1 U2365 ( .A1(n2429), .A2(n2430), .ZN(n2357) );
  NAND2_X1 U2366 ( .A1(n2431), .A2(n2339), .ZN(n2430) );
  NAND2_X1 U2367 ( .A1(n2331), .A2(n2432), .ZN(n2339) );
  NAND2_X1 U2368 ( .A1(n2330), .A2(n2328), .ZN(n2432) );
  NAND2_X1 U2369 ( .A1(n2433), .A2(n2434), .ZN(n2328) );
  NAND2_X1 U2370 ( .A1(n2435), .A2(n2310), .ZN(n2434) );
  INV_X1 U2371 ( .A(n2311), .ZN(n2310) );
  NOR2_X1 U2372 ( .A1(n2302), .A2(n2436), .ZN(n2311) );
  NOR2_X1 U2373 ( .A1(n2301), .A2(n2299), .ZN(n2436) );
  NOR2_X1 U2374 ( .A1(n2280), .A2(n2437), .ZN(n2299) );
  NOR2_X1 U2375 ( .A1(n2438), .A2(n2282), .ZN(n2437) );
  INV_X1 U2376 ( .A(n2281), .ZN(n2282) );
  NAND2_X1 U2377 ( .A1(n2273), .A2(n2439), .ZN(n2281) );
  NAND2_X1 U2378 ( .A1(n2272), .A2(n2270), .ZN(n2439) );
  NAND2_X1 U2379 ( .A1(n2252), .A2(n2440), .ZN(n2270) );
  NAND2_X1 U2380 ( .A1(n2441), .A2(n2251), .ZN(n2440) );
  NAND2_X1 U2381 ( .A1(n2242), .A2(n2442), .ZN(n2251) );
  NAND2_X1 U2382 ( .A1(n2243), .A2(n2241), .ZN(n2442) );
  NAND2_X1 U2383 ( .A1(n2443), .A2(n2444), .ZN(n2241) );
  NAND2_X1 U2384 ( .A1(n2445), .A2(n2221), .ZN(n2444) );
  NAND3_X1 U2385 ( .A1(n2446), .A2(n2447), .A3(n2448), .ZN(n2221) );
  NAND2_X1 U2386 ( .A1(a_14_), .A2(b_14_), .ZN(n2448) );
  NAND2_X1 U2387 ( .A1(n2449), .A2(a_15_), .ZN(n2447) );
  NAND2_X1 U2388 ( .A1(n2450), .A2(b_15_), .ZN(n2446) );
  NAND2_X1 U2389 ( .A1(n2225), .A2(n2223), .ZN(n2445) );
  NAND2_X1 U2390 ( .A1(n2451), .A2(n2238), .ZN(n2243) );
  NAND2_X1 U2391 ( .A1(n2256), .A2(n2254), .ZN(n2441) );
  NAND2_X1 U2392 ( .A1(n2452), .A2(n2453), .ZN(n2272) );
  NOR2_X1 U2393 ( .A1(b_9_), .A2(a_9_), .ZN(n2438) );
  NOR2_X1 U2394 ( .A1(b_8_), .A2(a_8_), .ZN(n2301) );
  NAND2_X1 U2395 ( .A1(n2314), .A2(n2312), .ZN(n2435) );
  NAND2_X1 U2396 ( .A1(n2454), .A2(n2455), .ZN(n2330) );
  NAND2_X1 U2397 ( .A1(n2343), .A2(n2341), .ZN(n2431) );
  NAND2_X1 U2398 ( .A1(n2456), .A2(n2457), .ZN(n2359) );
  INV_X1 U2399 ( .A(n2458), .ZN(n2360) );
  NAND2_X1 U2400 ( .A1(n2378), .A2(n2376), .ZN(n2427) );
  NAND2_X1 U2401 ( .A1(n2459), .A2(n2460), .ZN(n2394) );
  NOR2_X1 U2402 ( .A1(b_1_), .A2(a_1_), .ZN(n2410) );
  NOR2_X1 U2403 ( .A1(n2142), .A2(n2461), .ZN(Result_15_) );
  XNOR2_X1 U2404 ( .A(n2462), .B(n2463), .ZN(n2461) );
  NOR3_X1 U2405 ( .A1(n2464), .A2(n2142), .A3(n2465), .ZN(Result_14_) );
  NOR2_X1 U2406 ( .A1(n2466), .A2(n2467), .ZN(n2464) );
  XOR2_X1 U2407 ( .A(n2468), .B(n2469), .Z(n2467) );
  NOR2_X1 U2408 ( .A1(n2462), .A2(n2463), .ZN(n2466) );
  NOR2_X1 U2409 ( .A1(n2142), .A2(n2470), .ZN(Result_13_) );
  XNOR2_X1 U2410 ( .A(n2465), .B(n2471), .ZN(n2470) );
  NOR2_X1 U2411 ( .A1(n2472), .A2(n2473), .ZN(n2471) );
  INV_X1 U2412 ( .A(n2474), .ZN(n2473) );
  NAND2_X1 U2413 ( .A1(n2475), .A2(n2476), .ZN(n2474) );
  NOR2_X1 U2414 ( .A1(n2142), .A2(n2477), .ZN(Result_12_) );
  XNOR2_X1 U2415 ( .A(n2478), .B(n2479), .ZN(n2477) );
  NOR2_X1 U2416 ( .A1(n2142), .A2(n2480), .ZN(Result_11_) );
  XOR2_X1 U2417 ( .A(n2481), .B(n2482), .Z(n2480) );
  NOR2_X1 U2418 ( .A1(n2479), .A2(n2478), .ZN(n2482) );
  NAND2_X1 U2419 ( .A1(n2483), .A2(n2484), .ZN(n2481) );
  NAND2_X1 U2420 ( .A1(n2485), .A2(n2486), .ZN(n2483) );
  NAND2_X1 U2421 ( .A1(n2487), .A2(n2488), .ZN(n2486) );
  NOR2_X1 U2422 ( .A1(n2142), .A2(n2489), .ZN(Result_10_) );
  XNOR2_X1 U2423 ( .A(n2147), .B(n2146), .ZN(n2489) );
  NOR2_X1 U2424 ( .A1(n2142), .A2(n2490), .ZN(Result_0_) );
  NOR3_X1 U2425 ( .A1(n2491), .A2(n2492), .A3(n2364), .ZN(n2490) );
  INV_X1 U2426 ( .A(n2493), .ZN(n2364) );
  NAND4_X1 U2427 ( .A1(b_0_), .A2(n2494), .A3(n2495), .A4(n2496), .ZN(n2493)
         );
  INV_X1 U2428 ( .A(n2494), .ZN(n2492) );
  NOR2_X1 U2429 ( .A1(n2365), .A2(n2362), .ZN(n2491) );
  NAND2_X1 U2430 ( .A1(n2213), .A2(n2212), .ZN(n2362) );
  NAND3_X1 U2431 ( .A1(n2497), .A2(n2498), .A3(n2499), .ZN(n2212) );
  NAND3_X1 U2432 ( .A1(n2180), .A2(n2179), .A3(n2187), .ZN(n2499) );
  INV_X1 U2433 ( .A(n2500), .ZN(n2187) );
  NAND3_X1 U2434 ( .A1(n2501), .A2(n2502), .A3(n2503), .ZN(n2179) );
  NAND3_X1 U2435 ( .A1(n2168), .A2(n2167), .A3(n2175), .ZN(n2503) );
  INV_X1 U2436 ( .A(n2504), .ZN(n2175) );
  NAND3_X1 U2437 ( .A1(n2505), .A2(n2161), .A3(n2506), .ZN(n2167) );
  INV_X1 U2438 ( .A(n2507), .ZN(n2506) );
  NOR3_X1 U2439 ( .A1(n2156), .A2(n2155), .A3(n2162), .ZN(n2507) );
  NOR3_X1 U2440 ( .A1(n2508), .A2(n2509), .A3(n2510), .ZN(n2155) );
  NOR3_X1 U2441 ( .A1(n2150), .A2(n2146), .A3(n2147), .ZN(n2510) );
  XNOR2_X1 U2442 ( .A(n2152), .B(n2153), .ZN(n2147) );
  NOR3_X1 U2443 ( .A1(n2511), .A2(n2512), .A3(n2513), .ZN(n2146) );
  NOR3_X1 U2444 ( .A1(n2485), .A2(n2479), .A3(n2478), .ZN(n2513) );
  XNOR2_X1 U2445 ( .A(n2487), .B(n2488), .ZN(n2478) );
  NOR3_X1 U2446 ( .A1(n2514), .A2(n2472), .A3(n2515), .ZN(n2479) );
  NOR2_X1 U2447 ( .A1(n2516), .A2(n2476), .ZN(n2515) );
  INV_X1 U2448 ( .A(n2465), .ZN(n2516) );
  NOR4_X1 U2449 ( .A1(n2463), .A2(n2517), .A3(n2462), .A4(n2518), .ZN(n2465)
         );
  INV_X1 U2450 ( .A(n2475), .ZN(n2518) );
  NOR2_X1 U2451 ( .A1(n2519), .A2(n2520), .ZN(n2462) );
  NOR3_X1 U2452 ( .A1(n2192), .A2(n2521), .A3(n2420), .ZN(n2520) );
  NOR2_X1 U2453 ( .A1(n2418), .A2(n2417), .ZN(n2521) );
  INV_X1 U2454 ( .A(n2522), .ZN(n2519) );
  NAND2_X1 U2455 ( .A1(n2417), .A2(n2418), .ZN(n2522) );
  NAND2_X1 U2456 ( .A1(n2523), .A2(n2524), .ZN(n2418) );
  NAND3_X1 U2457 ( .A1(a_1_), .A2(n2525), .A3(b_15_), .ZN(n2524) );
  NAND2_X1 U2458 ( .A1(n2401), .A2(n2399), .ZN(n2525) );
  INV_X1 U2459 ( .A(n2526), .ZN(n2523) );
  NOR2_X1 U2460 ( .A1(n2399), .A2(n2401), .ZN(n2526) );
  NOR2_X1 U2461 ( .A1(n2527), .A2(n2528), .ZN(n2401) );
  NOR3_X1 U2462 ( .A1(n2192), .A2(n2529), .A3(n2460), .ZN(n2528) );
  NOR2_X1 U2463 ( .A1(n2389), .A2(n2387), .ZN(n2529) );
  INV_X1 U2464 ( .A(n2530), .ZN(n2527) );
  NAND2_X1 U2465 ( .A1(n2387), .A2(n2389), .ZN(n2530) );
  NAND2_X1 U2466 ( .A1(n2531), .A2(n2532), .ZN(n2389) );
  NAND2_X1 U2467 ( .A1(n2383), .A2(n2533), .ZN(n2532) );
  INV_X1 U2468 ( .A(n2534), .ZN(n2533) );
  NOR2_X1 U2469 ( .A1(n2382), .A2(n2381), .ZN(n2534) );
  NOR2_X1 U2470 ( .A1(n2376), .A2(n2192), .ZN(n2383) );
  NAND2_X1 U2471 ( .A1(n2381), .A2(n2382), .ZN(n2531) );
  NAND2_X1 U2472 ( .A1(n2535), .A2(n2536), .ZN(n2382) );
  NAND2_X1 U2473 ( .A1(n2355), .A2(n2537), .ZN(n2536) );
  INV_X1 U2474 ( .A(n2538), .ZN(n2537) );
  NOR2_X1 U2475 ( .A1(n2354), .A2(n2352), .ZN(n2538) );
  NOR2_X1 U2476 ( .A1(n2457), .A2(n2192), .ZN(n2355) );
  NAND2_X1 U2477 ( .A1(n2352), .A2(n2354), .ZN(n2535) );
  NAND2_X1 U2478 ( .A1(n2347), .A2(n2539), .ZN(n2354) );
  NAND2_X1 U2479 ( .A1(n2346), .A2(n2348), .ZN(n2539) );
  NAND2_X1 U2480 ( .A1(n2540), .A2(n2541), .ZN(n2348) );
  INV_X1 U2481 ( .A(n2542), .ZN(n2541) );
  NAND2_X1 U2482 ( .A1(a_5_), .A2(b_15_), .ZN(n2540) );
  XNOR2_X1 U2483 ( .A(n2543), .B(n2544), .ZN(n2346) );
  XNOR2_X1 U2484 ( .A(n2545), .B(n2546), .ZN(n2543) );
  NOR2_X1 U2485 ( .A1(n2207), .A2(n2455), .ZN(n2546) );
  NAND2_X1 U2486 ( .A1(n2542), .A2(a_5_), .ZN(n2347) );
  NOR2_X1 U2487 ( .A1(n2547), .A2(n2548), .ZN(n2542) );
  INV_X1 U2488 ( .A(n2549), .ZN(n2548) );
  NAND2_X1 U2489 ( .A1(n2550), .A2(n2325), .ZN(n2549) );
  NAND2_X1 U2490 ( .A1(a_6_), .A2(b_15_), .ZN(n2325) );
  NAND2_X1 U2491 ( .A1(n2323), .A2(n2326), .ZN(n2550) );
  NOR2_X1 U2492 ( .A1(n2326), .A2(n2323), .ZN(n2547) );
  XOR2_X1 U2493 ( .A(n2551), .B(n2552), .Z(n2323) );
  XNOR2_X1 U2494 ( .A(n2553), .B(n2554), .ZN(n2552) );
  NAND2_X1 U2495 ( .A1(a_7_), .A2(b_14_), .ZN(n2554) );
  NAND2_X1 U2496 ( .A1(n2318), .A2(n2555), .ZN(n2326) );
  NAND2_X1 U2497 ( .A1(n2317), .A2(n2319), .ZN(n2555) );
  NAND2_X1 U2498 ( .A1(n2556), .A2(n2557), .ZN(n2319) );
  INV_X1 U2499 ( .A(n2558), .ZN(n2557) );
  NAND2_X1 U2500 ( .A1(a_7_), .A2(b_15_), .ZN(n2556) );
  XNOR2_X1 U2501 ( .A(n2559), .B(n2560), .ZN(n2317) );
  XOR2_X1 U2502 ( .A(n2561), .B(n2562), .Z(n2560) );
  NAND2_X1 U2503 ( .A1(a_8_), .A2(b_14_), .ZN(n2562) );
  NAND2_X1 U2504 ( .A1(n2558), .A2(a_7_), .ZN(n2318) );
  NOR2_X1 U2505 ( .A1(n2563), .A2(n2564), .ZN(n2558) );
  INV_X1 U2506 ( .A(n2565), .ZN(n2564) );
  NAND2_X1 U2507 ( .A1(n2566), .A2(n2297), .ZN(n2565) );
  NAND2_X1 U2508 ( .A1(a_8_), .A2(b_15_), .ZN(n2297) );
  NAND2_X1 U2509 ( .A1(n2295), .A2(n2296), .ZN(n2566) );
  NOR2_X1 U2510 ( .A1(n2296), .A2(n2295), .ZN(n2563) );
  XNOR2_X1 U2511 ( .A(n2567), .B(n2568), .ZN(n2295) );
  NAND2_X1 U2512 ( .A1(n2569), .A2(n2570), .ZN(n2567) );
  NAND2_X1 U2513 ( .A1(n2571), .A2(n2572), .ZN(n2296) );
  NAND2_X1 U2514 ( .A1(n2290), .A2(n2573), .ZN(n2572) );
  NAND2_X1 U2515 ( .A1(n2289), .A2(n2288), .ZN(n2573) );
  NOR2_X1 U2516 ( .A1(n2283), .A2(n2192), .ZN(n2290) );
  INV_X1 U2517 ( .A(n2574), .ZN(n2571) );
  NOR2_X1 U2518 ( .A1(n2288), .A2(n2289), .ZN(n2574) );
  NOR2_X1 U2519 ( .A1(n2575), .A2(n2576), .ZN(n2289) );
  NOR2_X1 U2520 ( .A1(n2267), .A2(n2577), .ZN(n2576) );
  NOR2_X1 U2521 ( .A1(n2268), .A2(n2265), .ZN(n2577) );
  NAND2_X1 U2522 ( .A1(a_10_), .A2(b_15_), .ZN(n2267) );
  INV_X1 U2523 ( .A(n2578), .ZN(n2575) );
  NAND2_X1 U2524 ( .A1(n2265), .A2(n2268), .ZN(n2578) );
  NAND2_X1 U2525 ( .A1(n2579), .A2(n2580), .ZN(n2268) );
  NAND2_X1 U2526 ( .A1(n2261), .A2(n2581), .ZN(n2580) );
  NAND2_X1 U2527 ( .A1(n2260), .A2(n2259), .ZN(n2581) );
  NOR2_X1 U2528 ( .A1(n2254), .A2(n2192), .ZN(n2261) );
  INV_X1 U2529 ( .A(n2582), .ZN(n2579) );
  NOR2_X1 U2530 ( .A1(n2259), .A2(n2260), .ZN(n2582) );
  NOR2_X1 U2531 ( .A1(n2583), .A2(n2584), .ZN(n2260) );
  NOR3_X1 U2532 ( .A1(n2192), .A2(n2585), .A3(n2238), .ZN(n2584) );
  NOR2_X1 U2533 ( .A1(n2236), .A2(n2234), .ZN(n2585) );
  INV_X1 U2534 ( .A(n2586), .ZN(n2583) );
  NAND2_X1 U2535 ( .A1(n2234), .A2(n2236), .ZN(n2586) );
  NAND2_X1 U2536 ( .A1(n2587), .A2(n2588), .ZN(n2236) );
  NAND2_X1 U2537 ( .A1(n2229), .A2(n2589), .ZN(n2588) );
  INV_X1 U2538 ( .A(n2590), .ZN(n2589) );
  NOR2_X1 U2539 ( .A1(n2227), .A2(n2230), .ZN(n2590) );
  NOR2_X1 U2540 ( .A1(n2223), .A2(n2192), .ZN(n2229) );
  NAND2_X1 U2541 ( .A1(n2230), .A2(n2227), .ZN(n2587) );
  NAND2_X1 U2542 ( .A1(n2591), .A2(n2592), .ZN(n2227) );
  NAND2_X1 U2543 ( .A1(b_13_), .A2(n2593), .ZN(n2592) );
  NAND2_X1 U2544 ( .A1(n2202), .A2(n2594), .ZN(n2593) );
  NAND2_X1 U2545 ( .A1(a_15_), .A2(n2207), .ZN(n2594) );
  NAND2_X1 U2546 ( .A1(b_14_), .A2(n2595), .ZN(n2591) );
  NAND2_X1 U2547 ( .A1(n2205), .A2(n2596), .ZN(n2595) );
  NAND2_X1 U2548 ( .A1(a_14_), .A2(n2225), .ZN(n2596) );
  NOR2_X1 U2549 ( .A1(n2597), .A2(n2598), .ZN(n2230) );
  XOR2_X1 U2550 ( .A(n2599), .B(n2600), .Z(n2234) );
  XOR2_X1 U2551 ( .A(n2601), .B(n2602), .Z(n2599) );
  XOR2_X1 U2552 ( .A(n2603), .B(n2604), .Z(n2259) );
  XNOR2_X1 U2553 ( .A(n2605), .B(n2606), .ZN(n2603) );
  XNOR2_X1 U2554 ( .A(n2607), .B(n2608), .ZN(n2265) );
  XOR2_X1 U2555 ( .A(n2609), .B(n2610), .Z(n2607) );
  NAND2_X1 U2556 ( .A1(a_11_), .A2(b_14_), .ZN(n2609) );
  XNOR2_X1 U2557 ( .A(n2611), .B(n2612), .ZN(n2288) );
  XNOR2_X1 U2558 ( .A(n2613), .B(n2614), .ZN(n2612) );
  XNOR2_X1 U2559 ( .A(n2615), .B(n2616), .ZN(n2352) );
  NAND2_X1 U2560 ( .A1(n2617), .A2(n2618), .ZN(n2615) );
  XOR2_X1 U2561 ( .A(n2619), .B(n2620), .Z(n2381) );
  XOR2_X1 U2562 ( .A(n2621), .B(n2622), .Z(n2619) );
  NOR2_X1 U2563 ( .A1(n2207), .A2(n2457), .ZN(n2622) );
  XNOR2_X1 U2564 ( .A(n2623), .B(n2624), .ZN(n2387) );
  XNOR2_X1 U2565 ( .A(n2625), .B(n2626), .ZN(n2623) );
  NOR2_X1 U2566 ( .A1(n2207), .A2(n2376), .ZN(n2626) );
  XNOR2_X1 U2567 ( .A(n2627), .B(n2628), .ZN(n2399) );
  XNOR2_X1 U2568 ( .A(n2629), .B(n2630), .ZN(n2628) );
  NAND2_X1 U2569 ( .A1(a_2_), .A2(b_14_), .ZN(n2630) );
  XOR2_X1 U2570 ( .A(n2631), .B(n2632), .Z(n2417) );
  XNOR2_X1 U2571 ( .A(n2633), .B(n2634), .ZN(n2632) );
  NAND2_X1 U2572 ( .A1(b_14_), .A2(a_1_), .ZN(n2634) );
  NOR2_X1 U2573 ( .A1(n2468), .A2(n2469), .ZN(n2517) );
  XOR2_X1 U2574 ( .A(n2635), .B(n2636), .Z(n2463) );
  XNOR2_X1 U2575 ( .A(n2637), .B(n2638), .ZN(n2635) );
  NOR2_X1 U2576 ( .A1(n2207), .A2(n2420), .ZN(n2638) );
  NOR2_X1 U2577 ( .A1(n2475), .A2(n2476), .ZN(n2472) );
  XNOR2_X1 U2578 ( .A(n2639), .B(n2640), .ZN(n2476) );
  NAND2_X1 U2579 ( .A1(n2469), .A2(n2468), .ZN(n2475) );
  NAND2_X1 U2580 ( .A1(n2641), .A2(n2642), .ZN(n2468) );
  NAND3_X1 U2581 ( .A1(b_14_), .A2(n2643), .A3(a_0_), .ZN(n2642) );
  NAND2_X1 U2582 ( .A1(n2637), .A2(n2636), .ZN(n2643) );
  INV_X1 U2583 ( .A(n2644), .ZN(n2641) );
  NOR2_X1 U2584 ( .A1(n2636), .A2(n2637), .ZN(n2644) );
  NOR2_X1 U2585 ( .A1(n2645), .A2(n2646), .ZN(n2637) );
  NOR3_X1 U2586 ( .A1(n2647), .A2(n2648), .A3(n2207), .ZN(n2646) );
  INV_X1 U2587 ( .A(n2649), .ZN(n2648) );
  NAND2_X1 U2588 ( .A1(n2633), .A2(n2631), .ZN(n2649) );
  NOR2_X1 U2589 ( .A1(n2631), .A2(n2633), .ZN(n2645) );
  NOR2_X1 U2590 ( .A1(n2650), .A2(n2651), .ZN(n2633) );
  INV_X1 U2591 ( .A(n2652), .ZN(n2651) );
  NAND3_X1 U2592 ( .A1(b_14_), .A2(n2653), .A3(a_2_), .ZN(n2652) );
  NAND2_X1 U2593 ( .A1(n2629), .A2(n2627), .ZN(n2653) );
  NOR2_X1 U2594 ( .A1(n2627), .A2(n2629), .ZN(n2650) );
  NOR2_X1 U2595 ( .A1(n2654), .A2(n2655), .ZN(n2629) );
  NOR3_X1 U2596 ( .A1(n2207), .A2(n2656), .A3(n2376), .ZN(n2655) );
  INV_X1 U2597 ( .A(n2657), .ZN(n2656) );
  NAND2_X1 U2598 ( .A1(n2625), .A2(n2624), .ZN(n2657) );
  NOR2_X1 U2599 ( .A1(n2624), .A2(n2625), .ZN(n2654) );
  NOR2_X1 U2600 ( .A1(n2658), .A2(n2659), .ZN(n2625) );
  NOR3_X1 U2601 ( .A1(n2207), .A2(n2660), .A3(n2457), .ZN(n2659) );
  NOR2_X1 U2602 ( .A1(n2621), .A2(n2620), .ZN(n2660) );
  INV_X1 U2603 ( .A(n2661), .ZN(n2658) );
  NAND2_X1 U2604 ( .A1(n2620), .A2(n2621), .ZN(n2661) );
  NAND2_X1 U2605 ( .A1(n2617), .A2(n2662), .ZN(n2621) );
  NAND2_X1 U2606 ( .A1(n2616), .A2(n2618), .ZN(n2662) );
  NAND2_X1 U2607 ( .A1(n2663), .A2(n2664), .ZN(n2618) );
  NAND2_X1 U2608 ( .A1(a_5_), .A2(b_14_), .ZN(n2664) );
  XNOR2_X1 U2609 ( .A(n2665), .B(n2666), .ZN(n2616) );
  XOR2_X1 U2610 ( .A(n2667), .B(n2668), .Z(n2666) );
  NAND2_X1 U2611 ( .A1(a_6_), .A2(b_13_), .ZN(n2668) );
  INV_X1 U2612 ( .A(n2669), .ZN(n2617) );
  NOR2_X1 U2613 ( .A1(n2341), .A2(n2663), .ZN(n2669) );
  NOR2_X1 U2614 ( .A1(n2670), .A2(n2671), .ZN(n2663) );
  INV_X1 U2615 ( .A(n2672), .ZN(n2671) );
  NAND3_X1 U2616 ( .A1(b_14_), .A2(n2673), .A3(a_6_), .ZN(n2672) );
  NAND2_X1 U2617 ( .A1(n2545), .A2(n2544), .ZN(n2673) );
  NOR2_X1 U2618 ( .A1(n2544), .A2(n2545), .ZN(n2670) );
  NOR2_X1 U2619 ( .A1(n2674), .A2(n2675), .ZN(n2545) );
  INV_X1 U2620 ( .A(n2676), .ZN(n2675) );
  NAND3_X1 U2621 ( .A1(b_14_), .A2(n2677), .A3(a_7_), .ZN(n2676) );
  NAND2_X1 U2622 ( .A1(n2553), .A2(n2551), .ZN(n2677) );
  NOR2_X1 U2623 ( .A1(n2551), .A2(n2553), .ZN(n2674) );
  NOR2_X1 U2624 ( .A1(n2678), .A2(n2679), .ZN(n2553) );
  NOR3_X1 U2625 ( .A1(n2207), .A2(n2680), .A3(n2681), .ZN(n2679) );
  NOR2_X1 U2626 ( .A1(n2561), .A2(n2559), .ZN(n2680) );
  INV_X1 U2627 ( .A(n2682), .ZN(n2678) );
  NAND2_X1 U2628 ( .A1(n2559), .A2(n2561), .ZN(n2682) );
  NAND2_X1 U2629 ( .A1(n2569), .A2(n2683), .ZN(n2561) );
  NAND2_X1 U2630 ( .A1(n2568), .A2(n2570), .ZN(n2683) );
  NAND2_X1 U2631 ( .A1(n2684), .A2(n2685), .ZN(n2570) );
  NAND2_X1 U2632 ( .A1(a_9_), .A2(b_14_), .ZN(n2684) );
  XNOR2_X1 U2633 ( .A(n2686), .B(n2687), .ZN(n2568) );
  NAND2_X1 U2634 ( .A1(n2688), .A2(n2689), .ZN(n2686) );
  NAND2_X1 U2635 ( .A1(n2690), .A2(a_9_), .ZN(n2569) );
  INV_X1 U2636 ( .A(n2685), .ZN(n2690) );
  NAND2_X1 U2637 ( .A1(n2691), .A2(n2692), .ZN(n2685) );
  NAND2_X1 U2638 ( .A1(n2611), .A2(n2693), .ZN(n2692) );
  INV_X1 U2639 ( .A(n2694), .ZN(n2693) );
  NOR2_X1 U2640 ( .A1(n2614), .A2(n2613), .ZN(n2694) );
  XOR2_X1 U2641 ( .A(n2695), .B(n2696), .Z(n2611) );
  XNOR2_X1 U2642 ( .A(n2697), .B(n2698), .ZN(n2695) );
  NOR2_X1 U2643 ( .A1(n2225), .A2(n2254), .ZN(n2698) );
  NAND2_X1 U2644 ( .A1(n2613), .A2(n2614), .ZN(n2691) );
  NAND2_X1 U2645 ( .A1(a_10_), .A2(b_14_), .ZN(n2614) );
  NOR2_X1 U2646 ( .A1(n2699), .A2(n2700), .ZN(n2613) );
  NOR3_X1 U2647 ( .A1(n2207), .A2(n2701), .A3(n2254), .ZN(n2700) );
  INV_X1 U2648 ( .A(n2702), .ZN(n2701) );
  NAND2_X1 U2649 ( .A1(n2610), .A2(n2608), .ZN(n2702) );
  NOR2_X1 U2650 ( .A1(n2608), .A2(n2610), .ZN(n2699) );
  NOR2_X1 U2651 ( .A1(n2703), .A2(n2704), .ZN(n2610) );
  INV_X1 U2652 ( .A(n2705), .ZN(n2704) );
  NAND2_X1 U2653 ( .A1(n2605), .A2(n2706), .ZN(n2705) );
  NAND2_X1 U2654 ( .A1(n2606), .A2(n2604), .ZN(n2706) );
  NOR2_X1 U2655 ( .A1(n2238), .A2(n2207), .ZN(n2605) );
  NOR2_X1 U2656 ( .A1(n2604), .A2(n2606), .ZN(n2703) );
  NOR2_X1 U2657 ( .A1(n2707), .A2(n2708), .ZN(n2606) );
  INV_X1 U2658 ( .A(n2709), .ZN(n2708) );
  NAND2_X1 U2659 ( .A1(n2600), .A2(n2710), .ZN(n2709) );
  NAND2_X1 U2660 ( .A1(n2601), .A2(n2602), .ZN(n2710) );
  NOR2_X1 U2661 ( .A1(n2223), .A2(n2207), .ZN(n2600) );
  NOR2_X1 U2662 ( .A1(n2602), .A2(n2601), .ZN(n2707) );
  INV_X1 U2663 ( .A(n2711), .ZN(n2601) );
  NAND2_X1 U2664 ( .A1(n2712), .A2(n2713), .ZN(n2711) );
  NAND2_X1 U2665 ( .A1(b_12_), .A2(n2714), .ZN(n2713) );
  NAND2_X1 U2666 ( .A1(n2202), .A2(n2715), .ZN(n2714) );
  NAND2_X1 U2667 ( .A1(a_15_), .A2(n2225), .ZN(n2715) );
  NAND2_X1 U2668 ( .A1(b_13_), .A2(n2716), .ZN(n2712) );
  NAND2_X1 U2669 ( .A1(n2205), .A2(n2717), .ZN(n2716) );
  NAND2_X1 U2670 ( .A1(a_14_), .A2(n2451), .ZN(n2717) );
  NAND3_X1 U2671 ( .A1(b_13_), .A2(b_14_), .A3(n2450), .ZN(n2602) );
  XNOR2_X1 U2672 ( .A(n2718), .B(n2220), .ZN(n2604) );
  XNOR2_X1 U2673 ( .A(n2719), .B(n2720), .ZN(n2718) );
  XNOR2_X1 U2674 ( .A(n2721), .B(n2722), .ZN(n2608) );
  XOR2_X1 U2675 ( .A(n2723), .B(n2724), .Z(n2721) );
  NOR2_X1 U2676 ( .A1(n2225), .A2(n2238), .ZN(n2724) );
  XNOR2_X1 U2677 ( .A(n2725), .B(n2726), .ZN(n2559) );
  NAND2_X1 U2678 ( .A1(n2727), .A2(n2728), .ZN(n2725) );
  XOR2_X1 U2679 ( .A(n2729), .B(n2730), .Z(n2551) );
  XOR2_X1 U2680 ( .A(n2731), .B(n2732), .Z(n2730) );
  NAND2_X1 U2681 ( .A1(a_8_), .A2(b_13_), .ZN(n2732) );
  XNOR2_X1 U2682 ( .A(n2733), .B(n2734), .ZN(n2544) );
  XNOR2_X1 U2683 ( .A(n2735), .B(n2736), .ZN(n2734) );
  NAND2_X1 U2684 ( .A1(a_7_), .A2(b_13_), .ZN(n2736) );
  XNOR2_X1 U2685 ( .A(n2737), .B(n2738), .ZN(n2620) );
  NAND2_X1 U2686 ( .A1(n2739), .A2(n2740), .ZN(n2737) );
  XOR2_X1 U2687 ( .A(n2741), .B(n2742), .Z(n2624) );
  XOR2_X1 U2688 ( .A(n2743), .B(n2744), .Z(n2742) );
  NAND2_X1 U2689 ( .A1(a_4_), .A2(b_13_), .ZN(n2744) );
  XOR2_X1 U2690 ( .A(n2745), .B(n2746), .Z(n2627) );
  NAND2_X1 U2691 ( .A1(n2747), .A2(n2748), .ZN(n2745) );
  XOR2_X1 U2692 ( .A(n2749), .B(n2750), .Z(n2631) );
  XOR2_X1 U2693 ( .A(n2751), .B(n2752), .Z(n2750) );
  XOR2_X1 U2694 ( .A(n2753), .B(n2754), .Z(n2636) );
  XOR2_X1 U2695 ( .A(n2755), .B(n2756), .Z(n2753) );
  XNOR2_X1 U2696 ( .A(n2757), .B(n2758), .ZN(n2469) );
  XOR2_X1 U2697 ( .A(n2759), .B(n2760), .Z(n2757) );
  NOR2_X1 U2698 ( .A1(n2639), .A2(n2640), .ZN(n2514) );
  NOR2_X1 U2699 ( .A1(n2761), .A2(n2762), .ZN(n2640) );
  INV_X1 U2700 ( .A(n2763), .ZN(n2762) );
  NAND2_X1 U2701 ( .A1(n2760), .A2(n2764), .ZN(n2763) );
  NAND2_X1 U2702 ( .A1(n2765), .A2(n2758), .ZN(n2764) );
  NOR2_X1 U2703 ( .A1(n2420), .A2(n2225), .ZN(n2760) );
  NOR2_X1 U2704 ( .A1(n2758), .A2(n2765), .ZN(n2761) );
  INV_X1 U2705 ( .A(n2759), .ZN(n2765) );
  NAND2_X1 U2706 ( .A1(n2766), .A2(n2767), .ZN(n2759) );
  NAND2_X1 U2707 ( .A1(n2756), .A2(n2768), .ZN(n2767) );
  NAND2_X1 U2708 ( .A1(n2754), .A2(n2769), .ZN(n2768) );
  INV_X1 U2709 ( .A(n2755), .ZN(n2769) );
  NOR2_X1 U2710 ( .A1(n2225), .A2(n2647), .ZN(n2756) );
  NAND2_X1 U2711 ( .A1(n2770), .A2(n2755), .ZN(n2766) );
  NAND2_X1 U2712 ( .A1(n2771), .A2(n2772), .ZN(n2755) );
  INV_X1 U2713 ( .A(n2773), .ZN(n2772) );
  NOR2_X1 U2714 ( .A1(n2752), .A2(n2774), .ZN(n2773) );
  NOR2_X1 U2715 ( .A1(n2749), .A2(n2751), .ZN(n2774) );
  NAND2_X1 U2716 ( .A1(a_2_), .A2(b_13_), .ZN(n2752) );
  NAND2_X1 U2717 ( .A1(n2749), .A2(n2751), .ZN(n2771) );
  NAND2_X1 U2718 ( .A1(n2747), .A2(n2775), .ZN(n2751) );
  NAND2_X1 U2719 ( .A1(n2746), .A2(n2748), .ZN(n2775) );
  NAND2_X1 U2720 ( .A1(n2776), .A2(n2777), .ZN(n2748) );
  NAND2_X1 U2721 ( .A1(a_3_), .A2(b_13_), .ZN(n2777) );
  INV_X1 U2722 ( .A(n2778), .ZN(n2776) );
  XNOR2_X1 U2723 ( .A(n2779), .B(n2780), .ZN(n2746) );
  XOR2_X1 U2724 ( .A(n2781), .B(n2782), .Z(n2780) );
  NAND2_X1 U2725 ( .A1(a_4_), .A2(b_12_), .ZN(n2782) );
  NAND2_X1 U2726 ( .A1(a_3_), .A2(n2778), .ZN(n2747) );
  NAND2_X1 U2727 ( .A1(n2783), .A2(n2784), .ZN(n2778) );
  NAND3_X1 U2728 ( .A1(b_13_), .A2(n2785), .A3(a_4_), .ZN(n2784) );
  INV_X1 U2729 ( .A(n2786), .ZN(n2785) );
  NOR2_X1 U2730 ( .A1(n2743), .A2(n2741), .ZN(n2786) );
  NAND2_X1 U2731 ( .A1(n2741), .A2(n2743), .ZN(n2783) );
  NAND2_X1 U2732 ( .A1(n2739), .A2(n2787), .ZN(n2743) );
  NAND2_X1 U2733 ( .A1(n2738), .A2(n2740), .ZN(n2787) );
  NAND2_X1 U2734 ( .A1(n2788), .A2(n2789), .ZN(n2740) );
  NAND2_X1 U2735 ( .A1(a_5_), .A2(b_13_), .ZN(n2789) );
  XNOR2_X1 U2736 ( .A(n2790), .B(n2791), .ZN(n2738) );
  XOR2_X1 U2737 ( .A(n2792), .B(n2793), .Z(n2791) );
  NAND2_X1 U2738 ( .A1(a_6_), .A2(b_12_), .ZN(n2793) );
  NAND2_X1 U2739 ( .A1(a_5_), .A2(n2794), .ZN(n2739) );
  INV_X1 U2740 ( .A(n2788), .ZN(n2794) );
  NOR2_X1 U2741 ( .A1(n2795), .A2(n2796), .ZN(n2788) );
  NOR3_X1 U2742 ( .A1(n2225), .A2(n2797), .A3(n2455), .ZN(n2796) );
  NOR2_X1 U2743 ( .A1(n2665), .A2(n2667), .ZN(n2797) );
  INV_X1 U2744 ( .A(n2798), .ZN(n2795) );
  NAND2_X1 U2745 ( .A1(n2665), .A2(n2667), .ZN(n2798) );
  NAND2_X1 U2746 ( .A1(n2799), .A2(n2800), .ZN(n2667) );
  NAND3_X1 U2747 ( .A1(b_13_), .A2(n2801), .A3(a_7_), .ZN(n2800) );
  NAND2_X1 U2748 ( .A1(n2733), .A2(n2735), .ZN(n2801) );
  INV_X1 U2749 ( .A(n2802), .ZN(n2799) );
  NOR2_X1 U2750 ( .A1(n2733), .A2(n2735), .ZN(n2802) );
  NOR2_X1 U2751 ( .A1(n2803), .A2(n2804), .ZN(n2735) );
  NOR3_X1 U2752 ( .A1(n2225), .A2(n2805), .A3(n2681), .ZN(n2804) );
  NOR2_X1 U2753 ( .A1(n2731), .A2(n2729), .ZN(n2805) );
  INV_X1 U2754 ( .A(n2806), .ZN(n2803) );
  NAND2_X1 U2755 ( .A1(n2729), .A2(n2731), .ZN(n2806) );
  NAND2_X1 U2756 ( .A1(n2727), .A2(n2807), .ZN(n2731) );
  NAND2_X1 U2757 ( .A1(n2726), .A2(n2728), .ZN(n2807) );
  NAND2_X1 U2758 ( .A1(n2808), .A2(n2809), .ZN(n2728) );
  NAND2_X1 U2759 ( .A1(a_9_), .A2(b_13_), .ZN(n2809) );
  INV_X1 U2760 ( .A(n2810), .ZN(n2808) );
  XNOR2_X1 U2761 ( .A(n2811), .B(n2812), .ZN(n2726) );
  NAND2_X1 U2762 ( .A1(n2813), .A2(n2814), .ZN(n2811) );
  NAND2_X1 U2763 ( .A1(a_9_), .A2(n2810), .ZN(n2727) );
  NAND2_X1 U2764 ( .A1(n2688), .A2(n2815), .ZN(n2810) );
  NAND2_X1 U2765 ( .A1(n2687), .A2(n2689), .ZN(n2815) );
  NAND2_X1 U2766 ( .A1(n2816), .A2(n2817), .ZN(n2689) );
  NAND2_X1 U2767 ( .A1(a_10_), .A2(b_13_), .ZN(n2817) );
  XNOR2_X1 U2768 ( .A(n2818), .B(n2819), .ZN(n2687) );
  XOR2_X1 U2769 ( .A(n2820), .B(n2821), .Z(n2819) );
  NAND2_X1 U2770 ( .A1(a_11_), .A2(b_12_), .ZN(n2821) );
  NAND2_X1 U2771 ( .A1(a_10_), .A2(n2822), .ZN(n2688) );
  INV_X1 U2772 ( .A(n2816), .ZN(n2822) );
  NOR2_X1 U2773 ( .A1(n2823), .A2(n2824), .ZN(n2816) );
  INV_X1 U2774 ( .A(n2825), .ZN(n2824) );
  NAND3_X1 U2775 ( .A1(b_13_), .A2(n2826), .A3(a_11_), .ZN(n2825) );
  NAND2_X1 U2776 ( .A1(n2696), .A2(n2697), .ZN(n2826) );
  NOR2_X1 U2777 ( .A1(n2696), .A2(n2697), .ZN(n2823) );
  NOR2_X1 U2778 ( .A1(n2827), .A2(n2828), .ZN(n2697) );
  NOR3_X1 U2779 ( .A1(n2225), .A2(n2829), .A3(n2238), .ZN(n2828) );
  INV_X1 U2780 ( .A(n2830), .ZN(n2829) );
  NAND2_X1 U2781 ( .A1(n2722), .A2(n2723), .ZN(n2830) );
  NOR2_X1 U2782 ( .A1(n2722), .A2(n2723), .ZN(n2827) );
  NAND2_X1 U2783 ( .A1(n2831), .A2(n2832), .ZN(n2723) );
  NAND2_X1 U2784 ( .A1(n2833), .A2(n2720), .ZN(n2832) );
  NAND3_X1 U2785 ( .A1(b_12_), .A2(b_13_), .A3(n2450), .ZN(n2720) );
  NAND2_X1 U2786 ( .A1(n2220), .A2(n2719), .ZN(n2833) );
  INV_X1 U2787 ( .A(n2443), .ZN(n2220) );
  NAND2_X1 U2788 ( .A1(n2834), .A2(n2443), .ZN(n2831) );
  NAND2_X1 U2789 ( .A1(a_13_), .A2(b_13_), .ZN(n2443) );
  INV_X1 U2790 ( .A(n2719), .ZN(n2834) );
  NAND2_X1 U2791 ( .A1(n2835), .A2(n2836), .ZN(n2719) );
  NAND2_X1 U2792 ( .A1(b_11_), .A2(n2837), .ZN(n2836) );
  NAND2_X1 U2793 ( .A1(n2202), .A2(n2838), .ZN(n2837) );
  NAND2_X1 U2794 ( .A1(a_15_), .A2(n2451), .ZN(n2838) );
  NAND2_X1 U2795 ( .A1(b_12_), .A2(n2839), .ZN(n2835) );
  NAND2_X1 U2796 ( .A1(n2205), .A2(n2840), .ZN(n2839) );
  NAND2_X1 U2797 ( .A1(a_14_), .A2(n2256), .ZN(n2840) );
  XNOR2_X1 U2798 ( .A(n2841), .B(n2842), .ZN(n2722) );
  XOR2_X1 U2799 ( .A(n2843), .B(n2844), .Z(n2841) );
  XOR2_X1 U2800 ( .A(n2845), .B(n2846), .Z(n2696) );
  XOR2_X1 U2801 ( .A(n2242), .B(n2847), .Z(n2845) );
  XNOR2_X1 U2802 ( .A(n2848), .B(n2849), .ZN(n2729) );
  NAND2_X1 U2803 ( .A1(n2850), .A2(n2851), .ZN(n2848) );
  XNOR2_X1 U2804 ( .A(n2852), .B(n2853), .ZN(n2733) );
  XOR2_X1 U2805 ( .A(n2854), .B(n2855), .Z(n2852) );
  NOR2_X1 U2806 ( .A1(n2451), .A2(n2681), .ZN(n2855) );
  XNOR2_X1 U2807 ( .A(n2856), .B(n2857), .ZN(n2665) );
  XOR2_X1 U2808 ( .A(n2858), .B(n2859), .Z(n2857) );
  NAND2_X1 U2809 ( .A1(a_7_), .A2(b_12_), .ZN(n2859) );
  XNOR2_X1 U2810 ( .A(n2860), .B(n2861), .ZN(n2741) );
  NAND2_X1 U2811 ( .A1(n2862), .A2(n2863), .ZN(n2860) );
  XNOR2_X1 U2812 ( .A(n2864), .B(n2865), .ZN(n2749) );
  NAND2_X1 U2813 ( .A1(n2866), .A2(n2867), .ZN(n2864) );
  INV_X1 U2814 ( .A(n2754), .ZN(n2770) );
  XNOR2_X1 U2815 ( .A(n2868), .B(n2869), .ZN(n2754) );
  XNOR2_X1 U2816 ( .A(n2870), .B(n2871), .ZN(n2868) );
  NAND2_X1 U2817 ( .A1(a_2_), .A2(b_12_), .ZN(n2870) );
  XNOR2_X1 U2818 ( .A(n2872), .B(n2873), .ZN(n2758) );
  XOR2_X1 U2819 ( .A(n2874), .B(n2875), .Z(n2873) );
  XNOR2_X1 U2820 ( .A(n2876), .B(n2877), .ZN(n2639) );
  XOR2_X1 U2821 ( .A(n2878), .B(n2879), .Z(n2876) );
  INV_X1 U2822 ( .A(n2880), .ZN(n2485) );
  INV_X1 U2823 ( .A(n2484), .ZN(n2512) );
  NAND3_X1 U2824 ( .A1(n2487), .A2(n2488), .A3(n2880), .ZN(n2484) );
  NOR2_X1 U2825 ( .A1(n2511), .A2(n2881), .ZN(n2880) );
  INV_X1 U2826 ( .A(n2882), .ZN(n2881) );
  NAND2_X1 U2827 ( .A1(n2883), .A2(n2884), .ZN(n2882) );
  NAND2_X1 U2828 ( .A1(n2885), .A2(n2886), .ZN(n2488) );
  NAND2_X1 U2829 ( .A1(n2879), .A2(n2887), .ZN(n2886) );
  INV_X1 U2830 ( .A(n2888), .ZN(n2887) );
  NOR2_X1 U2831 ( .A1(n2878), .A2(n2877), .ZN(n2888) );
  NOR2_X1 U2832 ( .A1(n2420), .A2(n2451), .ZN(n2879) );
  NAND2_X1 U2833 ( .A1(n2877), .A2(n2878), .ZN(n2885) );
  NAND2_X1 U2834 ( .A1(n2889), .A2(n2890), .ZN(n2878) );
  NAND2_X1 U2835 ( .A1(n2875), .A2(n2891), .ZN(n2890) );
  NAND2_X1 U2836 ( .A1(n2874), .A2(n2872), .ZN(n2891) );
  NOR2_X1 U2837 ( .A1(n2451), .A2(n2647), .ZN(n2875) );
  INV_X1 U2838 ( .A(n2892), .ZN(n2889) );
  NOR2_X1 U2839 ( .A1(n2872), .A2(n2874), .ZN(n2892) );
  NOR2_X1 U2840 ( .A1(n2893), .A2(n2894), .ZN(n2874) );
  NOR3_X1 U2841 ( .A1(n2451), .A2(n2895), .A3(n2460), .ZN(n2894) );
  NOR2_X1 U2842 ( .A1(n2871), .A2(n2869), .ZN(n2895) );
  INV_X1 U2843 ( .A(n2896), .ZN(n2893) );
  NAND2_X1 U2844 ( .A1(n2869), .A2(n2871), .ZN(n2896) );
  NAND2_X1 U2845 ( .A1(n2866), .A2(n2897), .ZN(n2871) );
  NAND2_X1 U2846 ( .A1(n2865), .A2(n2867), .ZN(n2897) );
  NAND2_X1 U2847 ( .A1(n2898), .A2(n2899), .ZN(n2867) );
  NAND2_X1 U2848 ( .A1(a_3_), .A2(b_12_), .ZN(n2899) );
  XNOR2_X1 U2849 ( .A(n2900), .B(n2901), .ZN(n2865) );
  XOR2_X1 U2850 ( .A(n2902), .B(n2903), .Z(n2901) );
  NAND2_X1 U2851 ( .A1(a_4_), .A2(b_11_), .ZN(n2903) );
  NAND2_X1 U2852 ( .A1(a_3_), .A2(n2904), .ZN(n2866) );
  INV_X1 U2853 ( .A(n2898), .ZN(n2904) );
  NOR2_X1 U2854 ( .A1(n2905), .A2(n2906), .ZN(n2898) );
  NOR3_X1 U2855 ( .A1(n2451), .A2(n2907), .A3(n2457), .ZN(n2906) );
  NOR2_X1 U2856 ( .A1(n2781), .A2(n2779), .ZN(n2907) );
  INV_X1 U2857 ( .A(n2908), .ZN(n2905) );
  NAND2_X1 U2858 ( .A1(n2779), .A2(n2781), .ZN(n2908) );
  NAND2_X1 U2859 ( .A1(n2862), .A2(n2909), .ZN(n2781) );
  NAND2_X1 U2860 ( .A1(n2861), .A2(n2863), .ZN(n2909) );
  NAND2_X1 U2861 ( .A1(n2910), .A2(n2911), .ZN(n2863) );
  NAND2_X1 U2862 ( .A1(a_5_), .A2(b_12_), .ZN(n2911) );
  XOR2_X1 U2863 ( .A(n2912), .B(n2913), .Z(n2861) );
  XNOR2_X1 U2864 ( .A(n2914), .B(n2915), .ZN(n2913) );
  NAND2_X1 U2865 ( .A1(a_6_), .A2(b_11_), .ZN(n2915) );
  NAND2_X1 U2866 ( .A1(a_5_), .A2(n2916), .ZN(n2862) );
  INV_X1 U2867 ( .A(n2910), .ZN(n2916) );
  NOR2_X1 U2868 ( .A1(n2917), .A2(n2918), .ZN(n2910) );
  NOR3_X1 U2869 ( .A1(n2451), .A2(n2919), .A3(n2455), .ZN(n2918) );
  NOR2_X1 U2870 ( .A1(n2792), .A2(n2790), .ZN(n2919) );
  INV_X1 U2871 ( .A(n2920), .ZN(n2917) );
  NAND2_X1 U2872 ( .A1(n2790), .A2(n2792), .ZN(n2920) );
  NAND2_X1 U2873 ( .A1(n2921), .A2(n2922), .ZN(n2792) );
  INV_X1 U2874 ( .A(n2923), .ZN(n2922) );
  NOR3_X1 U2875 ( .A1(n2451), .A2(n2924), .A3(n2312), .ZN(n2923) );
  NOR2_X1 U2876 ( .A1(n2858), .A2(n2856), .ZN(n2924) );
  NAND2_X1 U2877 ( .A1(n2856), .A2(n2858), .ZN(n2921) );
  NAND2_X1 U2878 ( .A1(n2925), .A2(n2926), .ZN(n2858) );
  INV_X1 U2879 ( .A(n2927), .ZN(n2926) );
  NOR3_X1 U2880 ( .A1(n2451), .A2(n2928), .A3(n2681), .ZN(n2927) );
  NOR2_X1 U2881 ( .A1(n2854), .A2(n2853), .ZN(n2928) );
  NAND2_X1 U2882 ( .A1(n2853), .A2(n2854), .ZN(n2925) );
  NAND2_X1 U2883 ( .A1(n2850), .A2(n2929), .ZN(n2854) );
  NAND2_X1 U2884 ( .A1(n2849), .A2(n2851), .ZN(n2929) );
  NAND2_X1 U2885 ( .A1(n2930), .A2(n2931), .ZN(n2851) );
  NAND2_X1 U2886 ( .A1(a_9_), .A2(b_12_), .ZN(n2931) );
  INV_X1 U2887 ( .A(n2932), .ZN(n2930) );
  XNOR2_X1 U2888 ( .A(n2933), .B(n2934), .ZN(n2849) );
  NAND2_X1 U2889 ( .A1(n2935), .A2(n2936), .ZN(n2933) );
  NAND2_X1 U2890 ( .A1(a_9_), .A2(n2932), .ZN(n2850) );
  NAND2_X1 U2891 ( .A1(n2813), .A2(n2937), .ZN(n2932) );
  NAND2_X1 U2892 ( .A1(n2812), .A2(n2814), .ZN(n2937) );
  NAND2_X1 U2893 ( .A1(n2938), .A2(n2939), .ZN(n2814) );
  NAND2_X1 U2894 ( .A1(a_10_), .A2(b_12_), .ZN(n2939) );
  XOR2_X1 U2895 ( .A(n2940), .B(n2941), .Z(n2812) );
  XOR2_X1 U2896 ( .A(n2252), .B(n2942), .Z(n2940) );
  INV_X1 U2897 ( .A(n2943), .ZN(n2813) );
  NOR2_X1 U2898 ( .A1(n2453), .A2(n2938), .ZN(n2943) );
  NOR2_X1 U2899 ( .A1(n2944), .A2(n2945), .ZN(n2938) );
  INV_X1 U2900 ( .A(n2946), .ZN(n2945) );
  NAND3_X1 U2901 ( .A1(b_12_), .A2(n2947), .A3(a_11_), .ZN(n2946) );
  NAND2_X1 U2902 ( .A1(n2818), .A2(n2820), .ZN(n2947) );
  NOR2_X1 U2903 ( .A1(n2820), .A2(n2818), .ZN(n2944) );
  XOR2_X1 U2904 ( .A(n2948), .B(n2949), .Z(n2818) );
  XNOR2_X1 U2905 ( .A(n2950), .B(n2951), .ZN(n2948) );
  NAND2_X1 U2906 ( .A1(n2952), .A2(n2953), .ZN(n2820) );
  NAND2_X1 U2907 ( .A1(n2846), .A2(n2954), .ZN(n2953) );
  NAND2_X1 U2908 ( .A1(n2955), .A2(n2956), .ZN(n2954) );
  INV_X1 U2909 ( .A(n2242), .ZN(n2955) );
  XNOR2_X1 U2910 ( .A(n2957), .B(n2958), .ZN(n2846) );
  XOR2_X1 U2911 ( .A(n2959), .B(n2960), .Z(n2957) );
  NAND2_X1 U2912 ( .A1(n2847), .A2(n2242), .ZN(n2952) );
  NAND2_X1 U2913 ( .A1(b_12_), .A2(a_12_), .ZN(n2242) );
  INV_X1 U2914 ( .A(n2956), .ZN(n2847) );
  NAND2_X1 U2915 ( .A1(n2961), .A2(n2962), .ZN(n2956) );
  NAND2_X1 U2916 ( .A1(n2842), .A2(n2963), .ZN(n2962) );
  INV_X1 U2917 ( .A(n2964), .ZN(n2963) );
  NOR2_X1 U2918 ( .A1(n2843), .A2(n2844), .ZN(n2964) );
  NOR2_X1 U2919 ( .A1(n2451), .A2(n2223), .ZN(n2842) );
  NAND2_X1 U2920 ( .A1(n2844), .A2(n2843), .ZN(n2961) );
  NAND2_X1 U2921 ( .A1(n2965), .A2(n2966), .ZN(n2843) );
  NAND2_X1 U2922 ( .A1(b_10_), .A2(n2967), .ZN(n2966) );
  NAND2_X1 U2923 ( .A1(n2202), .A2(n2968), .ZN(n2967) );
  NAND2_X1 U2924 ( .A1(a_15_), .A2(n2256), .ZN(n2968) );
  NAND2_X1 U2925 ( .A1(b_11_), .A2(n2969), .ZN(n2965) );
  NAND2_X1 U2926 ( .A1(n2205), .A2(n2970), .ZN(n2969) );
  NAND2_X1 U2927 ( .A1(a_14_), .A2(n2452), .ZN(n2970) );
  NOR3_X1 U2928 ( .A1(n2451), .A2(n2256), .A3(n2598), .ZN(n2844) );
  XOR2_X1 U2929 ( .A(n2971), .B(n2972), .Z(n2853) );
  XNOR2_X1 U2930 ( .A(n2973), .B(n2974), .ZN(n2972) );
  XOR2_X1 U2931 ( .A(n2975), .B(n2976), .Z(n2856) );
  XOR2_X1 U2932 ( .A(n2977), .B(n2978), .Z(n2976) );
  NAND2_X1 U2933 ( .A1(a_8_), .A2(b_11_), .ZN(n2978) );
  XOR2_X1 U2934 ( .A(n2979), .B(n2980), .Z(n2790) );
  XOR2_X1 U2935 ( .A(n2981), .B(n2982), .Z(n2979) );
  NOR2_X1 U2936 ( .A1(n2256), .A2(n2312), .ZN(n2982) );
  XNOR2_X1 U2937 ( .A(n2983), .B(n2984), .ZN(n2779) );
  NAND2_X1 U2938 ( .A1(n2985), .A2(n2986), .ZN(n2983) );
  XNOR2_X1 U2939 ( .A(n2987), .B(n2988), .ZN(n2869) );
  NAND2_X1 U2940 ( .A1(n2989), .A2(n2990), .ZN(n2987) );
  XOR2_X1 U2941 ( .A(n2991), .B(n2992), .Z(n2872) );
  XOR2_X1 U2942 ( .A(n2993), .B(n2994), .Z(n2992) );
  NAND2_X1 U2943 ( .A1(a_2_), .A2(b_11_), .ZN(n2994) );
  XNOR2_X1 U2944 ( .A(n2995), .B(n2996), .ZN(n2877) );
  XOR2_X1 U2945 ( .A(n2997), .B(n2998), .Z(n2996) );
  NAND2_X1 U2946 ( .A1(b_11_), .A2(a_1_), .ZN(n2998) );
  XOR2_X1 U2947 ( .A(n2999), .B(n3000), .Z(n2487) );
  XOR2_X1 U2948 ( .A(n3001), .B(n3002), .Z(n2999) );
  NOR2_X1 U2949 ( .A1(n2256), .A2(n2420), .ZN(n3002) );
  NOR2_X1 U2950 ( .A1(n2884), .A2(n2883), .ZN(n2511) );
  NOR2_X1 U2951 ( .A1(n3003), .A2(n3004), .ZN(n2883) );
  NOR3_X1 U2952 ( .A1(n2256), .A2(n3005), .A3(n2420), .ZN(n3004) );
  NOR2_X1 U2953 ( .A1(n3001), .A2(n3000), .ZN(n3005) );
  INV_X1 U2954 ( .A(n3006), .ZN(n3003) );
  NAND2_X1 U2955 ( .A1(n3000), .A2(n3001), .ZN(n3006) );
  NAND2_X1 U2956 ( .A1(n3007), .A2(n3008), .ZN(n3001) );
  INV_X1 U2957 ( .A(n3009), .ZN(n3008) );
  NOR3_X1 U2958 ( .A1(n2647), .A2(n3010), .A3(n2256), .ZN(n3009) );
  NOR2_X1 U2959 ( .A1(n2995), .A2(n2997), .ZN(n3010) );
  NAND2_X1 U2960 ( .A1(n2995), .A2(n2997), .ZN(n3007) );
  NAND2_X1 U2961 ( .A1(n3011), .A2(n3012), .ZN(n2997) );
  INV_X1 U2962 ( .A(n3013), .ZN(n3012) );
  NOR3_X1 U2963 ( .A1(n2256), .A2(n3014), .A3(n2460), .ZN(n3013) );
  NOR2_X1 U2964 ( .A1(n2993), .A2(n2991), .ZN(n3014) );
  NAND2_X1 U2965 ( .A1(n2991), .A2(n2993), .ZN(n3011) );
  NAND2_X1 U2966 ( .A1(n2989), .A2(n3015), .ZN(n2993) );
  NAND2_X1 U2967 ( .A1(n2988), .A2(n2990), .ZN(n3015) );
  NAND2_X1 U2968 ( .A1(n3016), .A2(n3017), .ZN(n2990) );
  NAND2_X1 U2969 ( .A1(a_3_), .A2(b_11_), .ZN(n3017) );
  XNOR2_X1 U2970 ( .A(n3018), .B(n3019), .ZN(n2988) );
  XOR2_X1 U2971 ( .A(n3020), .B(n3021), .Z(n3019) );
  NAND2_X1 U2972 ( .A1(a_4_), .A2(b_10_), .ZN(n3021) );
  NAND2_X1 U2973 ( .A1(a_3_), .A2(n3022), .ZN(n2989) );
  INV_X1 U2974 ( .A(n3016), .ZN(n3022) );
  NOR2_X1 U2975 ( .A1(n3023), .A2(n3024), .ZN(n3016) );
  NOR3_X1 U2976 ( .A1(n2256), .A2(n3025), .A3(n2457), .ZN(n3024) );
  NOR2_X1 U2977 ( .A1(n2902), .A2(n2900), .ZN(n3025) );
  INV_X1 U2978 ( .A(n3026), .ZN(n3023) );
  NAND2_X1 U2979 ( .A1(n2900), .A2(n2902), .ZN(n3026) );
  NAND2_X1 U2980 ( .A1(n2985), .A2(n3027), .ZN(n2902) );
  NAND2_X1 U2981 ( .A1(n2984), .A2(n2986), .ZN(n3027) );
  NAND2_X1 U2982 ( .A1(n3028), .A2(n3029), .ZN(n2986) );
  NAND2_X1 U2983 ( .A1(a_5_), .A2(b_11_), .ZN(n3029) );
  INV_X1 U2984 ( .A(n3030), .ZN(n3028) );
  XNOR2_X1 U2985 ( .A(n3031), .B(n3032), .ZN(n2984) );
  XNOR2_X1 U2986 ( .A(n3033), .B(n3034), .ZN(n3031) );
  NOR2_X1 U2987 ( .A1(n2452), .A2(n2455), .ZN(n3034) );
  NAND2_X1 U2988 ( .A1(a_5_), .A2(n3030), .ZN(n2985) );
  NAND2_X1 U2989 ( .A1(n3035), .A2(n3036), .ZN(n3030) );
  NAND3_X1 U2990 ( .A1(b_11_), .A2(n3037), .A3(a_6_), .ZN(n3036) );
  NAND2_X1 U2991 ( .A1(n2912), .A2(n2914), .ZN(n3037) );
  INV_X1 U2992 ( .A(n3038), .ZN(n3035) );
  NOR2_X1 U2993 ( .A1(n2912), .A2(n2914), .ZN(n3038) );
  NOR2_X1 U2994 ( .A1(n3039), .A2(n3040), .ZN(n2914) );
  NOR3_X1 U2995 ( .A1(n2256), .A2(n3041), .A3(n2312), .ZN(n3040) );
  NOR2_X1 U2996 ( .A1(n2981), .A2(n2980), .ZN(n3041) );
  INV_X1 U2997 ( .A(n3042), .ZN(n3039) );
  NAND2_X1 U2998 ( .A1(n2980), .A2(n2981), .ZN(n3042) );
  NAND2_X1 U2999 ( .A1(n3043), .A2(n3044), .ZN(n2981) );
  NAND3_X1 U3000 ( .A1(b_11_), .A2(n3045), .A3(a_8_), .ZN(n3044) );
  NAND2_X1 U3001 ( .A1(n3046), .A2(n2977), .ZN(n3045) );
  INV_X1 U3002 ( .A(n2975), .ZN(n3046) );
  NAND2_X1 U3003 ( .A1(n2975), .A2(n3047), .ZN(n3043) );
  INV_X1 U3004 ( .A(n2977), .ZN(n3047) );
  NAND2_X1 U3005 ( .A1(n3048), .A2(n3049), .ZN(n2977) );
  NAND2_X1 U3006 ( .A1(n2971), .A2(n3050), .ZN(n3049) );
  NAND2_X1 U3007 ( .A1(n2974), .A2(n2973), .ZN(n3050) );
  XNOR2_X1 U3008 ( .A(n3051), .B(n3052), .ZN(n2971) );
  XNOR2_X1 U3009 ( .A(n3053), .B(n2273), .ZN(n3052) );
  INV_X1 U3010 ( .A(n3054), .ZN(n3048) );
  NOR2_X1 U3011 ( .A1(n2973), .A2(n2974), .ZN(n3054) );
  NOR2_X1 U3012 ( .A1(n2283), .A2(n2256), .ZN(n2974) );
  NAND2_X1 U3013 ( .A1(n2935), .A2(n3055), .ZN(n2973) );
  NAND2_X1 U3014 ( .A1(n2934), .A2(n2936), .ZN(n3055) );
  NAND2_X1 U3015 ( .A1(n3056), .A2(n3057), .ZN(n2936) );
  NAND2_X1 U3016 ( .A1(a_10_), .A2(b_11_), .ZN(n3056) );
  XNOR2_X1 U3017 ( .A(n3058), .B(n3059), .ZN(n2934) );
  XOR2_X1 U3018 ( .A(n3060), .B(n3061), .Z(n3058) );
  NAND2_X1 U3019 ( .A1(b_10_), .A2(a_11_), .ZN(n3060) );
  NAND2_X1 U3020 ( .A1(n3062), .A2(a_10_), .ZN(n2935) );
  INV_X1 U3021 ( .A(n3057), .ZN(n3062) );
  NAND2_X1 U3022 ( .A1(n3063), .A2(n3064), .ZN(n3057) );
  INV_X1 U3023 ( .A(n3065), .ZN(n3064) );
  NOR2_X1 U3024 ( .A1(n2941), .A2(n3066), .ZN(n3065) );
  NOR2_X1 U3025 ( .A1(n2252), .A2(n2942), .ZN(n3066) );
  XNOR2_X1 U3026 ( .A(n3067), .B(n3068), .ZN(n2941) );
  XNOR2_X1 U3027 ( .A(n3069), .B(n3070), .ZN(n3067) );
  NAND2_X1 U3028 ( .A1(n2942), .A2(n2252), .ZN(n3063) );
  NAND2_X1 U3029 ( .A1(a_11_), .A2(b_11_), .ZN(n2252) );
  NOR2_X1 U3030 ( .A1(n3071), .A2(n3072), .ZN(n2942) );
  INV_X1 U3031 ( .A(n3073), .ZN(n3072) );
  NAND2_X1 U3032 ( .A1(n2950), .A2(n3074), .ZN(n3073) );
  NAND2_X1 U3033 ( .A1(n2951), .A2(n2949), .ZN(n3074) );
  NOR2_X1 U3034 ( .A1(n2256), .A2(n2238), .ZN(n2950) );
  NOR2_X1 U3035 ( .A1(n2949), .A2(n2951), .ZN(n3071) );
  NOR2_X1 U3036 ( .A1(n3075), .A2(n3076), .ZN(n2951) );
  INV_X1 U3037 ( .A(n3077), .ZN(n3076) );
  NAND2_X1 U3038 ( .A1(n2958), .A2(n3078), .ZN(n3077) );
  NAND2_X1 U3039 ( .A1(n2959), .A2(n2960), .ZN(n3078) );
  NOR2_X1 U3040 ( .A1(n2256), .A2(n2223), .ZN(n2958) );
  NOR2_X1 U3041 ( .A1(n2960), .A2(n2959), .ZN(n3075) );
  INV_X1 U3042 ( .A(n3079), .ZN(n2959) );
  NAND2_X1 U3043 ( .A1(n3080), .A2(n3081), .ZN(n3079) );
  NAND2_X1 U3044 ( .A1(b_10_), .A2(n3082), .ZN(n3081) );
  NAND2_X1 U3045 ( .A1(n2205), .A2(n3083), .ZN(n3082) );
  NAND2_X1 U3046 ( .A1(a_14_), .A2(n2285), .ZN(n3083) );
  NAND2_X1 U3047 ( .A1(b_9_), .A2(n3084), .ZN(n3080) );
  NAND2_X1 U3048 ( .A1(n2202), .A2(n3085), .ZN(n3084) );
  NAND2_X1 U3049 ( .A1(a_15_), .A2(n2452), .ZN(n3085) );
  NAND3_X1 U3050 ( .A1(b_10_), .A2(b_11_), .A3(n2450), .ZN(n2960) );
  XNOR2_X1 U3051 ( .A(n3086), .B(n3087), .ZN(n2949) );
  XOR2_X1 U3052 ( .A(n3088), .B(n3089), .Z(n3086) );
  XNOR2_X1 U3053 ( .A(n3090), .B(n3091), .ZN(n2975) );
  NAND2_X1 U3054 ( .A1(n3092), .A2(n3093), .ZN(n3090) );
  XNOR2_X1 U3055 ( .A(n3094), .B(n3095), .ZN(n2980) );
  XOR2_X1 U3056 ( .A(n3096), .B(n3097), .Z(n3095) );
  NAND2_X1 U3057 ( .A1(a_8_), .A2(b_10_), .ZN(n3097) );
  XOR2_X1 U3058 ( .A(n3098), .B(n3099), .Z(n2912) );
  XOR2_X1 U3059 ( .A(n3100), .B(n3101), .Z(n3099) );
  NAND2_X1 U3060 ( .A1(a_7_), .A2(b_10_), .ZN(n3101) );
  XNOR2_X1 U3061 ( .A(n3102), .B(n3103), .ZN(n2900) );
  NAND2_X1 U3062 ( .A1(n3104), .A2(n3105), .ZN(n3102) );
  XNOR2_X1 U3063 ( .A(n3106), .B(n3107), .ZN(n2991) );
  XNOR2_X1 U3064 ( .A(n3108), .B(n3109), .ZN(n3106) );
  XOR2_X1 U3065 ( .A(n3110), .B(n3111), .Z(n2995) );
  XNOR2_X1 U3066 ( .A(n3112), .B(n3113), .ZN(n3111) );
  NAND2_X1 U3067 ( .A1(a_2_), .A2(b_10_), .ZN(n3113) );
  XNOR2_X1 U3068 ( .A(n3114), .B(n3115), .ZN(n3000) );
  NAND2_X1 U3069 ( .A1(n3116), .A2(n3117), .ZN(n3114) );
  XNOR2_X1 U3070 ( .A(n3118), .B(n3119), .ZN(n2884) );
  XNOR2_X1 U3071 ( .A(n3120), .B(n3121), .ZN(n3119) );
  INV_X1 U3072 ( .A(n3122), .ZN(n2150) );
  INV_X1 U3073 ( .A(n2149), .ZN(n2509) );
  NAND3_X1 U3074 ( .A1(n2153), .A2(n3122), .A3(n2152), .ZN(n2149) );
  NOR2_X1 U3075 ( .A1(n3123), .A2(n3124), .ZN(n2152) );
  INV_X1 U3076 ( .A(n3125), .ZN(n3124) );
  NAND2_X1 U3077 ( .A1(n3118), .A2(n3126), .ZN(n3125) );
  NAND2_X1 U3078 ( .A1(n3121), .A2(n3120), .ZN(n3126) );
  XOR2_X1 U3079 ( .A(n3127), .B(n3128), .Z(n3118) );
  XOR2_X1 U3080 ( .A(n3129), .B(n3130), .Z(n3128) );
  NAND2_X1 U3081 ( .A1(b_9_), .A2(a_1_), .ZN(n3130) );
  NOR2_X1 U3082 ( .A1(n3120), .A2(n3121), .ZN(n3123) );
  NOR2_X1 U3083 ( .A1(n2420), .A2(n2452), .ZN(n3121) );
  NAND2_X1 U3084 ( .A1(n3116), .A2(n3131), .ZN(n3120) );
  NAND2_X1 U3085 ( .A1(n3115), .A2(n3117), .ZN(n3131) );
  NAND2_X1 U3086 ( .A1(n3132), .A2(n3133), .ZN(n3117) );
  NAND2_X1 U3087 ( .A1(b_10_), .A2(a_1_), .ZN(n3133) );
  XNOR2_X1 U3088 ( .A(n3134), .B(n3135), .ZN(n3115) );
  XOR2_X1 U3089 ( .A(n3136), .B(n3137), .Z(n3135) );
  NAND2_X1 U3090 ( .A1(a_2_), .A2(b_9_), .ZN(n3137) );
  INV_X1 U3091 ( .A(n3138), .ZN(n3116) );
  NOR2_X1 U3092 ( .A1(n2647), .A2(n3132), .ZN(n3138) );
  NOR2_X1 U3093 ( .A1(n3139), .A2(n3140), .ZN(n3132) );
  INV_X1 U3094 ( .A(n3141), .ZN(n3140) );
  NAND3_X1 U3095 ( .A1(b_10_), .A2(n3142), .A3(a_2_), .ZN(n3141) );
  NAND2_X1 U3096 ( .A1(n3112), .A2(n3110), .ZN(n3142) );
  NOR2_X1 U3097 ( .A1(n3110), .A2(n3112), .ZN(n3139) );
  NOR2_X1 U3098 ( .A1(n3143), .A2(n3144), .ZN(n3112) );
  INV_X1 U3099 ( .A(n3145), .ZN(n3144) );
  NAND2_X1 U3100 ( .A1(n3109), .A2(n3146), .ZN(n3145) );
  NAND2_X1 U3101 ( .A1(n3108), .A2(n3107), .ZN(n3146) );
  NOR2_X1 U3102 ( .A1(n2376), .A2(n2452), .ZN(n3109) );
  NOR2_X1 U3103 ( .A1(n3107), .A2(n3108), .ZN(n3143) );
  NOR2_X1 U3104 ( .A1(n3147), .A2(n3148), .ZN(n3108) );
  NOR3_X1 U3105 ( .A1(n2452), .A2(n3149), .A3(n2457), .ZN(n3148) );
  NOR2_X1 U3106 ( .A1(n3020), .A2(n3018), .ZN(n3149) );
  INV_X1 U3107 ( .A(n3150), .ZN(n3147) );
  NAND2_X1 U3108 ( .A1(n3018), .A2(n3020), .ZN(n3150) );
  NAND2_X1 U3109 ( .A1(n3104), .A2(n3151), .ZN(n3020) );
  NAND2_X1 U3110 ( .A1(n3103), .A2(n3105), .ZN(n3151) );
  NAND2_X1 U3111 ( .A1(n3152), .A2(n3153), .ZN(n3105) );
  NAND2_X1 U3112 ( .A1(a_5_), .A2(b_10_), .ZN(n3153) );
  XOR2_X1 U3113 ( .A(n3154), .B(n3155), .Z(n3103) );
  XOR2_X1 U3114 ( .A(n3156), .B(n3157), .Z(n3154) );
  NOR2_X1 U3115 ( .A1(n2285), .A2(n2455), .ZN(n3157) );
  NAND2_X1 U3116 ( .A1(a_5_), .A2(n3158), .ZN(n3104) );
  INV_X1 U3117 ( .A(n3152), .ZN(n3158) );
  NOR2_X1 U3118 ( .A1(n3159), .A2(n3160), .ZN(n3152) );
  INV_X1 U3119 ( .A(n3161), .ZN(n3160) );
  NAND3_X1 U3120 ( .A1(b_10_), .A2(n3162), .A3(a_6_), .ZN(n3161) );
  NAND2_X1 U3121 ( .A1(n3033), .A2(n3032), .ZN(n3162) );
  NOR2_X1 U3122 ( .A1(n3032), .A2(n3033), .ZN(n3159) );
  NOR2_X1 U3123 ( .A1(n3163), .A2(n3164), .ZN(n3033) );
  NOR3_X1 U3124 ( .A1(n2452), .A2(n3165), .A3(n2312), .ZN(n3164) );
  NOR2_X1 U3125 ( .A1(n3100), .A2(n3098), .ZN(n3165) );
  INV_X1 U3126 ( .A(n3166), .ZN(n3163) );
  NAND2_X1 U3127 ( .A1(n3098), .A2(n3100), .ZN(n3166) );
  NAND2_X1 U3128 ( .A1(n3167), .A2(n3168), .ZN(n3100) );
  NAND3_X1 U3129 ( .A1(b_10_), .A2(n3169), .A3(a_8_), .ZN(n3168) );
  INV_X1 U3130 ( .A(n3170), .ZN(n3169) );
  NOR2_X1 U3131 ( .A1(n3096), .A2(n3094), .ZN(n3170) );
  NAND2_X1 U3132 ( .A1(n3094), .A2(n3096), .ZN(n3167) );
  NAND2_X1 U3133 ( .A1(n3092), .A2(n3171), .ZN(n3096) );
  NAND2_X1 U3134 ( .A1(n3091), .A2(n3093), .ZN(n3171) );
  NAND2_X1 U3135 ( .A1(n3172), .A2(n3173), .ZN(n3093) );
  NAND2_X1 U3136 ( .A1(a_9_), .A2(b_10_), .ZN(n3172) );
  XNOR2_X1 U3137 ( .A(n3174), .B(n3175), .ZN(n3091) );
  NAND2_X1 U3138 ( .A1(n3176), .A2(n3177), .ZN(n3174) );
  NAND2_X1 U3139 ( .A1(n3178), .A2(a_9_), .ZN(n3092) );
  INV_X1 U3140 ( .A(n3173), .ZN(n3178) );
  NAND2_X1 U3141 ( .A1(n3179), .A2(n3180), .ZN(n3173) );
  NAND2_X1 U3142 ( .A1(n3051), .A2(n3181), .ZN(n3180) );
  INV_X1 U3143 ( .A(n3182), .ZN(n3181) );
  NOR2_X1 U3144 ( .A1(n2273), .A2(n3053), .ZN(n3182) );
  XOR2_X1 U3145 ( .A(n3183), .B(n3184), .Z(n3051) );
  XOR2_X1 U3146 ( .A(n3185), .B(n3186), .Z(n3183) );
  NAND2_X1 U3147 ( .A1(b_9_), .A2(a_11_), .ZN(n3185) );
  NAND2_X1 U3148 ( .A1(n3053), .A2(n2273), .ZN(n3179) );
  NAND2_X1 U3149 ( .A1(b_10_), .A2(a_10_), .ZN(n2273) );
  NOR2_X1 U3150 ( .A1(n3187), .A2(n3188), .ZN(n3053) );
  INV_X1 U3151 ( .A(n3189), .ZN(n3188) );
  NAND3_X1 U3152 ( .A1(a_11_), .A2(n3190), .A3(b_10_), .ZN(n3189) );
  NAND2_X1 U3153 ( .A1(n3061), .A2(n3059), .ZN(n3190) );
  NOR2_X1 U3154 ( .A1(n3059), .A2(n3061), .ZN(n3187) );
  NOR2_X1 U3155 ( .A1(n3191), .A2(n3192), .ZN(n3061) );
  INV_X1 U3156 ( .A(n3193), .ZN(n3192) );
  NAND2_X1 U3157 ( .A1(n3069), .A2(n3194), .ZN(n3193) );
  NAND2_X1 U3158 ( .A1(n3070), .A2(n3068), .ZN(n3194) );
  NOR2_X1 U3159 ( .A1(n2452), .A2(n2238), .ZN(n3069) );
  NOR2_X1 U3160 ( .A1(n3068), .A2(n3070), .ZN(n3191) );
  NOR2_X1 U3161 ( .A1(n3195), .A2(n3196), .ZN(n3070) );
  INV_X1 U3162 ( .A(n3197), .ZN(n3196) );
  NAND2_X1 U3163 ( .A1(n3087), .A2(n3198), .ZN(n3197) );
  NAND2_X1 U3164 ( .A1(n3088), .A2(n3089), .ZN(n3198) );
  NOR2_X1 U3165 ( .A1(n2452), .A2(n2223), .ZN(n3087) );
  NOR2_X1 U3166 ( .A1(n3089), .A2(n3088), .ZN(n3195) );
  INV_X1 U3167 ( .A(n3199), .ZN(n3088) );
  NAND2_X1 U3168 ( .A1(n3200), .A2(n3201), .ZN(n3199) );
  NAND2_X1 U3169 ( .A1(b_8_), .A2(n3202), .ZN(n3201) );
  NAND2_X1 U3170 ( .A1(n2202), .A2(n3203), .ZN(n3202) );
  NAND2_X1 U3171 ( .A1(a_15_), .A2(n2285), .ZN(n3203) );
  NAND2_X1 U3172 ( .A1(b_9_), .A2(n3204), .ZN(n3200) );
  NAND2_X1 U3173 ( .A1(n2205), .A2(n3205), .ZN(n3204) );
  NAND2_X1 U3174 ( .A1(a_14_), .A2(n3206), .ZN(n3205) );
  NAND3_X1 U3175 ( .A1(b_9_), .A2(b_10_), .A3(n2450), .ZN(n3089) );
  XNOR2_X1 U3176 ( .A(n3207), .B(n3208), .ZN(n3068) );
  XOR2_X1 U3177 ( .A(n3209), .B(n3210), .Z(n3207) );
  XOR2_X1 U3178 ( .A(n3211), .B(n3212), .Z(n3059) );
  XNOR2_X1 U3179 ( .A(n3213), .B(n3214), .ZN(n3211) );
  XOR2_X1 U3180 ( .A(n3215), .B(n3216), .Z(n3094) );
  XNOR2_X1 U3181 ( .A(n3217), .B(n2280), .ZN(n3216) );
  XNOR2_X1 U3182 ( .A(n3218), .B(n3219), .ZN(n3098) );
  XOR2_X1 U3183 ( .A(n3220), .B(n3221), .Z(n3219) );
  NAND2_X1 U3184 ( .A1(a_8_), .A2(b_9_), .ZN(n3221) );
  XOR2_X1 U3185 ( .A(n3222), .B(n3223), .Z(n3032) );
  XOR2_X1 U3186 ( .A(n3224), .B(n3225), .Z(n3223) );
  NAND2_X1 U3187 ( .A1(a_7_), .A2(b_9_), .ZN(n3225) );
  XNOR2_X1 U3188 ( .A(n3226), .B(n3227), .ZN(n3018) );
  NAND2_X1 U3189 ( .A1(n3228), .A2(n3229), .ZN(n3226) );
  XOR2_X1 U3190 ( .A(n3230), .B(n3231), .Z(n3107) );
  XOR2_X1 U3191 ( .A(n3232), .B(n3233), .Z(n3230) );
  XNOR2_X1 U3192 ( .A(n3234), .B(n3235), .ZN(n3110) );
  XOR2_X1 U3193 ( .A(n3236), .B(n3237), .Z(n3235) );
  NAND2_X1 U3194 ( .A1(a_3_), .A2(b_9_), .ZN(n3237) );
  NOR2_X1 U3195 ( .A1(n2508), .A2(n3238), .ZN(n3122) );
  INV_X1 U3196 ( .A(n3239), .ZN(n3238) );
  NAND2_X1 U3197 ( .A1(n3240), .A2(n3241), .ZN(n3239) );
  XNOR2_X1 U3198 ( .A(n3242), .B(n3243), .ZN(n2153) );
  XOR2_X1 U3199 ( .A(n3244), .B(n3245), .Z(n3243) );
  NAND2_X1 U3200 ( .A1(a_0_), .A2(b_9_), .ZN(n3245) );
  NOR2_X1 U3201 ( .A1(n3241), .A2(n3240), .ZN(n2508) );
  NOR2_X1 U3202 ( .A1(n3246), .A2(n3247), .ZN(n3240) );
  NOR3_X1 U3203 ( .A1(n2285), .A2(n3248), .A3(n2420), .ZN(n3247) );
  NOR2_X1 U3204 ( .A1(n3244), .A2(n3242), .ZN(n3248) );
  INV_X1 U3205 ( .A(n3249), .ZN(n3246) );
  NAND2_X1 U3206 ( .A1(n3242), .A2(n3244), .ZN(n3249) );
  NAND2_X1 U3207 ( .A1(n3250), .A2(n3251), .ZN(n3244) );
  NAND3_X1 U3208 ( .A1(a_1_), .A2(n3252), .A3(b_9_), .ZN(n3251) );
  INV_X1 U3209 ( .A(n3253), .ZN(n3252) );
  NOR2_X1 U3210 ( .A1(n3127), .A2(n3129), .ZN(n3253) );
  NAND2_X1 U3211 ( .A1(n3127), .A2(n3129), .ZN(n3250) );
  NAND2_X1 U3212 ( .A1(n3254), .A2(n3255), .ZN(n3129) );
  INV_X1 U3213 ( .A(n3256), .ZN(n3255) );
  NOR3_X1 U3214 ( .A1(n2285), .A2(n3257), .A3(n2460), .ZN(n3256) );
  NOR2_X1 U3215 ( .A1(n3134), .A2(n3136), .ZN(n3257) );
  NAND2_X1 U3216 ( .A1(n3134), .A2(n3136), .ZN(n3254) );
  NAND2_X1 U3217 ( .A1(n3258), .A2(n3259), .ZN(n3136) );
  NAND3_X1 U3218 ( .A1(b_9_), .A2(n3260), .A3(a_3_), .ZN(n3259) );
  NAND2_X1 U3219 ( .A1(n3261), .A2(n3236), .ZN(n3260) );
  INV_X1 U3220 ( .A(n3234), .ZN(n3261) );
  NAND2_X1 U3221 ( .A1(n3234), .A2(n3262), .ZN(n3258) );
  INV_X1 U3222 ( .A(n3236), .ZN(n3262) );
  NAND2_X1 U3223 ( .A1(n3263), .A2(n3264), .ZN(n3236) );
  NAND2_X1 U3224 ( .A1(n3231), .A2(n3265), .ZN(n3264) );
  NAND2_X1 U3225 ( .A1(n3233), .A2(n3232), .ZN(n3265) );
  XNOR2_X1 U3226 ( .A(n3266), .B(n3267), .ZN(n3231) );
  XOR2_X1 U3227 ( .A(n3268), .B(n3269), .Z(n3267) );
  INV_X1 U3228 ( .A(n3270), .ZN(n3263) );
  NOR2_X1 U3229 ( .A1(n3232), .A2(n3233), .ZN(n3270) );
  NOR2_X1 U3230 ( .A1(n2457), .A2(n2285), .ZN(n3233) );
  NAND2_X1 U3231 ( .A1(n3228), .A2(n3271), .ZN(n3232) );
  NAND2_X1 U3232 ( .A1(n3227), .A2(n3229), .ZN(n3271) );
  NAND2_X1 U3233 ( .A1(n3272), .A2(n3273), .ZN(n3229) );
  NAND2_X1 U3234 ( .A1(a_5_), .A2(b_9_), .ZN(n3273) );
  XOR2_X1 U3235 ( .A(n3274), .B(n3275), .Z(n3227) );
  XOR2_X1 U3236 ( .A(n3276), .B(n3277), .Z(n3274) );
  NOR2_X1 U3237 ( .A1(n3206), .A2(n2455), .ZN(n3277) );
  NAND2_X1 U3238 ( .A1(a_5_), .A2(n3278), .ZN(n3228) );
  INV_X1 U3239 ( .A(n3272), .ZN(n3278) );
  NOR2_X1 U3240 ( .A1(n3279), .A2(n3280), .ZN(n3272) );
  NOR3_X1 U3241 ( .A1(n2285), .A2(n3281), .A3(n2455), .ZN(n3280) );
  NOR2_X1 U3242 ( .A1(n3155), .A2(n3156), .ZN(n3281) );
  INV_X1 U3243 ( .A(n3282), .ZN(n3279) );
  NAND2_X1 U3244 ( .A1(n3155), .A2(n3156), .ZN(n3282) );
  NAND2_X1 U3245 ( .A1(n3283), .A2(n3284), .ZN(n3156) );
  INV_X1 U3246 ( .A(n3285), .ZN(n3284) );
  NOR3_X1 U3247 ( .A1(n2285), .A2(n3286), .A3(n2312), .ZN(n3285) );
  NOR2_X1 U3248 ( .A1(n3222), .A2(n3224), .ZN(n3286) );
  NAND2_X1 U3249 ( .A1(n3222), .A2(n3224), .ZN(n3283) );
  NAND2_X1 U3250 ( .A1(n3287), .A2(n3288), .ZN(n3224) );
  NAND3_X1 U3251 ( .A1(b_9_), .A2(n3289), .A3(a_8_), .ZN(n3288) );
  NAND2_X1 U3252 ( .A1(n3218), .A2(n3220), .ZN(n3289) );
  INV_X1 U3253 ( .A(n3290), .ZN(n3287) );
  NOR2_X1 U3254 ( .A1(n3218), .A2(n3220), .ZN(n3290) );
  NAND2_X1 U3255 ( .A1(n3291), .A2(n3292), .ZN(n3220) );
  NAND2_X1 U3256 ( .A1(n3215), .A2(n3293), .ZN(n3292) );
  NAND2_X1 U3257 ( .A1(n2280), .A2(n3217), .ZN(n3293) );
  XOR2_X1 U3258 ( .A(n3294), .B(n3295), .Z(n3215) );
  NAND2_X1 U3259 ( .A1(n3296), .A2(n3297), .ZN(n3294) );
  INV_X1 U3260 ( .A(n3298), .ZN(n3291) );
  NOR2_X1 U3261 ( .A1(n3217), .A2(n2280), .ZN(n3298) );
  NOR2_X1 U3262 ( .A1(n2283), .A2(n2285), .ZN(n2280) );
  NAND2_X1 U3263 ( .A1(n3176), .A2(n3299), .ZN(n3217) );
  NAND2_X1 U3264 ( .A1(n3175), .A2(n3177), .ZN(n3299) );
  NAND2_X1 U3265 ( .A1(n3300), .A2(n3301), .ZN(n3177) );
  NAND2_X1 U3266 ( .A1(b_9_), .A2(a_10_), .ZN(n3301) );
  XNOR2_X1 U3267 ( .A(n3302), .B(n3303), .ZN(n3175) );
  XOR2_X1 U3268 ( .A(n3304), .B(n3305), .Z(n3302) );
  NAND2_X1 U3269 ( .A1(b_8_), .A2(a_11_), .ZN(n3304) );
  INV_X1 U3270 ( .A(n3306), .ZN(n3176) );
  NOR2_X1 U3271 ( .A1(n2453), .A2(n3300), .ZN(n3306) );
  NOR2_X1 U3272 ( .A1(n3307), .A2(n3308), .ZN(n3300) );
  INV_X1 U3273 ( .A(n3309), .ZN(n3308) );
  NAND3_X1 U3274 ( .A1(a_11_), .A2(n3310), .A3(b_9_), .ZN(n3309) );
  NAND2_X1 U3275 ( .A1(n3184), .A2(n3186), .ZN(n3310) );
  NOR2_X1 U3276 ( .A1(n3184), .A2(n3186), .ZN(n3307) );
  NOR2_X1 U3277 ( .A1(n3311), .A2(n3312), .ZN(n3186) );
  INV_X1 U3278 ( .A(n3313), .ZN(n3312) );
  NAND2_X1 U3279 ( .A1(n3213), .A2(n3314), .ZN(n3313) );
  NAND2_X1 U3280 ( .A1(n3214), .A2(n3212), .ZN(n3314) );
  NOR2_X1 U3281 ( .A1(n2285), .A2(n2238), .ZN(n3213) );
  NOR2_X1 U3282 ( .A1(n3212), .A2(n3214), .ZN(n3311) );
  NOR2_X1 U3283 ( .A1(n3315), .A2(n3316), .ZN(n3214) );
  INV_X1 U3284 ( .A(n3317), .ZN(n3316) );
  NAND2_X1 U3285 ( .A1(n3208), .A2(n3318), .ZN(n3317) );
  NAND2_X1 U3286 ( .A1(n3209), .A2(n3210), .ZN(n3318) );
  NOR2_X1 U3287 ( .A1(n2285), .A2(n2223), .ZN(n3208) );
  NOR2_X1 U3288 ( .A1(n3210), .A2(n3209), .ZN(n3315) );
  INV_X1 U3289 ( .A(n3319), .ZN(n3209) );
  NAND2_X1 U3290 ( .A1(n3320), .A2(n3321), .ZN(n3319) );
  NAND2_X1 U3291 ( .A1(b_7_), .A2(n3322), .ZN(n3321) );
  NAND2_X1 U3292 ( .A1(n2202), .A2(n3323), .ZN(n3322) );
  NAND2_X1 U3293 ( .A1(a_15_), .A2(n3206), .ZN(n3323) );
  NAND2_X1 U3294 ( .A1(b_8_), .A2(n3324), .ZN(n3320) );
  NAND2_X1 U3295 ( .A1(n2205), .A2(n3325), .ZN(n3324) );
  NAND2_X1 U3296 ( .A1(a_14_), .A2(n2314), .ZN(n3325) );
  NAND3_X1 U3297 ( .A1(b_8_), .A2(b_9_), .A3(n2450), .ZN(n3210) );
  XNOR2_X1 U3298 ( .A(n3326), .B(n3327), .ZN(n3212) );
  XOR2_X1 U3299 ( .A(n3328), .B(n3329), .Z(n3326) );
  XOR2_X1 U3300 ( .A(n3330), .B(n3331), .Z(n3184) );
  XNOR2_X1 U3301 ( .A(n3332), .B(n3333), .ZN(n3330) );
  XOR2_X1 U3302 ( .A(n3334), .B(n3335), .Z(n3218) );
  NAND2_X1 U3303 ( .A1(n3336), .A2(n3337), .ZN(n3334) );
  XOR2_X1 U3304 ( .A(n3338), .B(n3339), .Z(n3222) );
  XNOR2_X1 U3305 ( .A(n3340), .B(n2302), .ZN(n3339) );
  XNOR2_X1 U3306 ( .A(n3341), .B(n3342), .ZN(n3155) );
  XOR2_X1 U3307 ( .A(n3343), .B(n3344), .Z(n3342) );
  NAND2_X1 U3308 ( .A1(a_7_), .A2(b_8_), .ZN(n3344) );
  XOR2_X1 U3309 ( .A(n3345), .B(n3346), .Z(n3234) );
  XNOR2_X1 U3310 ( .A(n3347), .B(n3348), .ZN(n3345) );
  NAND2_X1 U3311 ( .A1(a_4_), .A2(b_8_), .ZN(n3347) );
  XNOR2_X1 U3312 ( .A(n3349), .B(n3350), .ZN(n3134) );
  NAND2_X1 U3313 ( .A1(n3351), .A2(n3352), .ZN(n3349) );
  XNOR2_X1 U3314 ( .A(n3353), .B(n3354), .ZN(n3127) );
  NAND2_X1 U3315 ( .A1(n3355), .A2(n3356), .ZN(n3353) );
  XNOR2_X1 U3316 ( .A(n3357), .B(n3358), .ZN(n3242) );
  NAND2_X1 U3317 ( .A1(n3359), .A2(n3360), .ZN(n3357) );
  XOR2_X1 U3318 ( .A(n3361), .B(n3362), .Z(n3241) );
  XNOR2_X1 U3319 ( .A(n3363), .B(n3364), .ZN(n3362) );
  XNOR2_X1 U3320 ( .A(n2165), .B(n2164), .ZN(n2156) );
  NAND3_X1 U3321 ( .A1(n2164), .A2(n2165), .A3(n3365), .ZN(n2161) );
  INV_X1 U3322 ( .A(n2162), .ZN(n3365) );
  NAND2_X1 U3323 ( .A1(n2505), .A2(n3366), .ZN(n2162) );
  INV_X1 U3324 ( .A(n3367), .ZN(n3366) );
  NOR2_X1 U3325 ( .A1(n3368), .A2(n3369), .ZN(n3367) );
  NAND2_X1 U3326 ( .A1(n3370), .A2(n3371), .ZN(n2165) );
  NAND2_X1 U3327 ( .A1(n3364), .A2(n3372), .ZN(n3371) );
  INV_X1 U3328 ( .A(n3373), .ZN(n3372) );
  NOR2_X1 U3329 ( .A1(n3363), .A2(n3361), .ZN(n3373) );
  NOR2_X1 U3330 ( .A1(n2420), .A2(n3206), .ZN(n3364) );
  NAND2_X1 U3331 ( .A1(n3361), .A2(n3363), .ZN(n3370) );
  NAND2_X1 U3332 ( .A1(n3359), .A2(n3374), .ZN(n3363) );
  NAND2_X1 U3333 ( .A1(n3358), .A2(n3360), .ZN(n3374) );
  NAND2_X1 U3334 ( .A1(n3375), .A2(n3376), .ZN(n3360) );
  NAND2_X1 U3335 ( .A1(b_8_), .A2(a_1_), .ZN(n3376) );
  INV_X1 U3336 ( .A(n3377), .ZN(n3375) );
  XOR2_X1 U3337 ( .A(n3378), .B(n3379), .Z(n3358) );
  XNOR2_X1 U3338 ( .A(n3380), .B(n3381), .ZN(n3379) );
  NAND2_X1 U3339 ( .A1(a_2_), .A2(b_7_), .ZN(n3381) );
  NAND2_X1 U3340 ( .A1(a_1_), .A2(n3377), .ZN(n3359) );
  NAND2_X1 U3341 ( .A1(n3355), .A2(n3382), .ZN(n3377) );
  NAND2_X1 U3342 ( .A1(n3354), .A2(n3356), .ZN(n3382) );
  NAND2_X1 U3343 ( .A1(n3383), .A2(n3384), .ZN(n3356) );
  NAND2_X1 U3344 ( .A1(a_2_), .A2(b_8_), .ZN(n3384) );
  INV_X1 U3345 ( .A(n3385), .ZN(n3383) );
  XNOR2_X1 U3346 ( .A(n3386), .B(n3387), .ZN(n3354) );
  XNOR2_X1 U3347 ( .A(n3388), .B(n3389), .ZN(n3386) );
  NOR2_X1 U3348 ( .A1(n2314), .A2(n2376), .ZN(n3389) );
  NAND2_X1 U3349 ( .A1(a_2_), .A2(n3385), .ZN(n3355) );
  NAND2_X1 U3350 ( .A1(n3351), .A2(n3390), .ZN(n3385) );
  NAND2_X1 U3351 ( .A1(n3350), .A2(n3352), .ZN(n3390) );
  NAND2_X1 U3352 ( .A1(n3391), .A2(n3392), .ZN(n3352) );
  NAND2_X1 U3353 ( .A1(a_3_), .A2(b_8_), .ZN(n3392) );
  XNOR2_X1 U3354 ( .A(n3393), .B(n3394), .ZN(n3350) );
  XOR2_X1 U3355 ( .A(n3395), .B(n3396), .Z(n3394) );
  NAND2_X1 U3356 ( .A1(a_4_), .A2(b_7_), .ZN(n3396) );
  NAND2_X1 U3357 ( .A1(a_3_), .A2(n3397), .ZN(n3351) );
  INV_X1 U3358 ( .A(n3391), .ZN(n3397) );
  NOR2_X1 U3359 ( .A1(n3398), .A2(n3399), .ZN(n3391) );
  NOR3_X1 U3360 ( .A1(n3206), .A2(n3400), .A3(n2457), .ZN(n3399) );
  NOR2_X1 U3361 ( .A1(n3346), .A2(n3348), .ZN(n3400) );
  INV_X1 U3362 ( .A(n3401), .ZN(n3398) );
  NAND2_X1 U3363 ( .A1(n3346), .A2(n3348), .ZN(n3401) );
  NAND2_X1 U3364 ( .A1(n3402), .A2(n3403), .ZN(n3348) );
  NAND2_X1 U3365 ( .A1(n3269), .A2(n3404), .ZN(n3403) );
  NAND2_X1 U3366 ( .A1(n3266), .A2(n3268), .ZN(n3404) );
  NOR2_X1 U3367 ( .A1(n2341), .A2(n3206), .ZN(n3269) );
  INV_X1 U3368 ( .A(n3405), .ZN(n3402) );
  NOR2_X1 U3369 ( .A1(n3266), .A2(n3268), .ZN(n3405) );
  NOR2_X1 U3370 ( .A1(n3406), .A2(n3407), .ZN(n3268) );
  NOR3_X1 U3371 ( .A1(n3206), .A2(n3408), .A3(n2455), .ZN(n3407) );
  NOR2_X1 U3372 ( .A1(n3276), .A2(n3275), .ZN(n3408) );
  INV_X1 U3373 ( .A(n3409), .ZN(n3406) );
  NAND2_X1 U3374 ( .A1(n3275), .A2(n3276), .ZN(n3409) );
  NAND2_X1 U3375 ( .A1(n3410), .A2(n3411), .ZN(n3276) );
  NAND3_X1 U3376 ( .A1(b_8_), .A2(n3412), .A3(a_7_), .ZN(n3411) );
  NAND2_X1 U3377 ( .A1(n3341), .A2(n3343), .ZN(n3412) );
  NAND2_X1 U3378 ( .A1(n3413), .A2(n3414), .ZN(n3410) );
  INV_X1 U3379 ( .A(n3341), .ZN(n3414) );
  XOR2_X1 U3380 ( .A(n3415), .B(n3416), .Z(n3341) );
  XOR2_X1 U3381 ( .A(n3417), .B(n3418), .Z(n3416) );
  INV_X1 U3382 ( .A(n3343), .ZN(n3413) );
  NAND2_X1 U3383 ( .A1(n3419), .A2(n3420), .ZN(n3343) );
  NAND2_X1 U3384 ( .A1(n3338), .A2(n3421), .ZN(n3420) );
  NAND2_X1 U3385 ( .A1(n2302), .A2(n3340), .ZN(n3421) );
  XOR2_X1 U3386 ( .A(n3422), .B(n3423), .Z(n3338) );
  NAND2_X1 U3387 ( .A1(n3424), .A2(n3425), .ZN(n3422) );
  INV_X1 U3388 ( .A(n3426), .ZN(n3419) );
  NOR2_X1 U3389 ( .A1(n3340), .A2(n2302), .ZN(n3426) );
  NOR2_X1 U3390 ( .A1(n3206), .A2(n2681), .ZN(n2302) );
  NAND2_X1 U3391 ( .A1(n3336), .A2(n3427), .ZN(n3340) );
  NAND2_X1 U3392 ( .A1(n3335), .A2(n3337), .ZN(n3427) );
  NAND2_X1 U3393 ( .A1(n3428), .A2(n3429), .ZN(n3337) );
  NAND2_X1 U3394 ( .A1(b_8_), .A2(a_9_), .ZN(n3429) );
  INV_X1 U3395 ( .A(n3430), .ZN(n3428) );
  XNOR2_X1 U3396 ( .A(n3431), .B(n3432), .ZN(n3335) );
  NAND2_X1 U3397 ( .A1(n3433), .A2(n3434), .ZN(n3431) );
  NAND2_X1 U3398 ( .A1(a_9_), .A2(n3430), .ZN(n3336) );
  NAND2_X1 U3399 ( .A1(n3296), .A2(n3435), .ZN(n3430) );
  NAND2_X1 U3400 ( .A1(n3295), .A2(n3297), .ZN(n3435) );
  NAND2_X1 U3401 ( .A1(n3436), .A2(n3437), .ZN(n3297) );
  NAND2_X1 U3402 ( .A1(b_8_), .A2(a_10_), .ZN(n3437) );
  XNOR2_X1 U3403 ( .A(n3438), .B(n3439), .ZN(n3295) );
  XOR2_X1 U3404 ( .A(n3440), .B(n3441), .Z(n3438) );
  NAND2_X1 U3405 ( .A1(b_7_), .A2(a_11_), .ZN(n3440) );
  INV_X1 U3406 ( .A(n3442), .ZN(n3296) );
  NOR2_X1 U3407 ( .A1(n2453), .A2(n3436), .ZN(n3442) );
  NOR2_X1 U3408 ( .A1(n3443), .A2(n3444), .ZN(n3436) );
  INV_X1 U3409 ( .A(n3445), .ZN(n3444) );
  NAND3_X1 U3410 ( .A1(a_11_), .A2(n3446), .A3(b_8_), .ZN(n3445) );
  NAND2_X1 U3411 ( .A1(n3303), .A2(n3305), .ZN(n3446) );
  NOR2_X1 U3412 ( .A1(n3303), .A2(n3305), .ZN(n3443) );
  NOR2_X1 U3413 ( .A1(n3447), .A2(n3448), .ZN(n3305) );
  INV_X1 U3414 ( .A(n3449), .ZN(n3448) );
  NAND2_X1 U3415 ( .A1(n3332), .A2(n3450), .ZN(n3449) );
  NAND2_X1 U3416 ( .A1(n3333), .A2(n3331), .ZN(n3450) );
  NOR2_X1 U3417 ( .A1(n3206), .A2(n2238), .ZN(n3332) );
  NOR2_X1 U3418 ( .A1(n3331), .A2(n3333), .ZN(n3447) );
  NOR2_X1 U3419 ( .A1(n3451), .A2(n3452), .ZN(n3333) );
  INV_X1 U3420 ( .A(n3453), .ZN(n3452) );
  NAND2_X1 U3421 ( .A1(n3327), .A2(n3454), .ZN(n3453) );
  NAND2_X1 U3422 ( .A1(n3328), .A2(n3329), .ZN(n3454) );
  NOR2_X1 U3423 ( .A1(n3206), .A2(n2223), .ZN(n3327) );
  NOR2_X1 U3424 ( .A1(n3329), .A2(n3328), .ZN(n3451) );
  INV_X1 U3425 ( .A(n3455), .ZN(n3328) );
  NAND2_X1 U3426 ( .A1(n3456), .A2(n3457), .ZN(n3455) );
  NAND2_X1 U3427 ( .A1(b_6_), .A2(n3458), .ZN(n3457) );
  NAND2_X1 U3428 ( .A1(n2202), .A2(n3459), .ZN(n3458) );
  NAND2_X1 U3429 ( .A1(a_15_), .A2(n2314), .ZN(n3459) );
  NAND2_X1 U3430 ( .A1(b_7_), .A2(n3460), .ZN(n3456) );
  NAND2_X1 U3431 ( .A1(n2205), .A2(n3461), .ZN(n3460) );
  NAND2_X1 U3432 ( .A1(a_14_), .A2(n2454), .ZN(n3461) );
  NAND3_X1 U3433 ( .A1(b_8_), .A2(b_7_), .A3(n2450), .ZN(n3329) );
  XNOR2_X1 U3434 ( .A(n3462), .B(n3463), .ZN(n3331) );
  XOR2_X1 U3435 ( .A(n3464), .B(n3465), .Z(n3462) );
  XOR2_X1 U3436 ( .A(n3466), .B(n3467), .Z(n3303) );
  XNOR2_X1 U3437 ( .A(n3468), .B(n3469), .ZN(n3466) );
  XNOR2_X1 U3438 ( .A(n3470), .B(n3471), .ZN(n3275) );
  XNOR2_X1 U3439 ( .A(n3472), .B(n2433), .ZN(n3470) );
  XNOR2_X1 U3440 ( .A(n3473), .B(n3474), .ZN(n3266) );
  NOR2_X1 U3441 ( .A1(n3475), .A2(n3476), .ZN(n3474) );
  NOR2_X1 U3442 ( .A1(n3477), .A2(n3478), .ZN(n3475) );
  NOR2_X1 U3443 ( .A1(n2314), .A2(n2455), .ZN(n3478) );
  INV_X1 U3444 ( .A(n3479), .ZN(n3477) );
  XNOR2_X1 U3445 ( .A(n3480), .B(n3481), .ZN(n3346) );
  XOR2_X1 U3446 ( .A(n3482), .B(n3483), .Z(n3481) );
  NAND2_X1 U3447 ( .A1(a_5_), .A2(b_7_), .ZN(n3483) );
  XNOR2_X1 U3448 ( .A(n3484), .B(n3485), .ZN(n3361) );
  XNOR2_X1 U3449 ( .A(n3486), .B(n3487), .ZN(n3484) );
  NOR2_X1 U3450 ( .A1(n2647), .A2(n2314), .ZN(n3487) );
  XNOR2_X1 U3451 ( .A(n3488), .B(n3489), .ZN(n2164) );
  XOR2_X1 U3452 ( .A(n3490), .B(n3491), .Z(n3489) );
  NAND2_X1 U3453 ( .A1(a_0_), .A2(b_7_), .ZN(n3491) );
  NAND2_X1 U3454 ( .A1(n3369), .A2(n3368), .ZN(n2505) );
  NAND2_X1 U3455 ( .A1(n3492), .A2(n3493), .ZN(n3368) );
  INV_X1 U3456 ( .A(n3494), .ZN(n3493) );
  NOR3_X1 U3457 ( .A1(n2314), .A2(n3495), .A3(n2420), .ZN(n3494) );
  NOR2_X1 U3458 ( .A1(n3490), .A2(n3488), .ZN(n3495) );
  NAND2_X1 U3459 ( .A1(n3488), .A2(n3490), .ZN(n3492) );
  NAND2_X1 U3460 ( .A1(n3496), .A2(n3497), .ZN(n3490) );
  NAND3_X1 U3461 ( .A1(a_1_), .A2(n3498), .A3(b_7_), .ZN(n3497) );
  NAND2_X1 U3462 ( .A1(n3485), .A2(n3486), .ZN(n3498) );
  INV_X1 U3463 ( .A(n3499), .ZN(n3496) );
  NOR2_X1 U3464 ( .A1(n3485), .A2(n3486), .ZN(n3499) );
  NOR2_X1 U3465 ( .A1(n3500), .A2(n3501), .ZN(n3486) );
  INV_X1 U3466 ( .A(n3502), .ZN(n3501) );
  NAND3_X1 U3467 ( .A1(b_7_), .A2(n3503), .A3(a_2_), .ZN(n3502) );
  NAND2_X1 U3468 ( .A1(n3380), .A2(n3378), .ZN(n3503) );
  NOR2_X1 U3469 ( .A1(n3378), .A2(n3380), .ZN(n3500) );
  NOR2_X1 U3470 ( .A1(n3504), .A2(n3505), .ZN(n3380) );
  NOR3_X1 U3471 ( .A1(n2314), .A2(n3506), .A3(n2376), .ZN(n3505) );
  INV_X1 U3472 ( .A(n3507), .ZN(n3506) );
  NAND2_X1 U3473 ( .A1(n3388), .A2(n3387), .ZN(n3507) );
  NOR2_X1 U3474 ( .A1(n3387), .A2(n3388), .ZN(n3504) );
  NOR2_X1 U3475 ( .A1(n3508), .A2(n3509), .ZN(n3388) );
  NOR3_X1 U3476 ( .A1(n2314), .A2(n3510), .A3(n2457), .ZN(n3509) );
  NOR2_X1 U3477 ( .A1(n3395), .A2(n3393), .ZN(n3510) );
  INV_X1 U3478 ( .A(n3511), .ZN(n3508) );
  NAND2_X1 U3479 ( .A1(n3393), .A2(n3395), .ZN(n3511) );
  NAND2_X1 U3480 ( .A1(n3512), .A2(n3513), .ZN(n3395) );
  NAND3_X1 U3481 ( .A1(b_7_), .A2(n3514), .A3(a_5_), .ZN(n3513) );
  INV_X1 U3482 ( .A(n3515), .ZN(n3514) );
  NOR2_X1 U3483 ( .A1(n3482), .A2(n3480), .ZN(n3515) );
  NAND2_X1 U3484 ( .A1(n3480), .A2(n3482), .ZN(n3512) );
  NAND2_X1 U3485 ( .A1(n3516), .A2(n3517), .ZN(n3482) );
  NAND2_X1 U3486 ( .A1(n3473), .A2(n3518), .ZN(n3517) );
  NAND2_X1 U3487 ( .A1(n3479), .A2(n3519), .ZN(n3518) );
  NAND2_X1 U3488 ( .A1(a_6_), .A2(b_7_), .ZN(n3519) );
  XNOR2_X1 U3489 ( .A(n3520), .B(n3521), .ZN(n3473) );
  XNOR2_X1 U3490 ( .A(n3522), .B(n3523), .ZN(n3521) );
  INV_X1 U3491 ( .A(n3476), .ZN(n3516) );
  NOR2_X1 U3492 ( .A1(n3479), .A2(n2455), .ZN(n3476) );
  NAND2_X1 U3493 ( .A1(n3524), .A2(n3525), .ZN(n3479) );
  NAND2_X1 U3494 ( .A1(n3471), .A2(n3526), .ZN(n3525) );
  NAND2_X1 U3495 ( .A1(n2309), .A2(n3472), .ZN(n3526) );
  XOR2_X1 U3496 ( .A(n3527), .B(n3528), .Z(n3471) );
  XOR2_X1 U3497 ( .A(n3529), .B(n3530), .Z(n3528) );
  NAND2_X1 U3498 ( .A1(b_6_), .A2(a_8_), .ZN(n3530) );
  NAND2_X1 U3499 ( .A1(n3531), .A2(n2433), .ZN(n3524) );
  INV_X1 U3500 ( .A(n2309), .ZN(n2433) );
  NOR2_X1 U3501 ( .A1(n2312), .A2(n2314), .ZN(n2309) );
  INV_X1 U3502 ( .A(n3472), .ZN(n3531) );
  NAND2_X1 U3503 ( .A1(n3532), .A2(n3533), .ZN(n3472) );
  INV_X1 U3504 ( .A(n3534), .ZN(n3533) );
  NOR2_X1 U3505 ( .A1(n3418), .A2(n3535), .ZN(n3534) );
  NOR2_X1 U3506 ( .A1(n3417), .A2(n3415), .ZN(n3535) );
  NAND2_X1 U3507 ( .A1(b_7_), .A2(a_8_), .ZN(n3418) );
  NAND2_X1 U3508 ( .A1(n3415), .A2(n3417), .ZN(n3532) );
  NAND2_X1 U3509 ( .A1(n3424), .A2(n3536), .ZN(n3417) );
  NAND2_X1 U3510 ( .A1(n3423), .A2(n3425), .ZN(n3536) );
  NAND2_X1 U3511 ( .A1(n3537), .A2(n3538), .ZN(n3425) );
  NAND2_X1 U3512 ( .A1(b_7_), .A2(a_9_), .ZN(n3538) );
  INV_X1 U3513 ( .A(n3539), .ZN(n3537) );
  XNOR2_X1 U3514 ( .A(n3540), .B(n3541), .ZN(n3423) );
  NAND2_X1 U3515 ( .A1(n3542), .A2(n3543), .ZN(n3540) );
  NAND2_X1 U3516 ( .A1(a_9_), .A2(n3539), .ZN(n3424) );
  NAND2_X1 U3517 ( .A1(n3433), .A2(n3544), .ZN(n3539) );
  NAND2_X1 U3518 ( .A1(n3432), .A2(n3434), .ZN(n3544) );
  NAND2_X1 U3519 ( .A1(n3545), .A2(n3546), .ZN(n3434) );
  NAND2_X1 U3520 ( .A1(b_7_), .A2(a_10_), .ZN(n3546) );
  XNOR2_X1 U3521 ( .A(n3547), .B(n3548), .ZN(n3432) );
  XOR2_X1 U3522 ( .A(n3549), .B(n3550), .Z(n3547) );
  NAND2_X1 U3523 ( .A1(b_6_), .A2(a_11_), .ZN(n3549) );
  INV_X1 U3524 ( .A(n3551), .ZN(n3433) );
  NOR2_X1 U3525 ( .A1(n2453), .A2(n3545), .ZN(n3551) );
  NOR2_X1 U3526 ( .A1(n3552), .A2(n3553), .ZN(n3545) );
  INV_X1 U3527 ( .A(n3554), .ZN(n3553) );
  NAND3_X1 U3528 ( .A1(a_11_), .A2(n3555), .A3(b_7_), .ZN(n3554) );
  NAND2_X1 U3529 ( .A1(n3439), .A2(n3441), .ZN(n3555) );
  NOR2_X1 U3530 ( .A1(n3439), .A2(n3441), .ZN(n3552) );
  NOR2_X1 U3531 ( .A1(n3556), .A2(n3557), .ZN(n3441) );
  INV_X1 U3532 ( .A(n3558), .ZN(n3557) );
  NAND2_X1 U3533 ( .A1(n3468), .A2(n3559), .ZN(n3558) );
  NAND2_X1 U3534 ( .A1(n3469), .A2(n3467), .ZN(n3559) );
  NOR2_X1 U3535 ( .A1(n2314), .A2(n2238), .ZN(n3468) );
  NOR2_X1 U3536 ( .A1(n3467), .A2(n3469), .ZN(n3556) );
  NOR2_X1 U3537 ( .A1(n3560), .A2(n3561), .ZN(n3469) );
  INV_X1 U3538 ( .A(n3562), .ZN(n3561) );
  NAND2_X1 U3539 ( .A1(n3463), .A2(n3563), .ZN(n3562) );
  NAND2_X1 U3540 ( .A1(n3464), .A2(n3465), .ZN(n3563) );
  NOR2_X1 U3541 ( .A1(n2314), .A2(n2223), .ZN(n3463) );
  NOR2_X1 U3542 ( .A1(n3465), .A2(n3464), .ZN(n3560) );
  INV_X1 U3543 ( .A(n3564), .ZN(n3464) );
  NAND2_X1 U3544 ( .A1(n3565), .A2(n3566), .ZN(n3564) );
  NAND2_X1 U3545 ( .A1(b_5_), .A2(n3567), .ZN(n3566) );
  NAND2_X1 U3546 ( .A1(n2202), .A2(n3568), .ZN(n3567) );
  NAND2_X1 U3547 ( .A1(a_15_), .A2(n2454), .ZN(n3568) );
  NAND2_X1 U3548 ( .A1(b_6_), .A2(n3569), .ZN(n3565) );
  NAND2_X1 U3549 ( .A1(n2205), .A2(n3570), .ZN(n3569) );
  NAND2_X1 U3550 ( .A1(a_14_), .A2(n2343), .ZN(n3570) );
  NAND3_X1 U3551 ( .A1(b_6_), .A2(b_7_), .A3(n2450), .ZN(n3465) );
  XNOR2_X1 U3552 ( .A(n3571), .B(n3572), .ZN(n3467) );
  XOR2_X1 U3553 ( .A(n3573), .B(n3574), .Z(n3571) );
  XOR2_X1 U3554 ( .A(n3575), .B(n3576), .Z(n3439) );
  XNOR2_X1 U3555 ( .A(n3577), .B(n3578), .ZN(n3575) );
  XNOR2_X1 U3556 ( .A(n3579), .B(n3580), .ZN(n3415) );
  NAND2_X1 U3557 ( .A1(n3581), .A2(n3582), .ZN(n3579) );
  XNOR2_X1 U3558 ( .A(n3583), .B(n3584), .ZN(n3480) );
  XOR2_X1 U3559 ( .A(n3585), .B(n3586), .Z(n3583) );
  XOR2_X1 U3560 ( .A(n3587), .B(n3588), .Z(n3393) );
  XOR2_X1 U3561 ( .A(n3589), .B(n3590), .Z(n3587) );
  XOR2_X1 U3562 ( .A(n3591), .B(n3592), .Z(n3387) );
  XNOR2_X1 U3563 ( .A(n3593), .B(n3594), .ZN(n3591) );
  XOR2_X1 U3564 ( .A(n3595), .B(n3596), .Z(n3378) );
  XNOR2_X1 U3565 ( .A(n3597), .B(n3598), .ZN(n3596) );
  XNOR2_X1 U3566 ( .A(n3599), .B(n3600), .ZN(n3485) );
  XOR2_X1 U3567 ( .A(n3601), .B(n3602), .Z(n3599) );
  XOR2_X1 U3568 ( .A(n3603), .B(n3604), .Z(n3488) );
  XOR2_X1 U3569 ( .A(n3605), .B(n3606), .Z(n3603) );
  XOR2_X1 U3570 ( .A(n3607), .B(n3608), .Z(n3369) );
  XOR2_X1 U3571 ( .A(n3609), .B(n3610), .Z(n3607) );
  XOR2_X1 U3572 ( .A(n2176), .B(n2177), .Z(n2168) );
  INV_X1 U3573 ( .A(n2172), .ZN(n2502) );
  NOR3_X1 U3574 ( .A1(n2177), .A2(n2176), .A3(n2504), .ZN(n2172) );
  NAND2_X1 U3575 ( .A1(n2501), .A2(n3611), .ZN(n2504) );
  NAND2_X1 U3576 ( .A1(n3612), .A2(n3613), .ZN(n3611) );
  INV_X1 U3577 ( .A(n3614), .ZN(n2176) );
  NAND2_X1 U3578 ( .A1(n3615), .A2(n3616), .ZN(n3614) );
  NAND2_X1 U3579 ( .A1(n3610), .A2(n3617), .ZN(n3616) );
  INV_X1 U3580 ( .A(n3618), .ZN(n3617) );
  NOR2_X1 U3581 ( .A1(n3609), .A2(n3608), .ZN(n3618) );
  NOR2_X1 U3582 ( .A1(n2420), .A2(n2454), .ZN(n3610) );
  NAND2_X1 U3583 ( .A1(n3608), .A2(n3609), .ZN(n3615) );
  NAND2_X1 U3584 ( .A1(n3619), .A2(n3620), .ZN(n3609) );
  NAND2_X1 U3585 ( .A1(n3606), .A2(n3621), .ZN(n3620) );
  INV_X1 U3586 ( .A(n3622), .ZN(n3621) );
  NOR2_X1 U3587 ( .A1(n3604), .A2(n3605), .ZN(n3622) );
  NOR2_X1 U3588 ( .A1(n2454), .A2(n2647), .ZN(n3606) );
  NAND2_X1 U3589 ( .A1(n3604), .A2(n3605), .ZN(n3619) );
  NAND2_X1 U3590 ( .A1(n3623), .A2(n3624), .ZN(n3605) );
  NAND2_X1 U3591 ( .A1(n3601), .A2(n3625), .ZN(n3624) );
  INV_X1 U3592 ( .A(n3626), .ZN(n3625) );
  NOR2_X1 U3593 ( .A1(n3602), .A2(n3600), .ZN(n3626) );
  NOR2_X1 U3594 ( .A1(n2460), .A2(n2454), .ZN(n3601) );
  NAND2_X1 U3595 ( .A1(n3600), .A2(n3602), .ZN(n3623) );
  NAND2_X1 U3596 ( .A1(n3627), .A2(n3628), .ZN(n3602) );
  NAND2_X1 U3597 ( .A1(n3598), .A2(n3629), .ZN(n3628) );
  INV_X1 U3598 ( .A(n3630), .ZN(n3629) );
  NOR2_X1 U3599 ( .A1(n3595), .A2(n3597), .ZN(n3630) );
  NOR2_X1 U3600 ( .A1(n2376), .A2(n2454), .ZN(n3598) );
  NAND2_X1 U3601 ( .A1(n3595), .A2(n3597), .ZN(n3627) );
  NAND2_X1 U3602 ( .A1(n3631), .A2(n3632), .ZN(n3597) );
  NAND2_X1 U3603 ( .A1(n3594), .A2(n3633), .ZN(n3632) );
  NAND2_X1 U3604 ( .A1(n3592), .A2(n3593), .ZN(n3633) );
  NOR2_X1 U3605 ( .A1(n2457), .A2(n2454), .ZN(n3594) );
  INV_X1 U3606 ( .A(n3634), .ZN(n3631) );
  NOR2_X1 U3607 ( .A1(n3592), .A2(n3593), .ZN(n3634) );
  NOR2_X1 U3608 ( .A1(n3635), .A2(n3636), .ZN(n3593) );
  INV_X1 U3609 ( .A(n3637), .ZN(n3636) );
  NAND2_X1 U3610 ( .A1(n3590), .A2(n3638), .ZN(n3637) );
  NAND2_X1 U3611 ( .A1(n3588), .A2(n3589), .ZN(n3638) );
  NOR2_X1 U3612 ( .A1(n2341), .A2(n2454), .ZN(n3590) );
  NOR2_X1 U3613 ( .A1(n3588), .A2(n3589), .ZN(n3635) );
  NAND2_X1 U3614 ( .A1(n3639), .A2(n3640), .ZN(n3589) );
  NAND2_X1 U3615 ( .A1(n3584), .A2(n3641), .ZN(n3640) );
  NAND2_X1 U3616 ( .A1(n3586), .A2(n3585), .ZN(n3641) );
  XOR2_X1 U3617 ( .A(n3642), .B(n3643), .Z(n3584) );
  XOR2_X1 U3618 ( .A(n3644), .B(n3645), .Z(n3643) );
  NAND2_X1 U3619 ( .A1(b_5_), .A2(a_7_), .ZN(n3645) );
  NAND2_X1 U3620 ( .A1(n3646), .A2(n2331), .ZN(n3639) );
  INV_X1 U3621 ( .A(n3586), .ZN(n2331) );
  NOR2_X1 U3622 ( .A1(n2454), .A2(n2455), .ZN(n3586) );
  INV_X1 U3623 ( .A(n3585), .ZN(n3646) );
  NAND2_X1 U3624 ( .A1(n3647), .A2(n3648), .ZN(n3585) );
  NAND2_X1 U3625 ( .A1(n3523), .A2(n3649), .ZN(n3648) );
  INV_X1 U3626 ( .A(n3650), .ZN(n3649) );
  NOR2_X1 U3627 ( .A1(n3522), .A2(n3520), .ZN(n3650) );
  NOR2_X1 U3628 ( .A1(n2454), .A2(n2312), .ZN(n3523) );
  NAND2_X1 U3629 ( .A1(n3520), .A2(n3522), .ZN(n3647) );
  NAND2_X1 U3630 ( .A1(n3651), .A2(n3652), .ZN(n3522) );
  NAND3_X1 U3631 ( .A1(a_8_), .A2(n3653), .A3(b_6_), .ZN(n3652) );
  INV_X1 U3632 ( .A(n3654), .ZN(n3653) );
  NOR2_X1 U3633 ( .A1(n3529), .A2(n3527), .ZN(n3654) );
  NAND2_X1 U3634 ( .A1(n3527), .A2(n3529), .ZN(n3651) );
  NAND2_X1 U3635 ( .A1(n3581), .A2(n3655), .ZN(n3529) );
  NAND2_X1 U3636 ( .A1(n3580), .A2(n3582), .ZN(n3655) );
  NAND2_X1 U3637 ( .A1(n3656), .A2(n3657), .ZN(n3582) );
  NAND2_X1 U3638 ( .A1(b_6_), .A2(a_9_), .ZN(n3657) );
  INV_X1 U3639 ( .A(n3658), .ZN(n3656) );
  XNOR2_X1 U3640 ( .A(n3659), .B(n3660), .ZN(n3580) );
  NAND2_X1 U3641 ( .A1(n3661), .A2(n3662), .ZN(n3659) );
  NAND2_X1 U3642 ( .A1(a_9_), .A2(n3658), .ZN(n3581) );
  NAND2_X1 U3643 ( .A1(n3542), .A2(n3663), .ZN(n3658) );
  NAND2_X1 U3644 ( .A1(n3541), .A2(n3543), .ZN(n3663) );
  NAND2_X1 U3645 ( .A1(n3664), .A2(n3665), .ZN(n3543) );
  NAND2_X1 U3646 ( .A1(b_6_), .A2(a_10_), .ZN(n3665) );
  XNOR2_X1 U3647 ( .A(n3666), .B(n3667), .ZN(n3541) );
  XOR2_X1 U3648 ( .A(n3668), .B(n3669), .Z(n3666) );
  NAND2_X1 U3649 ( .A1(b_5_), .A2(a_11_), .ZN(n3668) );
  INV_X1 U3650 ( .A(n3670), .ZN(n3542) );
  NOR2_X1 U3651 ( .A1(n2453), .A2(n3664), .ZN(n3670) );
  NOR2_X1 U3652 ( .A1(n3671), .A2(n3672), .ZN(n3664) );
  INV_X1 U3653 ( .A(n3673), .ZN(n3672) );
  NAND3_X1 U3654 ( .A1(a_11_), .A2(n3674), .A3(b_6_), .ZN(n3673) );
  NAND2_X1 U3655 ( .A1(n3548), .A2(n3550), .ZN(n3674) );
  NOR2_X1 U3656 ( .A1(n3548), .A2(n3550), .ZN(n3671) );
  NOR2_X1 U3657 ( .A1(n3675), .A2(n3676), .ZN(n3550) );
  INV_X1 U3658 ( .A(n3677), .ZN(n3676) );
  NAND2_X1 U3659 ( .A1(n3577), .A2(n3678), .ZN(n3677) );
  NAND2_X1 U3660 ( .A1(n3578), .A2(n3576), .ZN(n3678) );
  NOR2_X1 U3661 ( .A1(n2454), .A2(n2238), .ZN(n3577) );
  NOR2_X1 U3662 ( .A1(n3576), .A2(n3578), .ZN(n3675) );
  NOR2_X1 U3663 ( .A1(n3679), .A2(n3680), .ZN(n3578) );
  INV_X1 U3664 ( .A(n3681), .ZN(n3680) );
  NAND2_X1 U3665 ( .A1(n3572), .A2(n3682), .ZN(n3681) );
  NAND2_X1 U3666 ( .A1(n3573), .A2(n3574), .ZN(n3682) );
  NOR2_X1 U3667 ( .A1(n2454), .A2(n2223), .ZN(n3572) );
  NOR2_X1 U3668 ( .A1(n3574), .A2(n3573), .ZN(n3679) );
  INV_X1 U3669 ( .A(n3683), .ZN(n3573) );
  NAND2_X1 U3670 ( .A1(n3684), .A2(n3685), .ZN(n3683) );
  NAND2_X1 U3671 ( .A1(b_4_), .A2(n3686), .ZN(n3685) );
  NAND2_X1 U3672 ( .A1(n2202), .A2(n3687), .ZN(n3686) );
  NAND2_X1 U3673 ( .A1(a_15_), .A2(n2343), .ZN(n3687) );
  NAND2_X1 U3674 ( .A1(b_5_), .A2(n3688), .ZN(n3684) );
  NAND2_X1 U3675 ( .A1(n2205), .A2(n3689), .ZN(n3688) );
  NAND2_X1 U3676 ( .A1(a_14_), .A2(n2456), .ZN(n3689) );
  NAND3_X1 U3677 ( .A1(b_6_), .A2(b_5_), .A3(n2450), .ZN(n3574) );
  XNOR2_X1 U3678 ( .A(n3690), .B(n3691), .ZN(n3576) );
  XOR2_X1 U3679 ( .A(n3692), .B(n3693), .Z(n3690) );
  XOR2_X1 U3680 ( .A(n3694), .B(n3695), .Z(n3548) );
  XNOR2_X1 U3681 ( .A(n3696), .B(n3697), .ZN(n3694) );
  XNOR2_X1 U3682 ( .A(n3698), .B(n3699), .ZN(n3527) );
  NAND2_X1 U3683 ( .A1(n3700), .A2(n3701), .ZN(n3698) );
  XNOR2_X1 U3684 ( .A(n3702), .B(n3703), .ZN(n3520) );
  XOR2_X1 U3685 ( .A(n3704), .B(n3705), .Z(n3703) );
  NAND2_X1 U3686 ( .A1(b_5_), .A2(a_8_), .ZN(n3705) );
  XOR2_X1 U3687 ( .A(n3706), .B(n3707), .Z(n3588) );
  XOR2_X1 U3688 ( .A(n3708), .B(n3709), .Z(n3707) );
  NAND2_X1 U3689 ( .A1(b_5_), .A2(a_6_), .ZN(n3709) );
  XOR2_X1 U3690 ( .A(n3710), .B(n3711), .Z(n3592) );
  XOR2_X1 U3691 ( .A(n3712), .B(n2338), .Z(n3710) );
  XNOR2_X1 U3692 ( .A(n3713), .B(n3714), .ZN(n3595) );
  XOR2_X1 U3693 ( .A(n3715), .B(n3716), .Z(n3714) );
  NAND2_X1 U3694 ( .A1(a_4_), .A2(b_5_), .ZN(n3716) );
  XOR2_X1 U3695 ( .A(n3717), .B(n3718), .Z(n3600) );
  XNOR2_X1 U3696 ( .A(n3719), .B(n3720), .ZN(n3718) );
  NAND2_X1 U3697 ( .A1(a_3_), .A2(b_5_), .ZN(n3720) );
  XNOR2_X1 U3698 ( .A(n3721), .B(n3722), .ZN(n3604) );
  XOR2_X1 U3699 ( .A(n3723), .B(n3724), .Z(n3721) );
  NAND2_X1 U3700 ( .A1(a_2_), .A2(b_5_), .ZN(n3723) );
  XNOR2_X1 U3701 ( .A(n3725), .B(n3726), .ZN(n3608) );
  XNOR2_X1 U3702 ( .A(n3727), .B(n3728), .ZN(n3725) );
  NOR2_X1 U3703 ( .A1(n2647), .A2(n2343), .ZN(n3728) );
  XNOR2_X1 U3704 ( .A(n3729), .B(n3730), .ZN(n2177) );
  XNOR2_X1 U3705 ( .A(n3731), .B(n3732), .ZN(n3729) );
  NAND2_X1 U3706 ( .A1(a_0_), .A2(b_5_), .ZN(n3731) );
  INV_X1 U3707 ( .A(n3733), .ZN(n2501) );
  NOR2_X1 U3708 ( .A1(n3613), .A2(n3612), .ZN(n3733) );
  NOR2_X1 U3709 ( .A1(n3734), .A2(n3735), .ZN(n3612) );
  NOR3_X1 U3710 ( .A1(n2343), .A2(n3736), .A3(n2420), .ZN(n3735) );
  NOR2_X1 U3711 ( .A1(n3732), .A2(n3730), .ZN(n3736) );
  INV_X1 U3712 ( .A(n3737), .ZN(n3734) );
  NAND2_X1 U3713 ( .A1(n3730), .A2(n3732), .ZN(n3737) );
  NAND2_X1 U3714 ( .A1(n3738), .A2(n3739), .ZN(n3732) );
  NAND3_X1 U3715 ( .A1(a_1_), .A2(n3740), .A3(b_5_), .ZN(n3739) );
  NAND2_X1 U3716 ( .A1(n3726), .A2(n3727), .ZN(n3740) );
  INV_X1 U3717 ( .A(n3741), .ZN(n3738) );
  NOR2_X1 U3718 ( .A1(n3726), .A2(n3727), .ZN(n3741) );
  NOR2_X1 U3719 ( .A1(n3742), .A2(n3743), .ZN(n3727) );
  INV_X1 U3720 ( .A(n3744), .ZN(n3743) );
  NAND3_X1 U3721 ( .A1(b_5_), .A2(n3745), .A3(a_2_), .ZN(n3744) );
  NAND2_X1 U3722 ( .A1(n3724), .A2(n3722), .ZN(n3745) );
  NOR2_X1 U3723 ( .A1(n3722), .A2(n3724), .ZN(n3742) );
  NOR2_X1 U3724 ( .A1(n3746), .A2(n3747), .ZN(n3724) );
  NOR3_X1 U3725 ( .A1(n2343), .A2(n3748), .A3(n2376), .ZN(n3747) );
  INV_X1 U3726 ( .A(n3749), .ZN(n3748) );
  NAND2_X1 U3727 ( .A1(n3717), .A2(n3719), .ZN(n3749) );
  NOR2_X1 U3728 ( .A1(n3717), .A2(n3719), .ZN(n3746) );
  NOR2_X1 U3729 ( .A1(n3750), .A2(n3751), .ZN(n3719) );
  INV_X1 U3730 ( .A(n3752), .ZN(n3751) );
  NAND3_X1 U3731 ( .A1(b_5_), .A2(n3753), .A3(a_4_), .ZN(n3752) );
  NAND2_X1 U3732 ( .A1(n3713), .A2(n3715), .ZN(n3753) );
  NOR2_X1 U3733 ( .A1(n3715), .A2(n3713), .ZN(n3750) );
  XNOR2_X1 U3734 ( .A(n3754), .B(n3755), .ZN(n3713) );
  XOR2_X1 U3735 ( .A(n3756), .B(n3757), .Z(n3754) );
  NAND2_X1 U3736 ( .A1(n3758), .A2(n3759), .ZN(n3715) );
  NAND2_X1 U3737 ( .A1(n3711), .A2(n3760), .ZN(n3759) );
  NAND2_X1 U3738 ( .A1(n2338), .A2(n3712), .ZN(n3760) );
  INV_X1 U3739 ( .A(n2429), .ZN(n2338) );
  XNOR2_X1 U3740 ( .A(n3761), .B(n3762), .ZN(n3711) );
  XOR2_X1 U3741 ( .A(n3763), .B(n3764), .Z(n3761) );
  NAND2_X1 U3742 ( .A1(n3765), .A2(n2429), .ZN(n3758) );
  NAND2_X1 U3743 ( .A1(a_5_), .A2(b_5_), .ZN(n2429) );
  INV_X1 U3744 ( .A(n3712), .ZN(n3765) );
  NAND2_X1 U3745 ( .A1(n3766), .A2(n3767), .ZN(n3712) );
  NAND3_X1 U3746 ( .A1(a_6_), .A2(n3768), .A3(b_5_), .ZN(n3767) );
  INV_X1 U3747 ( .A(n3769), .ZN(n3768) );
  NOR2_X1 U3748 ( .A1(n3706), .A2(n3708), .ZN(n3769) );
  NAND2_X1 U3749 ( .A1(n3706), .A2(n3708), .ZN(n3766) );
  NAND2_X1 U3750 ( .A1(n3770), .A2(n3771), .ZN(n3708) );
  NAND3_X1 U3751 ( .A1(a_7_), .A2(n3772), .A3(b_5_), .ZN(n3771) );
  INV_X1 U3752 ( .A(n3773), .ZN(n3772) );
  NOR2_X1 U3753 ( .A1(n3644), .A2(n3642), .ZN(n3773) );
  NAND2_X1 U3754 ( .A1(n3642), .A2(n3644), .ZN(n3770) );
  NAND2_X1 U3755 ( .A1(n3774), .A2(n3775), .ZN(n3644) );
  INV_X1 U3756 ( .A(n3776), .ZN(n3775) );
  NOR3_X1 U3757 ( .A1(n2681), .A2(n3777), .A3(n2343), .ZN(n3776) );
  NOR2_X1 U3758 ( .A1(n3702), .A2(n3704), .ZN(n3777) );
  NAND2_X1 U3759 ( .A1(n3702), .A2(n3704), .ZN(n3774) );
  NAND2_X1 U3760 ( .A1(n3700), .A2(n3778), .ZN(n3704) );
  NAND2_X1 U3761 ( .A1(n3699), .A2(n3701), .ZN(n3778) );
  NAND2_X1 U3762 ( .A1(n3779), .A2(n3780), .ZN(n3701) );
  NAND2_X1 U3763 ( .A1(b_5_), .A2(a_9_), .ZN(n3780) );
  INV_X1 U3764 ( .A(n3781), .ZN(n3779) );
  XOR2_X1 U3765 ( .A(n3782), .B(n3783), .Z(n3699) );
  XNOR2_X1 U3766 ( .A(n3784), .B(n3785), .ZN(n3783) );
  NAND2_X1 U3767 ( .A1(a_9_), .A2(n3781), .ZN(n3700) );
  NAND2_X1 U3768 ( .A1(n3661), .A2(n3786), .ZN(n3781) );
  NAND2_X1 U3769 ( .A1(n3660), .A2(n3662), .ZN(n3786) );
  NAND2_X1 U3770 ( .A1(n3787), .A2(n3788), .ZN(n3662) );
  NAND2_X1 U3771 ( .A1(b_5_), .A2(a_10_), .ZN(n3788) );
  XNOR2_X1 U3772 ( .A(n3789), .B(n3790), .ZN(n3660) );
  XOR2_X1 U3773 ( .A(n3791), .B(n3792), .Z(n3789) );
  NAND2_X1 U3774 ( .A1(b_4_), .A2(a_11_), .ZN(n3791) );
  INV_X1 U3775 ( .A(n3793), .ZN(n3661) );
  NOR2_X1 U3776 ( .A1(n2453), .A2(n3787), .ZN(n3793) );
  NOR2_X1 U3777 ( .A1(n3794), .A2(n3795), .ZN(n3787) );
  INV_X1 U3778 ( .A(n3796), .ZN(n3795) );
  NAND3_X1 U3779 ( .A1(a_11_), .A2(n3797), .A3(b_5_), .ZN(n3796) );
  NAND2_X1 U3780 ( .A1(n3667), .A2(n3669), .ZN(n3797) );
  NOR2_X1 U3781 ( .A1(n3667), .A2(n3669), .ZN(n3794) );
  NOR2_X1 U3782 ( .A1(n3798), .A2(n3799), .ZN(n3669) );
  INV_X1 U3783 ( .A(n3800), .ZN(n3799) );
  NAND2_X1 U3784 ( .A1(n3696), .A2(n3801), .ZN(n3800) );
  NAND2_X1 U3785 ( .A1(n3697), .A2(n3695), .ZN(n3801) );
  NOR2_X1 U3786 ( .A1(n2343), .A2(n2238), .ZN(n3696) );
  NOR2_X1 U3787 ( .A1(n3695), .A2(n3697), .ZN(n3798) );
  NOR2_X1 U3788 ( .A1(n3802), .A2(n3803), .ZN(n3697) );
  INV_X1 U3789 ( .A(n3804), .ZN(n3803) );
  NAND2_X1 U3790 ( .A1(n3691), .A2(n3805), .ZN(n3804) );
  NAND2_X1 U3791 ( .A1(n3692), .A2(n3693), .ZN(n3805) );
  NOR2_X1 U3792 ( .A1(n2343), .A2(n2223), .ZN(n3691) );
  NOR2_X1 U3793 ( .A1(n3693), .A2(n3692), .ZN(n3802) );
  INV_X1 U3794 ( .A(n3806), .ZN(n3692) );
  NAND2_X1 U3795 ( .A1(n3807), .A2(n3808), .ZN(n3806) );
  NAND2_X1 U3796 ( .A1(b_3_), .A2(n3809), .ZN(n3808) );
  NAND2_X1 U3797 ( .A1(n2202), .A2(n3810), .ZN(n3809) );
  NAND2_X1 U3798 ( .A1(a_15_), .A2(n2456), .ZN(n3810) );
  NAND2_X1 U3799 ( .A1(b_4_), .A2(n3811), .ZN(n3807) );
  NAND2_X1 U3800 ( .A1(n2205), .A2(n3812), .ZN(n3811) );
  NAND2_X1 U3801 ( .A1(a_14_), .A2(n2378), .ZN(n3812) );
  NAND3_X1 U3802 ( .A1(b_4_), .A2(b_5_), .A3(n2450), .ZN(n3693) );
  XNOR2_X1 U3803 ( .A(n3813), .B(n3814), .ZN(n3695) );
  XOR2_X1 U3804 ( .A(n3815), .B(n3816), .Z(n3813) );
  XOR2_X1 U3805 ( .A(n3817), .B(n3818), .Z(n3667) );
  XNOR2_X1 U3806 ( .A(n3819), .B(n3820), .ZN(n3817) );
  XNOR2_X1 U3807 ( .A(n3821), .B(n3822), .ZN(n3702) );
  XNOR2_X1 U3808 ( .A(n3823), .B(n3824), .ZN(n3822) );
  XNOR2_X1 U3809 ( .A(n3825), .B(n3826), .ZN(n3642) );
  XNOR2_X1 U3810 ( .A(n3827), .B(n3828), .ZN(n3825) );
  XOR2_X1 U3811 ( .A(n3829), .B(n3830), .Z(n3706) );
  XOR2_X1 U3812 ( .A(n3831), .B(n3832), .Z(n3829) );
  XOR2_X1 U3813 ( .A(n3833), .B(n3834), .Z(n3717) );
  XOR2_X1 U3814 ( .A(n3835), .B(n2458), .Z(n3833) );
  XOR2_X1 U3815 ( .A(n3836), .B(n3837), .Z(n3722) );
  XNOR2_X1 U3816 ( .A(n3838), .B(n3839), .ZN(n3837) );
  XNOR2_X1 U3817 ( .A(n3840), .B(n3841), .ZN(n3726) );
  XOR2_X1 U3818 ( .A(n3842), .B(n3843), .Z(n3841) );
  XNOR2_X1 U3819 ( .A(n3844), .B(n3845), .ZN(n3730) );
  XNOR2_X1 U3820 ( .A(n3846), .B(n3847), .ZN(n3844) );
  XOR2_X1 U3821 ( .A(n3848), .B(n3849), .Z(n3613) );
  XNOR2_X1 U3822 ( .A(n3850), .B(n3851), .ZN(n3848) );
  XOR2_X1 U3823 ( .A(n2188), .B(n2189), .Z(n2180) );
  INV_X1 U3824 ( .A(n2184), .ZN(n2498) );
  NOR3_X1 U3825 ( .A1(n2189), .A2(n2188), .A3(n2500), .ZN(n2184) );
  NAND2_X1 U3826 ( .A1(n2497), .A2(n3852), .ZN(n2500) );
  NAND2_X1 U3827 ( .A1(n3853), .A2(n3854), .ZN(n3852) );
  NOR2_X1 U3828 ( .A1(n3855), .A2(n3856), .ZN(n2188) );
  INV_X1 U3829 ( .A(n3857), .ZN(n3856) );
  NAND2_X1 U3830 ( .A1(n3851), .A2(n3858), .ZN(n3857) );
  NAND2_X1 U3831 ( .A1(n3850), .A2(n3849), .ZN(n3858) );
  NOR2_X1 U3832 ( .A1(n2420), .A2(n2456), .ZN(n3851) );
  NOR2_X1 U3833 ( .A1(n3849), .A2(n3850), .ZN(n3855) );
  NOR2_X1 U3834 ( .A1(n3859), .A2(n3860), .ZN(n3850) );
  INV_X1 U3835 ( .A(n3861), .ZN(n3860) );
  NAND2_X1 U3836 ( .A1(n3846), .A2(n3862), .ZN(n3861) );
  NAND2_X1 U3837 ( .A1(n3845), .A2(n3847), .ZN(n3862) );
  NOR2_X1 U3838 ( .A1(n2456), .A2(n2647), .ZN(n3846) );
  NOR2_X1 U3839 ( .A1(n3845), .A2(n3847), .ZN(n3859) );
  NOR2_X1 U3840 ( .A1(n3863), .A2(n3864), .ZN(n3847) );
  INV_X1 U3841 ( .A(n3865), .ZN(n3864) );
  NAND2_X1 U3842 ( .A1(n3843), .A2(n3866), .ZN(n3865) );
  NAND2_X1 U3843 ( .A1(n3842), .A2(n3840), .ZN(n3866) );
  NOR2_X1 U3844 ( .A1(n2460), .A2(n2456), .ZN(n3843) );
  NOR2_X1 U3845 ( .A1(n3840), .A2(n3842), .ZN(n3863) );
  NOR2_X1 U3846 ( .A1(n3867), .A2(n3868), .ZN(n3842) );
  INV_X1 U3847 ( .A(n3869), .ZN(n3868) );
  NAND2_X1 U3848 ( .A1(n3839), .A2(n3870), .ZN(n3869) );
  NAND2_X1 U3849 ( .A1(n3836), .A2(n3838), .ZN(n3870) );
  NOR2_X1 U3850 ( .A1(n2376), .A2(n2456), .ZN(n3839) );
  NOR2_X1 U3851 ( .A1(n3836), .A2(n3838), .ZN(n3867) );
  NAND2_X1 U3852 ( .A1(n3871), .A2(n3872), .ZN(n3838) );
  NAND2_X1 U3853 ( .A1(n3834), .A2(n3873), .ZN(n3872) );
  NAND2_X1 U3854 ( .A1(n2458), .A2(n3835), .ZN(n3873) );
  XNOR2_X1 U3855 ( .A(n3874), .B(n3875), .ZN(n3834) );
  XNOR2_X1 U3856 ( .A(n3876), .B(n3877), .ZN(n3874) );
  NAND2_X1 U3857 ( .A1(b_3_), .A2(a_5_), .ZN(n3876) );
  INV_X1 U3858 ( .A(n3878), .ZN(n3871) );
  NOR2_X1 U3859 ( .A1(n3835), .A2(n2458), .ZN(n3878) );
  NOR2_X1 U3860 ( .A1(n2456), .A2(n2457), .ZN(n2458) );
  NAND2_X1 U3861 ( .A1(n3879), .A2(n3880), .ZN(n3835) );
  NAND2_X1 U3862 ( .A1(n3757), .A2(n3881), .ZN(n3880) );
  INV_X1 U3863 ( .A(n3882), .ZN(n3881) );
  NOR2_X1 U3864 ( .A1(n3756), .A2(n3755), .ZN(n3882) );
  NOR2_X1 U3865 ( .A1(n2456), .A2(n2341), .ZN(n3757) );
  NAND2_X1 U3866 ( .A1(n3755), .A2(n3756), .ZN(n3879) );
  NAND2_X1 U3867 ( .A1(n3883), .A2(n3884), .ZN(n3756) );
  NAND2_X1 U3868 ( .A1(n3764), .A2(n3885), .ZN(n3884) );
  INV_X1 U3869 ( .A(n3886), .ZN(n3885) );
  NOR2_X1 U3870 ( .A1(n3762), .A2(n3763), .ZN(n3886) );
  NOR2_X1 U3871 ( .A1(n2456), .A2(n2455), .ZN(n3764) );
  NAND2_X1 U3872 ( .A1(n3762), .A2(n3763), .ZN(n3883) );
  NAND2_X1 U3873 ( .A1(n3887), .A2(n3888), .ZN(n3763) );
  NAND2_X1 U3874 ( .A1(n3832), .A2(n3889), .ZN(n3888) );
  INV_X1 U3875 ( .A(n3890), .ZN(n3889) );
  NOR2_X1 U3876 ( .A1(n3831), .A2(n3830), .ZN(n3890) );
  NOR2_X1 U3877 ( .A1(n2456), .A2(n2312), .ZN(n3832) );
  NAND2_X1 U3878 ( .A1(n3830), .A2(n3831), .ZN(n3887) );
  NAND2_X1 U3879 ( .A1(n3891), .A2(n3892), .ZN(n3831) );
  NAND2_X1 U3880 ( .A1(n3828), .A2(n3893), .ZN(n3892) );
  NAND2_X1 U3881 ( .A1(n3826), .A2(n3827), .ZN(n3893) );
  NOR2_X1 U3882 ( .A1(n2456), .A2(n2681), .ZN(n3828) );
  INV_X1 U3883 ( .A(n3894), .ZN(n3891) );
  NOR2_X1 U3884 ( .A1(n3826), .A2(n3827), .ZN(n3894) );
  NOR2_X1 U3885 ( .A1(n3895), .A2(n3896), .ZN(n3827) );
  INV_X1 U3886 ( .A(n3897), .ZN(n3896) );
  NAND2_X1 U3887 ( .A1(n3824), .A2(n3898), .ZN(n3897) );
  NAND2_X1 U3888 ( .A1(n3821), .A2(n3823), .ZN(n3898) );
  NOR2_X1 U3889 ( .A1(n2456), .A2(n2283), .ZN(n3824) );
  NOR2_X1 U3890 ( .A1(n3823), .A2(n3821), .ZN(n3895) );
  XOR2_X1 U3891 ( .A(n3899), .B(n3900), .Z(n3821) );
  NAND2_X1 U3892 ( .A1(n3901), .A2(n3902), .ZN(n3899) );
  NAND2_X1 U3893 ( .A1(n3903), .A2(n3904), .ZN(n3823) );
  NAND2_X1 U3894 ( .A1(n3782), .A2(n3905), .ZN(n3904) );
  INV_X1 U3895 ( .A(n3906), .ZN(n3905) );
  NOR2_X1 U3896 ( .A1(n3785), .A2(n3784), .ZN(n3906) );
  XOR2_X1 U3897 ( .A(n3907), .B(n3908), .Z(n3782) );
  XOR2_X1 U3898 ( .A(n3909), .B(n3910), .Z(n3907) );
  NAND2_X1 U3899 ( .A1(b_3_), .A2(a_11_), .ZN(n3909) );
  NAND2_X1 U3900 ( .A1(n3784), .A2(n3785), .ZN(n3903) );
  NAND2_X1 U3901 ( .A1(b_4_), .A2(a_10_), .ZN(n3785) );
  NOR2_X1 U3902 ( .A1(n3911), .A2(n3912), .ZN(n3784) );
  NOR3_X1 U3903 ( .A1(n2254), .A2(n3913), .A3(n2456), .ZN(n3912) );
  INV_X1 U3904 ( .A(n3914), .ZN(n3913) );
  NAND2_X1 U3905 ( .A1(n3790), .A2(n3792), .ZN(n3914) );
  NOR2_X1 U3906 ( .A1(n3790), .A2(n3792), .ZN(n3911) );
  NOR2_X1 U3907 ( .A1(n3915), .A2(n3916), .ZN(n3792) );
  INV_X1 U3908 ( .A(n3917), .ZN(n3916) );
  NAND2_X1 U3909 ( .A1(n3819), .A2(n3918), .ZN(n3917) );
  NAND2_X1 U3910 ( .A1(n3820), .A2(n3818), .ZN(n3918) );
  NOR2_X1 U3911 ( .A1(n2456), .A2(n2238), .ZN(n3819) );
  NOR2_X1 U3912 ( .A1(n3818), .A2(n3820), .ZN(n3915) );
  NOR2_X1 U3913 ( .A1(n3919), .A2(n3920), .ZN(n3820) );
  INV_X1 U3914 ( .A(n3921), .ZN(n3920) );
  NAND2_X1 U3915 ( .A1(n3814), .A2(n3922), .ZN(n3921) );
  NAND2_X1 U3916 ( .A1(n3815), .A2(n3816), .ZN(n3922) );
  NOR2_X1 U3917 ( .A1(n2456), .A2(n2223), .ZN(n3814) );
  NOR2_X1 U3918 ( .A1(n3816), .A2(n3815), .ZN(n3919) );
  INV_X1 U3919 ( .A(n3923), .ZN(n3815) );
  NAND2_X1 U3920 ( .A1(n3924), .A2(n3925), .ZN(n3923) );
  NAND2_X1 U3921 ( .A1(b_2_), .A2(n3926), .ZN(n3925) );
  NAND2_X1 U3922 ( .A1(n2202), .A2(n3927), .ZN(n3926) );
  NAND2_X1 U3923 ( .A1(a_15_), .A2(n2378), .ZN(n3927) );
  NAND2_X1 U3924 ( .A1(b_3_), .A2(n3928), .ZN(n3924) );
  NAND2_X1 U3925 ( .A1(n2205), .A2(n3929), .ZN(n3928) );
  NAND2_X1 U3926 ( .A1(a_14_), .A2(n2459), .ZN(n3929) );
  NAND3_X1 U3927 ( .A1(b_4_), .A2(b_3_), .A3(n2450), .ZN(n3816) );
  XNOR2_X1 U3928 ( .A(n3930), .B(n3931), .ZN(n3818) );
  XOR2_X1 U3929 ( .A(n3932), .B(n3933), .Z(n3930) );
  XOR2_X1 U3930 ( .A(n3934), .B(n3935), .Z(n3790) );
  XNOR2_X1 U3931 ( .A(n3936), .B(n3937), .ZN(n3934) );
  XOR2_X1 U3932 ( .A(n3938), .B(n3939), .Z(n3826) );
  NAND2_X1 U3933 ( .A1(n3940), .A2(n3941), .ZN(n3938) );
  XOR2_X1 U3934 ( .A(n3942), .B(n3943), .Z(n3830) );
  XOR2_X1 U3935 ( .A(n3944), .B(n3945), .Z(n3942) );
  NOR2_X1 U3936 ( .A1(n2681), .A2(n2378), .ZN(n3945) );
  XNOR2_X1 U3937 ( .A(n3946), .B(n3947), .ZN(n3762) );
  NAND2_X1 U3938 ( .A1(n3948), .A2(n3949), .ZN(n3946) );
  XOR2_X1 U3939 ( .A(n3950), .B(n3951), .Z(n3755) );
  XOR2_X1 U3940 ( .A(n3952), .B(n3953), .Z(n3950) );
  NOR2_X1 U3941 ( .A1(n2455), .A2(n2378), .ZN(n3953) );
  XOR2_X1 U3942 ( .A(n3954), .B(n3955), .Z(n3836) );
  XNOR2_X1 U3943 ( .A(n3956), .B(n3957), .ZN(n3954) );
  NOR2_X1 U3944 ( .A1(n2457), .A2(n2378), .ZN(n3957) );
  XNOR2_X1 U3945 ( .A(n3958), .B(n3959), .ZN(n3840) );
  XOR2_X1 U3946 ( .A(n2374), .B(n3960), .Z(n3958) );
  XNOR2_X1 U3947 ( .A(n3961), .B(n3962), .ZN(n3845) );
  XNOR2_X1 U3948 ( .A(n3963), .B(n3964), .ZN(n3961) );
  NAND2_X1 U3949 ( .A1(a_2_), .A2(b_3_), .ZN(n3963) );
  XOR2_X1 U3950 ( .A(n3965), .B(n3966), .Z(n3849) );
  XNOR2_X1 U3951 ( .A(n3967), .B(n3968), .ZN(n3965) );
  NOR2_X1 U3952 ( .A1(n2647), .A2(n2378), .ZN(n3968) );
  XNOR2_X1 U3953 ( .A(n3969), .B(n3970), .ZN(n2189) );
  XNOR2_X1 U3954 ( .A(n3971), .B(n3972), .ZN(n3970) );
  NAND2_X1 U3955 ( .A1(a_0_), .A2(b_3_), .ZN(n3972) );
  INV_X1 U3956 ( .A(n3973), .ZN(n2497) );
  NOR2_X1 U3957 ( .A1(n3854), .A2(n3853), .ZN(n3973) );
  NOR2_X1 U3958 ( .A1(n3974), .A2(n3975), .ZN(n3853) );
  NOR3_X1 U3959 ( .A1(n2378), .A2(n3976), .A3(n2420), .ZN(n3975) );
  INV_X1 U3960 ( .A(n3977), .ZN(n3976) );
  NAND2_X1 U3961 ( .A1(n3971), .A2(n3969), .ZN(n3977) );
  NOR2_X1 U3962 ( .A1(n3969), .A2(n3971), .ZN(n3974) );
  NOR2_X1 U3963 ( .A1(n3978), .A2(n3979), .ZN(n3971) );
  NOR3_X1 U3964 ( .A1(n2647), .A2(n3980), .A3(n2378), .ZN(n3979) );
  INV_X1 U3965 ( .A(n3981), .ZN(n3980) );
  NAND2_X1 U3966 ( .A1(n3966), .A2(n3967), .ZN(n3981) );
  NOR2_X1 U3967 ( .A1(n3966), .A2(n3967), .ZN(n3978) );
  NOR2_X1 U3968 ( .A1(n3982), .A2(n3983), .ZN(n3967) );
  INV_X1 U3969 ( .A(n3984), .ZN(n3983) );
  NAND3_X1 U3970 ( .A1(b_3_), .A2(n3985), .A3(a_2_), .ZN(n3984) );
  NAND2_X1 U3971 ( .A1(n3962), .A2(n3964), .ZN(n3985) );
  NOR2_X1 U3972 ( .A1(n3964), .A2(n3962), .ZN(n3982) );
  XOR2_X1 U3973 ( .A(n3986), .B(n3987), .Z(n3962) );
  XNOR2_X1 U3974 ( .A(n3988), .B(n3989), .ZN(n3986) );
  NAND2_X1 U3975 ( .A1(n3990), .A2(n3991), .ZN(n3964) );
  INV_X1 U3976 ( .A(n3992), .ZN(n3991) );
  NOR2_X1 U3977 ( .A1(n3959), .A2(n3993), .ZN(n3992) );
  NOR2_X1 U3978 ( .A1(n2374), .A2(n3960), .ZN(n3993) );
  XNOR2_X1 U3979 ( .A(n3994), .B(n3995), .ZN(n3959) );
  XNOR2_X1 U3980 ( .A(n3996), .B(n3997), .ZN(n3994) );
  NAND2_X1 U3981 ( .A1(n3960), .A2(n2374), .ZN(n3990) );
  NAND2_X1 U3982 ( .A1(a_3_), .A2(b_3_), .ZN(n2374) );
  NOR2_X1 U3983 ( .A1(n3998), .A2(n3999), .ZN(n3960) );
  INV_X1 U3984 ( .A(n4000), .ZN(n3999) );
  NAND3_X1 U3985 ( .A1(a_4_), .A2(n4001), .A3(b_3_), .ZN(n4000) );
  NAND2_X1 U3986 ( .A1(n3955), .A2(n3956), .ZN(n4001) );
  NOR2_X1 U3987 ( .A1(n3955), .A2(n3956), .ZN(n3998) );
  NOR2_X1 U3988 ( .A1(n4002), .A2(n4003), .ZN(n3956) );
  NOR3_X1 U3989 ( .A1(n2341), .A2(n4004), .A3(n2378), .ZN(n4003) );
  NOR2_X1 U3990 ( .A1(n3875), .A2(n3877), .ZN(n4004) );
  INV_X1 U3991 ( .A(n4005), .ZN(n4002) );
  NAND2_X1 U3992 ( .A1(n3875), .A2(n3877), .ZN(n4005) );
  NAND2_X1 U3993 ( .A1(n4006), .A2(n4007), .ZN(n3877) );
  INV_X1 U3994 ( .A(n4008), .ZN(n4007) );
  NOR3_X1 U3995 ( .A1(n2455), .A2(n4009), .A3(n2378), .ZN(n4008) );
  NOR2_X1 U3996 ( .A1(n3951), .A2(n3952), .ZN(n4009) );
  NAND2_X1 U3997 ( .A1(n3951), .A2(n3952), .ZN(n4006) );
  NAND2_X1 U3998 ( .A1(n3948), .A2(n4010), .ZN(n3952) );
  NAND2_X1 U3999 ( .A1(n3947), .A2(n3949), .ZN(n4010) );
  NAND2_X1 U4000 ( .A1(n4011), .A2(n4012), .ZN(n3949) );
  NAND2_X1 U4001 ( .A1(b_3_), .A2(a_7_), .ZN(n4012) );
  XNOR2_X1 U4002 ( .A(n4013), .B(n4014), .ZN(n3947) );
  XNOR2_X1 U4003 ( .A(n4015), .B(n4016), .ZN(n4013) );
  NAND2_X1 U4004 ( .A1(a_7_), .A2(n4017), .ZN(n3948) );
  INV_X1 U4005 ( .A(n4011), .ZN(n4017) );
  NOR2_X1 U4006 ( .A1(n4018), .A2(n4019), .ZN(n4011) );
  NOR3_X1 U4007 ( .A1(n2681), .A2(n4020), .A3(n2378), .ZN(n4019) );
  NOR2_X1 U4008 ( .A1(n3943), .A2(n3944), .ZN(n4020) );
  INV_X1 U4009 ( .A(n4021), .ZN(n4018) );
  NAND2_X1 U4010 ( .A1(n3943), .A2(n3944), .ZN(n4021) );
  NAND2_X1 U4011 ( .A1(n3940), .A2(n4022), .ZN(n3944) );
  NAND2_X1 U4012 ( .A1(n3939), .A2(n3941), .ZN(n4022) );
  NAND2_X1 U4013 ( .A1(n4023), .A2(n4024), .ZN(n3941) );
  NAND2_X1 U4014 ( .A1(b_3_), .A2(a_9_), .ZN(n4024) );
  INV_X1 U4015 ( .A(n4025), .ZN(n4023) );
  XNOR2_X1 U4016 ( .A(n4026), .B(n4027), .ZN(n3939) );
  XOR2_X1 U4017 ( .A(n4028), .B(n4029), .Z(n4026) );
  NAND2_X1 U4018 ( .A1(a_9_), .A2(n4025), .ZN(n3940) );
  NAND2_X1 U4019 ( .A1(n3901), .A2(n4030), .ZN(n4025) );
  NAND2_X1 U4020 ( .A1(n3900), .A2(n3902), .ZN(n4030) );
  NAND2_X1 U4021 ( .A1(n4031), .A2(n4032), .ZN(n3902) );
  NAND2_X1 U4022 ( .A1(b_3_), .A2(a_10_), .ZN(n4032) );
  XNOR2_X1 U4023 ( .A(n4033), .B(n4034), .ZN(n3900) );
  XNOR2_X1 U4024 ( .A(n4035), .B(n4036), .ZN(n4034) );
  INV_X1 U4025 ( .A(n4037), .ZN(n3901) );
  NOR2_X1 U4026 ( .A1(n2453), .A2(n4031), .ZN(n4037) );
  NOR2_X1 U4027 ( .A1(n4038), .A2(n4039), .ZN(n4031) );
  INV_X1 U4028 ( .A(n4040), .ZN(n4039) );
  NAND3_X1 U4029 ( .A1(a_11_), .A2(n4041), .A3(b_3_), .ZN(n4040) );
  NAND2_X1 U4030 ( .A1(n3910), .A2(n3908), .ZN(n4041) );
  NOR2_X1 U4031 ( .A1(n3908), .A2(n3910), .ZN(n4038) );
  NOR2_X1 U4032 ( .A1(n4042), .A2(n4043), .ZN(n3910) );
  INV_X1 U4033 ( .A(n4044), .ZN(n4043) );
  NAND2_X1 U4034 ( .A1(n3936), .A2(n4045), .ZN(n4044) );
  NAND2_X1 U4035 ( .A1(n3937), .A2(n3935), .ZN(n4045) );
  NOR2_X1 U4036 ( .A1(n2378), .A2(n2238), .ZN(n3936) );
  NOR2_X1 U4037 ( .A1(n3935), .A2(n3937), .ZN(n4042) );
  NOR2_X1 U4038 ( .A1(n4046), .A2(n4047), .ZN(n3937) );
  INV_X1 U4039 ( .A(n4048), .ZN(n4047) );
  NAND2_X1 U4040 ( .A1(n3931), .A2(n4049), .ZN(n4048) );
  NAND2_X1 U4041 ( .A1(n3932), .A2(n3933), .ZN(n4049) );
  NOR2_X1 U4042 ( .A1(n2378), .A2(n2223), .ZN(n3931) );
  NOR2_X1 U4043 ( .A1(n3933), .A2(n3932), .ZN(n4046) );
  INV_X1 U4044 ( .A(n4050), .ZN(n3932) );
  NAND2_X1 U4045 ( .A1(n4051), .A2(n4052), .ZN(n4050) );
  NAND2_X1 U4046 ( .A1(b_1_), .A2(n4053), .ZN(n4052) );
  NAND2_X1 U4047 ( .A1(n2202), .A2(n4054), .ZN(n4053) );
  NAND2_X1 U4048 ( .A1(a_15_), .A2(n2459), .ZN(n4054) );
  NAND2_X1 U4049 ( .A1(b_2_), .A2(n4055), .ZN(n4051) );
  NAND2_X1 U4050 ( .A1(n2205), .A2(n4056), .ZN(n4055) );
  NAND2_X1 U4051 ( .A1(a_14_), .A2(n4057), .ZN(n4056) );
  NAND3_X1 U4052 ( .A1(b_2_), .A2(b_3_), .A3(n2450), .ZN(n3933) );
  XNOR2_X1 U4053 ( .A(n4058), .B(n4059), .ZN(n3935) );
  XOR2_X1 U4054 ( .A(n4060), .B(n4061), .Z(n4058) );
  XNOR2_X1 U4055 ( .A(n4062), .B(n4063), .ZN(n3908) );
  XNOR2_X1 U4056 ( .A(n4064), .B(n4065), .ZN(n4062) );
  XNOR2_X1 U4057 ( .A(n4066), .B(n4067), .ZN(n3943) );
  XNOR2_X1 U4058 ( .A(n4068), .B(n4069), .ZN(n4066) );
  XNOR2_X1 U4059 ( .A(n4070), .B(n4071), .ZN(n3951) );
  XNOR2_X1 U4060 ( .A(n4072), .B(n4073), .ZN(n4070) );
  XNOR2_X1 U4061 ( .A(n4074), .B(n4075), .ZN(n3875) );
  XNOR2_X1 U4062 ( .A(n4076), .B(n4077), .ZN(n4074) );
  XOR2_X1 U4063 ( .A(n4078), .B(n4079), .Z(n3955) );
  XNOR2_X1 U4064 ( .A(n4080), .B(n4081), .ZN(n4078) );
  XOR2_X1 U4065 ( .A(n4082), .B(n4083), .Z(n3966) );
  XOR2_X1 U4066 ( .A(n2395), .B(n4084), .Z(n4082) );
  XNOR2_X1 U4067 ( .A(n4085), .B(n4086), .ZN(n3969) );
  XOR2_X1 U4068 ( .A(n4087), .B(n4088), .Z(n4085) );
  XNOR2_X1 U4069 ( .A(n4089), .B(n4090), .ZN(n3854) );
  XNOR2_X1 U4070 ( .A(n4091), .B(n4092), .ZN(n4089) );
  NOR2_X1 U4071 ( .A1(n2459), .A2(n2420), .ZN(n4092) );
  XOR2_X1 U4072 ( .A(n2495), .B(n2496), .Z(n2213) );
  INV_X1 U4073 ( .A(n4093), .ZN(n2365) );
  NAND2_X1 U4074 ( .A1(n4094), .A2(n4095), .ZN(n4093) );
  NAND2_X1 U4075 ( .A1(b_0_), .A2(n2494), .ZN(n4095) );
  NAND2_X1 U4076 ( .A1(n4096), .A2(n4097), .ZN(n2494) );
  NAND2_X1 U4077 ( .A1(n2495), .A2(n2496), .ZN(n4094) );
  NAND3_X1 U4078 ( .A1(n4098), .A2(n4099), .A3(n4100), .ZN(n2496) );
  XNOR2_X1 U4079 ( .A(n4096), .B(n4097), .ZN(n4100) );
  NOR2_X1 U4080 ( .A1(n2647), .A2(n4101), .ZN(n4097) );
  NOR2_X1 U4081 ( .A1(n2420), .A2(n4057), .ZN(n4096) );
  NAND3_X1 U4082 ( .A1(a_2_), .A2(b_0_), .A3(n2409), .ZN(n4099) );
  NAND2_X1 U4083 ( .A1(n4091), .A2(n4102), .ZN(n2495) );
  NAND2_X1 U4084 ( .A1(n4090), .A2(b_2_), .ZN(n4102) );
  XNOR2_X1 U4085 ( .A(n4103), .B(n4104), .ZN(n4090) );
  NOR2_X1 U4086 ( .A1(n4101), .A2(n2460), .ZN(n4104) );
  NAND2_X1 U4087 ( .A1(n2409), .A2(n4098), .ZN(n4103) );
  NOR2_X1 U4088 ( .A1(n4105), .A2(n4106), .ZN(n4098) );
  INV_X1 U4089 ( .A(n4107), .ZN(n4106) );
  NAND3_X1 U4090 ( .A1(a_2_), .A2(n4108), .A3(b_1_), .ZN(n4107) );
  NAND2_X1 U4091 ( .A1(n4109), .A2(n4110), .ZN(n4108) );
  NOR2_X1 U4092 ( .A1(n4110), .A2(n4109), .ZN(n4105) );
  NOR2_X1 U4093 ( .A1(n4057), .A2(n2647), .ZN(n2409) );
  NOR2_X1 U4094 ( .A1(n4111), .A2(n4112), .ZN(n4091) );
  INV_X1 U4095 ( .A(n4113), .ZN(n4112) );
  NAND2_X1 U4096 ( .A1(n4087), .A2(n4114), .ZN(n4113) );
  NAND2_X1 U4097 ( .A1(n4086), .A2(n4088), .ZN(n4114) );
  NOR2_X1 U4098 ( .A1(n2459), .A2(n2647), .ZN(n4087) );
  NOR2_X1 U4099 ( .A1(n4086), .A2(n4088), .ZN(n4111) );
  NAND2_X1 U4100 ( .A1(n4115), .A2(n4116), .ZN(n4088) );
  NAND2_X1 U4101 ( .A1(n4083), .A2(n4117), .ZN(n4116) );
  INV_X1 U4102 ( .A(n4118), .ZN(n4117) );
  NOR2_X1 U4103 ( .A1(n2395), .A2(n4084), .ZN(n4118) );
  XNOR2_X1 U4104 ( .A(n4119), .B(n4120), .ZN(n4083) );
  NOR2_X1 U4105 ( .A1(n2376), .A2(n4057), .ZN(n4120) );
  XOR2_X1 U4106 ( .A(n4121), .B(n4122), .Z(n4119) );
  NAND2_X1 U4107 ( .A1(n4084), .A2(n2395), .ZN(n4115) );
  NAND2_X1 U4108 ( .A1(b_2_), .A2(a_2_), .ZN(n2395) );
  NOR2_X1 U4109 ( .A1(n4123), .A2(n4124), .ZN(n4084) );
  INV_X1 U4110 ( .A(n4125), .ZN(n4124) );
  NAND2_X1 U4111 ( .A1(n3989), .A2(n4126), .ZN(n4125) );
  NAND2_X1 U4112 ( .A1(n3988), .A2(n3987), .ZN(n4126) );
  NOR2_X1 U4113 ( .A1(n2459), .A2(n2376), .ZN(n3989) );
  NOR2_X1 U4114 ( .A1(n3987), .A2(n3988), .ZN(n4123) );
  NOR2_X1 U4115 ( .A1(n4127), .A2(n4128), .ZN(n3988) );
  INV_X1 U4116 ( .A(n4129), .ZN(n4128) );
  NAND2_X1 U4117 ( .A1(n3996), .A2(n4130), .ZN(n4129) );
  NAND2_X1 U4118 ( .A1(n3997), .A2(n3995), .ZN(n4130) );
  NOR2_X1 U4119 ( .A1(n2459), .A2(n2457), .ZN(n3996) );
  NOR2_X1 U4120 ( .A1(n3995), .A2(n3997), .ZN(n4127) );
  NOR2_X1 U4121 ( .A1(n4131), .A2(n4132), .ZN(n3997) );
  INV_X1 U4122 ( .A(n4133), .ZN(n4132) );
  NAND2_X1 U4123 ( .A1(n4081), .A2(n4134), .ZN(n4133) );
  NAND2_X1 U4124 ( .A1(n4080), .A2(n4079), .ZN(n4134) );
  NOR2_X1 U4125 ( .A1(n2459), .A2(n2341), .ZN(n4081) );
  NOR2_X1 U4126 ( .A1(n4079), .A2(n4080), .ZN(n4131) );
  NOR2_X1 U4127 ( .A1(n4135), .A2(n4136), .ZN(n4080) );
  INV_X1 U4128 ( .A(n4137), .ZN(n4136) );
  NAND2_X1 U4129 ( .A1(n4076), .A2(n4138), .ZN(n4137) );
  NAND2_X1 U4130 ( .A1(n4077), .A2(n4075), .ZN(n4138) );
  NOR2_X1 U4131 ( .A1(n2459), .A2(n2455), .ZN(n4076) );
  NOR2_X1 U4132 ( .A1(n4075), .A2(n4077), .ZN(n4135) );
  NOR2_X1 U4133 ( .A1(n4139), .A2(n4140), .ZN(n4077) );
  INV_X1 U4134 ( .A(n4141), .ZN(n4140) );
  NAND2_X1 U4135 ( .A1(n4073), .A2(n4142), .ZN(n4141) );
  NAND2_X1 U4136 ( .A1(n4072), .A2(n4071), .ZN(n4142) );
  NOR2_X1 U4137 ( .A1(n2459), .A2(n2312), .ZN(n4073) );
  NOR2_X1 U4138 ( .A1(n4071), .A2(n4072), .ZN(n4139) );
  NOR2_X1 U4139 ( .A1(n4143), .A2(n4144), .ZN(n4072) );
  INV_X1 U4140 ( .A(n4145), .ZN(n4144) );
  NAND2_X1 U4141 ( .A1(n4015), .A2(n4146), .ZN(n4145) );
  NAND2_X1 U4142 ( .A1(n4016), .A2(n4014), .ZN(n4146) );
  NOR2_X1 U4143 ( .A1(n2459), .A2(n2681), .ZN(n4015) );
  NOR2_X1 U4144 ( .A1(n4014), .A2(n4016), .ZN(n4143) );
  NOR2_X1 U4145 ( .A1(n4147), .A2(n4148), .ZN(n4016) );
  INV_X1 U4146 ( .A(n4149), .ZN(n4148) );
  NAND2_X1 U4147 ( .A1(n4069), .A2(n4150), .ZN(n4149) );
  NAND2_X1 U4148 ( .A1(n4068), .A2(n4067), .ZN(n4150) );
  NOR2_X1 U4149 ( .A1(n2459), .A2(n2283), .ZN(n4069) );
  NOR2_X1 U4150 ( .A1(n4067), .A2(n4068), .ZN(n4147) );
  NOR2_X1 U4151 ( .A1(n4151), .A2(n4152), .ZN(n4068) );
  INV_X1 U4152 ( .A(n4153), .ZN(n4152) );
  NAND2_X1 U4153 ( .A1(n4028), .A2(n4154), .ZN(n4153) );
  NAND2_X1 U4154 ( .A1(n4155), .A2(n4027), .ZN(n4154) );
  NOR2_X1 U4155 ( .A1(n2459), .A2(n2453), .ZN(n4028) );
  NOR2_X1 U4156 ( .A1(n4027), .A2(n4155), .ZN(n4151) );
  INV_X1 U4157 ( .A(n4029), .ZN(n4155) );
  NAND2_X1 U4158 ( .A1(n4156), .A2(n4157), .ZN(n4029) );
  NAND2_X1 U4159 ( .A1(n4036), .A2(n4158), .ZN(n4157) );
  INV_X1 U4160 ( .A(n4159), .ZN(n4158) );
  NOR2_X1 U4161 ( .A1(n4035), .A2(n4033), .ZN(n4159) );
  NOR2_X1 U4162 ( .A1(n2459), .A2(n2254), .ZN(n4036) );
  NAND2_X1 U4163 ( .A1(n4033), .A2(n4035), .ZN(n4156) );
  NAND2_X1 U4164 ( .A1(n4160), .A2(n4161), .ZN(n4035) );
  INV_X1 U4165 ( .A(n4162), .ZN(n4161) );
  NOR2_X1 U4166 ( .A1(n4064), .A2(n4163), .ZN(n4162) );
  NOR2_X1 U4167 ( .A1(n4063), .A2(n4065), .ZN(n4163) );
  NAND2_X1 U4168 ( .A1(b_2_), .A2(a_12_), .ZN(n4064) );
  NAND2_X1 U4169 ( .A1(n4063), .A2(n4065), .ZN(n4160) );
  NAND2_X1 U4170 ( .A1(n4164), .A2(n4165), .ZN(n4065) );
  NAND2_X1 U4171 ( .A1(n4059), .A2(n4166), .ZN(n4165) );
  INV_X1 U4172 ( .A(n4167), .ZN(n4166) );
  NOR2_X1 U4173 ( .A1(n4060), .A2(n4061), .ZN(n4167) );
  NOR2_X1 U4174 ( .A1(n2459), .A2(n2223), .ZN(n4059) );
  NAND2_X1 U4175 ( .A1(n4061), .A2(n4060), .ZN(n4164) );
  NAND2_X1 U4176 ( .A1(n4168), .A2(n4169), .ZN(n4060) );
  NAND2_X1 U4177 ( .A1(b_0_), .A2(n4170), .ZN(n4169) );
  NAND2_X1 U4178 ( .A1(n2202), .A2(n4171), .ZN(n4170) );
  NAND2_X1 U4179 ( .A1(a_15_), .A2(n4057), .ZN(n4171) );
  NAND2_X1 U4180 ( .A1(a_15_), .A2(n4172), .ZN(n2202) );
  NAND2_X1 U4181 ( .A1(b_1_), .A2(n4173), .ZN(n4168) );
  NAND2_X1 U4182 ( .A1(n2205), .A2(n4174), .ZN(n4173) );
  NAND2_X1 U4183 ( .A1(a_14_), .A2(n4101), .ZN(n4174) );
  NAND2_X1 U4184 ( .A1(a_14_), .A2(n2194), .ZN(n2205) );
  NOR3_X1 U4185 ( .A1(n2459), .A2(n4057), .A3(n2598), .ZN(n4061) );
  XNOR2_X1 U4186 ( .A(n4175), .B(n4176), .ZN(n4063) );
  XNOR2_X1 U4187 ( .A(n4177), .B(n4178), .ZN(n4176) );
  NAND2_X1 U4188 ( .A1(a_14_), .A2(b_0_), .ZN(n4175) );
  XNOR2_X1 U4189 ( .A(n4179), .B(n4180), .ZN(n4033) );
  NAND2_X1 U4190 ( .A1(n4181), .A2(n4182), .ZN(n4179) );
  NAND2_X1 U4191 ( .A1(n4183), .A2(n4184), .ZN(n4182) );
  NAND2_X1 U4192 ( .A1(b_1_), .A2(a_12_), .ZN(n4183) );
  XNOR2_X1 U4193 ( .A(n4185), .B(n4186), .ZN(n4027) );
  XOR2_X1 U4194 ( .A(n4187), .B(n4188), .Z(n4186) );
  NAND2_X1 U4195 ( .A1(b_1_), .A2(a_11_), .ZN(n4185) );
  XNOR2_X1 U4196 ( .A(n4189), .B(n4190), .ZN(n4067) );
  XNOR2_X1 U4197 ( .A(n4191), .B(n4192), .ZN(n4190) );
  NAND2_X1 U4198 ( .A1(b_1_), .A2(a_10_), .ZN(n4189) );
  XNOR2_X1 U4199 ( .A(n4193), .B(n4194), .ZN(n4014) );
  NOR2_X1 U4200 ( .A1(n2283), .A2(n4057), .ZN(n4194) );
  XOR2_X1 U4201 ( .A(n4195), .B(n4196), .Z(n4193) );
  XNOR2_X1 U4202 ( .A(n4197), .B(n4198), .ZN(n4071) );
  XNOR2_X1 U4203 ( .A(n4199), .B(n4200), .ZN(n4198) );
  NAND2_X1 U4204 ( .A1(b_1_), .A2(a_8_), .ZN(n4197) );
  XNOR2_X1 U4205 ( .A(n4201), .B(n4202), .ZN(n4075) );
  NOR2_X1 U4206 ( .A1(n2312), .A2(n4057), .ZN(n4202) );
  XOR2_X1 U4207 ( .A(n4203), .B(n4204), .Z(n4201) );
  XNOR2_X1 U4208 ( .A(n4205), .B(n4206), .ZN(n4079) );
  XNOR2_X1 U4209 ( .A(n4207), .B(n4208), .ZN(n4206) );
  NAND2_X1 U4210 ( .A1(b_1_), .A2(a_6_), .ZN(n4205) );
  XNOR2_X1 U4211 ( .A(n4209), .B(n4210), .ZN(n3995) );
  NOR2_X1 U4212 ( .A1(n2341), .A2(n4057), .ZN(n4210) );
  XOR2_X1 U4213 ( .A(n4211), .B(n4212), .Z(n4209) );
  XNOR2_X1 U4214 ( .A(n4213), .B(n4214), .ZN(n3987) );
  XNOR2_X1 U4215 ( .A(n4215), .B(n4216), .ZN(n4214) );
  NAND2_X1 U4216 ( .A1(b_1_), .A2(a_4_), .ZN(n4213) );
  XNOR2_X1 U4217 ( .A(n4217), .B(n4218), .ZN(n4086) );
  XNOR2_X1 U4218 ( .A(n4110), .B(n4109), .ZN(n4218) );
  NOR2_X1 U4219 ( .A1(n4219), .A2(n4220), .ZN(n4109) );
  NOR3_X1 U4220 ( .A1(n2376), .A2(n4221), .A3(n4057), .ZN(n4220) );
  INV_X1 U4221 ( .A(n4222), .ZN(n4221) );
  NAND2_X1 U4222 ( .A1(n4122), .A2(n4121), .ZN(n4222) );
  NOR2_X1 U4223 ( .A1(n4121), .A2(n4122), .ZN(n4219) );
  NOR2_X1 U4224 ( .A1(n4223), .A2(n4224), .ZN(n4122) );
  INV_X1 U4225 ( .A(n4225), .ZN(n4224) );
  NAND3_X1 U4226 ( .A1(a_4_), .A2(n4226), .A3(b_1_), .ZN(n4225) );
  NAND2_X1 U4227 ( .A1(n4216), .A2(n4215), .ZN(n4226) );
  NOR2_X1 U4228 ( .A1(n4215), .A2(n4216), .ZN(n4223) );
  NOR2_X1 U4229 ( .A1(n4227), .A2(n4228), .ZN(n4216) );
  NOR3_X1 U4230 ( .A1(n2341), .A2(n4229), .A3(n4057), .ZN(n4228) );
  INV_X1 U4231 ( .A(n4230), .ZN(n4229) );
  NAND2_X1 U4232 ( .A1(n4212), .A2(n4211), .ZN(n4230) );
  NOR2_X1 U4233 ( .A1(n4211), .A2(n4212), .ZN(n4227) );
  NOR2_X1 U4234 ( .A1(n4231), .A2(n4232), .ZN(n4212) );
  INV_X1 U4235 ( .A(n4233), .ZN(n4232) );
  NAND3_X1 U4236 ( .A1(a_6_), .A2(n4234), .A3(b_1_), .ZN(n4233) );
  NAND2_X1 U4237 ( .A1(n4208), .A2(n4207), .ZN(n4234) );
  NOR2_X1 U4238 ( .A1(n4207), .A2(n4208), .ZN(n4231) );
  NOR2_X1 U4239 ( .A1(n4235), .A2(n4236), .ZN(n4208) );
  NOR3_X1 U4240 ( .A1(n2312), .A2(n4237), .A3(n4057), .ZN(n4236) );
  INV_X1 U4241 ( .A(n4238), .ZN(n4237) );
  NAND2_X1 U4242 ( .A1(n4204), .A2(n4203), .ZN(n4238) );
  NOR2_X1 U4243 ( .A1(n4203), .A2(n4204), .ZN(n4235) );
  NOR2_X1 U4244 ( .A1(n4239), .A2(n4240), .ZN(n4204) );
  INV_X1 U4245 ( .A(n4241), .ZN(n4240) );
  NAND3_X1 U4246 ( .A1(a_8_), .A2(n4242), .A3(b_1_), .ZN(n4241) );
  NAND2_X1 U4247 ( .A1(n4200), .A2(n4199), .ZN(n4242) );
  NOR2_X1 U4248 ( .A1(n4199), .A2(n4200), .ZN(n4239) );
  NOR2_X1 U4249 ( .A1(n4243), .A2(n4244), .ZN(n4200) );
  NOR3_X1 U4250 ( .A1(n2283), .A2(n4245), .A3(n4057), .ZN(n4244) );
  INV_X1 U4251 ( .A(n4246), .ZN(n4245) );
  NAND2_X1 U4252 ( .A1(n4196), .A2(n4195), .ZN(n4246) );
  NOR2_X1 U4253 ( .A1(n4195), .A2(n4196), .ZN(n4243) );
  NOR2_X1 U4254 ( .A1(n4247), .A2(n4248), .ZN(n4196) );
  NOR3_X1 U4255 ( .A1(n2453), .A2(n4249), .A3(n4057), .ZN(n4248) );
  NOR2_X1 U4256 ( .A1(n4192), .A2(n4191), .ZN(n4249) );
  INV_X1 U4257 ( .A(n4250), .ZN(n4247) );
  NAND2_X1 U4258 ( .A1(n4191), .A2(n4192), .ZN(n4250) );
  NAND2_X1 U4259 ( .A1(n4251), .A2(n4252), .ZN(n4192) );
  NAND3_X1 U4260 ( .A1(a_11_), .A2(n4253), .A3(b_1_), .ZN(n4252) );
  NAND2_X1 U4261 ( .A1(n4188), .A2(n4254), .ZN(n4253) );
  INV_X1 U4262 ( .A(n4255), .ZN(n4188) );
  NAND2_X1 U4263 ( .A1(n4187), .A2(n4255), .ZN(n4251) );
  NAND2_X1 U4264 ( .A1(n4181), .A2(n4256), .ZN(n4255) );
  NAND2_X1 U4265 ( .A1(n4257), .A2(n4180), .ZN(n4256) );
  NAND2_X1 U4266 ( .A1(n4178), .A2(n4258), .ZN(n4180) );
  NAND3_X1 U4267 ( .A1(a_14_), .A2(b_0_), .A3(n4177), .ZN(n4258) );
  NOR2_X1 U4268 ( .A1(n4057), .A2(n2223), .ZN(n4177) );
  NAND3_X1 U4269 ( .A1(b_1_), .A2(b_0_), .A3(n2450), .ZN(n4178) );
  NAND2_X1 U4270 ( .A1(n4184), .A2(n2238), .ZN(n4257) );
  INV_X1 U4271 ( .A(n4259), .ZN(n4184) );
  NAND3_X1 U4272 ( .A1(b_1_), .A2(a_12_), .A3(n4259), .ZN(n4181) );
  NOR2_X1 U4273 ( .A1(n2223), .A2(n4101), .ZN(n4259) );
  INV_X1 U4274 ( .A(n4254), .ZN(n4187) );
  NAND2_X1 U4275 ( .A1(a_12_), .A2(b_0_), .ZN(n4254) );
  NOR2_X1 U4276 ( .A1(n2254), .A2(n4101), .ZN(n4191) );
  NAND2_X1 U4277 ( .A1(a_10_), .A2(b_0_), .ZN(n4195) );
  NAND2_X1 U4278 ( .A1(a_9_), .A2(b_0_), .ZN(n4199) );
  NAND2_X1 U4279 ( .A1(a_8_), .A2(b_0_), .ZN(n4203) );
  NAND2_X1 U4280 ( .A1(a_7_), .A2(b_0_), .ZN(n4207) );
  NAND2_X1 U4281 ( .A1(a_6_), .A2(b_0_), .ZN(n4211) );
  NAND2_X1 U4282 ( .A1(a_5_), .A2(b_0_), .ZN(n4215) );
  NAND2_X1 U4283 ( .A1(a_4_), .A2(b_0_), .ZN(n4121) );
  NAND2_X1 U4284 ( .A1(a_3_), .A2(b_0_), .ZN(n4110) );
  NAND2_X1 U4285 ( .A1(b_1_), .A2(a_2_), .ZN(n4217) );
  NAND2_X1 U4286 ( .A1(n4260), .A2(n4261), .ZN(n2195) );
  NAND2_X1 U4287 ( .A1(n4262), .A2(n2423), .ZN(n4261) );
  NAND2_X1 U4288 ( .A1(b_0_), .A2(n2420), .ZN(n2423) );
  INV_X1 U4289 ( .A(a_0_), .ZN(n2420) );
  NAND2_X1 U4290 ( .A1(n4263), .A2(n4264), .ZN(n4262) );
  NAND2_X1 U4291 ( .A1(a_1_), .A2(n4057), .ZN(n4264) );
  INV_X1 U4292 ( .A(b_1_), .ZN(n4057) );
  NAND3_X1 U4293 ( .A1(n4265), .A2(n4266), .A3(n4267), .ZN(n4263) );
  NAND2_X1 U4294 ( .A1(b_2_), .A2(n2460), .ZN(n4267) );
  INV_X1 U4295 ( .A(a_2_), .ZN(n2460) );
  NAND3_X1 U4296 ( .A1(n4268), .A2(n4269), .A3(n4270), .ZN(n4266) );
  NAND2_X1 U4297 ( .A1(a_3_), .A2(n2378), .ZN(n4270) );
  INV_X1 U4298 ( .A(b_3_), .ZN(n2378) );
  NAND3_X1 U4299 ( .A1(n4271), .A2(n4272), .A3(n4273), .ZN(n4269) );
  NAND2_X1 U4300 ( .A1(b_4_), .A2(n2457), .ZN(n4273) );
  INV_X1 U4301 ( .A(a_4_), .ZN(n2457) );
  NAND3_X1 U4302 ( .A1(n4274), .A2(n4275), .A3(n4276), .ZN(n4272) );
  NAND2_X1 U4303 ( .A1(a_5_), .A2(n2343), .ZN(n4276) );
  INV_X1 U4304 ( .A(b_5_), .ZN(n2343) );
  NAND3_X1 U4305 ( .A1(n4277), .A2(n4278), .A3(n4279), .ZN(n4275) );
  NAND2_X1 U4306 ( .A1(b_6_), .A2(n2455), .ZN(n4279) );
  INV_X1 U4307 ( .A(a_6_), .ZN(n2455) );
  NAND3_X1 U4308 ( .A1(n4280), .A2(n4281), .A3(n4282), .ZN(n4278) );
  NAND2_X1 U4309 ( .A1(a_7_), .A2(n2314), .ZN(n4282) );
  INV_X1 U4310 ( .A(b_7_), .ZN(n2314) );
  NAND3_X1 U4311 ( .A1(n4283), .A2(n4284), .A3(n4285), .ZN(n4281) );
  NAND2_X1 U4312 ( .A1(b_8_), .A2(n2681), .ZN(n4285) );
  INV_X1 U4313 ( .A(a_8_), .ZN(n2681) );
  NAND3_X1 U4314 ( .A1(n4286), .A2(n4287), .A3(n4288), .ZN(n4284) );
  NAND2_X1 U4315 ( .A1(a_9_), .A2(n2285), .ZN(n4288) );
  INV_X1 U4316 ( .A(b_9_), .ZN(n2285) );
  NAND3_X1 U4317 ( .A1(n4289), .A2(n4290), .A3(n4291), .ZN(n4287) );
  NAND2_X1 U4318 ( .A1(b_9_), .A2(n2283), .ZN(n4291) );
  INV_X1 U4319 ( .A(a_9_), .ZN(n2283) );
  NAND3_X1 U4320 ( .A1(n4292), .A2(n4293), .A3(n4294), .ZN(n4290) );
  NAND2_X1 U4321 ( .A1(a_11_), .A2(n2256), .ZN(n4294) );
  INV_X1 U4322 ( .A(b_11_), .ZN(n2256) );
  NAND3_X1 U4323 ( .A1(n4295), .A2(n4296), .A3(n4297), .ZN(n4293) );
  NAND2_X1 U4324 ( .A1(b_12_), .A2(n2238), .ZN(n4297) );
  INV_X1 U4325 ( .A(a_12_), .ZN(n2238) );
  NAND3_X1 U4326 ( .A1(n4298), .A2(n4299), .A3(n4300), .ZN(n4296) );
  NAND2_X1 U4327 ( .A1(a_13_), .A2(n2225), .ZN(n4300) );
  INV_X1 U4328 ( .A(b_13_), .ZN(n2225) );
  NAND4_X1 U4329 ( .A1(n4301), .A2(n4302), .A3(n4303), .A4(n2597), .ZN(n4299)
         );
  INV_X1 U4330 ( .A(n2449), .ZN(n2597) );
  NOR2_X1 U4331 ( .A1(n2192), .A2(n2207), .ZN(n2449) );
  INV_X1 U4332 ( .A(b_14_), .ZN(n2207) );
  NAND2_X1 U4333 ( .A1(n2203), .A2(n4172), .ZN(n4303) );
  NAND2_X1 U4334 ( .A1(a_15_), .A2(n2192), .ZN(n2203) );
  INV_X1 U4335 ( .A(b_15_), .ZN(n2192) );
  NAND2_X1 U4336 ( .A1(b_14_), .A2(n2598), .ZN(n4302) );
  INV_X1 U4337 ( .A(n2450), .ZN(n2598) );
  INV_X1 U4338 ( .A(a_15_), .ZN(n2194) );
  INV_X1 U4339 ( .A(a_14_), .ZN(n4172) );
  NAND2_X1 U4340 ( .A1(b_13_), .A2(n2223), .ZN(n4301) );
  INV_X1 U4341 ( .A(a_13_), .ZN(n2223) );
  NAND2_X1 U4342 ( .A1(a_12_), .A2(n2451), .ZN(n4298) );
  INV_X1 U4343 ( .A(b_12_), .ZN(n2451) );
  NAND2_X1 U4344 ( .A1(b_11_), .A2(n2254), .ZN(n4295) );
  INV_X1 U4345 ( .A(a_11_), .ZN(n2254) );
  NAND2_X1 U4346 ( .A1(a_10_), .A2(n2452), .ZN(n4292) );
  INV_X1 U4347 ( .A(b_10_), .ZN(n2452) );
  NAND2_X1 U4348 ( .A1(b_10_), .A2(n2453), .ZN(n4289) );
  INV_X1 U4349 ( .A(a_10_), .ZN(n2453) );
  NAND2_X1 U4350 ( .A1(a_8_), .A2(n3206), .ZN(n4286) );
  INV_X1 U4351 ( .A(b_8_), .ZN(n3206) );
  NAND2_X1 U4352 ( .A1(b_7_), .A2(n2312), .ZN(n4283) );
  INV_X1 U4353 ( .A(a_7_), .ZN(n2312) );
  NAND2_X1 U4354 ( .A1(a_6_), .A2(n2454), .ZN(n4280) );
  INV_X1 U4355 ( .A(b_6_), .ZN(n2454) );
  NAND2_X1 U4356 ( .A1(b_5_), .A2(n2341), .ZN(n4277) );
  INV_X1 U4357 ( .A(a_5_), .ZN(n2341) );
  NAND2_X1 U4358 ( .A1(a_4_), .A2(n2456), .ZN(n4274) );
  INV_X1 U4359 ( .A(b_4_), .ZN(n2456) );
  NAND2_X1 U4360 ( .A1(b_3_), .A2(n2376), .ZN(n4271) );
  INV_X1 U4361 ( .A(a_3_), .ZN(n2376) );
  NAND2_X1 U4362 ( .A1(a_2_), .A2(n2459), .ZN(n4268) );
  INV_X1 U4363 ( .A(b_2_), .ZN(n2459) );
  NAND2_X1 U4364 ( .A1(b_1_), .A2(n2647), .ZN(n4265) );
  INV_X1 U4365 ( .A(a_1_), .ZN(n2647) );
  NAND2_X1 U4366 ( .A1(a_0_), .A2(n4101), .ZN(n4260) );
  INV_X1 U4367 ( .A(b_0_), .ZN(n4101) );
endmodule

