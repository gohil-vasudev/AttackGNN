module locked_c1355 (  G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,  G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT  );
  input  G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n602_, new_n603_, new_n604_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n615_, new_n616_, new_n617_, new_n618_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_, new_n647_, new_n648_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n794_, new_n795_, new_n796_, new_n797_, new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n831_, new_n832_, new_n833_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_;
  NAND2_X1 g000 ( .A1(G141GAT), .A2(KEYINPUT2), .ZN(new_n138_) );
  INV_X1 g001 ( .A(G141GAT), .ZN(new_n139_) );
  INV_X1 g002 ( .A(KEYINPUT2), .ZN(new_n140_) );
  NAND2_X1 g003 ( .A1(new_n139_), .A2(new_n140_), .ZN(new_n141_) );
  NAND2_X1 g004 ( .A1(new_n141_), .A2(new_n138_), .ZN(new_n142_) );
  NAND2_X1 g005 ( .A1(G155GAT), .A2(KEYINPUT3), .ZN(new_n143_) );
  INV_X1 g006 ( .A(G155GAT), .ZN(new_n144_) );
  INV_X1 g007 ( .A(KEYINPUT3), .ZN(new_n145_) );
  NAND2_X1 g008 ( .A1(new_n144_), .A2(new_n145_), .ZN(new_n146_) );
  NAND2_X1 g009 ( .A1(new_n146_), .A2(new_n143_), .ZN(new_n147_) );
  NAND2_X1 g010 ( .A1(new_n142_), .A2(new_n147_), .ZN(new_n148_) );
  NAND4_X1 g011 ( .A1(new_n141_), .A2(new_n146_), .A3(new_n138_), .A4(new_n143_), .ZN(new_n149_) );
  NAND2_X1 g012 ( .A1(new_n148_), .A2(new_n149_), .ZN(new_n150_) );
  INV_X1 g013 ( .A(new_n150_), .ZN(new_n151_) );
  INV_X1 g014 ( .A(KEYINPUT1), .ZN(new_n152_) );
  NAND2_X1 g015 ( .A1(new_n152_), .A2(G57GAT), .ZN(new_n153_) );
  INV_X1 g016 ( .A(G57GAT), .ZN(new_n154_) );
  NAND2_X1 g017 ( .A1(new_n154_), .A2(KEYINPUT1), .ZN(new_n155_) );
  NAND2_X1 g018 ( .A1(new_n153_), .A2(new_n155_), .ZN(new_n156_) );
  NAND2_X1 g019 ( .A1(G225GAT), .A2(G233GAT), .ZN(new_n157_) );
  NAND2_X1 g020 ( .A1(new_n156_), .A2(new_n157_), .ZN(new_n158_) );
  NAND4_X1 g021 ( .A1(new_n153_), .A2(new_n155_), .A3(G225GAT), .A4(G233GAT), .ZN(new_n159_) );
  NAND2_X1 g022 ( .A1(new_n158_), .A2(new_n159_), .ZN(new_n160_) );
  NAND2_X1 g023 ( .A1(new_n151_), .A2(new_n160_), .ZN(new_n161_) );
  NAND3_X1 g024 ( .A1(new_n150_), .A2(new_n158_), .A3(new_n159_), .ZN(new_n162_) );
  NAND2_X1 g025 ( .A1(new_n161_), .A2(new_n162_), .ZN(new_n163_) );
  INV_X1 g026 ( .A(G1GAT), .ZN(new_n164_) );
  INV_X1 g027 ( .A(G127GAT), .ZN(new_n165_) );
  NAND2_X1 g028 ( .A1(new_n165_), .A2(G120GAT), .ZN(new_n166_) );
  INV_X1 g029 ( .A(G120GAT), .ZN(new_n167_) );
  NAND2_X1 g030 ( .A1(new_n167_), .A2(G127GAT), .ZN(new_n168_) );
  NAND2_X1 g031 ( .A1(new_n166_), .A2(new_n168_), .ZN(new_n169_) );
  NAND2_X1 g032 ( .A1(G113GAT), .A2(KEYINPUT0), .ZN(new_n170_) );
  INV_X1 g033 ( .A(G113GAT), .ZN(new_n171_) );
  INV_X1 g034 ( .A(KEYINPUT0), .ZN(new_n172_) );
  NAND2_X1 g035 ( .A1(new_n171_), .A2(new_n172_), .ZN(new_n173_) );
  NAND2_X1 g036 ( .A1(new_n173_), .A2(new_n170_), .ZN(new_n174_) );
  NAND2_X1 g037 ( .A1(new_n169_), .A2(new_n174_), .ZN(new_n175_) );
  NAND4_X1 g038 ( .A1(new_n173_), .A2(new_n166_), .A3(new_n168_), .A4(new_n170_), .ZN(new_n176_) );
  NAND2_X1 g039 ( .A1(new_n175_), .A2(new_n176_), .ZN(new_n177_) );
  NAND2_X1 g040 ( .A1(new_n177_), .A2(new_n164_), .ZN(new_n178_) );
  INV_X1 g041 ( .A(new_n177_), .ZN(new_n179_) );
  NAND2_X1 g042 ( .A1(new_n179_), .A2(G1GAT), .ZN(new_n180_) );
  NAND2_X1 g043 ( .A1(new_n180_), .A2(new_n178_), .ZN(new_n181_) );
  NAND2_X1 g044 ( .A1(new_n163_), .A2(new_n181_), .ZN(new_n182_) );
  NAND4_X1 g045 ( .A1(new_n161_), .A2(new_n180_), .A3(new_n162_), .A4(new_n178_), .ZN(new_n183_) );
  NAND2_X1 g046 ( .A1(new_n182_), .A2(new_n183_), .ZN(new_n184_) );
  NAND2_X1 g047 ( .A1(G29GAT), .A2(G134GAT), .ZN(new_n185_) );
  INV_X1 g048 ( .A(new_n185_), .ZN(new_n186_) );
  NOR2_X1 g049 ( .A1(G29GAT), .A2(G134GAT), .ZN(new_n187_) );
  NOR2_X1 g050 ( .A1(new_n186_), .A2(new_n187_), .ZN(new_n188_) );
  INV_X1 g051 ( .A(new_n188_), .ZN(new_n189_) );
  NAND2_X1 g052 ( .A1(new_n184_), .A2(new_n189_), .ZN(new_n190_) );
  NAND3_X1 g053 ( .A1(new_n182_), .A2(new_n183_), .A3(new_n188_), .ZN(new_n191_) );
  NAND2_X1 g054 ( .A1(new_n190_), .A2(new_n191_), .ZN(new_n192_) );
  NAND2_X1 g055 ( .A1(G85GAT), .A2(G162GAT), .ZN(new_n193_) );
  INV_X1 g056 ( .A(new_n193_), .ZN(new_n194_) );
  NOR2_X1 g057 ( .A1(G85GAT), .A2(G162GAT), .ZN(new_n195_) );
  NOR2_X1 g058 ( .A1(new_n194_), .A2(new_n195_), .ZN(new_n196_) );
  INV_X1 g059 ( .A(new_n196_), .ZN(new_n197_) );
  NAND2_X1 g060 ( .A1(new_n192_), .A2(new_n197_), .ZN(new_n198_) );
  NAND3_X1 g061 ( .A1(new_n190_), .A2(new_n191_), .A3(new_n196_), .ZN(new_n199_) );
  NAND2_X1 g062 ( .A1(new_n198_), .A2(new_n199_), .ZN(new_n200_) );
  NAND2_X1 g063 ( .A1(KEYINPUT5), .A2(KEYINPUT4), .ZN(new_n201_) );
  INV_X1 g064 ( .A(KEYINPUT5), .ZN(new_n202_) );
  INV_X1 g065 ( .A(KEYINPUT4), .ZN(new_n203_) );
  NAND2_X1 g066 ( .A1(new_n202_), .A2(new_n203_), .ZN(new_n204_) );
  NAND2_X1 g067 ( .A1(new_n204_), .A2(new_n201_), .ZN(new_n205_) );
  NAND2_X1 g068 ( .A1(G148GAT), .A2(KEYINPUT6), .ZN(new_n206_) );
  INV_X1 g069 ( .A(G148GAT), .ZN(new_n207_) );
  INV_X1 g070 ( .A(KEYINPUT6), .ZN(new_n208_) );
  NAND2_X1 g071 ( .A1(new_n207_), .A2(new_n208_), .ZN(new_n209_) );
  NAND2_X1 g072 ( .A1(new_n209_), .A2(new_n206_), .ZN(new_n210_) );
  NAND2_X1 g073 ( .A1(new_n205_), .A2(new_n210_), .ZN(new_n211_) );
  NAND4_X1 g074 ( .A1(new_n204_), .A2(new_n209_), .A3(new_n201_), .A4(new_n206_), .ZN(new_n212_) );
  NAND3_X1 g075 ( .A1(new_n200_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_) );
  NAND2_X1 g076 ( .A1(new_n211_), .A2(new_n212_), .ZN(new_n214_) );
  NAND3_X1 g077 ( .A1(new_n198_), .A2(new_n199_), .A3(new_n214_), .ZN(new_n215_) );
  NAND2_X1 g078 ( .A1(new_n213_), .A2(new_n215_), .ZN(new_n216_) );
  INV_X1 g079 ( .A(new_n216_), .ZN(new_n217_) );
  INV_X1 g080 ( .A(KEYINPUT25), .ZN(new_n218_) );
  INV_X1 g081 ( .A(G197GAT), .ZN(new_n219_) );
  INV_X1 g082 ( .A(G218GAT), .ZN(new_n220_) );
  NAND2_X1 g083 ( .A1(new_n220_), .A2(G211GAT), .ZN(new_n221_) );
  INV_X1 g084 ( .A(G211GAT), .ZN(new_n222_) );
  NAND2_X1 g085 ( .A1(new_n222_), .A2(G218GAT), .ZN(new_n223_) );
  NAND2_X1 g086 ( .A1(new_n221_), .A2(new_n223_), .ZN(new_n224_) );
  NAND2_X1 g087 ( .A1(G204GAT), .A2(KEYINPUT21), .ZN(new_n225_) );
  INV_X1 g088 ( .A(G204GAT), .ZN(new_n226_) );
  INV_X1 g089 ( .A(KEYINPUT21), .ZN(new_n227_) );
  NAND2_X1 g090 ( .A1(new_n226_), .A2(new_n227_), .ZN(new_n228_) );
  NAND2_X1 g091 ( .A1(new_n228_), .A2(new_n225_), .ZN(new_n229_) );
  NAND2_X1 g092 ( .A1(new_n224_), .A2(new_n229_), .ZN(new_n230_) );
  NAND4_X1 g093 ( .A1(new_n228_), .A2(new_n221_), .A3(new_n223_), .A4(new_n225_), .ZN(new_n231_) );
  NAND2_X1 g094 ( .A1(new_n230_), .A2(new_n231_), .ZN(new_n232_) );
  NAND2_X1 g095 ( .A1(new_n232_), .A2(new_n219_), .ZN(new_n233_) );
  NAND3_X1 g096 ( .A1(new_n230_), .A2(G197GAT), .A3(new_n231_), .ZN(new_n234_) );
  NAND2_X1 g097 ( .A1(new_n233_), .A2(new_n234_), .ZN(new_n235_) );
  INV_X1 g098 ( .A(new_n235_), .ZN(new_n236_) );
  NAND2_X1 g099 ( .A1(new_n236_), .A2(new_n150_), .ZN(new_n237_) );
  NAND2_X1 g100 ( .A1(new_n235_), .A2(new_n151_), .ZN(new_n238_) );
  NAND2_X1 g101 ( .A1(new_n237_), .A2(new_n238_), .ZN(new_n239_) );
  INV_X1 g102 ( .A(KEYINPUT23), .ZN(new_n240_) );
  NAND2_X1 g103 ( .A1(new_n240_), .A2(KEYINPUT24), .ZN(new_n241_) );
  INV_X1 g104 ( .A(KEYINPUT24), .ZN(new_n242_) );
  NAND2_X1 g105 ( .A1(new_n242_), .A2(KEYINPUT23), .ZN(new_n243_) );
  NAND2_X1 g106 ( .A1(new_n241_), .A2(new_n243_), .ZN(new_n244_) );
  NAND2_X1 g107 ( .A1(G22GAT), .A2(KEYINPUT22), .ZN(new_n245_) );
  INV_X1 g108 ( .A(G22GAT), .ZN(new_n246_) );
  INV_X1 g109 ( .A(KEYINPUT22), .ZN(new_n247_) );
  NAND2_X1 g110 ( .A1(new_n246_), .A2(new_n247_), .ZN(new_n248_) );
  NAND2_X1 g111 ( .A1(new_n248_), .A2(new_n245_), .ZN(new_n249_) );
  NAND2_X1 g112 ( .A1(new_n244_), .A2(new_n249_), .ZN(new_n250_) );
  NAND4_X1 g113 ( .A1(new_n248_), .A2(new_n241_), .A3(new_n243_), .A4(new_n245_), .ZN(new_n251_) );
  NAND2_X1 g114 ( .A1(new_n250_), .A2(new_n251_), .ZN(new_n252_) );
  INV_X1 g115 ( .A(G78GAT), .ZN(new_n253_) );
  INV_X1 g116 ( .A(G106GAT), .ZN(new_n254_) );
  NAND2_X1 g117 ( .A1(new_n253_), .A2(new_n254_), .ZN(new_n255_) );
  NAND2_X1 g118 ( .A1(G78GAT), .A2(G106GAT), .ZN(new_n256_) );
  NAND2_X1 g119 ( .A1(new_n255_), .A2(new_n256_), .ZN(new_n257_) );
  NAND2_X1 g120 ( .A1(new_n257_), .A2(G148GAT), .ZN(new_n258_) );
  NAND3_X1 g121 ( .A1(new_n255_), .A2(new_n207_), .A3(new_n256_), .ZN(new_n259_) );
  NAND2_X1 g122 ( .A1(new_n258_), .A2(new_n259_), .ZN(new_n260_) );
  NAND2_X1 g123 ( .A1(new_n252_), .A2(new_n260_), .ZN(new_n261_) );
  NAND4_X1 g124 ( .A1(new_n250_), .A2(new_n258_), .A3(new_n251_), .A4(new_n259_), .ZN(new_n262_) );
  NAND3_X1 g125 ( .A1(new_n239_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_) );
  NAND2_X1 g126 ( .A1(new_n261_), .A2(new_n262_), .ZN(new_n264_) );
  NAND3_X1 g127 ( .A1(new_n237_), .A2(new_n238_), .A3(new_n264_), .ZN(new_n265_) );
  NAND2_X1 g128 ( .A1(new_n263_), .A2(new_n265_), .ZN(new_n266_) );
  INV_X1 g129 ( .A(G50GAT), .ZN(new_n267_) );
  NOR2_X1 g130 ( .A1(new_n267_), .A2(G162GAT), .ZN(new_n268_) );
  INV_X1 g131 ( .A(G162GAT), .ZN(new_n269_) );
  NOR2_X1 g132 ( .A1(new_n269_), .A2(G50GAT), .ZN(new_n270_) );
  NOR2_X1 g133 ( .A1(new_n268_), .A2(new_n270_), .ZN(new_n271_) );
  NAND2_X1 g134 ( .A1(new_n266_), .A2(new_n271_), .ZN(new_n272_) );
  INV_X1 g135 ( .A(new_n271_), .ZN(new_n273_) );
  NAND3_X1 g136 ( .A1(new_n263_), .A2(new_n265_), .A3(new_n273_), .ZN(new_n274_) );
  NAND2_X1 g137 ( .A1(new_n272_), .A2(new_n274_), .ZN(new_n275_) );
  NAND3_X1 g138 ( .A1(new_n275_), .A2(G228GAT), .A3(G233GAT), .ZN(new_n276_) );
  NAND2_X1 g139 ( .A1(G228GAT), .A2(G233GAT), .ZN(new_n277_) );
  NAND3_X1 g140 ( .A1(new_n272_), .A2(new_n274_), .A3(new_n277_), .ZN(new_n278_) );
  NAND2_X1 g141 ( .A1(new_n276_), .A2(new_n278_), .ZN(new_n279_) );
  INV_X1 g142 ( .A(new_n279_), .ZN(new_n280_) );
  INV_X1 g143 ( .A(G15GAT), .ZN(new_n281_) );
  NAND2_X1 g144 ( .A1(new_n177_), .A2(new_n281_), .ZN(new_n282_) );
  NAND2_X1 g145 ( .A1(new_n179_), .A2(G15GAT), .ZN(new_n283_) );
  NAND2_X1 g146 ( .A1(new_n283_), .A2(new_n282_), .ZN(new_n284_) );
  NAND2_X1 g147 ( .A1(G227GAT), .A2(G233GAT), .ZN(new_n285_) );
  NAND2_X1 g148 ( .A1(new_n284_), .A2(new_n285_), .ZN(new_n286_) );
  NAND4_X1 g149 ( .A1(new_n283_), .A2(G227GAT), .A3(G233GAT), .A4(new_n282_), .ZN(new_n287_) );
  NAND2_X1 g150 ( .A1(G71GAT), .A2(KEYINPUT20), .ZN(new_n288_) );
  INV_X1 g151 ( .A(G71GAT), .ZN(new_n289_) );
  INV_X1 g152 ( .A(KEYINPUT20), .ZN(new_n290_) );
  NAND2_X1 g153 ( .A1(new_n289_), .A2(new_n290_), .ZN(new_n291_) );
  NAND2_X1 g154 ( .A1(new_n291_), .A2(new_n288_), .ZN(new_n292_) );
  NAND2_X1 g155 ( .A1(G176GAT), .A2(G183GAT), .ZN(new_n293_) );
  INV_X1 g156 ( .A(G176GAT), .ZN(new_n294_) );
  INV_X1 g157 ( .A(G183GAT), .ZN(new_n295_) );
  NAND2_X1 g158 ( .A1(new_n294_), .A2(new_n295_), .ZN(new_n296_) );
  NAND2_X1 g159 ( .A1(new_n296_), .A2(new_n293_), .ZN(new_n297_) );
  NAND2_X1 g160 ( .A1(new_n292_), .A2(new_n297_), .ZN(new_n298_) );
  NAND4_X1 g161 ( .A1(new_n291_), .A2(new_n296_), .A3(new_n288_), .A4(new_n293_), .ZN(new_n299_) );
  NAND4_X1 g162 ( .A1(new_n286_), .A2(new_n287_), .A3(new_n298_), .A4(new_n299_), .ZN(new_n300_) );
  NAND2_X1 g163 ( .A1(new_n286_), .A2(new_n287_), .ZN(new_n301_) );
  NAND2_X1 g164 ( .A1(new_n298_), .A2(new_n299_), .ZN(new_n302_) );
  NAND2_X1 g165 ( .A1(new_n301_), .A2(new_n302_), .ZN(new_n303_) );
  NAND2_X1 g166 ( .A1(new_n303_), .A2(new_n300_), .ZN(new_n304_) );
  NAND2_X1 g167 ( .A1(KEYINPUT18), .A2(KEYINPUT17), .ZN(new_n305_) );
  INV_X1 g168 ( .A(KEYINPUT18), .ZN(new_n306_) );
  INV_X1 g169 ( .A(KEYINPUT17), .ZN(new_n307_) );
  NAND2_X1 g170 ( .A1(new_n306_), .A2(new_n307_), .ZN(new_n308_) );
  NAND2_X1 g171 ( .A1(new_n308_), .A2(new_n305_), .ZN(new_n309_) );
  NAND2_X1 g172 ( .A1(G169GAT), .A2(KEYINPUT19), .ZN(new_n310_) );
  INV_X1 g173 ( .A(G169GAT), .ZN(new_n311_) );
  INV_X1 g174 ( .A(KEYINPUT19), .ZN(new_n312_) );
  NAND2_X1 g175 ( .A1(new_n311_), .A2(new_n312_), .ZN(new_n313_) );
  NAND2_X1 g176 ( .A1(new_n313_), .A2(new_n310_), .ZN(new_n314_) );
  NAND2_X1 g177 ( .A1(new_n309_), .A2(new_n314_), .ZN(new_n315_) );
  NAND4_X1 g178 ( .A1(new_n308_), .A2(new_n313_), .A3(new_n305_), .A4(new_n310_), .ZN(new_n316_) );
  NAND2_X1 g179 ( .A1(new_n315_), .A2(new_n316_), .ZN(new_n317_) );
  NAND2_X1 g180 ( .A1(G134GAT), .A2(G190GAT), .ZN(new_n318_) );
  INV_X1 g181 ( .A(G134GAT), .ZN(new_n319_) );
  INV_X1 g182 ( .A(G190GAT), .ZN(new_n320_) );
  NAND2_X1 g183 ( .A1(new_n319_), .A2(new_n320_), .ZN(new_n321_) );
  NAND2_X1 g184 ( .A1(new_n321_), .A2(new_n318_), .ZN(new_n322_) );
  NAND2_X1 g185 ( .A1(G43GAT), .A2(G99GAT), .ZN(new_n323_) );
  INV_X1 g186 ( .A(G43GAT), .ZN(new_n324_) );
  INV_X1 g187 ( .A(G99GAT), .ZN(new_n325_) );
  NAND2_X1 g188 ( .A1(new_n324_), .A2(new_n325_), .ZN(new_n326_) );
  NAND2_X1 g189 ( .A1(new_n326_), .A2(new_n323_), .ZN(new_n327_) );
  NAND2_X1 g190 ( .A1(new_n322_), .A2(new_n327_), .ZN(new_n328_) );
  NAND4_X1 g191 ( .A1(new_n321_), .A2(new_n326_), .A3(new_n318_), .A4(new_n323_), .ZN(new_n329_) );
  NAND2_X1 g192 ( .A1(new_n328_), .A2(new_n329_), .ZN(new_n330_) );
  NAND2_X1 g193 ( .A1(new_n317_), .A2(new_n330_), .ZN(new_n331_) );
  INV_X1 g194 ( .A(new_n317_), .ZN(new_n332_) );
  NAND3_X1 g195 ( .A1(new_n332_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n333_) );
  NAND2_X1 g196 ( .A1(new_n333_), .A2(new_n331_), .ZN(new_n334_) );
  NAND2_X1 g197 ( .A1(new_n304_), .A2(new_n334_), .ZN(new_n335_) );
  NAND4_X1 g198 ( .A1(new_n303_), .A2(new_n300_), .A3(new_n331_), .A4(new_n333_), .ZN(new_n336_) );
  NAND2_X1 g199 ( .A1(new_n335_), .A2(new_n336_), .ZN(new_n337_) );
  INV_X1 g200 ( .A(new_n337_), .ZN(new_n338_) );
  NAND2_X1 g201 ( .A1(G36GAT), .A2(G190GAT), .ZN(new_n339_) );
  INV_X1 g202 ( .A(new_n339_), .ZN(new_n340_) );
  NOR2_X1 g203 ( .A1(G36GAT), .A2(G190GAT), .ZN(new_n341_) );
  NOR2_X1 g204 ( .A1(new_n340_), .A2(new_n341_), .ZN(new_n342_) );
  NAND2_X1 g205 ( .A1(new_n236_), .A2(new_n342_), .ZN(new_n343_) );
  INV_X1 g206 ( .A(new_n342_), .ZN(new_n344_) );
  NAND2_X1 g207 ( .A1(new_n235_), .A2(new_n344_), .ZN(new_n345_) );
  NAND2_X1 g208 ( .A1(new_n343_), .A2(new_n345_), .ZN(new_n346_) );
  NAND2_X1 g209 ( .A1(G64GAT), .A2(G176GAT), .ZN(new_n347_) );
  INV_X1 g210 ( .A(new_n347_), .ZN(new_n348_) );
  NOR2_X1 g211 ( .A1(G64GAT), .A2(G176GAT), .ZN(new_n349_) );
  NOR2_X1 g212 ( .A1(new_n348_), .A2(new_n349_), .ZN(new_n350_) );
  INV_X1 g213 ( .A(new_n350_), .ZN(new_n351_) );
  NAND2_X1 g214 ( .A1(new_n351_), .A2(G92GAT), .ZN(new_n352_) );
  INV_X1 g215 ( .A(G92GAT), .ZN(new_n353_) );
  NAND2_X1 g216 ( .A1(new_n350_), .A2(new_n353_), .ZN(new_n354_) );
  NAND2_X1 g217 ( .A1(new_n352_), .A2(new_n354_), .ZN(new_n355_) );
  NAND2_X1 g218 ( .A1(G226GAT), .A2(G233GAT), .ZN(new_n356_) );
  NAND2_X1 g219 ( .A1(new_n355_), .A2(new_n356_), .ZN(new_n357_) );
  NAND4_X1 g220 ( .A1(new_n352_), .A2(G226GAT), .A3(G233GAT), .A4(new_n354_), .ZN(new_n358_) );
  NAND2_X1 g221 ( .A1(new_n357_), .A2(new_n358_), .ZN(new_n359_) );
  NAND2_X1 g222 ( .A1(G8GAT), .A2(G183GAT), .ZN(new_n360_) );
  INV_X1 g223 ( .A(new_n360_), .ZN(new_n361_) );
  NOR2_X1 g224 ( .A1(G8GAT), .A2(G183GAT), .ZN(new_n362_) );
  NOR2_X1 g225 ( .A1(new_n361_), .A2(new_n362_), .ZN(new_n363_) );
  NAND2_X1 g226 ( .A1(new_n359_), .A2(new_n363_), .ZN(new_n364_) );
  INV_X1 g227 ( .A(new_n363_), .ZN(new_n365_) );
  NAND3_X1 g228 ( .A1(new_n357_), .A2(new_n358_), .A3(new_n365_), .ZN(new_n366_) );
  NAND2_X1 g229 ( .A1(new_n364_), .A2(new_n366_), .ZN(new_n367_) );
  NAND2_X1 g230 ( .A1(new_n367_), .A2(new_n346_), .ZN(new_n368_) );
  NAND4_X1 g231 ( .A1(new_n364_), .A2(new_n343_), .A3(new_n345_), .A4(new_n366_), .ZN(new_n369_) );
  NAND2_X1 g232 ( .A1(new_n368_), .A2(new_n369_), .ZN(new_n370_) );
  NAND2_X1 g233 ( .A1(new_n370_), .A2(new_n317_), .ZN(new_n371_) );
  NAND3_X1 g234 ( .A1(new_n368_), .A2(new_n332_), .A3(new_n369_), .ZN(new_n372_) );
  NAND2_X1 g235 ( .A1(new_n371_), .A2(new_n372_), .ZN(new_n373_) );
  INV_X1 g236 ( .A(new_n373_), .ZN(new_n374_) );
  NAND2_X1 g237 ( .A1(new_n374_), .A2(new_n338_), .ZN(new_n375_) );
  NAND2_X1 g238 ( .A1(new_n280_), .A2(new_n375_), .ZN(new_n376_) );
  NAND2_X1 g239 ( .A1(new_n376_), .A2(new_n218_), .ZN(new_n377_) );
  NAND3_X1 g240 ( .A1(new_n280_), .A2(KEYINPUT25), .A3(new_n375_), .ZN(new_n378_) );
  NAND2_X1 g241 ( .A1(new_n377_), .A2(new_n378_), .ZN(new_n379_) );
  NAND2_X1 g242 ( .A1(new_n374_), .A2(KEYINPUT27), .ZN(new_n380_) );
  INV_X1 g243 ( .A(KEYINPUT27), .ZN(new_n381_) );
  NAND2_X1 g244 ( .A1(new_n373_), .A2(new_n381_), .ZN(new_n382_) );
  NAND2_X1 g245 ( .A1(new_n380_), .A2(new_n382_), .ZN(new_n383_) );
  INV_X1 g246 ( .A(KEYINPUT26), .ZN(new_n384_) );
  NAND2_X1 g247 ( .A1(new_n279_), .A2(new_n337_), .ZN(new_n385_) );
  NAND2_X1 g248 ( .A1(new_n385_), .A2(new_n384_), .ZN(new_n386_) );
  NAND3_X1 g249 ( .A1(new_n279_), .A2(KEYINPUT26), .A3(new_n337_), .ZN(new_n387_) );
  NAND2_X1 g250 ( .A1(new_n386_), .A2(new_n387_), .ZN(new_n388_) );
  NAND2_X1 g251 ( .A1(new_n388_), .A2(new_n383_), .ZN(new_n389_) );
  NAND2_X1 g252 ( .A1(new_n389_), .A2(new_n379_), .ZN(new_n390_) );
  NAND2_X1 g253 ( .A1(new_n390_), .A2(new_n216_), .ZN(new_n391_) );
  INV_X1 g254 ( .A(KEYINPUT28), .ZN(new_n392_) );
  NAND2_X1 g255 ( .A1(new_n279_), .A2(new_n392_), .ZN(new_n393_) );
  NAND2_X1 g256 ( .A1(new_n280_), .A2(KEYINPUT28), .ZN(new_n394_) );
  NAND2_X1 g257 ( .A1(new_n394_), .A2(new_n393_), .ZN(new_n395_) );
  INV_X1 g258 ( .A(new_n383_), .ZN(new_n396_) );
  NOR2_X1 g259 ( .A1(new_n396_), .A2(new_n216_), .ZN(new_n397_) );
  NAND3_X1 g260 ( .A1(new_n395_), .A2(new_n337_), .A3(new_n397_), .ZN(new_n398_) );
  NAND2_X1 g261 ( .A1(new_n391_), .A2(new_n398_), .ZN(new_n399_) );
  INV_X1 g262 ( .A(KEYINPUT16), .ZN(new_n400_) );
  INV_X1 g263 ( .A(KEYINPUT9), .ZN(new_n401_) );
  NAND2_X1 g264 ( .A1(KEYINPUT11), .A2(KEYINPUT10), .ZN(new_n402_) );
  INV_X1 g265 ( .A(KEYINPUT11), .ZN(new_n403_) );
  INV_X1 g266 ( .A(KEYINPUT10), .ZN(new_n404_) );
  NAND2_X1 g267 ( .A1(new_n403_), .A2(new_n404_), .ZN(new_n405_) );
  NAND2_X1 g268 ( .A1(new_n405_), .A2(new_n402_), .ZN(new_n406_) );
  NAND2_X1 g269 ( .A1(G232GAT), .A2(G233GAT), .ZN(new_n407_) );
  NAND2_X1 g270 ( .A1(new_n406_), .A2(new_n407_), .ZN(new_n408_) );
  NAND4_X1 g271 ( .A1(new_n405_), .A2(G232GAT), .A3(G233GAT), .A4(new_n402_), .ZN(new_n409_) );
  NAND2_X1 g272 ( .A1(new_n408_), .A2(new_n409_), .ZN(new_n410_) );
  NAND2_X1 g273 ( .A1(new_n410_), .A2(new_n401_), .ZN(new_n411_) );
  NAND3_X1 g274 ( .A1(new_n408_), .A2(KEYINPUT9), .A3(new_n409_), .ZN(new_n412_) );
  NAND2_X1 g275 ( .A1(new_n411_), .A2(new_n412_), .ZN(new_n413_) );
  INV_X1 g276 ( .A(KEYINPUT8), .ZN(new_n414_) );
  NAND2_X1 g277 ( .A1(new_n324_), .A2(new_n414_), .ZN(new_n415_) );
  NAND2_X1 g278 ( .A1(G43GAT), .A2(KEYINPUT8), .ZN(new_n416_) );
  NAND2_X1 g279 ( .A1(new_n415_), .A2(new_n416_), .ZN(new_n417_) );
  NAND2_X1 g280 ( .A1(new_n417_), .A2(KEYINPUT7), .ZN(new_n418_) );
  INV_X1 g281 ( .A(KEYINPUT7), .ZN(new_n419_) );
  NAND3_X1 g282 ( .A1(new_n415_), .A2(new_n419_), .A3(new_n416_), .ZN(new_n420_) );
  NAND2_X1 g283 ( .A1(new_n418_), .A2(new_n420_), .ZN(new_n421_) );
  INV_X1 g284 ( .A(G85GAT), .ZN(new_n422_) );
  NAND2_X1 g285 ( .A1(new_n422_), .A2(new_n325_), .ZN(new_n423_) );
  NAND2_X1 g286 ( .A1(G85GAT), .A2(G99GAT), .ZN(new_n424_) );
  NAND2_X1 g287 ( .A1(new_n423_), .A2(new_n424_), .ZN(new_n425_) );
  NAND2_X1 g288 ( .A1(new_n425_), .A2(G92GAT), .ZN(new_n426_) );
  NAND3_X1 g289 ( .A1(new_n423_), .A2(new_n353_), .A3(new_n424_), .ZN(new_n427_) );
  NAND2_X1 g290 ( .A1(new_n426_), .A2(new_n427_), .ZN(new_n428_) );
  NAND2_X1 g291 ( .A1(new_n421_), .A2(new_n428_), .ZN(new_n429_) );
  NAND4_X1 g292 ( .A1(new_n418_), .A2(new_n426_), .A3(new_n420_), .A4(new_n427_), .ZN(new_n430_) );
  NAND2_X1 g293 ( .A1(new_n429_), .A2(new_n430_), .ZN(new_n431_) );
  NAND2_X1 g294 ( .A1(new_n431_), .A2(new_n413_), .ZN(new_n432_) );
  NAND4_X1 g295 ( .A1(new_n429_), .A2(new_n411_), .A3(new_n412_), .A4(new_n430_), .ZN(new_n433_) );
  NAND2_X1 g296 ( .A1(new_n432_), .A2(new_n433_), .ZN(new_n434_) );
  NAND2_X1 g297 ( .A1(G106GAT), .A2(G218GAT), .ZN(new_n435_) );
  NAND2_X1 g298 ( .A1(new_n254_), .A2(new_n220_), .ZN(new_n436_) );
  NAND2_X1 g299 ( .A1(new_n436_), .A2(new_n435_), .ZN(new_n437_) );
  NAND2_X1 g300 ( .A1(new_n189_), .A2(new_n437_), .ZN(new_n438_) );
  NAND3_X1 g301 ( .A1(new_n188_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n439_) );
  NAND3_X1 g302 ( .A1(new_n434_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_) );
  NAND2_X1 g303 ( .A1(new_n438_), .A2(new_n439_), .ZN(new_n441_) );
  NAND3_X1 g304 ( .A1(new_n432_), .A2(new_n433_), .A3(new_n441_), .ZN(new_n442_) );
  NAND2_X1 g305 ( .A1(new_n440_), .A2(new_n442_), .ZN(new_n443_) );
  NAND2_X1 g306 ( .A1(new_n443_), .A2(new_n271_), .ZN(new_n444_) );
  NAND3_X1 g307 ( .A1(new_n440_), .A2(new_n273_), .A3(new_n442_), .ZN(new_n445_) );
  NAND2_X1 g308 ( .A1(new_n444_), .A2(new_n445_), .ZN(new_n446_) );
  NAND2_X1 g309 ( .A1(new_n446_), .A2(new_n342_), .ZN(new_n447_) );
  NAND3_X1 g310 ( .A1(new_n444_), .A2(new_n344_), .A3(new_n445_), .ZN(new_n448_) );
  NAND2_X1 g311 ( .A1(new_n447_), .A2(new_n448_), .ZN(new_n449_) );
  NAND2_X1 g312 ( .A1(new_n144_), .A2(G78GAT), .ZN(new_n450_) );
  NAND2_X1 g313 ( .A1(new_n253_), .A2(G155GAT), .ZN(new_n451_) );
  NAND2_X1 g314 ( .A1(new_n450_), .A2(new_n451_), .ZN(new_n452_) );
  NAND2_X1 g315 ( .A1(G127GAT), .A2(G211GAT), .ZN(new_n453_) );
  NAND2_X1 g316 ( .A1(new_n165_), .A2(new_n222_), .ZN(new_n454_) );
  NAND2_X1 g317 ( .A1(new_n454_), .A2(new_n453_), .ZN(new_n455_) );
  NAND2_X1 g318 ( .A1(new_n452_), .A2(new_n455_), .ZN(new_n456_) );
  NAND4_X1 g319 ( .A1(new_n454_), .A2(new_n450_), .A3(new_n451_), .A4(new_n453_), .ZN(new_n457_) );
  NAND2_X1 g320 ( .A1(new_n456_), .A2(new_n457_), .ZN(new_n458_) );
  INV_X1 g321 ( .A(KEYINPUT12), .ZN(new_n459_) );
  NAND2_X1 g322 ( .A1(new_n459_), .A2(KEYINPUT14), .ZN(new_n460_) );
  INV_X1 g323 ( .A(KEYINPUT14), .ZN(new_n461_) );
  NAND2_X1 g324 ( .A1(new_n461_), .A2(KEYINPUT12), .ZN(new_n462_) );
  NAND2_X1 g325 ( .A1(new_n460_), .A2(new_n462_), .ZN(new_n463_) );
  NAND2_X1 g326 ( .A1(G64GAT), .A2(KEYINPUT15), .ZN(new_n464_) );
  INV_X1 g327 ( .A(G64GAT), .ZN(new_n465_) );
  INV_X1 g328 ( .A(KEYINPUT15), .ZN(new_n466_) );
  NAND2_X1 g329 ( .A1(new_n465_), .A2(new_n466_), .ZN(new_n467_) );
  NAND2_X1 g330 ( .A1(new_n467_), .A2(new_n464_), .ZN(new_n468_) );
  NAND2_X1 g331 ( .A1(new_n463_), .A2(new_n468_), .ZN(new_n469_) );
  NAND4_X1 g332 ( .A1(new_n467_), .A2(new_n460_), .A3(new_n462_), .A4(new_n464_), .ZN(new_n470_) );
  NAND2_X1 g333 ( .A1(new_n469_), .A2(new_n470_), .ZN(new_n471_) );
  NAND2_X1 g334 ( .A1(new_n458_), .A2(new_n471_), .ZN(new_n472_) );
  NAND4_X1 g335 ( .A1(new_n456_), .A2(new_n469_), .A3(new_n457_), .A4(new_n470_), .ZN(new_n473_) );
  NAND2_X1 g336 ( .A1(G15GAT), .A2(G22GAT), .ZN(new_n474_) );
  INV_X1 g337 ( .A(new_n474_), .ZN(new_n475_) );
  NOR2_X1 g338 ( .A1(G15GAT), .A2(G22GAT), .ZN(new_n476_) );
  NOR2_X1 g339 ( .A1(new_n475_), .A2(new_n476_), .ZN(new_n477_) );
  NOR2_X1 g340 ( .A1(new_n477_), .A2(G1GAT), .ZN(new_n478_) );
  NAND2_X1 g341 ( .A1(new_n477_), .A2(G1GAT), .ZN(new_n479_) );
  INV_X1 g342 ( .A(new_n479_), .ZN(new_n480_) );
  NOR2_X1 g343 ( .A1(new_n480_), .A2(new_n478_), .ZN(new_n481_) );
  INV_X1 g344 ( .A(new_n481_), .ZN(new_n482_) );
  INV_X1 g345 ( .A(KEYINPUT13), .ZN(new_n483_) );
  NAND2_X1 g346 ( .A1(G57GAT), .A2(G71GAT), .ZN(new_n484_) );
  INV_X1 g347 ( .A(new_n484_), .ZN(new_n485_) );
  NOR2_X1 g348 ( .A1(G57GAT), .A2(G71GAT), .ZN(new_n486_) );
  NOR2_X1 g349 ( .A1(new_n485_), .A2(new_n486_), .ZN(new_n487_) );
  NOR2_X1 g350 ( .A1(new_n487_), .A2(new_n483_), .ZN(new_n488_) );
  NAND2_X1 g351 ( .A1(new_n487_), .A2(new_n483_), .ZN(new_n489_) );
  INV_X1 g352 ( .A(new_n489_), .ZN(new_n490_) );
  NOR2_X1 g353 ( .A1(new_n490_), .A2(new_n488_), .ZN(new_n491_) );
  INV_X1 g354 ( .A(new_n491_), .ZN(new_n492_) );
  NAND2_X1 g355 ( .A1(new_n492_), .A2(new_n482_), .ZN(new_n493_) );
  NAND2_X1 g356 ( .A1(new_n481_), .A2(new_n491_), .ZN(new_n494_) );
  NAND4_X1 g357 ( .A1(new_n493_), .A2(new_n472_), .A3(new_n473_), .A4(new_n494_), .ZN(new_n495_) );
  NAND2_X1 g358 ( .A1(new_n472_), .A2(new_n473_), .ZN(new_n496_) );
  NAND2_X1 g359 ( .A1(new_n493_), .A2(new_n494_), .ZN(new_n497_) );
  NAND2_X1 g360 ( .A1(new_n497_), .A2(new_n496_), .ZN(new_n498_) );
  NAND2_X1 g361 ( .A1(new_n498_), .A2(new_n495_), .ZN(new_n499_) );
  NAND2_X1 g362 ( .A1(new_n499_), .A2(new_n365_), .ZN(new_n500_) );
  NAND3_X1 g363 ( .A1(new_n498_), .A2(new_n363_), .A3(new_n495_), .ZN(new_n501_) );
  NAND2_X1 g364 ( .A1(new_n500_), .A2(new_n501_), .ZN(new_n502_) );
  NAND3_X1 g365 ( .A1(new_n502_), .A2(G231GAT), .A3(G233GAT), .ZN(new_n503_) );
  NAND2_X1 g366 ( .A1(G231GAT), .A2(G233GAT), .ZN(new_n504_) );
  NAND3_X1 g367 ( .A1(new_n500_), .A2(new_n501_), .A3(new_n504_), .ZN(new_n505_) );
  NAND2_X1 g368 ( .A1(new_n503_), .A2(new_n505_), .ZN(new_n506_) );
  INV_X1 g369 ( .A(new_n506_), .ZN(new_n507_) );
  NAND2_X1 g370 ( .A1(new_n507_), .A2(new_n449_), .ZN(new_n508_) );
  NAND2_X1 g371 ( .A1(new_n508_), .A2(new_n400_), .ZN(new_n509_) );
  NAND3_X1 g372 ( .A1(new_n507_), .A2(KEYINPUT16), .A3(new_n449_), .ZN(new_n510_) );
  NAND2_X1 g373 ( .A1(new_n509_), .A2(new_n510_), .ZN(new_n511_) );
  NAND2_X1 g374 ( .A1(new_n399_), .A2(new_n511_), .ZN(new_n512_) );
  INV_X1 g375 ( .A(new_n512_), .ZN(new_n513_) );
  NAND2_X1 g376 ( .A1(new_n260_), .A2(new_n428_), .ZN(new_n514_) );
  NAND4_X1 g377 ( .A1(new_n258_), .A2(new_n426_), .A3(new_n259_), .A4(new_n427_), .ZN(new_n515_) );
  NAND2_X1 g378 ( .A1(new_n514_), .A2(new_n515_), .ZN(new_n516_) );
  INV_X1 g379 ( .A(KEYINPUT32), .ZN(new_n517_) );
  INV_X1 g380 ( .A(KEYINPUT31), .ZN(new_n518_) );
  NAND2_X1 g381 ( .A1(new_n518_), .A2(KEYINPUT33), .ZN(new_n519_) );
  INV_X1 g382 ( .A(KEYINPUT33), .ZN(new_n520_) );
  NAND2_X1 g383 ( .A1(new_n520_), .A2(KEYINPUT31), .ZN(new_n521_) );
  NAND2_X1 g384 ( .A1(new_n519_), .A2(new_n521_), .ZN(new_n522_) );
  NAND2_X1 g385 ( .A1(G230GAT), .A2(G233GAT), .ZN(new_n523_) );
  NAND2_X1 g386 ( .A1(new_n522_), .A2(new_n523_), .ZN(new_n524_) );
  NAND4_X1 g387 ( .A1(new_n519_), .A2(new_n521_), .A3(G230GAT), .A4(G233GAT), .ZN(new_n525_) );
  NAND2_X1 g388 ( .A1(new_n524_), .A2(new_n525_), .ZN(new_n526_) );
  NAND2_X1 g389 ( .A1(new_n526_), .A2(new_n517_), .ZN(new_n527_) );
  NAND3_X1 g390 ( .A1(new_n524_), .A2(KEYINPUT32), .A3(new_n525_), .ZN(new_n528_) );
  NAND2_X1 g391 ( .A1(new_n527_), .A2(new_n528_), .ZN(new_n529_) );
  NAND2_X1 g392 ( .A1(new_n516_), .A2(new_n529_), .ZN(new_n530_) );
  NAND4_X1 g393 ( .A1(new_n514_), .A2(new_n527_), .A3(new_n515_), .A4(new_n528_), .ZN(new_n531_) );
  NAND2_X1 g394 ( .A1(new_n530_), .A2(new_n531_), .ZN(new_n532_) );
  NAND2_X1 g395 ( .A1(new_n532_), .A2(new_n351_), .ZN(new_n533_) );
  NAND3_X1 g396 ( .A1(new_n530_), .A2(new_n350_), .A3(new_n531_), .ZN(new_n534_) );
  NAND2_X1 g397 ( .A1(new_n533_), .A2(new_n534_), .ZN(new_n535_) );
  NAND2_X1 g398 ( .A1(G120GAT), .A2(G204GAT), .ZN(new_n536_) );
  INV_X1 g399 ( .A(new_n536_), .ZN(new_n537_) );
  NOR2_X1 g400 ( .A1(G120GAT), .A2(G204GAT), .ZN(new_n538_) );
  NOR2_X1 g401 ( .A1(new_n537_), .A2(new_n538_), .ZN(new_n539_) );
  NAND2_X1 g402 ( .A1(new_n535_), .A2(new_n539_), .ZN(new_n540_) );
  INV_X1 g403 ( .A(new_n539_), .ZN(new_n541_) );
  NAND3_X1 g404 ( .A1(new_n533_), .A2(new_n534_), .A3(new_n541_), .ZN(new_n542_) );
  NAND2_X1 g405 ( .A1(new_n540_), .A2(new_n542_), .ZN(new_n543_) );
  NAND2_X1 g406 ( .A1(new_n543_), .A2(new_n492_), .ZN(new_n544_) );
  NAND3_X1 g407 ( .A1(new_n540_), .A2(new_n491_), .A3(new_n542_), .ZN(new_n545_) );
  NAND2_X1 g408 ( .A1(new_n544_), .A2(new_n545_), .ZN(new_n546_) );
  INV_X1 g409 ( .A(KEYINPUT29), .ZN(new_n547_) );
  NAND2_X1 g410 ( .A1(new_n547_), .A2(KEYINPUT30), .ZN(new_n548_) );
  INV_X1 g411 ( .A(KEYINPUT30), .ZN(new_n549_) );
  NAND2_X1 g412 ( .A1(new_n549_), .A2(KEYINPUT29), .ZN(new_n550_) );
  NAND2_X1 g413 ( .A1(new_n548_), .A2(new_n550_), .ZN(new_n551_) );
  NAND2_X1 g414 ( .A1(G8GAT), .A2(G169GAT), .ZN(new_n552_) );
  INV_X1 g415 ( .A(G8GAT), .ZN(new_n553_) );
  NAND2_X1 g416 ( .A1(new_n553_), .A2(new_n311_), .ZN(new_n554_) );
  NAND2_X1 g417 ( .A1(new_n554_), .A2(new_n552_), .ZN(new_n555_) );
  NAND2_X1 g418 ( .A1(new_n551_), .A2(new_n555_), .ZN(new_n556_) );
  NAND4_X1 g419 ( .A1(new_n554_), .A2(new_n548_), .A3(new_n550_), .A4(new_n552_), .ZN(new_n557_) );
  NAND2_X1 g420 ( .A1(new_n556_), .A2(new_n557_), .ZN(new_n558_) );
  NAND2_X1 g421 ( .A1(new_n219_), .A2(G113GAT), .ZN(new_n559_) );
  NAND2_X1 g422 ( .A1(new_n171_), .A2(G197GAT), .ZN(new_n560_) );
  NAND2_X1 g423 ( .A1(new_n559_), .A2(new_n560_), .ZN(new_n561_) );
  NAND2_X1 g424 ( .A1(G29GAT), .A2(G141GAT), .ZN(new_n562_) );
  INV_X1 g425 ( .A(G29GAT), .ZN(new_n563_) );
  NAND2_X1 g426 ( .A1(new_n563_), .A2(new_n139_), .ZN(new_n564_) );
  NAND2_X1 g427 ( .A1(new_n564_), .A2(new_n562_), .ZN(new_n565_) );
  NAND2_X1 g428 ( .A1(new_n561_), .A2(new_n565_), .ZN(new_n566_) );
  NAND4_X1 g429 ( .A1(new_n564_), .A2(new_n559_), .A3(new_n560_), .A4(new_n562_), .ZN(new_n567_) );
  NAND2_X1 g430 ( .A1(new_n566_), .A2(new_n567_), .ZN(new_n568_) );
  NAND2_X1 g431 ( .A1(new_n558_), .A2(new_n568_), .ZN(new_n569_) );
  NAND4_X1 g432 ( .A1(new_n556_), .A2(new_n566_), .A3(new_n557_), .A4(new_n567_), .ZN(new_n570_) );
  NAND2_X1 g433 ( .A1(new_n569_), .A2(new_n570_), .ZN(new_n571_) );
  NAND2_X1 g434 ( .A1(new_n482_), .A2(new_n421_), .ZN(new_n572_) );
  NAND3_X1 g435 ( .A1(new_n481_), .A2(new_n418_), .A3(new_n420_), .ZN(new_n573_) );
  NAND2_X1 g436 ( .A1(new_n572_), .A2(new_n573_), .ZN(new_n574_) );
  NAND2_X1 g437 ( .A1(new_n574_), .A2(new_n571_), .ZN(new_n575_) );
  NAND4_X1 g438 ( .A1(new_n572_), .A2(new_n569_), .A3(new_n570_), .A4(new_n573_), .ZN(new_n576_) );
  NAND2_X1 g439 ( .A1(new_n575_), .A2(new_n576_), .ZN(new_n577_) );
  NAND2_X1 g440 ( .A1(new_n267_), .A2(G36GAT), .ZN(new_n578_) );
  INV_X1 g441 ( .A(G36GAT), .ZN(new_n579_) );
  NAND2_X1 g442 ( .A1(new_n579_), .A2(G50GAT), .ZN(new_n580_) );
  NAND2_X1 g443 ( .A1(new_n578_), .A2(new_n580_), .ZN(new_n581_) );
  NAND2_X1 g444 ( .A1(G229GAT), .A2(G233GAT), .ZN(new_n582_) );
  NAND2_X1 g445 ( .A1(new_n581_), .A2(new_n582_), .ZN(new_n583_) );
  NAND4_X1 g446 ( .A1(new_n578_), .A2(new_n580_), .A3(G229GAT), .A4(G233GAT), .ZN(new_n584_) );
  NAND2_X1 g447 ( .A1(new_n583_), .A2(new_n584_), .ZN(new_n585_) );
  NAND2_X1 g448 ( .A1(new_n577_), .A2(new_n585_), .ZN(new_n586_) );
  NAND4_X1 g449 ( .A1(new_n575_), .A2(new_n576_), .A3(new_n583_), .A4(new_n584_), .ZN(new_n587_) );
  NAND2_X1 g450 ( .A1(new_n586_), .A2(new_n587_), .ZN(new_n588_) );
  INV_X1 g451 ( .A(new_n588_), .ZN(new_n589_) );
  NAND2_X1 g452 ( .A1(new_n546_), .A2(new_n589_), .ZN(new_n590_) );
  INV_X1 g453 ( .A(new_n590_), .ZN(new_n591_) );
  NAND2_X1 g454 ( .A1(new_n513_), .A2(new_n591_), .ZN(new_n592_) );
  INV_X1 g455 ( .A(new_n592_), .ZN(new_n593_) );
  NAND2_X1 g456 ( .A1(new_n593_), .A2(new_n217_), .ZN(new_n594_) );
  NAND2_X1 g457 ( .A1(new_n594_), .A2(KEYINPUT34), .ZN(new_n595_) );
  INV_X1 g458 ( .A(KEYINPUT34), .ZN(new_n596_) );
  NAND3_X1 g459 ( .A1(new_n593_), .A2(new_n596_), .A3(new_n217_), .ZN(new_n597_) );
  NAND2_X1 g460 ( .A1(new_n595_), .A2(new_n597_), .ZN(new_n598_) );
  NAND2_X1 g461 ( .A1(new_n598_), .A2(G1GAT), .ZN(new_n599_) );
  NAND3_X1 g462 ( .A1(new_n595_), .A2(new_n164_), .A3(new_n597_), .ZN(new_n600_) );
  NAND2_X1 g463 ( .A1(new_n599_), .A2(new_n600_), .ZN(G1324GAT) );
  NAND2_X1 g464 ( .A1(new_n593_), .A2(new_n374_), .ZN(new_n602_) );
  NAND2_X1 g465 ( .A1(new_n602_), .A2(G8GAT), .ZN(new_n603_) );
  NAND3_X1 g466 ( .A1(new_n593_), .A2(new_n553_), .A3(new_n374_), .ZN(new_n604_) );
  NAND2_X1 g467 ( .A1(new_n603_), .A2(new_n604_), .ZN(G1325GAT) );
  NAND2_X1 g468 ( .A1(new_n593_), .A2(new_n338_), .ZN(new_n606_) );
  NOR2_X1 g469 ( .A1(new_n281_), .A2(KEYINPUT35), .ZN(new_n607_) );
  NAND2_X1 g470 ( .A1(new_n281_), .A2(KEYINPUT35), .ZN(new_n608_) );
  INV_X1 g471 ( .A(new_n608_), .ZN(new_n609_) );
  NOR2_X1 g472 ( .A1(new_n609_), .A2(new_n607_), .ZN(new_n610_) );
  INV_X1 g473 ( .A(new_n610_), .ZN(new_n611_) );
  NAND2_X1 g474 ( .A1(new_n606_), .A2(new_n611_), .ZN(new_n612_) );
  NAND3_X1 g475 ( .A1(new_n593_), .A2(new_n338_), .A3(new_n610_), .ZN(new_n613_) );
  NAND2_X1 g476 ( .A1(new_n612_), .A2(new_n613_), .ZN(G1326GAT) );
  INV_X1 g477 ( .A(new_n395_), .ZN(new_n615_) );
  NAND2_X1 g478 ( .A1(new_n593_), .A2(new_n615_), .ZN(new_n616_) );
  NAND2_X1 g479 ( .A1(new_n616_), .A2(G22GAT), .ZN(new_n617_) );
  NAND3_X1 g480 ( .A1(new_n593_), .A2(new_n246_), .A3(new_n615_), .ZN(new_n618_) );
  NAND2_X1 g481 ( .A1(new_n617_), .A2(new_n618_), .ZN(G1327GAT) );
  INV_X1 g482 ( .A(KEYINPUT38), .ZN(new_n620_) );
  NAND2_X1 g483 ( .A1(new_n449_), .A2(KEYINPUT36), .ZN(new_n621_) );
  INV_X1 g484 ( .A(KEYINPUT36), .ZN(new_n622_) );
  NAND3_X1 g485 ( .A1(new_n447_), .A2(new_n622_), .A3(new_n448_), .ZN(new_n623_) );
  NAND2_X1 g486 ( .A1(new_n621_), .A2(new_n623_), .ZN(new_n624_) );
  INV_X1 g487 ( .A(new_n624_), .ZN(new_n625_) );
  NAND2_X1 g488 ( .A1(new_n625_), .A2(new_n506_), .ZN(new_n626_) );
  INV_X1 g489 ( .A(new_n626_), .ZN(new_n627_) );
  NAND2_X1 g490 ( .A1(new_n399_), .A2(new_n627_), .ZN(new_n628_) );
  NAND2_X1 g491 ( .A1(new_n628_), .A2(KEYINPUT37), .ZN(new_n629_) );
  INV_X1 g492 ( .A(KEYINPUT37), .ZN(new_n630_) );
  NAND3_X1 g493 ( .A1(new_n399_), .A2(new_n630_), .A3(new_n627_), .ZN(new_n631_) );
  NAND2_X1 g494 ( .A1(new_n629_), .A2(new_n631_), .ZN(new_n632_) );
  NAND2_X1 g495 ( .A1(new_n632_), .A2(new_n591_), .ZN(new_n633_) );
  NAND2_X1 g496 ( .A1(new_n633_), .A2(new_n620_), .ZN(new_n634_) );
  NAND3_X1 g497 ( .A1(new_n632_), .A2(KEYINPUT38), .A3(new_n591_), .ZN(new_n635_) );
  NAND2_X1 g498 ( .A1(new_n634_), .A2(new_n635_), .ZN(new_n636_) );
  NAND2_X1 g499 ( .A1(new_n636_), .A2(new_n217_), .ZN(new_n637_) );
  NOR2_X1 g500 ( .A1(new_n563_), .A2(KEYINPUT39), .ZN(new_n638_) );
  NAND2_X1 g501 ( .A1(new_n563_), .A2(KEYINPUT39), .ZN(new_n639_) );
  INV_X1 g502 ( .A(new_n639_), .ZN(new_n640_) );
  NOR2_X1 g503 ( .A1(new_n640_), .A2(new_n638_), .ZN(new_n641_) );
  INV_X1 g504 ( .A(new_n641_), .ZN(new_n642_) );
  NAND2_X1 g505 ( .A1(new_n637_), .A2(new_n642_), .ZN(new_n643_) );
  NAND3_X1 g506 ( .A1(new_n636_), .A2(new_n217_), .A3(new_n641_), .ZN(new_n644_) );
  NAND2_X1 g507 ( .A1(new_n643_), .A2(new_n644_), .ZN(G1328GAT) );
  NAND2_X1 g508 ( .A1(new_n636_), .A2(new_n374_), .ZN(new_n646_) );
  NAND2_X1 g509 ( .A1(new_n646_), .A2(G36GAT), .ZN(new_n647_) );
  NAND3_X1 g510 ( .A1(new_n636_), .A2(new_n579_), .A3(new_n374_), .ZN(new_n648_) );
  NAND2_X1 g511 ( .A1(new_n647_), .A2(new_n648_), .ZN(G1329GAT) );
  NAND2_X1 g512 ( .A1(new_n636_), .A2(new_n338_), .ZN(new_n650_) );
  NAND2_X1 g513 ( .A1(new_n650_), .A2(KEYINPUT40), .ZN(new_n651_) );
  INV_X1 g514 ( .A(KEYINPUT40), .ZN(new_n652_) );
  NAND3_X1 g515 ( .A1(new_n636_), .A2(new_n652_), .A3(new_n338_), .ZN(new_n653_) );
  NAND2_X1 g516 ( .A1(new_n651_), .A2(new_n653_), .ZN(new_n654_) );
  NAND2_X1 g517 ( .A1(new_n654_), .A2(G43GAT), .ZN(new_n655_) );
  NAND3_X1 g518 ( .A1(new_n651_), .A2(new_n324_), .A3(new_n653_), .ZN(new_n656_) );
  NAND2_X1 g519 ( .A1(new_n655_), .A2(new_n656_), .ZN(G1330GAT) );
  NAND2_X1 g520 ( .A1(new_n636_), .A2(new_n615_), .ZN(new_n658_) );
  NAND2_X1 g521 ( .A1(new_n658_), .A2(G50GAT), .ZN(new_n659_) );
  NAND3_X1 g522 ( .A1(new_n636_), .A2(new_n267_), .A3(new_n615_), .ZN(new_n660_) );
  NAND2_X1 g523 ( .A1(new_n659_), .A2(new_n660_), .ZN(G1331GAT) );
  INV_X1 g524 ( .A(KEYINPUT41), .ZN(new_n662_) );
  NAND2_X1 g525 ( .A1(new_n546_), .A2(new_n662_), .ZN(new_n663_) );
  NAND3_X1 g526 ( .A1(new_n544_), .A2(KEYINPUT41), .A3(new_n545_), .ZN(new_n664_) );
  NAND2_X1 g527 ( .A1(new_n663_), .A2(new_n664_), .ZN(new_n665_) );
  INV_X1 g528 ( .A(new_n665_), .ZN(new_n666_) );
  NAND2_X1 g529 ( .A1(new_n666_), .A2(new_n588_), .ZN(new_n667_) );
  INV_X1 g530 ( .A(new_n667_), .ZN(new_n668_) );
  NAND2_X1 g531 ( .A1(new_n513_), .A2(new_n668_), .ZN(new_n669_) );
  INV_X1 g532 ( .A(new_n669_), .ZN(new_n670_) );
  NAND2_X1 g533 ( .A1(new_n670_), .A2(new_n217_), .ZN(new_n671_) );
  NAND2_X1 g534 ( .A1(G57GAT), .A2(KEYINPUT42), .ZN(new_n672_) );
  INV_X1 g535 ( .A(new_n672_), .ZN(new_n673_) );
  NOR2_X1 g536 ( .A1(G57GAT), .A2(KEYINPUT42), .ZN(new_n674_) );
  NOR2_X1 g537 ( .A1(new_n673_), .A2(new_n674_), .ZN(new_n675_) );
  INV_X1 g538 ( .A(new_n675_), .ZN(new_n676_) );
  NAND2_X1 g539 ( .A1(new_n671_), .A2(new_n676_), .ZN(new_n677_) );
  NAND3_X1 g540 ( .A1(new_n670_), .A2(new_n217_), .A3(new_n675_), .ZN(new_n678_) );
  NAND2_X1 g541 ( .A1(new_n677_), .A2(new_n678_), .ZN(G1332GAT) );
  NAND2_X1 g542 ( .A1(new_n670_), .A2(new_n374_), .ZN(new_n680_) );
  NAND2_X1 g543 ( .A1(new_n680_), .A2(G64GAT), .ZN(new_n681_) );
  NAND3_X1 g544 ( .A1(new_n670_), .A2(new_n465_), .A3(new_n374_), .ZN(new_n682_) );
  NAND2_X1 g545 ( .A1(new_n681_), .A2(new_n682_), .ZN(G1333GAT) );
  NAND2_X1 g546 ( .A1(new_n670_), .A2(new_n338_), .ZN(new_n684_) );
  NAND2_X1 g547 ( .A1(new_n684_), .A2(G71GAT), .ZN(new_n685_) );
  NAND3_X1 g548 ( .A1(new_n670_), .A2(new_n289_), .A3(new_n338_), .ZN(new_n686_) );
  NAND2_X1 g549 ( .A1(new_n685_), .A2(new_n686_), .ZN(G1334GAT) );
  NAND2_X1 g550 ( .A1(new_n670_), .A2(new_n615_), .ZN(new_n688_) );
  NOR2_X1 g551 ( .A1(new_n253_), .A2(KEYINPUT43), .ZN(new_n689_) );
  NAND2_X1 g552 ( .A1(new_n253_), .A2(KEYINPUT43), .ZN(new_n690_) );
  INV_X1 g553 ( .A(new_n690_), .ZN(new_n691_) );
  NOR2_X1 g554 ( .A1(new_n691_), .A2(new_n689_), .ZN(new_n692_) );
  INV_X1 g555 ( .A(new_n692_), .ZN(new_n693_) );
  NAND2_X1 g556 ( .A1(new_n688_), .A2(new_n693_), .ZN(new_n694_) );
  NAND3_X1 g557 ( .A1(new_n670_), .A2(new_n615_), .A3(new_n692_), .ZN(new_n695_) );
  NAND2_X1 g558 ( .A1(new_n694_), .A2(new_n695_), .ZN(G1335GAT) );
  NAND2_X1 g559 ( .A1(new_n632_), .A2(new_n668_), .ZN(new_n697_) );
  INV_X1 g560 ( .A(new_n697_), .ZN(new_n698_) );
  NAND2_X1 g561 ( .A1(new_n698_), .A2(new_n217_), .ZN(new_n699_) );
  NAND2_X1 g562 ( .A1(new_n699_), .A2(G85GAT), .ZN(new_n700_) );
  NAND3_X1 g563 ( .A1(new_n698_), .A2(new_n422_), .A3(new_n217_), .ZN(new_n701_) );
  NAND2_X1 g564 ( .A1(new_n700_), .A2(new_n701_), .ZN(G1336GAT) );
  NAND2_X1 g565 ( .A1(new_n698_), .A2(new_n374_), .ZN(new_n703_) );
  NAND2_X1 g566 ( .A1(new_n703_), .A2(G92GAT), .ZN(new_n704_) );
  NAND3_X1 g567 ( .A1(new_n698_), .A2(new_n353_), .A3(new_n374_), .ZN(new_n705_) );
  NAND2_X1 g568 ( .A1(new_n704_), .A2(new_n705_), .ZN(G1337GAT) );
  NAND2_X1 g569 ( .A1(new_n698_), .A2(new_n338_), .ZN(new_n707_) );
  NAND2_X1 g570 ( .A1(new_n707_), .A2(G99GAT), .ZN(new_n708_) );
  NAND3_X1 g571 ( .A1(new_n698_), .A2(new_n325_), .A3(new_n338_), .ZN(new_n709_) );
  NAND2_X1 g572 ( .A1(new_n708_), .A2(new_n709_), .ZN(G1338GAT) );
  NAND2_X1 g573 ( .A1(new_n698_), .A2(new_n615_), .ZN(new_n711_) );
  NAND2_X1 g574 ( .A1(new_n711_), .A2(KEYINPUT44), .ZN(new_n712_) );
  INV_X1 g575 ( .A(KEYINPUT44), .ZN(new_n713_) );
  NAND3_X1 g576 ( .A1(new_n698_), .A2(new_n713_), .A3(new_n615_), .ZN(new_n714_) );
  NAND2_X1 g577 ( .A1(new_n712_), .A2(new_n714_), .ZN(new_n715_) );
  NAND2_X1 g578 ( .A1(new_n715_), .A2(G106GAT), .ZN(new_n716_) );
  NAND3_X1 g579 ( .A1(new_n712_), .A2(new_n254_), .A3(new_n714_), .ZN(new_n717_) );
  NAND2_X1 g580 ( .A1(new_n716_), .A2(new_n717_), .ZN(G1339GAT) );
  INV_X1 g581 ( .A(KEYINPUT47), .ZN(new_n719_) );
  NAND4_X1 g582 ( .A1(new_n663_), .A2(KEYINPUT46), .A3(new_n589_), .A4(new_n664_), .ZN(new_n720_) );
  INV_X1 g583 ( .A(KEYINPUT46), .ZN(new_n721_) );
  NAND3_X1 g584 ( .A1(new_n663_), .A2(new_n589_), .A3(new_n664_), .ZN(new_n722_) );
  NAND2_X1 g585 ( .A1(new_n722_), .A2(new_n721_), .ZN(new_n723_) );
  NAND2_X1 g586 ( .A1(new_n449_), .A2(new_n506_), .ZN(new_n724_) );
  INV_X1 g587 ( .A(new_n724_), .ZN(new_n725_) );
  NAND4_X1 g588 ( .A1(new_n723_), .A2(new_n719_), .A3(new_n720_), .A4(new_n725_), .ZN(new_n726_) );
  NAND3_X1 g589 ( .A1(new_n723_), .A2(new_n720_), .A3(new_n725_), .ZN(new_n727_) );
  NAND2_X1 g590 ( .A1(new_n727_), .A2(KEYINPUT47), .ZN(new_n728_) );
  INV_X1 g591 ( .A(KEYINPUT45), .ZN(new_n729_) );
  NAND4_X1 g592 ( .A1(new_n621_), .A2(new_n507_), .A3(new_n729_), .A4(new_n623_), .ZN(new_n730_) );
  NAND3_X1 g593 ( .A1(new_n621_), .A2(new_n507_), .A3(new_n623_), .ZN(new_n731_) );
  NAND2_X1 g594 ( .A1(new_n731_), .A2(KEYINPUT45), .ZN(new_n732_) );
  NAND4_X1 g595 ( .A1(new_n732_), .A2(new_n546_), .A3(new_n588_), .A4(new_n730_), .ZN(new_n733_) );
  NAND4_X1 g596 ( .A1(new_n728_), .A2(KEYINPUT48), .A3(new_n733_), .A4(new_n726_), .ZN(new_n734_) );
  INV_X1 g597 ( .A(KEYINPUT48), .ZN(new_n735_) );
  NAND3_X1 g598 ( .A1(new_n728_), .A2(new_n726_), .A3(new_n733_), .ZN(new_n736_) );
  NAND2_X1 g599 ( .A1(new_n736_), .A2(new_n735_), .ZN(new_n737_) );
  NAND3_X1 g600 ( .A1(new_n737_), .A2(new_n397_), .A3(new_n734_), .ZN(new_n738_) );
  INV_X1 g601 ( .A(new_n738_), .ZN(new_n739_) );
  NAND3_X1 g602 ( .A1(new_n739_), .A2(new_n338_), .A3(new_n395_), .ZN(new_n740_) );
  NOR2_X1 g603 ( .A1(new_n740_), .A2(new_n588_), .ZN(new_n741_) );
  INV_X1 g604 ( .A(new_n741_), .ZN(new_n742_) );
  NAND2_X1 g605 ( .A1(new_n742_), .A2(G113GAT), .ZN(new_n743_) );
  NAND2_X1 g606 ( .A1(new_n741_), .A2(new_n171_), .ZN(new_n744_) );
  NAND2_X1 g607 ( .A1(new_n743_), .A2(new_n744_), .ZN(G1340GAT) );
  NOR2_X1 g608 ( .A1(new_n740_), .A2(new_n665_), .ZN(new_n746_) );
  INV_X1 g609 ( .A(new_n746_), .ZN(new_n747_) );
  NOR2_X1 g610 ( .A1(new_n167_), .A2(KEYINPUT49), .ZN(new_n748_) );
  NAND2_X1 g611 ( .A1(new_n167_), .A2(KEYINPUT49), .ZN(new_n749_) );
  INV_X1 g612 ( .A(new_n749_), .ZN(new_n750_) );
  NOR2_X1 g613 ( .A1(new_n750_), .A2(new_n748_), .ZN(new_n751_) );
  INV_X1 g614 ( .A(new_n751_), .ZN(new_n752_) );
  NAND2_X1 g615 ( .A1(new_n747_), .A2(new_n752_), .ZN(new_n753_) );
  NAND2_X1 g616 ( .A1(new_n746_), .A2(new_n751_), .ZN(new_n754_) );
  NAND2_X1 g617 ( .A1(new_n753_), .A2(new_n754_), .ZN(G1341GAT) );
  NOR2_X1 g618 ( .A1(new_n740_), .A2(new_n506_), .ZN(new_n756_) );
  NAND2_X1 g619 ( .A1(new_n756_), .A2(KEYINPUT50), .ZN(new_n757_) );
  INV_X1 g620 ( .A(KEYINPUT50), .ZN(new_n758_) );
  INV_X1 g621 ( .A(new_n756_), .ZN(new_n759_) );
  NAND2_X1 g622 ( .A1(new_n759_), .A2(new_n758_), .ZN(new_n760_) );
  NAND2_X1 g623 ( .A1(new_n760_), .A2(new_n757_), .ZN(new_n761_) );
  NAND2_X1 g624 ( .A1(new_n761_), .A2(new_n165_), .ZN(new_n762_) );
  NAND3_X1 g625 ( .A1(new_n760_), .A2(G127GAT), .A3(new_n757_), .ZN(new_n763_) );
  NAND2_X1 g626 ( .A1(new_n762_), .A2(new_n763_), .ZN(G1342GAT) );
  NOR2_X1 g627 ( .A1(new_n740_), .A2(new_n449_), .ZN(new_n765_) );
  NAND2_X1 g628 ( .A1(G134GAT), .A2(KEYINPUT51), .ZN(new_n766_) );
  INV_X1 g629 ( .A(new_n766_), .ZN(new_n767_) );
  NOR2_X1 g630 ( .A1(G134GAT), .A2(KEYINPUT51), .ZN(new_n768_) );
  NOR2_X1 g631 ( .A1(new_n767_), .A2(new_n768_), .ZN(new_n769_) );
  INV_X1 g632 ( .A(new_n769_), .ZN(new_n770_) );
  NAND2_X1 g633 ( .A1(new_n765_), .A2(new_n770_), .ZN(new_n771_) );
  INV_X1 g634 ( .A(new_n765_), .ZN(new_n772_) );
  NAND2_X1 g635 ( .A1(new_n772_), .A2(new_n769_), .ZN(new_n773_) );
  NAND2_X1 g636 ( .A1(new_n773_), .A2(new_n771_), .ZN(G1343GAT) );
  NAND2_X1 g637 ( .A1(new_n739_), .A2(new_n388_), .ZN(new_n775_) );
  NOR2_X1 g638 ( .A1(new_n775_), .A2(new_n588_), .ZN(new_n776_) );
  INV_X1 g639 ( .A(new_n776_), .ZN(new_n777_) );
  NAND2_X1 g640 ( .A1(new_n777_), .A2(G141GAT), .ZN(new_n778_) );
  NAND2_X1 g641 ( .A1(new_n776_), .A2(new_n139_), .ZN(new_n779_) );
  NAND2_X1 g642 ( .A1(new_n778_), .A2(new_n779_), .ZN(G1344GAT) );
  NOR2_X1 g643 ( .A1(new_n775_), .A2(new_n665_), .ZN(new_n781_) );
  INV_X1 g644 ( .A(new_n781_), .ZN(new_n782_) );
  NAND2_X1 g645 ( .A1(KEYINPUT53), .A2(KEYINPUT52), .ZN(new_n783_) );
  INV_X1 g646 ( .A(new_n783_), .ZN(new_n784_) );
  NOR2_X1 g647 ( .A1(KEYINPUT53), .A2(KEYINPUT52), .ZN(new_n785_) );
  NOR2_X1 g648 ( .A1(new_n784_), .A2(new_n785_), .ZN(new_n786_) );
  INV_X1 g649 ( .A(new_n786_), .ZN(new_n787_) );
  NAND2_X1 g650 ( .A1(new_n782_), .A2(new_n787_), .ZN(new_n788_) );
  NAND2_X1 g651 ( .A1(new_n781_), .A2(new_n786_), .ZN(new_n789_) );
  NAND2_X1 g652 ( .A1(new_n788_), .A2(new_n789_), .ZN(new_n790_) );
  NAND2_X1 g653 ( .A1(new_n790_), .A2(new_n207_), .ZN(new_n791_) );
  NAND3_X1 g654 ( .A1(new_n788_), .A2(G148GAT), .A3(new_n789_), .ZN(new_n792_) );
  NAND2_X1 g655 ( .A1(new_n791_), .A2(new_n792_), .ZN(G1345GAT) );
  NOR2_X1 g656 ( .A1(new_n775_), .A2(new_n506_), .ZN(new_n794_) );
  INV_X1 g657 ( .A(new_n794_), .ZN(new_n795_) );
  NAND2_X1 g658 ( .A1(new_n795_), .A2(G155GAT), .ZN(new_n796_) );
  NAND2_X1 g659 ( .A1(new_n794_), .A2(new_n144_), .ZN(new_n797_) );
  NAND2_X1 g660 ( .A1(new_n796_), .A2(new_n797_), .ZN(G1346GAT) );
  NOR2_X1 g661 ( .A1(new_n775_), .A2(new_n449_), .ZN(new_n799_) );
  INV_X1 g662 ( .A(new_n799_), .ZN(new_n800_) );
  NAND2_X1 g663 ( .A1(new_n800_), .A2(G162GAT), .ZN(new_n801_) );
  NAND2_X1 g664 ( .A1(new_n799_), .A2(new_n269_), .ZN(new_n802_) );
  NAND2_X1 g665 ( .A1(new_n801_), .A2(new_n802_), .ZN(G1347GAT) );
  INV_X1 g666 ( .A(KEYINPUT54), .ZN(new_n804_) );
  NAND4_X1 g667 ( .A1(new_n737_), .A2(new_n804_), .A3(new_n374_), .A4(new_n734_), .ZN(new_n805_) );
  NAND3_X1 g668 ( .A1(new_n737_), .A2(new_n374_), .A3(new_n734_), .ZN(new_n806_) );
  NAND2_X1 g669 ( .A1(new_n806_), .A2(KEYINPUT54), .ZN(new_n807_) );
  NAND4_X1 g670 ( .A1(new_n807_), .A2(new_n216_), .A3(new_n280_), .A4(new_n805_), .ZN(new_n808_) );
  NAND2_X1 g671 ( .A1(new_n808_), .A2(KEYINPUT55), .ZN(new_n809_) );
  INV_X1 g672 ( .A(KEYINPUT55), .ZN(new_n810_) );
  INV_X1 g673 ( .A(new_n808_), .ZN(new_n811_) );
  NAND2_X1 g674 ( .A1(new_n811_), .A2(new_n810_), .ZN(new_n812_) );
  NAND2_X1 g675 ( .A1(new_n812_), .A2(new_n809_), .ZN(new_n813_) );
  NAND3_X1 g676 ( .A1(new_n813_), .A2(new_n338_), .A3(new_n589_), .ZN(new_n814_) );
  NAND2_X1 g677 ( .A1(new_n814_), .A2(G169GAT), .ZN(new_n815_) );
  NAND4_X1 g678 ( .A1(new_n813_), .A2(new_n311_), .A3(new_n338_), .A4(new_n589_), .ZN(new_n816_) );
  NAND2_X1 g679 ( .A1(new_n815_), .A2(new_n816_), .ZN(G1348GAT) );
  NAND3_X1 g680 ( .A1(new_n813_), .A2(new_n338_), .A3(new_n666_), .ZN(new_n818_) );
  INV_X1 g681 ( .A(KEYINPUT57), .ZN(new_n819_) );
  NOR2_X1 g682 ( .A1(new_n819_), .A2(KEYINPUT56), .ZN(new_n820_) );
  NAND2_X1 g683 ( .A1(new_n819_), .A2(KEYINPUT56), .ZN(new_n821_) );
  INV_X1 g684 ( .A(new_n821_), .ZN(new_n822_) );
  NOR2_X1 g685 ( .A1(new_n822_), .A2(new_n820_), .ZN(new_n823_) );
  INV_X1 g686 ( .A(new_n823_), .ZN(new_n824_) );
  NAND2_X1 g687 ( .A1(new_n818_), .A2(new_n824_), .ZN(new_n825_) );
  NAND4_X1 g688 ( .A1(new_n813_), .A2(new_n338_), .A3(new_n666_), .A4(new_n823_), .ZN(new_n826_) );
  NAND2_X1 g689 ( .A1(new_n825_), .A2(new_n826_), .ZN(new_n827_) );
  NAND2_X1 g690 ( .A1(new_n827_), .A2(G176GAT), .ZN(new_n828_) );
  NAND3_X1 g691 ( .A1(new_n825_), .A2(new_n294_), .A3(new_n826_), .ZN(new_n829_) );
  NAND2_X1 g692 ( .A1(new_n828_), .A2(new_n829_), .ZN(G1349GAT) );
  NAND3_X1 g693 ( .A1(new_n813_), .A2(new_n338_), .A3(new_n507_), .ZN(new_n831_) );
  NAND2_X1 g694 ( .A1(new_n831_), .A2(G183GAT), .ZN(new_n832_) );
  NAND4_X1 g695 ( .A1(new_n813_), .A2(new_n295_), .A3(new_n338_), .A4(new_n507_), .ZN(new_n833_) );
  NAND2_X1 g696 ( .A1(new_n832_), .A2(new_n833_), .ZN(G1350GAT) );
  INV_X1 g697 ( .A(new_n449_), .ZN(new_n835_) );
  NAND3_X1 g698 ( .A1(new_n813_), .A2(new_n338_), .A3(new_n835_), .ZN(new_n836_) );
  NAND2_X1 g699 ( .A1(G190GAT), .A2(KEYINPUT58), .ZN(new_n837_) );
  INV_X1 g700 ( .A(new_n837_), .ZN(new_n838_) );
  NOR2_X1 g701 ( .A1(G190GAT), .A2(KEYINPUT58), .ZN(new_n839_) );
  NOR2_X1 g702 ( .A1(new_n838_), .A2(new_n839_), .ZN(new_n840_) );
  INV_X1 g703 ( .A(new_n840_), .ZN(new_n841_) );
  NAND2_X1 g704 ( .A1(new_n836_), .A2(new_n841_), .ZN(new_n842_) );
  NAND4_X1 g705 ( .A1(new_n813_), .A2(new_n338_), .A3(new_n835_), .A4(new_n840_), .ZN(new_n843_) );
  NAND2_X1 g706 ( .A1(new_n842_), .A2(new_n843_), .ZN(G1351GAT) );
  NAND3_X1 g707 ( .A1(new_n807_), .A2(new_n216_), .A3(new_n805_), .ZN(new_n845_) );
  INV_X1 g708 ( .A(new_n845_), .ZN(new_n846_) );
  NAND2_X1 g709 ( .A1(new_n846_), .A2(new_n388_), .ZN(new_n847_) );
  INV_X1 g710 ( .A(new_n847_), .ZN(new_n848_) );
  NAND2_X1 g711 ( .A1(new_n848_), .A2(new_n589_), .ZN(new_n849_) );
  NAND2_X1 g712 ( .A1(KEYINPUT60), .A2(KEYINPUT59), .ZN(new_n850_) );
  INV_X1 g713 ( .A(new_n850_), .ZN(new_n851_) );
  NOR2_X1 g714 ( .A1(KEYINPUT60), .A2(KEYINPUT59), .ZN(new_n852_) );
  NOR2_X1 g715 ( .A1(new_n851_), .A2(new_n852_), .ZN(new_n853_) );
  INV_X1 g716 ( .A(new_n853_), .ZN(new_n854_) );
  NAND2_X1 g717 ( .A1(new_n849_), .A2(new_n854_), .ZN(new_n855_) );
  NAND3_X1 g718 ( .A1(new_n848_), .A2(new_n589_), .A3(new_n853_), .ZN(new_n856_) );
  NAND2_X1 g719 ( .A1(new_n855_), .A2(new_n856_), .ZN(new_n857_) );
  NAND2_X1 g720 ( .A1(new_n857_), .A2(new_n219_), .ZN(new_n858_) );
  NAND3_X1 g721 ( .A1(new_n855_), .A2(G197GAT), .A3(new_n856_), .ZN(new_n859_) );
  NAND2_X1 g722 ( .A1(new_n858_), .A2(new_n859_), .ZN(G1352GAT) );
  NOR2_X1 g723 ( .A1(new_n847_), .A2(new_n546_), .ZN(new_n861_) );
  NAND2_X1 g724 ( .A1(G204GAT), .A2(KEYINPUT61), .ZN(new_n862_) );
  INV_X1 g725 ( .A(new_n862_), .ZN(new_n863_) );
  NOR2_X1 g726 ( .A1(G204GAT), .A2(KEYINPUT61), .ZN(new_n864_) );
  NOR2_X1 g727 ( .A1(new_n863_), .A2(new_n864_), .ZN(new_n865_) );
  INV_X1 g728 ( .A(new_n865_), .ZN(new_n866_) );
  NAND2_X1 g729 ( .A1(new_n861_), .A2(new_n866_), .ZN(new_n867_) );
  INV_X1 g730 ( .A(new_n861_), .ZN(new_n868_) );
  NAND2_X1 g731 ( .A1(new_n868_), .A2(new_n865_), .ZN(new_n869_) );
  NAND2_X1 g732 ( .A1(new_n869_), .A2(new_n867_), .ZN(G1353GAT) );
  NOR2_X1 g733 ( .A1(new_n847_), .A2(new_n506_), .ZN(new_n871_) );
  INV_X1 g734 ( .A(new_n871_), .ZN(new_n872_) );
  NAND2_X1 g735 ( .A1(new_n872_), .A2(G211GAT), .ZN(new_n873_) );
  NAND2_X1 g736 ( .A1(new_n871_), .A2(new_n222_), .ZN(new_n874_) );
  NAND2_X1 g737 ( .A1(new_n873_), .A2(new_n874_), .ZN(G1354GAT) );
  INV_X1 g738 ( .A(KEYINPUT62), .ZN(new_n876_) );
  NAND2_X1 g739 ( .A1(new_n848_), .A2(new_n625_), .ZN(new_n877_) );
  NAND2_X1 g740 ( .A1(new_n877_), .A2(new_n876_), .ZN(new_n878_) );
  NAND3_X1 g741 ( .A1(new_n848_), .A2(KEYINPUT62), .A3(new_n625_), .ZN(new_n879_) );
  NAND2_X1 g742 ( .A1(new_n878_), .A2(new_n879_), .ZN(new_n880_) );
  NAND2_X1 g743 ( .A1(new_n880_), .A2(new_n220_), .ZN(new_n881_) );
  NAND3_X1 g744 ( .A1(new_n878_), .A2(G218GAT), .A3(new_n879_), .ZN(new_n882_) );
  NAND2_X1 g745 ( .A1(new_n881_), .A2(new_n882_), .ZN(G1355GAT) );
endmodule


