module s38584 ( CK, g100, g10122, g10306, g10500, g10527, g113, g11349, g11388, 
        g114, g11418, g11447, g115, g116, g11678, g11770, g120, g12184, g12238, 
        g12300, g12350, g12368, g124, g12422, g12470, g125, g126, g127, g12832, 
        g12833, g12919, g12923, g13039, g13049, g13068, g13085, g13099, g13259, 
        g13272, g134, g135, g13865, g13881, g13895, g13906, g13926, g13966, 
        g14096, g14125, g14147, g14167, g14189, g14201, g14217, g14421, g14451, 
        g14518, g14597, g14635, g14662, g14673, g14694, g14705, g14738, g14749, 
        g14779, g14828, g16603, g16624, g16627, g16656, g16659, g16686, g16693, 
        g16718, g16722, g16744, g16748, g16775, g16874, g16924, g16955, g17291, 
        g17316, g17320, g17400, g17404, g17423, g17519, g17577, g17580, g17604, 
        g17607, g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711, 
        g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787, g17813, 
        g17819, g17845, g17871, g18092, g18094, g18095, g18096, g18097, g18098, 
        g18099, g18100, g18101, g18881, g19334, g19357, g20049, g20557, g20652, 
        g20654, g20763, g20899, g20901, g21176, g21245, g21270, g21292, g21698, 
        g21727, g23002, g23190, g23612, g23652, g23683, g23759, g24151, g24161, 
        g24162, g24163, g24164, g24165, g24166, g24167, g24168, g24169, g24170, 
        g24171, g24172, g24173, g24174, g24175, g24176, g24177, g24178, g24179, 
        g24180, g24181, g24182, g24183, g24184, g24185, g25114, g25167, g25219, 
        g25259, g25582, g25583, g25584, g25585, g25586, g25587, g25588, g25589, 
        g25590, g26801, g26875, g26876, g26877, g27831, g28030, g28041, g28042, 
        g28753, g29210, g29211, g29212, g29213, g29214, g29215, g29216, g29217, 
        g29218, g29219, g29220, g29221, g30327, g30329, g30330, g30331, g30332, 
        g31521, g31656, g31665, g31793, g31860, g31861, g31862, g31863, g32185, 
        g32429, g32454, g32975, g33079, g33435, g33533, g33636, g33659, g33874, 
        g33894, g33935, g33945, g33946, g33947, g33948, g33949, g33950, g33959, 
        g34201, g34221, g34232, g34233, g34234, g34235, g34236, g34237, g34238, 
        g34239, g34240, g34383, g34425, g34435, g34436, g34437, g34597, g34788, 
        g34839, g34913, g34915, g34917, g34919, g34921, g34923, g34925, g34927, 
        g34956, g34972, g35, g36, g44, g5, g53, g54, g56, g57, g64, g6744, 
        g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6752, g6753, g72, 
        g7243, g7245, g7257, g7260, g73, g7540, g7916, g7946, g8132, g8178, 
        g8215, g8235, g8277, g8279, g8283, g8291, g8342, g8344, g8353, g8358, 
        g8398, g84, g8403, g8416, g8475, g8719, g8783, g8784, g8785, g8786, 
        g8787, g8788, g8789, g8839, g8870, g8915, g8916, g8917, g8918, g8919, 
        g8920, g90, g9019, g9048, g91, g92, g9251, g9497, g9553, g9555, g9615, 
        g9617, g9680, g9682, g9741, g9743, g9817, g99, test_se, test_si1, 
        test_so1, test_si2, test_so2, test_si3, test_so3, test_si4, test_so4, 
        test_si5, test_so5, test_si6, test_so6, test_si7, test_so7, test_si8, 
        test_so8, test_si9, test_so9, test_si10, test_so10, test_si11, 
        test_so11, test_si12, test_so12, test_si13, test_so13, test_si14, 
        test_so14, test_si15, test_so15, test_si16, test_so16, test_si17, 
        test_so17, test_si18, test_so18, test_si19, test_so19, test_si20, 
        test_so20, test_si21, test_so21, test_si22, test_so22, test_si23, 
        test_so23, test_si24, test_so24, test_si25, test_so25, test_si26, 
        test_so26, test_si27, test_so27, test_si28, test_so28, test_si29, 
        test_so29, test_si30, test_so30, test_si31, test_so31, test_si32, 
        test_so32, test_si33, test_so33, test_si34, test_so34, test_si35, 
        test_so35, test_si36, test_so36, test_si37, test_so37, test_si38, 
        test_so38, test_si39, test_so39, test_si40, test_so40, test_si41, 
        test_so41, test_si42, test_so42, test_si43, test_so43, test_si44, 
        test_so44, test_si45, test_so45, test_si46, test_so46, test_si47, 
        test_so47, test_si48, test_so48, test_si49, test_so49, test_si50, 
        test_so50, test_si51, test_so51, test_si52, test_so52, test_si53, 
        test_so53, test_si54, test_so54, test_si55, test_so55, test_si56, 
        test_so56, test_si57, test_so57, test_si58, test_so58, test_si59, 
        test_so59, test_si60, test_so60, test_si61, test_so61, test_si62, 
        test_so62, test_si63, test_so63, test_si64, test_so64, test_si65, 
        test_so65, test_si66, test_so66, test_si67, test_so67, test_si68, 
        test_so68, test_si69, test_so69, test_si70, test_so70, test_si71, 
        test_so71, test_si72, test_so72, test_si73, test_so73, test_si74, 
        test_so74, test_si75, test_so75, test_si76, test_so76, test_si77, 
        test_so77, test_si78, test_so78, test_si79, test_so79, test_si80, 
        test_so80, test_si81, test_so81, test_si82, test_so82, test_si83, 
        test_so83, test_si84, test_so84, test_si85, test_so85, test_si86, 
        test_so86, test_si87, test_so87, test_si88, test_so88, test_si89, 
        test_so89, test_si90, test_so90, test_si91, test_so91, test_si92, 
        test_so92, test_si93, test_so93, test_si94, test_so94, test_si95, 
        test_so95, test_si96, test_so96, test_si97, test_so97, test_si98, 
        test_so98, test_si99, test_so99, test_si100, test_so100 );
  input CK, g100, g113, g114, g115, g116, g120, g124, g125, g126, g127, g134,
         g135, g35, g36, g44, g5, g53, g54, g56, g57, g64, g6744, g6745, g6746,
         g6747, g6748, g6749, g6750, g6751, g6752, g6753, g72, g73, g84, g90,
         g91, g92, g99, test_se, test_si1, test_si2, test_si3, test_si4,
         test_si5, test_si6, test_si7, test_si8, test_si9, test_si10,
         test_si11, test_si12, test_si13, test_si14, test_si15, test_si16,
         test_si17, test_si18, test_si19, test_si20, test_si21, test_si22,
         test_si23, test_si24, test_si25, test_si26, test_si27, test_si28,
         test_si29, test_si30, test_si31, test_si32, test_si33, test_si34,
         test_si35, test_si36, test_si37, test_si38, test_si39, test_si40,
         test_si41, test_si42, test_si43, test_si44, test_si45, test_si46,
         test_si47, test_si48, test_si49, test_si50, test_si51, test_si52,
         test_si53, test_si54, test_si55, test_si56, test_si57, test_si58,
         test_si59, test_si60, test_si61, test_si62, test_si63, test_si64,
         test_si65, test_si66, test_si67, test_si68, test_si69, test_si70,
         test_si71, test_si72, test_si73, test_si74, test_si75, test_si76,
         test_si77, test_si78, test_si79, test_si80, test_si81, test_si82,
         test_si83, test_si84, test_si85, test_si86, test_si87, test_si88,
         test_si89, test_si90, test_si91, test_si92, test_si93, test_si94,
         test_si95, test_si96, test_si97, test_si98, test_si99, test_si100;
  output g10122, g10306, g10500, g10527, g11349, g11388, g11418, g11447,
         g11678, g11770, g12184, g12238, g12300, g12350, g12368, g12422,
         g12470, g12832, g12833, g12919, g12923, g13039, g13049, g13068,
         g13085, g13099, g13259, g13272, g13865, g13881, g13895, g13906,
         g13926, g13966, g14096, g14125, g14147, g14167, g14189, g14201,
         g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673,
         g14694, g14705, g14738, g14749, g14779, g14828, g16603, g16624,
         g16627, g16656, g16659, g16686, g16693, g16718, g16722, g16744,
         g16748, g16775, g16874, g16924, g16955, g17291, g17316, g17320,
         g17400, g17404, g17423, g17519, g17577, g17580, g17604, g17607,
         g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711,
         g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787,
         g17813, g17819, g17845, g17871, g18092, g18094, g18095, g18096,
         g18097, g18098, g18099, g18100, g18101, g18881, g19334, g19357,
         g20049, g20557, g20652, g20654, g20763, g20899, g20901, g21176,
         g21245, g21270, g21292, g21698, g21727, g23002, g23190, g23612,
         g23652, g23683, g23759, g24151, g24161, g24162, g24163, g24164,
         g24165, g24166, g24167, g24168, g24169, g24170, g24171, g24172,
         g24173, g24174, g24175, g24176, g24177, g24178, g24179, g24180,
         g24181, g24182, g24183, g24184, g24185, g25114, g25167, g25219,
         g25259, g25582, g25583, g25584, g25585, g25586, g25587, g25588,
         g25589, g25590, g26801, g26875, g26876, g26877, g27831, g28030,
         g28041, g28042, g28753, g29210, g29211, g29212, g29213, g29214,
         g29215, g29216, g29217, g29218, g29219, g29220, g29221, g30327,
         g30329, g30330, g30331, g30332, g31521, g31656, g31665, g31793,
         g31860, g31861, g31862, g31863, g32185, g32429, g32454, g32975,
         g33079, g33435, g33533, g33636, g33659, g33874, g33894, g33935,
         g33945, g33946, g33947, g33948, g33949, g33950, g33959, g34201,
         g34221, g34232, g34233, g34234, g34235, g34236, g34237, g34238,
         g34239, g34240, g34383, g34425, g34435, g34436, g34437, g34597,
         g34788, g34839, g34913, g34915, g34917, g34919, g34921, g34923,
         g34925, g34927, g34956, g34972, g7243, g7245, g7257, g7260, g7540,
         g7916, g7946, g8132, g8178, g8215, g8235, g8277, g8279, g8283, g8291,
         g8342, g8344, g8353, g8358, g8398, g8403, g8416, g8475, g8719, g8783,
         g8784, g8785, g8786, g8787, g8788, g8789, g8839, g8870, g8915, g8916,
         g8917, g8918, g8919, g8920, g9019, g9048, g9251, g9497, g9553, g9555,
         g9615, g9617, g9680, g9682, g9741, g9743, g9817, test_so1, test_so2,
         test_so3, test_so4, test_so5, test_so6, test_so7, test_so8, test_so9,
         test_so10, test_so11, test_so12, test_so13, test_so14, test_so15,
         test_so16, test_so17, test_so18, test_so19, test_so20, test_so21,
         test_so22, test_so23, test_so24, test_so25, test_so26, test_so27,
         test_so28, test_so29, test_so30, test_so31, test_so32, test_so33,
         test_so34, test_so35, test_so36, test_so37, test_so38, test_so39,
         test_so40, test_so41, test_so42, test_so43, test_so44, test_so45,
         test_so46, test_so47, test_so48, test_so49, test_so50, test_so51,
         test_so52, test_so53, test_so54, test_so55, test_so56, test_so57,
         test_so58, test_so59, test_so60, test_so61, test_so62, test_so63,
         test_so64, test_so65, test_so66, test_so67, test_so68, test_so69,
         test_so70, test_so71, test_so72, test_so73, test_so74, test_so75,
         test_so76, test_so77, test_so78, test_so79, test_so80, test_so81,
         test_so82, test_so83, test_so84, test_so85, test_so86, test_so87,
         test_so88, test_so89, test_so90, test_so91, test_so92, test_so93,
         test_so94, test_so95, test_so96, test_so97, test_so98, test_so99,
         test_so100;
  wire   g100, g113, g114, g115, g116, g120, g124, g125, g126, g127, g134,
         g135, g18881, g23612, g23652, g73, g29211, g29212, g29213, g29214,
         g29215, g29216, g29217, g29219, g29220, g29221, g30327, g30331,
         g30332, g31656, g31665, g33533, g34435, g34788, g34839, g36, g44, g53,
         g54, g56, g57, g64, g6744, g6745, g6746, g6747, g6748, g6749, g6750,
         g6751, g6753, g84, g90, g91, g92, g99, test_so10, test_so26,
         test_so35, test_so39, test_so42, test_so44, test_so46, test_so80,
         test_so86, test_so92, test_so100, g34783, n2730, n4836, n4896, n4895,
         n4837, n4921, n4920, n2787, n4411, n5045, g559, n4959, g33046, g5057,
         n5615, g34441, g2771, n5544, g33982, g1882, n5854, g34007, g2299,
         g24276, g4040, n5530, g30381, g2547, n5782, g30405, g3243, g452,
         g30416, g3542, g30466, g5232, g25736, g5813, g34617, g33974, g1744,
         n5795, g30505, g5909, g33554, g1802, n5536, g30432, g3554, g33064,
         g6219, n5385, g34881, g807, n5479, g6031, g24216, g847, n5709, g24232,
         n9367, DFF_24_n1, g34733, g4172, g34882, g4372, g33026, g3512, g31867,
         n5471, g3490, n5454, g24344, n5432, g4235, g33966, g1600, n5811,
         g33550, g1714, n5460, g30393, g3155, n5366, g29248, g2236, g4571,
         g4555, g24274, g3698, g33973, g1736, n5817, g30360, g1968, n5664,
         g34460, g30494, g5607, g30384, g2657, n5316, g24340, n5439, g29223,
         g490, n5708, g26881, g311, n5317, g34252, g772, n5334, g30489, g5587,
         g29301, g6177, n5874, g6377, g33022, g3167, n5652, g30496, g5615,
         g33043, g4567, g29263, g30533, g6287, g24256, n5302, g34015, g2563,
         n5816, g34031, g4776, n5707, g34452, g4593, n5303, g34646, g6199,
         n5644, g34001, g2295, n5815, g25633, g1384, g24259, g1339, g33049,
         g5180, n5384, g34609, g2844, g31869, g1024, g30490, g30427, g3598,
         g21894, g4264, n5823, g33965, g767, n5333, g34645, g5853, n5499,
         n5580, g33571, g2089, g34267, g4933, n5878, g26971, g4521, n5752,
         g34644, g5507, n5643, g30534, g6291, g33535, g294, n5680, g30498,
         g25728, n5722, g25743, g25684, g3813, g25613, g562, g34438, g608,
         n5475, g24244, g1205, n5547, g30439, g3909, g30541, g6259, g30519,
         g5905, g25621, g921, g34807, g2955, g25599, g203, g24235, g34036,
         g4878, n5283, g30476, g5204, g30429, g3606, g32997, g1926, n5510,
         g33063, g6215, n5651, g30424, g3586, g32977, g291, n5679, g34026,
         g4674, n5440, g30420, g3570, g33560, g29226, g676, n5751, g25619,
         g843, g34455, g4332, n5540, g30457, g4153, g33625, g6336, n5592,
         g34790, g622, n5672, g30414, g3506, n5576, g26966, g4558, g25656,
         g3111, g30390, g25688, g34727, g939, n5415, g25594, g278, n5627,
         g26963, g4492, g34034, g4864, n5318, g33541, g1036, g28093, g24236,
         g1178, g30404, g3239, g28051, g718, g29303, g6195, g26917, g1135,
         n5328, g33624, g6395, n5396, g24337, g34911, g554, g33963, g496,
         g34627, g3853, n5641, g29282, g5134, n5807, g25676, n5721, g33013,
         g2485, n5509, g32981, g925, n5725, g34976, n9357, g30483, g5555,
         g32994, g1798, n5833, g28070, g34806, g2941, g30453, g3905, g33539,
         g763, n5332, g30526, g6255, g4375, g34035, g4871, n5443, g34636,
         g4722, g32978, g590, n5472, g30348, g1632, n5836, g24336, n5438,
         g3100, g24250, g29236, g1437, n5696, g29298, g6154, n5747, g1579,
         g30499, g5567, g33976, g1752, n5797, g32996, g1917, g30335, g744,
         n5470, g34637, g4737, n5867, g25694, g30528, g6267, g24251, g1442,
         g30521, g26960, g4477, n5849, g24239, g34259, g4643, n5382, g30474,
         g5264, n5703, g33016, g2610, g34643, g5160, n5498, g30510, g5933,
         g29239, g1454, n5866, g26897, g753, g34729, g1296, g34625, g3151,
         n5495, g34800, g24353, g6727, n5531, g33029, g3530, n5569, g33615,
         g4104, g24253, g1532, g24281, g33997, n9352, g34971, n9351, g34263,
         g4754, n5877, g24237, g1189, n5642, g33584, g2287, n5353, g24280,
         g4273, n5764, g26920, g1389, g33548, g29296, g5835, n5663, g30338,
         g1171, n5363, g21895, g4269, n5763, g2399, n5762, g34041, g4983,
         n5367, g30495, g5611, g29279, g4572, g25655, g3143, n5882, g34795,
         g2898, g24269, g3343, g30403, g3235, g33042, g30419, g3566, g34023,
         n9348, DFF_228_n1, g28090, g4961, n5770, g34642, g4927, n5879, g30370,
         g2259, n5419, g34448, g2819, n5609, g26946, g5802, g34610, g2852,
         g24209, g417, n5358, g28047, g681, g24206, g437, g26891, g30504,
         g5901, g34798, g2886, g25669, g3494, n5889, g30480, g5511, n5575,
         g33027, g3518, n5645, g33972, g1604, g25697, g5092, g28099, g4831,
         g26947, g4382, n5714, g24350, g6386, g24210, g479, g30455, g3965,
         g28084, g33993, g2008, g736, g30444, g3933, g33537, g222, g25650,
         g3050, g25625, g1052, g30366, g2122, n5784, g33593, g2465, n5523,
         g30502, g5889, g33036, g4495, g25595, g34462, g33024, g3179, n5390,
         g33552, g1728, n5352, g34014, g2433, g29273, g3835, n5662, g6187,
         n5453, g34638, g4917, n5408, g30341, g1070, g26899, g822, n5422,
         g30336, g914, n5560, g5339, g26940, g4164, g25622, g34447, g2807,
         n5379, g33613, g4054, n5395, g25749, g6191, n5888, g25704, g5077,
         n5455, g33053, g5523, n5647, g3680, g30555, g6637, g25601, g174,
         n5402, g33971, g1682, g26892, g355, g1087, g26915, g1105, n5478,
         g33008, g30538, g6307, g3802, g25750, g6159, g30369, g2255, n5414,
         g34446, g2815, n5404, g29230, g911, n5559, g43, g33975, g1748, g30497,
         g5551, g30418, g3558, g25721, g5499, g34622, g30438, g3901, g34266,
         g4888, n5863, g30540, g6251, g32986, g1373, g25648, n5723, g33960,
         g157, n5678, g34442, g2783, n5403, g4281, g30421, g3574, g33573,
         g2112, n5848, g34730, g1283, n5635, g24205, g10122_Tj, g4297, n5698,
         g32979, g758, n5331, g34025, g4639, n5727, g25763, g6537, g30481,
         g5543, g30517, g5961, g30539, g6243, g34880, n9340, g24242, n5654,
         g30436, g29265, g3476, n5786, g32990, g1664, n5407, g24245, g1246,
         n5756, g30553, g6629, g26907, g246, n6008, g24278, g4049, g26955,
         g24282, g2932, g4575, g31894, g4098, n5350, g33037, g4498, g26894,
         g528, n5327, g34977, n5477, g3139, n5447, g33962, g34451, g4584,
         n5539, g34250, g142, n5724, g29295, g5831, g26905, g239, g25629,
         g1216, n5442, g34792, g2848, g25703, g5022, g32983, g1030, g30402,
         g3231, g25757, g1430, n9336, g33999, g2241, g24262, g1564, g25729,
         g6148, g30558, g6649, g34781, g110, g26901, g225, n5597, g26961,
         g33039, g4504, g33059, g5873, n5388, g31899, g5037, n5611, g33007,
         g2319, n5375, g5495, n5446, g21891, g30462, g5208, g30487, g5579,
         g33058, g5869, n5649, g24261, g1589, n5755, g25730, g5752, g30531,
         g6279, g30506, g34804, g2975, n5750, g25747, g6167, n5430, n5701,
         g33601, g2599, n5524, g26922, g1448, n5343, g29250, g2370, g30459,
         g5164, n5570, g1333, n5616, g33534, g153, n5677, g30543, g6549, n5571,
         g29275, g4087, n5480, g34030, g34980, g2984, n5842, g30451, g3961,
         g25627, g962, n5630, g34657, g101, g30552, g6625, g34979, n9332,
         g30337, g1018, g24254, g24277, g4045, g29237, g1467, n5693, g30378,
         g2461, n5840, g33019, n5300, g33623, g5990, n5589, g29235, g1256,
         n5558, g31902, g5029, n5601, g6519, n5806, g25689, g4169, n5729,
         g33978, g1816, g26970, g4369, g4578, g34253, g4459, n5765, g29272,
         g3831, n5872, g33595, g2514, g33610, g3288, g33589, g34605, g2145,
         g30350, g1700, n5417, g25611, g513, g2841, n5963, g33619, g5297,
         n5588, g34022, g2763, g34033, g4793, n5368, g34726, g952, g31870,
         g1263, n5674, g33985, g1950, g29283, g5138, n5871, g34003, g2307,
         g25677, g34463, g4664, g33006, g2223, n5406, g29292, g5808, n5749,
         g30557, g6645, g33989, g2016, g33033, g3873, n5387, n5699, g34005,
         g2315, n5802, g26932, g2811, g30516, g5957, g33575, g2047, n5831,
         g33032, g30486, g5575, g34974, n9327, g25678, g3752, g30440, g3917,
         DFF_480_n1, g1585, n5757, g26949, g4388, g30530, g6275, g30542, g6311,
         g25624, g1041, g30383, g33597, g2537, n5411, g34598, g26957, g4430,
         g26967, n9325, g28102, g4826, g30524, g6239, g26903, g232, g30475,
         g5268, g34647, g6545, n5497, g30377, n9324, g33553, g1772, n5504,
         g31903, g5052, n5607, g25715, g33984, g1890, n5799, g33602, g2629,
         n5521, g28045, g572, n5337, g34603, g2130, n5487, g33035, g4108,
         g4308, g24208, g475, g990, n5622, g31, n5469, g34970, n9322, g33614,
         g3990, g33060, g30362, g1992, n5890, g33023, g3171, n5603, g26898,
         g812, n5733, g25618, g832, g30518, g5897, g4570, n5702, g26959, g4455,
         g34801, g2902, g26884, g333, g25600, g168, n5606, g26933, g28066,
         g3684, n5881, g33612, g3639, n5579, g24268, g3338, n5527, g25716,
         g5406, g26906, g269, g24203, g401, g24346, g6040, g24207, g441,
         g25701, n5690, g29269, g3808, n5745, g9, n5468, g34255, g30450, g3957,
         g30456, g4093, n5340, g32991, g1760, n5602, g24348, n5437, g34249,
         g160, n5843, g30371, g2279, n5778, g29268, g3498, g29224, g586, n5336,
         g33017, g2619, n5508, g30339, g1183, n5599, g33967, g1608, n5792,
         g33559, g1779, n5830, g2652, g30368, g2193, n5839, g30375, g2393,
         n5421, g28052, g661, g28089, g4950, n5772, g33055, g5535, n5566,
         g30392, g2834, g30343, g1361, g30523, g6235, g24233, g1146, n5851,
         g33018, g32976, g150, n5676, g30349, g1696, n5628, g33067, g6555,
         g26900, g33034, g3881, n5564, g30551, g6621, g25667, g3470, n5424,
         g30452, g3897, g34719, g518, g538, n5491, g33607, g2606, n5311,
         g26923, g1472, n5290, g24211, g33050, g5188, n5567, g24341, g5689,
         n5529, g24201, g405, g30463, g5216, g6494, g34464, g4669, g24243,
         g996, g24335, g4531, g34611, g2860, g34262, g4743, n5876, g30546,
         g6593, g25591, g4411, g30347, g1413, g30556, g6641, g6, g33562, g1936,
         n5534, g55, g25610, g504, n5519, g33015, g2587, n5372, g31896, g4480,
         g34004, n9314, g30428, g30485, g5571, g30422, g3578, g25714, g5827,
         n5809, g30423, g3582, g30529, g6271, g34028, g4688, n5656, g33587,
         g2380, g30460, g5196, g30401, g3227, g33990, n9312, g29309, g6541,
         g30411, g3203, g33546, g1668, n5598, g28085, g4760, n5775, g26904,
         g262, g1840, n5451, g25722, g5467, g25605, g460, g33062, g6209,
         g26893, n5704, g28050, g655, g33583, g2204, n5620, g30472, g5256,
         g34454, g4608, n5274, g34850, g794, n5291, n5583, g4423, g24272,
         g3689, n5532, g5685, g24214, g703, n5821, g26909, g862, n5682, g30406,
         g3247, g33569, g2040, g34628, g4146, n5981, g34458, g4633, n5844,
         g24240, n5304, g34634, g4732, n5296, g25700, n5689, g29293, g5817,
         g33009, g2351, n5511, g33603, g2648, g24355, g6736, g34268, g4944,
         n5875, g25691, g4072, g26890, g29264, g3466, g28072, g4116, g31900,
         g5041, n5605, g26956, g4434, g29271, g3827, n5808, g29304, g6500,
         n5748, g29261, g3133, n5661, g28063, g3333, g979, n5320, g34027,
         g4681, g33961, g298, n5675, g33604, g32995, g1894, n5374, g34624,
         g2988, g30415, g3538, g33536, g301, g26888, n9306, g28055, g827,
         n5728, g24238, g33600, g2555, n5351, g28105, g5011, g34721, g199,
         g29307, g6523, g30345, g34453, g4601, n5365, g32980, g854, n5754,
         g29238, g1484, n5865, g34639, g4922, n5346, g25695, g5080, n5893,
         g33057, g5863, g26969, g4581, n5670, g2518, g34021, g2567, g26895,
         g568, n5335, g30413, g3263, g30549, g6613, g24347, g25758, g6444,
         g34808, g2965, g30501, g5857, n5573, g33969, n9303, g34440, g890,
         n5305, g30433, g3562, g21900, g26921, g1404, g29270, g3817, n9302,
         n6010, g33038, g4501, g31865, g26926, g2724, n5301, g28083, g4704,
         n5771, g34797, g22, g2878, g30478, g5220, g34724, g617, n5339, g24212,
         g26883, g316, g32985, g1277, g25761, g6513, n5426, g26886, g336,
         n5824, g34796, g2882, g32982, g33561, g1906, n5503, g26880, g305,
         n5282, g34975, g8, g26931, g2799, g34641, g4912, n5297, g34629, g4157,
         n5983, g33598, g2541, n5461, g33576, g2153, n5356, g34720, g550,
         g26902, g255, g29244, g30468, g5240, g26924, g1478, n5289, g33031,
         g3863, g1959, g29266, g3480, n5868, g30559, g6653, g34794, g2864,
         g28087, g4894, n5774, g30435, g3857, n5572, g25609, g28057, g1002,
         g34439, g776, n5330, g28, n5324, g1236, g34260, g4646, n5712, g33012,
         g2476, g32989, g1657, n5525, g34006, g2375, g63, g358, g26910, g896,
         n5431, g33021, g3161, g2384, n5700, g34456, g4616, n5608, g26968,
         g4561, g33991, g2024, n5801, g3451, g26930, g2795, g34599, g613,
         n5474, g28082, g4527, g33557, g1844, n5847, g30511, g5937, g33045,
         g30379, g2523, n5281, g24267, n5436, g34020, g2643, g24249, g1489,
         n5850, g25592, g30382, n9295, g29285, g5156, n5526, n9294, g25662,
         n5717, g21896, g33563, g1955, g33622, g33582, g2273, n5458, n5584,
         g28086, g4771, n5769, g25744, g6098, g29262, g3147, g24270, g3347,
         g33581, g2269, n5410, g191, g24266, g2712, g34849, g626, n5288,
         g33618, g2729, g5357, n5393, g34038, g34032, g4709, n5518, g34803,
         g2927, g34459, g4340, n5653, g30509, g5929, g34640, g4907, n5295,
         g28069, g4035, g21899, g2946, g31868, g918, n5673, g26938, g4082,
         g25756, n5719, g30363, g30334, g577, n5294, g33970, g1620, n5791,
         g30391, g2831, g25615, g667, g33540, g930, n5731, g30445, g3937,
         g25617, g817, n5822, g24247, g1249, g24215, g837, n5562, g33964, g599,
         n5550, g25719, g5475, n5425, g29228, g30514, g5949, g33627, g6682,
         g24231, g904, g34615, g2873, n5488, g30356, g1854, n5785, g25696,
         g5084, n5681, g30493, g5603, n5726, g33594, g2495, n5522, g34009,
         g2437, n5789, g30365, g2102, n5666, g33004, g2208, g34018, g25685,
         g4064, n5416, g34040, g4899, n5517, g25639, g2719, n5465, g34029,
         g4785, n5361, g30488, g5583, g34600, g781, n5551, g29300, g6173,
         n5810, g34802, g2917, g25614, g686, g28058, g1252, n5554, g29225,
         g671, g33580, g30532, g6283, n5586, DFF_909_n1, g33054, g5527, n5389,
         g26962, g4489, g1974, n5450, g32984, g1270, n5716, g34039, g4966,
         n5706, g33065, g6227, n5568, g30443, g3929, g29291, g5503, g24279,
         g30508, g5925, g29232, g1124, n5692, g34269, g4955, n5614, g30464,
         g5224, g33988, g2012, n5790, g30522, g6203, n5574, g25708, g5120,
         g30374, g2389, n5631, g26953, g4438, g34008, g2429, n5814, g34444,
         g2787, n5610, g34731, g33606, g2675, n5457, g24334, n5541, g34265,
         g4836, n5713, g30340, g1199, g24257, g30482, g5547, g34604, g2138,
         n5275, g33591, g2338, n5310, g30525, g6247, g26929, g2791, g30448,
         g34602, g1291, n2549, g30513, g5945, g30469, g5244, g33608, g2759,
         g33626, g6741, n5398, g34725, g785, n5293, g30342, g1259, n5553,
         g29267, g3484, n5668, g25593, g209, n5595, g30548, g6609, g33052,
         g5517, g34012, g2449, n5798, g34017, n9281, g24263, g2715, n5299,
         g26912, g936, n5557, g30364, g2098, n5280, g34254, g4462, n5671,
         g34251, g604, n5473, g30560, g6589, g33983, n9280, g24204, g429,
         g33980, g1870, n5813, g34631, g1825, g25623, g1008, n5321, g26950,
         g4392, n5710, g30431, g3546, g30467, g5236, g30353, g1768, n5834,
         g34467, g4854, g30442, g3925, g29305, g6509, g25616, g732, n5732,
         g29252, g2504, g4519, g4520, g33003, g2185, n5376, g34613, g37, g4031,
         g33570, g2070, n5535, g34734, g4176, n5494, g24275, n5435, g4405,
         g872, g29302, g6181, n5667, g24349, g34264, g4765, n5613, g30484,
         g5563, g25634, g1395, g33567, g1913, n5828, g33585, g2331, n5513,
         g30527, g6263, g34978, n9276, g30447, g3945, g347, n5860, g34256,
         g4473, g25630, g1266, g29290, g5489, n5660, g29227, g31872, g2748,
         n5516, g29287, g5471, g31897, g4540, g6723, g30562, g6605, g34011,
         n9274, g33996, g2173, g21898, g33014, g2491, n5405, g34465, g4849,
         g33995, g2169, n5788, g30372, n9273, g30545, g30389, g33590, g2407,
         n5459, g34616, g2868, g26927, g2767, g32992, g1783, n5596, g25631,
         g1312, n5466, g30477, g5212, g34632, g4245, g28046, g645, g4291,
         g26896, n5657, g25602, g26916, g1129, n5329, g33578, g2227, n5538,
         g33579, g2246, g30354, g1830, n5413, g30425, g3590, g24200, g392,
         g33544, g1592, n5362, g25764, g6505, g24246, g1221, g30507, g5921,
         g26889, g30333, g218, g32998, g1932, n5829, g32987, g1624, n5370,
         g25702, g5062, g29286, g5462, n5744, g34606, g2689, n5347, g33070,
         g6573, n5563, g29240, g1677, g32999, g2028, n5371, g33605, g2671,
         n5278, g24255, g26945, g33558, g1848, n5464, g25699, n5669, g29289,
         g5485, g30388, g2741, n5349, n5482, g29254, g2638, g28074, g4122,
         g34450, g4322, n5506, g30512, g5941, g2108, n5452, g25, g33551,
         g33538, g595, n5476, g33005, g2217, n5512, g24248, n9267, DFF_1092_n1,
         g33002, g2066, n5832, g24234, g1152, n5618, g30471, g5252, g34000,
         g2165, g34016, g2571, n5787, g33048, g5176, n5650, n5581, g25628,
         g26934, g2827, g34468, g4859, g24202, g424, g33542, g1274, n5730,
         n9265, g34445, g2803, n5545, g33555, g1821, g34013, g2509, g28091,
         g5073, g26919, n5556, g30554, g6633, g29281, g5124, g30537, g6303,
         g28092, g5069, g34732, g2994, n5634, g28049, g650, g33545, g1636,
         n5549, g30441, g3921, g29247, g24354, g6732, g25636, g1306, n5796,
         g26914, g1061, g25670, g3462, g33998, g2181, n5803, g25626, g956,
         n5341, g33977, g1756, n5804, g29297, g5849, g28071, g4112, g30387,
         n9262, g33577, g2197, n5514, g33592, g26913, g1046, g28044, g482,
         n5820, g26948, g4401, g30344, g1514, n5364, g26885, g329, n5766,
         g33069, g6565, n5386, g34621, g2950, g28059, g1345, g6533, n5445,
         g34633, g4727, n5312, g24352, g26925, g1536, g30446, g3941, g25597,
         g370, g24342, g5694, g30357, g1858, n5892, g26908, g446, g30399,
         g3219, g29242, g1811, g30547, g6601, g34010, g2441, g33986, g1874,
         g34257, g30544, g6581, g30561, g6597, g5008, n5637, g30430, g3610,
         g34799, g2890, g33565, g1978, n5845, g33968, g1612, g34843, g112,
         g34793, g2856, g33566, g1982, n5462, g30465, g28073, g4119, g24351,
         g6390, g30346, g1542, g21893, g4258, g4818, g31904, g5033, g34635,
         g4717, n5344, g25637, g1554, n5768, g29274, g3849, g30396, g3199,
         g25735, g34037, g4975, n5360, g34791, g790, n5292, g30520, g5913,
         g30358, g1902, n5837, g29299, g6163, g25690, g4125, g28096, g4821,
         n5880, g28088, g4939, g24241, n5392, g30397, g3207, g4483, g30409,
         g29284, g5142, n5658, g30470, g5248, g30367, g2126, n5891, g24273,
         g3694, g5481, n5805, g30359, g1964, n5315, g25698, g5097, n5753,
         g30398, g3215, n9255, g26952, g4427, g26928, g2779, n5694, g26954,
         g30351, g1720, n5780, g31871, g1367, g5112, g19, g26939, g4145,
         g33994, g2161, n5812, g25596, g376, n5633, g33586, g2361, n5537,
         g21901, DFF_1234_n1, g31866, g582, n5552, g33000, g2051, g26918,
         g1193, g30373, g2327, n5841, g28056, g907, n5555, g34601, g947, n5286,
         g30355, g1834, n5665, g30426, g3594, g34805, g2999, g34002, g2303,
         n5794, g28053, g29229, g723, n5826, g33620, g5703, n5397, g34722,
         g546, n5492, g33599, g2472, n5619, g30515, g5953, g25649, g33979,
         g1740, g30417, g3550, g25683, g3845, g33574, g2116, n5463, n5582,
         g30410, g30454, g3913, g34024, g33547, g1687, g30386, g2681, n5777,
         g2533, n5761, g26887, g324, n5827, g34607, g2697, n5308, g31895,
         g4417, g33068, g6561, n5646, g29233, g1141, n5691, g24258, n5655,
         g30376, g33549, g1710, n5412, g29308, g6527, n5659, g30408, g3255,
         g1691, g34620, g2936, g33621, g5644, n5593, g25707, g5152, n5883,
         g24339, g5352, g34443, g2775, n5378, g34619, g2922, g29234, g30503,
         g5893, g30550, g6617, g33001, g2060, n5507, g33040, g4512, g30492,
         g5599, g25664, g3401, g26944, g4366, g34614, n5342, g29260, g3129,
         g33047, g5170, g24298, g25733, g5821, n5429, g30536, g6299, g29246,
         g2079, g34261, g4698, n5862, g33611, g3703, n5399, g25638, g1559,
         n5441, g34728, n9247, g29222, g411, n5629, g25742, n5718, g30449,
         g3953, g34608, g2704, n5377, g24345, g6035, n5528, n9245, g25635,
         g1300, n5483, g25686, g4057, n5711, g30461, g5200, g34466, g4843,
         g31901, g5046, n5578, g2250, g26882, n5456, g33041, g33011, g2453,
         n5373, g5841, n5449, n5705, g34618, g2912, g33010, g2357, n5276,
         g31864, g164, n5561, g34630, g4253, n5484, g31898, g5016, n5369,
         g25653, g3119, n5423, g25632, g1351, n5322, g32988, g33616, g29280,
         g5115, n5743, g33609, g3352, n5604, g30563, g6657, g33044, g4552,
         g30437, g3893, g30412, g3211, g30491, g5595, g30434, g3614, g34612,
         g29259, g3125, n5781, g25681, g3821, n5428, g25687, g4141, n5612,
         g33617, g30479, g5272, g29256, g2735, n5600, g28054, g728, g30535,
         g6295, g30385, g2661, n5418, g30361, g1988, n5783, g25705, g24260,
         g1548, n5546, g29257, g3106, n5742, g34461, g4659, g34258, g4358,
         n5348, g32993, g1792, n5359, g33992, g2084, g30394, g3187, g34449,
         g4311, n5323, g34019, g2583, n5800, g18597, n9240, DFF_1381_n1,
         g29231, g1094, n5697, g25682, g21897, g4284, g30395, g3191, g21892,
         g4239, g4180, n5380, g28048, g691, n5520, g34723, g534, n5490, g25598,
         g385, n5632, g33987, g2004, n5818, g30380, g2527, n5420, g5456,
         g26965, n6007, g25706, g30458, g4507, n5846, g24338, g5348, g30400,
         g3223, g34623, g2970, g24343, g5698, g30473, g5260, g24252, g1521,
         g33028, g3522, n5383, g29258, g3115, g30407, g3251, g26958, g34457,
         g33568, g1996, n5355, g25663, g26964, g4515, g34735, g4300, n5639,
         g30352, n9236, g33543, g1379, g24271, n5433, g33981, g1878, n5793,
         g30500, g5619, g34649, g71, g29277, g25612, n5287, g28060, n2505,
         n2499, n2461, n3141, n3122, g72, n5960, n4689, n5961, n4708, n3593,
         n3589, n3595, n3574, n3570, n3576, n3517, n3513, n3519, n3628, n3624,
         n3630, n3555, n3551, n3557, n3646, n3642, n3648, n3536, n3532, n3538,
         n3611, n3607, n3613, n3006, n3765, n3505, n3525, n3635, n4888, n3550,
         n2595, n2527, n3524, n3005, n3623, n3549, n3007, n3569, n3606, n3588,
         n3165, n3799, n3033, n3622, n3587, n3586, n3605, n3604, n3568, n3567,
         n3548, n3512, n3511, n3531, n3530, n3641, n3640, n3131, n3111, n3907,
         n3773, n3807, n3950, n3841, n3983, n3874, n4014, n4537, n4201, n3745,
         n3684, n3274, n2982, n2706, n2649, n2556, n2509, n2487, n2427, n2423,
         n2421, n4173, n4191, n4388, n4210, n3479, n3951, n3404, n3774, n3424,
         n3842, n3414, n3808, n3444, n3908, n3489, n3984, n3434, n3875, n4015,
         n3914, n3406, n3780, n3481, n3957, n3848, n3491, n3990, n3416, n3814,
         n3881, n3502, n4022, n3501, n4027, n3407, n3785, n3482, n3962, n3427,
         n3853, n3437, n3886, n3417, n3819, n3492, n3995, n3447, n3919, n3682,
         n3272, n2980, n2704, n2647, n2554, n2507, n2485, n2425, n2419, n3743,
         n2405, n2760, n2552, n4946, n4198, n2404, n4962, n4948, n2726, n2727,
         n3195, n2774, n3116, n4945, n4525, n4518, n3281, n3277, n3276, n2989,
         n2991, n2710, n2707, n3174, n3362, n3676, n2644, n3146, n3115, n3833,
         n3023, n3933, n2601, n3664, n3662, n3673, n3671, n2607, n3506, n2790,
         n4490, n4178, n4514, n4196, n3736, n3741, n2598, n4814, n4519, n2594,
         n3084, n2590, n3125, n3105, n3145, n3164, n3910, n3776, n3877, n3810,
         n3953, n3986, n3844, n3770, n3904, n3804, n3947, n3838, n3980, n4020,
         n3945, n3836, n3768, n3869, n3978, n3802, n3902, n2422, n4037, n4034,
         n4039, n3972, n3969, n3929, n3926, n3863, n3860, n4003, n4002, n4032,
         n4035, n3797, n3792, n3790, n3795, n3891, n3893, n3827, n3826, n3896,
         n4007, n3931, n3793, n3924, n3831, n3829, n3927, n3974, n3898, n3970,
         n4000, n3865, n3861, n3824, n3894, n3967, n3858, n4005, n3395, n4956,
         n5026, n3941, n3733, n4798, n4805, n4175, n3734, n4193, n3739, n3738,
         n4721, n4523, n4524, n4526, n2573, n2577, n2563, n2567, n4938, n4940,
         n4913, n4915, n4714, n4516, n4517, n5111, n4819, n3730, n4305, n4283,
         n2608, n4447, n4448, n4402, n4403, n4425, n4436, n4437, n4391, n4392,
         n4379, n4380, n4414, n4415, n4458, n4459, n5016, n5014, n3064, n3065,
         n4535, n5112, n3675, counter_31, counter_30, counter_29, counter_28,
         counter_27, counter_26, counter_25, counter_24, counter_23,
         counter_22, counter_21, counter_20, counter_19, counter_18,
         counter_17, counter_16, counter_15, counter_14, counter_13,
         counter_12, counter_11, counter_10, counter_9, counter_8, counter_7,
         counter_6, counter_5, counter_4, counter_3, counter_2, counter_1,
         counter_0, carry_31, carry_30, carry_29, carry_28, carry_27, carry_26,
         carry_25, carry_24, carry_23, carry_22, carry_21, carry_20, carry_19,
         carry_18, carry_17, carry_16, carry_15, carry_14, carry_13, carry_12,
         carry_11, carry_10, carry_9, carry_8, carry_7, carry_6, carry_5,
         carry_4, carry_3, carry_2, N31, N5, N6, N7, N8, N9, N10, N11, N12,
         N13, N14, N15, N23, N24, N25, N26, N2, N3, N4, N16, N17, N18, N19,
         N20, N21, N22, N27, N28, N29, N30, N1, N32, n37, n87, n73, n86, n85,
         n84, n83, n82, n81, n80, n79, n78, n77, n76, n75, n74, n58, n59, n60,
         n61, n62, n63, n64, Trigger_out, n65, n66, n67, n68, n69, n70, n71,
         n72, n2, n4, n5, n15, n29, n35, n45, n55, n92, n95, n97, n103, n120,
         n128, n132, n136, n154, n176, g33959, n198, n201, n227, n268, n290,
         n293, n315, n403, n418, n422, n450, n466, n473, n479, n503, n524,
         n552, n571, n580, n582, n591, n609, n623, n643, n735, n751, n755,
         n792, n831, n832, n864, n956, n978, n1052, n1101, g25167, n1192,
         n1249, n1269, n1363, n1418, n1426, n1432, n1436, n1545, n1688, n1730,
         n1770, n10087, n10088, n10089, n10090, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10126, n10127, n10128, n10129, n10130, n10131,
         n10133, n10134, n10135, n10136, n10138, n10139, n10141, n10142,
         n10144, n10148, n10149, n10152, n10153, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10169, n10170, n10171, n10172, n10173, n10174, n10176, n10178,
         n10180, n10181, n10182, n10183, n10184, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10207, n10208, n10209, n10210, n10212, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10240, n10242, n10243, n10244,
         n10245, n10246, n10247, n10249, n10250, n10251, n10252, n10253,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10270, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10346, n10347, n10349,
         n10350, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10403, n10404, n10406, n10408, n10409,
         n10411, n10412, n10414, n10415, n10417, n10418, n10420, n10421,
         n10423, n10424, n10426, n10427, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10442,
         n10443, n10445, n10447, n10448, n10450, n10452, n10454, n10455,
         n10457, n10458, n10460, n10462, n10463, n10464, n10465, n10467,
         n10468, n10469, n10470, n10472, n10473, n10474, n10476, n10477,
         n10479, n10481, n10482, n10483, n10484, n10486, n10487, n10488,
         n10489, n10491, n10492, n10493, n10495, n10496, n10499, n10500,
         n10503, n10504, n10506, n10507, n10508, n10511, n10512, n10515,
         n10516, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10550, n10551, n10552,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10598, n10606, n10609, n10610,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, g32975, n10626, n10627,
         n10628, n10629, n10630, n10631, g31860, n10633, g31862, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
         n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
         n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667,
         n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675,
         n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
         n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
         n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
         n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
         n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
         n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723,
         n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
         n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739,
         n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
         n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
         n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
         n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
         n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
         n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
         n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
         n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
         n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
         n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
         n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
         n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
         n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867,
         n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
         n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915,
         n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
         n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
         n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955,
         n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963,
         n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
         n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
         n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987,
         n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
         n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
         n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011,
         n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
         n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027,
         n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035,
         n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
         n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051,
         n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059,
         n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
         n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075,
         n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099,
         n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107,
         n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115,
         n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123,
         n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131,
         n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
         n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147,
         n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155,
         n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163,
         n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171,
         n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179,
         n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187,
         n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195,
         n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203,
         n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
         n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
         n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227,
         n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235,
         n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243,
         n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251,
         n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259,
         n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267,
         n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275,
         n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
         n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291,
         n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299,
         n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307,
         n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315,
         n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323,
         n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331,
         n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339,
         n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347,
         n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355,
         n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363,
         n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371,
         n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379,
         n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387,
         n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395,
         n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403,
         n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411,
         n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419,
         n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427,
         n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435,
         n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443,
         n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451,
         n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459,
         n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467,
         n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475,
         n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483,
         n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491,
         n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499,
         n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507,
         n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515,
         n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523,
         n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531,
         n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539,
         n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547,
         n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555,
         n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563,
         n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571,
         n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579,
         n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587,
         n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595,
         n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603,
         n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611,
         n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619,
         n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627,
         n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635,
         n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643,
         n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651,
         n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659,
         n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
         n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675,
         n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683,
         n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691,
         n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699,
         n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707,
         n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715,
         n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723,
         n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731,
         n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739,
         n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747,
         n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755,
         n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763,
         n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771,
         n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779,
         n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787,
         n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795,
         n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803,
         n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811,
         n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819,
         n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827,
         n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835,
         n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843,
         n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851,
         n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859,
         n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
         n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
         n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883,
         n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891,
         n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
         n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
         n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915,
         n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
         n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
         n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
         n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947,
         n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
         n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
         n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971,
         n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
         n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987,
         n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995,
         n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
         n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
         n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019,
         n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
         n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
         n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043,
         n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
         n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059,
         n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067,
         n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075,
         n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
         n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091,
         n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
         n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
         n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115,
         n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123,
         n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
         n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139,
         n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
         n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
         n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
         n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
         n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
         n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
         n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
         n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211,
         n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
         n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
         n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
         n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
         n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323,
         n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331,
         n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
         n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
         n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
         n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
         n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
         n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379,
         n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
         n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
         n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
         n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
         n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
         n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
         n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467,
         n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475,
         n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483,
         n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
         n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499,
         n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507,
         n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515,
         n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523,
         n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
         n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579,
         n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
         n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595,
         n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
         n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611,
         n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619,
         n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627,
         n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635,
         n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643,
         n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651,
         n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
         n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667,
         n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
         n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683,
         n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691,
         n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699,
         n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
         n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715,
         n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
         n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
         n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739,
         n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
         n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755,
         n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763,
         n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771,
         n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779,
         n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787,
         n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795,
         n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
         n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811,
         n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
         n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827,
         n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835,
         n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843,
         n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851,
         n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859,
         n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
         n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875,
         n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883,
         n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
         n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899,
         n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907,
         n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915,
         n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923,
         n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931,
         n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939,
         n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947,
         n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955,
         n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
         n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971,
         n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979,
         n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987,
         n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995,
         n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003,
         n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011,
         n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019,
         n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027,
         n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
         n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043,
         n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051,
         n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059,
         n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067,
         n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075,
         n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083,
         n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091,
         n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099,
         n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107,
         n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115,
         n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123,
         n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131,
         n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139,
         n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147,
         n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155,
         n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163,
         n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171,
         n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179,
         n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187,
         n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195,
         n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203,
         n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211,
         n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
         n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227,
         n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
         n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243,
         n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
         n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259,
         n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267,
         n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275,
         n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283,
         n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291,
         n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299,
         n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
         n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315,
         n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323,
         n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331,
         n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339,
         n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347,
         n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
         n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
         n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371,
         n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
         n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387,
         n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395,
         n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403,
         n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411,
         n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419,
         n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427,
         n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435,
         n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443,
         n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
         n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459,
         n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467,
         n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475,
         n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483,
         n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491,
         n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499,
         n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507,
         n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515,
         n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523,
         n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531,
         n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539,
         n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547,
         n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555,
         n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563,
         n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
         n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
         n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
         n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
         n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603,
         n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611,
         n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619,
         n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627,
         n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635,
         n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643,
         n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
         n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659,
         n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
         n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675,
         n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683,
         n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
         n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699,
         n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
         n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
         n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
         n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747,
         n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
         n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763,
         n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771,
         n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
         n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
         n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
         n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803,
         n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
         n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
         n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
         n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843,
         n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
         n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
         n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
         n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875,
         n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
         n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891,
         n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
         n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
         n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
         n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
         n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947,
         n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
         n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963,
         n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
         n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979,
         n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987,
         n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995,
         n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
         n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011,
         n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019,
         n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
         n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035,
         n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043,
         n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051,
         n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059,
         n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067,
         n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
         n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083,
         n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091,
         n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
         n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107,
         n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
         n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123,
         n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131,
         n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139,
         n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
         n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
         n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163,
         n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171,
         n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
         n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187,
         n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195,
         n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203,
         n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211,
         n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
         n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227,
         n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235,
         n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
         n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251,
         n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
         n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267,
         n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275,
         n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283,
         n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
         n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299,
         n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307,
         n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
         n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323,
         n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331,
         n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339,
         n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347,
         n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355,
         n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
         n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371,
         n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
         n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
         n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395,
         n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403,
         n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411,
         n19412, n19413, n19414, n19415, n19416, n19417, n19418, U5116_n1,
         U5126_n1, U5127_n1, U5128_n1, U5129_n1, U5353_n1, U5355_n1, U5961_n1,
         U5962_n1, U5963_n1, U5964_n1, U5965_n1, U5966_n1, U5967_n1, U5968_n1,
         U6100_n1, U6211_n1, U6212_n1, U6213_n1, U6214_n1, U6215_n1, U6216_n1,
         U6217_n1, U6218_n1, U6279_n1, U6280_n1, U6281_n1, U6282_n1, U6283_n1,
         U6284_n1, U6285_n1, U6286_n1, U6287_n1, U6288_n1, U6289_n1, U6290_n1,
         U6291_n1, U6292_n1, U6338_n1, U6341_n1, U6342_n1, U6343_n1, U6344_n1,
         U6345_n1, U6346_n1, U6347_n1, U6348_n1, U6349_n1, U6350_n1, U6351_n1,
         U6352_n1, U6353_n1, U6354_n1, U6355_n1, U6356_n1, U6357_n1, U6358_n1,
         U6359_n1, U6360_n1, U6361_n1, U6362_n1, U6363_n1, U6364_n1, U6365_n1,
         U6366_n1, U6367_n1, U6368_n1, U6369_n1, U6370_n1, U6371_n1, U6372_n1,
         U6373_n1, U6374_n1, U6375_n1, U6417_n1, U6446_n1, U6465_n1, U6497_n1,
         U6523_n1, U6542_n1, U6552_n1, U6553_n1, U6554_n1, U6555_n1, U6556_n1,
         U6559_n1, U6560_n1, U6561_n1, U6570_n1, U6911_n1, U6912_n1, U6917_n1,
         U6926_n1, U6927_n1, U6929_n1, U6931_n1, U6932_n1, U6933_n1, U6934_n1,
         U6935_n1, U6936_n1, U6937_n1, U6938_n1, U6939_n1, U6940_n1, U6941_n1,
         U6944_n1, U6950_n1, U6954_n1, U6955_n1, U6956_n1, U6957_n1, U7174_n1,
         U7248_n1, U7249_n1, U7402_n1, U7405_n1, U7413_n1, U7416_n1, U7427_n1,
         U7438_n1, U7449_n1, U7455_n1, U7464_n1, U7467_n1, U7482_n1, U7492_n1,
         U7513_n1, U7516_n1, U7549_n1, U7561_n1, U7574_n1, U7577_n1, U7585_n1,
         U7595_n1, U7614_n1, U7621_n1, U7629_n1, U7636_n1, U7639_n1, U7649_n1,
         U7652_n1, U7668_n1, U7673_n1, U7690_n1, U7707_n1, U7712_n1, U7792_n1,
         U7794_n1, U7895_n1, U7897_n1, U7977_n1, U8034_n1, U8036_n1, U8050_n1,
         U8055_n1, U8060_n1, U8070_n1, U8074_n1, U8088_n1, U8112_n1, U8113_n1,
         U8147_n1, U8165_n1, U8185_n1, U8192_n1, U8210_n1, U8223_n1, U8224_n1,
         U8281_n1, U8307_n1, U8974_n1, U8975_n1, U9065_n1, U9070_n1, U9075_n1,
         U9076_n1, U9080_n1, U9084_n1, U9085_n1, U9086_n1, U9090_n1, U9098_n1,
         U9099_n1, U9101_n1, U9107_n1, U9111_n1, U9116_n1, U9120_n1, U9124_n1,
         U9128_n1, U9132_n1, U9136_n1, U9315_n1, U9453_n1, U9825_n1, U9886_n1,
         U9927_n1, U9953_n1, U9957_n1, U9958_n1, U9968_n1, U9972_n1, U9992_n1,
         U10314_n1, U10318_n1;
  assign g34240 = 1'b1;
  assign g34239 = 1'b1;
  assign g34238 = 1'b1;
  assign g34237 = 1'b1;
  assign g34236 = 1'b1;
  assign g34235 = 1'b1;
  assign g34234 = 1'b1;
  assign g34233 = 1'b1;
  assign g34232 = 1'b1;
  assign g33950 = 1'b1;
  assign g33949 = 1'b1;
  assign g33948 = 1'b1;
  assign g33947 = 1'b1;
  assign g33946 = 1'b1;
  assign g33945 = 1'b1;
  assign g32454 = 1'b1;
  assign g32429 = 1'b1;
  assign g25590 = 1'b1;
  assign g25589 = 1'b1;
  assign g25588 = 1'b1;
  assign g25587 = 1'b1;
  assign g25586 = 1'b1;
  assign g25585 = 1'b1;
  assign g25584 = 1'b1;
  assign g25583 = 1'b1;
  assign g25582 = 1'b1;
  assign g24151 = 1'b1;
  assign g34597 = 1'b0;
  assign g24173 = g100;
  assign g24174 = g113;
  assign g24175 = g114;
  assign g24176 = g115;
  assign g24177 = g116;
  assign g24178 = g120;
  assign g24179 = g124;
  assign g24180 = g125;
  assign g24181 = g126;
  assign g24182 = g127;
  assign g24183 = g134;
  assign g24184 = g135;
  assign g29218 = g18881;
  assign g30329 = g23612;
  assign g30330 = g23652;
  assign g24167 = g73;
  assign g20763 = g29211;
  assign g20899 = g29212;
  assign g20557 = g29213;
  assign g20652 = g29214;
  assign g20901 = g29215;
  assign g21176 = g29216;
  assign g21270 = g29217;
  assign g20654 = g29219;
  assign g21245 = g29220;
  assign g21292 = g29221;
  assign g23002 = g30327;
  assign g23759 = g30331;
  assign g23683 = g30332;
  assign g34436 = g31656;
  assign g34437 = g31665;
  assign g27831 = g33533;
  assign g31521 = g34435;
  assign g33894 = g34788;
  assign g34956 = g34839;
  assign g21698 = g36;
  assign g24185 = g44;
  assign g24161 = g53;
  assign g24162 = g54;
  assign g24163 = g56;
  assign g24164 = g57;
  assign g24165 = g64;
  assign g18098 = g6744;
  assign g18099 = g6745;
  assign g18101 = g6746;
  assign g18097 = g6747;
  assign g18094 = g6748;
  assign g18095 = g6749;
  assign g18096 = g6750;
  assign g18100 = g6751;
  assign g18092 = g6753;
  assign g24168 = g84;
  assign g24169 = g90;
  assign g24170 = g91;
  assign g24171 = g92;
  assign g24172 = g99;
  assign g31861 = test_so10;
  assign g25219 = test_so10;
  assign g13881 = test_so26;
  assign g9615 = test_so35;
  assign g8785 = test_so39;
  assign g8291 = test_so42;
  assign g17316 = test_so44;
  assign g8178 = test_so46;
  assign g12470 = test_so80;
  assign g11447 = test_so86;
  assign g9682 = test_so92;
  assign g29210 = test_so100;
  assign g20049 = test_so100;
  assign g24166 = g72;
  assign g28753 = g33959;
  assign g31863 = g25167;
  assign g26801 = g32975;
  assign g25114 = g31860;
  assign g25259 = g31862;

  SDFFX1 DFF_0_Q_reg ( .D(g33046), .SI(test_si1), .SE(n10699), .CLK(n11082), 
        .Q(g5057), .QN(n5615) );
  SDFFX1 DFF_1_Q_reg ( .D(g34441), .SI(g5057), .SE(n10792), .CLK(n11175), .Q(
        g2771), .QN(n5544) );
  SDFFX1 DFF_2_Q_reg ( .D(g33982), .SI(g2771), .SE(n10758), .CLK(n11141), .Q(
        g1882), .QN(n5854) );
  SDFFX1 DFF_4_Q_reg ( .D(g34007), .SI(g1882), .SE(n10792), .CLK(n11175), .Q(
        g2299), .QN(n10152) );
  SDFFX1 DFF_5_Q_reg ( .D(g24276), .SI(g2299), .SE(n10802), .CLK(n11185), .Q(
        g4040), .QN(n5530) );
  SDFFX1 DFF_6_Q_reg ( .D(g30381), .SI(g4040), .SE(n10717), .CLK(n11100), .Q(
        g2547), .QN(n5782) );
  SDFFX1 DFF_7_Q_reg ( .D(g9048), .SI(g2547), .SE(n10750), .CLK(n11133), .Q(
        g559) );
  SDFFX1 DFF_9_Q_reg ( .D(g30405), .SI(g559), .SE(n10719), .CLK(n11102), .Q(
        g3243), .QN(n10334) );
  SDFFX1 DFF_10_Q_reg ( .D(n29), .SI(g3243), .SE(n10732), .CLK(n11115), .Q(
        g452), .QN(n10404) );
  SDFFX1 DFF_12_Q_reg ( .D(g30416), .SI(g452), .SE(n10732), .CLK(n11115), .Q(
        g3542), .QN(n10298) );
  SDFFX1 DFF_13_Q_reg ( .D(g30466), .SI(g3542), .SE(n10740), .CLK(n11123), .Q(
        g5232), .QN(n10411) );
  SDFFX1 DFF_14_Q_reg ( .D(g25736), .SI(g5232), .SE(n10740), .CLK(n11123), .Q(
        g5813) );
  SDFFX1 DFF_15_Q_reg ( .D(g34617), .SI(g5813), .SE(n10740), .CLK(n11123), .Q(
        test_so1), .QN(n10675) );
  SDFFX1 DFF_16_Q_reg ( .D(g33974), .SI(test_si2), .SE(n10771), .CLK(n11154), 
        .Q(g1744), .QN(n5795) );
  SDFFX1 DFF_17_Q_reg ( .D(g30505), .SI(g1744), .SE(n10742), .CLK(n11125), .Q(
        g5909), .QN(n10415) );
  SDFFX1 DFF_18_Q_reg ( .D(g33554), .SI(g5909), .SE(n10771), .CLK(n11154), .Q(
        g1802), .QN(n5536) );
  SDFFX1 DFF_19_Q_reg ( .D(g30432), .SI(g1802), .SE(n10732), .CLK(n11115), .Q(
        g3554), .QN(n10488) );
  SDFFX1 DFF_20_Q_reg ( .D(g33064), .SI(g3554), .SE(n10777), .CLK(n11160), .Q(
        g6219), .QN(n5385) );
  SDFFX1 DFF_21_Q_reg ( .D(g34881), .SI(g6219), .SE(n10767), .CLK(n11150), .Q(
        g807), .QN(n5479) );
  SDFFX1 DFF_22_Q_reg ( .D(g17715), .SI(g807), .SE(n10767), .CLK(n11150), .Q(
        g6031) );
  SDFFX1 DFF_23_Q_reg ( .D(g24216), .SI(g6031), .SE(n10767), .CLK(n11150), .Q(
        g847), .QN(n5709) );
  SDFFX1 DFF_24_Q_reg ( .D(g24232), .SI(g847), .SE(n10751), .CLK(n11134), .Q(
        n9367), .QN(DFF_24_n1) );
  SDFFX1 DFF_25_Q_reg ( .D(g34733), .SI(n9367), .SE(n10739), .CLK(n11122), .Q(
        g4172) );
  SDFFX1 DFF_26_Q_reg ( .D(g34882), .SI(g4172), .SE(n10719), .CLK(n11102), .Q(
        g4372) );
  SDFFX1 DFF_27_Q_reg ( .D(g33026), .SI(g4372), .SE(n10720), .CLK(n11103), .Q(
        g3512), .QN(n10587) );
  SDFFX1 DFF_28_Q_reg ( .D(g31867), .SI(g3512), .SE(n10765), .CLK(n11148), .Q(
        test_so2), .QN(n5471) );
  SDFFX1 DFF_29_Q_reg ( .D(n120), .SI(test_si3), .SE(n10777), .CLK(n11160), 
        .Q(g3490), .QN(n5454) );
  SDFFX1 DFF_30_Q_reg ( .D(g24344), .SI(g3490), .SE(n10725), .CLK(n11108), .Q(
        g12350), .QN(n5432) );
  SDFFX1 DFF_31_Q_reg ( .D(g8920), .SI(g12350), .SE(n10791), .CLK(n11174), .Q(
        g4235), .QN(n10325) );
  SDFFX1 DFF_32_Q_reg ( .D(g33966), .SI(g4235), .SE(n10737), .CLK(n11120), .Q(
        g1600), .QN(n5811) );
  SDFFX1 DFF_33_Q_reg ( .D(g33550), .SI(g1600), .SE(n10723), .CLK(n11106), .Q(
        g1714), .QN(n5460) );
  SDFFX1 DFF_34_Q_reg ( .D(g16656), .SI(g1714), .SE(n10789), .CLK(n11172), .Q(
        g14451), .QN(n10515) );
  SDFFX1 DFF_35_Q_reg ( .D(g30393), .SI(g14451), .SE(n10789), .CLK(n11172), 
        .Q(g3155), .QN(n5366) );
  SDFFX1 DFF_37_Q_reg ( .D(g29248), .SI(g3155), .SE(n10707), .CLK(n11090), .Q(
        g2236), .QN(n10315) );
  SDFFX1 DFF_38_Q_reg ( .D(g4571), .SI(g2236), .SE(n10782), .CLK(n11165), .Q(
        g4555) );
  SDFFX1 DFF_39_Q_reg ( .D(g24274), .SI(g4555), .SE(n10747), .CLK(n11130), .Q(
        g3698), .QN(n10392) );
  SDFFX1 DFF_41_Q_reg ( .D(g33973), .SI(g3698), .SE(n10708), .CLK(n11091), .Q(
        g1736), .QN(n5817) );
  SDFFX1 DFF_42_Q_reg ( .D(g30360), .SI(g1736), .SE(n10758), .CLK(n11141), .Q(
        g1968), .QN(n5664) );
  SDFFX1 DFF_43_Q_reg ( .D(g34460), .SI(g1968), .SE(n10758), .CLK(n11141), .Q(
        test_so3), .QN(n10667) );
  SDFFX1 DFF_44_Q_reg ( .D(g30494), .SI(test_si4), .SE(n10706), .CLK(n11089), 
        .Q(g5607), .QN(n10364) );
  SDFFX1 DFF_45_Q_reg ( .D(g30384), .SI(g5607), .SE(n10706), .CLK(n11089), .Q(
        g2657), .QN(n5316) );
  SDFFX1 DFF_46_Q_reg ( .D(g24340), .SI(g2657), .SE(n10713), .CLK(n11096), .Q(
        g12300), .QN(n5439) );
  SDFFX1 DFF_47_Q_reg ( .D(g29223), .SI(g12300), .SE(n10771), .CLK(n11154), 
        .Q(g490), .QN(n5708) );
  SDFFX1 DFF_48_Q_reg ( .D(g26881), .SI(g490), .SE(n10772), .CLK(n11155), .Q(
        g311), .QN(n5317) );
  SDFFX1 DFF_50_Q_reg ( .D(g34252), .SI(g311), .SE(n10766), .CLK(n11149), .Q(
        g772), .QN(n5334) );
  SDFFX1 DFF_51_Q_reg ( .D(g30489), .SI(g772), .SE(n10705), .CLK(n11088), .Q(
        g5587), .QN(n10434) );
  SDFFX1 DFF_52_Q_reg ( .D(g29301), .SI(g5587), .SE(n10705), .CLK(n11088), .Q(
        g6177), .QN(n5874) );
  SDFFX1 DFF_53_Q_reg ( .D(g17743), .SI(g6177), .SE(n10787), .CLK(n11170), .Q(
        g6377) );
  SDFFX1 DFF_54_Q_reg ( .D(g33022), .SI(g6377), .SE(n10789), .CLK(n11172), .Q(
        g3167), .QN(n5652) );
  SDFFX1 DFF_55_Q_reg ( .D(g30496), .SI(g3167), .SE(n10721), .CLK(n11104), .Q(
        g5615), .QN(n10342) );
  SDFFX1 DFF_56_Q_reg ( .D(g33043), .SI(g5615), .SE(n10784), .CLK(n11167), .Q(
        g4567) );
  SDFFX1 DFF_58_Q_reg ( .D(g29263), .SI(g4567), .SE(n10720), .CLK(n11103), .Q(
        test_so4), .QN(n10658) );
  SDFFX1 DFF_59_Q_reg ( .D(g30533), .SI(test_si5), .SE(n10762), .CLK(n11145), 
        .Q(g6287), .QN(n10489) );
  SDFFX1 DFF_60_Q_reg ( .D(g24256), .SI(g6287), .SE(n10762), .CLK(n11145), .Q(
        g7946), .QN(n5302) );
  SDFFX1 DFF_61_Q_reg ( .D(g34015), .SI(g7946), .SE(n10748), .CLK(n11131), .Q(
        g2563), .QN(n5816) );
  SDFFX1 DFF_62_Q_reg ( .D(g34031), .SI(g2563), .SE(n10748), .CLK(n11131), .Q(
        g4776), .QN(n5707) );
  SDFFX1 DFF_63_Q_reg ( .D(g34452), .SI(g4776), .SE(n10768), .CLK(n11151), .Q(
        g4593), .QN(n5303) );
  SDFFX1 DFF_64_Q_reg ( .D(g34646), .SI(g4593), .SE(n10768), .CLK(n11151), .Q(
        g6199), .QN(n5644) );
  SDFFX1 DFF_65_Q_reg ( .D(g34001), .SI(g6199), .SE(n10768), .CLK(n11151), .Q(
        g2295), .QN(n5815) );
  SDFFX1 DFF_66_Q_reg ( .D(g25633), .SI(g2295), .SE(n10723), .CLK(n11106), .Q(
        g1384), .QN(n10105) );
  SDFFX1 DFF_67_Q_reg ( .D(g24259), .SI(g1384), .SE(n10748), .CLK(n11131), .Q(
        g1339) );
  SDFFX1 DFF_68_Q_reg ( .D(g33049), .SI(g1339), .SE(n10779), .CLK(n11162), .Q(
        g5180), .QN(n5384) );
  SDFFX1 DFF_69_Q_reg ( .D(g34609), .SI(g5180), .SE(n10743), .CLK(n11126), .Q(
        g2844) );
  SDFFX1 DFF_70_Q_reg ( .D(g31869), .SI(g2844), .SE(n10704), .CLK(n11087), .Q(
        g1024), .QN(n10230) );
  SDFFX1 DFF_71_Q_reg ( .D(g30490), .SI(g1024), .SE(n10706), .CLK(n11089), .Q(
        test_so5), .QN(n10688) );
  SDFFX1 DFF_72_Q_reg ( .D(g30427), .SI(test_si6), .SE(n10763), .CLK(n11146), 
        .Q(g3598), .QN(n10296) );
  SDFFX1 DFF_73_Q_reg ( .D(g21894), .SI(g3598), .SE(n10763), .CLK(n11146), .Q(
        g4264), .QN(n5823) );
  SDFFX1 DFF_74_Q_reg ( .D(g33965), .SI(g4264), .SE(n10766), .CLK(n11149), .Q(
        g767), .QN(n5333) );
  SDFFX1 DFF_75_Q_reg ( .D(g34645), .SI(g767), .SE(n10766), .CLK(n11149), .Q(
        g5853), .QN(n5499) );
  SDFFX1 DFF_76_Q_reg ( .D(g16874), .SI(g5853), .SE(n10766), .CLK(n11149), .Q(
        g13865), .QN(n5580) );
  SDFFX1 DFF_77_Q_reg ( .D(g33571), .SI(g13865), .SE(n10744), .CLK(n11127), 
        .Q(g2089), .QN(n10161) );
  SDFFX1 DFF_78_Q_reg ( .D(g34267), .SI(g2089), .SE(n10721), .CLK(n11104), .Q(
        g4933), .QN(n5878) );
  SDFFX1 DFF_79_Q_reg ( .D(g26971), .SI(g4933), .SE(n10719), .CLK(n11102), .Q(
        g4521), .QN(n5752) );
  SDFFX1 DFF_80_Q_reg ( .D(g34644), .SI(g4521), .SE(n10719), .CLK(n11102), .Q(
        g5507), .QN(n5643) );
  SDFFX1 DFF_81_Q_reg ( .D(g16627), .SI(g5507), .SE(n10789), .CLK(n11172), .Q(
        g16656), .QN(n10487) );
  SDFFX1 DFF_82_Q_reg ( .D(g30534), .SI(g16656), .SE(n10760), .CLK(n11143), 
        .Q(g6291), .QN(n10355) );
  SDFFX1 DFF_83_Q_reg ( .D(g33535), .SI(g6291), .SE(n10711), .CLK(n11094), .Q(
        g294), .QN(n5680) );
  SDFFX1 DFF_84_Q_reg ( .D(g30498), .SI(g294), .SE(n10805), .CLK(n11188), .Q(
        test_so6) );
  SDFFX1 DFF_85_Q_reg ( .D(g25728), .SI(test_si7), .SE(n10786), .CLK(n11169), 
        .Q(g9617), .QN(n5722) );
  SDFFX1 DFF_86_Q_reg ( .D(g25743), .SI(g9617), .SE(n10749), .CLK(n11132), .Q(
        g9741) );
  SDFFX1 DFF_87_Q_reg ( .D(g25684), .SI(g9741), .SE(n10749), .CLK(n11132), .Q(
        g3813) );
  SDFFX1 DFF_88_Q_reg ( .D(g25613), .SI(g3813), .SE(n10749), .CLK(n11132), .Q(
        g562), .QN(n10098) );
  SDFFX1 DFF_89_Q_reg ( .D(g34438), .SI(g562), .SE(n10750), .CLK(n11133), .Q(
        g608), .QN(n5475) );
  SDFFX1 DFF_90_Q_reg ( .D(g24244), .SI(g608), .SE(n10770), .CLK(n11153), .Q(
        g1205), .QN(n5547) );
  SDFFX1 DFF_91_Q_reg ( .D(g30439), .SI(g1205), .SE(n10731), .CLK(n11114), .Q(
        g3909), .QN(n10421) );
  SDFFX1 DFF_92_Q_reg ( .D(g30541), .SI(g3909), .SE(n10800), .CLK(n11183), .Q(
        g6259) );
  SDFFX1 DFF_93_Q_reg ( .D(g30519), .SI(g6259), .SE(n10741), .CLK(n11124), .Q(
        g5905), .QN(n10469) );
  SDFFX1 DFF_94_Q_reg ( .D(g25621), .SI(g5905), .SE(n10730), .CLK(n11113), .Q(
        g921) );
  SDFFX1 DFF_95_Q_reg ( .D(g34807), .SI(g921), .SE(n10699), .CLK(n11082), .Q(
        g2955), .QN(n10232) );
  SDFFX1 DFF_96_Q_reg ( .D(g25599), .SI(g2955), .SE(n10785), .CLK(n11168), .Q(
        g203) );
  SDFFX1 DFF_98_Q_reg ( .D(g24235), .SI(g203), .SE(n10757), .CLK(n11140), .Q(
        test_so7) );
  SDFFX1 DFF_99_Q_reg ( .D(g34036), .SI(test_si8), .SE(n10759), .CLK(n11142), 
        .Q(g4878), .QN(n5283) );
  SDFFX1 DFF_100_Q_reg ( .D(g30476), .SI(g4878), .SE(n10774), .CLK(n11157), 
        .Q(g5204) );
  SDFFX1 DFF_101_Q_reg ( .D(g17580), .SI(g5204), .SE(n10774), .CLK(n11157), 
        .Q(g17604), .QN(n10473) );
  SDFFX1 DFF_102_Q_reg ( .D(g30429), .SI(g17604), .SE(n10733), .CLK(n11116), 
        .Q(g3606), .QN(n10486) );
  SDFFX1 DFF_103_Q_reg ( .D(g32997), .SI(g3606), .SE(n10760), .CLK(n11143), 
        .Q(g1926), .QN(n5510) );
  SDFFX1 DFF_104_Q_reg ( .D(g33063), .SI(g1926), .SE(n10760), .CLK(n11143), 
        .Q(g6215), .QN(n5651) );
  SDFFX1 DFF_105_Q_reg ( .D(g30424), .SI(g6215), .SE(n10732), .CLK(n11115), 
        .Q(g3586), .QN(n10384) );
  SDFFX1 DFF_106_Q_reg ( .D(g32977), .SI(g3586), .SE(n10711), .CLK(n11094), 
        .Q(g291), .QN(n5679) );
  SDFFX1 DFF_107_Q_reg ( .D(g34026), .SI(g291), .SE(n10796), .CLK(n11179), .Q(
        g4674), .QN(n5440) );
  SDFFX1 DFF_108_Q_reg ( .D(g30420), .SI(g4674), .SE(n10732), .CLK(n11115), 
        .Q(g3570), .QN(n10332) );
  SDFFX1 DFF_109_Q_reg ( .D(g12368), .SI(g3570), .SE(n10750), .CLK(n11133), 
        .Q(g9048), .QN(n10088) );
  SDFFX1 DFF_110_Q_reg ( .D(g17739), .SI(g9048), .SE(n10759), .CLK(n11142), 
        .Q(g17607), .QN(n10361) );
  SDFFX1 DFF_111_Q_reg ( .D(g33560), .SI(g17607), .SE(n10797), .CLK(n11180), 
        .Q(test_so8), .QN(n10657) );
  SDFFX1 DFF_112_Q_reg ( .D(g29226), .SI(test_si9), .SE(n10709), .CLK(n11092), 
        .Q(g676), .QN(n5751) );
  SDFFX1 DFF_113_Q_reg ( .D(g25619), .SI(g676), .SE(n10767), .CLK(n11150), .Q(
        g843), .QN(n10216) );
  SDFFX1 DFF_115_Q_reg ( .D(g34455), .SI(g843), .SE(n10767), .CLK(n11150), .Q(
        g4332), .QN(n5540) );
  SDFFX1 DFF_116_Q_reg ( .D(g30457), .SI(g4332), .SE(n10739), .CLK(n11122), 
        .Q(g4153) );
  SDFFX1 DFF_117_Q_reg ( .D(g14694), .SI(g4153), .SE(n10739), .CLK(n11122), 
        .Q(g17711), .QN(n10378) );
  SDFFX1 DFF_118_Q_reg ( .D(g33625), .SI(g17711), .SE(n10704), .CLK(n11087), 
        .Q(g6336), .QN(n5592) );
  SDFFX1 DFF_119_Q_reg ( .D(g34790), .SI(g6336), .SE(n10750), .CLK(n11133), 
        .Q(g622), .QN(n5672) );
  SDFFX1 DFF_120_Q_reg ( .D(g30414), .SI(g622), .SE(n10777), .CLK(n11160), .Q(
        g3506), .QN(n5576) );
  SDFFX1 DFF_121_Q_reg ( .D(g26966), .SI(g3506), .SE(n10782), .CLK(n11165), 
        .Q(g4558) );
  SDFFX1 DFF_123_Q_reg ( .D(g17649), .SI(g4558), .SE(n10782), .CLK(n11165), 
        .Q(g17685), .QN(n10492) );
  SDFFX1 DFF_124_Q_reg ( .D(g25656), .SI(g17685), .SE(n10787), .CLK(n11170), 
        .Q(g3111) );
  SDFFX1 DFF_125_Q_reg ( .D(g30390), .SI(g3111), .SE(n10787), .CLK(n11170), 
        .Q(g29217) );
  SDFFX1 DFF_126_Q_reg ( .D(g25688), .SI(g29217), .SE(n10787), .CLK(n11170), 
        .Q(test_so9), .QN(n19407) );
  SDFFX1 DFF_127_Q_reg ( .D(g34727), .SI(test_si10), .SE(n10804), .CLK(n11187), 
        .Q(g939), .QN(n5415) );
  SDFFX1 DFF_128_Q_reg ( .D(g25594), .SI(g939), .SE(n10726), .CLK(n11109), .Q(
        g278), .QN(n5627) );
  SDFFX1 DFF_129_Q_reg ( .D(g26963), .SI(g278), .SE(n10726), .CLK(n11109), .Q(
        g4492), .QN(n10541) );
  SDFFX1 DFF_130_Q_reg ( .D(g34034), .SI(g4492), .SE(n10759), .CLK(n11142), 
        .Q(g4864), .QN(n5318) );
  SDFFX1 DFF_131_Q_reg ( .D(g33541), .SI(g4864), .SE(n10764), .CLK(n11147), 
        .Q(g1036), .QN(n10191) );
  SDFFX1 DFF_132_Q_reg ( .D(g28093), .SI(g1036), .SE(n10715), .CLK(n11098), 
        .Q(g29220), .QN(n10172) );
  SDFFX1 DFF_133_Q_reg ( .D(g24236), .SI(g29220), .SE(n10757), .CLK(n11140), 
        .Q(g1178) );
  SDFFX1 DFF_134_Q_reg ( .D(g30404), .SI(g1178), .SE(n10718), .CLK(n11101), 
        .Q(g3239), .QN(n10455) );
  SDFFX1 DFF_135_Q_reg ( .D(g28051), .SI(g3239), .SE(n10718), .CLK(n11101), 
        .Q(g718), .QN(n10312) );
  SDFFX1 DFF_136_Q_reg ( .D(g29303), .SI(g718), .SE(n10778), .CLK(n11161), .Q(
        g6195) );
  SDFFX1 DFF_137_Q_reg ( .D(g26917), .SI(g6195), .SE(n10737), .CLK(n11120), 
        .Q(g1135), .QN(n5328) );
  SDFFX1 DFF_139_Q_reg ( .D(g33624), .SI(g1135), .SE(n10793), .CLK(n11176), 
        .Q(g6395), .QN(n5396) );
  SDFFX1 DFF_141_Q_reg ( .D(g24337), .SI(g6395), .SE(n10793), .CLK(n11176), 
        .Q(test_so10), .QN(n10641) );
  SDFFX1 DFF_142_Q_reg ( .D(g34911), .SI(test_si11), .SE(n10799), .CLK(n11182), 
        .Q(g554), .QN(n10212) );
  SDFFX1 DFF_143_Q_reg ( .D(g33963), .SI(g554), .SE(n10736), .CLK(n11119), .Q(
        g496) );
  SDFFX1 DFF_144_Q_reg ( .D(g34627), .SI(g496), .SE(n10736), .CLK(n11119), .Q(
        g3853), .QN(n5641) );
  SDFFX1 DFF_145_Q_reg ( .D(g29282), .SI(g3853), .SE(n10736), .CLK(n11119), 
        .Q(g5134), .QN(n5807) );
  SDFFX1 DFF_146_Q_reg ( .D(g17320), .SI(g5134), .SE(n10736), .CLK(n11119), 
        .Q(g17404), .QN(n10235) );
  SDFFX1 DFF_147_Q_reg ( .D(g25676), .SI(g17404), .SE(n10777), .CLK(n11160), 
        .Q(g8344), .QN(n5721) );
  SDFFX1 DFF_148_Q_reg ( .D(g33013), .SI(g8344), .SE(n10803), .CLK(n11186), 
        .Q(g2485), .QN(n5509) );
  SDFFX1 DFF_149_Q_reg ( .D(g32981), .SI(g2485), .SE(n10731), .CLK(n11114), 
        .Q(g925), .QN(n5725) );
  SDFFX1 DFF_150_Q_reg ( .D(g34976), .SI(g925), .SE(n10701), .CLK(n11084), .Q(
        n9357) );
  SDFFX1 DFF_151_Q_reg ( .D(g30483), .SI(n9357), .SE(n10701), .CLK(n11084), 
        .Q(g5555), .QN(n10504) );
  SDFFX1 DFF_152_Q_reg ( .D(g14217), .SI(g5555), .SE(n10753), .CLK(n11136), 
        .Q(g14096), .QN(n10107) );
  SDFFX1 DFF_153_Q_reg ( .D(g32994), .SI(g14096), .SE(n10775), .CLK(n11158), 
        .Q(g1798), .QN(n5833) );
  SDFFX1 DFF_154_Q_reg ( .D(g28070), .SI(g1798), .SE(n10775), .CLK(n11158), 
        .Q(test_so11), .QN(n10644) );
  SDFFX1 DFF_155_Q_reg ( .D(g34806), .SI(test_si12), .SE(n10803), .CLK(n11186), 
        .Q(g2941), .QN(n10562) );
  SDFFX1 DFF_156_Q_reg ( .D(g30453), .SI(g2941), .SE(n10731), .CLK(n11114), 
        .Q(g3905) );
  SDFFX1 DFF_157_Q_reg ( .D(g33539), .SI(g3905), .SE(n10765), .CLK(n11148), 
        .Q(g763), .QN(n5332) );
  SDFFX1 DFF_158_Q_reg ( .D(g30526), .SI(g763), .SE(n10760), .CLK(n11143), .Q(
        g6255), .QN(n10430) );
  SDFFX1 DFF_159_Q_reg ( .D(n1545), .SI(g6255), .SE(n10746), .CLK(n11129), .Q(
        g4375), .QN(n10621) );
  SDFFX1 DFF_160_Q_reg ( .D(g34035), .SI(g4375), .SE(n10759), .CLK(n11142), 
        .Q(g4871), .QN(n5443) );
  SDFFX1 DFF_161_Q_reg ( .D(g34636), .SI(g4871), .SE(n10769), .CLK(n11152), 
        .Q(g4722) );
  SDFFX1 DFF_162_Q_reg ( .D(g32978), .SI(g4722), .SE(n10749), .CLK(n11132), 
        .Q(g590), .QN(n5472) );
  SDFFX1 DFF_163_Q_reg ( .D(g17722), .SI(g590), .SE(n10800), .CLK(n11183), .Q(
        g13099), .QN(n10511) );
  SDFFX1 DFF_164_Q_reg ( .D(g30348), .SI(g13099), .SE(n10724), .CLK(n11107), 
        .Q(g1632), .QN(n5836) );
  SDFFX1 DFF_165_Q_reg ( .D(g24336), .SI(g1632), .SE(n10718), .CLK(n11101), 
        .Q(g12238), .QN(n5438) );
  SDFFX1 DFF_166_Q_reg ( .D(g8215), .SI(g12238), .SE(n10754), .CLK(n11137), 
        .Q(g3100) );
  SDFFX1 DFF_167_Q_reg ( .D(g24250), .SI(g3100), .SE(n10754), .CLK(n11137), 
        .Q(test_so12) );
  SDFFX1 DFF_169_Q_reg ( .D(g29236), .SI(test_si13), .SE(n10754), .CLK(n11137), 
        .Q(g1437), .QN(n5696) );
  SDFFX1 DFF_170_Q_reg ( .D(g29298), .SI(g1437), .SE(n10704), .CLK(n11087), 
        .Q(g6154), .QN(n5747) );
  SDFFX1 DFF_171_Q_reg ( .D(g10527), .SI(g6154), .SE(n10747), .CLK(n11130), 
        .Q(g1579) );
  SDFFX1 DFF_172_Q_reg ( .D(g30499), .SI(g1579), .SE(n10792), .CLK(n11175), 
        .Q(g5567) );
  SDFFX1 DFF_173_Q_reg ( .D(g33976), .SI(g5567), .SE(n10763), .CLK(n11146), 
        .Q(g1752), .QN(n5797) );
  SDFFX1 DFF_174_Q_reg ( .D(g32996), .SI(g1752), .SE(n10765), .CLK(n11148), 
        .Q(g1917), .QN(n10531) );
  SDFFX1 DFF_175_Q_reg ( .D(g30335), .SI(g1917), .SE(n10765), .CLK(n11148), 
        .Q(g744), .QN(n5470) );
  SDFFX1 DFF_177_Q_reg ( .D(g34637), .SI(g744), .SE(n10769), .CLK(n11152), .Q(
        g4737), .QN(n5867) );
  SDFFX1 DFF_178_Q_reg ( .D(g25694), .SI(g4737), .SE(n10769), .CLK(n11152), 
        .Q(g8132), .QN(n19398) );
  SDFFX1 DFF_179_Q_reg ( .D(g30528), .SI(g8132), .SE(n10761), .CLK(n11144), 
        .Q(g6267), .QN(n10333) );
  SDFFX1 DFF_181_Q_reg ( .D(g16775), .SI(g6267), .SE(n10761), .CLK(n11144), 
        .Q(g16659), .QN(n10365) );
  SDFFX1 DFF_182_Q_reg ( .D(g24251), .SI(g16659), .SE(n10761), .CLK(n11144), 
        .Q(g1442), .QN(n10536) );
  SDFFX1 DFF_183_Q_reg ( .D(g30521), .SI(g1442), .SE(n10742), .CLK(n11125), 
        .Q(test_so13), .QN(n10684) );
  SDFFX1 DFF_184_Q_reg ( .D(g26960), .SI(test_si14), .SE(n10781), .CLK(n11164), 
        .Q(g4477), .QN(n5849) );
  SDFFX1 DFF_185_Q_reg ( .D(g24239), .SI(g4477), .SE(n10756), .CLK(n11139), 
        .Q(g10500) );
  SDFFX1 DFF_186_Q_reg ( .D(g34259), .SI(g10500), .SE(n10756), .CLK(n11139), 
        .Q(g4643), .QN(n5382) );
  SDFFX1 DFF_187_Q_reg ( .D(g30474), .SI(g4643), .SE(n10714), .CLK(n11097), 
        .Q(g5264), .QN(n10462) );
  SDFFX1 DFF_188_Q_reg ( .D(g12422), .SI(g5264), .SE(n10793), .CLK(n11176), 
        .Q(g14779), .QN(n5703) );
  SDFFX1 DFF_189_Q_reg ( .D(g33016), .SI(g14779), .SE(n10729), .CLK(n11112), 
        .Q(g2610), .QN(n10529) );
  SDFFX1 DFF_190_Q_reg ( .D(g34643), .SI(g2610), .SE(n10729), .CLK(n11112), 
        .Q(g5160), .QN(n5498) );
  SDFFX1 DFF_192_Q_reg ( .D(g30510), .SI(g5160), .SE(n10752), .CLK(n11135), 
        .Q(g5933), .QN(n10433) );
  SDFFX1 DFF_193_Q_reg ( .D(g29239), .SI(g5933), .SE(n10707), .CLK(n11090), 
        .Q(g1454), .QN(n5866) );
  SDFFX1 DFF_194_Q_reg ( .D(g26897), .SI(g1454), .SE(n10802), .CLK(n11185), 
        .Q(g753), .QN(n10183) );
  SDFFX1 DFF_195_Q_reg ( .D(g34729), .SI(g753), .SE(n10802), .CLK(n11185), .Q(
        g1296), .QN(n10093) );
  SDFFX1 DFF_196_Q_reg ( .D(g34625), .SI(g1296), .SE(n10802), .CLK(n11185), 
        .Q(g3151), .QN(n5495) );
  SDFFX1 DFF_197_Q_reg ( .D(g34800), .SI(g3151), .SE(n10703), .CLK(n11086), 
        .Q(test_so14) );
  SDFFX1 DFF_198_Q_reg ( .D(g24353), .SI(test_si15), .SE(n10729), .CLK(n11112), 
        .Q(g6727), .QN(n5531) );
  SDFFX1 DFF_199_Q_reg ( .D(g33029), .SI(g6727), .SE(n10762), .CLK(n11145), 
        .Q(g3530), .QN(n5569) );
  SDFFX1 DFF_201_Q_reg ( .D(g33615), .SI(g3530), .SE(n10776), .CLK(n11159), 
        .Q(g4104), .QN(n10403) );
  SDFFX1 DFF_202_Q_reg ( .D(g24253), .SI(g4104), .SE(n10762), .CLK(n11145), 
        .Q(g1532), .QN(n10398) );
  SDFFX1 DFF_203_Q_reg ( .D(g24281), .SI(g1532), .SE(n10776), .CLK(n11159), 
        .Q(g9251) );
  SDFFX1 DFF_204_Q_reg ( .D(g33997), .SI(g9251), .SE(n10755), .CLK(n11138), 
        .Q(n9352), .QN(n19408) );
  SDFFX1 DFF_206_Q_reg ( .D(g34971), .SI(n9352), .SE(n10704), .CLK(n11087), 
        .Q(n9351) );
  SDFFX1 DFF_207_Q_reg ( .D(g34263), .SI(n9351), .SE(n10704), .CLK(n11087), 
        .Q(g4754), .QN(n5877) );
  SDFFX1 DFF_208_Q_reg ( .D(g24237), .SI(g4754), .SE(n10777), .CLK(n11160), 
        .Q(g1189), .QN(n5642) );
  SDFFX1 DFF_209_Q_reg ( .D(g33584), .SI(g1189), .SE(n10791), .CLK(n11174), 
        .Q(g2287), .QN(n5353) );
  SDFFX1 DFF_210_Q_reg ( .D(g24280), .SI(g2287), .SE(n10763), .CLK(n11146), 
        .Q(g4273), .QN(n5764) );
  SDFFX1 DFF_211_Q_reg ( .D(g26920), .SI(g4273), .SE(n10723), .CLK(n11106), 
        .Q(g1389), .QN(n10620) );
  SDFFX1 DFF_212_Q_reg ( .D(g33548), .SI(g1389), .SE(n10723), .CLK(n11106), 
        .Q(test_so15), .QN(n10678) );
  SDFFX1 DFF_213_Q_reg ( .D(g29296), .SI(test_si16), .SE(n10713), .CLK(n11096), 
        .Q(g5835), .QN(n5663) );
  SDFFX1 DFF_214_Q_reg ( .D(g30338), .SI(g5835), .SE(n10757), .CLK(n11140), 
        .Q(g1171), .QN(n5363) );
  SDFFX1 DFF_215_Q_reg ( .D(g21895), .SI(g1171), .SE(n10763), .CLK(n11146), 
        .Q(g4269), .QN(n5763) );
  SDFFX1 DFF_216_Q_reg ( .D(n403), .SI(g4269), .SE(n10708), .CLK(n11091), .Q(
        g2399), .QN(n5762) );
  SDFFX1 DFF_218_Q_reg ( .D(g34041), .SI(g2399), .SE(n10759), .CLK(n11142), 
        .Q(g4983), .QN(n5367) );
  SDFFX1 DFF_219_Q_reg ( .D(g30495), .SI(g4983), .SE(n10789), .CLK(n11172), 
        .Q(g5611), .QN(n10472) );
  SDFFX1 DFF_220_Q_reg ( .D(g16744), .SI(g5611), .SE(n10789), .CLK(n11172), 
        .Q(g16627), .QN(n10369) );
  SDFFX1 DFF_221_Q_reg ( .D(g29279), .SI(g16627), .SE(n10719), .CLK(n11102), 
        .Q(g4572), .QN(n10182) );
  SDFFX1 DFF_222_Q_reg ( .D(g25655), .SI(g4572), .SE(n10703), .CLK(n11086), 
        .Q(g3143), .QN(n5882) );
  SDFFX1 DFF_223_Q_reg ( .D(g34795), .SI(g3143), .SE(n10703), .CLK(n11086), 
        .Q(g2898), .QN(n10566) );
  SDFFX1 DFF_224_Q_reg ( .D(g24269), .SI(g2898), .SE(n10722), .CLK(n11105), 
        .Q(g3343), .QN(n10388) );
  SDFFX1 DFF_225_Q_reg ( .D(g30403), .SI(g3343), .SE(n10722), .CLK(n11105), 
        .Q(g3235), .QN(n10373) );
  SDFFX1 DFF_226_Q_reg ( .D(g33042), .SI(g3235), .SE(n10784), .CLK(n11167), 
        .Q(test_so16) );
  SDFFX1 DFF_227_Q_reg ( .D(g30419), .SI(test_si17), .SE(n10762), .CLK(n11145), 
        .Q(g3566), .QN(n10297) );
  SDFFX1 DFF_228_Q_reg ( .D(g34023), .SI(g3566), .SE(n10798), .CLK(n11181), 
        .Q(n9348), .QN(DFF_228_n1) );
  SDFFX1 DFF_229_Q_reg ( .D(g28090), .SI(n9348), .SE(n10702), .CLK(n11085), 
        .Q(g4961), .QN(n5770) );
  SDFFX1 DFF_231_Q_reg ( .D(g34642), .SI(g4961), .SE(n10734), .CLK(n11117), 
        .Q(g4927), .QN(n5879) );
  SDFFX1 DFF_232_Q_reg ( .D(g30370), .SI(g4927), .SE(n10734), .CLK(n11117), 
        .Q(g2259), .QN(n5419) );
  SDFFX1 DFF_233_Q_reg ( .D(g34448), .SI(g2259), .SE(n10728), .CLK(n11111), 
        .Q(g2819), .QN(n5609) );
  SDFFX1 DFF_234_Q_reg ( .D(g26946), .SI(g2819), .SE(n10772), .CLK(n11155), 
        .Q(g7257) );
  SDFFX1 DFF_235_Q_reg ( .D(g9617), .SI(g7257), .SE(n10786), .CLK(n11169), .Q(
        g5802) );
  SDFFX1 DFF_236_Q_reg ( .D(g34610), .SI(g5802), .SE(n10743), .CLK(n11126), 
        .Q(g2852) );
  SDFFX1 DFF_237_Q_reg ( .D(g24209), .SI(g2852), .SE(n10785), .CLK(n11168), 
        .Q(g417), .QN(n5358) );
  SDFFX1 DFF_238_Q_reg ( .D(g28047), .SI(g417), .SE(n10785), .CLK(n11168), .Q(
        g681), .QN(n10233) );
  SDFFX1 DFF_239_Q_reg ( .D(g24206), .SI(g681), .SE(n10770), .CLK(n11153), .Q(
        g437), .QN(n10246) );
  SDFFX1 DFF_240_Q_reg ( .D(g26891), .SI(g437), .SE(n10770), .CLK(n11153), .Q(
        test_so17), .QN(n10674) );
  SDFFX1 DFF_241_Q_reg ( .D(g30504), .SI(test_si18), .SE(n10741), .CLK(n11124), 
        .Q(g5901), .QN(n10500) );
  SDFFX1 DFF_242_Q_reg ( .D(g34798), .SI(g5901), .SE(n10703), .CLK(n11086), 
        .Q(g2886), .QN(n10564) );
  SDFFX1 DFF_243_Q_reg ( .D(g25669), .SI(g2886), .SE(n10720), .CLK(n11103), 
        .Q(g3494), .QN(n5889) );
  SDFFX1 DFF_244_Q_reg ( .D(g30480), .SI(g3494), .SE(n10720), .CLK(n11103), 
        .Q(g5511), .QN(n5575) );
  SDFFX1 DFF_245_Q_reg ( .D(g33027), .SI(g5511), .SE(n10777), .CLK(n11160), 
        .Q(g3518), .QN(n5645) );
  SDFFX1 DFF_246_Q_reg ( .D(g33972), .SI(g3518), .SE(n10737), .CLK(n11120), 
        .Q(g1604), .QN(n10135) );
  SDFFX1 DFF_248_Q_reg ( .D(g25697), .SI(g1604), .SE(n10699), .CLK(n11082), 
        .Q(g5092) );
  SDFFX1 DFF_249_Q_reg ( .D(g28099), .SI(g5092), .SE(n10742), .CLK(n11125), 
        .Q(g4831), .QN(n10173) );
  SDFFX1 DFF_250_Q_reg ( .D(g26947), .SI(g4831), .SE(n10742), .CLK(n11125), 
        .Q(g4382), .QN(n5714) );
  SDFFX1 DFF_251_Q_reg ( .D(g24350), .SI(g4382), .SE(n10794), .CLK(n11177), 
        .Q(g6386), .QN(n10390) );
  SDFFX1 DFF_252_Q_reg ( .D(g24210), .SI(g6386), .SE(n10735), .CLK(n11118), 
        .Q(g479), .QN(n10223) );
  SDFFX1 DFF_253_Q_reg ( .D(g30455), .SI(g479), .SE(n10800), .CLK(n11183), .Q(
        g3965), .QN(n10309) );
  SDFFX1 DFF_254_Q_reg ( .D(g28084), .SI(g3965), .SE(n10713), .CLK(n11096), 
        .Q(test_so18) );
  SDFFX1 DFF_255_Q_reg ( .D(g33993), .SI(test_si19), .SE(n10744), .CLK(n11127), 
        .Q(g2008), .QN(n10217) );
  SDFFX1 DFF_256_Q_reg ( .D(g11678), .SI(g2008), .SE(n10788), .CLK(n11171), 
        .Q(g736) );
  SDFFX1 DFF_257_Q_reg ( .D(g30444), .SI(g736), .SE(n10775), .CLK(n11158), .Q(
        g3933), .QN(n10435) );
  SDFFX1 DFF_258_Q_reg ( .D(g33537), .SI(g3933), .SE(n10775), .CLK(n11158), 
        .Q(g222), .QN(n10573) );
  SDFFX1 DFF_259_Q_reg ( .D(g25650), .SI(g222), .SE(n10801), .CLK(n11184), .Q(
        g3050) );
  SDFFX1 DFF_261_Q_reg ( .D(g25625), .SI(g3050), .SE(n10751), .CLK(n11134), 
        .Q(g1052), .QN(n10579) );
  SDFFX1 DFF_263_Q_reg ( .D(g17711), .SI(g1052), .SE(n10751), .CLK(n11134), 
        .Q(g17580), .QN(n10363) );
  SDFFX1 DFF_264_Q_reg ( .D(g30366), .SI(g17580), .SE(n10701), .CLK(n11084), 
        .Q(g2122), .QN(n5784) );
  SDFFX1 DFF_265_Q_reg ( .D(g33593), .SI(g2122), .SE(n10752), .CLK(n11135), 
        .Q(g2465), .QN(n5523) );
  SDFFX1 DFF_267_Q_reg ( .D(g30502), .SI(g2465), .SE(n10752), .CLK(n11135), 
        .Q(g5889), .QN(n10445) );
  SDFFX1 DFF_268_Q_reg ( .D(g33036), .SI(g5889), .SE(n10784), .CLK(n11167), 
        .Q(g4495) );
  SDFFX1 DFF_269_Q_reg ( .D(g25595), .SI(g4495), .SE(n10784), .CLK(n11167), 
        .Q(g8719), .QN(n10280) );
  SDFFX1 DFF_270_Q_reg ( .D(g34462), .SI(g8719), .SE(n10767), .CLK(n11150), 
        .Q(test_so19), .QN(n10645) );
  SDFFX1 DFF_271_Q_reg ( .D(g33024), .SI(test_si20), .SE(n10754), .CLK(n11137), 
        .Q(g3179), .QN(n5390) );
  SDFFX1 DFF_272_Q_reg ( .D(g33552), .SI(g3179), .SE(n10771), .CLK(n11154), 
        .Q(g1728), .QN(n5352) );
  SDFFX1 DFF_273_Q_reg ( .D(g34014), .SI(g1728), .SE(n10728), .CLK(n11111), 
        .Q(g2433), .QN(n10136) );
  SDFFX1 DFF_274_Q_reg ( .D(g29273), .SI(g2433), .SE(n10700), .CLK(n11083), 
        .Q(g3835), .QN(n5662) );
  SDFFX1 DFF_275_Q_reg ( .D(n55), .SI(g3835), .SE(n10778), .CLK(n11161), .Q(
        g6187), .QN(n5453) );
  SDFFX1 DFF_276_Q_reg ( .D(g34638), .SI(g6187), .SE(n10778), .CLK(n11161), 
        .Q(g4917), .QN(n5408) );
  SDFFX1 DFF_277_Q_reg ( .D(g30341), .SI(g4917), .SE(n10745), .CLK(n11128), 
        .Q(g1070), .QN(n10089) );
  SDFFX1 DFF_278_Q_reg ( .D(g26899), .SI(g1070), .SE(n10745), .CLK(n11128), 
        .Q(g822), .QN(n5422) );
  SDFFX1 DFF_279_Q_reg ( .D(g14673), .SI(g822), .SE(n10779), .CLK(n11162), .Q(
        g17715) );
  SDFFX1 DFF_280_Q_reg ( .D(g30336), .SI(g17715), .SE(n10730), .CLK(n11113), 
        .Q(g914), .QN(n5560) );
  SDFFX1 DFF_281_Q_reg ( .D(g17639), .SI(g914), .SE(n10786), .CLK(n11169), .Q(
        g5339) );
  SDFFX1 DFF_282_Q_reg ( .D(g26940), .SI(g5339), .SE(n10786), .CLK(n11169), 
        .Q(g4164), .QN(n10552) );
  SDFFX1 DFF_283_Q_reg ( .D(g25622), .SI(g4164), .SE(n10704), .CLK(n11087), 
        .Q(test_so20) );
  SDFFX1 DFF_284_Q_reg ( .D(g34447), .SI(test_si21), .SE(n10780), .CLK(n11163), 
        .Q(g2807), .QN(n5379) );
  SDFFX1 DFF_286_Q_reg ( .D(g33613), .SI(g2807), .SE(n10702), .CLK(n11085), 
        .Q(g4054), .QN(n5395) );
  SDFFX1 DFF_287_Q_reg ( .D(g25749), .SI(g4054), .SE(n10705), .CLK(n11088), 
        .Q(g6191), .QN(n5888) );
  SDFFX1 DFF_288_Q_reg ( .D(g25704), .SI(g6191), .SE(n10705), .CLK(n11088), 
        .Q(g5077), .QN(n5455) );
  SDFFX1 DFF_289_Q_reg ( .D(g33053), .SI(g5077), .SE(n10705), .CLK(n11088), 
        .Q(g5523), .QN(n5647) );
  SDFFX1 DFF_290_Q_reg ( .D(g16722), .SI(g5523), .SE(n10747), .CLK(n11130), 
        .Q(g3680) );
  SDFFX1 DFF_291_Q_reg ( .D(g30555), .SI(g3680), .SE(n10735), .CLK(n11118), 
        .Q(g6637), .QN(n10349) );
  SDFFX1 DFF_292_Q_reg ( .D(g25601), .SI(g6637), .SE(n10735), .CLK(n11118), 
        .Q(g174), .QN(n5402) );
  SDFFX1 DFF_293_Q_reg ( .D(g33971), .SI(g174), .SE(n10737), .CLK(n11120), .Q(
        g1682), .QN(n10201) );
  SDFFX1 DFF_294_Q_reg ( .D(g26892), .SI(g1682), .SE(n10770), .CLK(n11153), 
        .Q(g355) );
  SDFFX1 DFF_295_Q_reg ( .D(g17400), .SI(g355), .SE(n10770), .CLK(n11153), .Q(
        g1087), .QN(n10548) );
  SDFFX1 DFF_296_Q_reg ( .D(g26915), .SI(g1087), .SE(n10740), .CLK(n11123), 
        .Q(g1105), .QN(n5478) );
  SDFFX1 DFF_297_Q_reg ( .D(g33008), .SI(g1105), .SE(n10798), .CLK(n11181), 
        .Q(test_so21), .QN(n10640) );
  SDFFX1 DFF_298_Q_reg ( .D(g30538), .SI(test_si22), .SE(n10760), .CLK(n11143), 
        .Q(g6307), .QN(n10354) );
  SDFFX1 DFF_299_Q_reg ( .D(g8344), .SI(g6307), .SE(n10777), .CLK(n11160), .Q(
        g3802) );
  SDFFX1 DFF_300_Q_reg ( .D(g25750), .SI(g3802), .SE(n10778), .CLK(n11161), 
        .Q(g6159) );
  SDFFX1 DFF_301_Q_reg ( .D(g30369), .SI(g6159), .SE(n10803), .CLK(n11186), 
        .Q(g2255), .QN(n5414) );
  SDFFX1 DFF_302_Q_reg ( .D(g34446), .SI(g2255), .SE(n10717), .CLK(n11100), 
        .Q(g2815), .QN(n5404) );
  SDFFX1 DFF_303_Q_reg ( .D(g29230), .SI(g2815), .SE(n10730), .CLK(n11113), 
        .Q(g911), .QN(n5559) );
  SDFFX1 DFF_304_Q_reg ( .D(n10623), .SI(g911), .SE(n10727), .CLK(n11110), .Q(
        g43) );
  SDFFX1 DFF_305_Q_reg ( .D(g13966), .SI(g43), .SE(n10727), .CLK(n11110), .Q(
        g16775), .QN(n10379) );
  SDFFX1 DFF_306_Q_reg ( .D(g33975), .SI(g16775), .SE(n10763), .CLK(n11146), 
        .Q(g1748) );
  SDFFX1 DFF_307_Q_reg ( .D(g30497), .SI(g1748), .SE(n10705), .CLK(n11088), 
        .Q(g5551) );
  SDFFX1 DFF_309_Q_reg ( .D(g30418), .SI(g5551), .SE(n10804), .CLK(n11187), 
        .Q(g3558), .QN(n10427) );
  SDFFX1 DFF_310_Q_reg ( .D(g25721), .SI(g3558), .SE(n10699), .CLK(n11082), 
        .Q(g5499) );
  SDFFX1 DFF_311_Q_reg ( .D(g34622), .SI(g5499), .SE(n10803), .CLK(n11186), 
        .Q(test_so22), .QN(n10660) );
  SDFFX1 DFF_312_Q_reg ( .D(g30438), .SI(test_si23), .SE(n10731), .CLK(n11114), 
        .Q(g3901), .QN(n10508) );
  SDFFX1 DFF_313_Q_reg ( .D(g34266), .SI(g3901), .SE(n10730), .CLK(n11113), 
        .Q(g4888), .QN(n5863) );
  SDFFX1 DFF_314_Q_reg ( .D(g30540), .SI(g4888), .SE(n10761), .CLK(n11144), 
        .Q(g6251), .QN(n10493) );
  SDFFX1 DFF_315_Q_reg ( .D(g17760), .SI(g6251), .SE(n10793), .CLK(n11176), 
        .Q(g17649), .QN(n10370) );
  SDFFX1 DFF_316_Q_reg ( .D(g32986), .SI(g17649), .SE(n10724), .CLK(n11107), 
        .Q(g1373), .QN(n10259) );
  SDFFX1 DFF_317_Q_reg ( .D(g25648), .SI(g1373), .SE(n10754), .CLK(n11137), 
        .Q(g8215), .QN(n5723) );
  SDFFX1 DFF_318_Q_reg ( .D(g33960), .SI(g8215), .SE(n10711), .CLK(n11094), 
        .Q(g157), .QN(n5678) );
  SDFFX1 DFF_319_Q_reg ( .D(g34442), .SI(g157), .SE(n10792), .CLK(n11175), .Q(
        g2783), .QN(n5403) );
  SDFFX1 DFF_320_Q_reg ( .D(g8839), .SI(g2783), .SE(n10756), .CLK(n11139), .Q(
        g4281), .QN(n10576) );
  SDFFX1 DFF_321_Q_reg ( .D(g30421), .SI(g4281), .SE(n10732), .CLK(n11115), 
        .Q(g3574), .QN(n10426) );
  SDFFX1 DFF_322_Q_reg ( .D(g33573), .SI(g3574), .SE(n10804), .CLK(n11187), 
        .Q(g2112), .QN(n5848) );
  SDFFX1 DFF_323_Q_reg ( .D(g34730), .SI(g2112), .SE(n10710), .CLK(n11093), 
        .Q(g1283), .QN(n5635) );
  SDFFX1 DFF_324_Q_reg ( .D(g24205), .SI(g1283), .SE(n10710), .CLK(n11093), 
        .Q(test_so23), .QN(n10693) );
  SDFFX1 DFF_325_Q_reg ( .D(g10122_Tj), .SI(test_si24), .SE(n10733), .CLK(
        n11116), .Q(g4297) );
  SDFFX1 DFF_326_Q_reg ( .D(g12350), .SI(g4297), .SE(n10733), .CLK(n11116), 
        .Q(g14738), .QN(n5698) );
  SDFFX1 DFF_327_Q_reg ( .D(g19357), .SI(g14738), .SE(n10733), .CLK(n11116), 
        .Q(g13272), .QN(n10244) );
  SDFFX1 DFF_328_Q_reg ( .D(g32979), .SI(g13272), .SE(n10765), .CLK(n11148), 
        .Q(g758), .QN(n5331) );
  SDFFX1 DFF_331_Q_reg ( .D(g34025), .SI(g758), .SE(n10765), .CLK(n11148), .Q(
        g4639), .QN(n5727) );
  SDFFX1 DFF_332_Q_reg ( .D(g25763), .SI(g4639), .SE(n10804), .CLK(n11187), 
        .Q(g6537) );
  SDFFX1 DFF_333_Q_reg ( .D(g30481), .SI(g6537), .SE(n10705), .CLK(n11088), 
        .Q(g5543), .QN(n10447) );
  SDFFX1 DFF_334_Q_reg ( .D(g7946), .SI(g5543), .SE(n10762), .CLK(n11145), .Q(
        g8475), .QN(n10157) );
  SDFFX1 DFF_336_Q_reg ( .D(g30517), .SI(g8475), .SE(n10742), .CLK(n11125), 
        .Q(g5961), .QN(n10339) );
  SDFFX1 DFF_337_Q_reg ( .D(g30539), .SI(g5961), .SE(n10799), .CLK(n11182), 
        .Q(g6243) );
  SDFFX1 DFF_338_Q_reg ( .D(g34880), .SI(g6243), .SE(n10750), .CLK(n11133), 
        .Q(n9340), .QN(n19409) );
  SDFFX1 DFF_339_Q_reg ( .D(g24242), .SI(n9340), .SE(n10751), .CLK(n11134), 
        .Q(g12919), .QN(n5654) );
  SDFFX1 DFF_340_Q_reg ( .D(g30436), .SI(g12919), .SE(n10775), .CLK(n11158), 
        .Q(test_so24), .QN(n10686) );
  SDFFX1 DFF_341_Q_reg ( .D(g29265), .SI(test_si25), .SE(n10720), .CLK(n11103), 
        .Q(g3476), .QN(n5786) );
  SDFFX1 DFF_342_Q_reg ( .D(g32990), .SI(g3476), .SE(n10724), .CLK(n11107), 
        .Q(g1664), .QN(n5407) );
  SDFFX1 DFF_343_Q_reg ( .D(g24245), .SI(g1664), .SE(n10751), .CLK(n11134), 
        .Q(g1246), .QN(n5756) );
  SDFFX1 DFF_345_Q_reg ( .D(g30553), .SI(g1246), .SE(n10734), .CLK(n11117), 
        .Q(g6629), .QN(n10382) );
  SDFFX1 DFF_346_Q_reg ( .D(g26907), .SI(g6629), .SE(n10770), .CLK(n11153), 
        .Q(g246), .QN(n6008) );
  SDFFX1 DFF_347_Q_reg ( .D(g24278), .SI(g246), .SE(n10727), .CLK(n11110), .Q(
        g4049), .QN(n10396) );
  SDFFX1 DFF_348_Q_reg ( .D(g26955), .SI(g4049), .SE(n10742), .CLK(n11125), 
        .Q(g7260) );
  SDFFX1 DFF_349_Q_reg ( .D(g24282), .SI(g7260), .SE(n10742), .CLK(n11125), 
        .Q(g2932) );
  SDFFX1 DFF_350_Q_reg ( .D(n1688), .SI(g2932), .SE(n10742), .CLK(n11125), .Q(
        g4575) );
  SDFFX1 DFF_351_Q_reg ( .D(g31894), .SI(g4575), .SE(n10727), .CLK(n11110), 
        .Q(g4098), .QN(n5350) );
  SDFFX1 DFF_352_Q_reg ( .D(g33037), .SI(g4098), .SE(n10784), .CLK(n11167), 
        .Q(g4498) );
  SDFFX1 DFF_353_Q_reg ( .D(g26894), .SI(g4498), .SE(n10773), .CLK(n11156), 
        .Q(g528), .QN(n5327) );
  SDFFX1 DFF_355_Q_reg ( .D(g34977), .SI(g528), .SE(n10804), .CLK(n11187), .Q(
        test_so25), .QN(n5477) );
  SDFFX1 DFF_356_Q_reg ( .D(n176), .SI(test_si26), .SE(n10789), .CLK(n11172), 
        .Q(g3139), .QN(n5447) );
  SDFFX1 DFF_357_Q_reg ( .D(g33962), .SI(g3139), .SE(n10735), .CLK(n11118), 
        .Q(g29215) );
  SDFFX1 DFF_358_Q_reg ( .D(g34451), .SI(g29215), .SE(n10767), .CLK(n11150), 
        .Q(g4584), .QN(n5539) );
  SDFFX1 DFF_359_Q_reg ( .D(g34250), .SI(g4584), .SE(n10711), .CLK(n11094), 
        .Q(g142), .QN(n5724) );
  SDFFX1 DFF_360_Q_reg ( .D(g14597), .SI(g142), .SE(n10786), .CLK(n11169), .Q(
        g17639) );
  SDFFX1 DFF_361_Q_reg ( .D(g29295), .SI(g17639), .SE(n10713), .CLK(n11096), 
        .Q(g5831) );
  SDFFX1 DFF_362_Q_reg ( .D(g26905), .SI(g5831), .SE(n10753), .CLK(n11136), 
        .Q(g239), .QN(n10400) );
  SDFFX1 DFF_363_Q_reg ( .D(g25629), .SI(g239), .SE(n10756), .CLK(n11139), .Q(
        g1216), .QN(n5442) );
  SDFFX1 DFF_364_Q_reg ( .D(g34792), .SI(g1216), .SE(n10702), .CLK(n11085), 
        .Q(g2848), .QN(n10613) );
  SDFFX1 DFF_366_Q_reg ( .D(g25703), .SI(g2848), .SE(n10779), .CLK(n11162), 
        .Q(g5022), .QN(n10278) );
  SDFFX1 DFF_367_Q_reg ( .D(g14518), .SI(g5022), .SE(n10780), .CLK(n11163), 
        .Q(g16955) );
  SDFFX1 DFF_368_Q_reg ( .D(g32983), .SI(g16955), .SE(n10794), .CLK(n11177), 
        .Q(g1030), .QN(n10261) );
  SDFFX1 DFF_369_Q_reg ( .D(g16924), .SI(g1030), .SE(n10794), .CLK(n11177), 
        .Q(test_so26) );
  SDFFX1 DFF_370_Q_reg ( .D(g30402), .SI(test_si27), .SE(n10790), .CLK(n11173), 
        .Q(g3231), .QN(n10431) );
  SDFFX1 DFF_371_Q_reg ( .D(g25757), .SI(g3231), .SE(n10790), .CLK(n11173), 
        .Q(g9817) );
  SDFFX1 DFF_372_Q_reg ( .D(g17423), .SI(g9817), .SE(n10790), .CLK(n11173), 
        .Q(g1430), .QN(n10546) );
  SDFFX1 DFF_373_Q_reg ( .D(g7245), .SI(g1430), .SE(n10794), .CLK(n11177), .Q(
        n9336), .QN(n19410) );
  SDFFX1 DFF_374_Q_reg ( .D(g33999), .SI(n9336), .SE(n10736), .CLK(n11119), 
        .Q(g2241), .QN(n10200) );
  SDFFX1 DFF_375_Q_reg ( .D(g24262), .SI(g2241), .SE(n10790), .CLK(n11173), 
        .Q(g1564), .QN(n10545) );
  SDFFX1 DFF_376_Q_reg ( .D(g25729), .SI(g1564), .SE(n10799), .CLK(n11182), 
        .Q(g9680) );
  SDFFX1 DFF_377_Q_reg ( .D(test_so92), .SI(g9680), .SE(n10799), .CLK(n11182), 
        .Q(g6148) );
  SDFFX1 DFF_378_Q_reg ( .D(g30558), .SI(g6148), .SE(n10735), .CLK(n11118), 
        .Q(g6649), .QN(n10481) );
  SDFFX1 DFF_379_Q_reg ( .D(g34781), .SI(g6649), .SE(n10729), .CLK(n11112), 
        .Q(g110), .QN(n10087) );
  SDFFX1 DFF_380_Q_reg ( .D(g14125), .SI(g110), .SE(n10753), .CLK(n11136), .Q(
        g14147), .QN(n10110) );
  SDFFX1 DFF_382_Q_reg ( .D(g26901), .SI(g14147), .SE(n10753), .CLK(n11136), 
        .Q(g225), .QN(n5597) );
  SDFFX1 DFF_383_Q_reg ( .D(g26961), .SI(g225), .SE(n10753), .CLK(n11136), .Q(
        test_so27), .QN(n10692) );
  SDFFX1 DFF_384_Q_reg ( .D(g33039), .SI(test_si28), .SE(n10784), .CLK(n11167), 
        .Q(g4504) );
  SDFFX1 DFF_385_Q_reg ( .D(g33059), .SI(g4504), .SE(n10785), .CLK(n11168), 
        .Q(g5873), .QN(n5388) );
  SDFFX1 DFF_386_Q_reg ( .D(g31899), .SI(g5873), .SE(n10794), .CLK(n11177), 
        .Q(g5037), .QN(n5611) );
  SDFFX1 DFF_387_Q_reg ( .D(g33007), .SI(g5037), .SE(n10797), .CLK(n11180), 
        .Q(g2319), .QN(n5375) );
  SDFFX1 DFF_388_Q_reg ( .D(n623), .SI(g2319), .SE(n10798), .CLK(n11181), .Q(
        g5495), .QN(n5446) );
  SDFFX1 DFF_389_Q_reg ( .D(g21891), .SI(g5495), .SE(n10740), .CLK(n11123), 
        .Q(g11770) );
  SDFFX1 DFF_390_Q_reg ( .D(g30462), .SI(g11770), .SE(n10740), .CLK(n11123), 
        .Q(g5208), .QN(n10406) );
  SDFFX1 DFF_392_Q_reg ( .D(g30487), .SI(g5208), .SE(n10783), .CLK(n11166), 
        .Q(g5579), .QN(n10417) );
  SDFFX1 DFF_393_Q_reg ( .D(g33058), .SI(g5579), .SE(n10783), .CLK(n11166), 
        .Q(g5869), .QN(n5649) );
  SDFFX1 DFF_395_Q_reg ( .D(g24261), .SI(g5869), .SE(n10783), .CLK(n11166), 
        .Q(g1589), .QN(n5755) );
  SDFFX1 DFF_396_Q_reg ( .D(g25730), .SI(g1589), .SE(n10799), .CLK(n11182), 
        .Q(g5752) );
  SDFFX1 DFF_397_Q_reg ( .D(g30531), .SI(g5752), .SE(n10799), .CLK(n11182), 
        .Q(g6279), .QN(n10438) );
  SDFFX1 DFF_398_Q_reg ( .D(g30506), .SI(g6279), .SE(n10752), .CLK(n11135), 
        .Q(test_so28), .QN(n10685) );
  SDFFX1 DFF_399_Q_reg ( .D(g34804), .SI(test_si29), .SE(n10777), .CLK(n11160), 
        .Q(g2975), .QN(n5750) );
  SDFFX1 DFF_400_Q_reg ( .D(g25747), .SI(g2975), .SE(n10704), .CLK(n11087), 
        .Q(g6167), .QN(n5430) );
  SDFFX1 DFF_401_Q_reg ( .D(g11418), .SI(g6167), .SE(n10727), .CLK(n11110), 
        .Q(g13966), .QN(n5701) );
  SDFFX1 DFF_402_Q_reg ( .D(g33601), .SI(g13966), .SE(n10728), .CLK(n11111), 
        .Q(g2599), .QN(n5524) );
  SDFFX1 DFF_403_Q_reg ( .D(g26922), .SI(g2599), .SE(n10707), .CLK(n11090), 
        .Q(g1448), .QN(n5343) );
  SDFFX1 DFF_404_Q_reg ( .D(g14096), .SI(g1448), .SE(n10753), .CLK(n11136), 
        .Q(g14125), .QN(n10109) );
  SDFFX1 DFF_406_Q_reg ( .D(g29250), .SI(g14125), .SE(n10729), .CLK(n11112), 
        .Q(g2370), .QN(n10319) );
  SDFFX1 DFF_407_Q_reg ( .D(g30459), .SI(g2370), .SE(n10779), .CLK(n11162), 
        .Q(g5164), .QN(n5570) );
  SDFFX1 DFF_408_Q_reg ( .D(g8475), .SI(g5164), .SE(n10779), .CLK(n11162), .Q(
        g1333), .QN(n5616) );
  SDFFX1 DFF_409_Q_reg ( .D(g33534), .SI(g1333), .SE(n10711), .CLK(n11094), 
        .Q(g153), .QN(n5677) );
  SDFFX1 DFF_410_Q_reg ( .D(g30543), .SI(g153), .SE(n10776), .CLK(n11159), .Q(
        g6549), .QN(n5571) );
  SDFFX1 DFF_411_Q_reg ( .D(g29275), .SI(g6549), .SE(n10776), .CLK(n11159), 
        .Q(g4087), .QN(n5480) );
  SDFFX1 DFF_412_Q_reg ( .D(g34030), .SI(g4087), .SE(n10799), .CLK(n11182), 
        .Q(test_so29), .QN(n10661) );
  SDFFX1 DFF_413_Q_reg ( .D(g34980), .SI(test_si30), .SE(n10771), .CLK(n11154), 
        .Q(g2984), .QN(n5842) );
  SDFFX1 DFF_414_Q_reg ( .D(g30451), .SI(g2984), .SE(n10776), .CLK(n11159), 
        .Q(g3961) );
  SDFFX1 DFF_416_Q_reg ( .D(g25627), .SI(g3961), .SE(n10776), .CLK(n11159), 
        .Q(g962), .QN(n5630) );
  SDFFX1 DFF_417_Q_reg ( .D(g34657), .SI(g962), .SE(n10704), .CLK(n11087), .Q(
        g101), .QN(n19411) );
  SDFFX1 DFF_418_Q_reg ( .D(g8870), .SI(g101), .SE(n10716), .CLK(n11099), .Q(
        g8918) );
  SDFFX1 DFF_419_Q_reg ( .D(g30552), .SI(g8918), .SE(n10795), .CLK(n11178), 
        .Q(g6625), .QN(n10436) );
  SDFFX1 DFF_420_Q_reg ( .D(g34979), .SI(g6625), .SE(n10703), .CLK(n11086), 
        .Q(n9332) );
  SDFFX1 DFF_421_Q_reg ( .D(g30337), .SI(n9332), .SE(n10704), .CLK(n11087), 
        .Q(g1018), .QN(n10260) );
  SDFFX1 DFF_422_Q_reg ( .D(g24254), .SI(g1018), .SE(n10736), .CLK(n11119), 
        .Q(g17320), .QN(n10236) );
  SDFFX1 DFF_423_Q_reg ( .D(g24277), .SI(g17320), .SE(n10727), .CLK(n11110), 
        .Q(g4045), .QN(n10397) );
  SDFFX1 DFF_424_Q_reg ( .D(g29237), .SI(g4045), .SE(n10727), .CLK(n11110), 
        .Q(g1467), .QN(n5693) );
  SDFFX1 DFF_425_Q_reg ( .D(g30378), .SI(g1467), .SE(n10738), .CLK(n11121), 
        .Q(g2461), .QN(n5840) );
  SDFFX1 DFF_428_Q_reg ( .D(g33019), .SI(g2461), .SE(n10788), .CLK(n11171), 
        .Q(test_so30), .QN(n5300) );
  SDFFX1 DFF_429_Q_reg ( .D(g33623), .SI(test_si31), .SE(n10712), .CLK(n11095), 
        .Q(g5990), .QN(n5589) );
  SDFFX1 DFF_431_Q_reg ( .D(g29235), .SI(g5990), .SE(n10709), .CLK(n11092), 
        .Q(g1256), .QN(n5558) );
  SDFFX1 DFF_432_Q_reg ( .D(g31902), .SI(g1256), .SE(n10768), .CLK(n11151), 
        .Q(g5029), .QN(n5601) );
  SDFFX1 DFF_433_Q_reg ( .D(n479), .SI(g5029), .SE(n10727), .CLK(n11110), .Q(
        g6519), .QN(n5806) );
  SDFFX1 DFF_434_Q_reg ( .D(g25689), .SI(g6519), .SE(n10727), .CLK(n11110), 
        .Q(g4169), .QN(n5729) );
  SDFFX1 DFF_435_Q_reg ( .D(g33978), .SI(g4169), .SE(n10741), .CLK(n11124), 
        .Q(g1816), .QN(n10128) );
  SDFFX1 DFF_436_Q_reg ( .D(g26970), .SI(g1816), .SE(n10782), .CLK(n11165), 
        .Q(g4369), .QN(n10401) );
  SDFFX1 DFF_439_Q_reg ( .D(n524), .SI(g4369), .SE(n10782), .CLK(n11165), .Q(
        g4578) );
  SDFFX1 DFF_440_Q_reg ( .D(g34253), .SI(g4578), .SE(n10781), .CLK(n11164), 
        .Q(g4459), .QN(n5765) );
  SDFFX1 DFF_441_Q_reg ( .D(g29272), .SI(g4459), .SE(n10700), .CLK(n11083), 
        .Q(g3831), .QN(n5872) );
  SDFFX1 DFF_442_Q_reg ( .D(g33595), .SI(g3831), .SE(n10728), .CLK(n11111), 
        .Q(g2514), .QN(n10163) );
  SDFFX1 DFF_443_Q_reg ( .D(g33610), .SI(g2514), .SE(n10702), .CLK(n11085), 
        .Q(g3288) );
  SDFFX1 DFF_444_Q_reg ( .D(g33589), .SI(g3288), .SE(n10708), .CLK(n11091), 
        .Q(test_so31), .QN(n10671) );
  SDFFX1 DFF_445_Q_reg ( .D(g34605), .SI(test_si32), .SE(n10749), .CLK(n11132), 
        .Q(g2145) );
  SDFFX1 DFF_446_Q_reg ( .D(g30350), .SI(g2145), .SE(n10723), .CLK(n11106), 
        .Q(g1700), .QN(n5417) );
  SDFFX1 DFF_447_Q_reg ( .D(g25611), .SI(g1700), .SE(n10771), .CLK(n11154), 
        .Q(g513) );
  SDFFX1 DFF_448_Q_reg ( .D(test_so9), .SI(g513), .SE(n10787), .CLK(n11170), 
        .Q(g2841), .QN(n5963) );
  SDFFX1 DFF_449_Q_reg ( .D(g33619), .SI(g2841), .SE(n10714), .CLK(n11097), 
        .Q(g5297), .QN(n5588) );
  SDFFX1 DFF_451_Q_reg ( .D(g34022), .SI(g5297), .SE(n10792), .CLK(n11175), 
        .Q(g2763), .QN(n10100) );
  SDFFX1 DFF_452_Q_reg ( .D(g34033), .SI(g2763), .SE(n10798), .CLK(n11181), 
        .Q(g4793), .QN(n5368) );
  SDFFX1 DFF_453_Q_reg ( .D(g34726), .SI(g4793), .SE(n10798), .CLK(n11181), 
        .Q(g952), .QN(n10094) );
  SDFFX1 DFF_454_Q_reg ( .D(g31870), .SI(g952), .SE(n10710), .CLK(n11093), .Q(
        g1263), .QN(n5674) );
  SDFFX1 DFF_455_Q_reg ( .D(g33985), .SI(g1263), .SE(n10757), .CLK(n11140), 
        .Q(g1950), .QN(n10199) );
  SDFFX1 DFF_456_Q_reg ( .D(g29283), .SI(g1950), .SE(n10714), .CLK(n11097), 
        .Q(g5138), .QN(n5871) );
  SDFFX1 DFF_457_Q_reg ( .D(g34003), .SI(g5138), .SE(n10768), .CLK(n11151), 
        .Q(g2307) );
  SDFFX1 DFF_458_Q_reg ( .D(g9497), .SI(g2307), .SE(n10768), .CLK(n11151), .Q(
        test_so32) );
  SDFFX1 DFF_460_Q_reg ( .D(g25677), .SI(test_si33), .SE(n10712), .CLK(n11095), 
        .Q(g8398) );
  SDFFX1 DFF_461_Q_reg ( .D(g34463), .SI(g8398), .SE(n10712), .CLK(n11095), 
        .Q(g4664) );
  SDFFX1 DFF_462_Q_reg ( .D(g33006), .SI(g4664), .SE(n10792), .CLK(n11175), 
        .Q(g2223), .QN(n5406) );
  SDFFX1 DFF_463_Q_reg ( .D(g29292), .SI(g2223), .SE(n10712), .CLK(n11095), 
        .Q(g5808), .QN(n5749) );
  SDFFX1 DFF_464_Q_reg ( .D(g30557), .SI(g5808), .SE(n10734), .CLK(n11117), 
        .Q(g6645), .QN(n10368) );
  SDFFX1 DFF_465_Q_reg ( .D(g33989), .SI(g6645), .SE(n10744), .CLK(n11127), 
        .Q(g2016) );
  SDFFX1 DFF_467_Q_reg ( .D(g33033), .SI(g2016), .SE(n10776), .CLK(n11159), 
        .Q(g3873), .QN(n5387) );
  SDFFX1 DFF_468_Q_reg ( .D(g11388), .SI(g3873), .SE(n10791), .CLK(n11174), 
        .Q(g13926), .QN(n5699) );
  SDFFX1 DFF_469_Q_reg ( .D(g34005), .SI(g13926), .SE(n10768), .CLK(n11151), 
        .Q(g2315), .QN(n5802) );
  SDFFX1 DFF_470_Q_reg ( .D(g26932), .SI(g2315), .SE(n10717), .CLK(n11100), 
        .Q(g2811), .QN(n10121) );
  SDFFX1 DFF_471_Q_reg ( .D(g30516), .SI(g2811), .SE(n10742), .CLK(n11125), 
        .Q(g5957), .QN(n10467) );
  SDFFX1 DFF_472_Q_reg ( .D(g33575), .SI(g5957), .SE(n10764), .CLK(n11147), 
        .Q(g2047), .QN(n5831) );
  SDFFX1 DFF_473_Q_reg ( .D(g33032), .SI(g2047), .SE(n10764), .CLK(n11147), 
        .Q(test_so33), .QN(n10647) );
  SDFFX1 DFF_474_Q_reg ( .D(g14779), .SI(test_si34), .SE(n10793), .CLK(n11176), 
        .Q(g17760), .QN(n10385) );
  SDFFX1 DFF_476_Q_reg ( .D(g30486), .SI(g17760), .SE(n10706), .CLK(n11089), 
        .Q(g5575), .QN(n10329) );
  SDFFX1 DFF_477_Q_reg ( .D(g34974), .SI(g5575), .SE(n10712), .CLK(n11095), 
        .Q(n9327) );
  SDFFX1 DFF_478_Q_reg ( .D(g25678), .SI(n9327), .SE(n10712), .CLK(n11095), 
        .Q(g3752) );
  SDFFX1 DFF_479_Q_reg ( .D(g30440), .SI(g3752), .SE(n10775), .CLK(n11158), 
        .Q(g3917), .QN(n10310) );
  SDFFX1 DFF_480_Q_reg ( .D(test_so86), .SI(g3917), .SE(n10737), .CLK(n11120), 
        .Q(g8783), .QN(DFF_480_n1) );
  SDFFX1 DFF_481_Q_reg ( .D(g12923), .SI(g8783), .SE(n10738), .CLK(n11121), 
        .Q(g1585), .QN(n5757) );
  SDFFX1 DFF_482_Q_reg ( .D(g26949), .SI(g1585), .SE(n10773), .CLK(n11156), 
        .Q(g4388), .QN(n10181) );
  SDFFX1 DFF_483_Q_reg ( .D(g30530), .SI(g4388), .SE(n10760), .CLK(n11143), 
        .Q(g6275), .QN(n10356) );
  SDFFX1 DFF_484_Q_reg ( .D(g30542), .SI(g6275), .SE(n10761), .CLK(n11144), 
        .Q(g6311), .QN(n10299) );
  SDFFX1 DFF_485_Q_reg ( .D(g8915), .SI(g6311), .SE(n10761), .CLK(n11144), .Q(
        g8916), .QN(n19406) );
  SDFFX1 DFF_486_Q_reg ( .D(g25624), .SI(g8916), .SE(n10764), .CLK(n11147), 
        .Q(g1041), .QN(n10104) );
  SDFFX1 DFF_487_Q_reg ( .D(g30383), .SI(g1041), .SE(n10728), .CLK(n11111), 
        .Q(test_so34), .QN(n10679) );
  SDFFX1 DFF_488_Q_reg ( .D(g33597), .SI(test_si35), .SE(n10717), .CLK(n11100), 
        .Q(g2537), .QN(n5411) );
  SDFFX1 DFF_489_Q_reg ( .D(g34598), .SI(g2537), .SE(n10746), .CLK(n11129), 
        .Q(g29221), .QN(g23612) );
  SDFFX1 DFF_490_Q_reg ( .D(g26957), .SI(g29221), .SE(n10746), .CLK(n11129), 
        .Q(g4430), .QN(n10184) );
  SDFFX1 DFF_491_Q_reg ( .D(g26967), .SI(g4430), .SE(n10798), .CLK(n11181), 
        .Q(n9325), .QN(n19399) );
  SDFFX1 DFF_493_Q_reg ( .D(g28102), .SI(n9325), .SE(n10761), .CLK(n11144), 
        .Q(g4826) );
  SDFFX1 DFF_494_Q_reg ( .D(g30524), .SI(g4826), .SE(n10761), .CLK(n11144), 
        .Q(g6239), .QN(n10302) );
  SDFFX1 DFF_496_Q_reg ( .D(g26903), .SI(g6239), .SE(n10801), .CLK(n11184), 
        .Q(g232), .QN(n10399) );
  SDFFX1 DFF_497_Q_reg ( .D(g30475), .SI(g232), .SE(n10715), .CLK(n11098), .Q(
        g5268), .QN(n10336) );
  SDFFX1 DFF_498_Q_reg ( .D(g34647), .SI(g5268), .SE(n10715), .CLK(n11098), 
        .Q(g6545), .QN(n5497) );
  SDFFX1 DFF_499_Q_reg ( .D(g30377), .SI(g6545), .SE(n10708), .CLK(n11091), 
        .Q(n9324), .QN(n19403) );
  SDFFX1 DFF_500_Q_reg ( .D(g33553), .SI(n9324), .SE(n10708), .CLK(n11091), 
        .Q(g1772), .QN(n5504) );
  SDFFX1 DFF_502_Q_reg ( .D(g31903), .SI(g1772), .SE(n10769), .CLK(n11152), 
        .Q(g5052), .QN(n5607) );
  SDFFX1 DFF_503_Q_reg ( .D(g25715), .SI(g5052), .SE(n10769), .CLK(n11152), 
        .Q(test_so35) );
  SDFFX1 DFF_504_Q_reg ( .D(g33984), .SI(test_si36), .SE(n10758), .CLK(n11141), 
        .Q(g1890), .QN(n5799) );
  SDFFX1 DFF_505_Q_reg ( .D(g33602), .SI(g1890), .SE(n10797), .CLK(n11180), 
        .Q(g2629), .QN(n5521) );
  SDFFX1 DFF_506_Q_reg ( .D(g28045), .SI(g2629), .SE(n10749), .CLK(n11132), 
        .Q(g572), .QN(n5337) );
  SDFFX1 DFF_507_Q_reg ( .D(g34603), .SI(g572), .SE(n10749), .CLK(n11132), .Q(
        g2130), .QN(n5487) );
  SDFFX1 DFF_508_Q_reg ( .D(g33035), .SI(g2130), .SE(n10775), .CLK(n11158), 
        .Q(g4108) );
  SDFFX1 DFF_509_Q_reg ( .D(g9251), .SI(g4108), .SE(n10775), .CLK(n11158), .Q(
        g4308) );
  SDFFX1 DFF_510_Q_reg ( .D(g24208), .SI(g4308), .SE(n10770), .CLK(n11153), 
        .Q(g475), .QN(n10124) );
  SDFFX1 DFF_511_Q_reg ( .D(g8416), .SI(g475), .SE(n10770), .CLK(n11153), .Q(
        g990), .QN(n5622) );
  SDFFX1 DFF_512_Q_reg ( .D(g34971), .SI(g990), .SE(n10770), .CLK(n11153), .Q(
        g31), .QN(n5469) );
  SDFFX1 DFF_514_Q_reg ( .D(g34970), .SI(g31), .SE(n10702), .CLK(n11085), .Q(
        n9322) );
  SDFFX1 DFF_515_Q_reg ( .D(n473), .SI(n9322), .SE(n10702), .CLK(n11085), .Q(
        g12184) );
  SDFFX1 DFF_517_Q_reg ( .D(g33614), .SI(g12184), .SE(n10702), .CLK(n11085), 
        .Q(g3990) );
  SDFFX1 DFF_519_Q_reg ( .D(g33060), .SI(g3990), .SE(n10785), .CLK(n11168), 
        .Q(test_so36), .QN(n10651) );
  SDFFX1 DFF_520_Q_reg ( .D(g30362), .SI(test_si37), .SE(n10754), .CLK(n11137), 
        .Q(g1992), .QN(n5890) );
  SDFFX1 DFF_522_Q_reg ( .D(g33023), .SI(g1992), .SE(n10754), .CLK(n11137), 
        .Q(g3171), .QN(n5603) );
  SDFFX1 DFF_524_Q_reg ( .D(g26898), .SI(g3171), .SE(n10745), .CLK(n11128), 
        .Q(g812), .QN(n5733) );
  SDFFX1 DFF_525_Q_reg ( .D(g25618), .SI(g812), .SE(n10799), .CLK(n11182), .Q(
        g832), .QN(n10544) );
  SDFFX1 DFF_526_Q_reg ( .D(g30518), .SI(g832), .SE(n10752), .CLK(n11135), .Q(
        g5897) );
  SDFFX1 DFF_527_Q_reg ( .D(g25688), .SI(g5897), .SE(n10752), .CLK(n11135), 
        .Q(g25689), .QN(n10133) );
  SDFFX1 DFF_528_Q_reg ( .D(g4570), .SI(g25689), .SE(n10782), .CLK(n11165), 
        .Q(g4571) );
  SDFFX1 DFF_529_Q_reg ( .D(g11349), .SI(g4571), .SE(n10782), .CLK(n11165), 
        .Q(g13895), .QN(n5702) );
  SDFFX1 DFF_530_Q_reg ( .D(g26959), .SI(g13895), .SE(n10782), .CLK(n11165), 
        .Q(g4455) );
  SDFFX1 DFF_531_Q_reg ( .D(g34801), .SI(g4455), .SE(n10712), .CLK(n11095), 
        .Q(g2902), .QN(n10615) );
  SDFFX1 DFF_532_Q_reg ( .D(g26884), .SI(g2902), .SE(n10781), .CLK(n11164), 
        .Q(g333) );
  SDFFX1 DFF_533_Q_reg ( .D(g25600), .SI(g333), .SE(n10735), .CLK(n11118), .Q(
        g168), .QN(n5606) );
  SDFFX1 DFF_534_Q_reg ( .D(g26933), .SI(g168), .SE(n10717), .CLK(n11100), .Q(
        test_so37), .QN(n10666) );
  SDFFX1 DFF_535_Q_reg ( .D(g28066), .SI(test_si38), .SE(n10788), .CLK(n11171), 
        .Q(g3684), .QN(n5881) );
  SDFFX1 DFF_536_Q_reg ( .D(g33612), .SI(g3684), .SE(n10738), .CLK(n11121), 
        .Q(g3639) );
  SDFFX1 DFF_537_Q_reg ( .D(g17787), .SI(g3639), .SE(n10786), .CLK(n11169), 
        .Q(g14597), .QN(n5579) );
  SDFFX1 DFF_538_Q_reg ( .D(g24268), .SI(g14597), .SE(n10786), .CLK(n11169), 
        .Q(g3338), .QN(n5527) );
  SDFFX1 DFF_539_Q_reg ( .D(g25716), .SI(g3338), .SE(n10769), .CLK(n11152), 
        .Q(g5406) );
  SDFFX1 DFF_541_Q_reg ( .D(g26906), .SI(g5406), .SE(n10770), .CLK(n11153), 
        .Q(g269), .QN(n10277) );
  SDFFX1 DFF_542_Q_reg ( .D(g24203), .SI(g269), .SE(n10710), .CLK(n11093), .Q(
        g401), .QN(n10228) );
  SDFFX1 DFF_543_Q_reg ( .D(g24346), .SI(g401), .SE(n10725), .CLK(n11108), .Q(
        g6040), .QN(n10391) );
  SDFFX1 DFF_544_Q_reg ( .D(g24207), .SI(g6040), .SE(n10770), .CLK(n11153), 
        .Q(g441) );
  SDFFX1 DFF_545_Q_reg ( .D(g25701), .SI(g441), .SE(n10793), .CLK(n11176), .Q(
        g9553), .QN(n5690) );
  SDFFX1 DFF_546_Q_reg ( .D(g29269), .SI(g9553), .SE(n10700), .CLK(n11083), 
        .Q(g3808), .QN(n5745) );
  SDFFX1 DFF_547_Q_reg ( .D(g34976), .SI(g3808), .SE(n10701), .CLK(n11084), 
        .Q(g9), .QN(n5468) );
  SDFFX1 DFF_549_Q_reg ( .D(g34255), .SI(g9), .SE(n10781), .CLK(n11164), .Q(
        test_so38), .QN(n10656) );
  SDFFX1 DFF_550_Q_reg ( .D(g30450), .SI(test_si39), .SE(n10731), .CLK(n11114), 
        .Q(g3957), .QN(n10476) );
  SDFFX1 DFF_551_Q_reg ( .D(g30456), .SI(g3957), .SE(n10776), .CLK(n11159), 
        .Q(g4093), .QN(n5340) );
  SDFFX1 DFF_552_Q_reg ( .D(g32991), .SI(g4093), .SE(n10764), .CLK(n11147), 
        .Q(g1760), .QN(n5602) );
  SDFFX1 DFF_554_Q_reg ( .D(g24348), .SI(g1760), .SE(n10793), .CLK(n11176), 
        .Q(g12422), .QN(n5437) );
  SDFFX1 DFF_555_Q_reg ( .D(g34249), .SI(g12422), .SE(n10711), .CLK(n11094), 
        .Q(g160), .QN(n5843) );
  SDFFX1 DFF_558_Q_reg ( .D(g30371), .SI(g160), .SE(n10734), .CLK(n11117), .Q(
        g2279), .QN(n5778) );
  SDFFX1 DFF_559_Q_reg ( .D(g29268), .SI(g2279), .SE(n10777), .CLK(n11160), 
        .Q(g3498) );
  SDFFX1 DFF_560_Q_reg ( .D(g29224), .SI(g3498), .SE(n10749), .CLK(n11132), 
        .Q(g586), .QN(n5336) );
  SDFFX1 DFF_561_Q_reg ( .D(g14189), .SI(g586), .SE(n10753), .CLK(n11136), .Q(
        g14201), .QN(n10106) );
  SDFFX1 DFF_562_Q_reg ( .D(g33017), .SI(g14201), .SE(n10729), .CLK(n11112), 
        .Q(g2619), .QN(n5508) );
  SDFFX1 DFF_563_Q_reg ( .D(g30339), .SI(g2619), .SE(n10757), .CLK(n11140), 
        .Q(g1183), .QN(n5599) );
  SDFFX1 DFF_564_Q_reg ( .D(g33967), .SI(g1183), .SE(n10737), .CLK(n11120), 
        .Q(g1608), .QN(n5792) );
  SDFFX1 DFF_565_Q_reg ( .D(g8784), .SI(g1608), .SE(n10737), .CLK(n11120), .Q(
        test_so39), .QN(n10262) );
  SDFFX1 DFF_566_Q_reg ( .D(g17519), .SI(test_si40), .SE(n10786), .CLK(n11169), 
        .Q(g17577), .QN(n10463) );
  SDFFX1 DFF_567_Q_reg ( .D(g33559), .SI(g17577), .SE(n10787), .CLK(n11170), 
        .Q(g1779), .QN(n5830) );
  SDFFX1 DFF_568_Q_reg ( .D(n466), .SI(g1779), .SE(n10716), .CLK(n11099), .Q(
        g2652), .QN(n10324) );
  SDFFX1 DFF_570_Q_reg ( .D(g30368), .SI(g2652), .SE(n10716), .CLK(n11099), 
        .Q(g2193), .QN(n5839) );
  SDFFX1 DFF_571_Q_reg ( .D(g30375), .SI(g2193), .SE(n10708), .CLK(n11091), 
        .Q(g2393), .QN(n5421) );
  SDFFX1 DFF_573_Q_reg ( .D(g28052), .SI(g2393), .SE(n10718), .CLK(n11101), 
        .Q(g661), .QN(n10282) );
  SDFFX1 DFF_574_Q_reg ( .D(g28089), .SI(g661), .SE(n10738), .CLK(n11121), .Q(
        g4950), .QN(n5772) );
  SDFFX1 DFF_575_Q_reg ( .D(g33055), .SI(g4950), .SE(n10783), .CLK(n11166), 
        .Q(g5535), .QN(n5566) );
  SDFFX1 DFF_576_Q_reg ( .D(g30392), .SI(g5535), .SE(n10707), .CLK(n11090), 
        .Q(g2834), .QN(g23652) );
  SDFFX1 DFF_577_Q_reg ( .D(g30343), .SI(g2834), .SE(n10707), .CLK(n11090), 
        .Q(g1361), .QN(n10258) );
  SDFFX1 DFF_579_Q_reg ( .D(g30523), .SI(g1361), .SE(n10778), .CLK(n11161), 
        .Q(g6235), .QN(n10454) );
  SDFFX1 DFF_580_Q_reg ( .D(g24233), .SI(g6235), .SE(n10757), .CLK(n11140), 
        .Q(g1146), .QN(n5851) );
  SDFFX1 DFF_581_Q_reg ( .D(g33018), .SI(g1146), .SE(n10728), .CLK(n11111), 
        .Q(test_so40), .QN(n10653) );
  SDFFX1 DFF_582_Q_reg ( .D(g32976), .SI(test_si41), .SE(n10711), .CLK(n11094), 
        .Q(g150), .QN(n5676) );
  SDFFX1 DFF_583_Q_reg ( .D(g30349), .SI(g150), .SE(n10723), .CLK(n11106), .Q(
        g1696), .QN(n5628) );
  SDFFX1 DFF_584_Q_reg ( .D(g33067), .SI(g1696), .SE(n10776), .CLK(n11159), 
        .Q(g6555), .QN(n10592) );
  SDFFX1 DFF_585_Q_reg ( .D(g26900), .SI(g6555), .SE(n10753), .CLK(n11136), 
        .Q(g14189), .QN(n10112) );
  SDFFX1 DFF_587_Q_reg ( .D(g33034), .SI(g14189), .SE(n10776), .CLK(n11159), 
        .Q(g3881), .QN(n5564) );
  SDFFX1 DFF_588_Q_reg ( .D(g30551), .SI(g3881), .SE(n10735), .CLK(n11118), 
        .Q(g6621), .QN(n10350) );
  SDFFX1 DFF_589_Q_reg ( .D(g25667), .SI(g6621), .SE(n10720), .CLK(n11103), 
        .Q(g3470), .QN(n5424) );
  SDFFX1 DFF_590_Q_reg ( .D(g30452), .SI(g3470), .SE(n10795), .CLK(n11178), 
        .Q(g3897), .QN(n10448) );
  SDFFX1 DFF_593_Q_reg ( .D(g34719), .SI(g518), .SE(n10795), .CLK(n11178), .Q(
        g538), .QN(n5491) );
  SDFFX1 DFF_594_Q_reg ( .D(g33607), .SI(g538), .SE(n10728), .CLK(n11111), .Q(
        g2606), .QN(n5311) );
  SDFFX1 DFF_595_Q_reg ( .D(g26923), .SI(g2606), .SE(n10727), .CLK(n11110), 
        .Q(g1472), .QN(n5290) );
  SDFFX1 DFF_597_Q_reg ( .D(g24211), .SI(g1472), .SE(n10746), .CLK(n11129), 
        .Q(test_so41), .QN(n10670) );
  SDFFX1 DFF_598_Q_reg ( .D(g33050), .SI(test_si42), .SE(n10779), .CLK(n11162), 
        .Q(g5188), .QN(n5567) );
  SDFFX1 DFF_599_Q_reg ( .D(g24341), .SI(g5188), .SE(n10796), .CLK(n11179), 
        .Q(g5689), .QN(n5529) );
  SDFFX1 DFF_600_Q_reg ( .D(g19334), .SI(g5689), .SE(n10796), .CLK(n11179), 
        .Q(g13259), .QN(n10243) );
  SDFFX1 DFF_601_Q_reg ( .D(g24201), .SI(g13259), .SE(n10797), .CLK(n11180), 
        .Q(g405), .QN(n10247) );
  SDFFX1 DFF_602_Q_reg ( .D(g30463), .SI(g405), .SE(n10715), .CLK(n11098), .Q(
        g5216), .QN(n10412) );
  SDFFX1 DFF_603_Q_reg ( .D(g9743), .SI(g5216), .SE(n10781), .CLK(n11164), .Q(
        g6494) );
  SDFFX1 DFF_604_Q_reg ( .D(g34464), .SI(g6494), .SE(n10712), .CLK(n11095), 
        .Q(g4669), .QN(n10103) );
  SDFFX1 DFF_606_Q_reg ( .D(g24243), .SI(g4669), .SE(n10766), .CLK(n11149), 
        .Q(g996), .QN(n10255) );
  SDFFX1 DFF_607_Q_reg ( .D(g24335), .SI(g996), .SE(n10801), .CLK(n11184), .Q(
        g4531) );
  SDFFX1 DFF_608_Q_reg ( .D(g34611), .SI(g4531), .SE(n10743), .CLK(n11126), 
        .Q(g2860) );
  SDFFX1 DFF_609_Q_reg ( .D(g34262), .SI(g2860), .SE(n10713), .CLK(n11096), 
        .Q(g4743), .QN(n5876) );
  SDFFX1 DFF_610_Q_reg ( .D(g30546), .SI(g4743), .SE(n10735), .CLK(n11118), 
        .Q(g6593), .QN(n10512) );
  SDFFX1 DFF_612_Q_reg ( .D(g25591), .SI(g6593), .SE(n10795), .CLK(n11178), 
        .Q(test_so42) );
  SDFFX1 DFF_613_Q_reg ( .D(g7257), .SI(test_si43), .SE(n10772), .CLK(n11155), 
        .Q(g4411), .QN(n10095) );
  SDFFX1 DFF_614_Q_reg ( .D(g30347), .SI(g4411), .SE(n10748), .CLK(n11131), 
        .Q(g1413), .QN(n10090) );
  SDFFX1 DFF_615_Q_reg ( .D(test_so38), .SI(g1413), .SE(n10781), .CLK(n11164), 
        .Q(g26960), .QN(n10281) );
  SDFFX1 DFF_616_Q_reg ( .D(g17577), .SI(g26960), .SE(n10786), .CLK(n11169), 
        .Q(g13039), .QN(n10442) );
  SDFFX1 DFF_617_Q_reg ( .D(g30556), .SI(g13039), .SE(n10795), .CLK(n11178), 
        .Q(g6641), .QN(n10293) );
  SDFFX1 DFF_619_Q_reg ( .D(g34970), .SI(g6641), .SE(n10795), .CLK(n11178), 
        .Q(g6) );
  SDFFX1 DFF_620_Q_reg ( .D(g33562), .SI(g6), .SE(n10771), .CLK(n11154), .Q(
        g1936), .QN(n5534) );
  SDFFX1 DFF_621_Q_reg ( .D(n35), .SI(g1936), .SE(n10771), .CLK(n11154), .Q(
        g55) );
  SDFFX1 DFF_622_Q_reg ( .D(g25610), .SI(g55), .SE(n10771), .CLK(n11154), .Q(
        g504), .QN(n5519) );
  SDFFX1 DFF_623_Q_reg ( .D(g33015), .SI(g504), .SE(n10729), .CLK(n11112), .Q(
        g2587), .QN(n5372) );
  SDFFX1 DFF_624_Q_reg ( .D(g31896), .SI(g2587), .SE(n10784), .CLK(n11167), 
        .Q(g4480) );
  SDFFX1 DFF_625_Q_reg ( .D(g34004), .SI(g4480), .SE(n10768), .CLK(n11151), 
        .Q(n9314), .QN(n19412) );
  SDFFX1 DFF_626_Q_reg ( .D(g30428), .SI(n9314), .SE(n10732), .CLK(n11115), 
        .Q(test_so43), .QN(n10664) );
  SDFFX1 DFF_627_Q_reg ( .D(g30485), .SI(test_si44), .SE(n10705), .CLK(n11088), 
        .Q(g5571), .QN(n10290) );
  SDFFX1 DFF_628_Q_reg ( .D(g30422), .SI(g5571), .SE(n10720), .CLK(n11103), 
        .Q(g3578), .QN(n10353) );
  SDFFX1 DFF_630_Q_reg ( .D(g25714), .SI(g3578), .SE(n10783), .CLK(n11166), 
        .Q(g9555), .QN(n19405) );
  SDFFX1 DFF_632_Q_reg ( .D(n201), .SI(g9555), .SE(n10713), .CLK(n11096), .Q(
        g5827), .QN(n5809) );
  SDFFX1 DFF_633_Q_reg ( .D(g30423), .SI(g5827), .SE(n10763), .CLK(n11146), 
        .Q(g3582), .QN(n10437) );
  SDFFX1 DFF_634_Q_reg ( .D(g30529), .SI(g3582), .SE(n10762), .CLK(n11145), 
        .Q(g6271), .QN(n10429) );
  SDFFX1 DFF_635_Q_reg ( .D(g34028), .SI(g6271), .SE(n10796), .CLK(n11179), 
        .Q(g4688), .QN(n5656) );
  SDFFX1 DFF_637_Q_reg ( .D(g33587), .SI(g4688), .SE(n10707), .CLK(n11090), 
        .Q(g2380), .QN(n10162) );
  SDFFX1 DFF_638_Q_reg ( .D(g30460), .SI(g2380), .SE(n10779), .CLK(n11162), 
        .Q(g5196), .QN(n10443) );
  SDFFX1 DFF_640_Q_reg ( .D(g30401), .SI(g5196), .SE(n10719), .CLK(n11102), 
        .Q(g3227), .QN(n10335) );
  SDFFX1 DFF_641_Q_reg ( .D(g33990), .SI(g3227), .SE(n10744), .CLK(n11127), 
        .Q(n9312), .QN(n19413) );
  SDFFX1 DFF_642_Q_reg ( .D(g16693), .SI(n9312), .SE(n10774), .CLK(n11157), 
        .Q(g14518), .QN(n10507) );
  SDFFX1 DFF_643_Q_reg ( .D(g17291), .SI(g14518), .SE(n10756), .CLK(n11139), 
        .Q(test_so44) );
  SDFFX1 DFF_644_Q_reg ( .D(g29309), .SI(test_si45), .SE(n10756), .CLK(n11139), 
        .Q(g6541) );
  SDFFX1 DFF_645_Q_reg ( .D(g30411), .SI(g6541), .SE(n10722), .CLK(n11105), 
        .Q(g3203) );
  SDFFX1 DFF_646_Q_reg ( .D(g33546), .SI(g3203), .SE(n10722), .CLK(n11105), 
        .Q(g1668), .QN(n5598) );
  SDFFX1 DFF_647_Q_reg ( .D(g28085), .SI(g1668), .SE(n10726), .CLK(n11109), 
        .Q(g4760), .QN(n5775) );
  SDFFX1 DFF_648_Q_reg ( .D(g26904), .SI(g4760), .SE(n10726), .CLK(n11109), 
        .Q(g262), .QN(n10276) );
  SDFFX1 DFF_649_Q_reg ( .D(n45), .SI(g262), .SE(n10741), .CLK(n11124), .Q(
        g1840), .QN(n5451) );
  SDFFX1 DFF_651_Q_reg ( .D(g25722), .SI(g1840), .SE(n10732), .CLK(n11115), 
        .Q(g5467) );
  SDFFX1 DFF_652_Q_reg ( .D(g25605), .SI(g5467), .SE(n10732), .CLK(n11115), 
        .Q(g460), .QN(n10167) );
  SDFFX1 DFF_653_Q_reg ( .D(g33062), .SI(g460), .SE(n10777), .CLK(n11160), .Q(
        g6209), .QN(n10588) );
  SDFFX1 DFF_654_Q_reg ( .D(g26893), .SI(g6209), .SE(n10797), .CLK(n11180), 
        .Q(g29211) );
  SDFFX1 DFF_655_Q_reg ( .D(g12238), .SI(g29211), .SE(n10797), .CLK(n11180), 
        .Q(g14662), .QN(n5704) );
  SDFFX1 DFF_656_Q_reg ( .D(g28050), .SI(g14662), .SE(n10711), .CLK(n11094), 
        .Q(g655), .QN(n10313) );
  SDFFX1 DFF_657_Q_reg ( .D(n1052), .SI(g655), .SE(n10711), .CLK(n11094), .Q(
        test_so45), .QN(n10691) );
  SDFFX1 DFF_658_Q_reg ( .D(g33583), .SI(test_si46), .SE(n10774), .CLK(n11157), 
        .Q(g2204), .QN(n5620) );
  SDFFX1 DFF_659_Q_reg ( .D(g30472), .SI(g2204), .SE(n10774), .CLK(n11157), 
        .Q(g5256), .QN(n10304) );
  SDFFX1 DFF_660_Q_reg ( .D(g34454), .SI(g5256), .SE(n10798), .CLK(n11181), 
        .Q(g4608), .QN(n5274) );
  SDFFX1 DFF_661_Q_reg ( .D(g34850), .SI(g4608), .SE(n10767), .CLK(n11150), 
        .Q(g794), .QN(n5291) );
  SDFFX1 DFF_662_Q_reg ( .D(g16955), .SI(g794), .SE(n10780), .CLK(n11163), .Q(
        g13906), .QN(n5583) );
  SDFFX1 DFF_663_Q_reg ( .D(g10306), .SI(g13906), .SE(n10726), .CLK(n11109), 
        .Q(g4423), .QN(n10192) );
  SDFFX1 DFF_664_Q_reg ( .D(g24272), .SI(g4423), .SE(n10747), .CLK(n11130), 
        .Q(g3689), .QN(n5532) );
  SDFFX1 DFF_666_Q_reg ( .D(g17678), .SI(g3689), .SE(n10796), .CLK(n11179), 
        .Q(g5685) );
  SDFFX1 DFF_667_Q_reg ( .D(g24214), .SI(g5685), .SE(n10745), .CLK(n11128), 
        .Q(g703), .QN(n5821) );
  SDFFX1 DFF_669_Q_reg ( .D(g26909), .SI(g703), .SE(n10785), .CLK(n11168), .Q(
        g862), .QN(n5682) );
  SDFFX1 DFF_670_Q_reg ( .D(g30406), .SI(g862), .SE(n10790), .CLK(n11173), .Q(
        g3247), .QN(n10285) );
  SDFFX1 DFF_671_Q_reg ( .D(g33569), .SI(g3247), .SE(n10751), .CLK(n11134), 
        .Q(g2040) );
  SDFFX1 DFF_672_Q_reg ( .D(g25694), .SI(g2040), .SE(n10751), .CLK(n11134), 
        .Q(test_so46) );
  SDFFX1 DFF_673_Q_reg ( .D(g34628), .SI(test_si47), .SE(n10739), .CLK(n11122), 
        .Q(g4146), .QN(n5981) );
  SDFFX1 DFF_674_Q_reg ( .D(g34458), .SI(g4146), .SE(n10757), .CLK(n11140), 
        .Q(g4633), .QN(n5844) );
  SDFFX1 DFF_675_Q_reg ( .D(g24240), .SI(g4633), .SE(n10757), .CLK(n11140), 
        .Q(g7916), .QN(n5304) );
  SDFFX1 DFF_677_Q_reg ( .D(g34634), .SI(g7916), .SE(n10757), .CLK(n11140), 
        .Q(g4732), .QN(n5296) );
  SDFFX1 DFF_678_Q_reg ( .D(g25700), .SI(g4732), .SE(n10779), .CLK(n11162), 
        .Q(g9497), .QN(n5689) );
  SDFFX1 DFF_679_Q_reg ( .D(g29293), .SI(g9497), .SE(n10712), .CLK(n11095), 
        .Q(g5817), .QN(n10131) );
  SDFFX1 DFF_681_Q_reg ( .D(g33009), .SI(g5817), .SE(n10729), .CLK(n11112), 
        .Q(g2351), .QN(n5511) );
  SDFFX1 DFF_682_Q_reg ( .D(g33603), .SI(g2351), .SE(n10716), .CLK(n11099), 
        .Q(g2648), .QN(n10166) );
  SDFFX1 DFF_683_Q_reg ( .D(g24355), .SI(g2648), .SE(n10730), .CLK(n11113), 
        .Q(g6736), .QN(n10523) );
  SDFFX1 DFF_684_Q_reg ( .D(g34268), .SI(g6736), .SE(n10738), .CLK(n11121), 
        .Q(g4944), .QN(n5875) );
  SDFFX1 DFF_685_Q_reg ( .D(g25691), .SI(g4944), .SE(n10739), .CLK(n11122), 
        .Q(g4072), .QN(n10612) );
  SDFFX1 DFF_686_Q_reg ( .D(g26890), .SI(g4072), .SE(n10781), .CLK(n11164), 
        .Q(g7540), .QN(n10126) );
  SDFFX1 DFF_687_Q_reg ( .D(g7260), .SI(g7540), .SE(n10794), .CLK(n11177), .Q(
        test_so47) );
  SDFFX1 DFF_688_Q_reg ( .D(g29264), .SI(test_si48), .SE(n10720), .CLK(n11103), 
        .Q(g3466), .QN(n10149) );
  SDFFX1 DFF_689_Q_reg ( .D(g28072), .SI(g3466), .SE(n10786), .CLK(n11169), 
        .Q(g4116), .QN(n10102) );
  SDFFX1 DFF_690_Q_reg ( .D(g31900), .SI(g4116), .SE(n10769), .CLK(n11152), 
        .Q(g5041), .QN(n5605) );
  SDFFX1 DFF_692_Q_reg ( .D(g26956), .SI(g5041), .SE(n10794), .CLK(n11177), 
        .Q(g4434), .QN(n10180) );
  SDFFX1 DFF_693_Q_reg ( .D(g29271), .SI(g4434), .SE(n10700), .CLK(n11083), 
        .Q(g3827), .QN(n5808) );
  SDFFX1 DFF_694_Q_reg ( .D(g29304), .SI(g3827), .SE(n10726), .CLK(n11109), 
        .Q(g6500), .QN(n5748) );
  SDFFX1 DFF_695_Q_reg ( .D(g13049), .SI(g6500), .SE(n10774), .CLK(n11157), 
        .Q(g17813) );
  SDFFX1 DFF_696_Q_reg ( .D(g29261), .SI(g17813), .SE(n10703), .CLK(n11086), 
        .Q(g3133), .QN(n5661) );
  SDFFX1 DFF_697_Q_reg ( .D(g28063), .SI(g3133), .SE(n10719), .CLK(n11102), 
        .Q(g3333) );
  SDFFX1 DFF_698_Q_reg ( .D(g13259), .SI(g3333), .SE(n10796), .CLK(n11179), 
        .Q(g979), .QN(n5320) );
  SDFFX1 DFF_699_Q_reg ( .D(g34027), .SI(g979), .SE(n10796), .CLK(n11179), .Q(
        g4681), .QN(n10527) );
  SDFFX1 DFF_700_Q_reg ( .D(g33961), .SI(g4681), .SE(n10711), .CLK(n11094), 
        .Q(g298), .QN(n5675) );
  SDFFX1 DFF_702_Q_reg ( .D(g33604), .SI(g298), .SE(n10706), .CLK(n11089), .Q(
        test_so48), .QN(n10676) );
  SDFFX1 DFF_704_Q_reg ( .D(g8788), .SI(test_si49), .SE(n10773), .CLK(n11156), 
        .Q(g8789), .QN(n10264) );
  SDFFX1 DFF_705_Q_reg ( .D(g32995), .SI(g8789), .SE(n10758), .CLK(n11141), 
        .Q(g1894), .QN(n5374) );
  SDFFX1 DFF_706_Q_reg ( .D(g34624), .SI(g1894), .SE(n10743), .CLK(n11126), 
        .Q(g2988), .QN(n10582) );
  SDFFX1 DFF_707_Q_reg ( .D(g30415), .SI(g2988), .SE(n10762), .CLK(n11145), 
        .Q(g3538), .QN(n10452) );
  SDFFX1 DFF_708_Q_reg ( .D(g33536), .SI(g3538), .SE(n10712), .CLK(n11095), 
        .Q(g301), .QN(n10614) );
  SDFFX1 DFF_709_Q_reg ( .D(g26888), .SI(g301), .SE(n10802), .CLK(n11185), .Q(
        n9306) );
  SDFFX1 DFF_710_Q_reg ( .D(g28055), .SI(n9306), .SE(n10745), .CLK(n11128), 
        .Q(g827), .QN(n5728) );
  SDFFX1 DFF_711_Q_reg ( .D(g24238), .SI(g827), .SE(n10756), .CLK(n11139), .Q(
        g17291), .QN(n10218) );
  SDFFX1 DFF_713_Q_reg ( .D(g33600), .SI(g17291), .SE(n10797), .CLK(n11180), 
        .Q(g2555), .QN(n5351) );
  SDFFX1 DFF_714_Q_reg ( .D(g28105), .SI(g2555), .SE(n10721), .CLK(n11104), 
        .Q(g5011), .QN(n10174) );
  SDFFX1 DFF_715_Q_reg ( .D(g34721), .SI(g5011), .SE(n10721), .CLK(n11104), 
        .Q(g199), .QN(n10572) );
  SDFFX1 DFF_716_Q_reg ( .D(g29307), .SI(g199), .SE(n10721), .CLK(n11104), .Q(
        g6523) );
  SDFFX1 DFF_717_Q_reg ( .D(g30345), .SI(g6523), .SE(n10762), .CLK(n11145), 
        .Q(test_so49), .QN(n10662) );
  SDFFX1 DFF_718_Q_reg ( .D(g34453), .SI(test_si50), .SE(n10798), .CLK(n11181), 
        .Q(g4601), .QN(n5365) );
  SDFFX1 DFF_719_Q_reg ( .D(g32980), .SI(g4601), .SE(n10798), .CLK(n11181), 
        .Q(g854), .QN(n5754) );
  SDFFX1 DFF_720_Q_reg ( .D(g29238), .SI(g854), .SE(n10733), .CLK(n11116), .Q(
        g1484), .QN(n5865) );
  SDFFX1 DFF_721_Q_reg ( .D(g34639), .SI(g1484), .SE(n10733), .CLK(n11116), 
        .Q(g4922), .QN(n5346) );
  SDFFX1 DFF_722_Q_reg ( .D(g25695), .SI(g4922), .SE(n10699), .CLK(n11082), 
        .Q(g5080), .QN(n5893) );
  SDFFX1 DFF_723_Q_reg ( .D(g33057), .SI(g5080), .SE(n10784), .CLK(n11167), 
        .Q(g5863), .QN(n10590) );
  SDFFX1 DFF_724_Q_reg ( .D(g26969), .SI(g5863), .SE(n10784), .CLK(n11167), 
        .Q(g4581), .QN(n5670) );
  SDFFX1 DFF_726_Q_reg ( .D(n643), .SI(g4581), .SE(n10717), .CLK(n11100), .Q(
        g2518), .QN(n10323) );
  SDFFX1 DFF_727_Q_reg ( .D(g34021), .SI(g2518), .SE(n10716), .CLK(n11099), 
        .Q(g2567), .QN(n10134) );
  SDFFX1 DFF_728_Q_reg ( .D(g26895), .SI(g2567), .SE(n10750), .CLK(n11133), 
        .Q(g568), .QN(n5335) );
  SDFFX1 DFF_729_Q_reg ( .D(g30413), .SI(g568), .SE(n10719), .CLK(n11102), .Q(
        g3263), .QN(n10284) );
  SDFFX1 DFF_730_Q_reg ( .D(g30549), .SI(g3263), .SE(n10734), .CLK(n11117), 
        .Q(g6613), .QN(n10331) );
  SDFFX1 DFF_731_Q_reg ( .D(g24347), .SI(g6613), .SE(n10725), .CLK(n11108), 
        .Q(test_so50), .QN(n10694) );
  SDFFX1 DFF_732_Q_reg ( .D(g25758), .SI(test_si51), .SE(n10790), .CLK(n11173), 
        .Q(g6444) );
  SDFFX1 DFF_733_Q_reg ( .D(g34808), .SI(g6444), .SE(n10700), .CLK(n11083), 
        .Q(g2965), .QN(n10231) );
  SDFFX1 DFF_734_Q_reg ( .D(g30501), .SI(g2965), .SE(n10784), .CLK(n11167), 
        .Q(g5857), .QN(n5573) );
  SDFFX1 DFF_735_Q_reg ( .D(g33969), .SI(g5857), .SE(n10723), .CLK(n11106), 
        .Q(n9303), .QN(n19414) );
  SDFFX1 DFF_736_Q_reg ( .D(g34440), .SI(n9303), .SE(n10709), .CLK(n11092), 
        .Q(g890), .QN(n5305) );
  SDFFX1 DFF_737_Q_reg ( .D(g17607), .SI(g890), .SE(n10760), .CLK(n11143), .Q(
        g17646), .QN(n10468) );
  SDFFX1 DFF_738_Q_reg ( .D(g30433), .SI(g17646), .SE(n10733), .CLK(n11116), 
        .Q(g3562) );
  SDFFX1 DFF_739_Q_reg ( .D(g21900), .SI(g3562), .SE(n10733), .CLK(n11116), 
        .Q(g10122_Tj) );
  SDFFX1 DFF_740_Q_reg ( .D(g26921), .SI(g10122_Tj), .SE(n10707), .CLK(n11090), 
        .Q(g1404), .QN(n10251) );
  SDFFX1 DFF_742_Q_reg ( .D(g29270), .SI(g1404), .SE(n10700), .CLK(n11083), 
        .Q(g3817), .QN(n10130) );
  SDFFX1 DFF_743_Q_reg ( .D(n10626), .SI(g3817), .SE(n10702), .CLK(n11085), 
        .Q(n9302), .QN(n6010) );
  SDFFX1 DFF_744_Q_reg ( .D(g33038), .SI(n9302), .SE(n10784), .CLK(n11167), 
        .Q(g4501) );
  SDFFX1 DFF_745_Q_reg ( .D(g31865), .SI(g4501), .SE(n10804), .CLK(n11187), 
        .Q(test_so51), .QN(n10668) );
  SDFFX1 DFF_746_Q_reg ( .D(g26926), .SI(test_si52), .SE(n10787), .CLK(n11170), 
        .Q(g2724), .QN(n5301) );
  SDFFX1 DFF_747_Q_reg ( .D(g28083), .SI(g2724), .SE(n10714), .CLK(n11097), 
        .Q(g4704), .QN(n5771) );
  SDFFX1 DFF_749_Q_reg ( .D(g34797), .SI(g22), .SE(n10703), .CLK(n11086), .Q(
        g2878), .QN(n10563) );
  SDFFX1 DFF_750_Q_reg ( .D(g30478), .SI(g2878), .SE(n10714), .CLK(n11097), 
        .Q(g5220) );
  SDFFX1 DFF_751_Q_reg ( .D(g34724), .SI(g5220), .SE(n10750), .CLK(n11133), 
        .Q(g617), .QN(n5339) );
  SDFFX1 DFF_752_Q_reg ( .D(g24212), .SI(g617), .SE(n10750), .CLK(n11133), .Q(
        g12368) );
  SDFFX1 DFF_753_Q_reg ( .D(g26883), .SI(g12368), .SE(n10773), .CLK(n11156), 
        .Q(g316), .QN(n10169) );
  SDFFX1 DFF_754_Q_reg ( .D(g32985), .SI(g316), .SE(n10710), .CLK(n11093), .Q(
        g1277), .QN(n10570) );
  SDFFX1 DFF_755_Q_reg ( .D(g25761), .SI(g1277), .SE(n10726), .CLK(n11109), 
        .Q(g6513), .QN(n5426) );
  SDFFX1 DFF_756_Q_reg ( .D(g26886), .SI(g6513), .SE(n10772), .CLK(n11155), 
        .Q(g336), .QN(n5824) );
  SDFFX1 DFF_757_Q_reg ( .D(g34796), .SI(g336), .SE(n10703), .CLK(n11086), .Q(
        g2882), .QN(n10616) );
  SDFFX1 DFF_758_Q_reg ( .D(g32982), .SI(g2882), .SE(n10804), .CLK(n11187), 
        .Q(test_so52), .QN(n10574) );
  SDFFX1 DFF_759_Q_reg ( .D(g33561), .SI(test_si53), .SE(n10771), .CLK(n11154), 
        .Q(g1906), .QN(n5503) );
  SDFFX1 DFF_760_Q_reg ( .D(g26880), .SI(g1906), .SE(n10771), .CLK(n11154), 
        .Q(g305), .QN(n5282) );
  SDFFX1 DFF_761_Q_reg ( .D(g34975), .SI(g305), .SE(n10701), .CLK(n11084), .Q(
        g8), .QN(n10178) );
  SDFFX1 DFF_763_Q_reg ( .D(g26931), .SI(g8), .SE(n10716), .CLK(n11099), .Q(
        g2799), .QN(n10118) );
  SDFFX1 DFF_764_Q_reg ( .D(g14147), .SI(g2799), .SE(n10753), .CLK(n11136), 
        .Q(g14167), .QN(n10113) );
  SDFFX1 DFF_765_Q_reg ( .D(g13039), .SI(g14167), .SE(n10786), .CLK(n11169), 
        .Q(g17787) );
  SDFFX1 DFF_766_Q_reg ( .D(g34641), .SI(g17787), .SE(n10733), .CLK(n11116), 
        .Q(g4912), .QN(n5297) );
  SDFFX1 DFF_767_Q_reg ( .D(g34629), .SI(g4912), .SE(n10740), .CLK(n11123), 
        .Q(g4157), .QN(n5983) );
  SDFFX1 DFF_768_Q_reg ( .D(g33598), .SI(g4157), .SE(n10717), .CLK(n11100), 
        .Q(g2541), .QN(n5461) );
  SDFFX1 DFF_769_Q_reg ( .D(g33576), .SI(g2541), .SE(n10773), .CLK(n11156), 
        .Q(g2153), .QN(n5356) );
  SDFFX1 DFF_770_Q_reg ( .D(g34720), .SI(g2153), .SE(n10746), .CLK(n11129), 
        .Q(g550), .QN(n10571) );
  SDFFX1 DFF_771_Q_reg ( .D(g26902), .SI(g550), .SE(n10801), .CLK(n11184), .Q(
        g255), .QN(n10275) );
  SDFFX1 DFF_772_Q_reg ( .D(g29244), .SI(g255), .SE(n10801), .CLK(n11184), .Q(
        test_so53), .QN(n10669) );
  SDFFX1 DFF_773_Q_reg ( .D(g30468), .SI(test_si54), .SE(n10779), .CLK(n11162), 
        .Q(g5240), .QN(n10432) );
  SDFFX1 DFF_774_Q_reg ( .D(g26924), .SI(g5240), .SE(n10754), .CLK(n11137), 
        .Q(g1478), .QN(n5289) );
  SDFFX1 DFF_776_Q_reg ( .D(g33031), .SI(g1478), .SE(n10776), .CLK(n11159), 
        .Q(g3863), .QN(n10591) );
  SDFFX1 DFF_777_Q_reg ( .D(n450), .SI(g3863), .SE(n10801), .CLK(n11184), .Q(
        g1959), .QN(n10322) );
  SDFFX1 DFF_778_Q_reg ( .D(g29266), .SI(g1959), .SE(n10720), .CLK(n11103), 
        .Q(g3480), .QN(n5868) );
  SDFFX1 DFF_779_Q_reg ( .D(g30559), .SI(g3480), .SE(n10803), .CLK(n11186), 
        .Q(g6653) );
  SDFFX1 DFF_780_Q_reg ( .D(g14749), .SI(g6653), .SE(n10804), .CLK(n11187), 
        .Q(g17764) );
  SDFFX1 DFF_781_Q_reg ( .D(g34794), .SI(g17764), .SE(n10701), .CLK(n11084), 
        .Q(g2864) );
  SDFFX1 DFF_782_Q_reg ( .D(g28087), .SI(g2864), .SE(n10730), .CLK(n11113), 
        .Q(g4894), .QN(n5774) );
  SDFFX1 DFF_783_Q_reg ( .D(g14635), .SI(g4894), .SE(n10774), .CLK(n11157), 
        .Q(g17678) );
  SDFFX1 DFF_784_Q_reg ( .D(g30435), .SI(g17678), .SE(n10774), .CLK(n11157), 
        .Q(g3857), .QN(n5572) );
  SDFFX1 DFF_785_Q_reg ( .D(g16659), .SI(g3857), .SE(n10774), .CLK(n11157), 
        .Q(g16693), .QN(n10477) );
  SDFFX1 DFF_786_Q_reg ( .D(g25609), .SI(g16693), .SE(n10785), .CLK(n11168), 
        .Q(test_so54), .QN(n10649) );
  SDFFX1 DFF_788_Q_reg ( .D(g28057), .SI(test_si55), .SE(n10796), .CLK(n11179), 
        .Q(g1002), .QN(n10250) );
  SDFFX1 DFF_789_Q_reg ( .D(g34439), .SI(g1002), .SE(n10766), .CLK(n11149), 
        .Q(g776), .QN(n5330) );
  SDFFX1 DFF_790_Q_reg ( .D(g34979), .SI(g776), .SE(n10766), .CLK(n11149), .Q(
        g28), .QN(n5324) );
  SDFFX1 DFF_791_Q_reg ( .D(g10500), .SI(g28), .SE(n10766), .CLK(n11149), .Q(
        g1236), .QN(n10224) );
  SDFFX1 DFF_792_Q_reg ( .D(g34260), .SI(g1236), .SE(n10796), .CLK(n11179), 
        .Q(g4646), .QN(n5712) );
  SDFFX1 DFF_793_Q_reg ( .D(g33012), .SI(g4646), .SE(n10738), .CLK(n11121), 
        .Q(g2476), .QN(n10530) );
  SDFFX1 DFF_794_Q_reg ( .D(g32989), .SI(g2476), .SE(n10724), .CLK(n11107), 
        .Q(g1657), .QN(n5525) );
  SDFFX1 DFF_795_Q_reg ( .D(g34006), .SI(g1657), .SE(n10707), .CLK(n11090), 
        .Q(g2375), .QN(n10198) );
  SDFFX1 DFF_796_Q_reg ( .D(g34783), .SI(g2375), .SE(n10759), .CLK(n11142), 
        .Q(g63), .QN(n10237) );
  SDFFX1 DFF_797_Q_reg ( .D(g14738), .SI(g63), .SE(n10759), .CLK(n11142), .Q(
        g17739), .QN(n10376) );
  SDFFX1 DFF_798_Q_reg ( .D(g8719), .SI(g17739), .SE(n10784), .CLK(n11167), 
        .Q(g358), .QN(n10279) );
  SDFFX1 DFF_799_Q_reg ( .D(g26910), .SI(g358), .SE(n10785), .CLK(n11168), .Q(
        g896), .QN(n5431) );
  SDFFX1 DFF_802_Q_reg ( .D(n92), .SI(g896), .SE(n10804), .CLK(n11187), .Q(
        test_so55), .QN(n10655) );
  SDFFX1 DFF_803_Q_reg ( .D(g33021), .SI(test_si56), .SE(n10789), .CLK(n11172), 
        .Q(g3161), .QN(n10578) );
  SDFFX1 DFF_804_Q_reg ( .D(n609), .SI(g3161), .SE(n10729), .CLK(n11112), .Q(
        g2384), .QN(n10318) );
  SDFFX1 DFF_806_Q_reg ( .D(test_so80), .SI(g2384), .SE(n10729), .CLK(n11112), 
        .Q(g14828), .QN(n5700) );
  SDFFX1 DFF_807_Q_reg ( .D(g34456), .SI(g14828), .SE(n10798), .CLK(n11181), 
        .Q(g4616), .QN(n5608) );
  SDFFX1 DFF_808_Q_reg ( .D(g26968), .SI(g4616), .SE(n10798), .CLK(n11181), 
        .Q(g4561) );
  SDFFX1 DFF_809_Q_reg ( .D(g33991), .SI(g4561), .SE(n10744), .CLK(n11127), 
        .Q(g2024), .QN(n5801) );
  SDFFX1 DFF_810_Q_reg ( .D(g8279), .SI(g2024), .SE(n10800), .CLK(n11183), .Q(
        g3451) );
  SDFFX1 DFF_811_Q_reg ( .D(g26930), .SI(g3451), .SE(n10724), .CLK(n11107), 
        .Q(g2795), .QN(n10119) );
  SDFFX1 DFF_812_Q_reg ( .D(g34599), .SI(g2795), .SE(n10750), .CLK(n11133), 
        .Q(g613), .QN(n5474) );
  SDFFX1 DFF_813_Q_reg ( .D(g28082), .SI(g613), .SE(n10719), .CLK(n11102), .Q(
        g4527), .QN(n10550) );
  SDFFX1 DFF_814_Q_reg ( .D(g33557), .SI(g4527), .SE(n10741), .CLK(n11124), 
        .Q(g1844), .QN(n5847) );
  SDFFX1 DFF_815_Q_reg ( .D(g30511), .SI(g1844), .SE(n10741), .CLK(n11124), 
        .Q(g5937), .QN(n10377) );
  SDFFX1 DFF_816_Q_reg ( .D(g33045), .SI(g5937), .SE(n10782), .CLK(n11165), 
        .Q(test_so56) );
  SDFFX1 DFF_818_Q_reg ( .D(g30379), .SI(test_si57), .SE(n10717), .CLK(n11100), 
        .Q(g2523), .QN(n5281) );
  SDFFX1 DFF_819_Q_reg ( .D(g24267), .SI(g2523), .SE(n10722), .CLK(n11105), 
        .Q(g11349), .QN(n5436) );
  SDFFX1 DFF_820_Q_reg ( .D(g34020), .SI(g11349), .SE(n10716), .CLK(n11099), 
        .Q(g2643), .QN(n10197) );
  SDFFX1 DFF_822_Q_reg ( .D(g24249), .SI(g2643), .SE(n10754), .CLK(n11137), 
        .Q(g1489), .QN(n5850) );
  SDFFX1 DFF_824_Q_reg ( .D(g25592), .SI(g1489), .SE(n10775), .CLK(n11158), 
        .Q(g8358), .QN(n10256) );
  SDFFX1 DFF_825_Q_reg ( .D(g30382), .SI(g8358), .SE(n10717), .CLK(n11100), 
        .Q(n9295), .QN(n19401) );
  SDFFX1 DFF_826_Q_reg ( .D(g29285), .SI(n9295), .SE(n10717), .CLK(n11100), 
        .Q(g5156) );
  SDFFX1 DFF_828_Q_reg ( .D(g12919), .SI(g5156), .SE(n10751), .CLK(n11134), 
        .Q(g30332), .QN(n5526) );
  SDFFX1 DFF_829_Q_reg ( .D(g34975), .SI(g30332), .SE(n10751), .CLK(n11134), 
        .Q(n9294) );
  SDFFX1 DFF_830_Q_reg ( .D(g25662), .SI(n9294), .SE(n10800), .CLK(n11183), 
        .Q(g8279), .QN(n5717) );
  SDFFX1 DFF_831_Q_reg ( .D(g21896), .SI(g8279), .SE(n10755), .CLK(n11138), 
        .Q(g8839) );
  SDFFX1 DFF_832_Q_reg ( .D(g33563), .SI(g8839), .SE(n10758), .CLK(n11141), 
        .Q(g1955), .QN(n10159) );
  SDFFX1 DFF_833_Q_reg ( .D(g33622), .SI(g1955), .SE(n10767), .CLK(n11150), 
        .Q(test_so57), .QN(n10639) );
  SDFFX1 DFF_835_Q_reg ( .D(g33582), .SI(test_si58), .SE(n10734), .CLK(n11117), 
        .Q(g2273), .QN(n5458) );
  SDFFX1 DFF_836_Q_reg ( .D(g17871), .SI(g2273), .SE(n10800), .CLK(n11183), 
        .Q(g14749), .QN(n5584) );
  SDFFX1 DFF_837_Q_reg ( .D(g28086), .SI(g14749), .SE(n10748), .CLK(n11131), 
        .Q(g4771), .QN(n5769) );
  SDFFX1 DFF_838_Q_reg ( .D(g25744), .SI(g4771), .SE(n10748), .CLK(n11131), 
        .Q(g6098) );
  SDFFX1 DFF_839_Q_reg ( .D(g29262), .SI(g6098), .SE(n10789), .CLK(n11172), 
        .Q(g3147) );
  SDFFX1 DFF_840_Q_reg ( .D(g24270), .SI(g3147), .SE(n10722), .CLK(n11105), 
        .Q(g3347), .QN(n10387) );
  SDFFX1 DFF_841_Q_reg ( .D(g33581), .SI(g3347), .SE(n10734), .CLK(n11117), 
        .Q(g2269), .QN(n5410) );
  SDFFX1 DFF_842_Q_reg ( .D(g8358), .SI(g2269), .SE(n10775), .CLK(n11158), .Q(
        g191), .QN(n10257) );
  SDFFX1 DFF_843_Q_reg ( .D(g24266), .SI(g191), .SE(n10775), .CLK(n11158), .Q(
        g2712), .QN(n10142) );
  SDFFX1 DFF_844_Q_reg ( .D(g34849), .SI(g2712), .SE(n10750), .CLK(n11133), 
        .Q(g626), .QN(n5288) );
  SDFFX1 DFF_846_Q_reg ( .D(g33618), .SI(g2729), .SE(n10714), .CLK(n11097), 
        .Q(g5357), .QN(n5393) );
  SDFFX1 DFF_847_Q_reg ( .D(g34038), .SI(g5357), .SE(n10759), .CLK(n11142), 
        .Q(test_so58), .QN(n10652) );
  SDFFX1 DFF_848_Q_reg ( .D(g13068), .SI(test_si59), .SE(n10725), .CLK(n11108), 
        .Q(g17819) );
  SDFFX1 DFF_849_Q_reg ( .D(g34032), .SI(g17819), .SE(n10748), .CLK(n11131), 
        .Q(g4709), .QN(n5518) );
  SDFFX1 DFF_852_Q_reg ( .D(g34803), .SI(g4709), .SE(n10748), .CLK(n11131), 
        .Q(g2927), .QN(n10609) );
  SDFFX1 DFF_853_Q_reg ( .D(g34459), .SI(g2927), .SE(n10746), .CLK(n11129), 
        .Q(g4340), .QN(n5653) );
  SDFFX1 DFF_854_Q_reg ( .D(g30509), .SI(g4340), .SE(n10742), .CLK(n11125), 
        .Q(g5929), .QN(n10341) );
  SDFFX1 DFF_855_Q_reg ( .D(g34640), .SI(g5929), .SE(n10733), .CLK(n11116), 
        .Q(g4907), .QN(n5295) );
  SDFFX1 DFF_856_Q_reg ( .D(g14421), .SI(g4907), .SE(n10733), .CLK(n11116), 
        .Q(g16874) );
  SDFFX1 DFF_857_Q_reg ( .D(g28069), .SI(g16874), .SE(n10800), .CLK(n11183), 
        .Q(g4035), .QN(n10176) );
  SDFFX1 DFF_858_Q_reg ( .D(g21899), .SI(g4035), .SE(n10801), .CLK(n11184), 
        .Q(g2946), .QN(n10565) );
  SDFFX1 DFF_859_Q_reg ( .D(g31868), .SI(g2946), .SE(n10731), .CLK(n11114), 
        .Q(g918), .QN(n5673) );
  SDFFX1 DFF_860_Q_reg ( .D(g26938), .SI(g918), .SE(n10739), .CLK(n11122), .Q(
        g4082), .QN(n10238) );
  SDFFX1 DFF_861_Q_reg ( .D(g25756), .SI(g4082), .SE(n10781), .CLK(n11164), 
        .Q(g9743), .QN(n5719) );
  SDFFX1 DFF_862_Q_reg ( .D(g30363), .SI(g9743), .SE(n10744), .CLK(n11127), 
        .Q(test_so59), .QN(n10680) );
  SDFFX1 DFF_863_Q_reg ( .D(g30334), .SI(test_si60), .SE(n10749), .CLK(n11132), 
        .Q(g577), .QN(n5294) );
  SDFFX1 DFF_864_Q_reg ( .D(g33970), .SI(g577), .SE(n10803), .CLK(n11186), .Q(
        g1620), .QN(n5791) );
  SDFFX1 DFF_865_Q_reg ( .D(g30391), .SI(g1620), .SE(n10708), .CLK(n11091), 
        .Q(g2831), .QN(g30331) );
  SDFFX1 DFF_866_Q_reg ( .D(g25615), .SI(g2831), .SE(n10709), .CLK(n11092), 
        .Q(g667) );
  SDFFX1 DFF_867_Q_reg ( .D(g33540), .SI(g667), .SE(n10731), .CLK(n11114), .Q(
        g930), .QN(n5731) );
  SDFFX1 DFF_868_Q_reg ( .D(g30445), .SI(g930), .SE(n10731), .CLK(n11114), .Q(
        g3937), .QN(n10380) );
  SDFFX1 DFF_870_Q_reg ( .D(g25617), .SI(g3937), .SE(n10745), .CLK(n11128), 
        .Q(g817), .QN(n5822) );
  SDFFX1 DFF_871_Q_reg ( .D(g24247), .SI(g817), .SE(n10747), .CLK(n11130), .Q(
        g1249) );
  SDFFX1 DFF_872_Q_reg ( .D(g24215), .SI(g1249), .SE(n10745), .CLK(n11128), 
        .Q(g837), .QN(n5562) );
  SDFFX1 DFF_873_Q_reg ( .D(g14451), .SI(g837), .SE(n10789), .CLK(n11172), .Q(
        g16924) );
  SDFFX1 DFF_874_Q_reg ( .D(g33964), .SI(g16924), .SE(n10750), .CLK(n11133), 
        .Q(g599), .QN(n5550) );
  SDFFX1 DFF_875_Q_reg ( .D(g25719), .SI(g599), .SE(n10701), .CLK(n11084), .Q(
        g5475), .QN(n5425) );
  SDFFX1 DFF_876_Q_reg ( .D(g29228), .SI(g5475), .SE(n10788), .CLK(n11171), 
        .Q(test_so60) );
  SDFFX1 DFF_877_Q_reg ( .D(g30514), .SI(test_si61), .SE(n10752), .CLK(n11135), 
        .Q(g5949), .QN(n10307) );
  SDFFX1 DFF_878_Q_reg ( .D(g33627), .SI(g5949), .SE(n10730), .CLK(n11113), 
        .Q(g6682) );
  SDFFX1 DFF_880_Q_reg ( .D(g24231), .SI(g6682), .SE(n10730), .CLK(n11113), 
        .Q(g904), .QN(n10240) );
  SDFFX1 DFF_881_Q_reg ( .D(g34615), .SI(g904), .SE(n10743), .CLK(n11126), .Q(
        g2873), .QN(n5488) );
  SDFFX1 DFF_882_Q_reg ( .D(g30356), .SI(g2873), .SE(n10803), .CLK(n11186), 
        .Q(g1854), .QN(n5785) );
  SDFFX1 DFF_883_Q_reg ( .D(g25696), .SI(g1854), .SE(n10699), .CLK(n11082), 
        .Q(g5084), .QN(n5681) );
  SDFFX1 DFF_884_Q_reg ( .D(g30493), .SI(g5084), .SE(n10705), .CLK(n11088), 
        .Q(g5603), .QN(n10289) );
  SDFFX1 DFF_885_Q_reg ( .D(g8917), .SI(g5603), .SE(n10715), .CLK(n11098), .Q(
        g8870), .QN(n5726) );
  SDFFX1 DFF_886_Q_reg ( .D(g33594), .SI(g8870), .SE(n10802), .CLK(n11185), 
        .Q(g2495), .QN(n5522) );
  SDFFX1 DFF_887_Q_reg ( .D(g34009), .SI(g2495), .SE(n10802), .CLK(n11185), 
        .Q(g2437), .QN(n5789) );
  SDFFX1 DFF_888_Q_reg ( .D(g30365), .SI(g2437), .SE(n10725), .CLK(n11108), 
        .Q(g2102), .QN(n5666) );
  SDFFX1 DFF_889_Q_reg ( .D(g33004), .SI(g2102), .SE(n10793), .CLK(n11176), 
        .Q(g2208), .QN(n10532) );
  SDFFX1 DFF_890_Q_reg ( .D(g34018), .SI(g2208), .SE(n10728), .CLK(n11111), 
        .Q(test_so61), .QN(n10663) );
  SDFFX1 DFF_891_Q_reg ( .D(g25685), .SI(test_si62), .SE(n10739), .CLK(n11122), 
        .Q(g4064), .QN(n5416) );
  SDFFX1 DFF_892_Q_reg ( .D(g34040), .SI(g4064), .SE(n10760), .CLK(n11143), 
        .Q(g4899), .QN(n5517) );
  SDFFX1 DFF_893_Q_reg ( .D(g25639), .SI(g4899), .SE(n10760), .CLK(n11143), 
        .Q(g2719), .QN(n5465) );
  SDFFX1 DFF_894_Q_reg ( .D(g34029), .SI(g2719), .SE(n10748), .CLK(n11131), 
        .Q(g4785), .QN(n5361) );
  SDFFX1 DFF_895_Q_reg ( .D(g30488), .SI(g4785), .SE(n10720), .CLK(n11103), 
        .Q(g5583), .QN(n10344) );
  SDFFX1 DFF_896_Q_reg ( .D(g34600), .SI(g5583), .SE(n10766), .CLK(n11149), 
        .Q(g781), .QN(n5551) );
  SDFFX1 DFF_897_Q_reg ( .D(g29300), .SI(g781), .SE(n10705), .CLK(n11088), .Q(
        g6173), .QN(n5810) );
  SDFFX1 DFF_898_Q_reg ( .D(g14705), .SI(g6173), .SE(n10787), .CLK(n11170), 
        .Q(g17743) );
  SDFFX1 DFF_899_Q_reg ( .D(g34802), .SI(g17743), .SE(n10712), .CLK(n11095), 
        .Q(g2917), .QN(n10617) );
  SDFFX1 DFF_900_Q_reg ( .D(g25614), .SI(g2917), .SE(n10709), .CLK(n11092), 
        .Q(g686), .QN(n10141) );
  SDFFX1 DFF_901_Q_reg ( .D(g28058), .SI(g686), .SE(n10709), .CLK(n11092), .Q(
        g1252), .QN(n5554) );
  SDFFX1 DFF_902_Q_reg ( .D(g29225), .SI(g1252), .SE(n10709), .CLK(n11092), 
        .Q(g671), .QN(n10138) );
  SDFFX1 DFF_903_Q_reg ( .D(g33580), .SI(g671), .SE(n10734), .CLK(n11117), .Q(
        test_so62), .QN(n10677) );
  SDFFX1 DFF_904_Q_reg ( .D(g30532), .SI(test_si63), .SE(n10761), .CLK(n11144), 
        .Q(g6283), .QN(n10386) );
  SDFFX1 DFF_905_Q_reg ( .D(g17845), .SI(g6283), .SE(n10783), .CLK(n11166), 
        .Q(g14705), .QN(n5586) );
  SDFFX1 DFF_906_Q_reg ( .D(g17674), .SI(g14705), .SE(n10783), .CLK(n11166), 
        .Q(g17519), .QN(n10359) );
  SDFFX1 DFF_909_Q_reg ( .D(g8783), .SI(g17519), .SE(n10783), .CLK(n11166), 
        .Q(g8784), .QN(DFF_909_n1) );
  SDFFX1 DFF_910_Q_reg ( .D(g33054), .SI(g8784), .SE(n10783), .CLK(n11166), 
        .Q(g5527), .QN(n5389) );
  SDFFX1 DFF_911_Q_reg ( .D(g26962), .SI(g5527), .SE(n10753), .CLK(n11136), 
        .Q(g4489), .QN(n10540) );
  SDFFX1 DFF_912_Q_reg ( .D(n136), .SI(g4489), .SE(n10753), .CLK(n11136), .Q(
        g1974), .QN(n5450) );
  SDFFX1 DFF_913_Q_reg ( .D(g32984), .SI(g1974), .SE(n10710), .CLK(n11093), 
        .Q(g1270), .QN(n5716) );
  SDFFX1 DFF_914_Q_reg ( .D(g34039), .SI(g1270), .SE(n10760), .CLK(n11143), 
        .Q(g4966), .QN(n5706) );
  SDFFX1 DFF_916_Q_reg ( .D(g33065), .SI(g4966), .SE(n10778), .CLK(n11161), 
        .Q(g6227), .QN(n5568) );
  SDFFX1 DFF_917_Q_reg ( .D(g30443), .SI(g6227), .SE(n10732), .CLK(n11115), 
        .Q(g3929), .QN(n10347) );
  SDFFX1 DFF_918_Q_reg ( .D(g29291), .SI(g3929), .SE(n10732), .CLK(n11115), 
        .Q(g5503) );
  SDFFX1 DFF_919_Q_reg ( .D(g24279), .SI(g5503), .SE(n10716), .CLK(n11099), 
        .Q(test_so63), .QN(n10567) );
  SDFFX1 DFF_920_Q_reg ( .D(g30508), .SI(test_si64), .SE(n10741), .CLK(n11124), 
        .Q(g5925), .QN(n10414) );
  SDFFX1 DFF_921_Q_reg ( .D(g29232), .SI(g5925), .SE(n10757), .CLK(n11140), 
        .Q(g1124), .QN(n5692) );
  SDFFX1 DFF_922_Q_reg ( .D(g34269), .SI(g1124), .SE(n10702), .CLK(n11085), 
        .Q(g4955), .QN(n5614) );
  SDFFX1 DFF_923_Q_reg ( .D(g30464), .SI(g4955), .SE(n10779), .CLK(n11162), 
        .Q(g5224), .QN(n10305) );
  SDFFX1 DFF_924_Q_reg ( .D(g33988), .SI(g5224), .SE(n10744), .CLK(n11127), 
        .Q(g2012), .QN(n5790) );
  SDFFX1 DFF_925_Q_reg ( .D(g30522), .SI(g2012), .SE(n10777), .CLK(n11160), 
        .Q(g6203), .QN(n5574) );
  SDFFX1 DFF_926_Q_reg ( .D(g25708), .SI(g6203), .SE(n10718), .CLK(n11101), 
        .Q(g5120) );
  SDFFX1 DFF_927_Q_reg ( .D(g14662), .SI(g5120), .SE(n10718), .CLK(n11101), 
        .Q(g17674), .QN(n10374) );
  SDFFX1 DFF_928_Q_reg ( .D(g30374), .SI(g17674), .SE(n10708), .CLK(n11091), 
        .Q(g2389), .QN(n5631) );
  SDFFX1 DFF_929_Q_reg ( .D(g26953), .SI(g2389), .SE(n10726), .CLK(n11109), 
        .Q(g4438), .QN(n10538) );
  SDFFX1 DFF_930_Q_reg ( .D(g34008), .SI(g4438), .SE(n10802), .CLK(n11185), 
        .Q(g2429), .QN(n5814) );
  SDFFX1 DFF_931_Q_reg ( .D(g34444), .SI(g2429), .SE(n10724), .CLK(n11107), 
        .Q(g2787), .QN(n5610) );
  SDFFX1 DFF_932_Q_reg ( .D(g34731), .SI(g2787), .SE(n10805), .CLK(n11188), 
        .Q(test_so64) );
  SDFFX1 DFF_933_Q_reg ( .D(g33606), .SI(test_si65), .SE(n10706), .CLK(n11089), 
        .Q(g2675), .QN(n5457) );
  SDFFX1 DFF_934_Q_reg ( .D(g24334), .SI(g2675), .SE(n10758), .CLK(n11141), 
        .Q(g18881), .QN(n5541) );
  SDFFX1 DFF_935_Q_reg ( .D(g34265), .SI(g18881), .SE(n10759), .CLK(n11142), 
        .Q(g4836), .QN(n5713) );
  SDFFX1 DFF_936_Q_reg ( .D(g30340), .SI(g4836), .SE(n10745), .CLK(n11128), 
        .Q(g1199), .QN(n10583) );
  SDFFX1 DFF_937_Q_reg ( .D(g24257), .SI(g1199), .SE(n10707), .CLK(n11090), 
        .Q(g19357) );
  SDFFX1 DFF_938_Q_reg ( .D(g30482), .SI(g19357), .SE(n10705), .CLK(n11088), 
        .Q(g5547), .QN(n10291) );
  SDFFX1 DFF_941_Q_reg ( .D(g34604), .SI(g5547), .SE(n10749), .CLK(n11132), 
        .Q(g2138), .QN(n5275) );
  SDFFX1 DFF_942_Q_reg ( .D(g13926), .SI(g2138), .SE(n10791), .CLK(n11174), 
        .Q(g16744), .QN(n10383) );
  SDFFX1 DFF_943_Q_reg ( .D(g33591), .SI(g16744), .SE(n10791), .CLK(n11174), 
        .Q(g2338), .QN(n5310) );
  SDFFX1 DFF_944_Q_reg ( .D(g8918), .SI(g2338), .SE(n10791), .CLK(n11174), .Q(
        g8919) );
  SDFFX1 DFF_945_Q_reg ( .D(g30525), .SI(g8919), .SE(n10761), .CLK(n11144), 
        .Q(g6247), .QN(n10520) );
  SDFFX1 DFF_946_Q_reg ( .D(g26929), .SI(g6247), .SE(n10724), .CLK(n11107), 
        .Q(g2791), .QN(n10120) );
  SDFFX1 DFF_947_Q_reg ( .D(g30448), .SI(g2791), .SE(n10795), .CLK(n11178), 
        .Q(test_so65) );
  SDFFX1 DFF_948_Q_reg ( .D(g34602), .SI(test_si66), .SE(n10699), .CLK(n11082), 
        .Q(g1291), .QN(n2549) );
  SDFFX1 DFF_949_Q_reg ( .D(g30513), .SI(g1291), .SE(n10742), .CLK(n11125), 
        .Q(g5945), .QN(n10340) );
  SDFFX1 DFF_950_Q_reg ( .D(g30469), .SI(g5945), .SE(n10765), .CLK(n11148), 
        .Q(g5244), .QN(n10375) );
  SDFFX1 DFF_951_Q_reg ( .D(g33608), .SI(g5244), .SE(n10765), .CLK(n11148), 
        .Q(g2759), .QN(n10096) );
  SDFFX1 DFF_952_Q_reg ( .D(g33626), .SI(g2759), .SE(n10790), .CLK(n11173), 
        .Q(g6741), .QN(n5398) );
  SDFFX1 DFF_953_Q_reg ( .D(g34725), .SI(g6741), .SE(n10766), .CLK(n11149), 
        .Q(g785), .QN(n5293) );
  SDFFX1 DFF_954_Q_reg ( .D(g30342), .SI(g785), .SE(n10709), .CLK(n11092), .Q(
        g1259), .QN(n5553) );
  SDFFX1 DFF_955_Q_reg ( .D(g29267), .SI(g1259), .SE(n10720), .CLK(n11103), 
        .Q(g3484), .QN(n5668) );
  SDFFX1 DFF_956_Q_reg ( .D(g25593), .SI(g3484), .SE(n10795), .CLK(n11178), 
        .Q(g209), .QN(n5595) );
  SDFFX1 DFF_957_Q_reg ( .D(g30548), .SI(g209), .SE(n10795), .CLK(n11178), .Q(
        g6609), .QN(n10294) );
  SDFFX1 DFF_958_Q_reg ( .D(g33052), .SI(g6609), .SE(n10720), .CLK(n11103), 
        .Q(g5517), .QN(n10589) );
  SDFFX1 DFF_959_Q_reg ( .D(g34012), .SI(g5517), .SE(n10738), .CLK(n11121), 
        .Q(g2449), .QN(n5798) );
  SDFFX1 DFF_960_Q_reg ( .D(g34017), .SI(g2449), .SE(n10728), .CLK(n11111), 
        .Q(test_so66) );
  SDFFX1 DFF_961_Q_reg ( .D(g18881), .SI(test_si67), .SE(n10759), .CLK(n11142), 
        .Q(n9281) );
  SDFFX1 DFF_962_Q_reg ( .D(g24263), .SI(n9281), .SE(n10775), .CLK(n11158), 
        .Q(g2715), .QN(n5299) );
  SDFFX1 DFF_963_Q_reg ( .D(g26912), .SI(g2715), .SE(n10730), .CLK(n11113), 
        .Q(g936), .QN(n5557) );
  SDFFX1 DFF_964_Q_reg ( .D(g30364), .SI(g936), .SE(n10725), .CLK(n11108), .Q(
        g2098), .QN(n5280) );
  SDFFX1 DFF_965_Q_reg ( .D(g34254), .SI(g2098), .SE(n10781), .CLK(n11164), 
        .Q(g4462), .QN(n5671) );
  SDFFX1 DFF_966_Q_reg ( .D(g34251), .SI(g4462), .SE(n10750), .CLK(n11133), 
        .Q(g604), .QN(n5473) );
  SDFFX1 DFF_967_Q_reg ( .D(g30560), .SI(g604), .SE(n10795), .CLK(n11178), .Q(
        g6589) );
  SDFFX1 DFF_968_Q_reg ( .D(g33983), .SI(g6589), .SE(n10758), .CLK(n11141), 
        .Q(n9280), .QN(n19415) );
  SDFFX1 DFF_970_Q_reg ( .D(g13085), .SI(n9280), .SE(n10783), .CLK(n11166), 
        .Q(g17845) );
  SDFFX1 DFF_971_Q_reg ( .D(g13099), .SI(g17845), .SE(n10800), .CLK(n11183), 
        .Q(g17871) );
  SDFFX1 DFF_972_Q_reg ( .D(g24204), .SI(g17871), .SE(n10710), .CLK(n11093), 
        .Q(g429) );
  SDFFX1 DFF_973_Q_reg ( .D(g33980), .SI(g429), .SE(n10758), .CLK(n11141), .Q(
        g1870), .QN(n5813) );
  SDFFX1 DFF_974_Q_reg ( .D(g34631), .SI(g1870), .SE(n10755), .CLK(n11138), 
        .Q(test_so67) );
  SDFFX1 DFF_977_Q_reg ( .D(n956), .SI(test_si68), .SE(n10764), .CLK(n11147), 
        .Q(g1825), .QN(n10316) );
  SDFFX1 DFF_979_Q_reg ( .D(g25623), .SI(g1825), .SE(n10764), .CLK(n11147), 
        .Q(g1008), .QN(n5321) );
  SDFFX1 DFF_980_Q_reg ( .D(g26950), .SI(g1008), .SE(n10772), .CLK(n11155), 
        .Q(g4392), .QN(n5710) );
  SDFFX1 DFF_981_Q_reg ( .D(test_so46), .SI(g4392), .SE(n10772), .CLK(n11155), 
        .Q(g8283), .QN(n10219) );
  SDFFX1 DFF_982_Q_reg ( .D(g30431), .SI(g8283), .SE(n10800), .CLK(n11183), 
        .Q(g3546) );
  SDFFX1 DFF_983_Q_reg ( .D(g30467), .SI(g3546), .SE(n10715), .CLK(n11098), 
        .Q(g5236), .QN(n10338) );
  SDFFX1 DFF_984_Q_reg ( .D(g30353), .SI(g5236), .SE(n10763), .CLK(n11146), 
        .Q(g1768), .QN(n5834) );
  SDFFX1 DFF_985_Q_reg ( .D(g34467), .SI(g1768), .SE(n10763), .CLK(n11146), 
        .Q(g4854) );
  SDFFX1 DFF_986_Q_reg ( .D(g30442), .SI(g4854), .SE(n10731), .CLK(n11114), 
        .Q(g3925), .QN(n10420) );
  SDFFX1 DFF_987_Q_reg ( .D(g29305), .SI(g3925), .SE(n10726), .CLK(n11109), 
        .Q(g6509), .QN(n10171) );
  SDFFX1 DFF_988_Q_reg ( .D(g25616), .SI(g6509), .SE(n10801), .CLK(n11184), 
        .Q(g732), .QN(n5732) );
  SDFFX1 DFF_989_Q_reg ( .D(g29252), .SI(g732), .SE(n10728), .CLK(n11111), .Q(
        g2504), .QN(n10581) );
  SDFFX1 DFF_990_Q_reg ( .D(g13272), .SI(g2504), .SE(n10728), .CLK(n11111), 
        .Q(test_so68), .QN(n10650) );
  SDFFX1 DFF_991_Q_reg ( .D(g4519), .SI(test_si69), .SE(n10715), .CLK(n11098), 
        .Q(g4520) );
  SDFFX1 DFF_992_Q_reg ( .D(g8916), .SI(g4520), .SE(n10715), .CLK(n11098), .Q(
        g8917) );
  SDFFX1 DFF_993_Q_reg ( .D(g33003), .SI(g8917), .SE(n10793), .CLK(n11176), 
        .Q(g2185), .QN(n5376) );
  SDFFX1 DFF_994_Q_reg ( .D(g34613), .SI(g2185), .SE(n10743), .CLK(n11126), 
        .Q(g37), .QN(g30327) );
  SDFFX1 DFF_995_Q_reg ( .D(g16748), .SI(g37), .SE(n10743), .CLK(n11126), .Q(
        g4031) );
  SDFFX1 DFF_996_Q_reg ( .D(g33570), .SI(g4031), .SE(n10744), .CLK(n11127), 
        .Q(g2070), .QN(n5535) );
  SDFFX1 DFF_997_Q_reg ( .D(g8132), .SI(g2070), .SE(n10769), .CLK(n11152), .Q(
        g8235), .QN(n10221) );
  SDFFX1 DFF_1000_Q_reg ( .D(g34734), .SI(g8235), .SE(n10739), .CLK(n11122), 
        .Q(g4176), .QN(n5494) );
  SDFFX1 DFF_1001_Q_reg ( .D(g24275), .SI(g4176), .SE(n10727), .CLK(n11110), 
        .Q(g11418), .QN(n5435) );
  SDFFX1 DFF_1002_Q_reg ( .D(g7243), .SI(g11418), .SE(n10773), .CLK(n11156), 
        .Q(g4405), .QN(n10622) );
  SDFFX1 DFF_1003_Q_reg ( .D(g14167), .SI(g4405), .SE(n10773), .CLK(n11156), 
        .Q(g872), .QN(n10111) );
  SDFFX1 DFF_1004_Q_reg ( .D(g29302), .SI(g872), .SE(n10705), .CLK(n11088), 
        .Q(g6181), .QN(n5667) );
  SDFFX1 DFF_1005_Q_reg ( .D(g24349), .SI(g6181), .SE(n10793), .CLK(n11176), 
        .Q(test_so69), .QN(n10642) );
  SDFFX1 DFF_1006_Q_reg ( .D(g34264), .SI(test_si70), .SE(n10704), .CLK(n11087), .Q(g4765), .QN(n5613) );
  SDFFX1 DFF_1007_Q_reg ( .D(g30484), .SI(g4765), .SE(n10792), .CLK(n11175), 
        .Q(g5563), .QN(n10418) );
  SDFFX1 DFF_1008_Q_reg ( .D(g25634), .SI(g5563), .SE(n10792), .CLK(n11175), 
        .Q(g1395), .QN(n10580) );
  SDFFX1 DFF_1009_Q_reg ( .D(g33567), .SI(g1395), .SE(n10770), .CLK(n11153), 
        .Q(g1913), .QN(n5828) );
  SDFFX1 DFF_1010_Q_reg ( .D(g33585), .SI(g1913), .SE(n10791), .CLK(n11174), 
        .Q(g2331), .QN(n5513) );
  SDFFX1 DFF_1011_Q_reg ( .D(g30527), .SI(g2331), .SE(n10791), .CLK(n11174), 
        .Q(g6263), .QN(n10301) );
  SDFFX1 DFF_1012_Q_reg ( .D(g34978), .SI(g6263), .SE(n10700), .CLK(n11083), 
        .Q(n9276) );
  SDFFX1 DFF_1013_Q_reg ( .D(g30447), .SI(n9276), .SE(n10700), .CLK(n11083), 
        .Q(g3945), .QN(n10346) );
  SDFFX1 DFF_1014_Q_reg ( .D(g7540), .SI(g3945), .SE(n10781), .CLK(n11164), 
        .Q(g347), .QN(n5860) );
  SDFFX1 DFF_1016_Q_reg ( .D(g34256), .SI(g347), .SE(n10781), .CLK(n11164), 
        .Q(g4473), .QN(n10207) );
  SDFFX1 DFF_1017_Q_reg ( .D(g25630), .SI(g4473), .SE(n10781), .CLK(n11164), 
        .Q(g1266), .QN(n10242) );
  SDFFX1 DFF_1018_Q_reg ( .D(g29290), .SI(g1266), .SE(n10699), .CLK(n11082), 
        .Q(g5489), .QN(n5660) );
  SDFFX1 DFF_1019_Q_reg ( .D(g29227), .SI(g5489), .SE(n10709), .CLK(n11092), 
        .Q(test_so70) );
  SDFFX1 DFF_1020_Q_reg ( .D(g31872), .SI(test_si71), .SE(n10788), .CLK(n11171), .Q(g2748), .QN(n5516) );
  SDFFX1 DFF_1021_Q_reg ( .D(g29287), .SI(g2748), .SE(n10701), .CLK(n11084), 
        .Q(g5471), .QN(n10139) );
  SDFFX1 DFF_1022_Q_reg ( .D(g31897), .SI(g5471), .SE(n10726), .CLK(n11109), 
        .Q(g4540) );
  SDFFX1 DFF_1023_Q_reg ( .D(g17764), .SI(g4540), .SE(n10726), .CLK(n11109), 
        .Q(g6723) );
  SDFFX1 DFF_1024_Q_reg ( .D(g30562), .SI(g6723), .SE(n10735), .CLK(n11118), 
        .Q(g6605) );
  SDFFX1 DFF_1025_Q_reg ( .D(g34011), .SI(g6605), .SE(n10738), .CLK(n11121), 
        .Q(n9274), .QN(n19416) );
  SDFFX1 DFF_1026_Q_reg ( .D(g33996), .SI(n9274), .SE(n10755), .CLK(n11138), 
        .Q(g2173) );
  SDFFX1 DFF_1027_Q_reg ( .D(g21898), .SI(g2173), .SE(n10755), .CLK(n11138), 
        .Q(g9019) );
  SDFFX1 DFF_1028_Q_reg ( .D(g33014), .SI(g9019), .SE(n10738), .CLK(n11121), 
        .Q(g2491), .QN(n5405) );
  SDFFX1 DFF_1029_Q_reg ( .D(g34465), .SI(g2491), .SE(n10738), .CLK(n11121), 
        .Q(g4849), .QN(n10542) );
  SDFFX1 DFF_1030_Q_reg ( .D(g33995), .SI(g4849), .SE(n10774), .CLK(n11157), 
        .Q(g2169), .QN(n5788) );
  SDFFX1 DFF_1031_Q_reg ( .D(g30372), .SI(g2169), .SE(n10734), .CLK(n11117), 
        .Q(n9273), .QN(n19402) );
  SDFFX1 DFF_1032_Q_reg ( .D(g30545), .SI(n9273), .SE(n10734), .CLK(n11117), 
        .Q(test_so71), .QN(n10687) );
  SDFFX1 DFF_1033_Q_reg ( .D(g30389), .SI(test_si72), .SE(n10708), .CLK(n11091), .Q(g29219), .QN(n10101) );
  SDFFX1 DFF_1034_Q_reg ( .D(g33590), .SI(g29219), .SE(n10708), .CLK(n11091), 
        .Q(g2407), .QN(n5459) );
  SDFFX1 DFF_1035_Q_reg ( .D(g34616), .SI(g2407), .SE(n10743), .CLK(n11126), 
        .Q(g2868) );
  SDFFX1 DFF_1036_Q_reg ( .D(g26927), .SI(g2868), .SE(n10724), .CLK(n11107), 
        .Q(g2767), .QN(n10123) );
  SDFFX1 DFF_1037_Q_reg ( .D(g32992), .SI(g2767), .SE(n10788), .CLK(n11171), 
        .Q(g1783), .QN(n5596) );
  SDFFX1 DFF_1038_Q_reg ( .D(g13895), .SI(g1783), .SE(n10788), .CLK(n11171), 
        .Q(g16718), .QN(n10372) );
  SDFFX1 DFF_1039_Q_reg ( .D(g25631), .SI(g16718), .SE(n10707), .CLK(n11090), 
        .Q(g1312), .QN(n5466) );
  SDFFX1 DFF_1040_Q_reg ( .D(g30477), .SI(g1312), .SE(n10799), .CLK(n11182), 
        .Q(g5212), .QN(n10464) );
  SDFFX1 DFF_1041_Q_reg ( .D(g34632), .SI(g5212), .SE(n10755), .CLK(n11138), 
        .Q(g4245) );
  SDFFX1 DFF_1042_Q_reg ( .D(g28046), .SI(g4245), .SE(n10709), .CLK(n11092), 
        .Q(g645) );
  SDFFX1 DFF_1043_Q_reg ( .D(g9019), .SI(g645), .SE(n10755), .CLK(n11138), .Q(
        g4291), .QN(n10575) );
  SDFFX1 DFF_1044_Q_reg ( .D(g26896), .SI(g4291), .SE(n10755), .CLK(n11138), 
        .Q(g29212), .QN(n5657) );
  SDFFX1 DFF_1045_Q_reg ( .D(g25602), .SI(g29212), .SE(n10755), .CLK(n11138), 
        .Q(test_so72), .QN(n10672) );
  SDFFX1 DFF_1046_Q_reg ( .D(g26916), .SI(test_si73), .SE(n10757), .CLK(n11140), .Q(g1129), .QN(n5329) );
  SDFFX1 DFF_1047_Q_reg ( .D(g33578), .SI(g1129), .SE(n10773), .CLK(n11156), 
        .Q(g2227), .QN(n5538) );
  SDFFX1 DFF_1049_Q_reg ( .D(g8787), .SI(g2227), .SE(n10773), .CLK(n11156), 
        .Q(g8788), .QN(n10263) );
  SDFFX1 DFF_1050_Q_reg ( .D(g33579), .SI(g8788), .SE(n10736), .CLK(n11119), 
        .Q(g2246), .QN(n10165) );
  SDFFX1 DFF_1051_Q_reg ( .D(g30354), .SI(g2246), .SE(n10741), .CLK(n11124), 
        .Q(g1830), .QN(n5413) );
  SDFFX1 DFF_1052_Q_reg ( .D(g30425), .SI(g1830), .SE(n10733), .CLK(n11116), 
        .Q(g3590), .QN(n10484) );
  SDFFX1 DFF_1053_Q_reg ( .D(g24200), .SI(g3590), .SE(n10710), .CLK(n11093), 
        .Q(g392), .QN(n10272) );
  SDFFX1 DFF_1054_Q_reg ( .D(g33544), .SI(g392), .SE(n10801), .CLK(n11184), 
        .Q(g1592), .QN(n5362) );
  SDFFX1 DFF_1055_Q_reg ( .D(g25764), .SI(g1592), .SE(n10756), .CLK(n11139), 
        .Q(g6505) );
  SDFFX1 DFF_1057_Q_reg ( .D(g24246), .SI(g6505), .SE(n10756), .CLK(n11139), 
        .Q(g1221), .QN(n10547) );
  SDFFX1 DFF_1058_Q_reg ( .D(g30507), .SI(g1221), .SE(n10752), .CLK(n11135), 
        .Q(g5921), .QN(n10328) );
  SDFFX1 DFF_1059_Q_reg ( .D(g26889), .SI(g5921), .SE(n10752), .CLK(n11135), 
        .Q(g29216) );
  SDFFX1 DFF_1060_Q_reg ( .D(g30333), .SI(g29216), .SE(n10711), .CLK(n11094), 
        .Q(test_so73) );
  SDFFX1 DFF_1061_Q_reg ( .D(test_so42), .SI(test_si74), .SE(n10795), .CLK(
        n11178), .Q(g218), .QN(n10537) );
  SDFFX1 DFF_1063_Q_reg ( .D(g32998), .SI(g218), .SE(n10760), .CLK(n11143), 
        .Q(g1932), .QN(n5829) );
  SDFFX1 DFF_1064_Q_reg ( .D(g32987), .SI(g1932), .SE(n10792), .CLK(n11175), 
        .Q(g1624), .QN(n5370) );
  SDFFX1 DFF_1065_Q_reg ( .D(g25702), .SI(g1624), .SE(n10768), .CLK(n11151), 
        .Q(g5062), .QN(n10253) );
  SDFFX1 DFF_1066_Q_reg ( .D(g29286), .SI(g5062), .SE(n10701), .CLK(n11084), 
        .Q(g5462), .QN(n5744) );
  SDFFX1 DFF_1067_Q_reg ( .D(g34606), .SI(g5462), .SE(n10701), .CLK(n11084), 
        .Q(g2689), .QN(n5347) );
  SDFFX1 DFF_1068_Q_reg ( .D(g33070), .SI(g2689), .SE(n10780), .CLK(n11163), 
        .Q(g6573), .QN(n5563) );
  SDFFX1 DFF_1069_Q_reg ( .D(g29240), .SI(g6573), .SE(n10723), .CLK(n11106), 
        .Q(g1677), .QN(n10321) );
  SDFFX1 DFF_1070_Q_reg ( .D(g32999), .SI(g1677), .SE(n10744), .CLK(n11127), 
        .Q(g2028), .QN(n5371) );
  SDFFX1 DFF_1071_Q_reg ( .D(g33605), .SI(g2028), .SE(n10706), .CLK(n11089), 
        .Q(g2671), .QN(n5278) );
  SDFFX1 DFF_1072_Q_reg ( .D(g24255), .SI(g2671), .SE(n10747), .CLK(n11130), 
        .Q(g10527) );
  SDFFX1 DFF_1073_Q_reg ( .D(g26945), .SI(g10527), .SE(n10772), .CLK(n11155), 
        .Q(g7243) );
  SDFFX1 DFF_1074_Q_reg ( .D(n35), .SI(g7243), .SE(n10772), .CLK(n11155), .Q(
        test_so74) );
  SDFFX1 DFF_1075_Q_reg ( .D(g33558), .SI(test_si75), .SE(n10802), .CLK(n11185), .Q(g1848), .QN(n5464) );
  SDFFX1 DFF_1078_Q_reg ( .D(g25699), .SI(g1848), .SE(n10699), .CLK(n11082), 
        .Q(g29213), .QN(n5669) );
  SDFFX1 DFF_1079_Q_reg ( .D(g29289), .SI(g29213), .SE(n10699), .CLK(n11082), 
        .Q(g5485) );
  SDFFX1 DFF_1080_Q_reg ( .D(g30388), .SI(g5485), .SE(n10787), .CLK(n11170), 
        .Q(g2741), .QN(n5349) );
  SDFFX1 DFF_1081_Q_reg ( .D(g12184), .SI(g2741), .SE(n10788), .CLK(n11171), 
        .Q(g11678), .QN(n5482) );
  SDFFX1 DFF_1082_Q_reg ( .D(g29254), .SI(g11678), .SE(n10716), .CLK(n11099), 
        .Q(g2638), .QN(n10594) );
  SDFFX1 DFF_1083_Q_reg ( .D(g28074), .SI(g2638), .SE(n10739), .CLK(n11122), 
        .Q(g4122) );
  SDFFX1 DFF_1084_Q_reg ( .D(g34450), .SI(g4122), .SE(n10790), .CLK(n11173), 
        .Q(g4322), .QN(n5506) );
  SDFFX1 DFF_1085_Q_reg ( .D(g30512), .SI(g4322), .SE(n10741), .CLK(n11124), 
        .Q(g5941), .QN(n10465) );
  SDFFX1 DFF_1086_Q_reg ( .D(n290), .SI(g5941), .SE(n10725), .CLK(n11108), .Q(
        g2108), .QN(n5452) );
  SDFFX1 DFF_1087_Q_reg ( .D(g17646), .SI(g2108), .SE(n10725), .CLK(n11108), 
        .Q(g13068), .QN(n10499) );
  SDFFX1 DFF_1088_Q_reg ( .D(g25), .SI(g13068), .SE(n10725), .CLK(n11108), .Q(
        g25) );
  SDFFX1 DFF_1089_Q_reg ( .D(g33551), .SI(g25), .SE(n10722), .CLK(n11105), .Q(
        test_so75), .QN(n10646) );
  SDFFX1 DFF_1090_Q_reg ( .D(g33538), .SI(test_si76), .SE(n10749), .CLK(n11132), .Q(g595), .QN(n5476) );
  SDFFX1 DFF_1091_Q_reg ( .D(g33005), .SI(g595), .SE(n10792), .CLK(n11175), 
        .Q(g2217), .QN(n5512) );
  SDFFX1 DFF_1092_Q_reg ( .D(g24248), .SI(g2217), .SE(n10707), .CLK(n11090), 
        .Q(n9267), .QN(DFF_1092_n1) );
  SDFFX1 DFF_1093_Q_reg ( .D(g33002), .SI(n9267), .SE(n10724), .CLK(n11107), 
        .Q(g2066), .QN(n5832) );
  SDFFX1 DFF_1094_Q_reg ( .D(g24234), .SI(g2066), .SE(n10757), .CLK(n11140), 
        .Q(g1152), .QN(n5618) );
  SDFFX1 DFF_1095_Q_reg ( .D(g30471), .SI(g1152), .SE(n10715), .CLK(n11098), 
        .Q(g5252), .QN(n10337) );
  SDFFX1 DFF_1096_Q_reg ( .D(g34000), .SI(g5252), .SE(n10736), .CLK(n11119), 
        .Q(g2165), .QN(n10158) );
  SDFFX1 DFF_1097_Q_reg ( .D(g34016), .SI(g2165), .SE(n10736), .CLK(n11119), 
        .Q(g2571), .QN(n5787) );
  SDFFX1 DFF_1098_Q_reg ( .D(g33048), .SI(g2571), .SE(n10778), .CLK(n11161), 
        .Q(g5176), .QN(n5650) );
  SDFFX1 DFF_1100_Q_reg ( .D(g8283), .SI(g5176), .SE(n10778), .CLK(n11161), 
        .Q(g8403), .QN(n10220) );
  SDFFX1 DFF_1102_Q_reg ( .D(g17819), .SI(g8403), .SE(n10779), .CLK(n11162), 
        .Q(g14673), .QN(n5581) );
  SDFFX1 DFF_1103_Q_reg ( .D(g25628), .SI(g14673), .SE(n10756), .CLK(n11139), 
        .Q(test_so76), .QN(n10673) );
  SDFFX1 DFF_1104_Q_reg ( .D(g26934), .SI(test_si77), .SE(n10728), .CLK(n11111), .Q(g2827), .QN(n10122) );
  SDFFX1 DFF_1106_Q_reg ( .D(g14201), .SI(g2827), .SE(n10753), .CLK(n11136), 
        .Q(g14217), .QN(n10108) );
  SDFFX1 DFF_1107_Q_reg ( .D(g34468), .SI(g14217), .SE(n10764), .CLK(n11147), 
        .Q(g4859), .QN(n10099) );
  SDFFX1 DFF_1108_Q_reg ( .D(g24202), .SI(g4859), .SE(n10710), .CLK(n11093), 
        .Q(g424), .QN(n10245) );
  SDFFX1 DFF_1109_Q_reg ( .D(g33542), .SI(g424), .SE(n10710), .CLK(n11093), 
        .Q(g1274), .QN(n5730) );
  SDFFX1 DFF_1110_Q_reg ( .D(g17404), .SI(g1274), .SE(n10736), .CLK(n11119), 
        .Q(g17423), .QN(n10234) );
  SDFFX1 DFF_1111_Q_reg ( .D(g33435), .SI(g17423), .SE(n10792), .CLK(n11175), 
        .Q(n9265), .QN(n10690) );
  SDFFX1 DFF_1112_Q_reg ( .D(g34445), .SI(n9265), .SE(n10780), .CLK(n11163), 
        .Q(g2803), .QN(n5545) );
  SDFFX1 DFF_1114_Q_reg ( .D(g33555), .SI(g2803), .SE(n10741), .CLK(n11124), 
        .Q(g1821), .QN(n10160) );
  SDFFX1 DFF_1115_Q_reg ( .D(g34013), .SI(g1821), .SE(n10727), .CLK(n11110), 
        .Q(g2509), .QN(n10196) );
  SDFFX1 DFF_1116_Q_reg ( .D(g28091), .SI(g2509), .SE(n10769), .CLK(n11152), 
        .Q(g5073), .QN(n10194) );
  SDFFX1 DFF_1117_Q_reg ( .D(g26919), .SI(g5073), .SE(n10802), .CLK(n11185), 
        .Q(test_so77), .QN(n5556) );
  SDFFX1 DFF_1118_Q_reg ( .D(g8235), .SI(test_si78), .SE(n10769), .CLK(n11152), 
        .Q(g8353), .QN(n10222) );
  SDFFX1 DFF_1119_Q_reg ( .D(g17685), .SI(g8353), .SE(n10783), .CLK(n11166), 
        .Q(g13085), .QN(n10519) );
  SDFFX1 DFF_1120_Q_reg ( .D(g30554), .SI(g13085), .SE(n10735), .CLK(n11118), 
        .Q(g6633), .QN(n10479) );
  SDFFX1 DFF_1121_Q_reg ( .D(g29281), .SI(g6633), .SE(n10714), .CLK(n11097), 
        .Q(g5124), .QN(n10129) );
  SDFFX1 DFF_1122_Q_reg ( .D(test_so44), .SI(g5124), .SE(n10756), .CLK(n11139), 
        .Q(g17400), .QN(n10227) );
  SDFFX1 DFF_1123_Q_reg ( .D(g30537), .SI(g17400), .SE(n10800), .CLK(n11183), 
        .Q(g6303), .QN(n10491) );
  SDFFX1 DFF_1124_Q_reg ( .D(g28092), .SI(g6303), .SE(n10699), .CLK(n11082), 
        .Q(g5069), .QN(n10193) );
  SDFFX1 DFF_1125_Q_reg ( .D(g34732), .SI(g5069), .SE(n10743), .CLK(n11126), 
        .Q(g2994), .QN(n5634) );
  SDFFX1 DFF_1126_Q_reg ( .D(g28049), .SI(g2994), .SE(n10711), .CLK(n11094), 
        .Q(g650), .QN(n10270) );
  SDFFX1 DFF_1127_Q_reg ( .D(g33545), .SI(g650), .SE(n10722), .CLK(n11105), 
        .Q(g1636), .QN(n5549) );
  SDFFX1 DFF_1128_Q_reg ( .D(g30441), .SI(g1636), .SE(n10796), .CLK(n11179), 
        .Q(g3921), .QN(n10330) );
  SDFFX1 DFF_1129_Q_reg ( .D(g29247), .SI(g3921), .SE(n10725), .CLK(n11108), 
        .Q(test_so78) );
  SDFFX1 DFF_1130_Q_reg ( .D(g24354), .SI(test_si79), .SE(n10730), .CLK(n11113), .Q(g6732), .QN(n10524) );
  SDFFX1 DFF_1131_Q_reg ( .D(g25636), .SI(g6732), .SE(n10762), .CLK(n11145), 
        .Q(g1306), .QN(n5796) );
  SDFFX1 DFF_1133_Q_reg ( .D(g26914), .SI(g1306), .SE(n10797), .CLK(n11180), 
        .Q(g1061), .QN(n10252) );
  SDFFX1 DFF_1134_Q_reg ( .D(g25670), .SI(g1061), .SE(n10797), .CLK(n11180), 
        .Q(g3462) );
  SDFFX1 DFF_1135_Q_reg ( .D(g33998), .SI(g3462), .SE(n10755), .CLK(n11138), 
        .Q(g2181), .QN(n5803) );
  SDFFX1 DFF_1136_Q_reg ( .D(g25626), .SI(g2181), .SE(n10751), .CLK(n11134), 
        .Q(g956), .QN(n5341) );
  SDFFX1 DFF_1137_Q_reg ( .D(g33977), .SI(g956), .SE(n10763), .CLK(n11146), 
        .Q(g1756), .QN(n5804) );
  SDFFX1 DFF_1138_Q_reg ( .D(g29297), .SI(g1756), .SE(n10785), .CLK(n11168), 
        .Q(g5849) );
  SDFFX1 DFF_1139_Q_reg ( .D(g28071), .SI(g5849), .SE(n10786), .CLK(n11169), 
        .Q(g4112), .QN(n10522) );
  SDFFX1 DFF_1140_Q_reg ( .D(g30387), .SI(g4112), .SE(n10706), .CLK(n11089), 
        .Q(n9262), .QN(n19404) );
  SDFFX1 DFF_1141_Q_reg ( .D(g33577), .SI(n9262), .SE(n10706), .CLK(n11089), 
        .Q(g2197), .QN(n5514) );
  SDFFX1 DFF_1143_Q_reg ( .D(g33592), .SI(g2197), .SE(n10802), .CLK(n11185), 
        .Q(test_so79), .QN(n10648) );
  SDFFX1 DFF_1144_Q_reg ( .D(g26913), .SI(test_si80), .SE(n10764), .CLK(n11147), .Q(g1046), .QN(n10619) );
  SDFFX1 DFF_1145_Q_reg ( .D(g28044), .SI(g1046), .SE(n10764), .CLK(n11147), 
        .Q(g482), .QN(n5820) );
  SDFFX1 DFF_1146_Q_reg ( .D(g26948), .SI(g482), .SE(n10773), .CLK(n11156), 
        .Q(g4401) );
  SDFFX1 DFF_1148_Q_reg ( .D(g30344), .SI(g4401), .SE(n10773), .CLK(n11156), 
        .Q(g1514), .QN(n5364) );
  SDFFX1 DFF_1149_Q_reg ( .D(g26885), .SI(g1514), .SE(n10780), .CLK(n11163), 
        .Q(g329), .QN(n5766) );
  SDFFX1 DFF_1150_Q_reg ( .D(g33069), .SI(g329), .SE(n10780), .CLK(n11163), 
        .Q(g6565), .QN(n5386) );
  SDFFX1 DFF_1151_Q_reg ( .D(g34621), .SI(g6565), .SE(n10803), .CLK(n11186), 
        .Q(g2950), .QN(n10560) );
  SDFFX1 DFF_1153_Q_reg ( .D(g28059), .SI(g2950), .SE(n10804), .CLK(n11187), 
        .Q(g1345), .QN(n10249) );
  SDFFX1 DFF_1154_Q_reg ( .D(n1426), .SI(g1345), .SE(n10722), .CLK(n11105), 
        .Q(g6533), .QN(n5445) );
  SDFFX1 DFF_1155_Q_reg ( .D(g16624), .SI(g6533), .SE(n10722), .CLK(n11105), 
        .Q(g14421), .QN(n10495) );
  SDFFX1 DFF_1157_Q_reg ( .D(g34633), .SI(g14421), .SE(n10722), .CLK(n11105), 
        .Q(g4727), .QN(n5312) );
  SDFFX1 DFF_1158_Q_reg ( .D(g24352), .SI(g4727), .SE(n10729), .CLK(n11112), 
        .Q(test_so80) );
  SDFFX1 DFF_1159_Q_reg ( .D(g26925), .SI(test_si81), .SE(n10748), .CLK(n11131), .Q(g1536) );
  SDFFX1 DFF_1160_Q_reg ( .D(g30446), .SI(g1536), .SE(n10731), .CLK(n11114), 
        .Q(g3941), .QN(n10474) );
  SDFFX1 DFF_1161_Q_reg ( .D(g25597), .SI(g3941), .SE(n10785), .CLK(n11168), 
        .Q(g370), .QN(n10610) );
  SDFFX1 DFF_1162_Q_reg ( .D(g24342), .SI(g370), .SE(n10797), .CLK(n11180), 
        .Q(g5694), .QN(n10395) );
  SDFFX1 DFF_1163_Q_reg ( .D(g30357), .SI(g5694), .SE(n10803), .CLK(n11186), 
        .Q(g1858), .QN(n5892) );
  SDFFX1 DFF_1164_Q_reg ( .D(g26908), .SI(g1858), .SE(n10709), .CLK(n11092), 
        .Q(g446) );
  SDFFX1 DFF_1166_Q_reg ( .D(g30399), .SI(g446), .SE(n10791), .CLK(n11174), 
        .Q(g3219), .QN(n10327) );
  SDFFX1 DFF_1167_Q_reg ( .D(g29242), .SI(g3219), .SE(n10708), .CLK(n11091), 
        .Q(g1811), .QN(n10317) );
  SDFFX1 DFF_1169_Q_reg ( .D(g30547), .SI(g1811), .SE(n10735), .CLK(n11118), 
        .Q(g6601), .QN(n10424) );
  SDFFX1 DFF_1171_Q_reg ( .D(g34010), .SI(g6601), .SE(n10738), .CLK(n11121), 
        .Q(g2441) );
  SDFFX1 DFF_1172_Q_reg ( .D(g33986), .SI(g2441), .SE(n10758), .CLK(n11141), 
        .Q(g1874), .QN(n10144) );
  SDFFX1 DFF_1173_Q_reg ( .D(g34257), .SI(g1874), .SE(n10759), .CLK(n11142), 
        .Q(test_so81), .QN(n10643) );
  SDFFX1 DFF_1174_Q_reg ( .D(g30544), .SI(test_si82), .SE(n10780), .CLK(n11163), .Q(g6581), .QN(n10450) );
  SDFFX1 DFF_1175_Q_reg ( .D(g30561), .SI(g6581), .SE(n10734), .CLK(n11117), 
        .Q(g6597), .QN(n10483) );
  SDFFX1 DFF_1176_Q_reg ( .D(g8403), .SI(g6597), .SE(n10778), .CLK(n11161), 
        .Q(g5008), .QN(n5637) );
  SDFFX1 DFF_1177_Q_reg ( .D(g30430), .SI(g5008), .SE(n10779), .CLK(n11162), 
        .Q(g3610) );
  SDFFX1 DFF_1178_Q_reg ( .D(g34799), .SI(g3610), .SE(n10743), .CLK(n11126), 
        .Q(g2890), .QN(n10568) );
  SDFFX1 DFF_1179_Q_reg ( .D(g33565), .SI(g2890), .SE(n10754), .CLK(n11137), 
        .Q(g1978), .QN(n5845) );
  SDFFX1 DFF_1180_Q_reg ( .D(g33968), .SI(g1978), .SE(n10801), .CLK(n11184), 
        .Q(g1612) );
  SDFFX1 DFF_1181_Q_reg ( .D(g34843), .SI(g1612), .SE(n10751), .CLK(n11134), 
        .Q(g112), .QN(n10273) );
  SDFFX1 DFF_1182_Q_reg ( .D(g34793), .SI(g112), .SE(n10701), .CLK(n11084), 
        .Q(g2856), .QN(n10618) );
  SDFFX1 DFF_1184_Q_reg ( .D(g33566), .SI(g2856), .SE(n10754), .CLK(n11137), 
        .Q(g1982), .QN(n5462) );
  SDFFX1 DFF_1185_Q_reg ( .D(g17688), .SI(g1982), .SE(n10765), .CLK(n11148), 
        .Q(g17722), .QN(n10482) );
  SDFFX1 DFF_1186_Q_reg ( .D(g30465), .SI(g17722), .SE(n10765), .CLK(n11148), 
        .Q(test_so82), .QN(n10689) );
  SDFFX1 DFF_1187_Q_reg ( .D(g28073), .SI(test_si83), .SE(n10739), .CLK(n11122), .Q(g4119), .QN(n10114) );
  SDFFX1 DFF_1188_Q_reg ( .D(g24351), .SI(g4119), .SE(n10793), .CLK(n11176), 
        .Q(g6390), .QN(n10389) );
  SDFFX1 DFF_1189_Q_reg ( .D(g30346), .SI(g6390), .SE(n10748), .CLK(n11131), 
        .Q(g1542), .QN(n10584) );
  SDFFX1 DFF_1190_Q_reg ( .D(g21893), .SI(g1542), .SE(n10748), .CLK(n11131), 
        .Q(g4258), .QN(n10127) );
  SDFFX1 DFF_1191_Q_reg ( .D(g8353), .SI(g4258), .SE(n10769), .CLK(n11152), 
        .Q(g4818) );
  SDFFX1 DFF_1192_Q_reg ( .D(g31904), .SI(g4818), .SE(n10768), .CLK(n11151), 
        .Q(g5033), .QN(n10598) );
  SDFFX1 DFF_1193_Q_reg ( .D(g34635), .SI(g5033), .SE(n10768), .CLK(n11151), 
        .Q(g4717), .QN(n5344) );
  SDFFX1 DFF_1194_Q_reg ( .D(g25637), .SI(g4717), .SE(n10747), .CLK(n11130), 
        .Q(g1554), .QN(n5768) );
  SDFFX1 DFF_1195_Q_reg ( .D(g29274), .SI(g1554), .SE(n10764), .CLK(n11147), 
        .Q(g3849) );
  SDFFX1 DFF_1196_Q_reg ( .D(g14828), .SI(g3849), .SE(n10765), .CLK(n11148), 
        .Q(g17778), .QN(n10381) );
  SDFFX1 DFF_1197_Q_reg ( .D(g30396), .SI(g17778), .SE(n10804), .CLK(n11187), 
        .Q(g3199), .QN(n10496) );
  SDFFX1 DFF_1198_Q_reg ( .D(g25735), .SI(g3199), .SE(n10805), .CLK(n11188), 
        .Q(test_so83) );
  SDFFX1 DFF_1199_Q_reg ( .D(g34037), .SI(test_si84), .SE(n10760), .CLK(n11143), .Q(g4975), .QN(n5360) );
  SDFFX1 DFF_1200_Q_reg ( .D(g34791), .SI(g4975), .SE(n10767), .CLK(n11150), 
        .Q(g790), .QN(n5292) );
  SDFFX1 DFF_1201_Q_reg ( .D(g30520), .SI(g790), .SE(n10742), .CLK(n11125), 
        .Q(g5913) );
  SDFFX1 DFF_1202_Q_reg ( .D(g30358), .SI(g5913), .SE(n10758), .CLK(n11141), 
        .Q(g1902), .QN(n5837) );
  SDFFX1 DFF_1203_Q_reg ( .D(g29299), .SI(g1902), .SE(n10704), .CLK(n11087), 
        .Q(g6163), .QN(n10153) );
  SDFFX1 DFF_1204_Q_reg ( .D(g25690), .SI(g6163), .SE(n10752), .CLK(n11135), 
        .Q(g4125), .QN(n10521) );
  SDFFX1 DFF_1205_Q_reg ( .D(g28096), .SI(g4125), .SE(n10721), .CLK(n11104), 
        .Q(g4821), .QN(n5880) );
  SDFFX1 DFF_1206_Q_reg ( .D(g28088), .SI(g4821), .SE(n10721), .CLK(n11104), 
        .Q(g4939) );
  SDFFX1 DFF_1207_Q_reg ( .D(g24241), .SI(g4939), .SE(n10796), .CLK(n11179), 
        .Q(g19334), .QN(n5392) );
  SDFFX1 DFF_1208_Q_reg ( .D(g30397), .SI(g19334), .SE(n10718), .CLK(n11101), 
        .Q(g3207), .QN(n10409) );
  SDFFX1 DFF_1209_Q_reg ( .D(g4520), .SI(g3207), .SE(n10718), .CLK(n11101), 
        .Q(g4483), .QN(n10539) );
  SDFFX1 DFF_1210_Q_reg ( .D(g30409), .SI(g4483), .SE(n10719), .CLK(n11102), 
        .Q(test_so84) );
  SDFFX1 DFF_1211_Q_reg ( .D(g29284), .SI(test_si85), .SE(n10714), .CLK(n11097), .Q(g5142), .QN(n5658) );
  SDFFX1 DFF_1212_Q_reg ( .D(g30470), .SI(g5142), .SE(n10714), .CLK(n11097), 
        .Q(g5248), .QN(n10460) );
  SDFFX1 DFF_1213_Q_reg ( .D(g30367), .SI(g5248), .SE(n10701), .CLK(n11084), 
        .Q(g2126), .QN(n5891) );
  SDFFX1 DFF_1214_Q_reg ( .D(g24273), .SI(g2126), .SE(n10802), .CLK(n11185), 
        .Q(g3694), .QN(n10393) );
  SDFFX1 DFF_1215_Q_reg ( .D(n198), .SI(g3694), .SE(n10702), .CLK(n11085), .Q(
        g5481), .QN(n5805) );
  SDFFX1 DFF_1216_Q_reg ( .D(g30359), .SI(g5481), .SE(n10702), .CLK(n11085), 
        .Q(g1964), .QN(n5315) );
  SDFFX1 DFF_1217_Q_reg ( .D(g25698), .SI(g1964), .SE(n10699), .CLK(n11082), 
        .Q(g5097), .QN(n5753) );
  SDFFX1 DFF_1218_Q_reg ( .D(g30398), .SI(g5097), .SE(n10790), .CLK(n11173), 
        .Q(g3215), .QN(n10286) );
  SDFFX1 DFF_1219_Q_reg ( .D(g13906), .SI(g3215), .SE(n10780), .CLK(n11163), 
        .Q(g16748) );
  SDFFX1 DFF_1220_Q_reg ( .D(g33079), .SI(g16748), .SE(n10780), .CLK(n11163), 
        .Q(n9255) );
  SDFFX1 DFF_1221_Q_reg ( .D(g26952), .SI(n9255), .SE(n10746), .CLK(n11129), 
        .Q(g4427), .QN(n10266) );
  SDFFX1 DFF_1222_Q_reg ( .D(g34974), .SI(g4427), .SE(n10746), .CLK(n11129), 
        .Q(test_so85) );
  SDFFX1 DFF_1223_Q_reg ( .D(g26928), .SI(test_si86), .SE(n10724), .CLK(n11107), .Q(g2779), .QN(n10117) );
  SDFFX1 DFF_1224_Q_reg ( .D(test_so39), .SI(g2779), .SE(n10737), .CLK(n11120), 
        .Q(g8786), .QN(n5694) );
  SDFFX1 DFF_1225_Q_reg ( .D(g26954), .SI(g8786), .SE(n10794), .CLK(n11177), 
        .Q(g7245) );
  SDFFX1 DFF_1226_Q_reg ( .D(g30351), .SI(g7245), .SE(n10794), .CLK(n11177), 
        .Q(g1720), .QN(n5780) );
  SDFFX1 DFF_1227_Q_reg ( .D(g31871), .SI(g1720), .SE(n10707), .CLK(n11090), 
        .Q(g1367), .QN(n10229) );
  SDFFX1 DFF_1228_Q_reg ( .D(g9553), .SI(g1367), .SE(n10793), .CLK(n11176), 
        .Q(g5112) );
  SDFFX1 DFF_1229_Q_reg ( .D(g34978), .SI(g5112), .SE(n10794), .CLK(n11177), 
        .Q(g19), .QN(n10097) );
  SDFFX1 DFF_1230_Q_reg ( .D(g26939), .SI(g19), .SE(n10740), .CLK(n11123), .Q(
        g4145), .QN(n10551) );
  SDFFX1 DFF_1231_Q_reg ( .D(g33994), .SI(g4145), .SE(n10706), .CLK(n11089), 
        .Q(g2161), .QN(n5812) );
  SDFFX1 DFF_1232_Q_reg ( .D(g25596), .SI(g2161), .SE(n10785), .CLK(n11168), 
        .Q(g376), .QN(n5633) );
  SDFFX1 DFF_1233_Q_reg ( .D(g33586), .SI(g376), .SE(n10791), .CLK(n11174), 
        .Q(g2361), .QN(n5537) );
  SDFFX1 DFF_1234_Q_reg ( .D(g21901), .SI(g2361), .SE(n10737), .CLK(n11120), 
        .Q(test_so86), .QN(DFF_1234_n1) );
  SDFFX1 DFF_1235_Q_reg ( .D(g31866), .SI(test_si87), .SE(n10749), .CLK(n11132), .Q(g582), .QN(n5552) );
  SDFFX1 DFF_1236_Q_reg ( .D(g33000), .SI(g582), .SE(n10744), .CLK(n11127), 
        .Q(g2051), .QN(n10528) );
  SDFFX1 DFF_1237_Q_reg ( .D(g26918), .SI(g2051), .SE(n10745), .CLK(n11128), 
        .Q(g1193), .QN(n10606) );
  SDFFX1 DFF_1240_Q_reg ( .D(g30373), .SI(g1193), .SE(n10797), .CLK(n11180), 
        .Q(g2327), .QN(n5841) );
  SDFFX1 DFF_1241_Q_reg ( .D(g28056), .SI(g2327), .SE(n10730), .CLK(n11113), 
        .Q(g907), .QN(n5555) );
  SDFFX1 DFF_1242_Q_reg ( .D(g34601), .SI(g907), .SE(n10730), .CLK(n11113), 
        .Q(g947), .QN(n5286) );
  SDFFX1 DFF_1243_Q_reg ( .D(g30355), .SI(g947), .SE(n10741), .CLK(n11124), 
        .Q(g1834), .QN(n5665) );
  SDFFX1 DFF_1244_Q_reg ( .D(g30426), .SI(g1834), .SE(n10777), .CLK(n11160), 
        .Q(g3594), .QN(n10352) );
  SDFFX1 DFF_1245_Q_reg ( .D(g34805), .SI(g3594), .SE(n10743), .CLK(n11126), 
        .Q(g2999), .QN(n10569) );
  SDFFX1 DFF_1247_Q_reg ( .D(g34002), .SI(g2999), .SE(n10768), .CLK(n11151), 
        .Q(g2303), .QN(n5794) );
  SDFFX1 DFF_1248_Q_reg ( .D(g17778), .SI(g2303), .SE(n10765), .CLK(n11148), 
        .Q(g17688), .QN(n10367) );
  SDFFX1 DFF_1250_Q_reg ( .D(g28053), .SI(g17688), .SE(n10710), .CLK(n11093), 
        .Q(test_so87), .QN(n10659) );
  SDFFX1 DFF_1251_Q_reg ( .D(g29229), .SI(test_si88), .SE(n10745), .CLK(n11128), .Q(g723), .QN(n5826) );
  SDFFX1 DFF_1252_Q_reg ( .D(g33620), .SI(g723), .SE(n10745), .CLK(n11128), 
        .Q(g5703), .QN(n5397) );
  SDFFX1 DFF_1253_Q_reg ( .D(g34722), .SI(g5703), .SE(n10745), .CLK(n11128), 
        .Q(g546), .QN(n5492) );
  SDFFX1 DFF_1254_Q_reg ( .D(g33599), .SI(g546), .SE(n10752), .CLK(n11135), 
        .Q(g2472), .QN(n5619) );
  SDFFX1 DFF_1255_Q_reg ( .D(g30515), .SI(g2472), .SE(n10741), .CLK(n11124), 
        .Q(g5953), .QN(n10362) );
  SDFFX1 DFF_1256_Q_reg ( .D(g25649), .SI(g5953), .SE(n10801), .CLK(n11184), 
        .Q(g8277) );
  SDFFX1 DFF_1258_Q_reg ( .D(g33979), .SI(g8277), .SE(n10801), .CLK(n11184), 
        .Q(g1740), .QN(n10208) );
  SDFFX1 DFF_1259_Q_reg ( .D(g30417), .SI(g1740), .SE(n10732), .CLK(n11115), 
        .Q(g3550), .QN(n10516) );
  SDFFX1 DFF_1260_Q_reg ( .D(g25683), .SI(g3550), .SE(n10700), .CLK(n11083), 
        .Q(g3845) );
  SDFFX1 DFF_1261_Q_reg ( .D(g33574), .SI(g3845), .SE(n10700), .CLK(n11083), 
        .Q(g2116), .QN(n5463) );
  SDFFX1 DFF_1262_Q_reg ( .D(g17813), .SI(g2116), .SE(n10774), .CLK(n11157), 
        .Q(g14635), .QN(n5582) );
  SDFFX1 DFF_1263_Q_reg ( .D(g30410), .SI(g14635), .SE(n10790), .CLK(n11173), 
        .Q(test_so88) );
  SDFFX1 DFF_1264_Q_reg ( .D(g30454), .SI(test_si89), .SE(n10731), .CLK(n11114), .Q(g3913), .QN(n10506) );
  SDFFX1 DFF_1265_Q_reg ( .D(g34024), .SI(g3913), .SE(n10726), .CLK(n11109), 
        .Q(g10306) );
  SDFFX1 DFF_1266_Q_reg ( .D(g33547), .SI(g10306), .SE(n10737), .CLK(n11120), 
        .Q(g1687), .QN(n10164) );
  SDFFX1 DFF_1267_Q_reg ( .D(g30386), .SI(g1687), .SE(n10706), .CLK(n11089), 
        .Q(g2681), .QN(n5777) );
  SDFFX1 DFF_1268_Q_reg ( .D(n755), .SI(g2681), .SE(n10717), .CLK(n11100), .Q(
        g2533), .QN(n5761) );
  SDFFX1 DFF_1269_Q_reg ( .D(g26887), .SI(g2533), .SE(n10772), .CLK(n11155), 
        .Q(g324), .QN(n5827) );
  SDFFX1 DFF_1270_Q_reg ( .D(g34607), .SI(g324), .SE(n10772), .CLK(n11155), 
        .Q(g2697), .QN(n5308) );
  SDFFX1 DFF_1272_Q_reg ( .D(g31895), .SI(g2697), .SE(n10772), .CLK(n11155), 
        .Q(g4417) );
  SDFFX1 DFF_1273_Q_reg ( .D(g33068), .SI(g4417), .SE(n10776), .CLK(n11159), 
        .Q(g6561), .QN(n5646) );
  SDFFX1 DFF_1274_Q_reg ( .D(g29233), .SI(g6561), .SE(n10751), .CLK(n11134), 
        .Q(g1141), .QN(n5691) );
  SDFFX1 DFF_1275_Q_reg ( .D(g24258), .SI(g1141), .SE(n10747), .CLK(n11130), 
        .Q(g12923), .QN(n5655) );
  SDFFX1 DFF_1276_Q_reg ( .D(g30376), .SI(g12923), .SE(n10708), .CLK(n11091), 
        .Q(test_so89), .QN(n10681) );
  SDFFX1 DFF_1277_Q_reg ( .D(g33549), .SI(test_si90), .SE(n10723), .CLK(n11106), .Q(g1710), .QN(n5412) );
  SDFFX1 DFF_1278_Q_reg ( .D(g29308), .SI(g1710), .SE(n10721), .CLK(n11104), 
        .Q(g6527), .QN(n5659) );
  SDFFX1 DFF_1280_Q_reg ( .D(g30408), .SI(g6527), .SE(n10718), .CLK(n11101), 
        .Q(g3255), .QN(n10457) );
  SDFFX1 DFF_1281_Q_reg ( .D(n15), .SI(g3255), .SE(n10723), .CLK(n11106), .Q(
        g1691), .QN(n10320) );
  SDFFX1 DFF_1282_Q_reg ( .D(g34620), .SI(g1691), .SE(n10803), .CLK(n11186), 
        .Q(g2936), .QN(n10561) );
  SDFFX1 DFF_1283_Q_reg ( .D(g33621), .SI(g2936), .SE(n10713), .CLK(n11096), 
        .Q(g5644), .QN(n5593) );
  SDFFX1 DFF_1284_Q_reg ( .D(g25707), .SI(g5644), .SE(n10713), .CLK(n11096), 
        .Q(g5152), .QN(n5883) );
  SDFFX1 DFF_1285_Q_reg ( .D(g24339), .SI(g5152), .SE(n10713), .CLK(n11096), 
        .Q(g5352), .QN(n10525) );
  SDFFX1 DFF_1286_Q_reg ( .D(g11770), .SI(g5352), .SE(n10740), .CLK(n11123), 
        .Q(g8915) );
  SDFFX1 DFF_1288_Q_reg ( .D(g34443), .SI(g8915), .SE(n10792), .CLK(n11175), 
        .Q(g2775), .QN(n5378) );
  SDFFX1 DFF_1289_Q_reg ( .D(g34619), .SI(g2775), .SE(n10740), .CLK(n11123), 
        .Q(g2922), .QN(n10559) );
  SDFFX1 DFF_1290_Q_reg ( .D(g29234), .SI(g2922), .SE(n10740), .CLK(n11123), 
        .Q(test_so90), .QN(n10665) );
  SDFFX1 DFF_1291_Q_reg ( .D(g30503), .SI(test_si91), .SE(n10752), .CLK(n11135), .Q(g5893), .QN(n10308) );
  SDFFX1 DFF_1293_Q_reg ( .D(g16718), .SI(g5893), .SE(n10788), .CLK(n11171), 
        .Q(g16603), .QN(n10357) );
  SDFFX1 DFF_1294_Q_reg ( .D(g30550), .SI(g16603), .SE(n10735), .CLK(n11118), 
        .Q(g6617), .QN(n10423) );
  SDFFX1 DFF_1295_Q_reg ( .D(g33001), .SI(g6617), .SE(n10725), .CLK(n11108), 
        .Q(g2060), .QN(n5507) );
  SDFFX1 DFF_1296_Q_reg ( .D(g33040), .SI(g2060), .SE(n10719), .CLK(n11102), 
        .Q(g4512), .QN(n10265) );
  SDFFX1 DFF_1297_Q_reg ( .D(g30492), .SI(g4512), .SE(n10721), .CLK(n11104), 
        .Q(g5599), .QN(n10343) );
  SDFFX1 DFF_1298_Q_reg ( .D(g25664), .SI(g5599), .SE(n10800), .CLK(n11183), 
        .Q(g3401) );
  SDFFX1 DFF_1299_Q_reg ( .D(g26944), .SI(g3401), .SE(n10746), .CLK(n11129), 
        .Q(g4366) );
  SDFFX1 DFF_1300_Q_reg ( .D(test_so26), .SI(g4366), .SE(n10747), .CLK(n11130), 
        .Q(g16722) );
  SDFFX1 DFF_1301_Q_reg ( .D(g34614), .SI(g16722), .SE(n10747), .CLK(n11130), 
        .Q(g29214), .QN(n5342) );
  SDFFX1 DFF_1302_Q_reg ( .D(g29260), .SI(g29214), .SE(n10703), .CLK(n11086), 
        .Q(g3129) );
  SDFFX1 DFF_1303_Q_reg ( .D(g16686), .SI(g3129), .SE(n10766), .CLK(n11149), 
        .Q(test_so91) );
  SDFFX1 DFF_1304_Q_reg ( .D(g33047), .SI(test_si92), .SE(n10778), .CLK(n11161), .Q(g5170), .QN(n10586) );
  SDFFX1 DFF_1305_Q_reg ( .D(g24298), .SI(g5170), .SE(n10778), .CLK(n11161), 
        .Q(g26959) );
  SDFFX1 DFF_1306_Q_reg ( .D(g25733), .SI(g26959), .SE(n10712), .CLK(n11095), 
        .Q(g5821), .QN(n5429) );
  SDFFX1 DFF_1307_Q_reg ( .D(g30536), .SI(g5821), .SE(n10761), .CLK(n11144), 
        .Q(g6299), .QN(n10371) );
  SDFFX1 DFF_1308_Q_reg ( .D(g7916), .SI(g6299), .SE(n10761), .CLK(n11144), 
        .Q(g8416), .QN(n10148) );
  SDFFX1 DFF_1310_Q_reg ( .D(g29246), .SI(g8416), .SE(n10725), .CLK(n11108), 
        .Q(g2079), .QN(n10595) );
  SDFFX1 DFF_1311_Q_reg ( .D(g34261), .SI(g2079), .SE(n10714), .CLK(n11097), 
        .Q(g4698), .QN(n5862) );
  SDFFX1 DFF_1312_Q_reg ( .D(g33611), .SI(g4698), .SE(n10747), .CLK(n11130), 
        .Q(g3703), .QN(n5399) );
  SDFFX1 DFF_1313_Q_reg ( .D(g25638), .SI(g3703), .SE(n10747), .CLK(n11130), 
        .Q(g1559), .QN(n5441) );
  SDFFX1 DFF_1314_Q_reg ( .D(g34728), .SI(g1559), .SE(n10704), .CLK(n11087), 
        .Q(n9247), .QN(n19417) );
  SDFFX1 DFF_1315_Q_reg ( .D(g29222), .SI(n9247), .SE(n10710), .CLK(n11093), 
        .Q(g411), .QN(n5629) );
  SDFFX1 DFF_1316_Q_reg ( .D(g25742), .SI(g411), .SE(n10778), .CLK(n11161), 
        .Q(test_so92), .QN(n5718) );
  SDFFX1 DFF_1317_Q_reg ( .D(g30449), .SI(test_si93), .SE(n10731), .CLK(n11114), .Q(g3953), .QN(n10366) );
  SDFFX1 DFF_1319_Q_reg ( .D(g34608), .SI(g3953), .SE(n10773), .CLK(n11156), 
        .Q(g2704), .QN(n5377) );
  SDFFX1 DFF_1320_Q_reg ( .D(g24345), .SI(g2704), .SE(n10799), .CLK(n11182), 
        .Q(g6035), .QN(n5528) );
  SDFFX1 DFF_1322_Q_reg ( .D(g34977), .SI(g6035), .SE(n10716), .CLK(n11099), 
        .Q(n9245) );
  SDFFX1 DFF_1323_Q_reg ( .D(g25635), .SI(n9245), .SE(n10716), .CLK(n11099), 
        .Q(g1300), .QN(n5483) );
  SDFFX1 DFF_1324_Q_reg ( .D(g25686), .SI(g1300), .SE(n10739), .CLK(n11122), 
        .Q(g4057), .QN(n5711) );
  SDFFX1 DFF_1325_Q_reg ( .D(g30461), .SI(g4057), .SE(n10797), .CLK(n11180), 
        .Q(g5200), .QN(n10306) );
  SDFFX1 DFF_1326_Q_reg ( .D(g34466), .SI(g5200), .SE(n10759), .CLK(n11142), 
        .Q(g4843), .QN(n10209) );
  SDFFX1 DFF_1327_Q_reg ( .D(g31901), .SI(g4843), .SE(n10769), .CLK(n11152), 
        .Q(g5046), .QN(n5578) );
  SDFFX1 DFF_1328_Q_reg ( .D(n132), .SI(g5046), .SE(n10780), .CLK(n11163), .Q(
        g2250), .QN(n10314) );
  SDFFX1 DFF_1329_Q_reg ( .D(g26882), .SI(g2250), .SE(n10780), .CLK(n11163), 
        .Q(g26885), .QN(n5456) );
  SDFFX1 DFF_1330_Q_reg ( .D(g33041), .SI(g26885), .SE(n10782), .CLK(n11165), 
        .Q(test_so93) );
  SDFFX1 DFF_1331_Q_reg ( .D(g33011), .SI(test_si94), .SE(n10738), .CLK(n11121), .Q(g2453), .QN(n5373) );
  SDFFX1 DFF_1332_Q_reg ( .D(n503), .SI(g2453), .SE(n10713), .CLK(n11096), .Q(
        g5841), .QN(n5449) );
  SDFFX1 DFF_1335_Q_reg ( .D(g12300), .SI(g5841), .SE(n10713), .CLK(n11096), 
        .Q(g14694), .QN(n5705) );
  SDFFX1 DFF_1336_Q_reg ( .D(g34618), .SI(g14694), .SE(n10740), .CLK(n11123), 
        .Q(g2912), .QN(n10558) );
  SDFFX1 DFF_1337_Q_reg ( .D(g33010), .SI(g2912), .SE(n10729), .CLK(n11112), 
        .Q(g2357), .QN(n5276) );
  SDFFX1 DFF_1338_Q_reg ( .D(g8919), .SI(g2357), .SE(n10791), .CLK(n11174), 
        .Q(g8920) );
  SDFFX1 DFF_1339_Q_reg ( .D(g31864), .SI(g8920), .SE(n10755), .CLK(n11138), 
        .Q(g164), .QN(n5561) );
  SDFFX1 DFF_1340_Q_reg ( .D(g34630), .SI(g164), .SE(n10755), .CLK(n11138), 
        .Q(g4253), .QN(n5484) );
  SDFFX1 DFF_1341_Q_reg ( .D(g31898), .SI(g4253), .SE(n10794), .CLK(n11177), 
        .Q(g5016), .QN(n5369) );
  SDFFX1 DFF_1342_Q_reg ( .D(g25653), .SI(g5016), .SE(n10703), .CLK(n11086), 
        .Q(g3119), .QN(n5423) );
  SDFFX1 DFF_1343_Q_reg ( .D(g25632), .SI(g3119), .SE(n10724), .CLK(n11107), 
        .Q(g1351), .QN(n5322) );
  SDFFX1 DFF_1344_Q_reg ( .D(g32988), .SI(g1351), .SE(n10724), .CLK(n11107), 
        .Q(test_so94), .QN(n10638) );
  SDFFX1 DFF_1345_Q_reg ( .D(g33616), .SI(test_si95), .SE(n10715), .CLK(n11098), .Q(g4519) );
  SDFFX1 DFF_1346_Q_reg ( .D(g29280), .SI(g4519), .SE(n10714), .CLK(n11097), 
        .Q(g5115), .QN(n5743) );
  SDFFX1 DFF_1347_Q_reg ( .D(g33609), .SI(g5115), .SE(n10721), .CLK(n11104), 
        .Q(g3352), .QN(n5604) );
  SDFFX1 DFF_1348_Q_reg ( .D(g30563), .SI(g3352), .SE(n10721), .CLK(n11104), 
        .Q(g6657), .QN(n10292) );
  SDFFX1 DFF_1349_Q_reg ( .D(g33044), .SI(g6657), .SE(n10782), .CLK(n11165), 
        .Q(g4552) );
  SDFFX1 DFF_1350_Q_reg ( .D(g30437), .SI(g4552), .SE(n10796), .CLK(n11179), 
        .Q(g3893), .QN(n10311) );
  SDFFX1 DFF_1351_Q_reg ( .D(g30412), .SI(g3893), .SE(n10718), .CLK(n11101), 
        .Q(g3211) );
  SDFFX1 DFF_1352_Q_reg ( .D(g17604), .SI(g3211), .SE(n10774), .CLK(n11157), 
        .Q(g13049), .QN(n10503) );
  SDFFX1 DFF_1354_Q_reg ( .D(g16603), .SI(g13049), .SE(n10788), .CLK(n11171), 
        .Q(g16624), .QN(n10458) );
  SDFFX1 DFF_1355_Q_reg ( .D(g30491), .SI(g16624), .SE(n10788), .CLK(n11171), 
        .Q(g5595), .QN(n10470) );
  SDFFX1 DFF_1356_Q_reg ( .D(g30434), .SI(g5595), .SE(n10788), .CLK(n11171), 
        .Q(g3614), .QN(n10295) );
  SDFFX1 DFF_1357_Q_reg ( .D(g34612), .SI(g3614), .SE(n10743), .CLK(n11126), 
        .Q(test_so95) );
  SDFFX1 DFF_1358_Q_reg ( .D(g29259), .SI(test_si96), .SE(n10703), .CLK(n11086), .Q(g3125), .QN(n5781) );
  SDFFX1 DFF_1359_Q_reg ( .D(g13865), .SI(g3125), .SE(n10766), .CLK(n11149), 
        .Q(g16686) );
  SDFFX1 DFF_1360_Q_reg ( .D(g25681), .SI(g16686), .SE(n10700), .CLK(n11083), 
        .Q(g3821), .QN(n5428) );
  SDFFX1 DFF_1361_Q_reg ( .D(g25687), .SI(g3821), .SE(n10739), .CLK(n11122), 
        .Q(g4141), .QN(n5612) );
  SDFFX1 DFF_1362_Q_reg ( .D(g33617), .SI(g4141), .SE(n10782), .CLK(n11165), 
        .Q(g4570) );
  SDFFX1 DFF_1363_Q_reg ( .D(g30479), .SI(g4570), .SE(n10715), .CLK(n11098), 
        .Q(g5272), .QN(n10303) );
  SDFFX1 DFF_1364_Q_reg ( .D(g29256), .SI(g5272), .SE(n10787), .CLK(n11170), 
        .Q(g2735), .QN(n5600) );
  SDFFX1 DFF_1365_Q_reg ( .D(g28054), .SI(g2735), .SE(n10787), .CLK(n11170), 
        .Q(g728), .QN(n10283) );
  SDFFX1 DFF_1366_Q_reg ( .D(g30535), .SI(g728), .SE(n10799), .CLK(n11182), 
        .Q(g6295), .QN(n10300) );
  SDFFX1 DFF_1368_Q_reg ( .D(g30385), .SI(g6295), .SE(n10706), .CLK(n11089), 
        .Q(g2661), .QN(n5418) );
  SDFFX1 DFF_1369_Q_reg ( .D(g30361), .SI(g2661), .SE(n10754), .CLK(n11137), 
        .Q(g1988), .QN(n5783) );
  SDFFX1 DFF_1370_Q_reg ( .D(g25705), .SI(g1988), .SE(n10714), .CLK(n11097), 
        .Q(test_so96), .QN(n10654) );
  SDFFX1 DFF_1371_Q_reg ( .D(g24260), .SI(test_si97), .SE(n10790), .CLK(n11173), .Q(g1548), .QN(n5546) );
  SDFFX1 DFF_1372_Q_reg ( .D(g29257), .SI(g1548), .SE(n10702), .CLK(n11085), 
        .Q(g3106), .QN(n5742) );
  SDFFX1 DFF_1373_Q_reg ( .D(g34461), .SI(g3106), .SE(n10767), .CLK(n11150), 
        .Q(g4659), .QN(n10543) );
  SDFFX1 DFF_1374_Q_reg ( .D(g34258), .SI(g4659), .SE(n10767), .CLK(n11150), 
        .Q(g4358), .QN(n5348) );
  SDFFX1 DFF_1375_Q_reg ( .D(g32993), .SI(g4358), .SE(n10795), .CLK(n11178), 
        .Q(g1792), .QN(n5359) );
  SDFFX1 DFF_1376_Q_reg ( .D(g33992), .SI(g1792), .SE(n10744), .CLK(n11127), 
        .Q(g2084), .QN(n10195) );
  SDFFX1 DFF_1378_Q_reg ( .D(g30394), .SI(g2084), .SE(n10789), .CLK(n11172), 
        .Q(g3187), .QN(n10439) );
  SDFFX1 DFF_1379_Q_reg ( .D(g34449), .SI(g3187), .SE(n10789), .CLK(n11172), 
        .Q(g4311), .QN(n5323) );
  SDFFX1 DFF_1380_Q_reg ( .D(g34019), .SI(g4311), .SE(n10736), .CLK(n11119), 
        .Q(g2583), .QN(n5800) );
  SDFFX1 DFF_1381_Q_reg ( .D(g18597), .SI(g2583), .SE(n10736), .CLK(n11119), 
        .Q(n9240), .QN(DFF_1381_n1) );
  SDFFX1 DFF_1382_Q_reg ( .D(g29231), .SI(n9240), .SE(n10737), .CLK(n11120), 
        .Q(g1094), .QN(n5697) );
  SDFFX1 DFF_1383_Q_reg ( .D(g25682), .SI(g1094), .SE(n10700), .CLK(n11083), 
        .Q(test_so97), .QN(n10683) );
  SDFFX1 DFF_1384_Q_reg ( .D(g21897), .SI(test_si98), .SE(n10756), .CLK(n11139), .Q(g4284), .QN(n10593) );
  SDFFX1 DFF_1386_Q_reg ( .D(g30395), .SI(g4284), .SE(n10790), .CLK(n11173), 
        .Q(g3191), .QN(n10287) );
  SDFFX1 DFF_1387_Q_reg ( .D(g21892), .SI(g3191), .SE(n10763), .CLK(n11146), 
        .Q(g4239), .QN(n10210) );
  SDFFX1 DFF_1389_Q_reg ( .D(g8789), .SI(g4239), .SE(n10763), .CLK(n11146), 
        .Q(g4180), .QN(n5380) );
  SDFFX1 DFF_1390_Q_reg ( .D(g28048), .SI(g4180), .SE(n10709), .CLK(n11092), 
        .Q(g691), .QN(n5520) );
  SDFFX1 DFF_1391_Q_reg ( .D(g34723), .SI(g691), .SE(n10746), .CLK(n11129), 
        .Q(g534), .QN(n5490) );
  SDFFX1 DFF_1393_Q_reg ( .D(g25598), .SI(g534), .SE(n10785), .CLK(n11168), 
        .Q(g385), .QN(n5632) );
  SDFFX1 DFF_1394_Q_reg ( .D(g33987), .SI(g385), .SE(n10744), .CLK(n11127), 
        .Q(g2004), .QN(n5818) );
  SDFFX1 DFF_1395_Q_reg ( .D(g30380), .SI(g2004), .SE(n10717), .CLK(n11100), 
        .Q(g2527), .QN(n5420) );
  SDFFX1 DFF_1396_Q_reg ( .D(g9555), .SI(g2527), .SE(n10783), .CLK(n11166), 
        .Q(g5456) );
  SDFFX1 DFF_1397_Q_reg ( .D(g26965), .SI(g5456), .SE(n10798), .CLK(n11181), 
        .Q(n6007), .QN(n10695) );
  SDFFX1 DFF_1398_Q_reg ( .D(g25706), .SI(n6007), .SE(n10804), .CLK(n11187), 
        .Q(test_so98), .QN(n10682) );
  SDFFX1 DFF_1399_Q_reg ( .D(g30458), .SI(test_si99), .SE(n10794), .CLK(n11177), .Q(g4507), .QN(n5846) );
  SDFFX1 DFF_1400_Q_reg ( .D(g24338), .SI(g4507), .SE(n10718), .CLK(n11101), 
        .Q(g5348), .QN(n10526) );
  SDFFX1 DFF_1401_Q_reg ( .D(g30400), .SI(g5348), .SE(n10718), .CLK(n11101), 
        .Q(g3223), .QN(n10408) );
  SDFFX1 DFF_1403_Q_reg ( .D(g34623), .SI(g3223), .SE(n10803), .CLK(n11186), 
        .Q(g2970) );
  SDFFX1 DFF_1404_Q_reg ( .D(g24343), .SI(g2970), .SE(n10713), .CLK(n11096), 
        .Q(g5698), .QN(n10394) );
  SDFFX1 DFF_1406_Q_reg ( .D(g30473), .SI(g5698), .SE(n10799), .CLK(n11182), 
        .Q(g5260), .QN(n10360) );
  SDFFX1 DFF_1407_Q_reg ( .D(g24252), .SI(g5260), .SE(n10762), .CLK(n11145), 
        .Q(g1521) );
  SDFFX1 DFF_1408_Q_reg ( .D(g33028), .SI(g1521), .SE(n10762), .CLK(n11145), 
        .Q(g3522), .QN(n5383) );
  SDFFX1 DFF_1409_Q_reg ( .D(g29258), .SI(g3522), .SE(n10703), .CLK(n11086), 
        .Q(g3115), .QN(n10170) );
  SDFFX1 DFF_1410_Q_reg ( .D(g30407), .SI(g3115), .SE(n10722), .CLK(n11105), 
        .Q(g3251), .QN(n10358) );
  SDFFX1 DFF_1411_Q_reg ( .D(g26958), .SI(g3251), .SE(n10746), .CLK(n11129), 
        .Q(g12832) );
  SDFFX1 DFF_1412_Q_reg ( .D(g34457), .SI(g12832), .SE(n10746), .CLK(n11129), 
        .Q(test_so99) );
  SDFFX1 DFF_1413_Q_reg ( .D(g33568), .SI(test_si100), .SE(n10764), .CLK(
        n11147), .Q(g1996), .QN(n5355) );
  SDFFX1 DFF_1414_Q_reg ( .D(g25663), .SI(g1996), .SE(n10800), .CLK(n11183), 
        .Q(g8342) );
  SDFFX1 DFF_1415_Q_reg ( .D(g26964), .SI(g8342), .SE(n10719), .CLK(n11102), 
        .Q(g4515), .QN(n10533) );
  SDFFX1 DFF_1416_Q_reg ( .D(g8786), .SI(g4515), .SE(n10737), .CLK(n11120), 
        .Q(g8787) );
  SDFFX1 DFF_1417_Q_reg ( .D(g34735), .SI(g8787), .SE(n10716), .CLK(n11099), 
        .Q(g4300), .QN(n5639) );
  SDFFX1 DFF_1418_Q_reg ( .D(g30352), .SI(g4300), .SE(n10723), .CLK(n11106), 
        .Q(n9236), .QN(n19400) );
  SDFFX1 DFF_1419_Q_reg ( .D(g33543), .SI(n9236), .SE(n10723), .CLK(n11106), 
        .Q(g1379), .QN(n10190) );
  SDFFX1 DFF_1420_Q_reg ( .D(g24271), .SI(g1379), .SE(n10791), .CLK(n11174), 
        .Q(g11388), .QN(n5433) );
  SDFFX1 DFF_1422_Q_reg ( .D(g33981), .SI(g11388), .SE(n10758), .CLK(n11141), 
        .Q(g1878), .QN(n5793) );
  SDFFX1 DFF_1423_Q_reg ( .D(g30500), .SI(g1878), .SE(n10721), .CLK(n11104), 
        .Q(g5619), .QN(n10288) );
  SDFFX1 DFF_1424_Q_reg ( .D(g34649), .SI(g5619), .SE(n10803), .CLK(n11186), 
        .Q(g71), .QN(n19418) );
  SDFFX1 DFF_1425_Q_reg ( .D(g29277), .SI(g71), .SE(n10715), .CLK(n11098), .Q(
        test_so100) );
  SDFFX1 DFF_748_Q_reg ( .D(n1436), .SI(g4704), .SE(n10772), .CLK(n11155), .Q(
        g22), .QN(n10226) );
  SDFFX1 DFF_591_Q_reg ( .D(g25612), .SI(g3897), .SE(n10771), .CLK(n11154), 
        .Q(g518), .QN(n5287) );
  SDFFX1 DFF_845_Q_reg ( .D(g28060), .SI(g626), .SE(n10787), .CLK(n11170), .Q(
        g2729), .QN(n10274) );
  HADDX1 Trojan_U1_1_30 ( .A0(counter_30), .B0(carry_30), .C1(carry_31), .SO(
        N31) );
  HADDX1 Trojan_U1_1_4 ( .A0(counter_4), .B0(carry_4), .C1(carry_5), .SO(N5)
         );
  HADDX1 Trojan_U1_1_5 ( .A0(counter_5), .B0(carry_5), .C1(carry_6), .SO(N6)
         );
  HADDX1 Trojan_U1_1_6 ( .A0(counter_6), .B0(carry_6), .C1(carry_7), .SO(N7)
         );
  HADDX1 Trojan_U1_1_7 ( .A0(counter_7), .B0(carry_7), .C1(carry_8), .SO(N8)
         );
  HADDX1 Trojan_U1_1_8 ( .A0(counter_8), .B0(carry_8), .C1(carry_9), .SO(N9)
         );
  HADDX1 Trojan_U1_1_9 ( .A0(counter_9), .B0(carry_9), .C1(carry_10), .SO(N10)
         );
  HADDX1 Trojan_U1_1_10 ( .A0(counter_10), .B0(carry_10), .C1(carry_11), .SO(
        N11) );
  HADDX1 Trojan_U1_1_11 ( .A0(counter_11), .B0(carry_11), .C1(carry_12), .SO(
        N12) );
  HADDX1 Trojan_U1_1_12 ( .A0(counter_12), .B0(carry_12), .C1(carry_13), .SO(
        N13) );
  HADDX1 Trojan_U1_1_13 ( .A0(counter_13), .B0(carry_13), .C1(carry_14), .SO(
        N14) );
  HADDX1 Trojan_U1_1_14 ( .A0(counter_14), .B0(carry_14), .C1(carry_15), .SO(
        N15) );
  HADDX1 Trojan_U1_1_22 ( .A0(counter_22), .B0(carry_22), .C1(carry_23), .SO(
        N23) );
  HADDX1 Trojan_U1_1_23 ( .A0(counter_23), .B0(carry_23), .C1(carry_24), .SO(
        N24) );
  HADDX1 Trojan_U1_1_24 ( .A0(counter_24), .B0(carry_24), .C1(carry_25), .SO(
        N25) );
  HADDX1 Trojan_U1_1_25 ( .A0(counter_25), .B0(carry_25), .C1(carry_26), .SO(
        N26) );
  HADDX1 Trojan_U1_1_1 ( .A0(counter_1), .B0(counter_0), .C1(carry_2), .SO(N2)
         );
  HADDX1 Trojan_U1_1_2 ( .A0(counter_2), .B0(carry_2), .C1(carry_3), .SO(N3)
         );
  HADDX1 Trojan_U1_1_3 ( .A0(counter_3), .B0(carry_3), .C1(carry_4), .SO(N4)
         );
  HADDX1 Trojan_U1_1_15 ( .A0(counter_15), .B0(carry_15), .C1(carry_16), .SO(
        N16) );
  HADDX1 Trojan_U1_1_16 ( .A0(counter_16), .B0(carry_16), .C1(carry_17), .SO(
        N17) );
  HADDX1 Trojan_U1_1_17 ( .A0(counter_17), .B0(carry_17), .C1(carry_18), .SO(
        N18) );
  HADDX1 Trojan_U1_1_18 ( .A0(counter_18), .B0(carry_18), .C1(carry_19), .SO(
        N19) );
  HADDX1 Trojan_U1_1_19 ( .A0(counter_19), .B0(carry_19), .C1(carry_20), .SO(
        N20) );
  HADDX1 Trojan_U1_1_20 ( .A0(counter_20), .B0(carry_20), .C1(carry_21), .SO(
        N21) );
  HADDX1 Trojan_U1_1_21 ( .A0(counter_21), .B0(carry_21), .C1(carry_22), .SO(
        N22) );
  HADDX1 Trojan_U1_1_26 ( .A0(counter_26), .B0(carry_26), .C1(carry_27), .SO(
        N27) );
  HADDX1 Trojan_U1_1_27 ( .A0(counter_27), .B0(carry_27), .C1(carry_28), .SO(
        N28) );
  HADDX1 Trojan_U1_1_28 ( .A0(counter_28), .B0(carry_28), .C1(carry_29), .SO(
        N29) );
  HADDX1 Trojan_U1_1_29 ( .A0(counter_29), .B0(carry_29), .C1(carry_30), .SO(
        N30) );
  INVX0 Trojan_U1 ( .INP(counter_0), .ZN(N1) );
  XOR2X1 Trojan_U2 ( .IN1(carry_31), .IN2(counter_31), .Q(N32) );
  DFFARX1 Trojan_counter_reg_31_ ( .D(N32), .CLK(n37), .RSTB(n10698), .Q(
        counter_31), .QN(n73) );
  DFFARX1 Trojan_counter_reg_1_ ( .D(N2), .CLK(n37), .RSTB(n10697), .Q(
        counter_1) );
  DFFARX1 Trojan_counter_reg_2_ ( .D(N3), .CLK(n37), .RSTB(n87), .Q(counter_2)
         );
  DFFARX1 Trojan_counter_reg_3_ ( .D(N4), .CLK(n37), .RSTB(n10698), .Q(
        counter_3), .QN(n86) );
  DFFARX1 Trojan_counter_reg_15_ ( .D(N16), .CLK(n37), .RSTB(n10697), .Q(
        counter_15), .QN(n85) );
  DFFARX1 Trojan_counter_reg_16_ ( .D(N17), .CLK(n37), .RSTB(n87), .Q(
        counter_16), .QN(n84) );
  DFFARX1 Trojan_counter_reg_17_ ( .D(N18), .CLK(n37), .RSTB(n10698), .Q(
        counter_17), .QN(n83) );
  DFFARX1 Trojan_counter_reg_18_ ( .D(N19), .CLK(n37), .RSTB(n10697), .Q(
        counter_18), .QN(n82) );
  DFFARX1 Trojan_counter_reg_19_ ( .D(N20), .CLK(n37), .RSTB(n87), .Q(
        counter_19), .QN(n81) );
  DFFARX1 Trojan_counter_reg_20_ ( .D(N21), .CLK(n37), .RSTB(n10698), .Q(
        counter_20), .QN(n80) );
  DFFARX1 Trojan_counter_reg_21_ ( .D(N22), .CLK(n37), .RSTB(n10697), .Q(
        counter_21), .QN(n79) );
  DFFARX1 Trojan_counter_reg_26_ ( .D(N27), .CLK(n37), .RSTB(n87), .Q(
        counter_26), .QN(n78) );
  DFFARX1 Trojan_counter_reg_27_ ( .D(N28), .CLK(n37), .RSTB(n10698), .Q(
        counter_27), .QN(n77) );
  DFFARX1 Trojan_counter_reg_28_ ( .D(N29), .CLK(n37), .RSTB(n10697), .Q(
        counter_28), .QN(n76) );
  DFFARX1 Trojan_counter_reg_29_ ( .D(N30), .CLK(n37), .RSTB(n87), .Q(
        counter_29), .QN(n75) );
  DFFARX1 Trojan_counter_reg_30_ ( .D(N31), .CLK(n37), .RSTB(n10698), .Q(
        counter_30), .QN(n74) );
  DFFARX1 Trojan_counter_reg_7_ ( .D(N8), .CLK(n37), .RSTB(n10697), .Q(
        counter_7) );
  DFFARX1 Trojan_counter_reg_11_ ( .D(N12), .CLK(n37), .RSTB(n87), .Q(
        counter_11) );
  DFFARX1 Trojan_counter_reg_25_ ( .D(N26), .CLK(n37), .RSTB(n10698), .Q(
        counter_25) );
  DFFARX1 Trojan_counter_reg_6_ ( .D(N7), .CLK(n37), .RSTB(n10697), .Q(
        counter_6) );
  DFFARX1 Trojan_counter_reg_10_ ( .D(N11), .CLK(n37), .RSTB(n87), .Q(
        counter_10) );
  DFFARX1 Trojan_counter_reg_12_ ( .D(N13), .CLK(n37), .RSTB(n10698), .Q(
        counter_12) );
  DFFARX1 Trojan_counter_reg_24_ ( .D(N25), .CLK(n37), .RSTB(n10697), .Q(
        counter_24) );
  DFFARX1 Trojan_counter_reg_4_ ( .D(N5), .CLK(n37), .RSTB(n87), .Q(counter_4)
         );
  DFFARX1 Trojan_counter_reg_5_ ( .D(N6), .CLK(n37), .RSTB(n10698), .Q(
        counter_5) );
  DFFARX1 Trojan_counter_reg_9_ ( .D(N10), .CLK(n37), .RSTB(n10697), .Q(
        counter_9) );
  DFFARX1 Trojan_counter_reg_14_ ( .D(N15), .CLK(n37), .RSTB(n87), .Q(
        counter_14) );
  DFFARX1 Trojan_counter_reg_23_ ( .D(N24), .CLK(n37), .RSTB(n10698), .Q(
        counter_23) );
  DFFARX1 Trojan_counter_reg_8_ ( .D(N9), .CLK(n37), .RSTB(n10697), .Q(
        counter_8) );
  DFFARX1 Trojan_counter_reg_13_ ( .D(N14), .CLK(n37), .RSTB(n87), .Q(
        counter_13) );
  DFFARX1 Trojan_counter_reg_22_ ( .D(N23), .CLK(n37), .RSTB(n10698), .Q(
        counter_22) );
  DFFARX1 Trojan_counter_reg_0_ ( .D(N1), .CLK(n37), .RSTB(n10697), .Q(
        counter_0) );
  NAND4X0 Trojan_U14 ( .IN1(n293), .IN2(n571), .IN3(n2461), .IN4(n58), .QN(n87) );
  INVX0 Trojan_U15 ( .INP(n59), .ZN(n58) );
  NOR4X0 Trojan_U16 ( .IN1(n293), .IN2(n571), .IN3(n2461), .IN4(n59), .QN(n37)
         );
  NAND3X0 Trojan_U17 ( .IN1(n2601), .IN2(n5111), .IN3(n60), .QN(n59) );
  AND3X1 Trojan_U18 ( .IN1(n268), .IN2(n97), .IN3(n95), .Q(n60) );
  NOR4X0 Trojan_U19 ( .IN1(n61), .IN2(n62), .IN3(n63), .IN4(n64), .QN(
        Trigger_out) );
  NAND4X0 Trojan_U20 ( .IN1(n78), .IN2(n77), .IN3(n76), .IN4(n75), .QN(n64) );
  NAND4X0 Trojan_U21 ( .IN1(n74), .IN2(n73), .IN3(counter_6), .IN4(counter_5), 
        .QN(n63) );
  NAND4X0 Trojan_U22 ( .IN1(n80), .IN2(n79), .IN3(n81), .IN4(n65), .QN(n62) );
  NOR4X0 Trojan_U23 ( .IN1(counter_25), .IN2(counter_24), .IN3(counter_23), 
        .IN4(counter_22), .QN(n65) );
  NAND4X0 Trojan_U24 ( .IN1(n66), .IN2(n67), .IN3(n68), .IN4(n69), .QN(n61) );
  NOR4X0 Trojan_U25 ( .IN1(n70), .IN2(counter_12), .IN3(counter_14), .IN4(
        counter_13), .QN(n69) );
  NAND4X0 Trojan_U26 ( .IN1(n85), .IN2(n84), .IN3(n83), .IN4(n82), .QN(n70) );
  NOR4X0 Trojan_U27 ( .IN1(counter_11), .IN2(counter_10), .IN3(counter_9), 
        .IN4(counter_8), .QN(n68) );
  MUX21X1 Trojan_U28 ( .IN1(n71), .IN2(n72), .S(n86), .Q(n67) );
  OA21X1 Trojan_U29 ( .IN1(counter_1), .IN2(counter_0), .IN3(counter_2), .Q(
        n72) );
  NAND2X0 Trojan_U30 ( .IN1(counter_2), .IN2(counter_1), .QN(n71) );
  NOR2X0 Trojan_U31 ( .IN1(counter_7), .IN2(counter_4), .QN(n66) );
  MUX21X1 Trojan_Paylod ( .IN1(g10122_Tj), .IN2(g25715), .S(Trigger_out), .Q(
        g10122) );
  INVX0 U10583 ( .INP(n87), .ZN(n10696) );
  INVX0 U10584 ( .INP(n10696), .ZN(n10697) );
  INVX0 U10585 ( .INP(n10696), .ZN(n10698) );
  NBUFFX2 U10586 ( .INP(n10989), .Z(n10908) );
  NBUFFX2 U10587 ( .INP(n10983), .Z(n10937) );
  NBUFFX2 U10588 ( .INP(n10978), .Z(n10965) );
  NBUFFX2 U10589 ( .INP(n10977), .Z(n10967) );
  NBUFFX2 U10590 ( .INP(n10979), .Z(n10956) );
  NBUFFX2 U10591 ( .INP(n10981), .Z(n10948) );
  NBUFFX2 U10592 ( .INP(n10977), .Z(n10969) );
  NBUFFX2 U10593 ( .INP(n10978), .Z(n10962) );
  NBUFFX2 U10594 ( .INP(n10983), .Z(n10938) );
  NBUFFX2 U10595 ( .INP(n10977), .Z(n10970) );
  NBUFFX2 U10596 ( .INP(n10979), .Z(n10958) );
  NBUFFX2 U10597 ( .INP(n10979), .Z(n10960) );
  NBUFFX2 U10598 ( .INP(n10978), .Z(n10964) );
  NBUFFX2 U10599 ( .INP(n10979), .Z(n10957) );
  NBUFFX2 U10600 ( .INP(n10983), .Z(n10939) );
  NBUFFX2 U10601 ( .INP(n10981), .Z(n10947) );
  NBUFFX2 U10602 ( .INP(n10982), .Z(n10944) );
  NBUFFX2 U10603 ( .INP(n10982), .Z(n10941) );
  NBUFFX2 U10604 ( .INP(n10982), .Z(n10942) );
  NBUFFX2 U10605 ( .INP(n10979), .Z(n10959) );
  NBUFFX2 U10606 ( .INP(n10980), .Z(n10954) );
  NBUFFX2 U10607 ( .INP(n10981), .Z(n10950) );
  NBUFFX2 U10608 ( .INP(n10978), .Z(n10961) );
  NBUFFX2 U10609 ( .INP(n10977), .Z(n10968) );
  NBUFFX2 U10610 ( .INP(n10977), .Z(n10966) );
  NBUFFX2 U10611 ( .INP(n10980), .Z(n10953) );
  NBUFFX2 U10612 ( .INP(n10981), .Z(n10949) );
  NBUFFX2 U10613 ( .INP(n10982), .Z(n10943) );
  NBUFFX2 U10614 ( .INP(n10980), .Z(n10955) );
  NBUFFX2 U10615 ( .INP(n10982), .Z(n10945) );
  NBUFFX2 U10616 ( .INP(n10980), .Z(n10952) );
  NBUFFX2 U10617 ( .INP(n10978), .Z(n10963) );
  NBUFFX2 U10618 ( .INP(n10981), .Z(n10946) );
  NBUFFX2 U10619 ( .INP(n10983), .Z(n10940) );
  NBUFFX2 U10620 ( .INP(n10980), .Z(n10951) );
  NBUFFX2 U10621 ( .INP(n10990), .Z(n10904) );
  NBUFFX2 U10622 ( .INP(n10990), .Z(n10902) );
  NBUFFX2 U10623 ( .INP(n10989), .Z(n10906) );
  NBUFFX2 U10624 ( .INP(n10989), .Z(n10907) );
  NBUFFX2 U10625 ( .INP(n10990), .Z(n10903) );
  NBUFFX2 U10626 ( .INP(n10990), .Z(n10905) );
  NBUFFX2 U10627 ( .INP(n10984), .Z(n10932) );
  NBUFFX2 U10628 ( .INP(n10985), .Z(n10927) );
  NBUFFX2 U10629 ( .INP(n10985), .Z(n10930) );
  NBUFFX2 U10630 ( .INP(n10983), .Z(n10936) );
  NBUFFX2 U10631 ( .INP(n10986), .Z(n10922) );
  NBUFFX2 U10632 ( .INP(n10985), .Z(n10926) );
  NBUFFX2 U10633 ( .INP(n10984), .Z(n10935) );
  NBUFFX2 U10634 ( .INP(n10986), .Z(n10925) );
  NBUFFX2 U10635 ( .INP(n10984), .Z(n10933) );
  NBUFFX2 U10636 ( .INP(n10984), .Z(n10934) );
  NBUFFX2 U10637 ( .INP(n10984), .Z(n10931) );
  NBUFFX2 U10638 ( .INP(n10986), .Z(n10923) );
  NBUFFX2 U10639 ( .INP(n10985), .Z(n10928) );
  NBUFFX2 U10640 ( .INP(n10985), .Z(n10929) );
  NBUFFX2 U10641 ( .INP(n10987), .Z(n10920) );
  NBUFFX2 U10642 ( .INP(n10986), .Z(n10921) );
  NBUFFX2 U10643 ( .INP(n10986), .Z(n10924) );
  NBUFFX2 U10644 ( .INP(n11003), .Z(n10839) );
  NBUFFX2 U10645 ( .INP(n11003), .Z(n10840) );
  NBUFFX2 U10646 ( .INP(n10993), .Z(n10886) );
  NBUFFX2 U10647 ( .INP(n11002), .Z(n10843) );
  NBUFFX2 U10648 ( .INP(n10990), .Z(n10901) );
  NBUFFX2 U10649 ( .INP(n10995), .Z(n10880) );
  NBUFFX2 U10650 ( .INP(n10992), .Z(n10893) );
  NBUFFX2 U10651 ( .INP(n11001), .Z(n10849) );
  NBUFFX2 U10652 ( .INP(n10997), .Z(n10869) );
  NBUFFX2 U10653 ( .INP(n10991), .Z(n10898) );
  NBUFFX2 U10654 ( .INP(n10992), .Z(n10894) );
  NBUFFX2 U10655 ( .INP(n11001), .Z(n10848) );
  NBUFFX2 U10656 ( .INP(n10998), .Z(n10863) );
  NBUFFX2 U10657 ( .INP(n11000), .Z(n10851) );
  NBUFFX2 U10658 ( .INP(n10997), .Z(n10870) );
  NBUFFX2 U10659 ( .INP(n10996), .Z(n10874) );
  NBUFFX2 U10660 ( .INP(n10998), .Z(n10861) );
  NBUFFX2 U10661 ( .INP(n10994), .Z(n10883) );
  NBUFFX2 U10662 ( .INP(n11002), .Z(n10845) );
  NBUFFX2 U10663 ( .INP(n10992), .Z(n10891) );
  NBUFFX2 U10664 ( .INP(n10992), .Z(n10892) );
  NBUFFX2 U10665 ( .INP(n10993), .Z(n10888) );
  NBUFFX2 U10666 ( .INP(n10996), .Z(n10871) );
  NBUFFX2 U10667 ( .INP(n10998), .Z(n10865) );
  NBUFFX2 U10668 ( .INP(n11000), .Z(n10855) );
  NBUFFX2 U10669 ( .INP(n10998), .Z(n10862) );
  NBUFFX2 U10670 ( .INP(n11000), .Z(n10852) );
  NBUFFX2 U10671 ( .INP(n11001), .Z(n10850) );
  NBUFFX2 U10672 ( .INP(n10994), .Z(n10881) );
  NBUFFX2 U10673 ( .INP(n10993), .Z(n10887) );
  NBUFFX2 U10674 ( .INP(n10991), .Z(n10896) );
  NBUFFX2 U10675 ( .INP(n10994), .Z(n10885) );
  NBUFFX2 U10676 ( .INP(n10995), .Z(n10876) );
  NBUFFX2 U10677 ( .INP(n10994), .Z(n10882) );
  NBUFFX2 U10678 ( .INP(n10997), .Z(n10867) );
  NBUFFX2 U10679 ( .INP(n10991), .Z(n10899) );
  NBUFFX2 U10680 ( .INP(n10994), .Z(n10884) );
  NBUFFX2 U10681 ( .INP(n10995), .Z(n10879) );
  NBUFFX2 U10682 ( .INP(n10999), .Z(n10860) );
  NBUFFX2 U10683 ( .INP(n10991), .Z(n10900) );
  NBUFFX2 U10684 ( .INP(n11002), .Z(n10842) );
  NBUFFX2 U10685 ( .INP(n11002), .Z(n10841) );
  NBUFFX2 U10686 ( .INP(n10995), .Z(n10878) );
  NBUFFX2 U10687 ( .INP(n10996), .Z(n10875) );
  NBUFFX2 U10688 ( .INP(n10997), .Z(n10868) );
  NBUFFX2 U10689 ( .INP(n10998), .Z(n10864) );
  NBUFFX2 U10690 ( .INP(n10992), .Z(n10895) );
  NBUFFX2 U10691 ( .INP(n10999), .Z(n10857) );
  NBUFFX2 U10692 ( .INP(n10991), .Z(n10897) );
  NBUFFX2 U10693 ( .INP(n10993), .Z(n10890) );
  NBUFFX2 U10694 ( .INP(n10997), .Z(n10866) );
  NBUFFX2 U10695 ( .INP(n10996), .Z(n10872) );
  NBUFFX2 U10696 ( .INP(n10996), .Z(n10873) );
  NBUFFX2 U10697 ( .INP(n10999), .Z(n10858) );
  NBUFFX2 U10698 ( .INP(n11000), .Z(n10853) );
  NBUFFX2 U10699 ( .INP(n11001), .Z(n10846) );
  NBUFFX2 U10700 ( .INP(n11000), .Z(n10854) );
  NBUFFX2 U10701 ( .INP(n11001), .Z(n10847) );
  NBUFFX2 U10702 ( .INP(n10999), .Z(n10856) );
  NBUFFX2 U10703 ( .INP(n10995), .Z(n10877) );
  NBUFFX2 U10704 ( .INP(n11002), .Z(n10844) );
  NBUFFX2 U10705 ( .INP(n10999), .Z(n10859) );
  NBUFFX2 U10706 ( .INP(n10993), .Z(n10889) );
  NBUFFX2 U10707 ( .INP(n10988), .Z(n10912) );
  NBUFFX2 U10708 ( .INP(n10987), .Z(n10918) );
  NBUFFX2 U10709 ( .INP(n10988), .Z(n10913) );
  NBUFFX2 U10710 ( .INP(n10987), .Z(n10917) );
  NBUFFX2 U10711 ( .INP(n10988), .Z(n10911) );
  NBUFFX2 U10712 ( .INP(n10989), .Z(n10909) );
  NBUFFX2 U10713 ( .INP(n10987), .Z(n10919) );
  NBUFFX2 U10714 ( .INP(n10987), .Z(n10916) );
  NBUFFX2 U10715 ( .INP(n10988), .Z(n10914) );
  NBUFFX2 U10716 ( .INP(n10988), .Z(n10915) );
  NBUFFX2 U10717 ( .INP(n10989), .Z(n10910) );
  NBUFFX2 U10718 ( .INP(n10827), .Z(n10700) );
  NBUFFX2 U10719 ( .INP(n10827), .Z(n10699) );
  NBUFFX2 U10720 ( .INP(n10824), .Z(n10712) );
  NBUFFX2 U10721 ( .INP(n10819), .Z(n10738) );
  NBUFFX2 U10722 ( .INP(n10808), .Z(n10795) );
  NBUFFX2 U10723 ( .INP(n10823), .Z(n10716) );
  NBUFFX2 U10724 ( .INP(n10810), .Z(n10783) );
  NBUFFX2 U10725 ( .INP(n10809), .Z(n10790) );
  NBUFFX2 U10726 ( .INP(n10812), .Z(n10773) );
  NBUFFX2 U10727 ( .INP(n10825), .Z(n10710) );
  NBUFFX2 U10728 ( .INP(n10821), .Z(n10727) );
  NBUFFX2 U10729 ( .INP(n10811), .Z(n10780) );
  NBUFFX2 U10730 ( .INP(n10818), .Z(n10745) );
  NBUFFX2 U10731 ( .INP(n10809), .Z(n10788) );
  NBUFFX2 U10732 ( .INP(n10820), .Z(n10735) );
  NBUFFX2 U10733 ( .INP(n10808), .Z(n10794) );
  NBUFFX2 U10734 ( .INP(n10821), .Z(n10728) );
  NBUFFX2 U10735 ( .INP(n10820), .Z(n10734) );
  NBUFFX2 U10736 ( .INP(n10826), .Z(n10702) );
  NBUFFX2 U10737 ( .INP(n10807), .Z(n10798) );
  NBUFFX2 U10738 ( .INP(n10822), .Z(n10722) );
  NBUFFX2 U10739 ( .INP(n10816), .Z(n10755) );
  NBUFFX2 U10740 ( .INP(n10811), .Z(n10776) );
  NBUFFX2 U10741 ( .INP(n10826), .Z(n10703) );
  NBUFFX2 U10742 ( .INP(n10816), .Z(n10752) );
  NBUFFX2 U10743 ( .INP(n10821), .Z(n10729) );
  NBUFFX2 U10744 ( .INP(n10824), .Z(n10714) );
  NBUFFX2 U10745 ( .INP(n10815), .Z(n10756) );
  NBUFFX2 U10746 ( .INP(n10810), .Z(n10781) );
  NBUFFX2 U10747 ( .INP(n10814), .Z(n10761) );
  NBUFFX2 U10748 ( .INP(n10816), .Z(n10754) );
  NBUFFX2 U10749 ( .INP(n10822), .Z(n10724) );
  NBUFFX2 U10750 ( .INP(n10813), .Z(n10769) );
  NBUFFX2 U10751 ( .INP(n10817), .Z(n10746) );
  NBUFFX2 U10752 ( .INP(n10812), .Z(n10775) );
  NBUFFX2 U10753 ( .INP(n10816), .Z(n10753) );
  NBUFFX2 U10754 ( .INP(n10826), .Z(n10701) );
  NBUFFX2 U10755 ( .INP(n10819), .Z(n10736) );
  NBUFFX2 U10756 ( .INP(n10807), .Z(n10799) );
  NBUFFX2 U10757 ( .INP(n10808), .Z(n10793) );
  NBUFFX2 U10758 ( .INP(n10811), .Z(n10778) );
  NBUFFX2 U10759 ( .INP(n10823), .Z(n10718) );
  NBUFFX2 U10760 ( .INP(n10824), .Z(n10715) );
  NBUFFX2 U10761 ( .INP(n10814), .Z(n10764) );
  NBUFFX2 U10762 ( .INP(n10821), .Z(n10726) );
  NBUFFX2 U10763 ( .INP(n10825), .Z(n10709) );
  NBUFFX2 U10764 ( .INP(n10807), .Z(n10797) );
  NBUFFX2 U10765 ( .INP(n10807), .Z(n10796) );
  NBUFFX2 U10766 ( .INP(n10820), .Z(n10733) );
  NBUFFX2 U10767 ( .INP(n10812), .Z(n10774) );
  NBUFFX2 U10768 ( .INP(n10815), .Z(n10759) );
  NBUFFX2 U10769 ( .INP(n10815), .Z(n10757) );
  NBUFFX2 U10770 ( .INP(n10810), .Z(n10785) );
  NBUFFX2 U10771 ( .INP(n10821), .Z(n10730) );
  NBUFFX2 U10772 ( .INP(n10818), .Z(n10741) );
  NBUFFX2 U10773 ( .INP(n10807), .Z(n10800) );
  NBUFFX2 U10774 ( .INP(n10820), .Z(n10731) );
  NBUFFX2 U10775 ( .INP(n10813), .Z(n10770) );
  NBUFFX2 U10776 ( .INP(n10817), .Z(n10749) );
  NBUFFX2 U10777 ( .INP(n10809), .Z(n10786) );
  NBUFFX2 U10778 ( .INP(n10824), .Z(n10711) );
  NBUFFX2 U10779 ( .INP(n10815), .Z(n10760) );
  NBUFFX2 U10780 ( .INP(n10818), .Z(n10744) );
  NBUFFX2 U10781 ( .INP(n10814), .Z(n10763) );
  NBUFFX2 U10782 ( .INP(n10826), .Z(n10704) );
  NBUFFX2 U10783 ( .INP(n10818), .Z(n10743) );
  NBUFFX2 U10784 ( .INP(n10811), .Z(n10779) );
  NBUFFX2 U10785 ( .INP(n10813), .Z(n10768) );
  NBUFFX2 U10786 ( .INP(n10817), .Z(n10748) );
  NBUFFX2 U10787 ( .INP(n10814), .Z(n10762) );
  NBUFFX2 U10788 ( .INP(n10810), .Z(n10784) );
  NBUFFX2 U10789 ( .INP(n10822), .Z(n10721) );
  NBUFFX2 U10790 ( .INP(n10809), .Z(n10787) );
  NBUFFX2 U10791 ( .INP(n10826), .Z(n10705) );
  NBUFFX2 U10792 ( .INP(n10813), .Z(n10766) );
  NBUFFX2 U10793 ( .INP(n10812), .Z(n10772) );
  NBUFFX2 U10794 ( .INP(n10824), .Z(n10713) );
  NBUFFX2 U10795 ( .INP(n10825), .Z(n10706) );
  NBUFFX2 U10796 ( .INP(n10825), .Z(n10708) );
  NBUFFX2 U10797 ( .INP(n10817), .Z(n10747) );
  NBUFFX2 U10798 ( .INP(n10810), .Z(n10782) );
  NBUFFX2 U10799 ( .INP(n10825), .Z(n10707) );
  NBUFFX2 U10800 ( .INP(n10809), .Z(n10789) );
  NBUFFX2 U10801 ( .INP(n10822), .Z(n10723) );
  NBUFFX2 U10802 ( .INP(n10819), .Z(n10737) );
  NBUFFX2 U10803 ( .INP(n10808), .Z(n10791) );
  NBUFFX2 U10804 ( .INP(n10822), .Z(n10725) );
  NBUFFX2 U10805 ( .INP(n10814), .Z(n10765) );
  NBUFFX2 U10806 ( .INP(n10823), .Z(n10720) );
  NBUFFX2 U10807 ( .INP(n10819), .Z(n10739) );
  NBUFFX2 U10808 ( .INP(n10816), .Z(n10751) );
  NBUFFX2 U10809 ( .INP(n10813), .Z(n10767) );
  NBUFFX2 U10810 ( .INP(n10811), .Z(n10777) );
  NBUFFX2 U10811 ( .INP(n10818), .Z(n10742) );
  NBUFFX2 U10812 ( .INP(n10812), .Z(n10771) );
  NBUFFX2 U10813 ( .INP(n10819), .Z(n10740) );
  NBUFFX2 U10814 ( .INP(n10820), .Z(n10732) );
  NBUFFX2 U10815 ( .INP(n10823), .Z(n10719) );
  NBUFFX2 U10816 ( .INP(n10817), .Z(n10750) );
  NBUFFX2 U10817 ( .INP(n10823), .Z(n10717) );
  NBUFFX2 U10818 ( .INP(n10815), .Z(n10758) );
  NBUFFX2 U10819 ( .INP(n10808), .Z(n10792) );
  NBUFFX2 U10820 ( .INP(n11210), .Z(n11083) );
  NBUFFX2 U10821 ( .INP(n11210), .Z(n11082) );
  NBUFFX2 U10822 ( .INP(n11207), .Z(n11095) );
  NBUFFX2 U10823 ( .INP(n11202), .Z(n11121) );
  NBUFFX2 U10824 ( .INP(n11191), .Z(n11178) );
  NBUFFX2 U10825 ( .INP(n11206), .Z(n11099) );
  NBUFFX2 U10826 ( .INP(n11193), .Z(n11166) );
  NBUFFX2 U10827 ( .INP(n11192), .Z(n11173) );
  NBUFFX2 U10828 ( .INP(n11195), .Z(n11156) );
  NBUFFX2 U10829 ( .INP(n11208), .Z(n11093) );
  NBUFFX2 U10830 ( .INP(n11204), .Z(n11110) );
  NBUFFX2 U10831 ( .INP(n11194), .Z(n11163) );
  NBUFFX2 U10832 ( .INP(n11201), .Z(n11128) );
  NBUFFX2 U10833 ( .INP(n11192), .Z(n11171) );
  NBUFFX2 U10834 ( .INP(n11203), .Z(n11118) );
  NBUFFX2 U10835 ( .INP(n11191), .Z(n11177) );
  NBUFFX2 U10836 ( .INP(n11204), .Z(n11111) );
  NBUFFX2 U10837 ( .INP(n11203), .Z(n11117) );
  NBUFFX2 U10838 ( .INP(n11209), .Z(n11085) );
  NBUFFX2 U10839 ( .INP(n11190), .Z(n11181) );
  NBUFFX2 U10840 ( .INP(n11205), .Z(n11105) );
  NBUFFX2 U10841 ( .INP(n11199), .Z(n11138) );
  NBUFFX2 U10842 ( .INP(n11194), .Z(n11159) );
  NBUFFX2 U10843 ( .INP(n11209), .Z(n11086) );
  NBUFFX2 U10844 ( .INP(n11199), .Z(n11135) );
  NBUFFX2 U10845 ( .INP(n11204), .Z(n11112) );
  NBUFFX2 U10846 ( .INP(n11207), .Z(n11097) );
  NBUFFX2 U10847 ( .INP(n11198), .Z(n11139) );
  NBUFFX2 U10848 ( .INP(n11193), .Z(n11164) );
  NBUFFX2 U10849 ( .INP(n11197), .Z(n11144) );
  NBUFFX2 U10850 ( .INP(n11199), .Z(n11137) );
  NBUFFX2 U10851 ( .INP(n11205), .Z(n11107) );
  NBUFFX2 U10852 ( .INP(n11196), .Z(n11152) );
  NBUFFX2 U10853 ( .INP(n11200), .Z(n11129) );
  NBUFFX2 U10854 ( .INP(n11195), .Z(n11158) );
  NBUFFX2 U10855 ( .INP(n11199), .Z(n11136) );
  NBUFFX2 U10856 ( .INP(n11209), .Z(n11084) );
  NBUFFX2 U10857 ( .INP(n11202), .Z(n11119) );
  NBUFFX2 U10858 ( .INP(n11190), .Z(n11182) );
  NBUFFX2 U10859 ( .INP(n11191), .Z(n11176) );
  NBUFFX2 U10860 ( .INP(n11194), .Z(n11161) );
  NBUFFX2 U10861 ( .INP(n11206), .Z(n11101) );
  NBUFFX2 U10862 ( .INP(n11207), .Z(n11098) );
  NBUFFX2 U10863 ( .INP(n11197), .Z(n11147) );
  NBUFFX2 U10864 ( .INP(n11204), .Z(n11109) );
  NBUFFX2 U10865 ( .INP(n11208), .Z(n11092) );
  NBUFFX2 U10866 ( .INP(n11190), .Z(n11180) );
  NBUFFX2 U10867 ( .INP(n11190), .Z(n11179) );
  NBUFFX2 U10868 ( .INP(n11203), .Z(n11116) );
  NBUFFX2 U10869 ( .INP(n11195), .Z(n11157) );
  NBUFFX2 U10870 ( .INP(n11198), .Z(n11142) );
  NBUFFX2 U10871 ( .INP(n11198), .Z(n11140) );
  NBUFFX2 U10872 ( .INP(n11193), .Z(n11168) );
  NBUFFX2 U10873 ( .INP(n11204), .Z(n11113) );
  NBUFFX2 U10874 ( .INP(n11201), .Z(n11124) );
  NBUFFX2 U10875 ( .INP(n11190), .Z(n11183) );
  NBUFFX2 U10876 ( .INP(n11203), .Z(n11114) );
  NBUFFX2 U10877 ( .INP(n11196), .Z(n11153) );
  NBUFFX2 U10878 ( .INP(n11200), .Z(n11132) );
  NBUFFX2 U10879 ( .INP(n11192), .Z(n11169) );
  NBUFFX2 U10880 ( .INP(n11207), .Z(n11094) );
  NBUFFX2 U10881 ( .INP(n11198), .Z(n11143) );
  NBUFFX2 U10882 ( .INP(n11201), .Z(n11127) );
  NBUFFX2 U10883 ( .INP(n11197), .Z(n11146) );
  NBUFFX2 U10884 ( .INP(n11209), .Z(n11087) );
  NBUFFX2 U10885 ( .INP(n11201), .Z(n11126) );
  NBUFFX2 U10886 ( .INP(n11194), .Z(n11162) );
  NBUFFX2 U10887 ( .INP(n11196), .Z(n11151) );
  NBUFFX2 U10888 ( .INP(n11200), .Z(n11131) );
  NBUFFX2 U10889 ( .INP(n11197), .Z(n11145) );
  NBUFFX2 U10890 ( .INP(n11193), .Z(n11167) );
  NBUFFX2 U10891 ( .INP(n11205), .Z(n11104) );
  NBUFFX2 U10892 ( .INP(n11192), .Z(n11170) );
  NBUFFX2 U10893 ( .INP(n11209), .Z(n11088) );
  NBUFFX2 U10894 ( .INP(n11196), .Z(n11149) );
  NBUFFX2 U10895 ( .INP(n11195), .Z(n11155) );
  NBUFFX2 U10896 ( .INP(n11207), .Z(n11096) );
  NBUFFX2 U10897 ( .INP(n11208), .Z(n11089) );
  NBUFFX2 U10898 ( .INP(n11208), .Z(n11091) );
  NBUFFX2 U10899 ( .INP(n11200), .Z(n11130) );
  NBUFFX2 U10900 ( .INP(n11193), .Z(n11165) );
  NBUFFX2 U10901 ( .INP(n11208), .Z(n11090) );
  NBUFFX2 U10902 ( .INP(n11192), .Z(n11172) );
  NBUFFX2 U10903 ( .INP(n11205), .Z(n11106) );
  NBUFFX2 U10904 ( .INP(n11202), .Z(n11120) );
  NBUFFX2 U10905 ( .INP(n11191), .Z(n11174) );
  NBUFFX2 U10906 ( .INP(n11205), .Z(n11108) );
  NBUFFX2 U10907 ( .INP(n11197), .Z(n11148) );
  NBUFFX2 U10908 ( .INP(n11206), .Z(n11103) );
  NBUFFX2 U10909 ( .INP(n11202), .Z(n11122) );
  NBUFFX2 U10910 ( .INP(n11199), .Z(n11134) );
  NBUFFX2 U10911 ( .INP(n11196), .Z(n11150) );
  NBUFFX2 U10912 ( .INP(n11194), .Z(n11160) );
  NBUFFX2 U10913 ( .INP(n11201), .Z(n11125) );
  NBUFFX2 U10914 ( .INP(n11195), .Z(n11154) );
  NBUFFX2 U10915 ( .INP(n11202), .Z(n11123) );
  NBUFFX2 U10916 ( .INP(n11203), .Z(n11115) );
  NBUFFX2 U10917 ( .INP(n11206), .Z(n11102) );
  NBUFFX2 U10918 ( .INP(n11200), .Z(n11133) );
  NBUFFX2 U10919 ( .INP(n11206), .Z(n11100) );
  NBUFFX2 U10920 ( .INP(n11198), .Z(n11141) );
  NBUFFX2 U10921 ( .INP(n11191), .Z(n11175) );
  NBUFFX2 U10922 ( .INP(n10976), .Z(n10973) );
  NBUFFX2 U10923 ( .INP(n10976), .Z(n10974) );
  NBUFFX2 U10924 ( .INP(n10976), .Z(n10971) );
  NBUFFX2 U10925 ( .INP(n10976), .Z(n10972) );
  NBUFFX2 U10926 ( .INP(n10976), .Z(n10975) );
  NBUFFX2 U10927 ( .INP(n10806), .Z(n10801) );
  NBUFFX2 U10928 ( .INP(n10806), .Z(n10803) );
  NBUFFX2 U10929 ( .INP(n10806), .Z(n10804) );
  NBUFFX2 U10930 ( .INP(n10806), .Z(n10802) );
  NBUFFX2 U10931 ( .INP(n11189), .Z(n11184) );
  NBUFFX2 U10932 ( .INP(n11189), .Z(n11186) );
  NBUFFX2 U10933 ( .INP(n11189), .Z(n11187) );
  NBUFFX2 U10934 ( .INP(n11189), .Z(n11185) );
  NBUFFX2 U10935 ( .INP(n10806), .Z(n10805) );
  NBUFFX2 U10936 ( .INP(n11189), .Z(n11188) );
  INVX0 U10937 ( .INP(g35), .ZN(n11014) );
  NBUFFX2 U10938 ( .INP(n10835), .Z(n10806) );
  NBUFFX2 U10939 ( .INP(n10834), .Z(n10807) );
  NBUFFX2 U10940 ( .INP(n10834), .Z(n10808) );
  NBUFFX2 U10941 ( .INP(n10834), .Z(n10809) );
  NBUFFX2 U10942 ( .INP(n10833), .Z(n10810) );
  NBUFFX2 U10943 ( .INP(n10833), .Z(n10811) );
  NBUFFX2 U10944 ( .INP(n10833), .Z(n10812) );
  NBUFFX2 U10945 ( .INP(n10832), .Z(n10813) );
  NBUFFX2 U10946 ( .INP(n10832), .Z(n10814) );
  NBUFFX2 U10947 ( .INP(n10832), .Z(n10815) );
  NBUFFX2 U10948 ( .INP(n10831), .Z(n10816) );
  NBUFFX2 U10949 ( .INP(n10831), .Z(n10817) );
  NBUFFX2 U10950 ( .INP(n10831), .Z(n10818) );
  NBUFFX2 U10951 ( .INP(n10830), .Z(n10819) );
  NBUFFX2 U10952 ( .INP(n10830), .Z(n10820) );
  NBUFFX2 U10953 ( .INP(n10830), .Z(n10821) );
  NBUFFX2 U10954 ( .INP(n10829), .Z(n10822) );
  NBUFFX2 U10955 ( .INP(n10829), .Z(n10823) );
  NBUFFX2 U10956 ( .INP(n10829), .Z(n10824) );
  NBUFFX2 U10957 ( .INP(n10828), .Z(n10825) );
  NBUFFX2 U10958 ( .INP(n10828), .Z(n10826) );
  NBUFFX2 U10959 ( .INP(n10828), .Z(n10827) );
  NBUFFX2 U10960 ( .INP(n10838), .Z(n10828) );
  NBUFFX2 U10961 ( .INP(n10838), .Z(n10829) );
  NBUFFX2 U10962 ( .INP(n10837), .Z(n10830) );
  NBUFFX2 U10963 ( .INP(n10837), .Z(n10831) );
  NBUFFX2 U10964 ( .INP(n10837), .Z(n10832) );
  NBUFFX2 U10965 ( .INP(n10836), .Z(n10833) );
  NBUFFX2 U10966 ( .INP(n10836), .Z(n10834) );
  NBUFFX2 U10967 ( .INP(n10836), .Z(n10835) );
  NBUFFX2 U10968 ( .INP(test_se), .Z(n10836) );
  NBUFFX2 U10969 ( .INP(test_se), .Z(n10837) );
  NBUFFX2 U10970 ( .INP(test_se), .Z(n10838) );
  NBUFFX2 U10971 ( .INP(n11013), .Z(n10976) );
  NBUFFX2 U10972 ( .INP(n11012), .Z(n10977) );
  NBUFFX2 U10973 ( .INP(n11012), .Z(n10978) );
  NBUFFX2 U10974 ( .INP(n11012), .Z(n10979) );
  NBUFFX2 U10975 ( .INP(n11011), .Z(n10980) );
  NBUFFX2 U10976 ( .INP(n11011), .Z(n10981) );
  NBUFFX2 U10977 ( .INP(n11011), .Z(n10982) );
  NBUFFX2 U10978 ( .INP(n11010), .Z(n10983) );
  NBUFFX2 U10979 ( .INP(n11010), .Z(n10984) );
  NBUFFX2 U10980 ( .INP(n11010), .Z(n10985) );
  NBUFFX2 U10981 ( .INP(n11009), .Z(n10986) );
  NBUFFX2 U10982 ( .INP(n11009), .Z(n10987) );
  NBUFFX2 U10983 ( .INP(n11009), .Z(n10988) );
  NBUFFX2 U10984 ( .INP(n11008), .Z(n10989) );
  NBUFFX2 U10985 ( .INP(n11008), .Z(n10990) );
  NBUFFX2 U10986 ( .INP(n11008), .Z(n10991) );
  NBUFFX2 U10987 ( .INP(n11007), .Z(n10992) );
  NBUFFX2 U10988 ( .INP(n11007), .Z(n10993) );
  NBUFFX2 U10989 ( .INP(n11007), .Z(n10994) );
  NBUFFX2 U10990 ( .INP(n11006), .Z(n10995) );
  NBUFFX2 U10991 ( .INP(n11006), .Z(n10996) );
  NBUFFX2 U10992 ( .INP(n11006), .Z(n10997) );
  NBUFFX2 U10993 ( .INP(n11005), .Z(n10998) );
  NBUFFX2 U10994 ( .INP(n11005), .Z(n10999) );
  NBUFFX2 U10995 ( .INP(n11005), .Z(n11000) );
  NBUFFX2 U10996 ( .INP(n11004), .Z(n11001) );
  NBUFFX2 U10997 ( .INP(n11004), .Z(n11002) );
  NBUFFX2 U10998 ( .INP(n11004), .Z(n11003) );
  NBUFFX2 U10999 ( .INP(g35), .Z(n11004) );
  NBUFFX2 U11000 ( .INP(n11013), .Z(n11005) );
  NBUFFX2 U11001 ( .INP(g35), .Z(n11006) );
  NBUFFX2 U11002 ( .INP(n10975), .Z(n11007) );
  NBUFFX2 U11003 ( .INP(n11013), .Z(n11008) );
  NBUFFX2 U11004 ( .INP(n11003), .Z(n11009) );
  NBUFFX2 U11005 ( .INP(g35), .Z(n11010) );
  NBUFFX2 U11006 ( .INP(n11004), .Z(n11011) );
  NBUFFX2 U11007 ( .INP(n11003), .Z(n11012) );
  NBUFFX2 U11008 ( .INP(n11006), .Z(n11013) );
  INVX0 U11009 ( .INP(n10919), .ZN(n11015) );
  INVX0 U11010 ( .INP(n10919), .ZN(n11016) );
  INVX0 U11011 ( .INP(n10919), .ZN(n11017) );
  INVX0 U11012 ( .INP(n10919), .ZN(n11018) );
  INVX0 U11013 ( .INP(n10919), .ZN(n11019) );
  INVX0 U11014 ( .INP(n10919), .ZN(n11020) );
  INVX0 U11015 ( .INP(n10918), .ZN(n11021) );
  INVX0 U11016 ( .INP(n10918), .ZN(n11022) );
  INVX0 U11017 ( .INP(n10918), .ZN(n11023) );
  INVX0 U11018 ( .INP(n10918), .ZN(n11024) );
  INVX0 U11019 ( .INP(n10918), .ZN(n11025) );
  INVX0 U11020 ( .INP(n10917), .ZN(n11026) );
  INVX0 U11021 ( .INP(n10911), .ZN(n11027) );
  INVX0 U11022 ( .INP(n10908), .ZN(n11028) );
  INVX0 U11023 ( .INP(n10909), .ZN(n11029) );
  INVX0 U11024 ( .INP(n10908), .ZN(n11030) );
  INVX0 U11025 ( .INP(n10910), .ZN(n11031) );
  INVX0 U11026 ( .INP(n10908), .ZN(n11032) );
  INVX0 U11027 ( .INP(n10910), .ZN(n11033) );
  INVX0 U11028 ( .INP(n10909), .ZN(n11034) );
  INVX0 U11029 ( .INP(n10910), .ZN(n11035) );
  INVX0 U11030 ( .INP(n10909), .ZN(n11036) );
  INVX0 U11031 ( .INP(n10910), .ZN(n11037) );
  INVX0 U11032 ( .INP(n10909), .ZN(n11038) );
  INVX0 U11033 ( .INP(n10909), .ZN(n11039) );
  INVX0 U11034 ( .INP(n10910), .ZN(n11040) );
  INVX0 U11035 ( .INP(n10911), .ZN(n11041) );
  INVX0 U11036 ( .INP(n10910), .ZN(n11042) );
  INVX0 U11037 ( .INP(n10911), .ZN(n11043) );
  INVX0 U11038 ( .INP(n10911), .ZN(n11044) );
  INVX0 U11039 ( .INP(n10911), .ZN(n11045) );
  INVX0 U11040 ( .INP(n10912), .ZN(n11046) );
  INVX0 U11041 ( .INP(n10912), .ZN(n11047) );
  INVX0 U11042 ( .INP(n10912), .ZN(n11048) );
  INVX0 U11043 ( .INP(n10917), .ZN(n11049) );
  INVX0 U11044 ( .INP(n10912), .ZN(n11050) );
  INVX0 U11045 ( .INP(n10912), .ZN(n11051) );
  INVX0 U11046 ( .INP(n10912), .ZN(n11052) );
  INVX0 U11047 ( .INP(n10913), .ZN(n11053) );
  INVX0 U11048 ( .INP(n10913), .ZN(n11054) );
  INVX0 U11049 ( .INP(n10913), .ZN(n11055) );
  INVX0 U11050 ( .INP(n10913), .ZN(n11056) );
  INVX0 U11051 ( .INP(n10913), .ZN(n11057) );
  INVX0 U11052 ( .INP(n10913), .ZN(n11058) );
  INVX0 U11053 ( .INP(n10914), .ZN(n11059) );
  INVX0 U11054 ( .INP(n10914), .ZN(n11060) );
  INVX0 U11055 ( .INP(n10914), .ZN(n11061) );
  INVX0 U11056 ( .INP(n10914), .ZN(n11062) );
  INVX0 U11057 ( .INP(n10914), .ZN(n11063) );
  INVX0 U11058 ( .INP(n10914), .ZN(n11064) );
  INVX0 U11059 ( .INP(n10915), .ZN(n11065) );
  INVX0 U11060 ( .INP(n10915), .ZN(n11066) );
  INVX0 U11061 ( .INP(n10915), .ZN(n11067) );
  INVX0 U11062 ( .INP(n10915), .ZN(n11068) );
  INVX0 U11063 ( .INP(n10915), .ZN(n11069) );
  INVX0 U11064 ( .INP(n10915), .ZN(n11070) );
  INVX0 U11065 ( .INP(n10916), .ZN(n11071) );
  INVX0 U11066 ( .INP(n10916), .ZN(n11072) );
  INVX0 U11067 ( .INP(n10916), .ZN(n11073) );
  INVX0 U11068 ( .INP(n10916), .ZN(n11074) );
  INVX0 U11069 ( .INP(n10916), .ZN(n11075) );
  INVX0 U11070 ( .INP(n10916), .ZN(n11076) );
  INVX0 U11071 ( .INP(n10917), .ZN(n11077) );
  INVX0 U11072 ( .INP(n10917), .ZN(n11078) );
  INVX0 U11073 ( .INP(n10917), .ZN(n11079) );
  INVX0 U11074 ( .INP(n10917), .ZN(n11080) );
  INVX0 U11075 ( .INP(n10909), .ZN(n11081) );
  NBUFFX2 U11076 ( .INP(n11218), .Z(n11189) );
  NBUFFX2 U11077 ( .INP(n11217), .Z(n11190) );
  NBUFFX2 U11078 ( .INP(n11217), .Z(n11191) );
  NBUFFX2 U11079 ( .INP(n11217), .Z(n11192) );
  NBUFFX2 U11080 ( .INP(n11216), .Z(n11193) );
  NBUFFX2 U11081 ( .INP(n11216), .Z(n11194) );
  NBUFFX2 U11082 ( .INP(n11216), .Z(n11195) );
  NBUFFX2 U11083 ( .INP(n11215), .Z(n11196) );
  NBUFFX2 U11084 ( .INP(n11215), .Z(n11197) );
  NBUFFX2 U11085 ( .INP(n11215), .Z(n11198) );
  NBUFFX2 U11086 ( .INP(n11214), .Z(n11199) );
  NBUFFX2 U11087 ( .INP(n11214), .Z(n11200) );
  NBUFFX2 U11088 ( .INP(n11214), .Z(n11201) );
  NBUFFX2 U11089 ( .INP(n11213), .Z(n11202) );
  NBUFFX2 U11090 ( .INP(n11213), .Z(n11203) );
  NBUFFX2 U11091 ( .INP(n11213), .Z(n11204) );
  NBUFFX2 U11092 ( .INP(n11212), .Z(n11205) );
  NBUFFX2 U11093 ( .INP(n11212), .Z(n11206) );
  NBUFFX2 U11094 ( .INP(n11212), .Z(n11207) );
  NBUFFX2 U11095 ( .INP(n11211), .Z(n11208) );
  NBUFFX2 U11096 ( .INP(n11211), .Z(n11209) );
  NBUFFX2 U11097 ( .INP(n11211), .Z(n11210) );
  NBUFFX2 U11098 ( .INP(n11221), .Z(n11211) );
  NBUFFX2 U11099 ( .INP(n11221), .Z(n11212) );
  NBUFFX2 U11100 ( .INP(n11220), .Z(n11213) );
  NBUFFX2 U11101 ( .INP(n11220), .Z(n11214) );
  NBUFFX2 U11102 ( .INP(n11220), .Z(n11215) );
  NBUFFX2 U11103 ( .INP(n11219), .Z(n11216) );
  NBUFFX2 U11104 ( .INP(n11219), .Z(n11217) );
  NBUFFX2 U11105 ( .INP(n11219), .Z(n11218) );
  NBUFFX2 U11106 ( .INP(CK), .Z(n11219) );
  NBUFFX2 U11107 ( .INP(CK), .Z(n11220) );
  NBUFFX2 U11108 ( .INP(CK), .Z(n11221) );
  NAND2X0 U11109 ( .IN1(n11222), .IN2(n11223), .QN(n956) );
  NAND2X0 U11110 ( .IN1(n11224), .IN2(g1825), .QN(n11223) );
  NAND2X0 U11111 ( .IN1(n11225), .IN2(n11226), .QN(n11224) );
  NAND2X0 U11112 ( .IN1(n4447), .IN2(n10948), .QN(n11226) );
  NAND2X0 U11113 ( .IN1(n11227), .IN2(g1811), .QN(n11222) );
  INVX0 U11114 ( .INP(n11228), .ZN(n11227) );
  NOR2X0 U11115 ( .IN1(n11229), .IN2(n11022), .QN(n11228) );
  NOR2X0 U11116 ( .IN1(n11230), .IN2(n11231), .QN(n11229) );
  NAND2X0 U11117 ( .IN1(n11232), .IN2(n11233), .QN(n92) );
  NAND2X0 U11118 ( .IN1(n95), .IN2(n10655), .QN(n11233) );
  NAND2X0 U11119 ( .IN1(n11061), .IN2(g278), .QN(n11232) );
  NAND2X0 U11120 ( .IN1(n11234), .IN2(n11235), .QN(n755) );
  NAND2X0 U11121 ( .IN1(n11236), .IN2(g2533), .QN(n11235) );
  NAND2X0 U11122 ( .IN1(n11237), .IN2(g2527), .QN(n11234) );
  NAND2X0 U11123 ( .IN1(n11238), .IN2(n11239), .QN(n643) );
  NAND2X0 U11124 ( .IN1(n11240), .IN2(g2518), .QN(n11239) );
  NAND2X0 U11125 ( .IN1(n11241), .IN2(n11242), .QN(n11240) );
  NAND2X0 U11126 ( .IN1(n4391), .IN2(n10948), .QN(n11242) );
  NAND2X0 U11127 ( .IN1(n11243), .IN2(g2504), .QN(n11238) );
  INVX0 U11128 ( .INP(n11244), .ZN(n11243) );
  NOR2X0 U11129 ( .IN1(n11245), .IN2(n11022), .QN(n11244) );
  NOR2X0 U11130 ( .IN1(n11246), .IN2(n11247), .QN(n11245) );
  NAND2X0 U11131 ( .IN1(n11248), .IN2(n11249), .QN(n623) );
  NAND2X0 U11132 ( .IN1(n11250), .IN2(g5495), .QN(n11249) );
  NAND2X0 U11133 ( .IN1(n11251), .IN2(g5489), .QN(n11248) );
  NAND2X0 U11134 ( .IN1(n11252), .IN2(n11253), .QN(n609) );
  NAND2X0 U11135 ( .IN1(n11254), .IN2(g2384), .QN(n11253) );
  NAND2X0 U11136 ( .IN1(n11255), .IN2(n11256), .QN(n11254) );
  NAND2X0 U11137 ( .IN1(n4402), .IN2(n10948), .QN(n11256) );
  NAND2X0 U11138 ( .IN1(n11257), .IN2(g2370), .QN(n11252) );
  INVX0 U11139 ( .INP(n11258), .ZN(n11257) );
  NOR2X0 U11140 ( .IN1(n11259), .IN2(n11022), .QN(n11258) );
  NOR2X0 U11141 ( .IN1(n11260), .IN2(n11261), .QN(n11259) );
  NAND2X0 U11142 ( .IN1(n11262), .IN2(n11263), .QN(n5961) );
  NOR2X0 U11143 ( .IN1(n11264), .IN2(n11265), .QN(n11263) );
  NOR2X0 U11144 ( .IN1(n11266), .IN2(g5348), .QN(n11265) );
  NOR2X0 U11145 ( .IN1(n10526), .IN2(n11267), .QN(n11264) );
  NOR2X0 U11146 ( .IN1(n11268), .IN2(n11269), .QN(n11262) );
  NOR2X0 U11147 ( .IN1(n11270), .IN2(g5352), .QN(n11269) );
  NOR2X0 U11148 ( .IN1(n10525), .IN2(n11271), .QN(n11268) );
  NAND2X0 U11149 ( .IN1(n11272), .IN2(n11273), .QN(n5960) );
  NOR2X0 U11150 ( .IN1(n11274), .IN2(n11275), .QN(n11273) );
  INVX0 U11151 ( .INP(n11276), .ZN(n11275) );
  NAND2X0 U11152 ( .IN1(n11277), .IN2(n10524), .QN(n11276) );
  NOR2X0 U11153 ( .IN1(n10524), .IN2(n11278), .QN(n11274) );
  NOR2X0 U11154 ( .IN1(n11279), .IN2(n11280), .QN(n11272) );
  INVX0 U11155 ( .INP(n11281), .ZN(n11280) );
  NAND2X0 U11156 ( .IN1(n11282), .IN2(n10523), .QN(n11281) );
  NOR2X0 U11157 ( .IN1(n10523), .IN2(n11283), .QN(n11279) );
  NAND2X0 U11158 ( .IN1(n11284), .IN2(n11285), .QN(n55) );
  NAND2X0 U11159 ( .IN1(n11286), .IN2(g6187), .QN(n11285) );
  INVX0 U11160 ( .INP(n11287), .ZN(n11284) );
  NOR2X0 U11161 ( .IN1(n11286), .IN2(n5667), .QN(n11287) );
  INVX0 U11162 ( .INP(n11288), .ZN(n524) );
  NOR2X0 U11163 ( .IN1(n11289), .IN2(g29279), .QN(n11288) );
  NOR2X0 U11164 ( .IN1(n10182), .IN2(n10884), .QN(n11289) );
  NAND2X0 U11165 ( .IN1(n11290), .IN2(n11291), .QN(n503) );
  NAND2X0 U11166 ( .IN1(n11292), .IN2(g5841), .QN(n11291) );
  INVX0 U11167 ( .INP(n11293), .ZN(n11290) );
  NOR2X0 U11168 ( .IN1(n11292), .IN2(n5663), .QN(n11293) );
  INVX0 U11169 ( .INP(n11294), .ZN(n5) );
  NAND2X0 U11170 ( .IN1(n11295), .IN2(n11296), .QN(n479) );
  NAND2X0 U11171 ( .IN1(n11297), .IN2(g6519), .QN(n11296) );
  NAND2X0 U11172 ( .IN1(n11298), .IN2(g6513), .QN(n11295) );
  INVX0 U11173 ( .INP(n11299), .ZN(n473) );
  NOR2X0 U11174 ( .IN1(n11300), .IN2(g24212), .QN(n11299) );
  NOR2X0 U11175 ( .IN1(n10183), .IN2(n10884), .QN(n11300) );
  NAND2X0 U11176 ( .IN1(n11301), .IN2(n11302), .QN(n466) );
  NAND2X0 U11177 ( .IN1(n11303), .IN2(g2652), .QN(n11302) );
  NAND2X0 U11178 ( .IN1(n11304), .IN2(n11305), .QN(n11303) );
  NAND2X0 U11179 ( .IN1(n4379), .IN2(n10947), .QN(n11305) );
  NAND2X0 U11180 ( .IN1(n11306), .IN2(g2638), .QN(n11301) );
  INVX0 U11181 ( .INP(n11307), .ZN(n11306) );
  NOR2X0 U11182 ( .IN1(n11308), .IN2(n11022), .QN(n11307) );
  NOR2X0 U11183 ( .IN1(n11309), .IN2(n11310), .QN(n11308) );
  NAND2X0 U11184 ( .IN1(n11311), .IN2(n11312), .QN(n450) );
  NAND2X0 U11185 ( .IN1(n11313), .IN2(g1959), .QN(n11312) );
  NAND2X0 U11186 ( .IN1(n11314), .IN2(n11315), .QN(n11313) );
  NAND2X0 U11187 ( .IN1(n4436), .IN2(n10947), .QN(n11315) );
  NAND2X0 U11188 ( .IN1(test_so53), .IN2(n11316), .QN(n11311) );
  INVX0 U11189 ( .INP(n11317), .ZN(n11316) );
  NOR2X0 U11190 ( .IN1(n11318), .IN2(n11022), .QN(n11317) );
  NOR2X0 U11191 ( .IN1(n11319), .IN2(n11320), .QN(n11318) );
  NAND2X0 U11192 ( .IN1(n11321), .IN2(n11322), .QN(n45) );
  NAND2X0 U11193 ( .IN1(n11323), .IN2(g1840), .QN(n11322) );
  NAND2X0 U11194 ( .IN1(n11324), .IN2(g1834), .QN(n11321) );
  NAND2X0 U11195 ( .IN1(n11325), .IN2(g1677), .QN(n4459) );
  NAND2X0 U11196 ( .IN1(n11231), .IN2(g1811), .QN(n4448) );
  NOR2X0 U11197 ( .IN1(n10316), .IN2(n10633), .QN(n11231) );
  NAND2X0 U11198 ( .IN1(n11320), .IN2(test_so53), .QN(n4437) );
  NOR2X0 U11199 ( .IN1(n10322), .IN2(n10627), .QN(n11320) );
  NAND2X0 U11200 ( .IN1(n11326), .IN2(g2236), .QN(n4415) );
  NAND2X0 U11201 ( .IN1(n11261), .IN2(g2370), .QN(n4403) );
  NOR2X0 U11202 ( .IN1(n10318), .IN2(n10630), .QN(n11261) );
  NAND2X0 U11203 ( .IN1(n11247), .IN2(g2504), .QN(n4392) );
  NOR2X0 U11204 ( .IN1(n10323), .IN2(n10635), .QN(n11247) );
  NAND2X0 U11205 ( .IN1(n11310), .IN2(g2638), .QN(n4380) );
  NOR2X0 U11206 ( .IN1(n10324), .IN2(n10628), .QN(n11310) );
  NAND2X0 U11207 ( .IN1(n11327), .IN2(n11328), .QN(n4305) );
  NOR2X0 U11208 ( .IN1(n11329), .IN2(n11330), .QN(n11328) );
  NOR2X0 U11209 ( .IN1(n10527), .IN2(n10173), .QN(n11330) );
  NOR2X0 U11210 ( .IN1(n5712), .IN2(n10172), .QN(n11329) );
  NOR2X0 U11211 ( .IN1(n11331), .IN2(n11332), .QN(n11327) );
  NAND2X0 U11212 ( .IN1(n11333), .IN2(n11334), .QN(n11332) );
  NAND2X0 U11213 ( .IN1(n11335), .IN2(n5440), .QN(n11334) );
  NOR2X0 U11214 ( .IN1(n11336), .IN2(n11337), .QN(n11335) );
  NAND2X0 U11215 ( .IN1(n5712), .IN2(n5656), .QN(n11337) );
  NAND2X0 U11216 ( .IN1(n10527), .IN2(n11338), .QN(n11336) );
  NAND2X0 U11217 ( .IN1(n11339), .IN2(n11340), .QN(n11338) );
  NAND2X0 U11218 ( .IN1(n11341), .IN2(n11342), .QN(n11339) );
  NAND2X0 U11219 ( .IN1(n11343), .IN2(g4776), .QN(n11342) );
  NAND2X0 U11220 ( .IN1(n5368), .IN2(n11344), .QN(n11343) );
  XNOR2X1 U11221 ( .IN1(g34657), .IN2(n11345), .Q(n11344) );
  NOR2X0 U11222 ( .IN1(n11346), .IN2(n11347), .QN(n11345) );
  NAND2X0 U11223 ( .IN1(n11348), .IN2(n11349), .QN(n11347) );
  NAND2X0 U11224 ( .IN1(n11350), .IN2(g4727), .QN(n11349) );
  NAND2X0 U11225 ( .IN1(n11351), .IN2(g4722), .QN(n11348) );
  INVX0 U11226 ( .INP(n11352), .ZN(n11351) );
  INVX0 U11227 ( .INP(n11353), .ZN(n11346) );
  NOR2X0 U11228 ( .IN1(n11354), .IN2(n11355), .QN(n11353) );
  NOR2X0 U11229 ( .IN1(n11356), .IN2(n5296), .QN(n11355) );
  NOR2X0 U11230 ( .IN1(n11357), .IN2(n5344), .QN(n11354) );
  NOR2X0 U11231 ( .IN1(n11358), .IN2(n11359), .QN(n11341) );
  NOR2X0 U11232 ( .IN1(n11360), .IN2(g4793), .QN(n11359) );
  NOR2X0 U11233 ( .IN1(n11361), .IN2(test_so29), .QN(n11360) );
  NOR2X0 U11234 ( .IN1(n11362), .IN2(n11363), .QN(n11361) );
  NAND2X0 U11235 ( .IN1(n5707), .IN2(n11364), .QN(n11363) );
  NAND2X0 U11236 ( .IN1(n5867), .IN2(n11350), .QN(n11364) );
  INVX0 U11237 ( .INP(n11365), .ZN(n11350) );
  NAND2X0 U11238 ( .IN1(n11356), .IN2(n11357), .QN(n11362) );
  NOR2X0 U11239 ( .IN1(n5368), .IN2(g34657), .QN(n11358) );
  NAND2X0 U11240 ( .IN1(n5880), .IN2(g4674), .QN(n11333) );
  NOR2X0 U11241 ( .IN1(n5656), .IN2(g4826), .QN(n11331) );
  NAND2X0 U11242 ( .IN1(n11366), .IN2(n11367), .QN(n4283) );
  NOR2X0 U11243 ( .IN1(n11368), .IN2(n11369), .QN(n11367) );
  NOR2X0 U11244 ( .IN1(n5318), .IN2(g3333), .QN(n11369) );
  NOR2X0 U11245 ( .IN1(n5713), .IN2(n10174), .QN(n11368) );
  NOR2X0 U11246 ( .IN1(n11370), .IN2(n11371), .QN(n11366) );
  NAND2X0 U11247 ( .IN1(n11372), .IN2(n11373), .QN(n11371) );
  NAND2X0 U11248 ( .IN1(n10176), .IN2(g4878), .QN(n11373) );
  NAND2X0 U11249 ( .IN1(n11374), .IN2(n5283), .QN(n11372) );
  NOR2X0 U11250 ( .IN1(n11375), .IN2(n11376), .QN(n11374) );
  NOR2X0 U11251 ( .IN1(n11377), .IN2(n11378), .QN(n11375) );
  NOR2X0 U11252 ( .IN1(n11379), .IN2(n11380), .QN(n11378) );
  NAND2X0 U11253 ( .IN1(n11381), .IN2(n11382), .QN(n11380) );
  NAND2X0 U11254 ( .IN1(n11383), .IN2(g4983), .QN(n11382) );
  INVX0 U11255 ( .INP(g34649), .ZN(n11383) );
  NAND2X0 U11256 ( .IN1(n5367), .IN2(n11384), .QN(n11381) );
  NAND2X0 U11257 ( .IN1(n10652), .IN2(n11385), .QN(n11384) );
  NAND2X0 U11258 ( .IN1(n11386), .IN2(n11387), .QN(n11385) );
  NOR2X0 U11259 ( .IN1(n11388), .IN2(n11389), .QN(n11387) );
  NOR2X0 U11260 ( .IN1(n11390), .IN2(g4966), .QN(n11386) );
  NOR2X0 U11261 ( .IN1(n11391), .IN2(g4927), .QN(n11390) );
  NOR2X0 U11262 ( .IN1(n5706), .IN2(n11392), .QN(n11379) );
  NOR2X0 U11263 ( .IN1(n11393), .IN2(g4983), .QN(n11392) );
  XNOR2X1 U11264 ( .IN1(n11394), .IN2(g34649), .Q(n11393) );
  NAND2X0 U11265 ( .IN1(n11395), .IN2(n11396), .QN(n11394) );
  NOR2X0 U11266 ( .IN1(n11397), .IN2(n11398), .QN(n11396) );
  NOR2X0 U11267 ( .IN1(n5408), .IN2(n11391), .QN(n11398) );
  NOR2X0 U11268 ( .IN1(n5297), .IN2(n11399), .QN(n11397) );
  NOR2X0 U11269 ( .IN1(n11400), .IN2(n11401), .QN(n11395) );
  NOR2X0 U11270 ( .IN1(n5295), .IN2(n11402), .QN(n11401) );
  NOR2X0 U11271 ( .IN1(n5346), .IN2(n11403), .QN(n11400) );
  NOR2X0 U11272 ( .IN1(n5881), .IN2(n5443), .QN(n11370) );
  INVX0 U11273 ( .INP(n11404), .ZN(n4198) );
  NOR2X0 U11274 ( .IN1(g3167), .IN2(n11405), .QN(n4034) );
  NAND2X0 U11275 ( .IN1(n5366), .IN2(n10578), .QN(n11405) );
  NAND2X0 U11276 ( .IN1(n11406), .IN2(n11407), .QN(n403) );
  NAND2X0 U11277 ( .IN1(n11408), .IN2(g2399), .QN(n11407) );
  NAND2X0 U11278 ( .IN1(n11409), .IN2(g2393), .QN(n11406) );
  NOR2X0 U11279 ( .IN1(g3518), .IN2(n11410), .QN(n4002) );
  NAND2X0 U11280 ( .IN1(n5576), .IN2(n10587), .QN(n11410) );
  NOR2X0 U11281 ( .IN1(g3857), .IN2(n11411), .QN(n3969) );
  NAND2X0 U11282 ( .IN1(n10591), .IN2(n10647), .QN(n11411) );
  NOR2X0 U11283 ( .IN1(n11412), .IN2(n11413), .QN(n3933) );
  NAND2X0 U11284 ( .IN1(n2760), .IN2(g43), .QN(n11412) );
  NOR2X0 U11285 ( .IN1(g5176), .IN2(n11414), .QN(n3926) );
  NAND2X0 U11286 ( .IN1(n10586), .IN2(n5570), .QN(n11414) );
  NOR2X0 U11287 ( .IN1(g5523), .IN2(n11415), .QN(n3893) );
  NAND2X0 U11288 ( .IN1(n10589), .IN2(n5575), .QN(n11415) );
  NOR2X0 U11289 ( .IN1(g5869), .IN2(n11416), .QN(n3860) );
  NAND2X0 U11290 ( .IN1(n5573), .IN2(n10590), .QN(n11416) );
  NOR2X0 U11291 ( .IN1(g6215), .IN2(n11417), .QN(n3826) );
  NAND2X0 U11292 ( .IN1(n5574), .IN2(n10588), .QN(n11417) );
  NOR2X0 U11293 ( .IN1(g6561), .IN2(n11418), .QN(n3792) );
  NAND2X0 U11294 ( .IN1(n5571), .IN2(n10592), .QN(n11418) );
  INVX0 U11295 ( .INP(n11419), .ZN(n3743) );
  INVX0 U11296 ( .INP(n11420), .ZN(n3739) );
  INVX0 U11297 ( .INP(n11421), .ZN(n3734) );
  NAND2X0 U11298 ( .IN1(n11422), .IN2(n11423), .QN(n3675) );
  NOR2X0 U11299 ( .IN1(n11424), .IN2(n11425), .QN(n11423) );
  NOR2X0 U11300 ( .IN1(n10272), .IN2(n11426), .QN(n11425) );
  NOR2X0 U11301 ( .IN1(g441), .IN2(n11427), .QN(n11426) );
  XOR2X1 U11302 ( .IN1(test_so72), .IN2(n10404), .Q(n11427) );
  NOR2X0 U11303 ( .IN1(n11428), .IN2(g392), .QN(n11424) );
  NOR2X0 U11304 ( .IN1(g411), .IN2(n11429), .QN(n11428) );
  XOR2X1 U11305 ( .IN1(test_so72), .IN2(n5402), .Q(n11429) );
  NOR2X0 U11306 ( .IN1(g691), .IN2(g417), .QN(n11422) );
  NAND2X0 U11307 ( .IN1(n11430), .IN2(n5516), .QN(n3635) );
  NOR2X0 U11308 ( .IN1(test_so30), .IN2(n5349), .QN(n11430) );
  NOR2X0 U11309 ( .IN1(n11431), .IN2(n11432), .QN(n3174) );
  XOR2X1 U11310 ( .IN1(g482), .IN2(g72), .Q(n11432) );
  XOR2X1 U11311 ( .IN1(n5708), .IN2(n11433), .Q(n11431) );
  INVX0 U11312 ( .INP(n11434), .ZN(n315) );
  INVX0 U11313 ( .INP(n11435), .ZN(n3122) );
  NOR2X0 U11314 ( .IN1(n1770), .IN2(n6010), .QN(n3084) );
  NAND2X0 U11315 ( .IN1(n11436), .IN2(n11437), .QN(n3065) );
  NAND2X0 U11316 ( .IN1(n11438), .IN2(g4108), .QN(n11437) );
  NOR2X0 U11317 ( .IN1(n10403), .IN2(n11022), .QN(n11436) );
  INVX0 U11318 ( .INP(n11439), .ZN(n293) );
  NAND2X0 U11319 ( .IN1(n11440), .IN2(n11441), .QN(n290) );
  NAND2X0 U11320 ( .IN1(n11442), .IN2(g2108), .QN(n11441) );
  NAND2X0 U11321 ( .IN1(n11443), .IN2(g2102), .QN(n11440) );
  INVX0 U11322 ( .INP(n11444), .ZN(n29) );
  NOR2X0 U11323 ( .IN1(n11445), .IN2(n11446), .QN(n11444) );
  NOR2X0 U11324 ( .IN1(n11447), .IN2(n10404), .QN(n11446) );
  NOR2X0 U11325 ( .IN1(n11448), .IN2(n10167), .QN(n11445) );
  NOR2X0 U11326 ( .IN1(n11449), .IN2(n11450), .QN(n268) );
  XOR2X1 U11327 ( .IN1(n5323), .IN2(n2607), .Q(n2608) );
  NAND2X0 U11328 ( .IN1(n11451), .IN2(g34979), .QN(n2461) );
  NAND2X0 U11329 ( .IN1(n11452), .IN2(n11453), .QN(n201) );
  NAND2X0 U11330 ( .IN1(n11454), .IN2(g5827), .QN(n11453) );
  NAND2X0 U11331 ( .IN1(n11455), .IN2(g5821), .QN(n11452) );
  NAND2X0 U11332 ( .IN1(n11456), .IN2(n11457), .QN(n198) );
  NAND2X0 U11333 ( .IN1(n11458), .IN2(g5481), .QN(n11457) );
  NAND2X0 U11334 ( .IN1(n11459), .IN2(g5475), .QN(n11456) );
  NAND2X0 U11335 ( .IN1(n11460), .IN2(n11461), .QN(n176) );
  NAND2X0 U11336 ( .IN1(n11462), .IN2(g3139), .QN(n11461) );
  INVX0 U11337 ( .INP(n11463), .ZN(n11460) );
  NOR2X0 U11338 ( .IN1(n11462), .IN2(n5661), .QN(n11463) );
  NAND2X0 U11339 ( .IN1(n11464), .IN2(n11465), .QN(n1688) );
  INVX0 U11340 ( .INP(g29277), .ZN(n11465) );
  NAND2X0 U11341 ( .IN1(n11073), .IN2(test_so100), .QN(n11464) );
  INVX0 U11342 ( .INP(n11466), .ZN(n1545) );
  NOR2X0 U11343 ( .IN1(n11467), .IN2(g26953), .QN(n11466) );
  NOR2X0 U11344 ( .IN1(n10266), .IN2(n10884), .QN(n11467) );
  NAND2X0 U11345 ( .IN1(n11468), .IN2(n11469), .QN(n15) );
  NAND2X0 U11346 ( .IN1(n11470), .IN2(g1691), .QN(n11469) );
  NAND2X0 U11347 ( .IN1(n11471), .IN2(n11472), .QN(n11470) );
  NAND2X0 U11348 ( .IN1(n4458), .IN2(n10947), .QN(n11472) );
  NAND2X0 U11349 ( .IN1(n11473), .IN2(g1677), .QN(n11468) );
  INVX0 U11350 ( .INP(n11474), .ZN(n11473) );
  NOR2X0 U11351 ( .IN1(n11475), .IN2(n11021), .QN(n11474) );
  NOR2X0 U11352 ( .IN1(n11476), .IN2(n11325), .QN(n11475) );
  NOR2X0 U11353 ( .IN1(n10320), .IN2(n1418), .QN(n11325) );
  NAND2X0 U11354 ( .IN1(n11477), .IN2(g2079), .QN(n1432) );
  INVX0 U11355 ( .INP(n11478), .ZN(n11477) );
  NAND2X0 U11356 ( .IN1(n11479), .IN2(n11480), .QN(n1426) );
  NAND2X0 U11357 ( .IN1(n11481), .IN2(g6533), .QN(n11480) );
  INVX0 U11358 ( .INP(n11482), .ZN(n11479) );
  NOR2X0 U11359 ( .IN1(n11481), .IN2(n5659), .QN(n11482) );
  NAND2X0 U11360 ( .IN1(n11483), .IN2(n11484), .QN(n136) );
  NAND2X0 U11361 ( .IN1(n11485), .IN2(g1974), .QN(n11484) );
  NAND2X0 U11362 ( .IN1(n11486), .IN2(g1968), .QN(n11483) );
  NAND2X0 U11363 ( .IN1(n11487), .IN2(n11488), .QN(n132) );
  NAND2X0 U11364 ( .IN1(n11489), .IN2(g2250), .QN(n11488) );
  NAND2X0 U11365 ( .IN1(n11490), .IN2(n11491), .QN(n11489) );
  NAND2X0 U11366 ( .IN1(n4414), .IN2(n10947), .QN(n11491) );
  NAND2X0 U11367 ( .IN1(n11492), .IN2(g2236), .QN(n11487) );
  INVX0 U11368 ( .INP(n11493), .ZN(n11492) );
  NOR2X0 U11369 ( .IN1(n11494), .IN2(n11021), .QN(n11493) );
  NOR2X0 U11370 ( .IN1(n11495), .IN2(n11326), .QN(n11494) );
  NOR2X0 U11371 ( .IN1(n10314), .IN2(n10636), .QN(n11326) );
  NAND2X0 U11372 ( .IN1(n11496), .IN2(n11497), .QN(n120) );
  NAND2X0 U11373 ( .IN1(n11498), .IN2(g3490), .QN(n11497) );
  INVX0 U11374 ( .INP(n11499), .ZN(n11496) );
  NOR2X0 U11375 ( .IN1(n11498), .IN2(n5668), .QN(n11499) );
  NOR2X0 U11376 ( .IN1(n11500), .IN2(n11413), .QN(n10623) );
  INVX0 U11377 ( .INP(n11501), .ZN(n11500) );
  NOR2X0 U11378 ( .IN1(n11502), .IN2(n11503), .QN(n11501) );
  NOR2X0 U11379 ( .IN1(n11504), .IN2(n5350), .QN(n11503) );
  NOR2X0 U11380 ( .IN1(n11505), .IN2(g4098), .QN(n11502) );
  NOR2X0 U11381 ( .IN1(n11042), .IN2(n10691), .QN(n1052) );
  INVX0 U11382 ( .INP(n11506), .ZN(n103) );
  NAND2X0 U11383 ( .IN1(n11507), .IN2(n11508), .QN(g34980) );
  NAND2X0 U11384 ( .IN1(test_so14), .IN2(n11014), .QN(n11508) );
  NAND2X0 U11385 ( .IN1(n11509), .IN2(n10947), .QN(n11507) );
  NAND2X0 U11386 ( .IN1(n5842), .IN2(n11510), .QN(n11509) );
  NAND2X0 U11387 ( .IN1(n11511), .IN2(n11512), .QN(n11510) );
  NOR2X0 U11388 ( .IN1(g56), .IN2(g54), .QN(n11512) );
  NOR2X0 U11389 ( .IN1(g53), .IN2(n11513), .QN(n11511) );
  NAND2X0 U11390 ( .IN1(n11513), .IN2(g22), .QN(g34972) );
  INVX0 U11391 ( .INP(n35), .ZN(n11513) );
  XOR2X1 U11392 ( .IN1(n11514), .IN2(n11515), .Q(n35) );
  XOR2X1 U11393 ( .IN1(g34978), .IN2(g34977), .Q(n11515) );
  XOR2X1 U11394 ( .IN1(g34970), .IN2(n11516), .Q(n11514) );
  XOR2X1 U11395 ( .IN1(n11517), .IN2(n11518), .Q(n11516) );
  XNOR2X1 U11396 ( .IN1(n11519), .IN2(g34975), .Q(n11518) );
  XNOR2X1 U11397 ( .IN1(g34974), .IN2(g34976), .Q(n11519) );
  XOR2X1 U11398 ( .IN1(g34971), .IN2(n11520), .Q(n11517) );
  XOR2X1 U11399 ( .IN1(n11521), .IN2(g34979), .Q(n11520) );
  NAND2X0 U11400 ( .IN1(n11522), .IN2(g55), .QN(n11521) );
  INVX0 U11401 ( .INP(n11523), .ZN(g34927) );
  NOR2X0 U11402 ( .IN1(g34979), .IN2(n10226), .QN(n11523) );
  NAND2X0 U11403 ( .IN1(n11524), .IN2(n11525), .QN(g34979) );
  NOR2X0 U11404 ( .IN1(n11526), .IN2(n11527), .QN(n11525) );
  NAND2X0 U11405 ( .IN1(n11528), .IN2(n11529), .QN(n11527) );
  NAND2X0 U11406 ( .IN1(n1436), .IN2(n11530), .QN(n11529) );
  NAND2X0 U11407 ( .IN1(n11531), .IN2(n11532), .QN(n11530) );
  NOR2X0 U11408 ( .IN1(n11533), .IN2(n11534), .QN(n11532) );
  NAND2X0 U11409 ( .IN1(n11535), .IN2(n11536), .QN(n11534) );
  NAND2X0 U11410 ( .IN1(n11537), .IN2(g604), .QN(n11536) );
  NOR2X0 U11411 ( .IN1(n11538), .IN2(n11539), .QN(n11535) );
  NOR2X0 U11412 ( .IN1(n11540), .IN2(g23612), .QN(n11539) );
  NOR2X0 U11413 ( .IN1(n5293), .IN2(n11541), .QN(n11538) );
  NAND2X0 U11414 ( .IN1(n11542), .IN2(n11543), .QN(n11533) );
  INVX0 U11415 ( .INP(n11544), .ZN(n11543) );
  NAND2X0 U11416 ( .IN1(n11545), .IN2(n11546), .QN(n11544) );
  NAND2X0 U11417 ( .IN1(g92), .IN2(n11547), .QN(n11546) );
  INVX0 U11418 ( .INP(n11548), .ZN(n11547) );
  NAND2X0 U11419 ( .IN1(g127), .IN2(n11549), .QN(n11545) );
  NAND2X0 U11420 ( .IN1(n11451), .IN2(test_so14), .QN(n11542) );
  NOR2X0 U11421 ( .IN1(n11550), .IN2(n11551), .QN(n11531) );
  NAND2X0 U11422 ( .IN1(n11552), .IN2(n11553), .QN(n11551) );
  NAND2X0 U11423 ( .IN1(n11554), .IN2(g4146), .QN(n11553) );
  NOR2X0 U11424 ( .IN1(n11555), .IN2(n11556), .QN(n11552) );
  NOR2X0 U11425 ( .IN1(n5750), .IN2(n11557), .QN(n11556) );
  NOR2X0 U11426 ( .IN1(n10564), .IN2(n11558), .QN(n11555) );
  NAND2X0 U11427 ( .IN1(n11559), .IN2(n11560), .QN(n11550) );
  NAND2X0 U11428 ( .IN1(n11561), .IN2(g2970), .QN(n11560) );
  NOR2X0 U11429 ( .IN1(n11562), .IN2(n11563), .QN(n11559) );
  NOR2X0 U11430 ( .IN1(n5470), .IN2(n11564), .QN(n11563) );
  NOR2X0 U11431 ( .IN1(n5335), .IN2(n11565), .QN(n11562) );
  NAND2X0 U11432 ( .IN1(n11566), .IN2(g1283), .QN(n11528) );
  NAND2X0 U11433 ( .IN1(n11567), .IN2(n11568), .QN(n11526) );
  NAND2X0 U11434 ( .IN1(test_so67), .IN2(n11569), .QN(n11567) );
  NOR2X0 U11435 ( .IN1(n11570), .IN2(n11571), .QN(n11524) );
  NAND2X0 U11436 ( .IN1(n11572), .IN2(n11573), .QN(n11571) );
  NAND2X0 U11437 ( .IN1(n11574), .IN2(g2138), .QN(n11573) );
  NAND2X0 U11438 ( .IN1(n11575), .IN2(g2697), .QN(n11572) );
  NAND2X0 U11439 ( .IN1(n11576), .IN2(n11577), .QN(n11570) );
  NAND2X0 U11440 ( .IN1(n11578), .IN2(g939), .QN(n11577) );
  NAND2X0 U11441 ( .IN1(n11579), .IN2(n9332), .QN(n11576) );
  INVX0 U11442 ( .INP(n11580), .ZN(g34925) );
  NOR2X0 U11443 ( .IN1(g34978), .IN2(n10226), .QN(n11580) );
  NAND2X0 U11444 ( .IN1(n11581), .IN2(n11582), .QN(g34978) );
  NOR2X0 U11445 ( .IN1(n11583), .IN2(n11584), .QN(n11582) );
  NAND2X0 U11446 ( .IN1(n11585), .IN2(n11586), .QN(n11584) );
  NAND2X0 U11447 ( .IN1(n1436), .IN2(n11587), .QN(n11586) );
  NAND2X0 U11448 ( .IN1(n11588), .IN2(n11589), .QN(n11587) );
  NOR2X0 U11449 ( .IN1(n11590), .IN2(n11591), .QN(n11589) );
  NAND2X0 U11450 ( .IN1(n11592), .IN2(n11593), .QN(n11591) );
  NAND2X0 U11451 ( .IN1(n11594), .IN2(g572), .QN(n11593) );
  NOR2X0 U11452 ( .IN1(n11595), .IN2(n11596), .QN(n11592) );
  NOR2X0 U11453 ( .IN1(n5475), .IN2(n11597), .QN(n11596) );
  NOR2X0 U11454 ( .IN1(n11540), .IN2(g550), .QN(n11595) );
  NAND2X0 U11455 ( .IN1(n11598), .IN2(n11599), .QN(n11590) );
  NAND2X0 U11456 ( .IN1(n11600), .IN2(g790), .QN(n11599) );
  NOR2X0 U11457 ( .IN1(n11601), .IN2(n11602), .QN(n11598) );
  NOR2X0 U11458 ( .IN1(n5488), .IN2(n11603), .QN(n11602) );
  NOR2X0 U11459 ( .IN1(n5342), .IN2(n11548), .QN(n11601) );
  NOR2X0 U11460 ( .IN1(n11604), .IN2(n11605), .QN(n11588) );
  NAND2X0 U11461 ( .IN1(n11606), .IN2(n11607), .QN(n11605) );
  NAND2X0 U11462 ( .IN1(n11608), .IN2(g2965), .QN(n11607) );
  NAND2X0 U11463 ( .IN1(n11554), .IN2(g4176), .QN(n11606) );
  NAND2X0 U11464 ( .IN1(n11609), .IN2(n11610), .QN(n11604) );
  NAND2X0 U11465 ( .IN1(n11611), .IN2(g2878), .QN(n11610) );
  NOR2X0 U11466 ( .IN1(n11612), .IN2(n11613), .QN(n11609) );
  NOR2X0 U11467 ( .IN1(n11614), .IN2(n10660), .QN(n11613) );
  NOR2X0 U11468 ( .IN1(n11564), .IN2(n5471), .QN(n11612) );
  NAND2X0 U11469 ( .IN1(n10093), .IN2(n11566), .QN(n11585) );
  NAND2X0 U11470 ( .IN1(n11615), .IN2(n11568), .QN(n11583) );
  NAND2X0 U11471 ( .IN1(n11569), .IN2(g4253), .QN(n11615) );
  NOR2X0 U11472 ( .IN1(n11616), .IN2(n11617), .QN(n11581) );
  NAND2X0 U11473 ( .IN1(n11618), .IN2(n11619), .QN(n11617) );
  NAND2X0 U11474 ( .IN1(n11574), .IN2(g2130), .QN(n11619) );
  NAND2X0 U11475 ( .IN1(n11575), .IN2(g2689), .QN(n11618) );
  NAND2X0 U11476 ( .IN1(n11620), .IN2(n11621), .QN(n11616) );
  NAND2X0 U11477 ( .IN1(n10094), .IN2(n11578), .QN(n11621) );
  NAND2X0 U11478 ( .IN1(n11579), .IN2(n9276), .QN(n11620) );
  INVX0 U11479 ( .INP(n11622), .ZN(g34923) );
  NOR2X0 U11480 ( .IN1(g34977), .IN2(n10226), .QN(n11622) );
  NAND2X0 U11481 ( .IN1(n11623), .IN2(n11624), .QN(g34977) );
  NOR2X0 U11482 ( .IN1(n11625), .IN2(n11626), .QN(n11624) );
  NAND2X0 U11483 ( .IN1(n11627), .IN2(n11628), .QN(n11626) );
  NAND2X0 U11484 ( .IN1(n1436), .IN2(n11629), .QN(n11628) );
  NAND2X0 U11485 ( .IN1(n11630), .IN2(n11631), .QN(n11629) );
  NOR2X0 U11486 ( .IN1(n11632), .IN2(n11633), .QN(n11631) );
  NAND2X0 U11487 ( .IN1(n11634), .IN2(n11635), .QN(n11633) );
  NAND2X0 U11488 ( .IN1(n11537), .IN2(g613), .QN(n11635) );
  NOR2X0 U11489 ( .IN1(n11636), .IN2(n11637), .QN(n11634) );
  NOR2X0 U11490 ( .IN1(n5490), .IN2(n11540), .QN(n11637) );
  NOR2X0 U11491 ( .IN1(n5291), .IN2(n11541), .QN(n11636) );
  NAND2X0 U11492 ( .IN1(n11638), .IN2(n11639), .QN(n11632) );
  NAND2X0 U11493 ( .IN1(n11549), .IN2(g2868), .QN(n11639) );
  NOR2X0 U11494 ( .IN1(n11640), .IN2(n11641), .QN(n11638) );
  NOR2X0 U11495 ( .IN1(n11548), .IN2(g30327), .QN(n11641) );
  NOR2X0 U11496 ( .IN1(n11642), .IN2(n11643), .QN(n11630) );
  NAND2X0 U11497 ( .IN1(n11644), .IN2(n11645), .QN(n11643) );
  NAND2X0 U11498 ( .IN1(n11554), .IN2(g4172), .QN(n11645) );
  NOR2X0 U11499 ( .IN1(n11646), .IN2(n11647), .QN(n11644) );
  NOR2X0 U11500 ( .IN1(n10232), .IN2(n11557), .QN(n11647) );
  NOR2X0 U11501 ( .IN1(n10616), .IN2(n11558), .QN(n11646) );
  NAND2X0 U11502 ( .IN1(n11648), .IN2(n11649), .QN(n11642) );
  NAND2X0 U11503 ( .IN1(n11561), .IN2(g2950), .QN(n11649) );
  NOR2X0 U11504 ( .IN1(n11650), .IN2(n11651), .QN(n11648) );
  NOR2X0 U11505 ( .IN1(n5331), .IN2(n11564), .QN(n11651) );
  NOR2X0 U11506 ( .IN1(n5336), .IN2(n11565), .QN(n11650) );
  NAND2X0 U11507 ( .IN1(n11652), .IN2(n5879), .QN(n11627) );
  NAND2X0 U11508 ( .IN1(n11653), .IN2(n11568), .QN(n11625) );
  NAND2X0 U11509 ( .IN1(n11569), .IN2(g4300), .QN(n11653) );
  NOR2X0 U11510 ( .IN1(n11654), .IN2(n11655), .QN(n11623) );
  NAND2X0 U11511 ( .IN1(n11656), .IN2(n11657), .QN(n11655) );
  NAND2X0 U11512 ( .IN1(n11579), .IN2(n9245), .QN(n11657) );
  NAND2X0 U11513 ( .IN1(n11658), .IN2(n5867), .QN(n11656) );
  NAND2X0 U11514 ( .IN1(n11659), .IN2(n11660), .QN(n11654) );
  INVX0 U11515 ( .INP(n11661), .ZN(n11660) );
  NOR2X0 U11516 ( .IN1(n11662), .IN2(n2549), .QN(n11661) );
  NAND2X0 U11517 ( .IN1(n11578), .IN2(g947), .QN(n11659) );
  NAND2X0 U11518 ( .IN1(n11663), .IN2(g22), .QN(g34921) );
  INVX0 U11519 ( .INP(g34976), .ZN(n11663) );
  NAND2X0 U11520 ( .IN1(n11664), .IN2(n11665), .QN(g34976) );
  NOR2X0 U11521 ( .IN1(n11666), .IN2(n11667), .QN(n11665) );
  NAND2X0 U11522 ( .IN1(n11668), .IN2(n11669), .QN(n11667) );
  NAND2X0 U11523 ( .IN1(n1436), .IN2(n11670), .QN(n11669) );
  NAND2X0 U11524 ( .IN1(n11671), .IN2(n11672), .QN(n11670) );
  NOR2X0 U11525 ( .IN1(n11673), .IN2(n11674), .QN(n11672) );
  NAND2X0 U11526 ( .IN1(n11675), .IN2(n11676), .QN(n11674) );
  NAND2X0 U11527 ( .IN1(n11594), .IN2(g577), .QN(n11676) );
  NOR2X0 U11528 ( .IN1(n11677), .IN2(n11678), .QN(n11675) );
  NOR2X0 U11529 ( .IN1(n5339), .IN2(n11597), .QN(n11678) );
  NOR2X0 U11530 ( .IN1(n11540), .IN2(n10670), .QN(n11677) );
  NAND2X0 U11531 ( .IN1(n11679), .IN2(n11680), .QN(n11673) );
  NAND2X0 U11532 ( .IN1(n11600), .IN2(g807), .QN(n11680) );
  NOR2X0 U11533 ( .IN1(n11640), .IN2(n11681), .QN(n11679) );
  NOR2X0 U11534 ( .IN1(n10582), .IN2(n11603), .QN(n11681) );
  NOR2X0 U11535 ( .IN1(n11682), .IN2(n11683), .QN(n11671) );
  NAND2X0 U11536 ( .IN1(n11684), .IN2(n11685), .QN(n11683) );
  NAND2X0 U11537 ( .IN1(n11608), .IN2(g2941), .QN(n11685) );
  NAND2X0 U11538 ( .IN1(test_so95), .IN2(n11554), .QN(n11684) );
  NAND2X0 U11539 ( .IN1(n11686), .IN2(n11687), .QN(n11682) );
  NAND2X0 U11540 ( .IN1(n11611), .IN2(g2898), .QN(n11687) );
  NOR2X0 U11541 ( .IN1(n11688), .IN2(n11689), .QN(n11686) );
  NOR2X0 U11542 ( .IN1(n10561), .IN2(n11614), .QN(n11689) );
  NOR2X0 U11543 ( .IN1(n5332), .IN2(n11564), .QN(n11688) );
  NAND2X0 U11544 ( .IN1(n11652), .IN2(g4912), .QN(n11668) );
  NAND2X0 U11545 ( .IN1(n11690), .IN2(n11691), .QN(n11666) );
  NAND2X0 U11546 ( .IN1(n11692), .IN2(g1135), .QN(n11691) );
  NOR2X0 U11547 ( .IN1(n11693), .IN2(n11694), .QN(n11690) );
  NOR2X0 U11548 ( .IN1(n5289), .IN2(n11695), .QN(n11694) );
  NOR2X0 U11549 ( .IN1(n11696), .IN2(n11697), .QN(n11664) );
  NAND2X0 U11550 ( .IN1(n11698), .IN2(n11699), .QN(n11697) );
  NAND2X0 U11551 ( .IN1(n11658), .IN2(g4722), .QN(n11699) );
  NAND2X0 U11552 ( .IN1(n11575), .IN2(g6545), .QN(n11698) );
  NAND2X0 U11553 ( .IN1(n11700), .IN2(n11701), .QN(n11696) );
  NAND2X0 U11554 ( .IN1(n11579), .IN2(n9357), .QN(n11701) );
  NAND2X0 U11555 ( .IN1(n11574), .IN2(g5160), .QN(n11700) );
  NAND2X0 U11556 ( .IN1(n11702), .IN2(g22), .QN(g34919) );
  INVX0 U11557 ( .INP(g34975), .ZN(n11702) );
  NAND2X0 U11558 ( .IN1(n11703), .IN2(n11704), .QN(g34975) );
  NOR2X0 U11559 ( .IN1(n11705), .IN2(n11706), .QN(n11704) );
  NAND2X0 U11560 ( .IN1(n11707), .IN2(n11708), .QN(n11706) );
  NAND2X0 U11561 ( .IN1(n1436), .IN2(n11709), .QN(n11708) );
  NAND2X0 U11562 ( .IN1(n11710), .IN2(n11711), .QN(n11709) );
  NOR2X0 U11563 ( .IN1(n11712), .IN2(n11713), .QN(n11711) );
  NAND2X0 U11564 ( .IN1(n11714), .IN2(n11715), .QN(n11713) );
  NAND2X0 U11565 ( .IN1(n11537), .IN2(g622), .QN(n11715) );
  NAND2X0 U11566 ( .IN1(n11594), .IN2(g582), .QN(n11714) );
  NAND2X0 U11567 ( .IN1(n11716), .IN2(n11717), .QN(n11712) );
  NAND2X0 U11568 ( .IN1(n11718), .IN2(g546), .QN(n11717) );
  INVX0 U11569 ( .INP(n11540), .ZN(n11718) );
  NOR2X0 U11570 ( .IN1(n11719), .IN2(n11720), .QN(n11716) );
  NOR2X0 U11571 ( .IN1(n10212), .IN2(n11541), .QN(n11720) );
  NOR2X0 U11572 ( .IN1(n11603), .IN2(g2994), .QN(n11719) );
  NOR2X0 U11573 ( .IN1(n11721), .IN2(n11722), .QN(n11710) );
  NAND2X0 U11574 ( .IN1(n11723), .IN2(n11724), .QN(n11722) );
  NAND2X0 U11575 ( .IN1(n11608), .IN2(g2927), .QN(n11724) );
  NAND2X0 U11576 ( .IN1(n11554), .IN2(g2860), .QN(n11723) );
  NAND2X0 U11577 ( .IN1(n11725), .IN2(n11726), .QN(n11721) );
  NAND2X0 U11578 ( .IN1(n11611), .IN2(g2864), .QN(n11726) );
  NOR2X0 U11579 ( .IN1(n11727), .IN2(n11728), .QN(n11725) );
  NOR2X0 U11580 ( .IN1(n10559), .IN2(n11614), .QN(n11728) );
  NOR2X0 U11581 ( .IN1(n5333), .IN2(n11564), .QN(n11727) );
  NAND2X0 U11582 ( .IN1(n11652), .IN2(g4907), .QN(n11707) );
  NAND2X0 U11583 ( .IN1(n11729), .IN2(n11730), .QN(n11705) );
  NAND2X0 U11584 ( .IN1(n11692), .IN2(g1105), .QN(n11730) );
  NOR2X0 U11585 ( .IN1(n11693), .IN2(n11731), .QN(n11729) );
  NOR2X0 U11586 ( .IN1(n5343), .IN2(n11695), .QN(n11731) );
  INVX0 U11587 ( .INP(n11568), .ZN(n11693) );
  NOR2X0 U11588 ( .IN1(n11732), .IN2(n11733), .QN(n11703) );
  NAND2X0 U11589 ( .IN1(n11734), .IN2(n11735), .QN(n11733) );
  NAND2X0 U11590 ( .IN1(n11658), .IN2(g4717), .QN(n11735) );
  NAND2X0 U11591 ( .IN1(n11575), .IN2(g3151), .QN(n11734) );
  NAND2X0 U11592 ( .IN1(n11736), .IN2(n11737), .QN(n11732) );
  NAND2X0 U11593 ( .IN1(n11579), .IN2(n9294), .QN(n11737) );
  NAND2X0 U11594 ( .IN1(n11574), .IN2(g5507), .QN(n11736) );
  INVX0 U11595 ( .INP(n11738), .ZN(g34917) );
  NOR2X0 U11596 ( .IN1(g34974), .IN2(n10226), .QN(n11738) );
  NAND2X0 U11597 ( .IN1(n11739), .IN2(n11740), .QN(g34974) );
  NOR2X0 U11598 ( .IN1(n11741), .IN2(n11742), .QN(n11740) );
  NAND2X0 U11599 ( .IN1(n11743), .IN2(n11744), .QN(n11742) );
  NAND2X0 U11600 ( .IN1(n1436), .IN2(n11745), .QN(n11744) );
  NAND2X0 U11601 ( .IN1(n11746), .IN2(n11747), .QN(n11745) );
  NOR2X0 U11602 ( .IN1(n11748), .IN2(n11749), .QN(n11747) );
  NAND2X0 U11603 ( .IN1(n11750), .IN2(n11751), .QN(n11749) );
  NAND2X0 U11604 ( .IN1(n11594), .IN2(g590), .QN(n11751) );
  NAND2X0 U11605 ( .IN1(n11752), .IN2(g772), .QN(n11750) );
  NAND2X0 U11606 ( .IN1(n11753), .IN2(n11754), .QN(n11748) );
  NAND2X0 U11607 ( .IN1(n11537), .IN2(g626), .QN(n11754) );
  NOR2X0 U11608 ( .IN1(n11755), .IN2(n11756), .QN(n11753) );
  NOR2X0 U11609 ( .IN1(n10569), .IN2(n11603), .QN(n11756) );
  NOR2X0 U11610 ( .IN1(n11757), .IN2(n11758), .QN(n11746) );
  NAND2X0 U11611 ( .IN1(n11759), .IN2(n11760), .QN(n11758) );
  NAND2X0 U11612 ( .IN1(n11608), .IN2(g2917), .QN(n11760) );
  NAND2X0 U11613 ( .IN1(n11554), .IN2(g2852), .QN(n11759) );
  NAND2X0 U11614 ( .IN1(n11761), .IN2(n11762), .QN(n11757) );
  NAND2X0 U11615 ( .IN1(n11561), .IN2(g2912), .QN(n11762) );
  NAND2X0 U11616 ( .IN1(n11611), .IN2(g2856), .QN(n11761) );
  NAND2X0 U11617 ( .IN1(n11652), .IN2(g4922), .QN(n11743) );
  NAND2X0 U11618 ( .IN1(n11763), .IN2(n11764), .QN(n11741) );
  NAND2X0 U11619 ( .IN1(n11765), .IN2(g1472), .QN(n11764) );
  NAND2X0 U11620 ( .IN1(n11692), .IN2(g1129), .QN(n11763) );
  NOR2X0 U11621 ( .IN1(n11766), .IN2(n11767), .QN(n11739) );
  NAND2X0 U11622 ( .IN1(n11768), .IN2(n11769), .QN(n11767) );
  NAND2X0 U11623 ( .IN1(n11658), .IN2(g4732), .QN(n11769) );
  NAND2X0 U11624 ( .IN1(test_so45), .IN2(n11575), .QN(n11768) );
  NAND2X0 U11625 ( .IN1(n11770), .IN2(n11771), .QN(n11766) );
  NAND2X0 U11626 ( .IN1(n11579), .IN2(n9327), .QN(n11771) );
  NAND2X0 U11627 ( .IN1(n11574), .IN2(g5853), .QN(n11770) );
  NAND2X0 U11628 ( .IN1(n11449), .IN2(g22), .QN(g34915) );
  INVX0 U11629 ( .INP(g34971), .ZN(n11449) );
  NAND2X0 U11630 ( .IN1(n11772), .IN2(n11773), .QN(g34971) );
  NOR2X0 U11631 ( .IN1(n11774), .IN2(n11775), .QN(n11773) );
  NAND2X0 U11632 ( .IN1(n11776), .IN2(n11777), .QN(n11775) );
  NAND2X0 U11633 ( .IN1(n1436), .IN2(n11778), .QN(n11777) );
  NAND2X0 U11634 ( .IN1(n11779), .IN2(n11780), .QN(n11778) );
  NOR2X0 U11635 ( .IN1(n11781), .IN2(n11782), .QN(n11780) );
  NAND2X0 U11636 ( .IN1(n11783), .IN2(n11784), .QN(n11782) );
  NAND2X0 U11637 ( .IN1(n11451), .IN2(g2984), .QN(n11784) );
  INVX0 U11638 ( .INP(n11450), .ZN(n11451) );
  NAND2X0 U11639 ( .IN1(n11785), .IN2(n11786), .QN(n11450) );
  NOR2X0 U11640 ( .IN1(g28), .IN2(n11787), .QN(n11785) );
  NAND2X0 U11641 ( .IN1(n11600), .IN2(g781), .QN(n11783) );
  NAND2X0 U11642 ( .IN1(n11788), .IN2(n11789), .QN(n11781) );
  NAND2X0 U11643 ( .IN1(n11549), .IN2(g2890), .QN(n11789) );
  INVX0 U11644 ( .INP(n11603), .ZN(n11549) );
  NAND2X0 U11645 ( .IN1(n11790), .IN2(n11791), .QN(n11603) );
  INVX0 U11646 ( .INP(n11792), .ZN(n11791) );
  NOR2X0 U11647 ( .IN1(n11640), .IN2(n11793), .QN(n11788) );
  NOR2X0 U11648 ( .IN1(n11548), .IN2(n11794), .QN(n11793) );
  INVX0 U11649 ( .INP(g100), .ZN(n11794) );
  NAND2X0 U11650 ( .IN1(n11795), .IN2(n11796), .QN(n11548) );
  NOR2X0 U11651 ( .IN1(n5324), .IN2(n11787), .QN(n11796) );
  NOR2X0 U11652 ( .IN1(g9), .IN2(n11797), .QN(n11795) );
  NOR2X0 U11653 ( .IN1(n11798), .IN2(n11799), .QN(n11640) );
  NAND2X0 U11654 ( .IN1(n5477), .IN2(g28), .QN(n11799) );
  NAND2X0 U11655 ( .IN1(g19), .IN2(n11786), .QN(n11798) );
  NOR2X0 U11656 ( .IN1(n11800), .IN2(n11801), .QN(n11779) );
  NAND2X0 U11657 ( .IN1(n11802), .IN2(n11803), .QN(n11801) );
  NAND2X0 U11658 ( .IN1(n11752), .IN2(test_so60), .QN(n11803) );
  NAND2X0 U11659 ( .IN1(n11554), .IN2(g4157), .QN(n11802) );
  NAND2X0 U11660 ( .IN1(n11804), .IN2(n11805), .QN(n11800) );
  NAND2X0 U11661 ( .IN1(n11594), .IN2(g562), .QN(n11805) );
  NOR2X0 U11662 ( .IN1(n11806), .IN2(n11807), .QN(n11804) );
  NOR2X0 U11663 ( .IN1(n5550), .IN2(n11597), .QN(n11807) );
  NOR2X0 U11664 ( .IN1(n10572), .IN2(n11540), .QN(n11806) );
  NAND2X0 U11665 ( .IN1(test_so64), .IN2(n11566), .QN(n11776) );
  NAND2X0 U11666 ( .IN1(n11808), .IN2(n11568), .QN(n11774) );
  NAND2X0 U11667 ( .IN1(n11809), .IN2(n1436), .QN(n11568) );
  NOR2X0 U11668 ( .IN1(n10906), .IN2(n11810), .QN(n11809) );
  NOR2X0 U11669 ( .IN1(n11600), .IN2(n11811), .QN(n11810) );
  INVX0 U11670 ( .INP(n11541), .ZN(n11600) );
  NAND2X0 U11671 ( .IN1(n11812), .IN2(n11813), .QN(n11541) );
  NOR2X0 U11672 ( .IN1(g9), .IN2(n11792), .QN(n11812) );
  NAND2X0 U11673 ( .IN1(n11569), .IN2(g4245), .QN(n11808) );
  NOR2X0 U11674 ( .IN1(n11814), .IN2(n11792), .QN(n11569) );
  NOR2X0 U11675 ( .IN1(n11815), .IN2(n11816), .QN(n11772) );
  NAND2X0 U11676 ( .IN1(n11817), .IN2(n11818), .QN(n11816) );
  NAND2X0 U11677 ( .IN1(n11574), .IN2(g2145), .QN(n11818) );
  NAND2X0 U11678 ( .IN1(n11575), .IN2(g2704), .QN(n11817) );
  NAND2X0 U11679 ( .IN1(n11819), .IN2(n11820), .QN(n11815) );
  NAND2X0 U11680 ( .IN1(n11578), .IN2(n9247), .QN(n11820) );
  INVX0 U11681 ( .INP(n11821), .ZN(n11578) );
  NAND2X0 U11682 ( .IN1(n11579), .IN2(n9351), .QN(n11819) );
  INVX0 U11683 ( .INP(n11822), .ZN(g34913) );
  NOR2X0 U11684 ( .IN1(g34970), .IN2(n10226), .QN(n11822) );
  NAND2X0 U11685 ( .IN1(n11823), .IN2(n11824), .QN(g34970) );
  NOR2X0 U11686 ( .IN1(n11825), .IN2(n11826), .QN(n11824) );
  NAND2X0 U11687 ( .IN1(n11827), .IN2(n11828), .QN(n11826) );
  NAND2X0 U11688 ( .IN1(n1436), .IN2(n11829), .QN(n11828) );
  NAND2X0 U11689 ( .IN1(n11830), .IN2(n11831), .QN(n11829) );
  NOR2X0 U11690 ( .IN1(n11832), .IN2(n11833), .QN(n11831) );
  NAND2X0 U11691 ( .IN1(n11834), .IN2(n11835), .QN(n11833) );
  NAND2X0 U11692 ( .IN1(n11594), .IN2(g595), .QN(n11835) );
  NAND2X0 U11693 ( .IN1(n11752), .IN2(g776), .QN(n11834) );
  NAND2X0 U11694 ( .IN1(n11836), .IN2(n11837), .QN(n11832) );
  NAND2X0 U11695 ( .IN1(n11537), .IN2(n9340), .QN(n11837) );
  NOR2X0 U11696 ( .IN1(n11755), .IN2(n11838), .QN(n11836) );
  NOR2X0 U11697 ( .IN1(n5491), .IN2(n11540), .QN(n11838) );
  NAND2X0 U11698 ( .IN1(n11839), .IN2(n11813), .QN(n11540) );
  NOR2X0 U11699 ( .IN1(n11840), .IN2(g9), .QN(n11839) );
  NOR2X0 U11700 ( .IN1(n10906), .IN2(n11841), .QN(n11755) );
  INVX0 U11701 ( .INP(n11811), .ZN(n11841) );
  NAND2X0 U11702 ( .IN1(n11842), .IN2(n11565), .QN(n11811) );
  INVX0 U11703 ( .INP(n11594), .ZN(n11565) );
  NOR2X0 U11704 ( .IN1(n11843), .IN2(n11797), .QN(n11594) );
  NAND2X0 U11705 ( .IN1(n5324), .IN2(n2552), .QN(n11843) );
  NOR2X0 U11706 ( .IN1(n11537), .IN2(n11752), .QN(n11842) );
  INVX0 U11707 ( .INP(n11564), .ZN(n11752) );
  NAND2X0 U11708 ( .IN1(n11844), .IN2(n11845), .QN(n11564) );
  NOR2X0 U11709 ( .IN1(n5324), .IN2(g9), .QN(n11845) );
  NOR2X0 U11710 ( .IN1(n11846), .IN2(n11797), .QN(n11844) );
  INVX0 U11711 ( .INP(n11597), .ZN(n11537) );
  NAND2X0 U11712 ( .IN1(n2552), .IN2(n11847), .QN(n11597) );
  NOR2X0 U11713 ( .IN1(n11848), .IN2(n11849), .QN(n11830) );
  NAND2X0 U11714 ( .IN1(n11850), .IN2(n11851), .QN(n11849) );
  NAND2X0 U11715 ( .IN1(n11608), .IN2(g2902), .QN(n11851) );
  INVX0 U11716 ( .INP(n11557), .ZN(n11608) );
  NAND2X0 U11717 ( .IN1(n11852), .IN2(n11786), .QN(n11557) );
  NOR2X0 U11718 ( .IN1(g28), .IN2(n11846), .QN(n11852) );
  NAND2X0 U11719 ( .IN1(n11554), .IN2(g2844), .QN(n11850) );
  NOR2X0 U11720 ( .IN1(n11853), .IN2(n11846), .QN(n11554) );
  NAND2X0 U11721 ( .IN1(g9), .IN2(n11847), .QN(n11853) );
  INVX0 U11722 ( .INP(n11840), .ZN(n11847) );
  NAND2X0 U11723 ( .IN1(n11854), .IN2(n11855), .QN(n11848) );
  NAND2X0 U11724 ( .IN1(test_so1), .IN2(n11561), .QN(n11855) );
  INVX0 U11725 ( .INP(n11614), .ZN(n11561) );
  NAND2X0 U11726 ( .IN1(n11856), .IN2(n11786), .QN(n11614) );
  NOR2X0 U11727 ( .IN1(n11857), .IN2(n11858), .QN(n11786) );
  NAND2X0 U11728 ( .IN1(g9), .IN2(g8), .QN(n11858) );
  NAND2X0 U11729 ( .IN1(n3395), .IN2(test_so85), .QN(n11857) );
  NOR2X0 U11730 ( .IN1(n5324), .IN2(n11846), .QN(n11856) );
  NAND2X0 U11731 ( .IN1(n11611), .IN2(g2848), .QN(n11854) );
  INVX0 U11732 ( .INP(n11558), .ZN(n11611) );
  NAND2X0 U11733 ( .IN1(n11859), .IN2(n11813), .QN(n11558) );
  INVX0 U11734 ( .INP(n11846), .ZN(n11813) );
  NAND2X0 U11735 ( .IN1(n10097), .IN2(n5477), .QN(n11846) );
  NOR2X0 U11736 ( .IN1(n5468), .IN2(n11792), .QN(n11859) );
  NAND2X0 U11737 ( .IN1(n11652), .IN2(g4917), .QN(n11827) );
  INVX0 U11738 ( .INP(n11860), .ZN(n11652) );
  NAND2X0 U11739 ( .IN1(n11861), .IN2(n2527), .QN(n11860) );
  NAND2X0 U11740 ( .IN1(n11862), .IN2(n11863), .QN(n11825) );
  NAND2X0 U11741 ( .IN1(n11765), .IN2(g1300), .QN(n11863) );
  INVX0 U11742 ( .INP(n11695), .ZN(n11765) );
  NAND2X0 U11743 ( .IN1(n11566), .IN2(n2549), .QN(n11695) );
  INVX0 U11744 ( .INP(n11662), .ZN(n11566) );
  NAND2X0 U11745 ( .IN1(n11790), .IN2(n11864), .QN(n11662) );
  NOR2X0 U11746 ( .IN1(n11787), .IN2(g9), .QN(n11790) );
  NAND2X0 U11747 ( .IN1(test_so25), .IN2(n10097), .QN(n11787) );
  NAND2X0 U11748 ( .IN1(n11692), .IN2(g956), .QN(n11862) );
  NOR2X0 U11749 ( .IN1(n11821), .IN2(g947), .QN(n11692) );
  NAND2X0 U11750 ( .IN1(n11861), .IN2(n2552), .QN(n11821) );
  NOR2X0 U11751 ( .IN1(n11865), .IN2(n11792), .QN(n11861) );
  NAND2X0 U11752 ( .IN1(n11866), .IN2(g28), .QN(n11792) );
  NOR2X0 U11753 ( .IN1(n11867), .IN2(n11868), .QN(n11823) );
  NAND2X0 U11754 ( .IN1(n11869), .IN2(n11870), .QN(n11868) );
  NAND2X0 U11755 ( .IN1(n11658), .IN2(g4727), .QN(n11870) );
  INVX0 U11756 ( .INP(n11871), .ZN(n11658) );
  NAND2X0 U11757 ( .IN1(n11864), .IN2(n2527), .QN(n11871) );
  NOR2X0 U11758 ( .IN1(n11840), .IN2(n11865), .QN(n11864) );
  NAND2X0 U11759 ( .IN1(n11575), .IN2(g3853), .QN(n11869) );
  NOR2X0 U11760 ( .IN1(n11872), .IN2(n11814), .QN(n11575) );
  NAND2X0 U11761 ( .IN1(n5324), .IN2(n11873), .QN(n11872) );
  INVX0 U11762 ( .INP(n11797), .ZN(n11873) );
  NAND2X0 U11763 ( .IN1(n11874), .IN2(n11875), .QN(n11797) );
  NOR2X0 U11764 ( .IN1(test_so85), .IN2(n5469), .QN(n11875) );
  NOR2X0 U11765 ( .IN1(g6), .IN2(g8), .QN(n11874) );
  NAND2X0 U11766 ( .IN1(n11876), .IN2(n11877), .QN(n11867) );
  NAND2X0 U11767 ( .IN1(n11579), .IN2(n9322), .QN(n11877) );
  NOR2X0 U11768 ( .IN1(n1436), .IN2(g53), .QN(n11579) );
  INVX0 U11769 ( .INP(n11865), .ZN(n1436) );
  NAND2X0 U11770 ( .IN1(n11574), .IN2(g6199), .QN(n11876) );
  NOR2X0 U11771 ( .IN1(n11814), .IN2(n11840), .QN(n11574) );
  NAND2X0 U11772 ( .IN1(n5324), .IN2(n11866), .QN(n11840) );
  NOR2X0 U11773 ( .IN1(n11878), .IN2(n11879), .QN(n11866) );
  INVX0 U11774 ( .INP(n11880), .ZN(n11879) );
  NOR2X0 U11775 ( .IN1(test_so85), .IN2(g6), .QN(n11880) );
  NAND2X0 U11776 ( .IN1(n10178), .IN2(n5469), .QN(n11878) );
  NAND2X0 U11777 ( .IN1(n11881), .IN2(n11882), .QN(n11814) );
  NOR2X0 U11778 ( .IN1(test_so25), .IN2(n5468), .QN(n11882) );
  NOR2X0 U11779 ( .IN1(n10097), .IN2(n11865), .QN(n11881) );
  NAND2X0 U11780 ( .IN1(n11883), .IN2(n11884), .QN(n11865) );
  NOR2X0 U11781 ( .IN1(test_so74), .IN2(g57), .QN(n11884) );
  NOR2X0 U11782 ( .IN1(g53), .IN2(n11522), .QN(n11883) );
  NAND2X0 U11783 ( .IN1(g54), .IN2(n11885), .QN(n11522) );
  INVX0 U11784 ( .INP(g56), .ZN(n11885) );
  NAND2X0 U11785 ( .IN1(n11886), .IN2(n11887), .QN(g34911) );
  NAND2X0 U11786 ( .IN1(n11888), .IN2(g807), .QN(n11887) );
  NAND2X0 U11787 ( .IN1(n10920), .IN2(n11889), .QN(n11888) );
  NAND2X0 U11788 ( .IN1(n2404), .IN2(g554), .QN(n11886) );
  NAND2X0 U11789 ( .IN1(n11890), .IN2(n11891), .QN(g34882) );
  NAND2X0 U11790 ( .IN1(n11073), .IN2(g4366), .QN(n11891) );
  NAND2X0 U11791 ( .IN1(n11892), .IN2(n10946), .QN(n11890) );
  NAND2X0 U11792 ( .IN1(n11893), .IN2(n11894), .QN(n11892) );
  NAND2X0 U11793 ( .IN1(n11895), .IN2(n11896), .QN(n11894) );
  NOR2X0 U11794 ( .IN1(n11897), .IN2(g4340), .QN(n11895) );
  NOR2X0 U11795 ( .IN1(g4358), .IN2(n11898), .QN(n11897) );
  NOR2X0 U11796 ( .IN1(n11899), .IN2(n11900), .QN(n11893) );
  NOR2X0 U11797 ( .IN1(g4358), .IN2(n11901), .QN(n11900) );
  NAND2X0 U11798 ( .IN1(n11898), .IN2(n10643), .QN(n11901) );
  NAND2X0 U11799 ( .IN1(n11902), .IN2(n11903), .QN(n11898) );
  NOR2X0 U11800 ( .IN1(n11904), .IN2(n11905), .QN(n11903) );
  NOR2X0 U11801 ( .IN1(n5540), .IN2(n11906), .QN(n11905) );
  NAND2X0 U11802 ( .IN1(n5506), .IN2(g4311), .QN(n11906) );
  NOR2X0 U11803 ( .IN1(n11907), .IN2(g4332), .QN(n11904) );
  NOR2X0 U11804 ( .IN1(n11908), .IN2(n11909), .QN(n11907) );
  NAND2X0 U11805 ( .IN1(n11910), .IN2(n11911), .QN(n11909) );
  NAND2X0 U11806 ( .IN1(n10533), .IN2(g4322), .QN(n11911) );
  NAND2X0 U11807 ( .IN1(n11912), .IN2(n5506), .QN(n11910) );
  INVX0 U11808 ( .INP(n11913), .ZN(n11912) );
  NAND2X0 U11809 ( .IN1(n5634), .IN2(g90), .QN(n11913) );
  NOR2X0 U11810 ( .IN1(test_so81), .IN2(g4340), .QN(n11902) );
  NOR2X0 U11811 ( .IN1(n5348), .IN2(n11914), .QN(n11899) );
  NAND2X0 U11812 ( .IN1(test_so81), .IN2(g4340), .QN(n11914) );
  NAND2X0 U11813 ( .IN1(n11915), .IN2(n11916), .QN(g34881) );
  NAND2X0 U11814 ( .IN1(n11073), .IN2(g794), .QN(n11916) );
  NOR2X0 U11815 ( .IN1(n11917), .IN2(n11918), .QN(n11915) );
  NOR2X0 U11816 ( .IN1(g807), .IN2(n11889), .QN(n11918) );
  NOR2X0 U11817 ( .IN1(n5479), .IN2(n11919), .QN(n11917) );
  NAND2X0 U11818 ( .IN1(n2404), .IN2(n11889), .QN(n11919) );
  INVX0 U11819 ( .INP(n2405), .ZN(n11889) );
  NAND2X0 U11820 ( .IN1(n11920), .IN2(n11921), .QN(g34880) );
  NAND2X0 U11821 ( .IN1(n11073), .IN2(g626), .QN(n11921) );
  NOR2X0 U11822 ( .IN1(n11922), .IN2(n11923), .QN(n11920) );
  NOR2X0 U11823 ( .IN1(n9340), .IN2(n11924), .QN(n11923) );
  NOR2X0 U11824 ( .IN1(n19409), .IN2(n11925), .QN(n11922) );
  NAND2X0 U11825 ( .IN1(n2421), .IN2(n11924), .QN(n11925) );
  INVX0 U11826 ( .INP(n2422), .ZN(n11924) );
  NAND2X0 U11827 ( .IN1(n11926), .IN2(n11927), .QN(g34850) );
  NAND2X0 U11828 ( .IN1(n11073), .IN2(g790), .QN(n11927) );
  NOR2X0 U11829 ( .IN1(n11928), .IN2(n11929), .QN(n11926) );
  NOR2X0 U11830 ( .IN1(g794), .IN2(n11930), .QN(n11929) );
  NOR2X0 U11831 ( .IN1(n5291), .IN2(n11931), .QN(n11928) );
  NAND2X0 U11832 ( .IN1(n2404), .IN2(n11930), .QN(n11931) );
  INVX0 U11833 ( .INP(n2419), .ZN(n11930) );
  NAND2X0 U11834 ( .IN1(n11932), .IN2(n11933), .QN(g34849) );
  NAND2X0 U11835 ( .IN1(n11073), .IN2(g622), .QN(n11933) );
  NOR2X0 U11836 ( .IN1(n11934), .IN2(n11935), .QN(n11932) );
  NOR2X0 U11837 ( .IN1(g626), .IN2(n11936), .QN(n11935) );
  NOR2X0 U11838 ( .IN1(n5288), .IN2(n11937), .QN(n11934) );
  NAND2X0 U11839 ( .IN1(n2421), .IN2(n11936), .QN(n11937) );
  INVX0 U11840 ( .INP(n2423), .ZN(n11936) );
  NOR2X0 U11841 ( .IN1(n10401), .IN2(n11938), .QN(g34839) );
  NOR2X0 U11842 ( .IN1(g4366), .IN2(n11939), .QN(n11938) );
  NAND2X0 U11843 ( .IN1(n11940), .IN2(n11941), .QN(n11939) );
  NAND2X0 U11844 ( .IN1(n11942), .IN2(g4332), .QN(n11941) );
  NAND2X0 U11845 ( .IN1(n11943), .IN2(g73), .QN(n11942) );
  NOR2X0 U11846 ( .IN1(n11944), .IN2(g4311), .QN(n11943) );
  NAND2X0 U11847 ( .IN1(n5540), .IN2(n11945), .QN(n11940) );
  NAND2X0 U11848 ( .IN1(n11946), .IN2(n5323), .QN(n11945) );
  NOR2X0 U11849 ( .IN1(g73), .IN2(n11944), .QN(n11946) );
  INVX0 U11850 ( .INP(n11947), .ZN(g34808) );
  NOR2X0 U11851 ( .IN1(n11948), .IN2(n11949), .QN(n11947) );
  NOR2X0 U11852 ( .IN1(n10904), .IN2(n10232), .QN(n11949) );
  NOR2X0 U11853 ( .IN1(n11950), .IN2(n11021), .QN(n11948) );
  NOR2X0 U11854 ( .IN1(n11951), .IN2(g2965), .QN(n11950) );
  NAND2X0 U11855 ( .IN1(n11952), .IN2(g91), .QN(n11951) );
  NAND2X0 U11856 ( .IN1(n11953), .IN2(n11954), .QN(g34807) );
  NAND2X0 U11857 ( .IN1(n11073), .IN2(g2941), .QN(n11954) );
  NAND2X0 U11858 ( .IN1(n11955), .IN2(n10946), .QN(n11953) );
  NAND2X0 U11859 ( .IN1(n11956), .IN2(n11957), .QN(n11955) );
  NOR2X0 U11860 ( .IN1(n11958), .IN2(n11959), .QN(n11957) );
  INVX0 U11861 ( .INP(n11960), .ZN(n11959) );
  NOR2X0 U11862 ( .IN1(n11961), .IN2(n11962), .QN(n11960) );
  NAND2X0 U11863 ( .IN1(n11963), .IN2(n11964), .QN(n11958) );
  NOR2X0 U11864 ( .IN1(n11965), .IN2(n11966), .QN(n11956) );
  NAND2X0 U11865 ( .IN1(n10565), .IN2(n10232), .QN(n11966) );
  NAND2X0 U11866 ( .IN1(n10171), .IN2(n11967), .QN(n11965) );
  NAND2X0 U11867 ( .IN1(n11968), .IN2(n11969), .QN(g34806) );
  NAND2X0 U11868 ( .IN1(n11073), .IN2(g2927), .QN(n11969) );
  NAND2X0 U11869 ( .IN1(n11970), .IN2(n10946), .QN(n11968) );
  NAND2X0 U11870 ( .IN1(n11971), .IN2(n10612), .QN(n11970) );
  NOR2X0 U11871 ( .IN1(g2941), .IN2(g4153), .QN(n11971) );
  NOR2X0 U11872 ( .IN1(n11052), .IN2(n11972), .QN(g34805) );
  NOR2X0 U11873 ( .IN1(g2999), .IN2(g2932), .QN(n11972) );
  NAND2X0 U11874 ( .IN1(n11973), .IN2(n11974), .QN(g34804) );
  NAND2X0 U11875 ( .IN1(n11073), .IN2(g2965), .QN(n11974) );
  NAND2X0 U11876 ( .IN1(n11975), .IN2(n10946), .QN(n11973) );
  NAND2X0 U11877 ( .IN1(n11976), .IN2(n5750), .QN(n11975) );
  NOR2X0 U11878 ( .IN1(n5796), .IN2(n5630), .QN(n11976) );
  NAND2X0 U11879 ( .IN1(n11977), .IN2(n11978), .QN(g34803) );
  NAND2X0 U11880 ( .IN1(n11073), .IN2(g2917), .QN(n11978) );
  NAND2X0 U11881 ( .IN1(n11979), .IN2(n10946), .QN(n11977) );
  NAND2X0 U11882 ( .IN1(n11980), .IN2(n10609), .QN(n11979) );
  NOR2X0 U11883 ( .IN1(g2932), .IN2(n11981), .QN(n11980) );
  INVX0 U11884 ( .INP(g44), .ZN(n11981) );
  NAND2X0 U11885 ( .IN1(n11982), .IN2(n11983), .QN(g34802) );
  NAND2X0 U11886 ( .IN1(n11073), .IN2(g2902), .QN(n11983) );
  NAND2X0 U11887 ( .IN1(n11984), .IN2(n10946), .QN(n11982) );
  NAND2X0 U11888 ( .IN1(n11985), .IN2(n10617), .QN(n11984) );
  NOR2X0 U11889 ( .IN1(n11986), .IN2(n11987), .QN(n11985) );
  NAND2X0 U11890 ( .IN1(n11988), .IN2(n11989), .QN(g34801) );
  NAND2X0 U11891 ( .IN1(n11072), .IN2(g2970), .QN(n11989) );
  NAND2X0 U11892 ( .IN1(n11990), .IN2(n10945), .QN(n11988) );
  NAND2X0 U11893 ( .IN1(n11991), .IN2(n10615), .QN(n11990) );
  NOR2X0 U11894 ( .IN1(n11992), .IN2(g301), .QN(n11991) );
  INVX0 U11895 ( .INP(n11993), .ZN(g34800) );
  NOR2X0 U11896 ( .IN1(n11994), .IN2(n11995), .QN(n11993) );
  NOR2X0 U11897 ( .IN1(n10906), .IN2(n10564), .QN(n11995) );
  NOR2X0 U11898 ( .IN1(n11996), .IN2(n11020), .QN(n11994) );
  NOR2X0 U11899 ( .IN1(test_so74), .IN2(test_so14), .QN(n11996) );
  NAND2X0 U11900 ( .IN1(n11997), .IN2(n11998), .QN(g34799) );
  NAND2X0 U11901 ( .IN1(n11072), .IN2(g2873), .QN(n11998) );
  NAND2X0 U11902 ( .IN1(n11999), .IN2(n10945), .QN(n11997) );
  NAND2X0 U11903 ( .IN1(n10568), .IN2(g44), .QN(n11999) );
  NAND2X0 U11904 ( .IN1(n12000), .IN2(n12001), .QN(g34798) );
  NAND2X0 U11905 ( .IN1(n11072), .IN2(g2878), .QN(n12001) );
  NAND2X0 U11906 ( .IN1(n12002), .IN2(n10945), .QN(n12000) );
  NAND2X0 U11907 ( .IN1(n10564), .IN2(n10565), .QN(n12002) );
  NAND2X0 U11908 ( .IN1(n12003), .IN2(n12004), .QN(g34797) );
  NAND2X0 U11909 ( .IN1(n11072), .IN2(g2882), .QN(n12004) );
  NAND2X0 U11910 ( .IN1(n12005), .IN2(n10945), .QN(n12003) );
  NAND2X0 U11911 ( .IN1(n10563), .IN2(g91), .QN(n12005) );
  NAND2X0 U11912 ( .IN1(n12006), .IN2(n12007), .QN(g34796) );
  NAND2X0 U11913 ( .IN1(n11072), .IN2(g2898), .QN(n12007) );
  NAND2X0 U11914 ( .IN1(n12008), .IN2(n10945), .QN(n12006) );
  NAND2X0 U11915 ( .IN1(n10616), .IN2(n11952), .QN(n12008) );
  NOR2X0 U11916 ( .IN1(n12009), .IN2(n12010), .QN(n11952) );
  NAND2X0 U11917 ( .IN1(n12011), .IN2(n12012), .QN(g34795) );
  NAND2X0 U11918 ( .IN1(n11072), .IN2(g2864), .QN(n12012) );
  NAND2X0 U11919 ( .IN1(n12013), .IN2(n10945), .QN(n12011) );
  NAND2X0 U11920 ( .IN1(n10566), .IN2(n11963), .QN(n12013) );
  INVX0 U11921 ( .INP(n12014), .ZN(n11963) );
  NAND2X0 U11922 ( .IN1(n12015), .IN2(n12016), .QN(n12014) );
  NOR2X0 U11923 ( .IN1(n12017), .IN2(n12018), .QN(n12016) );
  NOR2X0 U11924 ( .IN1(g3129), .IN2(g3143), .QN(n12015) );
  NAND2X0 U11925 ( .IN1(n12019), .IN2(n12020), .QN(g34794) );
  INVX0 U11926 ( .INP(n12021), .ZN(n12020) );
  NOR2X0 U11927 ( .IN1(n12022), .IN2(n12023), .QN(n12019) );
  NOR2X0 U11928 ( .IN1(n11051), .IN2(n12024), .QN(n12023) );
  NOR2X0 U11929 ( .IN1(n11962), .IN2(g2864), .QN(n12024) );
  NAND2X0 U11930 ( .IN1(n12025), .IN2(n12026), .QN(n11962) );
  NOR2X0 U11931 ( .IN1(n12027), .IN2(n12028), .QN(n12025) );
  NOR2X0 U11932 ( .IN1(n10618), .IN2(n10884), .QN(n12022) );
  NAND2X0 U11933 ( .IN1(n12029), .IN2(n12030), .QN(g34793) );
  NAND2X0 U11934 ( .IN1(n11072), .IN2(g2848), .QN(n12030) );
  NAND2X0 U11935 ( .IN1(n12031), .IN2(n10944), .QN(n12029) );
  NAND2X0 U11936 ( .IN1(n12032), .IN2(n10618), .QN(n12031) );
  NOR2X0 U11937 ( .IN1(n11961), .IN2(n12033), .QN(n12032) );
  NAND2X0 U11938 ( .IN1(n12034), .IN2(n12035), .QN(g34792) );
  NAND2X0 U11939 ( .IN1(n11072), .IN2(g29214), .QN(n12035) );
  NAND2X0 U11940 ( .IN1(n12036), .IN2(n10944), .QN(n12034) );
  NAND2X0 U11941 ( .IN1(n10613), .IN2(n11964), .QN(n12036) );
  NOR2X0 U11942 ( .IN1(n12037), .IN2(n12038), .QN(n11964) );
  INVX0 U11943 ( .INP(n12039), .ZN(n12037) );
  NAND2X0 U11944 ( .IN1(n12040), .IN2(n12041), .QN(g34791) );
  NAND2X0 U11945 ( .IN1(n11072), .IN2(g785), .QN(n12041) );
  NOR2X0 U11946 ( .IN1(n12042), .IN2(n12043), .QN(n12040) );
  NOR2X0 U11947 ( .IN1(g790), .IN2(n12044), .QN(n12043) );
  NOR2X0 U11948 ( .IN1(n5292), .IN2(n12045), .QN(n12042) );
  NAND2X0 U11949 ( .IN1(n2404), .IN2(n12044), .QN(n12045) );
  INVX0 U11950 ( .INP(n2425), .ZN(n12044) );
  NAND2X0 U11951 ( .IN1(n12046), .IN2(n12047), .QN(g34790) );
  NAND2X0 U11952 ( .IN1(n11072), .IN2(g617), .QN(n12047) );
  NOR2X0 U11953 ( .IN1(n12048), .IN2(n12049), .QN(n12046) );
  NOR2X0 U11954 ( .IN1(g622), .IN2(n12050), .QN(n12049) );
  NOR2X0 U11955 ( .IN1(n5672), .IN2(n12051), .QN(n12048) );
  NAND2X0 U11956 ( .IN1(n2421), .IN2(n12050), .QN(n12051) );
  INVX0 U11957 ( .INP(n2427), .ZN(n12050) );
  NOR2X0 U11958 ( .IN1(n5305), .IN2(n12052), .QN(g34788) );
  NOR2X0 U11959 ( .IN1(n10223), .IN2(n12053), .QN(n12052) );
  NAND2X0 U11960 ( .IN1(n12054), .IN2(n12055), .QN(g34783) );
  NAND2X0 U11961 ( .IN1(n12056), .IN2(n12057), .QN(n12055) );
  NOR2X0 U11962 ( .IN1(n12058), .IN2(n12059), .QN(n12056) );
  NAND2X0 U11963 ( .IN1(n12060), .IN2(n12061), .QN(n12054) );
  NOR2X0 U11964 ( .IN1(n12062), .IN2(n12063), .QN(n12060) );
  NAND2X0 U11965 ( .IN1(n12064), .IN2(n12065), .QN(g34735) );
  NAND2X0 U11966 ( .IN1(n11072), .IN2(g4297), .QN(n12065) );
  NAND2X0 U11967 ( .IN1(n12066), .IN2(n10944), .QN(n12064) );
  NAND2X0 U11968 ( .IN1(n5639), .IN2(n10567), .QN(n12066) );
  NAND2X0 U11969 ( .IN1(n12067), .IN2(n12068), .QN(g34734) );
  NAND2X0 U11970 ( .IN1(n11072), .IN2(g4172), .QN(n12068) );
  NAND2X0 U11971 ( .IN1(n12069), .IN2(n10944), .QN(n12067) );
  NAND2X0 U11972 ( .IN1(n5494), .IN2(n10612), .QN(n12069) );
  NOR2X0 U11973 ( .IN1(n11051), .IN2(n12070), .QN(g34733) );
  NOR2X0 U11974 ( .IN1(g4153), .IN2(g4172), .QN(n12070) );
  NAND2X0 U11975 ( .IN1(n12071), .IN2(n12072), .QN(g34732) );
  NAND2X0 U11976 ( .IN1(n10920), .IN2(g2994), .QN(n12072) );
  NAND2X0 U11977 ( .IN1(n11072), .IN2(g2999), .QN(n12071) );
  NAND2X0 U11978 ( .IN1(n12073), .IN2(n12074), .QN(g34731) );
  NAND2X0 U11979 ( .IN1(n11072), .IN2(g1283), .QN(n12074) );
  NAND2X0 U11980 ( .IN1(n12075), .IN2(n10944), .QN(n12073) );
  INVX0 U11981 ( .INP(n12076), .ZN(n12075) );
  NOR2X0 U11982 ( .IN1(n11986), .IN2(test_so64), .QN(n12076) );
  NAND2X0 U11983 ( .IN1(n12077), .IN2(n12078), .QN(g34730) );
  NAND2X0 U11984 ( .IN1(n11072), .IN2(g1296), .QN(n12078) );
  NAND2X0 U11985 ( .IN1(n12079), .IN2(n10944), .QN(n12077) );
  NAND2X0 U11986 ( .IN1(n5635), .IN2(n10570), .QN(n12079) );
  NAND2X0 U11987 ( .IN1(n12080), .IN2(n12081), .QN(g34729) );
  INVX0 U11988 ( .INP(n2499), .ZN(n12081) );
  NOR2X0 U11989 ( .IN1(n12082), .IN2(n12083), .QN(n12080) );
  NOR2X0 U11990 ( .IN1(n2549), .IN2(n10885), .QN(n12083) );
  NAND2X0 U11991 ( .IN1(n12084), .IN2(n12085), .QN(g34728) );
  NAND2X0 U11992 ( .IN1(n11072), .IN2(g939), .QN(n12085) );
  NAND2X0 U11993 ( .IN1(n12086), .IN2(n10943), .QN(n12084) );
  NAND2X0 U11994 ( .IN1(n19417), .IN2(n12087), .QN(n12086) );
  NAND2X0 U11995 ( .IN1(n12088), .IN2(n12089), .QN(g34727) );
  NAND2X0 U11996 ( .IN1(n11072), .IN2(g952), .QN(n12089) );
  NAND2X0 U11997 ( .IN1(n12090), .IN2(n10943), .QN(n12088) );
  NAND2X0 U11998 ( .IN1(n5415), .IN2(n10574), .QN(n12090) );
  NAND2X0 U11999 ( .IN1(n12091), .IN2(n12092), .QN(g34726) );
  INVX0 U12000 ( .INP(n2505), .ZN(n12092) );
  NOR2X0 U12001 ( .IN1(n12093), .IN2(n12094), .QN(n12091) );
  NOR2X0 U12002 ( .IN1(n5286), .IN2(n10885), .QN(n12094) );
  NOR2X0 U12003 ( .IN1(n11051), .IN2(g962), .QN(n12093) );
  NAND2X0 U12004 ( .IN1(n12095), .IN2(n12096), .QN(g34725) );
  NAND2X0 U12005 ( .IN1(n11071), .IN2(g781), .QN(n12096) );
  NOR2X0 U12006 ( .IN1(n12097), .IN2(n12098), .QN(n12095) );
  NOR2X0 U12007 ( .IN1(g785), .IN2(n12099), .QN(n12098) );
  NOR2X0 U12008 ( .IN1(n5293), .IN2(n12100), .QN(n12097) );
  NAND2X0 U12009 ( .IN1(n2404), .IN2(n12099), .QN(n12100) );
  INVX0 U12010 ( .INP(n2485), .ZN(n12099) );
  NAND2X0 U12011 ( .IN1(n12101), .IN2(n12102), .QN(g34724) );
  NAND2X0 U12012 ( .IN1(n11071), .IN2(g613), .QN(n12102) );
  NOR2X0 U12013 ( .IN1(n12103), .IN2(n12104), .QN(n12101) );
  NOR2X0 U12014 ( .IN1(g617), .IN2(n12105), .QN(n12104) );
  NOR2X0 U12015 ( .IN1(n5339), .IN2(n12106), .QN(n12103) );
  NAND2X0 U12016 ( .IN1(n2421), .IN2(n12105), .QN(n12106) );
  INVX0 U12017 ( .INP(n2487), .ZN(n12105) );
  NAND2X0 U12018 ( .IN1(n12107), .IN2(n12108), .QN(g34723) );
  NAND2X0 U12019 ( .IN1(test_so41), .IN2(n11081), .QN(n12108) );
  NAND2X0 U12020 ( .IN1(n12109), .IN2(n10943), .QN(n12107) );
  NAND2X0 U12021 ( .IN1(n5490), .IN2(n10614), .QN(n12109) );
  NAND2X0 U12022 ( .IN1(n12110), .IN2(n12111), .QN(g34722) );
  NAND2X0 U12023 ( .IN1(n11071), .IN2(g538), .QN(n12111) );
  NAND2X0 U12024 ( .IN1(n12112), .IN2(n10943), .QN(n12110) );
  NAND2X0 U12025 ( .IN1(n5492), .IN2(g691), .QN(n12112) );
  NAND2X0 U12026 ( .IN1(n12113), .IN2(n12114), .QN(g34721) );
  NAND2X0 U12027 ( .IN1(g29221), .IN2(n11081), .QN(n12114) );
  NAND2X0 U12028 ( .IN1(n12115), .IN2(n10943), .QN(n12113) );
  NAND2X0 U12029 ( .IN1(n10573), .IN2(n10572), .QN(n12115) );
  NAND2X0 U12030 ( .IN1(n12116), .IN2(n12117), .QN(g34720) );
  NAND2X0 U12031 ( .IN1(n11071), .IN2(g534), .QN(n12117) );
  NAND2X0 U12032 ( .IN1(n12118), .IN2(n10943), .QN(n12116) );
  NAND2X0 U12033 ( .IN1(n10571), .IN2(g29212), .QN(n12118) );
  NOR2X0 U12034 ( .IN1(n11050), .IN2(n12119), .QN(g34719) );
  NOR2X0 U12035 ( .IN1(g209), .IN2(g538), .QN(n12119) );
  NOR2X0 U12036 ( .IN1(n5497), .IN2(n11018), .QN(g34647) );
  NOR2X0 U12037 ( .IN1(n5644), .IN2(n11018), .QN(g34646) );
  NOR2X0 U12038 ( .IN1(n5499), .IN2(n11017), .QN(g34645) );
  NOR2X0 U12039 ( .IN1(n5643), .IN2(n11017), .QN(g34644) );
  NOR2X0 U12040 ( .IN1(n5498), .IN2(n11017), .QN(g34643) );
  NAND2X0 U12041 ( .IN1(n12120), .IN2(n12121), .QN(g34642) );
  NAND2X0 U12042 ( .IN1(n10920), .IN2(g4927), .QN(n12121) );
  NAND2X0 U12043 ( .IN1(n11071), .IN2(g4912), .QN(n12120) );
  NAND2X0 U12044 ( .IN1(n12122), .IN2(n12123), .QN(g34641) );
  NAND2X0 U12045 ( .IN1(n10920), .IN2(g4912), .QN(n12123) );
  NAND2X0 U12046 ( .IN1(n11071), .IN2(g4907), .QN(n12122) );
  NAND2X0 U12047 ( .IN1(n12124), .IN2(n12125), .QN(g34640) );
  NAND2X0 U12048 ( .IN1(n10921), .IN2(g4907), .QN(n12125) );
  NAND2X0 U12049 ( .IN1(n11071), .IN2(g4922), .QN(n12124) );
  NAND2X0 U12050 ( .IN1(n12126), .IN2(n12127), .QN(g34639) );
  NAND2X0 U12051 ( .IN1(n10921), .IN2(g4922), .QN(n12127) );
  NAND2X0 U12052 ( .IN1(n11071), .IN2(g4917), .QN(n12126) );
  NOR2X0 U12053 ( .IN1(n5408), .IN2(n11017), .QN(g34638) );
  NAND2X0 U12054 ( .IN1(n12128), .IN2(n12129), .QN(g34637) );
  NAND2X0 U12055 ( .IN1(n10921), .IN2(g4737), .QN(n12129) );
  NAND2X0 U12056 ( .IN1(n11071), .IN2(g4722), .QN(n12128) );
  NAND2X0 U12057 ( .IN1(n12130), .IN2(n12131), .QN(g34636) );
  NAND2X0 U12058 ( .IN1(n10921), .IN2(g4722), .QN(n12131) );
  NAND2X0 U12059 ( .IN1(n11071), .IN2(g4717), .QN(n12130) );
  NAND2X0 U12060 ( .IN1(n12132), .IN2(n12133), .QN(g34635) );
  NAND2X0 U12061 ( .IN1(n10921), .IN2(g4717), .QN(n12133) );
  NAND2X0 U12062 ( .IN1(n11071), .IN2(g4732), .QN(n12132) );
  NAND2X0 U12063 ( .IN1(n12134), .IN2(n12135), .QN(g34634) );
  NAND2X0 U12064 ( .IN1(n10921), .IN2(g4732), .QN(n12135) );
  NAND2X0 U12065 ( .IN1(n11071), .IN2(g4727), .QN(n12134) );
  NOR2X0 U12066 ( .IN1(n5312), .IN2(n11016), .QN(g34633) );
  NAND2X0 U12067 ( .IN1(n12136), .IN2(n12137), .QN(g34632) );
  NAND2X0 U12068 ( .IN1(n10922), .IN2(g4245), .QN(n12137) );
  NAND2X0 U12069 ( .IN1(test_so67), .IN2(n11080), .QN(n12136) );
  NAND2X0 U12070 ( .IN1(n12138), .IN2(n12139), .QN(g34631) );
  NAND2X0 U12071 ( .IN1(test_so67), .IN2(n10941), .QN(n12139) );
  NAND2X0 U12072 ( .IN1(n11071), .IN2(g4253), .QN(n12138) );
  NAND2X0 U12073 ( .IN1(n12140), .IN2(n12141), .QN(g34630) );
  NAND2X0 U12074 ( .IN1(n10922), .IN2(g4253), .QN(n12141) );
  NAND2X0 U12075 ( .IN1(n11071), .IN2(g4300), .QN(n12140) );
  NAND2X0 U12076 ( .IN1(n12142), .IN2(n12143), .QN(g34629) );
  NAND2X0 U12077 ( .IN1(n10922), .IN2(g4157), .QN(n12143) );
  NAND2X0 U12078 ( .IN1(n11071), .IN2(g4146), .QN(n12142) );
  NAND2X0 U12079 ( .IN1(n12144), .IN2(n12145), .QN(g34628) );
  NAND2X0 U12080 ( .IN1(n10922), .IN2(g4146), .QN(n12145) );
  NAND2X0 U12081 ( .IN1(n11071), .IN2(g4176), .QN(n12144) );
  NOR2X0 U12082 ( .IN1(n5641), .IN2(n11016), .QN(g34627) );
  NOR2X0 U12083 ( .IN1(n5495), .IN2(n11016), .QN(g34625) );
  NAND2X0 U12084 ( .IN1(n12146), .IN2(n12147), .QN(g34624) );
  NAND2X0 U12085 ( .IN1(n11071), .IN2(g2994), .QN(n12146) );
  NAND2X0 U12086 ( .IN1(n12148), .IN2(n12149), .QN(g34623) );
  NAND2X0 U12087 ( .IN1(n10923), .IN2(g2970), .QN(n12149) );
  NAND2X0 U12088 ( .IN1(test_so22), .IN2(n11080), .QN(n12148) );
  NAND2X0 U12089 ( .IN1(n12150), .IN2(n12151), .QN(g34622) );
  NAND2X0 U12090 ( .IN1(test_so22), .IN2(n10941), .QN(n12151) );
  NAND2X0 U12091 ( .IN1(n11070), .IN2(g2950), .QN(n12150) );
  NAND2X0 U12092 ( .IN1(n12152), .IN2(n12153), .QN(g34621) );
  NAND2X0 U12093 ( .IN1(n10923), .IN2(g2950), .QN(n12153) );
  NAND2X0 U12094 ( .IN1(n11070), .IN2(g2936), .QN(n12152) );
  NAND2X0 U12095 ( .IN1(n12154), .IN2(n12155), .QN(g34620) );
  NAND2X0 U12096 ( .IN1(n10923), .IN2(g2936), .QN(n12155) );
  NAND2X0 U12097 ( .IN1(n11070), .IN2(g2922), .QN(n12154) );
  NAND2X0 U12098 ( .IN1(n12156), .IN2(n12157), .QN(g34619) );
  NAND2X0 U12099 ( .IN1(n10923), .IN2(g2922), .QN(n12157) );
  NAND2X0 U12100 ( .IN1(n11070), .IN2(g2912), .QN(n12156) );
  NAND2X0 U12101 ( .IN1(n12158), .IN2(n12159), .QN(g34618) );
  NAND2X0 U12102 ( .IN1(n10923), .IN2(g2912), .QN(n12159) );
  NAND2X0 U12103 ( .IN1(test_so1), .IN2(n11080), .QN(n12158) );
  NAND2X0 U12104 ( .IN1(n12160), .IN2(n12161), .QN(g34617) );
  NAND2X0 U12105 ( .IN1(test_so1), .IN2(n10940), .QN(n12161) );
  NAND2X0 U12106 ( .IN1(n11070), .IN2(g2984), .QN(n12160) );
  NAND2X0 U12107 ( .IN1(n12162), .IN2(n12163), .QN(g34616) );
  NAND2X0 U12108 ( .IN1(n10923), .IN2(g2868), .QN(n12163) );
  NAND2X0 U12109 ( .IN1(n11070), .IN2(g2988), .QN(n12162) );
  NAND2X0 U12110 ( .IN1(n12164), .IN2(n12165), .QN(g34615) );
  NAND2X0 U12111 ( .IN1(n10923), .IN2(g2873), .QN(n12165) );
  NAND2X0 U12112 ( .IN1(n11070), .IN2(g2868), .QN(n12164) );
  NAND2X0 U12113 ( .IN1(n12166), .IN2(n12167), .QN(g34614) );
  NAND2X0 U12114 ( .IN1(n10924), .IN2(g29214), .QN(n12167) );
  NAND2X0 U12115 ( .IN1(g37), .IN2(n11080), .QN(n12166) );
  NAND2X0 U12116 ( .IN1(n12168), .IN2(n12169), .QN(g34613) );
  NAND2X0 U12117 ( .IN1(test_so95), .IN2(n11081), .QN(n12169) );
  NAND2X0 U12118 ( .IN1(g37), .IN2(n10941), .QN(n12168) );
  NAND2X0 U12119 ( .IN1(n12170), .IN2(n12171), .QN(g34612) );
  NAND2X0 U12120 ( .IN1(test_so95), .IN2(n10939), .QN(n12171) );
  NAND2X0 U12121 ( .IN1(n11070), .IN2(g2860), .QN(n12170) );
  NAND2X0 U12122 ( .IN1(n12172), .IN2(n12173), .QN(g34611) );
  NAND2X0 U12123 ( .IN1(n10924), .IN2(g2860), .QN(n12173) );
  NAND2X0 U12124 ( .IN1(n11070), .IN2(g2852), .QN(n12172) );
  NAND2X0 U12125 ( .IN1(n12174), .IN2(n12175), .QN(g34610) );
  NAND2X0 U12126 ( .IN1(n10924), .IN2(g2852), .QN(n12175) );
  NAND2X0 U12127 ( .IN1(n11070), .IN2(g2844), .QN(n12174) );
  NAND2X0 U12128 ( .IN1(n12176), .IN2(n12177), .QN(g34609) );
  NAND2X0 U12129 ( .IN1(n10924), .IN2(g2844), .QN(n12177) );
  NAND2X0 U12130 ( .IN1(n11070), .IN2(g2890), .QN(n12176) );
  NAND2X0 U12131 ( .IN1(n12178), .IN2(n12179), .QN(g34608) );
  NAND2X0 U12132 ( .IN1(n10924), .IN2(g2704), .QN(n12179) );
  NAND2X0 U12133 ( .IN1(n11070), .IN2(g2697), .QN(n12178) );
  NAND2X0 U12134 ( .IN1(n12180), .IN2(n12181), .QN(g34607) );
  NAND2X0 U12135 ( .IN1(n10924), .IN2(g2697), .QN(n12181) );
  NAND2X0 U12136 ( .IN1(n11070), .IN2(g2689), .QN(n12180) );
  NOR2X0 U12137 ( .IN1(n5347), .IN2(n11015), .QN(g34606) );
  NAND2X0 U12138 ( .IN1(n12182), .IN2(n12183), .QN(g34605) );
  NAND2X0 U12139 ( .IN1(n10925), .IN2(g2145), .QN(n12183) );
  NAND2X0 U12140 ( .IN1(n11070), .IN2(g2138), .QN(n12182) );
  NAND2X0 U12141 ( .IN1(n12184), .IN2(n12185), .QN(g34604) );
  NAND2X0 U12142 ( .IN1(n10925), .IN2(g2138), .QN(n12185) );
  NAND2X0 U12143 ( .IN1(n11070), .IN2(g2130), .QN(n12184) );
  NOR2X0 U12144 ( .IN1(n5487), .IN2(n11015), .QN(g34603) );
  NOR2X0 U12145 ( .IN1(n2549), .IN2(n11015), .QN(g34602) );
  NOR2X0 U12146 ( .IN1(n5286), .IN2(n11015), .QN(g34601) );
  NAND2X0 U12147 ( .IN1(n12186), .IN2(n12187), .QN(g34600) );
  NAND2X0 U12148 ( .IN1(n11070), .IN2(g776), .QN(n12187) );
  NOR2X0 U12149 ( .IN1(n12188), .IN2(n12189), .QN(n12186) );
  NOR2X0 U12150 ( .IN1(g781), .IN2(n12190), .QN(n12189) );
  NOR2X0 U12151 ( .IN1(n5551), .IN2(n12191), .QN(n12188) );
  NAND2X0 U12152 ( .IN1(n2404), .IN2(n12190), .QN(n12191) );
  INVX0 U12153 ( .INP(n2507), .ZN(n12190) );
  NAND2X0 U12154 ( .IN1(n12192), .IN2(n12193), .QN(g34599) );
  NAND2X0 U12155 ( .IN1(n11070), .IN2(g608), .QN(n12193) );
  NOR2X0 U12156 ( .IN1(n12194), .IN2(n12195), .QN(n12192) );
  NOR2X0 U12157 ( .IN1(g613), .IN2(n12196), .QN(n12195) );
  NOR2X0 U12158 ( .IN1(n5474), .IN2(n12197), .QN(n12194) );
  NAND2X0 U12159 ( .IN1(n2421), .IN2(n12196), .QN(n12197) );
  INVX0 U12160 ( .INP(n2509), .ZN(n12196) );
  NAND2X0 U12161 ( .IN1(n12198), .IN2(n12199), .QN(g34598) );
  NAND2X0 U12162 ( .IN1(n11069), .IN2(g550), .QN(n12199) );
  NAND2X0 U12163 ( .IN1(g29221), .IN2(n10940), .QN(n12198) );
  NAND2X0 U12164 ( .IN1(n12200), .IN2(n12201), .QN(g34468) );
  NAND2X0 U12165 ( .IN1(n12202), .IN2(g4854), .QN(n12201) );
  NAND2X0 U12166 ( .IN1(n12203), .IN2(n10938), .QN(n12202) );
  NAND2X0 U12167 ( .IN1(n12204), .IN2(n12205), .QN(n12203) );
  NAND2X0 U12168 ( .IN1(n12206), .IN2(g4859), .QN(n12200) );
  NAND2X0 U12169 ( .IN1(n12207), .IN2(n12208), .QN(g34467) );
  NAND2X0 U12170 ( .IN1(n12209), .IN2(n12206), .QN(n12208) );
  INVX0 U12171 ( .INP(n12210), .ZN(n12206) );
  XOR2X1 U12172 ( .IN1(g4854), .IN2(n12205), .Q(n12209) );
  INVX0 U12173 ( .INP(n12211), .ZN(n12205) );
  NAND2X0 U12174 ( .IN1(n2563), .IN2(g4849), .QN(n12211) );
  NAND2X0 U12175 ( .IN1(n11069), .IN2(g4849), .QN(n12207) );
  NAND2X0 U12176 ( .IN1(n12212), .IN2(n12213), .QN(g34466) );
  NAND2X0 U12177 ( .IN1(n12214), .IN2(g4878), .QN(n12213) );
  NAND2X0 U12178 ( .IN1(n12215), .IN2(n10941), .QN(n12214) );
  NAND2X0 U12179 ( .IN1(n10209), .IN2(n12204), .QN(n12215) );
  NAND2X0 U12180 ( .IN1(n12216), .IN2(n5283), .QN(n12212) );
  NOR2X0 U12181 ( .IN1(n10209), .IN2(n12210), .QN(n12216) );
  NAND2X0 U12182 ( .IN1(n12217), .IN2(n12218), .QN(g34465) );
  NAND2X0 U12183 ( .IN1(n11069), .IN2(g4843), .QN(n12218) );
  NOR2X0 U12184 ( .IN1(n12219), .IN2(n12220), .QN(n12217) );
  NOR2X0 U12185 ( .IN1(n12210), .IN2(n12221), .QN(n12220) );
  INVX0 U12186 ( .INP(n2567), .ZN(n12221) );
  NOR2X0 U12187 ( .IN1(g4849), .IN2(n12222), .QN(n12219) );
  NAND2X0 U12188 ( .IN1(n12204), .IN2(n2563), .QN(n12222) );
  NAND2X0 U12189 ( .IN1(n12223), .IN2(n12224), .QN(g34464) );
  NAND2X0 U12190 ( .IN1(n12225), .IN2(g4664), .QN(n12224) );
  NAND2X0 U12191 ( .IN1(n12226), .IN2(n10938), .QN(n12225) );
  NAND2X0 U12192 ( .IN1(n12227), .IN2(n12228), .QN(n12226) );
  NAND2X0 U12193 ( .IN1(n12229), .IN2(g4669), .QN(n12223) );
  NAND2X0 U12194 ( .IN1(n12230), .IN2(n12231), .QN(g34463) );
  NAND2X0 U12195 ( .IN1(n12232), .IN2(n12229), .QN(n12231) );
  XOR2X1 U12196 ( .IN1(g4664), .IN2(n12228), .Q(n12232) );
  INVX0 U12197 ( .INP(n12233), .ZN(n12228) );
  NAND2X0 U12198 ( .IN1(n2573), .IN2(g4659), .QN(n12233) );
  NAND2X0 U12199 ( .IN1(n11069), .IN2(g4659), .QN(n12230) );
  NAND2X0 U12200 ( .IN1(n12234), .IN2(n12235), .QN(g34462) );
  NAND2X0 U12201 ( .IN1(n12236), .IN2(g4688), .QN(n12235) );
  NAND2X0 U12202 ( .IN1(n12237), .IN2(n10940), .QN(n12236) );
  NAND2X0 U12203 ( .IN1(n12227), .IN2(n10645), .QN(n12237) );
  NAND2X0 U12204 ( .IN1(n12238), .IN2(n5656), .QN(n12234) );
  NOR2X0 U12205 ( .IN1(n10645), .IN2(n12239), .QN(n12238) );
  NAND2X0 U12206 ( .IN1(n12240), .IN2(n12241), .QN(g34461) );
  NAND2X0 U12207 ( .IN1(test_so19), .IN2(n11080), .QN(n12241) );
  NOR2X0 U12208 ( .IN1(n12242), .IN2(n12243), .QN(n12240) );
  NOR2X0 U12209 ( .IN1(n12239), .IN2(n12244), .QN(n12243) );
  INVX0 U12210 ( .INP(n2577), .ZN(n12244) );
  NOR2X0 U12211 ( .IN1(g4659), .IN2(n12245), .QN(n12242) );
  NAND2X0 U12212 ( .IN1(n12227), .IN2(n2573), .QN(n12245) );
  NAND2X0 U12213 ( .IN1(n12246), .IN2(n12247), .QN(g34460) );
  NAND2X0 U12214 ( .IN1(n12248), .IN2(g4639), .QN(n12247) );
  NAND2X0 U12215 ( .IN1(n12249), .IN2(n10938), .QN(n12248) );
  NAND2X0 U12216 ( .IN1(n12250), .IN2(n10667), .QN(n12249) );
  NAND2X0 U12217 ( .IN1(g34025), .IN2(test_so3), .QN(n12246) );
  NAND2X0 U12218 ( .IN1(n12251), .IN2(n12252), .QN(g34459) );
  INVX0 U12219 ( .INP(n12253), .ZN(n12252) );
  NOR2X0 U12220 ( .IN1(n10905), .IN2(n5382), .QN(n12253) );
  NAND2X0 U12221 ( .IN1(n12254), .IN2(n10938), .QN(n12251) );
  NAND2X0 U12222 ( .IN1(n12255), .IN2(n12256), .QN(n12254) );
  NAND2X0 U12223 ( .IN1(n12257), .IN2(n12258), .QN(n12256) );
  NAND2X0 U12224 ( .IN1(n5653), .IN2(n12259), .QN(n12257) );
  NAND2X0 U12225 ( .IN1(test_so99), .IN2(n12260), .QN(n12259) );
  NAND2X0 U12226 ( .IN1(n12261), .IN2(n12262), .QN(g34458) );
  NAND2X0 U12227 ( .IN1(n12263), .IN2(g4633), .QN(n12262) );
  NAND2X0 U12228 ( .IN1(n12264), .IN2(n12265), .QN(n12263) );
  NAND2X0 U12229 ( .IN1(n12266), .IN2(n12250), .QN(n12265) );
  NOR2X0 U12230 ( .IN1(test_so99), .IN2(n11017), .QN(n12266) );
  INVX0 U12231 ( .INP(n12267), .ZN(n12264) );
  NAND2X0 U12232 ( .IN1(test_so99), .IN2(n12268), .QN(n12261) );
  NAND2X0 U12233 ( .IN1(n12269), .IN2(n10937), .QN(n12268) );
  NAND2X0 U12234 ( .IN1(n12270), .IN2(n12271), .QN(n12269) );
  NOR2X0 U12235 ( .IN1(n5727), .IN2(n10667), .QN(n12271) );
  NOR2X0 U12236 ( .IN1(n12272), .IN2(g4633), .QN(n12270) );
  NAND2X0 U12237 ( .IN1(n12273), .IN2(n12274), .QN(g34457) );
  NAND2X0 U12238 ( .IN1(test_so3), .IN2(n12275), .QN(n12274) );
  NAND2X0 U12239 ( .IN1(n12276), .IN2(n10940), .QN(n12275) );
  NAND2X0 U12240 ( .IN1(n12277), .IN2(n12250), .QN(n12276) );
  NOR2X0 U12241 ( .IN1(test_so99), .IN2(n5727), .QN(n12277) );
  NAND2X0 U12242 ( .IN1(test_so99), .IN2(n12267), .QN(n12273) );
  NAND2X0 U12243 ( .IN1(n12278), .IN2(n12279), .QN(n12267) );
  NAND2X0 U12244 ( .IN1(n12280), .IN2(n12250), .QN(n12279) );
  NOR2X0 U12245 ( .IN1(test_so3), .IN2(n11017), .QN(n12280) );
  NAND2X0 U12246 ( .IN1(n12281), .IN2(n12282), .QN(g34456) );
  NAND2X0 U12247 ( .IN1(n12283), .IN2(g4608), .QN(n12282) );
  NAND2X0 U12248 ( .IN1(n12284), .IN2(n10937), .QN(n12283) );
  NAND2X0 U12249 ( .IN1(n2590), .IN2(n12285), .QN(n12284) );
  NAND2X0 U12250 ( .IN1(n12286), .IN2(g4616), .QN(n12281) );
  NAND2X0 U12251 ( .IN1(n12287), .IN2(n12288), .QN(g34455) );
  NAND2X0 U12252 ( .IN1(n12289), .IN2(g4322), .QN(n12288) );
  NAND2X0 U12253 ( .IN1(n12290), .IN2(n10937), .QN(n12289) );
  NAND2X0 U12254 ( .IN1(n12291), .IN2(n2594), .QN(n12290) );
  NOR2X0 U12255 ( .IN1(n12292), .IN2(n12293), .QN(n12291) );
  NAND2X0 U12256 ( .IN1(n2595), .IN2(g4332), .QN(n12287) );
  INVX0 U12257 ( .INP(n12294), .ZN(n2595) );
  NAND2X0 U12258 ( .IN1(n12295), .IN2(n12296), .QN(g34454) );
  NAND2X0 U12259 ( .IN1(n12297), .IN2(n12286), .QN(n12296) );
  XOR2X1 U12260 ( .IN1(n2590), .IN2(g4608), .Q(n12297) );
  NAND2X0 U12261 ( .IN1(n11069), .IN2(g4601), .QN(n12295) );
  NAND2X0 U12262 ( .IN1(n12298), .IN2(n12299), .QN(g34453) );
  NAND2X0 U12263 ( .IN1(n11069), .IN2(g4593), .QN(n12299) );
  NOR2X0 U12264 ( .IN1(n12300), .IN2(n12301), .QN(n12298) );
  NOR2X0 U12265 ( .IN1(g4601), .IN2(n12302), .QN(n12301) );
  NAND2X0 U12266 ( .IN1(n2598), .IN2(n12285), .QN(n12302) );
  INVX0 U12267 ( .INP(n12303), .ZN(n12285) );
  NOR2X0 U12268 ( .IN1(n5365), .IN2(n12304), .QN(n12300) );
  NAND2X0 U12269 ( .IN1(n12286), .IN2(n12305), .QN(n12304) );
  INVX0 U12270 ( .INP(n2598), .ZN(n12305) );
  NAND2X0 U12271 ( .IN1(n12306), .IN2(n12307), .QN(g34452) );
  NAND2X0 U12272 ( .IN1(n12308), .IN2(n12286), .QN(n12307) );
  XNOR2X1 U12273 ( .IN1(n2601), .IN2(n5303), .Q(n12308) );
  NAND2X0 U12274 ( .IN1(n11069), .IN2(g4584), .QN(n12306) );
  NAND2X0 U12275 ( .IN1(n12309), .IN2(n12310), .QN(g34451) );
  NAND2X0 U12276 ( .IN1(n12311), .IN2(n12286), .QN(n12310) );
  NOR2X0 U12277 ( .IN1(n12303), .IN2(n11017), .QN(n12286) );
  NAND2X0 U12278 ( .IN1(n12255), .IN2(n12312), .QN(n12303) );
  NAND2X0 U12279 ( .IN1(n2601), .IN2(g4616), .QN(n12312) );
  NOR2X0 U12280 ( .IN1(n12313), .IN2(n5539), .QN(n2601) );
  XOR2X1 U12281 ( .IN1(g4584), .IN2(n12292), .Q(n12311) );
  INVX0 U12282 ( .INP(n12313), .ZN(n12292) );
  NAND2X0 U12283 ( .IN1(n11069), .IN2(g4332), .QN(n12309) );
  NAND2X0 U12284 ( .IN1(n12314), .IN2(n12315), .QN(g34450) );
  NAND2X0 U12285 ( .IN1(n11069), .IN2(g4311), .QN(n12315) );
  NOR2X0 U12286 ( .IN1(n12316), .IN2(n12317), .QN(n12314) );
  NOR2X0 U12287 ( .IN1(g4322), .IN2(n12318), .QN(n12317) );
  NAND2X0 U12288 ( .IN1(n2594), .IN2(n12255), .QN(n12318) );
  INVX0 U12289 ( .INP(n12319), .ZN(n12316) );
  NAND2X0 U12290 ( .IN1(g4322), .IN2(n12320), .QN(n12319) );
  NOR2X0 U12291 ( .IN1(n12294), .IN2(n2594), .QN(n12320) );
  NAND2X0 U12292 ( .IN1(n12321), .IN2(n12313), .QN(n12294) );
  NAND2X0 U12293 ( .IN1(n12322), .IN2(n2607), .QN(n12313) );
  NOR2X0 U12294 ( .IN1(n12323), .IN2(n5348), .QN(n2607) );
  NOR2X0 U12295 ( .IN1(n5540), .IN2(n5506), .QN(n12322) );
  NAND2X0 U12296 ( .IN1(n12324), .IN2(n12325), .QN(g34448) );
  NAND2X0 U12297 ( .IN1(n12326), .IN2(n12327), .QN(n12325) );
  INVX0 U12298 ( .INP(n12328), .ZN(n12327) );
  NOR2X0 U12299 ( .IN1(n12329), .IN2(n12330), .QN(n12326) );
  NOR2X0 U12300 ( .IN1(n10122), .IN2(n12331), .QN(n12329) );
  NOR2X0 U12301 ( .IN1(n12332), .IN2(n12333), .QN(n12324) );
  NOR2X0 U12302 ( .IN1(n10122), .IN2(n10887), .QN(n12333) );
  NOR2X0 U12303 ( .IN1(n11049), .IN2(n12334), .QN(n12332) );
  NAND2X0 U12304 ( .IN1(n12328), .IN2(g2819), .QN(n12334) );
  NAND2X0 U12305 ( .IN1(n12335), .IN2(n12336), .QN(g34447) );
  NAND2X0 U12306 ( .IN1(n12337), .IN2(n12338), .QN(n12336) );
  INVX0 U12307 ( .INP(n12339), .ZN(n12338) );
  NOR2X0 U12308 ( .IN1(n12340), .IN2(n12330), .QN(n12337) );
  NOR2X0 U12309 ( .IN1(n10121), .IN2(n12331), .QN(n12340) );
  NOR2X0 U12310 ( .IN1(n12341), .IN2(n12342), .QN(n12335) );
  NOR2X0 U12311 ( .IN1(n5404), .IN2(n10887), .QN(n12342) );
  NOR2X0 U12312 ( .IN1(n11049), .IN2(n12343), .QN(n12341) );
  NAND2X0 U12313 ( .IN1(n12339), .IN2(g2807), .QN(n12343) );
  NAND2X0 U12314 ( .IN1(n12344), .IN2(n12345), .QN(g34446) );
  NAND2X0 U12315 ( .IN1(n12346), .IN2(n12347), .QN(n12345) );
  INVX0 U12316 ( .INP(n12348), .ZN(n12347) );
  NOR2X0 U12317 ( .IN1(n12349), .IN2(n12330), .QN(n12346) );
  NOR2X0 U12318 ( .IN1(n12331), .IN2(n10666), .QN(n12349) );
  NOR2X0 U12319 ( .IN1(n12350), .IN2(n12351), .QN(n12344) );
  NOR2X0 U12320 ( .IN1(n5609), .IN2(n10887), .QN(n12351) );
  NOR2X0 U12321 ( .IN1(n11049), .IN2(n12352), .QN(n12350) );
  NAND2X0 U12322 ( .IN1(n12348), .IN2(g2815), .QN(n12352) );
  NAND2X0 U12323 ( .IN1(n12353), .IN2(n12354), .QN(g34445) );
  NAND2X0 U12324 ( .IN1(n12355), .IN2(n12356), .QN(n12354) );
  INVX0 U12325 ( .INP(n12357), .ZN(n12356) );
  NOR2X0 U12326 ( .IN1(n12358), .IN2(n12330), .QN(n12355) );
  NAND2X0 U12327 ( .IN1(n12359), .IN2(n10939), .QN(n12330) );
  NAND2X0 U12328 ( .IN1(n2760), .IN2(n9255), .QN(n12359) );
  NOR2X0 U12329 ( .IN1(n10118), .IN2(n12331), .QN(n12358) );
  NOR2X0 U12330 ( .IN1(n12360), .IN2(n12361), .QN(n12353) );
  NOR2X0 U12331 ( .IN1(n5379), .IN2(n10887), .QN(n12361) );
  NOR2X0 U12332 ( .IN1(n11049), .IN2(n12362), .QN(n12360) );
  NAND2X0 U12333 ( .IN1(n12357), .IN2(g2803), .QN(n12362) );
  NAND2X0 U12334 ( .IN1(n12363), .IN2(n12364), .QN(g34444) );
  NAND2X0 U12335 ( .IN1(n12365), .IN2(n12366), .QN(n12364) );
  NOR2X0 U12336 ( .IN1(n12367), .IN2(n12328), .QN(n12365) );
  NOR2X0 U12337 ( .IN1(n10119), .IN2(n12331), .QN(n12367) );
  NOR2X0 U12338 ( .IN1(n12368), .IN2(n12369), .QN(n12363) );
  NOR2X0 U12339 ( .IN1(n10119), .IN2(n10888), .QN(n12369) );
  NOR2X0 U12340 ( .IN1(n11049), .IN2(n12370), .QN(n12368) );
  NAND2X0 U12341 ( .IN1(n12328), .IN2(g2787), .QN(n12370) );
  NAND2X0 U12342 ( .IN1(n12371), .IN2(n12372), .QN(n12328) );
  NOR2X0 U12343 ( .IN1(n5301), .IN2(n10274), .QN(n12371) );
  NAND2X0 U12344 ( .IN1(n12373), .IN2(n12374), .QN(g34443) );
  NAND2X0 U12345 ( .IN1(n12375), .IN2(n12366), .QN(n12374) );
  NOR2X0 U12346 ( .IN1(n12376), .IN2(n12339), .QN(n12375) );
  NOR2X0 U12347 ( .IN1(n10117), .IN2(n12331), .QN(n12376) );
  NOR2X0 U12348 ( .IN1(n12377), .IN2(n12378), .QN(n12373) );
  NOR2X0 U12349 ( .IN1(n5403), .IN2(n10888), .QN(n12378) );
  NOR2X0 U12350 ( .IN1(n11049), .IN2(n12379), .QN(n12377) );
  NAND2X0 U12351 ( .IN1(n12339), .IN2(g2775), .QN(n12379) );
  NAND2X0 U12352 ( .IN1(n12380), .IN2(n12372), .QN(n12339) );
  NOR2X0 U12353 ( .IN1(n5301), .IN2(g2729), .QN(n12380) );
  NAND2X0 U12354 ( .IN1(n12381), .IN2(n12382), .QN(g34442) );
  NAND2X0 U12355 ( .IN1(n12383), .IN2(n12366), .QN(n12382) );
  NOR2X0 U12356 ( .IN1(n12384), .IN2(n12348), .QN(n12383) );
  NOR2X0 U12357 ( .IN1(n10120), .IN2(n12331), .QN(n12384) );
  NOR2X0 U12358 ( .IN1(n12385), .IN2(n12386), .QN(n12381) );
  NOR2X0 U12359 ( .IN1(n5610), .IN2(n10888), .QN(n12386) );
  NOR2X0 U12360 ( .IN1(n11048), .IN2(n12387), .QN(n12385) );
  NAND2X0 U12361 ( .IN1(n12348), .IN2(g2783), .QN(n12387) );
  NAND2X0 U12362 ( .IN1(n12388), .IN2(n12372), .QN(n12348) );
  INVX0 U12363 ( .INP(n12389), .ZN(n12388) );
  NAND2X0 U12364 ( .IN1(n12390), .IN2(n12391), .QN(g34441) );
  NAND2X0 U12365 ( .IN1(n12392), .IN2(n12366), .QN(n12391) );
  NOR2X0 U12366 ( .IN1(n12393), .IN2(n11018), .QN(n12366) );
  NOR2X0 U12367 ( .IN1(n1770), .IN2(n10690), .QN(n12393) );
  NOR2X0 U12368 ( .IN1(n12394), .IN2(n12357), .QN(n12392) );
  NOR2X0 U12369 ( .IN1(n10123), .IN2(n12331), .QN(n12394) );
  NOR2X0 U12370 ( .IN1(n12395), .IN2(n12396), .QN(n12390) );
  NOR2X0 U12371 ( .IN1(n5378), .IN2(n10889), .QN(n12396) );
  NOR2X0 U12372 ( .IN1(n11048), .IN2(n12397), .QN(n12395) );
  NAND2X0 U12373 ( .IN1(n12357), .IN2(g2771), .QN(n12397) );
  NAND2X0 U12374 ( .IN1(n12372), .IN2(n12398), .QN(n12357) );
  NAND2X0 U12375 ( .IN1(n12399), .IN2(n12400), .QN(g34440) );
  NAND2X0 U12376 ( .IN1(n11069), .IN2(g446), .QN(n12400) );
  NAND2X0 U12377 ( .IN1(n12401), .IN2(n10975), .QN(n12399) );
  NAND2X0 U12378 ( .IN1(n12402), .IN2(n12403), .QN(n12401) );
  NAND2X0 U12379 ( .IN1(n12404), .IN2(g862), .QN(n12403) );
  NAND2X0 U12380 ( .IN1(g896), .IN2(n12405), .QN(n12404) );
  NAND2X0 U12381 ( .IN1(n12406), .IN2(n12407), .QN(n12405) );
  NAND2X0 U12382 ( .IN1(n5821), .IN2(n12408), .QN(n12406) );
  NAND2X0 U12383 ( .IN1(g890), .IN2(g896), .QN(n12402) );
  NAND2X0 U12384 ( .IN1(n12409), .IN2(n12410), .QN(g34439) );
  NAND2X0 U12385 ( .IN1(n11069), .IN2(g772), .QN(n12410) );
  NOR2X0 U12386 ( .IN1(n12411), .IN2(n12412), .QN(n12409) );
  NOR2X0 U12387 ( .IN1(g776), .IN2(n12413), .QN(n12412) );
  NOR2X0 U12388 ( .IN1(n5330), .IN2(n12414), .QN(n12411) );
  NAND2X0 U12389 ( .IN1(n2404), .IN2(n12413), .QN(n12414) );
  INVX0 U12390 ( .INP(n2554), .ZN(n12413) );
  NAND2X0 U12391 ( .IN1(n12415), .IN2(n12416), .QN(g34438) );
  NAND2X0 U12392 ( .IN1(n11069), .IN2(g604), .QN(n12416) );
  NOR2X0 U12393 ( .IN1(n12417), .IN2(n12418), .QN(n12415) );
  NOR2X0 U12394 ( .IN1(g608), .IN2(n12419), .QN(n12418) );
  NOR2X0 U12395 ( .IN1(n5475), .IN2(n12420), .QN(n12417) );
  NAND2X0 U12396 ( .IN1(n2421), .IN2(n12419), .QN(n12420) );
  INVX0 U12397 ( .INP(n2556), .ZN(n12419) );
  NOR2X0 U12398 ( .IN1(n12421), .IN2(n12422), .QN(g34435) );
  NAND2X0 U12399 ( .IN1(n5711), .IN2(n5416), .QN(n12422) );
  NAND2X0 U12400 ( .IN1(n10521), .IN2(n12423), .QN(n12421) );
  NAND2X0 U12401 ( .IN1(n12424), .IN2(n12425), .QN(n12423) );
  NAND2X0 U12402 ( .IN1(n12426), .IN2(n12427), .QN(n12425) );
  NOR2X0 U12403 ( .IN1(n10522), .IN2(n12428), .QN(n12427) );
  NOR2X0 U12404 ( .IN1(g4098), .IN2(n10644), .QN(n12426) );
  NAND2X0 U12405 ( .IN1(n2730), .IN2(n12429), .QN(g34425) );
  INVX0 U12406 ( .INP(n10626), .ZN(n12429) );
  NAND2X0 U12407 ( .IN1(n12430), .IN2(n12431), .QN(n10626) );
  NAND2X0 U12408 ( .IN1(n5348), .IN2(n12432), .QN(n12431) );
  NAND2X0 U12409 ( .IN1(n12433), .IN2(n12434), .QN(n12432) );
  NOR2X0 U12410 ( .IN1(n12435), .IN2(n12436), .QN(n12434) );
  NOR2X0 U12411 ( .IN1(n11283), .IN2(n12437), .QN(n12436) );
  NOR2X0 U12412 ( .IN1(n11271), .IN2(n12438), .QN(n12435) );
  NOR2X0 U12413 ( .IN1(n12439), .IN2(n12440), .QN(n12433) );
  NOR2X0 U12414 ( .IN1(n12441), .IN2(n12442), .QN(n12440) );
  NOR2X0 U12415 ( .IN1(n12443), .IN2(n12444), .QN(n12439) );
  NAND2X0 U12416 ( .IN1(n12445), .IN2(g4358), .QN(n12430) );
  NAND2X0 U12417 ( .IN1(n12446), .IN2(n12447), .QN(n12445) );
  NOR2X0 U12418 ( .IN1(n12448), .IN2(n12449), .QN(n12447) );
  NOR2X0 U12419 ( .IN1(n12437), .IN2(n12450), .QN(n12449) );
  NOR2X0 U12420 ( .IN1(n12451), .IN2(n12438), .QN(n12448) );
  NOR2X0 U12421 ( .IN1(n12452), .IN2(n12453), .QN(n12446) );
  NOR2X0 U12422 ( .IN1(n12441), .IN2(n12454), .QN(n12453) );
  NOR2X0 U12423 ( .IN1(n12444), .IN2(n12455), .QN(n12452) );
  NOR2X0 U12424 ( .IN1(n12456), .IN2(n12457), .QN(n2730) );
  NOR2X0 U12425 ( .IN1(n12458), .IN2(n12459), .QN(n12457) );
  NAND2X0 U12426 ( .IN1(n12460), .IN2(n12461), .QN(g34383) );
  NOR2X0 U12427 ( .IN1(g34843), .IN2(n12462), .QN(n12460) );
  NOR2X0 U12428 ( .IN1(n12463), .IN2(n12464), .QN(n12462) );
  NAND2X0 U12429 ( .IN1(n12465), .IN2(n12466), .QN(n12464) );
  INVX0 U12430 ( .INP(n12467), .ZN(n12465) );
  NAND2X0 U12431 ( .IN1(n3146), .IN2(n12468), .QN(n12467) );
  NAND2X0 U12432 ( .IN1(n12469), .IN2(n12470), .QN(n12463) );
  NOR2X0 U12433 ( .IN1(n12471), .IN2(n12472), .QN(n12470) );
  NOR2X0 U12434 ( .IN1(n12473), .IN2(n12474), .QN(n12469) );
  INVX0 U12435 ( .INP(n3165), .ZN(n12474) );
  NAND2X0 U12436 ( .IN1(n12475), .IN2(n12476), .QN(g34843) );
  NOR2X0 U12437 ( .IN1(n12477), .IN2(n12478), .QN(n12476) );
  NAND2X0 U12438 ( .IN1(n12479), .IN2(n12480), .QN(n12478) );
  NAND2X0 U12439 ( .IN1(n12481), .IN2(n5513), .QN(n12480) );
  NAND2X0 U12440 ( .IN1(n12482), .IN2(n5514), .QN(n12479) );
  NAND2X0 U12441 ( .IN1(n12483), .IN2(n12484), .QN(n12477) );
  NAND2X0 U12442 ( .IN1(n12485), .IN2(n5504), .QN(n12484) );
  NOR2X0 U12443 ( .IN1(n5536), .IN2(n12468), .QN(n12485) );
  NAND2X0 U12444 ( .IN1(n12486), .IN2(n5524), .QN(n12483) );
  NOR2X0 U12445 ( .IN1(n12487), .IN2(n12488), .QN(n12475) );
  NAND2X0 U12446 ( .IN1(n12489), .IN2(n12490), .QN(n12488) );
  NAND2X0 U12447 ( .IN1(n12491), .IN2(n12472), .QN(n12490) );
  NAND2X0 U12448 ( .IN1(g31862), .IN2(n12471), .QN(n12489) );
  NAND2X0 U12449 ( .IN1(n12492), .IN2(n12493), .QN(n12487) );
  INVX0 U12450 ( .INP(n12494), .ZN(n12493) );
  NOR2X0 U12451 ( .IN1(n12466), .IN2(n12495), .QN(n12494) );
  NAND2X0 U12452 ( .IN1(n12496), .IN2(n12497), .QN(g34269) );
  NAND2X0 U12453 ( .IN1(n12498), .IN2(n12499), .QN(n12497) );
  NOR2X0 U12454 ( .IN1(n5614), .IN2(n12500), .QN(n12498) );
  NOR2X0 U12455 ( .IN1(n12501), .IN2(n12502), .QN(n12496) );
  NOR2X0 U12456 ( .IN1(n5770), .IN2(n12503), .QN(n12502) );
  NOR2X0 U12457 ( .IN1(n11048), .IN2(n12504), .QN(n12503) );
  NOR2X0 U12458 ( .IN1(n12505), .IN2(n12506), .QN(n12504) );
  NAND2X0 U12459 ( .IN1(n12507), .IN2(n12508), .QN(g34268) );
  NAND2X0 U12460 ( .IN1(n12509), .IN2(n12499), .QN(n12508) );
  NOR2X0 U12461 ( .IN1(n5875), .IN2(n12510), .QN(n12509) );
  NOR2X0 U12462 ( .IN1(n12501), .IN2(n12511), .QN(n12507) );
  NOR2X0 U12463 ( .IN1(n5772), .IN2(n12512), .QN(n12511) );
  NOR2X0 U12464 ( .IN1(n11048), .IN2(n12513), .QN(n12512) );
  NOR2X0 U12465 ( .IN1(n12505), .IN2(n12514), .QN(n12513) );
  NAND2X0 U12466 ( .IN1(n12515), .IN2(n12516), .QN(g34267) );
  NAND2X0 U12467 ( .IN1(n12517), .IN2(g4939), .QN(n12516) );
  NAND2X0 U12468 ( .IN1(n12518), .IN2(n10975), .QN(n12517) );
  NAND2X0 U12469 ( .IN1(n12519), .IN2(n12520), .QN(n12518) );
  NOR2X0 U12470 ( .IN1(n12501), .IN2(n12521), .QN(n12515) );
  INVX0 U12471 ( .INP(n12522), .ZN(n12521) );
  NAND2X0 U12472 ( .IN1(n12499), .IN2(n12523), .QN(n12522) );
  NOR2X0 U12473 ( .IN1(n12519), .IN2(n5878), .QN(n12523) );
  NAND2X0 U12474 ( .IN1(n12524), .IN2(n12525), .QN(g34266) );
  NAND2X0 U12475 ( .IN1(n12526), .IN2(n12499), .QN(n12525) );
  NOR2X0 U12476 ( .IN1(n12505), .IN2(n11018), .QN(n12499) );
  NOR2X0 U12477 ( .IN1(n5863), .IN2(n12527), .QN(n12526) );
  NOR2X0 U12478 ( .IN1(n12501), .IN2(n12528), .QN(n12524) );
  NOR2X0 U12479 ( .IN1(n5774), .IN2(n12529), .QN(n12528) );
  NOR2X0 U12480 ( .IN1(n11048), .IN2(n12530), .QN(n12529) );
  NOR2X0 U12481 ( .IN1(n12505), .IN2(n12063), .QN(n12530) );
  INVX0 U12482 ( .INP(n12531), .ZN(n12501) );
  NAND2X0 U12483 ( .IN1(n12532), .IN2(n12505), .QN(n12531) );
  INVX0 U12484 ( .INP(n12520), .ZN(n12505) );
  NAND2X0 U12485 ( .IN1(n12533), .IN2(n5637), .QN(n12520) );
  NOR2X0 U12486 ( .IN1(test_so46), .IN2(n12534), .QN(n12533) );
  NOR2X0 U12487 ( .IN1(n19418), .IN2(n11019), .QN(n12532) );
  NOR2X0 U12488 ( .IN1(n11376), .IN2(n12210), .QN(g34265) );
  NAND2X0 U12489 ( .IN1(n12204), .IN2(n10975), .QN(n12210) );
  NOR2X0 U12490 ( .IN1(n12535), .IN2(n12061), .QN(n12204) );
  NAND2X0 U12491 ( .IN1(n12536), .IN2(n5713), .QN(n11376) );
  NOR2X0 U12492 ( .IN1(g4864), .IN2(g4871), .QN(n12536) );
  NAND2X0 U12493 ( .IN1(n12537), .IN2(n12538), .QN(g34264) );
  NAND2X0 U12494 ( .IN1(n12539), .IN2(n12540), .QN(n12538) );
  NOR2X0 U12495 ( .IN1(n5613), .IN2(n12541), .QN(n12539) );
  NOR2X0 U12496 ( .IN1(n12542), .IN2(n12543), .QN(n12537) );
  NOR2X0 U12497 ( .IN1(n5769), .IN2(n12544), .QN(n12543) );
  NOR2X0 U12498 ( .IN1(n11048), .IN2(n12545), .QN(n12544) );
  NOR2X0 U12499 ( .IN1(n12546), .IN2(n12547), .QN(n12545) );
  INVX0 U12500 ( .INP(n12541), .ZN(n12547) );
  NAND2X0 U12501 ( .IN1(n12548), .IN2(n12549), .QN(g34263) );
  NAND2X0 U12502 ( .IN1(n12550), .IN2(n12540), .QN(n12549) );
  NOR2X0 U12503 ( .IN1(n5877), .IN2(n12551), .QN(n12550) );
  NOR2X0 U12504 ( .IN1(n12542), .IN2(n12552), .QN(n12548) );
  NOR2X0 U12505 ( .IN1(n5775), .IN2(n12553), .QN(n12552) );
  NOR2X0 U12506 ( .IN1(n11048), .IN2(n12554), .QN(n12553) );
  NOR2X0 U12507 ( .IN1(n12546), .IN2(n12555), .QN(n12554) );
  INVX0 U12508 ( .INP(n12551), .ZN(n12555) );
  NAND2X0 U12509 ( .IN1(n12556), .IN2(n12557), .QN(g34262) );
  NAND2X0 U12510 ( .IN1(test_so18), .IN2(n12558), .QN(n12557) );
  NAND2X0 U12511 ( .IN1(n12559), .IN2(n10974), .QN(n12558) );
  NAND2X0 U12512 ( .IN1(n12560), .IN2(n12561), .QN(n12559) );
  NOR2X0 U12513 ( .IN1(n12542), .IN2(n12562), .QN(n12556) );
  INVX0 U12514 ( .INP(n12563), .ZN(n12562) );
  NAND2X0 U12515 ( .IN1(n12540), .IN2(n12564), .QN(n12563) );
  NOR2X0 U12516 ( .IN1(n12560), .IN2(n5876), .QN(n12564) );
  NAND2X0 U12517 ( .IN1(n12565), .IN2(n12566), .QN(g34261) );
  NAND2X0 U12518 ( .IN1(n12567), .IN2(n12540), .QN(n12566) );
  NOR2X0 U12519 ( .IN1(n12546), .IN2(n11019), .QN(n12540) );
  NOR2X0 U12520 ( .IN1(n5862), .IN2(n12568), .QN(n12567) );
  NOR2X0 U12521 ( .IN1(n12542), .IN2(n12569), .QN(n12565) );
  NOR2X0 U12522 ( .IN1(n5771), .IN2(n12570), .QN(n12569) );
  NOR2X0 U12523 ( .IN1(n11048), .IN2(n12571), .QN(n12570) );
  NOR2X0 U12524 ( .IN1(n12546), .IN2(n12059), .QN(n12571) );
  INVX0 U12525 ( .INP(n12568), .ZN(n12059) );
  INVX0 U12526 ( .INP(n12572), .ZN(n12542) );
  NAND2X0 U12527 ( .IN1(n12573), .IN2(n12546), .QN(n12572) );
  INVX0 U12528 ( .INP(n12561), .ZN(n12546) );
  NAND2X0 U12529 ( .IN1(n12574), .IN2(n19398), .QN(n12561) );
  NOR2X0 U12530 ( .IN1(n12534), .IN2(g4818), .QN(n12574) );
  NOR2X0 U12531 ( .IN1(n19411), .IN2(n11019), .QN(n12573) );
  NOR2X0 U12532 ( .IN1(n12575), .IN2(n12576), .QN(g34260) );
  NAND2X0 U12533 ( .IN1(n12229), .IN2(n5712), .QN(n12576) );
  INVX0 U12534 ( .INP(n12239), .ZN(n12229) );
  NAND2X0 U12535 ( .IN1(n12227), .IN2(n10974), .QN(n12239) );
  NOR2X0 U12536 ( .IN1(n12577), .IN2(n12057), .QN(n12227) );
  NAND2X0 U12537 ( .IN1(n5440), .IN2(n10527), .QN(n12575) );
  NOR2X0 U12538 ( .IN1(n5844), .IN2(n12578), .QN(g34259) );
  NOR2X0 U12539 ( .IN1(n11048), .IN2(n12579), .QN(n12578) );
  NOR2X0 U12540 ( .IN1(n12580), .IN2(n12272), .QN(n12579) );
  NAND2X0 U12541 ( .IN1(n12581), .IN2(n12582), .QN(g34258) );
  NAND2X0 U12542 ( .IN1(test_so81), .IN2(n11081), .QN(n12582) );
  NOR2X0 U12543 ( .IN1(n12583), .IN2(n12584), .QN(n12581) );
  NOR2X0 U12544 ( .IN1(g4358), .IN2(n12585), .QN(n12584) );
  NAND2X0 U12545 ( .IN1(n12586), .IN2(n12255), .QN(n12585) );
  INVX0 U12546 ( .INP(n12323), .ZN(n12586) );
  NOR2X0 U12547 ( .IN1(n5348), .IN2(n12587), .QN(n12583) );
  NAND2X0 U12548 ( .IN1(n12321), .IN2(n12323), .QN(n12587) );
  NAND2X0 U12549 ( .IN1(test_so81), .IN2(n12588), .QN(n12323) );
  NAND2X0 U12550 ( .IN1(n12589), .IN2(n12590), .QN(g34257) );
  NAND2X0 U12551 ( .IN1(n11069), .IN2(g4340), .QN(n12590) );
  NOR2X0 U12552 ( .IN1(n12591), .IN2(n12592), .QN(n12589) );
  NOR2X0 U12553 ( .IN1(n12258), .IN2(n12593), .QN(n12592) );
  NAND2X0 U12554 ( .IN1(n12255), .IN2(n10643), .QN(n12593) );
  NOR2X0 U12555 ( .IN1(n12588), .IN2(n12594), .QN(n12591) );
  NAND2X0 U12556 ( .IN1(n12321), .IN2(test_so81), .QN(n12594) );
  NOR2X0 U12557 ( .IN1(n12293), .IN2(n11020), .QN(n12321) );
  INVX0 U12558 ( .INP(n12255), .ZN(n12293) );
  INVX0 U12559 ( .INP(n12258), .ZN(n12588) );
  NAND2X0 U12560 ( .IN1(n12595), .IN2(test_so99), .QN(n12258) );
  NOR2X0 U12561 ( .IN1(n5653), .IN2(n12580), .QN(n12595) );
  NAND2X0 U12562 ( .IN1(n12596), .IN2(n12597), .QN(g34256) );
  NAND2X0 U12563 ( .IN1(n11069), .IN2(g4369), .QN(n12597) );
  NAND2X0 U12564 ( .IN1(n12598), .IN2(n10974), .QN(n12596) );
  NAND2X0 U12565 ( .IN1(n12599), .IN2(n5765), .QN(n12598) );
  NOR2X0 U12566 ( .IN1(n12600), .IN2(n12601), .QN(n12599) );
  NOR2X0 U12567 ( .IN1(n10207), .IN2(g4462), .QN(n12601) );
  NAND2X0 U12568 ( .IN1(n12602), .IN2(n12603), .QN(g34255) );
  NOR2X0 U12569 ( .IN1(n11048), .IN2(n12600), .QN(n12603) );
  NOR2X0 U12570 ( .IN1(n12604), .IN2(g4462), .QN(n12602) );
  NOR2X0 U12571 ( .IN1(n10207), .IN2(n10656), .QN(n12604) );
  NAND2X0 U12572 ( .IN1(n12605), .IN2(n12606), .QN(g34254) );
  NAND2X0 U12573 ( .IN1(n12607), .IN2(g4473), .QN(n12606) );
  NAND2X0 U12574 ( .IN1(n12608), .IN2(n12609), .QN(n12607) );
  NOR2X0 U12575 ( .IN1(test_so38), .IN2(n5671), .QN(n12609) );
  NOR2X0 U12576 ( .IN1(n5382), .IN2(n11020), .QN(n12608) );
  NAND2X0 U12577 ( .IN1(n12600), .IN2(n10974), .QN(n12605) );
  INVX0 U12578 ( .INP(n12610), .ZN(n12600) );
  NOR2X0 U12579 ( .IN1(n11048), .IN2(n12611), .QN(g34253) );
  NOR2X0 U12580 ( .IN1(n10656), .IN2(n12612), .QN(n12611) );
  NAND2X0 U12581 ( .IN1(n12610), .IN2(g4462), .QN(n12612) );
  NAND2X0 U12582 ( .IN1(n12613), .IN2(n5849), .QN(n12610) );
  NOR2X0 U12583 ( .IN1(n10281), .IN2(n12614), .QN(n12613) );
  NOR2X0 U12584 ( .IN1(n12615), .IN2(n11908), .QN(n12614) );
  INVX0 U12585 ( .INP(n12616), .ZN(n12615) );
  NAND2X0 U12586 ( .IN1(n1363), .IN2(n5846), .QN(n12616) );
  NAND2X0 U12587 ( .IN1(n12617), .IN2(n12618), .QN(g34252) );
  NAND2X0 U12588 ( .IN1(n11069), .IN2(g767), .QN(n12618) );
  NOR2X0 U12589 ( .IN1(n12619), .IN2(n12620), .QN(n12617) );
  NOR2X0 U12590 ( .IN1(g772), .IN2(n12621), .QN(n12620) );
  NOR2X0 U12591 ( .IN1(n5334), .IN2(n12622), .QN(n12619) );
  NAND2X0 U12592 ( .IN1(n2404), .IN2(n12621), .QN(n12622) );
  INVX0 U12593 ( .INP(n2647), .ZN(n12621) );
  NAND2X0 U12594 ( .IN1(n12623), .IN2(n12624), .QN(g34251) );
  NAND2X0 U12595 ( .IN1(n11069), .IN2(g599), .QN(n12624) );
  NOR2X0 U12596 ( .IN1(n12625), .IN2(n12626), .QN(n12623) );
  NOR2X0 U12597 ( .IN1(g604), .IN2(n12627), .QN(n12626) );
  NOR2X0 U12598 ( .IN1(n5473), .IN2(n12628), .QN(n12625) );
  NAND2X0 U12599 ( .IN1(n2421), .IN2(n12627), .QN(n12628) );
  INVX0 U12600 ( .INP(n2649), .ZN(n12627) );
  NAND2X0 U12601 ( .IN1(n12629), .IN2(n12630), .QN(g34250) );
  NAND2X0 U12602 ( .IN1(n11068), .IN2(g298), .QN(n12630) );
  NOR2X0 U12603 ( .IN1(n12631), .IN2(n12632), .QN(n12629) );
  NOR2X0 U12604 ( .IN1(n12633), .IN2(g142), .QN(n12632) );
  NOR2X0 U12605 ( .IN1(n5724), .IN2(n12634), .QN(n12631) );
  NAND2X0 U12606 ( .IN1(n95), .IN2(n12633), .QN(n12634) );
  NAND2X0 U12607 ( .IN1(n12635), .IN2(n12636), .QN(g34249) );
  NAND2X0 U12608 ( .IN1(n11068), .IN2(g157), .QN(n12636) );
  NOR2X0 U12609 ( .IN1(n12637), .IN2(n12638), .QN(n12635) );
  NOR2X0 U12610 ( .IN1(g160), .IN2(n12639), .QN(n12638) );
  NOR2X0 U12611 ( .IN1(n5843), .IN2(n12640), .QN(n12637) );
  NAND2X0 U12612 ( .IN1(n12641), .IN2(n12639), .QN(n12640) );
  INVX0 U12613 ( .INP(n2710), .ZN(n12639) );
  NAND2X0 U12614 ( .IN1(n12642), .IN2(n12461), .QN(g34201) );
  INVX0 U12615 ( .INP(n12456), .ZN(n12461) );
  NOR2X0 U12616 ( .IN1(g34781), .IN2(n12643), .QN(n12642) );
  NOR2X0 U12617 ( .IN1(n12644), .IN2(n12645), .QN(n12643) );
  NAND2X0 U12618 ( .IN1(n12646), .IN2(n12647), .QN(n12645) );
  NOR2X0 U12619 ( .IN1(n12648), .IN2(n12649), .QN(n12647) );
  NOR2X0 U12620 ( .IN1(n12650), .IN2(n12651), .QN(n12646) );
  NAND2X0 U12621 ( .IN1(n12652), .IN2(n12653), .QN(n12644) );
  NOR2X0 U12622 ( .IN1(n3005), .IN2(n12654), .QN(n12653) );
  NOR2X0 U12623 ( .IN1(n12655), .IN2(n12656), .QN(n12652) );
  NAND2X0 U12624 ( .IN1(n12657), .IN2(n12658), .QN(g34781) );
  NOR2X0 U12625 ( .IN1(n12659), .IN2(n12660), .QN(n12658) );
  NAND2X0 U12626 ( .IN1(n12661), .IN2(n12662), .QN(n12660) );
  NAND2X0 U12627 ( .IN1(n12663), .IN2(n5511), .QN(n12662) );
  NOR2X0 U12628 ( .IN1(n3550), .IN2(n10640), .QN(n12663) );
  NAND2X0 U12629 ( .IN1(n12664), .IN2(n5512), .QN(n12661) );
  NOR2X0 U12630 ( .IN1(n10532), .IN2(n3569), .QN(n12664) );
  NAND2X0 U12631 ( .IN1(n12665), .IN2(n12666), .QN(n12659) );
  NAND2X0 U12632 ( .IN1(n12667), .IN2(n5508), .QN(n12666) );
  NOR2X0 U12633 ( .IN1(n10529), .IN2(n3006), .QN(n12667) );
  NAND2X0 U12634 ( .IN1(n12668), .IN2(n5509), .QN(n12665) );
  NOR2X0 U12635 ( .IN1(n10530), .IN2(n3007), .QN(n12668) );
  NOR2X0 U12636 ( .IN1(n12669), .IN2(n12670), .QN(n12657) );
  NAND2X0 U12637 ( .IN1(n12671), .IN2(n12672), .QN(n12670) );
  NAND2X0 U12638 ( .IN1(n12673), .IN2(n5359), .QN(n12672) );
  NOR2X0 U12639 ( .IN1(n5596), .IN2(n1730), .QN(n12673) );
  INVX0 U12640 ( .INP(n3005), .ZN(n1730) );
  NAND2X0 U12641 ( .IN1(g25167), .IN2(n12654), .QN(n12671) );
  NAND2X0 U12642 ( .IN1(n12674), .IN2(n12675), .QN(n12669) );
  NAND2X0 U12643 ( .IN1(n12676), .IN2(n5507), .QN(n12675) );
  NOR2X0 U12644 ( .IN1(n10528), .IN2(n3588), .QN(n12676) );
  NAND2X0 U12645 ( .IN1(n12677), .IN2(n5510), .QN(n12674) );
  NOR2X0 U12646 ( .IN1(n10531), .IN2(n3606), .QN(n12677) );
  NAND2X0 U12647 ( .IN1(n12678), .IN2(n12679), .QN(g34041) );
  NAND2X0 U12648 ( .IN1(n12680), .IN2(n12681), .QN(n12679) );
  XOR2X1 U12649 ( .IN1(n12682), .IN2(n5367), .Q(n12680) );
  NAND2X0 U12650 ( .IN1(n11068), .IN2(g5008), .QN(n12678) );
  NAND2X0 U12651 ( .IN1(n12683), .IN2(n12684), .QN(g34040) );
  NAND2X0 U12652 ( .IN1(n11068), .IN2(g4975), .QN(n12684) );
  NOR2X0 U12653 ( .IN1(n12685), .IN2(n12686), .QN(n12683) );
  NOR2X0 U12654 ( .IN1(n5517), .IN2(n12687), .QN(n12686) );
  NOR2X0 U12655 ( .IN1(n12535), .IN2(n12688), .QN(n12685) );
  NOR2X0 U12656 ( .IN1(n12689), .IN2(n12690), .QN(n12688) );
  NOR2X0 U12657 ( .IN1(n11047), .IN2(n11403), .QN(n12690) );
  NOR2X0 U12658 ( .IN1(n11402), .IN2(n12691), .QN(n12689) );
  NAND2X0 U12659 ( .IN1(n12692), .IN2(n12693), .QN(g34039) );
  NAND2X0 U12660 ( .IN1(test_so58), .IN2(n12694), .QN(n12693) );
  NAND2X0 U12661 ( .IN1(n12695), .IN2(n10974), .QN(n12694) );
  NAND2X0 U12662 ( .IN1(n12681), .IN2(g4966), .QN(n12692) );
  NAND2X0 U12663 ( .IN1(n12696), .IN2(n12697), .QN(g34038) );
  NAND2X0 U12664 ( .IN1(n11068), .IN2(g4983), .QN(n12697) );
  NOR2X0 U12665 ( .IN1(n12698), .IN2(n12699), .QN(n12696) );
  NOR2X0 U12666 ( .IN1(n10652), .IN2(n12700), .QN(n12699) );
  NAND2X0 U12667 ( .IN1(n12681), .IN2(n12701), .QN(n12700) );
  INVX0 U12668 ( .INP(n12687), .ZN(n12681) );
  NOR2X0 U12669 ( .IN1(test_so58), .IN2(n12695), .QN(n12698) );
  NAND2X0 U12670 ( .IN1(n12702), .IN2(n12703), .QN(n12695) );
  NOR2X0 U12671 ( .IN1(n12535), .IN2(n12704), .QN(n12702) );
  NAND2X0 U12672 ( .IN1(n12705), .IN2(n12706), .QN(g34037) );
  NAND2X0 U12673 ( .IN1(n11068), .IN2(g4966), .QN(n12706) );
  NOR2X0 U12674 ( .IN1(n12707), .IN2(n12708), .QN(n12705) );
  NOR2X0 U12675 ( .IN1(g4975), .IN2(n12709), .QN(n12708) );
  NAND2X0 U12676 ( .IN1(n12704), .IN2(n12710), .QN(n12709) );
  INVX0 U12677 ( .INP(n12691), .ZN(n12704) );
  NOR2X0 U12678 ( .IN1(n5360), .IN2(n12687), .QN(n12707) );
  NAND2X0 U12679 ( .IN1(n12711), .IN2(n12691), .QN(n12687) );
  NAND2X0 U12680 ( .IN1(n12703), .IN2(g4966), .QN(n12691) );
  INVX0 U12681 ( .INP(n12701), .ZN(n12703) );
  NAND2X0 U12682 ( .IN1(n12061), .IN2(g4983), .QN(n12701) );
  INVX0 U12683 ( .INP(n12682), .ZN(n12061) );
  NAND2X0 U12684 ( .IN1(n12712), .IN2(n12713), .QN(n12682) );
  NOR2X0 U12685 ( .IN1(n5283), .IN2(n10542), .QN(n12713) );
  NOR2X0 U12686 ( .IN1(n10209), .IN2(n10099), .QN(n12712) );
  NOR2X0 U12687 ( .IN1(n11047), .IN2(n12535), .QN(n12711) );
  INVX0 U12688 ( .INP(n12710), .ZN(n12535) );
  NOR2X0 U12689 ( .IN1(n5443), .IN2(n12714), .QN(g34036) );
  NOR2X0 U12690 ( .IN1(n5318), .IN2(n12714), .QN(g34035) );
  NOR2X0 U12691 ( .IN1(n5713), .IN2(n12714), .QN(g34034) );
  NOR2X0 U12692 ( .IN1(n12710), .IN2(n11022), .QN(n12714) );
  NAND2X0 U12693 ( .IN1(n12715), .IN2(n12458), .QN(n12710) );
  NAND2X0 U12694 ( .IN1(n12716), .IN2(n12717), .QN(g34033) );
  NAND2X0 U12695 ( .IN1(n12718), .IN2(n12719), .QN(n12717) );
  XOR2X1 U12696 ( .IN1(n12720), .IN2(n5368), .Q(n12718) );
  NAND2X0 U12697 ( .IN1(n11068), .IN2(g4818), .QN(n12716) );
  NAND2X0 U12698 ( .IN1(n12721), .IN2(n12722), .QN(g34032) );
  NAND2X0 U12699 ( .IN1(n11068), .IN2(g4785), .QN(n12722) );
  NOR2X0 U12700 ( .IN1(n12723), .IN2(n12724), .QN(n12721) );
  NOR2X0 U12701 ( .IN1(n5518), .IN2(n12725), .QN(n12724) );
  NOR2X0 U12702 ( .IN1(n12577), .IN2(n12726), .QN(n12723) );
  NOR2X0 U12703 ( .IN1(n12727), .IN2(n12728), .QN(n12726) );
  NOR2X0 U12704 ( .IN1(n11047), .IN2(n11356), .QN(n12728) );
  NOR2X0 U12705 ( .IN1(n11357), .IN2(n12729), .QN(n12727) );
  NAND2X0 U12706 ( .IN1(n12730), .IN2(n12731), .QN(g34031) );
  NAND2X0 U12707 ( .IN1(test_so29), .IN2(n12732), .QN(n12731) );
  NAND2X0 U12708 ( .IN1(n12733), .IN2(n10974), .QN(n12732) );
  NAND2X0 U12709 ( .IN1(n12719), .IN2(g4776), .QN(n12730) );
  NAND2X0 U12710 ( .IN1(n12734), .IN2(n12735), .QN(g34030) );
  NAND2X0 U12711 ( .IN1(n11068), .IN2(g4793), .QN(n12735) );
  NOR2X0 U12712 ( .IN1(n12736), .IN2(n12737), .QN(n12734) );
  NOR2X0 U12713 ( .IN1(n10661), .IN2(n12738), .QN(n12737) );
  NAND2X0 U12714 ( .IN1(n12719), .IN2(n12739), .QN(n12738) );
  INVX0 U12715 ( .INP(n12725), .ZN(n12719) );
  NOR2X0 U12716 ( .IN1(test_so29), .IN2(n12733), .QN(n12736) );
  NAND2X0 U12717 ( .IN1(n12740), .IN2(n12741), .QN(n12733) );
  NOR2X0 U12718 ( .IN1(n12577), .IN2(n12742), .QN(n12740) );
  NAND2X0 U12719 ( .IN1(n12743), .IN2(n12744), .QN(g34029) );
  NAND2X0 U12720 ( .IN1(n11068), .IN2(g4776), .QN(n12744) );
  NOR2X0 U12721 ( .IN1(n12745), .IN2(n12746), .QN(n12743) );
  NOR2X0 U12722 ( .IN1(g4785), .IN2(n12747), .QN(n12746) );
  NAND2X0 U12723 ( .IN1(n12742), .IN2(n12748), .QN(n12747) );
  INVX0 U12724 ( .INP(n12729), .ZN(n12742) );
  NOR2X0 U12725 ( .IN1(n5361), .IN2(n12725), .QN(n12745) );
  NAND2X0 U12726 ( .IN1(n12749), .IN2(n12729), .QN(n12725) );
  NAND2X0 U12727 ( .IN1(n12741), .IN2(g4776), .QN(n12729) );
  INVX0 U12728 ( .INP(n12739), .ZN(n12741) );
  NAND2X0 U12729 ( .IN1(n12057), .IN2(g4793), .QN(n12739) );
  INVX0 U12730 ( .INP(n12720), .ZN(n12057) );
  NAND2X0 U12731 ( .IN1(n12750), .IN2(n12751), .QN(n12720) );
  NOR2X0 U12732 ( .IN1(n5656), .IN2(n10543), .QN(n12751) );
  NOR2X0 U12733 ( .IN1(n10103), .IN2(n10645), .QN(n12750) );
  NOR2X0 U12734 ( .IN1(n11047), .IN2(n12577), .QN(n12749) );
  INVX0 U12735 ( .INP(n12748), .ZN(n12577) );
  NOR2X0 U12736 ( .IN1(n5440), .IN2(n2774), .QN(g34027) );
  NOR2X0 U12737 ( .IN1(n5712), .IN2(n2774), .QN(g34026) );
  NOR2X0 U12738 ( .IN1(n12748), .IN2(n11023), .QN(n2774) );
  NAND2X0 U12739 ( .IN1(n12715), .IN2(n12459), .QN(n12748) );
  NOR2X0 U12740 ( .IN1(n10237), .IN2(n1770), .QN(n12715) );
  INVX0 U12741 ( .INP(n12278), .ZN(g34025) );
  NAND2X0 U12742 ( .IN1(n12752), .IN2(n12250), .QN(n12278) );
  INVX0 U12743 ( .INP(n12272), .ZN(n12250) );
  NAND2X0 U12744 ( .IN1(n5382), .IN2(n12255), .QN(n12272) );
  NAND2X0 U12745 ( .IN1(n9281), .IN2(n12753), .QN(n12255) );
  NAND2X0 U12746 ( .IN1(n12754), .IN2(n1770), .QN(n12753) );
  NOR2X0 U12747 ( .IN1(n11047), .IN2(g4639), .QN(n12752) );
  NAND2X0 U12748 ( .IN1(n12755), .IN2(n12756), .QN(g34024) );
  NOR2X0 U12749 ( .IN1(n12757), .IN2(n12758), .QN(n12756) );
  NOR2X0 U12750 ( .IN1(n11047), .IN2(n12759), .QN(n12758) );
  NOR2X0 U12751 ( .IN1(n12760), .IN2(n12761), .QN(n12759) );
  NOR2X0 U12752 ( .IN1(n11908), .IN2(n12762), .QN(n12761) );
  NOR2X0 U12753 ( .IN1(n10265), .IN2(n12754), .QN(n12760) );
  NOR2X0 U12754 ( .IN1(n10541), .IN2(n10889), .QN(n12757) );
  NAND2X0 U12755 ( .IN1(n12763), .IN2(n12755), .QN(g34023) );
  NOR2X0 U12756 ( .IN1(n12764), .IN2(n12765), .QN(n12755) );
  NOR2X0 U12757 ( .IN1(n12147), .IN2(n11908), .QN(n12765) );
  NAND2X0 U12758 ( .IN1(g2988), .IN2(n10974), .QN(n12147) );
  NOR2X0 U12759 ( .IN1(n12766), .IN2(n12767), .QN(n12763) );
  NOR2X0 U12760 ( .IN1(n19399), .IN2(n12768), .QN(n12767) );
  NOR2X0 U12761 ( .IN1(n11047), .IN2(n12769), .QN(n12768) );
  NOR2X0 U12762 ( .IN1(n12770), .IN2(n12771), .QN(n12769) );
  NAND2X0 U12763 ( .IN1(n12754), .IN2(g4555), .QN(n12771) );
  NAND2X0 U12764 ( .IN1(g4558), .IN2(g4561), .QN(n12770) );
  NOR2X0 U12765 ( .IN1(n12754), .IN2(n12772), .QN(n12766) );
  NAND2X0 U12766 ( .IN1(n10926), .IN2(g4552), .QN(n12772) );
  NAND2X0 U12767 ( .IN1(n12773), .IN2(n12774), .QN(g34022) );
  NOR2X0 U12768 ( .IN1(n12775), .IN2(n12776), .QN(n12774) );
  NOR2X0 U12769 ( .IN1(n10096), .IN2(n10889), .QN(n12776) );
  NOR2X0 U12770 ( .IN1(n11046), .IN2(n12777), .QN(n12775) );
  NAND2X0 U12771 ( .IN1(n12778), .IN2(g2763), .QN(n12777) );
  NOR2X0 U12772 ( .IN1(n2787), .IN2(n12779), .QN(n12773) );
  NOR2X0 U12773 ( .IN1(g2763), .IN2(n12778), .QN(n12779) );
  INVX0 U12774 ( .INP(n12780), .ZN(n12778) );
  NOR2X0 U12775 ( .IN1(n12781), .IN2(n10096), .QN(n12780) );
  NAND2X0 U12776 ( .IN1(n12782), .IN2(n12783), .QN(g34021) );
  NAND2X0 U12777 ( .IN1(n11068), .IN2(g2648), .QN(n12783) );
  NOR2X0 U12778 ( .IN1(n12784), .IN2(n12785), .QN(n12782) );
  NOR2X0 U12779 ( .IN1(n10134), .IN2(n12786), .QN(n12785) );
  NOR2X0 U12780 ( .IN1(n12787), .IN2(n12788), .QN(n12784) );
  NAND2X0 U12781 ( .IN1(n12789), .IN2(n12790), .QN(g34020) );
  NAND2X0 U12782 ( .IN1(n12791), .IN2(n12792), .QN(n12790) );
  NOR2X0 U12783 ( .IN1(n10197), .IN2(n12793), .QN(n12792) );
  NOR2X0 U12784 ( .IN1(n12794), .IN2(n12795), .QN(n12791) );
  NOR2X0 U12785 ( .IN1(n12796), .IN2(g2629), .QN(n12794) );
  NOR2X0 U12786 ( .IN1(n12797), .IN2(n12798), .QN(n12789) );
  NOR2X0 U12787 ( .IN1(n11046), .IN2(n12799), .QN(n12798) );
  NOR2X0 U12788 ( .IN1(n12800), .IN2(n12801), .QN(n12799) );
  NOR2X0 U12789 ( .IN1(n10197), .IN2(n12802), .QN(n12801) );
  NOR2X0 U12790 ( .IN1(n12803), .IN2(n12804), .QN(n12800) );
  NOR2X0 U12791 ( .IN1(n12795), .IN2(n12793), .QN(n12804) );
  INVX0 U12792 ( .INP(n12805), .ZN(n12793) );
  NOR2X0 U12793 ( .IN1(g1589), .IN2(n12806), .QN(n12795) );
  NOR2X0 U12794 ( .IN1(n12807), .IN2(n12808), .QN(n12803) );
  NOR2X0 U12795 ( .IN1(n12809), .IN2(g2643), .QN(n12807) );
  NOR2X0 U12796 ( .IN1(n5521), .IN2(n10890), .QN(n12797) );
  NAND2X0 U12797 ( .IN1(n12810), .IN2(n12811), .QN(g34019) );
  NAND2X0 U12798 ( .IN1(n12812), .IN2(n12813), .QN(n12811) );
  INVX0 U12799 ( .INP(n12814), .ZN(n12812) );
  NOR2X0 U12800 ( .IN1(n12815), .IN2(n12816), .QN(n12810) );
  NOR2X0 U12801 ( .IN1(n5787), .IN2(n10890), .QN(n12816) );
  NOR2X0 U12802 ( .IN1(n11046), .IN2(n12817), .QN(n12815) );
  NAND2X0 U12803 ( .IN1(n12814), .IN2(g2583), .QN(n12817) );
  NAND2X0 U12804 ( .IN1(n12818), .IN2(g2629), .QN(n12814) );
  NAND2X0 U12805 ( .IN1(n12819), .IN2(n12820), .QN(g34018) );
  NAND2X0 U12806 ( .IN1(n12821), .IN2(n12813), .QN(n12820) );
  NOR2X0 U12807 ( .IN1(n12822), .IN2(n12823), .QN(n12819) );
  NOR2X0 U12808 ( .IN1(n5800), .IN2(n10890), .QN(n12823) );
  NOR2X0 U12809 ( .IN1(n11046), .IN2(n12824), .QN(n12822) );
  NAND2X0 U12810 ( .IN1(test_so61), .IN2(n12825), .QN(n12824) );
  INVX0 U12811 ( .INP(n12821), .ZN(n12825) );
  NOR2X0 U12812 ( .IN1(n12826), .IN2(g2555), .QN(n12821) );
  NAND2X0 U12813 ( .IN1(n12827), .IN2(n12828), .QN(g34017) );
  INVX0 U12814 ( .INP(n12829), .ZN(n12828) );
  NOR2X0 U12815 ( .IN1(n12830), .IN2(n12787), .QN(n12829) );
  NOR2X0 U12816 ( .IN1(n12831), .IN2(n12832), .QN(n12827) );
  NOR2X0 U12817 ( .IN1(n10903), .IN2(n10663), .QN(n12832) );
  NOR2X0 U12818 ( .IN1(n11046), .IN2(n12833), .QN(n12831) );
  NAND2X0 U12819 ( .IN1(test_so66), .IN2(n12830), .QN(n12833) );
  NAND2X0 U12820 ( .IN1(n12834), .IN2(n12802), .QN(n12830) );
  NOR2X0 U12821 ( .IN1(n5521), .IN2(n5351), .QN(n12834) );
  NAND2X0 U12822 ( .IN1(n12835), .IN2(n12836), .QN(g34016) );
  NAND2X0 U12823 ( .IN1(n12837), .IN2(n12813), .QN(n12836) );
  NOR2X0 U12824 ( .IN1(n12838), .IN2(n12839), .QN(n12835) );
  NOR2X0 U12825 ( .IN1(n5816), .IN2(n10890), .QN(n12839) );
  INVX0 U12826 ( .INP(n12840), .ZN(n12838) );
  NAND2X0 U12827 ( .IN1(n10925), .IN2(n12841), .QN(n12840) );
  NOR2X0 U12828 ( .IN1(n12837), .IN2(n5787), .QN(n12841) );
  NOR2X0 U12829 ( .IN1(n12826), .IN2(g2629), .QN(n12837) );
  NAND2X0 U12830 ( .IN1(n12842), .IN2(n12843), .QN(g34015) );
  NAND2X0 U12831 ( .IN1(n12844), .IN2(n12813), .QN(n12843) );
  INVX0 U12832 ( .INP(n12787), .ZN(n12813) );
  NAND2X0 U12833 ( .IN1(n12845), .IN2(n10973), .QN(n12787) );
  NAND2X0 U12834 ( .IN1(n12846), .IN2(n12805), .QN(n12845) );
  NAND2X0 U12835 ( .IN1(n12847), .IN2(n12848), .QN(n12805) );
  NAND2X0 U12836 ( .IN1(n5483), .IN2(n12849), .QN(n12848) );
  NOR2X0 U12837 ( .IN1(n12850), .IN2(n12851), .QN(n12847) );
  NAND2X0 U12838 ( .IN1(n5757), .IN2(n12851), .QN(n12846) );
  INVX0 U12839 ( .INP(n12852), .ZN(n12844) );
  NOR2X0 U12840 ( .IN1(n12853), .IN2(n12854), .QN(n12842) );
  NOR2X0 U12841 ( .IN1(n10134), .IN2(n10890), .QN(n12854) );
  NOR2X0 U12842 ( .IN1(n11046), .IN2(n12855), .QN(n12853) );
  NAND2X0 U12843 ( .IN1(n12852), .IN2(g2563), .QN(n12855) );
  NAND2X0 U12844 ( .IN1(n12818), .IN2(g2555), .QN(n12852) );
  NAND2X0 U12845 ( .IN1(n12856), .IN2(n12857), .QN(g34014) );
  NAND2X0 U12846 ( .IN1(n11068), .IN2(g2514), .QN(n12857) );
  NOR2X0 U12847 ( .IN1(n12858), .IN2(n12859), .QN(n12856) );
  NOR2X0 U12848 ( .IN1(n10136), .IN2(n11237), .QN(n12859) );
  NOR2X0 U12849 ( .IN1(n12860), .IN2(n12861), .QN(n12858) );
  NAND2X0 U12850 ( .IN1(n12862), .IN2(n12863), .QN(g34013) );
  NAND2X0 U12851 ( .IN1(n12864), .IN2(n12865), .QN(n12863) );
  NOR2X0 U12852 ( .IN1(n10196), .IN2(n12866), .QN(n12865) );
  NOR2X0 U12853 ( .IN1(n12867), .IN2(n12868), .QN(n12864) );
  NOR2X0 U12854 ( .IN1(n12869), .IN2(g2495), .QN(n12868) );
  NOR2X0 U12855 ( .IN1(n11046), .IN2(n10648), .QN(n12869) );
  NOR2X0 U12856 ( .IN1(n12870), .IN2(n12871), .QN(n12862) );
  NOR2X0 U12857 ( .IN1(n11046), .IN2(n12872), .QN(n12871) );
  NOR2X0 U12858 ( .IN1(n12873), .IN2(n12874), .QN(n12872) );
  NOR2X0 U12859 ( .IN1(n10196), .IN2(n12875), .QN(n12874) );
  NOR2X0 U12860 ( .IN1(n12876), .IN2(n12877), .QN(n12873) );
  NOR2X0 U12861 ( .IN1(n12867), .IN2(n12866), .QN(n12877) );
  INVX0 U12862 ( .INP(n12878), .ZN(n12866) );
  NOR2X0 U12863 ( .IN1(n12879), .IN2(n5755), .QN(n12867) );
  NOR2X0 U12864 ( .IN1(n12880), .IN2(n12881), .QN(n12876) );
  NOR2X0 U12865 ( .IN1(n12882), .IN2(g2509), .QN(n12880) );
  NOR2X0 U12866 ( .IN1(n5522), .IN2(n10892), .QN(n12870) );
  NAND2X0 U12867 ( .IN1(n12883), .IN2(n12884), .QN(g34012) );
  NAND2X0 U12868 ( .IN1(n12885), .IN2(n12886), .QN(n12884) );
  NOR2X0 U12869 ( .IN1(n12887), .IN2(n12888), .QN(n12883) );
  NOR2X0 U12870 ( .IN1(n5789), .IN2(n10892), .QN(n12888) );
  INVX0 U12871 ( .INP(n12889), .ZN(n12887) );
  NAND2X0 U12872 ( .IN1(n10922), .IN2(n12890), .QN(n12889) );
  NOR2X0 U12873 ( .IN1(n12885), .IN2(n5798), .QN(n12890) );
  NOR2X0 U12874 ( .IN1(n12891), .IN2(n12882), .QN(n12885) );
  NAND2X0 U12875 ( .IN1(n12892), .IN2(n12893), .QN(g34011) );
  NAND2X0 U12876 ( .IN1(n12894), .IN2(n12886), .QN(n12893) );
  NOR2X0 U12877 ( .IN1(n12895), .IN2(n12896), .QN(n12892) );
  NOR2X0 U12878 ( .IN1(n5798), .IN2(n10900), .QN(n12896) );
  NOR2X0 U12879 ( .IN1(n11046), .IN2(n12897), .QN(n12895) );
  INVX0 U12880 ( .INP(n12898), .ZN(n12897) );
  NOR2X0 U12881 ( .IN1(n12894), .IN2(n19416), .QN(n12898) );
  NOR2X0 U12882 ( .IN1(n12899), .IN2(test_so79), .QN(n12894) );
  NAND2X0 U12883 ( .IN1(n12900), .IN2(n12901), .QN(g34010) );
  NAND2X0 U12884 ( .IN1(n12902), .IN2(n12886), .QN(n12901) );
  NOR2X0 U12885 ( .IN1(n12903), .IN2(n12904), .QN(n12900) );
  NOR2X0 U12886 ( .IN1(n19416), .IN2(n10901), .QN(n12904) );
  NOR2X0 U12887 ( .IN1(n11046), .IN2(n12905), .QN(n12903) );
  NAND2X0 U12888 ( .IN1(n12906), .IN2(g2441), .QN(n12905) );
  INVX0 U12889 ( .INP(n12902), .ZN(n12906) );
  NOR2X0 U12890 ( .IN1(n12907), .IN2(n5522), .QN(n12902) );
  NAND2X0 U12891 ( .IN1(n12908), .IN2(n12909), .QN(g34009) );
  NAND2X0 U12892 ( .IN1(n12910), .IN2(n12886), .QN(n12909) );
  NOR2X0 U12893 ( .IN1(n12911), .IN2(n12912), .QN(n12908) );
  NOR2X0 U12894 ( .IN1(n5814), .IN2(n10901), .QN(n12912) );
  NOR2X0 U12895 ( .IN1(n11046), .IN2(n12913), .QN(n12911) );
  INVX0 U12896 ( .INP(n12914), .ZN(n12913) );
  NOR2X0 U12897 ( .IN1(n12910), .IN2(n5789), .QN(n12914) );
  NOR2X0 U12898 ( .IN1(n12899), .IN2(g2495), .QN(n12910) );
  NAND2X0 U12899 ( .IN1(n12915), .IN2(n12916), .QN(g34008) );
  NAND2X0 U12900 ( .IN1(n12917), .IN2(n12886), .QN(n12916) );
  INVX0 U12901 ( .INP(n12860), .ZN(n12886) );
  NAND2X0 U12902 ( .IN1(n12918), .IN2(n10972), .QN(n12860) );
  NAND2X0 U12903 ( .IN1(n12919), .IN2(n12878), .QN(n12918) );
  NAND2X0 U12904 ( .IN1(n12920), .IN2(n12921), .QN(n12878) );
  NAND2X0 U12905 ( .IN1(n5290), .IN2(n12849), .QN(n12921) );
  NOR2X0 U12906 ( .IN1(n12850), .IN2(n12922), .QN(n12920) );
  NAND2X0 U12907 ( .IN1(n12922), .IN2(g1585), .QN(n12919) );
  NOR2X0 U12908 ( .IN1(n12923), .IN2(n12924), .QN(n12915) );
  NOR2X0 U12909 ( .IN1(n10136), .IN2(n10898), .QN(n12924) );
  NOR2X0 U12910 ( .IN1(n11046), .IN2(n12925), .QN(n12923) );
  INVX0 U12911 ( .INP(n12926), .ZN(n12925) );
  NOR2X0 U12912 ( .IN1(n12917), .IN2(n5814), .QN(n12926) );
  NOR2X0 U12913 ( .IN1(n12907), .IN2(g2465), .QN(n12917) );
  NAND2X0 U12914 ( .IN1(n12927), .IN2(n12928), .QN(g34007) );
  NAND2X0 U12915 ( .IN1(n11068), .IN2(g2380), .QN(n12928) );
  NOR2X0 U12916 ( .IN1(n12929), .IN2(n12930), .QN(n12927) );
  NOR2X0 U12917 ( .IN1(n10152), .IN2(n11409), .QN(n12930) );
  NOR2X0 U12918 ( .IN1(n12931), .IN2(n12932), .QN(n12929) );
  NAND2X0 U12919 ( .IN1(n12933), .IN2(n12934), .QN(g34006) );
  NAND2X0 U12920 ( .IN1(n12935), .IN2(n12936), .QN(n12934) );
  NOR2X0 U12921 ( .IN1(n10198), .IN2(n12937), .QN(n12936) );
  NOR2X0 U12922 ( .IN1(n12938), .IN2(n12939), .QN(n12935) );
  NOR2X0 U12923 ( .IN1(n12940), .IN2(g2361), .QN(n12939) );
  NOR2X0 U12924 ( .IN1(n12941), .IN2(n12942), .QN(n12933) );
  NOR2X0 U12925 ( .IN1(n11045), .IN2(n12943), .QN(n12942) );
  NOR2X0 U12926 ( .IN1(n12944), .IN2(n12945), .QN(n12943) );
  NOR2X0 U12927 ( .IN1(n10198), .IN2(n12946), .QN(n12945) );
  NOR2X0 U12928 ( .IN1(n12947), .IN2(n12948), .QN(n12944) );
  NOR2X0 U12929 ( .IN1(n12938), .IN2(n12937), .QN(n12948) );
  INVX0 U12930 ( .INP(n12949), .ZN(n12937) );
  NOR2X0 U12931 ( .IN1(g1589), .IN2(n12950), .QN(n12938) );
  NOR2X0 U12932 ( .IN1(n12951), .IN2(n12952), .QN(n12947) );
  NOR2X0 U12933 ( .IN1(n12953), .IN2(g2375), .QN(n12951) );
  NOR2X0 U12934 ( .IN1(n5537), .IN2(n10898), .QN(n12941) );
  NAND2X0 U12935 ( .IN1(n12954), .IN2(n12955), .QN(g34005) );
  INVX0 U12936 ( .INP(n12956), .ZN(n12955) );
  NOR2X0 U12937 ( .IN1(n12957), .IN2(n12931), .QN(n12956) );
  NOR2X0 U12938 ( .IN1(n12958), .IN2(n12959), .QN(n12954) );
  NOR2X0 U12939 ( .IN1(n5794), .IN2(n10898), .QN(n12959) );
  NOR2X0 U12940 ( .IN1(n11045), .IN2(n12960), .QN(n12958) );
  NAND2X0 U12941 ( .IN1(n12957), .IN2(g2315), .QN(n12960) );
  NAND2X0 U12942 ( .IN1(n12961), .IN2(n5513), .QN(n12957) );
  NAND2X0 U12943 ( .IN1(n12962), .IN2(n12963), .QN(g34004) );
  NAND2X0 U12944 ( .IN1(n12964), .IN2(n12965), .QN(n12963) );
  NOR2X0 U12945 ( .IN1(n12966), .IN2(n12967), .QN(n12962) );
  NOR2X0 U12946 ( .IN1(n5802), .IN2(n10898), .QN(n12967) );
  INVX0 U12947 ( .INP(n12968), .ZN(n12966) );
  NAND2X0 U12948 ( .IN1(n10925), .IN2(n12969), .QN(n12968) );
  NOR2X0 U12949 ( .IN1(n12964), .IN2(n19412), .QN(n12969) );
  NOR2X0 U12950 ( .IN1(n12970), .IN2(g2287), .QN(n12964) );
  NAND2X0 U12951 ( .IN1(n12971), .IN2(n12972), .QN(g34003) );
  INVX0 U12952 ( .INP(n12973), .ZN(n12972) );
  NOR2X0 U12953 ( .IN1(n12974), .IN2(n12931), .QN(n12973) );
  NOR2X0 U12954 ( .IN1(n12975), .IN2(n12976), .QN(n12971) );
  NOR2X0 U12955 ( .IN1(n19412), .IN2(n10897), .QN(n12976) );
  NOR2X0 U12956 ( .IN1(n11045), .IN2(n12977), .QN(n12975) );
  NAND2X0 U12957 ( .IN1(n12974), .IN2(g2307), .QN(n12977) );
  NAND2X0 U12958 ( .IN1(n12961), .IN2(g2287), .QN(n12974) );
  NOR2X0 U12959 ( .IN1(n5537), .IN2(n12953), .QN(n12961) );
  NAND2X0 U12960 ( .IN1(n12978), .IN2(n12979), .QN(g34002) );
  NAND2X0 U12961 ( .IN1(n12980), .IN2(n12965), .QN(n12979) );
  NOR2X0 U12962 ( .IN1(n12981), .IN2(n12982), .QN(n12978) );
  NOR2X0 U12963 ( .IN1(n5815), .IN2(n10897), .QN(n12982) );
  INVX0 U12964 ( .INP(n12983), .ZN(n12981) );
  NAND2X0 U12965 ( .IN1(n10925), .IN2(n12984), .QN(n12983) );
  NOR2X0 U12966 ( .IN1(n12980), .IN2(n5794), .QN(n12984) );
  NOR2X0 U12967 ( .IN1(n12970), .IN2(g2361), .QN(n12980) );
  NAND2X0 U12968 ( .IN1(n12985), .IN2(n12986), .QN(g34001) );
  NAND2X0 U12969 ( .IN1(n12987), .IN2(n12965), .QN(n12986) );
  INVX0 U12970 ( .INP(n12931), .ZN(n12965) );
  NAND2X0 U12971 ( .IN1(n12988), .IN2(n10971), .QN(n12931) );
  NAND2X0 U12972 ( .IN1(n12989), .IN2(n12949), .QN(n12988) );
  NAND2X0 U12973 ( .IN1(n12990), .IN2(n12991), .QN(n12949) );
  NAND2X0 U12974 ( .IN1(n5343), .IN2(n12849), .QN(n12991) );
  NOR2X0 U12975 ( .IN1(n12850), .IN2(n12992), .QN(n12990) );
  NAND2X0 U12976 ( .IN1(n5757), .IN2(n12992), .QN(n12989) );
  INVX0 U12977 ( .INP(n12950), .ZN(n12992) );
  NOR2X0 U12978 ( .IN1(n12993), .IN2(n12994), .QN(n12985) );
  NOR2X0 U12979 ( .IN1(n10152), .IN2(n10897), .QN(n12994) );
  NOR2X0 U12980 ( .IN1(n11045), .IN2(n12995), .QN(n12993) );
  INVX0 U12981 ( .INP(n12996), .ZN(n12995) );
  NOR2X0 U12982 ( .IN1(n12987), .IN2(n5815), .QN(n12996) );
  NOR2X0 U12983 ( .IN1(n12997), .IN2(g2331), .QN(n12987) );
  NAND2X0 U12984 ( .IN1(g2287), .IN2(n12946), .QN(n12997) );
  NAND2X0 U12985 ( .IN1(n12998), .IN2(n12999), .QN(g34000) );
  NAND2X0 U12986 ( .IN1(n11068), .IN2(g2246), .QN(n12999) );
  NOR2X0 U12987 ( .IN1(n13000), .IN2(n13001), .QN(n12998) );
  NOR2X0 U12988 ( .IN1(n10158), .IN2(n13002), .QN(n13001) );
  NOR2X0 U12989 ( .IN1(n13003), .IN2(n13004), .QN(n13000) );
  NAND2X0 U12990 ( .IN1(n13005), .IN2(n13006), .QN(g33999) );
  NAND2X0 U12991 ( .IN1(n13007), .IN2(n13008), .QN(n13006) );
  NOR2X0 U12992 ( .IN1(n10200), .IN2(n13009), .QN(n13008) );
  NOR2X0 U12993 ( .IN1(n13010), .IN2(n13011), .QN(n13007) );
  NOR2X0 U12994 ( .IN1(n13012), .IN2(g2227), .QN(n13011) );
  NOR2X0 U12995 ( .IN1(n13013), .IN2(n13014), .QN(n13005) );
  NOR2X0 U12996 ( .IN1(n11045), .IN2(n13015), .QN(n13014) );
  NOR2X0 U12997 ( .IN1(n13016), .IN2(n13017), .QN(n13015) );
  NOR2X0 U12998 ( .IN1(n10200), .IN2(n13018), .QN(n13017) );
  NOR2X0 U12999 ( .IN1(n13019), .IN2(n13020), .QN(n13016) );
  NOR2X0 U13000 ( .IN1(n13010), .IN2(n13009), .QN(n13020) );
  INVX0 U13001 ( .INP(n13021), .ZN(n13009) );
  NOR2X0 U13002 ( .IN1(n13022), .IN2(n5755), .QN(n13010) );
  NOR2X0 U13003 ( .IN1(n13023), .IN2(n13024), .QN(n13019) );
  NOR2X0 U13004 ( .IN1(n13025), .IN2(g2241), .QN(n13023) );
  NOR2X0 U13005 ( .IN1(n5538), .IN2(n10897), .QN(n13013) );
  NAND2X0 U13006 ( .IN1(n13026), .IN2(n13027), .QN(g33998) );
  INVX0 U13007 ( .INP(n13028), .ZN(n13027) );
  NOR2X0 U13008 ( .IN1(n13029), .IN2(n13003), .QN(n13028) );
  NOR2X0 U13009 ( .IN1(n13030), .IN2(n13031), .QN(n13026) );
  NOR2X0 U13010 ( .IN1(n5788), .IN2(n10897), .QN(n13031) );
  NOR2X0 U13011 ( .IN1(n11045), .IN2(n13032), .QN(n13030) );
  NAND2X0 U13012 ( .IN1(n13029), .IN2(g2181), .QN(n13032) );
  NAND2X0 U13013 ( .IN1(n13033), .IN2(n5514), .QN(n13029) );
  NAND2X0 U13014 ( .IN1(n13034), .IN2(n13035), .QN(g33997) );
  NAND2X0 U13015 ( .IN1(n13036), .IN2(n13037), .QN(n13035) );
  NOR2X0 U13016 ( .IN1(n13038), .IN2(n13039), .QN(n13034) );
  NOR2X0 U13017 ( .IN1(n5803), .IN2(n10896), .QN(n13039) );
  INVX0 U13018 ( .INP(n13040), .ZN(n13038) );
  NAND2X0 U13019 ( .IN1(n10924), .IN2(n13041), .QN(n13040) );
  NOR2X0 U13020 ( .IN1(n13036), .IN2(n19408), .QN(n13041) );
  NOR2X0 U13021 ( .IN1(n13042), .IN2(g2153), .QN(n13036) );
  NAND2X0 U13022 ( .IN1(n13043), .IN2(n13044), .QN(g33996) );
  INVX0 U13023 ( .INP(n13045), .ZN(n13044) );
  NOR2X0 U13024 ( .IN1(n13046), .IN2(n13003), .QN(n13045) );
  NOR2X0 U13025 ( .IN1(n13047), .IN2(n13048), .QN(n13043) );
  NOR2X0 U13026 ( .IN1(n19408), .IN2(n10896), .QN(n13048) );
  NOR2X0 U13027 ( .IN1(n11045), .IN2(n13049), .QN(n13047) );
  NAND2X0 U13028 ( .IN1(n13046), .IN2(g2173), .QN(n13049) );
  NAND2X0 U13029 ( .IN1(n13033), .IN2(g2153), .QN(n13046) );
  NOR2X0 U13030 ( .IN1(n5538), .IN2(n13025), .QN(n13033) );
  NAND2X0 U13031 ( .IN1(n13050), .IN2(n13051), .QN(g33995) );
  NAND2X0 U13032 ( .IN1(n13052), .IN2(n13037), .QN(n13051) );
  NOR2X0 U13033 ( .IN1(n13053), .IN2(n13054), .QN(n13050) );
  NOR2X0 U13034 ( .IN1(n5812), .IN2(n10896), .QN(n13054) );
  INVX0 U13035 ( .INP(n13055), .ZN(n13053) );
  NAND2X0 U13036 ( .IN1(n10921), .IN2(n13056), .QN(n13055) );
  NOR2X0 U13037 ( .IN1(n13052), .IN2(n5788), .QN(n13056) );
  NOR2X0 U13038 ( .IN1(n13042), .IN2(g2227), .QN(n13052) );
  NAND2X0 U13039 ( .IN1(n13057), .IN2(n13058), .QN(g33994) );
  NAND2X0 U13040 ( .IN1(n13059), .IN2(n13037), .QN(n13058) );
  INVX0 U13041 ( .INP(n13003), .ZN(n13037) );
  NAND2X0 U13042 ( .IN1(n13060), .IN2(n10970), .QN(n13003) );
  NAND2X0 U13043 ( .IN1(n13061), .IN2(n13021), .QN(n13060) );
  NAND2X0 U13044 ( .IN1(n13062), .IN2(n13063), .QN(n13021) );
  NAND2X0 U13045 ( .IN1(n5289), .IN2(n12849), .QN(n13063) );
  NOR2X0 U13046 ( .IN1(n12850), .IN2(n13064), .QN(n13062) );
  NOR2X0 U13047 ( .IN1(n13065), .IN2(n2549), .QN(n12850) );
  INVX0 U13048 ( .INP(n12849), .ZN(n13065) );
  NOR2X0 U13049 ( .IN1(n13066), .IN2(n5380), .QN(n12849) );
  NAND2X0 U13050 ( .IN1(n13064), .IN2(g1585), .QN(n13061) );
  INVX0 U13051 ( .INP(n13022), .ZN(n13064) );
  NOR2X0 U13052 ( .IN1(n13067), .IN2(n13068), .QN(n13057) );
  NOR2X0 U13053 ( .IN1(n10158), .IN2(n10896), .QN(n13068) );
  NOR2X0 U13054 ( .IN1(n11045), .IN2(n13069), .QN(n13067) );
  INVX0 U13055 ( .INP(n13070), .ZN(n13069) );
  NOR2X0 U13056 ( .IN1(n13059), .IN2(n5812), .QN(n13070) );
  NOR2X0 U13057 ( .IN1(n13071), .IN2(g2197), .QN(n13059) );
  NAND2X0 U13058 ( .IN1(g2153), .IN2(n13018), .QN(n13071) );
  NAND2X0 U13059 ( .IN1(n13072), .IN2(n13073), .QN(g33993) );
  NAND2X0 U13060 ( .IN1(n11068), .IN2(g2089), .QN(n13073) );
  NOR2X0 U13061 ( .IN1(n13074), .IN2(n13075), .QN(n13072) );
  NOR2X0 U13062 ( .IN1(n10217), .IN2(n11443), .QN(n13075) );
  NOR2X0 U13063 ( .IN1(n13076), .IN2(n13077), .QN(n13074) );
  NAND2X0 U13064 ( .IN1(n13078), .IN2(n13079), .QN(g33992) );
  NAND2X0 U13065 ( .IN1(n13080), .IN2(n13081), .QN(n13079) );
  NOR2X0 U13066 ( .IN1(n10195), .IN2(n13082), .QN(n13081) );
  NOR2X0 U13067 ( .IN1(n13083), .IN2(n13084), .QN(n13080) );
  NOR2X0 U13068 ( .IN1(n13085), .IN2(g2070), .QN(n13083) );
  NOR2X0 U13069 ( .IN1(n5355), .IN2(n11014), .QN(n13085) );
  NOR2X0 U13070 ( .IN1(n13086), .IN2(n13087), .QN(n13078) );
  NOR2X0 U13071 ( .IN1(n11045), .IN2(n13088), .QN(n13087) );
  NOR2X0 U13072 ( .IN1(n13089), .IN2(n13090), .QN(n13088) );
  NOR2X0 U13073 ( .IN1(n10195), .IN2(n13091), .QN(n13090) );
  NOR2X0 U13074 ( .IN1(n13092), .IN2(n13093), .QN(n13089) );
  NOR2X0 U13075 ( .IN1(n13084), .IN2(n13082), .QN(n13093) );
  INVX0 U13076 ( .INP(n13094), .ZN(n13082) );
  NOR2X0 U13077 ( .IN1(g1246), .IN2(n13095), .QN(n13084) );
  NOR2X0 U13078 ( .IN1(n13096), .IN2(n13097), .QN(n13092) );
  NOR2X0 U13079 ( .IN1(n13098), .IN2(g2084), .QN(n13096) );
  NOR2X0 U13080 ( .IN1(n5535), .IN2(n10896), .QN(n13086) );
  NAND2X0 U13081 ( .IN1(n13099), .IN2(n13100), .QN(g33991) );
  INVX0 U13082 ( .INP(n13101), .ZN(n13100) );
  NOR2X0 U13083 ( .IN1(n13102), .IN2(n13076), .QN(n13101) );
  NOR2X0 U13084 ( .IN1(n13103), .IN2(n13104), .QN(n13099) );
  NOR2X0 U13085 ( .IN1(n5790), .IN2(n10895), .QN(n13104) );
  NOR2X0 U13086 ( .IN1(n11045), .IN2(n13105), .QN(n13103) );
  NAND2X0 U13087 ( .IN1(n13102), .IN2(g2024), .QN(n13105) );
  NAND2X0 U13088 ( .IN1(n12491), .IN2(n13091), .QN(n13102) );
  NAND2X0 U13089 ( .IN1(n13106), .IN2(n13107), .QN(g33990) );
  NAND2X0 U13090 ( .IN1(n13108), .IN2(n13109), .QN(n13107) );
  NOR2X0 U13091 ( .IN1(n13110), .IN2(n13111), .QN(n13106) );
  NOR2X0 U13092 ( .IN1(n5801), .IN2(n10895), .QN(n13111) );
  NOR2X0 U13093 ( .IN1(n11045), .IN2(n13112), .QN(n13110) );
  INVX0 U13094 ( .INP(n13113), .ZN(n13112) );
  NOR2X0 U13095 ( .IN1(n13108), .IN2(n19413), .QN(n13113) );
  NOR2X0 U13096 ( .IN1(n13114), .IN2(g1996), .QN(n13108) );
  NAND2X0 U13097 ( .IN1(n13115), .IN2(n13116), .QN(g33989) );
  NAND2X0 U13098 ( .IN1(n13117), .IN2(n13109), .QN(n13116) );
  NOR2X0 U13099 ( .IN1(n13118), .IN2(n13119), .QN(n13115) );
  NOR2X0 U13100 ( .IN1(n19413), .IN2(n10895), .QN(n13119) );
  NOR2X0 U13101 ( .IN1(n11045), .IN2(n13120), .QN(n13118) );
  NAND2X0 U13102 ( .IN1(n13121), .IN2(g2016), .QN(n13120) );
  INVX0 U13103 ( .INP(n13117), .ZN(n13121) );
  NOR2X0 U13104 ( .IN1(n13122), .IN2(n5535), .QN(n13117) );
  NAND2X0 U13105 ( .IN1(n13123), .IN2(n13124), .QN(g33988) );
  NAND2X0 U13106 ( .IN1(n13125), .IN2(n13109), .QN(n13124) );
  NOR2X0 U13107 ( .IN1(n13126), .IN2(n13127), .QN(n13123) );
  NOR2X0 U13108 ( .IN1(n5818), .IN2(n10895), .QN(n13127) );
  NOR2X0 U13109 ( .IN1(n11044), .IN2(n13128), .QN(n13126) );
  INVX0 U13110 ( .INP(n13129), .ZN(n13128) );
  NOR2X0 U13111 ( .IN1(n13125), .IN2(n5790), .QN(n13129) );
  NOR2X0 U13112 ( .IN1(n13114), .IN2(g2070), .QN(n13125) );
  NAND2X0 U13113 ( .IN1(n13130), .IN2(n13131), .QN(g33987) );
  NAND2X0 U13114 ( .IN1(n13132), .IN2(n13109), .QN(n13131) );
  INVX0 U13115 ( .INP(n13076), .ZN(n13109) );
  NAND2X0 U13116 ( .IN1(n13133), .IN2(n10969), .QN(n13076) );
  NAND2X0 U13117 ( .IN1(n13134), .IN2(n13094), .QN(n13133) );
  NAND2X0 U13118 ( .IN1(n13135), .IN2(n13136), .QN(n13094) );
  NAND2X0 U13119 ( .IN1(n5341), .IN2(n13137), .QN(n13136) );
  NOR2X0 U13120 ( .IN1(n13138), .IN2(n13139), .QN(n13135) );
  NAND2X0 U13121 ( .IN1(n5526), .IN2(n13139), .QN(n13134) );
  INVX0 U13122 ( .INP(n13095), .ZN(n13139) );
  NOR2X0 U13123 ( .IN1(n13140), .IN2(n13141), .QN(n13130) );
  NOR2X0 U13124 ( .IN1(n10217), .IN2(n10894), .QN(n13141) );
  NOR2X0 U13125 ( .IN1(n11044), .IN2(n13142), .QN(n13140) );
  INVX0 U13126 ( .INP(n13143), .ZN(n13142) );
  NOR2X0 U13127 ( .IN1(n13132), .IN2(n5818), .QN(n13143) );
  NOR2X0 U13128 ( .IN1(n13122), .IN2(g2040), .QN(n13132) );
  INVX0 U13129 ( .INP(n13144), .ZN(n13122) );
  NAND2X0 U13130 ( .IN1(n13145), .IN2(n13146), .QN(g33986) );
  NAND2X0 U13131 ( .IN1(n11068), .IN2(g1955), .QN(n13146) );
  NOR2X0 U13132 ( .IN1(n13147), .IN2(n13148), .QN(n13145) );
  NOR2X0 U13133 ( .IN1(n10144), .IN2(n11486), .QN(n13148) );
  NOR2X0 U13134 ( .IN1(n13149), .IN2(n13150), .QN(n13147) );
  NAND2X0 U13135 ( .IN1(n13151), .IN2(n13152), .QN(g33985) );
  NAND2X0 U13136 ( .IN1(n13153), .IN2(n13154), .QN(n13152) );
  NOR2X0 U13137 ( .IN1(n10199), .IN2(n13155), .QN(n13154) );
  NOR2X0 U13138 ( .IN1(n13156), .IN2(n13157), .QN(n13153) );
  NOR2X0 U13139 ( .IN1(n13158), .IN2(g1936), .QN(n13157) );
  NOR2X0 U13140 ( .IN1(n11044), .IN2(n10657), .QN(n13158) );
  NOR2X0 U13141 ( .IN1(n13159), .IN2(n13160), .QN(n13151) );
  NOR2X0 U13142 ( .IN1(n11044), .IN2(n13161), .QN(n13160) );
  NOR2X0 U13143 ( .IN1(n13162), .IN2(n13163), .QN(n13161) );
  NOR2X0 U13144 ( .IN1(n10199), .IN2(n13164), .QN(n13163) );
  NOR2X0 U13145 ( .IN1(n13165), .IN2(n13166), .QN(n13162) );
  NOR2X0 U13146 ( .IN1(n13156), .IN2(n13155), .QN(n13166) );
  INVX0 U13147 ( .INP(n13167), .ZN(n13155) );
  NOR2X0 U13148 ( .IN1(n13168), .IN2(n5756), .QN(n13156) );
  NOR2X0 U13149 ( .IN1(n13169), .IN2(n13170), .QN(n13165) );
  NOR2X0 U13150 ( .IN1(n13171), .IN2(g1950), .QN(n13169) );
  NOR2X0 U13151 ( .IN1(n5534), .IN2(n10894), .QN(n13159) );
  NAND2X0 U13152 ( .IN1(n13172), .IN2(n13173), .QN(g33984) );
  NAND2X0 U13153 ( .IN1(n13174), .IN2(n13175), .QN(n13173) );
  NOR2X0 U13154 ( .IN1(n13176), .IN2(n13177), .QN(n13172) );
  NOR2X0 U13155 ( .IN1(n5793), .IN2(n10860), .QN(n13177) );
  NOR2X0 U13156 ( .IN1(n11044), .IN2(n13178), .QN(n13176) );
  NAND2X0 U13157 ( .IN1(n13179), .IN2(g1890), .QN(n13178) );
  INVX0 U13158 ( .INP(n13174), .ZN(n13179) );
  NOR2X0 U13159 ( .IN1(n12495), .IN2(n13171), .QN(n13174) );
  NAND2X0 U13160 ( .IN1(n13180), .IN2(n13181), .QN(g33983) );
  NAND2X0 U13161 ( .IN1(n13182), .IN2(n13175), .QN(n13181) );
  NOR2X0 U13162 ( .IN1(n13183), .IN2(n13184), .QN(n13180) );
  NOR2X0 U13163 ( .IN1(n5799), .IN2(n10859), .QN(n13184) );
  NOR2X0 U13164 ( .IN1(n11044), .IN2(n13185), .QN(n13183) );
  INVX0 U13165 ( .INP(n13186), .ZN(n13185) );
  NOR2X0 U13166 ( .IN1(n13182), .IN2(n19415), .QN(n13186) );
  NOR2X0 U13167 ( .IN1(n13187), .IN2(test_so8), .QN(n13182) );
  NAND2X0 U13168 ( .IN1(n13188), .IN2(n13189), .QN(g33982) );
  NAND2X0 U13169 ( .IN1(n13190), .IN2(n13175), .QN(n13189) );
  NOR2X0 U13170 ( .IN1(n13191), .IN2(n13192), .QN(n13188) );
  NOR2X0 U13171 ( .IN1(n19415), .IN2(n10859), .QN(n13192) );
  INVX0 U13172 ( .INP(n13193), .ZN(n13191) );
  NAND2X0 U13173 ( .IN1(n10920), .IN2(n13194), .QN(n13193) );
  NOR2X0 U13174 ( .IN1(n13190), .IN2(n5854), .QN(n13194) );
  NOR2X0 U13175 ( .IN1(n13195), .IN2(n5534), .QN(n13190) );
  NAND2X0 U13176 ( .IN1(n13196), .IN2(n13197), .QN(g33981) );
  NAND2X0 U13177 ( .IN1(n13198), .IN2(n13175), .QN(n13197) );
  NOR2X0 U13178 ( .IN1(n13199), .IN2(n13200), .QN(n13196) );
  NOR2X0 U13179 ( .IN1(n5813), .IN2(n10859), .QN(n13200) );
  NOR2X0 U13180 ( .IN1(n11044), .IN2(n13201), .QN(n13199) );
  INVX0 U13181 ( .INP(n13202), .ZN(n13201) );
  NOR2X0 U13182 ( .IN1(n13198), .IN2(n5793), .QN(n13202) );
  NOR2X0 U13183 ( .IN1(n13187), .IN2(g1936), .QN(n13198) );
  NAND2X0 U13184 ( .IN1(n13203), .IN2(n13204), .QN(g33980) );
  NAND2X0 U13185 ( .IN1(n13205), .IN2(n13175), .QN(n13204) );
  INVX0 U13186 ( .INP(n13149), .ZN(n13175) );
  NAND2X0 U13187 ( .IN1(n13206), .IN2(n10968), .QN(n13149) );
  NAND2X0 U13188 ( .IN1(n13207), .IN2(n13167), .QN(n13206) );
  NAND2X0 U13189 ( .IN1(n13208), .IN2(n13209), .QN(n13167) );
  NAND2X0 U13190 ( .IN1(n5329), .IN2(n13137), .QN(n13209) );
  NOR2X0 U13191 ( .IN1(n13138), .IN2(n13210), .QN(n13208) );
  NAND2X0 U13192 ( .IN1(n13210), .IN2(g30332), .QN(n13207) );
  NOR2X0 U13193 ( .IN1(n13211), .IN2(n13212), .QN(n13203) );
  NOR2X0 U13194 ( .IN1(n10144), .IN2(n10859), .QN(n13212) );
  NOR2X0 U13195 ( .IN1(n11044), .IN2(n13213), .QN(n13211) );
  INVX0 U13196 ( .INP(n13214), .ZN(n13213) );
  NOR2X0 U13197 ( .IN1(n13205), .IN2(n5813), .QN(n13214) );
  NOR2X0 U13198 ( .IN1(n13195), .IN2(g1906), .QN(n13205) );
  NAND2X0 U13199 ( .IN1(n13215), .IN2(n13216), .QN(g33979) );
  NAND2X0 U13200 ( .IN1(n11068), .IN2(g1821), .QN(n13216) );
  NOR2X0 U13201 ( .IN1(n13217), .IN2(n13218), .QN(n13215) );
  NOR2X0 U13202 ( .IN1(n10208), .IN2(n11324), .QN(n13218) );
  NOR2X0 U13203 ( .IN1(n13219), .IN2(n13220), .QN(n13217) );
  NAND2X0 U13204 ( .IN1(n13221), .IN2(n13222), .QN(g33978) );
  NAND2X0 U13205 ( .IN1(n13223), .IN2(n13224), .QN(n13222) );
  NOR2X0 U13206 ( .IN1(n10128), .IN2(n13225), .QN(n13224) );
  NOR2X0 U13207 ( .IN1(n13226), .IN2(n13227), .QN(n13223) );
  NOR2X0 U13208 ( .IN1(n13228), .IN2(g1802), .QN(n13227) );
  NOR2X0 U13209 ( .IN1(n13229), .IN2(n13230), .QN(n13221) );
  NOR2X0 U13210 ( .IN1(n11044), .IN2(n13231), .QN(n13230) );
  NOR2X0 U13211 ( .IN1(n13232), .IN2(n13233), .QN(n13231) );
  NOR2X0 U13212 ( .IN1(n10128), .IN2(n13234), .QN(n13233) );
  NOR2X0 U13213 ( .IN1(n13235), .IN2(n13236), .QN(n13232) );
  NOR2X0 U13214 ( .IN1(n13226), .IN2(n13225), .QN(n13236) );
  INVX0 U13215 ( .INP(n13237), .ZN(n13225) );
  NOR2X0 U13216 ( .IN1(g1246), .IN2(n13238), .QN(n13226) );
  NOR2X0 U13217 ( .IN1(n13239), .IN2(n13240), .QN(n13235) );
  NOR2X0 U13218 ( .IN1(n13241), .IN2(g1816), .QN(n13239) );
  NOR2X0 U13219 ( .IN1(n5536), .IN2(n10858), .QN(n13229) );
  NAND2X0 U13220 ( .IN1(n13242), .IN2(n13243), .QN(g33977) );
  INVX0 U13221 ( .INP(n13244), .ZN(n13243) );
  NOR2X0 U13222 ( .IN1(n13245), .IN2(n13219), .QN(n13244) );
  NOR2X0 U13223 ( .IN1(n13246), .IN2(n13247), .QN(n13242) );
  NOR2X0 U13224 ( .IN1(n5795), .IN2(n10857), .QN(n13247) );
  NOR2X0 U13225 ( .IN1(n11044), .IN2(n13248), .QN(n13246) );
  NAND2X0 U13226 ( .IN1(n13245), .IN2(g1756), .QN(n13248) );
  NAND2X0 U13227 ( .IN1(n13249), .IN2(n5504), .QN(n13245) );
  NAND2X0 U13228 ( .IN1(n13250), .IN2(n13251), .QN(g33976) );
  NAND2X0 U13229 ( .IN1(n13252), .IN2(n13253), .QN(n13251) );
  NOR2X0 U13230 ( .IN1(n13254), .IN2(n13255), .QN(n13250) );
  NOR2X0 U13231 ( .IN1(n5804), .IN2(n10899), .QN(n13255) );
  INVX0 U13232 ( .INP(n13256), .ZN(n13254) );
  NAND2X0 U13233 ( .IN1(n10922), .IN2(n13257), .QN(n13256) );
  NOR2X0 U13234 ( .IN1(n13252), .IN2(n5797), .QN(n13257) );
  NOR2X0 U13235 ( .IN1(n13258), .IN2(g1728), .QN(n13252) );
  NAND2X0 U13236 ( .IN1(n13259), .IN2(n13260), .QN(g33975) );
  INVX0 U13237 ( .INP(n13261), .ZN(n13260) );
  NOR2X0 U13238 ( .IN1(n13262), .IN2(n13219), .QN(n13261) );
  NOR2X0 U13239 ( .IN1(n13263), .IN2(n13264), .QN(n13259) );
  NOR2X0 U13240 ( .IN1(n5797), .IN2(n10856), .QN(n13264) );
  NOR2X0 U13241 ( .IN1(n11044), .IN2(n13265), .QN(n13263) );
  NAND2X0 U13242 ( .IN1(n13262), .IN2(g1748), .QN(n13265) );
  NAND2X0 U13243 ( .IN1(n13249), .IN2(g1728), .QN(n13262) );
  NOR2X0 U13244 ( .IN1(n5536), .IN2(n13241), .QN(n13249) );
  NAND2X0 U13245 ( .IN1(n13266), .IN2(n13267), .QN(g33974) );
  NAND2X0 U13246 ( .IN1(n13268), .IN2(n13253), .QN(n13267) );
  NOR2X0 U13247 ( .IN1(n13269), .IN2(n13270), .QN(n13266) );
  NOR2X0 U13248 ( .IN1(n5817), .IN2(n10856), .QN(n13270) );
  INVX0 U13249 ( .INP(n13271), .ZN(n13269) );
  NAND2X0 U13250 ( .IN1(n10925), .IN2(n13272), .QN(n13271) );
  NOR2X0 U13251 ( .IN1(n13268), .IN2(n5795), .QN(n13272) );
  NOR2X0 U13252 ( .IN1(n13258), .IN2(g1802), .QN(n13268) );
  NAND2X0 U13253 ( .IN1(n13273), .IN2(n13274), .QN(g33973) );
  NAND2X0 U13254 ( .IN1(n13275), .IN2(n13253), .QN(n13274) );
  INVX0 U13255 ( .INP(n13219), .ZN(n13253) );
  NAND2X0 U13256 ( .IN1(n13276), .IN2(n10967), .QN(n13219) );
  NAND2X0 U13257 ( .IN1(n13277), .IN2(n13237), .QN(n13276) );
  NAND2X0 U13258 ( .IN1(n13278), .IN2(n13279), .QN(n13237) );
  NAND2X0 U13259 ( .IN1(n5478), .IN2(n13137), .QN(n13279) );
  NOR2X0 U13260 ( .IN1(n13138), .IN2(n13280), .QN(n13278) );
  NAND2X0 U13261 ( .IN1(n5526), .IN2(n13280), .QN(n13277) );
  NOR2X0 U13262 ( .IN1(n13281), .IN2(n13282), .QN(n13273) );
  NOR2X0 U13263 ( .IN1(n10208), .IN2(n10856), .QN(n13282) );
  NOR2X0 U13264 ( .IN1(n11043), .IN2(n13283), .QN(n13281) );
  INVX0 U13265 ( .INP(n13284), .ZN(n13283) );
  NOR2X0 U13266 ( .IN1(n13275), .IN2(n5817), .QN(n13284) );
  NOR2X0 U13267 ( .IN1(n13285), .IN2(g1772), .QN(n13275) );
  NAND2X0 U13268 ( .IN1(g1728), .IN2(n13234), .QN(n13285) );
  NAND2X0 U13269 ( .IN1(n13286), .IN2(n13287), .QN(g33972) );
  NAND2X0 U13270 ( .IN1(n11067), .IN2(g1687), .QN(n13287) );
  NOR2X0 U13271 ( .IN1(n13288), .IN2(n13289), .QN(n13286) );
  NOR2X0 U13272 ( .IN1(n10135), .IN2(n13290), .QN(n13289) );
  NOR2X0 U13273 ( .IN1(n13291), .IN2(n13292), .QN(n13288) );
  NAND2X0 U13274 ( .IN1(n13293), .IN2(n13294), .QN(g33971) );
  NAND2X0 U13275 ( .IN1(n13295), .IN2(n13296), .QN(n13294) );
  NOR2X0 U13276 ( .IN1(n10201), .IN2(n13297), .QN(n13296) );
  NOR2X0 U13277 ( .IN1(n13298), .IN2(n13299), .QN(n13295) );
  NOR2X0 U13278 ( .IN1(n13300), .IN2(g1668), .QN(n13299) );
  NOR2X0 U13279 ( .IN1(n5362), .IN2(n11015), .QN(n13300) );
  NOR2X0 U13280 ( .IN1(n13301), .IN2(n13302), .QN(n13293) );
  NOR2X0 U13281 ( .IN1(n11043), .IN2(n13303), .QN(n13302) );
  NOR2X0 U13282 ( .IN1(n13304), .IN2(n13305), .QN(n13303) );
  NOR2X0 U13283 ( .IN1(n10201), .IN2(n13306), .QN(n13305) );
  NOR2X0 U13284 ( .IN1(n13307), .IN2(n13308), .QN(n13304) );
  NOR2X0 U13285 ( .IN1(n13298), .IN2(n13297), .QN(n13308) );
  INVX0 U13286 ( .INP(n13309), .ZN(n13297) );
  NOR2X0 U13287 ( .IN1(n13310), .IN2(n5756), .QN(n13298) );
  NOR2X0 U13288 ( .IN1(n13311), .IN2(n13312), .QN(n13307) );
  NOR2X0 U13289 ( .IN1(n13313), .IN2(g1682), .QN(n13311) );
  NOR2X0 U13290 ( .IN1(n5598), .IN2(n10855), .QN(n13301) );
  NAND2X0 U13291 ( .IN1(n13314), .IN2(n13315), .QN(g33970) );
  NAND2X0 U13292 ( .IN1(n13316), .IN2(n13317), .QN(n13315) );
  INVX0 U13293 ( .INP(n13318), .ZN(n13316) );
  NOR2X0 U13294 ( .IN1(n13319), .IN2(n13320), .QN(n13314) );
  NOR2X0 U13295 ( .IN1(n5792), .IN2(n10855), .QN(n13320) );
  NOR2X0 U13296 ( .IN1(n11043), .IN2(n13321), .QN(n13319) );
  NAND2X0 U13297 ( .IN1(n13318), .IN2(g1620), .QN(n13321) );
  NAND2X0 U13298 ( .IN1(g31862), .IN2(n13306), .QN(n13318) );
  NAND2X0 U13299 ( .IN1(n13322), .IN2(n13323), .QN(g33969) );
  NAND2X0 U13300 ( .IN1(n13324), .IN2(n13317), .QN(n13323) );
  NOR2X0 U13301 ( .IN1(n13325), .IN2(n13326), .QN(n13322) );
  NOR2X0 U13302 ( .IN1(n5791), .IN2(n10855), .QN(n13326) );
  NOR2X0 U13303 ( .IN1(n11043), .IN2(n13327), .QN(n13325) );
  INVX0 U13304 ( .INP(n13328), .ZN(n13327) );
  NOR2X0 U13305 ( .IN1(n13324), .IN2(n19414), .QN(n13328) );
  NOR2X0 U13306 ( .IN1(n13329), .IN2(g1592), .QN(n13324) );
  NAND2X0 U13307 ( .IN1(n13330), .IN2(n13331), .QN(g33968) );
  NAND2X0 U13308 ( .IN1(n13332), .IN2(n13317), .QN(n13331) );
  INVX0 U13309 ( .INP(n13333), .ZN(n13332) );
  NOR2X0 U13310 ( .IN1(n13334), .IN2(n13335), .QN(n13330) );
  NOR2X0 U13311 ( .IN1(n19414), .IN2(n10854), .QN(n13335) );
  NOR2X0 U13312 ( .IN1(n11043), .IN2(n13336), .QN(n13334) );
  NAND2X0 U13313 ( .IN1(n13333), .IN2(g1612), .QN(n13336) );
  NAND2X0 U13314 ( .IN1(n13337), .IN2(g1668), .QN(n13333) );
  NAND2X0 U13315 ( .IN1(n13338), .IN2(n13339), .QN(g33967) );
  NAND2X0 U13316 ( .IN1(n13340), .IN2(n13317), .QN(n13339) );
  NOR2X0 U13317 ( .IN1(n13341), .IN2(n13342), .QN(n13338) );
  NOR2X0 U13318 ( .IN1(n5811), .IN2(n10854), .QN(n13342) );
  NOR2X0 U13319 ( .IN1(n11043), .IN2(n13343), .QN(n13341) );
  INVX0 U13320 ( .INP(n13344), .ZN(n13343) );
  NOR2X0 U13321 ( .IN1(n13340), .IN2(n5792), .QN(n13344) );
  NOR2X0 U13322 ( .IN1(n13329), .IN2(g1668), .QN(n13340) );
  NAND2X0 U13323 ( .IN1(n13345), .IN2(n13346), .QN(g33966) );
  NAND2X0 U13324 ( .IN1(n13347), .IN2(n13317), .QN(n13346) );
  INVX0 U13325 ( .INP(n13291), .ZN(n13317) );
  NAND2X0 U13326 ( .IN1(n13348), .IN2(n10966), .QN(n13291) );
  NAND2X0 U13327 ( .IN1(n13349), .IN2(n13309), .QN(n13348) );
  NAND2X0 U13328 ( .IN1(n13350), .IN2(n13351), .QN(n13309) );
  NAND2X0 U13329 ( .IN1(n5328), .IN2(n13137), .QN(n13351) );
  NOR2X0 U13330 ( .IN1(n13138), .IN2(n13352), .QN(n13350) );
  INVX0 U13331 ( .INP(n13353), .ZN(n13138) );
  NAND2X0 U13332 ( .IN1(n13137), .IN2(g947), .QN(n13353) );
  NOR2X0 U13333 ( .IN1(n13354), .IN2(n5380), .QN(n13137) );
  NAND2X0 U13334 ( .IN1(n13352), .IN2(g30332), .QN(n13349) );
  INVX0 U13335 ( .INP(n13310), .ZN(n13352) );
  INVX0 U13336 ( .INP(n13355), .ZN(n13347) );
  NOR2X0 U13337 ( .IN1(n13356), .IN2(n13357), .QN(n13345) );
  NOR2X0 U13338 ( .IN1(n10135), .IN2(n10854), .QN(n13357) );
  NOR2X0 U13339 ( .IN1(n11043), .IN2(n13358), .QN(n13356) );
  NAND2X0 U13340 ( .IN1(n13355), .IN2(g1600), .QN(n13358) );
  NAND2X0 U13341 ( .IN1(n13337), .IN2(n5549), .QN(n13355) );
  NAND2X0 U13342 ( .IN1(n13359), .IN2(n13360), .QN(g33965) );
  NAND2X0 U13343 ( .IN1(n11067), .IN2(g763), .QN(n13360) );
  NOR2X0 U13344 ( .IN1(n13361), .IN2(n13362), .QN(n13359) );
  NOR2X0 U13345 ( .IN1(g767), .IN2(n13363), .QN(n13362) );
  NOR2X0 U13346 ( .IN1(n5333), .IN2(n13364), .QN(n13361) );
  NAND2X0 U13347 ( .IN1(n2404), .IN2(n13363), .QN(n13364) );
  INVX0 U13348 ( .INP(n2704), .ZN(n13363) );
  NAND2X0 U13349 ( .IN1(n13365), .IN2(n13366), .QN(g33964) );
  NAND2X0 U13350 ( .IN1(n11067), .IN2(g595), .QN(n13366) );
  NOR2X0 U13351 ( .IN1(n13367), .IN2(n13368), .QN(n13365) );
  NOR2X0 U13352 ( .IN1(g599), .IN2(n13369), .QN(n13368) );
  NOR2X0 U13353 ( .IN1(n5550), .IN2(n13370), .QN(n13367) );
  NAND2X0 U13354 ( .IN1(n2421), .IN2(n13369), .QN(n13370) );
  INVX0 U13355 ( .INP(n2706), .ZN(n13369) );
  NAND2X0 U13356 ( .IN1(n13371), .IN2(n13372), .QN(g33963) );
  NAND2X0 U13357 ( .IN1(n11067), .IN2(g29215), .QN(n13372) );
  NAND2X0 U13358 ( .IN1(n13373), .IN2(n10966), .QN(n13371) );
  NOR2X0 U13359 ( .IN1(n13374), .IN2(n13375), .QN(n13373) );
  NOR2X0 U13360 ( .IN1(n13376), .IN2(n13377), .QN(n13375) );
  NOR2X0 U13361 ( .IN1(g72), .IN2(n10275), .QN(n13376) );
  NOR2X0 U13362 ( .IN1(n13378), .IN2(n13379), .QN(n13374) );
  NAND2X0 U13363 ( .IN1(n13380), .IN2(n11433), .QN(n13379) );
  NAND2X0 U13364 ( .IN1(n13381), .IN2(g269), .QN(n13380) );
  NOR2X0 U13365 ( .IN1(n10276), .IN2(n13382), .QN(n13378) );
  NAND2X0 U13366 ( .IN1(n13383), .IN2(n13384), .QN(g33962) );
  NAND2X0 U13367 ( .IN1(n11067), .IN2(g479), .QN(n13384) );
  NAND2X0 U13368 ( .IN1(n13385), .IN2(n10966), .QN(n13383) );
  NOR2X0 U13369 ( .IN1(n13386), .IN2(n13387), .QN(n13385) );
  NAND2X0 U13370 ( .IN1(n13388), .IN2(n13389), .QN(n13387) );
  NAND2X0 U13371 ( .IN1(n13390), .IN2(g73), .QN(n13389) );
  NOR2X0 U13372 ( .IN1(g225), .IN2(n13381), .QN(n13390) );
  NAND2X0 U13373 ( .IN1(n13391), .IN2(n13382), .QN(n13388) );
  NAND2X0 U13374 ( .IN1(n13392), .IN2(n13393), .QN(n13391) );
  NAND2X0 U13375 ( .IN1(g73), .IN2(n10399), .QN(n13393) );
  NOR2X0 U13376 ( .IN1(g239), .IN2(n13392), .QN(n13386) );
  NAND2X0 U13377 ( .IN1(n11433), .IN2(n13394), .QN(n13392) );
  NAND2X0 U13378 ( .IN1(n13381), .IN2(g246), .QN(n13394) );
  NAND2X0 U13379 ( .IN1(n13395), .IN2(n13396), .QN(g33961) );
  NAND2X0 U13380 ( .IN1(n11067), .IN2(g294), .QN(n13396) );
  NOR2X0 U13381 ( .IN1(n13397), .IN2(n13398), .QN(n13395) );
  NOR2X0 U13382 ( .IN1(g298), .IN2(n13399), .QN(n13398) );
  NOR2X0 U13383 ( .IN1(n5675), .IN2(n13400), .QN(n13397) );
  NAND2X0 U13384 ( .IN1(n95), .IN2(n13399), .QN(n13400) );
  INVX0 U13385 ( .INP(n2989), .ZN(n13399) );
  NAND2X0 U13386 ( .IN1(n13401), .IN2(n13402), .QN(g33960) );
  NAND2X0 U13387 ( .IN1(n11065), .IN2(g153), .QN(n13402) );
  NOR2X0 U13388 ( .IN1(n13403), .IN2(n13404), .QN(n13401) );
  NOR2X0 U13389 ( .IN1(g157), .IN2(n13405), .QN(n13404) );
  NOR2X0 U13390 ( .IN1(n5678), .IN2(n13406), .QN(n13403) );
  NAND2X0 U13391 ( .IN1(n12641), .IN2(n13405), .QN(n13406) );
  INVX0 U13392 ( .INP(n2991), .ZN(n13405) );
  NAND2X0 U13393 ( .IN1(n13407), .IN2(n13408), .QN(g33935) );
  NOR2X0 U13394 ( .IN1(n10220), .IN2(n10219), .QN(n13408) );
  NOR2X0 U13395 ( .IN1(g34649), .IN2(n12534), .QN(n13407) );
  NAND2X0 U13396 ( .IN1(n13409), .IN2(n13410), .QN(g34649) );
  NOR2X0 U13397 ( .IN1(n13411), .IN2(n13412), .QN(n13410) );
  NOR2X0 U13398 ( .IN1(n5614), .IN2(n11391), .QN(n13412) );
  NOR2X0 U13399 ( .IN1(n5863), .IN2(n11399), .QN(n13411) );
  NOR2X0 U13400 ( .IN1(n13413), .IN2(n13414), .QN(n13409) );
  NOR2X0 U13401 ( .IN1(n5878), .IN2(n11402), .QN(n13414) );
  NOR2X0 U13402 ( .IN1(n5875), .IN2(n11403), .QN(n13413) );
  NAND2X0 U13403 ( .IN1(n13415), .IN2(n5541), .QN(g33874) );
  NOR2X0 U13404 ( .IN1(n5846), .IN2(n12534), .QN(n13415) );
  NAND2X0 U13405 ( .IN1(n13416), .IN2(n13417), .QN(g33659) );
  INVX0 U13406 ( .INP(n11413), .ZN(n13417) );
  NAND2X0 U13407 ( .IN1(n13418), .IN2(n13419), .QN(n11413) );
  XOR2X1 U13408 ( .IN1(g4108), .IN2(n13382), .Q(n13419) );
  XOR2X1 U13409 ( .IN1(n10403), .IN2(g73), .Q(n13418) );
  NOR2X0 U13410 ( .IN1(n12456), .IN2(n13420), .QN(n13416) );
  NAND2X0 U13411 ( .IN1(n13421), .IN2(n13422), .QN(n13420) );
  NAND2X0 U13412 ( .IN1(n5350), .IN2(n11505), .QN(n13422) );
  NAND2X0 U13413 ( .IN1(n13423), .IN2(n13424), .QN(n11505) );
  NAND2X0 U13414 ( .IN1(n13425), .IN2(n13426), .QN(n13424) );
  NOR2X0 U13415 ( .IN1(n13427), .IN2(n13428), .QN(n13423) );
  NOR2X0 U13416 ( .IN1(n12428), .IN2(n13429), .QN(n13428) );
  NOR2X0 U13417 ( .IN1(n5340), .IN2(n13430), .QN(n13427) );
  NAND2X0 U13418 ( .IN1(n13431), .IN2(n13432), .QN(n13430) );
  NAND2X0 U13419 ( .IN1(n5480), .IN2(n13433), .QN(n13432) );
  NAND2X0 U13420 ( .IN1(n13434), .IN2(g4087), .QN(n13431) );
  NAND2X0 U13421 ( .IN1(n11504), .IN2(g4098), .QN(n13421) );
  NAND2X0 U13422 ( .IN1(n13435), .IN2(n13436), .QN(n11504) );
  NAND2X0 U13423 ( .IN1(n13437), .IN2(n13425), .QN(n13436) );
  NOR2X0 U13424 ( .IN1(n13438), .IN2(n13439), .QN(n13435) );
  NOR2X0 U13425 ( .IN1(n12428), .IN2(n13440), .QN(n13439) );
  NOR2X0 U13426 ( .IN1(n5340), .IN2(n13441), .QN(n13438) );
  NAND2X0 U13427 ( .IN1(n13442), .IN2(n13443), .QN(n13441) );
  NAND2X0 U13428 ( .IN1(n5480), .IN2(n13444), .QN(n13443) );
  NAND2X0 U13429 ( .IN1(n13445), .IN2(g4087), .QN(n13442) );
  NAND2X0 U13430 ( .IN1(g113), .IN2(n1363), .QN(n12456) );
  INVX0 U13431 ( .INP(n12534), .ZN(n1363) );
  NAND2X0 U13432 ( .IN1(n13446), .IN2(n13447), .QN(g33636) );
  NOR2X0 U13433 ( .IN1(n10222), .IN2(n10221), .QN(n13447) );
  NOR2X0 U13434 ( .IN1(g34657), .IN2(n12534), .QN(n13446) );
  NOR2X0 U13435 ( .IN1(n13448), .IN2(g134), .QN(n12534) );
  INVX0 U13436 ( .INP(n13449), .ZN(n13448) );
  NAND2X0 U13437 ( .IN1(g99), .IN2(g37), .QN(n13449) );
  NAND2X0 U13438 ( .IN1(n13450), .IN2(n13451), .QN(g34657) );
  NOR2X0 U13439 ( .IN1(n13452), .IN2(n13453), .QN(n13451) );
  NOR2X0 U13440 ( .IN1(n13454), .IN2(n13455), .QN(n13450) );
  NAND2X0 U13441 ( .IN1(n13456), .IN2(n13457), .QN(g33627) );
  NAND2X0 U13442 ( .IN1(n13458), .IN2(n13459), .QN(n13457) );
  NAND2X0 U13443 ( .IN1(n13460), .IN2(n13461), .QN(n13458) );
  NAND2X0 U13444 ( .IN1(n13462), .IN2(n10966), .QN(n13461) );
  NAND2X0 U13445 ( .IN1(n11278), .IN2(n13463), .QN(n13462) );
  NAND2X0 U13446 ( .IN1(n10629), .IN2(g6682), .QN(n13463) );
  NAND2X0 U13447 ( .IN1(n11282), .IN2(n13464), .QN(n13460) );
  NAND2X0 U13448 ( .IN1(n11067), .IN2(g6741), .QN(n13456) );
  NAND2X0 U13449 ( .IN1(n13465), .IN2(n13466), .QN(g33626) );
  NAND2X0 U13450 ( .IN1(n13467), .IN2(g6741), .QN(n13466) );
  NOR2X0 U13451 ( .IN1(n13468), .IN2(n13469), .QN(n13465) );
  NOR2X0 U13452 ( .IN1(n10523), .IN2(n10854), .QN(n13469) );
  NOR2X0 U13453 ( .IN1(n11047), .IN2(n13470), .QN(n13468) );
  NAND2X0 U13454 ( .IN1(n13471), .IN2(n5398), .QN(n13470) );
  NOR2X0 U13455 ( .IN1(n10629), .IN2(n13472), .QN(n13471) );
  INVX0 U13456 ( .INP(n13459), .ZN(n13472) );
  NAND2X0 U13457 ( .IN1(n13473), .IN2(n3023), .QN(n13459) );
  NOR2X0 U13458 ( .IN1(n10629), .IN2(n12437), .QN(n13473) );
  NAND2X0 U13459 ( .IN1(n13474), .IN2(n13475), .QN(g33625) );
  NAND2X0 U13460 ( .IN1(n13476), .IN2(n13477), .QN(n13475) );
  NAND2X0 U13461 ( .IN1(n13478), .IN2(n13479), .QN(n13476) );
  NAND2X0 U13462 ( .IN1(n13480), .IN2(n10966), .QN(n13479) );
  NAND2X0 U13463 ( .IN1(n13481), .IN2(n13482), .QN(n13480) );
  NAND2X0 U13464 ( .IN1(n13483), .IN2(g6336), .QN(n13482) );
  NAND2X0 U13465 ( .IN1(n13484), .IN2(n13485), .QN(n13478) );
  NAND2X0 U13466 ( .IN1(n11067), .IN2(g6395), .QN(n13474) );
  NAND2X0 U13467 ( .IN1(n13486), .IN2(n13487), .QN(g33624) );
  NAND2X0 U13468 ( .IN1(n13488), .IN2(g6395), .QN(n13487) );
  NOR2X0 U13469 ( .IN1(n13489), .IN2(n13490), .QN(n13486) );
  NOR2X0 U13470 ( .IN1(n10389), .IN2(n10853), .QN(n13490) );
  NOR2X0 U13471 ( .IN1(n11058), .IN2(n13491), .QN(n13489) );
  NAND2X0 U13472 ( .IN1(n13492), .IN2(n5396), .QN(n13491) );
  NOR2X0 U13473 ( .IN1(n13493), .IN2(n13483), .QN(n13492) );
  INVX0 U13474 ( .INP(n13477), .ZN(n13493) );
  NAND2X0 U13475 ( .IN1(n13494), .IN2(n3033), .QN(n13477) );
  NOR2X0 U13476 ( .IN1(n12444), .IN2(n13483), .QN(n13494) );
  NAND2X0 U13477 ( .IN1(n13495), .IN2(n13496), .QN(g33623) );
  NAND2X0 U13478 ( .IN1(n13497), .IN2(n13498), .QN(n13496) );
  NAND2X0 U13479 ( .IN1(n13499), .IN2(n13500), .QN(n13497) );
  NAND2X0 U13480 ( .IN1(n13501), .IN2(n10965), .QN(n13500) );
  NAND2X0 U13481 ( .IN1(n13502), .IN2(n13503), .QN(n13501) );
  NAND2X0 U13482 ( .IN1(n13504), .IN2(g5990), .QN(n13503) );
  NAND2X0 U13483 ( .IN1(n13505), .IN2(n13506), .QN(n13499) );
  NAND2X0 U13484 ( .IN1(test_so57), .IN2(n11081), .QN(n13495) );
  NAND2X0 U13485 ( .IN1(n13507), .IN2(n13508), .QN(g33622) );
  NAND2X0 U13486 ( .IN1(test_so50), .IN2(n11081), .QN(n13508) );
  NOR2X0 U13487 ( .IN1(n13509), .IN2(n13510), .QN(n13507) );
  NOR2X0 U13488 ( .IN1(n10639), .IN2(n13511), .QN(n13510) );
  NOR2X0 U13489 ( .IN1(test_so57), .IN2(n13512), .QN(n13509) );
  NAND2X0 U13490 ( .IN1(n13513), .IN2(n13498), .QN(n13512) );
  NAND2X0 U13491 ( .IN1(n13514), .IN2(n3033), .QN(n13498) );
  NOR2X0 U13492 ( .IN1(n13504), .IN2(n12438), .QN(n13514) );
  INVX0 U13493 ( .INP(n13515), .ZN(n13513) );
  NAND2X0 U13494 ( .IN1(n13516), .IN2(n13517), .QN(g33621) );
  NAND2X0 U13495 ( .IN1(n13518), .IN2(n13519), .QN(n13517) );
  NAND2X0 U13496 ( .IN1(n13520), .IN2(n13521), .QN(n13518) );
  NAND2X0 U13497 ( .IN1(n13522), .IN2(n10965), .QN(n13521) );
  NAND2X0 U13498 ( .IN1(n13523), .IN2(n13524), .QN(n13522) );
  NAND2X0 U13499 ( .IN1(n13525), .IN2(g5644), .QN(n13524) );
  NAND2X0 U13500 ( .IN1(n13526), .IN2(n13527), .QN(n13520) );
  NAND2X0 U13501 ( .IN1(n11067), .IN2(g5703), .QN(n13516) );
  NAND2X0 U13502 ( .IN1(n13528), .IN2(n13529), .QN(g33620) );
  NAND2X0 U13503 ( .IN1(n13530), .IN2(g5703), .QN(n13529) );
  NOR2X0 U13504 ( .IN1(n13531), .IN2(n13532), .QN(n13528) );
  NOR2X0 U13505 ( .IN1(n10394), .IN2(n10853), .QN(n13532) );
  NOR2X0 U13506 ( .IN1(n11058), .IN2(n13533), .QN(n13531) );
  NAND2X0 U13507 ( .IN1(n13534), .IN2(n5397), .QN(n13533) );
  NOR2X0 U13508 ( .IN1(n13535), .IN2(n13525), .QN(n13534) );
  INVX0 U13509 ( .INP(n13519), .ZN(n13535) );
  NAND2X0 U13510 ( .IN1(n13536), .IN2(n3023), .QN(n13519) );
  NOR2X0 U13511 ( .IN1(n13525), .IN2(n12444), .QN(n13536) );
  NAND2X0 U13512 ( .IN1(test_so81), .IN2(n12459), .QN(n12444) );
  NAND2X0 U13513 ( .IN1(n13537), .IN2(n13538), .QN(g33619) );
  NAND2X0 U13514 ( .IN1(n13539), .IN2(n13540), .QN(n13538) );
  NAND2X0 U13515 ( .IN1(n13541), .IN2(n13542), .QN(n13539) );
  NAND2X0 U13516 ( .IN1(n13543), .IN2(n10965), .QN(n13542) );
  NAND2X0 U13517 ( .IN1(n11267), .IN2(n13544), .QN(n13543) );
  NAND2X0 U13518 ( .IN1(n10624), .IN2(g5297), .QN(n13544) );
  NAND2X0 U13519 ( .IN1(n13545), .IN2(g33959), .QN(n13541) );
  NAND2X0 U13520 ( .IN1(n11067), .IN2(g5357), .QN(n13537) );
  NAND2X0 U13521 ( .IN1(n13546), .IN2(n13547), .QN(g33618) );
  NAND2X0 U13522 ( .IN1(n13548), .IN2(g5357), .QN(n13547) );
  NOR2X0 U13523 ( .IN1(n13549), .IN2(n13550), .QN(n13546) );
  NOR2X0 U13524 ( .IN1(n10525), .IN2(n10853), .QN(n13550) );
  NOR2X0 U13525 ( .IN1(n11058), .IN2(n13551), .QN(n13549) );
  NAND2X0 U13526 ( .IN1(n13552), .IN2(n5393), .QN(n13551) );
  NOR2X0 U13527 ( .IN1(n10624), .IN2(n13553), .QN(n13552) );
  INVX0 U13528 ( .INP(n13540), .ZN(n13553) );
  NAND2X0 U13529 ( .IN1(n13554), .IN2(n3023), .QN(n13540) );
  NOR2X0 U13530 ( .IN1(n10624), .IN2(n12438), .QN(n13554) );
  NAND2X0 U13531 ( .IN1(n12459), .IN2(n10643), .QN(n12438) );
  INVX0 U13532 ( .INP(n12058), .ZN(n12459) );
  NAND2X0 U13533 ( .IN1(n13555), .IN2(n5323), .QN(n12058) );
  NOR2X0 U13534 ( .IN1(n11944), .IN2(n13556), .QN(n13555) );
  INVX0 U13535 ( .INP(n13557), .ZN(n13556) );
  NAND2X0 U13536 ( .IN1(n13558), .IN2(n13559), .QN(g33617) );
  NAND2X0 U13537 ( .IN1(n13560), .IN2(g4552), .QN(n13559) );
  NOR2X0 U13538 ( .IN1(n12764), .IN2(n13561), .QN(n13558) );
  NAND2X0 U13539 ( .IN1(n13562), .IN2(n13563), .QN(g33616) );
  NOR2X0 U13540 ( .IN1(n12764), .IN2(n13564), .QN(n13563) );
  NOR2X0 U13541 ( .IN1(n13565), .IN2(n13566), .QN(n13562) );
  NOR2X0 U13542 ( .IN1(n10533), .IN2(n10852), .QN(n13566) );
  NOR2X0 U13543 ( .IN1(n10265), .IN2(n13567), .QN(n13565) );
  NAND2X0 U13544 ( .IN1(n3064), .IN2(n13568), .QN(g33615) );
  NAND2X0 U13545 ( .IN1(n13569), .IN2(g4108), .QN(n13568) );
  NAND2X0 U13546 ( .IN1(n13570), .IN2(n10965), .QN(n13569) );
  NAND2X0 U13547 ( .IN1(n11438), .IN2(n10403), .QN(n13570) );
  INVX0 U13548 ( .INP(n13571), .ZN(n11438) );
  NAND2X0 U13549 ( .IN1(n13572), .IN2(n13573), .QN(g33614) );
  NAND2X0 U13550 ( .IN1(n13574), .IN2(n13575), .QN(n13573) );
  NAND2X0 U13551 ( .IN1(n13576), .IN2(n13577), .QN(n13574) );
  NAND2X0 U13552 ( .IN1(n13578), .IN2(n10964), .QN(n13577) );
  NAND2X0 U13553 ( .IN1(n13579), .IN2(n13580), .QN(n13578) );
  NAND2X0 U13554 ( .IN1(n13581), .IN2(g3990), .QN(n13580) );
  NAND2X0 U13555 ( .IN1(n13582), .IN2(n13583), .QN(n13576) );
  NAND2X0 U13556 ( .IN1(n11067), .IN2(g4054), .QN(n13572) );
  NAND2X0 U13557 ( .IN1(n13584), .IN2(n13585), .QN(g33613) );
  NAND2X0 U13558 ( .IN1(n13586), .IN2(g4054), .QN(n13585) );
  NOR2X0 U13559 ( .IN1(n13587), .IN2(n13588), .QN(n13584) );
  NOR2X0 U13560 ( .IN1(n10396), .IN2(n10852), .QN(n13588) );
  NOR2X0 U13561 ( .IN1(n11058), .IN2(n13589), .QN(n13587) );
  NAND2X0 U13562 ( .IN1(n13590), .IN2(n5395), .QN(n13589) );
  NOR2X0 U13563 ( .IN1(n13591), .IN2(n13581), .QN(n13590) );
  INVX0 U13564 ( .INP(n13575), .ZN(n13591) );
  NAND2X0 U13565 ( .IN1(n13592), .IN2(n13583), .QN(n13575) );
  NOR2X0 U13566 ( .IN1(n12441), .IN2(n13593), .QN(n13592) );
  NAND2X0 U13567 ( .IN1(n13594), .IN2(n13595), .QN(g33612) );
  NAND2X0 U13568 ( .IN1(n13596), .IN2(n13597), .QN(n13595) );
  NAND2X0 U13569 ( .IN1(n13598), .IN2(n13599), .QN(n13596) );
  NAND2X0 U13570 ( .IN1(n13600), .IN2(n10964), .QN(n13599) );
  NAND2X0 U13571 ( .IN1(n13601), .IN2(n13602), .QN(n13600) );
  NAND2X0 U13572 ( .IN1(n13603), .IN2(g3639), .QN(n13602) );
  NAND2X0 U13573 ( .IN1(n13604), .IN2(n13605), .QN(n13598) );
  NAND2X0 U13574 ( .IN1(n11067), .IN2(g3703), .QN(n13594) );
  NAND2X0 U13575 ( .IN1(n13606), .IN2(n13607), .QN(g33611) );
  NAND2X0 U13576 ( .IN1(n13608), .IN2(g3703), .QN(n13607) );
  NOR2X0 U13577 ( .IN1(n13609), .IN2(n13610), .QN(n13606) );
  NOR2X0 U13578 ( .IN1(n10392), .IN2(n10852), .QN(n13610) );
  NOR2X0 U13579 ( .IN1(n11057), .IN2(n13611), .QN(n13609) );
  NAND2X0 U13580 ( .IN1(n13612), .IN2(n5399), .QN(n13611) );
  NOR2X0 U13581 ( .IN1(n13613), .IN2(n13603), .QN(n13612) );
  INVX0 U13582 ( .INP(n13597), .ZN(n13613) );
  NAND2X0 U13583 ( .IN1(n13614), .IN2(n13605), .QN(n13597) );
  NOR2X0 U13584 ( .IN1(n12437), .IN2(n13593), .QN(n13614) );
  INVX0 U13585 ( .INP(n3033), .ZN(n13593) );
  NAND2X0 U13586 ( .IN1(n12458), .IN2(n10643), .QN(n12437) );
  NAND2X0 U13587 ( .IN1(n13615), .IN2(n13616), .QN(g33610) );
  NAND2X0 U13588 ( .IN1(n11067), .IN2(g3352), .QN(n13616) );
  NAND2X0 U13589 ( .IN1(n13617), .IN2(n10964), .QN(n13615) );
  NOR2X0 U13590 ( .IN1(n13618), .IN2(n13619), .QN(n13617) );
  NOR2X0 U13591 ( .IN1(n13620), .IN2(n13621), .QN(n13619) );
  NAND2X0 U13592 ( .IN1(n13622), .IN2(n13623), .QN(n13621) );
  NAND2X0 U13593 ( .IN1(n13624), .IN2(n13625), .QN(n13623) );
  NAND2X0 U13594 ( .IN1(n13626), .IN2(g3288), .QN(n13622) );
  NAND2X0 U13595 ( .IN1(n13627), .IN2(n13628), .QN(g33609) );
  NAND2X0 U13596 ( .IN1(n13629), .IN2(g3352), .QN(n13628) );
  NOR2X0 U13597 ( .IN1(n13630), .IN2(n13631), .QN(n13627) );
  NOR2X0 U13598 ( .IN1(n10387), .IN2(n10852), .QN(n13631) );
  NOR2X0 U13599 ( .IN1(n11057), .IN2(n13632), .QN(n13630) );
  NAND2X0 U13600 ( .IN1(n13633), .IN2(n5604), .QN(n13632) );
  NOR2X0 U13601 ( .IN1(n13618), .IN2(n13626), .QN(n13633) );
  NOR2X0 U13602 ( .IN1(n13634), .IN2(n13626), .QN(n13618) );
  NAND2X0 U13603 ( .IN1(n13635), .IN2(n3023), .QN(n13634) );
  INVX0 U13604 ( .INP(n12441), .ZN(n13635) );
  NAND2X0 U13605 ( .IN1(n12458), .IN2(test_so81), .QN(n12441) );
  INVX0 U13606 ( .INP(n12062), .ZN(n12458) );
  NAND2X0 U13607 ( .IN1(n13636), .IN2(n13557), .QN(n12062) );
  XNOR2X1 U13608 ( .IN1(n11433), .IN2(n5540), .Q(n13557) );
  NOR2X0 U13609 ( .IN1(n5323), .IN2(n11944), .QN(n13636) );
  XOR2X1 U13610 ( .IN1(n13381), .IN2(n5506), .Q(n11944) );
  NAND2X0 U13611 ( .IN1(n13637), .IN2(n13638), .QN(g33608) );
  NOR2X0 U13612 ( .IN1(n13639), .IN2(n13640), .QN(n13638) );
  NOR2X0 U13613 ( .IN1(n10904), .IN2(n5300), .QN(n13640) );
  NOR2X0 U13614 ( .IN1(n11057), .IN2(n13641), .QN(n13639) );
  NAND2X0 U13615 ( .IN1(n12781), .IN2(g2759), .QN(n13641) );
  NOR2X0 U13616 ( .IN1(n2787), .IN2(n13642), .QN(n13637) );
  NOR2X0 U13617 ( .IN1(g2759), .IN2(n12781), .QN(n13642) );
  NAND2X0 U13618 ( .IN1(n2790), .IN2(test_so30), .QN(n12781) );
  NAND2X0 U13619 ( .IN1(n13643), .IN2(n13644), .QN(g33607) );
  NAND2X0 U13620 ( .IN1(n11067), .IN2(g2555), .QN(n13644) );
  NOR2X0 U13621 ( .IN1(n13645), .IN2(n13646), .QN(n13643) );
  NOR2X0 U13622 ( .IN1(n5311), .IN2(n13647), .QN(n13646) );
  NOR2X0 U13623 ( .IN1(n13648), .IN2(n13649), .QN(n13647) );
  NOR2X0 U13624 ( .IN1(n3105), .IN2(n11023), .QN(n13648) );
  NOR2X0 U13625 ( .IN1(n13650), .IN2(n13651), .QN(n13645) );
  NAND2X0 U13626 ( .IN1(n13652), .IN2(n13653), .QN(n13651) );
  NAND2X0 U13627 ( .IN1(n13654), .IN2(n13655), .QN(n13653) );
  NAND2X0 U13628 ( .IN1(n13656), .IN2(n12486), .QN(n13655) );
  NOR2X0 U13629 ( .IN1(n5521), .IN2(n2726), .QN(n12486) );
  NAND2X0 U13630 ( .IN1(n5519), .IN2(n12473), .QN(n2726) );
  NOR2X0 U13631 ( .IN1(n13657), .IN2(g2599), .QN(n13656) );
  NAND2X0 U13632 ( .IN1(n3111), .IN2(n10964), .QN(n13654) );
  NAND2X0 U13633 ( .IN1(n13658), .IN2(n5524), .QN(n13652) );
  NOR2X0 U13634 ( .IN1(n5521), .IN2(n10273), .QN(n13658) );
  NAND2X0 U13635 ( .IN1(n13659), .IN2(n13660), .QN(g33606) );
  NAND2X0 U13636 ( .IN1(n13661), .IN2(g2675), .QN(n13660) );
  NOR2X0 U13637 ( .IN1(n13662), .IN2(n13663), .QN(n13659) );
  NOR2X0 U13638 ( .IN1(n5278), .IN2(n10851), .QN(n13663) );
  NOR2X0 U13639 ( .IN1(n11058), .IN2(n13664), .QN(n13662) );
  NAND2X0 U13640 ( .IN1(n5457), .IN2(n12808), .QN(n13664) );
  INVX0 U13641 ( .INP(n12788), .ZN(n12808) );
  NAND2X0 U13642 ( .IN1(n13665), .IN2(n13666), .QN(g33605) );
  NAND2X0 U13643 ( .IN1(n13661), .IN2(g2671), .QN(n13666) );
  NOR2X0 U13644 ( .IN1(n13667), .IN2(n13668), .QN(n13665) );
  NOR2X0 U13645 ( .IN1(test_so48), .IN2(n13669), .QN(n13668) );
  NAND2X0 U13646 ( .IN1(n13670), .IN2(n5418), .QN(n13669) );
  NOR2X0 U13647 ( .IN1(n11057), .IN2(n12788), .QN(n13670) );
  NOR2X0 U13648 ( .IN1(n13671), .IN2(n10676), .QN(n13667) );
  NOR2X0 U13649 ( .IN1(n11057), .IN2(n13672), .QN(n13671) );
  NOR2X0 U13650 ( .IN1(n5418), .IN2(n12788), .QN(n13672) );
  NAND2X0 U13651 ( .IN1(n13673), .IN2(n13674), .QN(g33604) );
  NAND2X0 U13652 ( .IN1(test_so48), .IN2(n13661), .QN(n13674) );
  NAND2X0 U13653 ( .IN1(n12786), .IN2(g2661), .QN(n13673) );
  NAND2X0 U13654 ( .IN1(n13675), .IN2(n13676), .QN(g33603) );
  NAND2X0 U13655 ( .IN1(n13661), .IN2(g2648), .QN(n13676) );
  INVX0 U13656 ( .INP(n12786), .ZN(n13661) );
  NAND2X0 U13657 ( .IN1(n12786), .IN2(g2643), .QN(n13675) );
  NAND2X0 U13658 ( .IN1(n12788), .IN2(n10963), .QN(n12786) );
  NAND2X0 U13659 ( .IN1(n13677), .IN2(n5521), .QN(n12788) );
  NOR2X0 U13660 ( .IN1(n12809), .IN2(g2555), .QN(n13677) );
  NAND2X0 U13661 ( .IN1(n13678), .IN2(n13679), .QN(g33602) );
  INVX0 U13662 ( .INP(n13680), .ZN(n13679) );
  NOR2X0 U13663 ( .IN1(n12826), .IN2(n3111), .QN(n13680) );
  NAND2X0 U13664 ( .IN1(g2599), .IN2(n12802), .QN(n12826) );
  NOR2X0 U13665 ( .IN1(n13681), .IN2(n13682), .QN(n13678) );
  NOR2X0 U13666 ( .IN1(n11057), .IN2(n13683), .QN(n13682) );
  NAND2X0 U13667 ( .IN1(n12809), .IN2(g2629), .QN(n13683) );
  NOR2X0 U13668 ( .IN1(n5524), .IN2(n10851), .QN(n13681) );
  NAND2X0 U13669 ( .IN1(n13684), .IN2(n13685), .QN(g33601) );
  NAND2X0 U13670 ( .IN1(n13686), .IN2(n12796), .QN(n13685) );
  NOR2X0 U13671 ( .IN1(n3111), .IN2(n12809), .QN(n13686) );
  NOR2X0 U13672 ( .IN1(n13687), .IN2(n13688), .QN(n13684) );
  NOR2X0 U13673 ( .IN1(n5311), .IN2(n10851), .QN(n13688) );
  NOR2X0 U13674 ( .IN1(n11057), .IN2(n13689), .QN(n13687) );
  NAND2X0 U13675 ( .IN1(n12809), .IN2(g2599), .QN(n13689) );
  NAND2X0 U13676 ( .IN1(n13690), .IN2(n13691), .QN(g33600) );
  NAND2X0 U13677 ( .IN1(n13692), .IN2(n13693), .QN(n13691) );
  NOR2X0 U13678 ( .IN1(n3111), .IN2(n11023), .QN(n13693) );
  NOR2X0 U13679 ( .IN1(n13694), .IN2(g2629), .QN(n13692) );
  NOR2X0 U13680 ( .IN1(n12818), .IN2(g2555), .QN(n13694) );
  NOR2X0 U13681 ( .IN1(g2599), .IN2(n12809), .QN(n12818) );
  NAND2X0 U13682 ( .IN1(n12796), .IN2(n12809), .QN(n13690) );
  INVX0 U13683 ( .INP(n12802), .ZN(n12809) );
  NAND2X0 U13684 ( .IN1(n12851), .IN2(n13650), .QN(n12802) );
  INVX0 U13685 ( .INP(n735), .ZN(n13650) );
  NOR2X0 U13686 ( .IN1(n10546), .IN2(n13695), .QN(n735) );
  NOR2X0 U13687 ( .IN1(n13696), .IN2(g1514), .QN(n13695) );
  NAND2X0 U13688 ( .IN1(n10662), .IN2(n13697), .QN(n13696) );
  INVX0 U13689 ( .INP(n12806), .ZN(n12851) );
  NAND2X0 U13690 ( .IN1(n13698), .IN2(n13699), .QN(n12806) );
  NAND2X0 U13691 ( .IN1(n2549), .IN2(g1300), .QN(n13699) );
  NOR2X0 U13692 ( .IN1(n13066), .IN2(n13700), .QN(n13698) );
  NOR2X0 U13693 ( .IN1(n5308), .IN2(n13701), .QN(n13700) );
  NOR2X0 U13694 ( .IN1(n11057), .IN2(n5351), .QN(n12796) );
  NAND2X0 U13695 ( .IN1(n13702), .IN2(n13703), .QN(g33599) );
  NOR2X0 U13696 ( .IN1(n13704), .IN2(n13705), .QN(n13703) );
  NOR2X0 U13697 ( .IN1(n11056), .IN2(n13706), .QN(n13705) );
  NAND2X0 U13698 ( .IN1(n13707), .IN2(n3131), .QN(n13706) );
  NOR2X0 U13699 ( .IN1(n13708), .IN2(n11435), .QN(n13707) );
  NOR2X0 U13700 ( .IN1(n10273), .IN2(n12891), .QN(n13708) );
  NOR2X0 U13701 ( .IN1(n10908), .IN2(n10648), .QN(n13704) );
  NOR2X0 U13702 ( .IN1(n13709), .IN2(n13710), .QN(n13702) );
  NOR2X0 U13703 ( .IN1(n5619), .IN2(n13711), .QN(n13710) );
  NOR2X0 U13704 ( .IN1(n13712), .IN2(n13649), .QN(n13711) );
  NOR2X0 U13705 ( .IN1(n3125), .IN2(n11023), .QN(n13712) );
  INVX0 U13706 ( .INP(n571), .ZN(n13709) );
  NAND2X0 U13707 ( .IN1(n13713), .IN2(n13714), .QN(n571) );
  NOR2X0 U13708 ( .IN1(n13657), .IN2(n12492), .QN(n13714) );
  NAND2X0 U13709 ( .IN1(n13715), .IN2(n13716), .QN(n12492) );
  INVX0 U13710 ( .INP(n2727), .ZN(n13716) );
  NAND2X0 U13711 ( .IN1(n12473), .IN2(g504), .QN(n2727) );
  NOR2X0 U13712 ( .IN1(n13717), .IN2(n5287), .QN(n12473) );
  INVX0 U13713 ( .INP(n12891), .ZN(n13715) );
  NAND2X0 U13714 ( .IN1(n5523), .IN2(g2495), .QN(n12891) );
  NOR2X0 U13715 ( .IN1(n11435), .IN2(g112), .QN(n13713) );
  NAND2X0 U13716 ( .IN1(n13718), .IN2(n13719), .QN(g33598) );
  NAND2X0 U13717 ( .IN1(n11236), .IN2(g2541), .QN(n13719) );
  NOR2X0 U13718 ( .IN1(n13720), .IN2(n13721), .QN(n13718) );
  NOR2X0 U13719 ( .IN1(n5411), .IN2(n10850), .QN(n13721) );
  NOR2X0 U13720 ( .IN1(n11056), .IN2(n13722), .QN(n13720) );
  NAND2X0 U13721 ( .IN1(n5461), .IN2(n12881), .QN(n13722) );
  INVX0 U13722 ( .INP(n12861), .ZN(n12881) );
  NAND2X0 U13723 ( .IN1(n13723), .IN2(n13724), .QN(g33597) );
  NAND2X0 U13724 ( .IN1(n11236), .IN2(g2537), .QN(n13724) );
  NOR2X0 U13725 ( .IN1(n13725), .IN2(n13726), .QN(n13723) );
  NOR2X0 U13726 ( .IN1(g2533), .IN2(n13727), .QN(n13726) );
  NAND2X0 U13727 ( .IN1(n13728), .IN2(n5420), .QN(n13727) );
  NOR2X0 U13728 ( .IN1(n11057), .IN2(n12861), .QN(n13728) );
  NOR2X0 U13729 ( .IN1(n5761), .IN2(n13729), .QN(n13725) );
  NOR2X0 U13730 ( .IN1(n11056), .IN2(n13730), .QN(n13729) );
  NOR2X0 U13731 ( .IN1(n5420), .IN2(n12861), .QN(n13730) );
  NAND2X0 U13732 ( .IN1(n13731), .IN2(n13732), .QN(g33595) );
  NAND2X0 U13733 ( .IN1(n11236), .IN2(g2514), .QN(n13732) );
  INVX0 U13734 ( .INP(n11237), .ZN(n11236) );
  NAND2X0 U13735 ( .IN1(n11237), .IN2(g2509), .QN(n13731) );
  NAND2X0 U13736 ( .IN1(n12861), .IN2(n10963), .QN(n11237) );
  NAND2X0 U13737 ( .IN1(n13733), .IN2(n5522), .QN(n12861) );
  NOR2X0 U13738 ( .IN1(test_so79), .IN2(n12882), .QN(n13733) );
  NAND2X0 U13739 ( .IN1(n13734), .IN2(n13735), .QN(g33594) );
  NAND2X0 U13740 ( .IN1(n11067), .IN2(g2465), .QN(n13735) );
  NOR2X0 U13741 ( .IN1(n13736), .IN2(n13737), .QN(n13734) );
  NOR2X0 U13742 ( .IN1(n3131), .IN2(n12899), .QN(n13737) );
  NAND2X0 U13743 ( .IN1(g2465), .IN2(n12875), .QN(n12899) );
  NOR2X0 U13744 ( .IN1(n5522), .IN2(n13738), .QN(n13736) );
  INVX0 U13745 ( .INP(n13739), .ZN(n13738) );
  NAND2X0 U13746 ( .IN1(n13740), .IN2(n13741), .QN(g33593) );
  NAND2X0 U13747 ( .IN1(n13739), .IN2(g2465), .QN(n13741) );
  NOR2X0 U13748 ( .IN1(n13742), .IN2(n13743), .QN(n13740) );
  INVX0 U13749 ( .INP(n13744), .ZN(n13743) );
  NAND2X0 U13750 ( .IN1(n10925), .IN2(n13745), .QN(n13744) );
  NOR2X0 U13751 ( .IN1(n12907), .IN2(n3131), .QN(n13745) );
  NAND2X0 U13752 ( .IN1(test_so79), .IN2(n12875), .QN(n12907) );
  NOR2X0 U13753 ( .IN1(n5619), .IN2(n10850), .QN(n13742) );
  NAND2X0 U13754 ( .IN1(n13746), .IN2(n13747), .QN(g33592) );
  NAND2X0 U13755 ( .IN1(n13748), .IN2(n13749), .QN(n13747) );
  NOR2X0 U13756 ( .IN1(n3131), .IN2(n11023), .QN(n13749) );
  NOR2X0 U13757 ( .IN1(n13750), .IN2(g2495), .QN(n13748) );
  NOR2X0 U13758 ( .IN1(n13751), .IN2(test_so79), .QN(n13750) );
  NOR2X0 U13759 ( .IN1(n12882), .IN2(g2465), .QN(n13751) );
  INVX0 U13760 ( .INP(n12875), .ZN(n12882) );
  NAND2X0 U13761 ( .IN1(n13739), .IN2(test_so79), .QN(n13746) );
  NOR2X0 U13762 ( .IN1(n12875), .IN2(n11023), .QN(n13739) );
  NAND2X0 U13763 ( .IN1(n12922), .IN2(n11435), .QN(n12875) );
  NAND2X0 U13764 ( .IN1(n13752), .IN2(g17423), .QN(n11435) );
  NAND2X0 U13765 ( .IN1(n13697), .IN2(n13753), .QN(n13752) );
  INVX0 U13766 ( .INP(n13754), .ZN(n13697) );
  INVX0 U13767 ( .INP(n12879), .ZN(n12922) );
  NAND2X0 U13768 ( .IN1(n13755), .IN2(n13756), .QN(n12879) );
  NAND2X0 U13769 ( .IN1(n2549), .IN2(g1472), .QN(n13756) );
  NOR2X0 U13770 ( .IN1(n13066), .IN2(n13757), .QN(n13755) );
  NOR2X0 U13771 ( .IN1(g2704), .IN2(n13758), .QN(n13757) );
  NAND2X0 U13772 ( .IN1(g2697), .IN2(g2689), .QN(n13758) );
  NAND2X0 U13773 ( .IN1(n13759), .IN2(n13760), .QN(g33591) );
  NAND2X0 U13774 ( .IN1(n11067), .IN2(g2287), .QN(n13760) );
  NOR2X0 U13775 ( .IN1(n13761), .IN2(n13762), .QN(n13759) );
  NOR2X0 U13776 ( .IN1(n5310), .IN2(n13763), .QN(n13762) );
  NOR2X0 U13777 ( .IN1(n13764), .IN2(n13649), .QN(n13763) );
  NOR2X0 U13778 ( .IN1(n3145), .IN2(n11023), .QN(n13764) );
  NOR2X0 U13779 ( .IN1(n13765), .IN2(n13766), .QN(n13761) );
  NAND2X0 U13780 ( .IN1(n13767), .IN2(n13768), .QN(n13766) );
  NAND2X0 U13781 ( .IN1(n13769), .IN2(n13770), .QN(n13768) );
  NAND2X0 U13782 ( .IN1(n13771), .IN2(n12481), .QN(n13770) );
  NOR2X0 U13783 ( .IN1(n5537), .IN2(n3146), .QN(n12481) );
  NOR2X0 U13784 ( .IN1(n13657), .IN2(g2331), .QN(n13771) );
  NAND2X0 U13785 ( .IN1(n13772), .IN2(n10962), .QN(n13769) );
  NAND2X0 U13786 ( .IN1(n13773), .IN2(n5513), .QN(n13767) );
  NOR2X0 U13787 ( .IN1(n5537), .IN2(n10273), .QN(n13773) );
  INVX0 U13788 ( .INP(n3141), .ZN(n13765) );
  NAND2X0 U13789 ( .IN1(n13774), .IN2(n13775), .QN(g33590) );
  NAND2X0 U13790 ( .IN1(n11408), .IN2(g2407), .QN(n13775) );
  NOR2X0 U13791 ( .IN1(n13776), .IN2(n13777), .QN(n13774) );
  NOR2X0 U13792 ( .IN1(n10903), .IN2(n10671), .QN(n13777) );
  NOR2X0 U13793 ( .IN1(n11056), .IN2(n13778), .QN(n13776) );
  NAND2X0 U13794 ( .IN1(n5459), .IN2(n12952), .QN(n13778) );
  INVX0 U13795 ( .INP(n12932), .ZN(n12952) );
  NAND2X0 U13796 ( .IN1(n13779), .IN2(n13780), .QN(g33589) );
  NAND2X0 U13797 ( .IN1(test_so31), .IN2(n11408), .QN(n13780) );
  NOR2X0 U13798 ( .IN1(n13781), .IN2(n13782), .QN(n13779) );
  NOR2X0 U13799 ( .IN1(g2399), .IN2(n13783), .QN(n13782) );
  NAND2X0 U13800 ( .IN1(n13784), .IN2(n5421), .QN(n13783) );
  NOR2X0 U13801 ( .IN1(n11056), .IN2(n12932), .QN(n13784) );
  NOR2X0 U13802 ( .IN1(n5762), .IN2(n13785), .QN(n13781) );
  NOR2X0 U13803 ( .IN1(n11056), .IN2(n13786), .QN(n13785) );
  NOR2X0 U13804 ( .IN1(n5421), .IN2(n12932), .QN(n13786) );
  NAND2X0 U13805 ( .IN1(n13787), .IN2(n13788), .QN(g33587) );
  NAND2X0 U13806 ( .IN1(n11408), .IN2(g2380), .QN(n13788) );
  INVX0 U13807 ( .INP(n11409), .ZN(n11408) );
  NAND2X0 U13808 ( .IN1(n11409), .IN2(g2375), .QN(n13787) );
  NAND2X0 U13809 ( .IN1(n12932), .IN2(n10962), .QN(n11409) );
  NAND2X0 U13810 ( .IN1(n13789), .IN2(n5537), .QN(n12932) );
  NOR2X0 U13811 ( .IN1(n12953), .IN2(g2287), .QN(n13789) );
  NAND2X0 U13812 ( .IN1(n13790), .IN2(n13791), .QN(g33586) );
  INVX0 U13813 ( .INP(n13792), .ZN(n13791) );
  NOR2X0 U13814 ( .IN1(n12970), .IN2(n13772), .QN(n13792) );
  NAND2X0 U13815 ( .IN1(g2331), .IN2(n12946), .QN(n12970) );
  INVX0 U13816 ( .INP(n12953), .ZN(n12946) );
  NOR2X0 U13817 ( .IN1(n13793), .IN2(n13794), .QN(n13790) );
  NOR2X0 U13818 ( .IN1(n11056), .IN2(n13795), .QN(n13794) );
  NAND2X0 U13819 ( .IN1(n12953), .IN2(g2361), .QN(n13795) );
  NOR2X0 U13820 ( .IN1(n5513), .IN2(n10850), .QN(n13793) );
  NAND2X0 U13821 ( .IN1(n13796), .IN2(n13797), .QN(g33585) );
  NAND2X0 U13822 ( .IN1(n13798), .IN2(n12940), .QN(n13797) );
  NOR2X0 U13823 ( .IN1(n12953), .IN2(n13772), .QN(n13798) );
  NOR2X0 U13824 ( .IN1(n13799), .IN2(n13800), .QN(n13796) );
  NOR2X0 U13825 ( .IN1(n5310), .IN2(n10850), .QN(n13800) );
  NOR2X0 U13826 ( .IN1(n11056), .IN2(n13801), .QN(n13799) );
  NAND2X0 U13827 ( .IN1(n12953), .IN2(g2331), .QN(n13801) );
  NAND2X0 U13828 ( .IN1(n13802), .IN2(n13803), .QN(g33584) );
  NAND2X0 U13829 ( .IN1(n13804), .IN2(n13805), .QN(n13803) );
  NOR2X0 U13830 ( .IN1(n11056), .IN2(n13772), .QN(n13805) );
  NOR2X0 U13831 ( .IN1(n13806), .IN2(n3146), .QN(n13772) );
  NAND2X0 U13832 ( .IN1(n13807), .IN2(n3116), .QN(n3146) );
  NOR2X0 U13833 ( .IN1(n13808), .IN2(g2361), .QN(n13804) );
  NOR2X0 U13834 ( .IN1(n13809), .IN2(g2287), .QN(n13808) );
  NOR2X0 U13835 ( .IN1(n12953), .IN2(g2331), .QN(n13809) );
  NAND2X0 U13836 ( .IN1(n12940), .IN2(n12953), .QN(n13802) );
  NOR2X0 U13837 ( .IN1(n12950), .IN2(n3141), .QN(n12953) );
  NOR2X0 U13838 ( .IN1(n13810), .IN2(n10235), .QN(n3141) );
  NOR2X0 U13839 ( .IN1(n13811), .IN2(n13754), .QN(n13810) );
  NAND2X0 U13840 ( .IN1(n13812), .IN2(n13813), .QN(n12950) );
  NAND2X0 U13841 ( .IN1(n2549), .IN2(g1448), .QN(n13813) );
  NOR2X0 U13842 ( .IN1(n13066), .IN2(n13814), .QN(n13812) );
  NOR2X0 U13843 ( .IN1(g2697), .IN2(n13701), .QN(n13814) );
  NAND2X0 U13844 ( .IN1(g2689), .IN2(g2704), .QN(n13701) );
  NOR2X0 U13845 ( .IN1(n11056), .IN2(n5353), .QN(n12940) );
  NAND2X0 U13846 ( .IN1(n13815), .IN2(n13816), .QN(g33583) );
  NAND2X0 U13847 ( .IN1(n11066), .IN2(g2153), .QN(n13816) );
  NOR2X0 U13848 ( .IN1(n13817), .IN2(n13818), .QN(n13815) );
  NOR2X0 U13849 ( .IN1(n5620), .IN2(n13819), .QN(n13818) );
  NOR2X0 U13850 ( .IN1(n13820), .IN2(n13649), .QN(n13819) );
  NOR2X0 U13851 ( .IN1(n3164), .IN2(n11022), .QN(n13820) );
  NOR2X0 U13852 ( .IN1(n13821), .IN2(n13822), .QN(n13817) );
  NAND2X0 U13853 ( .IN1(n13823), .IN2(n13824), .QN(n13822) );
  NAND2X0 U13854 ( .IN1(n13825), .IN2(n13826), .QN(n13824) );
  NAND2X0 U13855 ( .IN1(n13827), .IN2(n12482), .QN(n13826) );
  NOR2X0 U13856 ( .IN1(n5538), .IN2(n3165), .QN(n12482) );
  NOR2X0 U13857 ( .IN1(n13657), .IN2(g2197), .QN(n13827) );
  NAND2X0 U13858 ( .IN1(n13828), .IN2(n10962), .QN(n13825) );
  NAND2X0 U13859 ( .IN1(n13829), .IN2(n5514), .QN(n13823) );
  NOR2X0 U13860 ( .IN1(n5538), .IN2(n10273), .QN(n13829) );
  INVX0 U13861 ( .INP(n751), .ZN(n13821) );
  NAND2X0 U13862 ( .IN1(n13830), .IN2(n13831), .QN(g33582) );
  NAND2X0 U13863 ( .IN1(n13832), .IN2(g2273), .QN(n13831) );
  NOR2X0 U13864 ( .IN1(n13833), .IN2(n13834), .QN(n13830) );
  NOR2X0 U13865 ( .IN1(n5410), .IN2(n10850), .QN(n13834) );
  NOR2X0 U13866 ( .IN1(n11056), .IN2(n13835), .QN(n13833) );
  NAND2X0 U13867 ( .IN1(n5458), .IN2(n13024), .QN(n13835) );
  INVX0 U13868 ( .INP(n13004), .ZN(n13024) );
  NAND2X0 U13869 ( .IN1(n13836), .IN2(n13837), .QN(g33581) );
  NAND2X0 U13870 ( .IN1(n13832), .IN2(g2269), .QN(n13837) );
  NOR2X0 U13871 ( .IN1(n13838), .IN2(n13839), .QN(n13836) );
  NOR2X0 U13872 ( .IN1(test_so62), .IN2(n13840), .QN(n13839) );
  NAND2X0 U13873 ( .IN1(n13841), .IN2(n5419), .QN(n13840) );
  NOR2X0 U13874 ( .IN1(n11056), .IN2(n13004), .QN(n13841) );
  NOR2X0 U13875 ( .IN1(n13842), .IN2(n10677), .QN(n13838) );
  NOR2X0 U13876 ( .IN1(n11055), .IN2(n13843), .QN(n13842) );
  NOR2X0 U13877 ( .IN1(n5419), .IN2(n13004), .QN(n13843) );
  NAND2X0 U13878 ( .IN1(n13844), .IN2(n13845), .QN(g33580) );
  NAND2X0 U13879 ( .IN1(test_so62), .IN2(n13832), .QN(n13845) );
  NAND2X0 U13880 ( .IN1(n13002), .IN2(g2259), .QN(n13844) );
  NAND2X0 U13881 ( .IN1(n13846), .IN2(n13847), .QN(g33579) );
  NAND2X0 U13882 ( .IN1(n13832), .IN2(g2246), .QN(n13847) );
  INVX0 U13883 ( .INP(n13002), .ZN(n13832) );
  NAND2X0 U13884 ( .IN1(n13002), .IN2(g2241), .QN(n13846) );
  NAND2X0 U13885 ( .IN1(n13004), .IN2(n10961), .QN(n13002) );
  NAND2X0 U13886 ( .IN1(n13848), .IN2(n5538), .QN(n13004) );
  NOR2X0 U13887 ( .IN1(n13025), .IN2(g2153), .QN(n13848) );
  NAND2X0 U13888 ( .IN1(n13849), .IN2(n13850), .QN(g33578) );
  INVX0 U13889 ( .INP(n13851), .ZN(n13850) );
  NOR2X0 U13890 ( .IN1(n13042), .IN2(n13828), .QN(n13851) );
  NAND2X0 U13891 ( .IN1(g2197), .IN2(n13018), .QN(n13042) );
  INVX0 U13892 ( .INP(n13025), .ZN(n13018) );
  NOR2X0 U13893 ( .IN1(n13852), .IN2(n13853), .QN(n13849) );
  NOR2X0 U13894 ( .IN1(n11055), .IN2(n13854), .QN(n13853) );
  NAND2X0 U13895 ( .IN1(n13025), .IN2(g2227), .QN(n13854) );
  NOR2X0 U13896 ( .IN1(n5514), .IN2(n10849), .QN(n13852) );
  NAND2X0 U13897 ( .IN1(n13855), .IN2(n13856), .QN(g33577) );
  NAND2X0 U13898 ( .IN1(n13857), .IN2(n13012), .QN(n13856) );
  NOR2X0 U13899 ( .IN1(n13025), .IN2(n13828), .QN(n13857) );
  NOR2X0 U13900 ( .IN1(n13858), .IN2(n13859), .QN(n13855) );
  NOR2X0 U13901 ( .IN1(n5620), .IN2(n10849), .QN(n13859) );
  NOR2X0 U13902 ( .IN1(n11055), .IN2(n13860), .QN(n13858) );
  NAND2X0 U13903 ( .IN1(n13025), .IN2(g2197), .QN(n13860) );
  NAND2X0 U13904 ( .IN1(n13861), .IN2(n13862), .QN(g33576) );
  NAND2X0 U13905 ( .IN1(n13863), .IN2(n13864), .QN(n13862) );
  NOR2X0 U13906 ( .IN1(n11055), .IN2(n13828), .QN(n13864) );
  NOR2X0 U13907 ( .IN1(n13806), .IN2(n3165), .QN(n13828) );
  NAND2X0 U13908 ( .IN1(n13865), .IN2(n5519), .QN(n3165) );
  NOR2X0 U13909 ( .IN1(g518), .IN2(n13717), .QN(n13865) );
  INVX0 U13910 ( .INP(n3116), .ZN(n13717) );
  NOR2X0 U13911 ( .IN1(n13866), .IN2(g2227), .QN(n13863) );
  NOR2X0 U13912 ( .IN1(n13867), .IN2(g2153), .QN(n13866) );
  NOR2X0 U13913 ( .IN1(n13025), .IN2(g2197), .QN(n13867) );
  NAND2X0 U13914 ( .IN1(n13012), .IN2(n13025), .QN(n13861) );
  NOR2X0 U13915 ( .IN1(n13022), .IN2(n751), .QN(n13025) );
  NOR2X0 U13916 ( .IN1(n10236), .IN2(n13868), .QN(n751) );
  NOR2X0 U13917 ( .IN1(n13869), .IN2(n13754), .QN(n13868) );
  NAND2X0 U13918 ( .IN1(n13870), .IN2(n13871), .QN(n13754) );
  NOR2X0 U13919 ( .IN1(g1559), .IN2(n13872), .QN(n13871) );
  NAND2X0 U13920 ( .IN1(n10545), .IN2(g1404), .QN(n13872) );
  NOR2X0 U13921 ( .IN1(n10650), .IN2(n13873), .QN(n13870) );
  NAND2X0 U13922 ( .IN1(n5768), .IN2(n5546), .QN(n13873) );
  NAND2X0 U13923 ( .IN1(n10662), .IN2(g1514), .QN(n13869) );
  NAND2X0 U13924 ( .IN1(n13874), .IN2(n13875), .QN(n13022) );
  NAND2X0 U13925 ( .IN1(n2549), .IN2(g1478), .QN(n13875) );
  NOR2X0 U13926 ( .IN1(n13066), .IN2(n13876), .QN(n13874) );
  NOR2X0 U13927 ( .IN1(g2697), .IN2(n13877), .QN(n13876) );
  NAND2X0 U13928 ( .IN1(n5377), .IN2(g2689), .QN(n13877) );
  NOR2X0 U13929 ( .IN1(n13878), .IN2(g134), .QN(n13066) );
  NOR2X0 U13930 ( .IN1(n11986), .IN2(n11992), .QN(n13878) );
  NOR2X0 U13931 ( .IN1(n11055), .IN2(n5356), .QN(n13012) );
  NAND2X0 U13932 ( .IN1(n13879), .IN2(n13880), .QN(g33575) );
  NOR2X0 U13933 ( .IN1(n13881), .IN2(n13882), .QN(n13880) );
  NOR2X0 U13934 ( .IN1(n11055), .IN2(n13883), .QN(n13882) );
  NAND2X0 U13935 ( .IN1(n13884), .IN2(n13885), .QN(n13883) );
  INVX0 U13936 ( .INP(n13886), .ZN(n13884) );
  NAND2X0 U13937 ( .IN1(n13887), .IN2(n13888), .QN(n13886) );
  NAND2X0 U13938 ( .IN1(g112), .IN2(n12491), .QN(n13887) );
  NOR2X0 U13939 ( .IN1(n5355), .IN2(n10849), .QN(n13881) );
  NOR2X0 U13940 ( .IN1(n11439), .IN2(n13889), .QN(n13879) );
  NOR2X0 U13941 ( .IN1(n5831), .IN2(n13890), .QN(n13889) );
  NOR2X0 U13942 ( .IN1(n13891), .IN2(n13649), .QN(n13890) );
  NOR2X0 U13943 ( .IN1(n11055), .IN2(n13892), .QN(n13891) );
  NOR2X0 U13944 ( .IN1(n13893), .IN2(n13894), .QN(n11439) );
  NAND2X0 U13945 ( .IN1(n12331), .IN2(n10273), .QN(n13894) );
  INVX0 U13946 ( .INP(n13657), .ZN(n12331) );
  NAND2X0 U13947 ( .IN1(n13892), .IN2(n12491), .QN(n13893) );
  NOR2X0 U13948 ( .IN1(g2040), .IN2(n5535), .QN(n12491) );
  INVX0 U13949 ( .INP(n13895), .ZN(n13892) );
  NAND2X0 U13950 ( .IN1(n13888), .IN2(n12472), .QN(n13895) );
  NAND2X0 U13951 ( .IN1(n13896), .IN2(n13897), .QN(g33574) );
  NAND2X0 U13952 ( .IN1(n11442), .IN2(g2116), .QN(n13897) );
  NOR2X0 U13953 ( .IN1(n13898), .IN2(n13899), .QN(n13896) );
  NOR2X0 U13954 ( .IN1(n5848), .IN2(n10849), .QN(n13899) );
  NOR2X0 U13955 ( .IN1(n11055), .IN2(n13900), .QN(n13898) );
  NAND2X0 U13956 ( .IN1(n5463), .IN2(n13097), .QN(n13900) );
  INVX0 U13957 ( .INP(n13077), .ZN(n13097) );
  NAND2X0 U13958 ( .IN1(n13901), .IN2(n13902), .QN(g33573) );
  NAND2X0 U13959 ( .IN1(n11442), .IN2(g2112), .QN(n13902) );
  NOR2X0 U13960 ( .IN1(n13903), .IN2(n13904), .QN(n13901) );
  NOR2X0 U13961 ( .IN1(g2108), .IN2(n13905), .QN(n13904) );
  NAND2X0 U13962 ( .IN1(n13906), .IN2(n5666), .QN(n13905) );
  NOR2X0 U13963 ( .IN1(n11055), .IN2(n13077), .QN(n13906) );
  NOR2X0 U13964 ( .IN1(n5452), .IN2(n13907), .QN(n13903) );
  NOR2X0 U13965 ( .IN1(n11055), .IN2(n13908), .QN(n13907) );
  NOR2X0 U13966 ( .IN1(n5666), .IN2(n13077), .QN(n13908) );
  NAND2X0 U13967 ( .IN1(n13909), .IN2(n13910), .QN(g33571) );
  NAND2X0 U13968 ( .IN1(n11442), .IN2(g2089), .QN(n13910) );
  INVX0 U13969 ( .INP(n11443), .ZN(n11442) );
  NAND2X0 U13970 ( .IN1(n11443), .IN2(g2084), .QN(n13909) );
  NAND2X0 U13971 ( .IN1(n13077), .IN2(n10961), .QN(n11443) );
  NAND2X0 U13972 ( .IN1(n13911), .IN2(n5535), .QN(n13077) );
  NOR2X0 U13973 ( .IN1(n13098), .IN2(g1996), .QN(n13911) );
  NAND2X0 U13974 ( .IN1(n13912), .IN2(n13913), .QN(g33570) );
  NAND2X0 U13975 ( .IN1(n11066), .IN2(g2040), .QN(n13913) );
  NOR2X0 U13976 ( .IN1(n13914), .IN2(n13915), .QN(n13912) );
  NOR2X0 U13977 ( .IN1(n13885), .IN2(n13114), .QN(n13915) );
  NAND2X0 U13978 ( .IN1(g2040), .IN2(n13091), .QN(n13114) );
  NOR2X0 U13979 ( .IN1(n5535), .IN2(n13916), .QN(n13914) );
  INVX0 U13980 ( .INP(n13917), .ZN(n13916) );
  NAND2X0 U13981 ( .IN1(n13918), .IN2(n13919), .QN(g33569) );
  NAND2X0 U13982 ( .IN1(n13917), .IN2(g2040), .QN(n13919) );
  NOR2X0 U13983 ( .IN1(n13920), .IN2(n13921), .QN(n13918) );
  NOR2X0 U13984 ( .IN1(n11054), .IN2(n13922), .QN(n13921) );
  NAND2X0 U13985 ( .IN1(n13144), .IN2(n13923), .QN(n13922) );
  NOR2X0 U13986 ( .IN1(n5355), .IN2(n13098), .QN(n13144) );
  NOR2X0 U13987 ( .IN1(n5831), .IN2(n10848), .QN(n13920) );
  NAND2X0 U13988 ( .IN1(n13924), .IN2(n13925), .QN(g33568) );
  NAND2X0 U13989 ( .IN1(n13926), .IN2(n13927), .QN(n13925) );
  NOR2X0 U13990 ( .IN1(n11054), .IN2(n13885), .QN(n13927) );
  INVX0 U13991 ( .INP(n13923), .ZN(n13885) );
  NAND2X0 U13992 ( .IN1(n3115), .IN2(n12472), .QN(n13923) );
  NOR2X0 U13993 ( .IN1(n13928), .IN2(n12053), .QN(n12472) );
  NAND2X0 U13994 ( .IN1(g518), .IN2(n5519), .QN(n13928) );
  NOR2X0 U13995 ( .IN1(n13929), .IN2(g2070), .QN(n13926) );
  NOR2X0 U13996 ( .IN1(n13930), .IN2(g1996), .QN(n13929) );
  NOR2X0 U13997 ( .IN1(n13098), .IN2(g2040), .QN(n13930) );
  NAND2X0 U13998 ( .IN1(n13917), .IN2(g1996), .QN(n13924) );
  NOR2X0 U13999 ( .IN1(n13091), .IN2(n11018), .QN(n13917) );
  INVX0 U14000 ( .INP(n13098), .ZN(n13091) );
  NOR2X0 U14001 ( .IN1(n13095), .IN2(n13888), .QN(n13098) );
  NOR2X0 U14002 ( .IN1(n13931), .IN2(n10548), .QN(n13888) );
  NOR2X0 U14003 ( .IN1(n13932), .IN2(g1171), .QN(n13931) );
  NAND2X0 U14004 ( .IN1(n13933), .IN2(n13934), .QN(n13095) );
  NAND2X0 U14005 ( .IN1(n5286), .IN2(g956), .QN(n13934) );
  NOR2X0 U14006 ( .IN1(n13354), .IN2(n13935), .QN(n13933) );
  NOR2X0 U14007 ( .IN1(n5275), .IN2(n13936), .QN(n13935) );
  NAND2X0 U14008 ( .IN1(n13937), .IN2(n13938), .QN(g33567) );
  NAND2X0 U14009 ( .IN1(test_so8), .IN2(n11081), .QN(n13938) );
  NOR2X0 U14010 ( .IN1(n13939), .IN2(n13940), .QN(n13937) );
  NOR2X0 U14011 ( .IN1(n5828), .IN2(n13941), .QN(n13940) );
  NOR2X0 U14012 ( .IN1(n13942), .IN2(n13649), .QN(n13941) );
  NOR2X0 U14013 ( .IN1(n11054), .IN2(n13943), .QN(n13942) );
  NOR2X0 U14014 ( .IN1(n12466), .IN2(n13944), .QN(n13943) );
  NOR2X0 U14015 ( .IN1(n13945), .IN2(n13944), .QN(n13939) );
  NOR2X0 U14016 ( .IN1(n13946), .IN2(n13947), .QN(n13945) );
  NOR2X0 U14017 ( .IN1(n13948), .IN2(g112), .QN(n13947) );
  NOR2X0 U14018 ( .IN1(n13949), .IN2(n13950), .QN(n13948) );
  NOR2X0 U14019 ( .IN1(n11054), .IN2(n13951), .QN(n13950) );
  NOR2X0 U14020 ( .IN1(n12466), .IN2(n13952), .QN(n13949) );
  INVX0 U14021 ( .INP(n13953), .ZN(n13952) );
  NOR2X0 U14022 ( .IN1(n12495), .IN2(n13657), .QN(n13953) );
  NOR2X0 U14023 ( .IN1(n13951), .IN2(n13954), .QN(n13946) );
  NAND2X0 U14024 ( .IN1(n12495), .IN2(n10961), .QN(n13954) );
  NAND2X0 U14025 ( .IN1(n5503), .IN2(g1936), .QN(n12495) );
  INVX0 U14026 ( .INP(n13955), .ZN(n13951) );
  NAND2X0 U14027 ( .IN1(n13956), .IN2(n13957), .QN(g33566) );
  NAND2X0 U14028 ( .IN1(n11485), .IN2(g1982), .QN(n13957) );
  NOR2X0 U14029 ( .IN1(n13958), .IN2(n13959), .QN(n13956) );
  NOR2X0 U14030 ( .IN1(n5845), .IN2(n10848), .QN(n13959) );
  NOR2X0 U14031 ( .IN1(n11054), .IN2(n13960), .QN(n13958) );
  NAND2X0 U14032 ( .IN1(n5462), .IN2(n13170), .QN(n13960) );
  INVX0 U14033 ( .INP(n13150), .ZN(n13170) );
  NAND2X0 U14034 ( .IN1(n13961), .IN2(n13962), .QN(g33565) );
  NAND2X0 U14035 ( .IN1(n11485), .IN2(g1978), .QN(n13962) );
  NOR2X0 U14036 ( .IN1(n13963), .IN2(n13964), .QN(n13961) );
  NOR2X0 U14037 ( .IN1(g1974), .IN2(n13965), .QN(n13964) );
  NAND2X0 U14038 ( .IN1(n13966), .IN2(n5664), .QN(n13965) );
  NOR2X0 U14039 ( .IN1(n11054), .IN2(n13150), .QN(n13966) );
  NOR2X0 U14040 ( .IN1(n5450), .IN2(n13967), .QN(n13963) );
  NOR2X0 U14041 ( .IN1(n11054), .IN2(n13968), .QN(n13967) );
  NOR2X0 U14042 ( .IN1(n5664), .IN2(n13150), .QN(n13968) );
  NAND2X0 U14043 ( .IN1(n13969), .IN2(n13970), .QN(g33563) );
  NAND2X0 U14044 ( .IN1(n11485), .IN2(g1955), .QN(n13970) );
  INVX0 U14045 ( .INP(n11486), .ZN(n11485) );
  NAND2X0 U14046 ( .IN1(n11486), .IN2(g1950), .QN(n13969) );
  NAND2X0 U14047 ( .IN1(n13150), .IN2(n10960), .QN(n11486) );
  NAND2X0 U14048 ( .IN1(n13971), .IN2(n5534), .QN(n13150) );
  NOR2X0 U14049 ( .IN1(test_so8), .IN2(n13171), .QN(n13971) );
  NAND2X0 U14050 ( .IN1(n13972), .IN2(n13973), .QN(g33562) );
  NAND2X0 U14051 ( .IN1(n11066), .IN2(g1906), .QN(n13973) );
  NOR2X0 U14052 ( .IN1(n13974), .IN2(n13975), .QN(n13972) );
  NOR2X0 U14053 ( .IN1(n13955), .IN2(n13187), .QN(n13975) );
  NAND2X0 U14054 ( .IN1(g1906), .IN2(n13164), .QN(n13187) );
  NOR2X0 U14055 ( .IN1(n5534), .IN2(n13976), .QN(n13974) );
  INVX0 U14056 ( .INP(n13977), .ZN(n13976) );
  NAND2X0 U14057 ( .IN1(n13978), .IN2(n13979), .QN(g33561) );
  NAND2X0 U14058 ( .IN1(n13977), .IN2(g1906), .QN(n13979) );
  NOR2X0 U14059 ( .IN1(n13980), .IN2(n13981), .QN(n13978) );
  INVX0 U14060 ( .INP(n13982), .ZN(n13981) );
  NAND2X0 U14061 ( .IN1(n10920), .IN2(n13983), .QN(n13982) );
  NOR2X0 U14062 ( .IN1(n13195), .IN2(n13955), .QN(n13983) );
  NAND2X0 U14063 ( .IN1(test_so8), .IN2(n13164), .QN(n13195) );
  NOR2X0 U14064 ( .IN1(n5828), .IN2(n10848), .QN(n13980) );
  NAND2X0 U14065 ( .IN1(n13984), .IN2(n13985), .QN(g33560) );
  NAND2X0 U14066 ( .IN1(n13986), .IN2(n13987), .QN(n13985) );
  NOR2X0 U14067 ( .IN1(n11054), .IN2(n13955), .QN(n13987) );
  NOR2X0 U14068 ( .IN1(n13806), .IN2(n12466), .QN(n13955) );
  NAND2X0 U14069 ( .IN1(n13988), .IN2(n3195), .QN(n12466) );
  NOR2X0 U14070 ( .IN1(n5519), .IN2(n5287), .QN(n13988) );
  NOR2X0 U14071 ( .IN1(n13989), .IN2(g1936), .QN(n13986) );
  NOR2X0 U14072 ( .IN1(n13990), .IN2(test_so8), .QN(n13989) );
  NOR2X0 U14073 ( .IN1(n13171), .IN2(g1906), .QN(n13990) );
  INVX0 U14074 ( .INP(n13164), .ZN(n13171) );
  NAND2X0 U14075 ( .IN1(n13977), .IN2(test_so8), .QN(n13984) );
  NOR2X0 U14076 ( .IN1(n13164), .IN2(n11016), .QN(n13977) );
  NAND2X0 U14077 ( .IN1(n13210), .IN2(n13944), .QN(n13164) );
  NAND2X0 U14078 ( .IN1(g17400), .IN2(n13991), .QN(n13944) );
  NAND2X0 U14079 ( .IN1(n13992), .IN2(n13993), .QN(n13991) );
  INVX0 U14080 ( .INP(n13168), .ZN(n13210) );
  NAND2X0 U14081 ( .IN1(n13994), .IN2(n13995), .QN(n13168) );
  NAND2X0 U14082 ( .IN1(n5286), .IN2(g1129), .QN(n13995) );
  NOR2X0 U14083 ( .IN1(n13354), .IN2(n13996), .QN(n13994) );
  NOR2X0 U14084 ( .IN1(g2145), .IN2(n13997), .QN(n13996) );
  NAND2X0 U14085 ( .IN1(g2138), .IN2(g2130), .QN(n13997) );
  NAND2X0 U14086 ( .IN1(n13998), .IN2(n13999), .QN(g33559) );
  NAND2X0 U14087 ( .IN1(n11066), .IN2(g1728), .QN(n13999) );
  NOR2X0 U14088 ( .IN1(n14000), .IN2(n14001), .QN(n13998) );
  NOR2X0 U14089 ( .IN1(n5830), .IN2(n14002), .QN(n14001) );
  NOR2X0 U14090 ( .IN1(n14003), .IN2(n13649), .QN(n14002) );
  INVX0 U14091 ( .INP(n14004), .ZN(n13649) );
  NOR2X0 U14092 ( .IN1(n11053), .IN2(n14005), .QN(n14003) );
  NOR2X0 U14093 ( .IN1(n12468), .IN2(n14006), .QN(n14005) );
  NOR2X0 U14094 ( .IN1(n14006), .IN2(n14007), .QN(n14000) );
  NAND2X0 U14095 ( .IN1(n14008), .IN2(n14009), .QN(n14007) );
  NAND2X0 U14096 ( .IN1(n14010), .IN2(n14011), .QN(n14009) );
  NAND2X0 U14097 ( .IN1(n14012), .IN2(n14013), .QN(n14011) );
  NOR2X0 U14098 ( .IN1(n5536), .IN2(n13657), .QN(n14013) );
  NOR2X0 U14099 ( .IN1(n12468), .IN2(g1772), .QN(n14012) );
  NAND2X0 U14100 ( .IN1(n14014), .IN2(n10960), .QN(n14010) );
  NAND2X0 U14101 ( .IN1(n14015), .IN2(n5504), .QN(n14008) );
  NOR2X0 U14102 ( .IN1(n5536), .IN2(n10273), .QN(n14015) );
  NAND2X0 U14103 ( .IN1(n14016), .IN2(n14017), .QN(g33558) );
  NAND2X0 U14104 ( .IN1(n11323), .IN2(g1848), .QN(n14017) );
  NOR2X0 U14105 ( .IN1(n14018), .IN2(n14019), .QN(n14016) );
  NOR2X0 U14106 ( .IN1(n5847), .IN2(n10847), .QN(n14019) );
  NOR2X0 U14107 ( .IN1(n11053), .IN2(n14020), .QN(n14018) );
  NAND2X0 U14108 ( .IN1(n5464), .IN2(n13240), .QN(n14020) );
  INVX0 U14109 ( .INP(n13220), .ZN(n13240) );
  NAND2X0 U14110 ( .IN1(n14021), .IN2(n14022), .QN(g33557) );
  NAND2X0 U14111 ( .IN1(n11323), .IN2(g1844), .QN(n14022) );
  NOR2X0 U14112 ( .IN1(n14023), .IN2(n14024), .QN(n14021) );
  NOR2X0 U14113 ( .IN1(g1840), .IN2(n14025), .QN(n14024) );
  NAND2X0 U14114 ( .IN1(n14026), .IN2(n5665), .QN(n14025) );
  NOR2X0 U14115 ( .IN1(n11053), .IN2(n13220), .QN(n14026) );
  NOR2X0 U14116 ( .IN1(n5451), .IN2(n14027), .QN(n14023) );
  NOR2X0 U14117 ( .IN1(n11053), .IN2(n14028), .QN(n14027) );
  NOR2X0 U14118 ( .IN1(n5665), .IN2(n13220), .QN(n14028) );
  NAND2X0 U14119 ( .IN1(n14029), .IN2(n14030), .QN(g33555) );
  NAND2X0 U14120 ( .IN1(n11323), .IN2(g1821), .QN(n14030) );
  INVX0 U14121 ( .INP(n11324), .ZN(n11323) );
  NAND2X0 U14122 ( .IN1(n11324), .IN2(g1816), .QN(n14029) );
  NAND2X0 U14123 ( .IN1(n13220), .IN2(n10960), .QN(n11324) );
  NAND2X0 U14124 ( .IN1(n14031), .IN2(n5536), .QN(n13220) );
  NOR2X0 U14125 ( .IN1(n13241), .IN2(g1728), .QN(n14031) );
  NAND2X0 U14126 ( .IN1(n14032), .IN2(n14033), .QN(g33554) );
  INVX0 U14127 ( .INP(n14034), .ZN(n14033) );
  NOR2X0 U14128 ( .IN1(n13258), .IN2(n14014), .QN(n14034) );
  NAND2X0 U14129 ( .IN1(g1772), .IN2(n13234), .QN(n13258) );
  NOR2X0 U14130 ( .IN1(n14035), .IN2(n14036), .QN(n14032) );
  NOR2X0 U14131 ( .IN1(n11053), .IN2(n14037), .QN(n14036) );
  NAND2X0 U14132 ( .IN1(n13241), .IN2(g1802), .QN(n14037) );
  NOR2X0 U14133 ( .IN1(n5504), .IN2(n10847), .QN(n14035) );
  NAND2X0 U14134 ( .IN1(n14038), .IN2(n14039), .QN(g33553) );
  NAND2X0 U14135 ( .IN1(n14040), .IN2(n13228), .QN(n14039) );
  NOR2X0 U14136 ( .IN1(n13241), .IN2(n14014), .QN(n14040) );
  NOR2X0 U14137 ( .IN1(n14041), .IN2(n14042), .QN(n14038) );
  NOR2X0 U14138 ( .IN1(n5830), .IN2(n10847), .QN(n14042) );
  NOR2X0 U14139 ( .IN1(n11053), .IN2(n14043), .QN(n14041) );
  NAND2X0 U14140 ( .IN1(n13241), .IN2(g1772), .QN(n14043) );
  NAND2X0 U14141 ( .IN1(n14044), .IN2(n14045), .QN(g33552) );
  NAND2X0 U14142 ( .IN1(n14046), .IN2(n14047), .QN(n14045) );
  NOR2X0 U14143 ( .IN1(n11053), .IN2(n14014), .QN(n14047) );
  NOR2X0 U14144 ( .IN1(n13806), .IN2(n12468), .QN(n14014) );
  NAND2X0 U14145 ( .IN1(n13807), .IN2(n3195), .QN(n12468) );
  NOR2X0 U14146 ( .IN1(n5519), .IN2(g518), .QN(n13807) );
  INVX0 U14147 ( .INP(n3115), .ZN(n13806) );
  NOR2X0 U14148 ( .IN1(n14048), .IN2(g1802), .QN(n14046) );
  NOR2X0 U14149 ( .IN1(n14049), .IN2(g1728), .QN(n14048) );
  NOR2X0 U14150 ( .IN1(n13241), .IN2(g1772), .QN(n14049) );
  NAND2X0 U14151 ( .IN1(n13228), .IN2(n13241), .QN(n14044) );
  INVX0 U14152 ( .INP(n13234), .ZN(n13241) );
  NAND2X0 U14153 ( .IN1(n13280), .IN2(n14006), .QN(n13234) );
  NAND2X0 U14154 ( .IN1(test_so44), .IN2(n14050), .QN(n14006) );
  NAND2X0 U14155 ( .IN1(n14051), .IN2(n13993), .QN(n14050) );
  INVX0 U14156 ( .INP(n13238), .ZN(n13280) );
  NAND2X0 U14157 ( .IN1(n14052), .IN2(n14053), .QN(n13238) );
  NAND2X0 U14158 ( .IN1(n5286), .IN2(g1105), .QN(n14053) );
  NOR2X0 U14159 ( .IN1(n13354), .IN2(n14054), .QN(n14052) );
  NOR2X0 U14160 ( .IN1(g2138), .IN2(n13936), .QN(n14054) );
  NAND2X0 U14161 ( .IN1(g2145), .IN2(g2130), .QN(n13936) );
  NOR2X0 U14162 ( .IN1(n11053), .IN2(n5352), .QN(n13228) );
  NAND2X0 U14163 ( .IN1(n14055), .IN2(n14056), .QN(g33551) );
  NOR2X0 U14164 ( .IN1(n14057), .IN2(n14058), .QN(n14056) );
  NOR2X0 U14165 ( .IN1(n11053), .IN2(n14059), .QN(n14058) );
  NOR2X0 U14166 ( .IN1(n14060), .IN2(n14061), .QN(n14059) );
  NOR2X0 U14167 ( .IN1(n14062), .IN2(n10646), .QN(n14061) );
  INVX0 U14168 ( .INP(n14063), .ZN(n14062) );
  NAND2X0 U14169 ( .IN1(n12471), .IN2(g33533), .QN(n14063) );
  NOR2X0 U14170 ( .IN1(n14064), .IN2(n14065), .QN(n14060) );
  NAND2X0 U14171 ( .IN1(g33533), .IN2(n14066), .QN(n14065) );
  NAND2X0 U14172 ( .IN1(g31862), .IN2(g112), .QN(n14066) );
  NOR2X0 U14173 ( .IN1(n5362), .IN2(n10847), .QN(n14057) );
  NOR2X0 U14174 ( .IN1(n14067), .IN2(n14068), .QN(n14055) );
  NOR2X0 U14175 ( .IN1(n14004), .IN2(n10646), .QN(n14068) );
  NOR2X0 U14176 ( .IN1(n14069), .IN2(n14070), .QN(n14067) );
  NAND2X0 U14177 ( .IN1(g33533), .IN2(g31862), .QN(n14070) );
  NAND2X0 U14178 ( .IN1(n14071), .IN2(n12471), .QN(n14069) );
  NOR2X0 U14179 ( .IN1(n13657), .IN2(g112), .QN(n14071) );
  NAND2X0 U14180 ( .IN1(n14072), .IN2(n14073), .QN(g33550) );
  NAND2X0 U14181 ( .IN1(n14074), .IN2(g1714), .QN(n14073) );
  NOR2X0 U14182 ( .IN1(n14075), .IN2(n14076), .QN(n14072) );
  NOR2X0 U14183 ( .IN1(n5412), .IN2(n10846), .QN(n14076) );
  NOR2X0 U14184 ( .IN1(n11053), .IN2(n14077), .QN(n14075) );
  NAND2X0 U14185 ( .IN1(n5460), .IN2(n13312), .QN(n14077) );
  INVX0 U14186 ( .INP(n13292), .ZN(n13312) );
  NAND2X0 U14187 ( .IN1(n14078), .IN2(n14079), .QN(g33549) );
  NAND2X0 U14188 ( .IN1(n14074), .IN2(g1710), .QN(n14079) );
  NOR2X0 U14189 ( .IN1(n14080), .IN2(n14081), .QN(n14078) );
  NOR2X0 U14190 ( .IN1(test_so15), .IN2(n14082), .QN(n14081) );
  NAND2X0 U14191 ( .IN1(n14083), .IN2(n5417), .QN(n14082) );
  NOR2X0 U14192 ( .IN1(n11052), .IN2(n13292), .QN(n14083) );
  NOR2X0 U14193 ( .IN1(n14084), .IN2(n10678), .QN(n14080) );
  NOR2X0 U14194 ( .IN1(n11052), .IN2(n14085), .QN(n14084) );
  NOR2X0 U14195 ( .IN1(n5417), .IN2(n13292), .QN(n14085) );
  NAND2X0 U14196 ( .IN1(n14086), .IN2(n14087), .QN(g33548) );
  NAND2X0 U14197 ( .IN1(test_so15), .IN2(n14074), .QN(n14087) );
  NAND2X0 U14198 ( .IN1(n13290), .IN2(g1700), .QN(n14086) );
  NAND2X0 U14199 ( .IN1(n14088), .IN2(n14089), .QN(g33547) );
  NAND2X0 U14200 ( .IN1(n14074), .IN2(g1687), .QN(n14089) );
  INVX0 U14201 ( .INP(n13290), .ZN(n14074) );
  NAND2X0 U14202 ( .IN1(n13290), .IN2(g1682), .QN(n14088) );
  NAND2X0 U14203 ( .IN1(n13292), .IN2(n10959), .QN(n13290) );
  NAND2X0 U14204 ( .IN1(n14090), .IN2(n5598), .QN(n13292) );
  NOR2X0 U14205 ( .IN1(n13313), .IN2(g1592), .QN(n14090) );
  NAND2X0 U14206 ( .IN1(n14091), .IN2(n14092), .QN(g33546) );
  NAND2X0 U14207 ( .IN1(n11066), .IN2(g1636), .QN(n14092) );
  NOR2X0 U14208 ( .IN1(n14093), .IN2(n14094), .QN(n14091) );
  NOR2X0 U14209 ( .IN1(n14095), .IN2(n13329), .QN(n14094) );
  NAND2X0 U14210 ( .IN1(g1636), .IN2(n13306), .QN(n13329) );
  NOR2X0 U14211 ( .IN1(n5598), .IN2(n14096), .QN(n14093) );
  INVX0 U14212 ( .INP(n14097), .ZN(n14096) );
  NAND2X0 U14213 ( .IN1(n14098), .IN2(n14099), .QN(g33545) );
  NAND2X0 U14214 ( .IN1(n14097), .IN2(g1636), .QN(n14099) );
  NOR2X0 U14215 ( .IN1(n14100), .IN2(n14101), .QN(n14098) );
  NOR2X0 U14216 ( .IN1(n11052), .IN2(n14102), .QN(n14101) );
  NAND2X0 U14217 ( .IN1(n13337), .IN2(n14064), .QN(n14102) );
  NOR2X0 U14218 ( .IN1(n5362), .IN2(n13313), .QN(n13337) );
  NOR2X0 U14219 ( .IN1(n10904), .IN2(n10646), .QN(n14100) );
  NAND2X0 U14220 ( .IN1(n14103), .IN2(n14104), .QN(g33544) );
  NAND2X0 U14221 ( .IN1(n14105), .IN2(n14106), .QN(n14104) );
  NOR2X0 U14222 ( .IN1(n11052), .IN2(n14095), .QN(n14106) );
  INVX0 U14223 ( .INP(n14064), .ZN(n14095) );
  NAND2X0 U14224 ( .IN1(n3115), .IN2(n12471), .QN(n14064) );
  NOR2X0 U14225 ( .IN1(n14107), .IN2(n12053), .QN(n12471) );
  INVX0 U14226 ( .INP(n3195), .ZN(n12053) );
  NAND2X0 U14227 ( .IN1(n5287), .IN2(n5519), .QN(n14107) );
  NOR2X0 U14228 ( .IN1(n14108), .IN2(g1668), .QN(n14105) );
  NOR2X0 U14229 ( .IN1(n14109), .IN2(g1592), .QN(n14108) );
  NOR2X0 U14230 ( .IN1(n13313), .IN2(g1636), .QN(n14109) );
  NAND2X0 U14231 ( .IN1(n14097), .IN2(g1592), .QN(n14103) );
  NOR2X0 U14232 ( .IN1(n13306), .IN2(n11016), .QN(n14097) );
  INVX0 U14233 ( .INP(n13313), .ZN(n13306) );
  NOR2X0 U14234 ( .IN1(n13310), .IN2(g33533), .QN(n13313) );
  NAND2X0 U14235 ( .IN1(n14110), .IN2(n14111), .QN(n13310) );
  NAND2X0 U14236 ( .IN1(n5286), .IN2(g1135), .QN(n14111) );
  NOR2X0 U14237 ( .IN1(n13354), .IN2(n14112), .QN(n14110) );
  NOR2X0 U14238 ( .IN1(g2145), .IN2(n14113), .QN(n14112) );
  NAND2X0 U14239 ( .IN1(n5275), .IN2(g2130), .QN(n14113) );
  NOR2X0 U14240 ( .IN1(n14114), .IN2(g134), .QN(n13354) );
  NOR2X0 U14241 ( .IN1(n11987), .IN2(n11992), .QN(n14114) );
  NAND2X0 U14242 ( .IN1(n5595), .IN2(g691), .QN(n11992) );
  NAND2X0 U14243 ( .IN1(n14115), .IN2(n14116), .QN(g33543) );
  NAND2X0 U14244 ( .IN1(n14117), .IN2(n14118), .QN(n14116) );
  NAND2X0 U14245 ( .IN1(n14119), .IN2(n14120), .QN(n14118) );
  NAND2X0 U14246 ( .IN1(n10259), .IN2(n14121), .QN(n14120) );
  INVX0 U14247 ( .INP(n14122), .ZN(n14119) );
  NOR2X0 U14248 ( .IN1(n10190), .IN2(n11016), .QN(n14117) );
  NAND2X0 U14249 ( .IN1(n14123), .IN2(g1373), .QN(n14115) );
  NAND2X0 U14250 ( .IN1(n14124), .IN2(n10959), .QN(n14123) );
  NAND2X0 U14251 ( .IN1(n14125), .IN2(n10190), .QN(n14124) );
  NOR2X0 U14252 ( .IN1(n14126), .IN2(n14122), .QN(n14125) );
  NAND2X0 U14253 ( .IN1(n14127), .IN2(n14128), .QN(g33542) );
  NAND2X0 U14254 ( .IN1(n11066), .IN2(g1270), .QN(n14128) );
  NOR2X0 U14255 ( .IN1(n14129), .IN2(n14130), .QN(n14127) );
  NOR2X0 U14256 ( .IN1(n14131), .IN2(g1274), .QN(n14130) );
  NOR2X0 U14257 ( .IN1(n5730), .IN2(n14132), .QN(n14129) );
  NAND2X0 U14258 ( .IN1(n14133), .IN2(n14131), .QN(n14132) );
  NAND2X0 U14259 ( .IN1(n14134), .IN2(n14135), .QN(g33541) );
  NAND2X0 U14260 ( .IN1(n14136), .IN2(n14137), .QN(n14135) );
  NAND2X0 U14261 ( .IN1(n14138), .IN2(n14139), .QN(n14137) );
  NAND2X0 U14262 ( .IN1(n10261), .IN2(n14140), .QN(n14139) );
  INVX0 U14263 ( .INP(n14141), .ZN(n14138) );
  NOR2X0 U14264 ( .IN1(n10191), .IN2(n11016), .QN(n14136) );
  NAND2X0 U14265 ( .IN1(n14142), .IN2(g1030), .QN(n14134) );
  NAND2X0 U14266 ( .IN1(n14143), .IN2(n10959), .QN(n14142) );
  NAND2X0 U14267 ( .IN1(n14144), .IN2(n10191), .QN(n14143) );
  NOR2X0 U14268 ( .IN1(n14145), .IN2(n14141), .QN(n14144) );
  NAND2X0 U14269 ( .IN1(n14146), .IN2(n14147), .QN(g33540) );
  NAND2X0 U14270 ( .IN1(n11066), .IN2(g925), .QN(n14147) );
  NOR2X0 U14271 ( .IN1(n14148), .IN2(n14149), .QN(n14146) );
  NOR2X0 U14272 ( .IN1(n14150), .IN2(g930), .QN(n14149) );
  NOR2X0 U14273 ( .IN1(n5731), .IN2(n14151), .QN(n14148) );
  NAND2X0 U14274 ( .IN1(n14152), .IN2(n14150), .QN(n14151) );
  NAND2X0 U14275 ( .IN1(n14153), .IN2(n14154), .QN(g33539) );
  NAND2X0 U14276 ( .IN1(n11066), .IN2(g758), .QN(n14154) );
  NOR2X0 U14277 ( .IN1(n14155), .IN2(n14156), .QN(n14153) );
  NOR2X0 U14278 ( .IN1(g763), .IN2(n14157), .QN(n14156) );
  NOR2X0 U14279 ( .IN1(n5332), .IN2(n14158), .QN(n14155) );
  NAND2X0 U14280 ( .IN1(n2404), .IN2(n14157), .QN(n14158) );
  INVX0 U14281 ( .INP(n2980), .ZN(n14157) );
  NAND2X0 U14282 ( .IN1(n14159), .IN2(n14160), .QN(g33538) );
  NAND2X0 U14283 ( .IN1(n11066), .IN2(g590), .QN(n14160) );
  NOR2X0 U14284 ( .IN1(n14161), .IN2(n14162), .QN(n14159) );
  NOR2X0 U14285 ( .IN1(g595), .IN2(n14163), .QN(n14162) );
  NOR2X0 U14286 ( .IN1(n5476), .IN2(n14164), .QN(n14161) );
  NAND2X0 U14287 ( .IN1(n2421), .IN2(n14163), .QN(n14164) );
  INVX0 U14288 ( .INP(n2982), .ZN(n14163) );
  NAND2X0 U14289 ( .IN1(n14165), .IN2(n14166), .QN(g33537) );
  NAND2X0 U14290 ( .IN1(n11066), .IN2(g301), .QN(n14166) );
  NAND2X0 U14291 ( .IN1(n14167), .IN2(n10959), .QN(n14165) );
  NOR2X0 U14292 ( .IN1(n5724), .IN2(n12633), .QN(n14167) );
  INVX0 U14293 ( .INP(n2707), .ZN(n12633) );
  NOR2X0 U14294 ( .IN1(n5843), .IN2(n14168), .QN(g33536) );
  NOR2X0 U14295 ( .IN1(n2710), .IN2(n11017), .QN(n14168) );
  NAND2X0 U14296 ( .IN1(n14169), .IN2(n14170), .QN(g33535) );
  NAND2X0 U14297 ( .IN1(n11066), .IN2(g291), .QN(n14170) );
  NOR2X0 U14298 ( .IN1(n14171), .IN2(n14172), .QN(n14169) );
  NOR2X0 U14299 ( .IN1(g294), .IN2(n14173), .QN(n14172) );
  NOR2X0 U14300 ( .IN1(n5680), .IN2(n14174), .QN(n14171) );
  NAND2X0 U14301 ( .IN1(n95), .IN2(n14173), .QN(n14174) );
  INVX0 U14302 ( .INP(n3276), .ZN(n14173) );
  NAND2X0 U14303 ( .IN1(n14175), .IN2(n14176), .QN(g33534) );
  NAND2X0 U14304 ( .IN1(n11066), .IN2(g150), .QN(n14176) );
  NOR2X0 U14305 ( .IN1(n14177), .IN2(n14178), .QN(n14175) );
  NOR2X0 U14306 ( .IN1(g153), .IN2(n14179), .QN(n14178) );
  NOR2X0 U14307 ( .IN1(n5677), .IN2(n14180), .QN(n14177) );
  NAND2X0 U14308 ( .IN1(n12641), .IN2(n14179), .QN(n14180) );
  INVX0 U14309 ( .INP(n3277), .ZN(n14179) );
  NOR2X0 U14310 ( .IN1(n14181), .IN2(n10218), .QN(g33533) );
  NOR2X0 U14311 ( .IN1(n13932), .IN2(n5363), .QN(n14181) );
  NAND2X0 U14312 ( .IN1(n5599), .IN2(n13993), .QN(n13932) );
  INVX0 U14313 ( .INP(n14182), .ZN(n13993) );
  NAND2X0 U14314 ( .IN1(n14183), .IN2(n14184), .QN(n14182) );
  NOR2X0 U14315 ( .IN1(n10252), .IN2(n14185), .QN(n14184) );
  NAND2X0 U14316 ( .IN1(g979), .IN2(n10673), .QN(n14185) );
  NOR2X0 U14317 ( .IN1(g1205), .IN2(n14186), .QN(n14183) );
  NAND2X0 U14318 ( .IN1(n5442), .IN2(n10547), .QN(n14186) );
  NOR2X0 U14319 ( .IN1(n14187), .IN2(n14188), .QN(g33435) );
  NAND2X0 U14320 ( .IN1(n14189), .IN2(n14190), .QN(n14188) );
  NAND2X0 U14321 ( .IN1(n14191), .IN2(g2724), .QN(n14190) );
  NOR2X0 U14322 ( .IN1(n14192), .IN2(n14193), .QN(n14191) );
  NOR2X0 U14323 ( .IN1(g2729), .IN2(g2775), .QN(n14193) );
  NOR2X0 U14324 ( .IN1(n10274), .IN2(g2787), .QN(n14192) );
  NAND2X0 U14325 ( .IN1(n12398), .IN2(g2771), .QN(n14189) );
  NOR2X0 U14326 ( .IN1(n5403), .IN2(n12389), .QN(n14187) );
  NOR2X0 U14327 ( .IN1(n14194), .IN2(n14195), .QN(g33079) );
  NAND2X0 U14328 ( .IN1(n14196), .IN2(n14197), .QN(n14195) );
  NAND2X0 U14329 ( .IN1(n14198), .IN2(g2724), .QN(n14197) );
  NOR2X0 U14330 ( .IN1(n14199), .IN2(n14200), .QN(n14198) );
  NOR2X0 U14331 ( .IN1(g2729), .IN2(g2807), .QN(n14200) );
  NOR2X0 U14332 ( .IN1(n10274), .IN2(g2819), .QN(n14199) );
  NAND2X0 U14333 ( .IN1(n12398), .IN2(g2803), .QN(n14196) );
  NOR2X0 U14334 ( .IN1(n5404), .IN2(n12389), .QN(n14194) );
  NAND2X0 U14335 ( .IN1(n5301), .IN2(g2729), .QN(n12389) );
  NAND2X0 U14336 ( .IN1(n14201), .IN2(n14202), .QN(g33070) );
  NAND2X0 U14337 ( .IN1(n14203), .IN2(n14204), .QN(n14202) );
  NAND2X0 U14338 ( .IN1(n14205), .IN2(n14206), .QN(n14203) );
  NAND2X0 U14339 ( .IN1(n10926), .IN2(n14207), .QN(n14206) );
  NOR2X0 U14340 ( .IN1(n14208), .IN2(n14209), .QN(n14205) );
  INVX0 U14341 ( .INP(n14210), .ZN(n14209) );
  NAND2X0 U14342 ( .IN1(n5646), .IN2(g25756), .QN(n14210) );
  NAND2X0 U14343 ( .IN1(n11066), .IN2(g6565), .QN(n14201) );
  NAND2X0 U14344 ( .IN1(n14211), .IN2(n14212), .QN(g33069) );
  NAND2X0 U14345 ( .IN1(n14213), .IN2(g6561), .QN(n14212) );
  NAND2X0 U14346 ( .IN1(n14214), .IN2(n10958), .QN(n14213) );
  NAND2X0 U14347 ( .IN1(n5386), .IN2(n14204), .QN(n14214) );
  NAND2X0 U14348 ( .IN1(n14215), .IN2(g6565), .QN(n14211) );
  INVX0 U14349 ( .INP(n14216), .ZN(n14215) );
  NAND2X0 U14350 ( .IN1(n14217), .IN2(n14218), .QN(g33068) );
  NAND2X0 U14351 ( .IN1(n14219), .IN2(n5646), .QN(n14218) );
  NOR2X0 U14352 ( .IN1(n3404), .IN2(n14220), .QN(n14219) );
  NAND2X0 U14353 ( .IN1(n11066), .IN2(g6555), .QN(n14217) );
  NAND2X0 U14354 ( .IN1(n14221), .IN2(n14222), .QN(g33067) );
  NAND2X0 U14355 ( .IN1(n14223), .IN2(n14204), .QN(n14222) );
  NAND2X0 U14356 ( .IN1(n3407), .IN2(n14224), .QN(n14223) );
  NAND2X0 U14357 ( .IN1(n10926), .IN2(n14225), .QN(n14224) );
  NAND2X0 U14358 ( .IN1(n11066), .IN2(g6549), .QN(n14221) );
  NAND2X0 U14359 ( .IN1(n14226), .IN2(n14227), .QN(g33065) );
  NAND2X0 U14360 ( .IN1(n14228), .IN2(n14229), .QN(n14227) );
  NAND2X0 U14361 ( .IN1(n14230), .IN2(n14231), .QN(n14228) );
  NAND2X0 U14362 ( .IN1(n10926), .IN2(n14232), .QN(n14231) );
  NOR2X0 U14363 ( .IN1(n14233), .IN2(n14234), .QN(n14230) );
  INVX0 U14364 ( .INP(n14235), .ZN(n14234) );
  NAND2X0 U14365 ( .IN1(n5651), .IN2(g25742), .QN(n14235) );
  NAND2X0 U14366 ( .IN1(n11066), .IN2(g6219), .QN(n14226) );
  NAND2X0 U14367 ( .IN1(n14236), .IN2(n14237), .QN(g33064) );
  NAND2X0 U14368 ( .IN1(n14238), .IN2(g6215), .QN(n14237) );
  NAND2X0 U14369 ( .IN1(n14239), .IN2(n10958), .QN(n14238) );
  NAND2X0 U14370 ( .IN1(n5385), .IN2(n14229), .QN(n14239) );
  NAND2X0 U14371 ( .IN1(n14240), .IN2(g6219), .QN(n14236) );
  INVX0 U14372 ( .INP(n14241), .ZN(n14240) );
  NAND2X0 U14373 ( .IN1(n14242), .IN2(n14243), .QN(g33063) );
  NAND2X0 U14374 ( .IN1(n14244), .IN2(n5651), .QN(n14243) );
  NOR2X0 U14375 ( .IN1(n3414), .IN2(n14245), .QN(n14244) );
  NAND2X0 U14376 ( .IN1(n11066), .IN2(g6209), .QN(n14242) );
  NAND2X0 U14377 ( .IN1(n14246), .IN2(n14247), .QN(g33062) );
  NAND2X0 U14378 ( .IN1(n14248), .IN2(n14229), .QN(n14247) );
  NAND2X0 U14379 ( .IN1(n3417), .IN2(n14249), .QN(n14248) );
  NAND2X0 U14380 ( .IN1(n10927), .IN2(n14250), .QN(n14249) );
  NAND2X0 U14381 ( .IN1(n11065), .IN2(g6203), .QN(n14246) );
  NAND2X0 U14382 ( .IN1(n14251), .IN2(n14252), .QN(g33060) );
  NAND2X0 U14383 ( .IN1(n14253), .IN2(n14254), .QN(n14252) );
  NAND2X0 U14384 ( .IN1(n14255), .IN2(n14256), .QN(n14253) );
  NAND2X0 U14385 ( .IN1(n10927), .IN2(n14257), .QN(n14256) );
  NOR2X0 U14386 ( .IN1(n14258), .IN2(n14259), .QN(n14255) );
  INVX0 U14387 ( .INP(n14260), .ZN(n14259) );
  NAND2X0 U14388 ( .IN1(n5649), .IN2(g25728), .QN(n14260) );
  NAND2X0 U14389 ( .IN1(n11065), .IN2(g5873), .QN(n14251) );
  NAND2X0 U14390 ( .IN1(n14261), .IN2(n14262), .QN(g33059) );
  NAND2X0 U14391 ( .IN1(n14263), .IN2(g5869), .QN(n14262) );
  NAND2X0 U14392 ( .IN1(n14264), .IN2(n10958), .QN(n14263) );
  NAND2X0 U14393 ( .IN1(n5388), .IN2(n14254), .QN(n14264) );
  NAND2X0 U14394 ( .IN1(n14265), .IN2(g5873), .QN(n14261) );
  INVX0 U14395 ( .INP(n14266), .ZN(n14265) );
  NAND2X0 U14396 ( .IN1(n14267), .IN2(n14268), .QN(g33058) );
  NAND2X0 U14397 ( .IN1(n14269), .IN2(n5649), .QN(n14268) );
  NOR2X0 U14398 ( .IN1(n3424), .IN2(n14270), .QN(n14269) );
  NAND2X0 U14399 ( .IN1(n11069), .IN2(g5863), .QN(n14267) );
  NAND2X0 U14400 ( .IN1(n14271), .IN2(n14272), .QN(g33057) );
  NAND2X0 U14401 ( .IN1(n14273), .IN2(n14254), .QN(n14272) );
  NAND2X0 U14402 ( .IN1(n3427), .IN2(n14274), .QN(n14273) );
  NAND2X0 U14403 ( .IN1(n14275), .IN2(n10957), .QN(n14274) );
  NAND2X0 U14404 ( .IN1(n11078), .IN2(g5857), .QN(n14271) );
  NAND2X0 U14405 ( .IN1(n14276), .IN2(n14277), .QN(g33055) );
  NAND2X0 U14406 ( .IN1(n14278), .IN2(n14279), .QN(n14277) );
  NAND2X0 U14407 ( .IN1(n14280), .IN2(n14281), .QN(n14278) );
  NAND2X0 U14408 ( .IN1(n10927), .IN2(n14282), .QN(n14281) );
  NOR2X0 U14409 ( .IN1(n14283), .IN2(n14284), .QN(n14280) );
  NOR2X0 U14410 ( .IN1(g5523), .IN2(n14285), .QN(n14284) );
  NAND2X0 U14411 ( .IN1(n11080), .IN2(g5527), .QN(n14276) );
  NAND2X0 U14412 ( .IN1(n14286), .IN2(n14287), .QN(g33054) );
  NAND2X0 U14413 ( .IN1(n14288), .IN2(g5523), .QN(n14287) );
  NAND2X0 U14414 ( .IN1(n14289), .IN2(n10957), .QN(n14288) );
  NAND2X0 U14415 ( .IN1(n5389), .IN2(n14279), .QN(n14289) );
  NAND2X0 U14416 ( .IN1(n14290), .IN2(g5527), .QN(n14286) );
  INVX0 U14417 ( .INP(n14291), .ZN(n14290) );
  NAND2X0 U14418 ( .IN1(n14292), .IN2(n14293), .QN(g33053) );
  NAND2X0 U14419 ( .IN1(n14294), .IN2(n5647), .QN(n14293) );
  NOR2X0 U14420 ( .IN1(n3434), .IN2(n14295), .QN(n14294) );
  NAND2X0 U14421 ( .IN1(n11079), .IN2(g5517), .QN(n14292) );
  NAND2X0 U14422 ( .IN1(n14296), .IN2(n14297), .QN(g33052) );
  NAND2X0 U14423 ( .IN1(n14298), .IN2(n14279), .QN(n14297) );
  NAND2X0 U14424 ( .IN1(n3437), .IN2(n14299), .QN(n14298) );
  NAND2X0 U14425 ( .IN1(n10927), .IN2(n14300), .QN(n14299) );
  NAND2X0 U14426 ( .IN1(n11080), .IN2(g5511), .QN(n14296) );
  NAND2X0 U14427 ( .IN1(n14301), .IN2(n14302), .QN(g33050) );
  NAND2X0 U14428 ( .IN1(n14303), .IN2(n14304), .QN(n14302) );
  NAND2X0 U14429 ( .IN1(n14305), .IN2(n14306), .QN(n14303) );
  NAND2X0 U14430 ( .IN1(n10927), .IN2(n14307), .QN(n14306) );
  NOR2X0 U14431 ( .IN1(n14308), .IN2(n14309), .QN(n14305) );
  INVX0 U14432 ( .INP(n14310), .ZN(n14309) );
  NAND2X0 U14433 ( .IN1(n5650), .IN2(g25700), .QN(n14310) );
  NAND2X0 U14434 ( .IN1(n11080), .IN2(g5180), .QN(n14301) );
  NAND2X0 U14435 ( .IN1(n14311), .IN2(n14312), .QN(g33049) );
  NAND2X0 U14436 ( .IN1(n14313), .IN2(g5176), .QN(n14312) );
  NAND2X0 U14437 ( .IN1(n14314), .IN2(n10957), .QN(n14313) );
  NAND2X0 U14438 ( .IN1(n5384), .IN2(n14304), .QN(n14314) );
  NAND2X0 U14439 ( .IN1(n14315), .IN2(g5180), .QN(n14311) );
  INVX0 U14440 ( .INP(n14316), .ZN(n14315) );
  NAND2X0 U14441 ( .IN1(n14317), .IN2(n14318), .QN(g33048) );
  NAND2X0 U14442 ( .IN1(n14319), .IN2(n5650), .QN(n14318) );
  NOR2X0 U14443 ( .IN1(n3444), .IN2(n14320), .QN(n14319) );
  NAND2X0 U14444 ( .IN1(n11079), .IN2(g5170), .QN(n14317) );
  NAND2X0 U14445 ( .IN1(n14321), .IN2(n14322), .QN(g33047) );
  NAND2X0 U14446 ( .IN1(n14323), .IN2(n14304), .QN(n14322) );
  NAND2X0 U14447 ( .IN1(n3447), .IN2(n14324), .QN(n14323) );
  NAND2X0 U14448 ( .IN1(n10927), .IN2(n14325), .QN(n14324) );
  NAND2X0 U14449 ( .IN1(n11080), .IN2(g5164), .QN(n14321) );
  NAND2X0 U14450 ( .IN1(n14326), .IN2(n14327), .QN(g33046) );
  NAND2X0 U14451 ( .IN1(n11079), .IN2(g5052), .QN(n14327) );
  NOR2X0 U14452 ( .IN1(n14328), .IN2(n14329), .QN(n14326) );
  NOR2X0 U14453 ( .IN1(n5615), .IN2(n14330), .QN(n14329) );
  NAND2X0 U14454 ( .IN1(n14331), .IN2(n14332), .QN(n14330) );
  INVX0 U14455 ( .INP(n14333), .ZN(n14332) );
  NOR2X0 U14456 ( .IN1(n14334), .IN2(g5057), .QN(n14328) );
  NOR2X0 U14457 ( .IN1(n14333), .IN2(n14335), .QN(n14334) );
  NOR2X0 U14458 ( .IN1(n14336), .IN2(n5607), .QN(n14333) );
  NAND2X0 U14459 ( .IN1(n14337), .IN2(n14338), .QN(g33045) );
  NAND2X0 U14460 ( .IN1(n13560), .IN2(g4567), .QN(n14338) );
  NOR2X0 U14461 ( .IN1(n14339), .IN2(n14340), .QN(n14337) );
  NAND2X0 U14462 ( .IN1(n14341), .IN2(n14342), .QN(g33044) );
  NAND2X0 U14463 ( .IN1(test_so93), .IN2(n13560), .QN(n14342) );
  NOR2X0 U14464 ( .IN1(n12764), .IN2(n14340), .QN(n14341) );
  NAND2X0 U14465 ( .IN1(n14343), .IN2(n14344), .QN(g33043) );
  NAND2X0 U14466 ( .IN1(test_so16), .IN2(n13560), .QN(n14344) );
  NOR2X0 U14467 ( .IN1(n14345), .IN2(n13561), .QN(n14343) );
  NAND2X0 U14468 ( .IN1(n14346), .IN2(n14347), .QN(g33042) );
  NAND2X0 U14469 ( .IN1(n13560), .IN2(g4540), .QN(n14347) );
  NOR2X0 U14470 ( .IN1(n14345), .IN2(n14340), .QN(n14346) );
  INVX0 U14471 ( .INP(n14348), .ZN(n14340) );
  NAND2X0 U14472 ( .IN1(n14349), .IN2(g4578), .QN(n14348) );
  NAND2X0 U14473 ( .IN1(n14350), .IN2(n14351), .QN(g33041) );
  NAND2X0 U14474 ( .IN1(test_so56), .IN2(n13560), .QN(n14351) );
  NOR2X0 U14475 ( .IN1(n14339), .IN2(n13561), .QN(n14350) );
  NAND2X0 U14476 ( .IN1(n14352), .IN2(n14353), .QN(g33040) );
  NAND2X0 U14477 ( .IN1(n13560), .IN2(g4504), .QN(n14353) );
  NOR2X0 U14478 ( .IN1(n12764), .IN2(n14354), .QN(n14352) );
  NOR2X0 U14479 ( .IN1(n13560), .IN2(n12754), .QN(n12764) );
  INVX0 U14480 ( .INP(n11908), .ZN(n12754) );
  NAND2X0 U14481 ( .IN1(n13377), .IN2(n13381), .QN(n11908) );
  INVX0 U14482 ( .INP(g72), .ZN(n13381) );
  INVX0 U14483 ( .INP(g73), .ZN(n13377) );
  NAND2X0 U14484 ( .IN1(n14355), .IN2(n14356), .QN(g33039) );
  NAND2X0 U14485 ( .IN1(n13560), .IN2(g4501), .QN(n14356) );
  NOR2X0 U14486 ( .IN1(n14339), .IN2(n13564), .QN(n14355) );
  NAND2X0 U14487 ( .IN1(n14357), .IN2(n14358), .QN(g33038) );
  NAND2X0 U14488 ( .IN1(n13560), .IN2(g4498), .QN(n14358) );
  NOR2X0 U14489 ( .IN1(n14339), .IN2(n14354), .QN(n14357) );
  NOR2X0 U14490 ( .IN1(n13560), .IN2(n14359), .QN(n14339) );
  NOR2X0 U14491 ( .IN1(n13382), .IN2(g73), .QN(n14359) );
  INVX0 U14492 ( .INP(g72), .ZN(n13382) );
  NAND2X0 U14493 ( .IN1(n14360), .IN2(n14361), .QN(g33037) );
  NAND2X0 U14494 ( .IN1(n13560), .IN2(g4495), .QN(n14361) );
  NOR2X0 U14495 ( .IN1(n14345), .IN2(n13564), .QN(n14360) );
  NAND2X0 U14496 ( .IN1(n14362), .IN2(n14363), .QN(g33036) );
  NAND2X0 U14497 ( .IN1(n13560), .IN2(g4480), .QN(n14363) );
  NOR2X0 U14498 ( .IN1(n14345), .IN2(n14354), .QN(n14362) );
  NOR2X0 U14499 ( .IN1(n13560), .IN2(n10182), .QN(n14354) );
  NOR2X0 U14500 ( .IN1(n13560), .IN2(n14364), .QN(n14345) );
  NOR2X0 U14501 ( .IN1(n11433), .IN2(g72), .QN(n14364) );
  INVX0 U14502 ( .INP(g73), .ZN(n11433) );
  INVX0 U14503 ( .INP(n14349), .ZN(n13560) );
  NAND2X0 U14504 ( .IN1(n14365), .IN2(n14366), .QN(g33035) );
  NOR2X0 U14505 ( .IN1(n14367), .IN2(n14368), .QN(n14366) );
  NOR2X0 U14506 ( .IN1(n5350), .IN2(n10846), .QN(n14368) );
  NOR2X0 U14507 ( .IN1(n11055), .IN2(n14369), .QN(n14367) );
  NAND2X0 U14508 ( .IN1(n13571), .IN2(g4108), .QN(n14369) );
  NOR2X0 U14509 ( .IN1(n10631), .IN2(n14370), .QN(n14365) );
  NOR2X0 U14510 ( .IN1(g4108), .IN2(n13571), .QN(n14370) );
  NAND2X0 U14511 ( .IN1(n14371), .IN2(g4098), .QN(n13571) );
  NAND2X0 U14512 ( .IN1(n14372), .IN2(n14373), .QN(g33034) );
  NAND2X0 U14513 ( .IN1(n14374), .IN2(n14375), .QN(n14373) );
  NAND2X0 U14514 ( .IN1(n14376), .IN2(n14377), .QN(n14374) );
  NAND2X0 U14515 ( .IN1(n10927), .IN2(n14378), .QN(n14377) );
  NOR2X0 U14516 ( .IN1(n14379), .IN2(n14380), .QN(n14376) );
  NOR2X0 U14517 ( .IN1(test_so33), .IN2(n14381), .QN(n14380) );
  INVX0 U14518 ( .INP(g25676), .ZN(n14381) );
  NAND2X0 U14519 ( .IN1(n11079), .IN2(g3873), .QN(n14372) );
  NAND2X0 U14520 ( .IN1(n14382), .IN2(n14383), .QN(g33033) );
  NAND2X0 U14521 ( .IN1(test_so33), .IN2(n14384), .QN(n14383) );
  NAND2X0 U14522 ( .IN1(n14385), .IN2(n10956), .QN(n14384) );
  NAND2X0 U14523 ( .IN1(n5387), .IN2(n14375), .QN(n14385) );
  NAND2X0 U14524 ( .IN1(n14386), .IN2(g3873), .QN(n14382) );
  INVX0 U14525 ( .INP(n14387), .ZN(n14386) );
  NAND2X0 U14526 ( .IN1(n14388), .IN2(n14389), .QN(g33032) );
  NAND2X0 U14527 ( .IN1(n14390), .IN2(n14375), .QN(n14389) );
  NOR2X0 U14528 ( .IN1(test_so33), .IN2(n3479), .QN(n14390) );
  NAND2X0 U14529 ( .IN1(n11080), .IN2(g3863), .QN(n14388) );
  NAND2X0 U14530 ( .IN1(n14391), .IN2(n14392), .QN(g33031) );
  NAND2X0 U14531 ( .IN1(n14393), .IN2(n14375), .QN(n14392) );
  NAND2X0 U14532 ( .IN1(n3482), .IN2(n14394), .QN(n14393) );
  NAND2X0 U14533 ( .IN1(n10926), .IN2(n14395), .QN(n14394) );
  NAND2X0 U14534 ( .IN1(n11079), .IN2(g3857), .QN(n14391) );
  NAND2X0 U14535 ( .IN1(n14396), .IN2(n14397), .QN(g33029) );
  NAND2X0 U14536 ( .IN1(n14398), .IN2(n14399), .QN(n14397) );
  NAND2X0 U14537 ( .IN1(n14400), .IN2(n14401), .QN(n14398) );
  NAND2X0 U14538 ( .IN1(n10926), .IN2(n14402), .QN(n14401) );
  NOR2X0 U14539 ( .IN1(n14403), .IN2(n14404), .QN(n14400) );
  INVX0 U14540 ( .INP(n14405), .ZN(n14404) );
  NAND2X0 U14541 ( .IN1(n5645), .IN2(g25662), .QN(n14405) );
  NAND2X0 U14542 ( .IN1(n11079), .IN2(g3522), .QN(n14396) );
  NAND2X0 U14543 ( .IN1(n14406), .IN2(n14407), .QN(g33028) );
  NAND2X0 U14544 ( .IN1(n14408), .IN2(g3518), .QN(n14407) );
  NAND2X0 U14545 ( .IN1(n14409), .IN2(n10956), .QN(n14408) );
  NAND2X0 U14546 ( .IN1(n5383), .IN2(n14399), .QN(n14409) );
  NAND2X0 U14547 ( .IN1(n14410), .IN2(g3522), .QN(n14406) );
  INVX0 U14548 ( .INP(n14411), .ZN(n14410) );
  NAND2X0 U14549 ( .IN1(n14412), .IN2(n14413), .QN(g33027) );
  NAND2X0 U14550 ( .IN1(n14414), .IN2(n5645), .QN(n14413) );
  NOR2X0 U14551 ( .IN1(n3489), .IN2(n14415), .QN(n14414) );
  NAND2X0 U14552 ( .IN1(n11079), .IN2(g3512), .QN(n14412) );
  NAND2X0 U14553 ( .IN1(n14416), .IN2(n14417), .QN(g33026) );
  NAND2X0 U14554 ( .IN1(n14418), .IN2(n14399), .QN(n14417) );
  NAND2X0 U14555 ( .IN1(n3492), .IN2(n14419), .QN(n14418) );
  NAND2X0 U14556 ( .IN1(n10926), .IN2(n14420), .QN(n14419) );
  NAND2X0 U14557 ( .IN1(n11079), .IN2(g3506), .QN(n14416) );
  NAND2X0 U14558 ( .IN1(n14421), .IN2(n14422), .QN(g33024) );
  NAND2X0 U14559 ( .IN1(n11078), .IN2(g3171), .QN(n14422) );
  NOR2X0 U14560 ( .IN1(n14423), .IN2(n14424), .QN(n14421) );
  NOR2X0 U14561 ( .IN1(n14425), .IN2(n14426), .QN(n14424) );
  INVX0 U14562 ( .INP(g25648), .ZN(n14426) );
  NOR2X0 U14563 ( .IN1(n14427), .IN2(n14428), .QN(n14423) );
  NOR2X0 U14564 ( .IN1(n14429), .IN2(n14430), .QN(n14427) );
  NAND2X0 U14565 ( .IN1(n14431), .IN2(n14432), .QN(g33023) );
  NAND2X0 U14566 ( .IN1(n14433), .IN2(n14434), .QN(n14432) );
  NOR2X0 U14567 ( .IN1(n5603), .IN2(n11021), .QN(n14433) );
  NAND2X0 U14568 ( .IN1(n14435), .IN2(g3167), .QN(n14431) );
  NAND2X0 U14569 ( .IN1(n14436), .IN2(n10956), .QN(n14435) );
  NAND2X0 U14570 ( .IN1(n5603), .IN2(n14437), .QN(n14436) );
  NAND2X0 U14571 ( .IN1(n14438), .IN2(n14439), .QN(g33022) );
  NAND2X0 U14572 ( .IN1(n14434), .IN2(n14440), .QN(n14439) );
  INVX0 U14573 ( .INP(n14425), .ZN(n14434) );
  NAND2X0 U14574 ( .IN1(n11079), .IN2(g3161), .QN(n14438) );
  NAND2X0 U14575 ( .IN1(n14441), .IN2(n14442), .QN(g33021) );
  NAND2X0 U14576 ( .IN1(n11079), .IN2(g3155), .QN(n14442) );
  NOR2X0 U14577 ( .IN1(n14443), .IN2(n14444), .QN(n14441) );
  NOR2X0 U14578 ( .IN1(n3502), .IN2(n14428), .QN(n14444) );
  NAND2X0 U14579 ( .IN1(n14437), .IN2(n10956), .QN(n14428) );
  INVX0 U14580 ( .INP(n14445), .ZN(n14443) );
  NAND2X0 U14581 ( .IN1(n14446), .IN2(n14437), .QN(n14445) );
  NAND2X0 U14582 ( .IN1(n14447), .IN2(n14448), .QN(g33019) );
  NOR2X0 U14583 ( .IN1(n14449), .IN2(n14450), .QN(n14447) );
  NOR2X0 U14584 ( .IN1(n11029), .IN2(n14451), .QN(n14450) );
  XOR2X1 U14585 ( .IN1(n2790), .IN2(n5300), .Q(n14451) );
  NOR2X0 U14586 ( .IN1(n5516), .IN2(n10846), .QN(n14449) );
  NAND2X0 U14587 ( .IN1(n14452), .IN2(n14453), .QN(g33018) );
  NOR2X0 U14588 ( .IN1(n14454), .IN2(n14455), .QN(n14453) );
  NOR2X0 U14589 ( .IN1(g2610), .IN2(n14456), .QN(n14455) );
  NAND2X0 U14590 ( .IN1(n14457), .IN2(n14458), .QN(n14456) );
  NOR2X0 U14591 ( .IN1(n5508), .IN2(n13657), .QN(n14458) );
  NOR2X0 U14592 ( .IN1(n11309), .IN2(n14459), .QN(n14457) );
  INVX0 U14593 ( .INP(n3511), .ZN(n14459) );
  NOR2X0 U14594 ( .IN1(n10529), .IN2(n10846), .QN(n14454) );
  NOR2X0 U14595 ( .IN1(n14460), .IN2(n14461), .QN(n14452) );
  NOR2X0 U14596 ( .IN1(n14462), .IN2(n10653), .QN(n14461) );
  NOR2X0 U14597 ( .IN1(n14463), .IN2(n14464), .QN(n14462) );
  NAND2X0 U14598 ( .IN1(n11304), .IN2(n14004), .QN(n14464) );
  NOR2X0 U14599 ( .IN1(n11029), .IN2(n12651), .QN(n14463) );
  NOR2X0 U14600 ( .IN1(n14465), .IN2(n14466), .QN(n14460) );
  NAND2X0 U14601 ( .IN1(n3512), .IN2(n14467), .QN(n14466) );
  INVX0 U14602 ( .INP(n3513), .ZN(n14467) );
  NAND2X0 U14603 ( .IN1(n3524), .IN2(n12651), .QN(n3513) );
  INVX0 U14604 ( .INP(n3006), .ZN(n12651) );
  NAND2X0 U14605 ( .IN1(n3525), .IN2(n3505), .QN(n3006) );
  NAND2X0 U14606 ( .IN1(n14468), .IN2(n10529), .QN(n3512) );
  NOR2X0 U14607 ( .IN1(n5508), .IN2(n10087), .QN(n14468) );
  NAND2X0 U14608 ( .IN1(n14469), .IN2(n14470), .QN(g33017) );
  NOR2X0 U14609 ( .IN1(n3519), .IN2(n14471), .QN(n14470) );
  NOR2X0 U14610 ( .IN1(n5508), .IN2(n11304), .QN(n14471) );
  NOR2X0 U14611 ( .IN1(n14472), .IN2(n14473), .QN(n14469) );
  NOR2X0 U14612 ( .IN1(n10903), .IN2(n10653), .QN(n14473) );
  NOR2X0 U14613 ( .IN1(n10529), .IN2(n14465), .QN(n14472) );
  NAND2X0 U14614 ( .IN1(n14474), .IN2(n14475), .QN(g33016) );
  INVX0 U14615 ( .INP(n3519), .ZN(n14475) );
  NOR2X0 U14616 ( .IN1(n14476), .IN2(n14477), .QN(n14474) );
  NOR2X0 U14617 ( .IN1(n5372), .IN2(n14478), .QN(n14477) );
  NOR2X0 U14618 ( .IN1(n10529), .IN2(n11304), .QN(n14476) );
  NAND2X0 U14619 ( .IN1(n14479), .IN2(n14480), .QN(g33015) );
  NOR2X0 U14620 ( .IN1(n3519), .IN2(n14481), .QN(n14480) );
  NOR2X0 U14621 ( .IN1(n14465), .IN2(n14482), .QN(n14481) );
  NAND2X0 U14622 ( .IN1(n5508), .IN2(n14483), .QN(n14482) );
  NOR2X0 U14623 ( .IN1(n14484), .IN2(n14485), .QN(n14479) );
  NOR2X0 U14624 ( .IN1(n10902), .IN2(n10679), .QN(n14485) );
  NOR2X0 U14625 ( .IN1(n5372), .IN2(n11304), .QN(n14484) );
  NAND2X0 U14626 ( .IN1(n14486), .IN2(n14487), .QN(g33014) );
  NOR2X0 U14627 ( .IN1(n14488), .IN2(n14489), .QN(n14487) );
  NOR2X0 U14628 ( .IN1(g2476), .IN2(n14490), .QN(n14489) );
  NAND2X0 U14629 ( .IN1(n14491), .IN2(n14492), .QN(n14490) );
  NOR2X0 U14630 ( .IN1(n5509), .IN2(n11246), .QN(n14492) );
  NOR2X0 U14631 ( .IN1(n13657), .IN2(n14493), .QN(n14491) );
  INVX0 U14632 ( .INP(n3530), .ZN(n14493) );
  NOR2X0 U14633 ( .IN1(n10530), .IN2(n10846), .QN(n14488) );
  NOR2X0 U14634 ( .IN1(n14494), .IN2(n14495), .QN(n14486) );
  NOR2X0 U14635 ( .IN1(n5405), .IN2(n14496), .QN(n14495) );
  NOR2X0 U14636 ( .IN1(n14497), .IN2(n14498), .QN(n14496) );
  NAND2X0 U14637 ( .IN1(n11241), .IN2(n14004), .QN(n14498) );
  NOR2X0 U14638 ( .IN1(n11029), .IN2(n12650), .QN(n14497) );
  NOR2X0 U14639 ( .IN1(n14499), .IN2(n14500), .QN(n14494) );
  NAND2X0 U14640 ( .IN1(n3531), .IN2(n14501), .QN(n14500) );
  INVX0 U14641 ( .INP(n3532), .ZN(n14501) );
  NAND2X0 U14642 ( .IN1(n3524), .IN2(n12650), .QN(n3532) );
  INVX0 U14643 ( .INP(n3007), .ZN(n12650) );
  NAND2X0 U14644 ( .IN1(n14502), .IN2(n3525), .QN(n3007) );
  NOR2X0 U14645 ( .IN1(n5516), .IN2(g2741), .QN(n14502) );
  NAND2X0 U14646 ( .IN1(n14503), .IN2(n10530), .QN(n3531) );
  NOR2X0 U14647 ( .IN1(n5509), .IN2(n10087), .QN(n14503) );
  NAND2X0 U14648 ( .IN1(n14504), .IN2(n14505), .QN(g33013) );
  NOR2X0 U14649 ( .IN1(n3538), .IN2(n14506), .QN(n14505) );
  NOR2X0 U14650 ( .IN1(n5509), .IN2(n11241), .QN(n14506) );
  NOR2X0 U14651 ( .IN1(n14507), .IN2(n14508), .QN(n14504) );
  NOR2X0 U14652 ( .IN1(n5405), .IN2(n10842), .QN(n14508) );
  NOR2X0 U14653 ( .IN1(n10530), .IN2(n14499), .QN(n14507) );
  NAND2X0 U14654 ( .IN1(n14509), .IN2(n14510), .QN(g33012) );
  INVX0 U14655 ( .INP(n3538), .ZN(n14510) );
  NOR2X0 U14656 ( .IN1(n14511), .IN2(n14512), .QN(n14509) );
  NOR2X0 U14657 ( .IN1(n5373), .IN2(n14513), .QN(n14512) );
  NOR2X0 U14658 ( .IN1(n10530), .IN2(n11241), .QN(n14511) );
  NAND2X0 U14659 ( .IN1(n14514), .IN2(n14515), .QN(g33011) );
  NOR2X0 U14660 ( .IN1(n3538), .IN2(n14516), .QN(n14515) );
  NOR2X0 U14661 ( .IN1(n14499), .IN2(n14517), .QN(n14516) );
  NAND2X0 U14662 ( .IN1(n5509), .IN2(n14518), .QN(n14517) );
  NOR2X0 U14663 ( .IN1(n14519), .IN2(n14520), .QN(n14514) );
  NOR2X0 U14664 ( .IN1(n5840), .IN2(n10842), .QN(n14520) );
  NOR2X0 U14665 ( .IN1(n5373), .IN2(n11241), .QN(n14519) );
  NAND2X0 U14666 ( .IN1(n14521), .IN2(n14522), .QN(g33010) );
  NOR2X0 U14667 ( .IN1(n14523), .IN2(n14524), .QN(n14522) );
  NOR2X0 U14668 ( .IN1(test_so21), .IN2(n14525), .QN(n14524) );
  NAND2X0 U14669 ( .IN1(n14526), .IN2(n14527), .QN(n14525) );
  NOR2X0 U14670 ( .IN1(n5511), .IN2(n11260), .QN(n14527) );
  NOR2X0 U14671 ( .IN1(n13657), .IN2(n14528), .QN(n14526) );
  INVX0 U14672 ( .INP(n3548), .ZN(n14528) );
  NOR2X0 U14673 ( .IN1(n10903), .IN2(n10640), .QN(n14523) );
  NOR2X0 U14674 ( .IN1(n14529), .IN2(n14530), .QN(n14521) );
  NOR2X0 U14675 ( .IN1(n5276), .IN2(n14531), .QN(n14530) );
  NOR2X0 U14676 ( .IN1(n14532), .IN2(n14533), .QN(n14531) );
  NAND2X0 U14677 ( .IN1(n11255), .IN2(n14004), .QN(n14533) );
  NOR2X0 U14678 ( .IN1(n11029), .IN2(n12649), .QN(n14532) );
  NOR2X0 U14679 ( .IN1(n14534), .IN2(n14535), .QN(n14529) );
  NAND2X0 U14680 ( .IN1(n3549), .IN2(n14536), .QN(n14535) );
  INVX0 U14681 ( .INP(n3551), .ZN(n14536) );
  NAND2X0 U14682 ( .IN1(n3524), .IN2(n12649), .QN(n3551) );
  INVX0 U14683 ( .INP(n3550), .ZN(n12649) );
  NAND2X0 U14684 ( .IN1(n14537), .IN2(n3525), .QN(n3550) );
  NOR2X0 U14685 ( .IN1(n5349), .IN2(g2748), .QN(n14537) );
  NAND2X0 U14686 ( .IN1(n14538), .IN2(g110), .QN(n3549) );
  NOR2X0 U14687 ( .IN1(test_so21), .IN2(n5511), .QN(n14538) );
  NAND2X0 U14688 ( .IN1(n14539), .IN2(n14540), .QN(g33009) );
  NOR2X0 U14689 ( .IN1(n3557), .IN2(n14541), .QN(n14540) );
  NOR2X0 U14690 ( .IN1(n5511), .IN2(n11255), .QN(n14541) );
  NOR2X0 U14691 ( .IN1(n14542), .IN2(n14543), .QN(n14539) );
  NOR2X0 U14692 ( .IN1(n5276), .IN2(n10842), .QN(n14543) );
  NOR2X0 U14693 ( .IN1(n10640), .IN2(n14534), .QN(n14542) );
  NAND2X0 U14694 ( .IN1(n14544), .IN2(n14545), .QN(g33008) );
  INVX0 U14695 ( .INP(n3557), .ZN(n14545) );
  NOR2X0 U14696 ( .IN1(n14546), .IN2(n14547), .QN(n14544) );
  NOR2X0 U14697 ( .IN1(n5375), .IN2(n14548), .QN(n14547) );
  NOR2X0 U14698 ( .IN1(n10640), .IN2(n11255), .QN(n14546) );
  NAND2X0 U14699 ( .IN1(n14549), .IN2(n14550), .QN(g33007) );
  NOR2X0 U14700 ( .IN1(n3557), .IN2(n14551), .QN(n14550) );
  NOR2X0 U14701 ( .IN1(n14534), .IN2(n14552), .QN(n14551) );
  NAND2X0 U14702 ( .IN1(n5511), .IN2(n14553), .QN(n14552) );
  NOR2X0 U14703 ( .IN1(n14554), .IN2(n14555), .QN(n14549) );
  NOR2X0 U14704 ( .IN1(n5841), .IN2(n10839), .QN(n14555) );
  NOR2X0 U14705 ( .IN1(n5375), .IN2(n11255), .QN(n14554) );
  NAND2X0 U14706 ( .IN1(n14556), .IN2(n14557), .QN(g33006) );
  NOR2X0 U14707 ( .IN1(n14558), .IN2(n14559), .QN(n14557) );
  NOR2X0 U14708 ( .IN1(g2208), .IN2(n14560), .QN(n14559) );
  NAND2X0 U14709 ( .IN1(n14561), .IN2(n14562), .QN(n14560) );
  NOR2X0 U14710 ( .IN1(n5512), .IN2(n13657), .QN(n14562) );
  NOR2X0 U14711 ( .IN1(n11495), .IN2(n14563), .QN(n14561) );
  INVX0 U14712 ( .INP(n3567), .ZN(n14563) );
  NOR2X0 U14713 ( .IN1(n10532), .IN2(n10839), .QN(n14558) );
  NOR2X0 U14714 ( .IN1(n14564), .IN2(n14565), .QN(n14556) );
  NOR2X0 U14715 ( .IN1(n5406), .IN2(n14566), .QN(n14565) );
  NOR2X0 U14716 ( .IN1(n14567), .IN2(n14568), .QN(n14566) );
  NAND2X0 U14717 ( .IN1(n11490), .IN2(n14004), .QN(n14568) );
  NOR2X0 U14718 ( .IN1(n11029), .IN2(n12648), .QN(n14567) );
  NOR2X0 U14719 ( .IN1(n14569), .IN2(n14570), .QN(n14564) );
  NAND2X0 U14720 ( .IN1(n3568), .IN2(n14571), .QN(n14570) );
  INVX0 U14721 ( .INP(n3570), .ZN(n14571) );
  NAND2X0 U14722 ( .IN1(n3524), .IN2(n12648), .QN(n3570) );
  INVX0 U14723 ( .INP(n3569), .ZN(n12648) );
  NAND2X0 U14724 ( .IN1(n14572), .IN2(n3525), .QN(n3569) );
  NOR2X0 U14725 ( .IN1(g2741), .IN2(g2748), .QN(n14572) );
  NAND2X0 U14726 ( .IN1(n14573), .IN2(n10532), .QN(n3568) );
  NOR2X0 U14727 ( .IN1(n5512), .IN2(n10087), .QN(n14573) );
  NAND2X0 U14728 ( .IN1(n14574), .IN2(n14575), .QN(g33005) );
  NOR2X0 U14729 ( .IN1(n3576), .IN2(n14576), .QN(n14575) );
  NOR2X0 U14730 ( .IN1(n5512), .IN2(n11490), .QN(n14576) );
  NOR2X0 U14731 ( .IN1(n14577), .IN2(n14578), .QN(n14574) );
  NOR2X0 U14732 ( .IN1(n5406), .IN2(n10849), .QN(n14578) );
  NOR2X0 U14733 ( .IN1(n10532), .IN2(n14569), .QN(n14577) );
  NAND2X0 U14734 ( .IN1(n14579), .IN2(n14580), .QN(g33004) );
  INVX0 U14735 ( .INP(n3576), .ZN(n14580) );
  NOR2X0 U14736 ( .IN1(n14581), .IN2(n14582), .QN(n14579) );
  NOR2X0 U14737 ( .IN1(n5376), .IN2(n14583), .QN(n14582) );
  NOR2X0 U14738 ( .IN1(n10532), .IN2(n11490), .QN(n14581) );
  NAND2X0 U14739 ( .IN1(n14584), .IN2(n14585), .QN(g33003) );
  NOR2X0 U14740 ( .IN1(n3576), .IN2(n14586), .QN(n14585) );
  NOR2X0 U14741 ( .IN1(n14569), .IN2(n14587), .QN(n14586) );
  NAND2X0 U14742 ( .IN1(n5512), .IN2(n14588), .QN(n14587) );
  NOR2X0 U14743 ( .IN1(n14589), .IN2(n14590), .QN(n14584) );
  NOR2X0 U14744 ( .IN1(n5839), .IN2(n10882), .QN(n14590) );
  NOR2X0 U14745 ( .IN1(n5376), .IN2(n11490), .QN(n14589) );
  NAND2X0 U14746 ( .IN1(n14591), .IN2(n14592), .QN(g33002) );
  NOR2X0 U14747 ( .IN1(n14593), .IN2(n14594), .QN(n14592) );
  NOR2X0 U14748 ( .IN1(g2051), .IN2(n14595), .QN(n14594) );
  NAND2X0 U14749 ( .IN1(n14596), .IN2(n14597), .QN(n14595) );
  NOR2X0 U14750 ( .IN1(n5507), .IN2(n13657), .QN(n14597) );
  NOR2X0 U14751 ( .IN1(n14598), .IN2(n14599), .QN(n14596) );
  INVX0 U14752 ( .INP(n3586), .ZN(n14599) );
  NOR2X0 U14753 ( .IN1(n10528), .IN2(n10879), .QN(n14593) );
  NOR2X0 U14754 ( .IN1(n14600), .IN2(n14601), .QN(n14591) );
  NOR2X0 U14755 ( .IN1(n5832), .IN2(n14602), .QN(n14601) );
  NOR2X0 U14756 ( .IN1(n14603), .IN2(n14604), .QN(n14602) );
  NAND2X0 U14757 ( .IN1(n14605), .IN2(n14004), .QN(n14604) );
  NOR2X0 U14758 ( .IN1(n11029), .IN2(n12656), .QN(n14603) );
  NOR2X0 U14759 ( .IN1(n14606), .IN2(n14607), .QN(n14600) );
  NAND2X0 U14760 ( .IN1(n3587), .IN2(n14608), .QN(n14607) );
  INVX0 U14761 ( .INP(n3589), .ZN(n14608) );
  NAND2X0 U14762 ( .IN1(n3524), .IN2(n12656), .QN(n3589) );
  INVX0 U14763 ( .INP(n3588), .ZN(n12656) );
  NAND2X0 U14764 ( .IN1(n14609), .IN2(n3505), .QN(n3588) );
  NOR2X0 U14765 ( .IN1(test_so30), .IN2(n14610), .QN(n14609) );
  NAND2X0 U14766 ( .IN1(n14611), .IN2(n10528), .QN(n3587) );
  NOR2X0 U14767 ( .IN1(n5507), .IN2(n10087), .QN(n14611) );
  NAND2X0 U14768 ( .IN1(n14612), .IN2(n14613), .QN(g33001) );
  NOR2X0 U14769 ( .IN1(n3595), .IN2(n14614), .QN(n14613) );
  NOR2X0 U14770 ( .IN1(n5507), .IN2(n14605), .QN(n14614) );
  NOR2X0 U14771 ( .IN1(n14615), .IN2(n14616), .QN(n14612) );
  NOR2X0 U14772 ( .IN1(n5832), .IN2(n10879), .QN(n14616) );
  NOR2X0 U14773 ( .IN1(n10528), .IN2(n14606), .QN(n14615) );
  NAND2X0 U14774 ( .IN1(n14617), .IN2(n14618), .QN(g33000) );
  INVX0 U14775 ( .INP(n3595), .ZN(n14618) );
  NOR2X0 U14776 ( .IN1(n14619), .IN2(n14620), .QN(n14617) );
  NOR2X0 U14777 ( .IN1(n5371), .IN2(n14621), .QN(n14620) );
  NOR2X0 U14778 ( .IN1(n10528), .IN2(n14605), .QN(n14619) );
  NAND2X0 U14779 ( .IN1(n14622), .IN2(n14623), .QN(g32999) );
  NOR2X0 U14780 ( .IN1(n3595), .IN2(n14624), .QN(n14623) );
  NOR2X0 U14781 ( .IN1(n14606), .IN2(n14625), .QN(n14624) );
  NAND2X0 U14782 ( .IN1(n5507), .IN2(n14626), .QN(n14625) );
  NOR2X0 U14783 ( .IN1(n14627), .IN2(n14628), .QN(n14622) );
  NOR2X0 U14784 ( .IN1(n10904), .IN2(n10680), .QN(n14628) );
  NOR2X0 U14785 ( .IN1(n5371), .IN2(n14605), .QN(n14627) );
  NAND2X0 U14786 ( .IN1(n14629), .IN2(n14630), .QN(g32998) );
  NOR2X0 U14787 ( .IN1(n14631), .IN2(n14632), .QN(n14630) );
  NOR2X0 U14788 ( .IN1(g1917), .IN2(n14633), .QN(n14632) );
  NAND2X0 U14789 ( .IN1(n14634), .IN2(n14635), .QN(n14633) );
  NOR2X0 U14790 ( .IN1(n5510), .IN2(n13657), .QN(n14635) );
  NOR2X0 U14791 ( .IN1(n11319), .IN2(n14636), .QN(n14634) );
  INVX0 U14792 ( .INP(n3604), .ZN(n14636) );
  NOR2X0 U14793 ( .IN1(n10531), .IN2(n10878), .QN(n14631) );
  NOR2X0 U14794 ( .IN1(n14637), .IN2(n14638), .QN(n14629) );
  NOR2X0 U14795 ( .IN1(n5829), .IN2(n14639), .QN(n14638) );
  NOR2X0 U14796 ( .IN1(n14640), .IN2(n14641), .QN(n14639) );
  NAND2X0 U14797 ( .IN1(n11314), .IN2(n14004), .QN(n14641) );
  NOR2X0 U14798 ( .IN1(n11029), .IN2(n12655), .QN(n14640) );
  NOR2X0 U14799 ( .IN1(n14642), .IN2(n14643), .QN(n14637) );
  NAND2X0 U14800 ( .IN1(n3605), .IN2(n14644), .QN(n14643) );
  INVX0 U14801 ( .INP(n3607), .ZN(n14644) );
  NAND2X0 U14802 ( .IN1(n3524), .IN2(n12655), .QN(n3607) );
  INVX0 U14803 ( .INP(n3606), .ZN(n12655) );
  NAND2X0 U14804 ( .IN1(n14645), .IN2(n14646), .QN(n3606) );
  NOR2X0 U14805 ( .IN1(test_so30), .IN2(n5516), .QN(n14646) );
  NOR2X0 U14806 ( .IN1(g2741), .IN2(n14610), .QN(n14645) );
  NAND2X0 U14807 ( .IN1(n14647), .IN2(n10531), .QN(n3605) );
  NOR2X0 U14808 ( .IN1(n5510), .IN2(n10087), .QN(n14647) );
  NAND2X0 U14809 ( .IN1(n14648), .IN2(n14649), .QN(g32997) );
  NOR2X0 U14810 ( .IN1(n3613), .IN2(n14650), .QN(n14649) );
  NOR2X0 U14811 ( .IN1(n5510), .IN2(n11314), .QN(n14650) );
  NOR2X0 U14812 ( .IN1(n14651), .IN2(n14652), .QN(n14648) );
  NOR2X0 U14813 ( .IN1(n5829), .IN2(n10878), .QN(n14652) );
  NOR2X0 U14814 ( .IN1(n10531), .IN2(n14642), .QN(n14651) );
  NAND2X0 U14815 ( .IN1(n14653), .IN2(n14654), .QN(g32996) );
  INVX0 U14816 ( .INP(n3613), .ZN(n14654) );
  NOR2X0 U14817 ( .IN1(n14655), .IN2(n14656), .QN(n14653) );
  NOR2X0 U14818 ( .IN1(n5374), .IN2(n14657), .QN(n14656) );
  NOR2X0 U14819 ( .IN1(n10531), .IN2(n11314), .QN(n14655) );
  NAND2X0 U14820 ( .IN1(n14658), .IN2(n14659), .QN(g32995) );
  NOR2X0 U14821 ( .IN1(n3613), .IN2(n14660), .QN(n14659) );
  NOR2X0 U14822 ( .IN1(n14642), .IN2(n14661), .QN(n14660) );
  NAND2X0 U14823 ( .IN1(n5510), .IN2(n14662), .QN(n14661) );
  NOR2X0 U14824 ( .IN1(n14663), .IN2(n14664), .QN(n14658) );
  NOR2X0 U14825 ( .IN1(n5837), .IN2(n10878), .QN(n14664) );
  NOR2X0 U14826 ( .IN1(n5374), .IN2(n11314), .QN(n14663) );
  NAND2X0 U14827 ( .IN1(n14665), .IN2(n14666), .QN(g32994) );
  NOR2X0 U14828 ( .IN1(n14667), .IN2(n14668), .QN(n14666) );
  NOR2X0 U14829 ( .IN1(g1783), .IN2(n14669), .QN(n14668) );
  NAND2X0 U14830 ( .IN1(n14670), .IN2(n14671), .QN(n14669) );
  NOR2X0 U14831 ( .IN1(n5359), .IN2(n11230), .QN(n14671) );
  NOR2X0 U14832 ( .IN1(n13657), .IN2(n14672), .QN(n14670) );
  INVX0 U14833 ( .INP(n3622), .ZN(n14672) );
  NOR2X0 U14834 ( .IN1(n5596), .IN2(n10878), .QN(n14667) );
  NOR2X0 U14835 ( .IN1(n14673), .IN2(n14674), .QN(n14665) );
  NOR2X0 U14836 ( .IN1(n5833), .IN2(n14675), .QN(n14674) );
  NOR2X0 U14837 ( .IN1(n14676), .IN2(n14677), .QN(n14675) );
  NAND2X0 U14838 ( .IN1(n11225), .IN2(n14004), .QN(n14677) );
  NOR2X0 U14839 ( .IN1(n3005), .IN2(n11019), .QN(n14676) );
  NOR2X0 U14840 ( .IN1(n14678), .IN2(n14679), .QN(n14673) );
  NAND2X0 U14841 ( .IN1(n3623), .IN2(n14680), .QN(n14679) );
  INVX0 U14842 ( .INP(n3624), .ZN(n14680) );
  NAND2X0 U14843 ( .IN1(n3524), .IN2(n3005), .QN(n3624) );
  NAND2X0 U14844 ( .IN1(n14681), .IN2(n5596), .QN(n3623) );
  NOR2X0 U14845 ( .IN1(n5359), .IN2(n10087), .QN(n14681) );
  NAND2X0 U14846 ( .IN1(n14682), .IN2(n14683), .QN(g32993) );
  NOR2X0 U14847 ( .IN1(n3630), .IN2(n14684), .QN(n14683) );
  NOR2X0 U14848 ( .IN1(n5359), .IN2(n11225), .QN(n14684) );
  NOR2X0 U14849 ( .IN1(n14685), .IN2(n14686), .QN(n14682) );
  NOR2X0 U14850 ( .IN1(n5833), .IN2(n10878), .QN(n14686) );
  NOR2X0 U14851 ( .IN1(n5596), .IN2(n14678), .QN(n14685) );
  NAND2X0 U14852 ( .IN1(n14687), .IN2(n14688), .QN(g32992) );
  INVX0 U14853 ( .INP(n3630), .ZN(n14688) );
  NOR2X0 U14854 ( .IN1(n14689), .IN2(n14690), .QN(n14687) );
  NOR2X0 U14855 ( .IN1(n5602), .IN2(n14691), .QN(n14690) );
  NOR2X0 U14856 ( .IN1(n5596), .IN2(n11225), .QN(n14689) );
  NAND2X0 U14857 ( .IN1(n14692), .IN2(n14693), .QN(g32991) );
  NOR2X0 U14858 ( .IN1(n3630), .IN2(n14694), .QN(n14693) );
  NOR2X0 U14859 ( .IN1(n14678), .IN2(n14695), .QN(n14694) );
  NAND2X0 U14860 ( .IN1(n5359), .IN2(n14696), .QN(n14695) );
  NOR2X0 U14861 ( .IN1(n14697), .IN2(n14698), .QN(n14692) );
  NOR2X0 U14862 ( .IN1(n5834), .IN2(n10875), .QN(n14698) );
  NOR2X0 U14863 ( .IN1(n5602), .IN2(n11225), .QN(n14697) );
  NAND2X0 U14864 ( .IN1(n14699), .IN2(n14700), .QN(g32990) );
  NOR2X0 U14865 ( .IN1(n14701), .IN2(n14702), .QN(n14700) );
  NOR2X0 U14866 ( .IN1(test_so94), .IN2(n14703), .QN(n14702) );
  NAND2X0 U14867 ( .IN1(n14704), .IN2(n14705), .QN(n14703) );
  NOR2X0 U14868 ( .IN1(n5525), .IN2(n13657), .QN(n14705) );
  NOR2X0 U14869 ( .IN1(n11476), .IN2(n14706), .QN(n14704) );
  INVX0 U14870 ( .INP(n3640), .ZN(n14706) );
  NOR2X0 U14871 ( .IN1(n10902), .IN2(n10638), .QN(n14701) );
  NOR2X0 U14872 ( .IN1(n14707), .IN2(n14708), .QN(n14699) );
  NOR2X0 U14873 ( .IN1(n5407), .IN2(n14709), .QN(n14708) );
  NOR2X0 U14874 ( .IN1(n14710), .IN2(n14711), .QN(n14709) );
  NAND2X0 U14875 ( .IN1(n14004), .IN2(n11471), .QN(n14711) );
  NAND2X0 U14876 ( .IN1(n10920), .IN2(n1770), .QN(n14004) );
  INVX0 U14877 ( .INP(n2760), .ZN(n1770) );
  NOR2X0 U14878 ( .IN1(n11029), .IN2(n12654), .QN(n14710) );
  NOR2X0 U14879 ( .IN1(n14712), .IN2(n14713), .QN(n14707) );
  NAND2X0 U14880 ( .IN1(n3641), .IN2(n14714), .QN(n14713) );
  INVX0 U14881 ( .INP(n3642), .ZN(n14714) );
  NAND2X0 U14882 ( .IN1(n3524), .IN2(n12654), .QN(n3642) );
  INVX0 U14883 ( .INP(n831), .ZN(n12654) );
  NAND2X0 U14884 ( .IN1(n832), .IN2(n864), .QN(n831) );
  INVX0 U14885 ( .INP(n14610), .ZN(n864) );
  NAND2X0 U14886 ( .IN1(n14715), .IN2(n14716), .QN(n14610) );
  XOR2X1 U14887 ( .IN1(n10100), .IN2(g73), .Q(n14716) );
  XOR2X1 U14888 ( .IN1(g72), .IN2(n10096), .Q(n14715) );
  INVX0 U14889 ( .INP(n14717), .ZN(n832) );
  NAND2X0 U14890 ( .IN1(n14718), .IN2(g110), .QN(n3641) );
  NOR2X0 U14891 ( .IN1(test_so94), .IN2(n5525), .QN(n14718) );
  NAND2X0 U14892 ( .IN1(n14719), .IN2(n14720), .QN(g32989) );
  NOR2X0 U14893 ( .IN1(n3648), .IN2(n14721), .QN(n14720) );
  NOR2X0 U14894 ( .IN1(n5525), .IN2(n11471), .QN(n14721) );
  NOR2X0 U14895 ( .IN1(n14722), .IN2(n14723), .QN(n14719) );
  NOR2X0 U14896 ( .IN1(n5407), .IN2(n10874), .QN(n14723) );
  NOR2X0 U14897 ( .IN1(n10638), .IN2(n14712), .QN(n14722) );
  NAND2X0 U14898 ( .IN1(n14724), .IN2(n14725), .QN(g32988) );
  INVX0 U14899 ( .INP(n3648), .ZN(n14725) );
  NOR2X0 U14900 ( .IN1(n14726), .IN2(n14727), .QN(n14724) );
  NOR2X0 U14901 ( .IN1(n5370), .IN2(n14728), .QN(n14727) );
  NOR2X0 U14902 ( .IN1(n10638), .IN2(n11471), .QN(n14726) );
  NAND2X0 U14903 ( .IN1(n14729), .IN2(n14730), .QN(g32987) );
  NOR2X0 U14904 ( .IN1(n3648), .IN2(n14731), .QN(n14730) );
  NOR2X0 U14905 ( .IN1(n14712), .IN2(n14732), .QN(n14731) );
  NAND2X0 U14906 ( .IN1(n5525), .IN2(n14733), .QN(n14732) );
  NOR2X0 U14907 ( .IN1(n14734), .IN2(n14735), .QN(n14729) );
  NOR2X0 U14908 ( .IN1(n5836), .IN2(n10871), .QN(n14735) );
  NOR2X0 U14909 ( .IN1(n5370), .IN2(n11471), .QN(n14734) );
  NAND2X0 U14910 ( .IN1(n14736), .IN2(n14737), .QN(g32986) );
  NAND2X0 U14911 ( .IN1(n14738), .IN2(n14739), .QN(n14737) );
  NOR2X0 U14912 ( .IN1(g1373), .IN2(n14122), .QN(n14738) );
  NOR2X0 U14913 ( .IN1(n14740), .IN2(n14741), .QN(n14736) );
  NOR2X0 U14914 ( .IN1(n10229), .IN2(n10871), .QN(n14741) );
  NOR2X0 U14915 ( .IN1(n11030), .IN2(n14742), .QN(n14740) );
  NAND2X0 U14916 ( .IN1(n14122), .IN2(g1373), .QN(n14742) );
  NAND2X0 U14917 ( .IN1(n227), .IN2(n14743), .QN(n14122) );
  NAND2X0 U14918 ( .IN1(n10229), .IN2(n14121), .QN(n14743) );
  NOR2X0 U14919 ( .IN1(n5730), .IN2(n14744), .QN(g32985) );
  NOR2X0 U14920 ( .IN1(n11030), .IN2(n14745), .QN(n14744) );
  NOR2X0 U14921 ( .IN1(n14746), .IN2(n14131), .QN(n14745) );
  NAND2X0 U14922 ( .IN1(n3662), .IN2(g1270), .QN(n14131) );
  NAND2X0 U14923 ( .IN1(n14747), .IN2(n14748), .QN(g32984) );
  NAND2X0 U14924 ( .IN1(n11079), .IN2(g1263), .QN(n14748) );
  NOR2X0 U14925 ( .IN1(n14749), .IN2(n14750), .QN(n14747) );
  NOR2X0 U14926 ( .IN1(n14751), .IN2(g1270), .QN(n14750) );
  NOR2X0 U14927 ( .IN1(n5716), .IN2(n14752), .QN(n14749) );
  NAND2X0 U14928 ( .IN1(n14133), .IN2(n14751), .QN(n14752) );
  INVX0 U14929 ( .INP(n3662), .ZN(n14751) );
  NAND2X0 U14930 ( .IN1(n14753), .IN2(n14754), .QN(g32983) );
  NAND2X0 U14931 ( .IN1(n14755), .IN2(n14756), .QN(n14754) );
  NOR2X0 U14932 ( .IN1(g1030), .IN2(n14141), .QN(n14755) );
  NOR2X0 U14933 ( .IN1(n14757), .IN2(n14758), .QN(n14753) );
  NOR2X0 U14934 ( .IN1(n10230), .IN2(n10871), .QN(n14758) );
  NOR2X0 U14935 ( .IN1(n11030), .IN2(n14759), .QN(n14757) );
  NAND2X0 U14936 ( .IN1(n14141), .IN2(g1030), .QN(n14759) );
  NAND2X0 U14937 ( .IN1(n591), .IN2(n14760), .QN(n14141) );
  NAND2X0 U14938 ( .IN1(n10230), .IN2(n14140), .QN(n14760) );
  NOR2X0 U14939 ( .IN1(n5731), .IN2(n14761), .QN(g32982) );
  NOR2X0 U14940 ( .IN1(n11030), .IN2(n14762), .QN(n14761) );
  NOR2X0 U14941 ( .IN1(n12087), .IN2(n14150), .QN(n14762) );
  NAND2X0 U14942 ( .IN1(n3671), .IN2(g925), .QN(n14150) );
  NAND2X0 U14943 ( .IN1(n14763), .IN2(n14764), .QN(g32981) );
  NAND2X0 U14944 ( .IN1(n11078), .IN2(g918), .QN(n14764) );
  NOR2X0 U14945 ( .IN1(n14765), .IN2(n14766), .QN(n14763) );
  NOR2X0 U14946 ( .IN1(n14767), .IN2(g925), .QN(n14766) );
  NOR2X0 U14947 ( .IN1(n5725), .IN2(n14768), .QN(n14765) );
  NAND2X0 U14948 ( .IN1(n14152), .IN2(n14767), .QN(n14768) );
  INVX0 U14949 ( .INP(n3671), .ZN(n14767) );
  NOR2X0 U14950 ( .IN1(n11030), .IN2(n14769), .QN(g32980) );
  NOR2X0 U14951 ( .IN1(n14770), .IN2(n12408), .QN(n14769) );
  NOR2X0 U14952 ( .IN1(n14771), .IN2(n2644), .QN(n12408) );
  NOR2X0 U14953 ( .IN1(n5754), .IN2(n14772), .QN(n14770) );
  INVX0 U14954 ( .INP(n14771), .ZN(n14772) );
  NAND2X0 U14955 ( .IN1(n14773), .IN2(n14774), .QN(n14771) );
  NOR2X0 U14956 ( .IN1(n5633), .IN2(n10610), .QN(n14774) );
  NOR2X0 U14957 ( .IN1(n10280), .IN2(g385), .QN(n14773) );
  NAND2X0 U14958 ( .IN1(n14775), .IN2(n14776), .QN(g32979) );
  NAND2X0 U14959 ( .IN1(test_so2), .IN2(n11081), .QN(n14776) );
  NOR2X0 U14960 ( .IN1(n14777), .IN2(n14778), .QN(n14775) );
  NOR2X0 U14961 ( .IN1(g758), .IN2(n14779), .QN(n14778) );
  NOR2X0 U14962 ( .IN1(n5331), .IN2(n14780), .QN(n14777) );
  NAND2X0 U14963 ( .IN1(n2404), .IN2(n14779), .QN(n14780) );
  INVX0 U14964 ( .INP(n3272), .ZN(n14779) );
  NAND2X0 U14965 ( .IN1(n14781), .IN2(n14782), .QN(g32978) );
  NAND2X0 U14966 ( .IN1(n11079), .IN2(g582), .QN(n14782) );
  NOR2X0 U14967 ( .IN1(n14783), .IN2(n14784), .QN(n14781) );
  NOR2X0 U14968 ( .IN1(g590), .IN2(n14785), .QN(n14784) );
  NOR2X0 U14969 ( .IN1(n5472), .IN2(n14786), .QN(n14783) );
  NAND2X0 U14970 ( .IN1(n2421), .IN2(n14785), .QN(n14786) );
  INVX0 U14971 ( .INP(n3274), .ZN(n14785) );
  NAND2X0 U14972 ( .IN1(n14787), .IN2(n14788), .QN(g32977) );
  NAND2X0 U14973 ( .IN1(test_so51), .IN2(n11081), .QN(n14788) );
  NOR2X0 U14974 ( .IN1(n14789), .IN2(n14790), .QN(n14787) );
  NOR2X0 U14975 ( .IN1(g291), .IN2(n14791), .QN(n14790) );
  NOR2X0 U14976 ( .IN1(n5679), .IN2(n14792), .QN(n14789) );
  NAND2X0 U14977 ( .IN1(n95), .IN2(n14791), .QN(n14792) );
  INVX0 U14978 ( .INP(n97), .ZN(n14791) );
  NOR2X0 U14979 ( .IN1(n14793), .IN2(n10655), .QN(n97) );
  NAND2X0 U14980 ( .IN1(n14794), .IN2(test_so51), .QN(n14793) );
  INVX0 U14981 ( .INP(n14795), .ZN(n95) );
  NAND2X0 U14982 ( .IN1(n14796), .IN2(n14797), .QN(g32976) );
  NAND2X0 U14983 ( .IN1(n11078), .IN2(g164), .QN(n14797) );
  NOR2X0 U14984 ( .IN1(n14798), .IN2(n14799), .QN(n14796) );
  NOR2X0 U14985 ( .IN1(g150), .IN2(n14800), .QN(n14799) );
  NOR2X0 U14986 ( .IN1(n5676), .IN2(n14801), .QN(n14798) );
  NAND2X0 U14987 ( .IN1(n12641), .IN2(n14800), .QN(n14801) );
  INVX0 U14988 ( .INP(n3281), .ZN(n14800) );
  NOR2X0 U14989 ( .IN1(n14802), .IN2(n14803), .QN(g32185) );
  NAND2X0 U14990 ( .IN1(n14804), .IN2(n14805), .QN(n14803) );
  NAND2X0 U14991 ( .IN1(g2970), .IN2(g2975), .QN(n14805) );
  NOR2X0 U14992 ( .IN1(n14806), .IN2(n14807), .QN(n14804) );
  NOR2X0 U14993 ( .IN1(n10560), .IN2(n10232), .QN(n14807) );
  NOR2X0 U14994 ( .IN1(n10231), .IN2(n10660), .QN(n14806) );
  NAND2X0 U14995 ( .IN1(n14808), .IN2(n14809), .QN(n14802) );
  NOR2X0 U14996 ( .IN1(n14810), .IN2(n14811), .QN(n14809) );
  NOR2X0 U14997 ( .IN1(n10609), .IN2(n10559), .QN(n14811) );
  NOR2X0 U14998 ( .IN1(n10617), .IN2(n10558), .QN(n14810) );
  NOR2X0 U14999 ( .IN1(n14812), .IN2(n14813), .QN(n14808) );
  NOR2X0 U15000 ( .IN1(n10615), .IN2(n10675), .QN(n14813) );
  NOR2X0 U15001 ( .IN1(n10562), .IN2(n10561), .QN(n14812) );
  NAND2X0 U15002 ( .IN1(n14814), .IN2(n14815), .QN(g31904) );
  NOR2X0 U15003 ( .IN1(n14816), .IN2(n14817), .QN(n14815) );
  NOR2X0 U15004 ( .IN1(n14818), .IN2(g5033), .QN(n14817) );
  NOR2X0 U15005 ( .IN1(n10598), .IN2(n14819), .QN(n14816) );
  NAND2X0 U15006 ( .IN1(n14820), .IN2(n14331), .QN(n14819) );
  NOR2X0 U15007 ( .IN1(n14821), .IN2(n14822), .QN(n14820) );
  NOR2X0 U15008 ( .IN1(n14823), .IN2(n14824), .QN(n14814) );
  NOR2X0 U15009 ( .IN1(n5601), .IN2(n10871), .QN(n14823) );
  NAND2X0 U15010 ( .IN1(n14825), .IN2(n14826), .QN(g31903) );
  NOR2X0 U15011 ( .IN1(n14827), .IN2(n14828), .QN(n14826) );
  NOR2X0 U15012 ( .IN1(n14336), .IN2(g5052), .QN(n14828) );
  INVX0 U15013 ( .INP(n14829), .ZN(n14336) );
  NOR2X0 U15014 ( .IN1(n5607), .IN2(n14830), .QN(n14827) );
  NAND2X0 U15015 ( .IN1(n14831), .IN2(n14331), .QN(n14830) );
  NOR2X0 U15016 ( .IN1(n14832), .IN2(n14829), .QN(n14831) );
  NOR2X0 U15017 ( .IN1(n14833), .IN2(n5578), .QN(n14829) );
  NOR2X0 U15018 ( .IN1(n14335), .IN2(n14834), .QN(n14825) );
  NOR2X0 U15019 ( .IN1(n5578), .IN2(n10868), .QN(n14834) );
  NOR2X0 U15020 ( .IN1(n14835), .IN2(g5052), .QN(n14335) );
  NAND2X0 U15021 ( .IN1(n14836), .IN2(n14837), .QN(g31902) );
  NAND2X0 U15022 ( .IN1(n14822), .IN2(n10955), .QN(n14837) );
  NOR2X0 U15023 ( .IN1(n14838), .IN2(n14839), .QN(n14836) );
  NOR2X0 U15024 ( .IN1(n5369), .IN2(n14840), .QN(n14839) );
  NOR2X0 U15025 ( .IN1(n11031), .IN2(n14841), .QN(n14840) );
  NOR2X0 U15026 ( .IN1(n10253), .IN2(g5029), .QN(n14841) );
  NOR2X0 U15027 ( .IN1(n14842), .IN2(n14843), .QN(n14838) );
  NAND2X0 U15028 ( .IN1(n14331), .IN2(g5029), .QN(n14843) );
  NAND2X0 U15029 ( .IN1(n14844), .IN2(n14845), .QN(n14842) );
  NAND2X0 U15030 ( .IN1(g5062), .IN2(g5016), .QN(n14844) );
  NAND2X0 U15031 ( .IN1(n14846), .IN2(n14847), .QN(g31901) );
  NOR2X0 U15032 ( .IN1(n14848), .IN2(n14849), .QN(n14847) );
  NOR2X0 U15033 ( .IN1(g5046), .IN2(n14833), .QN(n14849) );
  NOR2X0 U15034 ( .IN1(n5578), .IN2(n14850), .QN(n14848) );
  NAND2X0 U15035 ( .IN1(n14851), .IN2(n14331), .QN(n14850) );
  INVX0 U15036 ( .INP(n14852), .ZN(n14851) );
  NAND2X0 U15037 ( .IN1(n14833), .IN2(n14853), .QN(n14852) );
  NAND2X0 U15038 ( .IN1(n14854), .IN2(g5041), .QN(n14833) );
  NOR2X0 U15039 ( .IN1(n14855), .IN2(n14856), .QN(n14846) );
  INVX0 U15040 ( .INP(n14835), .ZN(n14856) );
  NAND2X0 U15041 ( .IN1(n10922), .IN2(n14832), .QN(n14835) );
  NOR2X0 U15042 ( .IN1(n14853), .IN2(g5046), .QN(n14832) );
  NAND2X0 U15043 ( .IN1(n14857), .IN2(n5611), .QN(n14853) );
  NOR2X0 U15044 ( .IN1(n14858), .IN2(g5041), .QN(n14857) );
  NOR2X0 U15045 ( .IN1(n5605), .IN2(n10867), .QN(n14855) );
  NAND2X0 U15046 ( .IN1(n14859), .IN2(n14860), .QN(g31900) );
  NAND2X0 U15047 ( .IN1(n5605), .IN2(n14861), .QN(n14860) );
  NAND2X0 U15048 ( .IN1(n14862), .IN2(n14863), .QN(n14861) );
  INVX0 U15049 ( .INP(n14854), .ZN(n14862) );
  NOR2X0 U15050 ( .IN1(n14864), .IN2(n14865), .QN(n14859) );
  NOR2X0 U15051 ( .IN1(n5611), .IN2(n10867), .QN(n14865) );
  NOR2X0 U15052 ( .IN1(n11031), .IN2(n14866), .QN(n14864) );
  NAND2X0 U15053 ( .IN1(n14867), .IN2(n14868), .QN(n14866) );
  NOR2X0 U15054 ( .IN1(n5605), .IN2(n14854), .QN(n14868) );
  NOR2X0 U15055 ( .IN1(n14869), .IN2(n5611), .QN(n14854) );
  NOR2X0 U15056 ( .IN1(n14870), .IN2(n14871), .QN(n14867) );
  NOR2X0 U15057 ( .IN1(n14858), .IN2(g5037), .QN(n14870) );
  NAND2X0 U15058 ( .IN1(n14872), .IN2(n14873), .QN(g31899) );
  NOR2X0 U15059 ( .IN1(n14874), .IN2(n14875), .QN(n14873) );
  NOR2X0 U15060 ( .IN1(n14869), .IN2(g5037), .QN(n14875) );
  NOR2X0 U15061 ( .IN1(n5611), .IN2(n14876), .QN(n14874) );
  INVX0 U15062 ( .INP(n14877), .ZN(n14876) );
  NOR2X0 U15063 ( .IN1(n14878), .IN2(n14879), .QN(n14877) );
  NAND2X0 U15064 ( .IN1(n14869), .IN2(n14858), .QN(n14878) );
  NAND2X0 U15065 ( .IN1(n14821), .IN2(g5033), .QN(n14869) );
  INVX0 U15066 ( .INP(n14818), .ZN(n14821) );
  NAND2X0 U15067 ( .IN1(n14880), .IN2(g5062), .QN(n14818) );
  NOR2X0 U15068 ( .IN1(n5601), .IN2(n5369), .QN(n14880) );
  NOR2X0 U15069 ( .IN1(n14881), .IN2(n14882), .QN(n14872) );
  NOR2X0 U15070 ( .IN1(n10598), .IN2(n10864), .QN(n14882) );
  INVX0 U15071 ( .INP(n14863), .ZN(n14881) );
  NAND2X0 U15072 ( .IN1(n14824), .IN2(n5611), .QN(n14863) );
  NOR2X0 U15073 ( .IN1(n11031), .IN2(n14858), .QN(n14824) );
  NAND2X0 U15074 ( .IN1(n10598), .IN2(n14822), .QN(n14858) );
  NOR2X0 U15075 ( .IN1(n14845), .IN2(g5029), .QN(n14822) );
  NAND2X0 U15076 ( .IN1(n5369), .IN2(g5022), .QN(n14845) );
  NAND2X0 U15077 ( .IN1(n14883), .IN2(n14884), .QN(g31898) );
  NAND2X0 U15078 ( .IN1(n14885), .IN2(n5369), .QN(n14884) );
  NOR2X0 U15079 ( .IN1(n14886), .IN2(n14879), .QN(n14885) );
  INVX0 U15080 ( .INP(n14331), .ZN(n14879) );
  NOR2X0 U15081 ( .IN1(n14871), .IN2(n11017), .QN(n14331) );
  NAND2X0 U15082 ( .IN1(n14887), .IN2(n14888), .QN(n14871) );
  NOR2X0 U15083 ( .IN1(n14889), .IN2(n14890), .QN(n14883) );
  NOR2X0 U15084 ( .IN1(n10278), .IN2(n10864), .QN(n14890) );
  NOR2X0 U15085 ( .IN1(n11031), .IN2(n14891), .QN(n14889) );
  NAND2X0 U15086 ( .IN1(n14886), .IN2(g5016), .QN(n14891) );
  NOR2X0 U15087 ( .IN1(g5022), .IN2(g5062), .QN(n14886) );
  NAND2X0 U15088 ( .IN1(n14892), .IN2(n14893), .QN(g31897) );
  NOR2X0 U15089 ( .IN1(n13561), .IN2(n14894), .QN(n14892) );
  NOR2X0 U15090 ( .IN1(n10192), .IN2(n10864), .QN(n14894) );
  INVX0 U15091 ( .INP(n14895), .ZN(n13561) );
  NAND2X0 U15092 ( .IN1(n14349), .IN2(g4575), .QN(n14895) );
  NAND2X0 U15093 ( .IN1(n14896), .IN2(n14893), .QN(g31896) );
  INVX0 U15094 ( .INP(n14897), .ZN(n14893) );
  NAND2X0 U15095 ( .IN1(n14898), .IN2(n14899), .QN(n14897) );
  NAND2X0 U15096 ( .IN1(n14349), .IN2(n14900), .QN(n14899) );
  NAND2X0 U15097 ( .IN1(g72), .IN2(g73), .QN(n14900) );
  NAND2X0 U15098 ( .IN1(n14901), .IN2(g4372), .QN(n14898) );
  INVX0 U15099 ( .INP(n13567), .ZN(n14901) );
  NOR2X0 U15100 ( .IN1(n13564), .IN2(n14902), .QN(n14896) );
  NOR2X0 U15101 ( .IN1(n5849), .IN2(n10863), .QN(n14902) );
  INVX0 U15102 ( .INP(n14903), .ZN(n13564) );
  NAND2X0 U15103 ( .IN1(n14349), .IN2(test_so100), .QN(n14903) );
  NOR2X0 U15104 ( .IN1(n11031), .IN2(n5670), .QN(n14349) );
  NAND2X0 U15105 ( .IN1(n13657), .IN2(n14904), .QN(g31895) );
  NAND2X0 U15106 ( .IN1(n11079), .IN2(g4382), .QN(n14904) );
  NAND2X0 U15107 ( .IN1(n2760), .IN2(n10955), .QN(n13657) );
  NAND2X0 U15108 ( .IN1(n14905), .IN2(n14906), .QN(g31894) );
  NOR2X0 U15109 ( .IN1(n14907), .IN2(n14908), .QN(n14905) );
  NOR2X0 U15110 ( .IN1(n11031), .IN2(n14909), .QN(n14908) );
  XOR2X1 U15111 ( .IN1(n5350), .IN2(n14371), .Q(n14909) );
  NOR2X0 U15112 ( .IN1(n418), .IN2(n5340), .QN(n14371) );
  NAND2X0 U15113 ( .IN1(n14910), .IN2(g4087), .QN(n418) );
  NOR2X0 U15114 ( .IN1(n5340), .IN2(n10860), .QN(n14907) );
  NAND2X0 U15115 ( .IN1(n14911), .IN2(n14912), .QN(g31872) );
  NAND2X0 U15116 ( .IN1(n14913), .IN2(n3730), .QN(n14912) );
  XOR2X1 U15117 ( .IN1(g2748), .IN2(n14914), .Q(n14913) );
  NOR2X0 U15118 ( .IN1(n5349), .IN2(n3506), .QN(n14914) );
  NAND2X0 U15119 ( .IN1(n11078), .IN2(g2741), .QN(n14911) );
  NAND2X0 U15120 ( .IN1(n14915), .IN2(n14916), .QN(g31871) );
  NAND2X0 U15121 ( .IN1(n3733), .IN2(n14739), .QN(n14916) );
  NOR2X0 U15122 ( .IN1(n14917), .IN2(n14918), .QN(n14915) );
  NOR2X0 U15123 ( .IN1(n11032), .IN2(n14919), .QN(n14918) );
  INVX0 U15124 ( .INP(n14920), .ZN(n14919) );
  NOR2X0 U15125 ( .IN1(n227), .IN2(n10229), .QN(n14920) );
  NOR2X0 U15126 ( .IN1(n11421), .IN2(n14921), .QN(n227) );
  NOR2X0 U15127 ( .IN1(g1361), .IN2(n14126), .QN(n14921) );
  NOR2X0 U15128 ( .IN1(n10258), .IN2(n10871), .QN(n14917) );
  NAND2X0 U15129 ( .IN1(n14922), .IN2(n14923), .QN(g31870) );
  NAND2X0 U15130 ( .IN1(n11079), .IN2(g1259), .QN(n14923) );
  NOR2X0 U15131 ( .IN1(n14924), .IN2(n14925), .QN(n14922) );
  NOR2X0 U15132 ( .IN1(g1263), .IN2(n14926), .QN(n14925) );
  NOR2X0 U15133 ( .IN1(n5674), .IN2(n14927), .QN(n14924) );
  NAND2X0 U15134 ( .IN1(n14133), .IN2(n14926), .QN(n14927) );
  INVX0 U15135 ( .INP(n3664), .ZN(n14926) );
  NAND2X0 U15136 ( .IN1(n14928), .IN2(n14929), .QN(g31869) );
  NAND2X0 U15137 ( .IN1(n3738), .IN2(n14756), .QN(n14929) );
  NOR2X0 U15138 ( .IN1(n14930), .IN2(n14931), .QN(n14928) );
  NOR2X0 U15139 ( .IN1(n11032), .IN2(n14932), .QN(n14931) );
  INVX0 U15140 ( .INP(n14933), .ZN(n14932) );
  NOR2X0 U15141 ( .IN1(n591), .IN2(n10230), .QN(n14933) );
  NOR2X0 U15142 ( .IN1(n11420), .IN2(n14934), .QN(n591) );
  NOR2X0 U15143 ( .IN1(g1018), .IN2(n14145), .QN(n14934) );
  NOR2X0 U15144 ( .IN1(n10260), .IN2(n10857), .QN(n14930) );
  NAND2X0 U15145 ( .IN1(n14935), .IN2(n14936), .QN(g31868) );
  NAND2X0 U15146 ( .IN1(n11078), .IN2(g914), .QN(n14936) );
  NOR2X0 U15147 ( .IN1(n14937), .IN2(n14938), .QN(n14935) );
  NOR2X0 U15148 ( .IN1(g918), .IN2(n14939), .QN(n14938) );
  NOR2X0 U15149 ( .IN1(n5673), .IN2(n14940), .QN(n14937) );
  NAND2X0 U15150 ( .IN1(n14152), .IN2(n14939), .QN(n14940) );
  INVX0 U15151 ( .INP(n3673), .ZN(n14939) );
  NAND2X0 U15152 ( .IN1(n14941), .IN2(n14942), .QN(g31867) );
  NAND2X0 U15153 ( .IN1(n11079), .IN2(g744), .QN(n14942) );
  NOR2X0 U15154 ( .IN1(n14943), .IN2(n14944), .QN(n14941) );
  INVX0 U15155 ( .INP(n14945), .ZN(n14944) );
  NAND2X0 U15156 ( .IN1(n5471), .IN2(n3682), .QN(n14945) );
  NOR2X0 U15157 ( .IN1(n3682), .IN2(n14946), .QN(n14943) );
  NAND2X0 U15158 ( .IN1(n2404), .IN2(test_so2), .QN(n14946) );
  NAND2X0 U15159 ( .IN1(n14947), .IN2(n14948), .QN(g31866) );
  NAND2X0 U15160 ( .IN1(n11079), .IN2(g577), .QN(n14948) );
  NOR2X0 U15161 ( .IN1(n14949), .IN2(n14950), .QN(n14947) );
  NOR2X0 U15162 ( .IN1(g582), .IN2(n14951), .QN(n14950) );
  NOR2X0 U15163 ( .IN1(n5552), .IN2(n14952), .QN(n14949) );
  NAND2X0 U15164 ( .IN1(n2421), .IN2(n14951), .QN(n14952) );
  INVX0 U15165 ( .INP(n3684), .ZN(n14951) );
  NAND2X0 U15166 ( .IN1(n14953), .IN2(n14954), .QN(g31865) );
  NAND2X0 U15167 ( .IN1(test_so55), .IN2(n14955), .QN(n14954) );
  NAND2X0 U15168 ( .IN1(n14956), .IN2(n10945), .QN(n14955) );
  NAND2X0 U15169 ( .IN1(n14794), .IN2(n10668), .QN(n14956) );
  NAND2X0 U15170 ( .IN1(n14957), .IN2(n10655), .QN(n14953) );
  NOR2X0 U15171 ( .IN1(n10668), .IN2(n14795), .QN(n14957) );
  NAND2X0 U15172 ( .IN1(n14794), .IN2(n10965), .QN(n14795) );
  NOR2X0 U15173 ( .IN1(n14958), .IN2(n14959), .QN(n14794) );
  NAND2X0 U15174 ( .IN1(g691), .IN2(n14960), .QN(n14959) );
  NAND2X0 U15175 ( .IN1(n14961), .IN2(n14962), .QN(n14958) );
  NAND2X0 U15176 ( .IN1(g278), .IN2(n14963), .QN(n14962) );
  NAND2X0 U15177 ( .IN1(n14964), .IN2(n14965), .QN(g31864) );
  NAND2X0 U15178 ( .IN1(test_so73), .IN2(n11081), .QN(n14965) );
  NOR2X0 U15179 ( .IN1(n14966), .IN2(n14967), .QN(n14964) );
  NOR2X0 U15180 ( .IN1(g164), .IN2(n11506), .QN(n14967) );
  NOR2X0 U15181 ( .IN1(n5561), .IN2(n14968), .QN(n14966) );
  NAND2X0 U15182 ( .IN1(n12641), .IN2(n11506), .QN(n14968) );
  NAND2X0 U15183 ( .IN1(n14969), .IN2(test_so73), .QN(n11506) );
  NOR2X0 U15184 ( .IN1(n14970), .IN2(n14971), .QN(n14969) );
  NOR2X0 U15185 ( .IN1(g1636), .IN2(n5598), .QN(g31862) );
  NAND2X0 U15186 ( .IN1(n14972), .IN2(n14973), .QN(g31793) );
  NAND2X0 U15187 ( .IN1(n14974), .IN2(n12026), .QN(n14973) );
  NOR2X0 U15188 ( .IN1(n12027), .IN2(n14975), .QN(n14974) );
  NOR2X0 U15189 ( .IN1(n14976), .IN2(n14977), .QN(n14975) );
  INVX0 U15190 ( .INP(n12028), .ZN(n14977) );
  NOR2X0 U15191 ( .IN1(n12021), .IN2(n14978), .QN(n14976) );
  NOR2X0 U15192 ( .IN1(n14979), .IN2(n14980), .QN(n14978) );
  NOR2X0 U15193 ( .IN1(n14981), .IN2(n14982), .QN(n14980) );
  NOR2X0 U15194 ( .IN1(g4427), .IN2(n14983), .QN(n14979) );
  NAND2X0 U15195 ( .IN1(n14984), .IN2(n10695), .QN(n14983) );
  NAND2X0 U15196 ( .IN1(n14982), .IN2(n14985), .QN(n14984) );
  NAND2X0 U15197 ( .IN1(n14986), .IN2(n14987), .QN(n14985) );
  INVX0 U15198 ( .INP(n14981), .ZN(n14987) );
  NAND2X0 U15199 ( .IN1(n14988), .IN2(n14989), .QN(n14986) );
  NAND2X0 U15200 ( .IN1(n10153), .IN2(n14990), .QN(n14989) );
  NAND2X0 U15201 ( .IN1(g5471), .IN2(g5817), .QN(n14990) );
  NAND2X0 U15202 ( .IN1(n10139), .IN2(n10131), .QN(n14988) );
  NAND2X0 U15203 ( .IN1(n14991), .IN2(n14992), .QN(n14972) );
  NOR2X0 U15204 ( .IN1(n14993), .IN2(n14994), .QN(n14992) );
  NOR2X0 U15205 ( .IN1(n12026), .IN2(n14995), .QN(n14994) );
  INVX0 U15206 ( .INP(n12027), .ZN(n14995) );
  NOR2X0 U15207 ( .IN1(n14996), .IN2(n14997), .QN(n12026) );
  NOR2X0 U15208 ( .IN1(n11032), .IN2(n10149), .QN(n14996) );
  NOR2X0 U15209 ( .IN1(n10149), .IN2(n14998), .QN(n14993) );
  INVX0 U15210 ( .INP(n14997), .ZN(n14998) );
  NOR2X0 U15211 ( .IN1(n12028), .IN2(g6509), .QN(n14991) );
  NAND2X0 U15212 ( .IN1(n14999), .IN2(n15000), .QN(n12028) );
  NOR2X0 U15213 ( .IN1(n6007), .IN2(n14981), .QN(n15000) );
  NOR2X0 U15214 ( .IN1(n14982), .IN2(g4427), .QN(n14999) );
  INVX0 U15215 ( .INP(n15001), .ZN(n14982) );
  NAND2X0 U15216 ( .IN1(n15002), .IN2(n10955), .QN(n15001) );
  NAND2X0 U15217 ( .IN1(n15003), .IN2(n10153), .QN(n15002) );
  NOR2X0 U15218 ( .IN1(g5817), .IN2(g5471), .QN(n15003) );
  NAND2X0 U15219 ( .IN1(g113), .IN2(g2868), .QN(g31665) );
  NAND2X0 U15220 ( .IN1(g113), .IN2(g2873), .QN(g31656) );
  NAND2X0 U15221 ( .IN1(n15004), .IN2(n15005), .QN(g30563) );
  NAND2X0 U15222 ( .IN1(n11078), .IN2(g6653), .QN(n15005) );
  NOR2X0 U15223 ( .IN1(n15006), .IN2(n15007), .QN(n15004) );
  NOR2X0 U15224 ( .IN1(n13440), .IN2(n15008), .QN(n15007) );
  NOR2X0 U15225 ( .IN1(n10292), .IN2(n15009), .QN(n15006) );
  NAND2X0 U15226 ( .IN1(n15010), .IN2(n15011), .QN(g30562) );
  NAND2X0 U15227 ( .IN1(n15012), .IN2(n3765), .QN(n15011) );
  NOR2X0 U15228 ( .IN1(n15013), .IN2(n15014), .QN(n15010) );
  NOR2X0 U15229 ( .IN1(n10481), .IN2(n10861), .QN(n15014) );
  NOR2X0 U15230 ( .IN1(n11032), .IN2(n15015), .QN(n15013) );
  NAND2X0 U15231 ( .IN1(n15016), .IN2(g6605), .QN(n15015) );
  INVX0 U15232 ( .INP(n15012), .ZN(n15016) );
  NOR2X0 U15233 ( .IN1(n3768), .IN2(n5646), .QN(n15012) );
  NAND2X0 U15234 ( .IN1(n15017), .IN2(n15018), .QN(g30561) );
  NAND2X0 U15235 ( .IN1(n14208), .IN2(n3765), .QN(n15018) );
  NOR2X0 U15236 ( .IN1(n15019), .IN2(n15020), .QN(n15017) );
  NOR2X0 U15237 ( .IN1(n10368), .IN2(n10861), .QN(n15020) );
  NOR2X0 U15238 ( .IN1(n11032), .IN2(n15021), .QN(n15019) );
  INVX0 U15239 ( .INP(n15022), .ZN(n15021) );
  NOR2X0 U15240 ( .IN1(n14208), .IN2(n10483), .QN(n15022) );
  NOR2X0 U15241 ( .IN1(n3770), .IN2(n5646), .QN(n14208) );
  NAND2X0 U15242 ( .IN1(n15023), .IN2(n15024), .QN(g30560) );
  NAND2X0 U15243 ( .IN1(n15025), .IN2(n3765), .QN(n15024) );
  NOR2X0 U15244 ( .IN1(n15026), .IN2(n15027), .QN(n15023) );
  NOR2X0 U15245 ( .IN1(n10293), .IN2(n10861), .QN(n15027) );
  NOR2X0 U15246 ( .IN1(n11032), .IN2(n15028), .QN(n15026) );
  NAND2X0 U15247 ( .IN1(n15029), .IN2(g6589), .QN(n15028) );
  INVX0 U15248 ( .INP(n15025), .ZN(n15029) );
  NOR2X0 U15249 ( .IN1(n3773), .IN2(n5646), .QN(n15025) );
  NAND2X0 U15250 ( .IN1(n15030), .IN2(n15031), .QN(g30559) );
  NAND2X0 U15251 ( .IN1(n3774), .IN2(n15032), .QN(n15031) );
  NOR2X0 U15252 ( .IN1(n15033), .IN2(n15034), .QN(n15030) );
  NOR2X0 U15253 ( .IN1(n11032), .IN2(n15035), .QN(n15034) );
  NAND2X0 U15254 ( .IN1(n15036), .IN2(g6653), .QN(n15035) );
  NAND2X0 U15255 ( .IN1(n15037), .IN2(n15032), .QN(n15036) );
  NOR2X0 U15256 ( .IN1(n10349), .IN2(n10861), .QN(n15033) );
  NAND2X0 U15257 ( .IN1(n15038), .IN2(n15039), .QN(g30558) );
  NAND2X0 U15258 ( .IN1(n3774), .IN2(n14207), .QN(n15039) );
  NOR2X0 U15259 ( .IN1(n15040), .IN2(n15041), .QN(n15038) );
  NOR2X0 U15260 ( .IN1(n11032), .IN2(n15042), .QN(n15041) );
  NAND2X0 U15261 ( .IN1(n15043), .IN2(g6649), .QN(n15042) );
  NAND2X0 U15262 ( .IN1(n15037), .IN2(n14207), .QN(n15043) );
  NOR2X0 U15263 ( .IN1(n10479), .IN2(n10861), .QN(n15040) );
  NAND2X0 U15264 ( .IN1(n15044), .IN2(n15045), .QN(g30557) );
  NAND2X0 U15265 ( .IN1(n3774), .IN2(n15046), .QN(n15045) );
  NOR2X0 U15266 ( .IN1(n15047), .IN2(n15048), .QN(n15044) );
  NOR2X0 U15267 ( .IN1(n11033), .IN2(n15049), .QN(n15048) );
  NAND2X0 U15268 ( .IN1(n15050), .IN2(g6645), .QN(n15049) );
  NAND2X0 U15269 ( .IN1(n15037), .IN2(n15046), .QN(n15050) );
  NOR2X0 U15270 ( .IN1(n10382), .IN2(n10862), .QN(n15047) );
  NAND2X0 U15271 ( .IN1(n15051), .IN2(n15052), .QN(g30556) );
  NAND2X0 U15272 ( .IN1(n3774), .IN2(n15053), .QN(n15052) );
  NOR2X0 U15273 ( .IN1(n15054), .IN2(n15055), .QN(n15051) );
  NOR2X0 U15274 ( .IN1(n11025), .IN2(n15056), .QN(n15055) );
  NAND2X0 U15275 ( .IN1(n15057), .IN2(g6641), .QN(n15056) );
  NAND2X0 U15276 ( .IN1(n15037), .IN2(n15053), .QN(n15057) );
  INVX0 U15277 ( .INP(n3404), .ZN(n15037) );
  NAND2X0 U15278 ( .IN1(g6549), .IN2(g6555), .QN(n3404) );
  NOR2X0 U15279 ( .IN1(n10436), .IN2(n10862), .QN(n15054) );
  NAND2X0 U15280 ( .IN1(n15058), .IN2(n15059), .QN(g30555) );
  NAND2X0 U15281 ( .IN1(n3780), .IN2(n15032), .QN(n15059) );
  NOR2X0 U15282 ( .IN1(n15060), .IN2(n15061), .QN(n15058) );
  NOR2X0 U15283 ( .IN1(n11032), .IN2(n15062), .QN(n15061) );
  NAND2X0 U15284 ( .IN1(n15063), .IN2(g6637), .QN(n15062) );
  NAND2X0 U15285 ( .IN1(n14225), .IN2(n15032), .QN(n15063) );
  NOR2X0 U15286 ( .IN1(n10350), .IN2(n10862), .QN(n15060) );
  NAND2X0 U15287 ( .IN1(n15064), .IN2(n15065), .QN(g30554) );
  NAND2X0 U15288 ( .IN1(n3780), .IN2(n14207), .QN(n15065) );
  NOR2X0 U15289 ( .IN1(n15066), .IN2(n15067), .QN(n15064) );
  NOR2X0 U15290 ( .IN1(n11032), .IN2(n15068), .QN(n15067) );
  NAND2X0 U15291 ( .IN1(n15069), .IN2(g6633), .QN(n15068) );
  NAND2X0 U15292 ( .IN1(n14225), .IN2(n14207), .QN(n15069) );
  NOR2X0 U15293 ( .IN1(n10423), .IN2(n10862), .QN(n15066) );
  NAND2X0 U15294 ( .IN1(n15070), .IN2(n15071), .QN(g30553) );
  NAND2X0 U15295 ( .IN1(n3780), .IN2(n15046), .QN(n15071) );
  NOR2X0 U15296 ( .IN1(n15072), .IN2(n15073), .QN(n15070) );
  NOR2X0 U15297 ( .IN1(n11032), .IN2(n15074), .QN(n15073) );
  NAND2X0 U15298 ( .IN1(n15075), .IN2(g6629), .QN(n15074) );
  NAND2X0 U15299 ( .IN1(n14225), .IN2(n15046), .QN(n15075) );
  NOR2X0 U15300 ( .IN1(n10331), .IN2(n10862), .QN(n15072) );
  NAND2X0 U15301 ( .IN1(n15076), .IN2(n15077), .QN(g30552) );
  NAND2X0 U15302 ( .IN1(n3780), .IN2(n15053), .QN(n15077) );
  NOR2X0 U15303 ( .IN1(n15078), .IN2(n15079), .QN(n15076) );
  NOR2X0 U15304 ( .IN1(n11032), .IN2(n15080), .QN(n15079) );
  NAND2X0 U15305 ( .IN1(n15081), .IN2(g6625), .QN(n15080) );
  NAND2X0 U15306 ( .IN1(n14225), .IN2(n15053), .QN(n15081) );
  INVX0 U15307 ( .INP(n3406), .ZN(n14225) );
  NAND2X0 U15308 ( .IN1(n5571), .IN2(g6555), .QN(n3406) );
  NOR2X0 U15309 ( .IN1(n10294), .IN2(n10863), .QN(n15078) );
  NAND2X0 U15310 ( .IN1(n15082), .IN2(n15083), .QN(g30551) );
  NAND2X0 U15311 ( .IN1(n3785), .IN2(n15032), .QN(n15083) );
  NOR2X0 U15312 ( .IN1(n15084), .IN2(n15085), .QN(n15082) );
  NOR2X0 U15313 ( .IN1(n11032), .IN2(n15086), .QN(n15085) );
  NAND2X0 U15314 ( .IN1(n15087), .IN2(g6621), .QN(n15086) );
  NAND2X0 U15315 ( .IN1(n15088), .IN2(n15032), .QN(n15087) );
  NOR2X0 U15316 ( .IN1(n10424), .IN2(n10863), .QN(n15084) );
  NAND2X0 U15317 ( .IN1(n15089), .IN2(n15090), .QN(g30550) );
  NAND2X0 U15318 ( .IN1(n3785), .IN2(n14207), .QN(n15090) );
  NOR2X0 U15319 ( .IN1(n15091), .IN2(n15092), .QN(n15089) );
  NOR2X0 U15320 ( .IN1(n11031), .IN2(n15093), .QN(n15092) );
  NAND2X0 U15321 ( .IN1(n15094), .IN2(g6617), .QN(n15093) );
  NAND2X0 U15322 ( .IN1(n15088), .IN2(n14207), .QN(n15094) );
  INVX0 U15323 ( .INP(n3768), .ZN(n14207) );
  NAND2X0 U15324 ( .IN1(n5386), .IN2(g6573), .QN(n3768) );
  NOR2X0 U15325 ( .IN1(n10512), .IN2(n10863), .QN(n15091) );
  NAND2X0 U15326 ( .IN1(n15095), .IN2(n15096), .QN(g30549) );
  NAND2X0 U15327 ( .IN1(n3785), .IN2(n15046), .QN(n15096) );
  NOR2X0 U15328 ( .IN1(n15097), .IN2(n15098), .QN(n15095) );
  NOR2X0 U15329 ( .IN1(n11031), .IN2(n15099), .QN(n15098) );
  NAND2X0 U15330 ( .IN1(n15100), .IN2(g6613), .QN(n15099) );
  NAND2X0 U15331 ( .IN1(n15088), .IN2(n15046), .QN(n15100) );
  INVX0 U15332 ( .INP(n3770), .ZN(n15046) );
  NAND2X0 U15333 ( .IN1(n5563), .IN2(g6565), .QN(n3770) );
  NOR2X0 U15334 ( .IN1(n10904), .IN2(n10687), .QN(n15097) );
  NAND2X0 U15335 ( .IN1(n15101), .IN2(n15102), .QN(g30548) );
  NAND2X0 U15336 ( .IN1(n3785), .IN2(n15053), .QN(n15102) );
  NOR2X0 U15337 ( .IN1(n15103), .IN2(n15104), .QN(n15101) );
  NOR2X0 U15338 ( .IN1(n11031), .IN2(n15105), .QN(n15104) );
  NAND2X0 U15339 ( .IN1(n15106), .IN2(g6609), .QN(n15105) );
  NAND2X0 U15340 ( .IN1(n15088), .IN2(n15053), .QN(n15106) );
  INVX0 U15341 ( .INP(n3773), .ZN(n15053) );
  NAND2X0 U15342 ( .IN1(n5563), .IN2(n5386), .QN(n3773) );
  INVX0 U15343 ( .INP(n3407), .ZN(n15088) );
  NAND2X0 U15344 ( .IN1(n10592), .IN2(g6549), .QN(n3407) );
  NOR2X0 U15345 ( .IN1(n10450), .IN2(n10863), .QN(n15103) );
  NAND2X0 U15346 ( .IN1(n15107), .IN2(n15108), .QN(g30547) );
  NAND2X0 U15347 ( .IN1(n11079), .IN2(g6605), .QN(n15108) );
  NOR2X0 U15348 ( .IN1(n15109), .IN2(n15110), .QN(n15107) );
  NOR2X0 U15349 ( .IN1(n15008), .IN2(n15111), .QN(n15110) );
  INVX0 U15350 ( .INP(n3790), .ZN(n15111) );
  NOR2X0 U15351 ( .IN1(n3790), .IN2(n15112), .QN(n15109) );
  NAND2X0 U15352 ( .IN1(n10934), .IN2(g6601), .QN(n15112) );
  NAND2X0 U15353 ( .IN1(n15113), .IN2(n15114), .QN(g30546) );
  NAND2X0 U15354 ( .IN1(n11077), .IN2(g6597), .QN(n15114) );
  NOR2X0 U15355 ( .IN1(n15115), .IN2(n15116), .QN(n15113) );
  NOR2X0 U15356 ( .IN1(n15008), .IN2(n15117), .QN(n15116) );
  INVX0 U15357 ( .INP(n3793), .ZN(n15117) );
  NOR2X0 U15358 ( .IN1(n3793), .IN2(n15118), .QN(n15115) );
  NAND2X0 U15359 ( .IN1(n10935), .IN2(g6593), .QN(n15118) );
  NAND2X0 U15360 ( .IN1(n15119), .IN2(n15120), .QN(g30545) );
  NAND2X0 U15361 ( .IN1(n11078), .IN2(g6589), .QN(n15120) );
  NOR2X0 U15362 ( .IN1(n15121), .IN2(n15122), .QN(n15119) );
  NOR2X0 U15363 ( .IN1(n15008), .IN2(n15123), .QN(n15122) );
  INVX0 U15364 ( .INP(n3795), .ZN(n15123) );
  NOR2X0 U15365 ( .IN1(n3795), .IN2(n15124), .QN(n15121) );
  NAND2X0 U15366 ( .IN1(test_so71), .IN2(n10955), .QN(n15124) );
  NAND2X0 U15367 ( .IN1(n15125), .IN2(n15126), .QN(g30544) );
  NAND2X0 U15368 ( .IN1(n11078), .IN2(g6573), .QN(n15126) );
  NOR2X0 U15369 ( .IN1(n15127), .IN2(n15128), .QN(n15125) );
  NOR2X0 U15370 ( .IN1(n15008), .IN2(n15129), .QN(n15128) );
  INVX0 U15371 ( .INP(n3797), .ZN(n15129) );
  NOR2X0 U15372 ( .IN1(n3797), .IN2(n15130), .QN(n15127) );
  NAND2X0 U15373 ( .IN1(n10936), .IN2(g6581), .QN(n15130) );
  NOR2X0 U15374 ( .IN1(g6549), .IN2(n14216), .QN(g30543) );
  NAND2X0 U15375 ( .IN1(n15131), .IN2(n5646), .QN(n14216) );
  NOR2X0 U15376 ( .IN1(n11031), .IN2(n14220), .QN(n15131) );
  INVX0 U15377 ( .INP(n14204), .ZN(n14220) );
  NAND2X0 U15378 ( .IN1(n3799), .IN2(n15132), .QN(n14204) );
  NAND2X0 U15379 ( .IN1(n15133), .IN2(n15134), .QN(g30542) );
  NAND2X0 U15380 ( .IN1(n11078), .IN2(g6307), .QN(n15134) );
  NOR2X0 U15381 ( .IN1(n15135), .IN2(n15136), .QN(n15133) );
  NOR2X0 U15382 ( .IN1(n15008), .IN2(n13434), .QN(n15136) );
  NOR2X0 U15383 ( .IN1(n10299), .IN2(n15137), .QN(n15135) );
  NAND2X0 U15384 ( .IN1(n15138), .IN2(n15139), .QN(g30541) );
  NAND2X0 U15385 ( .IN1(n15140), .IN2(n3765), .QN(n15139) );
  NOR2X0 U15386 ( .IN1(n15141), .IN2(n15142), .QN(n15138) );
  NOR2X0 U15387 ( .IN1(n10491), .IN2(n10864), .QN(n15142) );
  NOR2X0 U15388 ( .IN1(n11031), .IN2(n15143), .QN(n15141) );
  NAND2X0 U15389 ( .IN1(n15144), .IN2(g6259), .QN(n15143) );
  INVX0 U15390 ( .INP(n15140), .ZN(n15144) );
  NOR2X0 U15391 ( .IN1(n3802), .IN2(n5651), .QN(n15140) );
  NAND2X0 U15392 ( .IN1(n15145), .IN2(n15146), .QN(g30540) );
  NAND2X0 U15393 ( .IN1(n14233), .IN2(n3765), .QN(n15146) );
  NOR2X0 U15394 ( .IN1(n15147), .IN2(n15148), .QN(n15145) );
  NOR2X0 U15395 ( .IN1(n10371), .IN2(n10864), .QN(n15148) );
  NOR2X0 U15396 ( .IN1(n11031), .IN2(n15149), .QN(n15147) );
  INVX0 U15397 ( .INP(n15150), .ZN(n15149) );
  NOR2X0 U15398 ( .IN1(n14233), .IN2(n10493), .QN(n15150) );
  NOR2X0 U15399 ( .IN1(n3804), .IN2(n5651), .QN(n14233) );
  NAND2X0 U15400 ( .IN1(n15151), .IN2(n15152), .QN(g30539) );
  NAND2X0 U15401 ( .IN1(n15153), .IN2(n3765), .QN(n15152) );
  NOR2X0 U15402 ( .IN1(n15154), .IN2(n15155), .QN(n15151) );
  NOR2X0 U15403 ( .IN1(n10300), .IN2(n10865), .QN(n15155) );
  NOR2X0 U15404 ( .IN1(n11031), .IN2(n15156), .QN(n15154) );
  NAND2X0 U15405 ( .IN1(n15157), .IN2(g6243), .QN(n15156) );
  INVX0 U15406 ( .INP(n15153), .ZN(n15157) );
  NOR2X0 U15407 ( .IN1(n3807), .IN2(n5651), .QN(n15153) );
  NAND2X0 U15408 ( .IN1(n15158), .IN2(n15159), .QN(g30538) );
  NAND2X0 U15409 ( .IN1(n3808), .IN2(n15160), .QN(n15159) );
  NOR2X0 U15410 ( .IN1(n15161), .IN2(n15162), .QN(n15158) );
  NOR2X0 U15411 ( .IN1(n11030), .IN2(n15163), .QN(n15162) );
  NAND2X0 U15412 ( .IN1(n15164), .IN2(g6307), .QN(n15163) );
  NAND2X0 U15413 ( .IN1(n15165), .IN2(n15160), .QN(n15164) );
  NOR2X0 U15414 ( .IN1(n10355), .IN2(n10865), .QN(n15161) );
  NAND2X0 U15415 ( .IN1(n15166), .IN2(n15167), .QN(g30537) );
  NAND2X0 U15416 ( .IN1(n3808), .IN2(n14232), .QN(n15167) );
  NOR2X0 U15417 ( .IN1(n15168), .IN2(n15169), .QN(n15166) );
  NOR2X0 U15418 ( .IN1(n11030), .IN2(n15170), .QN(n15169) );
  NAND2X0 U15419 ( .IN1(n15171), .IN2(g6303), .QN(n15170) );
  NAND2X0 U15420 ( .IN1(n15165), .IN2(n14232), .QN(n15171) );
  NOR2X0 U15421 ( .IN1(n10489), .IN2(n10865), .QN(n15168) );
  NAND2X0 U15422 ( .IN1(n15172), .IN2(n15173), .QN(g30536) );
  NAND2X0 U15423 ( .IN1(n3808), .IN2(n15174), .QN(n15173) );
  NOR2X0 U15424 ( .IN1(n15175), .IN2(n15176), .QN(n15172) );
  NOR2X0 U15425 ( .IN1(n11030), .IN2(n15177), .QN(n15176) );
  NAND2X0 U15426 ( .IN1(n15178), .IN2(g6299), .QN(n15177) );
  NAND2X0 U15427 ( .IN1(n15165), .IN2(n15174), .QN(n15178) );
  NOR2X0 U15428 ( .IN1(n10386), .IN2(n10865), .QN(n15175) );
  NAND2X0 U15429 ( .IN1(n15179), .IN2(n15180), .QN(g30535) );
  NAND2X0 U15430 ( .IN1(n3808), .IN2(n15181), .QN(n15180) );
  NOR2X0 U15431 ( .IN1(n15182), .IN2(n15183), .QN(n15179) );
  NOR2X0 U15432 ( .IN1(n11030), .IN2(n15184), .QN(n15183) );
  NAND2X0 U15433 ( .IN1(n15185), .IN2(g6295), .QN(n15184) );
  NAND2X0 U15434 ( .IN1(n15165), .IN2(n15181), .QN(n15185) );
  INVX0 U15435 ( .INP(n3414), .ZN(n15165) );
  NAND2X0 U15436 ( .IN1(g6203), .IN2(g6209), .QN(n3414) );
  NOR2X0 U15437 ( .IN1(n10438), .IN2(n10865), .QN(n15182) );
  NAND2X0 U15438 ( .IN1(n15186), .IN2(n15187), .QN(g30534) );
  NAND2X0 U15439 ( .IN1(n3814), .IN2(n15160), .QN(n15187) );
  NOR2X0 U15440 ( .IN1(n15188), .IN2(n15189), .QN(n15186) );
  NOR2X0 U15441 ( .IN1(n11030), .IN2(n15190), .QN(n15189) );
  NAND2X0 U15442 ( .IN1(n15191), .IN2(g6291), .QN(n15190) );
  NAND2X0 U15443 ( .IN1(n14250), .IN2(n15160), .QN(n15191) );
  NOR2X0 U15444 ( .IN1(n10356), .IN2(n10866), .QN(n15188) );
  NAND2X0 U15445 ( .IN1(n15192), .IN2(n15193), .QN(g30533) );
  NAND2X0 U15446 ( .IN1(n3814), .IN2(n14232), .QN(n15193) );
  NOR2X0 U15447 ( .IN1(n15194), .IN2(n15195), .QN(n15192) );
  NOR2X0 U15448 ( .IN1(n11030), .IN2(n15196), .QN(n15195) );
  NAND2X0 U15449 ( .IN1(n15197), .IN2(g6287), .QN(n15196) );
  NAND2X0 U15450 ( .IN1(n14250), .IN2(n14232), .QN(n15197) );
  NOR2X0 U15451 ( .IN1(n10429), .IN2(n10866), .QN(n15194) );
  NAND2X0 U15452 ( .IN1(n15198), .IN2(n15199), .QN(g30532) );
  NAND2X0 U15453 ( .IN1(n3814), .IN2(n15174), .QN(n15199) );
  NOR2X0 U15454 ( .IN1(n15200), .IN2(n15201), .QN(n15198) );
  NOR2X0 U15455 ( .IN1(n11029), .IN2(n15202), .QN(n15201) );
  NAND2X0 U15456 ( .IN1(n15203), .IN2(g6283), .QN(n15202) );
  NAND2X0 U15457 ( .IN1(n14250), .IN2(n15174), .QN(n15203) );
  NOR2X0 U15458 ( .IN1(n10333), .IN2(n10866), .QN(n15200) );
  NAND2X0 U15459 ( .IN1(n15204), .IN2(n15205), .QN(g30531) );
  NAND2X0 U15460 ( .IN1(n3814), .IN2(n15181), .QN(n15205) );
  NOR2X0 U15461 ( .IN1(n15206), .IN2(n15207), .QN(n15204) );
  NOR2X0 U15462 ( .IN1(n11029), .IN2(n15208), .QN(n15207) );
  NAND2X0 U15463 ( .IN1(n15209), .IN2(g6279), .QN(n15208) );
  NAND2X0 U15464 ( .IN1(n14250), .IN2(n15181), .QN(n15209) );
  INVX0 U15465 ( .INP(n3416), .ZN(n14250) );
  NAND2X0 U15466 ( .IN1(n5574), .IN2(g6209), .QN(n3416) );
  NOR2X0 U15467 ( .IN1(n10301), .IN2(n10866), .QN(n15206) );
  NAND2X0 U15468 ( .IN1(n15210), .IN2(n15211), .QN(g30530) );
  NAND2X0 U15469 ( .IN1(n3819), .IN2(n15160), .QN(n15211) );
  NOR2X0 U15470 ( .IN1(n15212), .IN2(n15213), .QN(n15210) );
  NOR2X0 U15471 ( .IN1(n11029), .IN2(n15214), .QN(n15213) );
  NAND2X0 U15472 ( .IN1(n15215), .IN2(g6275), .QN(n15214) );
  NAND2X0 U15473 ( .IN1(n15216), .IN2(n15160), .QN(n15215) );
  NOR2X0 U15474 ( .IN1(n10430), .IN2(n10866), .QN(n15212) );
  NAND2X0 U15475 ( .IN1(n15217), .IN2(n15218), .QN(g30529) );
  NAND2X0 U15476 ( .IN1(n3819), .IN2(n14232), .QN(n15218) );
  NOR2X0 U15477 ( .IN1(n15219), .IN2(n15220), .QN(n15217) );
  NOR2X0 U15478 ( .IN1(n11029), .IN2(n15221), .QN(n15220) );
  NAND2X0 U15479 ( .IN1(n15222), .IN2(g6271), .QN(n15221) );
  NAND2X0 U15480 ( .IN1(n15216), .IN2(n14232), .QN(n15222) );
  INVX0 U15481 ( .INP(n3802), .ZN(n14232) );
  NAND2X0 U15482 ( .IN1(n5385), .IN2(g6227), .QN(n3802) );
  NOR2X0 U15483 ( .IN1(n10520), .IN2(n10867), .QN(n15219) );
  NAND2X0 U15484 ( .IN1(n15223), .IN2(n15224), .QN(g30528) );
  NAND2X0 U15485 ( .IN1(n3819), .IN2(n15174), .QN(n15224) );
  NOR2X0 U15486 ( .IN1(n15225), .IN2(n15226), .QN(n15223) );
  NOR2X0 U15487 ( .IN1(n11028), .IN2(n15227), .QN(n15226) );
  NAND2X0 U15488 ( .IN1(n15228), .IN2(g6267), .QN(n15227) );
  NAND2X0 U15489 ( .IN1(n15216), .IN2(n15174), .QN(n15228) );
  INVX0 U15490 ( .INP(n3804), .ZN(n15174) );
  NAND2X0 U15491 ( .IN1(n5568), .IN2(g6219), .QN(n3804) );
  NOR2X0 U15492 ( .IN1(n10302), .IN2(n10867), .QN(n15225) );
  NAND2X0 U15493 ( .IN1(n15229), .IN2(n15230), .QN(g30527) );
  NAND2X0 U15494 ( .IN1(n3819), .IN2(n15181), .QN(n15230) );
  NOR2X0 U15495 ( .IN1(n15231), .IN2(n15232), .QN(n15229) );
  NOR2X0 U15496 ( .IN1(n11028), .IN2(n15233), .QN(n15232) );
  NAND2X0 U15497 ( .IN1(n15234), .IN2(g6263), .QN(n15233) );
  NAND2X0 U15498 ( .IN1(n15216), .IN2(n15181), .QN(n15234) );
  INVX0 U15499 ( .INP(n3807), .ZN(n15181) );
  NAND2X0 U15500 ( .IN1(n5568), .IN2(n5385), .QN(n3807) );
  INVX0 U15501 ( .INP(n3417), .ZN(n15216) );
  NAND2X0 U15502 ( .IN1(n10588), .IN2(g6203), .QN(n3417) );
  NOR2X0 U15503 ( .IN1(n10454), .IN2(n10867), .QN(n15231) );
  NAND2X0 U15504 ( .IN1(n15235), .IN2(n15236), .QN(g30526) );
  NAND2X0 U15505 ( .IN1(n11077), .IN2(g6259), .QN(n15236) );
  NOR2X0 U15506 ( .IN1(n15237), .IN2(n15238), .QN(n15235) );
  NOR2X0 U15507 ( .IN1(n15008), .IN2(n15239), .QN(n15238) );
  INVX0 U15508 ( .INP(n3824), .ZN(n15239) );
  NOR2X0 U15509 ( .IN1(n3824), .IN2(n15240), .QN(n15237) );
  NAND2X0 U15510 ( .IN1(n10934), .IN2(g6255), .QN(n15240) );
  NAND2X0 U15511 ( .IN1(n15241), .IN2(n15242), .QN(g30525) );
  NAND2X0 U15512 ( .IN1(n11078), .IN2(g6251), .QN(n15242) );
  NOR2X0 U15513 ( .IN1(n15243), .IN2(n15244), .QN(n15241) );
  NOR2X0 U15514 ( .IN1(n15008), .IN2(n15245), .QN(n15244) );
  INVX0 U15515 ( .INP(n3827), .ZN(n15245) );
  NOR2X0 U15516 ( .IN1(n3827), .IN2(n15246), .QN(n15243) );
  NAND2X0 U15517 ( .IN1(n10934), .IN2(g6247), .QN(n15246) );
  NAND2X0 U15518 ( .IN1(n15247), .IN2(n15248), .QN(g30524) );
  NAND2X0 U15519 ( .IN1(n11078), .IN2(g6243), .QN(n15248) );
  NOR2X0 U15520 ( .IN1(n15249), .IN2(n15250), .QN(n15247) );
  NOR2X0 U15521 ( .IN1(n15008), .IN2(n15251), .QN(n15250) );
  INVX0 U15522 ( .INP(n3829), .ZN(n15251) );
  NOR2X0 U15523 ( .IN1(n3829), .IN2(n15252), .QN(n15249) );
  NAND2X0 U15524 ( .IN1(n10936), .IN2(g6239), .QN(n15252) );
  NAND2X0 U15525 ( .IN1(n15253), .IN2(n15254), .QN(g30523) );
  NAND2X0 U15526 ( .IN1(n11078), .IN2(g6227), .QN(n15254) );
  NOR2X0 U15527 ( .IN1(n15255), .IN2(n15256), .QN(n15253) );
  NOR2X0 U15528 ( .IN1(n15008), .IN2(n15257), .QN(n15256) );
  INVX0 U15529 ( .INP(n3831), .ZN(n15257) );
  NOR2X0 U15530 ( .IN1(n3831), .IN2(n15258), .QN(n15255) );
  NAND2X0 U15531 ( .IN1(n10935), .IN2(g6235), .QN(n15258) );
  NOR2X0 U15532 ( .IN1(g6203), .IN2(n14241), .QN(g30522) );
  NAND2X0 U15533 ( .IN1(n15259), .IN2(n5651), .QN(n14241) );
  NOR2X0 U15534 ( .IN1(n11028), .IN2(n14245), .QN(n15259) );
  INVX0 U15535 ( .INP(n14229), .ZN(n14245) );
  NAND2X0 U15536 ( .IN1(n15260), .IN2(n3833), .QN(n14229) );
  NAND2X0 U15537 ( .IN1(n15261), .IN2(n15262), .QN(g30521) );
  NAND2X0 U15538 ( .IN1(n11078), .IN2(g5961), .QN(n15262) );
  NOR2X0 U15539 ( .IN1(n15263), .IN2(n15264), .QN(n15261) );
  NOR2X0 U15540 ( .IN1(n15008), .IN2(n13433), .QN(n15264) );
  NOR2X0 U15541 ( .IN1(n15265), .IN2(n10684), .QN(n15263) );
  NAND2X0 U15542 ( .IN1(n15266), .IN2(n15267), .QN(g30520) );
  NAND2X0 U15543 ( .IN1(n15268), .IN2(n3765), .QN(n15267) );
  NOR2X0 U15544 ( .IN1(n15269), .IN2(n15270), .QN(n15266) );
  NOR2X0 U15545 ( .IN1(n10467), .IN2(n10868), .QN(n15270) );
  NOR2X0 U15546 ( .IN1(n11028), .IN2(n15271), .QN(n15269) );
  NAND2X0 U15547 ( .IN1(n15272), .IN2(g5913), .QN(n15271) );
  INVX0 U15548 ( .INP(n15268), .ZN(n15272) );
  NOR2X0 U15549 ( .IN1(n3836), .IN2(n5649), .QN(n15268) );
  NAND2X0 U15550 ( .IN1(n15273), .IN2(n15274), .QN(g30519) );
  NAND2X0 U15551 ( .IN1(n14258), .IN2(n3765), .QN(n15274) );
  NOR2X0 U15552 ( .IN1(n15275), .IN2(n15276), .QN(n15273) );
  NOR2X0 U15553 ( .IN1(n10362), .IN2(n10868), .QN(n15276) );
  NOR2X0 U15554 ( .IN1(n11028), .IN2(n15277), .QN(n15275) );
  INVX0 U15555 ( .INP(n15278), .ZN(n15277) );
  NOR2X0 U15556 ( .IN1(n14258), .IN2(n10469), .QN(n15278) );
  NOR2X0 U15557 ( .IN1(n3838), .IN2(n5649), .QN(n14258) );
  NAND2X0 U15558 ( .IN1(n15279), .IN2(n15280), .QN(g30518) );
  NAND2X0 U15559 ( .IN1(n15281), .IN2(n3765), .QN(n15280) );
  NOR2X0 U15560 ( .IN1(n15282), .IN2(n15283), .QN(n15279) );
  NOR2X0 U15561 ( .IN1(n10307), .IN2(n10868), .QN(n15283) );
  NOR2X0 U15562 ( .IN1(n11027), .IN2(n15284), .QN(n15282) );
  NAND2X0 U15563 ( .IN1(n15285), .IN2(g5897), .QN(n15284) );
  INVX0 U15564 ( .INP(n15281), .ZN(n15285) );
  NOR2X0 U15565 ( .IN1(n3841), .IN2(n5649), .QN(n15281) );
  NAND2X0 U15566 ( .IN1(n15286), .IN2(n15287), .QN(g30517) );
  NAND2X0 U15567 ( .IN1(n3842), .IN2(n15288), .QN(n15287) );
  NOR2X0 U15568 ( .IN1(n15289), .IN2(n15290), .QN(n15286) );
  NOR2X0 U15569 ( .IN1(n11028), .IN2(n15291), .QN(n15290) );
  NAND2X0 U15570 ( .IN1(n15292), .IN2(g5961), .QN(n15291) );
  NAND2X0 U15571 ( .IN1(n15293), .IN2(n15288), .QN(n15292) );
  NOR2X0 U15572 ( .IN1(n10340), .IN2(n10868), .QN(n15289) );
  NAND2X0 U15573 ( .IN1(n15294), .IN2(n15295), .QN(g30516) );
  NAND2X0 U15574 ( .IN1(n3842), .IN2(n14257), .QN(n15295) );
  NOR2X0 U15575 ( .IN1(n15296), .IN2(n15297), .QN(n15294) );
  NOR2X0 U15576 ( .IN1(n11027), .IN2(n15298), .QN(n15297) );
  NAND2X0 U15577 ( .IN1(n15299), .IN2(g5957), .QN(n15298) );
  NAND2X0 U15578 ( .IN1(n15293), .IN2(n14257), .QN(n15299) );
  NOR2X0 U15579 ( .IN1(n10465), .IN2(n10869), .QN(n15296) );
  NAND2X0 U15580 ( .IN1(n15300), .IN2(n15301), .QN(g30515) );
  NAND2X0 U15581 ( .IN1(n3842), .IN2(n15302), .QN(n15301) );
  NOR2X0 U15582 ( .IN1(n15303), .IN2(n15304), .QN(n15300) );
  NOR2X0 U15583 ( .IN1(n11027), .IN2(n15305), .QN(n15304) );
  NAND2X0 U15584 ( .IN1(n15306), .IN2(g5953), .QN(n15305) );
  NAND2X0 U15585 ( .IN1(n15293), .IN2(n15302), .QN(n15306) );
  NOR2X0 U15586 ( .IN1(n10377), .IN2(n10869), .QN(n15303) );
  NAND2X0 U15587 ( .IN1(n15307), .IN2(n15308), .QN(g30514) );
  NAND2X0 U15588 ( .IN1(n3842), .IN2(n15309), .QN(n15308) );
  NOR2X0 U15589 ( .IN1(n15310), .IN2(n15311), .QN(n15307) );
  NOR2X0 U15590 ( .IN1(n11027), .IN2(n15312), .QN(n15311) );
  NAND2X0 U15591 ( .IN1(n15313), .IN2(g5949), .QN(n15312) );
  NAND2X0 U15592 ( .IN1(n15293), .IN2(n15309), .QN(n15313) );
  INVX0 U15593 ( .INP(n3424), .ZN(n15293) );
  NAND2X0 U15594 ( .IN1(g5857), .IN2(g5863), .QN(n3424) );
  NOR2X0 U15595 ( .IN1(n10433), .IN2(n10869), .QN(n15310) );
  NAND2X0 U15596 ( .IN1(n15314), .IN2(n15315), .QN(g30513) );
  NAND2X0 U15597 ( .IN1(n3848), .IN2(n15288), .QN(n15315) );
  NOR2X0 U15598 ( .IN1(n15316), .IN2(n15317), .QN(n15314) );
  NOR2X0 U15599 ( .IN1(n11027), .IN2(n15318), .QN(n15317) );
  NAND2X0 U15600 ( .IN1(n15319), .IN2(g5945), .QN(n15318) );
  NAND2X0 U15601 ( .IN1(n14275), .IN2(n15288), .QN(n15319) );
  NOR2X0 U15602 ( .IN1(n10341), .IN2(n10869), .QN(n15316) );
  NAND2X0 U15603 ( .IN1(n15320), .IN2(n15321), .QN(g30512) );
  NAND2X0 U15604 ( .IN1(n3848), .IN2(n14257), .QN(n15321) );
  NOR2X0 U15605 ( .IN1(n15322), .IN2(n15323), .QN(n15320) );
  NOR2X0 U15606 ( .IN1(n11027), .IN2(n15324), .QN(n15323) );
  NAND2X0 U15607 ( .IN1(n15325), .IN2(g5941), .QN(n15324) );
  NAND2X0 U15608 ( .IN1(n14275), .IN2(n14257), .QN(n15325) );
  NOR2X0 U15609 ( .IN1(n10414), .IN2(n10869), .QN(n15322) );
  NAND2X0 U15610 ( .IN1(n15326), .IN2(n15327), .QN(g30511) );
  NAND2X0 U15611 ( .IN1(n3848), .IN2(n15302), .QN(n15327) );
  NOR2X0 U15612 ( .IN1(n15328), .IN2(n15329), .QN(n15326) );
  NOR2X0 U15613 ( .IN1(n11027), .IN2(n15330), .QN(n15329) );
  NAND2X0 U15614 ( .IN1(n15331), .IN2(g5937), .QN(n15330) );
  NAND2X0 U15615 ( .IN1(n14275), .IN2(n15302), .QN(n15331) );
  NOR2X0 U15616 ( .IN1(n10328), .IN2(n10870), .QN(n15328) );
  NAND2X0 U15617 ( .IN1(n15332), .IN2(n15333), .QN(g30510) );
  NAND2X0 U15618 ( .IN1(n3848), .IN2(n15309), .QN(n15333) );
  NOR2X0 U15619 ( .IN1(n15334), .IN2(n15335), .QN(n15332) );
  NOR2X0 U15620 ( .IN1(n11027), .IN2(n15336), .QN(n15335) );
  NAND2X0 U15621 ( .IN1(n15337), .IN2(g5933), .QN(n15336) );
  NAND2X0 U15622 ( .IN1(n14275), .IN2(n15309), .QN(n15337) );
  INVX0 U15623 ( .INP(n1101), .ZN(n14275) );
  NAND2X0 U15624 ( .IN1(n5573), .IN2(g5863), .QN(n1101) );
  NOR2X0 U15625 ( .IN1(n10907), .IN2(n10685), .QN(n15334) );
  NAND2X0 U15626 ( .IN1(n15338), .IN2(n15339), .QN(g30509) );
  NAND2X0 U15627 ( .IN1(n3853), .IN2(n15288), .QN(n15339) );
  NOR2X0 U15628 ( .IN1(n15340), .IN2(n15341), .QN(n15338) );
  NOR2X0 U15629 ( .IN1(n11027), .IN2(n15342), .QN(n15341) );
  NAND2X0 U15630 ( .IN1(n15343), .IN2(g5929), .QN(n15342) );
  NAND2X0 U15631 ( .IN1(n15344), .IN2(n15288), .QN(n15343) );
  NOR2X0 U15632 ( .IN1(n10415), .IN2(n10870), .QN(n15340) );
  NAND2X0 U15633 ( .IN1(n15345), .IN2(n15346), .QN(g30508) );
  NAND2X0 U15634 ( .IN1(n3853), .IN2(n14257), .QN(n15346) );
  NOR2X0 U15635 ( .IN1(n15347), .IN2(n15348), .QN(n15345) );
  NOR2X0 U15636 ( .IN1(n11026), .IN2(n15349), .QN(n15348) );
  NAND2X0 U15637 ( .IN1(n15350), .IN2(g5925), .QN(n15349) );
  NAND2X0 U15638 ( .IN1(n15344), .IN2(n14257), .QN(n15350) );
  INVX0 U15639 ( .INP(n3836), .ZN(n14257) );
  NAND2X0 U15640 ( .IN1(n5388), .IN2(test_so36), .QN(n3836) );
  NOR2X0 U15641 ( .IN1(n10500), .IN2(n10870), .QN(n15347) );
  NAND2X0 U15642 ( .IN1(n15351), .IN2(n15352), .QN(g30507) );
  NAND2X0 U15643 ( .IN1(n3853), .IN2(n15302), .QN(n15352) );
  NOR2X0 U15644 ( .IN1(n15353), .IN2(n15354), .QN(n15351) );
  NOR2X0 U15645 ( .IN1(n11028), .IN2(n15355), .QN(n15354) );
  NAND2X0 U15646 ( .IN1(n15356), .IN2(g5921), .QN(n15355) );
  NAND2X0 U15647 ( .IN1(n15344), .IN2(n15302), .QN(n15356) );
  INVX0 U15648 ( .INP(n3838), .ZN(n15302) );
  NAND2X0 U15649 ( .IN1(n10651), .IN2(g5873), .QN(n3838) );
  NOR2X0 U15650 ( .IN1(n10308), .IN2(n10870), .QN(n15353) );
  NAND2X0 U15651 ( .IN1(n15357), .IN2(n15358), .QN(g30506) );
  NAND2X0 U15652 ( .IN1(n3853), .IN2(n15309), .QN(n15358) );
  NOR2X0 U15653 ( .IN1(n15359), .IN2(n15360), .QN(n15357) );
  NOR2X0 U15654 ( .IN1(n11026), .IN2(n15361), .QN(n15360) );
  NAND2X0 U15655 ( .IN1(test_so28), .IN2(n15362), .QN(n15361) );
  NAND2X0 U15656 ( .IN1(n15344), .IN2(n15309), .QN(n15362) );
  INVX0 U15657 ( .INP(n3841), .ZN(n15309) );
  NAND2X0 U15658 ( .IN1(n5388), .IN2(n10651), .QN(n3841) );
  INVX0 U15659 ( .INP(n3427), .ZN(n15344) );
  NAND2X0 U15660 ( .IN1(n10590), .IN2(g5857), .QN(n3427) );
  NOR2X0 U15661 ( .IN1(n10445), .IN2(n10870), .QN(n15359) );
  NAND2X0 U15662 ( .IN1(n15363), .IN2(n15364), .QN(g30505) );
  NAND2X0 U15663 ( .IN1(n11078), .IN2(g5913), .QN(n15364) );
  NOR2X0 U15664 ( .IN1(n15365), .IN2(n15366), .QN(n15363) );
  NOR2X0 U15665 ( .IN1(n15008), .IN2(n15367), .QN(n15366) );
  INVX0 U15666 ( .INP(n3858), .ZN(n15367) );
  NOR2X0 U15667 ( .IN1(n3858), .IN2(n15368), .QN(n15365) );
  NAND2X0 U15668 ( .IN1(n10935), .IN2(g5909), .QN(n15368) );
  NAND2X0 U15669 ( .IN1(n15369), .IN2(n15370), .QN(g30504) );
  NAND2X0 U15670 ( .IN1(n11078), .IN2(g5905), .QN(n15370) );
  NOR2X0 U15671 ( .IN1(n15371), .IN2(n15372), .QN(n15369) );
  NOR2X0 U15672 ( .IN1(n15008), .IN2(n15373), .QN(n15372) );
  INVX0 U15673 ( .INP(n3861), .ZN(n15373) );
  NOR2X0 U15674 ( .IN1(n3861), .IN2(n15374), .QN(n15371) );
  NAND2X0 U15675 ( .IN1(n10936), .IN2(g5901), .QN(n15374) );
  NAND2X0 U15676 ( .IN1(n15375), .IN2(n15376), .QN(g30503) );
  NAND2X0 U15677 ( .IN1(n11078), .IN2(g5897), .QN(n15376) );
  NOR2X0 U15678 ( .IN1(n15377), .IN2(n15378), .QN(n15375) );
  NOR2X0 U15679 ( .IN1(n15008), .IN2(n15379), .QN(n15378) );
  INVX0 U15680 ( .INP(n3863), .ZN(n15379) );
  NOR2X0 U15681 ( .IN1(n3863), .IN2(n15380), .QN(n15377) );
  NAND2X0 U15682 ( .IN1(n10934), .IN2(g5893), .QN(n15380) );
  NAND2X0 U15683 ( .IN1(n15381), .IN2(n15382), .QN(g30502) );
  NAND2X0 U15684 ( .IN1(test_so36), .IN2(n11014), .QN(n15382) );
  NOR2X0 U15685 ( .IN1(n15383), .IN2(n15384), .QN(n15381) );
  NOR2X0 U15686 ( .IN1(n15008), .IN2(n15385), .QN(n15384) );
  INVX0 U15687 ( .INP(n3865), .ZN(n15385) );
  NOR2X0 U15688 ( .IN1(n3865), .IN2(n15386), .QN(n15383) );
  NAND2X0 U15689 ( .IN1(n10936), .IN2(g5889), .QN(n15386) );
  NOR2X0 U15690 ( .IN1(g5857), .IN2(n14266), .QN(g30501) );
  NAND2X0 U15691 ( .IN1(n15387), .IN2(n5649), .QN(n14266) );
  NOR2X0 U15692 ( .IN1(n11027), .IN2(n14270), .QN(n15387) );
  INVX0 U15693 ( .INP(n14254), .ZN(n14270) );
  NAND2X0 U15694 ( .IN1(n15388), .IN2(n3833), .QN(n14254) );
  NAND2X0 U15695 ( .IN1(n15389), .IN2(n15390), .QN(g30500) );
  NAND2X0 U15696 ( .IN1(n11077), .IN2(g5615), .QN(n15390) );
  NOR2X0 U15697 ( .IN1(n15391), .IN2(n15392), .QN(n15389) );
  NOR2X0 U15698 ( .IN1(n15393), .IN2(n15008), .QN(n15392) );
  NOR2X0 U15699 ( .IN1(n10288), .IN2(n11251), .QN(n15391) );
  NAND2X0 U15700 ( .IN1(n15394), .IN2(n15395), .QN(g30499) );
  NAND2X0 U15701 ( .IN1(n15396), .IN2(n3765), .QN(n15395) );
  NOR2X0 U15702 ( .IN1(n15397), .IN2(n15398), .QN(n15394) );
  NOR2X0 U15703 ( .IN1(n10472), .IN2(n10872), .QN(n15398) );
  NOR2X0 U15704 ( .IN1(n11027), .IN2(n15399), .QN(n15397) );
  NAND2X0 U15705 ( .IN1(n15400), .IN2(g5567), .QN(n15399) );
  INVX0 U15706 ( .INP(n15396), .ZN(n15400) );
  NOR2X0 U15707 ( .IN1(n3869), .IN2(n5647), .QN(n15396) );
  NAND2X0 U15708 ( .IN1(n15401), .IN2(n15402), .QN(g30498) );
  NAND2X0 U15709 ( .IN1(n14283), .IN2(n3765), .QN(n15402) );
  INVX0 U15710 ( .INP(n15403), .ZN(n14283) );
  NOR2X0 U15711 ( .IN1(n15404), .IN2(n15405), .QN(n15401) );
  NOR2X0 U15712 ( .IN1(n10364), .IN2(n10872), .QN(n15405) );
  NOR2X0 U15713 ( .IN1(n11026), .IN2(n15406), .QN(n15404) );
  NAND2X0 U15714 ( .IN1(test_so6), .IN2(n15403), .QN(n15406) );
  NAND2X0 U15715 ( .IN1(n15407), .IN2(g5523), .QN(n15403) );
  NAND2X0 U15716 ( .IN1(n15408), .IN2(n15409), .QN(g30497) );
  NAND2X0 U15717 ( .IN1(n15410), .IN2(n3765), .QN(n15409) );
  NOR2X0 U15718 ( .IN1(n15411), .IN2(n15412), .QN(n15408) );
  NOR2X0 U15719 ( .IN1(n10289), .IN2(n10872), .QN(n15412) );
  NOR2X0 U15720 ( .IN1(n11026), .IN2(n15413), .QN(n15411) );
  NAND2X0 U15721 ( .IN1(n15414), .IN2(g5551), .QN(n15413) );
  INVX0 U15722 ( .INP(n15410), .ZN(n15414) );
  NOR2X0 U15723 ( .IN1(n3874), .IN2(n5647), .QN(n15410) );
  NAND2X0 U15724 ( .IN1(n15415), .IN2(n15416), .QN(g30496) );
  NAND2X0 U15725 ( .IN1(n3875), .IN2(n15417), .QN(n15416) );
  NOR2X0 U15726 ( .IN1(n15418), .IN2(n15419), .QN(n15415) );
  NOR2X0 U15727 ( .IN1(n11025), .IN2(n15420), .QN(n15419) );
  NAND2X0 U15728 ( .IN1(n15421), .IN2(g5615), .QN(n15420) );
  NAND2X0 U15729 ( .IN1(n15422), .IN2(n15417), .QN(n15421) );
  NOR2X0 U15730 ( .IN1(n10343), .IN2(n10872), .QN(n15418) );
  NAND2X0 U15731 ( .IN1(n15423), .IN2(n15424), .QN(g30495) );
  NAND2X0 U15732 ( .IN1(n3875), .IN2(n14282), .QN(n15424) );
  NOR2X0 U15733 ( .IN1(n15425), .IN2(n15426), .QN(n15423) );
  NOR2X0 U15734 ( .IN1(n11026), .IN2(n15427), .QN(n15426) );
  NAND2X0 U15735 ( .IN1(n15428), .IN2(g5611), .QN(n15427) );
  NAND2X0 U15736 ( .IN1(n15422), .IN2(n14282), .QN(n15428) );
  NOR2X0 U15737 ( .IN1(n10470), .IN2(n10872), .QN(n15425) );
  NAND2X0 U15738 ( .IN1(n15429), .IN2(n15430), .QN(g30494) );
  NAND2X0 U15739 ( .IN1(n3875), .IN2(n15407), .QN(n15430) );
  NOR2X0 U15740 ( .IN1(n15431), .IN2(n15432), .QN(n15429) );
  NOR2X0 U15741 ( .IN1(n11025), .IN2(n15433), .QN(n15432) );
  NAND2X0 U15742 ( .IN1(n15434), .IN2(g5607), .QN(n15433) );
  NAND2X0 U15743 ( .IN1(n15422), .IN2(n15407), .QN(n15434) );
  NOR2X0 U15744 ( .IN1(n10905), .IN2(n10688), .QN(n15431) );
  NAND2X0 U15745 ( .IN1(n15435), .IN2(n15436), .QN(g30493) );
  NAND2X0 U15746 ( .IN1(n3875), .IN2(n15437), .QN(n15436) );
  NOR2X0 U15747 ( .IN1(n15438), .IN2(n15439), .QN(n15435) );
  NOR2X0 U15748 ( .IN1(n11026), .IN2(n15440), .QN(n15439) );
  NAND2X0 U15749 ( .IN1(n15441), .IN2(g5603), .QN(n15440) );
  NAND2X0 U15750 ( .IN1(n15422), .IN2(n15437), .QN(n15441) );
  INVX0 U15751 ( .INP(n3434), .ZN(n15422) );
  NAND2X0 U15752 ( .IN1(g5511), .IN2(g5517), .QN(n3434) );
  NOR2X0 U15753 ( .IN1(n10434), .IN2(n10873), .QN(n15438) );
  NAND2X0 U15754 ( .IN1(n15442), .IN2(n15443), .QN(g30492) );
  NAND2X0 U15755 ( .IN1(n3881), .IN2(n15417), .QN(n15443) );
  NOR2X0 U15756 ( .IN1(n15444), .IN2(n15445), .QN(n15442) );
  NOR2X0 U15757 ( .IN1(n11025), .IN2(n15446), .QN(n15445) );
  NAND2X0 U15758 ( .IN1(n15447), .IN2(g5599), .QN(n15446) );
  NAND2X0 U15759 ( .IN1(n15417), .IN2(n14300), .QN(n15447) );
  NOR2X0 U15760 ( .IN1(n10344), .IN2(n10873), .QN(n15444) );
  NAND2X0 U15761 ( .IN1(n15448), .IN2(n15449), .QN(g30491) );
  NAND2X0 U15762 ( .IN1(n3881), .IN2(n14282), .QN(n15449) );
  NOR2X0 U15763 ( .IN1(n15450), .IN2(n15451), .QN(n15448) );
  NOR2X0 U15764 ( .IN1(n11026), .IN2(n15452), .QN(n15451) );
  NAND2X0 U15765 ( .IN1(n15453), .IN2(g5595), .QN(n15452) );
  NAND2X0 U15766 ( .IN1(n14282), .IN2(n14300), .QN(n15453) );
  NOR2X0 U15767 ( .IN1(n10417), .IN2(n10873), .QN(n15450) );
  NAND2X0 U15768 ( .IN1(n15454), .IN2(n15455), .QN(g30490) );
  NAND2X0 U15769 ( .IN1(n3881), .IN2(n15407), .QN(n15455) );
  NOR2X0 U15770 ( .IN1(n15456), .IN2(n15457), .QN(n15454) );
  NOR2X0 U15771 ( .IN1(n11027), .IN2(n15458), .QN(n15457) );
  NAND2X0 U15772 ( .IN1(test_so5), .IN2(n15459), .QN(n15458) );
  NAND2X0 U15773 ( .IN1(n14300), .IN2(n15407), .QN(n15459) );
  NOR2X0 U15774 ( .IN1(n10329), .IN2(n10873), .QN(n15456) );
  NAND2X0 U15775 ( .IN1(n15460), .IN2(n15461), .QN(g30489) );
  NAND2X0 U15776 ( .IN1(n3881), .IN2(n15437), .QN(n15461) );
  NOR2X0 U15777 ( .IN1(n15462), .IN2(n15463), .QN(n15460) );
  NOR2X0 U15778 ( .IN1(n11026), .IN2(n15464), .QN(n15463) );
  NAND2X0 U15779 ( .IN1(n15465), .IN2(g5587), .QN(n15464) );
  NAND2X0 U15780 ( .IN1(n15437), .IN2(n14300), .QN(n15465) );
  INVX0 U15781 ( .INP(n552), .ZN(n14300) );
  NAND2X0 U15782 ( .IN1(n5575), .IN2(g5517), .QN(n552) );
  NOR2X0 U15783 ( .IN1(n10290), .IN2(n10873), .QN(n15462) );
  NAND2X0 U15784 ( .IN1(n15466), .IN2(n15467), .QN(g30488) );
  NAND2X0 U15785 ( .IN1(n3886), .IN2(n15417), .QN(n15467) );
  NOR2X0 U15786 ( .IN1(n15468), .IN2(n15469), .QN(n15466) );
  NOR2X0 U15787 ( .IN1(n11025), .IN2(n15470), .QN(n15469) );
  NAND2X0 U15788 ( .IN1(n15471), .IN2(g5583), .QN(n15470) );
  NAND2X0 U15789 ( .IN1(n15472), .IN2(n15417), .QN(n15471) );
  NOR2X0 U15790 ( .IN1(n10418), .IN2(n10874), .QN(n15468) );
  NAND2X0 U15791 ( .IN1(n15473), .IN2(n15474), .QN(g30487) );
  NAND2X0 U15792 ( .IN1(n3886), .IN2(n14282), .QN(n15474) );
  NOR2X0 U15793 ( .IN1(n15475), .IN2(n15476), .QN(n15473) );
  NOR2X0 U15794 ( .IN1(n11026), .IN2(n15477), .QN(n15476) );
  NAND2X0 U15795 ( .IN1(n15478), .IN2(g5579), .QN(n15477) );
  NAND2X0 U15796 ( .IN1(n15472), .IN2(n14282), .QN(n15478) );
  INVX0 U15797 ( .INP(n3869), .ZN(n14282) );
  NAND2X0 U15798 ( .IN1(n5389), .IN2(g5535), .QN(n3869) );
  NOR2X0 U15799 ( .IN1(n10504), .IN2(n10874), .QN(n15475) );
  NAND2X0 U15800 ( .IN1(n15479), .IN2(n15480), .QN(g30486) );
  NAND2X0 U15801 ( .IN1(n3886), .IN2(n15407), .QN(n15480) );
  NOR2X0 U15802 ( .IN1(n15481), .IN2(n15482), .QN(n15479) );
  NOR2X0 U15803 ( .IN1(n11026), .IN2(n15483), .QN(n15482) );
  NAND2X0 U15804 ( .IN1(n15484), .IN2(g5575), .QN(n15483) );
  NAND2X0 U15805 ( .IN1(n15472), .IN2(n15407), .QN(n15484) );
  INVX0 U15806 ( .INP(n978), .ZN(n15407) );
  NAND2X0 U15807 ( .IN1(n5566), .IN2(g5527), .QN(n978) );
  NOR2X0 U15808 ( .IN1(n10291), .IN2(n10874), .QN(n15481) );
  NAND2X0 U15809 ( .IN1(n15485), .IN2(n15486), .QN(g30485) );
  NAND2X0 U15810 ( .IN1(n3886), .IN2(n15437), .QN(n15486) );
  NOR2X0 U15811 ( .IN1(n15487), .IN2(n15488), .QN(n15485) );
  NOR2X0 U15812 ( .IN1(n11025), .IN2(n15489), .QN(n15488) );
  NAND2X0 U15813 ( .IN1(n15490), .IN2(g5571), .QN(n15489) );
  NAND2X0 U15814 ( .IN1(n15472), .IN2(n15437), .QN(n15490) );
  INVX0 U15815 ( .INP(n3874), .ZN(n15437) );
  NAND2X0 U15816 ( .IN1(n5389), .IN2(n5566), .QN(n3874) );
  INVX0 U15817 ( .INP(n3437), .ZN(n15472) );
  NAND2X0 U15818 ( .IN1(n10589), .IN2(g5511), .QN(n3437) );
  NOR2X0 U15819 ( .IN1(n10447), .IN2(n10874), .QN(n15487) );
  NAND2X0 U15820 ( .IN1(n15491), .IN2(n15492), .QN(g30484) );
  NAND2X0 U15821 ( .IN1(n11077), .IN2(g5567), .QN(n15492) );
  NOR2X0 U15822 ( .IN1(n15493), .IN2(n15494), .QN(n15491) );
  NOR2X0 U15823 ( .IN1(n15008), .IN2(n15495), .QN(n15494) );
  INVX0 U15824 ( .INP(n3891), .ZN(n15495) );
  NOR2X0 U15825 ( .IN1(n3891), .IN2(n15496), .QN(n15493) );
  NAND2X0 U15826 ( .IN1(n10937), .IN2(g5563), .QN(n15496) );
  NAND2X0 U15827 ( .IN1(n15497), .IN2(n15498), .QN(g30483) );
  NAND2X0 U15828 ( .IN1(test_so6), .IN2(n11080), .QN(n15498) );
  NOR2X0 U15829 ( .IN1(n15499), .IN2(n15500), .QN(n15497) );
  NOR2X0 U15830 ( .IN1(n15008), .IN2(n15501), .QN(n15500) );
  INVX0 U15831 ( .INP(n3894), .ZN(n15501) );
  NOR2X0 U15832 ( .IN1(n3894), .IN2(n15502), .QN(n15499) );
  NAND2X0 U15833 ( .IN1(n10937), .IN2(g5555), .QN(n15502) );
  NAND2X0 U15834 ( .IN1(n15503), .IN2(n15504), .QN(g30482) );
  NAND2X0 U15835 ( .IN1(n11077), .IN2(g5551), .QN(n15504) );
  NOR2X0 U15836 ( .IN1(n15505), .IN2(n15506), .QN(n15503) );
  NOR2X0 U15837 ( .IN1(n15008), .IN2(n15507), .QN(n15506) );
  INVX0 U15838 ( .INP(n3896), .ZN(n15507) );
  NOR2X0 U15839 ( .IN1(n3896), .IN2(n15508), .QN(n15505) );
  NAND2X0 U15840 ( .IN1(n10937), .IN2(g5547), .QN(n15508) );
  NAND2X0 U15841 ( .IN1(n15509), .IN2(n15510), .QN(g30481) );
  NAND2X0 U15842 ( .IN1(n11077), .IN2(g5535), .QN(n15510) );
  NOR2X0 U15843 ( .IN1(n15511), .IN2(n15512), .QN(n15509) );
  NOR2X0 U15844 ( .IN1(n15008), .IN2(n15513), .QN(n15512) );
  INVX0 U15845 ( .INP(n3898), .ZN(n15513) );
  NOR2X0 U15846 ( .IN1(n3898), .IN2(n15514), .QN(n15511) );
  NAND2X0 U15847 ( .IN1(n10936), .IN2(g5543), .QN(n15514) );
  NOR2X0 U15848 ( .IN1(g5511), .IN2(n14291), .QN(g30480) );
  NAND2X0 U15849 ( .IN1(n15515), .IN2(n5647), .QN(n14291) );
  NOR2X0 U15850 ( .IN1(n11026), .IN2(n14295), .QN(n15515) );
  INVX0 U15851 ( .INP(n14279), .ZN(n14295) );
  NAND2X0 U15852 ( .IN1(n3833), .IN2(n13425), .QN(n14279) );
  NAND2X0 U15853 ( .IN1(n15516), .IN2(n15517), .QN(g30479) );
  NAND2X0 U15854 ( .IN1(n11077), .IN2(g5268), .QN(n15517) );
  NOR2X0 U15855 ( .IN1(n15518), .IN2(n15519), .QN(n15516) );
  NOR2X0 U15856 ( .IN1(n13429), .IN2(n15008), .QN(n15519) );
  NOR2X0 U15857 ( .IN1(n10303), .IN2(n15520), .QN(n15518) );
  NAND2X0 U15858 ( .IN1(n15521), .IN2(n15522), .QN(g30478) );
  NAND2X0 U15859 ( .IN1(n15523), .IN2(n3765), .QN(n15522) );
  NOR2X0 U15860 ( .IN1(n15524), .IN2(n15525), .QN(n15521) );
  NOR2X0 U15861 ( .IN1(n10462), .IN2(n10875), .QN(n15525) );
  NOR2X0 U15862 ( .IN1(n11027), .IN2(n15526), .QN(n15524) );
  NAND2X0 U15863 ( .IN1(n15527), .IN2(g5220), .QN(n15526) );
  INVX0 U15864 ( .INP(n15523), .ZN(n15527) );
  NOR2X0 U15865 ( .IN1(n3902), .IN2(n5650), .QN(n15523) );
  NAND2X0 U15866 ( .IN1(n15528), .IN2(n15529), .QN(g30477) );
  NAND2X0 U15867 ( .IN1(n14308), .IN2(n3765), .QN(n15529) );
  NOR2X0 U15868 ( .IN1(n15530), .IN2(n15531), .QN(n15528) );
  NOR2X0 U15869 ( .IN1(n10360), .IN2(n10875), .QN(n15531) );
  NOR2X0 U15870 ( .IN1(n11025), .IN2(n15532), .QN(n15530) );
  INVX0 U15871 ( .INP(n15533), .ZN(n15532) );
  NOR2X0 U15872 ( .IN1(n14308), .IN2(n10464), .QN(n15533) );
  NOR2X0 U15873 ( .IN1(n3904), .IN2(n5650), .QN(n14308) );
  NAND2X0 U15874 ( .IN1(n15534), .IN2(n15535), .QN(g30476) );
  NAND2X0 U15875 ( .IN1(n15536), .IN2(n3765), .QN(n15535) );
  NOR2X0 U15876 ( .IN1(n15537), .IN2(n15538), .QN(n15534) );
  NOR2X0 U15877 ( .IN1(n10304), .IN2(n10875), .QN(n15538) );
  NOR2X0 U15878 ( .IN1(n11025), .IN2(n15539), .QN(n15537) );
  NAND2X0 U15879 ( .IN1(n15540), .IN2(g5204), .QN(n15539) );
  INVX0 U15880 ( .INP(n15536), .ZN(n15540) );
  NOR2X0 U15881 ( .IN1(n3907), .IN2(n5650), .QN(n15536) );
  NAND2X0 U15882 ( .IN1(n15541), .IN2(n15542), .QN(g30475) );
  NAND2X0 U15883 ( .IN1(n3908), .IN2(n15543), .QN(n15542) );
  NOR2X0 U15884 ( .IN1(n15544), .IN2(n15545), .QN(n15541) );
  NOR2X0 U15885 ( .IN1(n11025), .IN2(n15546), .QN(n15545) );
  NAND2X0 U15886 ( .IN1(n15547), .IN2(g5268), .QN(n15546) );
  NAND2X0 U15887 ( .IN1(n15548), .IN2(n15543), .QN(n15547) );
  NOR2X0 U15888 ( .IN1(n10337), .IN2(n10875), .QN(n15544) );
  NAND2X0 U15889 ( .IN1(n15549), .IN2(n15550), .QN(g30474) );
  NAND2X0 U15890 ( .IN1(n3908), .IN2(n14307), .QN(n15550) );
  NOR2X0 U15891 ( .IN1(n15551), .IN2(n15552), .QN(n15549) );
  NOR2X0 U15892 ( .IN1(n11025), .IN2(n15553), .QN(n15552) );
  NAND2X0 U15893 ( .IN1(n15554), .IN2(g5264), .QN(n15553) );
  NAND2X0 U15894 ( .IN1(n15548), .IN2(n14307), .QN(n15554) );
  NOR2X0 U15895 ( .IN1(n10460), .IN2(n10876), .QN(n15551) );
  NAND2X0 U15896 ( .IN1(n15555), .IN2(n15556), .QN(g30473) );
  NAND2X0 U15897 ( .IN1(n3908), .IN2(n15557), .QN(n15556) );
  NOR2X0 U15898 ( .IN1(n15558), .IN2(n15559), .QN(n15555) );
  NOR2X0 U15899 ( .IN1(n11028), .IN2(n15560), .QN(n15559) );
  NAND2X0 U15900 ( .IN1(n15561), .IN2(g5260), .QN(n15560) );
  NAND2X0 U15901 ( .IN1(n15548), .IN2(n15557), .QN(n15561) );
  NOR2X0 U15902 ( .IN1(n10375), .IN2(n10876), .QN(n15558) );
  NAND2X0 U15903 ( .IN1(n15562), .IN2(n15563), .QN(g30472) );
  NAND2X0 U15904 ( .IN1(n3908), .IN2(n15564), .QN(n15563) );
  NOR2X0 U15905 ( .IN1(n15565), .IN2(n15566), .QN(n15562) );
  NOR2X0 U15906 ( .IN1(n11042), .IN2(n15567), .QN(n15566) );
  NAND2X0 U15907 ( .IN1(n15568), .IN2(g5256), .QN(n15567) );
  NAND2X0 U15908 ( .IN1(n15548), .IN2(n15564), .QN(n15568) );
  INVX0 U15909 ( .INP(n3444), .ZN(n15548) );
  NAND2X0 U15910 ( .IN1(g5164), .IN2(g5170), .QN(n3444) );
  NOR2X0 U15911 ( .IN1(n10432), .IN2(n10876), .QN(n15565) );
  NAND2X0 U15912 ( .IN1(n15569), .IN2(n15570), .QN(g30471) );
  NAND2X0 U15913 ( .IN1(n3914), .IN2(n15543), .QN(n15570) );
  NOR2X0 U15914 ( .IN1(n15571), .IN2(n15572), .QN(n15569) );
  NOR2X0 U15915 ( .IN1(n11042), .IN2(n15573), .QN(n15572) );
  NAND2X0 U15916 ( .IN1(n15574), .IN2(g5252), .QN(n15573) );
  NAND2X0 U15917 ( .IN1(n15543), .IN2(n14325), .QN(n15574) );
  NOR2X0 U15918 ( .IN1(n10338), .IN2(n10876), .QN(n15571) );
  NAND2X0 U15919 ( .IN1(n15575), .IN2(n15576), .QN(g30470) );
  NAND2X0 U15920 ( .IN1(n3914), .IN2(n14307), .QN(n15576) );
  NOR2X0 U15921 ( .IN1(n15577), .IN2(n15578), .QN(n15575) );
  NOR2X0 U15922 ( .IN1(n11042), .IN2(n15579), .QN(n15578) );
  NAND2X0 U15923 ( .IN1(n15580), .IN2(g5248), .QN(n15579) );
  NAND2X0 U15924 ( .IN1(n14307), .IN2(n14325), .QN(n15580) );
  NOR2X0 U15925 ( .IN1(n10411), .IN2(n10876), .QN(n15577) );
  NAND2X0 U15926 ( .IN1(n15581), .IN2(n15582), .QN(g30469) );
  NAND2X0 U15927 ( .IN1(n3914), .IN2(n15557), .QN(n15582) );
  NOR2X0 U15928 ( .IN1(n15583), .IN2(n15584), .QN(n15581) );
  NOR2X0 U15929 ( .IN1(n11042), .IN2(n15585), .QN(n15584) );
  NAND2X0 U15930 ( .IN1(n15586), .IN2(g5244), .QN(n15585) );
  NAND2X0 U15931 ( .IN1(n15557), .IN2(n14325), .QN(n15586) );
  NOR2X0 U15932 ( .IN1(n10906), .IN2(n10689), .QN(n15583) );
  NAND2X0 U15933 ( .IN1(n15587), .IN2(n15588), .QN(g30468) );
  NAND2X0 U15934 ( .IN1(n3914), .IN2(n15564), .QN(n15588) );
  NOR2X0 U15935 ( .IN1(n15589), .IN2(n15590), .QN(n15587) );
  NOR2X0 U15936 ( .IN1(n11042), .IN2(n15591), .QN(n15590) );
  NAND2X0 U15937 ( .IN1(n15592), .IN2(g5240), .QN(n15591) );
  NAND2X0 U15938 ( .IN1(n15564), .IN2(n14325), .QN(n15592) );
  INVX0 U15939 ( .INP(n792), .ZN(n14325) );
  NAND2X0 U15940 ( .IN1(n5570), .IN2(g5170), .QN(n792) );
  NOR2X0 U15941 ( .IN1(n10305), .IN2(n10877), .QN(n15589) );
  NAND2X0 U15942 ( .IN1(n15593), .IN2(n15594), .QN(g30467) );
  NAND2X0 U15943 ( .IN1(n3919), .IN2(n15543), .QN(n15594) );
  NOR2X0 U15944 ( .IN1(n15595), .IN2(n15596), .QN(n15593) );
  NOR2X0 U15945 ( .IN1(n11042), .IN2(n15597), .QN(n15596) );
  NAND2X0 U15946 ( .IN1(n15598), .IN2(g5236), .QN(n15597) );
  NAND2X0 U15947 ( .IN1(n15599), .IN2(n15543), .QN(n15598) );
  NOR2X0 U15948 ( .IN1(n10412), .IN2(n10877), .QN(n15595) );
  NAND2X0 U15949 ( .IN1(n15600), .IN2(n15601), .QN(g30466) );
  NAND2X0 U15950 ( .IN1(n3919), .IN2(n14307), .QN(n15601) );
  NOR2X0 U15951 ( .IN1(n15602), .IN2(n15603), .QN(n15600) );
  NOR2X0 U15952 ( .IN1(n11042), .IN2(n15604), .QN(n15603) );
  NAND2X0 U15953 ( .IN1(n15605), .IN2(g5232), .QN(n15604) );
  NAND2X0 U15954 ( .IN1(n15599), .IN2(n14307), .QN(n15605) );
  INVX0 U15955 ( .INP(n3902), .ZN(n14307) );
  NAND2X0 U15956 ( .IN1(n5384), .IN2(g5188), .QN(n3902) );
  NOR2X0 U15957 ( .IN1(n10406), .IN2(n10877), .QN(n15602) );
  NAND2X0 U15958 ( .IN1(n15606), .IN2(n15607), .QN(g30465) );
  NAND2X0 U15959 ( .IN1(n3919), .IN2(n15557), .QN(n15607) );
  NOR2X0 U15960 ( .IN1(n15608), .IN2(n15609), .QN(n15606) );
  NOR2X0 U15961 ( .IN1(n11042), .IN2(n15610), .QN(n15609) );
  NAND2X0 U15962 ( .IN1(test_so82), .IN2(n15611), .QN(n15610) );
  NAND2X0 U15963 ( .IN1(n15599), .IN2(n15557), .QN(n15611) );
  INVX0 U15964 ( .INP(n3904), .ZN(n15557) );
  NAND2X0 U15965 ( .IN1(n5567), .IN2(g5180), .QN(n3904) );
  NOR2X0 U15966 ( .IN1(n10306), .IN2(n10877), .QN(n15608) );
  NAND2X0 U15967 ( .IN1(n15612), .IN2(n15613), .QN(g30464) );
  NAND2X0 U15968 ( .IN1(n3919), .IN2(n15564), .QN(n15613) );
  NOR2X0 U15969 ( .IN1(n15614), .IN2(n15615), .QN(n15612) );
  NOR2X0 U15970 ( .IN1(n11042), .IN2(n15616), .QN(n15615) );
  NAND2X0 U15971 ( .IN1(n15617), .IN2(g5224), .QN(n15616) );
  NAND2X0 U15972 ( .IN1(n15599), .IN2(n15564), .QN(n15617) );
  INVX0 U15973 ( .INP(n3907), .ZN(n15564) );
  NAND2X0 U15974 ( .IN1(n5567), .IN2(n5384), .QN(n3907) );
  INVX0 U15975 ( .INP(n3447), .ZN(n15599) );
  NAND2X0 U15976 ( .IN1(n10586), .IN2(g5164), .QN(n3447) );
  NOR2X0 U15977 ( .IN1(n10443), .IN2(n10877), .QN(n15614) );
  NAND2X0 U15978 ( .IN1(n15618), .IN2(n15619), .QN(g30463) );
  NAND2X0 U15979 ( .IN1(n11077), .IN2(g5220), .QN(n15619) );
  NOR2X0 U15980 ( .IN1(n15620), .IN2(n15621), .QN(n15618) );
  NOR2X0 U15981 ( .IN1(n15008), .IN2(n15622), .QN(n15621) );
  INVX0 U15982 ( .INP(n3924), .ZN(n15622) );
  NOR2X0 U15983 ( .IN1(n3924), .IN2(n15623), .QN(n15620) );
  NAND2X0 U15984 ( .IN1(n10936), .IN2(g5216), .QN(n15623) );
  NAND2X0 U15985 ( .IN1(n15624), .IN2(n15625), .QN(g30462) );
  NAND2X0 U15986 ( .IN1(n11077), .IN2(g5212), .QN(n15625) );
  NOR2X0 U15987 ( .IN1(n15626), .IN2(n15627), .QN(n15624) );
  NOR2X0 U15988 ( .IN1(n15008), .IN2(n15628), .QN(n15627) );
  INVX0 U15989 ( .INP(n3927), .ZN(n15628) );
  NOR2X0 U15990 ( .IN1(n3927), .IN2(n15629), .QN(n15626) );
  NAND2X0 U15991 ( .IN1(n10935), .IN2(g5208), .QN(n15629) );
  NAND2X0 U15992 ( .IN1(n15630), .IN2(n15631), .QN(g30461) );
  NAND2X0 U15993 ( .IN1(n11077), .IN2(g5204), .QN(n15631) );
  NOR2X0 U15994 ( .IN1(n15632), .IN2(n15633), .QN(n15630) );
  NOR2X0 U15995 ( .IN1(n15008), .IN2(n15634), .QN(n15633) );
  INVX0 U15996 ( .INP(n3929), .ZN(n15634) );
  NOR2X0 U15997 ( .IN1(n3929), .IN2(n15635), .QN(n15632) );
  NAND2X0 U15998 ( .IN1(n10936), .IN2(g5200), .QN(n15635) );
  NAND2X0 U15999 ( .IN1(n15636), .IN2(n15637), .QN(g30460) );
  NAND2X0 U16000 ( .IN1(n11077), .IN2(g5188), .QN(n15637) );
  NOR2X0 U16001 ( .IN1(n15638), .IN2(n15639), .QN(n15636) );
  NOR2X0 U16002 ( .IN1(n15008), .IN2(n15640), .QN(n15639) );
  INVX0 U16003 ( .INP(n3931), .ZN(n15640) );
  NOR2X0 U16004 ( .IN1(n3931), .IN2(n15641), .QN(n15638) );
  NAND2X0 U16005 ( .IN1(n10934), .IN2(g5196), .QN(n15641) );
  NOR2X0 U16006 ( .IN1(g5164), .IN2(n14316), .QN(g30459) );
  NAND2X0 U16007 ( .IN1(n15642), .IN2(n5650), .QN(n14316) );
  NOR2X0 U16008 ( .IN1(n11042), .IN2(n14320), .QN(n15642) );
  INVX0 U16009 ( .INP(n14304), .ZN(n14320) );
  NAND2X0 U16010 ( .IN1(n3833), .IN2(n15132), .QN(n14304) );
  NAND2X0 U16011 ( .IN1(n15643), .IN2(n10955), .QN(g30458) );
  NOR2X0 U16012 ( .IN1(n15644), .IN2(n15645), .QN(n15643) );
  NOR2X0 U16013 ( .IN1(n5846), .IN2(n15646), .QN(n15645) );
  INVX0 U16014 ( .INP(n15647), .ZN(n15644) );
  NAND2X0 U16015 ( .IN1(g113), .IN2(n15646), .QN(n15647) );
  NOR2X0 U16016 ( .IN1(g4459), .IN2(n10207), .QN(n15646) );
  NAND2X0 U16017 ( .IN1(n15648), .IN2(n15649), .QN(g30457) );
  NAND2X0 U16018 ( .IN1(n11077), .IN2(g4122), .QN(n15649) );
  NAND2X0 U16019 ( .IN1(n15650), .IN2(n10955), .QN(n15648) );
  NAND2X0 U16020 ( .IN1(n15651), .IN2(n15652), .QN(n15650) );
  NAND2X0 U16021 ( .IN1(n15653), .IN2(n5981), .QN(n15652) );
  XNOR2X1 U16022 ( .IN1(g126), .IN2(n15654), .Q(n15653) );
  NAND2X0 U16023 ( .IN1(n15655), .IN2(n5983), .QN(n15651) );
  XNOR2X1 U16024 ( .IN1(g115), .IN2(n15656), .Q(n15655) );
  NAND2X0 U16025 ( .IN1(n15657), .IN2(n15658), .QN(g30456) );
  NAND2X0 U16026 ( .IN1(n11077), .IN2(g4087), .QN(n15658) );
  NOR2X0 U16027 ( .IN1(n15659), .IN2(n15660), .QN(n15657) );
  NOR2X0 U16028 ( .IN1(n15661), .IN2(n15662), .QN(n15660) );
  INVX0 U16029 ( .INP(n3941), .ZN(n15662) );
  NOR2X0 U16030 ( .IN1(n15663), .IN2(n15664), .QN(n15659) );
  NAND2X0 U16031 ( .IN1(n14910), .IN2(g4169), .QN(n15664) );
  NAND2X0 U16032 ( .IN1(n15665), .IN2(n15666), .QN(g30455) );
  NAND2X0 U16033 ( .IN1(n11077), .IN2(g3961), .QN(n15666) );
  NOR2X0 U16034 ( .IN1(n15667), .IN2(n15668), .QN(n15665) );
  NOR2X0 U16035 ( .IN1(n15008), .IN2(n13445), .QN(n15668) );
  NOR2X0 U16036 ( .IN1(n10309), .IN2(n15669), .QN(n15667) );
  NAND2X0 U16037 ( .IN1(n15670), .IN2(n15671), .QN(g30454) );
  NAND2X0 U16038 ( .IN1(n15672), .IN2(n3765), .QN(n15671) );
  NOR2X0 U16039 ( .IN1(n15673), .IN2(n15674), .QN(n15670) );
  NOR2X0 U16040 ( .IN1(n10476), .IN2(n10879), .QN(n15674) );
  INVX0 U16041 ( .INP(n15675), .ZN(n15673) );
  NAND2X0 U16042 ( .IN1(n10935), .IN2(n15676), .QN(n15675) );
  NOR2X0 U16043 ( .IN1(n15672), .IN2(n10506), .QN(n15676) );
  NOR2X0 U16044 ( .IN1(n10647), .IN2(n3945), .QN(n15672) );
  NAND2X0 U16045 ( .IN1(n15677), .IN2(n15678), .QN(g30453) );
  NAND2X0 U16046 ( .IN1(n14379), .IN2(n3765), .QN(n15678) );
  INVX0 U16047 ( .INP(n15679), .ZN(n14379) );
  NOR2X0 U16048 ( .IN1(n15680), .IN2(n15681), .QN(n15677) );
  NOR2X0 U16049 ( .IN1(n10366), .IN2(n10879), .QN(n15681) );
  NOR2X0 U16050 ( .IN1(n11041), .IN2(n15682), .QN(n15680) );
  NAND2X0 U16051 ( .IN1(n15679), .IN2(g3905), .QN(n15682) );
  NAND2X0 U16052 ( .IN1(test_so33), .IN2(n15683), .QN(n15679) );
  NAND2X0 U16053 ( .IN1(n15684), .IN2(n15685), .QN(g30452) );
  NAND2X0 U16054 ( .IN1(n15686), .IN2(n3765), .QN(n15685) );
  INVX0 U16055 ( .INP(n15687), .ZN(n15684) );
  NAND2X0 U16056 ( .IN1(n15688), .IN2(n15689), .QN(n15687) );
  NAND2X0 U16057 ( .IN1(n11077), .IN2(test_so65), .QN(n15689) );
  NAND2X0 U16058 ( .IN1(n10933), .IN2(n15690), .QN(n15688) );
  NOR2X0 U16059 ( .IN1(n15686), .IN2(n10448), .QN(n15690) );
  NOR2X0 U16060 ( .IN1(n10647), .IN2(n3950), .QN(n15686) );
  NAND2X0 U16061 ( .IN1(n15691), .IN2(n15692), .QN(g30451) );
  NAND2X0 U16062 ( .IN1(n3951), .IN2(n15693), .QN(n15692) );
  NOR2X0 U16063 ( .IN1(n15694), .IN2(n15695), .QN(n15691) );
  NOR2X0 U16064 ( .IN1(n11041), .IN2(n15696), .QN(n15695) );
  NAND2X0 U16065 ( .IN1(n15697), .IN2(g3961), .QN(n15696) );
  NAND2X0 U16066 ( .IN1(n15698), .IN2(n15693), .QN(n15697) );
  NOR2X0 U16067 ( .IN1(n10346), .IN2(n10879), .QN(n15694) );
  NAND2X0 U16068 ( .IN1(n15699), .IN2(n15700), .QN(g30450) );
  NAND2X0 U16069 ( .IN1(n3951), .IN2(n14378), .QN(n15700) );
  NOR2X0 U16070 ( .IN1(n15701), .IN2(n15702), .QN(n15699) );
  NOR2X0 U16071 ( .IN1(n11041), .IN2(n15703), .QN(n15702) );
  NAND2X0 U16072 ( .IN1(n15704), .IN2(g3957), .QN(n15703) );
  NAND2X0 U16073 ( .IN1(n15698), .IN2(n14378), .QN(n15704) );
  NOR2X0 U16074 ( .IN1(n10474), .IN2(n10880), .QN(n15701) );
  NAND2X0 U16075 ( .IN1(n15705), .IN2(n15706), .QN(g30449) );
  NAND2X0 U16076 ( .IN1(n3951), .IN2(n15683), .QN(n15706) );
  NOR2X0 U16077 ( .IN1(n15707), .IN2(n15708), .QN(n15705) );
  NOR2X0 U16078 ( .IN1(n11041), .IN2(n15709), .QN(n15708) );
  NAND2X0 U16079 ( .IN1(n15710), .IN2(g3953), .QN(n15709) );
  NAND2X0 U16080 ( .IN1(n15698), .IN2(n15683), .QN(n15710) );
  NOR2X0 U16081 ( .IN1(n10380), .IN2(n10880), .QN(n15707) );
  NAND2X0 U16082 ( .IN1(n15711), .IN2(n15712), .QN(g30448) );
  NAND2X0 U16083 ( .IN1(n3951), .IN2(n15713), .QN(n15712) );
  NOR2X0 U16084 ( .IN1(n15714), .IN2(n15715), .QN(n15711) );
  NOR2X0 U16085 ( .IN1(n11041), .IN2(n15716), .QN(n15715) );
  NAND2X0 U16086 ( .IN1(test_so65), .IN2(n15717), .QN(n15716) );
  NAND2X0 U16087 ( .IN1(n15698), .IN2(n15713), .QN(n15717) );
  INVX0 U16088 ( .INP(n3479), .ZN(n15698) );
  NAND2X0 U16089 ( .IN1(g3857), .IN2(g3863), .QN(n3479) );
  NOR2X0 U16090 ( .IN1(n10435), .IN2(n10880), .QN(n15714) );
  NAND2X0 U16091 ( .IN1(n15718), .IN2(n15719), .QN(g30447) );
  NAND2X0 U16092 ( .IN1(n3957), .IN2(n15693), .QN(n15719) );
  NOR2X0 U16093 ( .IN1(n15720), .IN2(n15721), .QN(n15718) );
  NOR2X0 U16094 ( .IN1(n11041), .IN2(n15722), .QN(n15721) );
  NAND2X0 U16095 ( .IN1(n15723), .IN2(g3945), .QN(n15722) );
  NAND2X0 U16096 ( .IN1(n14395), .IN2(n15693), .QN(n15723) );
  NOR2X0 U16097 ( .IN1(n10347), .IN2(n10880), .QN(n15720) );
  NAND2X0 U16098 ( .IN1(n15724), .IN2(n15725), .QN(g30446) );
  NAND2X0 U16099 ( .IN1(n3957), .IN2(n14378), .QN(n15725) );
  NOR2X0 U16100 ( .IN1(n15726), .IN2(n15727), .QN(n15724) );
  NOR2X0 U16101 ( .IN1(n11041), .IN2(n15728), .QN(n15727) );
  NAND2X0 U16102 ( .IN1(n15729), .IN2(g3941), .QN(n15728) );
  NAND2X0 U16103 ( .IN1(n14395), .IN2(n14378), .QN(n15729) );
  NOR2X0 U16104 ( .IN1(n10420), .IN2(n10880), .QN(n15726) );
  NAND2X0 U16105 ( .IN1(n15730), .IN2(n15731), .QN(g30445) );
  NAND2X0 U16106 ( .IN1(n3957), .IN2(n15683), .QN(n15731) );
  NOR2X0 U16107 ( .IN1(n15732), .IN2(n15733), .QN(n15730) );
  NOR2X0 U16108 ( .IN1(n11041), .IN2(n15734), .QN(n15733) );
  NAND2X0 U16109 ( .IN1(n15735), .IN2(g3937), .QN(n15734) );
  NAND2X0 U16110 ( .IN1(n14395), .IN2(n15683), .QN(n15735) );
  NOR2X0 U16111 ( .IN1(n10330), .IN2(n10881), .QN(n15732) );
  NAND2X0 U16112 ( .IN1(n15736), .IN2(n15737), .QN(g30444) );
  NAND2X0 U16113 ( .IN1(n3957), .IN2(n15713), .QN(n15737) );
  NOR2X0 U16114 ( .IN1(n15738), .IN2(n15739), .QN(n15736) );
  NOR2X0 U16115 ( .IN1(n11041), .IN2(n15740), .QN(n15739) );
  NAND2X0 U16116 ( .IN1(n15741), .IN2(g3933), .QN(n15740) );
  NAND2X0 U16117 ( .IN1(n14395), .IN2(n15713), .QN(n15741) );
  INVX0 U16118 ( .INP(n3481), .ZN(n14395) );
  NAND2X0 U16119 ( .IN1(n5572), .IN2(g3863), .QN(n3481) );
  NOR2X0 U16120 ( .IN1(n10310), .IN2(n10881), .QN(n15738) );
  NAND2X0 U16121 ( .IN1(n15742), .IN2(n15743), .QN(g30443) );
  NAND2X0 U16122 ( .IN1(n3962), .IN2(n15693), .QN(n15743) );
  NOR2X0 U16123 ( .IN1(n15744), .IN2(n15745), .QN(n15742) );
  NOR2X0 U16124 ( .IN1(n11041), .IN2(n15746), .QN(n15745) );
  NAND2X0 U16125 ( .IN1(n15747), .IN2(g3929), .QN(n15746) );
  NAND2X0 U16126 ( .IN1(n15748), .IN2(n15693), .QN(n15747) );
  NOR2X0 U16127 ( .IN1(n10421), .IN2(n10881), .QN(n15744) );
  NAND2X0 U16128 ( .IN1(n15749), .IN2(n15750), .QN(g30442) );
  NAND2X0 U16129 ( .IN1(n3962), .IN2(n14378), .QN(n15750) );
  NOR2X0 U16130 ( .IN1(n15751), .IN2(n15752), .QN(n15749) );
  NOR2X0 U16131 ( .IN1(n11041), .IN2(n15753), .QN(n15752) );
  NAND2X0 U16132 ( .IN1(n15754), .IN2(g3925), .QN(n15753) );
  NAND2X0 U16133 ( .IN1(n15748), .IN2(n14378), .QN(n15754) );
  INVX0 U16134 ( .INP(n3945), .ZN(n14378) );
  NAND2X0 U16135 ( .IN1(n5387), .IN2(g3881), .QN(n3945) );
  NOR2X0 U16136 ( .IN1(n10508), .IN2(n10881), .QN(n15751) );
  NAND2X0 U16137 ( .IN1(n15755), .IN2(n15756), .QN(g30441) );
  NAND2X0 U16138 ( .IN1(n3962), .IN2(n15683), .QN(n15756) );
  NOR2X0 U16139 ( .IN1(n15757), .IN2(n15758), .QN(n15755) );
  NOR2X0 U16140 ( .IN1(n11041), .IN2(n15759), .QN(n15758) );
  NAND2X0 U16141 ( .IN1(n15760), .IN2(g3921), .QN(n15759) );
  NAND2X0 U16142 ( .IN1(n15748), .IN2(n15683), .QN(n15760) );
  INVX0 U16143 ( .INP(n3947), .ZN(n15683) );
  NAND2X0 U16144 ( .IN1(n5564), .IN2(g3873), .QN(n3947) );
  NOR2X0 U16145 ( .IN1(n10311), .IN2(n10881), .QN(n15757) );
  NAND2X0 U16146 ( .IN1(n15761), .IN2(n15762), .QN(g30440) );
  NAND2X0 U16147 ( .IN1(n3962), .IN2(n15713), .QN(n15762) );
  NOR2X0 U16148 ( .IN1(n15763), .IN2(n15764), .QN(n15761) );
  NOR2X0 U16149 ( .IN1(n11041), .IN2(n15765), .QN(n15764) );
  NAND2X0 U16150 ( .IN1(n15766), .IN2(g3917), .QN(n15765) );
  NAND2X0 U16151 ( .IN1(n15748), .IN2(n15713), .QN(n15766) );
  INVX0 U16152 ( .INP(n3950), .ZN(n15713) );
  NAND2X0 U16153 ( .IN1(n5564), .IN2(n5387), .QN(n3950) );
  INVX0 U16154 ( .INP(n3482), .ZN(n15748) );
  NAND2X0 U16155 ( .IN1(n10591), .IN2(g3857), .QN(n3482) );
  NOR2X0 U16156 ( .IN1(n10908), .IN2(n10686), .QN(n15763) );
  NAND2X0 U16157 ( .IN1(n15767), .IN2(n15768), .QN(g30439) );
  NAND2X0 U16158 ( .IN1(n11077), .IN2(g3913), .QN(n15768) );
  NOR2X0 U16159 ( .IN1(n15769), .IN2(n15770), .QN(n15767) );
  NOR2X0 U16160 ( .IN1(n15008), .IN2(n15771), .QN(n15770) );
  INVX0 U16161 ( .INP(n3967), .ZN(n15771) );
  NOR2X0 U16162 ( .IN1(n3967), .IN2(n15772), .QN(n15769) );
  NAND2X0 U16163 ( .IN1(n10934), .IN2(g3909), .QN(n15772) );
  NAND2X0 U16164 ( .IN1(n15773), .IN2(n15774), .QN(g30438) );
  NAND2X0 U16165 ( .IN1(n11076), .IN2(g3905), .QN(n15774) );
  NOR2X0 U16166 ( .IN1(n15775), .IN2(n15776), .QN(n15773) );
  NOR2X0 U16167 ( .IN1(n15008), .IN2(n15777), .QN(n15776) );
  INVX0 U16168 ( .INP(n3970), .ZN(n15777) );
  NOR2X0 U16169 ( .IN1(n3970), .IN2(n15778), .QN(n15775) );
  NAND2X0 U16170 ( .IN1(n10933), .IN2(g3901), .QN(n15778) );
  NAND2X0 U16171 ( .IN1(n15779), .IN2(n15780), .QN(g30437) );
  NAND2X0 U16172 ( .IN1(n11076), .IN2(g3897), .QN(n15780) );
  NOR2X0 U16173 ( .IN1(n15781), .IN2(n15782), .QN(n15779) );
  NOR2X0 U16174 ( .IN1(n15008), .IN2(n15783), .QN(n15782) );
  INVX0 U16175 ( .INP(n3972), .ZN(n15783) );
  NOR2X0 U16176 ( .IN1(n3972), .IN2(n15784), .QN(n15781) );
  NAND2X0 U16177 ( .IN1(n10933), .IN2(g3893), .QN(n15784) );
  NAND2X0 U16178 ( .IN1(n15785), .IN2(n15786), .QN(g30436) );
  NAND2X0 U16179 ( .IN1(n11076), .IN2(g3881), .QN(n15786) );
  NOR2X0 U16180 ( .IN1(n15787), .IN2(n15788), .QN(n15785) );
  NOR2X0 U16181 ( .IN1(n15008), .IN2(n15789), .QN(n15788) );
  INVX0 U16182 ( .INP(n3974), .ZN(n15789) );
  NOR2X0 U16183 ( .IN1(n3974), .IN2(n15790), .QN(n15787) );
  NAND2X0 U16184 ( .IN1(test_so24), .IN2(n10955), .QN(n15790) );
  NOR2X0 U16185 ( .IN1(g3857), .IN2(n14387), .QN(g30435) );
  NAND2X0 U16186 ( .IN1(n15791), .IN2(n14375), .QN(n14387) );
  NAND2X0 U16187 ( .IN1(n15260), .IN2(n3799), .QN(n14375) );
  NOR2X0 U16188 ( .IN1(n5480), .IN2(n5340), .QN(n15260) );
  NOR2X0 U16189 ( .IN1(test_so33), .IN2(n11023), .QN(n15791) );
  NAND2X0 U16190 ( .IN1(n15792), .IN2(n15793), .QN(g30434) );
  NAND2X0 U16191 ( .IN1(n11076), .IN2(g3610), .QN(n15793) );
  NOR2X0 U16192 ( .IN1(n15794), .IN2(n15795), .QN(n15792) );
  NOR2X0 U16193 ( .IN1(n15008), .IN2(n13444), .QN(n15795) );
  NOR2X0 U16194 ( .IN1(n10295), .IN2(n15796), .QN(n15794) );
  NAND2X0 U16195 ( .IN1(n15797), .IN2(n15798), .QN(g30433) );
  NAND2X0 U16196 ( .IN1(n15799), .IN2(n3765), .QN(n15798) );
  NOR2X0 U16197 ( .IN1(n15800), .IN2(n15801), .QN(n15797) );
  NOR2X0 U16198 ( .IN1(n10486), .IN2(n10839), .QN(n15801) );
  NOR2X0 U16199 ( .IN1(n11040), .IN2(n15802), .QN(n15800) );
  NAND2X0 U16200 ( .IN1(n15803), .IN2(g3562), .QN(n15802) );
  INVX0 U16201 ( .INP(n15799), .ZN(n15803) );
  NOR2X0 U16202 ( .IN1(n3978), .IN2(n5645), .QN(n15799) );
  NAND2X0 U16203 ( .IN1(n15804), .IN2(n15805), .QN(g30432) );
  NAND2X0 U16204 ( .IN1(n14403), .IN2(n3765), .QN(n15805) );
  NOR2X0 U16205 ( .IN1(n15806), .IN2(n15807), .QN(n15804) );
  NOR2X0 U16206 ( .IN1(n10905), .IN2(n10664), .QN(n15807) );
  NOR2X0 U16207 ( .IN1(n11040), .IN2(n15808), .QN(n15806) );
  INVX0 U16208 ( .INP(n15809), .ZN(n15808) );
  NOR2X0 U16209 ( .IN1(n14403), .IN2(n10488), .QN(n15809) );
  NOR2X0 U16210 ( .IN1(n3980), .IN2(n5645), .QN(n14403) );
  NAND2X0 U16211 ( .IN1(n15810), .IN2(n15811), .QN(g30431) );
  NAND2X0 U16212 ( .IN1(n15812), .IN2(n3765), .QN(n15811) );
  NOR2X0 U16213 ( .IN1(n15813), .IN2(n15814), .QN(n15810) );
  NOR2X0 U16214 ( .IN1(n10296), .IN2(n10839), .QN(n15814) );
  NOR2X0 U16215 ( .IN1(n11040), .IN2(n15815), .QN(n15813) );
  NAND2X0 U16216 ( .IN1(n15816), .IN2(g3546), .QN(n15815) );
  INVX0 U16217 ( .INP(n15812), .ZN(n15816) );
  NOR2X0 U16218 ( .IN1(n3983), .IN2(n5645), .QN(n15812) );
  NAND2X0 U16219 ( .IN1(n15817), .IN2(n15818), .QN(g30430) );
  NAND2X0 U16220 ( .IN1(n3984), .IN2(n15819), .QN(n15818) );
  NOR2X0 U16221 ( .IN1(n15820), .IN2(n15821), .QN(n15817) );
  NOR2X0 U16222 ( .IN1(n11040), .IN2(n15822), .QN(n15821) );
  NAND2X0 U16223 ( .IN1(n15823), .IN2(g3610), .QN(n15822) );
  NAND2X0 U16224 ( .IN1(n15824), .IN2(n15819), .QN(n15823) );
  NOR2X0 U16225 ( .IN1(n10352), .IN2(n10840), .QN(n15820) );
  NAND2X0 U16226 ( .IN1(n15825), .IN2(n15826), .QN(g30429) );
  NAND2X0 U16227 ( .IN1(n3984), .IN2(n14402), .QN(n15826) );
  NOR2X0 U16228 ( .IN1(n15827), .IN2(n15828), .QN(n15825) );
  NOR2X0 U16229 ( .IN1(n11040), .IN2(n15829), .QN(n15828) );
  NAND2X0 U16230 ( .IN1(n15830), .IN2(g3606), .QN(n15829) );
  NAND2X0 U16231 ( .IN1(n15824), .IN2(n14402), .QN(n15830) );
  NOR2X0 U16232 ( .IN1(n10484), .IN2(n10840), .QN(n15827) );
  NAND2X0 U16233 ( .IN1(n15831), .IN2(n15832), .QN(g30428) );
  NAND2X0 U16234 ( .IN1(n3984), .IN2(n15833), .QN(n15832) );
  NOR2X0 U16235 ( .IN1(n15834), .IN2(n15835), .QN(n15831) );
  NOR2X0 U16236 ( .IN1(n11040), .IN2(n15836), .QN(n15835) );
  NAND2X0 U16237 ( .IN1(test_so43), .IN2(n15837), .QN(n15836) );
  NAND2X0 U16238 ( .IN1(n15824), .IN2(n15833), .QN(n15837) );
  NOR2X0 U16239 ( .IN1(n10384), .IN2(n10840), .QN(n15834) );
  NAND2X0 U16240 ( .IN1(n15838), .IN2(n15839), .QN(g30427) );
  NAND2X0 U16241 ( .IN1(n3984), .IN2(n15840), .QN(n15839) );
  NOR2X0 U16242 ( .IN1(n15841), .IN2(n15842), .QN(n15838) );
  NOR2X0 U16243 ( .IN1(n11040), .IN2(n15843), .QN(n15842) );
  NAND2X0 U16244 ( .IN1(n15844), .IN2(g3598), .QN(n15843) );
  NAND2X0 U16245 ( .IN1(n15824), .IN2(n15840), .QN(n15844) );
  INVX0 U16246 ( .INP(n3489), .ZN(n15824) );
  NAND2X0 U16247 ( .IN1(g3506), .IN2(g3512), .QN(n3489) );
  NOR2X0 U16248 ( .IN1(n10437), .IN2(n10840), .QN(n15841) );
  NAND2X0 U16249 ( .IN1(n15845), .IN2(n15846), .QN(g30426) );
  NAND2X0 U16250 ( .IN1(n3990), .IN2(n15819), .QN(n15846) );
  NOR2X0 U16251 ( .IN1(n15847), .IN2(n15848), .QN(n15845) );
  NOR2X0 U16252 ( .IN1(n11040), .IN2(n15849), .QN(n15848) );
  NAND2X0 U16253 ( .IN1(n15850), .IN2(g3594), .QN(n15849) );
  NAND2X0 U16254 ( .IN1(n14420), .IN2(n15819), .QN(n15850) );
  NOR2X0 U16255 ( .IN1(n10353), .IN2(n10840), .QN(n15847) );
  NAND2X0 U16256 ( .IN1(n15851), .IN2(n15852), .QN(g30425) );
  NAND2X0 U16257 ( .IN1(n3990), .IN2(n14402), .QN(n15852) );
  NOR2X0 U16258 ( .IN1(n15853), .IN2(n15854), .QN(n15851) );
  NOR2X0 U16259 ( .IN1(n11040), .IN2(n15855), .QN(n15854) );
  NAND2X0 U16260 ( .IN1(n15856), .IN2(g3590), .QN(n15855) );
  NAND2X0 U16261 ( .IN1(n14420), .IN2(n14402), .QN(n15856) );
  NOR2X0 U16262 ( .IN1(n10426), .IN2(n10841), .QN(n15853) );
  NAND2X0 U16263 ( .IN1(n15857), .IN2(n15858), .QN(g30424) );
  NAND2X0 U16264 ( .IN1(n3990), .IN2(n15833), .QN(n15858) );
  NOR2X0 U16265 ( .IN1(n15859), .IN2(n15860), .QN(n15857) );
  NOR2X0 U16266 ( .IN1(n11040), .IN2(n15861), .QN(n15860) );
  NAND2X0 U16267 ( .IN1(n15862), .IN2(g3586), .QN(n15861) );
  NAND2X0 U16268 ( .IN1(n14420), .IN2(n15833), .QN(n15862) );
  NOR2X0 U16269 ( .IN1(n10332), .IN2(n10841), .QN(n15859) );
  NAND2X0 U16270 ( .IN1(n15863), .IN2(n15864), .QN(g30423) );
  NAND2X0 U16271 ( .IN1(n3990), .IN2(n15840), .QN(n15864) );
  NOR2X0 U16272 ( .IN1(n15865), .IN2(n15866), .QN(n15863) );
  NOR2X0 U16273 ( .IN1(n11040), .IN2(n15867), .QN(n15866) );
  NAND2X0 U16274 ( .IN1(n15868), .IN2(g3582), .QN(n15867) );
  NAND2X0 U16275 ( .IN1(n14420), .IN2(n15840), .QN(n15868) );
  INVX0 U16276 ( .INP(n3491), .ZN(n14420) );
  NAND2X0 U16277 ( .IN1(n5576), .IN2(g3512), .QN(n3491) );
  NOR2X0 U16278 ( .IN1(n10297), .IN2(n10841), .QN(n15865) );
  NAND2X0 U16279 ( .IN1(n15869), .IN2(n15870), .QN(g30422) );
  NAND2X0 U16280 ( .IN1(n3995), .IN2(n15819), .QN(n15870) );
  NOR2X0 U16281 ( .IN1(n15871), .IN2(n15872), .QN(n15869) );
  NOR2X0 U16282 ( .IN1(n11040), .IN2(n15873), .QN(n15872) );
  NAND2X0 U16283 ( .IN1(n15874), .IN2(g3578), .QN(n15873) );
  NAND2X0 U16284 ( .IN1(n15875), .IN2(n15819), .QN(n15874) );
  NOR2X0 U16285 ( .IN1(n10427), .IN2(n10841), .QN(n15871) );
  NAND2X0 U16286 ( .IN1(n15876), .IN2(n15877), .QN(g30421) );
  NAND2X0 U16287 ( .IN1(n3995), .IN2(n14402), .QN(n15877) );
  NOR2X0 U16288 ( .IN1(n15878), .IN2(n15879), .QN(n15876) );
  NOR2X0 U16289 ( .IN1(n11040), .IN2(n15880), .QN(n15879) );
  NAND2X0 U16290 ( .IN1(n15881), .IN2(g3574), .QN(n15880) );
  NAND2X0 U16291 ( .IN1(n15875), .IN2(n14402), .QN(n15881) );
  INVX0 U16292 ( .INP(n3978), .ZN(n14402) );
  NAND2X0 U16293 ( .IN1(n5383), .IN2(g3530), .QN(n3978) );
  NOR2X0 U16294 ( .IN1(n10516), .IN2(n10841), .QN(n15878) );
  NAND2X0 U16295 ( .IN1(n15882), .IN2(n15883), .QN(g30420) );
  NAND2X0 U16296 ( .IN1(n3995), .IN2(n15833), .QN(n15883) );
  NOR2X0 U16297 ( .IN1(n15884), .IN2(n15885), .QN(n15882) );
  NOR2X0 U16298 ( .IN1(n11039), .IN2(n15886), .QN(n15885) );
  NAND2X0 U16299 ( .IN1(n15887), .IN2(g3570), .QN(n15886) );
  NAND2X0 U16300 ( .IN1(n15875), .IN2(n15833), .QN(n15887) );
  INVX0 U16301 ( .INP(n3980), .ZN(n15833) );
  NAND2X0 U16302 ( .IN1(n5569), .IN2(g3522), .QN(n3980) );
  NOR2X0 U16303 ( .IN1(n10298), .IN2(n10842), .QN(n15884) );
  NAND2X0 U16304 ( .IN1(n15888), .IN2(n15889), .QN(g30419) );
  NAND2X0 U16305 ( .IN1(n3995), .IN2(n15840), .QN(n15889) );
  NOR2X0 U16306 ( .IN1(n15890), .IN2(n15891), .QN(n15888) );
  NOR2X0 U16307 ( .IN1(n11039), .IN2(n15892), .QN(n15891) );
  NAND2X0 U16308 ( .IN1(n15893), .IN2(g3566), .QN(n15892) );
  NAND2X0 U16309 ( .IN1(n15875), .IN2(n15840), .QN(n15893) );
  INVX0 U16310 ( .INP(n3983), .ZN(n15840) );
  NAND2X0 U16311 ( .IN1(n5569), .IN2(n5383), .QN(n3983) );
  INVX0 U16312 ( .INP(n3492), .ZN(n15875) );
  NAND2X0 U16313 ( .IN1(n10587), .IN2(g3506), .QN(n3492) );
  NOR2X0 U16314 ( .IN1(n10452), .IN2(n10842), .QN(n15890) );
  NAND2X0 U16315 ( .IN1(n15894), .IN2(n15895), .QN(g30418) );
  NAND2X0 U16316 ( .IN1(n11076), .IN2(g3562), .QN(n15895) );
  NOR2X0 U16317 ( .IN1(n15896), .IN2(n15897), .QN(n15894) );
  NOR2X0 U16318 ( .IN1(n15008), .IN2(n15898), .QN(n15897) );
  INVX0 U16319 ( .INP(n4000), .ZN(n15898) );
  NOR2X0 U16320 ( .IN1(n4000), .IN2(n15899), .QN(n15896) );
  NAND2X0 U16321 ( .IN1(n10933), .IN2(g3558), .QN(n15899) );
  NAND2X0 U16322 ( .IN1(n15900), .IN2(n15901), .QN(g30417) );
  NAND2X0 U16323 ( .IN1(n11076), .IN2(g3554), .QN(n15901) );
  NOR2X0 U16324 ( .IN1(n15902), .IN2(n15903), .QN(n15900) );
  NOR2X0 U16325 ( .IN1(n15008), .IN2(n15904), .QN(n15903) );
  INVX0 U16326 ( .INP(n4003), .ZN(n15904) );
  NOR2X0 U16327 ( .IN1(n4003), .IN2(n15905), .QN(n15902) );
  NAND2X0 U16328 ( .IN1(n10933), .IN2(g3550), .QN(n15905) );
  NAND2X0 U16329 ( .IN1(n15906), .IN2(n15907), .QN(g30416) );
  NAND2X0 U16330 ( .IN1(n11076), .IN2(g3546), .QN(n15907) );
  NOR2X0 U16331 ( .IN1(n15908), .IN2(n15909), .QN(n15906) );
  NOR2X0 U16332 ( .IN1(n15008), .IN2(n15910), .QN(n15909) );
  INVX0 U16333 ( .INP(n4005), .ZN(n15910) );
  NOR2X0 U16334 ( .IN1(n4005), .IN2(n15911), .QN(n15908) );
  NAND2X0 U16335 ( .IN1(n10933), .IN2(g3542), .QN(n15911) );
  NAND2X0 U16336 ( .IN1(n15912), .IN2(n15913), .QN(g30415) );
  NAND2X0 U16337 ( .IN1(n11076), .IN2(g3530), .QN(n15913) );
  NOR2X0 U16338 ( .IN1(n15914), .IN2(n15915), .QN(n15912) );
  NOR2X0 U16339 ( .IN1(n15008), .IN2(n15916), .QN(n15915) );
  INVX0 U16340 ( .INP(n4007), .ZN(n15916) );
  NOR2X0 U16341 ( .IN1(n4007), .IN2(n15917), .QN(n15914) );
  NAND2X0 U16342 ( .IN1(n10932), .IN2(g3538), .QN(n15917) );
  NOR2X0 U16343 ( .IN1(g3506), .IN2(n14411), .QN(g30414) );
  NAND2X0 U16344 ( .IN1(n15918), .IN2(n5645), .QN(n14411) );
  NOR2X0 U16345 ( .IN1(n11039), .IN2(n14415), .QN(n15918) );
  INVX0 U16346 ( .INP(n14399), .ZN(n14415) );
  NAND2X0 U16347 ( .IN1(n15388), .IN2(n3799), .QN(n14399) );
  NOR2X0 U16348 ( .IN1(n5340), .IN2(g4087), .QN(n15388) );
  NAND2X0 U16349 ( .IN1(n15919), .IN2(n15920), .QN(g30413) );
  NAND2X0 U16350 ( .IN1(test_so84), .IN2(n11080), .QN(n15920) );
  NOR2X0 U16351 ( .IN1(n15921), .IN2(n15922), .QN(n15919) );
  NOR2X0 U16352 ( .IN1(n15923), .IN2(n15008), .QN(n15922) );
  NOR2X0 U16353 ( .IN1(n10284), .IN2(n15924), .QN(n15921) );
  NAND2X0 U16354 ( .IN1(n15925), .IN2(n15926), .QN(g30412) );
  NAND2X0 U16355 ( .IN1(n15927), .IN2(n3765), .QN(n15926) );
  NOR2X0 U16356 ( .IN1(n15928), .IN2(n15929), .QN(n15925) );
  NOR2X0 U16357 ( .IN1(n10457), .IN2(n10843), .QN(n15929) );
  NOR2X0 U16358 ( .IN1(n11039), .IN2(n15930), .QN(n15928) );
  NAND2X0 U16359 ( .IN1(n15931), .IN2(g3211), .QN(n15930) );
  INVX0 U16360 ( .INP(n15927), .ZN(n15931) );
  NOR2X0 U16361 ( .IN1(n580), .IN2(n5652), .QN(n15927) );
  NAND2X0 U16362 ( .IN1(n15932), .IN2(n15933), .QN(g30411) );
  NAND2X0 U16363 ( .IN1(n14429), .IN2(n3765), .QN(n15933) );
  INVX0 U16364 ( .INP(n15934), .ZN(n14429) );
  NOR2X0 U16365 ( .IN1(n15935), .IN2(n15936), .QN(n15932) );
  NOR2X0 U16366 ( .IN1(n10358), .IN2(n10843), .QN(n15936) );
  NOR2X0 U16367 ( .IN1(n11039), .IN2(n15937), .QN(n15935) );
  NAND2X0 U16368 ( .IN1(n15934), .IN2(g3203), .QN(n15937) );
  NAND2X0 U16369 ( .IN1(n15938), .IN2(g3167), .QN(n15934) );
  NAND2X0 U16370 ( .IN1(n15939), .IN2(n15940), .QN(g30410) );
  INVX0 U16371 ( .INP(n15941), .ZN(n15940) );
  NOR2X0 U16372 ( .IN1(n15942), .IN2(n15008), .QN(n15941) );
  NOR2X0 U16373 ( .IN1(n15943), .IN2(n15944), .QN(n15939) );
  NOR2X0 U16374 ( .IN1(n10285), .IN2(n10843), .QN(n15944) );
  NOR2X0 U16375 ( .IN1(n11039), .IN2(n15945), .QN(n15943) );
  NAND2X0 U16376 ( .IN1(test_so88), .IN2(n15942), .QN(n15945) );
  NAND2X0 U16377 ( .IN1(n15946), .IN2(g3167), .QN(n15942) );
  NAND2X0 U16378 ( .IN1(n15947), .IN2(n15948), .QN(g30409) );
  NAND2X0 U16379 ( .IN1(n4015), .IN2(n15949), .QN(n15948) );
  NOR2X0 U16380 ( .IN1(n15950), .IN2(n15951), .QN(n15947) );
  NOR2X0 U16381 ( .IN1(n11039), .IN2(n15952), .QN(n15951) );
  NAND2X0 U16382 ( .IN1(test_so84), .IN2(n15953), .QN(n15952) );
  NAND2X0 U16383 ( .IN1(n14440), .IN2(n15949), .QN(n15953) );
  NOR2X0 U16384 ( .IN1(n10334), .IN2(n10843), .QN(n15950) );
  NAND2X0 U16385 ( .IN1(n15954), .IN2(n15955), .QN(g30408) );
  NAND2X0 U16386 ( .IN1(n4015), .IN2(n14430), .QN(n15955) );
  NOR2X0 U16387 ( .IN1(n15956), .IN2(n15957), .QN(n15954) );
  NOR2X0 U16388 ( .IN1(n11039), .IN2(n15958), .QN(n15957) );
  NAND2X0 U16389 ( .IN1(n15959), .IN2(g3255), .QN(n15958) );
  NAND2X0 U16390 ( .IN1(n14440), .IN2(n14430), .QN(n15959) );
  NOR2X0 U16391 ( .IN1(n10455), .IN2(n10843), .QN(n15956) );
  NAND2X0 U16392 ( .IN1(n15960), .IN2(n15961), .QN(g30407) );
  NAND2X0 U16393 ( .IN1(n4015), .IN2(n15938), .QN(n15961) );
  NOR2X0 U16394 ( .IN1(n15962), .IN2(n15963), .QN(n15960) );
  NOR2X0 U16395 ( .IN1(n11039), .IN2(n15964), .QN(n15963) );
  NAND2X0 U16396 ( .IN1(n15965), .IN2(g3251), .QN(n15964) );
  NAND2X0 U16397 ( .IN1(n14440), .IN2(n15938), .QN(n15965) );
  NOR2X0 U16398 ( .IN1(n10373), .IN2(n10844), .QN(n15962) );
  NAND2X0 U16399 ( .IN1(n15966), .IN2(n15967), .QN(g30406) );
  NAND2X0 U16400 ( .IN1(n4015), .IN2(n15946), .QN(n15967) );
  NOR2X0 U16401 ( .IN1(n15968), .IN2(n15969), .QN(n15966) );
  NOR2X0 U16402 ( .IN1(n11039), .IN2(n15970), .QN(n15969) );
  NAND2X0 U16403 ( .IN1(n15971), .IN2(g3247), .QN(n15970) );
  NAND2X0 U16404 ( .IN1(n14440), .IN2(n15946), .QN(n15971) );
  INVX0 U16405 ( .INP(n128), .ZN(n14440) );
  NAND2X0 U16406 ( .IN1(g3161), .IN2(g3155), .QN(n128) );
  NOR2X0 U16407 ( .IN1(n10431), .IN2(n10844), .QN(n15968) );
  NAND2X0 U16408 ( .IN1(n15972), .IN2(n15973), .QN(g30405) );
  NAND2X0 U16409 ( .IN1(n4022), .IN2(n15949), .QN(n15973) );
  NOR2X0 U16410 ( .IN1(n15974), .IN2(n15975), .QN(n15972) );
  NOR2X0 U16411 ( .IN1(n11039), .IN2(n15976), .QN(n15975) );
  NAND2X0 U16412 ( .IN1(n15977), .IN2(g3243), .QN(n15976) );
  NAND2X0 U16413 ( .IN1(n15978), .IN2(n15949), .QN(n15977) );
  NOR2X0 U16414 ( .IN1(n10335), .IN2(n10844), .QN(n15974) );
  NAND2X0 U16415 ( .IN1(n15979), .IN2(n15980), .QN(g30404) );
  NAND2X0 U16416 ( .IN1(n4022), .IN2(n14430), .QN(n15980) );
  NOR2X0 U16417 ( .IN1(n15981), .IN2(n15982), .QN(n15979) );
  NOR2X0 U16418 ( .IN1(n11038), .IN2(n15983), .QN(n15982) );
  NAND2X0 U16419 ( .IN1(n15984), .IN2(g3239), .QN(n15983) );
  NAND2X0 U16420 ( .IN1(n15978), .IN2(n14430), .QN(n15984) );
  NOR2X0 U16421 ( .IN1(n10408), .IN2(n10844), .QN(n15981) );
  NAND2X0 U16422 ( .IN1(n15985), .IN2(n15986), .QN(g30403) );
  NAND2X0 U16423 ( .IN1(n4022), .IN2(n15938), .QN(n15986) );
  NOR2X0 U16424 ( .IN1(n15987), .IN2(n15988), .QN(n15985) );
  NOR2X0 U16425 ( .IN1(n11038), .IN2(n15989), .QN(n15988) );
  NAND2X0 U16426 ( .IN1(n15990), .IN2(g3235), .QN(n15989) );
  NAND2X0 U16427 ( .IN1(n15978), .IN2(n15938), .QN(n15990) );
  NOR2X0 U16428 ( .IN1(n10327), .IN2(n10844), .QN(n15987) );
  NAND2X0 U16429 ( .IN1(n15991), .IN2(n15992), .QN(g30402) );
  NAND2X0 U16430 ( .IN1(n4022), .IN2(n15946), .QN(n15992) );
  NOR2X0 U16431 ( .IN1(n15993), .IN2(n15994), .QN(n15991) );
  NOR2X0 U16432 ( .IN1(n11038), .IN2(n15995), .QN(n15994) );
  NAND2X0 U16433 ( .IN1(n15996), .IN2(g3231), .QN(n15995) );
  NAND2X0 U16434 ( .IN1(n15978), .IN2(n15946), .QN(n15996) );
  INVX0 U16435 ( .INP(n3502), .ZN(n15978) );
  NAND2X0 U16436 ( .IN1(n5366), .IN2(g3161), .QN(n3502) );
  NOR2X0 U16437 ( .IN1(n10286), .IN2(n10845), .QN(n15993) );
  NAND2X0 U16438 ( .IN1(n15997), .IN2(n15998), .QN(g30401) );
  NAND2X0 U16439 ( .IN1(n4027), .IN2(n15949), .QN(n15998) );
  NOR2X0 U16440 ( .IN1(n15999), .IN2(n16000), .QN(n15997) );
  NOR2X0 U16441 ( .IN1(n11038), .IN2(n16001), .QN(n16000) );
  NAND2X0 U16442 ( .IN1(n16002), .IN2(g3227), .QN(n16001) );
  NAND2X0 U16443 ( .IN1(n14446), .IN2(n15949), .QN(n16002) );
  NOR2X0 U16444 ( .IN1(n10409), .IN2(n10845), .QN(n15999) );
  NAND2X0 U16445 ( .IN1(n16003), .IN2(n16004), .QN(g30400) );
  NAND2X0 U16446 ( .IN1(n4027), .IN2(n14430), .QN(n16004) );
  NOR2X0 U16447 ( .IN1(n16005), .IN2(n16006), .QN(n16003) );
  NOR2X0 U16448 ( .IN1(n11038), .IN2(n16007), .QN(n16006) );
  NAND2X0 U16449 ( .IN1(n16008), .IN2(g3223), .QN(n16007) );
  NAND2X0 U16450 ( .IN1(n14446), .IN2(n14430), .QN(n16008) );
  INVX0 U16451 ( .INP(n580), .ZN(n14430) );
  NAND2X0 U16452 ( .IN1(n5603), .IN2(g3179), .QN(n580) );
  NOR2X0 U16453 ( .IN1(n10496), .IN2(n10845), .QN(n16005) );
  NAND2X0 U16454 ( .IN1(n16009), .IN2(n16010), .QN(g30399) );
  NAND2X0 U16455 ( .IN1(n4027), .IN2(n15938), .QN(n16010) );
  NOR2X0 U16456 ( .IN1(n16011), .IN2(n16012), .QN(n16009) );
  NOR2X0 U16457 ( .IN1(n11038), .IN2(n16013), .QN(n16012) );
  NAND2X0 U16458 ( .IN1(n16014), .IN2(g3219), .QN(n16013) );
  NAND2X0 U16459 ( .IN1(n14446), .IN2(n15938), .QN(n16014) );
  INVX0 U16460 ( .INP(n4020), .ZN(n15938) );
  NAND2X0 U16461 ( .IN1(n5390), .IN2(g3171), .QN(n4020) );
  NOR2X0 U16462 ( .IN1(n10287), .IN2(n10845), .QN(n16011) );
  NAND2X0 U16463 ( .IN1(n16015), .IN2(n16016), .QN(g30398) );
  NAND2X0 U16464 ( .IN1(n4027), .IN2(n15946), .QN(n16016) );
  NOR2X0 U16465 ( .IN1(n16017), .IN2(n16018), .QN(n16015) );
  NOR2X0 U16466 ( .IN1(n11038), .IN2(n16019), .QN(n16018) );
  NAND2X0 U16467 ( .IN1(n16020), .IN2(g3215), .QN(n16019) );
  NAND2X0 U16468 ( .IN1(n14446), .IN2(n15946), .QN(n16020) );
  INVX0 U16469 ( .INP(n4014), .ZN(n15946) );
  NAND2X0 U16470 ( .IN1(n5390), .IN2(n5603), .QN(n4014) );
  INVX0 U16471 ( .INP(n3501), .ZN(n14446) );
  NAND2X0 U16472 ( .IN1(n10578), .IN2(g3155), .QN(n3501) );
  NOR2X0 U16473 ( .IN1(n10439), .IN2(n10845), .QN(n16017) );
  NAND2X0 U16474 ( .IN1(n16021), .IN2(n16022), .QN(g30397) );
  NAND2X0 U16475 ( .IN1(n11076), .IN2(g3211), .QN(n16022) );
  NOR2X0 U16476 ( .IN1(n16023), .IN2(n16024), .QN(n16021) );
  NOR2X0 U16477 ( .IN1(n15008), .IN2(n16025), .QN(n16024) );
  INVX0 U16478 ( .INP(n4032), .ZN(n16025) );
  NOR2X0 U16479 ( .IN1(n4032), .IN2(n16026), .QN(n16023) );
  NAND2X0 U16480 ( .IN1(n10932), .IN2(g3207), .QN(n16026) );
  NAND2X0 U16481 ( .IN1(n16027), .IN2(n16028), .QN(g30396) );
  NAND2X0 U16482 ( .IN1(n11076), .IN2(g3203), .QN(n16028) );
  NOR2X0 U16483 ( .IN1(n16029), .IN2(n16030), .QN(n16027) );
  NOR2X0 U16484 ( .IN1(n15008), .IN2(n16031), .QN(n16030) );
  INVX0 U16485 ( .INP(n4035), .ZN(n16031) );
  NOR2X0 U16486 ( .IN1(n4035), .IN2(n16032), .QN(n16029) );
  NAND2X0 U16487 ( .IN1(n10932), .IN2(g3199), .QN(n16032) );
  NAND2X0 U16488 ( .IN1(n16033), .IN2(n16034), .QN(g30395) );
  NAND2X0 U16489 ( .IN1(test_so88), .IN2(n11080), .QN(n16034) );
  NOR2X0 U16490 ( .IN1(n16035), .IN2(n16036), .QN(n16033) );
  NOR2X0 U16491 ( .IN1(n15008), .IN2(n16037), .QN(n16036) );
  INVX0 U16492 ( .INP(n4037), .ZN(n16037) );
  NOR2X0 U16493 ( .IN1(n4037), .IN2(n16038), .QN(n16035) );
  NAND2X0 U16494 ( .IN1(n10932), .IN2(g3191), .QN(n16038) );
  NAND2X0 U16495 ( .IN1(n16039), .IN2(n16040), .QN(g30394) );
  NAND2X0 U16496 ( .IN1(n11076), .IN2(g3179), .QN(n16040) );
  NOR2X0 U16497 ( .IN1(n16041), .IN2(n16042), .QN(n16039) );
  NOR2X0 U16498 ( .IN1(n15008), .IN2(n16043), .QN(n16042) );
  INVX0 U16499 ( .INP(n4039), .ZN(n16043) );
  NOR2X0 U16500 ( .IN1(n4039), .IN2(n16044), .QN(n16041) );
  NAND2X0 U16501 ( .IN1(n10932), .IN2(g3187), .QN(n16044) );
  NOR2X0 U16502 ( .IN1(n14425), .IN2(n16045), .QN(g30393) );
  NAND2X0 U16503 ( .IN1(n5366), .IN2(n10956), .QN(n16045) );
  NAND2X0 U16504 ( .IN1(n5652), .IN2(n14437), .QN(n14425) );
  NAND2X0 U16505 ( .IN1(n3799), .IN2(n13425), .QN(n14437) );
  NAND2X0 U16506 ( .IN1(n16046), .IN2(n16047), .QN(g30392) );
  NAND2X0 U16507 ( .IN1(n11076), .IN2(g2803), .QN(n16047) );
  NAND2X0 U16508 ( .IN1(n16048), .IN2(n16049), .QN(g30391) );
  NAND2X0 U16509 ( .IN1(n11076), .IN2(g2771), .QN(n16049) );
  NAND2X0 U16510 ( .IN1(n16046), .IN2(n16050), .QN(g30390) );
  NAND2X0 U16511 ( .IN1(g2834), .IN2(n11080), .QN(n16050) );
  NAND2X0 U16512 ( .IN1(n16051), .IN2(n10956), .QN(n16046) );
  NAND2X0 U16513 ( .IN1(n16052), .IN2(n16053), .QN(n16051) );
  NAND2X0 U16514 ( .IN1(n16054), .IN2(n16055), .QN(n16053) );
  NOR2X0 U16515 ( .IN1(n16056), .IN2(n16057), .QN(n16054) );
  NAND2X0 U16516 ( .IN1(n16058), .IN2(n16059), .QN(n16057) );
  NAND2X0 U16517 ( .IN1(n10581), .IN2(n16060), .QN(n16059) );
  NAND2X0 U16518 ( .IN1(n10319), .IN2(n16061), .QN(n16058) );
  NAND2X0 U16519 ( .IN1(n16062), .IN2(n16063), .QN(n16056) );
  NAND2X0 U16520 ( .IN1(n10315), .IN2(n16064), .QN(n16063) );
  NAND2X0 U16521 ( .IN1(n10594), .IN2(n16065), .QN(n16062) );
  NAND2X0 U16522 ( .IN1(n16066), .IN2(n16067), .QN(n16052) );
  NOR2X0 U16523 ( .IN1(n16068), .IN2(n16069), .QN(n16066) );
  NAND2X0 U16524 ( .IN1(n16070), .IN2(n16071), .QN(n16069) );
  NAND2X0 U16525 ( .IN1(n16060), .IN2(g2815), .QN(n16071) );
  NAND2X0 U16526 ( .IN1(n16061), .IN2(g2807), .QN(n16070) );
  NAND2X0 U16527 ( .IN1(n16072), .IN2(n16073), .QN(n16068) );
  NAND2X0 U16528 ( .IN1(n16064), .IN2(g2803), .QN(n16073) );
  NAND2X0 U16529 ( .IN1(n16065), .IN2(g2819), .QN(n16072) );
  NAND2X0 U16530 ( .IN1(n16048), .IN2(n16074), .QN(g30389) );
  NAND2X0 U16531 ( .IN1(g2831), .IN2(n11081), .QN(n16074) );
  NAND2X0 U16532 ( .IN1(n16075), .IN2(n10956), .QN(n16048) );
  NAND2X0 U16533 ( .IN1(n16076), .IN2(n16077), .QN(n16075) );
  NAND2X0 U16534 ( .IN1(n16078), .IN2(n16055), .QN(n16077) );
  NOR2X0 U16535 ( .IN1(n16079), .IN2(n16080), .QN(n16078) );
  NAND2X0 U16536 ( .IN1(n16081), .IN2(n16082), .QN(n16080) );
  NAND2X0 U16537 ( .IN1(n16060), .IN2(n10669), .QN(n16082) );
  NAND2X0 U16538 ( .IN1(n10317), .IN2(n16061), .QN(n16081) );
  NAND2X0 U16539 ( .IN1(n16083), .IN2(n16084), .QN(n16079) );
  NAND2X0 U16540 ( .IN1(n10321), .IN2(n16064), .QN(n16084) );
  NAND2X0 U16541 ( .IN1(n10595), .IN2(n16065), .QN(n16083) );
  NAND2X0 U16542 ( .IN1(n16085), .IN2(n16067), .QN(n16076) );
  INVX0 U16543 ( .INP(n16055), .ZN(n16067) );
  NAND2X0 U16544 ( .IN1(n16086), .IN2(n5600), .QN(n16055) );
  NOR2X0 U16545 ( .IN1(n16087), .IN2(n14717), .QN(n16086) );
  NAND2X0 U16546 ( .IN1(n16088), .IN2(n5516), .QN(n14717) );
  NOR2X0 U16547 ( .IN1(test_so30), .IN2(g2741), .QN(n16088) );
  NOR2X0 U16548 ( .IN1(n16089), .IN2(n16090), .QN(n16085) );
  NAND2X0 U16549 ( .IN1(n16091), .IN2(n16092), .QN(n16090) );
  NAND2X0 U16550 ( .IN1(n16060), .IN2(g2783), .QN(n16092) );
  NAND2X0 U16551 ( .IN1(n16061), .IN2(g2775), .QN(n16091) );
  INVX0 U16552 ( .INP(n4411), .ZN(n16061) );
  NAND2X0 U16553 ( .IN1(n16093), .IN2(n16094), .QN(n16089) );
  NAND2X0 U16554 ( .IN1(n16064), .IN2(g2771), .QN(n16094) );
  NAND2X0 U16555 ( .IN1(n16065), .IN2(g2787), .QN(n16093) );
  NAND2X0 U16556 ( .IN1(n16095), .IN2(n16096), .QN(g30388) );
  NAND2X0 U16557 ( .IN1(n16097), .IN2(n3730), .QN(n16096) );
  XOR2X1 U16558 ( .IN1(n3506), .IN2(n5349), .Q(n16097) );
  NAND2X0 U16559 ( .IN1(n16098), .IN2(g2735), .QN(n3506) );
  NAND2X0 U16560 ( .IN1(n11076), .IN2(g2735), .QN(n16095) );
  NAND2X0 U16561 ( .IN1(n16099), .IN2(n16100), .QN(g30387) );
  INVX0 U16562 ( .INP(n16101), .ZN(n16100) );
  NOR2X0 U16563 ( .IN1(n16102), .IN2(n19404), .QN(n16101) );
  NOR2X0 U16564 ( .IN1(n16103), .IN2(n16104), .QN(n16099) );
  NOR2X0 U16565 ( .IN1(g2681), .IN2(n16105), .QN(n16104) );
  NAND2X0 U16566 ( .IN1(n16106), .IN2(n5457), .QN(n16105) );
  NOR2X0 U16567 ( .IN1(n5777), .IN2(n16107), .QN(n16103) );
  NOR2X0 U16568 ( .IN1(n11038), .IN2(n16108), .QN(n16107) );
  NOR2X0 U16569 ( .IN1(n5457), .IN2(n16109), .QN(n16108) );
  NAND2X0 U16570 ( .IN1(n16110), .IN2(n16111), .QN(g30386) );
  NAND2X0 U16571 ( .IN1(n16112), .IN2(g2681), .QN(n16111) );
  INVX0 U16572 ( .INP(n16102), .ZN(n16112) );
  NAND2X0 U16573 ( .IN1(n16102), .IN2(g2675), .QN(n16110) );
  NAND2X0 U16574 ( .IN1(n16113), .IN2(n16114), .QN(g30385) );
  NAND2X0 U16575 ( .IN1(n11076), .IN2(g2657), .QN(n16114) );
  NOR2X0 U16576 ( .IN1(n16115), .IN2(n16116), .QN(n16113) );
  NOR2X0 U16577 ( .IN1(g2661), .IN2(n16117), .QN(n16116) );
  NOR2X0 U16578 ( .IN1(n5418), .IN2(n16102), .QN(n16115) );
  NAND2X0 U16579 ( .IN1(n16109), .IN2(n10956), .QN(n16102) );
  NAND2X0 U16580 ( .IN1(n16118), .IN2(n16119), .QN(g30384) );
  NAND2X0 U16581 ( .IN1(n11076), .IN2(g2652), .QN(n16119) );
  NOR2X0 U16582 ( .IN1(n16120), .IN2(n16121), .QN(n16118) );
  NOR2X0 U16583 ( .IN1(n5316), .IN2(n16122), .QN(n16121) );
  NOR2X0 U16584 ( .IN1(n16123), .IN2(n14478), .QN(n16122) );
  INVX0 U16585 ( .INP(n11304), .ZN(n14478) );
  NOR2X0 U16586 ( .IN1(n11038), .IN2(n10628), .QN(n16123) );
  INVX0 U16587 ( .INP(n14483), .ZN(n10628) );
  NOR2X0 U16588 ( .IN1(n14483), .IN2(n16124), .QN(n16120) );
  NAND2X0 U16589 ( .IN1(n3517), .IN2(n16125), .QN(n16124) );
  XOR2X1 U16590 ( .IN1(n10324), .IN2(n10166), .Q(n16125) );
  INVX0 U16591 ( .INP(n14465), .ZN(n3517) );
  NAND2X0 U16592 ( .IN1(n16126), .IN2(n16127), .QN(g30383) );
  NAND2X0 U16593 ( .IN1(test_so66), .IN2(n11080), .QN(n16127) );
  NAND2X0 U16594 ( .IN1(n16128), .IN2(n10957), .QN(n16126) );
  NAND2X0 U16595 ( .IN1(n16129), .IN2(n16130), .QN(n16128) );
  NAND2X0 U16596 ( .IN1(test_so34), .IN2(n16131), .QN(n16130) );
  NAND2X0 U16597 ( .IN1(n16132), .IN2(n16133), .QN(n16129) );
  NAND2X0 U16598 ( .IN1(n5351), .IN2(g2599), .QN(n16133) );
  INVX0 U16599 ( .INP(n16131), .ZN(n16132) );
  NAND2X0 U16600 ( .IN1(n16134), .IN2(n5508), .QN(n16131) );
  NOR2X0 U16601 ( .IN1(n10529), .IN2(n11309), .QN(n16134) );
  NAND2X0 U16602 ( .IN1(n16135), .IN2(n16136), .QN(g30382) );
  INVX0 U16603 ( .INP(n16137), .ZN(n16136) );
  NOR2X0 U16604 ( .IN1(n16138), .IN2(n19401), .QN(n16137) );
  NOR2X0 U16605 ( .IN1(n16139), .IN2(n16140), .QN(n16135) );
  NOR2X0 U16606 ( .IN1(g2547), .IN2(n16141), .QN(n16140) );
  NAND2X0 U16607 ( .IN1(n16142), .IN2(n5461), .QN(n16141) );
  NOR2X0 U16608 ( .IN1(n5782), .IN2(n16143), .QN(n16139) );
  NOR2X0 U16609 ( .IN1(n11038), .IN2(n16144), .QN(n16143) );
  NOR2X0 U16610 ( .IN1(n5461), .IN2(n16145), .QN(n16144) );
  NAND2X0 U16611 ( .IN1(n16146), .IN2(n16147), .QN(g30381) );
  NAND2X0 U16612 ( .IN1(n16148), .IN2(g2547), .QN(n16147) );
  INVX0 U16613 ( .INP(n16138), .ZN(n16148) );
  NAND2X0 U16614 ( .IN1(n16138), .IN2(g2541), .QN(n16146) );
  NAND2X0 U16615 ( .IN1(n16149), .IN2(n16150), .QN(g30380) );
  NAND2X0 U16616 ( .IN1(n11076), .IN2(g2523), .QN(n16150) );
  NOR2X0 U16617 ( .IN1(n16151), .IN2(n16152), .QN(n16149) );
  NOR2X0 U16618 ( .IN1(g2527), .IN2(n16153), .QN(n16152) );
  NOR2X0 U16619 ( .IN1(n5420), .IN2(n16138), .QN(n16151) );
  NAND2X0 U16620 ( .IN1(n16145), .IN2(n10957), .QN(n16138) );
  NAND2X0 U16621 ( .IN1(n16154), .IN2(n16155), .QN(g30379) );
  NAND2X0 U16622 ( .IN1(n11075), .IN2(g2518), .QN(n16155) );
  NOR2X0 U16623 ( .IN1(n16156), .IN2(n16157), .QN(n16154) );
  NOR2X0 U16624 ( .IN1(n5281), .IN2(n16158), .QN(n16157) );
  NOR2X0 U16625 ( .IN1(n16159), .IN2(n14513), .QN(n16158) );
  INVX0 U16626 ( .INP(n11241), .ZN(n14513) );
  NOR2X0 U16627 ( .IN1(n11037), .IN2(n10635), .QN(n16159) );
  INVX0 U16628 ( .INP(n14518), .ZN(n10635) );
  NOR2X0 U16629 ( .IN1(n14518), .IN2(n16160), .QN(n16156) );
  NAND2X0 U16630 ( .IN1(n3536), .IN2(n16161), .QN(n16160) );
  XOR2X1 U16631 ( .IN1(n10323), .IN2(n10163), .Q(n16161) );
  INVX0 U16632 ( .INP(n14499), .ZN(n3536) );
  NAND2X0 U16633 ( .IN1(n16162), .IN2(n16163), .QN(g30378) );
  NAND2X0 U16634 ( .IN1(n11075), .IN2(g2441), .QN(n16163) );
  NAND2X0 U16635 ( .IN1(n16164), .IN2(n10957), .QN(n16162) );
  NAND2X0 U16636 ( .IN1(n16165), .IN2(n16166), .QN(n16164) );
  NAND2X0 U16637 ( .IN1(n16167), .IN2(g2461), .QN(n16166) );
  NAND2X0 U16638 ( .IN1(n16168), .IN2(n16169), .QN(n16165) );
  NAND2X0 U16639 ( .IN1(g2465), .IN2(n10648), .QN(n16169) );
  INVX0 U16640 ( .INP(n16167), .ZN(n16168) );
  NAND2X0 U16641 ( .IN1(n16170), .IN2(n5509), .QN(n16167) );
  NOR2X0 U16642 ( .IN1(n10530), .IN2(n11246), .QN(n16170) );
  NAND2X0 U16643 ( .IN1(n16171), .IN2(n16172), .QN(g30377) );
  INVX0 U16644 ( .INP(n16173), .ZN(n16172) );
  NOR2X0 U16645 ( .IN1(n16174), .IN2(n19403), .QN(n16173) );
  NOR2X0 U16646 ( .IN1(n16175), .IN2(n16176), .QN(n16171) );
  NOR2X0 U16647 ( .IN1(test_so89), .IN2(n16177), .QN(n16176) );
  NAND2X0 U16648 ( .IN1(n16178), .IN2(n5459), .QN(n16177) );
  NOR2X0 U16649 ( .IN1(n16179), .IN2(n10681), .QN(n16175) );
  NOR2X0 U16650 ( .IN1(n11037), .IN2(n16180), .QN(n16179) );
  NOR2X0 U16651 ( .IN1(n5459), .IN2(n16181), .QN(n16180) );
  NAND2X0 U16652 ( .IN1(n16182), .IN2(n16183), .QN(g30376) );
  NAND2X0 U16653 ( .IN1(test_so89), .IN2(n16184), .QN(n16183) );
  INVX0 U16654 ( .INP(n16174), .ZN(n16184) );
  NAND2X0 U16655 ( .IN1(n16174), .IN2(g2407), .QN(n16182) );
  NAND2X0 U16656 ( .IN1(n16185), .IN2(n16186), .QN(g30375) );
  NAND2X0 U16657 ( .IN1(n11075), .IN2(g2389), .QN(n16186) );
  NOR2X0 U16658 ( .IN1(n16187), .IN2(n16188), .QN(n16185) );
  NOR2X0 U16659 ( .IN1(g2393), .IN2(n16189), .QN(n16188) );
  NOR2X0 U16660 ( .IN1(n5421), .IN2(n16174), .QN(n16187) );
  NAND2X0 U16661 ( .IN1(n16181), .IN2(n10957), .QN(n16174) );
  NAND2X0 U16662 ( .IN1(n16190), .IN2(n16191), .QN(g30374) );
  NAND2X0 U16663 ( .IN1(n11075), .IN2(g2384), .QN(n16191) );
  NOR2X0 U16664 ( .IN1(n16192), .IN2(n16193), .QN(n16190) );
  NOR2X0 U16665 ( .IN1(n5631), .IN2(n16194), .QN(n16193) );
  NOR2X0 U16666 ( .IN1(n16195), .IN2(n14548), .QN(n16194) );
  INVX0 U16667 ( .INP(n11255), .ZN(n14548) );
  NOR2X0 U16668 ( .IN1(n11037), .IN2(n10630), .QN(n16195) );
  INVX0 U16669 ( .INP(n14553), .ZN(n10630) );
  NOR2X0 U16670 ( .IN1(n14553), .IN2(n16196), .QN(n16192) );
  NAND2X0 U16671 ( .IN1(n3555), .IN2(n16197), .QN(n16196) );
  XOR2X1 U16672 ( .IN1(n10318), .IN2(n10162), .Q(n16197) );
  INVX0 U16673 ( .INP(n14534), .ZN(n3555) );
  NAND2X0 U16674 ( .IN1(n16198), .IN2(n16199), .QN(g30373) );
  NAND2X0 U16675 ( .IN1(n11075), .IN2(g2307), .QN(n16199) );
  NAND2X0 U16676 ( .IN1(n16200), .IN2(n10957), .QN(n16198) );
  NAND2X0 U16677 ( .IN1(n16201), .IN2(n16202), .QN(n16200) );
  NAND2X0 U16678 ( .IN1(n16203), .IN2(g2327), .QN(n16202) );
  NAND2X0 U16679 ( .IN1(n16204), .IN2(n16205), .QN(n16201) );
  NAND2X0 U16680 ( .IN1(n5353), .IN2(g2331), .QN(n16205) );
  INVX0 U16681 ( .INP(n16203), .ZN(n16204) );
  NAND2X0 U16682 ( .IN1(n16206), .IN2(n5511), .QN(n16203) );
  NOR2X0 U16683 ( .IN1(n10640), .IN2(n11260), .QN(n16206) );
  NAND2X0 U16684 ( .IN1(n16207), .IN2(n16208), .QN(g30372) );
  INVX0 U16685 ( .INP(n16209), .ZN(n16208) );
  NOR2X0 U16686 ( .IN1(n16210), .IN2(n19402), .QN(n16209) );
  NOR2X0 U16687 ( .IN1(n16211), .IN2(n16212), .QN(n16207) );
  NOR2X0 U16688 ( .IN1(g2279), .IN2(n16213), .QN(n16212) );
  NAND2X0 U16689 ( .IN1(n16214), .IN2(n5458), .QN(n16213) );
  NOR2X0 U16690 ( .IN1(n5778), .IN2(n16215), .QN(n16211) );
  NOR2X0 U16691 ( .IN1(n11037), .IN2(n16216), .QN(n16215) );
  NOR2X0 U16692 ( .IN1(n5458), .IN2(n16217), .QN(n16216) );
  NAND2X0 U16693 ( .IN1(n16218), .IN2(n16219), .QN(g30371) );
  NAND2X0 U16694 ( .IN1(n16220), .IN2(g2279), .QN(n16219) );
  INVX0 U16695 ( .INP(n16210), .ZN(n16220) );
  NAND2X0 U16696 ( .IN1(n16210), .IN2(g2273), .QN(n16218) );
  NAND2X0 U16697 ( .IN1(n16221), .IN2(n16222), .QN(g30370) );
  NAND2X0 U16698 ( .IN1(n11075), .IN2(g2255), .QN(n16222) );
  NOR2X0 U16699 ( .IN1(n16223), .IN2(n16224), .QN(n16221) );
  NOR2X0 U16700 ( .IN1(g2259), .IN2(n16225), .QN(n16224) );
  NOR2X0 U16701 ( .IN1(n5419), .IN2(n16210), .QN(n16223) );
  NAND2X0 U16702 ( .IN1(n16217), .IN2(n10958), .QN(n16210) );
  NAND2X0 U16703 ( .IN1(n16226), .IN2(n16227), .QN(g30369) );
  NAND2X0 U16704 ( .IN1(n11075), .IN2(g2250), .QN(n16227) );
  NOR2X0 U16705 ( .IN1(n16228), .IN2(n16229), .QN(n16226) );
  NOR2X0 U16706 ( .IN1(n5414), .IN2(n16230), .QN(n16229) );
  NOR2X0 U16707 ( .IN1(n16231), .IN2(n14583), .QN(n16230) );
  INVX0 U16708 ( .INP(n11490), .ZN(n14583) );
  NOR2X0 U16709 ( .IN1(n11037), .IN2(n10636), .QN(n16231) );
  INVX0 U16710 ( .INP(n14588), .ZN(n10636) );
  NOR2X0 U16711 ( .IN1(n14588), .IN2(n16232), .QN(n16228) );
  NAND2X0 U16712 ( .IN1(n3574), .IN2(n16233), .QN(n16232) );
  XOR2X1 U16713 ( .IN1(n10314), .IN2(n10165), .Q(n16233) );
  INVX0 U16714 ( .INP(n14569), .ZN(n3574) );
  NAND2X0 U16715 ( .IN1(n16234), .IN2(n16235), .QN(g30368) );
  NAND2X0 U16716 ( .IN1(n11075), .IN2(g2173), .QN(n16235) );
  NAND2X0 U16717 ( .IN1(n16236), .IN2(n10958), .QN(n16234) );
  NAND2X0 U16718 ( .IN1(n16237), .IN2(n16238), .QN(n16236) );
  NAND2X0 U16719 ( .IN1(n16239), .IN2(g2193), .QN(n16238) );
  NAND2X0 U16720 ( .IN1(n16240), .IN2(n16241), .QN(n16237) );
  NAND2X0 U16721 ( .IN1(n5356), .IN2(g2197), .QN(n16241) );
  INVX0 U16722 ( .INP(n16239), .ZN(n16240) );
  NAND2X0 U16723 ( .IN1(n16242), .IN2(n5512), .QN(n16239) );
  NOR2X0 U16724 ( .IN1(n10532), .IN2(n11495), .QN(n16242) );
  NAND2X0 U16725 ( .IN1(n16243), .IN2(n16244), .QN(g30367) );
  INVX0 U16726 ( .INP(n16245), .ZN(n16244) );
  NOR2X0 U16727 ( .IN1(n16246), .IN2(n5891), .QN(n16245) );
  NOR2X0 U16728 ( .IN1(n16247), .IN2(n16248), .QN(n16243) );
  NOR2X0 U16729 ( .IN1(g2122), .IN2(n16249), .QN(n16248) );
  NAND2X0 U16730 ( .IN1(n16250), .IN2(n5463), .QN(n16249) );
  NOR2X0 U16731 ( .IN1(n5784), .IN2(n16251), .QN(n16247) );
  NOR2X0 U16732 ( .IN1(n11037), .IN2(n16252), .QN(n16251) );
  NOR2X0 U16733 ( .IN1(n5463), .IN2(n16253), .QN(n16252) );
  NAND2X0 U16734 ( .IN1(n16254), .IN2(n16255), .QN(g30366) );
  NAND2X0 U16735 ( .IN1(n16256), .IN2(g2122), .QN(n16255) );
  INVX0 U16736 ( .INP(n16246), .ZN(n16256) );
  NAND2X0 U16737 ( .IN1(n16246), .IN2(g2116), .QN(n16254) );
  NAND2X0 U16738 ( .IN1(n16257), .IN2(n16258), .QN(g30365) );
  INVX0 U16739 ( .INP(n16259), .ZN(n16258) );
  NOR2X0 U16740 ( .IN1(n10902), .IN2(n5280), .QN(n16259) );
  NOR2X0 U16741 ( .IN1(n16260), .IN2(n16261), .QN(n16257) );
  NOR2X0 U16742 ( .IN1(g2102), .IN2(n16262), .QN(n16261) );
  NOR2X0 U16743 ( .IN1(n5666), .IN2(n16246), .QN(n16260) );
  NAND2X0 U16744 ( .IN1(n16253), .IN2(n10958), .QN(n16246) );
  NAND2X0 U16745 ( .IN1(n16263), .IN2(n16264), .QN(g30364) );
  NAND2X0 U16746 ( .IN1(test_so78), .IN2(n11081), .QN(n16264) );
  NOR2X0 U16747 ( .IN1(n16265), .IN2(n16266), .QN(n16263) );
  NOR2X0 U16748 ( .IN1(n5280), .IN2(n16267), .QN(n16266) );
  NOR2X0 U16749 ( .IN1(n16268), .IN2(n14621), .QN(n16267) );
  INVX0 U16750 ( .INP(n14605), .ZN(n14621) );
  NOR2X0 U16751 ( .IN1(n11037), .IN2(n10637), .QN(n16268) );
  NOR2X0 U16752 ( .IN1(n16269), .IN2(n16270), .QN(n16265) );
  NAND2X0 U16753 ( .IN1(n10637), .IN2(n3593), .QN(n16270) );
  INVX0 U16754 ( .INP(n14606), .ZN(n3593) );
  INVX0 U16755 ( .INP(n14626), .ZN(n10637) );
  XOR2X1 U16756 ( .IN1(test_so78), .IN2(n10161), .Q(n16269) );
  NAND2X0 U16757 ( .IN1(n16271), .IN2(n16272), .QN(g30363) );
  NAND2X0 U16758 ( .IN1(n11075), .IN2(g2016), .QN(n16272) );
  NAND2X0 U16759 ( .IN1(n16273), .IN2(n10958), .QN(n16271) );
  NAND2X0 U16760 ( .IN1(n16274), .IN2(n16275), .QN(n16273) );
  NAND2X0 U16761 ( .IN1(test_so59), .IN2(n16276), .QN(n16275) );
  NAND2X0 U16762 ( .IN1(n16277), .IN2(n16278), .QN(n16274) );
  NAND2X0 U16763 ( .IN1(n5355), .IN2(g2040), .QN(n16278) );
  INVX0 U16764 ( .INP(n16276), .ZN(n16277) );
  NAND2X0 U16765 ( .IN1(n16279), .IN2(n5507), .QN(n16276) );
  NOR2X0 U16766 ( .IN1(n10528), .IN2(n14598), .QN(n16279) );
  NAND2X0 U16767 ( .IN1(n16280), .IN2(n16281), .QN(g30362) );
  INVX0 U16768 ( .INP(n16282), .ZN(n16281) );
  NOR2X0 U16769 ( .IN1(n16283), .IN2(n5890), .QN(n16282) );
  NOR2X0 U16770 ( .IN1(n16284), .IN2(n16285), .QN(n16280) );
  NOR2X0 U16771 ( .IN1(g1988), .IN2(n16286), .QN(n16285) );
  NAND2X0 U16772 ( .IN1(n16287), .IN2(n5462), .QN(n16286) );
  NOR2X0 U16773 ( .IN1(n5783), .IN2(n16288), .QN(n16284) );
  NOR2X0 U16774 ( .IN1(n11037), .IN2(n16289), .QN(n16288) );
  NOR2X0 U16775 ( .IN1(n5462), .IN2(n16290), .QN(n16289) );
  NAND2X0 U16776 ( .IN1(n16291), .IN2(n16292), .QN(g30361) );
  NAND2X0 U16777 ( .IN1(n16293), .IN2(g1988), .QN(n16292) );
  INVX0 U16778 ( .INP(n16283), .ZN(n16293) );
  NAND2X0 U16779 ( .IN1(n16283), .IN2(g1982), .QN(n16291) );
  NAND2X0 U16780 ( .IN1(n16294), .IN2(n16295), .QN(g30360) );
  INVX0 U16781 ( .INP(n16296), .ZN(n16295) );
  NOR2X0 U16782 ( .IN1(n10903), .IN2(n5315), .QN(n16296) );
  NOR2X0 U16783 ( .IN1(n16297), .IN2(n16298), .QN(n16294) );
  NOR2X0 U16784 ( .IN1(g1968), .IN2(n16299), .QN(n16298) );
  NOR2X0 U16785 ( .IN1(n5664), .IN2(n16283), .QN(n16297) );
  NAND2X0 U16786 ( .IN1(n16290), .IN2(n10958), .QN(n16283) );
  NAND2X0 U16787 ( .IN1(n16300), .IN2(n16301), .QN(g30359) );
  NAND2X0 U16788 ( .IN1(n11075), .IN2(g1959), .QN(n16301) );
  NOR2X0 U16789 ( .IN1(n16302), .IN2(n16303), .QN(n16300) );
  NOR2X0 U16790 ( .IN1(n5315), .IN2(n16304), .QN(n16303) );
  NOR2X0 U16791 ( .IN1(n16305), .IN2(n14657), .QN(n16304) );
  INVX0 U16792 ( .INP(n11314), .ZN(n14657) );
  NOR2X0 U16793 ( .IN1(n11036), .IN2(n10627), .QN(n16305) );
  INVX0 U16794 ( .INP(n14662), .ZN(n10627) );
  NOR2X0 U16795 ( .IN1(n14662), .IN2(n16306), .QN(n16302) );
  NAND2X0 U16796 ( .IN1(n3611), .IN2(n16307), .QN(n16306) );
  XOR2X1 U16797 ( .IN1(n10322), .IN2(n10159), .Q(n16307) );
  INVX0 U16798 ( .INP(n14642), .ZN(n3611) );
  NAND2X0 U16799 ( .IN1(n16308), .IN2(n16309), .QN(g30358) );
  NAND2X0 U16800 ( .IN1(n11075), .IN2(g1882), .QN(n16309) );
  NAND2X0 U16801 ( .IN1(n16310), .IN2(n10959), .QN(n16308) );
  NAND2X0 U16802 ( .IN1(n16311), .IN2(n16312), .QN(n16310) );
  NAND2X0 U16803 ( .IN1(n16313), .IN2(g1902), .QN(n16312) );
  NAND2X0 U16804 ( .IN1(n16314), .IN2(n16315), .QN(n16311) );
  NAND2X0 U16805 ( .IN1(g1906), .IN2(n10657), .QN(n16315) );
  INVX0 U16806 ( .INP(n16313), .ZN(n16314) );
  NAND2X0 U16807 ( .IN1(n16316), .IN2(n5510), .QN(n16313) );
  NOR2X0 U16808 ( .IN1(n10531), .IN2(n11319), .QN(n16316) );
  NAND2X0 U16809 ( .IN1(n16317), .IN2(n16318), .QN(g30357) );
  INVX0 U16810 ( .INP(n16319), .ZN(n16318) );
  NOR2X0 U16811 ( .IN1(n16320), .IN2(n5892), .QN(n16319) );
  NOR2X0 U16812 ( .IN1(n16321), .IN2(n16322), .QN(n16317) );
  NOR2X0 U16813 ( .IN1(g1854), .IN2(n16323), .QN(n16322) );
  NAND2X0 U16814 ( .IN1(n16324), .IN2(n5464), .QN(n16323) );
  NOR2X0 U16815 ( .IN1(n5785), .IN2(n16325), .QN(n16321) );
  NOR2X0 U16816 ( .IN1(n11036), .IN2(n16326), .QN(n16325) );
  NOR2X0 U16817 ( .IN1(n5464), .IN2(n16327), .QN(n16326) );
  NAND2X0 U16818 ( .IN1(n16328), .IN2(n16329), .QN(g30356) );
  NAND2X0 U16819 ( .IN1(n16330), .IN2(g1854), .QN(n16329) );
  INVX0 U16820 ( .INP(n16320), .ZN(n16330) );
  NAND2X0 U16821 ( .IN1(n16320), .IN2(g1848), .QN(n16328) );
  NAND2X0 U16822 ( .IN1(n16331), .IN2(n16332), .QN(g30355) );
  NAND2X0 U16823 ( .IN1(n11075), .IN2(g1830), .QN(n16332) );
  NOR2X0 U16824 ( .IN1(n16333), .IN2(n16334), .QN(n16331) );
  NOR2X0 U16825 ( .IN1(g1834), .IN2(n16335), .QN(n16334) );
  NOR2X0 U16826 ( .IN1(n5665), .IN2(n16320), .QN(n16333) );
  NAND2X0 U16827 ( .IN1(n16327), .IN2(n10959), .QN(n16320) );
  NAND2X0 U16828 ( .IN1(n16336), .IN2(n16337), .QN(g30354) );
  NAND2X0 U16829 ( .IN1(n11075), .IN2(g1825), .QN(n16337) );
  NOR2X0 U16830 ( .IN1(n16338), .IN2(n16339), .QN(n16336) );
  NOR2X0 U16831 ( .IN1(n5413), .IN2(n16340), .QN(n16339) );
  NOR2X0 U16832 ( .IN1(n16341), .IN2(n14691), .QN(n16340) );
  INVX0 U16833 ( .INP(n11225), .ZN(n14691) );
  NOR2X0 U16834 ( .IN1(n11036), .IN2(n10633), .QN(n16341) );
  INVX0 U16835 ( .INP(n14696), .ZN(n10633) );
  NOR2X0 U16836 ( .IN1(n14696), .IN2(n16342), .QN(n16338) );
  NAND2X0 U16837 ( .IN1(n3628), .IN2(n16343), .QN(n16342) );
  XOR2X1 U16838 ( .IN1(n10316), .IN2(n10160), .Q(n16343) );
  INVX0 U16839 ( .INP(n14678), .ZN(n3628) );
  NAND2X0 U16840 ( .IN1(n16344), .IN2(n16345), .QN(g30353) );
  NAND2X0 U16841 ( .IN1(n11075), .IN2(g1748), .QN(n16345) );
  NAND2X0 U16842 ( .IN1(n16346), .IN2(n10959), .QN(n16344) );
  NAND2X0 U16843 ( .IN1(n16347), .IN2(n16348), .QN(n16346) );
  NAND2X0 U16844 ( .IN1(n16349), .IN2(g1768), .QN(n16348) );
  NAND2X0 U16845 ( .IN1(n16350), .IN2(n16351), .QN(n16347) );
  NAND2X0 U16846 ( .IN1(n5352), .IN2(g1772), .QN(n16351) );
  INVX0 U16847 ( .INP(n16349), .ZN(n16350) );
  NAND2X0 U16848 ( .IN1(n16352), .IN2(n5359), .QN(n16349) );
  NOR2X0 U16849 ( .IN1(n5596), .IN2(n11230), .QN(n16352) );
  NAND2X0 U16850 ( .IN1(n16353), .IN2(n16354), .QN(g30352) );
  NAND2X0 U16851 ( .IN1(n16355), .IN2(n9236), .QN(n16354) );
  NOR2X0 U16852 ( .IN1(n16356), .IN2(n16357), .QN(n16353) );
  NOR2X0 U16853 ( .IN1(g1720), .IN2(n16358), .QN(n16357) );
  NAND2X0 U16854 ( .IN1(n16359), .IN2(n16360), .QN(n16358) );
  NOR2X0 U16855 ( .IN1(n11036), .IN2(g1714), .QN(n16359) );
  NOR2X0 U16856 ( .IN1(n5780), .IN2(n16361), .QN(n16356) );
  NOR2X0 U16857 ( .IN1(n11036), .IN2(n16362), .QN(n16361) );
  NOR2X0 U16858 ( .IN1(n5460), .IN2(n16363), .QN(n16362) );
  NAND2X0 U16859 ( .IN1(n16364), .IN2(n16365), .QN(g30351) );
  NAND2X0 U16860 ( .IN1(n16355), .IN2(g1720), .QN(n16365) );
  NAND2X0 U16861 ( .IN1(n16366), .IN2(g1714), .QN(n16364) );
  NAND2X0 U16862 ( .IN1(n16367), .IN2(n16368), .QN(g30350) );
  NAND2X0 U16863 ( .IN1(n16355), .IN2(g1700), .QN(n16368) );
  INVX0 U16864 ( .INP(n16366), .ZN(n16355) );
  NAND2X0 U16865 ( .IN1(n16363), .IN2(n10959), .QN(n16366) );
  NOR2X0 U16866 ( .IN1(n16369), .IN2(n16370), .QN(n16367) );
  NOR2X0 U16867 ( .IN1(n5628), .IN2(n10847), .QN(n16370) );
  NOR2X0 U16868 ( .IN1(n11036), .IN2(n16371), .QN(n16369) );
  NAND2X0 U16869 ( .IN1(n16360), .IN2(n5417), .QN(n16371) );
  INVX0 U16870 ( .INP(n16363), .ZN(n16360) );
  NAND2X0 U16871 ( .IN1(n16372), .IN2(n16373), .QN(g30349) );
  NAND2X0 U16872 ( .IN1(n11075), .IN2(g1691), .QN(n16373) );
  NOR2X0 U16873 ( .IN1(n16374), .IN2(n16375), .QN(n16372) );
  NOR2X0 U16874 ( .IN1(n5628), .IN2(n16376), .QN(n16375) );
  NOR2X0 U16875 ( .IN1(n16377), .IN2(n14728), .QN(n16376) );
  NOR2X0 U16876 ( .IN1(n11036), .IN2(n1418), .QN(n16377) );
  NOR2X0 U16877 ( .IN1(n14733), .IN2(n16378), .QN(n16374) );
  NAND2X0 U16878 ( .IN1(n3646), .IN2(n16379), .QN(n16378) );
  XOR2X1 U16879 ( .IN1(n10320), .IN2(n10164), .Q(n16379) );
  INVX0 U16880 ( .INP(n14712), .ZN(n3646) );
  NAND2X0 U16881 ( .IN1(n16380), .IN2(n16381), .QN(g30348) );
  NAND2X0 U16882 ( .IN1(n11075), .IN2(g1612), .QN(n16381) );
  NOR2X0 U16883 ( .IN1(n16382), .IN2(n16383), .QN(n16380) );
  NOR2X0 U16884 ( .IN1(n5836), .IN2(n16384), .QN(n16383) );
  NOR2X0 U16885 ( .IN1(n16385), .IN2(n14728), .QN(n16384) );
  INVX0 U16886 ( .INP(n11471), .ZN(n14728) );
  NOR2X0 U16887 ( .IN1(n11036), .IN2(g25167), .QN(n16385) );
  NOR2X0 U16888 ( .IN1(n14712), .IN2(n16386), .QN(n16382) );
  NAND2X0 U16889 ( .IN1(g25167), .IN2(n16387), .QN(n16386) );
  NAND2X0 U16890 ( .IN1(n5362), .IN2(g1636), .QN(n16387) );
  NAND2X0 U16891 ( .IN1(n16388), .IN2(n16389), .QN(g30347) );
  NAND2X0 U16892 ( .IN1(n16390), .IN2(n16391), .QN(n16389) );
  NOR2X0 U16893 ( .IN1(n16392), .IN2(n16393), .QN(n16390) );
  NOR2X0 U16894 ( .IN1(n16394), .IN2(n16395), .QN(n16393) );
  NOR2X0 U16895 ( .IN1(n10090), .IN2(n11015), .QN(n16395) );
  INVX0 U16896 ( .INP(n16396), .ZN(n16388) );
  NOR2X0 U16897 ( .IN1(n10905), .IN2(n10584), .QN(n16396) );
  NAND2X0 U16898 ( .IN1(n16397), .IN2(n16398), .QN(g30346) );
  NAND2X0 U16899 ( .IN1(n11075), .IN2(g1536), .QN(n16398) );
  NAND2X0 U16900 ( .IN1(n16399), .IN2(n10960), .QN(n16397) );
  NOR2X0 U16901 ( .IN1(n16400), .IN2(n16401), .QN(n16399) );
  NAND2X0 U16902 ( .IN1(n16402), .IN2(n16403), .QN(n16401) );
  NAND2X0 U16903 ( .IN1(n10584), .IN2(n16404), .QN(n16402) );
  NAND2X0 U16904 ( .IN1(n16405), .IN2(n16406), .QN(g30345) );
  NAND2X0 U16905 ( .IN1(n16407), .IN2(n10960), .QN(n16406) );
  NAND2X0 U16906 ( .IN1(n16391), .IN2(n13811), .QN(n16407) );
  INVX0 U16907 ( .INP(n16400), .ZN(n16391) );
  NAND2X0 U16908 ( .IN1(n16408), .IN2(g1514), .QN(n16405) );
  NAND2X0 U16909 ( .IN1(n16409), .IN2(n10960), .QN(n16408) );
  XOR2X1 U16910 ( .IN1(test_so49), .IN2(n5302), .Q(n16409) );
  NOR2X0 U16911 ( .IN1(n11035), .IN2(n16410), .QN(g30344) );
  NOR2X0 U16912 ( .IN1(n16400), .IN2(n16411), .QN(n16410) );
  XOR2X1 U16913 ( .IN1(n5364), .IN2(n5302), .Q(n16411) );
  NAND2X0 U16914 ( .IN1(n16412), .IN2(n16413), .QN(n16400) );
  NAND2X0 U16915 ( .IN1(n2), .IN2(n16414), .QN(n16412) );
  NOR2X0 U16916 ( .IN1(n16415), .IN2(n16416), .QN(n2) );
  NAND2X0 U16917 ( .IN1(n4895), .IN2(n10398), .QN(n16416) );
  NAND2X0 U16918 ( .IN1(n16417), .IN2(g1521), .QN(n16415) );
  NAND2X0 U16919 ( .IN1(n16418), .IN2(n16419), .QN(g30343) );
  NAND2X0 U16920 ( .IN1(n4175), .IN2(n14739), .QN(n16419) );
  NOR2X0 U16921 ( .IN1(n16420), .IN2(n16421), .QN(n16418) );
  NOR2X0 U16922 ( .IN1(n11035), .IN2(n16422), .QN(n16421) );
  NAND2X0 U16923 ( .IN1(n11421), .IN2(g1361), .QN(n16422) );
  NAND2X0 U16924 ( .IN1(n16423), .IN2(n16424), .QN(n11421) );
  NAND2X0 U16925 ( .IN1(n10249), .IN2(n14121), .QN(n16423) );
  INVX0 U16926 ( .INP(n14126), .ZN(n14121) );
  NOR2X0 U16927 ( .IN1(n10249), .IN2(n10848), .QN(n16420) );
  NAND2X0 U16928 ( .IN1(n16425), .IN2(n16426), .QN(g30342) );
  NAND2X0 U16929 ( .IN1(n11074), .IN2(g1256), .QN(n16426) );
  NOR2X0 U16930 ( .IN1(n16427), .IN2(n16428), .QN(n16425) );
  NOR2X0 U16931 ( .IN1(g1259), .IN2(n16429), .QN(n16428) );
  NOR2X0 U16932 ( .IN1(n5553), .IN2(n16430), .QN(n16427) );
  NAND2X0 U16933 ( .IN1(n14133), .IN2(n16429), .QN(n16430) );
  INVX0 U16934 ( .INP(n3736), .ZN(n16429) );
  NAND2X0 U16935 ( .IN1(n16431), .IN2(n16432), .QN(g30341) );
  NAND2X0 U16936 ( .IN1(n16433), .IN2(n16434), .QN(n16432) );
  NOR2X0 U16937 ( .IN1(n16435), .IN2(n16436), .QN(n16433) );
  NOR2X0 U16938 ( .IN1(n16437), .IN2(n16438), .QN(n16436) );
  NOR2X0 U16939 ( .IN1(n10089), .IN2(n11015), .QN(n16438) );
  INVX0 U16940 ( .INP(n16439), .ZN(n16431) );
  NOR2X0 U16941 ( .IN1(n10906), .IN2(n10583), .QN(n16439) );
  NAND2X0 U16942 ( .IN1(n16440), .IN2(n16441), .QN(g30340) );
  INVX0 U16943 ( .INP(n16442), .ZN(n16441) );
  NOR2X0 U16944 ( .IN1(n10907), .IN2(n10606), .QN(n16442) );
  NAND2X0 U16945 ( .IN1(n16443), .IN2(n10960), .QN(n16440) );
  NOR2X0 U16946 ( .IN1(n16444), .IN2(n16445), .QN(n16443) );
  NAND2X0 U16947 ( .IN1(n16446), .IN2(n16447), .QN(n16445) );
  NAND2X0 U16948 ( .IN1(n10583), .IN2(n16448), .QN(n16446) );
  NAND2X0 U16949 ( .IN1(n16449), .IN2(n16450), .QN(g30339) );
  NAND2X0 U16950 ( .IN1(n16451), .IN2(n10960), .QN(n16450) );
  NAND2X0 U16951 ( .IN1(n16434), .IN2(n16452), .QN(n16451) );
  NAND2X0 U16952 ( .IN1(n16453), .IN2(g1171), .QN(n16449) );
  NAND2X0 U16953 ( .IN1(n16454), .IN2(n10961), .QN(n16453) );
  XOR2X1 U16954 ( .IN1(g7916), .IN2(n5599), .Q(n16454) );
  NOR2X0 U16955 ( .IN1(n11035), .IN2(n16455), .QN(g30338) );
  NOR2X0 U16956 ( .IN1(n16444), .IN2(n16456), .QN(n16455) );
  XOR2X1 U16957 ( .IN1(n5363), .IN2(n5304), .Q(n16456) );
  INVX0 U16958 ( .INP(n16434), .ZN(n16444) );
  NOR2X0 U16959 ( .IN1(n16457), .IN2(n4191), .QN(n16434) );
  NOR2X0 U16960 ( .IN1(n16458), .IN2(n16452), .QN(n16457) );
  INVX0 U16961 ( .INP(n4), .ZN(n16458) );
  NOR2X0 U16962 ( .IN1(n16459), .IN2(n16460), .QN(n4) );
  NAND2X0 U16963 ( .IN1(n5642), .IN2(n4920), .QN(n16460) );
  NAND2X0 U16964 ( .IN1(n16461), .IN2(g1178), .QN(n16459) );
  NOR2X0 U16965 ( .IN1(n5304), .IN2(n10255), .QN(n16461) );
  NAND2X0 U16966 ( .IN1(n16462), .IN2(n16463), .QN(g30337) );
  NAND2X0 U16967 ( .IN1(n4193), .IN2(n14756), .QN(n16463) );
  NOR2X0 U16968 ( .IN1(n16464), .IN2(n16465), .QN(n16462) );
  NOR2X0 U16969 ( .IN1(n11035), .IN2(n16466), .QN(n16465) );
  NAND2X0 U16970 ( .IN1(n11420), .IN2(g1018), .QN(n16466) );
  NAND2X0 U16971 ( .IN1(n16467), .IN2(n16468), .QN(n11420) );
  NAND2X0 U16972 ( .IN1(n10250), .IN2(n14140), .QN(n16467) );
  INVX0 U16973 ( .INP(n14145), .ZN(n14140) );
  NOR2X0 U16974 ( .IN1(n10250), .IN2(n10848), .QN(n16464) );
  NAND2X0 U16975 ( .IN1(n16469), .IN2(n16470), .QN(g30336) );
  NAND2X0 U16976 ( .IN1(n11074), .IN2(g911), .QN(n16470) );
  NOR2X0 U16977 ( .IN1(n16471), .IN2(n16472), .QN(n16469) );
  NOR2X0 U16978 ( .IN1(g914), .IN2(n16473), .QN(n16472) );
  NOR2X0 U16979 ( .IN1(n5560), .IN2(n16474), .QN(n16471) );
  NAND2X0 U16980 ( .IN1(n14152), .IN2(n16473), .QN(n16474) );
  INVX0 U16981 ( .INP(n3741), .ZN(n16473) );
  NAND2X0 U16982 ( .IN1(n16475), .IN2(n16476), .QN(g30335) );
  NAND2X0 U16983 ( .IN1(test_so60), .IN2(n11081), .QN(n16476) );
  NOR2X0 U16984 ( .IN1(n16477), .IN2(n16478), .QN(n16475) );
  NOR2X0 U16985 ( .IN1(g744), .IN2(n11419), .QN(n16478) );
  NOR2X0 U16986 ( .IN1(n5470), .IN2(n16479), .QN(n16477) );
  NAND2X0 U16987 ( .IN1(n2404), .IN2(n11419), .QN(n16479) );
  NAND2X0 U16988 ( .IN1(n16480), .IN2(test_so60), .QN(n11419) );
  NOR2X0 U16989 ( .IN1(n11404), .IN2(n16481), .QN(n16480) );
  NOR2X0 U16990 ( .IN1(g736), .IN2(n5482), .QN(n11404) );
  NAND2X0 U16991 ( .IN1(n16482), .IN2(n16483), .QN(g30334) );
  NAND2X0 U16992 ( .IN1(n11074), .IN2(g586), .QN(n16483) );
  NOR2X0 U16993 ( .IN1(n16484), .IN2(n16485), .QN(n16482) );
  NOR2X0 U16994 ( .IN1(g577), .IN2(n16486), .QN(n16485) );
  NOR2X0 U16995 ( .IN1(n5294), .IN2(n16487), .QN(n16484) );
  NAND2X0 U16996 ( .IN1(n2421), .IN2(n16486), .QN(n16487) );
  INVX0 U16997 ( .INP(n3745), .ZN(n16486) );
  NAND2X0 U16998 ( .IN1(n16488), .IN2(n16489), .QN(g30333) );
  NAND2X0 U16999 ( .IN1(n12641), .IN2(n16490), .QN(n16489) );
  XNOR2X1 U17000 ( .IN1(test_so73), .IN2(n14970), .Q(n16490) );
  NOR2X0 U17001 ( .IN1(n14971), .IN2(n11016), .QN(n12641) );
  NAND2X0 U17002 ( .IN1(n16491), .IN2(n16492), .QN(n14971) );
  INVX0 U17003 ( .INP(n16493), .ZN(n16492) );
  NOR2X0 U17004 ( .IN1(n14970), .IN2(n16494), .QN(n16493) );
  NOR2X0 U17005 ( .IN1(n16495), .IN2(test_so72), .QN(n16494) );
  NOR2X0 U17006 ( .IN1(n5520), .IN2(n16496), .QN(n16491) );
  NAND2X0 U17007 ( .IN1(n11074), .IN2(g142), .QN(n16488) );
  NAND2X0 U17008 ( .IN1(n16497), .IN2(n16498), .QN(g29309) );
  NAND2X0 U17009 ( .IN1(n3765), .IN2(n16499), .QN(n16498) );
  NAND2X0 U17010 ( .IN1(g6541), .IN2(n13440), .QN(n16499) );
  NOR2X0 U17011 ( .IN1(n16500), .IN2(n16501), .QN(n16497) );
  NOR2X0 U17012 ( .IN1(n15009), .IN2(n16502), .QN(n16501) );
  NAND2X0 U17013 ( .IN1(n16503), .IN2(g6541), .QN(n16502) );
  NAND2X0 U17014 ( .IN1(n16504), .IN2(n16505), .QN(g29308) );
  NAND2X0 U17015 ( .IN1(n11074), .IN2(g6523), .QN(n16505) );
  NOR2X0 U17016 ( .IN1(n16506), .IN2(n16507), .QN(n16504) );
  INVX0 U17017 ( .INP(n16508), .ZN(n16507) );
  NAND2X0 U17018 ( .IN1(n16509), .IN2(n5659), .QN(n16508) );
  NOR2X0 U17019 ( .IN1(n5659), .IN2(n11298), .QN(n16506) );
  NAND2X0 U17020 ( .IN1(n16510), .IN2(n16511), .QN(g29307) );
  NAND2X0 U17021 ( .IN1(n11297), .IN2(g6523), .QN(n16511) );
  INVX0 U17022 ( .INP(n11298), .ZN(n11297) );
  NAND2X0 U17023 ( .IN1(n16512), .IN2(n10961), .QN(n11298) );
  NOR2X0 U17024 ( .IN1(n16513), .IN2(n16514), .QN(n16510) );
  NOR2X0 U17025 ( .IN1(g6519), .IN2(n16515), .QN(n16514) );
  NAND2X0 U17026 ( .IN1(n5426), .IN2(n16509), .QN(n16515) );
  NOR2X0 U17027 ( .IN1(n5806), .IN2(n16516), .QN(n16513) );
  NOR2X0 U17028 ( .IN1(n11035), .IN2(n16517), .QN(n16516) );
  NOR2X0 U17029 ( .IN1(n5426), .IN2(n16512), .QN(n16517) );
  NAND2X0 U17030 ( .IN1(n16518), .IN2(n16519), .QN(g29305) );
  NAND2X0 U17031 ( .IN1(n12021), .IN2(n16512), .QN(n16519) );
  NOR2X0 U17032 ( .IN1(n11035), .IN2(n10171), .QN(n12021) );
  NOR2X0 U17033 ( .IN1(n16520), .IN2(n16521), .QN(n16518) );
  NOR2X0 U17034 ( .IN1(g6500), .IN2(n16522), .QN(n16521) );
  NAND2X0 U17035 ( .IN1(n16509), .IN2(g6505), .QN(n16522) );
  NOR2X0 U17036 ( .IN1(n16512), .IN2(n11017), .QN(n16509) );
  NOR2X0 U17037 ( .IN1(n5748), .IN2(n16523), .QN(n16520) );
  NOR2X0 U17038 ( .IN1(n11035), .IN2(n16524), .QN(n16523) );
  NOR2X0 U17039 ( .IN1(n16512), .IN2(g6505), .QN(n16524) );
  NAND2X0 U17040 ( .IN1(n16525), .IN2(n13464), .QN(n16512) );
  NAND2X0 U17041 ( .IN1(n16526), .IN2(n16527), .QN(g29304) );
  NAND2X0 U17042 ( .IN1(n11074), .IN2(g6505), .QN(n16527) );
  NAND2X0 U17043 ( .IN1(n16528), .IN2(n10961), .QN(n16526) );
  NAND2X0 U17044 ( .IN1(n16529), .IN2(n16530), .QN(n16528) );
  NAND2X0 U17045 ( .IN1(n10629), .IN2(g6500), .QN(n16530) );
  INVX0 U17046 ( .INP(n13464), .ZN(n10629) );
  NAND2X0 U17047 ( .IN1(n16531), .IN2(n13464), .QN(n16529) );
  XOR2X1 U17048 ( .IN1(n16532), .IN2(n16533), .Q(n16531) );
  NOR2X0 U17049 ( .IN1(n16525), .IN2(n5748), .QN(n16533) );
  NOR2X0 U17050 ( .IN1(n16534), .IN2(n11283), .QN(n16525) );
  NAND2X0 U17051 ( .IN1(g6727), .IN2(g17722), .QN(n16534) );
  NAND2X0 U17052 ( .IN1(n16535), .IN2(n16536), .QN(g29303) );
  NAND2X0 U17053 ( .IN1(n3765), .IN2(n16537), .QN(n16536) );
  NAND2X0 U17054 ( .IN1(g6195), .IN2(n13434), .QN(n16537) );
  NOR2X0 U17055 ( .IN1(n16500), .IN2(n16538), .QN(n16535) );
  NOR2X0 U17056 ( .IN1(n15137), .IN2(n16539), .QN(n16538) );
  NAND2X0 U17057 ( .IN1(n16503), .IN2(g6195), .QN(n16539) );
  NAND2X0 U17058 ( .IN1(n16540), .IN2(n16541), .QN(g29302) );
  NAND2X0 U17059 ( .IN1(n11074), .IN2(g6177), .QN(n16541) );
  NOR2X0 U17060 ( .IN1(n16542), .IN2(n16543), .QN(n16540) );
  INVX0 U17061 ( .INP(n16544), .ZN(n16543) );
  NAND2X0 U17062 ( .IN1(n16545), .IN2(n5667), .QN(n16544) );
  NOR2X0 U17063 ( .IN1(n5667), .IN2(n16546), .QN(n16542) );
  NAND2X0 U17064 ( .IN1(n16547), .IN2(n16548), .QN(g29301) );
  NAND2X0 U17065 ( .IN1(n16549), .IN2(g6177), .QN(n16548) );
  NOR2X0 U17066 ( .IN1(n16550), .IN2(n16551), .QN(n16547) );
  NOR2X0 U17067 ( .IN1(g6173), .IN2(n16552), .QN(n16551) );
  NAND2X0 U17068 ( .IN1(n5430), .IN2(n16545), .QN(n16552) );
  NOR2X0 U17069 ( .IN1(n5810), .IN2(n16553), .QN(n16550) );
  NOR2X0 U17070 ( .IN1(n11035), .IN2(n16554), .QN(n16553) );
  NOR2X0 U17071 ( .IN1(n5430), .IN2(n16555), .QN(n16554) );
  NAND2X0 U17072 ( .IN1(n16556), .IN2(n16557), .QN(g29300) );
  NAND2X0 U17073 ( .IN1(n16549), .IN2(g6173), .QN(n16557) );
  NAND2X0 U17074 ( .IN1(n16546), .IN2(g6167), .QN(n16556) );
  NAND2X0 U17075 ( .IN1(n16558), .IN2(n16559), .QN(g29299) );
  NAND2X0 U17076 ( .IN1(n16549), .IN2(g6163), .QN(n16559) );
  INVX0 U17077 ( .INP(n16546), .ZN(n16549) );
  NAND2X0 U17078 ( .IN1(n16555), .IN2(n10961), .QN(n16546) );
  NOR2X0 U17079 ( .IN1(n16560), .IN2(n16561), .QN(n16558) );
  NOR2X0 U17080 ( .IN1(g6154), .IN2(n16562), .QN(n16561) );
  NAND2X0 U17081 ( .IN1(n16545), .IN2(g6159), .QN(n16562) );
  NOR2X0 U17082 ( .IN1(n16555), .IN2(n11017), .QN(n16545) );
  NOR2X0 U17083 ( .IN1(n5747), .IN2(n16563), .QN(n16560) );
  NOR2X0 U17084 ( .IN1(n11034), .IN2(n16564), .QN(n16563) );
  NOR2X0 U17085 ( .IN1(n16555), .IN2(g6159), .QN(n16564) );
  NAND2X0 U17086 ( .IN1(n16565), .IN2(n13485), .QN(n16555) );
  NAND2X0 U17087 ( .IN1(n16566), .IN2(n16567), .QN(g29298) );
  NAND2X0 U17088 ( .IN1(n11074), .IN2(g6159), .QN(n16567) );
  NAND2X0 U17089 ( .IN1(n16568), .IN2(n10961), .QN(n16566) );
  NAND2X0 U17090 ( .IN1(n16569), .IN2(n16570), .QN(n16568) );
  NAND2X0 U17091 ( .IN1(n13483), .IN2(g6154), .QN(n16570) );
  NAND2X0 U17092 ( .IN1(n16571), .IN2(n13485), .QN(n16569) );
  XOR2X1 U17093 ( .IN1(n16572), .IN2(n16573), .Q(n16571) );
  NOR2X0 U17094 ( .IN1(n16565), .IN2(n5747), .QN(n16573) );
  NOR2X0 U17095 ( .IN1(n16574), .IN2(n10642), .QN(n16565) );
  NAND2X0 U17096 ( .IN1(g17685), .IN2(n16575), .QN(n16574) );
  NAND2X0 U17097 ( .IN1(n16576), .IN2(n16577), .QN(g29297) );
  NAND2X0 U17098 ( .IN1(n3765), .IN2(n16578), .QN(n16577) );
  NAND2X0 U17099 ( .IN1(g5849), .IN2(n13433), .QN(n16578) );
  NOR2X0 U17100 ( .IN1(n16500), .IN2(n16579), .QN(n16576) );
  NOR2X0 U17101 ( .IN1(n15265), .IN2(n16580), .QN(n16579) );
  NAND2X0 U17102 ( .IN1(n16503), .IN2(g5849), .QN(n16580) );
  NAND2X0 U17103 ( .IN1(n16581), .IN2(n16582), .QN(g29296) );
  NAND2X0 U17104 ( .IN1(n11074), .IN2(g5831), .QN(n16582) );
  NOR2X0 U17105 ( .IN1(n16583), .IN2(n16584), .QN(n16581) );
  INVX0 U17106 ( .INP(n16585), .ZN(n16584) );
  NAND2X0 U17107 ( .IN1(n16586), .IN2(n5663), .QN(n16585) );
  NOR2X0 U17108 ( .IN1(n5663), .IN2(n11455), .QN(n16583) );
  NAND2X0 U17109 ( .IN1(n16587), .IN2(n16588), .QN(g29295) );
  NAND2X0 U17110 ( .IN1(n11454), .IN2(g5831), .QN(n16588) );
  NOR2X0 U17111 ( .IN1(n16589), .IN2(n16590), .QN(n16587) );
  NOR2X0 U17112 ( .IN1(g5827), .IN2(n16591), .QN(n16590) );
  NAND2X0 U17113 ( .IN1(n5429), .IN2(n16586), .QN(n16591) );
  NOR2X0 U17114 ( .IN1(n5809), .IN2(n16592), .QN(n16589) );
  NOR2X0 U17115 ( .IN1(n11034), .IN2(n16593), .QN(n16592) );
  NOR2X0 U17116 ( .IN1(n5429), .IN2(n16594), .QN(n16593) );
  NAND2X0 U17117 ( .IN1(n16595), .IN2(n16596), .QN(g29293) );
  NAND2X0 U17118 ( .IN1(n11454), .IN2(g5817), .QN(n16596) );
  INVX0 U17119 ( .INP(n11455), .ZN(n11454) );
  NAND2X0 U17120 ( .IN1(n16594), .IN2(n10962), .QN(n11455) );
  NOR2X0 U17121 ( .IN1(n16597), .IN2(n16598), .QN(n16595) );
  NOR2X0 U17122 ( .IN1(g5808), .IN2(n16599), .QN(n16598) );
  NAND2X0 U17123 ( .IN1(n16586), .IN2(g5813), .QN(n16599) );
  NOR2X0 U17124 ( .IN1(n16594), .IN2(n11018), .QN(n16586) );
  NOR2X0 U17125 ( .IN1(n5749), .IN2(n16600), .QN(n16597) );
  NOR2X0 U17126 ( .IN1(n11034), .IN2(n16601), .QN(n16600) );
  NOR2X0 U17127 ( .IN1(n16594), .IN2(g5813), .QN(n16601) );
  NAND2X0 U17128 ( .IN1(n13506), .IN2(n16602), .QN(n16594) );
  NAND2X0 U17129 ( .IN1(n16603), .IN2(n16604), .QN(g29292) );
  NAND2X0 U17130 ( .IN1(n11074), .IN2(g5813), .QN(n16604) );
  NOR2X0 U17131 ( .IN1(n16605), .IN2(n16606), .QN(n16603) );
  NOR2X0 U17132 ( .IN1(n5749), .IN2(n13511), .QN(n16606) );
  NOR2X0 U17133 ( .IN1(n13515), .IN2(n16607), .QN(n16605) );
  XNOR2X1 U17134 ( .IN1(n16608), .IN2(n16609), .Q(n16607) );
  NOR2X0 U17135 ( .IN1(n16602), .IN2(n5749), .QN(n16609) );
  NOR2X0 U17136 ( .IN1(n16610), .IN2(n12451), .QN(n16602) );
  NAND2X0 U17137 ( .IN1(g6035), .IN2(g17646), .QN(n16610) );
  NAND2X0 U17138 ( .IN1(n16611), .IN2(n16612), .QN(g29291) );
  NAND2X0 U17139 ( .IN1(n3765), .IN2(n16613), .QN(n16612) );
  NAND2X0 U17140 ( .IN1(g5503), .IN2(n15393), .QN(n16613) );
  NOR2X0 U17141 ( .IN1(n16500), .IN2(n16614), .QN(n16611) );
  NOR2X0 U17142 ( .IN1(n11251), .IN2(n16615), .QN(n16614) );
  NAND2X0 U17143 ( .IN1(n16503), .IN2(g5503), .QN(n16615) );
  NAND2X0 U17144 ( .IN1(n16616), .IN2(n16617), .QN(g29290) );
  NAND2X0 U17145 ( .IN1(n11074), .IN2(g5485), .QN(n16617) );
  NOR2X0 U17146 ( .IN1(n16618), .IN2(n16619), .QN(n16616) );
  NOR2X0 U17147 ( .IN1(n16620), .IN2(g5489), .QN(n16619) );
  NOR2X0 U17148 ( .IN1(n5660), .IN2(n11459), .QN(n16618) );
  NAND2X0 U17149 ( .IN1(n16621), .IN2(n16622), .QN(g29289) );
  NAND2X0 U17150 ( .IN1(n11458), .IN2(g5485), .QN(n16622) );
  NOR2X0 U17151 ( .IN1(n16623), .IN2(n16624), .QN(n16621) );
  NOR2X0 U17152 ( .IN1(g5481), .IN2(n16625), .QN(n16624) );
  NAND2X0 U17153 ( .IN1(n5425), .IN2(n16626), .QN(n16625) );
  NOR2X0 U17154 ( .IN1(n5805), .IN2(n16627), .QN(n16623) );
  NOR2X0 U17155 ( .IN1(n11034), .IN2(n16628), .QN(n16627) );
  NOR2X0 U17156 ( .IN1(n5425), .IN2(n16629), .QN(n16628) );
  NAND2X0 U17157 ( .IN1(n16630), .IN2(n16631), .QN(g29287) );
  NAND2X0 U17158 ( .IN1(n11458), .IN2(g5471), .QN(n16631) );
  INVX0 U17159 ( .INP(n11459), .ZN(n11458) );
  NAND2X0 U17160 ( .IN1(n16629), .IN2(n10962), .QN(n11459) );
  NOR2X0 U17161 ( .IN1(n16632), .IN2(n16633), .QN(n16630) );
  NOR2X0 U17162 ( .IN1(g5462), .IN2(n16634), .QN(n16633) );
  NAND2X0 U17163 ( .IN1(n16626), .IN2(g5467), .QN(n16634) );
  INVX0 U17164 ( .INP(n16620), .ZN(n16626) );
  NAND2X0 U17165 ( .IN1(n16635), .IN2(n10962), .QN(n16620) );
  NOR2X0 U17166 ( .IN1(n5744), .IN2(n16636), .QN(n16632) );
  NOR2X0 U17167 ( .IN1(n11034), .IN2(n16637), .QN(n16636) );
  NOR2X0 U17168 ( .IN1(n16629), .IN2(g5467), .QN(n16637) );
  INVX0 U17169 ( .INP(n16635), .ZN(n16629) );
  NOR2X0 U17170 ( .IN1(n16638), .IN2(n13525), .QN(n16635) );
  NAND2X0 U17171 ( .IN1(n16639), .IN2(n16640), .QN(g29286) );
  NAND2X0 U17172 ( .IN1(n11074), .IN2(g5467), .QN(n16640) );
  NAND2X0 U17173 ( .IN1(n16641), .IN2(n10962), .QN(n16639) );
  NAND2X0 U17174 ( .IN1(n16642), .IN2(n16643), .QN(n16641) );
  NAND2X0 U17175 ( .IN1(n13525), .IN2(g5462), .QN(n16643) );
  NAND2X0 U17176 ( .IN1(n16644), .IN2(n13527), .QN(n16642) );
  XNOR2X1 U17177 ( .IN1(n16645), .IN2(n16646), .Q(n16644) );
  NAND2X0 U17178 ( .IN1(g5462), .IN2(n16638), .QN(n16645) );
  NAND2X0 U17179 ( .IN1(n16647), .IN2(n16648), .QN(n16638) );
  NOR2X0 U17180 ( .IN1(n5529), .IN2(n10473), .QN(n16647) );
  NAND2X0 U17181 ( .IN1(n16649), .IN2(n16650), .QN(g29285) );
  NAND2X0 U17182 ( .IN1(n3765), .IN2(n16651), .QN(n16650) );
  NAND2X0 U17183 ( .IN1(g5156), .IN2(n13429), .QN(n16651) );
  NOR2X0 U17184 ( .IN1(n16500), .IN2(n16652), .QN(n16649) );
  NOR2X0 U17185 ( .IN1(n15520), .IN2(n16653), .QN(n16652) );
  NAND2X0 U17186 ( .IN1(n16503), .IN2(g5156), .QN(n16653) );
  NAND2X0 U17187 ( .IN1(n16654), .IN2(n16655), .QN(g29284) );
  NAND2X0 U17188 ( .IN1(n11074), .IN2(g5138), .QN(n16655) );
  NOR2X0 U17189 ( .IN1(n16656), .IN2(n16657), .QN(n16654) );
  INVX0 U17190 ( .INP(n16658), .ZN(n16657) );
  NAND2X0 U17191 ( .IN1(n16659), .IN2(n5658), .QN(n16658) );
  NOR2X0 U17192 ( .IN1(n5658), .IN2(n16660), .QN(n16656) );
  NAND2X0 U17193 ( .IN1(n16661), .IN2(n16662), .QN(g29283) );
  NAND2X0 U17194 ( .IN1(n16663), .IN2(g5138), .QN(n16662) );
  NOR2X0 U17195 ( .IN1(n16664), .IN2(n16665), .QN(n16661) );
  NOR2X0 U17196 ( .IN1(g5134), .IN2(n16666), .QN(n16665) );
  NAND2X0 U17197 ( .IN1(n16659), .IN2(n10654), .QN(n16666) );
  NOR2X0 U17198 ( .IN1(n5807), .IN2(n16667), .QN(n16664) );
  NOR2X0 U17199 ( .IN1(n11034), .IN2(n16668), .QN(n16667) );
  NOR2X0 U17200 ( .IN1(n16669), .IN2(n10654), .QN(n16668) );
  NAND2X0 U17201 ( .IN1(n16670), .IN2(n16671), .QN(g29282) );
  NAND2X0 U17202 ( .IN1(n16663), .IN2(g5134), .QN(n16671) );
  INVX0 U17203 ( .INP(n16660), .ZN(n16663) );
  NAND2X0 U17204 ( .IN1(test_so96), .IN2(n16660), .QN(n16670) );
  NAND2X0 U17205 ( .IN1(n16669), .IN2(n10962), .QN(n16660) );
  NAND2X0 U17206 ( .IN1(n16672), .IN2(n16673), .QN(g29281) );
  NAND2X0 U17207 ( .IN1(n14981), .IN2(n16669), .QN(n16673) );
  NOR2X0 U17208 ( .IN1(n11034), .IN2(n10129), .QN(n14981) );
  NOR2X0 U17209 ( .IN1(n16674), .IN2(n16675), .QN(n16672) );
  NOR2X0 U17210 ( .IN1(g5115), .IN2(n16676), .QN(n16675) );
  NAND2X0 U17211 ( .IN1(n16659), .IN2(g5120), .QN(n16676) );
  NOR2X0 U17212 ( .IN1(n16669), .IN2(n11019), .QN(n16659) );
  NOR2X0 U17213 ( .IN1(n5743), .IN2(n16677), .QN(n16674) );
  NOR2X0 U17214 ( .IN1(n11034), .IN2(n16678), .QN(n16677) );
  NOR2X0 U17215 ( .IN1(n16669), .IN2(g5120), .QN(n16678) );
  NAND2X0 U17216 ( .IN1(n16679), .IN2(g33959), .QN(n16669) );
  NAND2X0 U17217 ( .IN1(n16680), .IN2(n16681), .QN(g29280) );
  NAND2X0 U17218 ( .IN1(n11074), .IN2(g5120), .QN(n16681) );
  NAND2X0 U17219 ( .IN1(n16682), .IN2(n10963), .QN(n16680) );
  NAND2X0 U17220 ( .IN1(n16683), .IN2(n16684), .QN(n16682) );
  NAND2X0 U17221 ( .IN1(n10624), .IN2(g5115), .QN(n16684) );
  NAND2X0 U17222 ( .IN1(n16685), .IN2(g33959), .QN(n16683) );
  XOR2X1 U17223 ( .IN1(n16686), .IN2(n16687), .Q(n16685) );
  NOR2X0 U17224 ( .IN1(n16679), .IN2(n5743), .QN(n16687) );
  NOR2X0 U17225 ( .IN1(n16688), .IN2(n10641), .QN(n16679) );
  NAND2X0 U17226 ( .IN1(g17577), .IN2(g31860), .QN(n16688) );
  NAND2X0 U17227 ( .IN1(n16689), .IN2(n16690), .QN(g29275) );
  NAND2X0 U17228 ( .IN1(n16691), .IN2(n16692), .QN(n16690) );
  XOR2X1 U17229 ( .IN1(n14910), .IN2(g4087), .Q(n16691) );
  NOR2X0 U17230 ( .IN1(n10644), .IN2(n16693), .QN(n14910) );
  NAND2X0 U17231 ( .IN1(test_so11), .IN2(n11081), .QN(n16689) );
  NAND2X0 U17232 ( .IN1(n16694), .IN2(n16695), .QN(g29274) );
  NAND2X0 U17233 ( .IN1(n3765), .IN2(n16696), .QN(n16695) );
  NAND2X0 U17234 ( .IN1(g3849), .IN2(n13445), .QN(n16696) );
  NOR2X0 U17235 ( .IN1(n16500), .IN2(n16697), .QN(n16694) );
  NOR2X0 U17236 ( .IN1(n15669), .IN2(n16698), .QN(n16697) );
  NAND2X0 U17237 ( .IN1(n16503), .IN2(g3849), .QN(n16698) );
  NAND2X0 U17238 ( .IN1(n16699), .IN2(n16700), .QN(g29273) );
  NAND2X0 U17239 ( .IN1(n11074), .IN2(g3831), .QN(n16700) );
  NOR2X0 U17240 ( .IN1(n16701), .IN2(n16702), .QN(n16699) );
  INVX0 U17241 ( .INP(n16703), .ZN(n16702) );
  NAND2X0 U17242 ( .IN1(n16704), .IN2(n5662), .QN(n16703) );
  NOR2X0 U17243 ( .IN1(n5662), .IN2(n16705), .QN(n16701) );
  NAND2X0 U17244 ( .IN1(n16706), .IN2(n16707), .QN(g29272) );
  NAND2X0 U17245 ( .IN1(n16708), .IN2(g3831), .QN(n16707) );
  NOR2X0 U17246 ( .IN1(n16709), .IN2(n16710), .QN(n16706) );
  NOR2X0 U17247 ( .IN1(g3827), .IN2(n16711), .QN(n16710) );
  NAND2X0 U17248 ( .IN1(n5428), .IN2(n16704), .QN(n16711) );
  NOR2X0 U17249 ( .IN1(n5808), .IN2(n16712), .QN(n16709) );
  NOR2X0 U17250 ( .IN1(n11033), .IN2(n16713), .QN(n16712) );
  NOR2X0 U17251 ( .IN1(n5428), .IN2(n16714), .QN(n16713) );
  NAND2X0 U17252 ( .IN1(n16715), .IN2(n16716), .QN(g29271) );
  NAND2X0 U17253 ( .IN1(n16708), .IN2(g3827), .QN(n16716) );
  INVX0 U17254 ( .INP(n16705), .ZN(n16708) );
  NAND2X0 U17255 ( .IN1(n16705), .IN2(g3821), .QN(n16715) );
  NAND2X0 U17256 ( .IN1(n16714), .IN2(n10963), .QN(n16705) );
  NAND2X0 U17257 ( .IN1(n16717), .IN2(n16718), .QN(g29270) );
  NAND2X0 U17258 ( .IN1(n14997), .IN2(n16714), .QN(n16718) );
  NOR2X0 U17259 ( .IN1(n11033), .IN2(n10130), .QN(n14997) );
  NOR2X0 U17260 ( .IN1(n16719), .IN2(n16720), .QN(n16717) );
  NOR2X0 U17261 ( .IN1(g3808), .IN2(n16721), .QN(n16720) );
  NAND2X0 U17262 ( .IN1(n16704), .IN2(g3813), .QN(n16721) );
  NOR2X0 U17263 ( .IN1(n16714), .IN2(n11019), .QN(n16704) );
  NOR2X0 U17264 ( .IN1(n5745), .IN2(n16722), .QN(n16719) );
  NOR2X0 U17265 ( .IN1(n11033), .IN2(n16723), .QN(n16722) );
  NOR2X0 U17266 ( .IN1(n16714), .IN2(g3813), .QN(n16723) );
  NAND2X0 U17267 ( .IN1(n16724), .IN2(n13583), .QN(n16714) );
  NAND2X0 U17268 ( .IN1(n16725), .IN2(n16726), .QN(g29269) );
  NAND2X0 U17269 ( .IN1(n11074), .IN2(g3813), .QN(n16726) );
  NAND2X0 U17270 ( .IN1(n16727), .IN2(n10963), .QN(n16725) );
  NAND2X0 U17271 ( .IN1(n16728), .IN2(n16729), .QN(n16727) );
  NAND2X0 U17272 ( .IN1(n13581), .IN2(g3808), .QN(n16729) );
  NAND2X0 U17273 ( .IN1(n16730), .IN2(n13583), .QN(n16728) );
  XOR2X1 U17274 ( .IN1(n16731), .IN2(n16732), .Q(n16730) );
  NOR2X0 U17275 ( .IN1(n16724), .IN2(n5745), .QN(n16732) );
  NOR2X0 U17276 ( .IN1(n16733), .IN2(n12454), .QN(n16724) );
  NAND2X0 U17277 ( .IN1(g4040), .IN2(g16693), .QN(n16733) );
  NAND2X0 U17278 ( .IN1(n16734), .IN2(n16735), .QN(g29268) );
  NAND2X0 U17279 ( .IN1(n3765), .IN2(n16736), .QN(n16735) );
  NAND2X0 U17280 ( .IN1(g3498), .IN2(n13444), .QN(n16736) );
  NOR2X0 U17281 ( .IN1(n16500), .IN2(n16737), .QN(n16734) );
  NOR2X0 U17282 ( .IN1(n15796), .IN2(n16738), .QN(n16737) );
  NAND2X0 U17283 ( .IN1(n16503), .IN2(g3498), .QN(n16738) );
  NAND2X0 U17284 ( .IN1(n16739), .IN2(n16740), .QN(g29267) );
  NAND2X0 U17285 ( .IN1(n11074), .IN2(g3480), .QN(n16740) );
  NOR2X0 U17286 ( .IN1(n16741), .IN2(n16742), .QN(n16739) );
  INVX0 U17287 ( .INP(n16743), .ZN(n16742) );
  NAND2X0 U17288 ( .IN1(n16744), .IN2(n5668), .QN(n16743) );
  NOR2X0 U17289 ( .IN1(n5668), .IN2(n16745), .QN(n16741) );
  NAND2X0 U17290 ( .IN1(n16746), .IN2(n16747), .QN(g29266) );
  NAND2X0 U17291 ( .IN1(n16748), .IN2(g3480), .QN(n16747) );
  NOR2X0 U17292 ( .IN1(n16749), .IN2(n16750), .QN(n16746) );
  NOR2X0 U17293 ( .IN1(g3476), .IN2(n16751), .QN(n16750) );
  NAND2X0 U17294 ( .IN1(n5424), .IN2(n16744), .QN(n16751) );
  NOR2X0 U17295 ( .IN1(n5786), .IN2(n16752), .QN(n16749) );
  NOR2X0 U17296 ( .IN1(n11033), .IN2(n16753), .QN(n16752) );
  NOR2X0 U17297 ( .IN1(n5424), .IN2(n16754), .QN(n16753) );
  NAND2X0 U17298 ( .IN1(n16755), .IN2(n16756), .QN(g29265) );
  NAND2X0 U17299 ( .IN1(n16748), .IN2(g3476), .QN(n16756) );
  INVX0 U17300 ( .INP(n16745), .ZN(n16748) );
  NAND2X0 U17301 ( .IN1(n16745), .IN2(g3470), .QN(n16755) );
  NAND2X0 U17302 ( .IN1(n16757), .IN2(n16758), .QN(g29264) );
  INVX0 U17303 ( .INP(n16759), .ZN(n16758) );
  NOR2X0 U17304 ( .IN1(n16745), .IN2(n10149), .QN(n16759) );
  NAND2X0 U17305 ( .IN1(n16754), .IN2(n10963), .QN(n16745) );
  NOR2X0 U17306 ( .IN1(n16760), .IN2(n16761), .QN(n16757) );
  NOR2X0 U17307 ( .IN1(test_so4), .IN2(n16762), .QN(n16761) );
  NAND2X0 U17308 ( .IN1(n16744), .IN2(g3462), .QN(n16762) );
  NOR2X0 U17309 ( .IN1(n16754), .IN2(n11019), .QN(n16744) );
  NOR2X0 U17310 ( .IN1(n16763), .IN2(n10658), .QN(n16760) );
  NOR2X0 U17311 ( .IN1(n11033), .IN2(n16764), .QN(n16763) );
  NOR2X0 U17312 ( .IN1(n16754), .IN2(g3462), .QN(n16764) );
  NAND2X0 U17313 ( .IN1(n16765), .IN2(n13605), .QN(n16754) );
  NAND2X0 U17314 ( .IN1(n16766), .IN2(n16767), .QN(g29263) );
  NAND2X0 U17315 ( .IN1(n11073), .IN2(g3462), .QN(n16767) );
  NAND2X0 U17316 ( .IN1(n16768), .IN2(n10963), .QN(n16766) );
  NAND2X0 U17317 ( .IN1(n16769), .IN2(n16770), .QN(n16768) );
  NAND2X0 U17318 ( .IN1(test_so4), .IN2(n13603), .QN(n16770) );
  NAND2X0 U17319 ( .IN1(n16771), .IN2(n13605), .QN(n16769) );
  XOR2X1 U17320 ( .IN1(n16772), .IN2(n16773), .Q(n16771) );
  NOR2X0 U17321 ( .IN1(n16765), .IN2(n10658), .QN(n16773) );
  NOR2X0 U17322 ( .IN1(n16774), .IN2(n12450), .QN(n16765) );
  NAND2X0 U17323 ( .IN1(g3689), .IN2(g16656), .QN(n16774) );
  NAND2X0 U17324 ( .IN1(n16775), .IN2(n16776), .QN(g29262) );
  NAND2X0 U17325 ( .IN1(n3765), .IN2(n16777), .QN(n16776) );
  NAND2X0 U17326 ( .IN1(g3147), .IN2(n15923), .QN(n16777) );
  NOR2X0 U17327 ( .IN1(n16500), .IN2(n16778), .QN(n16775) );
  NOR2X0 U17328 ( .IN1(n15924), .IN2(n16779), .QN(n16778) );
  NAND2X0 U17329 ( .IN1(n16503), .IN2(g3147), .QN(n16779) );
  INVX0 U17330 ( .INP(n4210), .ZN(n16503) );
  NOR2X0 U17331 ( .IN1(n15008), .IN2(n4210), .QN(n16500) );
  NAND2X0 U17332 ( .IN1(n10593), .IN2(g4180), .QN(n4210) );
  INVX0 U17333 ( .INP(n3765), .ZN(n15008) );
  NAND2X0 U17334 ( .IN1(n16780), .IN2(n16781), .QN(g29261) );
  NAND2X0 U17335 ( .IN1(n11073), .IN2(g3129), .QN(n16781) );
  NOR2X0 U17336 ( .IN1(n16782), .IN2(n16783), .QN(n16780) );
  INVX0 U17337 ( .INP(n16784), .ZN(n16783) );
  NAND2X0 U17338 ( .IN1(n16785), .IN2(n5661), .QN(n16784) );
  NOR2X0 U17339 ( .IN1(n5661), .IN2(n16786), .QN(n16782) );
  NAND2X0 U17340 ( .IN1(n16787), .IN2(n16788), .QN(g29260) );
  NAND2X0 U17341 ( .IN1(n16789), .IN2(g3129), .QN(n16788) );
  NOR2X0 U17342 ( .IN1(n16790), .IN2(n16791), .QN(n16787) );
  NOR2X0 U17343 ( .IN1(g3125), .IN2(n16792), .QN(n16791) );
  NAND2X0 U17344 ( .IN1(n5423), .IN2(n16785), .QN(n16792) );
  NOR2X0 U17345 ( .IN1(n5781), .IN2(n16793), .QN(n16790) );
  NOR2X0 U17346 ( .IN1(n11033), .IN2(n16794), .QN(n16793) );
  NOR2X0 U17347 ( .IN1(n5423), .IN2(n16795), .QN(n16794) );
  NAND2X0 U17348 ( .IN1(n16796), .IN2(n16797), .QN(g29259) );
  NAND2X0 U17349 ( .IN1(n16789), .IN2(g3125), .QN(n16797) );
  INVX0 U17350 ( .INP(n16786), .ZN(n16789) );
  NAND2X0 U17351 ( .IN1(n16786), .IN2(g3119), .QN(n16796) );
  NAND2X0 U17352 ( .IN1(n16795), .IN2(n10963), .QN(n16786) );
  NAND2X0 U17353 ( .IN1(n16798), .IN2(n16799), .QN(g29258) );
  NAND2X0 U17354 ( .IN1(n12027), .IN2(n16795), .QN(n16799) );
  NOR2X0 U17355 ( .IN1(n11033), .IN2(n10170), .QN(n12027) );
  NOR2X0 U17356 ( .IN1(n16800), .IN2(n16801), .QN(n16798) );
  NOR2X0 U17357 ( .IN1(g3106), .IN2(n16802), .QN(n16801) );
  NAND2X0 U17358 ( .IN1(n16785), .IN2(g3111), .QN(n16802) );
  NOR2X0 U17359 ( .IN1(n16795), .IN2(n11020), .QN(n16785) );
  NOR2X0 U17360 ( .IN1(n5742), .IN2(n16803), .QN(n16800) );
  NOR2X0 U17361 ( .IN1(n11033), .IN2(n16804), .QN(n16803) );
  NOR2X0 U17362 ( .IN1(n16795), .IN2(g3111), .QN(n16804) );
  NAND2X0 U17363 ( .IN1(n16805), .IN2(n13625), .QN(n16795) );
  NAND2X0 U17364 ( .IN1(n16806), .IN2(n16807), .QN(g29257) );
  NAND2X0 U17365 ( .IN1(n11073), .IN2(g3111), .QN(n16807) );
  NAND2X0 U17366 ( .IN1(n16808), .IN2(n10964), .QN(n16806) );
  NAND2X0 U17367 ( .IN1(n16809), .IN2(n16810), .QN(n16808) );
  NAND2X0 U17368 ( .IN1(n13626), .IN2(g3106), .QN(n16810) );
  NAND2X0 U17369 ( .IN1(n16811), .IN2(n13625), .QN(n16809) );
  XOR2X1 U17370 ( .IN1(n16812), .IN2(n16813), .Q(n16811) );
  NOR2X0 U17371 ( .IN1(n16805), .IN2(n5742), .QN(n16813) );
  NOR2X0 U17372 ( .IN1(n16814), .IN2(n12442), .QN(n16805) );
  NAND2X0 U17373 ( .IN1(g3338), .IN2(g16624), .QN(n16814) );
  NAND2X0 U17374 ( .IN1(n16815), .IN2(n16816), .QN(g29256) );
  NOR2X0 U17375 ( .IN1(n16817), .IN2(n16818), .QN(n16816) );
  NOR2X0 U17376 ( .IN1(n10274), .IN2(n10851), .QN(n16818) );
  NOR2X0 U17377 ( .IN1(n11033), .IN2(n16819), .QN(n16817) );
  NAND2X0 U17378 ( .IN1(n16820), .IN2(g2735), .QN(n16819) );
  NOR2X0 U17379 ( .IN1(n2787), .IN2(n16821), .QN(n16815) );
  NOR2X0 U17380 ( .IN1(n16820), .IN2(g2735), .QN(n16821) );
  INVX0 U17381 ( .INP(n16098), .ZN(n16820) );
  NOR2X0 U17382 ( .IN1(n16822), .IN2(n10274), .QN(n16098) );
  NAND2X0 U17383 ( .IN1(n16823), .IN2(n16824), .QN(g29254) );
  NOR2X0 U17384 ( .IN1(n16825), .IN2(n16826), .QN(n16824) );
  NOR2X0 U17385 ( .IN1(n16827), .IN2(n14465), .QN(n16826) );
  NAND2X0 U17386 ( .IN1(n16828), .IN2(n10964), .QN(n14465) );
  NOR2X0 U17387 ( .IN1(n16829), .IN2(n16830), .QN(n16827) );
  NAND2X0 U17388 ( .IN1(n16831), .IN2(n16832), .QN(n16830) );
  NAND2X0 U17389 ( .IN1(n10529), .IN2(n16833), .QN(n16832) );
  INVX0 U17390 ( .INP(n16834), .ZN(n16833) );
  NOR2X0 U17391 ( .IN1(n16835), .IN2(n16836), .QN(n16834) );
  NOR2X0 U17392 ( .IN1(n10663), .IN2(n5372), .QN(n16836) );
  NOR2X0 U17393 ( .IN1(n5508), .IN2(n5787), .QN(n16835) );
  NAND2X0 U17394 ( .IN1(n5508), .IN2(n16837), .QN(n16831) );
  NAND2X0 U17395 ( .IN1(n16838), .IN2(n16839), .QN(n16837) );
  NAND2X0 U17396 ( .IN1(g2610), .IN2(g2583), .QN(n16839) );
  NAND2X0 U17397 ( .IN1(test_so66), .IN2(n5372), .QN(n16838) );
  NOR2X0 U17398 ( .IN1(n5816), .IN2(n14483), .QN(n16829) );
  NAND2X0 U17399 ( .IN1(n5372), .IN2(g2610), .QN(n14483) );
  NOR2X0 U17400 ( .IN1(n10134), .IN2(n16117), .QN(n16825) );
  INVX0 U17401 ( .INP(n16106), .ZN(n16117) );
  NOR2X0 U17402 ( .IN1(n16109), .IN2(n11020), .QN(n16106) );
  NAND2X0 U17403 ( .IN1(n16840), .IN2(n16828), .QN(n16109) );
  INVX0 U17404 ( .INP(n11309), .ZN(n16828) );
  NOR2X0 U17405 ( .IN1(n5508), .IN2(n5372), .QN(n16840) );
  NOR2X0 U17406 ( .IN1(n16841), .IN2(n16842), .QN(n16823) );
  NOR2X0 U17407 ( .IN1(n5508), .IN2(n10851), .QN(n16842) );
  NOR2X0 U17408 ( .IN1(n10594), .IN2(n11304), .QN(n16841) );
  NAND2X0 U17409 ( .IN1(n11309), .IN2(n10964), .QN(n11304) );
  NAND2X0 U17410 ( .IN1(n16843), .IN2(n16065), .QN(n11309) );
  NOR2X0 U17411 ( .IN1(n16844), .IN2(n16845), .QN(n16843) );
  NOR2X0 U17412 ( .IN1(n5609), .IN2(n16087), .QN(n16845) );
  NAND2X0 U17413 ( .IN1(n16846), .IN2(n16847), .QN(g29252) );
  NOR2X0 U17414 ( .IN1(n16848), .IN2(n16849), .QN(n16847) );
  NOR2X0 U17415 ( .IN1(n16850), .IN2(n14499), .QN(n16849) );
  NAND2X0 U17416 ( .IN1(n16851), .IN2(n10964), .QN(n14499) );
  NOR2X0 U17417 ( .IN1(n16852), .IN2(n16853), .QN(n16850) );
  NAND2X0 U17418 ( .IN1(n16854), .IN2(n16855), .QN(n16853) );
  NAND2X0 U17419 ( .IN1(n10530), .IN2(n16856), .QN(n16855) );
  INVX0 U17420 ( .INP(n16857), .ZN(n16856) );
  NOR2X0 U17421 ( .IN1(n16858), .IN2(n16859), .QN(n16857) );
  NOR2X0 U17422 ( .IN1(n5373), .IN2(n19416), .QN(n16859) );
  NOR2X0 U17423 ( .IN1(n5509), .IN2(n5789), .QN(n16858) );
  NAND2X0 U17424 ( .IN1(n5509), .IN2(n16860), .QN(n16854) );
  NAND2X0 U17425 ( .IN1(n16861), .IN2(n16862), .QN(n16860) );
  INVX0 U17426 ( .INP(n16863), .ZN(n16862) );
  NOR2X0 U17427 ( .IN1(n10530), .IN2(n5798), .QN(n16863) );
  NAND2X0 U17428 ( .IN1(n5373), .IN2(g2441), .QN(n16861) );
  NOR2X0 U17429 ( .IN1(n5814), .IN2(n14518), .QN(n16852) );
  NAND2X0 U17430 ( .IN1(n5373), .IN2(g2476), .QN(n14518) );
  NOR2X0 U17431 ( .IN1(n10136), .IN2(n16153), .QN(n16848) );
  INVX0 U17432 ( .INP(n16142), .ZN(n16153) );
  NOR2X0 U17433 ( .IN1(n16145), .IN2(n11020), .QN(n16142) );
  NAND2X0 U17434 ( .IN1(n16864), .IN2(n16851), .QN(n16145) );
  INVX0 U17435 ( .INP(n11246), .ZN(n16851) );
  NOR2X0 U17436 ( .IN1(n5509), .IN2(n5373), .QN(n16864) );
  NOR2X0 U17437 ( .IN1(n16865), .IN2(n16866), .QN(n16846) );
  NOR2X0 U17438 ( .IN1(n5509), .IN2(n10852), .QN(n16866) );
  NOR2X0 U17439 ( .IN1(n10581), .IN2(n11241), .QN(n16865) );
  NAND2X0 U17440 ( .IN1(n11246), .IN2(n10965), .QN(n11241) );
  NAND2X0 U17441 ( .IN1(n16867), .IN2(n16060), .QN(n11246) );
  NOR2X0 U17442 ( .IN1(n16844), .IN2(n16868), .QN(n16867) );
  NOR2X0 U17443 ( .IN1(n5404), .IN2(n16087), .QN(n16868) );
  NAND2X0 U17444 ( .IN1(n16869), .IN2(n16870), .QN(g29250) );
  NOR2X0 U17445 ( .IN1(n16871), .IN2(n16872), .QN(n16870) );
  NOR2X0 U17446 ( .IN1(n16873), .IN2(n14534), .QN(n16872) );
  NAND2X0 U17447 ( .IN1(n16874), .IN2(n10965), .QN(n14534) );
  NOR2X0 U17448 ( .IN1(n16875), .IN2(n16876), .QN(n16873) );
  NAND2X0 U17449 ( .IN1(n16877), .IN2(n16878), .QN(n16876) );
  NAND2X0 U17450 ( .IN1(n5511), .IN2(n16879), .QN(n16878) );
  NAND2X0 U17451 ( .IN1(n16880), .IN2(n16881), .QN(n16879) );
  NAND2X0 U17452 ( .IN1(n5375), .IN2(g2307), .QN(n16881) );
  NAND2X0 U17453 ( .IN1(test_so21), .IN2(g2315), .QN(n16880) );
  NAND2X0 U17454 ( .IN1(n16882), .IN2(n10640), .QN(n16877) );
  INVX0 U17455 ( .INP(n16883), .ZN(n16882) );
  NOR2X0 U17456 ( .IN1(n16884), .IN2(n16885), .QN(n16883) );
  NOR2X0 U17457 ( .IN1(n5375), .IN2(n19412), .QN(n16885) );
  NOR2X0 U17458 ( .IN1(n5511), .IN2(n5794), .QN(n16884) );
  NOR2X0 U17459 ( .IN1(n5815), .IN2(n14553), .QN(n16875) );
  NAND2X0 U17460 ( .IN1(test_so21), .IN2(n5375), .QN(n14553) );
  NOR2X0 U17461 ( .IN1(n10152), .IN2(n16189), .QN(n16871) );
  INVX0 U17462 ( .INP(n16178), .ZN(n16189) );
  NOR2X0 U17463 ( .IN1(n16181), .IN2(n11021), .QN(n16178) );
  NAND2X0 U17464 ( .IN1(n16886), .IN2(n16874), .QN(n16181) );
  INVX0 U17465 ( .INP(n11260), .ZN(n16874) );
  NOR2X0 U17466 ( .IN1(n5511), .IN2(n5375), .QN(n16886) );
  NOR2X0 U17467 ( .IN1(n16887), .IN2(n16888), .QN(n16869) );
  NOR2X0 U17468 ( .IN1(n5511), .IN2(n10853), .QN(n16888) );
  NOR2X0 U17469 ( .IN1(n10319), .IN2(n11255), .QN(n16887) );
  NAND2X0 U17470 ( .IN1(n11260), .IN2(n10965), .QN(n11255) );
  NAND2X0 U17471 ( .IN1(n16889), .IN2(n16890), .QN(n11260) );
  NAND2X0 U17472 ( .IN1(n12398), .IN2(g2807), .QN(n16890) );
  NAND2X0 U17473 ( .IN1(n16891), .IN2(n16892), .QN(g29248) );
  NOR2X0 U17474 ( .IN1(n16893), .IN2(n16894), .QN(n16892) );
  NOR2X0 U17475 ( .IN1(n16895), .IN2(n14569), .QN(n16894) );
  NAND2X0 U17476 ( .IN1(n16896), .IN2(n10966), .QN(n14569) );
  NOR2X0 U17477 ( .IN1(n16897), .IN2(n16898), .QN(n16895) );
  NAND2X0 U17478 ( .IN1(n16899), .IN2(n16900), .QN(n16898) );
  NAND2X0 U17479 ( .IN1(n10532), .IN2(n16901), .QN(n16900) );
  INVX0 U17480 ( .INP(n16902), .ZN(n16901) );
  NOR2X0 U17481 ( .IN1(n16903), .IN2(n16904), .QN(n16902) );
  NOR2X0 U17482 ( .IN1(n5376), .IN2(n19408), .QN(n16904) );
  NOR2X0 U17483 ( .IN1(n5512), .IN2(n5788), .QN(n16903) );
  NAND2X0 U17484 ( .IN1(n5512), .IN2(n16905), .QN(n16899) );
  NAND2X0 U17485 ( .IN1(n16906), .IN2(n16907), .QN(n16905) );
  NAND2X0 U17486 ( .IN1(g2208), .IN2(g2181), .QN(n16907) );
  NAND2X0 U17487 ( .IN1(n5376), .IN2(g2173), .QN(n16906) );
  NOR2X0 U17488 ( .IN1(n5812), .IN2(n14588), .QN(n16897) );
  NAND2X0 U17489 ( .IN1(n5376), .IN2(g2208), .QN(n14588) );
  NOR2X0 U17490 ( .IN1(n10158), .IN2(n16225), .QN(n16893) );
  INVX0 U17491 ( .INP(n16214), .ZN(n16225) );
  NOR2X0 U17492 ( .IN1(n16217), .IN2(n11021), .QN(n16214) );
  NAND2X0 U17493 ( .IN1(n16908), .IN2(n16896), .QN(n16217) );
  INVX0 U17494 ( .INP(n11495), .ZN(n16896) );
  NOR2X0 U17495 ( .IN1(n5512), .IN2(n5376), .QN(n16908) );
  NOR2X0 U17496 ( .IN1(n16909), .IN2(n16910), .QN(n16891) );
  NOR2X0 U17497 ( .IN1(n5512), .IN2(n10853), .QN(n16910) );
  NOR2X0 U17498 ( .IN1(n10315), .IN2(n11490), .QN(n16909) );
  NAND2X0 U17499 ( .IN1(n11495), .IN2(n10966), .QN(n11490) );
  NAND2X0 U17500 ( .IN1(n16911), .IN2(n16064), .QN(n11495) );
  NOR2X0 U17501 ( .IN1(n16844), .IN2(n16912), .QN(n16911) );
  NOR2X0 U17502 ( .IN1(n5545), .IN2(n16087), .QN(n16912) );
  NAND2X0 U17503 ( .IN1(n16913), .IN2(n16914), .QN(g29247) );
  NAND2X0 U17504 ( .IN1(n16915), .IN2(g2079), .QN(n16914) );
  NAND2X0 U17505 ( .IN1(n16916), .IN2(n10966), .QN(n16915) );
  NAND2X0 U17506 ( .IN1(n16917), .IN2(n11478), .QN(n16916) );
  NAND2X0 U17507 ( .IN1(test_so78), .IN2(n14626), .QN(n11478) );
  NAND2X0 U17508 ( .IN1(test_so78), .IN2(n16918), .QN(n16913) );
  NAND2X0 U17509 ( .IN1(n14605), .IN2(n16919), .QN(n16918) );
  NAND2X0 U17510 ( .IN1(n4425), .IN2(n10967), .QN(n16919) );
  NAND2X0 U17511 ( .IN1(n16920), .IN2(n16921), .QN(g29246) );
  NOR2X0 U17512 ( .IN1(n16922), .IN2(n16923), .QN(n16921) );
  NOR2X0 U17513 ( .IN1(n16924), .IN2(n14606), .QN(n16923) );
  NAND2X0 U17514 ( .IN1(n16917), .IN2(n10967), .QN(n14606) );
  NOR2X0 U17515 ( .IN1(n16925), .IN2(n16926), .QN(n16924) );
  NAND2X0 U17516 ( .IN1(n16927), .IN2(n16928), .QN(n16926) );
  NAND2X0 U17517 ( .IN1(n10528), .IN2(n16929), .QN(n16928) );
  INVX0 U17518 ( .INP(n16930), .ZN(n16929) );
  NOR2X0 U17519 ( .IN1(n16931), .IN2(n16932), .QN(n16930) );
  NOR2X0 U17520 ( .IN1(n5371), .IN2(n19413), .QN(n16932) );
  NOR2X0 U17521 ( .IN1(n5507), .IN2(n5790), .QN(n16931) );
  NAND2X0 U17522 ( .IN1(n5507), .IN2(n16933), .QN(n16927) );
  NAND2X0 U17523 ( .IN1(n16934), .IN2(n16935), .QN(n16933) );
  NAND2X0 U17524 ( .IN1(g2051), .IN2(g2024), .QN(n16935) );
  NAND2X0 U17525 ( .IN1(n5371), .IN2(g2016), .QN(n16934) );
  NOR2X0 U17526 ( .IN1(n5818), .IN2(n14626), .QN(n16925) );
  NAND2X0 U17527 ( .IN1(n5371), .IN2(g2051), .QN(n14626) );
  NOR2X0 U17528 ( .IN1(n10217), .IN2(n16262), .QN(n16922) );
  INVX0 U17529 ( .INP(n16250), .ZN(n16262) );
  NOR2X0 U17530 ( .IN1(n16253), .IN2(n11021), .QN(n16250) );
  NAND2X0 U17531 ( .IN1(n16936), .IN2(n16917), .QN(n16253) );
  INVX0 U17532 ( .INP(n14598), .ZN(n16917) );
  NOR2X0 U17533 ( .IN1(n5507), .IN2(n5371), .QN(n16936) );
  NOR2X0 U17534 ( .IN1(n16937), .IN2(n16938), .QN(n16920) );
  NOR2X0 U17535 ( .IN1(n5507), .IN2(n10854), .QN(n16938) );
  NOR2X0 U17536 ( .IN1(n10595), .IN2(n14605), .QN(n16937) );
  NAND2X0 U17537 ( .IN1(n14598), .IN2(n10967), .QN(n14605) );
  NAND2X0 U17538 ( .IN1(n16939), .IN2(n16065), .QN(n14598) );
  NOR2X0 U17539 ( .IN1(n16844), .IN2(n16940), .QN(n16939) );
  NOR2X0 U17540 ( .IN1(n5610), .IN2(n16087), .QN(n16940) );
  NAND2X0 U17541 ( .IN1(n16941), .IN2(n16942), .QN(g29244) );
  NOR2X0 U17542 ( .IN1(n16943), .IN2(n16944), .QN(n16942) );
  NOR2X0 U17543 ( .IN1(n16945), .IN2(n14642), .QN(n16944) );
  NAND2X0 U17544 ( .IN1(n16946), .IN2(n10967), .QN(n14642) );
  NOR2X0 U17545 ( .IN1(n16947), .IN2(n16948), .QN(n16945) );
  NAND2X0 U17546 ( .IN1(n16949), .IN2(n16950), .QN(n16948) );
  NAND2X0 U17547 ( .IN1(n10531), .IN2(n16951), .QN(n16950) );
  INVX0 U17548 ( .INP(n16952), .ZN(n16951) );
  NOR2X0 U17549 ( .IN1(n16953), .IN2(n16954), .QN(n16952) );
  NOR2X0 U17550 ( .IN1(n5374), .IN2(n19415), .QN(n16954) );
  NOR2X0 U17551 ( .IN1(n5510), .IN2(n5793), .QN(n16953) );
  NAND2X0 U17552 ( .IN1(n5510), .IN2(n16955), .QN(n16949) );
  NAND2X0 U17553 ( .IN1(n16956), .IN2(n16957), .QN(n16955) );
  NAND2X0 U17554 ( .IN1(g1917), .IN2(g1890), .QN(n16957) );
  NAND2X0 U17555 ( .IN1(n5374), .IN2(g1882), .QN(n16956) );
  NOR2X0 U17556 ( .IN1(n5813), .IN2(n14662), .QN(n16947) );
  NAND2X0 U17557 ( .IN1(n5374), .IN2(g1917), .QN(n14662) );
  NOR2X0 U17558 ( .IN1(n10144), .IN2(n16299), .QN(n16943) );
  INVX0 U17559 ( .INP(n16287), .ZN(n16299) );
  NOR2X0 U17560 ( .IN1(n16290), .IN2(n11021), .QN(n16287) );
  NAND2X0 U17561 ( .IN1(n16958), .IN2(n16946), .QN(n16290) );
  INVX0 U17562 ( .INP(n11319), .ZN(n16946) );
  NOR2X0 U17563 ( .IN1(n5510), .IN2(n5374), .QN(n16958) );
  NOR2X0 U17564 ( .IN1(n16959), .IN2(n16960), .QN(n16941) );
  NOR2X0 U17565 ( .IN1(n5510), .IN2(n10855), .QN(n16960) );
  NOR2X0 U17566 ( .IN1(n10669), .IN2(n11314), .QN(n16959) );
  NAND2X0 U17567 ( .IN1(n11319), .IN2(n10967), .QN(n11314) );
  NAND2X0 U17568 ( .IN1(n16961), .IN2(n16060), .QN(n11319) );
  NOR2X0 U17569 ( .IN1(n16844), .IN2(n16962), .QN(n16961) );
  NOR2X0 U17570 ( .IN1(n5403), .IN2(n16087), .QN(n16962) );
  NAND2X0 U17571 ( .IN1(n16963), .IN2(n16964), .QN(g29242) );
  NOR2X0 U17572 ( .IN1(n16965), .IN2(n16966), .QN(n16964) );
  NOR2X0 U17573 ( .IN1(n16967), .IN2(n14678), .QN(n16966) );
  NAND2X0 U17574 ( .IN1(n16968), .IN2(n10967), .QN(n14678) );
  NOR2X0 U17575 ( .IN1(n16969), .IN2(n16970), .QN(n16967) );
  NAND2X0 U17576 ( .IN1(n16971), .IN2(n16972), .QN(n16970) );
  NAND2X0 U17577 ( .IN1(n5359), .IN2(n16973), .QN(n16972) );
  NAND2X0 U17578 ( .IN1(n16974), .IN2(n16975), .QN(n16973) );
  NAND2X0 U17579 ( .IN1(g1783), .IN2(g1756), .QN(n16975) );
  NAND2X0 U17580 ( .IN1(n5602), .IN2(g1748), .QN(n16974) );
  NAND2X0 U17581 ( .IN1(n5596), .IN2(n16976), .QN(n16971) );
  INVX0 U17582 ( .INP(n16977), .ZN(n16976) );
  NOR2X0 U17583 ( .IN1(n16978), .IN2(n16979), .QN(n16977) );
  NOR2X0 U17584 ( .IN1(n5359), .IN2(n5795), .QN(n16979) );
  NOR2X0 U17585 ( .IN1(n5602), .IN2(n5797), .QN(n16978) );
  NOR2X0 U17586 ( .IN1(n5817), .IN2(n14696), .QN(n16969) );
  NAND2X0 U17587 ( .IN1(n5602), .IN2(g1783), .QN(n14696) );
  NOR2X0 U17588 ( .IN1(n10208), .IN2(n16335), .QN(n16965) );
  INVX0 U17589 ( .INP(n16324), .ZN(n16335) );
  NOR2X0 U17590 ( .IN1(n16327), .IN2(n11021), .QN(n16324) );
  NAND2X0 U17591 ( .IN1(n16980), .IN2(n16968), .QN(n16327) );
  INVX0 U17592 ( .INP(n11230), .ZN(n16968) );
  NOR2X0 U17593 ( .IN1(n5602), .IN2(n5359), .QN(n16980) );
  NOR2X0 U17594 ( .IN1(n16981), .IN2(n16982), .QN(n16963) );
  NOR2X0 U17595 ( .IN1(n5359), .IN2(n10855), .QN(n16982) );
  NOR2X0 U17596 ( .IN1(n10317), .IN2(n11225), .QN(n16981) );
  NAND2X0 U17597 ( .IN1(n11230), .IN2(n10967), .QN(n11225) );
  NAND2X0 U17598 ( .IN1(n16889), .IN2(n16983), .QN(n11230) );
  NAND2X0 U17599 ( .IN1(n12398), .IN2(g2775), .QN(n16983) );
  INVX0 U17600 ( .INP(n16087), .ZN(n12398) );
  NOR2X0 U17601 ( .IN1(n4411), .IN2(n16844), .QN(n16889) );
  NAND2X0 U17602 ( .IN1(n5465), .IN2(g2715), .QN(n4411) );
  NAND2X0 U17603 ( .IN1(n16984), .IN2(n16985), .QN(g29240) );
  NOR2X0 U17604 ( .IN1(n16986), .IN2(n16987), .QN(n16985) );
  NOR2X0 U17605 ( .IN1(n10321), .IN2(n11471), .QN(n16987) );
  NAND2X0 U17606 ( .IN1(n11476), .IN2(n10968), .QN(n11471) );
  NOR2X0 U17607 ( .IN1(n16988), .IN2(n14712), .QN(n16986) );
  NAND2X0 U17608 ( .IN1(n16989), .IN2(n10968), .QN(n14712) );
  NOR2X0 U17609 ( .IN1(n16990), .IN2(n16991), .QN(n16988) );
  NAND2X0 U17610 ( .IN1(n16992), .IN2(n16993), .QN(n16991) );
  NAND2X0 U17611 ( .IN1(n1418), .IN2(g1600), .QN(n16993) );
  INVX0 U17612 ( .INP(n14733), .ZN(n1418) );
  NAND2X0 U17613 ( .IN1(test_so94), .IN2(n5370), .QN(n14733) );
  NAND2X0 U17614 ( .IN1(g25167), .IN2(g1620), .QN(n16992) );
  INVX0 U17615 ( .INP(n16994), .ZN(n16990) );
  NOR2X0 U17616 ( .IN1(n16995), .IN2(n16996), .QN(n16994) );
  NOR2X0 U17617 ( .IN1(n16997), .IN2(g1657), .QN(n16996) );
  NAND2X0 U17618 ( .IN1(g1612), .IN2(n5370), .QN(n16997) );
  NOR2X0 U17619 ( .IN1(n16998), .IN2(test_so94), .QN(n16995) );
  NOR2X0 U17620 ( .IN1(n16999), .IN2(n17000), .QN(n16998) );
  NOR2X0 U17621 ( .IN1(n5370), .IN2(n19414), .QN(n17000) );
  NOR2X0 U17622 ( .IN1(n5525), .IN2(n5792), .QN(n16999) );
  NOR2X0 U17623 ( .IN1(n17001), .IN2(n17002), .QN(n16984) );
  NOR2X0 U17624 ( .IN1(n5525), .IN2(n10856), .QN(n17002) );
  NOR2X0 U17625 ( .IN1(n10135), .IN2(n16363), .QN(n17001) );
  NAND2X0 U17626 ( .IN1(n17003), .IN2(n16989), .QN(n16363) );
  INVX0 U17627 ( .INP(n11476), .ZN(n16989) );
  NAND2X0 U17628 ( .IN1(n17004), .IN2(n16064), .QN(n11476) );
  NOR2X0 U17629 ( .IN1(g2715), .IN2(g2719), .QN(n16064) );
  NOR2X0 U17630 ( .IN1(n16844), .IN2(n17005), .QN(n17004) );
  NOR2X0 U17631 ( .IN1(n5544), .IN2(n16087), .QN(n17005) );
  NOR2X0 U17632 ( .IN1(n4388), .IN2(n16087), .QN(n16844) );
  NAND2X0 U17633 ( .IN1(n5301), .IN2(n10274), .QN(n16087) );
  NOR2X0 U17634 ( .IN1(n5525), .IN2(n5370), .QN(n17003) );
  NAND2X0 U17635 ( .IN1(n17006), .IN2(n17007), .QN(g29239) );
  NAND2X0 U17636 ( .IN1(n11073), .IN2(g1478), .QN(n17007) );
  NAND2X0 U17637 ( .IN1(n17008), .IN2(n10968), .QN(n17006) );
  NAND2X0 U17638 ( .IN1(n17009), .IN2(n17010), .QN(n17008) );
  NAND2X0 U17639 ( .IN1(n17011), .IN2(n17012), .QN(n17010) );
  NOR2X0 U17640 ( .IN1(n17013), .IN2(n17014), .QN(n17011) );
  NAND2X0 U17641 ( .IN1(n17015), .IN2(g1454), .QN(n17009) );
  NAND2X0 U17642 ( .IN1(n17016), .IN2(n17014), .QN(n17015) );
  XOR2X1 U17643 ( .IN1(n5343), .IN2(n17017), .Q(n17014) );
  INVX0 U17644 ( .INP(n17013), .ZN(n17016) );
  NAND2X0 U17645 ( .IN1(n17018), .IN2(n17019), .QN(g29238) );
  NAND2X0 U17646 ( .IN1(n17020), .IN2(g1484), .QN(n17019) );
  NOR2X0 U17647 ( .IN1(n17021), .IN2(n17022), .QN(n17018) );
  NOR2X0 U17648 ( .IN1(n11033), .IN2(n17023), .QN(n17022) );
  NAND2X0 U17649 ( .IN1(n17024), .IN2(n17025), .QN(n17023) );
  NAND2X0 U17650 ( .IN1(n5865), .IN2(n17026), .QN(n17025) );
  NAND2X0 U17651 ( .IN1(n17027), .IN2(n17012), .QN(n17026) );
  XOR2X1 U17652 ( .IN1(g1300), .IN2(n17017), .Q(n17024) );
  NOR2X0 U17653 ( .IN1(n5290), .IN2(n10856), .QN(n17021) );
  NAND2X0 U17654 ( .IN1(n17028), .IN2(n17029), .QN(g29237) );
  NAND2X0 U17655 ( .IN1(n11073), .IN2(g1448), .QN(n17029) );
  NAND2X0 U17656 ( .IN1(n17030), .IN2(n10968), .QN(n17028) );
  NAND2X0 U17657 ( .IN1(n17031), .IN2(n17032), .QN(n17030) );
  NAND2X0 U17658 ( .IN1(n17033), .IN2(n17034), .QN(n17032) );
  NOR2X0 U17659 ( .IN1(n10244), .IN2(n17035), .QN(n17034) );
  NOR2X0 U17660 ( .IN1(n17036), .IN2(n17037), .QN(n17033) );
  NAND2X0 U17661 ( .IN1(n17038), .IN2(g1467), .QN(n17031) );
  INVX0 U17662 ( .INP(n17039), .ZN(n17038) );
  NOR2X0 U17663 ( .IN1(n17040), .IN2(n17035), .QN(n17039) );
  NAND2X0 U17664 ( .IN1(g13272), .IN2(n17037), .QN(n17040) );
  XNOR2X1 U17665 ( .IN1(g1472), .IN2(n17017), .Q(n17037) );
  NAND2X0 U17666 ( .IN1(n17041), .IN2(n17042), .QN(g29236) );
  NAND2X0 U17667 ( .IN1(n11073), .IN2(g1442), .QN(n17042) );
  NAND2X0 U17668 ( .IN1(n17043), .IN2(n10968), .QN(n17041) );
  NAND2X0 U17669 ( .IN1(n17044), .IN2(n17045), .QN(n17043) );
  NAND2X0 U17670 ( .IN1(n17046), .IN2(n17047), .QN(n17045) );
  NAND2X0 U17671 ( .IN1(n5696), .IN2(n17048), .QN(n17047) );
  NAND2X0 U17672 ( .IN1(n17049), .IN2(n17012), .QN(n17048) );
  INVX0 U17673 ( .INP(n17036), .ZN(n17012) );
  NAND2X0 U17674 ( .IN1(n5850), .IN2(n10536), .QN(n17036) );
  INVX0 U17675 ( .INP(n17050), .ZN(n17049) );
  XOR2X1 U17676 ( .IN1(g1478), .IN2(n17017), .Q(n17046) );
  INVX0 U17677 ( .INP(n17051), .ZN(n17017) );
  NAND2X0 U17678 ( .IN1(n14746), .IN2(DFF_1092_n1), .QN(n17051) );
  NAND2X0 U17679 ( .IN1(n17050), .IN2(g1437), .QN(n17044) );
  NAND2X0 U17680 ( .IN1(n17052), .IN2(n17053), .QN(g29235) );
  NAND2X0 U17681 ( .IN1(n11077), .IN2(g1252), .QN(n17053) );
  NOR2X0 U17682 ( .IN1(n17054), .IN2(n17055), .QN(n17052) );
  NOR2X0 U17683 ( .IN1(g1256), .IN2(n17056), .QN(n17055) );
  NOR2X0 U17684 ( .IN1(n5558), .IN2(n17057), .QN(n17054) );
  NAND2X0 U17685 ( .IN1(n14133), .IN2(n17056), .QN(n17057) );
  INVX0 U17686 ( .INP(n4178), .ZN(n17056) );
  NAND2X0 U17687 ( .IN1(n17058), .IN2(n17059), .QN(g29234) );
  NAND2X0 U17688 ( .IN1(n17060), .IN2(n17061), .QN(n17059) );
  INVX0 U17689 ( .INP(n17062), .ZN(n17061) );
  NOR2X0 U17690 ( .IN1(n17063), .IN2(n17064), .QN(n17060) );
  NOR2X0 U17691 ( .IN1(n17065), .IN2(n17066), .QN(n17058) );
  NOR2X0 U17692 ( .IN1(n11052), .IN2(n17067), .QN(n17066) );
  NAND2X0 U17693 ( .IN1(test_so90), .IN2(n17068), .QN(n17067) );
  NAND2X0 U17694 ( .IN1(n17069), .IN2(n17064), .QN(n17068) );
  XOR2X1 U17695 ( .IN1(n17070), .IN2(g1105), .Q(n17064) );
  INVX0 U17696 ( .INP(n17063), .ZN(n17069) );
  NOR2X0 U17697 ( .IN1(n5328), .IN2(n10857), .QN(n17065) );
  NAND2X0 U17698 ( .IN1(n17071), .IN2(n17072), .QN(g29233) );
  NAND2X0 U17699 ( .IN1(n17073), .IN2(g1141), .QN(n17072) );
  NOR2X0 U17700 ( .IN1(n17074), .IN2(n17075), .QN(n17071) );
  NOR2X0 U17701 ( .IN1(n11028), .IN2(n17076), .QN(n17075) );
  NAND2X0 U17702 ( .IN1(n17077), .IN2(n17078), .QN(n17076) );
  NAND2X0 U17703 ( .IN1(n5691), .IN2(n17079), .QN(n17078) );
  NAND2X0 U17704 ( .IN1(n17080), .IN2(n17081), .QN(n17079) );
  NOR2X0 U17705 ( .IN1(test_so7), .IN2(g1146), .QN(n17080) );
  XOR2X1 U17706 ( .IN1(n17070), .IN2(n5341), .Q(n17077) );
  NOR2X0 U17707 ( .IN1(n5329), .IN2(n10857), .QN(n17074) );
  NAND2X0 U17708 ( .IN1(n17082), .IN2(n17083), .QN(g29232) );
  NAND2X0 U17709 ( .IN1(n17084), .IN2(n17085), .QN(n17083) );
  NOR2X0 U17710 ( .IN1(n5599), .IN2(n17062), .QN(n17085) );
  NOR2X0 U17711 ( .IN1(n17086), .IN2(n17087), .QN(n17084) );
  NOR2X0 U17712 ( .IN1(n17088), .IN2(n17089), .QN(n17082) );
  NOR2X0 U17713 ( .IN1(n11038), .IN2(n17090), .QN(n17089) );
  INVX0 U17714 ( .INP(n17091), .ZN(n17090) );
  NOR2X0 U17715 ( .IN1(n17092), .IN2(n5692), .QN(n17091) );
  NOR2X0 U17716 ( .IN1(n17093), .IN2(n17086), .QN(n17092) );
  NAND2X0 U17717 ( .IN1(g1183), .IN2(n17087), .QN(n17093) );
  XNOR2X1 U17718 ( .IN1(n17070), .IN2(n5329), .Q(n17087) );
  NOR2X0 U17719 ( .IN1(n5478), .IN2(n10857), .QN(n17088) );
  NAND2X0 U17720 ( .IN1(n17094), .IN2(n17095), .QN(g29231) );
  NAND2X0 U17721 ( .IN1(n17096), .IN2(n17097), .QN(n17095) );
  NOR2X0 U17722 ( .IN1(g1183), .IN2(n17062), .QN(n17097) );
  NAND2X0 U17723 ( .IN1(n17098), .IN2(n5851), .QN(n17062) );
  NOR2X0 U17724 ( .IN1(n17086), .IN2(n17099), .QN(n17096) );
  INVX0 U17725 ( .INP(n17100), .ZN(n17094) );
  NAND2X0 U17726 ( .IN1(n17101), .IN2(n17102), .QN(n17100) );
  NAND2X0 U17727 ( .IN1(n10930), .IN2(n17103), .QN(n17102) );
  NOR2X0 U17728 ( .IN1(n17104), .IN2(n5697), .QN(n17103) );
  NOR2X0 U17729 ( .IN1(n17105), .IN2(n17086), .QN(n17104) );
  NAND2X0 U17730 ( .IN1(n17099), .IN2(n5599), .QN(n17105) );
  XNOR2X1 U17731 ( .IN1(n17070), .IN2(n5328), .Q(n17099) );
  NAND2X0 U17732 ( .IN1(n12087), .IN2(DFF_24_n1), .QN(n17070) );
  NAND2X0 U17733 ( .IN1(n11061), .IN2(test_so7), .QN(n17101) );
  NAND2X0 U17734 ( .IN1(n17106), .IN2(n17107), .QN(g29230) );
  NAND2X0 U17735 ( .IN1(n11060), .IN2(g907), .QN(n17107) );
  NOR2X0 U17736 ( .IN1(n17108), .IN2(n17109), .QN(n17106) );
  NOR2X0 U17737 ( .IN1(g911), .IN2(n17110), .QN(n17109) );
  NOR2X0 U17738 ( .IN1(n5559), .IN2(n17111), .QN(n17108) );
  NAND2X0 U17739 ( .IN1(n14152), .IN2(n17110), .QN(n17111) );
  INVX0 U17740 ( .INP(n4196), .ZN(n17110) );
  NAND2X0 U17741 ( .IN1(n17112), .IN2(n17113), .QN(g29229) );
  NAND2X0 U17742 ( .IN1(n11060), .IN2(g827), .QN(n17113) );
  NOR2X0 U17743 ( .IN1(n17114), .IN2(n17115), .QN(n17112) );
  NOR2X0 U17744 ( .IN1(g723), .IN2(n17116), .QN(n17115) );
  NAND2X0 U17745 ( .IN1(n4516), .IN2(n17117), .QN(n17116) );
  NOR2X0 U17746 ( .IN1(n5826), .IN2(n17118), .QN(n17114) );
  INVX0 U17747 ( .INP(n4517), .ZN(n17118) );
  NAND2X0 U17748 ( .IN1(n17119), .IN2(n17120), .QN(g29228) );
  NAND2X0 U17749 ( .IN1(n2404), .IN2(n17121), .QN(n17120) );
  XNOR2X1 U17750 ( .IN1(test_so60), .IN2(n16481), .Q(n17121) );
  NAND2X0 U17751 ( .IN1(n16496), .IN2(n17122), .QN(n16481) );
  NAND2X0 U17752 ( .IN1(n5482), .IN2(g12184), .QN(n17122) );
  INVX0 U17753 ( .INP(n14961), .ZN(n16496) );
  NAND2X0 U17754 ( .IN1(n17123), .IN2(n17124), .QN(n14961) );
  NOR2X0 U17755 ( .IN1(n17125), .IN2(n17126), .QN(n17124) );
  NOR2X0 U17756 ( .IN1(g655), .IN2(n17127), .QN(n17126) );
  NAND2X0 U17757 ( .IN1(n10312), .IN2(n10183), .QN(n17127) );
  NOR2X0 U17758 ( .IN1(n10313), .IN2(n17128), .QN(n17125) );
  NAND2X0 U17759 ( .IN1(g753), .IN2(g718), .QN(n17128) );
  NOR2X0 U17760 ( .IN1(n17129), .IN2(n17130), .QN(n17123) );
  NOR2X0 U17761 ( .IN1(n5479), .IN2(n10212), .QN(n17129) );
  NAND2X0 U17762 ( .IN1(n11060), .IN2(g736), .QN(n17119) );
  NAND2X0 U17763 ( .IN1(n17131), .IN2(n17132), .QN(g29227) );
  NAND2X0 U17764 ( .IN1(n11058), .IN2(g676), .QN(n17132) );
  NOR2X0 U17765 ( .IN1(n17133), .IN2(n17134), .QN(n17131) );
  INVX0 U17766 ( .INP(n17135), .ZN(n17134) );
  NAND2X0 U17767 ( .IN1(test_so70), .IN2(n4524), .QN(n17135) );
  NOR2X0 U17768 ( .IN1(test_so70), .IN2(n17136), .QN(n17133) );
  NAND2X0 U17769 ( .IN1(n4523), .IN2(n17137), .QN(n17136) );
  NAND2X0 U17770 ( .IN1(n17138), .IN2(n17139), .QN(g29226) );
  NAND2X0 U17771 ( .IN1(n11058), .IN2(g671), .QN(n17139) );
  NOR2X0 U17772 ( .IN1(n17140), .IN2(n17141), .QN(n17138) );
  NOR2X0 U17773 ( .IN1(g676), .IN2(n17142), .QN(n17141) );
  NAND2X0 U17774 ( .IN1(n4526), .IN2(n17137), .QN(n17142) );
  INVX0 U17775 ( .INP(n17143), .ZN(n17137) );
  NOR2X0 U17776 ( .IN1(n5751), .IN2(n17144), .QN(n17140) );
  NAND2X0 U17777 ( .IN1(n4525), .IN2(n17145), .QN(n17144) );
  INVX0 U17778 ( .INP(n4526), .ZN(n17145) );
  NAND2X0 U17779 ( .IN1(n17146), .IN2(n17147), .QN(g29225) );
  NAND2X0 U17780 ( .IN1(n17148), .IN2(n4525), .QN(n17147) );
  NOR2X0 U17781 ( .IN1(n17143), .IN2(n11019), .QN(n4525) );
  NAND2X0 U17782 ( .IN1(g703), .IN2(n17149), .QN(n17143) );
  NAND2X0 U17783 ( .IN1(n17150), .IN2(n17151), .QN(n17149) );
  NOR2X0 U17784 ( .IN1(n10233), .IN2(n154), .QN(n17151) );
  NOR2X0 U17785 ( .IN1(n17152), .IN2(n4535), .QN(n17150) );
  XOR2X1 U17786 ( .IN1(n10312), .IN2(n10313), .Q(n4535) );
  XOR2X1 U17787 ( .IN1(n154), .IN2(n10138), .Q(n17148) );
  NAND2X0 U17788 ( .IN1(n11059), .IN2(g667), .QN(n17146) );
  NAND2X0 U17789 ( .IN1(n17153), .IN2(n17154), .QN(g29224) );
  NAND2X0 U17790 ( .IN1(n11060), .IN2(g572), .QN(n17154) );
  NOR2X0 U17791 ( .IN1(n17155), .IN2(n17156), .QN(n17153) );
  NOR2X0 U17792 ( .IN1(g586), .IN2(n17157), .QN(n17156) );
  NOR2X0 U17793 ( .IN1(n5336), .IN2(n17158), .QN(n17155) );
  NAND2X0 U17794 ( .IN1(n2421), .IN2(n17157), .QN(n17158) );
  INVX0 U17795 ( .INP(n4201), .ZN(n17157) );
  NAND2X0 U17796 ( .IN1(n17159), .IN2(n17160), .QN(g29223) );
  NAND2X0 U17797 ( .IN1(n17161), .IN2(n5708), .QN(n17160) );
  NOR2X0 U17798 ( .IN1(n17162), .IN2(n17163), .QN(n17159) );
  NOR2X0 U17799 ( .IN1(n11033), .IN2(n17164), .QN(n17163) );
  NOR2X0 U17800 ( .IN1(n17165), .IN2(n4962), .QN(n17164) );
  NOR2X0 U17801 ( .IN1(n5708), .IN2(n17161), .QN(n17165) );
  INVX0 U17802 ( .INP(n17166), .ZN(n17161) );
  NAND2X0 U17803 ( .IN1(n17167), .IN2(g482), .QN(n17166) );
  NOR2X0 U17804 ( .IN1(n5820), .IN2(n10858), .QN(n17162) );
  NAND2X0 U17805 ( .IN1(n17168), .IN2(n17169), .QN(g29222) );
  NAND2X0 U17806 ( .IN1(n17170), .IN2(g411), .QN(n17169) );
  NOR2X0 U17807 ( .IN1(n17171), .IN2(n17172), .QN(n17168) );
  NOR2X0 U17808 ( .IN1(g417), .IN2(n17173), .QN(n17172) );
  NAND2X0 U17809 ( .IN1(n17174), .IN2(n3676), .QN(n17173) );
  NOR2X0 U17810 ( .IN1(n5358), .IN2(n17175), .QN(n17171) );
  NOR2X0 U17811 ( .IN1(n11034), .IN2(n17176), .QN(n17175) );
  NOR2X0 U17812 ( .IN1(n3676), .IN2(n17177), .QN(n17176) );
  XOR2X1 U17813 ( .IN1(g417), .IN2(n17178), .Q(n3676) );
  NOR2X0 U17814 ( .IN1(n17179), .IN2(n17180), .QN(n17178) );
  NOR2X0 U17815 ( .IN1(g392), .IN2(n17181), .QN(n17180) );
  NOR2X0 U17816 ( .IN1(n17182), .IN2(n17183), .QN(n17181) );
  NOR2X0 U17817 ( .IN1(n10245), .IN2(g405), .QN(n17183) );
  NOR2X0 U17818 ( .IN1(n10247), .IN2(n10246), .QN(n17182) );
  NOR2X0 U17819 ( .IN1(n10272), .IN2(n17184), .QN(n17179) );
  NOR2X0 U17820 ( .IN1(n17185), .IN2(n17186), .QN(n17184) );
  NOR2X0 U17821 ( .IN1(n10247), .IN2(n10228), .QN(n17186) );
  NOR2X0 U17822 ( .IN1(n10246), .IN2(g405), .QN(n17185) );
  NAND2X0 U17823 ( .IN1(n17187), .IN2(n17188), .QN(g28105) );
  NAND2X0 U17824 ( .IN1(n13467), .IN2(g5011), .QN(n17188) );
  NOR2X0 U17825 ( .IN1(n17189), .IN2(n17190), .QN(n17187) );
  NOR2X0 U17826 ( .IN1(n11034), .IN2(n17191), .QN(n17190) );
  NAND2X0 U17827 ( .IN1(n13464), .IN2(n16532), .QN(n17191) );
  NAND2X0 U17828 ( .IN1(n17192), .IN2(n17193), .QN(n16532) );
  NOR2X0 U17829 ( .IN1(n17194), .IN2(n17195), .QN(n17193) );
  NOR2X0 U17830 ( .IN1(n17196), .IN2(n17197), .QN(n17195) );
  NOR2X0 U17831 ( .IN1(n17198), .IN2(n17199), .QN(n17196) );
  NAND2X0 U17832 ( .IN1(n17200), .IN2(n17201), .QN(n17199) );
  NAND2X0 U17833 ( .IN1(n17202), .IN2(n11277), .QN(n17201) );
  NOR2X0 U17834 ( .IN1(n5700), .IN2(n10350), .QN(n17202) );
  NAND2X0 U17835 ( .IN1(n17203), .IN2(n11282), .QN(n17200) );
  NOR2X0 U17836 ( .IN1(n10381), .IN2(n10349), .QN(n17203) );
  NOR2X0 U17837 ( .IN1(n11278), .IN2(n17204), .QN(n17198) );
  NAND2X0 U17838 ( .IN1(g6653), .IN2(g17688), .QN(n17204) );
  NOR2X0 U17839 ( .IN1(n17205), .IN2(n17206), .QN(n17194) );
  INVX0 U17840 ( .INP(n17197), .ZN(n17206) );
  XOR2X1 U17841 ( .IN1(test_so80), .IN2(n5531), .Q(n17197) );
  NOR2X0 U17842 ( .IN1(n17207), .IN2(n17208), .QN(n17205) );
  NAND2X0 U17843 ( .IN1(n17209), .IN2(n17210), .QN(n17208) );
  NAND2X0 U17844 ( .IN1(n17211), .IN2(n11277), .QN(n17210) );
  NOR2X0 U17845 ( .IN1(n10368), .IN2(n10367), .QN(n17211) );
  NAND2X0 U17846 ( .IN1(n17212), .IN2(n17213), .QN(n17209) );
  NOR2X0 U17847 ( .IN1(n5700), .IN2(n10331), .QN(n17212) );
  NOR2X0 U17848 ( .IN1(n11283), .IN2(n17214), .QN(n17207) );
  NAND2X0 U17849 ( .IN1(g17778), .IN2(g6629), .QN(n17214) );
  NOR2X0 U17850 ( .IN1(n17215), .IN2(n17216), .QN(n17192) );
  NOR2X0 U17851 ( .IN1(n5531), .IN2(n17217), .QN(n17216) );
  NOR2X0 U17852 ( .IN1(n17218), .IN2(n17219), .QN(n17217) );
  NAND2X0 U17853 ( .IN1(n17220), .IN2(n17221), .QN(n17219) );
  NAND2X0 U17854 ( .IN1(n11282), .IN2(n17222), .QN(n17221) );
  NAND2X0 U17855 ( .IN1(n17223), .IN2(n17224), .QN(n17222) );
  NAND2X0 U17856 ( .IN1(g6609), .IN2(g17871), .QN(n17224) );
  NAND2X0 U17857 ( .IN1(test_so80), .IN2(test_so71), .QN(n17223) );
  NAND2X0 U17858 ( .IN1(n17225), .IN2(n17226), .QN(n17220) );
  NAND2X0 U17859 ( .IN1(n17227), .IN2(n17228), .QN(n17226) );
  NAND2X0 U17860 ( .IN1(g6657), .IN2(g17722), .QN(n17228) );
  NAND2X0 U17861 ( .IN1(g6641), .IN2(g17764), .QN(n17227) );
  NAND2X0 U17862 ( .IN1(n17229), .IN2(n17230), .QN(n17218) );
  NAND2X0 U17863 ( .IN1(n17231), .IN2(n17213), .QN(n17230) );
  NOR2X0 U17864 ( .IN1(n5584), .IN2(n10436), .QN(n17231) );
  NAND2X0 U17865 ( .IN1(n11277), .IN2(n17232), .QN(n17229) );
  NAND2X0 U17866 ( .IN1(n17233), .IN2(n17234), .QN(n17232) );
  NAND2X0 U17867 ( .IN1(g6589), .IN2(g6723), .QN(n17234) );
  NAND2X0 U17868 ( .IN1(g6581), .IN2(g13099), .QN(n17233) );
  NOR2X0 U17869 ( .IN1(n17235), .IN2(g6727), .QN(n17215) );
  NOR2X0 U17870 ( .IN1(n17236), .IN2(n17237), .QN(n17235) );
  NAND2X0 U17871 ( .IN1(n17238), .IN2(n17239), .QN(n17237) );
  NAND2X0 U17872 ( .IN1(n17213), .IN2(n17240), .QN(n17239) );
  NAND2X0 U17873 ( .IN1(n17241), .IN2(n17242), .QN(n17240) );
  NAND2X0 U17874 ( .IN1(g6723), .IN2(g6605), .QN(n17242) );
  NAND2X0 U17875 ( .IN1(g13099), .IN2(g6593), .QN(n17241) );
  INVX0 U17876 ( .INP(n11278), .ZN(n17213) );
  NAND2X0 U17877 ( .IN1(n5398), .IN2(g6682), .QN(n11278) );
  NAND2X0 U17878 ( .IN1(n17225), .IN2(n17243), .QN(n17238) );
  NAND2X0 U17879 ( .IN1(n17244), .IN2(n17245), .QN(n17243) );
  NAND2X0 U17880 ( .IN1(g17871), .IN2(g6617), .QN(n17245) );
  NAND2X0 U17881 ( .IN1(test_so80), .IN2(g6601), .QN(n17244) );
  INVX0 U17882 ( .INP(n11283), .ZN(n17225) );
  NAND2X0 U17883 ( .IN1(g6741), .IN2(g6682), .QN(n11283) );
  NAND2X0 U17884 ( .IN1(n17246), .IN2(n17247), .QN(n17236) );
  NAND2X0 U17885 ( .IN1(n17248), .IN2(n11277), .QN(n17247) );
  NOR2X0 U17886 ( .IN1(g6682), .IN2(g6741), .QN(n11277) );
  NOR2X0 U17887 ( .IN1(n5584), .IN2(n10479), .QN(n17248) );
  NAND2X0 U17888 ( .IN1(n11282), .IN2(n17249), .QN(n17246) );
  NAND2X0 U17889 ( .IN1(n17250), .IN2(n17251), .QN(n17249) );
  NAND2X0 U17890 ( .IN1(g17764), .IN2(g6649), .QN(n17251) );
  NAND2X0 U17891 ( .IN1(g17722), .IN2(g6597), .QN(n17250) );
  NOR2X0 U17892 ( .IN1(g6682), .IN2(n5398), .QN(n11282) );
  NOR2X0 U17893 ( .IN1(n10292), .IN2(n10858), .QN(n17189) );
  NAND2X0 U17894 ( .IN1(n17252), .IN2(n17253), .QN(g28102) );
  NAND2X0 U17895 ( .IN1(n13488), .IN2(g4826), .QN(n17253) );
  NOR2X0 U17896 ( .IN1(n17254), .IN2(n17255), .QN(n17252) );
  NOR2X0 U17897 ( .IN1(n11034), .IN2(n17256), .QN(n17255) );
  NAND2X0 U17898 ( .IN1(n13485), .IN2(n16572), .QN(n17256) );
  NAND2X0 U17899 ( .IN1(n17257), .IN2(n17258), .QN(n16572) );
  NOR2X0 U17900 ( .IN1(n17259), .IN2(n17260), .QN(n17258) );
  NOR2X0 U17901 ( .IN1(n17261), .IN2(n17262), .QN(n17260) );
  NOR2X0 U17902 ( .IN1(n17263), .IN2(n17264), .QN(n17261) );
  NAND2X0 U17903 ( .IN1(n17265), .IN2(n17266), .QN(n17264) );
  NAND2X0 U17904 ( .IN1(n17267), .IN2(n17268), .QN(n17266) );
  NOR2X0 U17905 ( .IN1(n10370), .IN2(n10354), .QN(n17267) );
  NAND2X0 U17906 ( .IN1(n17269), .IN2(n13484), .QN(n17265) );
  NOR2X0 U17907 ( .IN1(n10385), .IN2(n10355), .QN(n17269) );
  NOR2X0 U17908 ( .IN1(n17270), .IN2(n17271), .QN(n17263) );
  NAND2X0 U17909 ( .IN1(g6275), .IN2(g14779), .QN(n17271) );
  NOR2X0 U17910 ( .IN1(n17272), .IN2(n17273), .QN(n17259) );
  INVX0 U17911 ( .INP(n17262), .ZN(n17273) );
  XNOR2X1 U17912 ( .IN1(g12422), .IN2(test_so69), .Q(n17262) );
  NOR2X0 U17913 ( .IN1(n17274), .IN2(n17275), .QN(n17272) );
  NAND2X0 U17914 ( .IN1(n17276), .IN2(n17277), .QN(n17275) );
  NAND2X0 U17915 ( .IN1(n17278), .IN2(n17268), .QN(n17277) );
  NOR2X0 U17916 ( .IN1(n5703), .IN2(n10333), .QN(n17278) );
  NAND2X0 U17917 ( .IN1(n17279), .IN2(n16575), .QN(n17276) );
  NOR2X0 U17918 ( .IN1(n10386), .IN2(n10385), .QN(n17279) );
  NOR2X0 U17919 ( .IN1(n17270), .IN2(n17280), .QN(n17274) );
  NAND2X0 U17920 ( .IN1(g17649), .IN2(g6299), .QN(n17280) );
  NOR2X0 U17921 ( .IN1(n17281), .IN2(n17282), .QN(n17257) );
  NOR2X0 U17922 ( .IN1(test_so69), .IN2(n17283), .QN(n17282) );
  NOR2X0 U17923 ( .IN1(n17284), .IN2(n17285), .QN(n17283) );
  NAND2X0 U17924 ( .IN1(n17286), .IN2(n17287), .QN(n17285) );
  NAND2X0 U17925 ( .IN1(n16575), .IN2(n17288), .QN(n17287) );
  NAND2X0 U17926 ( .IN1(n17289), .IN2(n17290), .QN(n17288) );
  NAND2X0 U17927 ( .IN1(g17845), .IN2(g6271), .QN(n17290) );
  NAND2X0 U17928 ( .IN1(g6255), .IN2(g12422), .QN(n17289) );
  NAND2X0 U17929 ( .IN1(n13484), .IN2(n17291), .QN(n17286) );
  NAND2X0 U17930 ( .IN1(n17292), .IN2(n17293), .QN(n17291) );
  NAND2X0 U17931 ( .IN1(g17743), .IN2(g6303), .QN(n17293) );
  NAND2X0 U17932 ( .IN1(g17685), .IN2(g6251), .QN(n17292) );
  NAND2X0 U17933 ( .IN1(n17294), .IN2(n17295), .QN(n17284) );
  NAND2X0 U17934 ( .IN1(n17296), .IN2(n17297), .QN(n17295) );
  NOR2X0 U17935 ( .IN1(n5586), .IN2(n10489), .QN(n17296) );
  NAND2X0 U17936 ( .IN1(n17268), .IN2(n17298), .QN(n17294) );
  NAND2X0 U17937 ( .IN1(n17299), .IN2(n17300), .QN(n17298) );
  NAND2X0 U17938 ( .IN1(g6377), .IN2(g6259), .QN(n17300) );
  NAND2X0 U17939 ( .IN1(g13085), .IN2(g6247), .QN(n17299) );
  NOR2X0 U17940 ( .IN1(n17301), .IN2(n10642), .QN(n17281) );
  NOR2X0 U17941 ( .IN1(n17302), .IN2(n17303), .QN(n17301) );
  NAND2X0 U17942 ( .IN1(n17304), .IN2(n17305), .QN(n17303) );
  NAND2X0 U17943 ( .IN1(n13484), .IN2(n17306), .QN(n17305) );
  NAND2X0 U17944 ( .IN1(n17307), .IN2(n17308), .QN(n17306) );
  NAND2X0 U17945 ( .IN1(g6263), .IN2(g17845), .QN(n17308) );
  NAND2X0 U17946 ( .IN1(g6239), .IN2(g12422), .QN(n17307) );
  NAND2X0 U17947 ( .IN1(n17297), .IN2(n17309), .QN(n17304) );
  NAND2X0 U17948 ( .IN1(n17310), .IN2(n17311), .QN(n17309) );
  NAND2X0 U17949 ( .IN1(g6243), .IN2(g6377), .QN(n17311) );
  NAND2X0 U17950 ( .IN1(g6235), .IN2(g13085), .QN(n17310) );
  NAND2X0 U17951 ( .IN1(n17312), .IN2(n17313), .QN(n17302) );
  NAND2X0 U17952 ( .IN1(n17314), .IN2(n17268), .QN(n17313) );
  NOR2X0 U17953 ( .IN1(n5586), .IN2(n10438), .QN(n17314) );
  NAND2X0 U17954 ( .IN1(n16575), .IN2(n17315), .QN(n17312) );
  NAND2X0 U17955 ( .IN1(n17316), .IN2(n17317), .QN(n17315) );
  NAND2X0 U17956 ( .IN1(g6311), .IN2(g17685), .QN(n17317) );
  NAND2X0 U17957 ( .IN1(g6295), .IN2(g17743), .QN(n17316) );
  NOR2X0 U17958 ( .IN1(n10299), .IN2(n10858), .QN(n17254) );
  NAND2X0 U17959 ( .IN1(n17318), .IN2(n17319), .QN(g28099) );
  NAND2X0 U17960 ( .IN1(test_so13), .IN2(n11014), .QN(n17319) );
  NOR2X0 U17961 ( .IN1(n17320), .IN2(n17321), .QN(n17318) );
  NOR2X0 U17962 ( .IN1(n10173), .IN2(n13511), .QN(n17321) );
  NOR2X0 U17963 ( .IN1(n17322), .IN2(n13515), .QN(n17320) );
  NAND2X0 U17964 ( .IN1(n13506), .IN2(n10968), .QN(n13515) );
  INVX0 U17965 ( .INP(n16608), .ZN(n17322) );
  NAND2X0 U17966 ( .IN1(n17323), .IN2(n17324), .QN(n16608) );
  NOR2X0 U17967 ( .IN1(n17325), .IN2(n17326), .QN(n17324) );
  NOR2X0 U17968 ( .IN1(n17327), .IN2(n17328), .QN(n17326) );
  NOR2X0 U17969 ( .IN1(n17329), .IN2(n17330), .QN(n17327) );
  NAND2X0 U17970 ( .IN1(n17331), .IN2(n17332), .QN(n17330) );
  NAND2X0 U17971 ( .IN1(n17333), .IN2(n17334), .QN(n17332) );
  NOR2X0 U17972 ( .IN1(n5698), .IN2(n10328), .QN(n17333) );
  NAND2X0 U17973 ( .IN1(n17335), .IN2(n17336), .QN(n17331) );
  NOR2X0 U17974 ( .IN1(n10377), .IN2(n10376), .QN(n17335) );
  NOR2X0 U17975 ( .IN1(n17337), .IN2(n17338), .QN(n17329) );
  NAND2X0 U17976 ( .IN1(g17607), .IN2(g5953), .QN(n17338) );
  NOR2X0 U17977 ( .IN1(n17339), .IN2(n17340), .QN(n17325) );
  INVX0 U17978 ( .INP(n17328), .ZN(n17340) );
  XNOR2X1 U17979 ( .IN1(g12350), .IN2(n5528), .Q(n17328) );
  NOR2X0 U17980 ( .IN1(n17341), .IN2(n17342), .QN(n17339) );
  NAND2X0 U17981 ( .IN1(n17343), .IN2(n17344), .QN(n17342) );
  NAND2X0 U17982 ( .IN1(n17345), .IN2(n17334), .QN(n17344) );
  NOR2X0 U17983 ( .IN1(n10361), .IN2(n10339), .QN(n17345) );
  NAND2X0 U17984 ( .IN1(n17346), .IN2(n13505), .QN(n17343) );
  NOR2X0 U17985 ( .IN1(n10376), .IN2(n10340), .QN(n17346) );
  NOR2X0 U17986 ( .IN1(n17337), .IN2(n17347), .QN(n17341) );
  NAND2X0 U17987 ( .IN1(g5929), .IN2(g14738), .QN(n17347) );
  NOR2X0 U17988 ( .IN1(n17348), .IN2(n17349), .QN(n17323) );
  NOR2X0 U17989 ( .IN1(n5528), .IN2(n17350), .QN(n17349) );
  NOR2X0 U17990 ( .IN1(n17351), .IN2(n17352), .QN(n17350) );
  NAND2X0 U17991 ( .IN1(n17353), .IN2(n17354), .QN(n17352) );
  NAND2X0 U17992 ( .IN1(n13505), .IN2(n17355), .QN(n17354) );
  NAND2X0 U17993 ( .IN1(n17356), .IN2(n17357), .QN(n17355) );
  NAND2X0 U17994 ( .IN1(g5893), .IN2(g12350), .QN(n17357) );
  NAND2X0 U17995 ( .IN1(test_so28), .IN2(g17819), .QN(n17356) );
  NAND2X0 U17996 ( .IN1(n17358), .IN2(n17359), .QN(n17353) );
  NAND2X0 U17997 ( .IN1(n17360), .IN2(n17361), .QN(n17359) );
  NAND2X0 U17998 ( .IN1(g5897), .IN2(g6031), .QN(n17361) );
  NAND2X0 U17999 ( .IN1(g5889), .IN2(g13068), .QN(n17360) );
  NAND2X0 U18000 ( .IN1(n17362), .IN2(n17363), .QN(n17351) );
  NAND2X0 U18001 ( .IN1(n17364), .IN2(n17334), .QN(n17363) );
  NOR2X0 U18002 ( .IN1(n5581), .IN2(n10433), .QN(n17364) );
  NAND2X0 U18003 ( .IN1(n17336), .IN2(n17365), .QN(n17362) );
  NAND2X0 U18004 ( .IN1(n17366), .IN2(n17367), .QN(n17365) );
  NAND2X0 U18005 ( .IN1(g5949), .IN2(g17715), .QN(n17367) );
  NAND2X0 U18006 ( .IN1(test_so13), .IN2(g17646), .QN(n17366) );
  NOR2X0 U18007 ( .IN1(n17368), .IN2(g6035), .QN(n17348) );
  NOR2X0 U18008 ( .IN1(n17369), .IN2(n17370), .QN(n17368) );
  NAND2X0 U18009 ( .IN1(n17371), .IN2(n17372), .QN(n17370) );
  NAND2X0 U18010 ( .IN1(n17336), .IN2(n17373), .QN(n17372) );
  NAND2X0 U18011 ( .IN1(n17374), .IN2(n17375), .QN(n17373) );
  NAND2X0 U18012 ( .IN1(g17819), .IN2(g5925), .QN(n17375) );
  NAND2X0 U18013 ( .IN1(g5909), .IN2(g12350), .QN(n17374) );
  NAND2X0 U18014 ( .IN1(n13505), .IN2(n17376), .QN(n17371) );
  NAND2X0 U18015 ( .IN1(n17377), .IN2(n17378), .QN(n17376) );
  NAND2X0 U18016 ( .IN1(g17715), .IN2(g5957), .QN(n17378) );
  NAND2X0 U18017 ( .IN1(g17646), .IN2(g5905), .QN(n17377) );
  NAND2X0 U18018 ( .IN1(n17379), .IN2(n17380), .QN(n17369) );
  NAND2X0 U18019 ( .IN1(n17381), .IN2(n17358), .QN(n17380) );
  NOR2X0 U18020 ( .IN1(n5581), .IN2(n10465), .QN(n17381) );
  NAND2X0 U18021 ( .IN1(n17334), .IN2(n17382), .QN(n17379) );
  NAND2X0 U18022 ( .IN1(n17383), .IN2(n17384), .QN(n17382) );
  NAND2X0 U18023 ( .IN1(g6031), .IN2(g5913), .QN(n17384) );
  NAND2X0 U18024 ( .IN1(g13068), .IN2(g5901), .QN(n17383) );
  NAND2X0 U18025 ( .IN1(n17385), .IN2(n17386), .QN(g28096) );
  NAND2X0 U18026 ( .IN1(n13530), .IN2(g4821), .QN(n17386) );
  NOR2X0 U18027 ( .IN1(n17387), .IN2(n17388), .QN(n17385) );
  NOR2X0 U18028 ( .IN1(n11034), .IN2(n17389), .QN(n17388) );
  NAND2X0 U18029 ( .IN1(n13527), .IN2(n16646), .QN(n17389) );
  NAND2X0 U18030 ( .IN1(n17390), .IN2(n17391), .QN(n16646) );
  NOR2X0 U18031 ( .IN1(n17392), .IN2(n17393), .QN(n17391) );
  NOR2X0 U18032 ( .IN1(n17394), .IN2(n17395), .QN(n17393) );
  NOR2X0 U18033 ( .IN1(n17396), .IN2(n17397), .QN(n17394) );
  NAND2X0 U18034 ( .IN1(n17398), .IN2(n17399), .QN(n17397) );
  NAND2X0 U18035 ( .IN1(n17400), .IN2(n17401), .QN(n17399) );
  NOR2X0 U18036 ( .IN1(n5705), .IN2(n10329), .QN(n17400) );
  NAND2X0 U18037 ( .IN1(n17402), .IN2(test_so5), .QN(n17398) );
  NOR2X0 U18038 ( .IN1(n10378), .IN2(n12443), .QN(n17402) );
  NOR2X0 U18039 ( .IN1(n17403), .IN2(n17404), .QN(n17396) );
  NAND2X0 U18040 ( .IN1(g17580), .IN2(g5607), .QN(n17404) );
  NOR2X0 U18041 ( .IN1(n17405), .IN2(n17406), .QN(n17392) );
  INVX0 U18042 ( .INP(n17395), .ZN(n17406) );
  XNOR2X1 U18043 ( .IN1(g12300), .IN2(n5529), .Q(n17395) );
  NOR2X0 U18044 ( .IN1(n17407), .IN2(n17408), .QN(n17405) );
  NAND2X0 U18045 ( .IN1(n17409), .IN2(n17410), .QN(n17408) );
  NAND2X0 U18046 ( .IN1(n17411), .IN2(n17401), .QN(n17410) );
  NOR2X0 U18047 ( .IN1(n10363), .IN2(n10342), .QN(n17411) );
  NAND2X0 U18048 ( .IN1(n17412), .IN2(n13526), .QN(n17409) );
  NOR2X0 U18049 ( .IN1(n10378), .IN2(n10343), .QN(n17412) );
  NOR2X0 U18050 ( .IN1(n17403), .IN2(n17413), .QN(n17407) );
  NAND2X0 U18051 ( .IN1(g5583), .IN2(g14694), .QN(n17413) );
  NOR2X0 U18052 ( .IN1(n17414), .IN2(n17415), .QN(n17390) );
  NOR2X0 U18053 ( .IN1(n5529), .IN2(n17416), .QN(n17415) );
  NOR2X0 U18054 ( .IN1(n17417), .IN2(n17418), .QN(n17416) );
  NAND2X0 U18055 ( .IN1(n17419), .IN2(n17420), .QN(n17418) );
  NAND2X0 U18056 ( .IN1(n13526), .IN2(n17421), .QN(n17420) );
  NAND2X0 U18057 ( .IN1(n17422), .IN2(n17423), .QN(n17421) );
  NAND2X0 U18058 ( .IN1(g5571), .IN2(g17813), .QN(n17423) );
  NAND2X0 U18059 ( .IN1(g5547), .IN2(g12300), .QN(n17422) );
  NAND2X0 U18060 ( .IN1(n17424), .IN2(n17425), .QN(n17419) );
  NAND2X0 U18061 ( .IN1(n17426), .IN2(n17427), .QN(n17425) );
  NAND2X0 U18062 ( .IN1(g5551), .IN2(g5685), .QN(n17427) );
  NAND2X0 U18063 ( .IN1(g5543), .IN2(g13049), .QN(n17426) );
  NAND2X0 U18064 ( .IN1(n17428), .IN2(n17429), .QN(n17417) );
  NAND2X0 U18065 ( .IN1(n17430), .IN2(n17401), .QN(n17429) );
  NOR2X0 U18066 ( .IN1(n5582), .IN2(n10434), .QN(n17430) );
  NAND2X0 U18067 ( .IN1(n16648), .IN2(n17431), .QN(n17428) );
  NAND2X0 U18068 ( .IN1(n17432), .IN2(n17433), .QN(n17431) );
  NAND2X0 U18069 ( .IN1(g5619), .IN2(g17604), .QN(n17433) );
  NAND2X0 U18070 ( .IN1(g5603), .IN2(g17678), .QN(n17432) );
  NOR2X0 U18071 ( .IN1(n17434), .IN2(g5689), .QN(n17414) );
  NOR2X0 U18072 ( .IN1(n17435), .IN2(n17436), .QN(n17434) );
  NAND2X0 U18073 ( .IN1(n17437), .IN2(n17438), .QN(n17436) );
  NAND2X0 U18074 ( .IN1(n16648), .IN2(n17439), .QN(n17438) );
  NAND2X0 U18075 ( .IN1(n17440), .IN2(n17441), .QN(n17439) );
  NAND2X0 U18076 ( .IN1(g17813), .IN2(g5579), .QN(n17441) );
  NAND2X0 U18077 ( .IN1(g5563), .IN2(g12300), .QN(n17440) );
  NAND2X0 U18078 ( .IN1(n13526), .IN2(n17442), .QN(n17437) );
  NAND2X0 U18079 ( .IN1(n17443), .IN2(n17444), .QN(n17442) );
  NAND2X0 U18080 ( .IN1(g17678), .IN2(g5611), .QN(n17444) );
  NAND2X0 U18081 ( .IN1(test_so6), .IN2(g17604), .QN(n17443) );
  NAND2X0 U18082 ( .IN1(n17445), .IN2(n17446), .QN(n17435) );
  NAND2X0 U18083 ( .IN1(n17447), .IN2(n17424), .QN(n17446) );
  NOR2X0 U18084 ( .IN1(n5582), .IN2(n10470), .QN(n17447) );
  NAND2X0 U18085 ( .IN1(n17401), .IN2(n17448), .QN(n17445) );
  NAND2X0 U18086 ( .IN1(n17449), .IN2(n17450), .QN(n17448) );
  NAND2X0 U18087 ( .IN1(g5685), .IN2(g5567), .QN(n17450) );
  NAND2X0 U18088 ( .IN1(g13049), .IN2(g5555), .QN(n17449) );
  NOR2X0 U18089 ( .IN1(n10288), .IN2(n10858), .QN(n17387) );
  NAND2X0 U18090 ( .IN1(n17451), .IN2(n17452), .QN(g28093) );
  NAND2X0 U18091 ( .IN1(n13548), .IN2(g29220), .QN(n17452) );
  NOR2X0 U18092 ( .IN1(n17453), .IN2(n17454), .QN(n17451) );
  NOR2X0 U18093 ( .IN1(n11034), .IN2(n17455), .QN(n17454) );
  NAND2X0 U18094 ( .IN1(g33959), .IN2(n16686), .QN(n17455) );
  NAND2X0 U18095 ( .IN1(n17456), .IN2(n17457), .QN(n16686) );
  NOR2X0 U18096 ( .IN1(n17458), .IN2(n17459), .QN(n17457) );
  NOR2X0 U18097 ( .IN1(n17460), .IN2(n17461), .QN(n17459) );
  NOR2X0 U18098 ( .IN1(n17462), .IN2(n17463), .QN(n17460) );
  NAND2X0 U18099 ( .IN1(n17464), .IN2(n17465), .QN(n17463) );
  NAND2X0 U18100 ( .IN1(n17466), .IN2(n17467), .QN(n17465) );
  NOR2X0 U18101 ( .IN1(n10359), .IN2(n10336), .QN(n17466) );
  NAND2X0 U18102 ( .IN1(n17468), .IN2(n13545), .QN(n17464) );
  NOR2X0 U18103 ( .IN1(n10374), .IN2(n10337), .QN(n17468) );
  NOR2X0 U18104 ( .IN1(n11266), .IN2(n17469), .QN(n17462) );
  NAND2X0 U18105 ( .IN1(g5236), .IN2(g14662), .QN(n17469) );
  NOR2X0 U18106 ( .IN1(n17470), .IN2(n17471), .QN(n17458) );
  INVX0 U18107 ( .INP(n17461), .ZN(n17471) );
  XNOR2X1 U18108 ( .IN1(g12238), .IN2(test_so10), .Q(n17461) );
  NOR2X0 U18109 ( .IN1(n17472), .IN2(n17473), .QN(n17470) );
  NAND2X0 U18110 ( .IN1(n17474), .IN2(n17475), .QN(n17473) );
  NAND2X0 U18111 ( .IN1(n17476), .IN2(test_so82), .QN(n17475) );
  NOR2X0 U18112 ( .IN1(n5704), .IN2(n11267), .QN(n17476) );
  NAND2X0 U18113 ( .IN1(n17477), .IN2(n17478), .QN(n17474) );
  NOR2X0 U18114 ( .IN1(n10360), .IN2(n10359), .QN(n17477) );
  NOR2X0 U18115 ( .IN1(n11271), .IN2(n17479), .QN(n17472) );
  INVX0 U18116 ( .INP(n17480), .ZN(n17479) );
  NOR2X0 U18117 ( .IN1(n10374), .IN2(n10375), .QN(n17480) );
  NOR2X0 U18118 ( .IN1(n17481), .IN2(n17482), .QN(n17456) );
  NOR2X0 U18119 ( .IN1(test_so10), .IN2(n17483), .QN(n17482) );
  NOR2X0 U18120 ( .IN1(n17484), .IN2(n17485), .QN(n17483) );
  NAND2X0 U18121 ( .IN1(n17486), .IN2(n17487), .QN(n17485) );
  NAND2X0 U18122 ( .IN1(n13545), .IN2(n17488), .QN(n17487) );
  NAND2X0 U18123 ( .IN1(n17489), .IN2(n17490), .QN(n17488) );
  NAND2X0 U18124 ( .IN1(g17639), .IN2(g5264), .QN(n17490) );
  NAND2X0 U18125 ( .IN1(g17577), .IN2(g5212), .QN(n17489) );
  NAND2X0 U18126 ( .IN1(g31860), .IN2(n17491), .QN(n17486) );
  NAND2X0 U18127 ( .IN1(n17492), .IN2(n17493), .QN(n17491) );
  NAND2X0 U18128 ( .IN1(g17787), .IN2(g5232), .QN(n17493) );
  NAND2X0 U18129 ( .IN1(g5216), .IN2(g12238), .QN(n17492) );
  NAND2X0 U18130 ( .IN1(n17494), .IN2(n17495), .QN(n17484) );
  NAND2X0 U18131 ( .IN1(n17496), .IN2(n17478), .QN(n17495) );
  NOR2X0 U18132 ( .IN1(n5579), .IN2(n10460), .QN(n17496) );
  NAND2X0 U18133 ( .IN1(n17467), .IN2(n17497), .QN(n17494) );
  NAND2X0 U18134 ( .IN1(n17498), .IN2(n17499), .QN(n17497) );
  NAND2X0 U18135 ( .IN1(g5220), .IN2(g5339), .QN(n17499) );
  NAND2X0 U18136 ( .IN1(g5208), .IN2(g13039), .QN(n17498) );
  NOR2X0 U18137 ( .IN1(n17500), .IN2(n10641), .QN(n17481) );
  NOR2X0 U18138 ( .IN1(n17501), .IN2(n17502), .QN(n17500) );
  NAND2X0 U18139 ( .IN1(n17503), .IN2(n17504), .QN(n17502) );
  NAND2X0 U18140 ( .IN1(n17478), .IN2(n17505), .QN(n17504) );
  NAND2X0 U18141 ( .IN1(n17506), .IN2(n17507), .QN(n17505) );
  NAND2X0 U18142 ( .IN1(g5339), .IN2(g5204), .QN(n17507) );
  NAND2X0 U18143 ( .IN1(g13039), .IN2(g5196), .QN(n17506) );
  INVX0 U18144 ( .INP(n11266), .ZN(n17478) );
  NAND2X0 U18145 ( .IN1(n5588), .IN2(n5393), .QN(n11266) );
  NAND2X0 U18146 ( .IN1(g31860), .IN2(n17508), .QN(n17503) );
  NAND2X0 U18147 ( .IN1(n17509), .IN2(n17510), .QN(n17508) );
  NAND2X0 U18148 ( .IN1(g5272), .IN2(g17577), .QN(n17510) );
  NAND2X0 U18149 ( .IN1(g5256), .IN2(g17639), .QN(n17509) );
  INVX0 U18150 ( .INP(n11271), .ZN(g31860) );
  NAND2X0 U18151 ( .IN1(g5357), .IN2(g5297), .QN(n11271) );
  NAND2X0 U18152 ( .IN1(n17511), .IN2(n17512), .QN(n17501) );
  NAND2X0 U18153 ( .IN1(n17513), .IN2(n17467), .QN(n17512) );
  INVX0 U18154 ( .INP(n11267), .ZN(n17467) );
  NAND2X0 U18155 ( .IN1(n5393), .IN2(g5297), .QN(n11267) );
  NOR2X0 U18156 ( .IN1(n5579), .IN2(n10432), .QN(n17513) );
  NAND2X0 U18157 ( .IN1(n13545), .IN2(n17514), .QN(n17511) );
  NAND2X0 U18158 ( .IN1(n17515), .IN2(n17516), .QN(n17514) );
  NAND2X0 U18159 ( .IN1(g5224), .IN2(g17787), .QN(n17516) );
  NAND2X0 U18160 ( .IN1(g5200), .IN2(g12238), .QN(n17515) );
  INVX0 U18161 ( .INP(n11270), .ZN(n13545) );
  NAND2X0 U18162 ( .IN1(n5588), .IN2(g5357), .QN(n11270) );
  NOR2X0 U18163 ( .IN1(n10303), .IN2(n10859), .QN(n17453) );
  NAND2X0 U18164 ( .IN1(n17517), .IN2(n17518), .QN(g28092) );
  NAND2X0 U18165 ( .IN1(n11060), .IN2(g5057), .QN(n17518) );
  NAND2X0 U18166 ( .IN1(n14887), .IN2(n10968), .QN(n17517) );
  NAND2X0 U18167 ( .IN1(n17519), .IN2(n17520), .QN(n14887) );
  NOR2X0 U18168 ( .IN1(n5615), .IN2(n10278), .QN(n17520) );
  NOR2X0 U18169 ( .IN1(g5046), .IN2(n17521), .QN(n17519) );
  NAND2X0 U18170 ( .IN1(n17522), .IN2(n17523), .QN(g28091) );
  NAND2X0 U18171 ( .IN1(n11060), .IN2(g5069), .QN(n17523) );
  NAND2X0 U18172 ( .IN1(n14888), .IN2(n10969), .QN(n17522) );
  NAND2X0 U18173 ( .IN1(n17524), .IN2(n17525), .QN(n14888) );
  NOR2X0 U18174 ( .IN1(n5578), .IN2(n10253), .QN(n17525) );
  NOR2X0 U18175 ( .IN1(n17526), .IN2(g5057), .QN(n17524) );
  INVX0 U18176 ( .INP(n17521), .ZN(n17526) );
  NAND2X0 U18177 ( .IN1(n17527), .IN2(n17528), .QN(n17521) );
  NAND2X0 U18178 ( .IN1(g84), .IN2(g5041), .QN(n17528) );
  NAND2X0 U18179 ( .IN1(n17529), .IN2(g5052), .QN(n17527) );
  INVX0 U18180 ( .INP(g84), .ZN(n17529) );
  NAND2X0 U18181 ( .IN1(n17530), .IN2(n17531), .QN(g28090) );
  NAND2X0 U18182 ( .IN1(n17532), .IN2(n12500), .QN(n17531) );
  INVX0 U18183 ( .INP(n12506), .ZN(n12500) );
  NAND2X0 U18184 ( .IN1(n11377), .IN2(n11389), .QN(n12506) );
  NOR2X0 U18185 ( .IN1(n11035), .IN2(n17533), .QN(n17532) );
  NOR2X0 U18186 ( .IN1(n17534), .IN2(g4961), .QN(n17533) );
  NOR2X0 U18187 ( .IN1(n17535), .IN2(n13581), .QN(n17534) );
  NOR2X0 U18188 ( .IN1(n17536), .IN2(n17537), .QN(n17535) );
  NAND2X0 U18189 ( .IN1(n17538), .IN2(n17539), .QN(n17537) );
  NAND2X0 U18190 ( .IN1(n17540), .IN2(g4049), .QN(n17539) );
  NAND2X0 U18191 ( .IN1(n10396), .IN2(n13582), .QN(n17538) );
  NAND2X0 U18192 ( .IN1(n17541), .IN2(n17542), .QN(n17536) );
  NAND2X0 U18193 ( .IN1(n17543), .IN2(g4045), .QN(n17542) );
  NAND2X0 U18194 ( .IN1(n10397), .IN2(n17544), .QN(n17541) );
  NAND2X0 U18195 ( .IN1(n13586), .IN2(g4961), .QN(n17530) );
  NAND2X0 U18196 ( .IN1(n17545), .IN2(n17546), .QN(g28089) );
  NAND2X0 U18197 ( .IN1(n17547), .IN2(n12510), .QN(n17546) );
  INVX0 U18198 ( .INP(n12514), .ZN(n12510) );
  NAND2X0 U18199 ( .IN1(n11377), .IN2(n11388), .QN(n12514) );
  NOR2X0 U18200 ( .IN1(n11035), .IN2(n17548), .QN(n17547) );
  NOR2X0 U18201 ( .IN1(n17549), .IN2(g4950), .QN(n17548) );
  NOR2X0 U18202 ( .IN1(n17550), .IN2(n13603), .QN(n17549) );
  NOR2X0 U18203 ( .IN1(n17551), .IN2(n17552), .QN(n17550) );
  NAND2X0 U18204 ( .IN1(n17553), .IN2(n17554), .QN(n17552) );
  NAND2X0 U18205 ( .IN1(n17555), .IN2(g3698), .QN(n17554) );
  NAND2X0 U18206 ( .IN1(n10392), .IN2(n13604), .QN(n17553) );
  NAND2X0 U18207 ( .IN1(n17556), .IN2(n17557), .QN(n17551) );
  NAND2X0 U18208 ( .IN1(n17558), .IN2(g3694), .QN(n17557) );
  NAND2X0 U18209 ( .IN1(n10393), .IN2(n17559), .QN(n17556) );
  NAND2X0 U18210 ( .IN1(n13608), .IN2(g4950), .QN(n17545) );
  NAND2X0 U18211 ( .IN1(n17560), .IN2(n17561), .QN(g28088) );
  NAND2X0 U18212 ( .IN1(n17562), .IN2(n12519), .QN(n17561) );
  NOR2X0 U18213 ( .IN1(n17563), .IN2(n11399), .QN(n12519) );
  INVX0 U18214 ( .INP(n11377), .ZN(n17563) );
  NOR2X0 U18215 ( .IN1(n11035), .IN2(n17564), .QN(n17562) );
  NOR2X0 U18216 ( .IN1(n17565), .IN2(g4939), .QN(n17564) );
  NOR2X0 U18217 ( .IN1(n17566), .IN2(n13626), .QN(n17565) );
  NOR2X0 U18218 ( .IN1(n17567), .IN2(n17568), .QN(n17566) );
  NAND2X0 U18219 ( .IN1(n17569), .IN2(n17570), .QN(n17568) );
  NAND2X0 U18220 ( .IN1(n17571), .IN2(g3347), .QN(n17570) );
  NAND2X0 U18221 ( .IN1(n10387), .IN2(n13624), .QN(n17569) );
  NAND2X0 U18222 ( .IN1(n17572), .IN2(n17573), .QN(n17567) );
  NAND2X0 U18223 ( .IN1(n13620), .IN2(g3343), .QN(n17573) );
  NAND2X0 U18224 ( .IN1(n10388), .IN2(n17574), .QN(n17572) );
  NAND2X0 U18225 ( .IN1(n13629), .IN2(g4939), .QN(n17560) );
  NAND2X0 U18226 ( .IN1(n17575), .IN2(n17576), .QN(g28087) );
  NAND2X0 U18227 ( .IN1(n17577), .IN2(n12527), .QN(n17576) );
  INVX0 U18228 ( .INP(n12063), .ZN(n12527) );
  NAND2X0 U18229 ( .IN1(n11377), .IN2(n17578), .QN(n12063) );
  NOR2X0 U18230 ( .IN1(n17579), .IN2(n5367), .QN(n11377) );
  NOR2X0 U18231 ( .IN1(n11035), .IN2(n17580), .QN(n17577) );
  NOR2X0 U18232 ( .IN1(n4689), .IN2(g4894), .QN(n17580) );
  NAND2X0 U18233 ( .IN1(n13467), .IN2(g4894), .QN(n17575) );
  NOR2X0 U18234 ( .IN1(n13464), .IN2(n11016), .QN(n13467) );
  NOR2X0 U18235 ( .IN1(n5713), .IN2(n17581), .QN(n13464) );
  NOR2X0 U18236 ( .IN1(n17582), .IN2(n11399), .QN(n17581) );
  NAND2X0 U18237 ( .IN1(n5517), .IN2(n5360), .QN(n11399) );
  INVX0 U18238 ( .INP(n17583), .ZN(n17582) );
  NOR2X0 U18239 ( .IN1(n5863), .IN2(n17584), .QN(n17583) );
  NAND2X0 U18240 ( .IN1(n17585), .IN2(n17586), .QN(g28086) );
  NAND2X0 U18241 ( .IN1(n17587), .IN2(n12541), .QN(n17586) );
  NOR2X0 U18242 ( .IN1(n11340), .IN2(n11356), .QN(n12541) );
  NOR2X0 U18243 ( .IN1(n11035), .IN2(n17588), .QN(n17587) );
  NOR2X0 U18244 ( .IN1(n17589), .IN2(g4771), .QN(n17588) );
  NOR2X0 U18245 ( .IN1(n17590), .IN2(n13483), .QN(n17589) );
  NOR2X0 U18246 ( .IN1(n17591), .IN2(n17592), .QN(n17590) );
  NAND2X0 U18247 ( .IN1(n17593), .IN2(n17594), .QN(n17592) );
  NAND2X0 U18248 ( .IN1(n16575), .IN2(g6390), .QN(n17594) );
  INVX0 U18249 ( .INP(n12455), .ZN(n16575) );
  NAND2X0 U18250 ( .IN1(g6395), .IN2(g6336), .QN(n12455) );
  NAND2X0 U18251 ( .IN1(n10389), .IN2(n13484), .QN(n17593) );
  NOR2X0 U18252 ( .IN1(g6336), .IN2(n5396), .QN(n13484) );
  NAND2X0 U18253 ( .IN1(n17595), .IN2(n17596), .QN(n17591) );
  NAND2X0 U18254 ( .IN1(n17268), .IN2(g6386), .QN(n17596) );
  INVX0 U18255 ( .INP(n13481), .ZN(n17268) );
  NAND2X0 U18256 ( .IN1(n5396), .IN2(g6336), .QN(n13481) );
  NAND2X0 U18257 ( .IN1(n10390), .IN2(n17297), .QN(n17595) );
  INVX0 U18258 ( .INP(n17270), .ZN(n17297) );
  NAND2X0 U18259 ( .IN1(n5592), .IN2(n5396), .QN(n17270) );
  NAND2X0 U18260 ( .IN1(n13488), .IN2(g4771), .QN(n17585) );
  NOR2X0 U18261 ( .IN1(n13485), .IN2(n11015), .QN(n13488) );
  INVX0 U18262 ( .INP(n13483), .ZN(n13485) );
  NAND2X0 U18263 ( .IN1(g4688), .IN2(n17597), .QN(n13483) );
  NAND2X0 U18264 ( .IN1(n13454), .IN2(n17598), .QN(n17597) );
  NOR2X0 U18265 ( .IN1(n5613), .IN2(n11365), .QN(n13454) );
  NAND2X0 U18266 ( .IN1(n17599), .IN2(n17600), .QN(g28085) );
  NAND2X0 U18267 ( .IN1(n17601), .IN2(n12551), .QN(n17600) );
  NOR2X0 U18268 ( .IN1(n11340), .IN2(n11357), .QN(n12551) );
  NOR2X0 U18269 ( .IN1(n11036), .IN2(n17602), .QN(n17601) );
  NOR2X0 U18270 ( .IN1(n17603), .IN2(g4760), .QN(n17602) );
  NOR2X0 U18271 ( .IN1(n17604), .IN2(n13504), .QN(n17603) );
  NOR2X0 U18272 ( .IN1(n17605), .IN2(n17606), .QN(n17604) );
  NAND2X0 U18273 ( .IN1(n17607), .IN2(n17608), .QN(n17606) );
  NAND2X0 U18274 ( .IN1(n13505), .IN2(n10694), .QN(n17608) );
  NOR2X0 U18275 ( .IN1(g5990), .IN2(n10639), .QN(n13505) );
  NAND2X0 U18276 ( .IN1(test_so50), .IN2(n17336), .QN(n17607) );
  INVX0 U18277 ( .INP(n12451), .ZN(n17336) );
  NAND2X0 U18278 ( .IN1(test_so57), .IN2(g5990), .QN(n12451) );
  NAND2X0 U18279 ( .IN1(n17609), .IN2(n17610), .QN(n17605) );
  NAND2X0 U18280 ( .IN1(n17334), .IN2(g6040), .QN(n17610) );
  INVX0 U18281 ( .INP(n13502), .ZN(n17334) );
  NAND2X0 U18282 ( .IN1(g5990), .IN2(n10639), .QN(n13502) );
  NAND2X0 U18283 ( .IN1(n10391), .IN2(n17358), .QN(n17609) );
  INVX0 U18284 ( .INP(n17337), .ZN(n17358) );
  NAND2X0 U18285 ( .IN1(n5589), .IN2(n10639), .QN(n17337) );
  INVX0 U18286 ( .INP(n17611), .ZN(n17599) );
  NOR2X0 U18287 ( .IN1(n13511), .IN2(n5775), .QN(n17611) );
  NAND2X0 U18288 ( .IN1(n13504), .IN2(n10969), .QN(n13511) );
  INVX0 U18289 ( .INP(n13506), .ZN(n13504) );
  NOR2X0 U18290 ( .IN1(n10527), .IN2(n17612), .QN(n13506) );
  INVX0 U18291 ( .INP(n17613), .ZN(n17612) );
  NAND2X0 U18292 ( .IN1(n13452), .IN2(n17598), .QN(n17613) );
  NOR2X0 U18293 ( .IN1(n5877), .IN2(n11356), .QN(n13452) );
  NAND2X0 U18294 ( .IN1(n5361), .IN2(g4709), .QN(n11356) );
  NAND2X0 U18295 ( .IN1(n17614), .IN2(n17615), .QN(g28084) );
  NAND2X0 U18296 ( .IN1(n17616), .IN2(n12560), .QN(n17615) );
  NOR2X0 U18297 ( .IN1(n11340), .IN2(n11352), .QN(n12560) );
  NOR2X0 U18298 ( .IN1(n11036), .IN2(n17617), .QN(n17616) );
  NOR2X0 U18299 ( .IN1(n17618), .IN2(test_so18), .QN(n17617) );
  NOR2X0 U18300 ( .IN1(n17619), .IN2(n13525), .QN(n17618) );
  NOR2X0 U18301 ( .IN1(n17620), .IN2(n17621), .QN(n17619) );
  NAND2X0 U18302 ( .IN1(n17622), .IN2(n17623), .QN(n17621) );
  NAND2X0 U18303 ( .IN1(n16648), .IN2(g5698), .QN(n17623) );
  INVX0 U18304 ( .INP(n12443), .ZN(n16648) );
  NAND2X0 U18305 ( .IN1(g5703), .IN2(g5644), .QN(n12443) );
  NAND2X0 U18306 ( .IN1(n10394), .IN2(n13526), .QN(n17622) );
  NOR2X0 U18307 ( .IN1(g5644), .IN2(n5397), .QN(n13526) );
  NAND2X0 U18308 ( .IN1(n17624), .IN2(n17625), .QN(n17620) );
  NAND2X0 U18309 ( .IN1(n17401), .IN2(g5694), .QN(n17625) );
  INVX0 U18310 ( .INP(n13523), .ZN(n17401) );
  NAND2X0 U18311 ( .IN1(n5397), .IN2(g5644), .QN(n13523) );
  NAND2X0 U18312 ( .IN1(n10395), .IN2(n17424), .QN(n17624) );
  INVX0 U18313 ( .INP(n17403), .ZN(n17424) );
  NAND2X0 U18314 ( .IN1(n5593), .IN2(n5397), .QN(n17403) );
  NAND2X0 U18315 ( .IN1(n13530), .IN2(test_so18), .QN(n17614) );
  NOR2X0 U18316 ( .IN1(n13527), .IN2(n11019), .QN(n13530) );
  INVX0 U18317 ( .INP(n13525), .ZN(n13527) );
  NAND2X0 U18318 ( .IN1(g4674), .IN2(n17626), .QN(n13525) );
  NAND2X0 U18319 ( .IN1(n13453), .IN2(n17598), .QN(n17626) );
  NOR2X0 U18320 ( .IN1(n5876), .IN2(n11357), .QN(n13453) );
  NAND2X0 U18321 ( .IN1(n5518), .IN2(g4785), .QN(n11357) );
  NAND2X0 U18322 ( .IN1(n17627), .IN2(n17628), .QN(g28083) );
  NAND2X0 U18323 ( .IN1(n17629), .IN2(n12568), .QN(n17628) );
  NOR2X0 U18324 ( .IN1(n11340), .IN2(n11365), .QN(n12568) );
  NAND2X0 U18325 ( .IN1(g4785), .IN2(g4709), .QN(n11365) );
  NAND2X0 U18326 ( .IN1(n17630), .IN2(g4793), .QN(n11340) );
  NOR2X0 U18327 ( .IN1(test_so29), .IN2(n5707), .QN(n17630) );
  NOR2X0 U18328 ( .IN1(n11036), .IN2(n17631), .QN(n17629) );
  NOR2X0 U18329 ( .IN1(n4708), .IN2(g4704), .QN(n17631) );
  NAND2X0 U18330 ( .IN1(n13548), .IN2(g4704), .QN(n17627) );
  NOR2X0 U18331 ( .IN1(g33959), .IN2(n11015), .QN(n13548) );
  INVX0 U18332 ( .INP(n10624), .ZN(g33959) );
  NAND2X0 U18333 ( .IN1(g4646), .IN2(n17632), .QN(n10624) );
  NAND2X0 U18334 ( .IN1(n13455), .IN2(n17598), .QN(n17632) );
  INVX0 U18335 ( .INP(n17633), .ZN(n17598) );
  NAND2X0 U18336 ( .IN1(n17634), .IN2(n17635), .QN(n17633) );
  NOR2X0 U18337 ( .IN1(n10543), .IN2(n17636), .QN(n17635) );
  NAND2X0 U18338 ( .IN1(g4776), .IN2(n10661), .QN(n17636) );
  NOR2X0 U18339 ( .IN1(n10645), .IN2(n17637), .QN(n17634) );
  NAND2X0 U18340 ( .IN1(n5368), .IN2(g4669), .QN(n17637) );
  NOR2X0 U18341 ( .IN1(n5862), .IN2(n11352), .QN(n13455) );
  NAND2X0 U18342 ( .IN1(n5518), .IN2(n5361), .QN(n11352) );
  NAND2X0 U18343 ( .IN1(n17638), .IN2(n17639), .QN(g28082) );
  NAND2X0 U18344 ( .IN1(n17640), .IN2(g4521), .QN(n17639) );
  NAND2X0 U18345 ( .IN1(n17641), .IN2(n10969), .QN(n17640) );
  NAND2X0 U18346 ( .IN1(n17642), .IN2(n5752), .QN(n17638) );
  NOR2X0 U18347 ( .IN1(n11036), .IN2(n17643), .QN(n17642) );
  NAND2X0 U18348 ( .IN1(n17644), .IN2(n17645), .QN(g28074) );
  NAND2X0 U18349 ( .IN1(n11062), .IN2(g4119), .QN(n17645) );
  NOR2X0 U18350 ( .IN1(n17646), .IN2(n17647), .QN(n17644) );
  INVX0 U18351 ( .INP(n17648), .ZN(n17647) );
  NAND2X0 U18352 ( .IN1(n4721), .IN2(n4714), .QN(n17648) );
  NOR2X0 U18353 ( .IN1(n4714), .IN2(n17649), .QN(n17646) );
  NAND2X0 U18354 ( .IN1(n10930), .IN2(g4122), .QN(n17649) );
  NAND2X0 U18355 ( .IN1(n17650), .IN2(n17651), .QN(g28073) );
  NAND2X0 U18356 ( .IN1(n17652), .IN2(n4721), .QN(n17651) );
  NOR2X0 U18357 ( .IN1(n17653), .IN2(n17654), .QN(n17650) );
  NOR2X0 U18358 ( .IN1(n10102), .IN2(n10860), .QN(n17654) );
  INVX0 U18359 ( .INP(n17655), .ZN(n17653) );
  NAND2X0 U18360 ( .IN1(n10930), .IN2(n17656), .QN(n17655) );
  NOR2X0 U18361 ( .IN1(n17652), .IN2(n10114), .QN(n17656) );
  NOR2X0 U18362 ( .IN1(n17657), .IN2(n5711), .QN(n17652) );
  NAND2X0 U18363 ( .IN1(n17658), .IN2(n17659), .QN(g28072) );
  NAND2X0 U18364 ( .IN1(n17660), .IN2(n4721), .QN(n17659) );
  NOR2X0 U18365 ( .IN1(n17661), .IN2(n17662), .QN(n17658) );
  NOR2X0 U18366 ( .IN1(n10522), .IN2(n10860), .QN(n17662) );
  NOR2X0 U18367 ( .IN1(n11036), .IN2(n17663), .QN(n17661) );
  INVX0 U18368 ( .INP(n17664), .ZN(n17663) );
  NOR2X0 U18369 ( .IN1(n17660), .IN2(n10102), .QN(n17664) );
  INVX0 U18370 ( .INP(n17665), .ZN(n17660) );
  NAND2X0 U18371 ( .IN1(n17666), .IN2(n422), .QN(n17665) );
  NOR2X0 U18372 ( .IN1(n5416), .IN2(g4057), .QN(n17666) );
  INVX0 U18373 ( .INP(n17667), .ZN(g28071) );
  NOR2X0 U18374 ( .IN1(n17668), .IN2(n17669), .QN(n17667) );
  NOR2X0 U18375 ( .IN1(n17670), .IN2(n10522), .QN(n17669) );
  INVX0 U18376 ( .INP(n17671), .ZN(n17670) );
  NOR2X0 U18377 ( .IN1(n17671), .IN2(n10551), .QN(n17668) );
  NOR2X0 U18378 ( .IN1(n17672), .IN2(n11017), .QN(n17671) );
  NOR2X0 U18379 ( .IN1(n17657), .IN2(g4057), .QN(n17672) );
  NAND2X0 U18380 ( .IN1(n422), .IN2(n5416), .QN(n17657) );
  NOR2X0 U18381 ( .IN1(n17673), .IN2(n17674), .QN(n422) );
  NAND2X0 U18382 ( .IN1(n10644), .IN2(n12424), .QN(n17674) );
  NAND2X0 U18383 ( .IN1(n15132), .IN2(n5350), .QN(n17673) );
  INVX0 U18384 ( .INP(n12428), .ZN(n15132) );
  NAND2X0 U18385 ( .IN1(n5480), .IN2(n5340), .QN(n12428) );
  NAND2X0 U18386 ( .IN1(n17675), .IN2(n17676), .QN(g28070) );
  NOR2X0 U18387 ( .IN1(n17677), .IN2(n17678), .QN(n17676) );
  NOR2X0 U18388 ( .IN1(n10238), .IN2(n10860), .QN(n17678) );
  NOR2X0 U18389 ( .IN1(n11037), .IN2(n17679), .QN(n17677) );
  NAND2X0 U18390 ( .IN1(test_so11), .IN2(n16693), .QN(n17679) );
  NOR2X0 U18391 ( .IN1(n10631), .IN2(n17680), .QN(n17675) );
  NOR2X0 U18392 ( .IN1(test_so11), .IN2(n16693), .QN(n17680) );
  NAND2X0 U18393 ( .IN1(n17681), .IN2(g4082), .QN(n16693) );
  NAND2X0 U18394 ( .IN1(n17682), .IN2(n17683), .QN(g28069) );
  NAND2X0 U18395 ( .IN1(n13586), .IN2(g4035), .QN(n17683) );
  NOR2X0 U18396 ( .IN1(n13583), .IN2(n11018), .QN(n13586) );
  NOR2X0 U18397 ( .IN1(n17684), .IN2(n17685), .QN(n17682) );
  NOR2X0 U18398 ( .IN1(n11037), .IN2(n17686), .QN(n17685) );
  NAND2X0 U18399 ( .IN1(n13583), .IN2(n16731), .QN(n17686) );
  NAND2X0 U18400 ( .IN1(n17687), .IN2(n17688), .QN(n16731) );
  NOR2X0 U18401 ( .IN1(n17689), .IN2(n17690), .QN(n17688) );
  NOR2X0 U18402 ( .IN1(n17691), .IN2(n17692), .QN(n17690) );
  NOR2X0 U18403 ( .IN1(n17693), .IN2(n17694), .QN(n17691) );
  NAND2X0 U18404 ( .IN1(n17695), .IN2(n17696), .QN(n17694) );
  NAND2X0 U18405 ( .IN1(n17697), .IN2(n17544), .QN(n17696) );
  NOR2X0 U18406 ( .IN1(n10366), .IN2(n10365), .QN(n17697) );
  NAND2X0 U18407 ( .IN1(n17698), .IN2(n17543), .QN(n17695) );
  NOR2X0 U18408 ( .IN1(n5701), .IN2(n10330), .QN(n17698) );
  NOR2X0 U18409 ( .IN1(n12454), .IN2(n17699), .QN(n17693) );
  NAND2X0 U18410 ( .IN1(g16775), .IN2(g3937), .QN(n17699) );
  NOR2X0 U18411 ( .IN1(n17700), .IN2(n17701), .QN(n17689) );
  INVX0 U18412 ( .INP(n17692), .ZN(n17701) );
  XNOR2X1 U18413 ( .IN1(g11418), .IN2(n5530), .Q(n17692) );
  NOR2X0 U18414 ( .IN1(n17702), .IN2(n17703), .QN(n17700) );
  NAND2X0 U18415 ( .IN1(n17704), .IN2(n17705), .QN(n17703) );
  NAND2X0 U18416 ( .IN1(n17706), .IN2(n17544), .QN(n17705) );
  NOR2X0 U18417 ( .IN1(n5701), .IN2(n10347), .QN(n17706) );
  NAND2X0 U18418 ( .IN1(n17707), .IN2(n13582), .QN(n17704) );
  NOR2X0 U18419 ( .IN1(n10379), .IN2(n10346), .QN(n17707) );
  NOR2X0 U18420 ( .IN1(n13579), .IN2(n17708), .QN(n17702) );
  NAND2X0 U18421 ( .IN1(g3961), .IN2(g16659), .QN(n17708) );
  NOR2X0 U18422 ( .IN1(n17709), .IN2(n17710), .QN(n17687) );
  NOR2X0 U18423 ( .IN1(n5530), .IN2(n17711), .QN(n17710) );
  NOR2X0 U18424 ( .IN1(n17712), .IN2(n17713), .QN(n17711) );
  NAND2X0 U18425 ( .IN1(n17714), .IN2(n17715), .QN(n17713) );
  NAND2X0 U18426 ( .IN1(n13582), .IN2(n17716), .QN(n17715) );
  NAND2X0 U18427 ( .IN1(n17717), .IN2(n17718), .QN(n17716) );
  NAND2X0 U18428 ( .IN1(g3917), .IN2(g16955), .QN(n17718) );
  NAND2X0 U18429 ( .IN1(g3893), .IN2(g11418), .QN(n17717) );
  NAND2X0 U18430 ( .IN1(n17540), .IN2(n17719), .QN(n17714) );
  NAND2X0 U18431 ( .IN1(n17720), .IN2(n17721), .QN(n17719) );
  NAND2X0 U18432 ( .IN1(g3965), .IN2(g16693), .QN(n17721) );
  NAND2X0 U18433 ( .IN1(test_so65), .IN2(g16748), .QN(n17720) );
  NAND2X0 U18434 ( .IN1(n17722), .IN2(n17723), .QN(n17712) );
  NAND2X0 U18435 ( .IN1(n17724), .IN2(n17543), .QN(n17723) );
  NOR2X0 U18436 ( .IN1(n5583), .IN2(n10435), .QN(n17724) );
  NAND2X0 U18437 ( .IN1(n17544), .IN2(n17725), .QN(n17722) );
  NAND2X0 U18438 ( .IN1(n17726), .IN2(n17727), .QN(n17725) );
  NAND2X0 U18439 ( .IN1(g3897), .IN2(g4031), .QN(n17727) );
  NAND2X0 U18440 ( .IN1(test_so24), .IN2(g14518), .QN(n17726) );
  NOR2X0 U18441 ( .IN1(n17728), .IN2(g4040), .QN(n17709) );
  NOR2X0 U18442 ( .IN1(n17729), .IN2(n17730), .QN(n17728) );
  NAND2X0 U18443 ( .IN1(n17731), .IN2(n17732), .QN(n17730) );
  NAND2X0 U18444 ( .IN1(n17543), .IN2(n17733), .QN(n17732) );
  NAND2X0 U18445 ( .IN1(n17734), .IN2(n17735), .QN(n17733) );
  NAND2X0 U18446 ( .IN1(g4031), .IN2(g3913), .QN(n17735) );
  NAND2X0 U18447 ( .IN1(g14518), .IN2(g3901), .QN(n17734) );
  INVX0 U18448 ( .INP(n13579), .ZN(n17543) );
  NAND2X0 U18449 ( .IN1(n5395), .IN2(g3990), .QN(n13579) );
  NAND2X0 U18450 ( .IN1(n17540), .IN2(n17736), .QN(n17731) );
  NAND2X0 U18451 ( .IN1(n17737), .IN2(n17738), .QN(n17736) );
  NAND2X0 U18452 ( .IN1(g16955), .IN2(g3925), .QN(n17738) );
  NAND2X0 U18453 ( .IN1(g3909), .IN2(g11418), .QN(n17737) );
  INVX0 U18454 ( .INP(n12454), .ZN(n17540) );
  NAND2X0 U18455 ( .IN1(g4054), .IN2(g3990), .QN(n12454) );
  NAND2X0 U18456 ( .IN1(n17739), .IN2(n17740), .QN(n17729) );
  NAND2X0 U18457 ( .IN1(n17741), .IN2(n17544), .QN(n17740) );
  NOR2X0 U18458 ( .IN1(g3990), .IN2(g4054), .QN(n17544) );
  NOR2X0 U18459 ( .IN1(n5583), .IN2(n10474), .QN(n17741) );
  NAND2X0 U18460 ( .IN1(n13582), .IN2(n17742), .QN(n17739) );
  NAND2X0 U18461 ( .IN1(n17743), .IN2(n17744), .QN(n17742) );
  NAND2X0 U18462 ( .IN1(g16748), .IN2(g3957), .QN(n17744) );
  NAND2X0 U18463 ( .IN1(g16693), .IN2(g3905), .QN(n17743) );
  NOR2X0 U18464 ( .IN1(g3990), .IN2(n5395), .QN(n13582) );
  INVX0 U18465 ( .INP(n13581), .ZN(n13583) );
  NAND2X0 U18466 ( .IN1(g4878), .IN2(n17745), .QN(n13581) );
  NAND2X0 U18467 ( .IN1(n17746), .IN2(n17578), .QN(n17745) );
  INVX0 U18468 ( .INP(n11391), .ZN(n17578) );
  NAND2X0 U18469 ( .IN1(g4975), .IN2(g4899), .QN(n11391) );
  NOR2X0 U18470 ( .IN1(n5614), .IN2(n17584), .QN(n17746) );
  NOR2X0 U18471 ( .IN1(n10309), .IN2(n10893), .QN(n17684) );
  NAND2X0 U18472 ( .IN1(n17747), .IN2(n17748), .QN(g28066) );
  NAND2X0 U18473 ( .IN1(n13608), .IN2(g3684), .QN(n17748) );
  NOR2X0 U18474 ( .IN1(n13605), .IN2(n11018), .QN(n13608) );
  NOR2X0 U18475 ( .IN1(n17749), .IN2(n17750), .QN(n17747) );
  NOR2X0 U18476 ( .IN1(n11037), .IN2(n17751), .QN(n17750) );
  NAND2X0 U18477 ( .IN1(n13605), .IN2(n16772), .QN(n17751) );
  NAND2X0 U18478 ( .IN1(n17752), .IN2(n17753), .QN(n16772) );
  NOR2X0 U18479 ( .IN1(n17754), .IN2(n17755), .QN(n17753) );
  NOR2X0 U18480 ( .IN1(n17756), .IN2(n17757), .QN(n17755) );
  NOR2X0 U18481 ( .IN1(n17758), .IN2(n17759), .QN(n17756) );
  NAND2X0 U18482 ( .IN1(n17760), .IN2(n17761), .QN(n17759) );
  NAND2X0 U18483 ( .IN1(n17762), .IN2(n17559), .QN(n17761) );
  NOR2X0 U18484 ( .IN1(n10369), .IN2(n10664), .QN(n17762) );
  NAND2X0 U18485 ( .IN1(n17763), .IN2(n17558), .QN(n17760) );
  NOR2X0 U18486 ( .IN1(n5699), .IN2(n10332), .QN(n17763) );
  NOR2X0 U18487 ( .IN1(n12450), .IN2(n17764), .QN(n17758) );
  NAND2X0 U18488 ( .IN1(g16744), .IN2(g3586), .QN(n17764) );
  NOR2X0 U18489 ( .IN1(n17765), .IN2(n17766), .QN(n17754) );
  INVX0 U18490 ( .INP(n17757), .ZN(n17766) );
  XNOR2X1 U18491 ( .IN1(g11388), .IN2(n5532), .Q(n17757) );
  NOR2X0 U18492 ( .IN1(n17767), .IN2(n17768), .QN(n17765) );
  NAND2X0 U18493 ( .IN1(n17769), .IN2(n17770), .QN(n17768) );
  NAND2X0 U18494 ( .IN1(n17771), .IN2(n17559), .QN(n17770) );
  NOR2X0 U18495 ( .IN1(n5699), .IN2(n10353), .QN(n17771) );
  NAND2X0 U18496 ( .IN1(n17772), .IN2(n13604), .QN(n17769) );
  NOR2X0 U18497 ( .IN1(n10383), .IN2(n10352), .QN(n17772) );
  NOR2X0 U18498 ( .IN1(n13601), .IN2(n17773), .QN(n17767) );
  NAND2X0 U18499 ( .IN1(g3610), .IN2(g16627), .QN(n17773) );
  NOR2X0 U18500 ( .IN1(n17774), .IN2(n17775), .QN(n17752) );
  NOR2X0 U18501 ( .IN1(n5532), .IN2(n17776), .QN(n17775) );
  NOR2X0 U18502 ( .IN1(n17777), .IN2(n17778), .QN(n17776) );
  NAND2X0 U18503 ( .IN1(n17779), .IN2(n17780), .QN(n17778) );
  NAND2X0 U18504 ( .IN1(n13604), .IN2(n17781), .QN(n17780) );
  NAND2X0 U18505 ( .IN1(n17782), .IN2(n17783), .QN(n17781) );
  NAND2X0 U18506 ( .IN1(g3566), .IN2(g16924), .QN(n17783) );
  NAND2X0 U18507 ( .IN1(g3542), .IN2(g11388), .QN(n17782) );
  NAND2X0 U18508 ( .IN1(n17555), .IN2(n17784), .QN(n17779) );
  NAND2X0 U18509 ( .IN1(n17785), .IN2(n17786), .QN(n17784) );
  NAND2X0 U18510 ( .IN1(g3614), .IN2(g16656), .QN(n17786) );
  NAND2X0 U18511 ( .IN1(g3598), .IN2(g16722), .QN(n17785) );
  NAND2X0 U18512 ( .IN1(n17787), .IN2(n17788), .QN(n17777) );
  NAND2X0 U18513 ( .IN1(n17789), .IN2(test_so26), .QN(n17788) );
  NOR2X0 U18514 ( .IN1(n10437), .IN2(n13601), .QN(n17789) );
  NAND2X0 U18515 ( .IN1(n17559), .IN2(n17790), .QN(n17787) );
  NAND2X0 U18516 ( .IN1(n17791), .IN2(n17792), .QN(n17790) );
  NAND2X0 U18517 ( .IN1(g3546), .IN2(g3680), .QN(n17792) );
  NAND2X0 U18518 ( .IN1(g3538), .IN2(g14451), .QN(n17791) );
  NOR2X0 U18519 ( .IN1(n17793), .IN2(g3689), .QN(n17774) );
  NOR2X0 U18520 ( .IN1(n17794), .IN2(n17795), .QN(n17793) );
  NAND2X0 U18521 ( .IN1(n17796), .IN2(n17797), .QN(n17795) );
  NAND2X0 U18522 ( .IN1(n17558), .IN2(n17798), .QN(n17797) );
  NAND2X0 U18523 ( .IN1(n17799), .IN2(n17800), .QN(n17798) );
  NAND2X0 U18524 ( .IN1(g3680), .IN2(g3562), .QN(n17800) );
  NAND2X0 U18525 ( .IN1(g14451), .IN2(g3550), .QN(n17799) );
  INVX0 U18526 ( .INP(n13601), .ZN(n17558) );
  NAND2X0 U18527 ( .IN1(n5399), .IN2(g3639), .QN(n13601) );
  NAND2X0 U18528 ( .IN1(n17555), .IN2(n17801), .QN(n17796) );
  NAND2X0 U18529 ( .IN1(n17802), .IN2(n17803), .QN(n17801) );
  NAND2X0 U18530 ( .IN1(g16924), .IN2(g3574), .QN(n17803) );
  NAND2X0 U18531 ( .IN1(g3558), .IN2(g11388), .QN(n17802) );
  INVX0 U18532 ( .INP(n12450), .ZN(n17555) );
  NAND2X0 U18533 ( .IN1(g3703), .IN2(g3639), .QN(n12450) );
  NAND2X0 U18534 ( .IN1(n17804), .IN2(n17805), .QN(n17794) );
  NAND2X0 U18535 ( .IN1(n17806), .IN2(test_so26), .QN(n17805) );
  NOR2X0 U18536 ( .IN1(n10484), .IN2(n17807), .QN(n17806) );
  INVX0 U18537 ( .INP(n17559), .ZN(n17807) );
  NOR2X0 U18538 ( .IN1(g3639), .IN2(g3703), .QN(n17559) );
  NAND2X0 U18539 ( .IN1(n13604), .IN2(n17808), .QN(n17804) );
  NAND2X0 U18540 ( .IN1(n17809), .IN2(n17810), .QN(n17808) );
  NAND2X0 U18541 ( .IN1(g16722), .IN2(g3606), .QN(n17810) );
  NAND2X0 U18542 ( .IN1(g16656), .IN2(g3554), .QN(n17809) );
  NOR2X0 U18543 ( .IN1(g3639), .IN2(n5399), .QN(n13604) );
  INVX0 U18544 ( .INP(n13603), .ZN(n13605) );
  NAND2X0 U18545 ( .IN1(g4871), .IN2(n17811), .QN(n13603) );
  NAND2X0 U18546 ( .IN1(n17812), .IN2(n11389), .QN(n17811) );
  INVX0 U18547 ( .INP(n11403), .ZN(n11389) );
  NAND2X0 U18548 ( .IN1(n5360), .IN2(g4899), .QN(n11403) );
  NOR2X0 U18549 ( .IN1(n5875), .IN2(n17584), .QN(n17812) );
  NOR2X0 U18550 ( .IN1(n10295), .IN2(n10893), .QN(n17749) );
  NAND2X0 U18551 ( .IN1(n17813), .IN2(n17814), .QN(g28063) );
  NAND2X0 U18552 ( .IN1(n13629), .IN2(g3333), .QN(n17814) );
  NOR2X0 U18553 ( .IN1(n13625), .IN2(n11018), .QN(n13629) );
  NOR2X0 U18554 ( .IN1(n17815), .IN2(n17816), .QN(n17813) );
  NOR2X0 U18555 ( .IN1(n11037), .IN2(n17817), .QN(n17816) );
  NAND2X0 U18556 ( .IN1(n13625), .IN2(n16812), .QN(n17817) );
  NAND2X0 U18557 ( .IN1(n17818), .IN2(n17819), .QN(n16812) );
  NOR2X0 U18558 ( .IN1(n17820), .IN2(n17821), .QN(n17819) );
  NOR2X0 U18559 ( .IN1(n17822), .IN2(n17823), .QN(n17821) );
  NOR2X0 U18560 ( .IN1(n17824), .IN2(n17825), .QN(n17822) );
  NAND2X0 U18561 ( .IN1(n17826), .IN2(n17827), .QN(n17825) );
  NAND2X0 U18562 ( .IN1(n17828), .IN2(n17574), .QN(n17827) );
  NOR2X0 U18563 ( .IN1(n10358), .IN2(n10357), .QN(n17828) );
  NAND2X0 U18564 ( .IN1(n17829), .IN2(n13620), .QN(n17826) );
  NOR2X0 U18565 ( .IN1(n5702), .IN2(n10327), .QN(n17829) );
  NOR2X0 U18566 ( .IN1(n12442), .IN2(n17830), .QN(n17824) );
  NAND2X0 U18567 ( .IN1(g16718), .IN2(g3235), .QN(n17830) );
  NOR2X0 U18568 ( .IN1(n17831), .IN2(n17832), .QN(n17820) );
  INVX0 U18569 ( .INP(n17823), .ZN(n17832) );
  XNOR2X1 U18570 ( .IN1(g11349), .IN2(n5527), .Q(n17823) );
  NOR2X0 U18571 ( .IN1(n17833), .IN2(n17834), .QN(n17831) );
  NAND2X0 U18572 ( .IN1(n17835), .IN2(n17836), .QN(n17834) );
  NAND2X0 U18573 ( .IN1(n17837), .IN2(n17574), .QN(n17836) );
  NOR2X0 U18574 ( .IN1(n5702), .IN2(n10335), .QN(n17837) );
  NAND2X0 U18575 ( .IN1(n17838), .IN2(n13624), .QN(n17835) );
  NOR2X0 U18576 ( .IN1(n10372), .IN2(n10334), .QN(n17838) );
  NOR2X0 U18577 ( .IN1(n17839), .IN2(n17840), .QN(n17833) );
  NAND2X0 U18578 ( .IN1(test_so84), .IN2(g16603), .QN(n17840) );
  NOR2X0 U18579 ( .IN1(n17841), .IN2(n17842), .QN(n17818) );
  NOR2X0 U18580 ( .IN1(n5527), .IN2(n17843), .QN(n17842) );
  NOR2X0 U18581 ( .IN1(n17844), .IN2(n17845), .QN(n17843) );
  NAND2X0 U18582 ( .IN1(n17846), .IN2(n17847), .QN(n17845) );
  NAND2X0 U18583 ( .IN1(n13624), .IN2(n17848), .QN(n17847) );
  NAND2X0 U18584 ( .IN1(n17849), .IN2(n17850), .QN(n17848) );
  NAND2X0 U18585 ( .IN1(g3215), .IN2(g16874), .QN(n17850) );
  NAND2X0 U18586 ( .IN1(g3191), .IN2(g11349), .QN(n17849) );
  NAND2X0 U18587 ( .IN1(n17571), .IN2(n17851), .QN(n17846) );
  NAND2X0 U18588 ( .IN1(n17852), .IN2(n17853), .QN(n17851) );
  NAND2X0 U18589 ( .IN1(g3263), .IN2(g16624), .QN(n17853) );
  NAND2X0 U18590 ( .IN1(g3247), .IN2(g16686), .QN(n17852) );
  NAND2X0 U18591 ( .IN1(n17854), .IN2(n17855), .QN(n17844) );
  NAND2X0 U18592 ( .IN1(n17856), .IN2(n13620), .QN(n17855) );
  NOR2X0 U18593 ( .IN1(n5580), .IN2(n10431), .QN(n17856) );
  NAND2X0 U18594 ( .IN1(n17574), .IN2(n17857), .QN(n17854) );
  NAND2X0 U18595 ( .IN1(n17858), .IN2(n17859), .QN(n17857) );
  NAND2X0 U18596 ( .IN1(g3187), .IN2(g14421), .QN(n17859) );
  NAND2X0 U18597 ( .IN1(test_so91), .IN2(test_so88), .QN(n17858) );
  NOR2X0 U18598 ( .IN1(n17860), .IN2(g3338), .QN(n17841) );
  NOR2X0 U18599 ( .IN1(n17861), .IN2(n17862), .QN(n17860) );
  NAND2X0 U18600 ( .IN1(n17863), .IN2(n17864), .QN(n17862) );
  NAND2X0 U18601 ( .IN1(n13620), .IN2(n17865), .QN(n17864) );
  NAND2X0 U18602 ( .IN1(n17866), .IN2(n17867), .QN(n17865) );
  NAND2X0 U18603 ( .IN1(test_so91), .IN2(g3211), .QN(n17867) );
  NAND2X0 U18604 ( .IN1(g14421), .IN2(g3199), .QN(n17866) );
  INVX0 U18605 ( .INP(n17839), .ZN(n13620) );
  NAND2X0 U18606 ( .IN1(n5604), .IN2(g3288), .QN(n17839) );
  NAND2X0 U18607 ( .IN1(n17571), .IN2(n17868), .QN(n17863) );
  NAND2X0 U18608 ( .IN1(n17869), .IN2(n17870), .QN(n17868) );
  NAND2X0 U18609 ( .IN1(g16874), .IN2(g3223), .QN(n17870) );
  NAND2X0 U18610 ( .IN1(g3207), .IN2(g11349), .QN(n17869) );
  INVX0 U18611 ( .INP(n12442), .ZN(n17571) );
  NAND2X0 U18612 ( .IN1(g3288), .IN2(g3352), .QN(n12442) );
  NAND2X0 U18613 ( .IN1(n17871), .IN2(n17872), .QN(n17861) );
  NAND2X0 U18614 ( .IN1(n17873), .IN2(n17574), .QN(n17872) );
  NOR2X0 U18615 ( .IN1(g3288), .IN2(g3352), .QN(n17574) );
  NOR2X0 U18616 ( .IN1(n5580), .IN2(n10455), .QN(n17873) );
  NAND2X0 U18617 ( .IN1(n13624), .IN2(n17874), .QN(n17871) );
  NAND2X0 U18618 ( .IN1(n17875), .IN2(n17876), .QN(n17874) );
  NAND2X0 U18619 ( .IN1(g16686), .IN2(g3255), .QN(n17876) );
  NAND2X0 U18620 ( .IN1(g16624), .IN2(g3203), .QN(n17875) );
  NOR2X0 U18621 ( .IN1(g3288), .IN2(n5604), .QN(n13624) );
  INVX0 U18622 ( .INP(n13626), .ZN(n13625) );
  NAND2X0 U18623 ( .IN1(g4864), .IN2(n17877), .QN(n13626) );
  NAND2X0 U18624 ( .IN1(n17878), .IN2(n11388), .QN(n17877) );
  INVX0 U18625 ( .INP(n11402), .ZN(n11388) );
  NAND2X0 U18626 ( .IN1(n5517), .IN2(g4975), .QN(n11402) );
  NOR2X0 U18627 ( .IN1(n5878), .IN2(n17584), .QN(n17878) );
  NAND2X0 U18628 ( .IN1(n17879), .IN2(n17880), .QN(n17584) );
  NOR2X0 U18629 ( .IN1(n10542), .IN2(n17579), .QN(n17880) );
  NAND2X0 U18630 ( .IN1(n10652), .IN2(g4966), .QN(n17579) );
  NOR2X0 U18631 ( .IN1(g4983), .IN2(n17881), .QN(n17879) );
  NAND2X0 U18632 ( .IN1(g4859), .IN2(g4843), .QN(n17881) );
  NOR2X0 U18633 ( .IN1(n10284), .IN2(n10893), .QN(n17815) );
  NAND2X0 U18634 ( .IN1(n17882), .IN2(n17883), .QN(g28060) );
  NOR2X0 U18635 ( .IN1(n17884), .IN2(n17885), .QN(n17883) );
  NOR2X0 U18636 ( .IN1(n5301), .IN2(n10894), .QN(n17885) );
  NOR2X0 U18637 ( .IN1(n11037), .IN2(n17886), .QN(n17884) );
  NAND2X0 U18638 ( .IN1(n16822), .IN2(g2729), .QN(n17886) );
  NOR2X0 U18639 ( .IN1(n2787), .IN2(n17887), .QN(n17882) );
  NOR2X0 U18640 ( .IN1(g2729), .IN2(n16822), .QN(n17887) );
  NAND2X0 U18641 ( .IN1(n16065), .IN2(g2724), .QN(n16822) );
  INVX0 U18642 ( .INP(n14448), .ZN(n2787) );
  INVX0 U18643 ( .INP(n17888), .ZN(g28059) );
  NOR2X0 U18644 ( .IN1(n17889), .IN2(n17890), .QN(n17888) );
  NAND2X0 U18645 ( .IN1(n17891), .IN2(n17892), .QN(n17890) );
  NAND2X0 U18646 ( .IN1(n17893), .IN2(n16424), .QN(n17892) );
  INVX0 U18647 ( .INP(n17894), .ZN(n17893) );
  NAND2X0 U18648 ( .IN1(n10249), .IN2(n14739), .QN(n17894) );
  NOR2X0 U18649 ( .IN1(n14126), .IN2(n11019), .QN(n14739) );
  NAND2X0 U18650 ( .IN1(n17895), .IN2(n17896), .QN(n14126) );
  NOR2X0 U18651 ( .IN1(n17897), .IN2(n17898), .QN(n17896) );
  NOR2X0 U18652 ( .IN1(n17899), .IN2(n17900), .QN(n17898) );
  NOR2X0 U18653 ( .IN1(g1351), .IN2(n17901), .QN(n17897) );
  NOR2X0 U18654 ( .IN1(n17902), .IN2(g1312), .QN(n17895) );
  NAND2X0 U18655 ( .IN1(n4798), .IN2(n17903), .QN(n17891) );
  NOR2X0 U18656 ( .IN1(n5322), .IN2(n10894), .QN(n17889) );
  NAND2X0 U18657 ( .IN1(n17904), .IN2(n17905), .QN(g28058) );
  NAND2X0 U18658 ( .IN1(test_so77), .IN2(n11081), .QN(n17905) );
  NOR2X0 U18659 ( .IN1(n17906), .IN2(n17907), .QN(n17904) );
  NOR2X0 U18660 ( .IN1(g1252), .IN2(n17908), .QN(n17907) );
  NOR2X0 U18661 ( .IN1(n5554), .IN2(n17909), .QN(n17906) );
  NAND2X0 U18662 ( .IN1(n14133), .IN2(n17908), .QN(n17909) );
  INVX0 U18663 ( .INP(n4490), .ZN(n17908) );
  INVX0 U18664 ( .INP(n17910), .ZN(g28057) );
  NOR2X0 U18665 ( .IN1(n17911), .IN2(n17912), .QN(n17910) );
  NAND2X0 U18666 ( .IN1(n17913), .IN2(n17914), .QN(n17912) );
  NAND2X0 U18667 ( .IN1(n17915), .IN2(n16468), .QN(n17914) );
  INVX0 U18668 ( .INP(n17916), .ZN(n17915) );
  NAND2X0 U18669 ( .IN1(n10250), .IN2(n14756), .QN(n17916) );
  NOR2X0 U18670 ( .IN1(n14145), .IN2(n11019), .QN(n14756) );
  NAND2X0 U18671 ( .IN1(n17917), .IN2(n17918), .QN(n14145) );
  NOR2X0 U18672 ( .IN1(n17919), .IN2(n17920), .QN(n17918) );
  NOR2X0 U18673 ( .IN1(n17921), .IN2(g1008), .QN(n17920) );
  NOR2X0 U18674 ( .IN1(n17922), .IN2(n17923), .QN(n17919) );
  NOR2X0 U18675 ( .IN1(test_so20), .IN2(n17924), .QN(n17917) );
  NAND2X0 U18676 ( .IN1(n4805), .IN2(n17925), .QN(n17913) );
  NOR2X0 U18677 ( .IN1(n5321), .IN2(n10894), .QN(n17911) );
  NAND2X0 U18678 ( .IN1(n17926), .IN2(n17927), .QN(g28056) );
  NAND2X0 U18679 ( .IN1(n11063), .IN2(g936), .QN(n17927) );
  NOR2X0 U18680 ( .IN1(n17928), .IN2(n17929), .QN(n17926) );
  NOR2X0 U18681 ( .IN1(g907), .IN2(n17930), .QN(n17929) );
  NOR2X0 U18682 ( .IN1(n5555), .IN2(n17931), .QN(n17928) );
  NAND2X0 U18683 ( .IN1(n14152), .IN2(n17930), .QN(n17931) );
  INVX0 U18684 ( .INP(n4514), .ZN(n17930) );
  NAND2X0 U18685 ( .IN1(n17932), .IN2(n17933), .QN(g28055) );
  NAND2X0 U18686 ( .IN1(n11063), .IN2(g822), .QN(n17933) );
  NOR2X0 U18687 ( .IN1(n17934), .IN2(n17935), .QN(n17932) );
  NOR2X0 U18688 ( .IN1(g827), .IN2(n17936), .QN(n17935) );
  NAND2X0 U18689 ( .IN1(n4519), .IN2(n17117), .QN(n17936) );
  NOR2X0 U18690 ( .IN1(n5728), .IN2(n17937), .QN(n17934) );
  NAND2X0 U18691 ( .IN1(n4518), .IN2(n17938), .QN(n17937) );
  INVX0 U18692 ( .INP(n4519), .ZN(n17938) );
  NAND2X0 U18693 ( .IN1(n17939), .IN2(n17940), .QN(g28054) );
  NAND2X0 U18694 ( .IN1(n17941), .IN2(g728), .QN(n17940) );
  NAND2X0 U18695 ( .IN1(n17942), .IN2(g661), .QN(n17939) );
  NAND2X0 U18696 ( .IN1(n17943), .IN2(n17944), .QN(g28053) );
  NAND2X0 U18697 ( .IN1(n11063), .IN2(g681), .QN(n17944) );
  NOR2X0 U18698 ( .IN1(n17945), .IN2(n17946), .QN(n17943) );
  NOR2X0 U18699 ( .IN1(n10659), .IN2(n17947), .QN(n17946) );
  NAND2X0 U18700 ( .IN1(n17948), .IN2(n17949), .QN(g28052) );
  NAND2X0 U18701 ( .IN1(n17941), .IN2(g661), .QN(n17949) );
  NAND2X0 U18702 ( .IN1(n17942), .IN2(g718), .QN(n17948) );
  NAND2X0 U18703 ( .IN1(n17950), .IN2(n17951), .QN(g28051) );
  NAND2X0 U18704 ( .IN1(n17941), .IN2(g718), .QN(n17951) );
  NAND2X0 U18705 ( .IN1(n17942), .IN2(g655), .QN(n17950) );
  NAND2X0 U18706 ( .IN1(n17952), .IN2(n17953), .QN(g28050) );
  NAND2X0 U18707 ( .IN1(n17941), .IN2(g655), .QN(n17953) );
  NAND2X0 U18708 ( .IN1(n17942), .IN2(g650), .QN(n17952) );
  NAND2X0 U18709 ( .IN1(n17954), .IN2(n17955), .QN(g28049) );
  NAND2X0 U18710 ( .IN1(test_so87), .IN2(n11080), .QN(n17955) );
  NOR2X0 U18711 ( .IN1(n17956), .IN2(n17957), .QN(n17954) );
  NOR2X0 U18712 ( .IN1(n10270), .IN2(n17942), .QN(n17957) );
  NOR2X0 U18713 ( .IN1(n10233), .IN2(n17958), .QN(n17956) );
  INVX0 U18714 ( .INP(n17945), .ZN(n17958) );
  NAND2X0 U18715 ( .IN1(n17959), .IN2(n17960), .QN(g28048) );
  NAND2X0 U18716 ( .IN1(n11063), .IN2(g29212), .QN(n17960) );
  NOR2X0 U18717 ( .IN1(n17961), .IN2(n17962), .QN(n17959) );
  NOR2X0 U18718 ( .IN1(n4819), .IN2(n17963), .QN(n17962) );
  NAND2X0 U18719 ( .IN1(n17964), .IN2(n17965), .QN(n4819) );
  NOR2X0 U18720 ( .IN1(n5821), .IN2(n17152), .QN(n17965) );
  NAND2X0 U18721 ( .IN1(n17966), .IN2(n17967), .QN(n17152) );
  NOR2X0 U18722 ( .IN1(g645), .IN2(g650), .QN(n17967) );
  NOR2X0 U18723 ( .IN1(n10659), .IN2(n17968), .QN(n17966) );
  XOR2X1 U18724 ( .IN1(n10283), .IN2(n10282), .Q(n17968) );
  NOR2X0 U18725 ( .IN1(n17969), .IN2(g691), .QN(n17964) );
  INVX0 U18726 ( .INP(n5112), .ZN(n17969) );
  NOR2X0 U18727 ( .IN1(n5520), .IN2(n17970), .QN(n17961) );
  INVX0 U18728 ( .INP(n17971), .ZN(n17970) );
  NAND2X0 U18729 ( .IN1(n17972), .IN2(n17973), .QN(n17971) );
  NAND2X0 U18730 ( .IN1(n10928), .IN2(n17974), .QN(n17972) );
  NOR2X0 U18731 ( .IN1(n5821), .IN2(test_so70), .QN(n17974) );
  NAND2X0 U18732 ( .IN1(n17975), .IN2(n17976), .QN(g28047) );
  NAND2X0 U18733 ( .IN1(n17941), .IN2(g681), .QN(n17976) );
  NAND2X0 U18734 ( .IN1(n17942), .IN2(g645), .QN(n17975) );
  NAND2X0 U18735 ( .IN1(n17977), .IN2(n17978), .QN(g28046) );
  NAND2X0 U18736 ( .IN1(n17945), .IN2(g446), .QN(n17978) );
  NOR2X0 U18737 ( .IN1(n17979), .IN2(n11020), .QN(n17945) );
  NAND2X0 U18738 ( .IN1(n17941), .IN2(g645), .QN(n17977) );
  INVX0 U18739 ( .INP(n17942), .ZN(n17941) );
  NAND2X0 U18740 ( .IN1(n17979), .IN2(n10969), .QN(n17942) );
  NAND2X0 U18741 ( .IN1(n17980), .IN2(n17981), .QN(n17979) );
  NOR2X0 U18742 ( .IN1(n17982), .IN2(n17983), .QN(n17981) );
  NOR2X0 U18743 ( .IN1(n17984), .IN2(g691), .QN(n17983) );
  NOR2X0 U18744 ( .IN1(g424), .IN2(n17985), .QN(n17984) );
  NAND2X0 U18745 ( .IN1(n5629), .IN2(g417), .QN(n17985) );
  NOR2X0 U18746 ( .IN1(n5520), .IN2(n17986), .QN(n17982) );
  NOR2X0 U18747 ( .IN1(n1192), .IN2(g370), .QN(n17980) );
  NAND2X0 U18748 ( .IN1(n17987), .IN2(n17988), .QN(g28045) );
  NAND2X0 U18749 ( .IN1(n11063), .IN2(g568), .QN(n17988) );
  NOR2X0 U18750 ( .IN1(n17989), .IN2(n17990), .QN(n17987) );
  NOR2X0 U18751 ( .IN1(g572), .IN2(n17991), .QN(n17990) );
  NOR2X0 U18752 ( .IN1(n5337), .IN2(n17992), .QN(n17989) );
  NAND2X0 U18753 ( .IN1(n2421), .IN2(n17991), .QN(n17992) );
  INVX0 U18754 ( .INP(n4537), .ZN(n17991) );
  NAND2X0 U18755 ( .IN1(n17993), .IN2(n17994), .QN(g28044) );
  NAND2X0 U18756 ( .IN1(n11063), .IN2(g528), .QN(n17994) );
  NAND2X0 U18757 ( .IN1(n17995), .IN2(n10969), .QN(n17993) );
  NAND2X0 U18758 ( .IN1(n17996), .IN2(n17997), .QN(n17995) );
  XOR2X1 U18759 ( .IN1(n5820), .IN2(n17167), .Q(n17996) );
  NOR2X0 U18760 ( .IN1(n17998), .IN2(n17999), .QN(n17167) );
  NAND2X0 U18761 ( .IN1(n18000), .IN2(n18001), .QN(n17998) );
  NAND2X0 U18762 ( .IN1(n18002), .IN2(n5327), .QN(n18000) );
  NAND2X0 U18763 ( .IN1(n12082), .IN2(n5630), .QN(g28042) );
  NOR2X0 U18764 ( .IN1(n11038), .IN2(g1306), .QN(n12082) );
  NAND2X0 U18765 ( .IN1(n18003), .IN2(n11987), .QN(g28041) );
  INVX0 U18766 ( .INP(n12087), .ZN(n11987) );
  NOR2X0 U18767 ( .IN1(n10606), .IN2(n18004), .QN(n12087) );
  NOR2X0 U18768 ( .IN1(n11038), .IN2(n14746), .QN(n18003) );
  INVX0 U18769 ( .INP(n11986), .ZN(n14746) );
  NAND2X0 U18770 ( .IN1(n4836), .IN2(g1536), .QN(n11986) );
  NAND2X0 U18771 ( .IN1(n18005), .IN2(n18006), .QN(g28030) );
  NAND2X0 U18772 ( .IN1(n18007), .IN2(n5882), .QN(n18006) );
  NOR2X0 U18773 ( .IN1(n18008), .IN2(g3129), .QN(n18007) );
  NOR2X0 U18774 ( .IN1(n18009), .IN2(n18010), .QN(n18008) );
  NOR2X0 U18775 ( .IN1(n12017), .IN2(n18011), .QN(n18009) );
  NOR2X0 U18776 ( .IN1(n18012), .IN2(n18013), .QN(n18011) );
  NOR2X0 U18777 ( .IN1(n18014), .IN2(n18015), .QN(n18013) );
  NOR2X0 U18778 ( .IN1(g3845), .IN2(n18016), .QN(n18012) );
  NAND2X0 U18779 ( .IN1(n5872), .IN2(n18017), .QN(n18016) );
  NAND2X0 U18780 ( .IN1(n18018), .IN2(n18015), .QN(n18017) );
  INVX0 U18781 ( .INP(n18019), .ZN(n18015) );
  NAND2X0 U18782 ( .IN1(n18020), .IN2(n18021), .QN(n18018) );
  NAND2X0 U18783 ( .IN1(n18022), .IN2(n18023), .QN(n18021) );
  NAND2X0 U18784 ( .IN1(n18024), .IN2(n18025), .QN(n18022) );
  NOR2X0 U18785 ( .IN1(n18026), .IN2(n18027), .QN(n18024) );
  INVX0 U18786 ( .INP(n18028), .ZN(n18027) );
  NAND2X0 U18787 ( .IN1(n18029), .IN2(n18030), .QN(n18028) );
  NOR2X0 U18788 ( .IN1(n18031), .IN2(n18032), .QN(n18026) );
  INVX0 U18789 ( .INP(n18033), .ZN(n12017) );
  NAND2X0 U18790 ( .IN1(n18010), .IN2(n18033), .QN(n18005) );
  NAND2X0 U18791 ( .IN1(n18034), .IN2(n10969), .QN(n18033) );
  NAND2X0 U18792 ( .IN1(n5889), .IN2(n5868), .QN(n18034) );
  INVX0 U18793 ( .INP(n12018), .ZN(n18010) );
  NAND2X0 U18794 ( .IN1(n18035), .IN2(n18019), .QN(n12018) );
  NOR2X0 U18795 ( .IN1(n18023), .IN2(n18036), .QN(n18019) );
  NOR2X0 U18796 ( .IN1(n18025), .IN2(n11021), .QN(n18036) );
  NOR2X0 U18797 ( .IN1(g5499), .IN2(g5485), .QN(n18025) );
  NAND2X0 U18798 ( .IN1(n18031), .IN2(n18032), .QN(n18023) );
  NAND2X0 U18799 ( .IN1(n18037), .IN2(n10969), .QN(n18032) );
  NAND2X0 U18800 ( .IN1(n5888), .IN2(n5874), .QN(n18037) );
  NOR2X0 U18801 ( .IN1(n18030), .IN2(n18029), .QN(n18031) );
  NOR2X0 U18802 ( .IN1(n18038), .IN2(n11022), .QN(n18029) );
  NOR2X0 U18803 ( .IN1(g6537), .IN2(g6523), .QN(n18038) );
  NOR2X0 U18804 ( .IN1(n18039), .IN2(n11022), .QN(n18030) );
  NOR2X0 U18805 ( .IN1(g5831), .IN2(test_so83), .QN(n18039) );
  NOR2X0 U18806 ( .IN1(n18014), .IN2(n18040), .QN(n18035) );
  NOR2X0 U18807 ( .IN1(n11039), .IN2(n18041), .QN(n18040) );
  NOR2X0 U18808 ( .IN1(g3831), .IN2(g3845), .QN(n18041) );
  INVX0 U18809 ( .INP(n18020), .ZN(n18014) );
  NAND2X0 U18810 ( .IN1(n18042), .IN2(n10970), .QN(n18020) );
  NAND2X0 U18811 ( .IN1(n5883), .IN2(n5871), .QN(n18042) );
  NAND2X0 U18812 ( .IN1(n18043), .IN2(n13567), .QN(g26971) );
  NAND2X0 U18813 ( .IN1(n5670), .IN2(n10970), .QN(n13567) );
  NOR2X0 U18814 ( .IN1(n18044), .IN2(n18045), .QN(n18043) );
  NOR2X0 U18815 ( .IN1(n10265), .IN2(n10895), .QN(n18045) );
  NOR2X0 U18816 ( .IN1(n11039), .IN2(g4531), .QN(n18044) );
  NAND2X0 U18817 ( .IN1(n18046), .IN2(n18047), .QN(g26970) );
  NAND2X0 U18818 ( .IN1(n10929), .IN2(g4473), .QN(n18047) );
  NAND2X0 U18819 ( .IN1(n11064), .IN2(g4459), .QN(n18046) );
  NAND2X0 U18820 ( .IN1(n18048), .IN2(n18049), .QN(g26969) );
  NAND2X0 U18821 ( .IN1(n11064), .IN2(g4462), .QN(n18049) );
  NAND2X0 U18822 ( .IN1(n18050), .IN2(n10970), .QN(n18048) );
  NOR2X0 U18823 ( .IN1(test_so38), .IN2(g4473), .QN(n18050) );
  NAND2X0 U18824 ( .IN1(n18051), .IN2(n18052), .QN(g26968) );
  NAND2X0 U18825 ( .IN1(n11064), .IN2(g4558), .QN(n18051) );
  NAND2X0 U18826 ( .IN1(n18053), .IN2(n18054), .QN(g26967) );
  NAND2X0 U18827 ( .IN1(n11064), .IN2(g4561), .QN(n18053) );
  NAND2X0 U18828 ( .IN1(n18055), .IN2(n18056), .QN(g26966) );
  NAND2X0 U18829 ( .IN1(n11064), .IN2(g4555), .QN(n18055) );
  XOR2X1 U18830 ( .IN1(DFF_228_n1), .IN2(n18057), .Q(g26965) );
  NAND2X0 U18831 ( .IN1(n10929), .IN2(g10306), .QN(n18057) );
  INVX0 U18832 ( .INP(n18058), .ZN(g26964) );
  NOR2X0 U18833 ( .IN1(n18059), .IN2(n18060), .QN(n18058) );
  NOR2X0 U18834 ( .IN1(n10907), .IN2(n10550), .QN(n18060) );
  NOR2X0 U18835 ( .IN1(n18061), .IN2(n11014), .QN(n18059) );
  NOR2X0 U18836 ( .IN1(n18062), .IN2(n18063), .QN(n18061) );
  NOR2X0 U18837 ( .IN1(n10533), .IN2(n5752), .QN(n18063) );
  NOR2X0 U18838 ( .IN1(g4521), .IN2(n17641), .QN(n18062) );
  XNOR2X1 U18839 ( .IN1(n12762), .IN2(n10550), .Q(n17641) );
  NAND2X0 U18840 ( .IN1(n18064), .IN2(n18065), .QN(n12762) );
  NOR2X0 U18841 ( .IN1(n10541), .IN2(n10540), .QN(n18065) );
  NOR2X0 U18842 ( .IN1(n10539), .IN2(n10692), .QN(n18064) );
  NAND2X0 U18843 ( .IN1(n18066), .IN2(n18054), .QN(g26963) );
  NAND2X0 U18844 ( .IN1(g6750), .IN2(n10970), .QN(n18054) );
  NAND2X0 U18845 ( .IN1(n11064), .IN2(g4489), .QN(n18066) );
  NAND2X0 U18846 ( .IN1(n18052), .IN2(n18067), .QN(g26962) );
  NAND2X0 U18847 ( .IN1(test_so27), .IN2(n11080), .QN(n18067) );
  NAND2X0 U18848 ( .IN1(g6749), .IN2(n10970), .QN(n18052) );
  NAND2X0 U18849 ( .IN1(n18068), .IN2(n18056), .QN(g26961) );
  NAND2X0 U18850 ( .IN1(g6748), .IN2(n10970), .QN(n18056) );
  INVX0 U18851 ( .INP(n18069), .ZN(n18068) );
  NOR2X0 U18852 ( .IN1(n10905), .IN2(n10539), .QN(n18069) );
  NAND2X0 U18853 ( .IN1(n18070), .IN2(n18071), .QN(g26958) );
  NAND2X0 U18854 ( .IN1(n11064), .IN2(g4455), .QN(n18071) );
  NAND2X0 U18855 ( .IN1(n18072), .IN2(n18073), .QN(g26957) );
  NAND2X0 U18856 ( .IN1(n18074), .IN2(g4434), .QN(n18073) );
  NAND2X0 U18857 ( .IN1(n18075), .IN2(n10970), .QN(n18074) );
  NAND2X0 U18858 ( .IN1(n18076), .IN2(g4392), .QN(n18075) );
  NAND2X0 U18859 ( .IN1(test_so47), .IN2(n10971), .QN(n18072) );
  NAND2X0 U18860 ( .IN1(n19410), .IN2(n18077), .QN(g26956) );
  NAND2X0 U18861 ( .IN1(n18078), .IN2(n18079), .QN(n18077) );
  NOR2X0 U18862 ( .IN1(n10184), .IN2(n18080), .QN(n18078) );
  NAND2X0 U18863 ( .IN1(n18081), .IN2(n18082), .QN(g26955) );
  NAND2X0 U18864 ( .IN1(n18083), .IN2(n18076), .QN(n18082) );
  INVX0 U18865 ( .INP(n18080), .ZN(n18076) );
  NAND2X0 U18866 ( .IN1(n18084), .IN2(g4438), .QN(n18081) );
  NAND2X0 U18867 ( .IN1(n18085), .IN2(n18086), .QN(g26954) );
  NAND2X0 U18868 ( .IN1(test_so47), .IN2(n11081), .QN(n18086) );
  NOR2X0 U18869 ( .IN1(n18087), .IN2(n18088), .QN(n18085) );
  NOR2X0 U18870 ( .IN1(n10538), .IN2(n18084), .QN(n18088) );
  NOR2X0 U18871 ( .IN1(n18080), .IN2(n18089), .QN(n18087) );
  NAND2X0 U18872 ( .IN1(n18090), .IN2(n18091), .QN(n18080) );
  INVX0 U18873 ( .INP(n18092), .ZN(n18091) );
  NAND2X0 U18874 ( .IN1(n19410), .IN2(n18093), .QN(n18092) );
  NOR2X0 U18875 ( .IN1(g4438), .IN2(test_so47), .QN(n18093) );
  NOR2X0 U18876 ( .IN1(g7245), .IN2(g7260), .QN(n18090) );
  NAND2X0 U18877 ( .IN1(n18094), .IN2(n18095), .QN(g26952) );
  NAND2X0 U18878 ( .IN1(n18096), .IN2(g4430), .QN(n18095) );
  NAND2X0 U18879 ( .IN1(n10929), .IN2(g4388), .QN(n18096) );
  NAND2X0 U18880 ( .IN1(n18097), .IN2(n10971), .QN(n18094) );
  NAND2X0 U18881 ( .IN1(n18098), .IN2(n18099), .QN(n18097) );
  NAND2X0 U18882 ( .IN1(n10184), .IN2(g4388), .QN(n18099) );
  XOR2X1 U18883 ( .IN1(g4401), .IN2(n10180), .Q(n18098) );
  NAND2X0 U18884 ( .IN1(n18070), .IN2(n18100), .QN(g26950) );
  NAND2X0 U18885 ( .IN1(n11064), .IN2(g4417), .QN(n18100) );
  NAND2X0 U18886 ( .IN1(n18101), .IN2(n10971), .QN(n18070) );
  NAND2X0 U18887 ( .IN1(n18102), .IN2(n18103), .QN(n18101) );
  NAND2X0 U18888 ( .IN1(n18104), .IN2(g4392), .QN(n18103) );
  NAND2X0 U18889 ( .IN1(n18105), .IN2(n18106), .QN(g26949) );
  NAND2X0 U18890 ( .IN1(n18107), .IN2(g4401), .QN(n18106) );
  NAND2X0 U18891 ( .IN1(n18108), .IN2(n10971), .QN(n18107) );
  NAND2X0 U18892 ( .IN1(n18109), .IN2(g4392), .QN(n18108) );
  NAND2X0 U18893 ( .IN1(n10929), .IN2(g4411), .QN(n18105) );
  NAND2X0 U18894 ( .IN1(n10622), .IN2(n18110), .QN(g26948) );
  NAND2X0 U18895 ( .IN1(n18111), .IN2(n18079), .QN(n18110) );
  INVX0 U18896 ( .INP(n18089), .ZN(n18079) );
  NOR2X0 U18897 ( .IN1(n10181), .IN2(n18104), .QN(n18111) );
  NAND2X0 U18898 ( .IN1(n18112), .IN2(n18113), .QN(g26947) );
  NAND2X0 U18899 ( .IN1(n11064), .IN2(g4388), .QN(n18113) );
  NAND2X0 U18900 ( .IN1(n18114), .IN2(n10971), .QN(n18112) );
  NAND2X0 U18901 ( .IN1(n18102), .IN2(n18115), .QN(n18114) );
  NAND2X0 U18902 ( .IN1(n18116), .IN2(n18104), .QN(n18115) );
  XOR2X1 U18903 ( .IN1(n5714), .IN2(n10621), .Q(n18116) );
  NAND2X0 U18904 ( .IN1(n18117), .IN2(n5710), .QN(n18102) );
  NOR2X0 U18905 ( .IN1(n18104), .IN2(g4417), .QN(n18117) );
  NAND2X0 U18906 ( .IN1(n18118), .IN2(n18119), .QN(g26946) );
  NAND2X0 U18907 ( .IN1(n18083), .IN2(n18109), .QN(n18119) );
  INVX0 U18908 ( .INP(n18104), .ZN(n18109) );
  NOR2X0 U18909 ( .IN1(n5710), .IN2(n11014), .QN(n18083) );
  NAND2X0 U18910 ( .IN1(n18084), .IN2(g4375), .QN(n18118) );
  NAND2X0 U18911 ( .IN1(n18120), .IN2(n18121), .QN(g26945) );
  NAND2X0 U18912 ( .IN1(n11065), .IN2(g4411), .QN(n18121) );
  NOR2X0 U18913 ( .IN1(n18122), .IN2(n18123), .QN(n18120) );
  NOR2X0 U18914 ( .IN1(n10621), .IN2(n18084), .QN(n18123) );
  NAND2X0 U18915 ( .IN1(n5714), .IN2(n10971), .QN(n18084) );
  NOR2X0 U18916 ( .IN1(n18104), .IN2(n18089), .QN(n18122) );
  NAND2X0 U18917 ( .IN1(n5710), .IN2(n10971), .QN(n18089) );
  NAND2X0 U18918 ( .IN1(n18124), .IN2(n18125), .QN(n18104) );
  NOR2X0 U18919 ( .IN1(g4405), .IN2(n18126), .QN(n18125) );
  NAND2X0 U18920 ( .IN1(n10621), .IN2(n10095), .QN(n18126) );
  NOR2X0 U18921 ( .IN1(g7257), .IN2(g7243), .QN(n18124) );
  NOR2X0 U18922 ( .IN1(n11042), .IN2(n18127), .QN(g26944) );
  NOR2X0 U18923 ( .IN1(n18128), .IN2(n18129), .QN(n18127) );
  NAND2X0 U18924 ( .IN1(n18130), .IN2(n11896), .QN(n18129) );
  INVX0 U18925 ( .INP(n17643), .ZN(n11896) );
  NAND2X0 U18926 ( .IN1(n18131), .IN2(n18132), .QN(n17643) );
  INVX0 U18927 ( .INP(g135), .ZN(n18132) );
  NAND2X0 U18928 ( .IN1(n18133), .IN2(n18134), .QN(n18131) );
  NAND2X0 U18929 ( .IN1(n18135), .IN2(n18136), .QN(n18134) );
  XOR2X1 U18930 ( .IN1(g4608), .IN2(n5539), .Q(n18136) );
  NOR2X0 U18931 ( .IN1(g4616), .IN2(n18137), .QN(n18135) );
  XOR2X1 U18932 ( .IN1(n5365), .IN2(n5303), .Q(n18137) );
  NOR2X0 U18933 ( .IN1(n18138), .IN2(n18139), .QN(n18133) );
  NOR2X0 U18934 ( .IN1(g4584), .IN2(n18140), .QN(n18139) );
  NAND2X0 U18935 ( .IN1(n5303), .IN2(g4608), .QN(n18140) );
  NOR2X0 U18936 ( .IN1(n5539), .IN2(n18141), .QN(n18138) );
  NAND2X0 U18937 ( .IN1(n18142), .IN2(n5274), .QN(n18141) );
  NOR2X0 U18938 ( .IN1(n5303), .IN2(g4601), .QN(n18142) );
  NOR2X0 U18939 ( .IN1(n12580), .IN2(n10643), .QN(n18130) );
  NAND2X0 U18940 ( .IN1(n18143), .IN2(g4358), .QN(n18128) );
  NAND2X0 U18941 ( .IN1(n18144), .IN2(n18145), .QN(g26940) );
  NAND2X0 U18942 ( .IN1(n11065), .IN2(g4153), .QN(n18145) );
  NAND2X0 U18943 ( .IN1(n15656), .IN2(n10972), .QN(n18144) );
  NAND2X0 U18944 ( .IN1(n18146), .IN2(n18147), .QN(n15656) );
  NAND2X0 U18945 ( .IN1(g116), .IN2(g4157), .QN(n18147) );
  NAND2X0 U18946 ( .IN1(g114), .IN2(n5983), .QN(n18146) );
  NAND2X0 U18947 ( .IN1(n18148), .IN2(n18149), .QN(g26939) );
  NAND2X0 U18948 ( .IN1(n11065), .IN2(g4104), .QN(n18149) );
  NAND2X0 U18949 ( .IN1(n15654), .IN2(n10972), .QN(n18148) );
  NAND2X0 U18950 ( .IN1(n18150), .IN2(n18151), .QN(n15654) );
  NAND2X0 U18951 ( .IN1(g124), .IN2(g4146), .QN(n18151) );
  NAND2X0 U18952 ( .IN1(g120), .IN2(n5981), .QN(n18150) );
  NAND2X0 U18953 ( .IN1(n18152), .IN2(n14906), .QN(g26938) );
  NOR2X0 U18954 ( .IN1(n18153), .IN2(n18154), .QN(n18152) );
  NOR2X0 U18955 ( .IN1(n11042), .IN2(n18155), .QN(n18154) );
  XNOR2X1 U18956 ( .IN1(g4082), .IN2(n17681), .Q(n18155) );
  NOR2X0 U18957 ( .IN1(n1269), .IN2(n5612), .QN(n17681) );
  NOR2X0 U18958 ( .IN1(n5612), .IN2(n10898), .QN(n18153) );
  NAND2X0 U18959 ( .IN1(n18156), .IN2(n18157), .QN(g26934) );
  NAND2X0 U18960 ( .IN1(n4888), .IN2(g2827), .QN(n18157) );
  NOR2X0 U18961 ( .IN1(n18158), .IN2(n18159), .QN(n18156) );
  NOR2X0 U18962 ( .IN1(n10902), .IN2(n10666), .QN(n18159) );
  NOR2X0 U18963 ( .IN1(test_so34), .IN2(n18160), .QN(n18158) );
  NAND2X0 U18964 ( .IN1(n18161), .IN2(n18162), .QN(g26933) );
  NAND2X0 U18965 ( .IN1(n4888), .IN2(test_so37), .QN(n18162) );
  NOR2X0 U18966 ( .IN1(n18163), .IN2(n18164), .QN(n18161) );
  NOR2X0 U18967 ( .IN1(n10121), .IN2(n10899), .QN(n18164) );
  NOR2X0 U18968 ( .IN1(n18160), .IN2(g2461), .QN(n18163) );
  NAND2X0 U18969 ( .IN1(n18165), .IN2(n18166), .QN(g26932) );
  NAND2X0 U18970 ( .IN1(n4888), .IN2(g2811), .QN(n18166) );
  NOR2X0 U18971 ( .IN1(n18167), .IN2(n18168), .QN(n18165) );
  NOR2X0 U18972 ( .IN1(n10118), .IN2(n10899), .QN(n18168) );
  NOR2X0 U18973 ( .IN1(n18160), .IN2(g2327), .QN(n18167) );
  NAND2X0 U18974 ( .IN1(n18169), .IN2(n18170), .QN(g26931) );
  NAND2X0 U18975 ( .IN1(n4888), .IN2(g2799), .QN(n18170) );
  NOR2X0 U18976 ( .IN1(n18171), .IN2(n18172), .QN(n18169) );
  NOR2X0 U18977 ( .IN1(n10101), .IN2(n10901), .QN(n18172) );
  NOR2X0 U18978 ( .IN1(n18160), .IN2(g2193), .QN(n18171) );
  NAND2X0 U18979 ( .IN1(n18173), .IN2(n18174), .QN(g26930) );
  NAND2X0 U18980 ( .IN1(n4888), .IN2(g2795), .QN(n18174) );
  NOR2X0 U18981 ( .IN1(n18175), .IN2(n18176), .QN(n18173) );
  NOR2X0 U18982 ( .IN1(n10120), .IN2(n10899), .QN(n18176) );
  NOR2X0 U18983 ( .IN1(test_so59), .IN2(n18160), .QN(n18175) );
  NAND2X0 U18984 ( .IN1(n18177), .IN2(n18178), .QN(g26929) );
  NAND2X0 U18985 ( .IN1(n4888), .IN2(g2791), .QN(n18178) );
  NOR2X0 U18986 ( .IN1(n18179), .IN2(n18180), .QN(n18177) );
  NOR2X0 U18987 ( .IN1(n10117), .IN2(n10900), .QN(n18180) );
  NOR2X0 U18988 ( .IN1(n18160), .IN2(g1902), .QN(n18179) );
  NAND2X0 U18989 ( .IN1(n18181), .IN2(n18182), .QN(g26928) );
  NAND2X0 U18990 ( .IN1(n4888), .IN2(g2779), .QN(n18182) );
  NOR2X0 U18991 ( .IN1(n18183), .IN2(n18184), .QN(n18181) );
  NOR2X0 U18992 ( .IN1(n10123), .IN2(n10900), .QN(n18184) );
  NOR2X0 U18993 ( .IN1(n18160), .IN2(g1768), .QN(n18183) );
  NAND2X0 U18994 ( .IN1(n18185), .IN2(n18186), .QN(g26927) );
  NAND2X0 U18995 ( .IN1(n4888), .IN2(g2767), .QN(n18186) );
  NOR2X0 U18996 ( .IN1(n18187), .IN2(n18188), .QN(n18185) );
  NOR2X0 U18997 ( .IN1(n10100), .IN2(n10900), .QN(n18188) );
  NOR2X0 U18998 ( .IN1(n18160), .IN2(g1632), .QN(n18187) );
  NAND2X0 U18999 ( .IN1(n18189), .IN2(n4888), .QN(n18160) );
  NOR2X0 U19000 ( .IN1(n12372), .IN2(n18190), .QN(n18189) );
  NOR2X0 U19001 ( .IN1(test_so30), .IN2(g2748), .QN(n18190) );
  NOR2X0 U19002 ( .IN1(n18191), .IN2(n5300), .QN(n12372) );
  NAND2X0 U19003 ( .IN1(g2735), .IN2(n3505), .QN(n18191) );
  NOR2X0 U19004 ( .IN1(n5349), .IN2(n5516), .QN(n3505) );
  NAND2X0 U19005 ( .IN1(n18192), .IN2(n18193), .QN(g26926) );
  NAND2X0 U19006 ( .IN1(n18194), .IN2(n3730), .QN(n18193) );
  XOR2X1 U19007 ( .IN1(g2724), .IN2(n16065), .Q(n18194) );
  NOR2X0 U19008 ( .IN1(n5299), .IN2(n5465), .QN(n16065) );
  NAND2X0 U19009 ( .IN1(n11065), .IN2(g2719), .QN(n18192) );
  NAND2X0 U19010 ( .IN1(n18195), .IN2(n18196), .QN(g26925) );
  NAND2X0 U19011 ( .IN1(n11065), .IN2(g1532), .QN(n18196) );
  NAND2X0 U19012 ( .IN1(n18197), .IN2(n10972), .QN(n18195) );
  NAND2X0 U19013 ( .IN1(n16413), .IN2(n18198), .QN(n18197) );
  NAND2X0 U19014 ( .IN1(n18199), .IN2(g1536), .QN(n18198) );
  INVX0 U19015 ( .INP(n16392), .ZN(n18199) );
  NOR2X0 U19016 ( .IN1(n16403), .IN2(n10090), .QN(n16392) );
  INVX0 U19017 ( .INP(n16394), .ZN(n16403) );
  NOR2X0 U19018 ( .IN1(n16404), .IN2(n10584), .QN(n16394) );
  NAND2X0 U19019 ( .IN1(n18200), .IN2(n16414), .QN(n16404) );
  NOR2X0 U19020 ( .IN1(n5302), .IN2(n18201), .QN(n18200) );
  NOR2X0 U19021 ( .IN1(g1532), .IN2(n18202), .QN(n18201) );
  NAND2X0 U19022 ( .IN1(g1339), .IN2(g1521), .QN(n18202) );
  INVX0 U19023 ( .INP(n4173), .ZN(n16413) );
  NAND2X0 U19024 ( .IN1(n18203), .IN2(n18204), .QN(g26924) );
  NAND2X0 U19025 ( .IN1(n18205), .IN2(n5289), .QN(n18204) );
  INVX0 U19026 ( .INP(n18206), .ZN(n18205) );
  NOR2X0 U19027 ( .IN1(n18207), .IN2(n18208), .QN(n18203) );
  NOR2X0 U19028 ( .IN1(n5696), .IN2(n10901), .QN(n18208) );
  NOR2X0 U19029 ( .IN1(n11026), .IN2(n18209), .QN(n18207) );
  NAND2X0 U19030 ( .IN1(n18206), .IN2(g1478), .QN(n18209) );
  NAND2X0 U19031 ( .IN1(n18210), .IN2(n18211), .QN(n18206) );
  NOR2X0 U19032 ( .IN1(n5696), .IN2(n17050), .QN(n18210) );
  NAND2X0 U19033 ( .IN1(n18212), .IN2(g13272), .QN(n17050) );
  NOR2X0 U19034 ( .IN1(test_so49), .IN2(n5364), .QN(n18212) );
  NAND2X0 U19035 ( .IN1(n18213), .IN2(n18214), .QN(g26923) );
  NAND2X0 U19036 ( .IN1(n18215), .IN2(n5290), .QN(n18214) );
  NOR2X0 U19037 ( .IN1(n18216), .IN2(n18217), .QN(n18213) );
  NOR2X0 U19038 ( .IN1(n5693), .IN2(n10901), .QN(n18217) );
  NOR2X0 U19039 ( .IN1(n11025), .IN2(n18218), .QN(n18216) );
  INVX0 U19040 ( .INP(n18219), .ZN(n18218) );
  NOR2X0 U19041 ( .IN1(n18215), .IN2(n5290), .QN(n18219) );
  NOR2X0 U19042 ( .IN1(n18220), .IN2(n18221), .QN(n18215) );
  NAND2X0 U19043 ( .IN1(g1467), .IN2(g13272), .QN(n18221) );
  NAND2X0 U19044 ( .IN1(n13753), .IN2(n18211), .QN(n18220) );
  NAND2X0 U19045 ( .IN1(n18222), .IN2(n18223), .QN(g26922) );
  NAND2X0 U19046 ( .IN1(n18224), .IN2(n5343), .QN(n18223) );
  INVX0 U19047 ( .INP(n18225), .ZN(n18224) );
  NOR2X0 U19048 ( .IN1(n18226), .IN2(n18227), .QN(n18222) );
  NOR2X0 U19049 ( .IN1(n5866), .IN2(n10899), .QN(n18227) );
  NOR2X0 U19050 ( .IN1(n11026), .IN2(n18228), .QN(n18226) );
  NAND2X0 U19051 ( .IN1(n18225), .IN2(g1448), .QN(n18228) );
  NAND2X0 U19052 ( .IN1(n18229), .IN2(n18211), .QN(n18225) );
  NOR2X0 U19053 ( .IN1(n5866), .IN2(n17013), .QN(n18229) );
  NAND2X0 U19054 ( .IN1(n16414), .IN2(g13272), .QN(n17013) );
  INVX0 U19055 ( .INP(n13811), .ZN(n16414) );
  NAND2X0 U19056 ( .IN1(n5364), .IN2(test_so49), .QN(n13811) );
  NAND2X0 U19057 ( .IN1(n18230), .IN2(n18231), .QN(g26921) );
  NAND2X0 U19058 ( .IN1(n11065), .IN2(g1395), .QN(n18231) );
  NAND2X0 U19059 ( .IN1(n18232), .IN2(n10972), .QN(n18230) );
  NOR2X0 U19060 ( .IN1(test_so68), .IN2(n18233), .QN(n18232) );
  XNOR2X1 U19061 ( .IN1(n10251), .IN2(n18234), .Q(n18233) );
  NAND2X0 U19062 ( .IN1(n18235), .IN2(n18236), .QN(g26920) );
  NAND2X0 U19063 ( .IN1(n11065), .IN2(g1384), .QN(n18236) );
  NAND2X0 U19064 ( .IN1(n18237), .IN2(n10972), .QN(n18235) );
  NAND2X0 U19065 ( .IN1(n18238), .IN2(n18239), .QN(n18237) );
  INVX0 U19066 ( .INP(n18240), .ZN(n18239) );
  NOR2X0 U19067 ( .IN1(n4915), .IN2(n10620), .QN(n18240) );
  NOR2X0 U19068 ( .IN1(n18241), .IN2(n18242), .QN(n4915) );
  NOR2X0 U19069 ( .IN1(g1384), .IN2(n5322), .QN(n18242) );
  NAND2X0 U19070 ( .IN1(n4913), .IN2(g1351), .QN(n18238) );
  NAND2X0 U19071 ( .IN1(n18243), .IN2(n18244), .QN(g26919) );
  NAND2X0 U19072 ( .IN1(n11065), .IN2(g1266), .QN(n18244) );
  NOR2X0 U19073 ( .IN1(n18245), .IN2(n18246), .QN(n18243) );
  NOR2X0 U19074 ( .IN1(test_so77), .IN2(n18247), .QN(n18246) );
  NOR2X0 U19075 ( .IN1(n1249), .IN2(n18248), .QN(n18245) );
  NAND2X0 U19076 ( .IN1(test_so77), .IN2(n14133), .QN(n18248) );
  INVX0 U19077 ( .INP(n18247), .ZN(n1249) );
  NAND2X0 U19078 ( .IN1(n18249), .IN2(g1249), .QN(n18247) );
  NOR2X0 U19079 ( .IN1(n5655), .IN2(n10242), .QN(n18249) );
  NAND2X0 U19080 ( .IN1(n18250), .IN2(n18251), .QN(g26918) );
  NAND2X0 U19081 ( .IN1(n11064), .IN2(g1189), .QN(n18251) );
  INVX0 U19082 ( .INP(n18252), .ZN(n18250) );
  NOR2X0 U19083 ( .IN1(n18253), .IN2(n11023), .QN(n18252) );
  NOR2X0 U19084 ( .IN1(n4191), .IN2(n18254), .QN(n18253) );
  NOR2X0 U19085 ( .IN1(n16435), .IN2(n10606), .QN(n18254) );
  NOR2X0 U19086 ( .IN1(n16447), .IN2(n10089), .QN(n16435) );
  INVX0 U19087 ( .INP(n16437), .ZN(n16447) );
  NOR2X0 U19088 ( .IN1(n16448), .IN2(n10583), .QN(n16437) );
  NAND2X0 U19089 ( .IN1(n18255), .IN2(n14051), .QN(n16448) );
  NOR2X0 U19090 ( .IN1(n5304), .IN2(n18256), .QN(n18255) );
  NOR2X0 U19091 ( .IN1(g1189), .IN2(n18257), .QN(n18256) );
  NAND2X0 U19092 ( .IN1(g1178), .IN2(g996), .QN(n18257) );
  NAND2X0 U19093 ( .IN1(n18258), .IN2(n18259), .QN(g26917) );
  NAND2X0 U19094 ( .IN1(n18260), .IN2(n5328), .QN(n18259) );
  INVX0 U19095 ( .INP(n18261), .ZN(n18260) );
  NOR2X0 U19096 ( .IN1(n18262), .IN2(n18263), .QN(n18258) );
  NOR2X0 U19097 ( .IN1(n5697), .IN2(n10900), .QN(n18263) );
  NOR2X0 U19098 ( .IN1(n11028), .IN2(n18264), .QN(n18262) );
  NAND2X0 U19099 ( .IN1(n18261), .IN2(g1135), .QN(n18264) );
  NAND2X0 U19100 ( .IN1(n18265), .IN2(n18266), .QN(n18261) );
  NOR2X0 U19101 ( .IN1(n5697), .IN2(g1183), .QN(n18266) );
  NAND2X0 U19102 ( .IN1(n18267), .IN2(n18268), .QN(g26916) );
  NAND2X0 U19103 ( .IN1(n18269), .IN2(n5329), .QN(n18268) );
  INVX0 U19104 ( .INP(n18270), .ZN(n18269) );
  NOR2X0 U19105 ( .IN1(n18271), .IN2(n18272), .QN(n18267) );
  NOR2X0 U19106 ( .IN1(n5692), .IN2(n10893), .QN(n18272) );
  NOR2X0 U19107 ( .IN1(n11028), .IN2(n18273), .QN(n18271) );
  NAND2X0 U19108 ( .IN1(n18270), .IN2(g1129), .QN(n18273) );
  NAND2X0 U19109 ( .IN1(n18265), .IN2(n18274), .QN(n18270) );
  NOR2X0 U19110 ( .IN1(n5692), .IN2(n5599), .QN(n18274) );
  NOR2X0 U19111 ( .IN1(n17086), .IN2(n18275), .QN(n18265) );
  NAND2X0 U19112 ( .IN1(g1171), .IN2(g13259), .QN(n17086) );
  NAND2X0 U19113 ( .IN1(n18276), .IN2(n18277), .QN(g26915) );
  NAND2X0 U19114 ( .IN1(n18278), .IN2(n5478), .QN(n18277) );
  INVX0 U19115 ( .INP(n18279), .ZN(n18278) );
  NOR2X0 U19116 ( .IN1(n18280), .IN2(n18281), .QN(n18276) );
  NOR2X0 U19117 ( .IN1(n10907), .IN2(n10665), .QN(n18281) );
  NOR2X0 U19118 ( .IN1(n11028), .IN2(n18282), .QN(n18280) );
  NAND2X0 U19119 ( .IN1(n18279), .IN2(g1105), .QN(n18282) );
  NAND2X0 U19120 ( .IN1(n18283), .IN2(n18284), .QN(n18279) );
  NOR2X0 U19121 ( .IN1(n17063), .IN2(n10665), .QN(n18283) );
  NAND2X0 U19122 ( .IN1(n14051), .IN2(g13259), .QN(n17063) );
  INVX0 U19123 ( .INP(n16452), .ZN(n14051) );
  NAND2X0 U19124 ( .IN1(n5363), .IN2(g1183), .QN(n16452) );
  NAND2X0 U19125 ( .IN1(n18285), .IN2(n18286), .QN(g26914) );
  NAND2X0 U19126 ( .IN1(n11064), .IN2(g1052), .QN(n18286) );
  NAND2X0 U19127 ( .IN1(n18287), .IN2(n10972), .QN(n18285) );
  NOR2X0 U19128 ( .IN1(n18288), .IN2(g979), .QN(n18287) );
  XNOR2X1 U19129 ( .IN1(n10252), .IN2(n18289), .Q(n18288) );
  NAND2X0 U19130 ( .IN1(n18290), .IN2(n18291), .QN(g26913) );
  NAND2X0 U19131 ( .IN1(n4938), .IN2(n18292), .QN(n18291) );
  NOR2X0 U19132 ( .IN1(n18293), .IN2(n18294), .QN(n18290) );
  NOR2X0 U19133 ( .IN1(n11028), .IN2(n18295), .QN(n18294) );
  INVX0 U19134 ( .INP(n18296), .ZN(n18295) );
  NOR2X0 U19135 ( .IN1(n4940), .IN2(n10619), .QN(n18296) );
  NOR2X0 U19136 ( .IN1(n18297), .IN2(n18298), .QN(n4940) );
  NOR2X0 U19137 ( .IN1(g1041), .IN2(n5321), .QN(n18298) );
  NOR2X0 U19138 ( .IN1(n10104), .IN2(n10893), .QN(n18293) );
  NAND2X0 U19139 ( .IN1(n18299), .IN2(n18300), .QN(g26912) );
  NAND2X0 U19140 ( .IN1(n11063), .IN2(g921), .QN(n18300) );
  NOR2X0 U19141 ( .IN1(n18301), .IN2(n18302), .QN(n18299) );
  NOR2X0 U19142 ( .IN1(g936), .IN2(n11434), .QN(n18302) );
  NOR2X0 U19143 ( .IN1(n5557), .IN2(n18303), .QN(n18301) );
  NAND2X0 U19144 ( .IN1(n14152), .IN2(n11434), .QN(n18303) );
  NAND2X0 U19145 ( .IN1(n18304), .IN2(g921), .QN(n11434) );
  NOR2X0 U19146 ( .IN1(n5654), .IN2(n10240), .QN(n18304) );
  XOR2X1 U19147 ( .IN1(n18305), .IN2(n5682), .Q(g26910) );
  NAND2X0 U19148 ( .IN1(n5305), .IN2(n10972), .QN(n18305) );
  NAND2X0 U19149 ( .IN1(n18306), .IN2(n18307), .QN(g26909) );
  NAND2X0 U19150 ( .IN1(n11063), .IN2(g890), .QN(n18307) );
  NAND2X0 U19151 ( .IN1(n18308), .IN2(n10973), .QN(n18306) );
  NAND2X0 U19152 ( .IN1(n18309), .IN2(n18310), .QN(n18308) );
  NAND2X0 U19153 ( .IN1(n5431), .IN2(g862), .QN(n18310) );
  NAND2X0 U19154 ( .IN1(n5305), .IN2(g896), .QN(n18309) );
  NAND2X0 U19155 ( .IN1(n18311), .IN2(n18312), .QN(g26908) );
  NAND2X0 U19156 ( .IN1(n4945), .IN2(g446), .QN(n18312) );
  NOR2X0 U19157 ( .IN1(n18313), .IN2(n18314), .QN(n18311) );
  NOR2X0 U19158 ( .IN1(n6008), .IN2(n10892), .QN(n18314) );
  NOR2X0 U19159 ( .IN1(n10111), .IN2(n18315), .QN(n18313) );
  NAND2X0 U19160 ( .IN1(n18316), .IN2(n18317), .QN(g26907) );
  NAND2X0 U19161 ( .IN1(n4945), .IN2(g246), .QN(n18317) );
  NOR2X0 U19162 ( .IN1(n18318), .IN2(n18319), .QN(n18316) );
  NOR2X0 U19163 ( .IN1(n10277), .IN2(n10892), .QN(n18319) );
  NOR2X0 U19164 ( .IN1(n10113), .IN2(n18315), .QN(n18318) );
  NAND2X0 U19165 ( .IN1(n18320), .IN2(n18321), .QN(g26906) );
  NAND2X0 U19166 ( .IN1(n4945), .IN2(g269), .QN(n18321) );
  NOR2X0 U19167 ( .IN1(n18322), .IN2(n18323), .QN(n18320) );
  NOR2X0 U19168 ( .IN1(n10400), .IN2(n10892), .QN(n18323) );
  NOR2X0 U19169 ( .IN1(n10110), .IN2(n18315), .QN(n18322) );
  NAND2X0 U19170 ( .IN1(n18324), .IN2(n18325), .QN(g26905) );
  NAND2X0 U19171 ( .IN1(n4945), .IN2(g239), .QN(n18325) );
  NOR2X0 U19172 ( .IN1(n18326), .IN2(n18327), .QN(n18324) );
  NOR2X0 U19173 ( .IN1(n10276), .IN2(n10891), .QN(n18327) );
  NOR2X0 U19174 ( .IN1(n10109), .IN2(n18315), .QN(n18326) );
  NAND2X0 U19175 ( .IN1(n18328), .IN2(n18329), .QN(g26904) );
  NAND2X0 U19176 ( .IN1(n4945), .IN2(g262), .QN(n18329) );
  NOR2X0 U19177 ( .IN1(n18330), .IN2(n18331), .QN(n18328) );
  NOR2X0 U19178 ( .IN1(n10399), .IN2(n10891), .QN(n18331) );
  NOR2X0 U19179 ( .IN1(n10107), .IN2(n18315), .QN(n18330) );
  NAND2X0 U19180 ( .IN1(n18332), .IN2(n18333), .QN(g26903) );
  NAND2X0 U19181 ( .IN1(n4945), .IN2(g232), .QN(n18333) );
  NOR2X0 U19182 ( .IN1(n18334), .IN2(n18335), .QN(n18332) );
  NOR2X0 U19183 ( .IN1(n10275), .IN2(n10891), .QN(n18335) );
  NOR2X0 U19184 ( .IN1(n10108), .IN2(n18315), .QN(n18334) );
  NAND2X0 U19185 ( .IN1(n18336), .IN2(n18337), .QN(g26902) );
  NAND2X0 U19186 ( .IN1(n4945), .IN2(g255), .QN(n18337) );
  NOR2X0 U19187 ( .IN1(n18338), .IN2(n18339), .QN(n18336) );
  NOR2X0 U19188 ( .IN1(n5597), .IN2(n10891), .QN(n18339) );
  NOR2X0 U19189 ( .IN1(n10106), .IN2(n18315), .QN(n18338) );
  NAND2X0 U19190 ( .IN1(n18340), .IN2(n18341), .QN(g26901) );
  NAND2X0 U19191 ( .IN1(n4945), .IN2(g225), .QN(n18341) );
  NOR2X0 U19192 ( .IN1(n18342), .IN2(n18343), .QN(n18340) );
  NOR2X0 U19193 ( .IN1(n10111), .IN2(n10891), .QN(n18343) );
  NOR2X0 U19194 ( .IN1(n10112), .IN2(n18315), .QN(n18342) );
  NAND2X0 U19195 ( .IN1(n10928), .IN2(n18344), .QN(n18315) );
  INVX0 U19196 ( .INP(n4946), .ZN(n18344) );
  NAND2X0 U19197 ( .IN1(n18345), .IN2(n5682), .QN(n4946) );
  NOR2X0 U19198 ( .IN1(n5305), .IN2(g896), .QN(n18345) );
  NAND2X0 U19199 ( .IN1(n18346), .IN2(n18347), .QN(g26899) );
  NAND2X0 U19200 ( .IN1(n18348), .IN2(n4518), .QN(n18347) );
  XOR2X1 U19201 ( .IN1(n4814), .IN2(g822), .Q(n18348) );
  NOR2X0 U19202 ( .IN1(n18349), .IN2(n17177), .QN(n4814) );
  NAND2X0 U19203 ( .IN1(g817), .IN2(g832), .QN(n18349) );
  NAND2X0 U19204 ( .IN1(n11063), .IN2(g832), .QN(n18346) );
  NAND2X0 U19205 ( .IN1(n18350), .IN2(n18351), .QN(g26898) );
  NAND2X0 U19206 ( .IN1(n18352), .IN2(n18353), .QN(n18351) );
  NAND2X0 U19207 ( .IN1(n18354), .IN2(n18355), .QN(n18353) );
  NAND2X0 U19208 ( .IN1(n10216), .IN2(n10973), .QN(n18355) );
  NAND2X0 U19209 ( .IN1(n18356), .IN2(g843), .QN(n18350) );
  NAND2X0 U19210 ( .IN1(n18357), .IN2(n10973), .QN(n18356) );
  NAND2X0 U19211 ( .IN1(n18358), .IN2(n18359), .QN(n18357) );
  NOR2X0 U19212 ( .IN1(n5562), .IN2(g812), .QN(n18358) );
  NAND2X0 U19213 ( .IN1(n18360), .IN2(n18361), .QN(g26897) );
  NAND2X0 U19214 ( .IN1(n18362), .IN2(g753), .QN(n18361) );
  NAND2X0 U19215 ( .IN1(n18363), .IN2(g732), .QN(n18360) );
  INVX0 U19216 ( .INP(n18362), .ZN(n18363) );
  NOR2X0 U19217 ( .IN1(n18364), .IN2(n11018), .QN(n18362) );
  NAND2X0 U19218 ( .IN1(n18365), .IN2(n18366), .QN(g26896) );
  NAND2X0 U19219 ( .IN1(n4956), .IN2(n18367), .QN(n18366) );
  INVX0 U19220 ( .INP(n154), .ZN(n18367) );
  NOR2X0 U19221 ( .IN1(n18368), .IN2(n18369), .QN(n18365) );
  NOR2X0 U19222 ( .IN1(n10283), .IN2(n18370), .QN(n18369) );
  INVX0 U19223 ( .INP(n18371), .ZN(n18370) );
  NOR2X0 U19224 ( .IN1(n5657), .IN2(n18371), .QN(n18368) );
  NAND2X0 U19225 ( .IN1(n154), .IN2(n10973), .QN(n18371) );
  NAND2X0 U19226 ( .IN1(n18372), .IN2(n18373), .QN(n154) );
  NOR2X0 U19227 ( .IN1(n17177), .IN2(n18002), .QN(n18373) );
  NOR2X0 U19228 ( .IN1(g504), .IN2(n10649), .QN(n18372) );
  NAND2X0 U19229 ( .IN1(n18374), .IN2(n18375), .QN(g26895) );
  NAND2X0 U19230 ( .IN1(n11063), .IN2(g562), .QN(n18375) );
  NOR2X0 U19231 ( .IN1(n18376), .IN2(n18377), .QN(n18374) );
  NOR2X0 U19232 ( .IN1(g568), .IN2(n11294), .QN(n18377) );
  NOR2X0 U19233 ( .IN1(n5335), .IN2(n18378), .QN(n18376) );
  NAND2X0 U19234 ( .IN1(n2421), .IN2(n11294), .QN(n18378) );
  NAND2X0 U19235 ( .IN1(n18379), .IN2(n4959), .QN(n11294) );
  NOR2X0 U19236 ( .IN1(n10098), .IN2(n18380), .QN(n18379) );
  NAND2X0 U19237 ( .IN1(n18381), .IN2(n18382), .QN(g26894) );
  NAND2X0 U19238 ( .IN1(n18383), .IN2(n17997), .QN(n18382) );
  NOR2X0 U19239 ( .IN1(n18384), .IN2(n18385), .QN(n18383) );
  NOR2X0 U19240 ( .IN1(n5327), .IN2(n18386), .QN(n18385) );
  NAND2X0 U19241 ( .IN1(n18387), .IN2(n17973), .QN(n18386) );
  INVX0 U19242 ( .INP(n18388), .ZN(n18387) );
  NOR2X0 U19243 ( .IN1(n18001), .IN2(n11015), .QN(n18388) );
  NOR2X0 U19244 ( .IN1(n18389), .IN2(g528), .QN(n18384) );
  NOR2X0 U19245 ( .IN1(n17999), .IN2(n18390), .QN(n18389) );
  NAND2X0 U19246 ( .IN1(n18001), .IN2(n18002), .QN(n18390) );
  NAND2X0 U19247 ( .IN1(n18391), .IN2(n5327), .QN(n18002) );
  NOR2X0 U19248 ( .IN1(n5820), .IN2(n5708), .QN(n18391) );
  NAND2X0 U19249 ( .IN1(n11063), .IN2(g518), .QN(n18381) );
  NAND2X0 U19250 ( .IN1(n18392), .IN2(n18393), .QN(g26893) );
  NAND2X0 U19251 ( .IN1(n11062), .IN2(g355), .QN(n18393) );
  NAND2X0 U19252 ( .IN1(n18394), .IN2(n10973), .QN(n18392) );
  NAND2X0 U19253 ( .IN1(n18395), .IN2(n18396), .QN(n18394) );
  NAND2X0 U19254 ( .IN1(g29211), .IN2(n10674), .QN(n18396) );
  NAND2X0 U19255 ( .IN1(test_so17), .IN2(n18397), .QN(n18395) );
  INVX0 U19256 ( .INP(n18398), .ZN(n18397) );
  NAND2X0 U19257 ( .IN1(n18399), .IN2(n18400), .QN(g26892) );
  NAND2X0 U19258 ( .IN1(n18401), .IN2(n10674), .QN(n18400) );
  NOR2X0 U19259 ( .IN1(n18398), .IN2(n11015), .QN(n18401) );
  NOR2X0 U19260 ( .IN1(g355), .IN2(g333), .QN(n18398) );
  NAND2X0 U19261 ( .IN1(test_so17), .IN2(n11081), .QN(n18399) );
  NAND2X0 U19262 ( .IN1(n18402), .IN2(n18403), .QN(g26891) );
  NAND2X0 U19263 ( .IN1(n11062), .IN2(g347), .QN(n18403) );
  NAND2X0 U19264 ( .IN1(n18404), .IN2(n5860), .QN(n18402) );
  NOR2X0 U19265 ( .IN1(n10126), .IN2(n11016), .QN(n18404) );
  NAND2X0 U19266 ( .IN1(n18405), .IN2(n18406), .QN(g26890) );
  NAND2X0 U19267 ( .IN1(n5860), .IN2(n10973), .QN(n18406) );
  NAND2X0 U19268 ( .IN1(n11062), .IN2(g333), .QN(n18405) );
  NAND2X0 U19269 ( .IN1(n18407), .IN2(n18408), .QN(g26889) );
  NAND2X0 U19270 ( .IN1(n11062), .IN2(g29211), .QN(n18408) );
  NAND2X0 U19271 ( .IN1(n18409), .IN2(n10973), .QN(n18407) );
  NOR2X0 U19272 ( .IN1(n9306), .IN2(n18410), .QN(n18409) );
  NAND2X0 U19273 ( .IN1(n18411), .IN2(g329), .QN(n18410) );
  NAND2X0 U19274 ( .IN1(n18412), .IN2(n18413), .QN(g26888) );
  NAND2X0 U19275 ( .IN1(n10928), .IN2(g316), .QN(n18413) );
  NAND2X0 U19276 ( .IN1(n11060), .IN2(g29216), .QN(n18412) );
  NAND2X0 U19277 ( .IN1(n18414), .IN2(n18415), .QN(g26887) );
  NOR2X0 U19278 ( .IN1(n18416), .IN2(n18417), .QN(n18414) );
  NOR2X0 U19279 ( .IN1(n11030), .IN2(n18418), .QN(n18417) );
  NAND2X0 U19280 ( .IN1(n5317), .IN2(g324), .QN(n18418) );
  NOR2X0 U19281 ( .IN1(n5824), .IN2(n10889), .QN(n18416) );
  NAND2X0 U19282 ( .IN1(n18419), .IN2(n18420), .QN(g26886) );
  NAND2X0 U19283 ( .IN1(n18421), .IN2(n18422), .QN(n18420) );
  INVX0 U19284 ( .INP(n18415), .ZN(n18421) );
  NOR2X0 U19285 ( .IN1(n18423), .IN2(n18424), .QN(n18419) );
  NOR2X0 U19286 ( .IN1(n5317), .IN2(n10889), .QN(n18424) );
  NOR2X0 U19287 ( .IN1(n11030), .IN2(n18425), .QN(n18423) );
  NAND2X0 U19288 ( .IN1(n18411), .IN2(g336), .QN(n18425) );
  NAND2X0 U19289 ( .IN1(n18426), .IN2(n18427), .QN(g26884) );
  NAND2X0 U19290 ( .IN1(n11060), .IN2(g329), .QN(n18427) );
  NAND2X0 U19291 ( .IN1(n18428), .IN2(n10974), .QN(n18426) );
  NAND2X0 U19292 ( .IN1(n18429), .IN2(n18430), .QN(n18428) );
  INVX0 U19293 ( .INP(n18431), .ZN(n18430) );
  NOR2X0 U19294 ( .IN1(n18432), .IN2(n18433), .QN(n18431) );
  NAND2X0 U19295 ( .IN1(n5317), .IN2(n5282), .QN(n18433) );
  NAND2X0 U19296 ( .IN1(n5456), .IN2(n5766), .QN(n18432) );
  NAND2X0 U19297 ( .IN1(n18422), .IN2(n18434), .QN(n18429) );
  NAND2X0 U19298 ( .IN1(n18435), .IN2(n5456), .QN(n18434) );
  NOR2X0 U19299 ( .IN1(n18436), .IN2(n18437), .QN(n18435) );
  NOR2X0 U19300 ( .IN1(n5824), .IN2(n5282), .QN(n18437) );
  NOR2X0 U19301 ( .IN1(n5317), .IN2(g336), .QN(n18436) );
  NAND2X0 U19302 ( .IN1(n18438), .IN2(n18439), .QN(g26883) );
  NAND2X0 U19303 ( .IN1(n11059), .IN2(g324), .QN(n18439) );
  NAND2X0 U19304 ( .IN1(n18422), .IN2(n10975), .QN(n18438) );
  INVX0 U19305 ( .INP(n18411), .ZN(n18422) );
  NAND2X0 U19306 ( .IN1(n18440), .IN2(n18441), .QN(n18411) );
  NAND2X0 U19307 ( .IN1(n5282), .IN2(g324), .QN(n18441) );
  NAND2X0 U19308 ( .IN1(n5827), .IN2(n5317), .QN(n18440) );
  NAND2X0 U19309 ( .IN1(n18442), .IN2(n18415), .QN(g26882) );
  NAND2X0 U19310 ( .IN1(n10933), .IN2(g305), .QN(n18415) );
  NOR2X0 U19311 ( .IN1(n18443), .IN2(n18444), .QN(n18442) );
  NOR2X0 U19312 ( .IN1(n10169), .IN2(n10888), .QN(n18444) );
  NOR2X0 U19313 ( .IN1(n5317), .IN2(n11019), .QN(n18443) );
  NAND2X0 U19314 ( .IN1(n18445), .IN2(n18446), .QN(g26881) );
  NAND2X0 U19315 ( .IN1(g6744), .IN2(n10937), .QN(n18446) );
  NAND2X0 U19316 ( .IN1(n11059), .IN2(g305), .QN(n18445) );
  NAND2X0 U19317 ( .IN1(n18447), .IN2(n12010), .QN(g26877) );
  NAND2X0 U19318 ( .IN1(n18448), .IN2(n18449), .QN(n12010) );
  NOR2X0 U19319 ( .IN1(n18450), .IN2(n18451), .QN(n18449) );
  NAND2X0 U19320 ( .IN1(n5311), .IN2(n5310), .QN(n18451) );
  NAND2X0 U19321 ( .IN1(n5276), .IN2(n10653), .QN(n18450) );
  NOR2X0 U19322 ( .IN1(n18452), .IN2(n18453), .QN(n18448) );
  NAND2X0 U19323 ( .IN1(n5620), .IN2(n5619), .QN(n18453) );
  NAND2X0 U19324 ( .IN1(n5406), .IN2(n5405), .QN(n18452) );
  NOR2X0 U19325 ( .IN1(n11029), .IN2(n18454), .QN(n18447) );
  INVX0 U19326 ( .INP(n12009), .ZN(n18454) );
  NAND2X0 U19327 ( .IN1(n18455), .IN2(n18456), .QN(n12009) );
  NOR2X0 U19328 ( .IN1(n18457), .IN2(n18458), .QN(n18456) );
  NAND2X0 U19329 ( .IN1(n5829), .IN2(n5828), .QN(n18458) );
  NAND2X0 U19330 ( .IN1(n5407), .IN2(n10646), .QN(n18457) );
  NOR2X0 U19331 ( .IN1(n18459), .IN2(n18460), .QN(n18455) );
  NAND2X0 U19332 ( .IN1(n5833), .IN2(n5832), .QN(n18460) );
  NAND2X0 U19333 ( .IN1(n5831), .IN2(n5830), .QN(n18459) );
  NAND2X0 U19334 ( .IN1(n18461), .IN2(n11961), .QN(g26876) );
  NAND2X0 U19335 ( .IN1(n18462), .IN2(n18463), .QN(n11961) );
  NOR2X0 U19336 ( .IN1(n18464), .IN2(n18465), .QN(n18463) );
  NAND2X0 U19337 ( .IN1(n5848), .IN2(n5847), .QN(n18465) );
  NAND2X0 U19338 ( .IN1(n5845), .IN2(n5412), .QN(n18464) );
  NOR2X0 U19339 ( .IN1(n18466), .IN2(n18467), .QN(n18462) );
  NAND2X0 U19340 ( .IN1(n19400), .IN2(n5892), .QN(n18467) );
  NAND2X0 U19341 ( .IN1(n5891), .IN2(n5890), .QN(n18466) );
  NOR2X0 U19342 ( .IN1(n11033), .IN2(n11967), .QN(n18461) );
  INVX0 U19343 ( .INP(n12033), .ZN(n11967) );
  NAND2X0 U19344 ( .IN1(n18468), .IN2(n18469), .QN(n12033) );
  NOR2X0 U19345 ( .IN1(n18470), .IN2(n18471), .QN(n18469) );
  NAND2X0 U19346 ( .IN1(n5411), .IN2(n5410), .QN(n18471) );
  NAND2X0 U19347 ( .IN1(n5278), .IN2(n10671), .QN(n18470) );
  NOR2X0 U19348 ( .IN1(n18472), .IN2(n18473), .QN(n18468) );
  NAND2X0 U19349 ( .IN1(n19401), .IN2(n19402), .QN(n18473) );
  NAND2X0 U19350 ( .IN1(n19403), .IN2(n19404), .QN(n18472) );
  NAND2X0 U19351 ( .IN1(n18474), .IN2(n12038), .QN(g26875) );
  NAND2X0 U19352 ( .IN1(n18475), .IN2(n18476), .QN(n12038) );
  NOR2X0 U19353 ( .IN1(g2523), .IN2(g2657), .QN(n18476) );
  NOR2X0 U19354 ( .IN1(g2255), .IN2(g2389), .QN(n18475) );
  NOR2X0 U19355 ( .IN1(n11057), .IN2(n12039), .QN(n18474) );
  NOR2X0 U19356 ( .IN1(n18477), .IN2(n18478), .QN(n12039) );
  NAND2X0 U19357 ( .IN1(n5280), .IN2(n5315), .QN(n18478) );
  NAND2X0 U19358 ( .IN1(n5413), .IN2(n5628), .QN(n18477) );
  NAND2X0 U19359 ( .IN1(n18479), .IN2(n18480), .QN(g25764) );
  NAND2X0 U19360 ( .IN1(n11481), .IN2(g6505), .QN(n18480) );
  NAND2X0 U19361 ( .IN1(n15009), .IN2(g6541), .QN(n18479) );
  NAND2X0 U19362 ( .IN1(n18481), .IN2(n18482), .QN(g25763) );
  NAND2X0 U19363 ( .IN1(n11481), .IN2(g6537), .QN(n18482) );
  NOR2X0 U19364 ( .IN1(n18483), .IN2(n18484), .QN(n18481) );
  NOR2X0 U19365 ( .IN1(g6533), .IN2(n18485), .QN(n18484) );
  NAND2X0 U19366 ( .IN1(n18486), .IN2(n5659), .QN(n18485) );
  NOR2X0 U19367 ( .IN1(n11057), .IN2(n13440), .QN(n18486) );
  NOR2X0 U19368 ( .IN1(n5445), .IN2(n18487), .QN(n18483) );
  NOR2X0 U19369 ( .IN1(n11058), .IN2(n18488), .QN(n18487) );
  NOR2X0 U19370 ( .IN1(n5659), .IN2(n13440), .QN(n18488) );
  NAND2X0 U19371 ( .IN1(n18489), .IN2(n18490), .QN(g25761) );
  NAND2X0 U19372 ( .IN1(n11481), .IN2(g6513), .QN(n18490) );
  INVX0 U19373 ( .INP(n15009), .ZN(n11481) );
  NAND2X0 U19374 ( .IN1(n13440), .IN2(n10939), .QN(n15009) );
  NOR2X0 U19375 ( .IN1(n18491), .IN2(n18492), .QN(n18489) );
  NOR2X0 U19376 ( .IN1(n10171), .IN2(n10888), .QN(n18492) );
  NOR2X0 U19377 ( .IN1(n11057), .IN2(n18493), .QN(n18491) );
  NAND2X0 U19378 ( .IN1(n5426), .IN2(n18494), .QN(n18493) );
  INVX0 U19379 ( .INP(n13440), .ZN(n18494) );
  NAND2X0 U19380 ( .IN1(n15032), .IN2(g6561), .QN(n13440) );
  INVX0 U19381 ( .INP(n3776), .ZN(n15032) );
  NAND2X0 U19382 ( .IN1(g6573), .IN2(g6565), .QN(n3776) );
  NAND2X0 U19383 ( .IN1(n18495), .IN2(n18496), .QN(g25758) );
  NAND2X0 U19384 ( .IN1(n11059), .IN2(g6494), .QN(n18496) );
  NAND2X0 U19385 ( .IN1(n18497), .IN2(n10940), .QN(n18495) );
  NOR2X0 U19386 ( .IN1(n18498), .IN2(g9817), .QN(n18497) );
  NOR2X0 U19387 ( .IN1(n18499), .IN2(g6444), .QN(n18498) );
  NOR2X0 U19388 ( .IN1(n5719), .IN2(g6494), .QN(n18499) );
  NAND2X0 U19389 ( .IN1(n18500), .IN2(n18501), .QN(g25757) );
  NAND2X0 U19390 ( .IN1(n10928), .IN2(g6727), .QN(n18501) );
  NAND2X0 U19391 ( .IN1(n11059), .IN2(g6444), .QN(n18500) );
  NOR2X0 U19392 ( .IN1(n11055), .IN2(n5563), .QN(g25756) );
  NAND2X0 U19393 ( .IN1(n18502), .IN2(n18503), .QN(g25750) );
  NAND2X0 U19394 ( .IN1(n11286), .IN2(g6159), .QN(n18503) );
  NAND2X0 U19395 ( .IN1(n15137), .IN2(g6195), .QN(n18502) );
  NAND2X0 U19396 ( .IN1(n18504), .IN2(n18505), .QN(g25749) );
  NAND2X0 U19397 ( .IN1(n11286), .IN2(g6191), .QN(n18505) );
  NOR2X0 U19398 ( .IN1(n18506), .IN2(n18507), .QN(n18504) );
  NOR2X0 U19399 ( .IN1(g6187), .IN2(n18508), .QN(n18507) );
  NAND2X0 U19400 ( .IN1(n18509), .IN2(n5667), .QN(n18508) );
  NOR2X0 U19401 ( .IN1(n11055), .IN2(n13434), .QN(n18509) );
  NOR2X0 U19402 ( .IN1(n5453), .IN2(n18510), .QN(n18506) );
  NOR2X0 U19403 ( .IN1(n11054), .IN2(n18511), .QN(n18510) );
  NOR2X0 U19404 ( .IN1(n5667), .IN2(n13434), .QN(n18511) );
  NAND2X0 U19405 ( .IN1(n18512), .IN2(n18513), .QN(g25747) );
  NAND2X0 U19406 ( .IN1(n11286), .IN2(g6167), .QN(n18513) );
  INVX0 U19407 ( .INP(n15137), .ZN(n11286) );
  NAND2X0 U19408 ( .IN1(n13434), .IN2(n10937), .QN(n15137) );
  NOR2X0 U19409 ( .IN1(n18514), .IN2(n18515), .QN(n18512) );
  NOR2X0 U19410 ( .IN1(n10153), .IN2(n10887), .QN(n18515) );
  NOR2X0 U19411 ( .IN1(n11054), .IN2(n18516), .QN(n18514) );
  NAND2X0 U19412 ( .IN1(n5430), .IN2(n18517), .QN(n18516) );
  INVX0 U19413 ( .INP(n13434), .ZN(n18517) );
  NAND2X0 U19414 ( .IN1(n15160), .IN2(g6215), .QN(n13434) );
  INVX0 U19415 ( .INP(n3810), .ZN(n15160) );
  NAND2X0 U19416 ( .IN1(g6227), .IN2(g6219), .QN(n3810) );
  NAND2X0 U19417 ( .IN1(n18518), .IN2(n18519), .QN(g25744) );
  NAND2X0 U19418 ( .IN1(n11059), .IN2(g6148), .QN(n18519) );
  NAND2X0 U19419 ( .IN1(n18520), .IN2(n10939), .QN(n18518) );
  NOR2X0 U19420 ( .IN1(n18521), .IN2(g9741), .QN(n18520) );
  NOR2X0 U19421 ( .IN1(n18522), .IN2(g6098), .QN(n18521) );
  NOR2X0 U19422 ( .IN1(g6148), .IN2(n5718), .QN(n18522) );
  NAND2X0 U19423 ( .IN1(n18523), .IN2(n18524), .QN(g25743) );
  NAND2X0 U19424 ( .IN1(test_so69), .IN2(n10938), .QN(n18524) );
  NAND2X0 U19425 ( .IN1(n11060), .IN2(g6098), .QN(n18523) );
  NOR2X0 U19426 ( .IN1(n11054), .IN2(n5568), .QN(g25742) );
  NAND2X0 U19427 ( .IN1(n18525), .IN2(n18526), .QN(g25736) );
  NAND2X0 U19428 ( .IN1(n11292), .IN2(g5813), .QN(n18526) );
  NAND2X0 U19429 ( .IN1(n15265), .IN2(g5849), .QN(n18525) );
  NAND2X0 U19430 ( .IN1(n18527), .IN2(n18528), .QN(g25735) );
  NAND2X0 U19431 ( .IN1(test_so83), .IN2(n11292), .QN(n18528) );
  NOR2X0 U19432 ( .IN1(n18529), .IN2(n18530), .QN(n18527) );
  NOR2X0 U19433 ( .IN1(g5841), .IN2(n18531), .QN(n18530) );
  NAND2X0 U19434 ( .IN1(n18532), .IN2(n5663), .QN(n18531) );
  NOR2X0 U19435 ( .IN1(n11053), .IN2(n13433), .QN(n18532) );
  NOR2X0 U19436 ( .IN1(n5449), .IN2(n18533), .QN(n18529) );
  NOR2X0 U19437 ( .IN1(n11053), .IN2(n18534), .QN(n18533) );
  NOR2X0 U19438 ( .IN1(n5663), .IN2(n13433), .QN(n18534) );
  NAND2X0 U19439 ( .IN1(n18535), .IN2(n18536), .QN(g25733) );
  NAND2X0 U19440 ( .IN1(n11292), .IN2(g5821), .QN(n18536) );
  INVX0 U19441 ( .INP(n15265), .ZN(n11292) );
  NAND2X0 U19442 ( .IN1(n13433), .IN2(n10938), .QN(n15265) );
  NOR2X0 U19443 ( .IN1(n18537), .IN2(n18538), .QN(n18535) );
  NOR2X0 U19444 ( .IN1(n10131), .IN2(n10886), .QN(n18538) );
  NOR2X0 U19445 ( .IN1(n11053), .IN2(n18539), .QN(n18537) );
  NAND2X0 U19446 ( .IN1(n5429), .IN2(n18540), .QN(n18539) );
  INVX0 U19447 ( .INP(n13433), .ZN(n18540) );
  NAND2X0 U19448 ( .IN1(n15288), .IN2(g5869), .QN(n13433) );
  INVX0 U19449 ( .INP(n3844), .ZN(n15288) );
  NAND2X0 U19450 ( .IN1(test_so36), .IN2(g5873), .QN(n3844) );
  NAND2X0 U19451 ( .IN1(n18541), .IN2(n18542), .QN(g25730) );
  NAND2X0 U19452 ( .IN1(n11060), .IN2(g5802), .QN(n18542) );
  NAND2X0 U19453 ( .IN1(n18543), .IN2(n10939), .QN(n18541) );
  NOR2X0 U19454 ( .IN1(n18544), .IN2(g9680), .QN(n18543) );
  NOR2X0 U19455 ( .IN1(n18545), .IN2(g5752), .QN(n18544) );
  NOR2X0 U19456 ( .IN1(n5722), .IN2(g5802), .QN(n18545) );
  NAND2X0 U19457 ( .IN1(n18546), .IN2(n18547), .QN(g25729) );
  NAND2X0 U19458 ( .IN1(n10928), .IN2(g6035), .QN(n18547) );
  NAND2X0 U19459 ( .IN1(n11060), .IN2(g5752), .QN(n18546) );
  NOR2X0 U19460 ( .IN1(n10651), .IN2(n11018), .QN(g25728) );
  NAND2X0 U19461 ( .IN1(n18548), .IN2(n18549), .QN(g25722) );
  NAND2X0 U19462 ( .IN1(n11250), .IN2(g5467), .QN(n18549) );
  NAND2X0 U19463 ( .IN1(n11251), .IN2(g5503), .QN(n18548) );
  NAND2X0 U19464 ( .IN1(n18550), .IN2(n18551), .QN(g25721) );
  NAND2X0 U19465 ( .IN1(n11250), .IN2(g5499), .QN(n18551) );
  NOR2X0 U19466 ( .IN1(n18552), .IN2(n18553), .QN(n18550) );
  NOR2X0 U19467 ( .IN1(g5495), .IN2(n18554), .QN(n18553) );
  NAND2X0 U19468 ( .IN1(n18555), .IN2(n5660), .QN(n18554) );
  NOR2X0 U19469 ( .IN1(n11052), .IN2(n15393), .QN(n18555) );
  NOR2X0 U19470 ( .IN1(n5446), .IN2(n18556), .QN(n18552) );
  NOR2X0 U19471 ( .IN1(n11052), .IN2(n18557), .QN(n18556) );
  NOR2X0 U19472 ( .IN1(n5660), .IN2(n15393), .QN(n18557) );
  NAND2X0 U19473 ( .IN1(n18558), .IN2(n18559), .QN(g25719) );
  NAND2X0 U19474 ( .IN1(n11250), .IN2(g5475), .QN(n18559) );
  INVX0 U19475 ( .INP(n11251), .ZN(n11250) );
  NAND2X0 U19476 ( .IN1(n15393), .IN2(n10940), .QN(n11251) );
  NOR2X0 U19477 ( .IN1(n18560), .IN2(n18561), .QN(n18558) );
  NOR2X0 U19478 ( .IN1(n10139), .IN2(n10886), .QN(n18561) );
  NOR2X0 U19479 ( .IN1(n11052), .IN2(n18562), .QN(n18560) );
  NAND2X0 U19480 ( .IN1(n5425), .IN2(n13426), .QN(n18562) );
  INVX0 U19481 ( .INP(n15393), .ZN(n13426) );
  NAND2X0 U19482 ( .IN1(n15417), .IN2(g5523), .QN(n15393) );
  INVX0 U19483 ( .INP(n3877), .ZN(n15417) );
  NAND2X0 U19484 ( .IN1(g5535), .IN2(g5527), .QN(n3877) );
  NAND2X0 U19485 ( .IN1(n18563), .IN2(n18564), .QN(g25716) );
  NAND2X0 U19486 ( .IN1(n11061), .IN2(g5456), .QN(n18564) );
  NAND2X0 U19487 ( .IN1(n18565), .IN2(n10939), .QN(n18563) );
  NOR2X0 U19488 ( .IN1(test_so35), .IN2(n18566), .QN(n18565) );
  NOR2X0 U19489 ( .IN1(n18567), .IN2(g5406), .QN(n18566) );
  NOR2X0 U19490 ( .IN1(n19405), .IN2(g5456), .QN(n18567) );
  NAND2X0 U19491 ( .IN1(n18568), .IN2(n18569), .QN(g25715) );
  NAND2X0 U19492 ( .IN1(n10928), .IN2(g5689), .QN(n18569) );
  NAND2X0 U19493 ( .IN1(n11061), .IN2(g5406), .QN(n18568) );
  INVX0 U19494 ( .INP(n14285), .ZN(g25714) );
  NAND2X0 U19495 ( .IN1(n10928), .IN2(g5535), .QN(n14285) );
  NAND2X0 U19496 ( .IN1(n18570), .IN2(n18571), .QN(g25708) );
  NAND2X0 U19497 ( .IN1(n18572), .IN2(g5120), .QN(n18571) );
  NAND2X0 U19498 ( .IN1(n15520), .IN2(g5156), .QN(n18570) );
  NAND2X0 U19499 ( .IN1(n18573), .IN2(n18574), .QN(g25707) );
  NAND2X0 U19500 ( .IN1(n18572), .IN2(g5152), .QN(n18574) );
  NOR2X0 U19501 ( .IN1(n18575), .IN2(n18576), .QN(n18573) );
  NOR2X0 U19502 ( .IN1(test_so98), .IN2(n18577), .QN(n18576) );
  NAND2X0 U19503 ( .IN1(n18578), .IN2(n5658), .QN(n18577) );
  NOR2X0 U19504 ( .IN1(n11056), .IN2(n13429), .QN(n18578) );
  NOR2X0 U19505 ( .IN1(n18579), .IN2(n10682), .QN(n18575) );
  NOR2X0 U19506 ( .IN1(n11052), .IN2(n18580), .QN(n18579) );
  NOR2X0 U19507 ( .IN1(n5658), .IN2(n13429), .QN(n18580) );
  NAND2X0 U19508 ( .IN1(n18581), .IN2(n18582), .QN(g25706) );
  NAND2X0 U19509 ( .IN1(test_so98), .IN2(n18572), .QN(n18582) );
  NAND2X0 U19510 ( .IN1(n15520), .IN2(g5142), .QN(n18581) );
  NAND2X0 U19511 ( .IN1(n18583), .IN2(n18584), .QN(g25705) );
  NAND2X0 U19512 ( .IN1(test_so96), .IN2(n18572), .QN(n18584) );
  INVX0 U19513 ( .INP(n15520), .ZN(n18572) );
  NAND2X0 U19514 ( .IN1(n13429), .IN2(n10940), .QN(n15520) );
  NOR2X0 U19515 ( .IN1(n18585), .IN2(n18586), .QN(n18583) );
  NOR2X0 U19516 ( .IN1(n10129), .IN2(n10886), .QN(n18586) );
  NOR2X0 U19517 ( .IN1(n11052), .IN2(n18587), .QN(n18585) );
  NAND2X0 U19518 ( .IN1(g32975), .IN2(n10654), .QN(n18587) );
  INVX0 U19519 ( .INP(n13429), .ZN(g32975) );
  NAND2X0 U19520 ( .IN1(n15543), .IN2(g5176), .QN(n13429) );
  INVX0 U19521 ( .INP(n3910), .ZN(n15543) );
  NAND2X0 U19522 ( .IN1(g5188), .IN2(g5180), .QN(n3910) );
  NOR2X0 U19523 ( .IN1(n10194), .IN2(n18588), .QN(g25704) );
  NOR2X0 U19524 ( .IN1(n11052), .IN2(g5069), .QN(n18588) );
  NAND2X0 U19525 ( .IN1(n18589), .IN2(n18590), .QN(g25703) );
  NAND2X0 U19526 ( .IN1(n11062), .IN2(g5112), .QN(n18590) );
  NAND2X0 U19527 ( .IN1(n18591), .IN2(n10940), .QN(n18589) );
  NOR2X0 U19528 ( .IN1(n18592), .IN2(g9497), .QN(n18591) );
  NOR2X0 U19529 ( .IN1(n18593), .IN2(g5022), .QN(n18592) );
  NOR2X0 U19530 ( .IN1(n5690), .IN2(g5112), .QN(n18593) );
  NAND2X0 U19531 ( .IN1(n18594), .IN2(n18595), .QN(g25702) );
  NAND2X0 U19532 ( .IN1(test_so32), .IN2(n11081), .QN(n18595) );
  NAND2X0 U19533 ( .IN1(n18596), .IN2(n10941), .QN(n18594) );
  NOR2X0 U19534 ( .IN1(n18597), .IN2(g9553), .QN(n18596) );
  NOR2X0 U19535 ( .IN1(n18598), .IN2(g5062), .QN(n18597) );
  NOR2X0 U19536 ( .IN1(test_so32), .IN2(n5689), .QN(n18598) );
  NAND2X0 U19537 ( .IN1(n18599), .IN2(n18600), .QN(g25701) );
  NAND2X0 U19538 ( .IN1(test_so10), .IN2(n10941), .QN(n18600) );
  NAND2X0 U19539 ( .IN1(n11063), .IN2(g5062), .QN(n18599) );
  NOR2X0 U19540 ( .IN1(n11054), .IN2(n5567), .QN(g25700) );
  NAND2X0 U19541 ( .IN1(n18601), .IN2(n18602), .QN(g25699) );
  NAND2X0 U19542 ( .IN1(n11063), .IN2(g5097), .QN(n18602) );
  NOR2X0 U19543 ( .IN1(n18603), .IN2(n18604), .QN(n18601) );
  INVX0 U19544 ( .INP(n18605), .ZN(n18604) );
  NAND2X0 U19545 ( .IN1(n5669), .IN2(n5014), .QN(n18605) );
  NOR2X0 U19546 ( .IN1(n5669), .IN2(n18606), .QN(n18603) );
  INVX0 U19547 ( .INP(n18607), .ZN(n18606) );
  NOR2X0 U19548 ( .IN1(n11054), .IN2(n5014), .QN(n18607) );
  NAND2X0 U19549 ( .IN1(n18608), .IN2(n18609), .QN(g25698) );
  NAND2X0 U19550 ( .IN1(n11064), .IN2(g5092), .QN(n18609) );
  NOR2X0 U19551 ( .IN1(n18610), .IN2(n18611), .QN(n18608) );
  NOR2X0 U19552 ( .IN1(g5097), .IN2(n18612), .QN(n18611) );
  NOR2X0 U19553 ( .IN1(n5753), .IN2(n18613), .QN(n18610) );
  NAND2X0 U19554 ( .IN1(n10929), .IN2(n18612), .QN(n18613) );
  INVX0 U19555 ( .INP(n5016), .ZN(n18612) );
  XOR2X1 U19556 ( .IN1(n18614), .IN2(n5681), .Q(g25697) );
  NAND2X0 U19557 ( .IN1(n10929), .IN2(g5092), .QN(n18614) );
  NAND2X0 U19558 ( .IN1(n18615), .IN2(n18616), .QN(g25696) );
  NAND2X0 U19559 ( .IN1(n18617), .IN2(n10194), .QN(n18616) );
  NOR2X0 U19560 ( .IN1(n5455), .IN2(n11022), .QN(n18617) );
  NOR2X0 U19561 ( .IN1(n18618), .IN2(n18619), .QN(n18615) );
  NOR2X0 U19562 ( .IN1(g5080), .IN2(n18620), .QN(n18619) );
  NAND2X0 U19563 ( .IN1(n18621), .IN2(n18622), .QN(n18620) );
  NAND2X0 U19564 ( .IN1(n10193), .IN2(g5077), .QN(n18622) );
  NOR2X0 U19565 ( .IN1(n5893), .IN2(n18621), .QN(n18618) );
  NOR2X0 U19566 ( .IN1(g5084), .IN2(n11023), .QN(n18621) );
  NOR2X0 U19567 ( .IN1(n5455), .IN2(n18623), .QN(g25695) );
  NOR2X0 U19568 ( .IN1(n11057), .IN2(n18624), .QN(n18623) );
  NAND2X0 U19569 ( .IN1(n18625), .IN2(n18626), .QN(n18624) );
  NAND2X0 U19570 ( .IN1(n10193), .IN2(g5084), .QN(n18626) );
  NAND2X0 U19571 ( .IN1(n10194), .IN2(n5681), .QN(n18625) );
  NAND2X0 U19572 ( .IN1(n18627), .IN2(n18628), .QN(g25691) );
  NAND2X0 U19573 ( .IN1(n10631), .IN2(n18629), .QN(n18628) );
  NAND2X0 U19574 ( .IN1(n18630), .IN2(n18631), .QN(n18629) );
  NOR2X0 U19575 ( .IN1(n10644), .IN2(n18632), .QN(n18631) );
  NAND2X0 U19576 ( .IN1(n12424), .IN2(g4098), .QN(n18632) );
  NOR2X0 U19577 ( .IN1(g4141), .IN2(g4082), .QN(n12424) );
  NOR2X0 U19578 ( .IN1(g4057), .IN2(n18633), .QN(n18630) );
  NAND2X0 U19579 ( .IN1(n5416), .IN2(n13425), .QN(n18633) );
  INVX0 U19580 ( .INP(n15663), .ZN(n13425) );
  NAND2X0 U19581 ( .IN1(n5340), .IN2(g4087), .QN(n15663) );
  INVX0 U19582 ( .INP(n14906), .ZN(n10631) );
  NAND2X0 U19583 ( .IN1(n11065), .IN2(g4125), .QN(n18627) );
  NAND2X0 U19584 ( .IN1(n18634), .IN2(n18635), .QN(g25690) );
  NAND2X0 U19585 ( .IN1(n11065), .IN2(g4169), .QN(n18635) );
  NAND2X0 U19586 ( .IN1(n18636), .IN2(n10941), .QN(n18634) );
  NOR2X0 U19587 ( .IN1(n10133), .IN2(g4125), .QN(n18636) );
  NAND2X0 U19588 ( .IN1(n18637), .IN2(n18638), .QN(g25687) );
  NAND2X0 U19589 ( .IN1(n11065), .IN2(g4057), .QN(n18638) );
  INVX0 U19590 ( .INP(n18639), .ZN(n18637) );
  NAND2X0 U19591 ( .IN1(n18640), .IN2(n18641), .QN(n18639) );
  NAND2X0 U19592 ( .IN1(n16692), .IN2(n5026), .QN(n18641) );
  INVX0 U19593 ( .INP(n15661), .ZN(n16692) );
  NAND2X0 U19594 ( .IN1(n5612), .IN2(n18642), .QN(n18640) );
  NOR2X0 U19595 ( .IN1(n1269), .IN2(n5729), .QN(n18642) );
  NAND2X0 U19596 ( .IN1(g4057), .IN2(g4064), .QN(n1269) );
  NAND2X0 U19597 ( .IN1(n18643), .IN2(n18644), .QN(g25686) );
  NAND2X0 U19598 ( .IN1(n18645), .IN2(g4064), .QN(n18644) );
  NAND2X0 U19599 ( .IN1(n18646), .IN2(n10942), .QN(n18645) );
  NAND2X0 U19600 ( .IN1(n5711), .IN2(g4169), .QN(n18646) );
  NAND2X0 U19601 ( .IN1(n18647), .IN2(n5416), .QN(n18643) );
  NOR2X0 U19602 ( .IN1(n5711), .IN2(n15661), .QN(n18647) );
  NAND2X0 U19603 ( .IN1(n10929), .IN2(g4169), .QN(n15661) );
  NAND2X0 U19604 ( .IN1(n18648), .IN2(n14906), .QN(g25685) );
  NAND2X0 U19605 ( .IN1(n5729), .IN2(n10941), .QN(n14906) );
  NOR2X0 U19606 ( .IN1(n18649), .IN2(n18650), .QN(n18648) );
  NOR2X0 U19607 ( .IN1(n10612), .IN2(n10886), .QN(n18650) );
  NOR2X0 U19608 ( .IN1(n11058), .IN2(g4064), .QN(n18649) );
  NAND2X0 U19609 ( .IN1(n18651), .IN2(n18652), .QN(g25684) );
  NAND2X0 U19610 ( .IN1(n18653), .IN2(g3813), .QN(n18652) );
  NAND2X0 U19611 ( .IN1(n15669), .IN2(g3849), .QN(n18651) );
  NAND2X0 U19612 ( .IN1(n18654), .IN2(n18655), .QN(g25683) );
  NAND2X0 U19613 ( .IN1(n18653), .IN2(g3845), .QN(n18655) );
  NOR2X0 U19614 ( .IN1(n18656), .IN2(n18657), .QN(n18654) );
  NOR2X0 U19615 ( .IN1(test_so97), .IN2(n18658), .QN(n18657) );
  NAND2X0 U19616 ( .IN1(n18659), .IN2(n5662), .QN(n18658) );
  NOR2X0 U19617 ( .IN1(n11058), .IN2(n13445), .QN(n18659) );
  NOR2X0 U19618 ( .IN1(n18660), .IN2(n10683), .QN(n18656) );
  NOR2X0 U19619 ( .IN1(n11058), .IN2(n18661), .QN(n18660) );
  NOR2X0 U19620 ( .IN1(n5662), .IN2(n13445), .QN(n18661) );
  NAND2X0 U19621 ( .IN1(n18662), .IN2(n18663), .QN(g25682) );
  NAND2X0 U19622 ( .IN1(test_so97), .IN2(n18653), .QN(n18663) );
  NAND2X0 U19623 ( .IN1(n15669), .IN2(g3835), .QN(n18662) );
  NAND2X0 U19624 ( .IN1(n18664), .IN2(n18665), .QN(g25681) );
  NAND2X0 U19625 ( .IN1(n18653), .IN2(g3821), .QN(n18665) );
  INVX0 U19626 ( .INP(n15669), .ZN(n18653) );
  NAND2X0 U19627 ( .IN1(n13445), .IN2(n10942), .QN(n15669) );
  NOR2X0 U19628 ( .IN1(n18666), .IN2(n18667), .QN(n18664) );
  NOR2X0 U19629 ( .IN1(n10130), .IN2(n10886), .QN(n18667) );
  NOR2X0 U19630 ( .IN1(n11058), .IN2(n18668), .QN(n18666) );
  NAND2X0 U19631 ( .IN1(n5428), .IN2(n18669), .QN(n18668) );
  INVX0 U19632 ( .INP(n13445), .ZN(n18669) );
  NAND2X0 U19633 ( .IN1(test_so33), .IN2(n15693), .QN(n13445) );
  INVX0 U19634 ( .INP(n3953), .ZN(n15693) );
  NAND2X0 U19635 ( .IN1(g3881), .IN2(g3873), .QN(n3953) );
  NAND2X0 U19636 ( .IN1(n18670), .IN2(n18671), .QN(g25678) );
  NAND2X0 U19637 ( .IN1(n11065), .IN2(g3802), .QN(n18671) );
  NAND2X0 U19638 ( .IN1(n18672), .IN2(n10942), .QN(n18670) );
  NOR2X0 U19639 ( .IN1(n18673), .IN2(g8398), .QN(n18672) );
  NOR2X0 U19640 ( .IN1(n18674), .IN2(g3752), .QN(n18673) );
  NOR2X0 U19641 ( .IN1(n5721), .IN2(g3802), .QN(n18674) );
  NAND2X0 U19642 ( .IN1(n18675), .IN2(n18676), .QN(g25677) );
  NAND2X0 U19643 ( .IN1(n10930), .IN2(g4040), .QN(n18676) );
  NAND2X0 U19644 ( .IN1(n11061), .IN2(g3752), .QN(n18675) );
  NOR2X0 U19645 ( .IN1(n11043), .IN2(n5564), .QN(g25676) );
  NAND2X0 U19646 ( .IN1(n18677), .IN2(n18678), .QN(g25670) );
  NAND2X0 U19647 ( .IN1(n11498), .IN2(g3462), .QN(n18678) );
  NAND2X0 U19648 ( .IN1(n15796), .IN2(g3498), .QN(n18677) );
  NAND2X0 U19649 ( .IN1(n18679), .IN2(n18680), .QN(g25669) );
  NAND2X0 U19650 ( .IN1(n11498), .IN2(g3494), .QN(n18680) );
  NOR2X0 U19651 ( .IN1(n18681), .IN2(n18682), .QN(n18679) );
  NOR2X0 U19652 ( .IN1(g3490), .IN2(n18683), .QN(n18682) );
  NAND2X0 U19653 ( .IN1(n18684), .IN2(n5668), .QN(n18683) );
  NOR2X0 U19654 ( .IN1(n11043), .IN2(n13444), .QN(n18684) );
  NOR2X0 U19655 ( .IN1(n5454), .IN2(n18685), .QN(n18681) );
  NOR2X0 U19656 ( .IN1(n11043), .IN2(n18686), .QN(n18685) );
  NOR2X0 U19657 ( .IN1(n5668), .IN2(n13444), .QN(n18686) );
  NAND2X0 U19658 ( .IN1(n18687), .IN2(n18688), .QN(g25667) );
  NAND2X0 U19659 ( .IN1(n11498), .IN2(g3470), .QN(n18688) );
  INVX0 U19660 ( .INP(n15796), .ZN(n11498) );
  NAND2X0 U19661 ( .IN1(n13444), .IN2(n10942), .QN(n15796) );
  NOR2X0 U19662 ( .IN1(n18689), .IN2(n18690), .QN(n18687) );
  NOR2X0 U19663 ( .IN1(n10149), .IN2(n10885), .QN(n18690) );
  NOR2X0 U19664 ( .IN1(n11043), .IN2(n18691), .QN(n18689) );
  NAND2X0 U19665 ( .IN1(n5424), .IN2(n18692), .QN(n18691) );
  INVX0 U19666 ( .INP(n13444), .ZN(n18692) );
  NAND2X0 U19667 ( .IN1(n15819), .IN2(g3518), .QN(n13444) );
  INVX0 U19668 ( .INP(n3986), .ZN(n15819) );
  NAND2X0 U19669 ( .IN1(g3530), .IN2(g3522), .QN(n3986) );
  NAND2X0 U19670 ( .IN1(n18693), .IN2(n18694), .QN(g25664) );
  NAND2X0 U19671 ( .IN1(n11065), .IN2(g3451), .QN(n18694) );
  NAND2X0 U19672 ( .IN1(n18695), .IN2(n10942), .QN(n18693) );
  NOR2X0 U19673 ( .IN1(n18696), .IN2(g8342), .QN(n18695) );
  NOR2X0 U19674 ( .IN1(n18697), .IN2(g3401), .QN(n18696) );
  NOR2X0 U19675 ( .IN1(n5717), .IN2(g3451), .QN(n18697) );
  NAND2X0 U19676 ( .IN1(n18698), .IN2(n18699), .QN(g25663) );
  NAND2X0 U19677 ( .IN1(n10930), .IN2(g3689), .QN(n18699) );
  NAND2X0 U19678 ( .IN1(n11065), .IN2(g3401), .QN(n18698) );
  NOR2X0 U19679 ( .IN1(n11043), .IN2(n5569), .QN(g25662) );
  NAND2X0 U19680 ( .IN1(n18700), .IN2(n18701), .QN(g25656) );
  NAND2X0 U19681 ( .IN1(n11462), .IN2(g3111), .QN(n18701) );
  NAND2X0 U19682 ( .IN1(n15924), .IN2(g3147), .QN(n18700) );
  NAND2X0 U19683 ( .IN1(n18702), .IN2(n18703), .QN(g25655) );
  NAND2X0 U19684 ( .IN1(n11462), .IN2(g3143), .QN(n18703) );
  NOR2X0 U19685 ( .IN1(n18704), .IN2(n18705), .QN(n18702) );
  NOR2X0 U19686 ( .IN1(g3139), .IN2(n18706), .QN(n18705) );
  NAND2X0 U19687 ( .IN1(n18707), .IN2(n5661), .QN(n18706) );
  NOR2X0 U19688 ( .IN1(n11043), .IN2(n15923), .QN(n18707) );
  NOR2X0 U19689 ( .IN1(n5447), .IN2(n18708), .QN(n18704) );
  NOR2X0 U19690 ( .IN1(n11044), .IN2(n18709), .QN(n18708) );
  NOR2X0 U19691 ( .IN1(n5661), .IN2(n15923), .QN(n18709) );
  NAND2X0 U19692 ( .IN1(n18710), .IN2(n18711), .QN(g25653) );
  NAND2X0 U19693 ( .IN1(n11462), .IN2(g3119), .QN(n18711) );
  INVX0 U19694 ( .INP(n15924), .ZN(n11462) );
  NAND2X0 U19695 ( .IN1(n15923), .IN2(n10942), .QN(n15924) );
  NOR2X0 U19696 ( .IN1(n18712), .IN2(n18713), .QN(n18710) );
  NOR2X0 U19697 ( .IN1(n10170), .IN2(n10885), .QN(n18713) );
  NOR2X0 U19698 ( .IN1(n11044), .IN2(n18714), .QN(n18712) );
  NAND2X0 U19699 ( .IN1(n5423), .IN2(n13437), .QN(n18714) );
  INVX0 U19700 ( .INP(n15923), .ZN(n13437) );
  NAND2X0 U19701 ( .IN1(n15949), .IN2(g3167), .QN(n15923) );
  INVX0 U19702 ( .INP(n582), .ZN(n15949) );
  NAND2X0 U19703 ( .IN1(g3179), .IN2(g3171), .QN(n582) );
  NAND2X0 U19704 ( .IN1(n18715), .IN2(n18716), .QN(g25650) );
  NAND2X0 U19705 ( .IN1(n11064), .IN2(g3100), .QN(n18716) );
  NAND2X0 U19706 ( .IN1(n18717), .IN2(n10942), .QN(n18715) );
  NOR2X0 U19707 ( .IN1(n18718), .IN2(g8277), .QN(n18717) );
  NOR2X0 U19708 ( .IN1(n18719), .IN2(g3050), .QN(n18718) );
  NOR2X0 U19709 ( .IN1(n5723), .IN2(g3100), .QN(n18719) );
  NAND2X0 U19710 ( .IN1(n18720), .IN2(n18721), .QN(g25649) );
  NAND2X0 U19711 ( .IN1(n10930), .IN2(g3338), .QN(n18721) );
  NAND2X0 U19712 ( .IN1(n11064), .IN2(g3050), .QN(n18720) );
  NOR2X0 U19713 ( .IN1(n11045), .IN2(n5390), .QN(g25648) );
  NAND2X0 U19714 ( .IN1(n18722), .IN2(n18723), .QN(g25639) );
  INVX0 U19715 ( .INP(n5045), .ZN(n18723) );
  NOR2X0 U19716 ( .IN1(n18724), .IN2(n18725), .QN(n18722) );
  NOR2X0 U19717 ( .IN1(n11046), .IN2(n18726), .QN(n18725) );
  INVX0 U19718 ( .INP(n16060), .ZN(n18726) );
  NOR2X0 U19719 ( .IN1(g2715), .IN2(n5465), .QN(n16060) );
  NOR2X0 U19720 ( .IN1(n5299), .IN2(n10885), .QN(n18724) );
  NAND2X0 U19721 ( .IN1(n18727), .IN2(n18728), .QN(g25638) );
  NAND2X0 U19722 ( .IN1(n11064), .IN2(g1564), .QN(n18728) );
  NAND2X0 U19723 ( .IN1(n18729), .IN2(n10942), .QN(n18727) );
  NAND2X0 U19724 ( .IN1(n18730), .IN2(n18731), .QN(n18729) );
  NAND2X0 U19725 ( .IN1(n18732), .IN2(g1559), .QN(n18731) );
  NAND2X0 U19726 ( .IN1(n18733), .IN2(n5441), .QN(n18730) );
  NAND2X0 U19727 ( .IN1(n18734), .IN2(n18735), .QN(g25637) );
  NAND2X0 U19728 ( .IN1(n18736), .IN2(n18732), .QN(n18735) );
  NOR2X0 U19729 ( .IN1(n5768), .IN2(n11023), .QN(n18736) );
  NAND2X0 U19730 ( .IN1(n18737), .IN2(g1559), .QN(n18734) );
  NAND2X0 U19731 ( .IN1(n18738), .IN2(n10943), .QN(n18737) );
  INVX0 U19732 ( .INP(n18733), .ZN(n18738) );
  NOR2X0 U19733 ( .IN1(n18732), .IN2(g1554), .QN(n18733) );
  NAND2X0 U19734 ( .IN1(n18739), .IN2(n18740), .QN(g25636) );
  NAND2X0 U19735 ( .IN1(n11064), .IN2(g1521), .QN(n18740) );
  NAND2X0 U19736 ( .IN1(n18741), .IN2(n10943), .QN(n18739) );
  NAND2X0 U19737 ( .IN1(n18742), .IN2(n18743), .QN(n18741) );
  NAND2X0 U19738 ( .IN1(n16417), .IN2(n13753), .QN(n18743) );
  INVX0 U19739 ( .INP(n18744), .ZN(n16417) );
  NAND2X0 U19740 ( .IN1(n18745), .IN2(g1306), .QN(n18742) );
  NAND2X0 U19741 ( .IN1(n13753), .IN2(g7946), .QN(n18745) );
  INVX0 U19742 ( .INP(n17035), .ZN(n13753) );
  NAND2X0 U19743 ( .IN1(test_so49), .IN2(g1514), .QN(n17035) );
  NAND2X0 U19744 ( .IN1(n18746), .IN2(n18747), .QN(g25635) );
  NAND2X0 U19745 ( .IN1(n18748), .IN2(g1484), .QN(n18747) );
  NAND2X0 U19746 ( .IN1(n18749), .IN2(n10944), .QN(n18748) );
  NAND2X0 U19747 ( .IN1(n18750), .IN2(n18211), .QN(n18749) );
  NOR2X0 U19748 ( .IN1(g1300), .IN2(n18751), .QN(n18750) );
  NAND2X0 U19749 ( .IN1(n18752), .IN2(g1300), .QN(n18746) );
  NAND2X0 U19750 ( .IN1(n18753), .IN2(n18754), .QN(n18752) );
  NAND2X0 U19751 ( .IN1(n18755), .IN2(n10944), .QN(n18754) );
  NAND2X0 U19752 ( .IN1(n18211), .IN2(g1484), .QN(n18755) );
  NOR2X0 U19753 ( .IN1(n10536), .IN2(test_so12), .QN(n18211) );
  NOR2X0 U19754 ( .IN1(n18756), .IN2(n18757), .QN(g25634) );
  NAND2X0 U19755 ( .IN1(n18234), .IN2(n10650), .QN(n18757) );
  NAND2X0 U19756 ( .IN1(n18758), .IN2(n18759), .QN(n18234) );
  INVX0 U19757 ( .INP(n18760), .ZN(n18759) );
  NOR2X0 U19758 ( .IN1(n5655), .IN2(n10580), .QN(n18758) );
  NOR2X0 U19759 ( .IN1(n18761), .IN2(n18762), .QN(n18756) );
  NOR2X0 U19760 ( .IN1(n10580), .IN2(n11023), .QN(n18762) );
  NOR2X0 U19761 ( .IN1(n18760), .IN2(n18763), .QN(n18761) );
  NAND2X0 U19762 ( .IN1(n18764), .IN2(n18765), .QN(g25633) );
  NAND2X0 U19763 ( .IN1(n11064), .IN2(g1379), .QN(n18765) );
  NAND2X0 U19764 ( .IN1(n18766), .IN2(n10945), .QN(n18764) );
  NAND2X0 U19765 ( .IN1(n18767), .IN2(n18768), .QN(n18766) );
  NAND2X0 U19766 ( .IN1(n18241), .IN2(g1384), .QN(n18768) );
  NAND2X0 U19767 ( .IN1(n18769), .IN2(n10105), .QN(n18767) );
  NOR2X0 U19768 ( .IN1(n5322), .IN2(n18241), .QN(n18769) );
  NAND2X0 U19769 ( .IN1(n18770), .IN2(n18771), .QN(g25632) );
  NAND2X0 U19770 ( .IN1(n18772), .IN2(g1312), .QN(n18771) );
  NAND2X0 U19771 ( .IN1(n18241), .IN2(n10946), .QN(n18772) );
  NAND2X0 U19772 ( .IN1(n18773), .IN2(n18774), .QN(n18770) );
  NOR2X0 U19773 ( .IN1(n5322), .IN2(n11022), .QN(n18774) );
  NOR2X0 U19774 ( .IN1(n18775), .IN2(n18776), .QN(n18773) );
  NOR2X0 U19775 ( .IN1(n10620), .IN2(n18241), .QN(n18776) );
  NOR2X0 U19776 ( .IN1(n17903), .IN2(n18777), .QN(n18775) );
  NAND2X0 U19777 ( .IN1(g1361), .IN2(g1373), .QN(n18777) );
  NOR2X0 U19778 ( .IN1(n11047), .IN2(n18778), .QN(g25631) );
  NOR2X0 U19779 ( .IN1(n18779), .IN2(n18780), .QN(n18778) );
  INVX0 U19780 ( .INP(n18781), .ZN(n18780) );
  NAND2X0 U19781 ( .IN1(g1312), .IN2(n18241), .QN(n18781) );
  NOR2X0 U19782 ( .IN1(n17903), .IN2(n18782), .QN(n18779) );
  NOR2X0 U19783 ( .IN1(n18783), .IN2(n18784), .QN(n18782) );
  NOR2X0 U19784 ( .IN1(n4896), .IN2(g1351), .QN(n18784) );
  NAND2X0 U19785 ( .IN1(n18785), .IN2(n18786), .QN(n4896) );
  NOR2X0 U19786 ( .IN1(n10249), .IN2(n10229), .QN(n18786) );
  NOR2X0 U19787 ( .IN1(n10190), .IN2(n17899), .QN(n18785) );
  NOR2X0 U19788 ( .IN1(n17902), .IN2(n17900), .QN(n18783) );
  NAND2X0 U19789 ( .IN1(n18787), .IN2(g1361), .QN(n17900) );
  NOR2X0 U19790 ( .IN1(n5322), .IN2(n10259), .QN(n18787) );
  NOR2X0 U19791 ( .IN1(n17901), .IN2(n10620), .QN(n17902) );
  INVX0 U19792 ( .INP(n16424), .ZN(n17903) );
  NAND2X0 U19793 ( .IN1(n18788), .IN2(n18789), .QN(g25630) );
  NAND2X0 U19794 ( .IN1(n18790), .IN2(g1249), .QN(n18789) );
  NAND2X0 U19795 ( .IN1(n18791), .IN2(n10946), .QN(n18790) );
  INVX0 U19796 ( .INP(n18792), .ZN(n18791) );
  NOR2X0 U19797 ( .IN1(g1266), .IN2(n5655), .QN(n18792) );
  NAND2X0 U19798 ( .IN1(g24247), .IN2(g1266), .QN(n18788) );
  NAND2X0 U19799 ( .IN1(n18793), .IN2(n18794), .QN(g25629) );
  NAND2X0 U19800 ( .IN1(n11063), .IN2(g1221), .QN(n18794) );
  NAND2X0 U19801 ( .IN1(n18795), .IN2(n10947), .QN(n18793) );
  NAND2X0 U19802 ( .IN1(n18796), .IN2(n18797), .QN(n18795) );
  NAND2X0 U19803 ( .IN1(n18798), .IN2(g1216), .QN(n18797) );
  NAND2X0 U19804 ( .IN1(n18799), .IN2(n5442), .QN(n18796) );
  NOR2X0 U19805 ( .IN1(test_so76), .IN2(n18798), .QN(n18799) );
  NAND2X0 U19806 ( .IN1(n18800), .IN2(n18801), .QN(g25628) );
  NAND2X0 U19807 ( .IN1(n18802), .IN2(test_so76), .QN(n18801) );
  NOR2X0 U19808 ( .IN1(n11047), .IN2(n18803), .QN(n18802) );
  NAND2X0 U19809 ( .IN1(n18804), .IN2(g1216), .QN(n18800) );
  NAND2X0 U19810 ( .IN1(n18805), .IN2(n10947), .QN(n18804) );
  NAND2X0 U19811 ( .IN1(n18803), .IN2(n10673), .QN(n18805) );
  INVX0 U19812 ( .INP(n18798), .ZN(n18803) );
  NAND2X0 U19813 ( .IN1(n18806), .IN2(n18807), .QN(g25627) );
  NAND2X0 U19814 ( .IN1(n11063), .IN2(g1178), .QN(n18807) );
  NAND2X0 U19815 ( .IN1(n18808), .IN2(n10947), .QN(n18806) );
  NAND2X0 U19816 ( .IN1(n18809), .IN2(n18810), .QN(n18808) );
  NAND2X0 U19817 ( .IN1(n18811), .IN2(g996), .QN(n18810) );
  INVX0 U19818 ( .INP(n18812), .ZN(n18811) );
  NAND2X0 U19819 ( .IN1(n18812), .IN2(g962), .QN(n18809) );
  NAND2X0 U19820 ( .IN1(n13992), .IN2(g7916), .QN(n18812) );
  NOR2X0 U19821 ( .IN1(n5599), .IN2(n5363), .QN(n13992) );
  NAND2X0 U19822 ( .IN1(n18813), .IN2(n18814), .QN(g25626) );
  NAND2X0 U19823 ( .IN1(n18815), .IN2(g1141), .QN(n18814) );
  NAND2X0 U19824 ( .IN1(n18816), .IN2(n10948), .QN(n18815) );
  NAND2X0 U19825 ( .IN1(n18817), .IN2(n18284), .QN(n18816) );
  NOR2X0 U19826 ( .IN1(g956), .IN2(n18818), .QN(n18817) );
  NAND2X0 U19827 ( .IN1(n18819), .IN2(g956), .QN(n18813) );
  NAND2X0 U19828 ( .IN1(n18820), .IN2(n18821), .QN(n18819) );
  NAND2X0 U19829 ( .IN1(n18822), .IN2(n10948), .QN(n18821) );
  NAND2X0 U19830 ( .IN1(n18284), .IN2(g1141), .QN(n18822) );
  INVX0 U19831 ( .INP(n18275), .ZN(n18284) );
  NAND2X0 U19832 ( .IN1(n5618), .IN2(test_so7), .QN(n18275) );
  NOR2X0 U19833 ( .IN1(g979), .IN2(n18823), .QN(g25625) );
  NAND2X0 U19834 ( .IN1(n18824), .IN2(n18289), .QN(n18823) );
  NAND2X0 U19835 ( .IN1(n18825), .IN2(n18826), .QN(n18289) );
  NOR2X0 U19836 ( .IN1(n5654), .IN2(n10579), .QN(n18825) );
  NAND2X0 U19837 ( .IN1(n18827), .IN2(n18828), .QN(n18824) );
  NAND2X0 U19838 ( .IN1(n14152), .IN2(n18826), .QN(n18828) );
  NAND2X0 U19839 ( .IN1(n10930), .IN2(g1052), .QN(n18827) );
  NAND2X0 U19840 ( .IN1(n18829), .IN2(n18830), .QN(g25624) );
  NAND2X0 U19841 ( .IN1(n18831), .IN2(n18292), .QN(n18830) );
  NOR2X0 U19842 ( .IN1(g1041), .IN2(n18297), .QN(n18831) );
  NOR2X0 U19843 ( .IN1(n18832), .IN2(n18833), .QN(n18829) );
  NOR2X0 U19844 ( .IN1(n10191), .IN2(n10884), .QN(n18833) );
  NOR2X0 U19845 ( .IN1(n11047), .IN2(n18834), .QN(n18832) );
  NAND2X0 U19846 ( .IN1(n18297), .IN2(g1041), .QN(n18834) );
  NAND2X0 U19847 ( .IN1(n18835), .IN2(n18836), .QN(g25623) );
  NAND2X0 U19848 ( .IN1(test_so20), .IN2(n18837), .QN(n18836) );
  NAND2X0 U19849 ( .IN1(n18297), .IN2(n10948), .QN(n18837) );
  NAND2X0 U19850 ( .IN1(n18292), .IN2(n18838), .QN(n18835) );
  NAND2X0 U19851 ( .IN1(n16468), .IN2(n18839), .QN(n18838) );
  NAND2X0 U19852 ( .IN1(n18840), .IN2(n18841), .QN(n18839) );
  INVX0 U19853 ( .INP(n17924), .ZN(n18841) );
  NAND2X0 U19854 ( .IN1(g1030), .IN2(g1018), .QN(n18840) );
  NOR2X0 U19855 ( .IN1(n11047), .IN2(n5321), .QN(n18292) );
  NOR2X0 U19856 ( .IN1(n11047), .IN2(n18842), .QN(g25622) );
  NOR2X0 U19857 ( .IN1(n18843), .IN2(n18844), .QN(n18842) );
  INVX0 U19858 ( .INP(n18845), .ZN(n18844) );
  NAND2X0 U19859 ( .IN1(n18297), .IN2(test_so20), .QN(n18845) );
  NOR2X0 U19860 ( .IN1(n17925), .IN2(n18846), .QN(n18843) );
  NOR2X0 U19861 ( .IN1(n18847), .IN2(n18848), .QN(n18846) );
  NOR2X0 U19862 ( .IN1(n4921), .IN2(g1008), .QN(n18848) );
  NAND2X0 U19863 ( .IN1(n18849), .IN2(n18850), .QN(n4921) );
  NOR2X0 U19864 ( .IN1(n10250), .IN2(n10230), .QN(n18850) );
  NOR2X0 U19865 ( .IN1(n10191), .IN2(n17923), .QN(n18849) );
  NOR2X0 U19866 ( .IN1(n17924), .IN2(n17922), .QN(n18847) );
  NAND2X0 U19867 ( .IN1(n18851), .IN2(g1018), .QN(n17922) );
  NOR2X0 U19868 ( .IN1(n5321), .IN2(n10261), .QN(n18851) );
  NOR2X0 U19869 ( .IN1(n17921), .IN2(n10619), .QN(n17924) );
  INVX0 U19870 ( .INP(n17923), .ZN(n17921) );
  INVX0 U19871 ( .INP(n16468), .ZN(n17925) );
  NAND2X0 U19872 ( .IN1(n18852), .IN2(n18853), .QN(g25621) );
  INVX0 U19873 ( .INP(n18854), .ZN(n18853) );
  NOR2X0 U19874 ( .IN1(n18855), .IN2(n10240), .QN(n18854) );
  NOR2X0 U19875 ( .IN1(n18856), .IN2(n11020), .QN(n18855) );
  NOR2X0 U19876 ( .IN1(g921), .IN2(n5654), .QN(n18856) );
  NAND2X0 U19877 ( .IN1(g24231), .IN2(g921), .QN(n18852) );
  NOR2X0 U19878 ( .IN1(n5562), .IN2(n18857), .QN(g25619) );
  NOR2X0 U19879 ( .IN1(n11048), .IN2(n18858), .QN(n18857) );
  XOR2X1 U19880 ( .IN1(n18359), .IN2(g843), .Q(n18858) );
  NAND2X0 U19881 ( .IN1(n18859), .IN2(n18860), .QN(g25618) );
  NAND2X0 U19882 ( .IN1(n18861), .IN2(g832), .QN(n18860) );
  NAND2X0 U19883 ( .IN1(n18862), .IN2(n18863), .QN(n18861) );
  NAND2X0 U19884 ( .IN1(n17170), .IN2(n17117), .QN(n18863) );
  NAND2X0 U19885 ( .IN1(n5822), .IN2(n4518), .QN(n18862) );
  NOR2X0 U19886 ( .IN1(n18864), .IN2(n11020), .QN(n4518) );
  NAND2X0 U19887 ( .IN1(n18865), .IN2(g817), .QN(n18859) );
  NAND2X0 U19888 ( .IN1(n18866), .IN2(n10948), .QN(n18865) );
  NAND2X0 U19889 ( .IN1(n18867), .IN2(n10544), .QN(n18866) );
  NOR2X0 U19890 ( .IN1(n18864), .IN2(n17177), .QN(n18867) );
  INVX0 U19891 ( .INP(n17117), .ZN(n18864) );
  NAND2X0 U19892 ( .IN1(n18868), .IN2(n18869), .QN(g25617) );
  NAND2X0 U19893 ( .IN1(n18870), .IN2(n17117), .QN(n18869) );
  NAND2X0 U19894 ( .IN1(g847), .IN2(n18871), .QN(n17117) );
  NAND2X0 U19895 ( .IN1(n5733), .IN2(g837), .QN(n18871) );
  NOR2X0 U19896 ( .IN1(n18872), .IN2(n18873), .QN(n18870) );
  NOR2X0 U19897 ( .IN1(n5822), .IN2(n17170), .QN(n18873) );
  NOR2X0 U19898 ( .IN1(n17174), .IN2(g817), .QN(n18872) );
  NAND2X0 U19899 ( .IN1(n11063), .IN2(g812), .QN(n18868) );
  NOR2X0 U19900 ( .IN1(n11048), .IN2(n18874), .QN(g25616) );
  NOR2X0 U19901 ( .IN1(n18875), .IN2(n18876), .QN(n18874) );
  NAND2X0 U19902 ( .IN1(n18877), .IN2(n18878), .QN(n18876) );
  NAND2X0 U19903 ( .IN1(n18879), .IN2(g732), .QN(n18878) );
  NOR2X0 U19904 ( .IN1(n18364), .IN2(n18880), .QN(n18879) );
  INVX0 U19905 ( .INP(n17130), .ZN(n18364) );
  NAND2X0 U19906 ( .IN1(n18880), .IN2(n5732), .QN(n18877) );
  INVX0 U19907 ( .INP(n18881), .ZN(n18880) );
  NOR2X0 U19908 ( .IN1(n17130), .IN2(n18881), .QN(n18875) );
  XNOR2X1 U19909 ( .IN1(n18882), .IN2(n18883), .Q(n18881) );
  XOR2X1 U19910 ( .IN1(n18884), .IN2(n18885), .Q(n18883) );
  XOR2X1 U19911 ( .IN1(n10400), .IN2(n10399), .Q(n18885) );
  XOR2X1 U19912 ( .IN1(n6008), .IN2(n5597), .Q(n18884) );
  XOR2X1 U19913 ( .IN1(g255), .IN2(n18886), .Q(n18882) );
  XOR2X1 U19914 ( .IN1(n10277), .IN2(n10276), .Q(n18886) );
  NAND2X0 U19915 ( .IN1(n18887), .IN2(n18888), .QN(n17130) );
  NOR2X0 U19916 ( .IN1(g370), .IN2(n18889), .QN(n18888) );
  NAND2X0 U19917 ( .IN1(n17986), .IN2(n18890), .QN(n18889) );
  NOR2X0 U19918 ( .IN1(g518), .IN2(test_so54), .QN(n17986) );
  NOR2X0 U19919 ( .IN1(g482), .IN2(n18891), .QN(n18887) );
  NAND2X0 U19920 ( .IN1(n5708), .IN2(n5327), .QN(n18891) );
  NAND2X0 U19921 ( .IN1(n18892), .IN2(n18893), .QN(g25615) );
  NAND2X0 U19922 ( .IN1(n18894), .IN2(g667), .QN(n18893) );
  NAND2X0 U19923 ( .IN1(n17973), .IN2(g686), .QN(n18892) );
  NAND2X0 U19924 ( .IN1(n18895), .IN2(n18896), .QN(g25614) );
  NAND2X0 U19925 ( .IN1(n11063), .IN2(g691), .QN(n18896) );
  NOR2X0 U19926 ( .IN1(n18897), .IN2(n18898), .QN(n18895) );
  NOR2X0 U19927 ( .IN1(n17999), .IN2(n18899), .QN(n18898) );
  INVX0 U19928 ( .INP(n5111), .ZN(n18899) );
  NOR2X0 U19929 ( .IN1(n10141), .IN2(n17973), .QN(n18897) );
  NAND2X0 U19930 ( .IN1(n18900), .IN2(n18901), .QN(g25613) );
  NAND2X0 U19931 ( .IN1(n11062), .IN2(g559), .QN(n18901) );
  NAND2X0 U19932 ( .IN1(n18902), .IN2(n18903), .QN(n18900) );
  XOR2X1 U19933 ( .IN1(n10098), .IN2(n18380), .Q(n18903) );
  NAND2X0 U19934 ( .IN1(g29211), .IN2(n18904), .QN(n18380) );
  NAND2X0 U19935 ( .IN1(n10088), .IN2(g12368), .QN(n18904) );
  NOR2X0 U19936 ( .IN1(n18905), .IN2(n18906), .QN(n18902) );
  INVX0 U19937 ( .INP(n2421), .ZN(n18906) );
  NOR2X0 U19938 ( .IN1(n19409), .IN2(n5288), .QN(n18905) );
  NAND2X0 U19939 ( .IN1(n18907), .IN2(n18908), .QN(g25612) );
  NAND2X0 U19940 ( .IN1(n18909), .IN2(g513), .QN(n18908) );
  NAND2X0 U19941 ( .IN1(n18894), .IN2(g518), .QN(n18907) );
  NAND2X0 U19942 ( .IN1(n18910), .IN2(n18911), .QN(g25611) );
  NAND2X0 U19943 ( .IN1(n18909), .IN2(g504), .QN(n18911) );
  NAND2X0 U19944 ( .IN1(n18912), .IN2(n10948), .QN(n18909) );
  NAND2X0 U19945 ( .IN1(n18913), .IN2(n17997), .QN(n18912) );
  INVX0 U19946 ( .INP(n4962), .ZN(n17997) );
  NAND2X0 U19947 ( .IN1(n18894), .IN2(g513), .QN(n18910) );
  NAND2X0 U19948 ( .IN1(n18914), .IN2(n18915), .QN(g25610) );
  NOR2X0 U19949 ( .IN1(n18916), .IN2(n18917), .QN(n18914) );
  NOR2X0 U19950 ( .IN1(n18894), .IN2(n10649), .QN(n18917) );
  NOR2X0 U19951 ( .IN1(n5519), .IN2(n17973), .QN(n18916) );
  NAND2X0 U19952 ( .IN1(n18918), .IN2(n18919), .QN(g25609) );
  NAND2X0 U19953 ( .IN1(n18920), .IN2(n5287), .QN(n18919) );
  NOR2X0 U19954 ( .IN1(n18921), .IN2(n18922), .QN(n18918) );
  NOR2X0 U19955 ( .IN1(n18923), .IN2(n10649), .QN(n18922) );
  NOR2X0 U19956 ( .IN1(n18924), .IN2(n18894), .QN(n18923) );
  INVX0 U19957 ( .INP(n17973), .ZN(n18894) );
  NAND2X0 U19958 ( .IN1(n17999), .IN2(n10949), .QN(n17973) );
  NOR2X0 U19959 ( .IN1(n11049), .IN2(g513), .QN(n18924) );
  INVX0 U19960 ( .INP(n18915), .ZN(n18921) );
  NAND2X0 U19961 ( .IN1(n4962), .IN2(n18920), .QN(n18915) );
  INVX0 U19962 ( .INP(n17963), .ZN(n18920) );
  NAND2X0 U19963 ( .IN1(n18913), .IN2(n10949), .QN(n17963) );
  INVX0 U19964 ( .INP(n17999), .ZN(n18913) );
  NAND2X0 U19965 ( .IN1(n18925), .IN2(n5633), .QN(n17999) );
  NOR2X0 U19966 ( .IN1(n5632), .IN2(n10279), .QN(n18925) );
  NAND2X0 U19967 ( .IN1(n18926), .IN2(n18927), .QN(g25605) );
  NAND2X0 U19968 ( .IN1(n11062), .IN2(g168), .QN(n18927) );
  NOR2X0 U19969 ( .IN1(n18928), .IN2(n18929), .QN(n18926) );
  NOR2X0 U19970 ( .IN1(n10167), .IN2(n11447), .QN(n18929) );
  NOR2X0 U19971 ( .IN1(n18930), .IN2(n18931), .QN(n18928) );
  NAND2X0 U19972 ( .IN1(n18890), .IN2(g246), .QN(n18931) );
  NAND2X0 U19973 ( .IN1(n18932), .IN2(n18933), .QN(g25602) );
  NAND2X0 U19974 ( .IN1(n11062), .IN2(g405), .QN(n18933) );
  NOR2X0 U19975 ( .IN1(n18934), .IN2(n18935), .QN(n18932) );
  NOR2X0 U19976 ( .IN1(n10672), .IN2(n11447), .QN(n18935) );
  NOR2X0 U19977 ( .IN1(n18930), .IN2(n18936), .QN(n18934) );
  NAND2X0 U19978 ( .IN1(n18890), .IN2(g446), .QN(n18936) );
  NAND2X0 U19979 ( .IN1(n18937), .IN2(n18938), .QN(g25601) );
  NAND2X0 U19980 ( .IN1(n11448), .IN2(g174), .QN(n18938) );
  NAND2X0 U19981 ( .IN1(test_so72), .IN2(n11447), .QN(n18937) );
  NAND2X0 U19982 ( .IN1(n18939), .IN2(n18940), .QN(g25600) );
  NAND2X0 U19983 ( .IN1(n11448), .IN2(g168), .QN(n18940) );
  INVX0 U19984 ( .INP(n11447), .ZN(n11448) );
  NAND2X0 U19985 ( .IN1(n11447), .IN2(g174), .QN(n18939) );
  NAND2X0 U19986 ( .IN1(n18941), .IN2(n10949), .QN(n11447) );
  NAND2X0 U19987 ( .IN1(n10610), .IN2(n18890), .QN(n18941) );
  INVX0 U19988 ( .INP(n1192), .ZN(n18890) );
  NAND2X0 U19989 ( .IN1(n12407), .IN2(n18942), .QN(g25599) );
  NAND2X0 U19990 ( .IN1(n11062), .IN2(g385), .QN(n18942) );
  NAND2X0 U19991 ( .IN1(n18943), .IN2(n18944), .QN(g25598) );
  NAND2X0 U19992 ( .IN1(n18945), .IN2(n1192), .QN(n18944) );
  NOR2X0 U19993 ( .IN1(n5632), .IN2(n11016), .QN(n18945) );
  NAND2X0 U19994 ( .IN1(n18946), .IN2(g376), .QN(n18943) );
  NAND2X0 U19995 ( .IN1(n18947), .IN2(n10949), .QN(n18946) );
  NAND2X0 U19996 ( .IN1(n1192), .IN2(g358), .QN(n18947) );
  NAND2X0 U19997 ( .IN1(n18948), .IN2(g358), .QN(n1192) );
  NAND2X0 U19998 ( .IN1(n18949), .IN2(n18950), .QN(g25597) );
  INVX0 U19999 ( .INP(n18951), .ZN(n18950) );
  NOR2X0 U20000 ( .IN1(n12407), .IN2(n18930), .QN(n18951) );
  NAND2X0 U20001 ( .IN1(n10610), .IN2(n10949), .QN(n18930) );
  NOR2X0 U20002 ( .IN1(n18952), .IN2(n18953), .QN(n18949) );
  NOR2X0 U20003 ( .IN1(n10279), .IN2(n10883), .QN(n18953) );
  NOR2X0 U20004 ( .IN1(n11049), .IN2(n18954), .QN(n18952) );
  NAND2X0 U20005 ( .IN1(n12407), .IN2(g370), .QN(n18954) );
  NAND2X0 U20006 ( .IN1(n18948), .IN2(g8719), .QN(n12407) );
  NOR2X0 U20007 ( .IN1(n5633), .IN2(n5632), .QN(n18948) );
  NAND2X0 U20008 ( .IN1(n18955), .IN2(n18956), .QN(g25596) );
  NAND2X0 U20009 ( .IN1(n11062), .IN2(g370), .QN(n18956) );
  NAND2X0 U20010 ( .IN1(n18957), .IN2(n10949), .QN(n18955) );
  XOR2X1 U20011 ( .IN1(n5633), .IN2(n10279), .Q(n18957) );
  NOR2X0 U20012 ( .IN1(g8719), .IN2(n18958), .QN(g25595) );
  NAND2X0 U20013 ( .IN1(n10279), .IN2(n10949), .QN(n18958) );
  NOR2X0 U20014 ( .IN1(n18959), .IN2(n18960), .QN(g25594) );
  NAND2X0 U20015 ( .IN1(n14960), .IN2(n10949), .QN(n18960) );
  NAND2X0 U20016 ( .IN1(n5627), .IN2(n18961), .QN(n14960) );
  NAND2X0 U20017 ( .IN1(n18962), .IN2(n18963), .QN(n18961) );
  NOR2X0 U20018 ( .IN1(n18964), .IN2(n18965), .QN(n18963) );
  NAND2X0 U20019 ( .IN1(n10399), .IN2(g255), .QN(n18965) );
  NAND2X0 U20020 ( .IN1(g262), .IN2(g269), .QN(n18964) );
  NOR2X0 U20021 ( .IN1(g246), .IN2(n18966), .QN(n18962) );
  NAND2X0 U20022 ( .IN1(n5597), .IN2(n10400), .QN(n18966) );
  INVX0 U20023 ( .INP(n14963), .ZN(n18959) );
  NAND2X0 U20024 ( .IN1(n18967), .IN2(n18968), .QN(n14963) );
  NOR2X0 U20025 ( .IN1(n18969), .IN2(n18970), .QN(n18968) );
  NAND2X0 U20026 ( .IN1(g232), .IN2(g239), .QN(n18970) );
  NAND2X0 U20027 ( .IN1(g225), .IN2(g246), .QN(n18969) );
  NOR2X0 U20028 ( .IN1(g269), .IN2(n18971), .QN(n18967) );
  NAND2X0 U20029 ( .IN1(n10276), .IN2(n10275), .QN(n18971) );
  NAND2X0 U20030 ( .IN1(n18972), .IN2(n18973), .QN(g25593) );
  NAND2X0 U20031 ( .IN1(n11062), .IN2(g191), .QN(n18973) );
  NAND2X0 U20032 ( .IN1(n18974), .IN2(n10950), .QN(n18972) );
  NAND2X0 U20033 ( .IN1(n18975), .IN2(n18976), .QN(n18974) );
  NAND2X0 U20034 ( .IN1(n18977), .IN2(g209), .QN(n18976) );
  NAND2X0 U20035 ( .IN1(n18978), .IN2(n18979), .QN(n18975) );
  INVX0 U20036 ( .INP(n18977), .ZN(n18979) );
  NAND2X0 U20037 ( .IN1(n18980), .IN2(n18981), .QN(g25592) );
  NAND2X0 U20038 ( .IN1(n11062), .IN2(g222), .QN(n18981) );
  NAND2X0 U20039 ( .IN1(n18982), .IN2(n10950), .QN(n18980) );
  XNOR2X1 U20040 ( .IN1(n10256), .IN2(n18983), .Q(n18982) );
  NOR2X0 U20041 ( .IN1(n18977), .IN2(n18978), .QN(n18983) );
  XOR2X1 U20042 ( .IN1(n10256), .IN2(n10257), .Q(n18978) );
  NAND2X0 U20043 ( .IN1(test_so42), .IN2(g218), .QN(n18977) );
  NAND2X0 U20044 ( .IN1(n18984), .IN2(n18985), .QN(g25591) );
  NAND2X0 U20045 ( .IN1(n10537), .IN2(n10950), .QN(n18985) );
  NAND2X0 U20046 ( .IN1(n11062), .IN2(g209), .QN(n18984) );
  NOR2X0 U20047 ( .IN1(g1657), .IN2(n10638), .QN(g25167) );
  NOR2X0 U20048 ( .IN1(n10524), .IN2(n18986), .QN(g24355) );
  NOR2X0 U20049 ( .IN1(n11049), .IN2(n18987), .QN(n18986) );
  NAND2X0 U20050 ( .IN1(n18988), .IN2(n18989), .QN(g24354) );
  NAND2X0 U20051 ( .IN1(n11062), .IN2(g6727), .QN(n18989) );
  INVX0 U20052 ( .INP(n18990), .ZN(n18988) );
  NOR2X0 U20053 ( .IN1(n18991), .IN2(n11015), .QN(n18990) );
  NAND2X0 U20054 ( .IN1(n18987), .IN2(n10523), .QN(n18991) );
  NAND2X0 U20055 ( .IN1(n18992), .IN2(g6727), .QN(n18987) );
  NAND2X0 U20056 ( .IN1(n18993), .IN2(n18994), .QN(g24353) );
  NAND2X0 U20057 ( .IN1(n11062), .IN2(g6723), .QN(n18994) );
  NAND2X0 U20058 ( .IN1(n18995), .IN2(n10950), .QN(n18993) );
  XOR2X1 U20059 ( .IN1(n18992), .IN2(g6727), .Q(n18995) );
  NOR2X0 U20060 ( .IN1(n18996), .IN2(n18997), .QN(n18992) );
  NAND2X0 U20061 ( .IN1(g14828), .IN2(g17778), .QN(n18997) );
  NAND2X0 U20062 ( .IN1(g17688), .IN2(test_so80), .QN(n18996) );
  NOR2X0 U20063 ( .IN1(n18998), .IN2(n18999), .QN(g24352) );
  NAND2X0 U20064 ( .IN1(n19000), .IN2(n10511), .QN(n18999) );
  NOR2X0 U20065 ( .IN1(n19001), .IN2(n19002), .QN(n19000) );
  NOR2X0 U20066 ( .IN1(n10381), .IN2(g14828), .QN(n19002) );
  NOR2X0 U20067 ( .IN1(test_so80), .IN2(n5700), .QN(n19001) );
  NAND2X0 U20068 ( .IN1(n19003), .IN2(n10482), .QN(n18998) );
  NOR2X0 U20069 ( .IN1(n11049), .IN2(g17688), .QN(n19003) );
  NOR2X0 U20070 ( .IN1(n10390), .IN2(n19004), .QN(g24351) );
  NOR2X0 U20071 ( .IN1(n11049), .IN2(n19005), .QN(n19004) );
  INVX0 U20072 ( .INP(n19006), .ZN(n19005) );
  NAND2X0 U20073 ( .IN1(n19007), .IN2(n19008), .QN(g24350) );
  NAND2X0 U20074 ( .IN1(test_so69), .IN2(n11080), .QN(n19008) );
  NAND2X0 U20075 ( .IN1(n19009), .IN2(n10950), .QN(n19007) );
  NOR2X0 U20076 ( .IN1(n19006), .IN2(g6390), .QN(n19009) );
  NOR2X0 U20077 ( .IN1(n19010), .IN2(n10642), .QN(n19006) );
  NAND2X0 U20078 ( .IN1(n19011), .IN2(n19012), .QN(g24349) );
  NAND2X0 U20079 ( .IN1(n11062), .IN2(g6377), .QN(n19012) );
  NAND2X0 U20080 ( .IN1(n19013), .IN2(n10950), .QN(n19011) );
  XOR2X1 U20081 ( .IN1(n10642), .IN2(n19010), .Q(n19013) );
  NAND2X0 U20082 ( .IN1(n19014), .IN2(n19015), .QN(n19010) );
  NOR2X0 U20083 ( .IN1(n5703), .IN2(n5437), .QN(n19015) );
  NOR2X0 U20084 ( .IN1(n10385), .IN2(n10370), .QN(n19014) );
  NOR2X0 U20085 ( .IN1(n19016), .IN2(n19017), .QN(g24348) );
  NAND2X0 U20086 ( .IN1(n19018), .IN2(n10519), .QN(n19017) );
  NOR2X0 U20087 ( .IN1(n19019), .IN2(n19020), .QN(n19018) );
  NOR2X0 U20088 ( .IN1(n10385), .IN2(g14779), .QN(n19020) );
  NOR2X0 U20089 ( .IN1(n5703), .IN2(g12422), .QN(n19019) );
  NAND2X0 U20090 ( .IN1(n19021), .IN2(n10492), .QN(n19016) );
  NOR2X0 U20091 ( .IN1(n11049), .IN2(g17649), .QN(n19021) );
  NOR2X0 U20092 ( .IN1(n10391), .IN2(n19022), .QN(g24347) );
  NOR2X0 U20093 ( .IN1(n11049), .IN2(n19023), .QN(n19022) );
  INVX0 U20094 ( .INP(n19024), .ZN(n19023) );
  NAND2X0 U20095 ( .IN1(n19025), .IN2(n19026), .QN(g24346) );
  NAND2X0 U20096 ( .IN1(n11061), .IN2(g6035), .QN(n19026) );
  NAND2X0 U20097 ( .IN1(n19027), .IN2(n10950), .QN(n19025) );
  NOR2X0 U20098 ( .IN1(test_so50), .IN2(n19024), .QN(n19027) );
  NOR2X0 U20099 ( .IN1(n19028), .IN2(n5528), .QN(n19024) );
  NAND2X0 U20100 ( .IN1(n19029), .IN2(n19030), .QN(g24345) );
  NAND2X0 U20101 ( .IN1(n11061), .IN2(g6031), .QN(n19030) );
  NAND2X0 U20102 ( .IN1(n19031), .IN2(n10950), .QN(n19029) );
  XOR2X1 U20103 ( .IN1(n19028), .IN2(n5528), .Q(n19031) );
  NAND2X0 U20104 ( .IN1(n19032), .IN2(n19033), .QN(n19028) );
  NOR2X0 U20105 ( .IN1(n5698), .IN2(n5432), .QN(n19033) );
  NOR2X0 U20106 ( .IN1(n10376), .IN2(n10361), .QN(n19032) );
  NOR2X0 U20107 ( .IN1(n19034), .IN2(n19035), .QN(g24344) );
  NAND2X0 U20108 ( .IN1(n19036), .IN2(n10499), .QN(n19035) );
  NOR2X0 U20109 ( .IN1(n19037), .IN2(n19038), .QN(n19036) );
  NOR2X0 U20110 ( .IN1(n10376), .IN2(g14738), .QN(n19038) );
  NOR2X0 U20111 ( .IN1(n5698), .IN2(g12350), .QN(n19037) );
  NAND2X0 U20112 ( .IN1(n19039), .IN2(n10468), .QN(n19034) );
  NOR2X0 U20113 ( .IN1(n11050), .IN2(g17607), .QN(n19039) );
  NOR2X0 U20114 ( .IN1(n10395), .IN2(n19040), .QN(g24343) );
  NOR2X0 U20115 ( .IN1(n11050), .IN2(n19041), .QN(n19040) );
  INVX0 U20116 ( .INP(n19042), .ZN(n19041) );
  NAND2X0 U20117 ( .IN1(n19043), .IN2(n19044), .QN(g24342) );
  NAND2X0 U20118 ( .IN1(n11061), .IN2(g5689), .QN(n19044) );
  NAND2X0 U20119 ( .IN1(n19045), .IN2(n10951), .QN(n19043) );
  NOR2X0 U20120 ( .IN1(n19042), .IN2(g5698), .QN(n19045) );
  NOR2X0 U20121 ( .IN1(n19046), .IN2(n5529), .QN(n19042) );
  NAND2X0 U20122 ( .IN1(n19047), .IN2(n19048), .QN(g24341) );
  NAND2X0 U20123 ( .IN1(n11061), .IN2(g5685), .QN(n19048) );
  NAND2X0 U20124 ( .IN1(n19049), .IN2(n10951), .QN(n19047) );
  XOR2X1 U20125 ( .IN1(n19046), .IN2(n5529), .Q(n19049) );
  NAND2X0 U20126 ( .IN1(n19050), .IN2(n19051), .QN(n19046) );
  NOR2X0 U20127 ( .IN1(n5705), .IN2(n5439), .QN(n19051) );
  NOR2X0 U20128 ( .IN1(n10378), .IN2(n10363), .QN(n19050) );
  NOR2X0 U20129 ( .IN1(n19052), .IN2(n19053), .QN(g24340) );
  NAND2X0 U20130 ( .IN1(n19054), .IN2(n10503), .QN(n19053) );
  NOR2X0 U20131 ( .IN1(n19055), .IN2(n19056), .QN(n19054) );
  NOR2X0 U20132 ( .IN1(n10378), .IN2(g14694), .QN(n19056) );
  NOR2X0 U20133 ( .IN1(n5705), .IN2(g12300), .QN(n19055) );
  NAND2X0 U20134 ( .IN1(n19057), .IN2(n10473), .QN(n19052) );
  NOR2X0 U20135 ( .IN1(n11050), .IN2(g17580), .QN(n19057) );
  NOR2X0 U20136 ( .IN1(n10526), .IN2(n19058), .QN(g24339) );
  NOR2X0 U20137 ( .IN1(n11050), .IN2(n19059), .QN(n19058) );
  INVX0 U20138 ( .INP(n19060), .ZN(n19059) );
  NAND2X0 U20139 ( .IN1(n19061), .IN2(n19062), .QN(g24338) );
  NAND2X0 U20140 ( .IN1(test_so10), .IN2(n11014), .QN(n19062) );
  NAND2X0 U20141 ( .IN1(n19063), .IN2(n10951), .QN(n19061) );
  NOR2X0 U20142 ( .IN1(n19060), .IN2(g5352), .QN(n19063) );
  NOR2X0 U20143 ( .IN1(n19064), .IN2(n10641), .QN(n19060) );
  NAND2X0 U20144 ( .IN1(n19065), .IN2(n19066), .QN(g24337) );
  NAND2X0 U20145 ( .IN1(n11061), .IN2(g5339), .QN(n19066) );
  NAND2X0 U20146 ( .IN1(n19067), .IN2(n10951), .QN(n19065) );
  XOR2X1 U20147 ( .IN1(n10641), .IN2(n19064), .Q(n19067) );
  NAND2X0 U20148 ( .IN1(n19068), .IN2(n19069), .QN(n19064) );
  NOR2X0 U20149 ( .IN1(n5704), .IN2(n5438), .QN(n19069) );
  NOR2X0 U20150 ( .IN1(n10374), .IN2(n10359), .QN(n19068) );
  NOR2X0 U20151 ( .IN1(n19070), .IN2(n19071), .QN(g24336) );
  NAND2X0 U20152 ( .IN1(n19072), .IN2(n10463), .QN(n19071) );
  NOR2X0 U20153 ( .IN1(n19073), .IN2(n19074), .QN(n19072) );
  NOR2X0 U20154 ( .IN1(n10374), .IN2(g14662), .QN(n19074) );
  NOR2X0 U20155 ( .IN1(n5704), .IN2(g12238), .QN(n19073) );
  NAND2X0 U20156 ( .IN1(n19075), .IN2(n10442), .QN(n19070) );
  INVX0 U20157 ( .INP(n19076), .ZN(n19075) );
  NAND2X0 U20158 ( .IN1(n10931), .IN2(n10359), .QN(n19076) );
  NAND2X0 U20159 ( .IN1(n19077), .IN2(n19078), .QN(g24335) );
  NAND2X0 U20160 ( .IN1(n19079), .IN2(n19080), .QN(n19078) );
  NOR2X0 U20161 ( .IN1(n5382), .IN2(g4340), .QN(n19079) );
  NAND2X0 U20162 ( .IN1(n11061), .IN2(g18881), .QN(n19077) );
  NAND2X0 U20163 ( .IN1(n19081), .IN2(n19082), .QN(g24334) );
  NAND2X0 U20164 ( .IN1(n19083), .IN2(n19084), .QN(n19082) );
  NOR2X0 U20165 ( .IN1(n19085), .IN2(n19086), .QN(n19084) );
  NAND2X0 U20166 ( .IN1(n5303), .IN2(n5365), .QN(n19086) );
  NAND2X0 U20167 ( .IN1(n18143), .IN2(n12260), .QN(n19085) );
  INVX0 U20168 ( .INP(n12580), .ZN(n12260) );
  NAND2X0 U20169 ( .IN1(test_so3), .IN2(n5727), .QN(n12580) );
  NOR2X0 U20170 ( .IN1(n5844), .IN2(n5653), .QN(n18143) );
  NOR2X0 U20171 ( .IN1(n19087), .IN2(n19088), .QN(n19083) );
  NAND2X0 U20172 ( .IN1(n19080), .IN2(n5608), .QN(n19088) );
  INVX0 U20173 ( .INP(n19089), .ZN(n19080) );
  NAND2X0 U20174 ( .IN1(n19090), .IN2(n19091), .QN(n19089) );
  NOR2X0 U20175 ( .IN1(g4322), .IN2(n19092), .QN(n19091) );
  NAND2X0 U20176 ( .IN1(n10931), .IN2(n10643), .QN(n19092) );
  NOR2X0 U20177 ( .IN1(g4358), .IN2(n19093), .QN(n19090) );
  NAND2X0 U20178 ( .IN1(n5323), .IN2(n5540), .QN(n19093) );
  NAND2X0 U20179 ( .IN1(n5274), .IN2(n5539), .QN(n19087) );
  NAND2X0 U20180 ( .IN1(n11061), .IN2(g4358), .QN(n19081) );
  NOR2X0 U20181 ( .IN1(n5710), .IN2(n10883), .QN(g24298) );
  NAND2X0 U20182 ( .IN1(n19094), .IN2(n19095), .QN(g24282) );
  NAND2X0 U20183 ( .IN1(n19096), .IN2(g4308), .QN(n19095) );
  NAND2X0 U20184 ( .IN1(n10931), .IN2(g9251), .QN(n19096) );
  NAND2X0 U20185 ( .IN1(g24281), .IN2(g9251), .QN(n19094) );
  NOR2X0 U20186 ( .IN1(g4308), .IN2(n11016), .QN(g24281) );
  NAND2X0 U20187 ( .IN1(n19097), .IN2(n19098), .QN(g24280) );
  NAND2X0 U20188 ( .IN1(n19099), .IN2(g4269), .QN(n19098) );
  NAND2X0 U20189 ( .IN1(n19100), .IN2(n10951), .QN(n19099) );
  NAND2X0 U20190 ( .IN1(n19101), .IN2(n5764), .QN(n19100) );
  NOR2X0 U20191 ( .IN1(n5823), .IN2(n10127), .QN(n19101) );
  NAND2X0 U20192 ( .IN1(n19102), .IN2(g4273), .QN(n19097) );
  NAND2X0 U20193 ( .IN1(n19103), .IN2(n19104), .QN(n19102) );
  NAND2X0 U20194 ( .IN1(n5763), .IN2(n10951), .QN(n19104) );
  NAND2X0 U20195 ( .IN1(n19105), .IN2(n19106), .QN(g24279) );
  NAND2X0 U20196 ( .IN1(n19107), .IN2(n19108), .QN(n19106) );
  NOR2X0 U20197 ( .IN1(n19109), .IN2(n19110), .QN(n19105) );
  NOR2X0 U20198 ( .IN1(n11050), .IN2(n19111), .QN(n19110) );
  NOR2X0 U20199 ( .IN1(n19112), .IN2(n19113), .QN(n19111) );
  NOR2X0 U20200 ( .IN1(n19114), .IN2(n19115), .QN(n19113) );
  INVX0 U20201 ( .INP(n19108), .ZN(n19114) );
  INVX0 U20202 ( .INP(n19116), .ZN(n19112) );
  NAND2X0 U20203 ( .IN1(n19115), .IN2(n19117), .QN(n19116) );
  NOR2X0 U20204 ( .IN1(n19108), .IN2(n19107), .QN(n19117) );
  NOR2X0 U20205 ( .IN1(n5726), .IN2(n10325), .QN(n19107) );
  NAND2X0 U20206 ( .IN1(n19118), .IN2(n5726), .QN(n19115) );
  NOR2X0 U20207 ( .IN1(n19119), .IN2(g4235), .QN(n19118) );
  NOR2X0 U20208 ( .IN1(n19120), .IN2(n19121), .QN(n19119) );
  NAND2X0 U20209 ( .IN1(n19122), .IN2(n19406), .QN(n19121) );
  NOR2X0 U20210 ( .IN1(g8919), .IN2(g11770), .QN(n19122) );
  NAND2X0 U20211 ( .IN1(n19123), .IN2(n19124), .QN(n19120) );
  NOR2X0 U20212 ( .IN1(g8915), .IN2(g8918), .QN(n19124) );
  NOR2X0 U20213 ( .IN1(g8917), .IN2(g8920), .QN(n19123) );
  NOR2X0 U20214 ( .IN1(n10325), .IN2(n10883), .QN(n19109) );
  NOR2X0 U20215 ( .IN1(n10397), .IN2(n19125), .QN(g24278) );
  NOR2X0 U20216 ( .IN1(n11050), .IN2(n19126), .QN(n19125) );
  INVX0 U20217 ( .INP(n19127), .ZN(n19126) );
  NAND2X0 U20218 ( .IN1(n19128), .IN2(n19129), .QN(g24277) );
  NAND2X0 U20219 ( .IN1(n11061), .IN2(g4040), .QN(n19129) );
  NAND2X0 U20220 ( .IN1(n19130), .IN2(n10951), .QN(n19128) );
  NOR2X0 U20221 ( .IN1(n19127), .IN2(g4049), .QN(n19130) );
  NOR2X0 U20222 ( .IN1(n19131), .IN2(n5530), .QN(n19127) );
  NAND2X0 U20223 ( .IN1(n19132), .IN2(n19133), .QN(g24276) );
  NAND2X0 U20224 ( .IN1(n11061), .IN2(g4031), .QN(n19133) );
  NAND2X0 U20225 ( .IN1(n19134), .IN2(n10951), .QN(n19132) );
  XOR2X1 U20226 ( .IN1(n19131), .IN2(n5530), .Q(n19134) );
  NAND2X0 U20227 ( .IN1(n19135), .IN2(n19136), .QN(n19131) );
  NOR2X0 U20228 ( .IN1(n5701), .IN2(n5435), .QN(n19136) );
  NOR2X0 U20229 ( .IN1(n10379), .IN2(n10365), .QN(n19135) );
  NOR2X0 U20230 ( .IN1(n19137), .IN2(n19138), .QN(g24275) );
  NAND2X0 U20231 ( .IN1(n19139), .IN2(n10507), .QN(n19138) );
  NOR2X0 U20232 ( .IN1(n19140), .IN2(n19141), .QN(n19139) );
  NOR2X0 U20233 ( .IN1(n10379), .IN2(g13966), .QN(n19141) );
  NOR2X0 U20234 ( .IN1(n5701), .IN2(g11418), .QN(n19140) );
  NAND2X0 U20235 ( .IN1(n19142), .IN2(n10477), .QN(n19137) );
  NOR2X0 U20236 ( .IN1(n11050), .IN2(g16659), .QN(n19142) );
  NOR2X0 U20237 ( .IN1(n10393), .IN2(n19143), .QN(g24274) );
  NOR2X0 U20238 ( .IN1(n11050), .IN2(n19144), .QN(n19143) );
  INVX0 U20239 ( .INP(n19145), .ZN(n19144) );
  NAND2X0 U20240 ( .IN1(n19146), .IN2(n19147), .QN(g24273) );
  NAND2X0 U20241 ( .IN1(n11061), .IN2(g3689), .QN(n19147) );
  NAND2X0 U20242 ( .IN1(n19148), .IN2(n10952), .QN(n19146) );
  NOR2X0 U20243 ( .IN1(n19145), .IN2(g3698), .QN(n19148) );
  NOR2X0 U20244 ( .IN1(n19149), .IN2(n5532), .QN(n19145) );
  NAND2X0 U20245 ( .IN1(n19150), .IN2(n19151), .QN(g24272) );
  NAND2X0 U20246 ( .IN1(n11060), .IN2(g3680), .QN(n19151) );
  NAND2X0 U20247 ( .IN1(n19152), .IN2(n10952), .QN(n19150) );
  XOR2X1 U20248 ( .IN1(n19149), .IN2(n5532), .Q(n19152) );
  NAND2X0 U20249 ( .IN1(n19153), .IN2(n19154), .QN(n19149) );
  NOR2X0 U20250 ( .IN1(n5699), .IN2(n5433), .QN(n19154) );
  NOR2X0 U20251 ( .IN1(n10383), .IN2(n10369), .QN(n19153) );
  NOR2X0 U20252 ( .IN1(n19155), .IN2(n19156), .QN(g24271) );
  NAND2X0 U20253 ( .IN1(n19157), .IN2(n10515), .QN(n19156) );
  NOR2X0 U20254 ( .IN1(n19158), .IN2(n19159), .QN(n19157) );
  NOR2X0 U20255 ( .IN1(n10383), .IN2(g13926), .QN(n19159) );
  NOR2X0 U20256 ( .IN1(n5699), .IN2(g11388), .QN(n19158) );
  NAND2X0 U20257 ( .IN1(n19160), .IN2(n10487), .QN(n19155) );
  NOR2X0 U20258 ( .IN1(n11050), .IN2(g16627), .QN(n19160) );
  NOR2X0 U20259 ( .IN1(n10388), .IN2(n19161), .QN(g24270) );
  NOR2X0 U20260 ( .IN1(n11050), .IN2(n19162), .QN(n19161) );
  INVX0 U20261 ( .INP(n19163), .ZN(n19162) );
  NAND2X0 U20262 ( .IN1(n19164), .IN2(n19165), .QN(g24269) );
  NAND2X0 U20263 ( .IN1(n11060), .IN2(g3338), .QN(n19165) );
  NAND2X0 U20264 ( .IN1(n19166), .IN2(n10952), .QN(n19164) );
  NOR2X0 U20265 ( .IN1(n19163), .IN2(g3347), .QN(n19166) );
  NOR2X0 U20266 ( .IN1(n19167), .IN2(n5527), .QN(n19163) );
  NAND2X0 U20267 ( .IN1(n19168), .IN2(n19169), .QN(g24268) );
  NAND2X0 U20268 ( .IN1(test_so91), .IN2(n11014), .QN(n19169) );
  NAND2X0 U20269 ( .IN1(n19170), .IN2(n10952), .QN(n19168) );
  XOR2X1 U20270 ( .IN1(n19167), .IN2(n5527), .Q(n19170) );
  NAND2X0 U20271 ( .IN1(n19171), .IN2(n19172), .QN(n19167) );
  NOR2X0 U20272 ( .IN1(n5702), .IN2(n5436), .QN(n19172) );
  NOR2X0 U20273 ( .IN1(n10372), .IN2(n10357), .QN(n19171) );
  NOR2X0 U20274 ( .IN1(n19173), .IN2(n19174), .QN(g24267) );
  NAND2X0 U20275 ( .IN1(n19175), .IN2(n10495), .QN(n19174) );
  NOR2X0 U20276 ( .IN1(n19176), .IN2(n19177), .QN(n19175) );
  NOR2X0 U20277 ( .IN1(n10372), .IN2(g13895), .QN(n19177) );
  NOR2X0 U20278 ( .IN1(n5702), .IN2(g11349), .QN(n19176) );
  NAND2X0 U20279 ( .IN1(n19178), .IN2(n10458), .QN(n19173) );
  NOR2X0 U20280 ( .IN1(n11050), .IN2(g16603), .QN(n19178) );
  NAND2X0 U20281 ( .IN1(n19179), .IN2(n19180), .QN(g24266) );
  INVX0 U20282 ( .INP(n19181), .ZN(n19180) );
  NOR2X0 U20283 ( .IN1(n10908), .IN2(n5963), .QN(n19181) );
  NAND2X0 U20284 ( .IN1(n19182), .IN2(n10952), .QN(n19179) );
  NOR2X0 U20285 ( .IN1(g2712), .IN2(n19407), .QN(n19182) );
  NAND2X0 U20286 ( .IN1(n19183), .IN2(n14448), .QN(g24263) );
  NAND2X0 U20287 ( .IN1(n5963), .IN2(n10952), .QN(n14448) );
  NOR2X0 U20288 ( .IN1(n19184), .IN2(n19185), .QN(n19183) );
  NOR2X0 U20289 ( .IN1(n10142), .IN2(n10883), .QN(n19185) );
  NOR2X0 U20290 ( .IN1(n11050), .IN2(g2715), .QN(n19184) );
  NAND2X0 U20291 ( .IN1(n19186), .IN2(n19187), .QN(g24262) );
  NAND2X0 U20292 ( .IN1(n19188), .IN2(n10545), .QN(n19187) );
  NOR2X0 U20293 ( .IN1(n19189), .IN2(n19190), .QN(n19186) );
  NOR2X0 U20294 ( .IN1(n5546), .IN2(n10883), .QN(n19190) );
  INVX0 U20295 ( .INP(n19191), .ZN(n19189) );
  NAND2X0 U20296 ( .IN1(n10931), .IN2(n19192), .QN(n19191) );
  NOR2X0 U20297 ( .IN1(n19188), .IN2(n10545), .QN(n19192) );
  NAND2X0 U20298 ( .IN1(n18763), .IN2(n19193), .QN(g24261) );
  NAND2X0 U20299 ( .IN1(n11059), .IN2(g1585), .QN(n19193) );
  XNOR2X1 U20300 ( .IN1(n19194), .IN2(n10546), .Q(g24260) );
  NOR2X0 U20301 ( .IN1(n11051), .IN2(n5546), .QN(n19194) );
  NAND2X0 U20302 ( .IN1(n18763), .IN2(n19195), .QN(g24259) );
  NAND2X0 U20303 ( .IN1(n11060), .IN2(g1579), .QN(n19195) );
  NAND2X0 U20304 ( .IN1(n19196), .IN2(n19197), .QN(g24258) );
  NAND2X0 U20305 ( .IN1(n10931), .IN2(g496), .QN(n19197) );
  NAND2X0 U20306 ( .IN1(n11059), .IN2(g1554), .QN(n19196) );
  XNOR2X1 U20307 ( .IN1(n19198), .IN2(n5616), .Q(g24257) );
  NOR2X0 U20308 ( .IN1(n19199), .IN2(n11018), .QN(n19198) );
  NAND2X0 U20309 ( .IN1(n19200), .IN2(n19201), .QN(g24256) );
  NAND2X0 U20310 ( .IN1(n11060), .IN2(g1339), .QN(n19201) );
  NAND2X0 U20311 ( .IN1(n19202), .IN2(n10952), .QN(n19200) );
  XNOR2X1 U20312 ( .IN1(n19199), .IN2(n19203), .Q(n19202) );
  NOR2X0 U20313 ( .IN1(g13272), .IN2(n19204), .QN(n19203) );
  NAND2X0 U20314 ( .IN1(n10157), .IN2(n18760), .QN(n19204) );
  NOR2X0 U20315 ( .IN1(n19205), .IN2(g19357), .QN(n18760) );
  NAND2X0 U20316 ( .IN1(n5616), .IN2(n5302), .QN(n19205) );
  NAND2X0 U20317 ( .IN1(n19206), .IN2(n19207), .QN(n19199) );
  XOR2X1 U20318 ( .IN1(g1579), .IN2(test_so68), .Q(n19207) );
  NAND2X0 U20319 ( .IN1(n19208), .IN2(n19209), .QN(g24255) );
  NAND2X0 U20320 ( .IN1(n14133), .IN2(g17423), .QN(n19209) );
  NOR2X0 U20321 ( .IN1(n19210), .IN2(n19211), .QN(n19208) );
  NOR2X0 U20322 ( .IN1(n5755), .IN2(n10882), .QN(n19211) );
  NOR2X0 U20323 ( .IN1(n11051), .IN2(n19212), .QN(n19210) );
  NAND2X0 U20324 ( .IN1(n10234), .IN2(g10527), .QN(n19212) );
  NOR2X0 U20325 ( .IN1(n19213), .IN2(n19214), .QN(g24254) );
  NAND2X0 U20326 ( .IN1(n10236), .IN2(n10235), .QN(n19214) );
  NAND2X0 U20327 ( .IN1(n19215), .IN2(n10234), .QN(n19213) );
  NOR2X0 U20328 ( .IN1(n11051), .IN2(n19216), .QN(n19215) );
  NOR2X0 U20329 ( .IN1(n18732), .IN2(n19217), .QN(n19216) );
  INVX0 U20330 ( .INP(n19218), .ZN(n19217) );
  NOR2X0 U20331 ( .IN1(n19206), .IN2(n5768), .QN(n19218) );
  NOR2X0 U20332 ( .IN1(n18241), .IN2(n4836), .QN(n19206) );
  NAND2X0 U20333 ( .IN1(n5466), .IN2(n5322), .QN(n4836) );
  NAND2X0 U20334 ( .IN1(n17899), .IN2(n16424), .QN(n18241) );
  NAND2X0 U20335 ( .IN1(n5616), .IN2(n10650), .QN(n16424) );
  INVX0 U20336 ( .INP(n17901), .ZN(n17899) );
  XNOR2X1 U20337 ( .IN1(g1339), .IN2(test_so68), .Q(n17901) );
  NAND2X0 U20338 ( .IN1(n19188), .IN2(g1564), .QN(n18732) );
  NOR2X0 U20339 ( .IN1(n5546), .IN2(n10546), .QN(n19188) );
  NAND2X0 U20340 ( .IN1(n19219), .IN2(n19220), .QN(g24253) );
  NAND2X0 U20341 ( .IN1(n11059), .IN2(g1306), .QN(n19220) );
  NAND2X0 U20342 ( .IN1(n19221), .IN2(n10953), .QN(n19219) );
  NAND2X0 U20343 ( .IN1(n19222), .IN2(n19223), .QN(n19221) );
  NAND2X0 U20344 ( .IN1(g7946), .IN2(g1521), .QN(n19223) );
  NAND2X0 U20345 ( .IN1(n5302), .IN2(g1532), .QN(n19222) );
  NAND2X0 U20346 ( .IN1(n19224), .IN2(n19225), .QN(g24252) );
  NAND2X0 U20347 ( .IN1(test_so49), .IN2(n11081), .QN(n19225) );
  NAND2X0 U20348 ( .IN1(n19226), .IN2(n10953), .QN(n19224) );
  NAND2X0 U20349 ( .IN1(n18744), .IN2(n19227), .QN(n19226) );
  NAND2X0 U20350 ( .IN1(n5302), .IN2(g1521), .QN(n19227) );
  NAND2X0 U20351 ( .IN1(g7946), .IN2(g1339), .QN(n18744) );
  NAND2X0 U20352 ( .IN1(n19228), .IN2(n19229), .QN(g24251) );
  NAND2X0 U20353 ( .IN1(n17020), .IN2(g1442), .QN(n19229) );
  NAND2X0 U20354 ( .IN1(test_so12), .IN2(n18753), .QN(n19228) );
  NAND2X0 U20355 ( .IN1(n19230), .IN2(n19231), .QN(g24250) );
  NAND2X0 U20356 ( .IN1(test_so12), .IN2(n17020), .QN(n19231) );
  NAND2X0 U20357 ( .IN1(n18753), .IN2(g1489), .QN(n19230) );
  NAND2X0 U20358 ( .IN1(n19232), .IN2(n19233), .QN(g24249) );
  NAND2X0 U20359 ( .IN1(n19234), .IN2(n17027), .QN(n19233) );
  INVX0 U20360 ( .INP(n18751), .ZN(n17027) );
  NOR2X0 U20361 ( .IN1(n11051), .IN2(g1442), .QN(n19234) );
  NAND2X0 U20362 ( .IN1(n19235), .IN2(g1489), .QN(n19232) );
  INVX0 U20363 ( .INP(n19236), .ZN(n19235) );
  NOR2X0 U20364 ( .IN1(n17020), .IN2(n19237), .QN(n19236) );
  NOR2X0 U20365 ( .IN1(n11051), .IN2(test_so12), .QN(n19237) );
  INVX0 U20366 ( .INP(n18753), .ZN(n17020) );
  NAND2X0 U20367 ( .IN1(n18751), .IN2(n10953), .QN(n18753) );
  NAND2X0 U20368 ( .IN1(n19238), .IN2(n5364), .QN(n18751) );
  NOR2X0 U20369 ( .IN1(test_so49), .IN2(n10244), .QN(n19238) );
  NAND2X0 U20370 ( .IN1(n19239), .IN2(n19240), .QN(g24248) );
  XNOR2X1 U20371 ( .IN1(n10251), .IN2(n19241), .Q(n19240) );
  NAND2X0 U20372 ( .IN1(n5655), .IN2(n10953), .QN(n19241) );
  NOR2X0 U20373 ( .IN1(n19242), .IN2(n19243), .QN(n19239) );
  NOR2X0 U20374 ( .IN1(n11051), .IN2(g19357), .QN(n19243) );
  NOR2X0 U20375 ( .IN1(n10580), .IN2(n18763), .QN(n19242) );
  NOR2X0 U20376 ( .IN1(g1249), .IN2(n18763), .QN(g24247) );
  INVX0 U20377 ( .INP(n14133), .ZN(n18763) );
  NOR2X0 U20378 ( .IN1(n11051), .IN2(n5655), .QN(n14133) );
  NAND2X0 U20379 ( .IN1(n19244), .IN2(n19245), .QN(g24246) );
  NAND2X0 U20380 ( .IN1(n19246), .IN2(n10547), .QN(n19245) );
  NOR2X0 U20381 ( .IN1(n19247), .IN2(n19248), .QN(n19244) );
  NOR2X0 U20382 ( .IN1(n5547), .IN2(n10882), .QN(n19248) );
  INVX0 U20383 ( .INP(n19249), .ZN(n19247) );
  NAND2X0 U20384 ( .IN1(n10931), .IN2(n19250), .QN(n19249) );
  NOR2X0 U20385 ( .IN1(n19246), .IN2(n10547), .QN(n19250) );
  NAND2X0 U20386 ( .IN1(n19251), .IN2(n19252), .QN(g24245) );
  NAND2X0 U20387 ( .IN1(n11058), .IN2(g30332), .QN(n19252) );
  XOR2X1 U20388 ( .IN1(n19253), .IN2(n10548), .Q(g24244) );
  NAND2X0 U20389 ( .IN1(n10931), .IN2(g1205), .QN(n19253) );
  NAND2X0 U20390 ( .IN1(n19251), .IN2(n19254), .QN(g24243) );
  NAND2X0 U20391 ( .IN1(n11059), .IN2(g1236), .QN(n19254) );
  NAND2X0 U20392 ( .IN1(n19255), .IN2(n19256), .QN(g24242) );
  NAND2X0 U20393 ( .IN1(n10932), .IN2(g29215), .QN(n19256) );
  NAND2X0 U20394 ( .IN1(test_so76), .IN2(n11014), .QN(n19255) );
  XOR2X1 U20395 ( .IN1(n19257), .IN2(n5622), .Q(g24241) );
  NAND2X0 U20396 ( .IN1(n19258), .IN2(n10953), .QN(n19257) );
  NAND2X0 U20397 ( .IN1(n19259), .IN2(n19260), .QN(g24240) );
  NAND2X0 U20398 ( .IN1(n11059), .IN2(g996), .QN(n19260) );
  NAND2X0 U20399 ( .IN1(n19261), .IN2(n10953), .QN(n19259) );
  XOR2X1 U20400 ( .IN1(n19258), .IN2(n19262), .Q(n19261) );
  NOR2X0 U20401 ( .IN1(g13259), .IN2(n19263), .QN(n19262) );
  NAND2X0 U20402 ( .IN1(n10148), .IN2(n19264), .QN(n19263) );
  INVX0 U20403 ( .INP(n18826), .ZN(n19264) );
  NAND2X0 U20404 ( .IN1(n19265), .IN2(n5392), .QN(n18826) );
  NOR2X0 U20405 ( .IN1(g990), .IN2(g7916), .QN(n19265) );
  NOR2X0 U20406 ( .IN1(n19266), .IN2(n18297), .QN(n19258) );
  NAND2X0 U20407 ( .IN1(n18004), .IN2(n19267), .QN(n19266) );
  XOR2X1 U20408 ( .IN1(n10224), .IN2(n5320), .Q(n19267) );
  NAND2X0 U20409 ( .IN1(n19268), .IN2(n19269), .QN(g24239) );
  NAND2X0 U20410 ( .IN1(n14152), .IN2(g17400), .QN(n19269) );
  NOR2X0 U20411 ( .IN1(n19270), .IN2(n19271), .QN(n19268) );
  NOR2X0 U20412 ( .IN1(n5756), .IN2(n10882), .QN(n19271) );
  NOR2X0 U20413 ( .IN1(n11051), .IN2(n19272), .QN(n19270) );
  NAND2X0 U20414 ( .IN1(n10227), .IN2(g10500), .QN(n19272) );
  NOR2X0 U20415 ( .IN1(n19273), .IN2(n19274), .QN(g24238) );
  NAND2X0 U20416 ( .IN1(n10218), .IN2(n10227), .QN(n19274) );
  NAND2X0 U20417 ( .IN1(n19275), .IN2(n19276), .QN(n19273) );
  NAND2X0 U20418 ( .IN1(n19277), .IN2(test_so76), .QN(n19276) );
  NOR2X0 U20419 ( .IN1(n19278), .IN2(n18798), .QN(n19277) );
  NAND2X0 U20420 ( .IN1(n19246), .IN2(g1221), .QN(n18798) );
  NOR2X0 U20421 ( .IN1(n5547), .IN2(n10548), .QN(n19246) );
  NOR2X0 U20422 ( .IN1(n4837), .IN2(n18297), .QN(n19278) );
  NAND2X0 U20423 ( .IN1(n17923), .IN2(n16468), .QN(n18297) );
  NAND2X0 U20424 ( .IN1(n5622), .IN2(n5320), .QN(n16468) );
  XNOR2X1 U20425 ( .IN1(g996), .IN2(n5320), .Q(n17923) );
  INVX0 U20426 ( .INP(n18004), .ZN(n4837) );
  NOR2X0 U20427 ( .IN1(g1008), .IN2(test_so20), .QN(n18004) );
  NOR2X0 U20428 ( .IN1(test_so44), .IN2(n11020), .QN(n19275) );
  NAND2X0 U20429 ( .IN1(n19279), .IN2(n19280), .QN(g24237) );
  NAND2X0 U20430 ( .IN1(n11059), .IN2(g962), .QN(n19280) );
  NAND2X0 U20431 ( .IN1(n19281), .IN2(n10953), .QN(n19279) );
  NAND2X0 U20432 ( .IN1(n19282), .IN2(n19283), .QN(n19281) );
  NAND2X0 U20433 ( .IN1(n5304), .IN2(g1189), .QN(n19283) );
  NAND2X0 U20434 ( .IN1(g1178), .IN2(g7916), .QN(n19282) );
  NAND2X0 U20435 ( .IN1(n19284), .IN2(n19285), .QN(g24236) );
  NAND2X0 U20436 ( .IN1(n11059), .IN2(g1183), .QN(n19285) );
  NAND2X0 U20437 ( .IN1(n19286), .IN2(n10953), .QN(n19284) );
  NAND2X0 U20438 ( .IN1(n19287), .IN2(n19288), .QN(n19286) );
  NAND2X0 U20439 ( .IN1(g996), .IN2(g7916), .QN(n19288) );
  NAND2X0 U20440 ( .IN1(n5304), .IN2(g1178), .QN(n19287) );
  NAND2X0 U20441 ( .IN1(n19289), .IN2(n19290), .QN(g24235) );
  NAND2X0 U20442 ( .IN1(test_so7), .IN2(n17073), .QN(n19290) );
  NAND2X0 U20443 ( .IN1(n18820), .IN2(g1152), .QN(n19289) );
  NAND2X0 U20444 ( .IN1(n19291), .IN2(n19292), .QN(g24234) );
  NAND2X0 U20445 ( .IN1(n17073), .IN2(g1152), .QN(n19292) );
  INVX0 U20446 ( .INP(n18820), .ZN(n17073) );
  NAND2X0 U20447 ( .IN1(n18820), .IN2(g1146), .QN(n19291) );
  NAND2X0 U20448 ( .IN1(n19293), .IN2(n19294), .QN(g24233) );
  NAND2X0 U20449 ( .IN1(n17098), .IN2(n17081), .QN(n19294) );
  INVX0 U20450 ( .INP(n18818), .ZN(n17081) );
  NOR2X0 U20451 ( .IN1(test_so7), .IN2(n11020), .QN(n17098) );
  NAND2X0 U20452 ( .IN1(n19295), .IN2(g1146), .QN(n19293) );
  NAND2X0 U20453 ( .IN1(n18820), .IN2(n19296), .QN(n19295) );
  NAND2X0 U20454 ( .IN1(n5618), .IN2(n10954), .QN(n19296) );
  NAND2X0 U20455 ( .IN1(n18818), .IN2(n10954), .QN(n18820) );
  NAND2X0 U20456 ( .IN1(n19297), .IN2(n5599), .QN(n18818) );
  NOR2X0 U20457 ( .IN1(n10243), .IN2(g1171), .QN(n19297) );
  NAND2X0 U20458 ( .IN1(n19298), .IN2(n19299), .QN(g24232) );
  XNOR2X1 U20459 ( .IN1(n10252), .IN2(n19300), .Q(n19299) );
  NAND2X0 U20460 ( .IN1(n5654), .IN2(n10954), .QN(n19300) );
  NOR2X0 U20461 ( .IN1(n19301), .IN2(n19302), .QN(n19298) );
  NOR2X0 U20462 ( .IN1(n11051), .IN2(g19334), .QN(n19302) );
  NOR2X0 U20463 ( .IN1(n10579), .IN2(n19251), .QN(n19301) );
  INVX0 U20464 ( .INP(n14152), .ZN(n19251) );
  INVX0 U20465 ( .INP(n19303), .ZN(g24231) );
  NAND2X0 U20466 ( .IN1(n10240), .IN2(n14152), .QN(n19303) );
  NOR2X0 U20467 ( .IN1(n11051), .IN2(n5654), .QN(n14152) );
  NAND2X0 U20468 ( .IN1(n19304), .IN2(n19305), .QN(g24216) );
  NAND2X0 U20469 ( .IN1(n17170), .IN2(g847), .QN(n19305) );
  NAND2X0 U20470 ( .IN1(n17947), .IN2(g854), .QN(n19304) );
  NAND2X0 U20471 ( .IN1(n19306), .IN2(n19307), .QN(g24215) );
  NAND2X0 U20472 ( .IN1(n19308), .IN2(g837), .QN(n19307) );
  NAND2X0 U20473 ( .IN1(n17947), .IN2(n19309), .QN(n19308) );
  NAND2X0 U20474 ( .IN1(n19310), .IN2(n19311), .QN(n19309) );
  NAND2X0 U20475 ( .IN1(g847), .IN2(g812), .QN(n19311) );
  NOR2X0 U20476 ( .IN1(n11052), .IN2(n19312), .QN(n19310) );
  NOR2X0 U20477 ( .IN1(n5728), .IN2(n10544), .QN(n19312) );
  NAND2X0 U20478 ( .IN1(n19313), .IN2(g703), .QN(n19306) );
  NAND2X0 U20479 ( .IN1(n19314), .IN2(n10954), .QN(n19313) );
  NAND2X0 U20480 ( .IN1(n5562), .IN2(n18359), .QN(n19314) );
  NOR2X0 U20481 ( .IN1(n17177), .IN2(n5709), .QN(n18359) );
  NAND2X0 U20482 ( .IN1(n19315), .IN2(n19316), .QN(g24214) );
  NAND2X0 U20483 ( .IN1(n19317), .IN2(g703), .QN(n19316) );
  NAND2X0 U20484 ( .IN1(n18354), .IN2(n19318), .QN(n19317) );
  NAND2X0 U20485 ( .IN1(n19319), .IN2(n10954), .QN(n19318) );
  INVX0 U20486 ( .INP(n18352), .ZN(n19319) );
  NOR2X0 U20487 ( .IN1(n5733), .IN2(n5562), .QN(n18352) );
  NOR2X0 U20488 ( .IN1(n17170), .IN2(n19320), .QN(n18354) );
  NOR2X0 U20489 ( .IN1(g847), .IN2(n11020), .QN(n19320) );
  NOR2X0 U20490 ( .IN1(n19321), .IN2(n19322), .QN(n19315) );
  NOR2X0 U20491 ( .IN1(g847), .IN2(n19323), .QN(n19322) );
  NAND2X0 U20492 ( .IN1(n19324), .IN2(n19325), .QN(n19323) );
  NOR2X0 U20493 ( .IN1(n5826), .IN2(n5822), .QN(n19325) );
  NOR2X0 U20494 ( .IN1(n5422), .IN2(n19326), .QN(n19324) );
  NOR2X0 U20495 ( .IN1(n5709), .IN2(n10882), .QN(n19321) );
  NAND2X0 U20496 ( .IN1(n19327), .IN2(n19328), .QN(g24211) );
  NAND2X0 U20497 ( .IN1(n2404), .IN2(n19329), .QN(n19328) );
  NAND2X0 U20498 ( .IN1(n10670), .IN2(g691), .QN(n19329) );
  NAND2X0 U20499 ( .IN1(n11059), .IN2(g546), .QN(n19327) );
  NOR2X0 U20500 ( .IN1(n14970), .IN2(n19330), .QN(g24210) );
  NAND2X0 U20501 ( .IN1(n19331), .IN2(n10954), .QN(n19330) );
  NAND2X0 U20502 ( .IN1(n19332), .IN2(n19333), .QN(n19331) );
  NAND2X0 U20503 ( .IN1(test_so72), .IN2(n16495), .QN(n19333) );
  NAND2X0 U20504 ( .IN1(n5606), .IN2(n5402), .QN(n16495) );
  NAND2X0 U20505 ( .IN1(g174), .IN2(g168), .QN(n19332) );
  NAND2X0 U20506 ( .IN1(n18001), .IN2(g203), .QN(n14970) );
  NOR2X0 U20507 ( .IN1(g513), .IN2(n5287), .QN(n18001) );
  NAND2X0 U20508 ( .IN1(n19334), .IN2(n19335), .QN(g24209) );
  NAND2X0 U20509 ( .IN1(n17170), .IN2(g417), .QN(n19335) );
  NAND2X0 U20510 ( .IN1(n17174), .IN2(g446), .QN(n19334) );
  INVX0 U20511 ( .INP(n19326), .ZN(n17174) );
  NAND2X0 U20512 ( .IN1(n19336), .IN2(n19337), .QN(g24208) );
  NAND2X0 U20513 ( .IN1(n11059), .IN2(g424), .QN(n19337) );
  NOR2X0 U20514 ( .IN1(n19338), .IN2(n19339), .QN(n19336) );
  NOR2X0 U20515 ( .IN1(n6008), .IN2(n19326), .QN(n19339) );
  NOR2X0 U20516 ( .IN1(n10124), .IN2(n17947), .QN(n19338) );
  NAND2X0 U20517 ( .IN1(n19340), .IN2(n19341), .QN(g24207) );
  NAND2X0 U20518 ( .IN1(n17170), .IN2(g441), .QN(n19341) );
  NAND2X0 U20519 ( .IN1(n17947), .IN2(g475), .QN(n19340) );
  NAND2X0 U20520 ( .IN1(n19342), .IN2(n19343), .QN(g24206) );
  NAND2X0 U20521 ( .IN1(n17170), .IN2(g437), .QN(n19343) );
  NAND2X0 U20522 ( .IN1(n17947), .IN2(g441), .QN(n19342) );
  NAND2X0 U20523 ( .IN1(n19344), .IN2(n19345), .QN(g24205) );
  NAND2X0 U20524 ( .IN1(n11060), .IN2(g437), .QN(n19345) );
  NOR2X0 U20525 ( .IN1(n19346), .IN2(n19347), .QN(n19344) );
  NOR2X0 U20526 ( .IN1(n10277), .IN2(n19326), .QN(n19347) );
  NOR2X0 U20527 ( .IN1(n17947), .IN2(n10693), .QN(n19346) );
  NAND2X0 U20528 ( .IN1(n19348), .IN2(n19349), .QN(g24204) );
  NAND2X0 U20529 ( .IN1(n17170), .IN2(g429), .QN(n19349) );
  NAND2X0 U20530 ( .IN1(test_so23), .IN2(n17947), .QN(n19348) );
  NAND2X0 U20531 ( .IN1(n19350), .IN2(n19351), .QN(g24203) );
  NAND2X0 U20532 ( .IN1(n17170), .IN2(g401), .QN(n19351) );
  NAND2X0 U20533 ( .IN1(n17947), .IN2(g429), .QN(n19350) );
  NAND2X0 U20534 ( .IN1(n19352), .IN2(n19353), .QN(g24202) );
  NAND2X0 U20535 ( .IN1(n17170), .IN2(g424), .QN(n19353) );
  NAND2X0 U20536 ( .IN1(n17947), .IN2(g411), .QN(n19352) );
  NAND2X0 U20537 ( .IN1(n19354), .IN2(n19355), .QN(g24201) );
  NAND2X0 U20538 ( .IN1(n17170), .IN2(g405), .QN(n19355) );
  INVX0 U20539 ( .INP(n17947), .ZN(n17170) );
  NAND2X0 U20540 ( .IN1(n17947), .IN2(g392), .QN(n19354) );
  NAND2X0 U20541 ( .IN1(n19356), .IN2(n19357), .QN(g24200) );
  NAND2X0 U20542 ( .IN1(n11059), .IN2(g401), .QN(n19357) );
  NOR2X0 U20543 ( .IN1(n19358), .IN2(n19359), .QN(n19356) );
  NOR2X0 U20544 ( .IN1(n10272), .IN2(n17947), .QN(n19359) );
  NAND2X0 U20545 ( .IN1(n10932), .IN2(n17177), .QN(n17947) );
  INVX0 U20546 ( .INP(n4948), .ZN(n17177) );
  NOR2X0 U20547 ( .IN1(n19326), .IN2(n19360), .QN(n19358) );
  NAND2X0 U20548 ( .IN1(n5821), .IN2(g854), .QN(n19360) );
  NAND2X0 U20549 ( .IN1(n4948), .IN2(n10954), .QN(n19326) );
  NOR2X0 U20550 ( .IN1(g22), .IN2(g25), .QN(g23190) );
  NAND2X0 U20551 ( .IN1(n19361), .IN2(n19362), .QN(g21901) );
  NAND2X0 U20552 ( .IN1(n11059), .IN2(g2946), .QN(n19362) );
  NAND2X0 U20553 ( .IN1(n19363), .IN2(n10954), .QN(n19361) );
  NAND2X0 U20554 ( .IN1(n19364), .IN2(n19365), .QN(n19363) );
  NAND2X0 U20555 ( .IN1(n5694), .IN2(g4180), .QN(n19365) );
  NAND2X0 U20556 ( .IN1(n5380), .IN2(n19366), .QN(n19364) );
  NAND2X0 U20557 ( .IN1(n5694), .IN2(n19367), .QN(n19366) );
  NAND2X0 U20558 ( .IN1(n19368), .IN2(n19369), .QN(n19367) );
  NOR2X0 U20559 ( .IN1(n19370), .IN2(n19371), .QN(n19369) );
  NAND2X0 U20560 ( .IN1(DFF_480_n1), .IN2(DFF_909_n1), .QN(n19371) );
  NAND2X0 U20561 ( .IN1(n10262), .IN2(DFF_1234_n1), .QN(n19370) );
  NOR2X0 U20562 ( .IN1(g8787), .IN2(n19372), .QN(n19368) );
  NAND2X0 U20563 ( .IN1(n10264), .IN2(n10263), .QN(n19372) );
  NAND2X0 U20564 ( .IN1(n19373), .IN2(n19374), .QN(g21900) );
  NAND2X0 U20565 ( .IN1(n11060), .IN2(g4239), .QN(n19374) );
  NAND2X0 U20566 ( .IN1(n19375), .IN2(n10938), .QN(n19373) );
  NOR2X0 U20567 ( .IN1(g10122_Tj), .IN2(g4297), .QN(n19375) );
  XOR2X1 U20568 ( .IN1(n19376), .IN2(n10575), .Q(g21899) );
  NAND2X0 U20569 ( .IN1(n10935), .IN2(g9019), .QN(n19376) );
  NAND2X0 U20570 ( .IN1(n19377), .IN2(n19378), .QN(g21898) );
  NAND2X0 U20571 ( .IN1(n10575), .IN2(n10952), .QN(n19378) );
  INVX0 U20572 ( .INP(n19379), .ZN(n19377) );
  NOR2X0 U20573 ( .IN1(n10902), .IN2(n10593), .QN(n19379) );
  XOR2X1 U20574 ( .IN1(n19380), .IN2(n10576), .Q(g21897) );
  NAND2X0 U20575 ( .IN1(n10935), .IN2(g8839), .QN(n19380) );
  NAND2X0 U20576 ( .IN1(n19381), .IN2(n19382), .QN(g21896) );
  NAND2X0 U20577 ( .IN1(n10576), .IN2(n10939), .QN(n19382) );
  NAND2X0 U20578 ( .IN1(n11061), .IN2(g4245), .QN(n19381) );
  NAND2X0 U20579 ( .IN1(n19383), .IN2(n19384), .QN(g21895) );
  NAND2X0 U20580 ( .IN1(n19385), .IN2(g4264), .QN(n19384) );
  NAND2X0 U20581 ( .IN1(n19386), .IN2(n10938), .QN(n19385) );
  NAND2X0 U20582 ( .IN1(n5763), .IN2(g4258), .QN(n19386) );
  NAND2X0 U20583 ( .IN1(n19387), .IN2(g4269), .QN(n19383) );
  INVX0 U20584 ( .INP(n19103), .ZN(n19387) );
  NOR2X0 U20585 ( .IN1(g21893), .IN2(n19388), .QN(n19103) );
  NOR2X0 U20586 ( .IN1(g4264), .IN2(n11021), .QN(n19388) );
  NAND2X0 U20587 ( .IN1(n19389), .IN2(n19390), .QN(g21894) );
  NAND2X0 U20588 ( .IN1(n19391), .IN2(g4258), .QN(n19390) );
  NAND2X0 U20589 ( .IN1(n10934), .IN2(g4264), .QN(n19391) );
  NAND2X0 U20590 ( .IN1(g21893), .IN2(g4264), .QN(n19389) );
  NOR2X0 U20591 ( .IN1(g4258), .IN2(n11021), .QN(g21893) );
  NAND2X0 U20592 ( .IN1(n19392), .IN2(n19393), .QN(g21892) );
  NAND2X0 U20593 ( .IN1(n10210), .IN2(n10939), .QN(n19393) );
  NAND2X0 U20594 ( .IN1(n11061), .IN2(g4273), .QN(n19392) );
  NAND2X0 U20595 ( .IN1(n19394), .IN2(n19395), .QN(g21891) );
  NAND2X0 U20596 ( .IN1(n11067), .IN2(g4180), .QN(n19395) );
  NAND2X0 U20597 ( .IN1(n19108), .IN2(n10955), .QN(n19394) );
  NAND2X0 U20598 ( .IN1(n19396), .IN2(n19397), .QN(n19108) );
  NAND2X0 U20599 ( .IN1(n10552), .IN2(g4253), .QN(n19397) );
  NAND2X0 U20600 ( .IN1(n5484), .IN2(n10551), .QN(n19396) );
  NOR2X0 U20601 ( .IN1(n10907), .IN2(DFF_1381_n1), .QN(g21727) );
  NOR2X0 U20602 ( .IN1(n5750), .IN2(n10839), .QN(g18597) );
  INVX0 U20603 ( .INP(g5), .ZN(g12833) );
  NOR2X0 U5116_U2 ( .IN1(g34783), .IN2(n2730), .QN(U5116_n1) );
  INVX0 U5116_U1 ( .INP(U5116_n1), .ZN(g34221) );
  NOR2X0 U5126_U2 ( .IN1(n4836), .IN2(n4896), .QN(U5126_n1) );
  INVX0 U5126_U1 ( .INP(U5126_n1), .ZN(n4895) );
  NOR2X0 U5127_U2 ( .IN1(n4837), .IN2(n4921), .QN(U5127_n1) );
  INVX0 U5127_U1 ( .INP(U5127_n1), .ZN(n4920) );
  NOR2X0 U5128_U2 ( .IN1(n2787), .IN2(n4411), .QN(U5128_n1) );
  INVX0 U5128_U1 ( .INP(U5128_n1), .ZN(n5045) );
  NOR2X0 U5129_U2 ( .IN1(g559), .IN2(g9048), .QN(U5129_n1) );
  INVX0 U5129_U1 ( .INP(U5129_n1), .ZN(n4959) );
  INVX0 U5353_U2 ( .INP(n5960), .ZN(U5353_n1) );
  NOR2X0 U5353_U1 ( .IN1(n10629), .IN2(U5353_n1), .QN(n4689) );
  INVX0 U5355_U2 ( .INP(n5961), .ZN(U5355_n1) );
  NOR2X0 U5355_U1 ( .IN1(n10624), .IN2(U5355_n1), .QN(n4708) );
  INVX0 U5961_U2 ( .INP(n3593), .ZN(U5961_n1) );
  NOR2X0 U5961_U1 ( .IN1(n3589), .IN2(U5961_n1), .QN(n3595) );
  INVX0 U5962_U2 ( .INP(n3574), .ZN(U5962_n1) );
  NOR2X0 U5962_U1 ( .IN1(n3570), .IN2(U5962_n1), .QN(n3576) );
  INVX0 U5963_U2 ( .INP(n3517), .ZN(U5963_n1) );
  NOR2X0 U5963_U1 ( .IN1(n3513), .IN2(U5963_n1), .QN(n3519) );
  INVX0 U5964_U2 ( .INP(n3628), .ZN(U5964_n1) );
  NOR2X0 U5964_U1 ( .IN1(n3624), .IN2(U5964_n1), .QN(n3630) );
  INVX0 U5965_U2 ( .INP(n3555), .ZN(U5965_n1) );
  NOR2X0 U5965_U1 ( .IN1(n3551), .IN2(U5965_n1), .QN(n3557) );
  INVX0 U5966_U2 ( .INP(n3646), .ZN(U5966_n1) );
  NOR2X0 U5966_U1 ( .IN1(n3642), .IN2(U5966_n1), .QN(n3648) );
  INVX0 U5967_U2 ( .INP(n3536), .ZN(U5967_n1) );
  NOR2X0 U5967_U1 ( .IN1(n3532), .IN2(U5967_n1), .QN(n3538) );
  INVX0 U5968_U2 ( .INP(n3611), .ZN(U5968_n1) );
  NOR2X0 U5968_U1 ( .IN1(n3607), .IN2(U5968_n1), .QN(n3613) );
  INVX0 U6100_U2 ( .INP(n3635), .ZN(U6100_n1) );
  NOR2X0 U6100_U1 ( .IN1(n11014), .IN2(U6100_n1), .QN(n4888) );
  INVX0 U6211_U2 ( .INP(n3623), .ZN(U6211_n1) );
  NOR2X0 U6211_U1 ( .IN1(n1730), .IN2(U6211_n1), .QN(n3622) );
  INVX0 U6212_U2 ( .INP(n3587), .ZN(U6212_n1) );
  NOR2X0 U6212_U1 ( .IN1(n3588), .IN2(U6212_n1), .QN(n3586) );
  INVX0 U6213_U2 ( .INP(n3605), .ZN(U6213_n1) );
  NOR2X0 U6213_U1 ( .IN1(n3606), .IN2(U6213_n1), .QN(n3604) );
  INVX0 U6214_U2 ( .INP(n3568), .ZN(U6214_n1) );
  NOR2X0 U6214_U1 ( .IN1(n3569), .IN2(U6214_n1), .QN(n3567) );
  INVX0 U6215_U2 ( .INP(n3549), .ZN(U6215_n1) );
  NOR2X0 U6215_U1 ( .IN1(n3550), .IN2(U6215_n1), .QN(n3548) );
  INVX0 U6216_U2 ( .INP(n3512), .ZN(U6216_n1) );
  NOR2X0 U6216_U1 ( .IN1(n3006), .IN2(U6216_n1), .QN(n3511) );
  INVX0 U6217_U2 ( .INP(n3531), .ZN(U6217_n1) );
  NOR2X0 U6217_U1 ( .IN1(n3007), .IN2(U6217_n1), .QN(n3530) );
  INVX0 U6218_U2 ( .INP(n3641), .ZN(U6218_n1) );
  NOR2X0 U6218_U1 ( .IN1(n831), .IN2(U6218_n1), .QN(n3640) );
  INVX0 U6279_U2 ( .INP(n4537), .ZN(U6279_n1) );
  NOR2X0 U6279_U1 ( .IN1(n5337), .IN2(U6279_n1), .QN(n4201) );
  INVX0 U6280_U2 ( .INP(n4201), .ZN(U6280_n1) );
  NOR2X0 U6280_U1 ( .IN1(n5336), .IN2(U6280_n1), .QN(n3745) );
  INVX0 U6281_U2 ( .INP(n3745), .ZN(U6281_n1) );
  NOR2X0 U6281_U1 ( .IN1(n5294), .IN2(U6281_n1), .QN(n3684) );
  INVX0 U6282_U2 ( .INP(n3684), .ZN(U6282_n1) );
  NOR2X0 U6282_U1 ( .IN1(n5552), .IN2(U6282_n1), .QN(n3274) );
  INVX0 U6283_U2 ( .INP(n3274), .ZN(U6283_n1) );
  NOR2X0 U6283_U1 ( .IN1(n5472), .IN2(U6283_n1), .QN(n2982) );
  INVX0 U6284_U2 ( .INP(n2982), .ZN(U6284_n1) );
  NOR2X0 U6284_U1 ( .IN1(n5476), .IN2(U6284_n1), .QN(n2706) );
  INVX0 U6285_U2 ( .INP(n2706), .ZN(U6285_n1) );
  NOR2X0 U6285_U1 ( .IN1(n5550), .IN2(U6285_n1), .QN(n2649) );
  INVX0 U6286_U2 ( .INP(n2649), .ZN(U6286_n1) );
  NOR2X0 U6286_U1 ( .IN1(n5473), .IN2(U6286_n1), .QN(n2556) );
  INVX0 U6287_U2 ( .INP(n2556), .ZN(U6287_n1) );
  NOR2X0 U6287_U1 ( .IN1(n5475), .IN2(U6287_n1), .QN(n2509) );
  INVX0 U6288_U2 ( .INP(n2509), .ZN(U6288_n1) );
  NOR2X0 U6288_U1 ( .IN1(n5474), .IN2(U6288_n1), .QN(n2487) );
  INVX0 U6289_U2 ( .INP(n2487), .ZN(U6289_n1) );
  NOR2X0 U6289_U1 ( .IN1(n5339), .IN2(U6289_n1), .QN(n2427) );
  INVX0 U6290_U2 ( .INP(n2427), .ZN(U6290_n1) );
  NOR2X0 U6290_U1 ( .IN1(n5672), .IN2(U6290_n1), .QN(n2423) );
  INVX0 U6291_U2 ( .INP(n5), .ZN(U6291_n1) );
  NOR2X0 U6291_U1 ( .IN1(n5335), .IN2(U6291_n1), .QN(n4537) );
  INVX0 U6292_U2 ( .INP(n4959), .ZN(U6292_n1) );
  NOR2X0 U6292_U1 ( .IN1(n11014), .IN2(U6292_n1), .QN(n2421) );
  INVX0 U6338_U2 ( .INP(n4210), .ZN(U6338_n1) );
  NOR2X0 U6338_U1 ( .IN1(n11024), .IN2(U6338_n1), .QN(n3765) );
  INVX0 U6341_U2 ( .INP(n3765), .ZN(U6341_n1) );
  NOR2X0 U6341_U1 ( .IN1(n3479), .IN2(U6341_n1), .QN(n3951) );
  INVX0 U6342_U2 ( .INP(n3765), .ZN(U6342_n1) );
  NOR2X0 U6342_U1 ( .IN1(n3404), .IN2(U6342_n1), .QN(n3774) );
  INVX0 U6343_U2 ( .INP(n3765), .ZN(U6343_n1) );
  NOR2X0 U6343_U1 ( .IN1(n3424), .IN2(U6343_n1), .QN(n3842) );
  INVX0 U6344_U2 ( .INP(n3765), .ZN(U6344_n1) );
  NOR2X0 U6344_U1 ( .IN1(n3414), .IN2(U6344_n1), .QN(n3808) );
  INVX0 U6345_U2 ( .INP(n3765), .ZN(U6345_n1) );
  NOR2X0 U6345_U1 ( .IN1(n3444), .IN2(U6345_n1), .QN(n3908) );
  INVX0 U6346_U2 ( .INP(n3765), .ZN(U6346_n1) );
  NOR2X0 U6346_U1 ( .IN1(n3489), .IN2(U6346_n1), .QN(n3984) );
  INVX0 U6347_U2 ( .INP(n3765), .ZN(U6347_n1) );
  NOR2X0 U6347_U1 ( .IN1(n3434), .IN2(U6347_n1), .QN(n3875) );
  INVX0 U6348_U2 ( .INP(n3765), .ZN(U6348_n1) );
  NOR2X0 U6348_U1 ( .IN1(n128), .IN2(U6348_n1), .QN(n4015) );
  INVX0 U6349_U2 ( .INP(n3765), .ZN(U6349_n1) );
  NOR2X0 U6349_U1 ( .IN1(n792), .IN2(U6349_n1), .QN(n3914) );
  INVX0 U6350_U2 ( .INP(n3765), .ZN(U6350_n1) );
  NOR2X0 U6350_U1 ( .IN1(n3406), .IN2(U6350_n1), .QN(n3780) );
  INVX0 U6351_U2 ( .INP(n3765), .ZN(U6351_n1) );
  NOR2X0 U6351_U1 ( .IN1(n3481), .IN2(U6351_n1), .QN(n3957) );
  INVX0 U6352_U2 ( .INP(n3765), .ZN(U6352_n1) );
  NOR2X0 U6352_U1 ( .IN1(n1101), .IN2(U6352_n1), .QN(n3848) );
  INVX0 U6353_U2 ( .INP(n3765), .ZN(U6353_n1) );
  NOR2X0 U6353_U1 ( .IN1(n3491), .IN2(U6353_n1), .QN(n3990) );
  INVX0 U6354_U2 ( .INP(n3765), .ZN(U6354_n1) );
  NOR2X0 U6354_U1 ( .IN1(n3416), .IN2(U6354_n1), .QN(n3814) );
  INVX0 U6355_U2 ( .INP(n3765), .ZN(U6355_n1) );
  NOR2X0 U6355_U1 ( .IN1(n552), .IN2(U6355_n1), .QN(n3881) );
  INVX0 U6356_U2 ( .INP(n3765), .ZN(U6356_n1) );
  NOR2X0 U6356_U1 ( .IN1(n3502), .IN2(U6356_n1), .QN(n4022) );
  INVX0 U6357_U2 ( .INP(n3765), .ZN(U6357_n1) );
  NOR2X0 U6357_U1 ( .IN1(n3501), .IN2(U6357_n1), .QN(n4027) );
  INVX0 U6358_U2 ( .INP(n3765), .ZN(U6358_n1) );
  NOR2X0 U6358_U1 ( .IN1(n3407), .IN2(U6358_n1), .QN(n3785) );
  INVX0 U6359_U2 ( .INP(n3765), .ZN(U6359_n1) );
  NOR2X0 U6359_U1 ( .IN1(n3482), .IN2(U6359_n1), .QN(n3962) );
  INVX0 U6360_U2 ( .INP(n3765), .ZN(U6360_n1) );
  NOR2X0 U6360_U1 ( .IN1(n3427), .IN2(U6360_n1), .QN(n3853) );
  INVX0 U6361_U2 ( .INP(n3765), .ZN(U6361_n1) );
  NOR2X0 U6361_U1 ( .IN1(n3437), .IN2(U6361_n1), .QN(n3886) );
  INVX0 U6362_U2 ( .INP(n3765), .ZN(U6362_n1) );
  NOR2X0 U6362_U1 ( .IN1(n3417), .IN2(U6362_n1), .QN(n3819) );
  INVX0 U6363_U2 ( .INP(n3765), .ZN(U6363_n1) );
  NOR2X0 U6363_U1 ( .IN1(n3492), .IN2(U6363_n1), .QN(n3995) );
  INVX0 U6364_U2 ( .INP(n3765), .ZN(U6364_n1) );
  NOR2X0 U6364_U1 ( .IN1(n3447), .IN2(U6364_n1), .QN(n3919) );
  INVX0 U6365_U2 ( .INP(n3682), .ZN(U6365_n1) );
  NOR2X0 U6365_U1 ( .IN1(n5471), .IN2(U6365_n1), .QN(n3272) );
  INVX0 U6366_U2 ( .INP(n3272), .ZN(U6366_n1) );
  NOR2X0 U6366_U1 ( .IN1(n5331), .IN2(U6366_n1), .QN(n2980) );
  INVX0 U6367_U2 ( .INP(n2980), .ZN(U6367_n1) );
  NOR2X0 U6367_U1 ( .IN1(n5332), .IN2(U6367_n1), .QN(n2704) );
  INVX0 U6368_U2 ( .INP(n2704), .ZN(U6368_n1) );
  NOR2X0 U6368_U1 ( .IN1(n5333), .IN2(U6368_n1), .QN(n2647) );
  INVX0 U6369_U2 ( .INP(n2647), .ZN(U6369_n1) );
  NOR2X0 U6369_U1 ( .IN1(n5334), .IN2(U6369_n1), .QN(n2554) );
  INVX0 U6370_U2 ( .INP(n2554), .ZN(U6370_n1) );
  NOR2X0 U6370_U1 ( .IN1(n5330), .IN2(U6370_n1), .QN(n2507) );
  INVX0 U6371_U2 ( .INP(n2507), .ZN(U6371_n1) );
  NOR2X0 U6371_U1 ( .IN1(n5551), .IN2(U6371_n1), .QN(n2485) );
  INVX0 U6372_U2 ( .INP(n2485), .ZN(U6372_n1) );
  NOR2X0 U6372_U1 ( .IN1(n5293), .IN2(U6372_n1), .QN(n2425) );
  INVX0 U6373_U2 ( .INP(n2425), .ZN(U6373_n1) );
  NOR2X0 U6373_U1 ( .IN1(n5292), .IN2(U6373_n1), .QN(n2419) );
  INVX0 U6374_U2 ( .INP(n3743), .ZN(U6374_n1) );
  NOR2X0 U6374_U1 ( .IN1(n5470), .IN2(U6374_n1), .QN(n3682) );
  INVX0 U6375_U2 ( .INP(n2419), .ZN(U6375_n1) );
  NOR2X0 U6375_U1 ( .IN1(n5291), .IN2(U6375_n1), .QN(n2405) );
  INVX0 U6417_U2 ( .INP(n4198), .ZN(U6417_n1) );
  NOR2X0 U6417_U1 ( .IN1(n11014), .IN2(U6417_n1), .QN(n2404) );
  INVX0 U6446_U2 ( .INP(g110), .ZN(U6446_n1) );
  NOR2X0 U6446_U1 ( .IN1(n1770), .IN2(U6446_n1), .QN(n3524) );
  INVX0 U6465_U2 ( .INP(n832), .ZN(U6465_n1) );
  NOR2X0 U6465_U1 ( .IN1(n5600), .IN2(U6465_n1), .QN(n4388) );
  INVX0 U6497_U2 ( .INP(n864), .ZN(U6497_n1) );
  NOR2X0 U6497_U1 ( .IN1(n3635), .IN2(U6497_n1), .QN(n3005) );
  INVX0 U6523_U2 ( .INP(n4946), .ZN(U6523_n1) );
  NOR2X0 U6523_U1 ( .IN1(n11014), .IN2(U6523_n1), .QN(n4945) );
  INVX0 U6542_U2 ( .INP(n864), .ZN(U6542_n1) );
  NOR2X0 U6542_U1 ( .IN1(n5300), .IN2(U6542_n1), .QN(n3525) );
  INVX0 U6552_U2 ( .INP(n3281), .ZN(U6552_n1) );
  NOR2X0 U6552_U1 ( .IN1(n5676), .IN2(U6552_n1), .QN(n3277) );
  INVX0 U6553_U2 ( .INP(n3276), .ZN(U6553_n1) );
  NOR2X0 U6553_U1 ( .IN1(n5680), .IN2(U6553_n1), .QN(n2989) );
  INVX0 U6554_U2 ( .INP(n3277), .ZN(U6554_n1) );
  NOR2X0 U6554_U1 ( .IN1(n5677), .IN2(U6554_n1), .QN(n2991) );
  INVX0 U6555_U2 ( .INP(n103), .ZN(U6555_n1) );
  NOR2X0 U6555_U1 ( .IN1(n5561), .IN2(U6555_n1), .QN(n3281) );
  INVX0 U6556_U2 ( .INP(n97), .ZN(U6556_n1) );
  NOR2X0 U6556_U1 ( .IN1(n5679), .IN2(U6556_n1), .QN(n3276) );
  INVX0 U6559_U2 ( .INP(n2991), .ZN(U6559_n1) );
  NOR2X0 U6559_U1 ( .IN1(n5678), .IN2(U6559_n1), .QN(n2710) );
  INVX0 U6560_U2 ( .INP(n2989), .ZN(U6560_n1) );
  NOR2X0 U6560_U1 ( .IN1(n5675), .IN2(U6560_n1), .QN(n2707) );
  INVX0 U6561_U2 ( .INP(n3174), .ZN(U6561_n1) );
  NOR2X0 U6561_U1 ( .IN1(n5327), .IN2(U6561_n1), .QN(n3116) );
  INVX0 U6570_U2 ( .INP(n3362), .ZN(U6570_n1) );
  NOR2X0 U6570_U1 ( .IN1(n5477), .IN2(U6570_n1), .QN(n2527) );
  INVX0 U6911_U2 ( .INP(n3115), .ZN(U6911_n1) );
  NOR2X0 U6911_U1 ( .IN1(n2726), .IN2(U6911_n1), .QN(n3111) );
  INVX0 U6912_U2 ( .INP(n3115), .ZN(U6912_n1) );
  NOR2X0 U6912_U1 ( .IN1(n2727), .IN2(U6912_n1), .QN(n3131) );
  INVX0 U6917_U2 ( .INP(n3933), .ZN(U6917_n1) );
  NOR2X0 U6917_U1 ( .IN1(n5350), .IN2(U6917_n1), .QN(n3799) );
  INVX0 U6926_U2 ( .INP(n3664), .ZN(U6926_n1) );
  NOR2X0 U6926_U1 ( .IN1(n5674), .IN2(U6926_n1), .QN(n3662) );
  INVX0 U6927_U2 ( .INP(n3673), .ZN(U6927_n1) );
  NOR2X0 U6927_U1 ( .IN1(n5673), .IN2(U6927_n1), .QN(n3671) );
  INVX0 U6929_U2 ( .INP(n3505), .ZN(U6929_n1) );
  NOR2X0 U6929_U1 ( .IN1(n3506), .IN2(U6929_n1), .QN(n2790) );
  INVX0 U6931_U2 ( .INP(n4490), .ZN(U6931_n1) );
  NOR2X0 U6931_U1 ( .IN1(n5554), .IN2(U6931_n1), .QN(n4178) );
  INVX0 U6932_U2 ( .INP(n4514), .ZN(U6932_n1) );
  NOR2X0 U6932_U1 ( .IN1(n5555), .IN2(U6932_n1), .QN(n4196) );
  INVX0 U6933_U2 ( .INP(n4178), .ZN(U6933_n1) );
  NOR2X0 U6933_U1 ( .IN1(n5558), .IN2(U6933_n1), .QN(n3736) );
  INVX0 U6934_U2 ( .INP(n4196), .ZN(U6934_n1) );
  NOR2X0 U6934_U1 ( .IN1(n5559), .IN2(U6934_n1), .QN(n3741) );
  INVX0 U6935_U2 ( .INP(n3736), .ZN(U6935_n1) );
  NOR2X0 U6935_U1 ( .IN1(n5553), .IN2(U6935_n1), .QN(n3664) );
  INVX0 U6936_U2 ( .INP(n3741), .ZN(U6936_n1) );
  NOR2X0 U6936_U1 ( .IN1(n5560), .IN2(U6936_n1), .QN(n3673) );
  INVX0 U6937_U2 ( .INP(n2601), .ZN(U6937_n1) );
  NOR2X0 U6937_U1 ( .IN1(n5303), .IN2(U6937_n1), .QN(n2598) );
  INVX0 U6938_U2 ( .INP(n1249), .ZN(U6938_n1) );
  NOR2X0 U6938_U1 ( .IN1(n5556), .IN2(U6938_n1), .QN(n4490) );
  INVX0 U6939_U2 ( .INP(n315), .ZN(U6939_n1) );
  NOR2X0 U6939_U1 ( .IN1(n5557), .IN2(U6939_n1), .QN(n4514) );
  INVX0 U6940_U2 ( .INP(n4814), .ZN(U6940_n1) );
  NOR2X0 U6940_U1 ( .IN1(n5422), .IN2(U6940_n1), .QN(n4519) );
  INVX0 U6941_U2 ( .INP(n2607), .ZN(U6941_n1) );
  NOR2X0 U6941_U1 ( .IN1(n5323), .IN2(U6941_n1), .QN(n2594) );
  INVX0 U6944_U2 ( .INP(n3084), .ZN(U6944_n1) );
  NOR2X0 U6944_U1 ( .IN1(n5348), .IN2(U6944_n1), .QN(n3033) );
  INVX0 U6950_U2 ( .INP(n2598), .ZN(U6950_n1) );
  NOR2X0 U6950_U1 ( .IN1(n5365), .IN2(U6950_n1), .QN(n2590) );
  INVX0 U6954_U2 ( .INP(n3122), .ZN(U6954_n1) );
  NOR2X0 U6954_U1 ( .IN1(n2727), .IN2(U6954_n1), .QN(n3125) );
  INVX0 U6955_U2 ( .INP(n735), .ZN(U6955_n1) );
  NOR2X0 U6955_U1 ( .IN1(n2726), .IN2(U6955_n1), .QN(n3105) );
  INVX0 U6956_U2 ( .INP(n3141), .ZN(U6956_n1) );
  NOR2X0 U6956_U1 ( .IN1(n3146), .IN2(U6956_n1), .QN(n3145) );
  INVX0 U6957_U2 ( .INP(n751), .ZN(U6957_n1) );
  NOR2X0 U6957_U1 ( .IN1(n3165), .IN2(U6957_n1), .QN(n3164) );
  INVX0 U7174_U2 ( .INP(n2423), .ZN(U7174_n1) );
  NOR2X0 U7174_U1 ( .IN1(n5288), .IN2(U7174_n1), .QN(n2422) );
  INVX0 U7248_U2 ( .INP(n2), .ZN(U7248_n1) );
  NOR2X0 U7248_U1 ( .IN1(g1536), .IN2(U7248_n1), .QN(n4173) );
  INVX0 U7249_U2 ( .INP(n4), .ZN(U7249_n1) );
  NOR2X0 U7249_U1 ( .IN1(g1193), .IN2(U7249_n1), .QN(n4191) );
  INVX0 U7402_U2 ( .INP(n4034), .ZN(U7402_n1) );
  NOR2X0 U7402_U1 ( .IN1(n4020), .IN2(U7402_n1), .QN(n4037) );
  INVX0 U7405_U2 ( .INP(n4034), .ZN(U7405_n1) );
  NOR2X0 U7405_U1 ( .IN1(n4014), .IN2(U7405_n1), .QN(n4039) );
  INVX0 U7413_U2 ( .INP(n3969), .ZN(U7413_n1) );
  NOR2X0 U7413_U1 ( .IN1(n3947), .IN2(U7413_n1), .QN(n3972) );
  INVX0 U7416_U2 ( .INP(n3926), .ZN(U7416_n1) );
  NOR2X0 U7416_U1 ( .IN1(n3904), .IN2(U7416_n1), .QN(n3929) );
  INVX0 U7427_U2 ( .INP(n3860), .ZN(U7427_n1) );
  NOR2X0 U7427_U1 ( .IN1(n3838), .IN2(U7427_n1), .QN(n3863) );
  INVX0 U7438_U2 ( .INP(n4002), .ZN(U7438_n1) );
  NOR2X0 U7438_U1 ( .IN1(n3978), .IN2(U7438_n1), .QN(n4003) );
  INVX0 U7449_U2 ( .INP(n4034), .ZN(U7449_n1) );
  NOR2X0 U7449_U1 ( .IN1(n582), .IN2(U7449_n1), .QN(n4032) );
  INVX0 U7455_U2 ( .INP(n4034), .ZN(U7455_n1) );
  NOR2X0 U7455_U1 ( .IN1(n580), .IN2(U7455_n1), .QN(n4035) );
  INVX0 U7464_U2 ( .INP(n3792), .ZN(U7464_n1) );
  NOR2X0 U7464_U1 ( .IN1(n3773), .IN2(U7464_n1), .QN(n3797) );
  INVX0 U7467_U2 ( .INP(n3792), .ZN(U7467_n1) );
  NOR2X0 U7467_U1 ( .IN1(n3776), .IN2(U7467_n1), .QN(n3790) );
  INVX0 U7482_U2 ( .INP(n3792), .ZN(U7482_n1) );
  NOR2X0 U7482_U1 ( .IN1(n3770), .IN2(U7482_n1), .QN(n3795) );
  INVX0 U7492_U2 ( .INP(n3893), .ZN(U7492_n1) );
  NOR2X0 U7492_U1 ( .IN1(n3877), .IN2(U7492_n1), .QN(n3891) );
  INVX0 U7513_U2 ( .INP(n3826), .ZN(U7513_n1) );
  NOR2X0 U7513_U1 ( .IN1(n3802), .IN2(U7513_n1), .QN(n3827) );
  INVX0 U7516_U2 ( .INP(n3893), .ZN(U7516_n1) );
  NOR2X0 U7516_U1 ( .IN1(n978), .IN2(U7516_n1), .QN(n3896) );
  INVX0 U7549_U2 ( .INP(n4002), .ZN(U7549_n1) );
  NOR2X0 U7549_U1 ( .IN1(n3983), .IN2(U7549_n1), .QN(n4007) );
  INVX0 U7561_U2 ( .INP(n3926), .ZN(U7561_n1) );
  NOR2X0 U7561_U1 ( .IN1(n3907), .IN2(U7561_n1), .QN(n3931) );
  INVX0 U7574_U2 ( .INP(n3792), .ZN(U7574_n1) );
  NOR2X0 U7574_U1 ( .IN1(n3768), .IN2(U7574_n1), .QN(n3793) );
  INVX0 U7577_U2 ( .INP(n3926), .ZN(U7577_n1) );
  NOR2X0 U7577_U1 ( .IN1(n3910), .IN2(U7577_n1), .QN(n3924) );
  INVX0 U7585_U2 ( .INP(n3826), .ZN(U7585_n1) );
  NOR2X0 U7585_U1 ( .IN1(n3807), .IN2(U7585_n1), .QN(n3831) );
  INVX0 U7595_U2 ( .INP(n3826), .ZN(U7595_n1) );
  NOR2X0 U7595_U1 ( .IN1(n3804), .IN2(U7595_n1), .QN(n3829) );
  INVX0 U7614_U2 ( .INP(n3926), .ZN(U7614_n1) );
  NOR2X0 U7614_U1 ( .IN1(n3902), .IN2(U7614_n1), .QN(n3927) );
  INVX0 U7621_U2 ( .INP(n3969), .ZN(U7621_n1) );
  NOR2X0 U7621_U1 ( .IN1(n3950), .IN2(U7621_n1), .QN(n3974) );
  INVX0 U7629_U2 ( .INP(n3893), .ZN(U7629_n1) );
  NOR2X0 U7629_U1 ( .IN1(n3874), .IN2(U7629_n1), .QN(n3898) );
  INVX0 U7636_U2 ( .INP(n3969), .ZN(U7636_n1) );
  NOR2X0 U7636_U1 ( .IN1(n3945), .IN2(U7636_n1), .QN(n3970) );
  INVX0 U7639_U2 ( .INP(n4002), .ZN(U7639_n1) );
  NOR2X0 U7639_U1 ( .IN1(n3986), .IN2(U7639_n1), .QN(n4000) );
  INVX0 U7649_U2 ( .INP(n3860), .ZN(U7649_n1) );
  NOR2X0 U7649_U1 ( .IN1(n3841), .IN2(U7649_n1), .QN(n3865) );
  INVX0 U7652_U2 ( .INP(n3860), .ZN(U7652_n1) );
  NOR2X0 U7652_U1 ( .IN1(n3836), .IN2(U7652_n1), .QN(n3861) );
  INVX0 U7668_U2 ( .INP(n3826), .ZN(U7668_n1) );
  NOR2X0 U7668_U1 ( .IN1(n3810), .IN2(U7668_n1), .QN(n3824) );
  INVX0 U7673_U2 ( .INP(n3893), .ZN(U7673_n1) );
  NOR2X0 U7673_U1 ( .IN1(n3869), .IN2(U7673_n1), .QN(n3894) );
  INVX0 U7690_U2 ( .INP(n3969), .ZN(U7690_n1) );
  NOR2X0 U7690_U1 ( .IN1(n3953), .IN2(U7690_n1), .QN(n3967) );
  INVX0 U7707_U2 ( .INP(n3860), .ZN(U7707_n1) );
  NOR2X0 U7707_U1 ( .IN1(n3844), .IN2(U7707_n1), .QN(n3858) );
  INVX0 U7712_U2 ( .INP(n4002), .ZN(U7712_n1) );
  NOR2X0 U7712_U1 ( .IN1(n3980), .IN2(U7712_n1), .QN(n4005) );
  INVX0 U7792_U2 ( .INP(g952), .ZN(U7792_n1) );
  NOR2X0 U7792_U1 ( .IN1(n11024), .IN2(U7792_n1), .QN(n2505) );
  INVX0 U7794_U2 ( .INP(g1296), .ZN(U7794_n1) );
  NOR2X0 U7794_U1 ( .IN1(n11024), .IN2(U7794_n1), .QN(n2499) );
  INVX0 U7895_U2 ( .INP(n1363), .ZN(U7895_n1) );
  NOR2X0 U7895_U1 ( .IN1(g113), .IN2(U7895_n1), .QN(n2760) );
  INVX0 U7897_U2 ( .INP(g6), .ZN(U7897_n1) );
  NOR2X0 U7897_U1 ( .IN1(g31), .IN2(U7897_n1), .QN(n3395) );
  INVX0 U7977_U2 ( .INP(g661), .ZN(U7977_n1) );
  NOR2X0 U7977_U1 ( .IN1(n11024), .IN2(U7977_n1), .QN(n4956) );
  INVX0 U8034_U2 ( .INP(n1269), .ZN(U8034_n1) );
  NOR2X0 U8034_U1 ( .IN1(n5612), .IN2(U8034_n1), .QN(n5026) );
  INVX0 U8036_U2 ( .INP(n418), .ZN(U8036_n1) );
  NOR2X0 U8036_U1 ( .IN1(n5340), .IN2(U8036_n1), .QN(n3941) );
  INVX0 U8050_U2 ( .INP(n227), .ZN(U8050_n1) );
  NOR2X0 U8050_U1 ( .IN1(g1367), .IN2(U8050_n1), .QN(n3733) );
  INVX0 U8055_U2 ( .INP(g1345), .ZN(U8055_n1) );
  NOR2X0 U8055_U1 ( .IN1(n11014), .IN2(U8055_n1), .QN(n4798) );
  INVX0 U8060_U2 ( .INP(g1002), .ZN(U8060_n1) );
  NOR2X0 U8060_U1 ( .IN1(n11024), .IN2(U8060_n1), .QN(n4805) );
  INVX0 U8070_U2 ( .INP(n3734), .ZN(U8070_n1) );
  NOR2X0 U8070_U1 ( .IN1(g1361), .IN2(U8070_n1), .QN(n4175) );
  INVX0 U8074_U2 ( .INP(n3739), .ZN(U8074_n1) );
  NOR2X0 U8074_U1 ( .IN1(g1018), .IN2(U8074_n1), .QN(n4193) );
  INVX0 U8088_U2 ( .INP(n591), .ZN(U8088_n1) );
  NOR2X0 U8088_U1 ( .IN1(g1024), .IN2(U8088_n1), .QN(n3738) );
  INVX0 U8112_U2 ( .INP(n4525), .ZN(U8112_n1) );
  NOR2X0 U8112_U1 ( .IN1(n4523), .IN2(U8112_n1), .QN(n4524) );
  INVX0 U8113_U2 ( .INP(n4526), .ZN(U8113_n1) );
  NOR2X0 U8113_U1 ( .IN1(n5751), .IN2(U8113_n1), .QN(n4523) );
  INVX0 U8147_U2 ( .INP(g4659), .ZN(U8147_n1) );
  NOR2X0 U8147_U1 ( .IN1(n2573), .IN2(U8147_n1), .QN(n2577) );
  INVX0 U8165_U2 ( .INP(g4849), .ZN(U8165_n1) );
  NOR2X0 U8165_U1 ( .IN1(n2563), .IN2(U8165_n1), .QN(n2567) );
  INVX0 U8185_U2 ( .INP(n4940), .ZN(U8185_n1) );
  NOR2X0 U8185_U1 ( .IN1(g1046), .IN2(U8185_n1), .QN(n4938) );
  INVX0 U8192_U2 ( .INP(n4915), .ZN(U8192_n1) );
  NOR2X0 U8192_U1 ( .IN1(g1389), .IN2(U8192_n1), .QN(n4913) );
  INVX0 U8210_U2 ( .INP(n422), .ZN(U8210_n1) );
  NOR2X0 U8210_U1 ( .IN1(n1269), .IN2(U8210_n1), .QN(n4714) );
  INVX0 U8223_U2 ( .INP(n4518), .ZN(U8223_n1) );
  NOR2X0 U8223_U1 ( .IN1(n4516), .IN2(U8223_n1), .QN(n4517) );
  INVX0 U8224_U2 ( .INP(n4519), .ZN(U8224_n1) );
  NOR2X0 U8224_U1 ( .IN1(n5728), .IN2(U8224_n1), .QN(n4516) );
  INVX0 U8281_U2 ( .INP(n4819), .ZN(U8281_n1) );
  NOR2X0 U8281_U1 ( .IN1(n11024), .IN2(U8281_n1), .QN(n5111) );
  INVX0 U8307_U2 ( .INP(g29216), .ZN(U8307_n1) );
  NOR2X0 U8307_U1 ( .IN1(n11024), .IN2(U8307_n1), .QN(g26900) );
  INVX0 U8974_U2 ( .INP(n3362), .ZN(U8974_n1) );
  NOR2X0 U8974_U1 ( .IN1(test_so25), .IN2(U8974_n1), .QN(n2552) );
  INVX0 U8975_U2 ( .INP(n3174), .ZN(U8975_n1) );
  NOR2X0 U8975_U1 ( .IN1(g528), .IN2(U8975_n1), .QN(n3195) );
  INVX0 U9065_U2 ( .INP(g4145), .ZN(U9065_n1) );
  NOR2X0 U9065_U1 ( .IN1(n11014), .IN2(U9065_n1), .QN(n4721) );
  INVX0 U9070_U2 ( .INP(g2841), .ZN(U9070_n1) );
  NOR2X0 U9070_U1 ( .IN1(n11024), .IN2(U9070_n1), .QN(n3730) );
  INVX0 U9075_U2 ( .INP(g19), .ZN(U9075_n1) );
  NOR2X0 U9075_U1 ( .IN1(g9), .IN2(U9075_n1), .QN(n3362) );
  INVX0 U9076_U2 ( .INP(g113), .ZN(U9076_n1) );
  NOR2X0 U9076_U1 ( .IN1(n11024), .IN2(U9076_n1), .QN(g25694) );
  INVX0 U9080_U2 ( .INP(n4305), .ZN(U9080_n1) );
  NOR2X0 U9080_U1 ( .IN1(n11024), .IN2(U9080_n1), .QN(g29277) );
  INVX0 U9084_U2 ( .INP(g4423), .ZN(U9084_n1) );
  NOR2X0 U9084_U1 ( .IN1(n11024), .IN2(U9084_n1), .QN(g26953) );
  INVX0 U9085_U2 ( .INP(g64), .ZN(U9085_n1) );
  NOR2X0 U9085_U1 ( .IN1(n11025), .IN2(U9085_n1), .QN(g24212) );
  INVX0 U9086_U2 ( .INP(n4283), .ZN(U9086_n1) );
  NOR2X0 U9086_U1 ( .IN1(n11024), .IN2(U9086_n1), .QN(g29279) );
  INVX0 U9090_U2 ( .INP(g125), .ZN(U9090_n1) );
  NOR2X0 U9090_U1 ( .IN1(n11025), .IN2(U9090_n1), .QN(g25688) );
  INVX0 U9098_U2 ( .INP(g4681), .ZN(U9098_n1) );
  NOR2X0 U9098_U1 ( .IN1(n2774), .IN2(U9098_n1), .QN(g34028) );
  INVX0 U9099_U2 ( .INP(n2595), .ZN(U9099_n1) );
  NOR2X0 U9099_U1 ( .IN1(n2608), .IN2(U9099_n1), .QN(g34449) );
  INVX0 U9101_U2 ( .INP(g6745), .ZN(U9101_n1) );
  NOR2X0 U9101_U1 ( .IN1(n11024), .IN2(U9101_n1), .QN(g26880) );
  INVX0 U9107_U2 ( .INP(n4448), .ZN(U9107_n1) );
  NOR2X0 U9107_U1 ( .IN1(n10633), .IN2(U9107_n1), .QN(n4447) );
  INVX0 U9111_U2 ( .INP(n4403), .ZN(U9111_n1) );
  NOR2X0 U9111_U1 ( .IN1(n10630), .IN2(U9111_n1), .QN(n4402) );
  INVX0 U9116_U2 ( .INP(n1432), .ZN(U9116_n1) );
  NOR2X0 U9116_U1 ( .IN1(n10637), .IN2(U9116_n1), .QN(n4425) );
  INVX0 U9120_U2 ( .INP(n4437), .ZN(U9120_n1) );
  NOR2X0 U9120_U1 ( .IN1(n10627), .IN2(U9120_n1), .QN(n4436) );
  INVX0 U9124_U2 ( .INP(n4392), .ZN(U9124_n1) );
  NOR2X0 U9124_U1 ( .IN1(n10635), .IN2(U9124_n1), .QN(n4391) );
  INVX0 U9128_U2 ( .INP(n4380), .ZN(U9128_n1) );
  NOR2X0 U9128_U1 ( .IN1(n10628), .IN2(U9128_n1), .QN(n4379) );
  INVX0 U9132_U2 ( .INP(n4415), .ZN(U9132_n1) );
  NOR2X0 U9132_U1 ( .IN1(n10636), .IN2(U9132_n1), .QN(n4414) );
  INVX0 U9136_U2 ( .INP(n4459), .ZN(U9136_n1) );
  NOR2X0 U9136_U1 ( .IN1(n1418), .IN2(U9136_n1), .QN(n4458) );
  INVX0 U9315_U2 ( .INP(n5016), .ZN(U9315_n1) );
  NOR2X0 U9315_U1 ( .IN1(n5753), .IN2(U9315_n1), .QN(n5014) );
  INVX0 U9453_U2 ( .INP(n3065), .ZN(U9453_n1) );
  NOR2X0 U9453_U1 ( .IN1(n10631), .IN2(U9453_n1), .QN(n3064) );
  INVX0 U9825_U2 ( .INP(g112), .ZN(U9825_n1) );
  NOR2X0 U9825_U1 ( .IN1(n1770), .IN2(U9825_n1), .QN(n3115) );
  INVX0 U9886_U2 ( .INP(g370), .ZN(U9886_n1) );
  NOR2X0 U9886_U1 ( .IN1(n1192), .IN2(U9886_n1), .QN(n4948) );
  INVX0 U9927_U2 ( .INP(n3933), .ZN(U9927_n1) );
  NOR2X0 U9927_U1 ( .IN1(g4098), .IN2(U9927_n1), .QN(n3833) );
  INVX0 U9953_U2 ( .INP(g671), .ZN(U9953_n1) );
  NOR2X0 U9953_U1 ( .IN1(n154), .IN2(U9953_n1), .QN(n4526) );
  INVX0 U9957_U2 ( .INP(g4843), .ZN(U9957_n1) );
  NOR2X0 U9957_U1 ( .IN1(n5283), .IN2(U9957_n1), .QN(n2563) );
  INVX0 U9958_U2 ( .INP(test_so19), .ZN(U9958_n1) );
  NOR2X0 U9958_U1 ( .IN1(n5656), .IN2(U9958_n1), .QN(n2573) );
  INVX0 U9968_U2 ( .INP(n3084), .ZN(U9968_n1) );
  NOR2X0 U9968_U1 ( .IN1(g4358), .IN2(U9968_n1), .QN(n3023) );
  INVX0 U9972_U2 ( .INP(g681), .ZN(U9972_n1) );
  NOR2X0 U9972_U1 ( .IN1(n4535), .IN2(U9972_n1), .QN(n5112) );
  INVX0 U9992_U2 ( .INP(n3675), .ZN(U9992_n1) );
  NOR2X0 U9992_U1 ( .IN1(n3676), .IN2(U9992_n1), .QN(n2644) );
  INVX0 U10314_U2 ( .INP(g667), .ZN(U10314_n1) );
  NOR2X0 U10314_U1 ( .IN1(g686), .IN2(U10314_n1), .QN(n4962) );
  INVX0 U10318_U2 ( .INP(g5092), .ZN(U10318_n1) );
  NOR2X0 U10318_U1 ( .IN1(n5681), .IN2(U10318_n1), .QN(n5016) );
endmodule

