module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n1359_, new_n595_, new_n1233_, new_n445_, new_n1009_, new_n238_, new_n479_, new_n1105_, new_n1215_, new_n1448_, new_n608_, new_n501_, new_n1157_, new_n1442_, new_n1345_, new_n421_, new_n777_, new_n1433_, new_n1517_, new_n1472_, new_n1048_, new_n885_, new_n439_, new_n1532_, new_n283_, new_n223_, new_n390_, new_n743_, new_n1327_, new_n241_, new_n1535_, new_n566_, new_n641_, new_n339_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n1351_, new_n556_, new_n636_, new_n691_, new_n1024_, new_n670_, new_n456_, new_n1125_, new_n246_, new_n911_, new_n679_, new_n937_, new_n667_, new_n367_, new_n1237_, new_n728_, new_n1479_, new_n1071_, new_n1294_, new_n214_, new_n894_, new_n853_, new_n695_, new_n660_, new_n1311_, new_n526_, new_n908_, new_n552_, new_n678_, new_n342_, new_n706_, new_n649_, new_n1119_, new_n1213_, new_n752_, new_n1524_, new_n1305_, new_n500_, new_n1163_, new_n786_, new_n317_, new_n1188_, new_n1415_, new_n1390_, new_n721_, new_n504_, new_n1414_, new_n742_, new_n892_, new_n1368_, new_n234_, new_n472_, new_n873_, new_n1167_, new_n1530_, new_n1300_, new_n1490_, new_n774_, new_n792_, new_n953_, new_n257_, new_n481_, new_n1265_, new_n1110_, new_n449_, new_n580_, new_n639_, new_n484_, new_n766_, new_n272_, new_n282_, new_n1262_, new_n1212_, new_n1059_, new_n634_, new_n1332_, new_n635_, new_n685_, new_n326_, new_n648_, new_n903_, new_n983_, new_n822_, new_n1406_, new_n1082_, new_n1018_, new_n606_, new_n796_, new_n1054_, new_n655_, new_n1288_, new_n630_, new_n385_, new_n1049_, new_n1330_, new_n694_, new_n461_, new_n1323_, new_n297_, new_n565_, new_n1196_, new_n1366_, new_n511_, new_n303_, new_n325_, new_n1285_, new_n1031_, new_n1216_, new_n1281_, new_n629_, new_n1214_, new_n883_, new_n1005_, new_n321_, new_n324_, new_n960_, new_n1377_, new_n1522_, new_n549_, new_n491_, new_n676_, new_n995_, new_n271_, new_n674_, new_n274_, new_n991_, new_n1044_, new_n1362_, new_n1404_, new_n1443_, new_n1484_, new_n1512_, new_n497_, new_n816_, new_n1355_, new_n568_, new_n420_, new_n876_, new_n423_, new_n498_, new_n496_, new_n1217_, new_n1046_, new_n1182_, new_n708_, new_n206_, new_n1463_, new_n429_, new_n1222_, new_n353_, new_n734_, new_n912_, new_n1424_, new_n1062_, new_n680_, new_n981_, new_n506_, new_n872_, new_n1527_, new_n1275_, new_n1277_, new_n1198_, new_n1428_, new_n1440_, new_n656_, new_n1127_, new_n388_, new_n1028_, new_n483_, new_n1004_, new_n1152_, new_n394_, new_n299_, new_n935_, new_n657_, new_n1150_, new_n652_, new_n582_, new_n1020_, new_n363_, new_n1266_, new_n1113_, new_n785_, new_n1501_, new_n441_, new_n477_, new_n664_, new_n600_, new_n280_, new_n1041_, new_n426_, new_n1036_, new_n235_, new_n398_, new_n301_, new_n1333_, new_n1132_, new_n395_, new_n383_, new_n343_, new_n854_, new_n458_, new_n207_, new_n267_, new_n473_, new_n1147_, new_n1373_, new_n1229_, new_n1422_, new_n1523_, new_n1468_, new_n969_, new_n334_, new_n331_, new_n1234_, new_n835_, new_n1360_, new_n378_, new_n621_, new_n1423_, new_n244_, new_n705_, new_n943_, new_n874_, new_n402_, new_n1321_, new_n1209_, new_n335_, new_n347_, new_n659_, new_n700_, new_n1419_, new_n921_, new_n346_, new_n396_, new_n1315_, new_n1003_, new_n696_, new_n208_, new_n1039_, new_n1507_, new_n1439_, new_n1365_, new_n1239_, new_n528_, new_n952_, new_n1158_, new_n729_, new_n1111_, new_n1413_, new_n1218_, new_n1346_, new_n1201_, new_n559_, new_n1282_, new_n762_, new_n1193_, new_n1437_, new_n1187_, new_n1205_, new_n1154_, new_n1253_, new_n295_, new_n1453_, new_n1256_, new_n628_, new_n1513_, new_n409_, new_n1090_, new_n745_, new_n1489_, new_n553_, new_n1114_, new_n1084_, new_n1061_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n1171_, new_n867_, new_n1032_, new_n901_, new_n276_, new_n688_, new_n1255_, new_n410_, new_n985_, new_n851_, new_n1518_, new_n932_, new_n878_, new_n543_, new_n886_, new_n371_, new_n509_, new_n202_, new_n296_, new_n661_, new_n797_, new_n232_, new_n1358_, new_n724_, new_n1070_, new_n1416_, new_n1109_, new_n261_, new_n672_, new_n1496_, new_n1269_, new_n616_, new_n529_, new_n323_, new_n914_, new_n884_, new_n938_, new_n362_, new_n809_, new_n1142_, new_n604_, new_n1461_, new_n1104_, new_n1511_, new_n571_, new_n1504_, new_n758_, new_n460_, new_n1267_, new_n328_, new_n268_, new_n1466_, new_n1516_, new_n1299_, new_n380_, new_n1477_, new_n1079_, new_n861_, new_n1252_, new_n352_, new_n931_, new_n575_, new_n1493_, new_n562_, new_n944_, new_n1064_, new_n1065_, new_n1118_, new_n493_, new_n547_, new_n1480_, new_n264_, new_n379_, new_n273_, new_n224_, new_n586_, new_n963_, new_n1481_, new_n1325_, new_n993_, new_n1191_, new_n1357_, new_n824_, new_n717_, new_n1455_, new_n403_, new_n868_, new_n1242_, new_n475_, new_n237_, new_n858_, new_n1384_, new_n1343_, new_n936_, new_n1459_, new_n1434_, new_n1016_, new_n411_, new_n673_, new_n1144_, new_n666_, new_n1290_, new_n407_, new_n1519_, new_n1407_, new_n879_, new_n1417_, new_n736_, new_n513_, new_n558_, new_n219_, new_n382_, new_n313_, new_n1370_, new_n239_, new_n718_, new_n1310_, new_n1398_, new_n1126_, new_n546_, new_n612_, new_n1015_, new_n919_, new_n302_, new_n755_, new_n1040_, new_n1509_, new_n544_, new_n615_, new_n722_, new_n856_, new_n415_, new_n1324_, new_n1293_, new_n537_, new_n1336_, new_n345_, new_n499_, new_n533_, new_n255_, new_n1130_, new_n795_, new_n459_, new_n1441_, new_n1122_, new_n1185_, new_n1240_, new_n1510_, new_n354_, new_n1174_, new_n968_, new_n1464_, new_n613_, new_n1508_, new_n337_, new_n1195_, new_n417_, new_n658_, new_n837_, new_n591_, new_n801_, new_n1458_, new_n631_, new_n453_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n1521_, new_n1334_, new_n531_, new_n593_, new_n974_, new_n252_, new_n1248_, new_n751_, new_n1038_, new_n372_, new_n852_, new_n1454_, new_n1474_, new_n1328_, new_n978_, new_n1308_, new_n408_, new_n1430_, new_n470_, new_n213_, new_n769_, new_n433_, new_n871_, new_n1450_, new_n992_, new_n1098_, new_n265_, new_n732_, new_n689_, new_n933_, new_n584_, new_n815_, new_n1492_, new_n1367_, new_n278_, new_n304_, new_n1052_, new_n1425_, new_n857_, new_n1379_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n269_, new_n512_, new_n1471_, new_n1220_, new_n989_, new_n1117_, new_n644_, new_n836_, new_n1116_, new_n904_, new_n1392_, new_n1276_, new_n1444_, new_n913_, new_n327_, new_n681_, new_n594_, new_n561_, new_n495_, new_n927_, new_n431_, new_n1206_, new_n1427_, new_n818_, new_n881_, new_n1268_, new_n1376_, new_n1381_, new_n1534_, new_n684_, new_n640_, new_n1274_, new_n754_, new_n653_, new_n905_, new_n377_, new_n1258_, new_n375_, new_n962_, new_n760_, new_n627_, new_n1391_, new_n1436_, new_n567_, new_n1353_, new_n1033_, new_n576_, new_n831_, new_n791_, new_n1153_, new_n357_, new_n320_, new_n780_, new_n1183_, new_n245_, new_n643_, new_n1316_, new_n1194_, new_n1338_, new_n1460_, new_n1230_, new_n1027_, new_n348_, new_n610_, new_n1369_, new_n843_, new_n322_, new_n703_, new_n698_, new_n1165_, new_n1401_, new_n1259_, new_n226_, new_n1208_, new_n697_, new_n1099_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n1235_, new_n1320_, new_n540_, new_n1149_, new_n1066_, new_n434_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n686_, new_n293_, new_n934_, new_n770_, new_n1389_, new_n1400_, new_n757_, new_n1225_, new_n521_, new_n793_, new_n406_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n1089_, new_n1192_, new_n405_, new_n942_, new_n614_, new_n895_, new_n958_, new_n976_, new_n699_, new_n236_, new_n1405_, new_n1249_, new_n1354_, new_n955_, new_n847_, new_n250_, new_n888_, new_n1505_, new_n288_, new_n1340_, new_n798_, new_n1180_, new_n817_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1361_, new_n941_, new_n1410_, new_n738_, new_n827_, new_n1356_, new_n1363_, new_n1317_, new_n366_, new_n779_, new_n1232_, new_n365_, new_n859_, new_n1211_, new_n1412_, new_n1207_, new_n1176_, new_n1374_, new_n601_, new_n842_, new_n1057_, new_n682_, new_n1075_, new_n812_, new_n266_, new_n821_, new_n542_, new_n548_, new_n669_, new_n1397_, new_n220_, new_n1402_, new_n1313_, new_n1172_, new_n419_, new_n624_, new_n534_, new_n1131_, new_n1120_, new_n819_, new_n637_, new_n451_, new_n489_, new_n804_, new_n1342_, new_n424_, new_n602_, new_n1210_, new_n1060_, new_n1303_, new_n240_, new_n413_, new_n1382_, new_n442_, new_n677_, new_n1487_, new_n642_, new_n211_, new_n1418_, new_n462_, new_n603_, new_n564_, new_n1528_, new_n761_, new_n840_, new_n735_, new_n1283_, new_n898_, new_n799_, new_n1304_, new_n1537_, new_n946_, new_n344_, new_n287_, new_n1108_, new_n1469_, new_n862_, new_n427_, new_n532_, new_n393_, new_n418_, new_n746_, new_n1221_, new_n292_, new_n1264_, new_n215_, new_n1319_, new_n626_, new_n1473_, new_n959_, new_n990_, new_n716_, new_n701_, new_n1238_, new_n1058_, new_n1162_, new_n212_, new_n1278_, new_n902_, new_n364_, new_n832_, new_n414_, new_n1101_, new_n1250_, new_n315_, new_n1482_, new_n1050_, new_n554_, new_n230_, new_n1151_, new_n844_, new_n1302_, new_n281_, new_n430_, new_n482_, new_n849_, new_n1203_, new_n855_, new_n1037_, new_n589_, new_n248_, new_n350_, new_n759_, new_n1083_, new_n1297_, new_n829_, new_n1257_, new_n1306_, new_n988_, new_n478_, new_n1307_, new_n1228_, new_n710_, new_n971_, new_n1486_, new_n361_, new_n764_, new_n906_, new_n683_, new_n1409_, new_n1429_, new_n463_, new_n1372_, new_n510_, new_n966_, new_n351_, new_n1292_, new_n1426_, new_n517_, new_n609_, new_n961_, new_n530_, new_n890_, new_n318_, new_n1006_, new_n622_, new_n702_, new_n833_, new_n715_, new_n811_, new_n1445_, new_n1371_, new_n443_, new_n1086_, new_n956_, new_n763_, new_n486_, new_n466_, new_n262_, new_n218_, new_n1170_, new_n845_, new_n768_, new_n773_, new_n305_, new_n1452_, new_n1051_, new_n899_, new_n1053_, new_n205_, new_n492_, new_n1200_, new_n1533_, new_n650_, new_n750_, new_n887_, new_n254_, new_n355_, new_n926_, new_n432_, new_n925_, new_n875_, new_n256_, new_n1226_, new_n778_, new_n452_, new_n381_, new_n1483_, new_n1219_, new_n920_, new_n1121_, new_n1495_, new_n1341_, new_n820_, new_n1386_, new_n771_, new_n979_, new_n508_, new_n1435_, new_n714_, new_n1280_, new_n1007_, new_n1241_, new_n882_, new_n1145_, new_n929_, new_n986_, new_n1159_, new_n314_, new_n1337_, new_n216_, new_n1348_, new_n917_, new_n1322_, new_n1133_, new_n1177_, new_n646_, new_n538_, new_n1026_, new_n541_, new_n210_, new_n447_, new_n1388_, new_n790_, new_n1081_, new_n311_, new_n587_, new_n1247_, new_n465_, new_n783_, new_n1380_, new_n739_, new_n263_, new_n341_, new_n996_, new_n1318_, new_n846_, new_n915_, new_n488_, new_n524_, new_n349_, new_n848_, new_n277_, new_n1245_, new_n663_, new_n1499_, new_n1497_, new_n579_, new_n286_, new_n1375_, new_n1254_, new_n438_, new_n1344_, new_n939_, new_n1393_, new_n632_, new_n1335_, new_n1364_, new_n671_, new_n965_, new_n1514_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n1202_, new_n1526_, new_n397_, new_n1446_, new_n975_, new_n1199_, new_n399_, new_n596_, new_n945_, new_n870_, new_n805_, new_n1420_, new_n1403_, new_n1115_, new_n1383_, new_n1231_, new_n948_, new_n1055_, new_n1431_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n437_, new_n1085_, new_n359_, new_n794_, new_n457_, new_n1301_, new_n1128_, new_n1002_, new_n1169_, new_n448_, new_n384_, new_n900_, new_n1161_, new_n924_, new_n775_, new_n454_, new_n1034_, new_n1124_, new_n1000_, new_n308_, new_n633_, new_n784_, new_n1273_, new_n1396_, new_n1491_, new_n258_, new_n860_, new_n306_, new_n494_, new_n291_, new_n309_, new_n1160_, new_n1166_, new_n259_, new_n1536_, new_n654_, new_n1456_, new_n713_, new_n880_, new_n1102_, new_n227_, new_n690_, new_n416_, new_n1043_, new_n222_, new_n744_, new_n400_, new_n1175_, new_n1136_, new_n1272_, new_n693_, new_n1287_, new_n1485_, new_n505_, new_n1462_, new_n619_, new_n471_, new_n967_, new_n577_, new_n374_, new_n1135_, new_n376_, new_n1538_, new_n1289_, new_n1271_, new_n1251_, new_n747_, new_n749_, new_n1091_, new_n1095_, new_n310_, new_n275_, new_n998_, new_n1056_, new_n1331_, new_n1094_, new_n839_, new_n485_, new_n578_, new_n525_, new_n918_, new_n940_, new_n810_, new_n808_, new_n1284_, new_n907_, new_n665_, new_n800_, new_n897_, new_n1012_, new_n1387_, new_n719_, new_n869_, new_n1178_, new_n1525_, new_n270_, new_n570_, new_n598_, new_n893_, new_n1063_, new_n520_, new_n1347_, new_n1001_, new_n253_, new_n825_, new_n557_, new_n260_, new_n251_, new_n300_, new_n507_, new_n741_, new_n806_, new_n605_, new_n1224_, new_n1074_, new_n748_, new_n1137_, new_n1286_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n1141_, new_n807_, new_n1326_, new_n592_, new_n726_, new_n1263_, new_n1123_, new_n231_, new_n1080_, new_n583_, new_n617_, new_n1279_, new_n1467_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n916_, new_n428_, new_n487_, new_n675_, new_n1155_, new_n360_, new_n1186_, new_n1261_, new_n225_, new_n1246_, new_n1488_, new_n922_, new_n387_, new_n476_, new_n987_, new_n949_, new_n221_, new_n450_, new_n1394_, new_n243_, new_n1179_, new_n298_, new_n1088_, new_n1146_, new_n569_, new_n555_, new_n468_, new_n977_, new_n1139_, new_n782_, new_n444_, new_n392_, new_n518_, new_n950_, new_n737_, new_n1022_, new_n340_, new_n285_, new_n692_, new_n502_, new_n209_, new_n623_, new_n446_, new_n316_, new_n203_, new_n590_, new_n826_, new_n789_, new_n1476_, new_n515_, new_n332_, new_n972_, new_n1067_, new_n891_, new_n516_, new_n1227_, new_n1352_, new_n733_, new_n1021_, new_n1076_, new_n585_, new_n1350_, new_n312_, new_n535_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n1244_, new_n307_, new_n1378_, new_n1478_, new_n1181_, new_n1093_, new_n597_, new_n1451_, new_n1092_, new_n1143_, new_n1072_, new_n1190_, new_n1097_, new_n1069_, new_n651_, new_n1164_, new_n1296_, new_n435_, new_n1309_, new_n1010_, new_n776_, new_n687_, new_n1029_, new_n370_, new_n1515_, new_n638_, new_n523_, new_n909_, new_n217_, new_n788_, new_n841_, new_n1457_, new_n1204_, new_n1112_, new_n711_, new_n1156_, new_n1298_, new_n731_, new_n599_, new_n930_, new_n1475_, new_n1260_, new_n973_, new_n412_, new_n607_, new_n645_, new_n723_, new_n756_, new_n823_, new_n574_, new_n1500_, new_n928_, new_n319_, new_n1008_, new_n338_, new_n707_, new_n740_, new_n957_, new_n1047_, new_n787_, new_n1134_, new_n336_, new_n1291_, new_n247_, new_n539_, new_n1399_, new_n803_, new_n330_, new_n1270_, new_n727_, new_n1531_, new_n294_, new_n1295_, new_n1173_, new_n704_, new_n1432_, new_n1189_, new_n1197_, new_n1502_, new_n474_, new_n1223_, new_n1129_, new_n1013_, new_n467_, new_n404_, new_n1243_, new_n1077_, new_n490_, new_n560_, new_n1100_, new_n865_, new_n358_, new_n877_, new_n1506_, new_n545_, new_n228_, new_n611_, new_n289_, new_n1011_, new_n425_, new_n896_, new_n802_, new_n1236_, new_n866_, new_n947_, new_n994_, new_n982_, new_n1494_, new_n1449_, new_n964_, new_n1078_, new_n551_, new_n1408_, new_n279_, new_n455_, new_n618_, new_n1140_, new_n1042_, new_n863_, new_n828_, new_n980_, new_n464_, new_n1498_, new_n204_, new_n573_, new_n765_, new_n1314_, new_n1103_;

not g0000 ( new_n202_, keyIn_0_107 );
not g0001 ( new_n203_, N1 );
not g0002 ( new_n204_, keyIn_0_36 );
not g0003 ( new_n205_, N85 );
nand g0004 ( new_n206_, new_n205_, N81 );
not g0005 ( new_n207_, N81 );
nand g0006 ( new_n208_, new_n207_, N85 );
nand g0007 ( new_n209_, new_n206_, new_n208_ );
nand g0008 ( new_n210_, new_n209_, keyIn_0_5 );
not g0009 ( new_n211_, keyIn_0_5 );
not g0010 ( new_n212_, new_n209_ );
nand g0011 ( new_n213_, new_n212_, new_n211_ );
nand g0012 ( new_n214_, new_n213_, new_n210_ );
not g0013 ( new_n215_, keyIn_0_6 );
not g0014 ( new_n216_, N93 );
nand g0015 ( new_n217_, new_n216_, N89 );
not g0016 ( new_n218_, N89 );
nand g0017 ( new_n219_, new_n218_, N93 );
nand g0018 ( new_n220_, new_n217_, new_n219_ );
nor g0019 ( new_n221_, new_n220_, new_n215_ );
nand g0020 ( new_n222_, new_n220_, new_n215_ );
not g0021 ( new_n223_, new_n222_ );
nor g0022 ( new_n224_, new_n223_, new_n221_ );
nand g0023 ( new_n225_, new_n224_, new_n214_ );
not g0024 ( new_n226_, new_n210_ );
nor g0025 ( new_n227_, new_n209_, keyIn_0_5 );
nor g0026 ( new_n228_, new_n226_, new_n227_ );
not g0027 ( new_n229_, new_n220_ );
nand g0028 ( new_n230_, new_n229_, keyIn_0_6 );
nand g0029 ( new_n231_, new_n230_, new_n222_ );
nand g0030 ( new_n232_, new_n228_, new_n231_ );
nand g0031 ( new_n233_, new_n225_, new_n232_ );
nand g0032 ( new_n234_, new_n233_, keyIn_0_28 );
not g0033 ( new_n235_, keyIn_0_28 );
not g0034 ( new_n236_, new_n233_ );
nand g0035 ( new_n237_, new_n236_, new_n235_ );
nand g0036 ( new_n238_, new_n237_, new_n234_ );
not g0037 ( new_n239_, N65 );
nor g0038 ( new_n240_, new_n239_, N69 );
not g0039 ( new_n241_, N69 );
nor g0040 ( new_n242_, new_n241_, N65 );
nor g0041 ( new_n243_, new_n240_, new_n242_ );
not g0042 ( new_n244_, N73 );
nor g0043 ( new_n245_, new_n244_, N77 );
not g0044 ( new_n246_, N77 );
nor g0045 ( new_n247_, new_n246_, N73 );
nor g0046 ( new_n248_, new_n245_, new_n247_ );
not g0047 ( new_n249_, new_n248_ );
nor g0048 ( new_n250_, new_n249_, new_n243_ );
nand g0049 ( new_n251_, new_n249_, new_n243_ );
not g0050 ( new_n252_, new_n251_ );
nor g0051 ( new_n253_, new_n252_, new_n250_ );
not g0052 ( new_n254_, new_n253_ );
nand g0053 ( new_n255_, new_n238_, new_n254_ );
not g0054 ( new_n256_, new_n234_ );
nor g0055 ( new_n257_, new_n233_, keyIn_0_28 );
nor g0056 ( new_n258_, new_n256_, new_n257_ );
nand g0057 ( new_n259_, new_n258_, new_n253_ );
nand g0058 ( new_n260_, new_n259_, new_n255_ );
nand g0059 ( new_n261_, new_n260_, keyIn_0_34 );
not g0060 ( new_n262_, keyIn_0_34 );
nor g0061 ( new_n263_, new_n258_, new_n253_ );
nor g0062 ( new_n264_, new_n238_, new_n254_ );
nor g0063 ( new_n265_, new_n263_, new_n264_ );
nand g0064 ( new_n266_, new_n265_, new_n262_ );
nand g0065 ( new_n267_, new_n266_, new_n261_ );
nand g0066 ( new_n268_, N129, N137 );
nand g0067 ( new_n269_, new_n268_, keyIn_0_9 );
not g0068 ( new_n270_, N129 );
nor g0069 ( new_n271_, new_n270_, keyIn_0_9 );
nand g0070 ( new_n272_, new_n271_, N137 );
nand g0071 ( new_n273_, new_n272_, new_n269_ );
not g0072 ( new_n274_, new_n273_ );
nand g0073 ( new_n275_, new_n267_, new_n274_ );
nor g0074 ( new_n276_, new_n265_, new_n262_ );
nor g0075 ( new_n277_, new_n260_, keyIn_0_34 );
nor g0076 ( new_n278_, new_n276_, new_n277_ );
nand g0077 ( new_n279_, new_n278_, new_n273_ );
nand g0078 ( new_n280_, new_n279_, new_n275_ );
nand g0079 ( new_n281_, new_n280_, new_n204_ );
nor g0080 ( new_n282_, new_n278_, new_n273_ );
nor g0081 ( new_n283_, new_n267_, new_n274_ );
nor g0082 ( new_n284_, new_n282_, new_n283_ );
nand g0083 ( new_n285_, new_n284_, keyIn_0_36 );
nand g0084 ( new_n286_, new_n285_, new_n281_ );
not g0085 ( new_n287_, N33 );
nor g0086 ( new_n288_, new_n287_, N49 );
not g0087 ( new_n289_, N49 );
nor g0088 ( new_n290_, new_n289_, N33 );
nor g0089 ( new_n291_, new_n288_, new_n290_ );
not g0090 ( new_n292_, new_n291_ );
nand g0091 ( new_n293_, new_n292_, keyIn_0_16 );
not g0092 ( new_n294_, new_n293_ );
nor g0093 ( new_n295_, new_n292_, keyIn_0_16 );
nor g0094 ( new_n296_, new_n294_, new_n295_ );
nor g0095 ( new_n297_, new_n203_, N17 );
not g0096 ( new_n298_, N17 );
nor g0097 ( new_n299_, new_n298_, N1 );
nor g0098 ( new_n300_, new_n297_, new_n299_ );
nor g0099 ( new_n301_, new_n296_, new_n300_ );
nand g0100 ( new_n302_, new_n296_, new_n300_ );
not g0101 ( new_n303_, new_n302_ );
nor g0102 ( new_n304_, new_n303_, new_n301_ );
nand g0103 ( new_n305_, new_n286_, new_n304_ );
nor g0104 ( new_n306_, new_n284_, keyIn_0_36 );
nor g0105 ( new_n307_, new_n280_, new_n204_ );
nor g0106 ( new_n308_, new_n306_, new_n307_ );
not g0107 ( new_n309_, new_n304_ );
nand g0108 ( new_n310_, new_n308_, new_n309_ );
nand g0109 ( new_n311_, new_n310_, new_n305_ );
nand g0110 ( new_n312_, new_n311_, keyIn_0_40 );
not g0111 ( new_n313_, keyIn_0_40 );
nor g0112 ( new_n314_, new_n308_, new_n309_ );
nor g0113 ( new_n315_, new_n286_, new_n304_ );
nor g0114 ( new_n316_, new_n314_, new_n315_ );
nand g0115 ( new_n317_, new_n316_, new_n313_ );
nand g0116 ( new_n318_, new_n317_, new_n312_ );
not g0117 ( new_n319_, keyIn_0_72 );
nand g0118 ( new_n320_, new_n318_, keyIn_0_46 );
nor g0119 ( new_n321_, new_n318_, keyIn_0_46 );
not g0120 ( new_n322_, new_n321_ );
nand g0121 ( new_n323_, new_n322_, new_n320_ );
not g0122 ( new_n324_, keyIn_0_35 );
not g0123 ( new_n325_, keyIn_0_7 );
not g0124 ( new_n326_, N109 );
nand g0125 ( new_n327_, new_n326_, N105 );
not g0126 ( new_n328_, N105 );
nand g0127 ( new_n329_, new_n328_, N109 );
nand g0128 ( new_n330_, new_n327_, new_n329_ );
nand g0129 ( new_n331_, new_n330_, new_n325_ );
not g0130 ( new_n332_, new_n331_ );
nor g0131 ( new_n333_, new_n330_, new_n325_ );
nor g0132 ( new_n334_, new_n332_, new_n333_ );
not g0133 ( new_n335_, N97 );
nor g0134 ( new_n336_, new_n335_, N101 );
not g0135 ( new_n337_, N101 );
nor g0136 ( new_n338_, new_n337_, N97 );
nor g0137 ( new_n339_, new_n336_, new_n338_ );
nor g0138 ( new_n340_, new_n334_, new_n339_ );
nand g0139 ( new_n341_, new_n334_, new_n339_ );
not g0140 ( new_n342_, new_n341_ );
nor g0141 ( new_n343_, new_n342_, new_n340_ );
not g0142 ( new_n344_, new_n343_ );
not g0143 ( new_n345_, keyIn_0_8 );
not g0144 ( new_n346_, N125 );
nand g0145 ( new_n347_, new_n346_, N121 );
not g0146 ( new_n348_, N121 );
nand g0147 ( new_n349_, new_n348_, N125 );
nand g0148 ( new_n350_, new_n347_, new_n349_ );
nand g0149 ( new_n351_, new_n350_, new_n345_ );
not g0150 ( new_n352_, new_n351_ );
nor g0151 ( new_n353_, new_n350_, new_n345_ );
nor g0152 ( new_n354_, new_n352_, new_n353_ );
not g0153 ( new_n355_, new_n354_ );
not g0154 ( new_n356_, N113 );
nor g0155 ( new_n357_, new_n356_, N117 );
not g0156 ( new_n358_, N117 );
nor g0157 ( new_n359_, new_n358_, N113 );
nor g0158 ( new_n360_, new_n357_, new_n359_ );
nor g0159 ( new_n361_, new_n355_, new_n360_ );
nand g0160 ( new_n362_, new_n355_, new_n360_ );
not g0161 ( new_n363_, new_n362_ );
nor g0162 ( new_n364_, new_n363_, new_n361_ );
nand g0163 ( new_n365_, new_n364_, new_n344_ );
not g0164 ( new_n366_, new_n364_ );
nand g0165 ( new_n367_, new_n366_, new_n343_ );
nand g0166 ( new_n368_, new_n367_, new_n365_ );
nand g0167 ( new_n369_, new_n368_, new_n324_ );
nor g0168 ( new_n370_, new_n368_, new_n324_ );
not g0169 ( new_n371_, new_n370_ );
nand g0170 ( new_n372_, new_n371_, new_n369_ );
nand g0171 ( new_n373_, new_n372_, keyIn_0_10 );
not g0172 ( new_n374_, keyIn_0_10 );
not g0173 ( new_n375_, new_n369_ );
nor g0174 ( new_n376_, new_n375_, new_n370_ );
nand g0175 ( new_n377_, new_n376_, new_n374_ );
nand g0176 ( new_n378_, new_n377_, new_n373_ );
nand g0177 ( new_n379_, N130, N137 );
nand g0178 ( new_n380_, new_n378_, new_n379_ );
not g0179 ( new_n381_, new_n378_ );
not g0180 ( new_n382_, new_n379_ );
nand g0181 ( new_n383_, new_n381_, new_n382_ );
nand g0182 ( new_n384_, new_n383_, new_n380_ );
not g0183 ( new_n385_, N5 );
nor g0184 ( new_n386_, new_n385_, N21 );
not g0185 ( new_n387_, N21 );
nor g0186 ( new_n388_, new_n387_, N5 );
nor g0187 ( new_n389_, new_n386_, new_n388_ );
not g0188 ( new_n390_, new_n389_ );
nand g0189 ( new_n391_, new_n390_, keyIn_0_17 );
not g0190 ( new_n392_, new_n391_ );
nor g0191 ( new_n393_, new_n390_, keyIn_0_17 );
nor g0192 ( new_n394_, new_n392_, new_n393_ );
not g0193 ( new_n395_, N37 );
nor g0194 ( new_n396_, new_n395_, N53 );
not g0195 ( new_n397_, N53 );
nor g0196 ( new_n398_, new_n397_, N37 );
nor g0197 ( new_n399_, new_n396_, new_n398_ );
not g0198 ( new_n400_, new_n399_ );
nand g0199 ( new_n401_, new_n400_, keyIn_0_18 );
not g0200 ( new_n402_, new_n401_ );
nor g0201 ( new_n403_, new_n400_, keyIn_0_18 );
nor g0202 ( new_n404_, new_n402_, new_n403_ );
not g0203 ( new_n405_, new_n404_ );
nor g0204 ( new_n406_, new_n405_, new_n394_ );
nand g0205 ( new_n407_, new_n405_, new_n394_ );
not g0206 ( new_n408_, new_n407_ );
nor g0207 ( new_n409_, new_n408_, new_n406_ );
nand g0208 ( new_n410_, new_n384_, new_n409_ );
not g0209 ( new_n411_, new_n380_ );
nor g0210 ( new_n412_, new_n378_, new_n379_ );
nor g0211 ( new_n413_, new_n411_, new_n412_ );
not g0212 ( new_n414_, new_n409_ );
nand g0213 ( new_n415_, new_n413_, new_n414_ );
nand g0214 ( new_n416_, new_n415_, new_n410_ );
not g0215 ( new_n417_, new_n416_ );
nor g0216 ( new_n418_, new_n417_, keyIn_0_47 );
nand g0217 ( new_n419_, new_n417_, keyIn_0_47 );
not g0218 ( new_n420_, new_n419_ );
nor g0219 ( new_n421_, new_n420_, new_n418_ );
nand g0220 ( new_n422_, new_n238_, new_n366_ );
nand g0221 ( new_n423_, new_n258_, new_n364_ );
nand g0222 ( new_n424_, new_n423_, new_n422_ );
nand g0223 ( new_n425_, N132, N137 );
nand g0224 ( new_n426_, new_n425_, keyIn_0_12 );
not g0225 ( new_n427_, N132 );
nor g0226 ( new_n428_, new_n427_, keyIn_0_12 );
nand g0227 ( new_n429_, new_n428_, N137 );
nand g0228 ( new_n430_, new_n429_, new_n426_ );
nand g0229 ( new_n431_, new_n424_, new_n430_ );
nor g0230 ( new_n432_, new_n258_, new_n364_ );
nor g0231 ( new_n433_, new_n238_, new_n366_ );
nor g0232 ( new_n434_, new_n432_, new_n433_ );
not g0233 ( new_n435_, new_n430_ );
nand g0234 ( new_n436_, new_n434_, new_n435_ );
nand g0235 ( new_n437_, new_n436_, new_n431_ );
nand g0236 ( new_n438_, new_n437_, keyIn_0_37 );
not g0237 ( new_n439_, keyIn_0_37 );
not g0238 ( new_n440_, new_n431_ );
nor g0239 ( new_n441_, new_n424_, new_n430_ );
nor g0240 ( new_n442_, new_n440_, new_n441_ );
nand g0241 ( new_n443_, new_n442_, new_n439_ );
nand g0242 ( new_n444_, new_n443_, new_n438_ );
not g0243 ( new_n445_, keyIn_0_30 );
not g0244 ( new_n446_, N13 );
nor g0245 ( new_n447_, new_n446_, N29 );
not g0246 ( new_n448_, N29 );
nor g0247 ( new_n449_, new_n448_, N13 );
nor g0248 ( new_n450_, new_n447_, new_n449_ );
not g0249 ( new_n451_, new_n450_ );
nand g0250 ( new_n452_, new_n451_, keyIn_0_20 );
not g0251 ( new_n453_, new_n452_ );
nor g0252 ( new_n454_, new_n451_, keyIn_0_20 );
nor g0253 ( new_n455_, new_n453_, new_n454_ );
not g0254 ( new_n456_, N45 );
nor g0255 ( new_n457_, new_n456_, N61 );
not g0256 ( new_n458_, N61 );
nor g0257 ( new_n459_, new_n458_, N45 );
nor g0258 ( new_n460_, new_n457_, new_n459_ );
not g0259 ( new_n461_, new_n460_ );
nor g0260 ( new_n462_, new_n455_, new_n461_ );
nand g0261 ( new_n463_, new_n455_, new_n461_ );
not g0262 ( new_n464_, new_n463_ );
nor g0263 ( new_n465_, new_n464_, new_n462_ );
nor g0264 ( new_n466_, new_n465_, new_n445_ );
nand g0265 ( new_n467_, new_n465_, new_n445_ );
not g0266 ( new_n468_, new_n467_ );
nor g0267 ( new_n469_, new_n468_, new_n466_ );
nand g0268 ( new_n470_, new_n444_, new_n469_ );
not g0269 ( new_n471_, new_n438_ );
nor g0270 ( new_n472_, new_n437_, keyIn_0_37 );
nor g0271 ( new_n473_, new_n471_, new_n472_ );
not g0272 ( new_n474_, new_n469_ );
nand g0273 ( new_n475_, new_n473_, new_n474_ );
nand g0274 ( new_n476_, new_n475_, new_n470_ );
nand g0275 ( new_n477_, new_n476_, keyIn_0_41 );
not g0276 ( new_n478_, keyIn_0_41 );
not g0277 ( new_n479_, new_n470_ );
nor g0278 ( new_n480_, new_n444_, new_n469_ );
nor g0279 ( new_n481_, new_n479_, new_n480_ );
nand g0280 ( new_n482_, new_n481_, new_n478_ );
nand g0281 ( new_n483_, new_n482_, new_n477_ );
not g0282 ( new_n484_, new_n483_ );
not g0283 ( new_n485_, keyIn_0_48 );
not g0284 ( new_n486_, keyIn_0_11 );
nor g0285 ( new_n487_, new_n343_, new_n254_ );
nor g0286 ( new_n488_, new_n344_, new_n253_ );
nor g0287 ( new_n489_, new_n488_, new_n487_ );
nor g0288 ( new_n490_, new_n489_, new_n486_ );
nand g0289 ( new_n491_, new_n489_, new_n486_ );
not g0290 ( new_n492_, new_n491_ );
nor g0291 ( new_n493_, new_n492_, new_n490_ );
not g0292 ( new_n494_, new_n493_ );
nand g0293 ( new_n495_, N131, N137 );
nand g0294 ( new_n496_, new_n494_, new_n495_ );
not g0295 ( new_n497_, new_n495_ );
nand g0296 ( new_n498_, new_n493_, new_n497_ );
nand g0297 ( new_n499_, new_n496_, new_n498_ );
not g0298 ( new_n500_, N41 );
nor g0299 ( new_n501_, new_n500_, N57 );
not g0300 ( new_n502_, N57 );
nor g0301 ( new_n503_, new_n502_, N41 );
nor g0302 ( new_n504_, new_n501_, new_n503_ );
not g0303 ( new_n505_, new_n504_ );
nand g0304 ( new_n506_, new_n505_, keyIn_0_19 );
not g0305 ( new_n507_, new_n506_ );
nor g0306 ( new_n508_, new_n505_, keyIn_0_19 );
nor g0307 ( new_n509_, new_n507_, new_n508_ );
not g0308 ( new_n510_, N9 );
nor g0309 ( new_n511_, new_n510_, N25 );
not g0310 ( new_n512_, N25 );
nor g0311 ( new_n513_, new_n512_, N9 );
nor g0312 ( new_n514_, new_n511_, new_n513_ );
not g0313 ( new_n515_, new_n514_ );
nor g0314 ( new_n516_, new_n509_, new_n515_ );
nand g0315 ( new_n517_, new_n509_, new_n515_ );
not g0316 ( new_n518_, new_n517_ );
nor g0317 ( new_n519_, new_n518_, new_n516_ );
nor g0318 ( new_n520_, new_n519_, keyIn_0_29 );
nand g0319 ( new_n521_, new_n519_, keyIn_0_29 );
not g0320 ( new_n522_, new_n521_ );
nor g0321 ( new_n523_, new_n522_, new_n520_ );
not g0322 ( new_n524_, new_n523_ );
nand g0323 ( new_n525_, new_n499_, new_n524_ );
nor g0324 ( new_n526_, new_n499_, new_n524_ );
not g0325 ( new_n527_, new_n526_ );
nand g0326 ( new_n528_, new_n527_, new_n525_ );
nor g0327 ( new_n529_, new_n528_, new_n485_ );
not g0328 ( new_n530_, new_n525_ );
nor g0329 ( new_n531_, new_n530_, new_n526_ );
nor g0330 ( new_n532_, new_n531_, keyIn_0_48 );
nor g0331 ( new_n533_, new_n532_, new_n529_ );
not g0332 ( new_n534_, new_n533_ );
nand g0333 ( new_n535_, new_n534_, new_n484_ );
nor g0334 ( new_n536_, new_n421_, new_n535_ );
nand g0335 ( new_n537_, new_n323_, new_n536_ );
nand g0336 ( new_n538_, new_n537_, new_n319_ );
nor g0337 ( new_n539_, new_n537_, new_n319_ );
not g0338 ( new_n540_, new_n539_ );
nand g0339 ( new_n541_, new_n540_, new_n538_ );
not g0340 ( new_n542_, keyIn_0_73 );
nand g0341 ( new_n543_, new_n318_, keyIn_0_49 );
not g0342 ( new_n544_, keyIn_0_49 );
nor g0343 ( new_n545_, new_n316_, new_n313_ );
nor g0344 ( new_n546_, new_n311_, keyIn_0_40 );
nor g0345 ( new_n547_, new_n545_, new_n546_ );
nand g0346 ( new_n548_, new_n547_, new_n544_ );
nand g0347 ( new_n549_, new_n548_, new_n543_ );
nand g0348 ( new_n550_, new_n483_, new_n528_ );
not g0349 ( new_n551_, keyIn_0_50 );
nor g0350 ( new_n552_, new_n416_, new_n551_ );
nor g0351 ( new_n553_, new_n417_, keyIn_0_50 );
nor g0352 ( new_n554_, new_n553_, new_n552_ );
nor g0353 ( new_n555_, new_n554_, new_n550_ );
nand g0354 ( new_n556_, new_n549_, new_n555_ );
nand g0355 ( new_n557_, new_n556_, new_n542_ );
not g0356 ( new_n558_, new_n557_ );
nor g0357 ( new_n559_, new_n556_, new_n542_ );
nor g0358 ( new_n560_, new_n558_, new_n559_ );
nand g0359 ( new_n561_, new_n318_, new_n416_ );
not g0360 ( new_n562_, new_n561_ );
nand g0361 ( new_n563_, new_n483_, keyIn_0_52 );
not g0362 ( new_n564_, new_n563_ );
not g0363 ( new_n565_, keyIn_0_51 );
nor g0364 ( new_n566_, new_n528_, new_n565_ );
nor g0365 ( new_n567_, new_n531_, keyIn_0_51 );
nor g0366 ( new_n568_, new_n567_, new_n566_ );
not g0367 ( new_n569_, new_n568_ );
not g0368 ( new_n570_, keyIn_0_52 );
nand g0369 ( new_n571_, new_n484_, new_n570_ );
nand g0370 ( new_n572_, new_n571_, new_n569_ );
nor g0371 ( new_n573_, new_n572_, new_n564_ );
nand g0372 ( new_n574_, new_n562_, new_n573_ );
nor g0373 ( new_n575_, new_n574_, keyIn_0_74 );
not g0374 ( new_n576_, new_n575_ );
not g0375 ( new_n577_, keyIn_0_74 );
nor g0376 ( new_n578_, new_n483_, keyIn_0_52 );
nor g0377 ( new_n579_, new_n578_, new_n568_ );
nand g0378 ( new_n580_, new_n579_, new_n563_ );
nor g0379 ( new_n581_, new_n580_, new_n561_ );
nor g0380 ( new_n582_, new_n581_, new_n577_ );
not g0381 ( new_n583_, keyIn_0_75 );
nor g0382 ( new_n584_, new_n416_, new_n528_ );
nand g0383 ( new_n585_, new_n584_, new_n483_ );
nor g0384 ( new_n586_, new_n318_, new_n585_ );
nor g0385 ( new_n587_, new_n586_, new_n583_ );
not g0386 ( new_n588_, new_n585_ );
nand g0387 ( new_n589_, new_n547_, new_n588_ );
nor g0388 ( new_n590_, new_n589_, keyIn_0_75 );
nor g0389 ( new_n591_, new_n590_, new_n587_ );
nor g0390 ( new_n592_, new_n591_, new_n582_ );
nand g0391 ( new_n593_, new_n592_, new_n576_ );
nor g0392 ( new_n594_, new_n560_, new_n593_ );
nand g0393 ( new_n595_, new_n594_, new_n541_ );
nand g0394 ( new_n596_, new_n595_, keyIn_0_78 );
not g0395 ( new_n597_, keyIn_0_78 );
not g0396 ( new_n598_, new_n538_ );
nor g0397 ( new_n599_, new_n598_, new_n539_ );
not g0398 ( new_n600_, new_n556_ );
nand g0399 ( new_n601_, new_n600_, keyIn_0_73 );
nand g0400 ( new_n602_, new_n601_, new_n557_ );
nand g0401 ( new_n603_, new_n574_, keyIn_0_74 );
nand g0402 ( new_n604_, new_n589_, keyIn_0_75 );
nand g0403 ( new_n605_, new_n586_, new_n583_ );
nand g0404 ( new_n606_, new_n604_, new_n605_ );
nand g0405 ( new_n607_, new_n603_, new_n606_ );
nor g0406 ( new_n608_, new_n607_, new_n575_ );
nand g0407 ( new_n609_, new_n602_, new_n608_ );
nor g0408 ( new_n610_, new_n609_, new_n599_ );
nand g0409 ( new_n611_, new_n610_, new_n597_ );
nand g0410 ( new_n612_, new_n596_, new_n611_ );
not g0411 ( new_n613_, keyIn_0_53 );
not g0412 ( new_n614_, keyIn_0_43 );
not g0413 ( new_n615_, keyIn_0_1 );
nor g0414 ( new_n616_, new_n287_, N37 );
nor g0415 ( new_n617_, new_n395_, N33 );
nor g0416 ( new_n618_, new_n616_, new_n617_ );
not g0417 ( new_n619_, new_n618_ );
nand g0418 ( new_n620_, new_n619_, new_n615_ );
nand g0419 ( new_n621_, new_n618_, keyIn_0_1 );
nand g0420 ( new_n622_, new_n620_, new_n621_ );
not g0421 ( new_n623_, keyIn_0_2 );
nor g0422 ( new_n624_, new_n500_, N45 );
not g0423 ( new_n625_, new_n624_ );
nor g0424 ( new_n626_, new_n456_, N41 );
not g0425 ( new_n627_, new_n626_ );
nand g0426 ( new_n628_, new_n625_, new_n627_ );
nand g0427 ( new_n629_, new_n628_, new_n623_ );
nor g0428 ( new_n630_, new_n628_, new_n623_ );
not g0429 ( new_n631_, new_n630_ );
nand g0430 ( new_n632_, new_n631_, new_n629_ );
nand g0431 ( new_n633_, new_n632_, new_n622_ );
not g0432 ( new_n634_, new_n622_ );
not g0433 ( new_n635_, new_n629_ );
nor g0434 ( new_n636_, new_n635_, new_n630_ );
nand g0435 ( new_n637_, new_n634_, new_n636_ );
nand g0436 ( new_n638_, new_n637_, new_n633_ );
nand g0437 ( new_n639_, new_n638_, keyIn_0_26 );
not g0438 ( new_n640_, new_n639_ );
nor g0439 ( new_n641_, new_n638_, keyIn_0_26 );
nor g0440 ( new_n642_, new_n640_, new_n641_ );
not g0441 ( new_n643_, keyIn_0_27 );
nor g0442 ( new_n644_, new_n502_, N61 );
not g0443 ( new_n645_, new_n644_ );
nor g0444 ( new_n646_, new_n458_, N57 );
not g0445 ( new_n647_, new_n646_ );
nand g0446 ( new_n648_, new_n645_, new_n647_ );
nand g0447 ( new_n649_, new_n648_, keyIn_0_4 );
nor g0448 ( new_n650_, new_n648_, keyIn_0_4 );
not g0449 ( new_n651_, new_n650_ );
nand g0450 ( new_n652_, new_n651_, new_n649_ );
not g0451 ( new_n653_, keyIn_0_3 );
nor g0452 ( new_n654_, new_n289_, N53 );
not g0453 ( new_n655_, new_n654_ );
nor g0454 ( new_n656_, new_n397_, N49 );
not g0455 ( new_n657_, new_n656_ );
nand g0456 ( new_n658_, new_n655_, new_n657_ );
nand g0457 ( new_n659_, new_n658_, new_n653_ );
not g0458 ( new_n660_, new_n658_ );
nand g0459 ( new_n661_, new_n660_, keyIn_0_3 );
nand g0460 ( new_n662_, new_n661_, new_n659_ );
nand g0461 ( new_n663_, new_n652_, new_n662_ );
not g0462 ( new_n664_, new_n649_ );
nor g0463 ( new_n665_, new_n664_, new_n650_ );
not g0464 ( new_n666_, new_n659_ );
nor g0465 ( new_n667_, new_n658_, new_n653_ );
nor g0466 ( new_n668_, new_n666_, new_n667_ );
nand g0467 ( new_n669_, new_n665_, new_n668_ );
nand g0468 ( new_n670_, new_n669_, new_n663_ );
nand g0469 ( new_n671_, new_n670_, new_n643_ );
not g0470 ( new_n672_, new_n670_ );
nand g0471 ( new_n673_, new_n672_, keyIn_0_27 );
nand g0472 ( new_n674_, new_n673_, new_n671_ );
nand g0473 ( new_n675_, new_n642_, new_n674_ );
not g0474 ( new_n676_, keyIn_0_26 );
not g0475 ( new_n677_, new_n638_ );
nand g0476 ( new_n678_, new_n677_, new_n676_ );
nand g0477 ( new_n679_, new_n678_, new_n639_ );
not g0478 ( new_n680_, new_n671_ );
nor g0479 ( new_n681_, new_n670_, new_n643_ );
nor g0480 ( new_n682_, new_n680_, new_n681_ );
nand g0481 ( new_n683_, new_n682_, new_n679_ );
nand g0482 ( new_n684_, new_n675_, new_n683_ );
nand g0483 ( new_n685_, new_n684_, keyIn_0_33 );
not g0484 ( new_n686_, new_n685_ );
nor g0485 ( new_n687_, new_n684_, keyIn_0_33 );
nor g0486 ( new_n688_, new_n686_, new_n687_ );
not g0487 ( new_n689_, keyIn_0_14 );
nand g0488 ( new_n690_, N134, N137 );
nand g0489 ( new_n691_, new_n690_, new_n689_ );
not g0490 ( new_n692_, new_n691_ );
not g0491 ( new_n693_, N137 );
nand g0492 ( new_n694_, keyIn_0_14, N134 );
nor g0493 ( new_n695_, new_n694_, new_n693_ );
nor g0494 ( new_n696_, new_n692_, new_n695_ );
nor g0495 ( new_n697_, new_n688_, new_n696_ );
not g0496 ( new_n698_, keyIn_0_33 );
not g0497 ( new_n699_, new_n684_ );
nand g0498 ( new_n700_, new_n699_, new_n698_ );
nand g0499 ( new_n701_, new_n700_, new_n685_ );
not g0500 ( new_n702_, new_n696_ );
nor g0501 ( new_n703_, new_n701_, new_n702_ );
nor g0502 ( new_n704_, new_n697_, new_n703_ );
nor g0503 ( new_n705_, new_n704_, keyIn_0_39 );
not g0504 ( new_n706_, keyIn_0_39 );
nand g0505 ( new_n707_, new_n701_, new_n702_ );
nand g0506 ( new_n708_, new_n688_, new_n696_ );
nand g0507 ( new_n709_, new_n708_, new_n707_ );
nor g0508 ( new_n710_, new_n709_, new_n706_ );
nor g0509 ( new_n711_, new_n705_, new_n710_ );
not g0510 ( new_n712_, keyIn_0_23 );
nor g0511 ( new_n713_, new_n241_, N85 );
nor g0512 ( new_n714_, new_n205_, N69 );
nor g0513 ( new_n715_, new_n713_, new_n714_ );
not g0514 ( new_n716_, new_n715_ );
nand g0515 ( new_n717_, new_n716_, new_n712_ );
not g0516 ( new_n718_, new_n717_ );
nor g0517 ( new_n719_, new_n716_, new_n712_ );
nor g0518 ( new_n720_, new_n718_, new_n719_ );
not g0519 ( new_n721_, keyIn_0_24 );
nor g0520 ( new_n722_, new_n337_, N117 );
nor g0521 ( new_n723_, new_n358_, N101 );
nor g0522 ( new_n724_, new_n722_, new_n723_ );
not g0523 ( new_n725_, new_n724_ );
nand g0524 ( new_n726_, new_n725_, new_n721_ );
not g0525 ( new_n727_, new_n726_ );
nor g0526 ( new_n728_, new_n725_, new_n721_ );
nor g0527 ( new_n729_, new_n727_, new_n728_ );
nor g0528 ( new_n730_, new_n720_, new_n729_ );
nand g0529 ( new_n731_, new_n720_, new_n729_ );
not g0530 ( new_n732_, new_n731_ );
nor g0531 ( new_n733_, new_n732_, new_n730_ );
not g0532 ( new_n734_, new_n733_ );
nand g0533 ( new_n735_, new_n711_, new_n734_ );
nand g0534 ( new_n736_, new_n709_, new_n706_ );
nand g0535 ( new_n737_, new_n704_, keyIn_0_39 );
nand g0536 ( new_n738_, new_n737_, new_n736_ );
nand g0537 ( new_n739_, new_n738_, new_n733_ );
nand g0538 ( new_n740_, new_n735_, new_n739_ );
nand g0539 ( new_n741_, new_n740_, new_n614_ );
nor g0540 ( new_n742_, new_n738_, new_n733_ );
nor g0541 ( new_n743_, new_n711_, new_n734_ );
nor g0542 ( new_n744_, new_n743_, new_n742_ );
nand g0543 ( new_n745_, new_n744_, keyIn_0_43 );
nand g0544 ( new_n746_, new_n745_, new_n741_ );
nor g0545 ( new_n747_, new_n746_, new_n613_ );
not g0546 ( new_n748_, new_n741_ );
nor g0547 ( new_n749_, new_n740_, new_n614_ );
nor g0548 ( new_n750_, new_n748_, new_n749_ );
nor g0549 ( new_n751_, new_n750_, keyIn_0_53 );
nor g0550 ( new_n752_, new_n751_, new_n747_ );
not g0551 ( new_n753_, keyIn_0_25 );
nor g0552 ( new_n754_, new_n298_, N21 );
not g0553 ( new_n755_, new_n754_ );
nor g0554 ( new_n756_, new_n387_, N17 );
not g0555 ( new_n757_, new_n756_ );
nand g0556 ( new_n758_, new_n755_, new_n757_ );
nand g0557 ( new_n759_, new_n758_, keyIn_0_0 );
not g0558 ( new_n760_, keyIn_0_0 );
not g0559 ( new_n761_, new_n758_ );
nand g0560 ( new_n762_, new_n761_, new_n760_ );
nand g0561 ( new_n763_, new_n762_, new_n759_ );
nor g0562 ( new_n764_, new_n512_, N29 );
nor g0563 ( new_n765_, new_n448_, N25 );
nor g0564 ( new_n766_, new_n764_, new_n765_ );
nand g0565 ( new_n767_, new_n763_, new_n766_ );
not g0566 ( new_n768_, new_n759_ );
nor g0567 ( new_n769_, new_n758_, keyIn_0_0 );
nor g0568 ( new_n770_, new_n768_, new_n769_ );
not g0569 ( new_n771_, new_n766_ );
nand g0570 ( new_n772_, new_n770_, new_n771_ );
nand g0571 ( new_n773_, new_n772_, new_n767_ );
nand g0572 ( new_n774_, new_n773_, new_n753_ );
nor g0573 ( new_n775_, new_n770_, new_n771_ );
nor g0574 ( new_n776_, new_n763_, new_n766_ );
nor g0575 ( new_n777_, new_n775_, new_n776_ );
nand g0576 ( new_n778_, new_n777_, keyIn_0_25 );
nand g0577 ( new_n779_, new_n778_, new_n774_ );
nand g0578 ( new_n780_, new_n674_, new_n779_ );
not g0579 ( new_n781_, new_n774_ );
nor g0580 ( new_n782_, new_n773_, new_n753_ );
nor g0581 ( new_n783_, new_n781_, new_n782_ );
nand g0582 ( new_n784_, new_n682_, new_n783_ );
nand g0583 ( new_n785_, new_n784_, new_n780_ );
nand g0584 ( new_n786_, new_n785_, keyIn_0_15 );
not g0585 ( new_n787_, keyIn_0_15 );
nor g0586 ( new_n788_, new_n682_, new_n783_ );
nor g0587 ( new_n789_, new_n674_, new_n779_ );
nor g0588 ( new_n790_, new_n788_, new_n789_ );
nand g0589 ( new_n791_, new_n790_, new_n787_ );
nand g0590 ( new_n792_, new_n791_, new_n786_ );
nand g0591 ( new_n793_, N136, N137 );
nand g0592 ( new_n794_, new_n792_, new_n793_ );
not g0593 ( new_n795_, new_n786_ );
nor g0594 ( new_n796_, new_n785_, keyIn_0_15 );
nor g0595 ( new_n797_, new_n795_, new_n796_ );
not g0596 ( new_n798_, new_n793_ );
nand g0597 ( new_n799_, new_n797_, new_n798_ );
nand g0598 ( new_n800_, new_n799_, new_n794_ );
not g0599 ( new_n801_, keyIn_0_32 );
nor g0600 ( new_n802_, new_n246_, N93 );
nor g0601 ( new_n803_, new_n216_, N77 );
nor g0602 ( new_n804_, new_n802_, new_n803_ );
nor g0603 ( new_n805_, new_n326_, N125 );
nor g0604 ( new_n806_, new_n346_, N109 );
nor g0605 ( new_n807_, new_n805_, new_n806_ );
not g0606 ( new_n808_, new_n807_ );
nor g0607 ( new_n809_, new_n808_, new_n804_ );
nand g0608 ( new_n810_, new_n808_, new_n804_ );
not g0609 ( new_n811_, new_n810_ );
nor g0610 ( new_n812_, new_n811_, new_n809_ );
not g0611 ( new_n813_, new_n812_ );
nand g0612 ( new_n814_, new_n813_, new_n801_ );
not g0613 ( new_n815_, new_n814_ );
nor g0614 ( new_n816_, new_n813_, new_n801_ );
nor g0615 ( new_n817_, new_n815_, new_n816_ );
not g0616 ( new_n818_, new_n817_ );
nand g0617 ( new_n819_, new_n800_, new_n818_ );
nor g0618 ( new_n820_, new_n797_, new_n798_ );
nor g0619 ( new_n821_, new_n792_, new_n793_ );
nor g0620 ( new_n822_, new_n820_, new_n821_ );
nand g0621 ( new_n823_, new_n822_, new_n817_ );
nand g0622 ( new_n824_, new_n823_, new_n819_ );
nand g0623 ( new_n825_, new_n824_, keyIn_0_45 );
not g0624 ( new_n826_, new_n825_ );
nor g0625 ( new_n827_, new_n824_, keyIn_0_45 );
nor g0626 ( new_n828_, new_n826_, new_n827_ );
nor g0627 ( new_n829_, new_n828_, keyIn_0_54 );
nand g0628 ( new_n830_, new_n828_, keyIn_0_54 );
not g0629 ( new_n831_, keyIn_0_38 );
nor g0630 ( new_n832_, new_n203_, N5 );
nor g0631 ( new_n833_, new_n385_, N1 );
nor g0632 ( new_n834_, new_n832_, new_n833_ );
nor g0633 ( new_n835_, new_n510_, N13 );
nor g0634 ( new_n836_, new_n446_, N9 );
nor g0635 ( new_n837_, new_n835_, new_n836_ );
not g0636 ( new_n838_, new_n837_ );
nor g0637 ( new_n839_, new_n838_, new_n834_ );
nand g0638 ( new_n840_, new_n838_, new_n834_ );
not g0639 ( new_n841_, new_n840_ );
nor g0640 ( new_n842_, new_n841_, new_n839_ );
not g0641 ( new_n843_, new_n842_ );
nand g0642 ( new_n844_, new_n779_, new_n843_ );
nor g0643 ( new_n845_, new_n779_, new_n843_ );
not g0644 ( new_n846_, new_n845_ );
nand g0645 ( new_n847_, new_n846_, new_n844_ );
not g0646 ( new_n848_, keyIn_0_13 );
nand g0647 ( new_n849_, N133, N137 );
nand g0648 ( new_n850_, new_n849_, new_n848_ );
not g0649 ( new_n851_, new_n850_ );
nand g0650 ( new_n852_, keyIn_0_13, N133 );
nor g0651 ( new_n853_, new_n852_, new_n693_ );
nor g0652 ( new_n854_, new_n851_, new_n853_ );
not g0653 ( new_n855_, new_n854_ );
nand g0654 ( new_n856_, new_n847_, new_n855_ );
not g0655 ( new_n857_, new_n844_ );
nor g0656 ( new_n858_, new_n857_, new_n845_ );
nand g0657 ( new_n859_, new_n858_, new_n854_ );
nand g0658 ( new_n860_, new_n859_, new_n856_ );
nand g0659 ( new_n861_, new_n860_, new_n831_ );
nor g0660 ( new_n862_, new_n858_, new_n854_ );
nor g0661 ( new_n863_, new_n847_, new_n855_ );
nor g0662 ( new_n864_, new_n862_, new_n863_ );
nand g0663 ( new_n865_, new_n864_, keyIn_0_38 );
nand g0664 ( new_n866_, new_n865_, new_n861_ );
not g0665 ( new_n867_, keyIn_0_21 );
nor g0666 ( new_n868_, new_n239_, N81 );
nor g0667 ( new_n869_, new_n207_, N65 );
nor g0668 ( new_n870_, new_n868_, new_n869_ );
not g0669 ( new_n871_, new_n870_ );
nand g0670 ( new_n872_, new_n871_, new_n867_ );
not g0671 ( new_n873_, new_n872_ );
nor g0672 ( new_n874_, new_n871_, new_n867_ );
nor g0673 ( new_n875_, new_n873_, new_n874_ );
nor g0674 ( new_n876_, new_n335_, N113 );
nor g0675 ( new_n877_, new_n356_, N97 );
nor g0676 ( new_n878_, new_n876_, new_n877_ );
not g0677 ( new_n879_, new_n878_ );
nand g0678 ( new_n880_, new_n879_, keyIn_0_22 );
not g0679 ( new_n881_, new_n880_ );
nor g0680 ( new_n882_, new_n879_, keyIn_0_22 );
nor g0681 ( new_n883_, new_n881_, new_n882_ );
nor g0682 ( new_n884_, new_n875_, new_n883_ );
nand g0683 ( new_n885_, new_n875_, new_n883_ );
not g0684 ( new_n886_, new_n885_ );
nor g0685 ( new_n887_, new_n886_, new_n884_ );
not g0686 ( new_n888_, new_n887_ );
nand g0687 ( new_n889_, new_n866_, new_n888_ );
not g0688 ( new_n890_, new_n861_ );
nor g0689 ( new_n891_, new_n860_, new_n831_ );
nor g0690 ( new_n892_, new_n890_, new_n891_ );
nand g0691 ( new_n893_, new_n892_, new_n887_ );
nand g0692 ( new_n894_, new_n893_, new_n889_ );
nand g0693 ( new_n895_, new_n894_, keyIn_0_42 );
not g0694 ( new_n896_, keyIn_0_42 );
nor g0695 ( new_n897_, new_n892_, new_n887_ );
nor g0696 ( new_n898_, new_n866_, new_n888_ );
nor g0697 ( new_n899_, new_n897_, new_n898_ );
nand g0698 ( new_n900_, new_n899_, new_n896_ );
nand g0699 ( new_n901_, new_n900_, new_n895_ );
nor g0700 ( new_n902_, new_n679_, new_n842_ );
not g0701 ( new_n903_, new_n902_ );
nand g0702 ( new_n904_, new_n679_, new_n842_ );
nand g0703 ( new_n905_, new_n903_, new_n904_ );
nand g0704 ( new_n906_, N135, N137 );
nand g0705 ( new_n907_, new_n905_, new_n906_ );
not g0706 ( new_n908_, new_n904_ );
nor g0707 ( new_n909_, new_n908_, new_n902_ );
not g0708 ( new_n910_, new_n906_ );
nand g0709 ( new_n911_, new_n909_, new_n910_ );
nand g0710 ( new_n912_, new_n911_, new_n907_ );
not g0711 ( new_n913_, keyIn_0_31 );
nor g0712 ( new_n914_, new_n244_, N89 );
nor g0713 ( new_n915_, new_n218_, N73 );
nor g0714 ( new_n916_, new_n914_, new_n915_ );
nor g0715 ( new_n917_, new_n328_, N121 );
nor g0716 ( new_n918_, new_n348_, N105 );
nor g0717 ( new_n919_, new_n917_, new_n918_ );
not g0718 ( new_n920_, new_n919_ );
nor g0719 ( new_n921_, new_n920_, new_n916_ );
nand g0720 ( new_n922_, new_n920_, new_n916_ );
not g0721 ( new_n923_, new_n922_ );
nor g0722 ( new_n924_, new_n923_, new_n921_ );
not g0723 ( new_n925_, new_n924_ );
nor g0724 ( new_n926_, new_n925_, new_n913_ );
nand g0725 ( new_n927_, new_n925_, new_n913_ );
not g0726 ( new_n928_, new_n927_ );
nor g0727 ( new_n929_, new_n928_, new_n926_ );
nor g0728 ( new_n930_, new_n912_, new_n929_ );
nand g0729 ( new_n931_, new_n912_, new_n929_ );
not g0730 ( new_n932_, new_n931_ );
nor g0731 ( new_n933_, new_n932_, new_n930_ );
nor g0732 ( new_n934_, new_n933_, keyIn_0_44 );
not g0733 ( new_n935_, keyIn_0_44 );
not g0734 ( new_n936_, new_n930_ );
nand g0735 ( new_n937_, new_n936_, new_n931_ );
nor g0736 ( new_n938_, new_n937_, new_n935_ );
nor g0737 ( new_n939_, new_n934_, new_n938_ );
nor g0738 ( new_n940_, new_n901_, new_n939_ );
nand g0739 ( new_n941_, new_n830_, new_n940_ );
nor g0740 ( new_n942_, new_n941_, new_n829_ );
not g0741 ( new_n943_, new_n942_ );
nor g0742 ( new_n944_, new_n752_, new_n943_ );
nand g0743 ( new_n945_, new_n612_, new_n944_ );
nor g0744 ( new_n946_, new_n945_, new_n318_ );
nor g0745 ( new_n947_, new_n946_, new_n203_ );
nand g0746 ( new_n948_, new_n946_, new_n203_ );
not g0747 ( new_n949_, new_n948_ );
nor g0748 ( new_n950_, new_n949_, new_n947_ );
nor g0749 ( new_n951_, new_n950_, new_n202_ );
not g0750 ( new_n952_, new_n950_ );
nor g0751 ( new_n953_, new_n952_, keyIn_0_107 );
nor g0752 ( N724, new_n953_, new_n951_ );
not g0753 ( new_n955_, keyIn_0_86 );
nor g0754 ( new_n956_, new_n945_, new_n417_ );
nor g0755 ( new_n957_, new_n956_, new_n955_ );
nand g0756 ( new_n958_, new_n956_, new_n955_ );
not g0757 ( new_n959_, new_n958_ );
nor g0758 ( new_n960_, new_n959_, new_n957_ );
not g0759 ( new_n961_, new_n960_ );
nand g0760 ( new_n962_, new_n961_, N5 );
not g0761 ( new_n963_, new_n962_ );
nor g0762 ( new_n964_, new_n961_, N5 );
nor g0763 ( new_n965_, new_n963_, new_n964_ );
nor g0764 ( new_n966_, new_n965_, keyIn_0_108 );
not g0765 ( new_n967_, keyIn_0_108 );
not g0766 ( new_n968_, new_n965_ );
nor g0767 ( new_n969_, new_n968_, new_n967_ );
nor g0768 ( N725, new_n969_, new_n966_ );
nor g0769 ( new_n971_, new_n945_, new_n531_ );
nor g0770 ( new_n972_, new_n971_, keyIn_0_87 );
nand g0771 ( new_n973_, new_n971_, keyIn_0_87 );
not g0772 ( new_n974_, new_n973_ );
nor g0773 ( new_n975_, new_n974_, new_n972_ );
not g0774 ( new_n976_, new_n975_ );
nand g0775 ( new_n977_, new_n976_, N9 );
nand g0776 ( new_n978_, new_n975_, new_n510_ );
nand g0777 ( new_n979_, new_n977_, new_n978_ );
nand g0778 ( new_n980_, new_n979_, keyIn_0_109 );
not g0779 ( new_n981_, keyIn_0_109 );
not g0780 ( new_n982_, new_n979_ );
nand g0781 ( new_n983_, new_n982_, new_n981_ );
nand g0782 ( N726, new_n983_, new_n980_ );
not g0783 ( new_n985_, keyIn_0_88 );
nor g0784 ( new_n986_, new_n945_, new_n483_ );
nor g0785 ( new_n987_, new_n986_, new_n985_ );
nand g0786 ( new_n988_, new_n986_, new_n985_ );
not g0787 ( new_n989_, new_n988_ );
nor g0788 ( new_n990_, new_n989_, new_n987_ );
not g0789 ( new_n991_, new_n990_ );
nand g0790 ( new_n992_, new_n991_, new_n446_ );
nand g0791 ( new_n993_, new_n990_, N13 );
nand g0792 ( new_n994_, new_n992_, new_n993_ );
nand g0793 ( new_n995_, new_n994_, keyIn_0_110 );
not g0794 ( new_n996_, keyIn_0_110 );
not g0795 ( new_n997_, new_n994_ );
nand g0796 ( new_n998_, new_n997_, new_n996_ );
nand g0797 ( N727, new_n998_, new_n995_ );
nor g0798 ( new_n1000_, new_n746_, keyIn_0_55 );
nand g0799 ( new_n1001_, new_n746_, keyIn_0_55 );
not g0800 ( new_n1002_, new_n1001_ );
nor g0801 ( new_n1003_, new_n1002_, new_n1000_ );
not g0802 ( new_n1004_, keyIn_0_45 );
not g0803 ( new_n1005_, new_n819_ );
nor g0804 ( new_n1006_, new_n800_, new_n818_ );
nor g0805 ( new_n1007_, new_n1005_, new_n1006_ );
nand g0806 ( new_n1008_, new_n1007_, new_n1004_ );
nand g0807 ( new_n1009_, new_n1008_, new_n825_ );
nand g0808 ( new_n1010_, new_n937_, new_n935_ );
nand g0809 ( new_n1011_, new_n933_, keyIn_0_44 );
nand g0810 ( new_n1012_, new_n1011_, new_n1010_ );
nor g0811 ( new_n1013_, new_n901_, new_n1012_ );
nand g0812 ( new_n1014_, new_n1013_, new_n1009_ );
nor g0813 ( new_n1015_, new_n1003_, new_n1014_ );
nand g0814 ( new_n1016_, new_n612_, new_n1015_ );
nand g0815 ( new_n1017_, new_n1016_, keyIn_0_80 );
not g0816 ( new_n1018_, new_n1017_ );
nor g0817 ( new_n1019_, new_n1016_, keyIn_0_80 );
nor g0818 ( new_n1020_, new_n1018_, new_n1019_ );
nor g0819 ( new_n1021_, new_n1020_, new_n318_ );
not g0820 ( new_n1022_, new_n1021_ );
nand g0821 ( new_n1023_, new_n1022_, N17 );
nand g0822 ( new_n1024_, new_n1021_, new_n298_ );
nand g0823 ( N728, new_n1023_, new_n1024_ );
nor g0824 ( new_n1026_, new_n1020_, new_n417_ );
not g0825 ( new_n1027_, new_n1026_ );
nand g0826 ( new_n1028_, new_n1027_, N21 );
nand g0827 ( new_n1029_, new_n1026_, new_n387_ );
nand g0828 ( N729, new_n1028_, new_n1029_ );
nor g0829 ( new_n1031_, new_n1020_, new_n531_ );
not g0830 ( new_n1032_, new_n1031_ );
nand g0831 ( new_n1033_, new_n1032_, N25 );
nand g0832 ( new_n1034_, new_n1031_, new_n512_ );
nand g0833 ( N730, new_n1033_, new_n1034_ );
nor g0834 ( new_n1036_, new_n1020_, new_n483_ );
nor g0835 ( new_n1037_, new_n1036_, new_n448_ );
nand g0836 ( new_n1038_, new_n1036_, new_n448_ );
not g0837 ( new_n1039_, new_n1038_ );
nor g0838 ( new_n1040_, new_n1039_, new_n1037_ );
nor g0839 ( new_n1041_, new_n1040_, keyIn_0_111 );
not g0840 ( new_n1042_, keyIn_0_111 );
not g0841 ( new_n1043_, new_n1040_ );
nor g0842 ( new_n1044_, new_n1043_, new_n1042_ );
nor g0843 ( N731, new_n1044_, new_n1041_ );
not g0844 ( new_n1046_, keyIn_0_56 );
nor g0845 ( new_n1047_, new_n901_, new_n1046_ );
not g0846 ( new_n1048_, new_n895_ );
nor g0847 ( new_n1049_, new_n894_, keyIn_0_42 );
nor g0848 ( new_n1050_, new_n1048_, new_n1049_ );
nor g0849 ( new_n1051_, new_n1050_, keyIn_0_56 );
nor g0850 ( new_n1052_, new_n1009_, new_n939_ );
not g0851 ( new_n1053_, new_n1052_ );
nor g0852 ( new_n1054_, new_n1053_, new_n1051_ );
not g0853 ( new_n1055_, new_n1054_ );
nor g0854 ( new_n1056_, new_n1055_, new_n1047_ );
nand g0855 ( new_n1057_, new_n1056_, new_n750_ );
not g0856 ( new_n1058_, new_n1057_ );
nand g0857 ( new_n1059_, new_n612_, new_n1058_ );
nor g0858 ( new_n1060_, new_n1059_, new_n318_ );
nor g0859 ( new_n1061_, new_n1060_, keyIn_0_89 );
nand g0860 ( new_n1062_, new_n1060_, keyIn_0_89 );
not g0861 ( new_n1063_, new_n1062_ );
nor g0862 ( new_n1064_, new_n1063_, new_n1061_ );
not g0863 ( new_n1065_, new_n1064_ );
nand g0864 ( new_n1066_, new_n1065_, new_n287_ );
nand g0865 ( new_n1067_, new_n1064_, N33 );
nand g0866 ( new_n1068_, new_n1066_, new_n1067_ );
nand g0867 ( new_n1069_, new_n1068_, keyIn_0_112 );
not g0868 ( new_n1070_, keyIn_0_112 );
not g0869 ( new_n1071_, new_n1068_ );
nand g0870 ( new_n1072_, new_n1071_, new_n1070_ );
nand g0871 ( N732, new_n1072_, new_n1069_ );
not g0872 ( new_n1074_, keyIn_0_113 );
nor g0873 ( new_n1075_, new_n1059_, new_n417_ );
nor g0874 ( new_n1076_, new_n1075_, keyIn_0_90 );
nand g0875 ( new_n1077_, new_n1075_, keyIn_0_90 );
not g0876 ( new_n1078_, new_n1077_ );
nor g0877 ( new_n1079_, new_n1078_, new_n1076_ );
not g0878 ( new_n1080_, new_n1079_ );
nand g0879 ( new_n1081_, new_n1080_, new_n395_ );
nand g0880 ( new_n1082_, new_n1079_, N37 );
nand g0881 ( new_n1083_, new_n1081_, new_n1082_ );
nand g0882 ( new_n1084_, new_n1083_, new_n1074_ );
not g0883 ( new_n1085_, new_n1083_ );
nand g0884 ( new_n1086_, new_n1085_, keyIn_0_113 );
nand g0885 ( N733, new_n1086_, new_n1084_ );
nor g0886 ( new_n1088_, new_n1059_, new_n531_ );
nor g0887 ( new_n1089_, new_n1088_, keyIn_0_91 );
nand g0888 ( new_n1090_, new_n1088_, keyIn_0_91 );
not g0889 ( new_n1091_, new_n1090_ );
nor g0890 ( new_n1092_, new_n1091_, new_n1089_ );
not g0891 ( new_n1093_, new_n1092_ );
nand g0892 ( new_n1094_, new_n1093_, new_n500_ );
nand g0893 ( new_n1095_, new_n1092_, N41 );
nand g0894 ( N734, new_n1094_, new_n1095_ );
not g0895 ( new_n1097_, keyIn_0_114 );
nor g0896 ( new_n1098_, new_n1059_, new_n483_ );
nor g0897 ( new_n1099_, new_n1098_, new_n456_ );
nand g0898 ( new_n1100_, new_n1098_, new_n456_ );
not g0899 ( new_n1101_, new_n1100_ );
nor g0900 ( new_n1102_, new_n1101_, new_n1099_ );
not g0901 ( new_n1103_, new_n1102_ );
nand g0902 ( new_n1104_, new_n1103_, new_n1097_ );
nand g0903 ( new_n1105_, new_n1102_, keyIn_0_114 );
nand g0904 ( N735, new_n1104_, new_n1105_ );
not g0905 ( new_n1107_, keyIn_0_92 );
nor g0906 ( new_n1108_, new_n901_, keyIn_0_57 );
nand g0907 ( new_n1109_, new_n901_, keyIn_0_57 );
not g0908 ( new_n1110_, new_n1109_ );
nor g0909 ( new_n1111_, new_n1110_, new_n1108_ );
not g0910 ( new_n1112_, keyIn_0_58 );
nand g0911 ( new_n1113_, new_n939_, new_n1112_ );
nand g0912 ( new_n1114_, new_n1012_, keyIn_0_58 );
nand g0913 ( new_n1115_, new_n1113_, new_n1114_ );
nand g0914 ( new_n1116_, new_n1115_, new_n1009_ );
nor g0915 ( new_n1117_, new_n746_, new_n1116_ );
not g0916 ( new_n1118_, new_n1117_ );
nor g0917 ( new_n1119_, new_n1118_, new_n1111_ );
nand g0918 ( new_n1120_, new_n612_, new_n1119_ );
nand g0919 ( new_n1121_, new_n1120_, keyIn_0_81 );
not g0920 ( new_n1122_, keyIn_0_81 );
nor g0921 ( new_n1123_, new_n610_, new_n597_ );
nor g0922 ( new_n1124_, new_n595_, keyIn_0_78 );
nor g0923 ( new_n1125_, new_n1124_, new_n1123_ );
not g0924 ( new_n1126_, new_n1119_ );
nor g0925 ( new_n1127_, new_n1125_, new_n1126_ );
nand g0926 ( new_n1128_, new_n1127_, new_n1122_ );
nand g0927 ( new_n1129_, new_n1128_, new_n1121_ );
nor g0928 ( new_n1130_, new_n1129_, new_n318_ );
nor g0929 ( new_n1131_, new_n1130_, new_n1107_ );
nand g0930 ( new_n1132_, new_n1130_, new_n1107_ );
not g0931 ( new_n1133_, new_n1132_ );
nor g0932 ( new_n1134_, new_n1133_, new_n1131_ );
not g0933 ( new_n1135_, new_n1134_ );
nand g0934 ( new_n1136_, new_n1135_, N49 );
nand g0935 ( new_n1137_, new_n1134_, new_n289_ );
nand g0936 ( N736, new_n1136_, new_n1137_ );
not g0937 ( new_n1139_, keyIn_0_93 );
nor g0938 ( new_n1140_, new_n1129_, new_n417_ );
nor g0939 ( new_n1141_, new_n1140_, new_n1139_ );
nand g0940 ( new_n1142_, new_n1140_, new_n1139_ );
not g0941 ( new_n1143_, new_n1142_ );
nor g0942 ( new_n1144_, new_n1143_, new_n1141_ );
not g0943 ( new_n1145_, new_n1144_ );
nand g0944 ( new_n1146_, new_n1145_, N53 );
nand g0945 ( new_n1147_, new_n1144_, new_n397_ );
nand g0946 ( N737, new_n1146_, new_n1147_ );
not g0947 ( new_n1149_, new_n1121_ );
nor g0948 ( new_n1150_, new_n1120_, keyIn_0_81 );
nor g0949 ( new_n1151_, new_n1149_, new_n1150_ );
nand g0950 ( new_n1152_, new_n1151_, new_n528_ );
nand g0951 ( new_n1153_, new_n1152_, keyIn_0_94 );
not g0952 ( new_n1154_, keyIn_0_94 );
nor g0953 ( new_n1155_, new_n1129_, new_n531_ );
nand g0954 ( new_n1156_, new_n1155_, new_n1154_ );
nand g0955 ( new_n1157_, new_n1153_, new_n1156_ );
nand g0956 ( new_n1158_, new_n1157_, N57 );
not g0957 ( new_n1159_, new_n1158_ );
nor g0958 ( new_n1160_, new_n1157_, N57 );
nor g0959 ( new_n1161_, new_n1159_, new_n1160_ );
nor g0960 ( new_n1162_, new_n1161_, keyIn_0_115 );
not g0961 ( new_n1163_, keyIn_0_115 );
not g0962 ( new_n1164_, new_n1157_ );
nand g0963 ( new_n1165_, new_n1164_, new_n502_ );
nand g0964 ( new_n1166_, new_n1165_, new_n1158_ );
nor g0965 ( new_n1167_, new_n1166_, new_n1163_ );
nor g0966 ( N738, new_n1162_, new_n1167_ );
nand g0967 ( new_n1169_, new_n1151_, new_n484_ );
nand g0968 ( new_n1170_, new_n1169_, keyIn_0_95 );
not g0969 ( new_n1171_, keyIn_0_95 );
nor g0970 ( new_n1172_, new_n1129_, new_n483_ );
nand g0971 ( new_n1173_, new_n1172_, new_n1171_ );
nand g0972 ( new_n1174_, new_n1170_, new_n1173_ );
nand g0973 ( new_n1175_, new_n1174_, new_n458_ );
nor g0974 ( new_n1176_, new_n1174_, new_n458_ );
not g0975 ( new_n1177_, new_n1176_ );
nand g0976 ( new_n1178_, new_n1177_, new_n1175_ );
nand g0977 ( new_n1179_, new_n1178_, keyIn_0_116 );
not g0978 ( new_n1180_, keyIn_0_116 );
not g0979 ( new_n1181_, new_n1175_ );
nor g0980 ( new_n1182_, new_n1181_, new_n1176_ );
nand g0981 ( new_n1183_, new_n1182_, new_n1180_ );
nand g0982 ( N739, new_n1183_, new_n1179_ );
not g0983 ( new_n1185_, keyIn_0_96 );
nor g0984 ( new_n1186_, new_n746_, keyIn_0_59 );
not g0985 ( new_n1187_, new_n1186_ );
nand g0986 ( new_n1188_, new_n746_, keyIn_0_59 );
nor g0987 ( new_n1189_, new_n1012_, keyIn_0_60 );
not g0988 ( new_n1190_, keyIn_0_60 );
nor g0989 ( new_n1191_, new_n939_, new_n1190_ );
nor g0990 ( new_n1192_, new_n1191_, new_n1189_ );
nand g0991 ( new_n1193_, new_n1009_, new_n901_ );
nor g0992 ( new_n1194_, new_n1193_, new_n1192_ );
nand g0993 ( new_n1195_, new_n1188_, new_n1194_ );
not g0994 ( new_n1196_, new_n1195_ );
nand g0995 ( new_n1197_, new_n1196_, new_n1187_ );
nand g0996 ( new_n1198_, new_n1197_, keyIn_0_76 );
not g0997 ( new_n1199_, keyIn_0_76 );
nor g0998 ( new_n1200_, new_n1195_, new_n1186_ );
nand g0999 ( new_n1201_, new_n1200_, new_n1199_ );
nand g1000 ( new_n1202_, new_n1198_, new_n1201_ );
not g1001 ( new_n1203_, keyIn_0_77 );
nor g1002 ( new_n1204_, new_n1009_, keyIn_0_66 );
nand g1003 ( new_n1205_, new_n1009_, keyIn_0_66 );
not g1004 ( new_n1206_, new_n1205_ );
nor g1005 ( new_n1207_, new_n1206_, new_n1204_ );
not g1006 ( new_n1208_, new_n1207_ );
not g1007 ( new_n1209_, keyIn_0_65 );
nand g1008 ( new_n1210_, new_n1012_, new_n1209_ );
nand g1009 ( new_n1211_, new_n939_, keyIn_0_65 );
nand g1010 ( new_n1212_, new_n1211_, new_n1210_ );
nor g1011 ( new_n1213_, new_n1212_, new_n901_ );
nand g1012 ( new_n1214_, new_n746_, new_n1213_ );
not g1013 ( new_n1215_, new_n1214_ );
nand g1014 ( new_n1216_, new_n1215_, new_n1208_ );
nor g1015 ( new_n1217_, new_n1216_, new_n1203_ );
nand g1016 ( new_n1218_, new_n1216_, new_n1203_ );
nor g1017 ( new_n1219_, new_n1009_, keyIn_0_61 );
not g1018 ( new_n1220_, new_n1219_ );
not g1019 ( new_n1221_, keyIn_0_61 );
nor g1020 ( new_n1222_, new_n828_, new_n1221_ );
nand g1021 ( new_n1223_, new_n901_, new_n1012_ );
nor g1022 ( new_n1224_, new_n1222_, new_n1223_ );
nand g1023 ( new_n1225_, new_n1224_, new_n1220_ );
nor g1024 ( new_n1226_, new_n1225_, new_n750_ );
nor g1025 ( new_n1227_, new_n1009_, keyIn_0_64 );
not g1026 ( new_n1228_, new_n1227_ );
not g1027 ( new_n1229_, keyIn_0_62 );
nand g1028 ( new_n1230_, new_n901_, new_n1229_ );
not g1029 ( new_n1231_, new_n1230_ );
nor g1030 ( new_n1232_, new_n901_, new_n1229_ );
nor g1031 ( new_n1233_, new_n1231_, new_n1232_ );
nand g1032 ( new_n1234_, new_n1233_, new_n1228_ );
nand g1033 ( new_n1235_, new_n1009_, keyIn_0_64 );
not g1034 ( new_n1236_, keyIn_0_63 );
nor g1035 ( new_n1237_, new_n939_, new_n1236_ );
nor g1036 ( new_n1238_, new_n1012_, keyIn_0_63 );
nor g1037 ( new_n1239_, new_n1237_, new_n1238_ );
nand g1038 ( new_n1240_, new_n1239_, new_n1235_ );
not g1039 ( new_n1241_, new_n1240_ );
nand g1040 ( new_n1242_, new_n750_, new_n1241_ );
nor g1041 ( new_n1243_, new_n1242_, new_n1234_ );
nor g1042 ( new_n1244_, new_n1243_, new_n1226_ );
nand g1043 ( new_n1245_, new_n1244_, new_n1218_ );
nor g1044 ( new_n1246_, new_n1245_, new_n1217_ );
nand g1045 ( new_n1247_, new_n1246_, new_n1202_ );
nand g1046 ( new_n1248_, new_n1247_, keyIn_0_79 );
not g1047 ( new_n1249_, keyIn_0_79 );
nor g1048 ( new_n1250_, new_n1200_, new_n1199_ );
not g1049 ( new_n1251_, new_n1201_ );
nor g1050 ( new_n1252_, new_n1251_, new_n1250_ );
not g1051 ( new_n1253_, new_n1217_ );
nor g1052 ( new_n1254_, new_n1214_, new_n1207_ );
nor g1053 ( new_n1255_, new_n1254_, keyIn_0_77 );
nand g1054 ( new_n1256_, new_n1009_, keyIn_0_61 );
not g1055 ( new_n1257_, new_n1223_ );
nand g1056 ( new_n1258_, new_n1257_, new_n1256_ );
nor g1057 ( new_n1259_, new_n1258_, new_n1219_ );
nand g1058 ( new_n1260_, new_n1259_, new_n746_ );
nand g1059 ( new_n1261_, new_n1050_, keyIn_0_62 );
nand g1060 ( new_n1262_, new_n1261_, new_n1230_ );
nor g1061 ( new_n1263_, new_n1262_, new_n1227_ );
nor g1062 ( new_n1264_, new_n746_, new_n1240_ );
nand g1063 ( new_n1265_, new_n1264_, new_n1263_ );
nand g1064 ( new_n1266_, new_n1260_, new_n1265_ );
nor g1065 ( new_n1267_, new_n1255_, new_n1266_ );
nand g1066 ( new_n1268_, new_n1267_, new_n1253_ );
nor g1067 ( new_n1269_, new_n1252_, new_n1268_ );
nand g1068 ( new_n1270_, new_n1269_, new_n1249_ );
nand g1069 ( new_n1271_, new_n1270_, new_n1248_ );
not g1070 ( new_n1272_, keyIn_0_68 );
nor g1071 ( new_n1273_, new_n483_, new_n1272_ );
nor g1072 ( new_n1274_, new_n484_, keyIn_0_68 );
nor g1073 ( new_n1275_, new_n417_, keyIn_0_67 );
nand g1074 ( new_n1276_, new_n417_, keyIn_0_67 );
nand g1075 ( new_n1277_, new_n1276_, new_n528_ );
nor g1076 ( new_n1278_, new_n1277_, new_n1275_ );
not g1077 ( new_n1279_, new_n1278_ );
nor g1078 ( new_n1280_, new_n1279_, new_n1274_ );
not g1079 ( new_n1281_, new_n1280_ );
nor g1080 ( new_n1282_, new_n1281_, new_n1273_ );
nand g1081 ( new_n1283_, new_n1282_, new_n547_ );
not g1082 ( new_n1284_, new_n1283_ );
nand g1083 ( new_n1285_, new_n1271_, new_n1284_ );
nand g1084 ( new_n1286_, new_n1285_, keyIn_0_82 );
not g1085 ( new_n1287_, new_n1286_ );
nor g1086 ( new_n1288_, new_n1285_, keyIn_0_82 );
nor g1087 ( new_n1289_, new_n1287_, new_n1288_ );
nand g1088 ( new_n1290_, new_n1289_, new_n1050_ );
nand g1089 ( new_n1291_, new_n1290_, new_n1185_ );
not g1090 ( new_n1292_, keyIn_0_82 );
nor g1091 ( new_n1293_, new_n1269_, new_n1249_ );
nor g1092 ( new_n1294_, new_n1247_, keyIn_0_79 );
nor g1093 ( new_n1295_, new_n1293_, new_n1294_ );
nor g1094 ( new_n1296_, new_n1295_, new_n1283_ );
nand g1095 ( new_n1297_, new_n1296_, new_n1292_ );
nand g1096 ( new_n1298_, new_n1297_, new_n1286_ );
nor g1097 ( new_n1299_, new_n1298_, new_n901_ );
nand g1098 ( new_n1300_, new_n1299_, keyIn_0_96 );
nand g1099 ( new_n1301_, new_n1291_, new_n1300_ );
nand g1100 ( new_n1302_, new_n1301_, N65 );
not g1101 ( new_n1303_, new_n1302_ );
nor g1102 ( new_n1304_, new_n1301_, N65 );
nor g1103 ( new_n1305_, new_n1303_, new_n1304_ );
nor g1104 ( new_n1306_, new_n1305_, keyIn_0_117 );
not g1105 ( new_n1307_, keyIn_0_117 );
not g1106 ( new_n1308_, new_n1301_ );
nand g1107 ( new_n1309_, new_n1308_, new_n239_ );
nand g1108 ( new_n1310_, new_n1309_, new_n1302_ );
nor g1109 ( new_n1311_, new_n1310_, new_n1307_ );
nor g1110 ( N740, new_n1306_, new_n1311_ );
not g1111 ( new_n1313_, keyIn_0_97 );
nand g1112 ( new_n1314_, new_n1289_, new_n750_ );
nand g1113 ( new_n1315_, new_n1314_, new_n1313_ );
nor g1114 ( new_n1316_, new_n1298_, new_n746_ );
nand g1115 ( new_n1317_, new_n1316_, keyIn_0_97 );
nand g1116 ( new_n1318_, new_n1315_, new_n1317_ );
nand g1117 ( new_n1319_, new_n1318_, new_n241_ );
not g1118 ( new_n1320_, new_n1319_ );
nor g1119 ( new_n1321_, new_n1318_, new_n241_ );
nor g1120 ( new_n1322_, new_n1320_, new_n1321_ );
nor g1121 ( new_n1323_, new_n1322_, keyIn_0_118 );
not g1122 ( new_n1324_, keyIn_0_118 );
not g1123 ( new_n1325_, new_n1318_ );
nand g1124 ( new_n1326_, new_n1325_, N69 );
nand g1125 ( new_n1327_, new_n1326_, new_n1319_ );
nor g1126 ( new_n1328_, new_n1327_, new_n1324_ );
nor g1127 ( N741, new_n1323_, new_n1328_ );
not g1128 ( new_n1330_, keyIn_0_98 );
nor g1129 ( new_n1331_, new_n1298_, new_n939_ );
nor g1130 ( new_n1332_, new_n1331_, new_n1330_ );
nand g1131 ( new_n1333_, new_n1331_, new_n1330_ );
not g1132 ( new_n1334_, new_n1333_ );
nor g1133 ( new_n1335_, new_n1334_, new_n1332_ );
not g1134 ( new_n1336_, new_n1335_ );
nand g1135 ( new_n1337_, new_n1336_, new_n244_ );
nand g1136 ( new_n1338_, new_n1335_, N73 );
nand g1137 ( N742, new_n1337_, new_n1338_ );
not g1138 ( new_n1340_, keyIn_0_119 );
nor g1139 ( new_n1341_, new_n1298_, new_n828_ );
nor g1140 ( new_n1342_, new_n1341_, new_n246_ );
nand g1141 ( new_n1343_, new_n1341_, new_n246_ );
not g1142 ( new_n1344_, new_n1343_ );
nor g1143 ( new_n1345_, new_n1344_, new_n1342_ );
not g1144 ( new_n1346_, new_n1345_ );
nand g1145 ( new_n1347_, new_n1346_, new_n1340_ );
nand g1146 ( new_n1348_, new_n1345_, keyIn_0_119 );
nand g1147 ( N743, new_n1347_, new_n1348_ );
not g1148 ( new_n1350_, keyIn_0_120 );
nor g1149 ( new_n1351_, new_n416_, keyIn_0_69 );
nand g1150 ( new_n1352_, new_n416_, keyIn_0_69 );
not g1151 ( new_n1353_, new_n1352_ );
nor g1152 ( new_n1354_, new_n1353_, new_n1351_ );
nor g1153 ( new_n1355_, new_n528_, keyIn_0_70 );
nand g1154 ( new_n1356_, new_n528_, keyIn_0_70 );
not g1155 ( new_n1357_, new_n1356_ );
nor g1156 ( new_n1358_, new_n1357_, new_n1355_ );
nor g1157 ( new_n1359_, new_n1358_, new_n483_ );
not g1158 ( new_n1360_, new_n1359_ );
nor g1159 ( new_n1361_, new_n1360_, new_n1354_ );
nand g1160 ( new_n1362_, new_n1361_, new_n547_ );
not g1161 ( new_n1363_, new_n1362_ );
nand g1162 ( new_n1364_, new_n1271_, new_n1363_ );
nand g1163 ( new_n1365_, new_n1364_, keyIn_0_83 );
nor g1164 ( new_n1366_, new_n1364_, keyIn_0_83 );
not g1165 ( new_n1367_, new_n1366_ );
nand g1166 ( new_n1368_, new_n1367_, new_n1365_ );
nand g1167 ( new_n1369_, new_n1368_, new_n1050_ );
nand g1168 ( new_n1370_, new_n1369_, keyIn_0_99 );
not g1169 ( new_n1371_, keyIn_0_99 );
not g1170 ( new_n1372_, new_n1365_ );
nor g1171 ( new_n1373_, new_n1372_, new_n1366_ );
nor g1172 ( new_n1374_, new_n1373_, new_n901_ );
nand g1173 ( new_n1375_, new_n1374_, new_n1371_ );
nand g1174 ( new_n1376_, new_n1375_, new_n1370_ );
nand g1175 ( new_n1377_, new_n1376_, N81 );
nor g1176 ( new_n1378_, new_n1376_, N81 );
not g1177 ( new_n1379_, new_n1378_ );
nand g1178 ( new_n1380_, new_n1379_, new_n1377_ );
nand g1179 ( new_n1381_, new_n1380_, new_n1350_ );
not g1180 ( new_n1382_, new_n1377_ );
nor g1181 ( new_n1383_, new_n1382_, new_n1378_ );
nand g1182 ( new_n1384_, new_n1383_, keyIn_0_120 );
nand g1183 ( N744, new_n1384_, new_n1381_ );
nor g1184 ( new_n1386_, new_n1373_, new_n746_ );
nor g1185 ( new_n1387_, new_n1386_, new_n205_ );
nand g1186 ( new_n1388_, new_n1386_, new_n205_ );
not g1187 ( new_n1389_, new_n1388_ );
nor g1188 ( new_n1390_, new_n1389_, new_n1387_ );
nor g1189 ( new_n1391_, new_n1390_, keyIn_0_121 );
not g1190 ( new_n1392_, keyIn_0_121 );
not g1191 ( new_n1393_, new_n1390_ );
nor g1192 ( new_n1394_, new_n1393_, new_n1392_ );
nor g1193 ( N745, new_n1394_, new_n1391_ );
not g1194 ( new_n1396_, keyIn_0_122 );
nand g1195 ( new_n1397_, new_n1368_, new_n1012_ );
nand g1196 ( new_n1398_, new_n1397_, keyIn_0_100 );
not g1197 ( new_n1399_, keyIn_0_100 );
nor g1198 ( new_n1400_, new_n1373_, new_n939_ );
nand g1199 ( new_n1401_, new_n1400_, new_n1399_ );
nand g1200 ( new_n1402_, new_n1401_, new_n1398_ );
nand g1201 ( new_n1403_, new_n1402_, N89 );
nor g1202 ( new_n1404_, new_n1402_, N89 );
not g1203 ( new_n1405_, new_n1404_ );
nand g1204 ( new_n1406_, new_n1405_, new_n1403_ );
nand g1205 ( new_n1407_, new_n1406_, new_n1396_ );
not g1206 ( new_n1408_, new_n1403_ );
nor g1207 ( new_n1409_, new_n1408_, new_n1404_ );
nand g1208 ( new_n1410_, new_n1409_, keyIn_0_122 );
nand g1209 ( N746, new_n1410_, new_n1407_ );
not g1210 ( new_n1412_, keyIn_0_101 );
nor g1211 ( new_n1413_, new_n1373_, new_n828_ );
nor g1212 ( new_n1414_, new_n1413_, new_n1412_ );
nand g1213 ( new_n1415_, new_n1413_, new_n1412_ );
not g1214 ( new_n1416_, new_n1415_ );
nor g1215 ( new_n1417_, new_n1416_, new_n1414_ );
not g1216 ( new_n1418_, new_n1417_ );
nand g1217 ( new_n1419_, new_n1418_, new_n216_ );
nand g1218 ( new_n1420_, new_n1417_, N93 );
nand g1219 ( N747, new_n1419_, new_n1420_ );
not g1220 ( new_n1422_, keyIn_0_102 );
not g1221 ( new_n1423_, keyIn_0_84 );
nor g1222 ( new_n1424_, new_n561_, new_n550_ );
nand g1223 ( new_n1425_, new_n1271_, new_n1424_ );
nand g1224 ( new_n1426_, new_n1425_, new_n1423_ );
not g1225 ( new_n1427_, new_n1426_ );
nor g1226 ( new_n1428_, new_n1425_, new_n1423_ );
nor g1227 ( new_n1429_, new_n1427_, new_n1428_ );
nor g1228 ( new_n1430_, new_n1429_, new_n901_ );
nor g1229 ( new_n1431_, new_n1430_, new_n1422_ );
nand g1230 ( new_n1432_, new_n1430_, new_n1422_ );
not g1231 ( new_n1433_, new_n1432_ );
nor g1232 ( new_n1434_, new_n1433_, new_n1431_ );
not g1233 ( new_n1435_, new_n1434_ );
nand g1234 ( new_n1436_, new_n1435_, new_n335_ );
nand g1235 ( new_n1437_, new_n1434_, N97 );
nand g1236 ( N748, new_n1436_, new_n1437_ );
nor g1237 ( new_n1439_, new_n1429_, new_n746_ );
nor g1238 ( new_n1440_, new_n1439_, keyIn_0_103 );
nand g1239 ( new_n1441_, new_n1439_, keyIn_0_103 );
not g1240 ( new_n1442_, new_n1441_ );
nor g1241 ( new_n1443_, new_n1442_, new_n1440_ );
not g1242 ( new_n1444_, new_n1443_ );
nand g1243 ( new_n1445_, new_n1444_, N101 );
nand g1244 ( new_n1446_, new_n1443_, new_n337_ );
nand g1245 ( N749, new_n1445_, new_n1446_ );
not g1246 ( new_n1448_, keyIn_0_123 );
not g1247 ( new_n1449_, keyIn_0_104 );
not g1248 ( new_n1450_, new_n1428_ );
nand g1249 ( new_n1451_, new_n1450_, new_n1426_ );
nand g1250 ( new_n1452_, new_n1451_, new_n1012_ );
nand g1251 ( new_n1453_, new_n1452_, new_n1449_ );
nor g1252 ( new_n1454_, new_n1429_, new_n939_ );
nand g1253 ( new_n1455_, new_n1454_, keyIn_0_104 );
nand g1254 ( new_n1456_, new_n1455_, new_n1453_ );
nand g1255 ( new_n1457_, new_n1456_, new_n328_ );
nor g1256 ( new_n1458_, new_n1456_, new_n328_ );
not g1257 ( new_n1459_, new_n1458_ );
nand g1258 ( new_n1460_, new_n1459_, new_n1457_ );
nand g1259 ( new_n1461_, new_n1460_, new_n1448_ );
not g1260 ( new_n1462_, new_n1457_ );
nor g1261 ( new_n1463_, new_n1462_, new_n1458_ );
nand g1262 ( new_n1464_, new_n1463_, keyIn_0_123 );
nand g1263 ( N750, new_n1464_, new_n1461_ );
nor g1264 ( new_n1466_, new_n1429_, new_n828_ );
not g1265 ( new_n1467_, new_n1466_ );
nand g1266 ( new_n1468_, new_n1467_, N109 );
nand g1267 ( new_n1469_, new_n1466_, new_n326_ );
nand g1268 ( N751, new_n1468_, new_n1469_ );
not g1269 ( new_n1471_, keyIn_0_105 );
not g1270 ( new_n1472_, keyIn_0_85 );
not g1271 ( new_n1473_, keyIn_0_71 );
nor g1272 ( new_n1474_, new_n528_, new_n1473_ );
nor g1273 ( new_n1475_, new_n531_, keyIn_0_71 );
nor g1274 ( new_n1476_, new_n1475_, new_n1474_ );
nor g1275 ( new_n1477_, new_n1476_, new_n483_ );
nand g1276 ( new_n1478_, new_n562_, new_n1477_ );
not g1277 ( new_n1479_, new_n1478_ );
nand g1278 ( new_n1480_, new_n1271_, new_n1479_ );
nand g1279 ( new_n1481_, new_n1480_, new_n1472_ );
not g1280 ( new_n1482_, new_n1481_ );
nor g1281 ( new_n1483_, new_n1480_, new_n1472_ );
nor g1282 ( new_n1484_, new_n1482_, new_n1483_ );
nand g1283 ( new_n1485_, new_n1484_, new_n1050_ );
nand g1284 ( new_n1486_, new_n1485_, new_n1471_ );
nor g1285 ( new_n1487_, new_n1295_, new_n1478_ );
nand g1286 ( new_n1488_, new_n1487_, keyIn_0_85 );
nand g1287 ( new_n1489_, new_n1488_, new_n1481_ );
nor g1288 ( new_n1490_, new_n1489_, new_n901_ );
nand g1289 ( new_n1491_, new_n1490_, keyIn_0_105 );
nand g1290 ( new_n1492_, new_n1486_, new_n1491_ );
nand g1291 ( new_n1493_, new_n1492_, new_n356_ );
not g1292 ( new_n1494_, new_n1493_ );
nor g1293 ( new_n1495_, new_n1492_, new_n356_ );
nor g1294 ( new_n1496_, new_n1494_, new_n1495_ );
nor g1295 ( new_n1497_, new_n1496_, keyIn_0_124 );
not g1296 ( new_n1498_, keyIn_0_124 );
not g1297 ( new_n1499_, new_n1492_ );
nand g1298 ( new_n1500_, new_n1499_, N113 );
nand g1299 ( new_n1501_, new_n1500_, new_n1493_ );
nor g1300 ( new_n1502_, new_n1501_, new_n1498_ );
nor g1301 ( N752, new_n1497_, new_n1502_ );
not g1302 ( new_n1504_, keyIn_0_106 );
nand g1303 ( new_n1505_, new_n1484_, new_n750_ );
nand g1304 ( new_n1506_, new_n1505_, new_n1504_ );
nor g1305 ( new_n1507_, new_n1489_, new_n746_ );
nand g1306 ( new_n1508_, new_n1507_, keyIn_0_106 );
nand g1307 ( new_n1509_, new_n1506_, new_n1508_ );
nand g1308 ( new_n1510_, new_n1509_, new_n358_ );
not g1309 ( new_n1511_, new_n1510_ );
nor g1310 ( new_n1512_, new_n1509_, new_n358_ );
nor g1311 ( new_n1513_, new_n1511_, new_n1512_ );
nor g1312 ( new_n1514_, new_n1513_, keyIn_0_125 );
not g1313 ( new_n1515_, keyIn_0_125 );
not g1314 ( new_n1516_, new_n1509_ );
nand g1315 ( new_n1517_, new_n1516_, N117 );
nand g1316 ( new_n1518_, new_n1517_, new_n1510_ );
nor g1317 ( new_n1519_, new_n1518_, new_n1515_ );
nor g1318 ( N753, new_n1514_, new_n1519_ );
nor g1319 ( new_n1521_, new_n1489_, new_n939_ );
not g1320 ( new_n1522_, new_n1521_ );
nand g1321 ( new_n1523_, new_n1522_, N121 );
nand g1322 ( new_n1524_, new_n1521_, new_n348_ );
nand g1323 ( new_n1525_, new_n1523_, new_n1524_ );
nand g1324 ( new_n1526_, new_n1525_, keyIn_0_126 );
not g1325 ( new_n1527_, new_n1526_ );
nor g1326 ( new_n1528_, new_n1525_, keyIn_0_126 );
nor g1327 ( N754, new_n1527_, new_n1528_ );
not g1328 ( new_n1530_, keyIn_0_127 );
nor g1329 ( new_n1531_, new_n1489_, new_n828_ );
nor g1330 ( new_n1532_, new_n1531_, new_n346_ );
nand g1331 ( new_n1533_, new_n1531_, new_n346_ );
not g1332 ( new_n1534_, new_n1533_ );
nor g1333 ( new_n1535_, new_n1534_, new_n1532_ );
not g1334 ( new_n1536_, new_n1535_ );
nand g1335 ( new_n1537_, new_n1536_, new_n1530_ );
nand g1336 ( new_n1538_, new_n1535_, keyIn_0_127 );
nand g1337 ( N755, new_n1537_, new_n1538_ );
endmodule