module add_mul_sub_8_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, operation_0_, 
        operation_1_, Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, 
        Result_5_, Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, 
        Result_11_, Result_12_, Result_13_, Result_14_, Result_15_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_,
         b_4_, b_5_, b_6_, b_7_, operation_0_, operation_1_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_;
  wire   n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255;

  NOR2_X2 U606 ( .A1(operation_0_), .A2(operation_1_), .ZN(n606) );
  NOR2_X2 U607 ( .A1(n1216), .A2(operation_0_), .ZN(n608) );
  NAND2_X1 U608 ( .A1(n590), .A2(n591), .ZN(Result_9_) );
  NAND2_X1 U609 ( .A1(n592), .A2(n593), .ZN(n591) );
  XNOR2_X1 U610 ( .A(n594), .B(n595), .ZN(n593) );
  XNOR2_X1 U611 ( .A(n596), .B(n597), .ZN(n595) );
  NOR2_X1 U612 ( .A1(n598), .A2(n599), .ZN(n590) );
  NOR2_X1 U613 ( .A1(n600), .A2(n601), .ZN(n599) );
  NOR2_X1 U614 ( .A1(n602), .A2(n603), .ZN(n600) );
  NAND2_X1 U615 ( .A1(n604), .A2(n605), .ZN(n603) );
  NAND2_X1 U616 ( .A1(n606), .A2(n607), .ZN(n605) );
  NAND2_X1 U617 ( .A1(n608), .A2(n609), .ZN(n604) );
  NOR2_X1 U618 ( .A1(n610), .A2(n611), .ZN(n602) );
  NOR2_X1 U619 ( .A1(n612), .A2(n613), .ZN(n598) );
  INV_X1 U620 ( .A(n601), .ZN(n613) );
  XNOR2_X1 U621 ( .A(n614), .B(a_1_), .ZN(n601) );
  NOR2_X1 U622 ( .A1(n615), .A2(n616), .ZN(n612) );
  NAND2_X1 U623 ( .A1(n617), .A2(n618), .ZN(n616) );
  NAND2_X1 U624 ( .A1(n619), .A2(n606), .ZN(n618) );
  NAND2_X1 U625 ( .A1(n608), .A2(n620), .ZN(n617) );
  NOR2_X1 U626 ( .A1(n621), .A2(n610), .ZN(n615) );
  NAND2_X1 U627 ( .A1(n622), .A2(n623), .ZN(Result_8_) );
  NAND2_X1 U628 ( .A1(n624), .A2(n592), .ZN(n623) );
  XOR2_X1 U629 ( .A(n625), .B(n626), .Z(n624) );
  XOR2_X1 U630 ( .A(n627), .B(n628), .Z(n625) );
  NOR2_X1 U631 ( .A1(n629), .A2(n630), .ZN(n622) );
  NOR2_X1 U632 ( .A1(n631), .A2(n632), .ZN(n630) );
  NOR2_X1 U633 ( .A1(n633), .A2(n634), .ZN(n631) );
  NAND2_X1 U634 ( .A1(n635), .A2(n636), .ZN(n634) );
  NAND2_X1 U635 ( .A1(n637), .A2(n606), .ZN(n636) );
  INV_X1 U636 ( .A(n638), .ZN(n637) );
  NAND2_X1 U637 ( .A1(n639), .A2(n608), .ZN(n635) );
  NOR2_X1 U638 ( .A1(n610), .A2(n640), .ZN(n633) );
  NOR2_X1 U639 ( .A1(n641), .A2(n642), .ZN(n629) );
  INV_X1 U640 ( .A(n632), .ZN(n642) );
  XNOR2_X1 U641 ( .A(n643), .B(a_0_), .ZN(n632) );
  NOR2_X1 U642 ( .A1(n644), .A2(n645), .ZN(n641) );
  NAND2_X1 U643 ( .A1(n646), .A2(n647), .ZN(n645) );
  NAND2_X1 U644 ( .A1(n606), .A2(n638), .ZN(n647) );
  NAND2_X1 U645 ( .A1(n648), .A2(n649), .ZN(n638) );
  OR2_X1 U646 ( .A1(n607), .A2(n650), .ZN(n649) );
  INV_X1 U647 ( .A(n619), .ZN(n607) );
  NOR2_X1 U648 ( .A1(n651), .A2(n652), .ZN(n619) );
  AND2_X1 U649 ( .A1(n653), .A2(n654), .ZN(n652) );
  NAND2_X1 U650 ( .A1(n655), .A2(n656), .ZN(n653) );
  NAND2_X1 U651 ( .A1(n614), .A2(n657), .ZN(n648) );
  NAND2_X1 U652 ( .A1(n608), .A2(n658), .ZN(n646) );
  NOR2_X1 U653 ( .A1(n659), .A2(n610), .ZN(n644) );
  NAND2_X1 U654 ( .A1(n660), .A2(n661), .ZN(Result_7_) );
  NAND2_X1 U655 ( .A1(n662), .A2(n592), .ZN(n661) );
  XOR2_X1 U656 ( .A(n663), .B(n664), .Z(n662) );
  NAND2_X1 U657 ( .A1(n660), .A2(n665), .ZN(Result_6_) );
  NAND2_X1 U658 ( .A1(n666), .A2(n592), .ZN(n665) );
  NOR2_X1 U659 ( .A1(n667), .A2(n668), .ZN(n666) );
  NOR2_X1 U660 ( .A1(n669), .A2(n670), .ZN(n668) );
  NAND2_X1 U661 ( .A1(n660), .A2(n671), .ZN(Result_5_) );
  NAND2_X1 U662 ( .A1(n592), .A2(n672), .ZN(n671) );
  XNOR2_X1 U663 ( .A(n667), .B(n673), .ZN(n672) );
  NAND2_X1 U664 ( .A1(n674), .A2(n675), .ZN(n673) );
  NAND2_X1 U665 ( .A1(n676), .A2(n677), .ZN(n675) );
  INV_X1 U666 ( .A(n678), .ZN(n677) );
  NAND2_X1 U667 ( .A1(n679), .A2(n680), .ZN(n676) );
  NAND2_X1 U668 ( .A1(n660), .A2(n681), .ZN(Result_4_) );
  NAND2_X1 U669 ( .A1(n682), .A2(n592), .ZN(n681) );
  XOR2_X1 U670 ( .A(n683), .B(n684), .Z(n682) );
  NAND2_X1 U671 ( .A1(n660), .A2(n685), .ZN(Result_3_) );
  NAND2_X1 U672 ( .A1(n592), .A2(n686), .ZN(n685) );
  XOR2_X1 U673 ( .A(n687), .B(n688), .Z(n686) );
  AND2_X1 U674 ( .A1(n689), .A2(n690), .ZN(n687) );
  NAND2_X1 U675 ( .A1(n660), .A2(n691), .ZN(Result_2_) );
  NAND2_X1 U676 ( .A1(n692), .A2(n592), .ZN(n691) );
  XOR2_X1 U677 ( .A(n693), .B(n694), .Z(n692) );
  AND2_X1 U678 ( .A1(n695), .A2(n696), .ZN(n694) );
  NAND2_X1 U679 ( .A1(n660), .A2(n697), .ZN(Result_1_) );
  NAND2_X1 U680 ( .A1(n698), .A2(n592), .ZN(n697) );
  XNOR2_X1 U681 ( .A(n699), .B(n700), .ZN(n698) );
  NOR2_X1 U682 ( .A1(n701), .A2(n702), .ZN(n700) );
  NAND2_X1 U683 ( .A1(n703), .A2(n704), .ZN(Result_15_) );
  NAND2_X1 U684 ( .A1(n592), .A2(n705), .ZN(n704) );
  NAND2_X1 U685 ( .A1(n706), .A2(n707), .ZN(n703) );
  NAND2_X1 U686 ( .A1(n708), .A2(n610), .ZN(n707) );
  NOR2_X1 U687 ( .A1(n608), .A2(n606), .ZN(n708) );
  NAND2_X1 U688 ( .A1(n709), .A2(n710), .ZN(n706) );
  NAND2_X1 U689 ( .A1(n711), .A2(n712), .ZN(Result_14_) );
  NAND2_X1 U690 ( .A1(n592), .A2(n713), .ZN(n712) );
  NAND2_X1 U691 ( .A1(n714), .A2(n715), .ZN(n713) );
  NOR2_X1 U692 ( .A1(n716), .A2(n717), .ZN(n715) );
  NOR2_X1 U693 ( .A1(n718), .A2(n719), .ZN(n717) );
  NOR2_X1 U694 ( .A1(n720), .A2(n721), .ZN(n716) );
  NOR2_X1 U695 ( .A1(n722), .A2(n723), .ZN(n714) );
  NOR2_X1 U696 ( .A1(n724), .A2(n710), .ZN(n723) );
  NOR2_X1 U697 ( .A1(n725), .A2(n709), .ZN(n722) );
  NOR2_X1 U698 ( .A1(n726), .A2(n727), .ZN(n711) );
  NOR2_X1 U699 ( .A1(n728), .A2(n729), .ZN(n727) );
  NOR2_X1 U700 ( .A1(n730), .A2(n731), .ZN(n728) );
  NAND2_X1 U701 ( .A1(n732), .A2(n733), .ZN(n731) );
  NAND2_X1 U702 ( .A1(n606), .A2(n705), .ZN(n733) );
  NAND2_X1 U703 ( .A1(n734), .A2(n608), .ZN(n732) );
  INV_X1 U704 ( .A(n709), .ZN(n734) );
  NOR2_X1 U705 ( .A1(n610), .A2(n710), .ZN(n730) );
  NOR2_X1 U706 ( .A1(n735), .A2(n736), .ZN(n726) );
  NOR2_X1 U707 ( .A1(n737), .A2(n738), .ZN(n736) );
  NAND2_X1 U708 ( .A1(n739), .A2(n740), .ZN(n738) );
  NAND2_X1 U709 ( .A1(n606), .A2(n741), .ZN(n740) );
  NAND2_X1 U710 ( .A1(n608), .A2(n709), .ZN(n739) );
  AND2_X1 U711 ( .A1(n710), .A2(n742), .ZN(n737) );
  INV_X1 U712 ( .A(n729), .ZN(n735) );
  NAND2_X1 U713 ( .A1(n719), .A2(n721), .ZN(n729) );
  NAND2_X1 U714 ( .A1(n743), .A2(n744), .ZN(Result_13_) );
  NAND2_X1 U715 ( .A1(n592), .A2(n745), .ZN(n744) );
  XNOR2_X1 U716 ( .A(n746), .B(n747), .ZN(n745) );
  NAND2_X1 U717 ( .A1(n748), .A2(n749), .ZN(n746) );
  NOR2_X1 U718 ( .A1(n750), .A2(n751), .ZN(n743) );
  NOR2_X1 U719 ( .A1(n752), .A2(n753), .ZN(n751) );
  NOR2_X1 U720 ( .A1(n754), .A2(n755), .ZN(n752) );
  NAND2_X1 U721 ( .A1(n756), .A2(n757), .ZN(n755) );
  NAND2_X1 U722 ( .A1(n606), .A2(n758), .ZN(n757) );
  NAND2_X1 U723 ( .A1(n608), .A2(n759), .ZN(n756) );
  NOR2_X1 U724 ( .A1(n760), .A2(n610), .ZN(n754) );
  NOR2_X1 U725 ( .A1(n761), .A2(n762), .ZN(n750) );
  INV_X1 U726 ( .A(n753), .ZN(n762) );
  XNOR2_X1 U727 ( .A(n763), .B(a_5_), .ZN(n753) );
  NOR2_X1 U728 ( .A1(n764), .A2(n765), .ZN(n761) );
  NAND2_X1 U729 ( .A1(n766), .A2(n767), .ZN(n765) );
  NAND2_X1 U730 ( .A1(n768), .A2(n606), .ZN(n767) );
  INV_X1 U731 ( .A(n758), .ZN(n768) );
  NAND2_X1 U732 ( .A1(n608), .A2(n769), .ZN(n766) );
  NOR2_X1 U733 ( .A1(n770), .A2(n610), .ZN(n764) );
  NAND2_X1 U734 ( .A1(n771), .A2(n772), .ZN(Result_12_) );
  NAND2_X1 U735 ( .A1(n773), .A2(n592), .ZN(n772) );
  XNOR2_X1 U736 ( .A(n774), .B(n775), .ZN(n773) );
  XNOR2_X1 U737 ( .A(n776), .B(n777), .ZN(n775) );
  NOR2_X1 U738 ( .A1(n778), .A2(n779), .ZN(n771) );
  NOR2_X1 U739 ( .A1(n780), .A2(n781), .ZN(n779) );
  NOR2_X1 U740 ( .A1(n782), .A2(n783), .ZN(n780) );
  NAND2_X1 U741 ( .A1(n784), .A2(n785), .ZN(n783) );
  NAND2_X1 U742 ( .A1(n606), .A2(n786), .ZN(n785) );
  NAND2_X1 U743 ( .A1(n608), .A2(n787), .ZN(n784) );
  NOR2_X1 U744 ( .A1(n788), .A2(n610), .ZN(n782) );
  NOR2_X1 U745 ( .A1(n789), .A2(n790), .ZN(n778) );
  INV_X1 U746 ( .A(n781), .ZN(n790) );
  XNOR2_X1 U747 ( .A(n791), .B(a_4_), .ZN(n781) );
  NOR2_X1 U748 ( .A1(n792), .A2(n793), .ZN(n789) );
  NAND2_X1 U749 ( .A1(n794), .A2(n795), .ZN(n793) );
  NAND2_X1 U750 ( .A1(n796), .A2(n606), .ZN(n795) );
  INV_X1 U751 ( .A(n786), .ZN(n796) );
  NAND2_X1 U752 ( .A1(n608), .A2(n797), .ZN(n794) );
  NOR2_X1 U753 ( .A1(n798), .A2(n610), .ZN(n792) );
  NAND2_X1 U754 ( .A1(n799), .A2(n800), .ZN(Result_11_) );
  NAND2_X1 U755 ( .A1(n801), .A2(n592), .ZN(n800) );
  XNOR2_X1 U756 ( .A(n802), .B(n803), .ZN(n801) );
  XOR2_X1 U757 ( .A(n804), .B(n805), .Z(n803) );
  NAND2_X1 U758 ( .A1(b_7_), .A2(a_3_), .ZN(n805) );
  NOR2_X1 U759 ( .A1(n806), .A2(n807), .ZN(n799) );
  NOR2_X1 U760 ( .A1(n808), .A2(n809), .ZN(n807) );
  NOR2_X1 U761 ( .A1(n810), .A2(n811), .ZN(n808) );
  NAND2_X1 U762 ( .A1(n812), .A2(n813), .ZN(n811) );
  NAND2_X1 U763 ( .A1(n606), .A2(n814), .ZN(n813) );
  NAND2_X1 U764 ( .A1(n608), .A2(n815), .ZN(n812) );
  NOR2_X1 U765 ( .A1(n816), .A2(n610), .ZN(n810) );
  NOR2_X1 U766 ( .A1(n817), .A2(n818), .ZN(n806) );
  INV_X1 U767 ( .A(n809), .ZN(n818) );
  XNOR2_X1 U768 ( .A(n819), .B(a_3_), .ZN(n809) );
  NOR2_X1 U769 ( .A1(n820), .A2(n821), .ZN(n817) );
  NAND2_X1 U770 ( .A1(n822), .A2(n823), .ZN(n821) );
  NAND2_X1 U771 ( .A1(n824), .A2(n606), .ZN(n823) );
  INV_X1 U772 ( .A(n814), .ZN(n824) );
  NAND2_X1 U773 ( .A1(n608), .A2(n825), .ZN(n822) );
  NOR2_X1 U774 ( .A1(n826), .A2(n610), .ZN(n820) );
  NAND2_X1 U775 ( .A1(n827), .A2(n828), .ZN(Result_10_) );
  NAND2_X1 U776 ( .A1(n592), .A2(n829), .ZN(n828) );
  XNOR2_X1 U777 ( .A(n830), .B(n831), .ZN(n829) );
  XOR2_X1 U778 ( .A(n832), .B(n833), .Z(n831) );
  NAND2_X1 U779 ( .A1(b_7_), .A2(a_2_), .ZN(n833) );
  NOR2_X1 U780 ( .A1(n834), .A2(n835), .ZN(n827) );
  NOR2_X1 U781 ( .A1(n836), .A2(n837), .ZN(n835) );
  NOR2_X1 U782 ( .A1(n838), .A2(n839), .ZN(n836) );
  NAND2_X1 U783 ( .A1(n840), .A2(n841), .ZN(n839) );
  NAND2_X1 U784 ( .A1(n606), .A2(n654), .ZN(n841) );
  INV_X1 U785 ( .A(n842), .ZN(n654) );
  NAND2_X1 U786 ( .A1(n608), .A2(n843), .ZN(n840) );
  NOR2_X1 U787 ( .A1(n844), .A2(n610), .ZN(n838) );
  NOR2_X1 U788 ( .A1(n845), .A2(n846), .ZN(n834) );
  INV_X1 U789 ( .A(n837), .ZN(n846) );
  XNOR2_X1 U790 ( .A(n655), .B(a_2_), .ZN(n837) );
  NOR2_X1 U791 ( .A1(n847), .A2(n848), .ZN(n845) );
  NAND2_X1 U792 ( .A1(n849), .A2(n850), .ZN(n848) );
  NAND2_X1 U793 ( .A1(n842), .A2(n606), .ZN(n850) );
  NOR2_X1 U794 ( .A1(n851), .A2(n852), .ZN(n842) );
  AND2_X1 U795 ( .A1(n853), .A2(n814), .ZN(n852) );
  NAND2_X1 U796 ( .A1(n854), .A2(n855), .ZN(n814) );
  NAND2_X1 U797 ( .A1(n856), .A2(n786), .ZN(n855) );
  NAND2_X1 U798 ( .A1(n857), .A2(n858), .ZN(n786) );
  NAND2_X1 U799 ( .A1(n859), .A2(n758), .ZN(n858) );
  NAND2_X1 U800 ( .A1(n860), .A2(n861), .ZN(n758) );
  NAND2_X1 U801 ( .A1(n705), .A2(n862), .ZN(n861) );
  NAND2_X1 U802 ( .A1(n724), .A2(n725), .ZN(n862) );
  NAND2_X1 U803 ( .A1(n763), .A2(n863), .ZN(n859) );
  NAND2_X1 U804 ( .A1(n791), .A2(n864), .ZN(n856) );
  NAND2_X1 U805 ( .A1(n819), .A2(n865), .ZN(n853) );
  NAND2_X1 U806 ( .A1(n608), .A2(n866), .ZN(n849) );
  NOR2_X1 U807 ( .A1(n867), .A2(n610), .ZN(n847) );
  NAND2_X1 U808 ( .A1(n660), .A2(n868), .ZN(Result_0_) );
  NAND2_X1 U809 ( .A1(n592), .A2(n869), .ZN(n868) );
  NAND2_X1 U810 ( .A1(n870), .A2(n871), .ZN(n869) );
  NAND2_X1 U811 ( .A1(a_0_), .A2(n872), .ZN(n871) );
  NOR2_X1 U812 ( .A1(n702), .A2(n873), .ZN(n870) );
  NOR2_X1 U813 ( .A1(n699), .A2(n701), .ZN(n873) );
  AND2_X1 U814 ( .A1(n874), .A2(n875), .ZN(n701) );
  OR2_X1 U815 ( .A1(n876), .A2(n877), .ZN(n875) );
  XOR2_X1 U816 ( .A(n872), .B(n878), .Z(n874) );
  AND2_X1 U817 ( .A1(n696), .A2(n879), .ZN(n699) );
  NAND2_X1 U818 ( .A1(n695), .A2(n693), .ZN(n879) );
  NAND2_X1 U819 ( .A1(n690), .A2(n880), .ZN(n693) );
  NAND2_X1 U820 ( .A1(n688), .A2(n689), .ZN(n880) );
  NAND2_X1 U821 ( .A1(n881), .A2(n882), .ZN(n689) );
  NAND2_X1 U822 ( .A1(n883), .A2(n884), .ZN(n882) );
  AND2_X1 U823 ( .A1(n683), .A2(n684), .ZN(n688) );
  NAND2_X1 U824 ( .A1(n885), .A2(n886), .ZN(n684) );
  NAND2_X1 U825 ( .A1(n667), .A2(n678), .ZN(n886) );
  AND2_X1 U826 ( .A1(n669), .A2(n670), .ZN(n667) );
  XOR2_X1 U827 ( .A(n680), .B(n679), .Z(n670) );
  NOR2_X1 U828 ( .A1(n663), .A2(n664), .ZN(n669) );
  XOR2_X1 U829 ( .A(n887), .B(n888), .Z(n664) );
  NAND2_X1 U830 ( .A1(n889), .A2(n890), .ZN(n887) );
  AND2_X1 U831 ( .A1(n891), .A2(n892), .ZN(n663) );
  NAND2_X1 U832 ( .A1(n628), .A2(n893), .ZN(n892) );
  OR2_X1 U833 ( .A1(n626), .A2(n627), .ZN(n893) );
  NOR2_X1 U834 ( .A1(n894), .A2(n720), .ZN(n628) );
  NAND2_X1 U835 ( .A1(n626), .A2(n627), .ZN(n891) );
  NAND2_X1 U836 ( .A1(n895), .A2(n896), .ZN(n627) );
  NAND2_X1 U837 ( .A1(n597), .A2(n897), .ZN(n896) );
  OR2_X1 U838 ( .A1(n596), .A2(n594), .ZN(n897) );
  NOR2_X1 U839 ( .A1(n657), .A2(n720), .ZN(n597) );
  NAND2_X1 U840 ( .A1(n594), .A2(n596), .ZN(n895) );
  NAND2_X1 U841 ( .A1(n898), .A2(n899), .ZN(n596) );
  NAND2_X1 U842 ( .A1(n900), .A2(b_7_), .ZN(n899) );
  NOR2_X1 U843 ( .A1(n901), .A2(n656), .ZN(n900) );
  NOR2_X1 U844 ( .A1(n830), .A2(n832), .ZN(n901) );
  NAND2_X1 U845 ( .A1(n830), .A2(n832), .ZN(n898) );
  NAND2_X1 U846 ( .A1(n902), .A2(n903), .ZN(n832) );
  NAND2_X1 U847 ( .A1(n904), .A2(b_7_), .ZN(n903) );
  NOR2_X1 U848 ( .A1(n905), .A2(n865), .ZN(n904) );
  NOR2_X1 U849 ( .A1(n802), .A2(n804), .ZN(n905) );
  NAND2_X1 U850 ( .A1(n802), .A2(n804), .ZN(n902) );
  NAND2_X1 U851 ( .A1(n906), .A2(n907), .ZN(n804) );
  NAND2_X1 U852 ( .A1(n777), .A2(n908), .ZN(n907) );
  OR2_X1 U853 ( .A1(n776), .A2(n774), .ZN(n908) );
  NOR2_X1 U854 ( .A1(n720), .A2(n864), .ZN(n777) );
  NAND2_X1 U855 ( .A1(n774), .A2(n776), .ZN(n906) );
  NAND2_X1 U856 ( .A1(n748), .A2(n909), .ZN(n776) );
  NAND2_X1 U857 ( .A1(n747), .A2(n749), .ZN(n909) );
  NAND2_X1 U858 ( .A1(n910), .A2(n911), .ZN(n749) );
  NAND2_X1 U859 ( .A1(b_7_), .A2(a_5_), .ZN(n910) );
  XNOR2_X1 U860 ( .A(n860), .B(n912), .ZN(n747) );
  OR2_X1 U861 ( .A1(n911), .A2(n863), .ZN(n748) );
  NAND2_X1 U862 ( .A1(n705), .A2(n913), .ZN(n911) );
  INV_X1 U863 ( .A(n741), .ZN(n705) );
  NAND2_X1 U864 ( .A1(b_7_), .A2(a_7_), .ZN(n741) );
  XNOR2_X1 U865 ( .A(n914), .B(n915), .ZN(n774) );
  NAND2_X1 U866 ( .A1(n916), .A2(n917), .ZN(n914) );
  XNOR2_X1 U867 ( .A(n918), .B(n919), .ZN(n802) );
  NAND2_X1 U868 ( .A1(n920), .A2(n921), .ZN(n918) );
  XOR2_X1 U869 ( .A(n922), .B(n923), .Z(n830) );
  XNOR2_X1 U870 ( .A(n924), .B(n925), .ZN(n922) );
  NAND2_X1 U871 ( .A1(b_6_), .A2(a_3_), .ZN(n924) );
  XNOR2_X1 U872 ( .A(n926), .B(n927), .ZN(n594) );
  XOR2_X1 U873 ( .A(n928), .B(n929), .Z(n927) );
  NAND2_X1 U874 ( .A1(a_2_), .A2(b_6_), .ZN(n929) );
  XOR2_X1 U875 ( .A(n930), .B(n931), .Z(n626) );
  XOR2_X1 U876 ( .A(n932), .B(n933), .Z(n931) );
  NOR2_X1 U877 ( .A1(n934), .A2(n935), .ZN(n885) );
  INV_X1 U878 ( .A(n674), .ZN(n934) );
  NAND2_X1 U879 ( .A1(n936), .A2(n678), .ZN(n674) );
  NOR2_X1 U880 ( .A1(n935), .A2(n937), .ZN(n678) );
  AND2_X1 U881 ( .A1(n938), .A2(n939), .ZN(n937) );
  NOR2_X1 U882 ( .A1(n939), .A2(n938), .ZN(n935) );
  AND2_X1 U883 ( .A1(n940), .A2(n941), .ZN(n938) );
  NAND2_X1 U884 ( .A1(n942), .A2(n943), .ZN(n941) );
  XNOR2_X1 U885 ( .A(n944), .B(n945), .ZN(n939) );
  XNOR2_X1 U886 ( .A(n946), .B(n947), .ZN(n944) );
  AND2_X1 U887 ( .A1(n680), .A2(n679), .ZN(n936) );
  XNOR2_X1 U888 ( .A(n948), .B(n942), .ZN(n679) );
  XNOR2_X1 U889 ( .A(n949), .B(n950), .ZN(n942) );
  NAND2_X1 U890 ( .A1(n951), .A2(n952), .ZN(n949) );
  NAND2_X1 U891 ( .A1(n940), .A2(n943), .ZN(n948) );
  NAND2_X1 U892 ( .A1(n953), .A2(n954), .ZN(n943) );
  NAND2_X1 U893 ( .A1(a_0_), .A2(b_5_), .ZN(n954) );
  INV_X1 U894 ( .A(n955), .ZN(n953) );
  NAND2_X1 U895 ( .A1(a_0_), .A2(n955), .ZN(n940) );
  NAND2_X1 U896 ( .A1(n956), .A2(n957), .ZN(n955) );
  NAND2_X1 U897 ( .A1(n958), .A2(n959), .ZN(n957) );
  OR2_X1 U898 ( .A1(n960), .A2(n961), .ZN(n959) );
  NAND2_X1 U899 ( .A1(n961), .A2(n960), .ZN(n956) );
  NAND2_X1 U900 ( .A1(n889), .A2(n962), .ZN(n680) );
  NAND2_X1 U901 ( .A1(n888), .A2(n890), .ZN(n962) );
  NAND2_X1 U902 ( .A1(n963), .A2(n964), .ZN(n890) );
  NAND2_X1 U903 ( .A1(a_0_), .A2(b_6_), .ZN(n964) );
  INV_X1 U904 ( .A(n965), .ZN(n963) );
  XNOR2_X1 U905 ( .A(n961), .B(n966), .ZN(n888) );
  XNOR2_X1 U906 ( .A(n960), .B(n958), .ZN(n966) );
  NOR2_X1 U907 ( .A1(n657), .A2(n763), .ZN(n958) );
  NAND2_X1 U908 ( .A1(n967), .A2(n968), .ZN(n960) );
  NAND2_X1 U909 ( .A1(n969), .A2(a_2_), .ZN(n968) );
  NOR2_X1 U910 ( .A1(n970), .A2(n763), .ZN(n969) );
  NOR2_X1 U911 ( .A1(n971), .A2(n972), .ZN(n970) );
  NAND2_X1 U912 ( .A1(n972), .A2(n971), .ZN(n967) );
  XOR2_X1 U913 ( .A(n973), .B(n974), .Z(n961) );
  NOR2_X1 U914 ( .A1(n975), .A2(n976), .ZN(n974) );
  NOR2_X1 U915 ( .A1(n977), .A2(n978), .ZN(n975) );
  NOR2_X1 U916 ( .A1(n791), .A2(n656), .ZN(n978) );
  INV_X1 U917 ( .A(n979), .ZN(n977) );
  NAND2_X1 U918 ( .A1(a_0_), .A2(n965), .ZN(n889) );
  NAND2_X1 U919 ( .A1(n980), .A2(n981), .ZN(n965) );
  NAND2_X1 U920 ( .A1(n933), .A2(n982), .ZN(n981) );
  NAND2_X1 U921 ( .A1(n932), .A2(n930), .ZN(n982) );
  NOR2_X1 U922 ( .A1(n657), .A2(n724), .ZN(n933) );
  OR2_X1 U923 ( .A1(n930), .A2(n932), .ZN(n980) );
  AND2_X1 U924 ( .A1(n983), .A2(n984), .ZN(n932) );
  NAND2_X1 U925 ( .A1(n985), .A2(a_2_), .ZN(n984) );
  NOR2_X1 U926 ( .A1(n986), .A2(n724), .ZN(n985) );
  NOR2_X1 U927 ( .A1(n928), .A2(n926), .ZN(n986) );
  NAND2_X1 U928 ( .A1(n926), .A2(n928), .ZN(n983) );
  NAND2_X1 U929 ( .A1(n987), .A2(n988), .ZN(n928) );
  NAND2_X1 U930 ( .A1(n989), .A2(b_6_), .ZN(n988) );
  NOR2_X1 U931 ( .A1(n990), .A2(n865), .ZN(n989) );
  NOR2_X1 U932 ( .A1(n923), .A2(n925), .ZN(n990) );
  NAND2_X1 U933 ( .A1(n923), .A2(n925), .ZN(n987) );
  NAND2_X1 U934 ( .A1(n920), .A2(n991), .ZN(n925) );
  NAND2_X1 U935 ( .A1(n919), .A2(n921), .ZN(n991) );
  NAND2_X1 U936 ( .A1(n992), .A2(n993), .ZN(n921) );
  NAND2_X1 U937 ( .A1(b_6_), .A2(a_4_), .ZN(n993) );
  INV_X1 U938 ( .A(n994), .ZN(n992) );
  XOR2_X1 U939 ( .A(n995), .B(n996), .Z(n919) );
  XOR2_X1 U940 ( .A(n857), .B(n997), .Z(n995) );
  NAND2_X1 U941 ( .A1(a_4_), .A2(n994), .ZN(n920) );
  NAND2_X1 U942 ( .A1(n916), .A2(n998), .ZN(n994) );
  NAND2_X1 U943 ( .A1(n915), .A2(n917), .ZN(n998) );
  NAND2_X1 U944 ( .A1(n999), .A2(n1000), .ZN(n917) );
  NAND2_X1 U945 ( .A1(b_6_), .A2(a_5_), .ZN(n999) );
  XOR2_X1 U946 ( .A(n1001), .B(n1002), .Z(n915) );
  OR2_X1 U947 ( .A1(n1000), .A2(n863), .ZN(n916) );
  NAND2_X1 U948 ( .A1(n912), .A2(n913), .ZN(n1000) );
  INV_X1 U949 ( .A(n860), .ZN(n913) );
  NAND2_X1 U950 ( .A1(b_6_), .A2(a_6_), .ZN(n860) );
  NOR2_X1 U951 ( .A1(n718), .A2(n763), .ZN(n912) );
  XNOR2_X1 U952 ( .A(n1003), .B(n1004), .ZN(n923) );
  NAND2_X1 U953 ( .A1(n1005), .A2(n1006), .ZN(n1003) );
  XOR2_X1 U954 ( .A(n1007), .B(n1008), .Z(n926) );
  XOR2_X1 U955 ( .A(n1009), .B(n1010), .Z(n1007) );
  NOR2_X1 U956 ( .A1(n763), .A2(n865), .ZN(n1010) );
  XOR2_X1 U957 ( .A(n972), .B(n1011), .Z(n930) );
  XOR2_X1 U958 ( .A(n971), .B(n1012), .Z(n1011) );
  NAND2_X1 U959 ( .A1(a_2_), .A2(b_5_), .ZN(n1012) );
  NAND2_X1 U960 ( .A1(n1013), .A2(n1014), .ZN(n971) );
  NAND2_X1 U961 ( .A1(n1015), .A2(a_3_), .ZN(n1014) );
  NOR2_X1 U962 ( .A1(n1016), .A2(n763), .ZN(n1015) );
  NOR2_X1 U963 ( .A1(n1008), .A2(n1009), .ZN(n1016) );
  NAND2_X1 U964 ( .A1(n1008), .A2(n1009), .ZN(n1013) );
  NAND2_X1 U965 ( .A1(n1005), .A2(n1017), .ZN(n1009) );
  NAND2_X1 U966 ( .A1(n1004), .A2(n1006), .ZN(n1017) );
  NAND2_X1 U967 ( .A1(n1018), .A2(n1019), .ZN(n1006) );
  NAND2_X1 U968 ( .A1(b_5_), .A2(a_4_), .ZN(n1019) );
  INV_X1 U969 ( .A(n1020), .ZN(n1018) );
  XNOR2_X1 U970 ( .A(n1021), .B(n1022), .ZN(n1004) );
  NAND2_X1 U971 ( .A1(n1023), .A2(n1024), .ZN(n1021) );
  NAND2_X1 U972 ( .A1(a_4_), .A2(n1020), .ZN(n1005) );
  NAND2_X1 U973 ( .A1(n1025), .A2(n1026), .ZN(n1020) );
  NAND2_X1 U974 ( .A1(n997), .A2(n1027), .ZN(n1026) );
  NAND2_X1 U975 ( .A1(n996), .A2(n857), .ZN(n1027) );
  AND2_X1 U976 ( .A1(n1001), .A2(n1002), .ZN(n997) );
  NOR2_X1 U977 ( .A1(n763), .A2(n725), .ZN(n1001) );
  OR2_X1 U978 ( .A1(n857), .A2(n996), .ZN(n1025) );
  NAND2_X1 U979 ( .A1(n1028), .A2(n1029), .ZN(n996) );
  NAND2_X1 U980 ( .A1(n1030), .A2(n1031), .ZN(n1029) );
  NAND2_X1 U981 ( .A1(b_3_), .A2(a_7_), .ZN(n1031) );
  NAND2_X1 U982 ( .A1(b_4_), .A2(a_6_), .ZN(n1030) );
  NAND2_X1 U983 ( .A1(b_5_), .A2(a_5_), .ZN(n857) );
  XOR2_X1 U984 ( .A(n1032), .B(n1033), .Z(n1008) );
  XOR2_X1 U985 ( .A(n854), .B(n1034), .Z(n1033) );
  XNOR2_X1 U986 ( .A(n1035), .B(n1036), .ZN(n972) );
  XOR2_X1 U987 ( .A(n1037), .B(n1038), .Z(n1036) );
  XOR2_X1 U988 ( .A(n883), .B(n884), .Z(n683) );
  INV_X1 U989 ( .A(n1039), .ZN(n884) );
  NAND2_X1 U990 ( .A1(n1040), .A2(n883), .ZN(n690) );
  AND2_X1 U991 ( .A1(n1041), .A2(n1042), .ZN(n883) );
  NAND2_X1 U992 ( .A1(n946), .A2(n1043), .ZN(n1042) );
  NAND2_X1 U993 ( .A1(n945), .A2(n947), .ZN(n1043) );
  AND2_X1 U994 ( .A1(n951), .A2(n1044), .ZN(n946) );
  NAND2_X1 U995 ( .A1(n950), .A2(n952), .ZN(n1044) );
  NAND2_X1 U996 ( .A1(n1045), .A2(n1046), .ZN(n952) );
  NAND2_X1 U997 ( .A1(a_1_), .A2(b_4_), .ZN(n1046) );
  XNOR2_X1 U998 ( .A(n1047), .B(n1048), .ZN(n950) );
  XOR2_X1 U999 ( .A(n1049), .B(n1050), .Z(n1047) );
  NAND2_X1 U1000 ( .A1(a_2_), .A2(b_3_), .ZN(n1049) );
  OR2_X1 U1001 ( .A1(n657), .A2(n1045), .ZN(n951) );
  NOR2_X1 U1002 ( .A1(n976), .A2(n1051), .ZN(n1045) );
  AND2_X1 U1003 ( .A1(n973), .A2(n1052), .ZN(n1051) );
  NAND2_X1 U1004 ( .A1(n979), .A2(n1053), .ZN(n1052) );
  NAND2_X1 U1005 ( .A1(a_2_), .A2(b_4_), .ZN(n1053) );
  XNOR2_X1 U1006 ( .A(n1054), .B(n1055), .ZN(n973) );
  XOR2_X1 U1007 ( .A(n851), .B(n1056), .Z(n1055) );
  NOR2_X1 U1008 ( .A1(n979), .A2(n656), .ZN(n976) );
  NAND2_X1 U1009 ( .A1(n1057), .A2(n1058), .ZN(n979) );
  NAND2_X1 U1010 ( .A1(n1035), .A2(n1059), .ZN(n1058) );
  OR2_X1 U1011 ( .A1(n1038), .A2(n1037), .ZN(n1059) );
  XOR2_X1 U1012 ( .A(n1060), .B(n1061), .Z(n1035) );
  NAND2_X1 U1013 ( .A1(n1062), .A2(n1063), .ZN(n1060) );
  NAND2_X1 U1014 ( .A1(n1038), .A2(n1037), .ZN(n1057) );
  NAND2_X1 U1015 ( .A1(n1064), .A2(n1065), .ZN(n1037) );
  NAND2_X1 U1016 ( .A1(n1032), .A2(n1066), .ZN(n1065) );
  NAND2_X1 U1017 ( .A1(n1067), .A2(n1034), .ZN(n1066) );
  XOR2_X1 U1018 ( .A(n1068), .B(n1069), .Z(n1032) );
  NAND2_X1 U1019 ( .A1(n1070), .A2(n1071), .ZN(n1068) );
  OR2_X1 U1020 ( .A1(n1034), .A2(n1067), .ZN(n1064) );
  INV_X1 U1021 ( .A(n854), .ZN(n1067) );
  NAND2_X1 U1022 ( .A1(b_4_), .A2(a_4_), .ZN(n854) );
  NAND2_X1 U1023 ( .A1(n1023), .A2(n1072), .ZN(n1034) );
  NAND2_X1 U1024 ( .A1(n1022), .A2(n1024), .ZN(n1072) );
  NAND2_X1 U1025 ( .A1(n1028), .A2(n1073), .ZN(n1024) );
  NAND2_X1 U1026 ( .A1(b_4_), .A2(a_5_), .ZN(n1073) );
  AND2_X1 U1027 ( .A1(n1074), .A2(n1075), .ZN(n1022) );
  NAND2_X1 U1028 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
  OR2_X1 U1029 ( .A1(n1028), .A2(n863), .ZN(n1023) );
  NAND2_X1 U1030 ( .A1(n1002), .A2(n1078), .ZN(n1028) );
  INV_X1 U1031 ( .A(n1076), .ZN(n1078) );
  NOR2_X1 U1032 ( .A1(n791), .A2(n718), .ZN(n1002) );
  NAND2_X1 U1033 ( .A1(a_3_), .A2(b_4_), .ZN(n1038) );
  OR2_X1 U1034 ( .A1(n945), .A2(n947), .ZN(n1041) );
  NOR2_X1 U1035 ( .A1(n894), .A2(n791), .ZN(n947) );
  XOR2_X1 U1036 ( .A(n1079), .B(n1080), .Z(n945) );
  XNOR2_X1 U1037 ( .A(n1081), .B(n1082), .ZN(n1079) );
  NOR2_X1 U1038 ( .A1(n1039), .A2(n881), .ZN(n1040) );
  XOR2_X1 U1039 ( .A(n1083), .B(n1084), .Z(n881) );
  XNOR2_X1 U1040 ( .A(n1085), .B(n1086), .ZN(n1039) );
  XNOR2_X1 U1041 ( .A(n1087), .B(n1088), .ZN(n1086) );
  NAND2_X1 U1042 ( .A1(a_0_), .A2(b_3_), .ZN(n1088) );
  NAND2_X1 U1043 ( .A1(n1089), .A2(n1090), .ZN(n695) );
  NAND2_X1 U1044 ( .A1(n1083), .A2(n1091), .ZN(n1090) );
  NAND2_X1 U1045 ( .A1(n1092), .A2(n1083), .ZN(n696) );
  XNOR2_X1 U1046 ( .A(n1093), .B(n1094), .ZN(n1083) );
  NAND2_X1 U1047 ( .A1(n1095), .A2(n1096), .ZN(n1093) );
  NOR2_X1 U1048 ( .A1(n1084), .A2(n1089), .ZN(n1092) );
  XNOR2_X1 U1049 ( .A(n877), .B(n876), .ZN(n1089) );
  INV_X1 U1050 ( .A(n1091), .ZN(n1084) );
  NAND2_X1 U1051 ( .A1(n1097), .A2(n1098), .ZN(n1091) );
  NAND2_X1 U1052 ( .A1(n1099), .A2(a_0_), .ZN(n1098) );
  NOR2_X1 U1053 ( .A1(n1100), .A2(n819), .ZN(n1099) );
  NOR2_X1 U1054 ( .A1(n1087), .A2(n1085), .ZN(n1100) );
  NAND2_X1 U1055 ( .A1(n1087), .A2(n1085), .ZN(n1097) );
  XOR2_X1 U1056 ( .A(n1101), .B(n1102), .Z(n1085) );
  XOR2_X1 U1057 ( .A(n1103), .B(n1104), .Z(n1101) );
  AND2_X1 U1058 ( .A1(n1105), .A2(n1106), .ZN(n1087) );
  NAND2_X1 U1059 ( .A1(n1082), .A2(n1107), .ZN(n1106) );
  NAND2_X1 U1060 ( .A1(n1081), .A2(n1080), .ZN(n1107) );
  AND2_X1 U1061 ( .A1(n1108), .A2(n1109), .ZN(n1082) );
  NAND2_X1 U1062 ( .A1(n1110), .A2(a_2_), .ZN(n1109) );
  NOR2_X1 U1063 ( .A1(n1111), .A2(n819), .ZN(n1110) );
  NOR2_X1 U1064 ( .A1(n1050), .A2(n1048), .ZN(n1111) );
  NAND2_X1 U1065 ( .A1(n1050), .A2(n1048), .ZN(n1108) );
  XOR2_X1 U1066 ( .A(n1112), .B(n1113), .Z(n1048) );
  XOR2_X1 U1067 ( .A(n1114), .B(n1115), .Z(n1112) );
  NOR2_X1 U1068 ( .A1(n655), .A2(n865), .ZN(n1115) );
  AND2_X1 U1069 ( .A1(n1116), .A2(n1117), .ZN(n1050) );
  NAND2_X1 U1070 ( .A1(n1056), .A2(n1118), .ZN(n1117) );
  NAND2_X1 U1071 ( .A1(n851), .A2(n1054), .ZN(n1118) );
  AND2_X1 U1072 ( .A1(n1062), .A2(n1119), .ZN(n1056) );
  NAND2_X1 U1073 ( .A1(n1061), .A2(n1063), .ZN(n1119) );
  NAND2_X1 U1074 ( .A1(n1120), .A2(n1121), .ZN(n1063) );
  NAND2_X1 U1075 ( .A1(a_4_), .A2(b_3_), .ZN(n1121) );
  INV_X1 U1076 ( .A(n1122), .ZN(n1120) );
  XNOR2_X1 U1077 ( .A(n1123), .B(n1124), .ZN(n1061) );
  NAND2_X1 U1078 ( .A1(n1125), .A2(n1126), .ZN(n1123) );
  NAND2_X1 U1079 ( .A1(a_4_), .A2(n1122), .ZN(n1062) );
  NAND2_X1 U1080 ( .A1(n1070), .A2(n1127), .ZN(n1122) );
  NAND2_X1 U1081 ( .A1(n1069), .A2(n1071), .ZN(n1127) );
  NAND2_X1 U1082 ( .A1(n1074), .A2(n1128), .ZN(n1071) );
  NAND2_X1 U1083 ( .A1(a_5_), .A2(b_3_), .ZN(n1128) );
  INV_X1 U1084 ( .A(n1129), .ZN(n1074) );
  XOR2_X1 U1085 ( .A(n1130), .B(n1131), .Z(n1069) );
  NAND2_X1 U1086 ( .A1(n1129), .A2(a_5_), .ZN(n1070) );
  NOR2_X1 U1087 ( .A1(n1077), .A2(n1076), .ZN(n1129) );
  NAND2_X1 U1088 ( .A1(b_3_), .A2(a_6_), .ZN(n1076) );
  NAND2_X1 U1089 ( .A1(b_2_), .A2(a_7_), .ZN(n1077) );
  OR2_X1 U1090 ( .A1(n1054), .A2(n851), .ZN(n1116) );
  NOR2_X1 U1091 ( .A1(n865), .A2(n819), .ZN(n851) );
  XNOR2_X1 U1092 ( .A(n1132), .B(n1133), .ZN(n1054) );
  NAND2_X1 U1093 ( .A1(n1134), .A2(n1135), .ZN(n1132) );
  OR2_X1 U1094 ( .A1(n1080), .A2(n1081), .ZN(n1105) );
  NOR2_X1 U1095 ( .A1(n657), .A2(n819), .ZN(n1081) );
  XOR2_X1 U1096 ( .A(n1136), .B(n1137), .Z(n1080) );
  XOR2_X1 U1097 ( .A(n1138), .B(n651), .Z(n1136) );
  AND2_X1 U1098 ( .A1(n1139), .A2(n1140), .ZN(n702) );
  NOR2_X1 U1099 ( .A1(n877), .A2(n876), .ZN(n1140) );
  XOR2_X1 U1100 ( .A(n1141), .B(n1142), .Z(n876) );
  NAND2_X1 U1101 ( .A1(n1143), .A2(n1144), .ZN(n1141) );
  NAND2_X1 U1102 ( .A1(n1145), .A2(n1146), .ZN(n1144) );
  NAND2_X1 U1103 ( .A1(a_0_), .A2(b_1_), .ZN(n1145) );
  AND2_X1 U1104 ( .A1(n1095), .A2(n1147), .ZN(n877) );
  NAND2_X1 U1105 ( .A1(n1094), .A2(n1096), .ZN(n1147) );
  NAND2_X1 U1106 ( .A1(n1148), .A2(n1149), .ZN(n1096) );
  NAND2_X1 U1107 ( .A1(a_0_), .A2(b_2_), .ZN(n1149) );
  INV_X1 U1108 ( .A(n1150), .ZN(n1148) );
  XOR2_X1 U1109 ( .A(n1151), .B(n1152), .Z(n1094) );
  XNOR2_X1 U1110 ( .A(n650), .B(n1153), .ZN(n1152) );
  NAND2_X1 U1111 ( .A1(b_0_), .A2(a_2_), .ZN(n1151) );
  NAND2_X1 U1112 ( .A1(a_0_), .A2(n1150), .ZN(n1095) );
  NAND2_X1 U1113 ( .A1(n1154), .A2(n1155), .ZN(n1150) );
  NAND2_X1 U1114 ( .A1(n1104), .A2(n1156), .ZN(n1155) );
  OR2_X1 U1115 ( .A1(n1103), .A2(n1102), .ZN(n1156) );
  NOR2_X1 U1116 ( .A1(n657), .A2(n655), .ZN(n1104) );
  NAND2_X1 U1117 ( .A1(n1102), .A2(n1103), .ZN(n1154) );
  NAND2_X1 U1118 ( .A1(n1157), .A2(n1158), .ZN(n1103) );
  NAND2_X1 U1119 ( .A1(n651), .A2(n1159), .ZN(n1158) );
  OR2_X1 U1120 ( .A1(n1138), .A2(n1137), .ZN(n1159) );
  NOR2_X1 U1121 ( .A1(n656), .A2(n655), .ZN(n651) );
  NAND2_X1 U1122 ( .A1(n1137), .A2(n1138), .ZN(n1157) );
  NAND2_X1 U1123 ( .A1(n1160), .A2(n1161), .ZN(n1138) );
  NAND2_X1 U1124 ( .A1(n1162), .A2(a_3_), .ZN(n1161) );
  NOR2_X1 U1125 ( .A1(n1163), .A2(n655), .ZN(n1162) );
  NOR2_X1 U1126 ( .A1(n1113), .A2(n1114), .ZN(n1163) );
  NAND2_X1 U1127 ( .A1(n1113), .A2(n1114), .ZN(n1160) );
  NAND2_X1 U1128 ( .A1(n1134), .A2(n1164), .ZN(n1114) );
  NAND2_X1 U1129 ( .A1(n1133), .A2(n1135), .ZN(n1164) );
  NAND2_X1 U1130 ( .A1(n1165), .A2(n1166), .ZN(n1135) );
  NAND2_X1 U1131 ( .A1(a_4_), .A2(b_2_), .ZN(n1166) );
  INV_X1 U1132 ( .A(n1167), .ZN(n1165) );
  XNOR2_X1 U1133 ( .A(n1168), .B(n1169), .ZN(n1133) );
  XOR2_X1 U1134 ( .A(n1170), .B(n1171), .Z(n1168) );
  NAND2_X1 U1135 ( .A1(a_4_), .A2(n1167), .ZN(n1134) );
  NAND2_X1 U1136 ( .A1(n1125), .A2(n1172), .ZN(n1167) );
  NAND2_X1 U1137 ( .A1(n1124), .A2(n1126), .ZN(n1172) );
  NAND2_X1 U1138 ( .A1(n1173), .A2(n1174), .ZN(n1126) );
  NAND2_X1 U1139 ( .A1(a_5_), .A2(b_2_), .ZN(n1174) );
  AND2_X1 U1140 ( .A1(n1171), .A2(n1175), .ZN(n1124) );
  NAND2_X1 U1141 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
  OR2_X1 U1142 ( .A1(n1173), .A2(n863), .ZN(n1125) );
  NAND2_X1 U1143 ( .A1(n1130), .A2(n1131), .ZN(n1173) );
  NOR2_X1 U1144 ( .A1(n725), .A2(n655), .ZN(n1131) );
  NOR2_X1 U1145 ( .A1(n614), .A2(n718), .ZN(n1130) );
  XOR2_X1 U1146 ( .A(n1178), .B(n1179), .Z(n1113) );
  NOR2_X1 U1147 ( .A1(n863), .A2(n643), .ZN(n1179) );
  XOR2_X1 U1148 ( .A(n1180), .B(n1181), .Z(n1178) );
  XOR2_X1 U1149 ( .A(n1182), .B(n1183), .Z(n1137) );
  XNOR2_X1 U1150 ( .A(n1184), .B(n1185), .ZN(n1183) );
  NAND2_X1 U1151 ( .A1(b_0_), .A2(a_4_), .ZN(n1182) );
  XNOR2_X1 U1152 ( .A(n1186), .B(n1187), .ZN(n1102) );
  NAND2_X1 U1153 ( .A1(n1188), .A2(n1189), .ZN(n1186) );
  NAND2_X1 U1154 ( .A1(n1190), .A2(n1191), .ZN(n1189) );
  NAND2_X1 U1155 ( .A1(a_2_), .A2(b_1_), .ZN(n1190) );
  NOR2_X1 U1156 ( .A1(n872), .A2(n878), .ZN(n1139) );
  NAND2_X1 U1157 ( .A1(a_0_), .A2(b_0_), .ZN(n878) );
  NAND2_X1 U1158 ( .A1(n1143), .A2(n1192), .ZN(n872) );
  NAND2_X1 U1159 ( .A1(n1193), .A2(n1142), .ZN(n1192) );
  NAND2_X1 U1160 ( .A1(n1194), .A2(n1195), .ZN(n1142) );
  NAND2_X1 U1161 ( .A1(n1196), .A2(b_0_), .ZN(n1195) );
  NOR2_X1 U1162 ( .A1(n1197), .A2(n656), .ZN(n1196) );
  NOR2_X1 U1163 ( .A1(n650), .A2(n1153), .ZN(n1197) );
  NAND2_X1 U1164 ( .A1(n650), .A2(n1153), .ZN(n1194) );
  NAND2_X1 U1165 ( .A1(n1188), .A2(n1198), .ZN(n1153) );
  NAND2_X1 U1166 ( .A1(n1199), .A2(n1187), .ZN(n1198) );
  NAND2_X1 U1167 ( .A1(n1200), .A2(n1201), .ZN(n1187) );
  NAND2_X1 U1168 ( .A1(n1202), .A2(b_0_), .ZN(n1201) );
  NOR2_X1 U1169 ( .A1(n1203), .A2(n864), .ZN(n1202) );
  NOR2_X1 U1170 ( .A1(n1184), .A2(n1185), .ZN(n1203) );
  NAND2_X1 U1171 ( .A1(n1184), .A2(n1185), .ZN(n1200) );
  NAND2_X1 U1172 ( .A1(n1204), .A2(n1205), .ZN(n1185) );
  NAND2_X1 U1173 ( .A1(n1206), .A2(b_0_), .ZN(n1205) );
  NOR2_X1 U1174 ( .A1(n1207), .A2(n863), .ZN(n1206) );
  NOR2_X1 U1175 ( .A1(n1180), .A2(n1181), .ZN(n1207) );
  NAND2_X1 U1176 ( .A1(n1180), .A2(n1181), .ZN(n1204) );
  NAND2_X1 U1177 ( .A1(n1171), .A2(n1208), .ZN(n1181) );
  NAND2_X1 U1178 ( .A1(n1169), .A2(n1170), .ZN(n1208) );
  NOR2_X1 U1179 ( .A1(n614), .A2(n863), .ZN(n1170) );
  NOR2_X1 U1180 ( .A1(n725), .A2(n643), .ZN(n1169) );
  OR2_X1 U1181 ( .A1(n1177), .A2(n1176), .ZN(n1171) );
  NAND2_X1 U1182 ( .A1(b_1_), .A2(a_6_), .ZN(n1176) );
  NAND2_X1 U1183 ( .A1(b_0_), .A2(a_7_), .ZN(n1177) );
  NOR2_X1 U1184 ( .A1(n864), .A2(n614), .ZN(n1180) );
  NOR2_X1 U1185 ( .A1(n865), .A2(n614), .ZN(n1184) );
  NAND2_X1 U1186 ( .A1(n1191), .A2(n656), .ZN(n1199) );
  NAND2_X1 U1187 ( .A1(n1209), .A2(n1210), .ZN(n1188) );
  INV_X1 U1188 ( .A(n1191), .ZN(n1210) );
  NAND2_X1 U1189 ( .A1(b_0_), .A2(a_3_), .ZN(n1191) );
  NOR2_X1 U1190 ( .A1(n614), .A2(n656), .ZN(n1209) );
  NOR2_X1 U1191 ( .A1(n657), .A2(n614), .ZN(n650) );
  NAND2_X1 U1192 ( .A1(n1146), .A2(n894), .ZN(n1193) );
  NAND2_X1 U1193 ( .A1(n1211), .A2(n1212), .ZN(n1143) );
  INV_X1 U1194 ( .A(n1146), .ZN(n1212) );
  NAND2_X1 U1195 ( .A1(b_0_), .A2(a_1_), .ZN(n1146) );
  NOR2_X1 U1196 ( .A1(n614), .A2(n894), .ZN(n1211) );
  AND2_X1 U1197 ( .A1(operation_1_), .A2(operation_0_), .ZN(n592) );
  AND2_X1 U1198 ( .A1(n1213), .A2(n1214), .ZN(n660) );
  NAND2_X1 U1199 ( .A1(n1215), .A2(n608), .ZN(n1214) );
  NOR2_X1 U1200 ( .A1(n1217), .A2(n1218), .ZN(n1215) );
  NOR2_X1 U1201 ( .A1(n639), .A2(n894), .ZN(n1218) );
  INV_X1 U1202 ( .A(n658), .ZN(n639) );
  NOR2_X1 U1203 ( .A1(b_0_), .A2(n1219), .ZN(n1217) );
  NOR2_X1 U1204 ( .A1(a_0_), .A2(n658), .ZN(n1219) );
  NAND2_X1 U1205 ( .A1(n1220), .A2(n1221), .ZN(n658) );
  NAND2_X1 U1206 ( .A1(n1222), .A2(n614), .ZN(n1221) );
  INV_X1 U1207 ( .A(b_1_), .ZN(n614) );
  NAND2_X1 U1208 ( .A1(n609), .A2(n657), .ZN(n1222) );
  INV_X1 U1209 ( .A(n620), .ZN(n609) );
  NAND2_X1 U1210 ( .A1(a_1_), .A2(n620), .ZN(n1220) );
  NAND2_X1 U1211 ( .A1(n1223), .A2(n1224), .ZN(n620) );
  NAND2_X1 U1212 ( .A1(n1225), .A2(n655), .ZN(n1224) );
  INV_X1 U1213 ( .A(b_2_), .ZN(n655) );
  NAND2_X1 U1214 ( .A1(n843), .A2(n656), .ZN(n1225) );
  INV_X1 U1215 ( .A(n866), .ZN(n843) );
  NAND2_X1 U1216 ( .A1(a_2_), .A2(n866), .ZN(n1223) );
  NAND2_X1 U1217 ( .A1(n1226), .A2(n1227), .ZN(n866) );
  NAND2_X1 U1218 ( .A1(n1228), .A2(n819), .ZN(n1227) );
  INV_X1 U1219 ( .A(b_3_), .ZN(n819) );
  NAND2_X1 U1220 ( .A1(n815), .A2(n865), .ZN(n1228) );
  INV_X1 U1221 ( .A(n825), .ZN(n815) );
  NAND2_X1 U1222 ( .A1(a_3_), .A2(n825), .ZN(n1226) );
  NAND2_X1 U1223 ( .A1(n1229), .A2(n1230), .ZN(n825) );
  NAND2_X1 U1224 ( .A1(n1231), .A2(n791), .ZN(n1230) );
  INV_X1 U1225 ( .A(b_4_), .ZN(n791) );
  NAND2_X1 U1226 ( .A1(n787), .A2(n864), .ZN(n1231) );
  INV_X1 U1227 ( .A(n797), .ZN(n787) );
  NAND2_X1 U1228 ( .A1(a_4_), .A2(n797), .ZN(n1229) );
  NAND2_X1 U1229 ( .A1(n1232), .A2(n1233), .ZN(n797) );
  NAND2_X1 U1230 ( .A1(n1234), .A2(n763), .ZN(n1233) );
  INV_X1 U1231 ( .A(b_5_), .ZN(n763) );
  NAND2_X1 U1232 ( .A1(n759), .A2(n863), .ZN(n1234) );
  INV_X1 U1233 ( .A(n769), .ZN(n759) );
  NAND2_X1 U1234 ( .A1(a_5_), .A2(n769), .ZN(n1232) );
  NAND2_X1 U1235 ( .A1(n721), .A2(n1235), .ZN(n769) );
  NAND2_X1 U1236 ( .A1(n709), .A2(n719), .ZN(n1235) );
  NAND2_X1 U1237 ( .A1(b_7_), .A2(n718), .ZN(n709) );
  INV_X1 U1238 ( .A(a_7_), .ZN(n718) );
  NAND2_X1 U1239 ( .A1(n1236), .A2(n742), .ZN(n1213) );
  INV_X1 U1240 ( .A(n610), .ZN(n742) );
  NAND2_X1 U1241 ( .A1(operation_0_), .A2(n1216), .ZN(n610) );
  INV_X1 U1242 ( .A(operation_1_), .ZN(n1216) );
  NOR2_X1 U1243 ( .A1(n1237), .A2(n1238), .ZN(n1236) );
  NOR2_X1 U1244 ( .A1(a_0_), .A2(n659), .ZN(n1238) );
  INV_X1 U1245 ( .A(n640), .ZN(n659) );
  NOR2_X1 U1246 ( .A1(n1239), .A2(n643), .ZN(n1237) );
  INV_X1 U1247 ( .A(b_0_), .ZN(n643) );
  NOR2_X1 U1248 ( .A1(n894), .A2(n640), .ZN(n1239) );
  NAND2_X1 U1249 ( .A1(n1240), .A2(n1241), .ZN(n640) );
  NAND2_X1 U1250 ( .A1(b_1_), .A2(n1242), .ZN(n1241) );
  NAND2_X1 U1251 ( .A1(n621), .A2(a_1_), .ZN(n1242) );
  INV_X1 U1252 ( .A(n611), .ZN(n621) );
  NAND2_X1 U1253 ( .A1(n611), .A2(n657), .ZN(n1240) );
  INV_X1 U1254 ( .A(a_1_), .ZN(n657) );
  NAND2_X1 U1255 ( .A1(n1243), .A2(n1244), .ZN(n611) );
  NAND2_X1 U1256 ( .A1(b_2_), .A2(n1245), .ZN(n1244) );
  NAND2_X1 U1257 ( .A1(n867), .A2(a_2_), .ZN(n1245) );
  INV_X1 U1258 ( .A(n844), .ZN(n867) );
  NAND2_X1 U1259 ( .A1(n844), .A2(n656), .ZN(n1243) );
  INV_X1 U1260 ( .A(a_2_), .ZN(n656) );
  NAND2_X1 U1261 ( .A1(n1246), .A2(n1247), .ZN(n844) );
  NAND2_X1 U1262 ( .A1(b_3_), .A2(n1248), .ZN(n1247) );
  NAND2_X1 U1263 ( .A1(n826), .A2(a_3_), .ZN(n1248) );
  INV_X1 U1264 ( .A(n816), .ZN(n826) );
  NAND2_X1 U1265 ( .A1(n816), .A2(n865), .ZN(n1246) );
  INV_X1 U1266 ( .A(a_3_), .ZN(n865) );
  NAND2_X1 U1267 ( .A1(n1249), .A2(n1250), .ZN(n816) );
  NAND2_X1 U1268 ( .A1(b_4_), .A2(n1251), .ZN(n1250) );
  NAND2_X1 U1269 ( .A1(n798), .A2(a_4_), .ZN(n1251) );
  INV_X1 U1270 ( .A(n788), .ZN(n798) );
  NAND2_X1 U1271 ( .A1(n788), .A2(n864), .ZN(n1249) );
  INV_X1 U1272 ( .A(a_4_), .ZN(n864) );
  NAND2_X1 U1273 ( .A1(n1252), .A2(n1253), .ZN(n788) );
  NAND2_X1 U1274 ( .A1(b_5_), .A2(n1254), .ZN(n1253) );
  NAND2_X1 U1275 ( .A1(n770), .A2(a_5_), .ZN(n1254) );
  INV_X1 U1276 ( .A(n760), .ZN(n770) );
  NAND2_X1 U1277 ( .A1(n760), .A2(n863), .ZN(n1252) );
  INV_X1 U1278 ( .A(a_5_), .ZN(n863) );
  NAND2_X1 U1279 ( .A1(n719), .A2(n1255), .ZN(n760) );
  NAND2_X1 U1280 ( .A1(n710), .A2(n721), .ZN(n1255) );
  NAND2_X1 U1281 ( .A1(a_6_), .A2(n724), .ZN(n721) );
  INV_X1 U1282 ( .A(b_6_), .ZN(n724) );
  NAND2_X1 U1283 ( .A1(a_7_), .A2(n720), .ZN(n710) );
  INV_X1 U1284 ( .A(b_7_), .ZN(n720) );
  NAND2_X1 U1285 ( .A1(b_6_), .A2(n725), .ZN(n719) );
  INV_X1 U1286 ( .A(a_6_), .ZN(n725) );
  INV_X1 U1287 ( .A(a_0_), .ZN(n894) );
endmodule

