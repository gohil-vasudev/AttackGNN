module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n614_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n847_, new_n250_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n636_, new_n670_, new_n456_, new_n170_, new_n246_, new_n682_, new_n812_, new_n679_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n602_, new_n188_, new_n695_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n500_, new_n786_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n742_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n774_, new_n157_, new_n716_, new_n153_, new_n701_, new_n792_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n606_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n167_, new_n385_, new_n829_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n764_, new_n150_, new_n683_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n180_, new_n530_, new_n318_, new_n622_, new_n629_, new_n702_, new_n833_, new_n321_, new_n443_, new_n324_, new_n158_, new_n763_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n816_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n650_, new_n708_, new_n750_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n506_, new_n680_, new_n256_, new_n778_, new_n452_, new_n381_, new_n656_, new_n820_, new_n771_, new_n388_, new_n508_, new_n714_, new_n194_, new_n483_, new_n394_, new_n299_, new_n142_, new_n139_, new_n657_, new_n652_, new_n314_, new_n363_, new_n165_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n790_, new_n187_, new_n311_, new_n465_, new_n739_, new_n783_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n846_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n208_, new_n632_, new_n671_, new_n179_, new_n850_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n805_, new_n559_, new_n762_, new_n838_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n794_, new_n628_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n448_, new_n276_, new_n688_, new_n155_, new_n384_, new_n410_, new_n851_, new_n775_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n809_, new_n654_, new_n713_, new_n227_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n376_, new_n380_, new_n747_, new_n138_, new_n749_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n839_, new_n485_, new_n525_, new_n562_, new_n578_, new_n810_, new_n808_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n800_, new_n379_, new_n719_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n824_, new_n143_, new_n520_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n237_, new_n825_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n748_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n191_, new_n755_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n737_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n662_, new_n440_, new_n733_, new_n531_, new_n593_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n651_, new_n433_, new_n435_, new_n776_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n815_, new_n278_, new_n304_, new_n523_, new_n638_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n711_, new_n644_, new_n731_, new_n836_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n723_, new_n756_, new_n495_, new_n431_, new_n196_, new_n818_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n754_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n803_, new_n330_, new_n375_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n357_, new_n320_, new_n780_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n358_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n802_, new_n697_, new_n185_, new_n709_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n168_, new_n279_, new_n455_, new_n770_, new_n618_, new_n521_, new_n793_, new_n406_, new_n828_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n573_, new_n765_, new_n405_;

not g000 ( new_n138_, N85 );
nand g001 ( new_n139_, new_n138_, N81 );
not g002 ( new_n140_, N81 );
nand g003 ( new_n141_, new_n140_, N85 );
nand g004 ( new_n142_, new_n139_, new_n141_ );
not g005 ( new_n143_, N89 );
not g006 ( new_n144_, N93 );
nand g007 ( new_n145_, new_n143_, new_n144_ );
nand g008 ( new_n146_, N89, N93 );
nand g009 ( new_n147_, new_n145_, new_n146_ );
nand g010 ( new_n148_, new_n142_, new_n147_ );
nand g011 ( new_n149_, new_n145_, new_n139_, new_n141_, new_n146_ );
nand g012 ( new_n150_, new_n148_, new_n149_ );
not g013 ( new_n151_, new_n150_ );
not g014 ( new_n152_, N69 );
nand g015 ( new_n153_, new_n152_, N65 );
not g016 ( new_n154_, N65 );
nand g017 ( new_n155_, new_n154_, N69 );
nand g018 ( new_n156_, new_n153_, new_n155_ );
not g019 ( new_n157_, N73 );
not g020 ( new_n158_, N77 );
nand g021 ( new_n159_, new_n157_, new_n158_ );
nand g022 ( new_n160_, N73, N77 );
nand g023 ( new_n161_, new_n159_, new_n160_ );
nand g024 ( new_n162_, new_n156_, new_n161_ );
nand g025 ( new_n163_, new_n159_, new_n153_, new_n155_, new_n160_ );
nand g026 ( new_n164_, new_n162_, new_n163_ );
nand g027 ( new_n165_, new_n151_, new_n164_ );
not g028 ( new_n166_, new_n164_ );
nand g029 ( new_n167_, new_n166_, new_n150_ );
nand g030 ( new_n168_, new_n165_, new_n167_ );
nand g031 ( new_n169_, N129, N137 );
nand g032 ( new_n170_, new_n168_, new_n169_ );
nand g033 ( new_n171_, new_n165_, new_n167_, N129, N137 );
nand g034 ( new_n172_, new_n170_, new_n171_ );
not g035 ( new_n173_, N1 );
not g036 ( new_n174_, N17 );
nand g037 ( new_n175_, new_n173_, new_n174_ );
nand g038 ( new_n176_, N1, N17 );
nand g039 ( new_n177_, new_n175_, new_n176_ );
not g040 ( new_n178_, N33 );
not g041 ( new_n179_, N49 );
nand g042 ( new_n180_, new_n178_, new_n179_ );
nand g043 ( new_n181_, N33, N49 );
nand g044 ( new_n182_, new_n180_, new_n181_ );
nand g045 ( new_n183_, new_n177_, new_n182_ );
nand g046 ( new_n184_, new_n175_, new_n180_, new_n176_, new_n181_ );
nand g047 ( new_n185_, new_n183_, new_n184_ );
nand g048 ( new_n186_, new_n172_, new_n185_ );
nand g049 ( new_n187_, new_n170_, new_n171_, new_n183_, new_n184_ );
nand g050 ( new_n188_, new_n186_, new_n187_ );
not g051 ( new_n189_, new_n188_ );
not g052 ( new_n190_, keyIn_0_22 );
not g053 ( new_n191_, keyIn_0_20 );
not g054 ( new_n192_, keyIn_0_18 );
not g055 ( new_n193_, keyIn_0_0 );
not g056 ( new_n194_, N5 );
nand g057 ( new_n195_, new_n173_, new_n194_ );
nand g058 ( new_n196_, N1, N5 );
nand g059 ( new_n197_, new_n195_, new_n196_ );
nand g060 ( new_n198_, new_n197_, new_n193_ );
nand g061 ( new_n199_, new_n195_, keyIn_0_0, new_n196_ );
nand g062 ( new_n200_, new_n198_, new_n199_ );
not g063 ( new_n201_, N9 );
not g064 ( new_n202_, N13 );
nand g065 ( new_n203_, new_n201_, new_n202_ );
nand g066 ( new_n204_, N9, N13 );
nand g067 ( new_n205_, new_n203_, new_n204_ );
nand g068 ( new_n206_, new_n205_, keyIn_0_1 );
not g069 ( new_n207_, keyIn_0_1 );
nand g070 ( new_n208_, new_n203_, new_n207_, new_n204_ );
nand g071 ( new_n209_, new_n206_, new_n208_ );
nand g072 ( new_n210_, new_n200_, new_n209_ );
nand g073 ( new_n211_, new_n198_, new_n206_, new_n199_, new_n208_ );
nand g074 ( new_n212_, new_n210_, new_n211_ );
nand g075 ( new_n213_, new_n212_, keyIn_0_12 );
not g076 ( new_n214_, keyIn_0_12 );
nand g077 ( new_n215_, new_n210_, new_n214_, new_n211_ );
nand g078 ( new_n216_, new_n213_, new_n215_ );
not g079 ( new_n217_, keyIn_0_13 );
not g080 ( new_n218_, N25 );
not g081 ( new_n219_, N29 );
nand g082 ( new_n220_, new_n218_, new_n219_ );
nand g083 ( new_n221_, N25, N29 );
nand g084 ( new_n222_, new_n220_, new_n221_ );
nand g085 ( new_n223_, new_n222_, keyIn_0_3 );
not g086 ( new_n224_, keyIn_0_3 );
nand g087 ( new_n225_, new_n220_, new_n224_, new_n221_ );
nand g088 ( new_n226_, new_n223_, new_n225_ );
not g089 ( new_n227_, keyIn_0_2 );
not g090 ( new_n228_, N21 );
nand g091 ( new_n229_, new_n174_, new_n228_ );
nand g092 ( new_n230_, N17, N21 );
nand g093 ( new_n231_, new_n229_, new_n230_ );
nand g094 ( new_n232_, new_n231_, new_n227_ );
nand g095 ( new_n233_, new_n229_, keyIn_0_2, new_n230_ );
nand g096 ( new_n234_, new_n232_, new_n233_ );
nand g097 ( new_n235_, new_n226_, new_n234_ );
nand g098 ( new_n236_, new_n223_, new_n232_, new_n225_, new_n233_ );
nand g099 ( new_n237_, new_n235_, new_n236_ );
nand g100 ( new_n238_, new_n237_, new_n217_ );
nand g101 ( new_n239_, new_n235_, keyIn_0_13, new_n236_ );
nand g102 ( new_n240_, new_n238_, new_n239_ );
nand g103 ( new_n241_, new_n216_, new_n240_ );
nand g104 ( new_n242_, new_n213_, new_n238_, new_n215_, new_n239_ );
nand g105 ( new_n243_, new_n241_, new_n242_ );
nand g106 ( new_n244_, new_n243_, new_n192_ );
nand g107 ( new_n245_, new_n241_, keyIn_0_18, new_n242_ );
nand g108 ( new_n246_, new_n244_, new_n245_ );
nand g109 ( new_n247_, N133, N137 );
nand g110 ( new_n248_, new_n247_, keyIn_0_6 );
not g111 ( new_n249_, keyIn_0_6 );
nand g112 ( new_n250_, new_n249_, N133, N137 );
nand g113 ( new_n251_, new_n248_, new_n250_ );
nand g114 ( new_n252_, new_n246_, new_n251_ );
nand g115 ( new_n253_, new_n244_, new_n245_, new_n248_, new_n250_ );
nand g116 ( new_n254_, new_n252_, new_n253_ );
nand g117 ( new_n255_, new_n254_, new_n191_ );
nand g118 ( new_n256_, new_n252_, keyIn_0_20, new_n253_ );
nand g119 ( new_n257_, new_n255_, new_n256_ );
not g120 ( new_n258_, keyIn_0_16 );
nor g121 ( new_n259_, N97, N113 );
not g122 ( new_n260_, new_n259_ );
nand g123 ( new_n261_, N97, N113 );
nand g124 ( new_n262_, new_n260_, new_n261_ );
nand g125 ( new_n263_, new_n262_, keyIn_0_9 );
not g126 ( new_n264_, new_n263_ );
nor g127 ( new_n265_, new_n262_, keyIn_0_9 );
nor g128 ( new_n266_, new_n264_, new_n265_ );
not g129 ( new_n267_, new_n266_ );
nand g130 ( new_n268_, new_n140_, N65 );
nand g131 ( new_n269_, new_n154_, N81 );
nand g132 ( new_n270_, new_n268_, new_n269_ );
nand g133 ( new_n271_, new_n270_, keyIn_0_8 );
not g134 ( new_n272_, keyIn_0_8 );
nand g135 ( new_n273_, new_n268_, new_n269_, new_n272_ );
nand g136 ( new_n274_, new_n271_, new_n273_ );
nand g137 ( new_n275_, new_n267_, new_n274_ );
nand g138 ( new_n276_, new_n266_, new_n271_, new_n273_ );
nand g139 ( new_n277_, new_n275_, new_n276_ );
nand g140 ( new_n278_, new_n277_, new_n258_ );
nand g141 ( new_n279_, new_n275_, keyIn_0_16, new_n276_ );
nand g142 ( new_n280_, new_n278_, new_n279_ );
not g143 ( new_n281_, new_n280_ );
nand g144 ( new_n282_, new_n257_, new_n281_ );
nand g145 ( new_n283_, new_n255_, new_n256_, new_n280_ );
nand g146 ( new_n284_, new_n282_, new_n283_ );
nand g147 ( new_n285_, new_n284_, new_n190_ );
nand g148 ( new_n286_, new_n282_, keyIn_0_22, new_n283_ );
nand g149 ( new_n287_, new_n285_, new_n286_ );
not g150 ( new_n288_, new_n287_ );
not g151 ( new_n289_, keyIn_0_4 );
not g152 ( new_n290_, N37 );
nand g153 ( new_n291_, new_n178_, new_n290_ );
nand g154 ( new_n292_, N33, N37 );
nand g155 ( new_n293_, new_n291_, new_n292_ );
nand g156 ( new_n294_, new_n293_, new_n289_ );
nand g157 ( new_n295_, new_n291_, keyIn_0_4, new_n292_ );
nand g158 ( new_n296_, new_n294_, new_n295_ );
not g159 ( new_n297_, N41 );
not g160 ( new_n298_, N45 );
nand g161 ( new_n299_, new_n297_, new_n298_ );
nand g162 ( new_n300_, N41, N45 );
nand g163 ( new_n301_, new_n299_, new_n300_ );
nand g164 ( new_n302_, new_n301_, keyIn_0_5 );
not g165 ( new_n303_, keyIn_0_5 );
nand g166 ( new_n304_, new_n299_, new_n303_, new_n300_ );
nand g167 ( new_n305_, new_n302_, new_n304_ );
nand g168 ( new_n306_, new_n296_, new_n305_ );
nand g169 ( new_n307_, new_n294_, new_n302_, new_n295_, new_n304_ );
nand g170 ( new_n308_, new_n306_, new_n307_ );
nand g171 ( new_n309_, new_n308_, keyIn_0_14 );
not g172 ( new_n310_, keyIn_0_14 );
nand g173 ( new_n311_, new_n306_, new_n310_, new_n307_ );
nand g174 ( new_n312_, new_n309_, new_n311_ );
not g175 ( new_n313_, N53 );
nand g176 ( new_n314_, new_n313_, N49 );
nand g177 ( new_n315_, new_n179_, N53 );
nand g178 ( new_n316_, new_n314_, new_n315_ );
not g179 ( new_n317_, N57 );
not g180 ( new_n318_, N61 );
nand g181 ( new_n319_, new_n317_, new_n318_ );
nand g182 ( new_n320_, N57, N61 );
nand g183 ( new_n321_, new_n319_, new_n320_ );
nand g184 ( new_n322_, new_n316_, new_n321_ );
nand g185 ( new_n323_, new_n319_, new_n314_, new_n315_, new_n320_ );
nand g186 ( new_n324_, new_n322_, new_n323_ );
not g187 ( new_n325_, new_n324_ );
nand g188 ( new_n326_, new_n312_, new_n325_ );
nand g189 ( new_n327_, new_n309_, new_n311_, new_n324_ );
nand g190 ( new_n328_, new_n326_, new_n327_ );
nand g191 ( new_n329_, N134, N137 );
nand g192 ( new_n330_, new_n328_, new_n329_ );
nand g193 ( new_n331_, new_n326_, N134, N137, new_n327_ );
nand g194 ( new_n332_, new_n330_, new_n331_ );
nand g195 ( new_n333_, new_n152_, new_n138_ );
nand g196 ( new_n334_, N69, N85 );
nand g197 ( new_n335_, new_n333_, new_n334_ );
not g198 ( new_n336_, N101 );
not g199 ( new_n337_, N117 );
nand g200 ( new_n338_, new_n336_, new_n337_ );
nand g201 ( new_n339_, N101, N117 );
nand g202 ( new_n340_, new_n338_, new_n339_ );
nand g203 ( new_n341_, new_n335_, new_n340_ );
nand g204 ( new_n342_, new_n333_, new_n338_, new_n334_, new_n339_ );
nand g205 ( new_n343_, new_n341_, new_n342_ );
nand g206 ( new_n344_, new_n332_, new_n343_ );
nand g207 ( new_n345_, new_n330_, new_n331_, new_n341_, new_n342_ );
nand g208 ( new_n346_, new_n344_, new_n345_ );
not g209 ( new_n347_, new_n346_ );
nand g210 ( new_n348_, new_n288_, new_n347_ );
not g211 ( new_n349_, keyIn_0_23 );
not g212 ( new_n350_, keyIn_0_21 );
nand g213 ( new_n351_, new_n216_, new_n312_ );
nand g214 ( new_n352_, new_n213_, new_n309_, new_n215_, new_n311_ );
nand g215 ( new_n353_, new_n351_, new_n352_ );
nand g216 ( new_n354_, new_n353_, keyIn_0_19 );
not g217 ( new_n355_, keyIn_0_19 );
nand g218 ( new_n356_, new_n351_, new_n355_, new_n352_ );
nand g219 ( new_n357_, new_n354_, new_n356_ );
nand g220 ( new_n358_, N135, N137 );
nand g221 ( new_n359_, new_n358_, keyIn_0_7 );
not g222 ( new_n360_, keyIn_0_7 );
nand g223 ( new_n361_, new_n360_, N135, N137 );
nand g224 ( new_n362_, new_n359_, new_n361_ );
not g225 ( new_n363_, new_n362_ );
nand g226 ( new_n364_, new_n357_, new_n363_ );
nand g227 ( new_n365_, new_n354_, new_n356_, new_n362_ );
nand g228 ( new_n366_, new_n364_, new_n365_ );
nand g229 ( new_n367_, new_n366_, new_n350_ );
nand g230 ( new_n368_, new_n364_, keyIn_0_21, new_n365_ );
nand g231 ( new_n369_, new_n367_, new_n368_ );
nand g232 ( new_n370_, new_n143_, N73 );
nand g233 ( new_n371_, new_n157_, N89 );
nand g234 ( new_n372_, new_n370_, new_n371_ );
nand g235 ( new_n373_, new_n372_, keyIn_0_10 );
not g236 ( new_n374_, keyIn_0_10 );
nand g237 ( new_n375_, new_n370_, new_n371_, new_n374_ );
nand g238 ( new_n376_, new_n373_, new_n375_ );
not g239 ( new_n377_, N121 );
nand g240 ( new_n378_, new_n377_, N105 );
not g241 ( new_n379_, N105 );
nand g242 ( new_n380_, new_n379_, N121 );
nand g243 ( new_n381_, new_n378_, new_n380_ );
nand g244 ( new_n382_, new_n381_, keyIn_0_11 );
not g245 ( new_n383_, keyIn_0_11 );
nand g246 ( new_n384_, new_n378_, new_n380_, new_n383_ );
nand g247 ( new_n385_, new_n382_, new_n384_ );
nand g248 ( new_n386_, new_n376_, new_n385_ );
nand g249 ( new_n387_, new_n373_, new_n382_, new_n375_, new_n384_ );
nand g250 ( new_n388_, new_n386_, new_n387_ );
nand g251 ( new_n389_, new_n388_, keyIn_0_17 );
not g252 ( new_n390_, keyIn_0_17 );
nand g253 ( new_n391_, new_n386_, new_n390_, new_n387_ );
nand g254 ( new_n392_, new_n389_, new_n391_ );
not g255 ( new_n393_, new_n392_ );
nand g256 ( new_n394_, new_n369_, new_n393_ );
nand g257 ( new_n395_, new_n367_, new_n368_, new_n392_ );
nand g258 ( new_n396_, new_n394_, new_n395_ );
nand g259 ( new_n397_, new_n396_, new_n349_ );
nand g260 ( new_n398_, new_n394_, keyIn_0_23, new_n395_ );
nand g261 ( new_n399_, new_n397_, new_n398_ );
nand g262 ( new_n400_, new_n336_, N97 );
not g263 ( new_n401_, N97 );
nand g264 ( new_n402_, new_n401_, N101 );
nand g265 ( new_n403_, new_n400_, new_n402_ );
not g266 ( new_n404_, N109 );
nand g267 ( new_n405_, new_n379_, new_n404_ );
nand g268 ( new_n406_, N105, N109 );
nand g269 ( new_n407_, new_n405_, new_n406_ );
nand g270 ( new_n408_, new_n403_, new_n407_ );
nand g271 ( new_n409_, new_n405_, new_n400_, new_n402_, new_n406_ );
nand g272 ( new_n410_, new_n408_, new_n409_ );
not g273 ( new_n411_, new_n410_ );
nand g274 ( new_n412_, new_n411_, new_n164_ );
nand g275 ( new_n413_, new_n166_, new_n410_ );
nand g276 ( new_n414_, new_n412_, new_n413_ );
nand g277 ( new_n415_, N131, N137 );
nand g278 ( new_n416_, new_n414_, new_n415_ );
nand g279 ( new_n417_, new_n412_, new_n413_, N131, N137 );
nand g280 ( new_n418_, new_n416_, new_n417_ );
nand g281 ( new_n419_, new_n201_, new_n218_ );
nand g282 ( new_n420_, N9, N25 );
nand g283 ( new_n421_, new_n419_, new_n420_ );
nand g284 ( new_n422_, new_n297_, new_n317_ );
nand g285 ( new_n423_, N41, N57 );
nand g286 ( new_n424_, new_n422_, new_n423_ );
nand g287 ( new_n425_, new_n421_, new_n424_ );
nand g288 ( new_n426_, new_n419_, new_n422_, new_n420_, new_n423_ );
nand g289 ( new_n427_, new_n425_, new_n426_ );
nand g290 ( new_n428_, new_n418_, new_n427_ );
nand g291 ( new_n429_, new_n416_, new_n417_, new_n425_, new_n426_ );
nand g292 ( new_n430_, new_n428_, new_n429_ );
not g293 ( new_n431_, new_n430_ );
nand g294 ( new_n432_, new_n189_, new_n431_ );
not g295 ( new_n433_, new_n432_ );
nand g296 ( new_n434_, new_n337_, N113 );
not g297 ( new_n435_, N113 );
nand g298 ( new_n436_, new_n435_, N117 );
nand g299 ( new_n437_, new_n434_, new_n436_ );
not g300 ( new_n438_, N125 );
nand g301 ( new_n439_, new_n377_, new_n438_ );
nand g302 ( new_n440_, N121, N125 );
nand g303 ( new_n441_, new_n439_, new_n440_ );
nand g304 ( new_n442_, new_n437_, new_n441_ );
nand g305 ( new_n443_, new_n439_, new_n434_, new_n436_, new_n440_ );
nand g306 ( new_n444_, new_n442_, new_n443_ );
nand g307 ( new_n445_, new_n411_, new_n444_ );
not g308 ( new_n446_, new_n444_ );
nand g309 ( new_n447_, new_n446_, new_n410_ );
nand g310 ( new_n448_, new_n445_, new_n447_ );
nand g311 ( new_n449_, N130, N137 );
nand g312 ( new_n450_, new_n448_, new_n449_ );
nand g313 ( new_n451_, new_n445_, new_n447_, N130, N137 );
nand g314 ( new_n452_, new_n450_, new_n451_ );
nand g315 ( new_n453_, new_n194_, new_n228_ );
nand g316 ( new_n454_, N5, N21 );
nand g317 ( new_n455_, new_n453_, new_n454_ );
nand g318 ( new_n456_, new_n290_, new_n313_ );
nand g319 ( new_n457_, N37, N53 );
nand g320 ( new_n458_, new_n456_, new_n457_ );
nand g321 ( new_n459_, new_n455_, new_n458_ );
nand g322 ( new_n460_, new_n453_, new_n456_, new_n454_, new_n457_ );
nand g323 ( new_n461_, new_n459_, new_n460_ );
nand g324 ( new_n462_, new_n452_, new_n461_ );
nand g325 ( new_n463_, new_n450_, new_n451_, new_n459_, new_n460_ );
nand g326 ( new_n464_, new_n462_, new_n463_ );
nand g327 ( new_n465_, new_n433_, new_n464_ );
not g328 ( new_n466_, new_n464_ );
nand g329 ( new_n467_, new_n188_, new_n430_, keyIn_0_24 );
nand g330 ( new_n468_, new_n430_, keyIn_0_24 );
nand g331 ( new_n469_, new_n468_, new_n189_ );
nand g332 ( new_n470_, new_n469_, new_n466_, new_n467_ );
nand g333 ( new_n471_, new_n465_, new_n470_ );
nand g334 ( new_n472_, new_n446_, new_n150_ );
nand g335 ( new_n473_, new_n151_, new_n444_ );
nand g336 ( new_n474_, new_n472_, new_n473_ );
nand g337 ( new_n475_, N132, N137 );
nand g338 ( new_n476_, new_n474_, new_n475_ );
nand g339 ( new_n477_, new_n472_, new_n473_, N132, N137 );
nand g340 ( new_n478_, new_n476_, new_n477_ );
not g341 ( new_n479_, keyIn_0_15 );
nand g342 ( new_n480_, new_n219_, N13 );
nand g343 ( new_n481_, new_n202_, N29 );
nand g344 ( new_n482_, new_n480_, new_n481_ );
nand g345 ( new_n483_, new_n298_, new_n318_ );
nand g346 ( new_n484_, N45, N61 );
nand g347 ( new_n485_, new_n483_, new_n484_ );
nand g348 ( new_n486_, new_n482_, new_n485_ );
nand g349 ( new_n487_, new_n483_, new_n480_, new_n481_, new_n484_ );
nand g350 ( new_n488_, new_n486_, new_n487_ );
nand g351 ( new_n489_, new_n488_, new_n479_ );
nand g352 ( new_n490_, new_n486_, keyIn_0_15, new_n487_ );
nand g353 ( new_n491_, new_n489_, new_n490_ );
nand g354 ( new_n492_, new_n478_, new_n491_ );
nand g355 ( new_n493_, new_n476_, new_n477_, new_n489_, new_n490_ );
nand g356 ( new_n494_, new_n492_, new_n493_ );
not g357 ( new_n495_, new_n494_ );
nand g358 ( new_n496_, new_n471_, new_n495_ );
nand g359 ( new_n497_, new_n433_, new_n466_, new_n494_ );
nand g360 ( new_n498_, new_n496_, new_n497_ );
nand g361 ( new_n499_, new_n240_, new_n325_ );
nand g362 ( new_n500_, new_n238_, new_n239_, new_n324_ );
nand g363 ( new_n501_, new_n499_, new_n500_ );
nand g364 ( new_n502_, N136, N137 );
nand g365 ( new_n503_, new_n501_, new_n502_ );
nand g366 ( new_n504_, new_n499_, N136, N137, new_n500_ );
nand g367 ( new_n505_, new_n503_, new_n504_ );
nand g368 ( new_n506_, new_n158_, new_n144_ );
nand g369 ( new_n507_, N77, N93 );
nand g370 ( new_n508_, new_n506_, new_n507_ );
nand g371 ( new_n509_, new_n404_, new_n438_ );
nand g372 ( new_n510_, N109, N125 );
nand g373 ( new_n511_, new_n509_, new_n510_ );
nand g374 ( new_n512_, new_n508_, new_n511_ );
nand g375 ( new_n513_, new_n506_, new_n509_, new_n507_, new_n510_ );
nand g376 ( new_n514_, new_n512_, new_n513_ );
nand g377 ( new_n515_, new_n505_, new_n514_ );
nand g378 ( new_n516_, new_n503_, new_n504_, new_n512_, new_n513_ );
nand g379 ( new_n517_, new_n515_, new_n516_ );
not g380 ( new_n518_, new_n517_ );
nand g381 ( new_n519_, new_n498_, new_n518_ );
not g382 ( new_n520_, new_n519_ );
nand g383 ( new_n521_, new_n399_, new_n520_ );
nor g384 ( new_n522_, new_n348_, new_n521_ );
not g385 ( new_n523_, new_n522_ );
nor g386 ( new_n524_, new_n523_, new_n189_ );
not g387 ( new_n525_, new_n524_ );
nand g388 ( new_n526_, new_n525_, N1 );
nand g389 ( new_n527_, new_n524_, new_n173_ );
nand g390 ( N724, new_n526_, new_n527_ );
nor g391 ( new_n529_, new_n523_, new_n466_ );
not g392 ( new_n530_, new_n529_ );
nand g393 ( new_n531_, new_n530_, N5 );
nand g394 ( new_n532_, new_n529_, new_n194_ );
nand g395 ( N725, new_n531_, new_n532_ );
nor g396 ( new_n534_, new_n523_, new_n431_ );
not g397 ( new_n535_, new_n534_ );
nand g398 ( new_n536_, new_n535_, N9 );
nand g399 ( new_n537_, new_n534_, new_n201_ );
nand g400 ( N726, new_n536_, new_n537_ );
nor g401 ( new_n539_, new_n523_, new_n495_ );
not g402 ( new_n540_, new_n539_ );
nand g403 ( new_n541_, new_n540_, N13 );
nand g404 ( new_n542_, new_n539_, new_n202_ );
nand g405 ( N727, new_n541_, new_n542_ );
nand g406 ( new_n544_, new_n397_, new_n398_, new_n498_, new_n517_ );
nor g407 ( new_n545_, new_n348_, new_n544_ );
not g408 ( new_n546_, new_n545_ );
nor g409 ( new_n547_, new_n546_, new_n189_ );
not g410 ( new_n548_, new_n547_ );
nand g411 ( new_n549_, new_n548_, N17 );
nand g412 ( new_n550_, new_n547_, new_n174_ );
nand g413 ( N728, new_n549_, new_n550_ );
nor g414 ( new_n552_, new_n546_, new_n466_ );
not g415 ( new_n553_, new_n552_ );
nand g416 ( new_n554_, new_n553_, N21 );
nand g417 ( new_n555_, new_n552_, new_n228_ );
nand g418 ( N729, new_n554_, new_n555_ );
nor g419 ( new_n557_, new_n546_, new_n431_ );
not g420 ( new_n558_, new_n557_ );
nand g421 ( new_n559_, new_n558_, N25 );
nand g422 ( new_n560_, new_n557_, new_n218_ );
nand g423 ( N730, new_n559_, new_n560_ );
nor g424 ( new_n562_, new_n546_, new_n495_ );
not g425 ( new_n563_, new_n562_ );
nand g426 ( new_n564_, new_n563_, N29 );
nand g427 ( new_n565_, new_n562_, new_n219_ );
nand g428 ( N731, new_n564_, new_n565_ );
nand g429 ( new_n567_, new_n287_, new_n399_, new_n346_, new_n520_ );
nor g430 ( new_n568_, new_n567_, new_n189_ );
not g431 ( new_n569_, new_n568_ );
nand g432 ( new_n570_, new_n569_, N33 );
nand g433 ( new_n571_, new_n568_, new_n178_ );
nand g434 ( N732, new_n570_, new_n571_ );
nor g435 ( new_n573_, new_n567_, new_n466_ );
not g436 ( new_n574_, new_n573_ );
nand g437 ( new_n575_, new_n574_, N37 );
nand g438 ( new_n576_, new_n573_, new_n290_ );
nand g439 ( N733, new_n575_, new_n576_ );
nor g440 ( new_n578_, new_n567_, new_n431_ );
not g441 ( new_n579_, new_n578_ );
nand g442 ( new_n580_, new_n579_, N41 );
nand g443 ( new_n581_, new_n578_, new_n297_ );
nand g444 ( N734, new_n580_, new_n581_ );
nor g445 ( new_n583_, new_n567_, new_n495_ );
not g446 ( new_n584_, new_n583_ );
nand g447 ( new_n585_, new_n584_, N45 );
nand g448 ( new_n586_, new_n583_, new_n298_ );
nand g449 ( N735, new_n585_, new_n586_ );
nor g450 ( new_n588_, new_n288_, new_n544_, new_n347_ );
not g451 ( new_n589_, new_n588_ );
nor g452 ( new_n590_, new_n589_, new_n189_ );
not g453 ( new_n591_, new_n590_ );
nand g454 ( new_n592_, new_n591_, N49 );
nand g455 ( new_n593_, new_n590_, new_n179_ );
nand g456 ( N736, new_n592_, new_n593_ );
nor g457 ( new_n595_, new_n589_, new_n466_ );
not g458 ( new_n596_, new_n595_ );
nand g459 ( new_n597_, new_n596_, N53 );
nand g460 ( new_n598_, new_n595_, new_n313_ );
nand g461 ( N737, new_n597_, new_n598_ );
nor g462 ( new_n600_, new_n589_, new_n431_ );
not g463 ( new_n601_, new_n600_ );
nand g464 ( new_n602_, new_n601_, N57 );
nand g465 ( new_n603_, new_n600_, new_n317_ );
nand g466 ( N738, new_n602_, new_n603_ );
nor g467 ( new_n605_, new_n589_, new_n495_ );
not g468 ( new_n606_, new_n605_ );
nand g469 ( new_n607_, new_n606_, N61 );
nand g470 ( new_n608_, new_n605_, new_n318_ );
nand g471 ( N739, new_n607_, new_n608_ );
not g472 ( new_n610_, keyIn_0_52 );
not g473 ( new_n611_, keyIn_0_32 );
nand g474 ( new_n612_, new_n399_, keyIn_0_27 );
not g475 ( new_n613_, keyIn_0_27 );
nand g476 ( new_n614_, new_n397_, new_n613_, new_n398_ );
nand g477 ( new_n615_, new_n612_, new_n614_ );
not g478 ( new_n616_, keyIn_0_25 );
nand g479 ( new_n617_, new_n288_, new_n616_ );
nand g480 ( new_n618_, new_n287_, keyIn_0_25 );
not g481 ( new_n619_, keyIn_0_26 );
nand g482 ( new_n620_, new_n347_, new_n619_ );
nand g483 ( new_n621_, new_n346_, keyIn_0_26 );
nand g484 ( new_n622_, new_n620_, new_n517_, new_n621_ );
not g485 ( new_n623_, new_n622_ );
nand g486 ( new_n624_, new_n615_, new_n617_, new_n618_, new_n623_ );
nand g487 ( new_n625_, new_n624_, new_n611_ );
nand g488 ( new_n626_, new_n618_, new_n623_ );
not g489 ( new_n627_, new_n626_ );
nand g490 ( new_n628_, new_n627_, keyIn_0_32, new_n615_, new_n617_ );
nand g491 ( new_n629_, new_n625_, new_n628_ );
not g492 ( new_n630_, new_n629_ );
nand g493 ( new_n631_, new_n399_, keyIn_0_30 );
nor g494 ( new_n632_, new_n347_, new_n517_ );
nand g495 ( new_n633_, new_n631_, new_n632_ );
not g496 ( new_n634_, keyIn_0_29 );
nand g497 ( new_n635_, new_n287_, new_n634_ );
not g498 ( new_n636_, keyIn_0_30 );
nand g499 ( new_n637_, new_n397_, new_n636_, new_n398_ );
nand g500 ( new_n638_, new_n285_, keyIn_0_29, new_n286_ );
nand g501 ( new_n639_, new_n635_, new_n637_, new_n638_ );
nor g502 ( new_n640_, new_n639_, new_n633_ );
nor g503 ( new_n641_, new_n640_, keyIn_0_34 );
not g504 ( new_n642_, keyIn_0_34 );
nor g505 ( new_n643_, new_n639_, new_n633_, new_n642_ );
nor g506 ( new_n644_, new_n641_, new_n643_ );
not g507 ( new_n645_, keyIn_0_31 );
nand g508 ( new_n646_, new_n399_, new_n645_ );
nand g509 ( new_n647_, new_n397_, keyIn_0_31, new_n398_ );
nand g510 ( new_n648_, new_n646_, new_n647_ );
nand g511 ( new_n649_, new_n285_, new_n286_, new_n347_, new_n518_ );
not g512 ( new_n650_, new_n649_ );
nand g513 ( new_n651_, new_n648_, new_n650_ );
nand g514 ( new_n652_, new_n651_, keyIn_0_35 );
not g515 ( new_n653_, keyIn_0_35 );
nand g516 ( new_n654_, new_n648_, new_n653_, new_n650_ );
nand g517 ( new_n655_, new_n652_, new_n654_ );
not g518 ( new_n656_, keyIn_0_33 );
nand g519 ( new_n657_, new_n288_, keyIn_0_28 );
not g520 ( new_n658_, keyIn_0_28 );
nand g521 ( new_n659_, new_n287_, new_n658_ );
nand g522 ( new_n660_, new_n399_, new_n347_, new_n518_ );
not g523 ( new_n661_, new_n660_ );
nand g524 ( new_n662_, new_n661_, new_n657_, new_n659_ );
nand g525 ( new_n663_, new_n662_, new_n656_ );
nand g526 ( new_n664_, new_n661_, new_n657_, keyIn_0_33, new_n659_ );
nand g527 ( new_n665_, new_n663_, new_n664_ );
nand g528 ( new_n666_, new_n630_, new_n644_, new_n655_, new_n665_ );
nand g529 ( new_n667_, new_n666_, keyIn_0_36 );
not g530 ( new_n668_, keyIn_0_36 );
nand g531 ( new_n669_, new_n665_, new_n655_ );
not g532 ( new_n670_, new_n669_ );
nand g533 ( new_n671_, new_n670_, new_n668_, new_n630_, new_n644_ );
nand g534 ( new_n672_, new_n667_, new_n671_ );
nand g535 ( new_n673_, new_n495_, new_n430_ );
nand g536 ( new_n674_, new_n466_, new_n188_ );
nor g537 ( new_n675_, new_n673_, new_n674_ );
nand g538 ( new_n676_, new_n672_, new_n675_ );
nand g539 ( new_n677_, new_n676_, keyIn_0_37 );
not g540 ( new_n678_, keyIn_0_37 );
nand g541 ( new_n679_, new_n672_, new_n678_, new_n675_ );
nand g542 ( new_n680_, new_n677_, new_n679_ );
nand g543 ( new_n681_, new_n680_, new_n288_ );
nand g544 ( new_n682_, new_n681_, keyIn_0_40 );
not g545 ( new_n683_, keyIn_0_40 );
nand g546 ( new_n684_, new_n680_, new_n683_, new_n288_ );
nand g547 ( new_n685_, new_n682_, new_n684_ );
nand g548 ( new_n686_, new_n685_, N65 );
nand g549 ( new_n687_, new_n682_, new_n154_, new_n684_ );
nand g550 ( new_n688_, new_n686_, new_n687_ );
nand g551 ( new_n689_, new_n688_, new_n610_ );
nand g552 ( new_n690_, new_n686_, keyIn_0_52, new_n687_ );
nand g553 ( N740, new_n689_, new_n690_ );
not g554 ( new_n692_, keyIn_0_53 );
not g555 ( new_n693_, keyIn_0_41 );
nand g556 ( new_n694_, new_n680_, new_n346_ );
nand g557 ( new_n695_, new_n694_, new_n693_ );
nand g558 ( new_n696_, new_n680_, keyIn_0_41, new_n346_ );
nand g559 ( new_n697_, new_n695_, new_n696_ );
nand g560 ( new_n698_, new_n697_, new_n152_ );
nand g561 ( new_n699_, new_n695_, N69, new_n696_ );
nand g562 ( new_n700_, new_n698_, new_n699_ );
nand g563 ( new_n701_, new_n700_, new_n692_ );
nand g564 ( new_n702_, new_n698_, keyIn_0_53, new_n699_ );
nand g565 ( N741, new_n701_, new_n702_ );
nand g566 ( new_n704_, new_n680_, new_n399_ );
nand g567 ( new_n705_, new_n704_, keyIn_0_42 );
not g568 ( new_n706_, keyIn_0_42 );
nand g569 ( new_n707_, new_n680_, new_n706_, new_n399_ );
nand g570 ( new_n708_, new_n705_, new_n707_ );
nand g571 ( new_n709_, new_n708_, new_n157_ );
nand g572 ( new_n710_, new_n705_, N73, new_n707_ );
nand g573 ( new_n711_, new_n709_, new_n710_ );
nand g574 ( new_n712_, new_n711_, keyIn_0_54 );
not g575 ( new_n713_, keyIn_0_54 );
nand g576 ( new_n714_, new_n709_, new_n713_, new_n710_ );
nand g577 ( N742, new_n712_, new_n714_ );
not g578 ( new_n716_, keyIn_0_55 );
nand g579 ( new_n717_, new_n680_, new_n517_ );
nand g580 ( new_n718_, new_n717_, keyIn_0_43 );
not g581 ( new_n719_, keyIn_0_43 );
nand g582 ( new_n720_, new_n680_, new_n719_, new_n517_ );
nand g583 ( new_n721_, new_n718_, new_n720_ );
nand g584 ( new_n722_, new_n721_, N77 );
nand g585 ( new_n723_, new_n718_, new_n158_, new_n720_ );
nand g586 ( new_n724_, new_n722_, new_n723_ );
nand g587 ( new_n725_, new_n724_, new_n716_ );
nand g588 ( new_n726_, new_n722_, keyIn_0_55, new_n723_ );
nand g589 ( N743, new_n725_, new_n726_ );
not g590 ( new_n728_, keyIn_0_44 );
not g591 ( new_n729_, keyIn_0_38 );
nor g592 ( new_n730_, new_n674_, new_n430_, new_n495_ );
nand g593 ( new_n731_, new_n672_, new_n730_ );
nand g594 ( new_n732_, new_n731_, new_n729_ );
nand g595 ( new_n733_, new_n672_, keyIn_0_38, new_n730_ );
nand g596 ( new_n734_, new_n732_, new_n733_ );
nand g597 ( new_n735_, new_n734_, new_n288_ );
nand g598 ( new_n736_, new_n735_, new_n728_ );
nand g599 ( new_n737_, new_n734_, keyIn_0_44, new_n288_ );
nand g600 ( new_n738_, new_n736_, new_n737_ );
nand g601 ( new_n739_, new_n738_, new_n140_ );
nand g602 ( new_n740_, new_n736_, N81, new_n737_ );
nand g603 ( new_n741_, new_n739_, new_n740_ );
nand g604 ( new_n742_, new_n741_, keyIn_0_56 );
not g605 ( new_n743_, keyIn_0_56 );
nand g606 ( new_n744_, new_n739_, new_n743_, new_n740_ );
nand g607 ( N744, new_n742_, new_n744_ );
not g608 ( new_n746_, keyIn_0_57 );
nand g609 ( new_n747_, new_n734_, new_n346_ );
nand g610 ( new_n748_, new_n747_, keyIn_0_45 );
not g611 ( new_n749_, keyIn_0_45 );
nand g612 ( new_n750_, new_n734_, new_n749_, new_n346_ );
nand g613 ( new_n751_, new_n748_, new_n750_ );
nand g614 ( new_n752_, new_n751_, N85 );
nand g615 ( new_n753_, new_n748_, new_n138_, new_n750_ );
nand g616 ( new_n754_, new_n752_, new_n753_ );
nand g617 ( new_n755_, new_n754_, new_n746_ );
nand g618 ( new_n756_, new_n752_, keyIn_0_57, new_n753_ );
nand g619 ( N745, new_n755_, new_n756_ );
nand g620 ( new_n758_, new_n734_, new_n399_ );
nand g621 ( new_n759_, new_n758_, keyIn_0_46 );
not g622 ( new_n760_, keyIn_0_46 );
nand g623 ( new_n761_, new_n734_, new_n760_, new_n399_ );
nand g624 ( new_n762_, new_n759_, new_n761_ );
nand g625 ( new_n763_, new_n762_, N89 );
nand g626 ( new_n764_, new_n759_, new_n143_, new_n761_ );
nand g627 ( new_n765_, new_n763_, new_n764_ );
nand g628 ( new_n766_, new_n765_, keyIn_0_58 );
not g629 ( new_n767_, keyIn_0_58 );
nand g630 ( new_n768_, new_n763_, new_n767_, new_n764_ );
nand g631 ( N746, new_n766_, new_n768_ );
not g632 ( new_n770_, keyIn_0_59 );
nand g633 ( new_n771_, new_n734_, new_n517_ );
nand g634 ( new_n772_, new_n771_, keyIn_0_47 );
not g635 ( new_n773_, keyIn_0_47 );
nand g636 ( new_n774_, new_n734_, new_n773_, new_n517_ );
nand g637 ( new_n775_, new_n772_, new_n774_ );
nand g638 ( new_n776_, new_n775_, N93 );
nand g639 ( new_n777_, new_n772_, new_n144_, new_n774_ );
nand g640 ( new_n778_, new_n776_, new_n777_ );
nand g641 ( new_n779_, new_n778_, new_n770_ );
nand g642 ( new_n780_, new_n776_, keyIn_0_59, new_n777_ );
nand g643 ( N747, new_n779_, new_n780_ );
nor g644 ( new_n782_, new_n673_, new_n188_, new_n466_ );
nand g645 ( new_n783_, new_n672_, new_n782_ );
nand g646 ( new_n784_, new_n783_, keyIn_0_39 );
not g647 ( new_n785_, keyIn_0_39 );
nand g648 ( new_n786_, new_n672_, new_n785_, new_n782_ );
nand g649 ( new_n787_, new_n784_, new_n786_ );
nand g650 ( new_n788_, new_n787_, new_n288_ );
nand g651 ( new_n789_, new_n788_, keyIn_0_48 );
not g652 ( new_n790_, keyIn_0_48 );
nand g653 ( new_n791_, new_n787_, new_n790_, new_n288_ );
nand g654 ( new_n792_, new_n789_, new_n791_ );
nand g655 ( new_n793_, new_n792_, N97 );
nand g656 ( new_n794_, new_n789_, new_n401_, new_n791_ );
nand g657 ( new_n795_, new_n793_, new_n794_ );
nand g658 ( new_n796_, new_n795_, keyIn_0_60 );
not g659 ( new_n797_, keyIn_0_60 );
nand g660 ( new_n798_, new_n793_, new_n797_, new_n794_ );
nand g661 ( N748, new_n796_, new_n798_ );
not g662 ( new_n800_, keyIn_0_49 );
nand g663 ( new_n801_, new_n787_, new_n346_ );
nand g664 ( new_n802_, new_n801_, new_n800_ );
nand g665 ( new_n803_, new_n787_, keyIn_0_49, new_n346_ );
nand g666 ( new_n804_, new_n802_, new_n803_ );
nand g667 ( new_n805_, new_n804_, new_n336_ );
nand g668 ( new_n806_, new_n802_, N101, new_n803_ );
nand g669 ( new_n807_, new_n805_, new_n806_ );
nand g670 ( new_n808_, new_n807_, keyIn_0_61 );
not g671 ( new_n809_, keyIn_0_61 );
nand g672 ( new_n810_, new_n805_, new_n809_, new_n806_ );
nand g673 ( N749, new_n808_, new_n810_ );
not g674 ( new_n812_, keyIn_0_50 );
nand g675 ( new_n813_, new_n787_, new_n399_ );
nand g676 ( new_n814_, new_n813_, new_n812_ );
nand g677 ( new_n815_, new_n787_, keyIn_0_50, new_n399_ );
nand g678 ( new_n816_, new_n814_, new_n815_ );
nand g679 ( new_n817_, new_n816_, new_n379_ );
nand g680 ( new_n818_, new_n814_, N105, new_n815_ );
nand g681 ( new_n819_, new_n817_, new_n818_ );
nand g682 ( new_n820_, new_n819_, keyIn_0_62 );
not g683 ( new_n821_, keyIn_0_62 );
nand g684 ( new_n822_, new_n817_, new_n821_, new_n818_ );
nand g685 ( N750, new_n820_, new_n822_ );
not g686 ( new_n824_, keyIn_0_63 );
nand g687 ( new_n825_, new_n787_, new_n517_ );
nand g688 ( new_n826_, new_n825_, keyIn_0_51 );
not g689 ( new_n827_, keyIn_0_51 );
nand g690 ( new_n828_, new_n787_, new_n827_, new_n517_ );
nand g691 ( new_n829_, new_n826_, new_n828_ );
nand g692 ( new_n830_, new_n829_, new_n404_ );
nand g693 ( new_n831_, new_n826_, N109, new_n828_ );
nand g694 ( new_n832_, new_n830_, new_n831_ );
nand g695 ( new_n833_, new_n832_, new_n824_ );
nand g696 ( new_n834_, new_n830_, keyIn_0_63, new_n831_ );
nand g697 ( N751, new_n833_, new_n834_ );
not g698 ( new_n836_, new_n672_ );
nor g699 ( new_n837_, new_n836_, new_n465_, new_n495_ );
nand g700 ( new_n838_, new_n837_, new_n288_ );
nand g701 ( new_n839_, new_n838_, N113 );
nand g702 ( new_n840_, new_n837_, new_n435_, new_n288_ );
nand g703 ( N752, new_n839_, new_n840_ );
nand g704 ( new_n842_, new_n837_, new_n346_ );
nand g705 ( new_n843_, new_n842_, N117 );
nand g706 ( new_n844_, new_n837_, new_n337_, new_n346_ );
nand g707 ( N753, new_n843_, new_n844_ );
nand g708 ( new_n846_, new_n837_, new_n399_ );
nand g709 ( new_n847_, new_n846_, N121 );
nand g710 ( new_n848_, new_n837_, new_n377_, new_n399_ );
nand g711 ( N754, new_n847_, new_n848_ );
nand g712 ( new_n850_, new_n837_, new_n517_ );
nand g713 ( new_n851_, new_n850_, N125 );
nand g714 ( new_n852_, new_n837_, new_n438_, new_n517_ );
nand g715 ( N755, new_n851_, new_n852_ );
endmodule