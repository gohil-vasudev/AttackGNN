module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n236_, new_n976_, new_n1009_, new_n479_, new_n955_, new_n608_, new_n888_, new_n847_, new_n250_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1048_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n1025_, new_n566_, new_n641_, new_n339_, new_n365_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n1057_, new_n670_, new_n1024_, new_n456_, new_n691_, new_n682_, new_n812_, new_n911_, new_n679_, new_n937_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n419_, new_n728_, new_n624_, new_n534_, new_n819_, new_n637_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n695_, new_n240_, new_n660_, new_n413_, new_n1060_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n1045_, new_n500_, new_n898_, new_n786_, new_n799_, new_n946_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n862_, new_n742_, new_n892_, new_n427_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n959_, new_n990_, new_n774_, new_n716_, new_n701_, new_n792_, new_n1058_, new_n257_, new_n481_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n1059_, new_n634_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n1050_, new_n903_, new_n230_, new_n983_, new_n281_, new_n430_, new_n822_, new_n844_, new_n1018_, new_n855_, new_n606_, new_n1037_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n1054_, new_n385_, new_n1049_, new_n829_, new_n988_, new_n478_, new_n461_, new_n710_, new_n971_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n683_, new_n511_, new_n463_, new_n303_, new_n510_, new_n966_, new_n351_, new_n517_, new_n325_, new_n609_, new_n1031_, new_n961_, new_n890_, new_n530_, new_n318_, new_n1006_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n1005_, new_n999_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n956_, new_n763_, new_n960_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n970_, new_n995_, new_n1035_, new_n271_, new_n274_, new_n991_, new_n1044_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n1051_, new_n1053_, new_n423_, new_n498_, new_n492_, new_n496_, new_n1046_, new_n650_, new_n708_, new_n750_, new_n887_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n734_, new_n912_, new_n925_, new_n1062_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n820_, new_n771_, new_n388_, new_n979_, new_n1028_, new_n508_, new_n714_, new_n483_, new_n1004_, new_n394_, new_n299_, new_n1007_, new_n935_, new_n882_, new_n657_, new_n929_, new_n652_, new_n314_, new_n582_, new_n986_, new_n1020_, new_n363_, new_n441_, new_n785_, new_n477_, new_n664_, new_n600_, new_n280_, new_n917_, new_n1041_, new_n426_, new_n1036_, new_n235_, new_n398_, new_n301_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n541_, new_n458_, new_n854_, new_n447_, new_n1026_, new_n267_, new_n473_, new_n790_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n969_, new_n263_, new_n334_, new_n835_, new_n341_, new_n378_, new_n996_, new_n621_, new_n846_, new_n915_, new_n349_, new_n244_, new_n488_, new_n524_, new_n705_, new_n277_, new_n848_, new_n943_, new_n874_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n632_, new_n1039_, new_n671_, new_n965_, new_n528_, new_n952_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n397_, new_n729_, new_n975_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n559_, new_n948_, new_n762_, new_n1055_, new_n838_, new_n923_, new_n469_, new_n391_, new_n437_, new_n295_, new_n359_, new_n794_, new_n628_, new_n409_, new_n745_, new_n457_, new_n553_, new_n1061_, new_n668_, new_n333_, new_n1002_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n1032_, new_n276_, new_n688_, new_n384_, new_n900_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n1034_, new_n296_, new_n661_, new_n308_, new_n1000_, new_n633_, new_n797_, new_n784_, new_n258_, new_n724_, new_n860_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n938_, new_n809_, new_n654_, new_n713_, new_n880_, new_n604_, new_n227_, new_n690_, new_n416_, new_n1043_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n967_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n749_, new_n861_, new_n310_, new_n275_, new_n998_, new_n1056_, new_n352_, new_n931_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n1064_, new_n1065_, new_n493_, new_n547_, new_n907_, new_n264_, new_n665_, new_n800_, new_n379_, new_n897_, new_n1012_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n963_, new_n270_, new_n570_, new_n598_, new_n893_, new_n993_, new_n1063_, new_n824_, new_n520_, new_n1001_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n825_, new_n858_, new_n557_, new_n260_, new_n936_, new_n251_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1016_, new_n748_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n879_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n313_, new_n382_, new_n583_, new_n239_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n428_, new_n916_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n302_, new_n755_, new_n225_, new_n1040_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n221_, new_n450_, new_n345_, new_n298_, new_n499_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n468_, new_n977_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n337_, new_n623_, new_n446_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n972_, new_n1067_, new_n891_, new_n631_, new_n453_, new_n516_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n252_, new_n585_, new_n751_, new_n312_, new_n535_, new_n1038_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n597_, new_n978_, new_n408_, new_n470_, new_n769_, new_n1069_, new_n651_, new_n433_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n992_, new_n265_, new_n732_, new_n687_, new_n370_, new_n1029_, new_n689_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n1052_, new_n1017_, new_n550_, new_n1068_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n989_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n319_, new_n1008_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n957_, new_n754_, new_n1047_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n330_, new_n727_, new_n375_, new_n962_, new_n760_, new_n627_, new_n704_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n357_, new_n320_, new_n780_, new_n984_, new_n245_, new_n643_, new_n474_, new_n467_, new_n1013_, new_n404_, new_n490_, new_n560_, new_n865_, new_n1027_, new_n358_, new_n877_, new_n348_, new_n610_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n1011_, new_n425_, new_n896_, new_n802_, new_n697_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n866_, new_n540_, new_n1066_, new_n434_, new_n947_, new_n994_, new_n982_, new_n422_, new_n964_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n551_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n521_, new_n1042_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n573_, new_n765_, new_n405_;

nand g000 ( new_n215_, N29, N42, N75 );
not g001 ( N388, new_n215_ );
nand g002 ( new_n217_, N29, N36, N80 );
not g003 ( N389, new_n217_ );
nand g004 ( new_n219_, N29, N36, N42 );
not g005 ( N390, new_n219_ );
nand g006 ( new_n221_, N85, N86 );
not g007 ( N391, new_n221_ );
nand g008 ( new_n223_, N1, N8 );
not g009 ( new_n224_, new_n223_ );
nand g010 ( new_n225_, new_n224_, N13, N17 );
not g011 ( N418, new_n225_ );
not g012 ( new_n227_, N13 );
not g013 ( new_n228_, N17 );
nand g014 ( new_n229_, N1, N26 );
nor g015 ( new_n230_, new_n229_, new_n227_, new_n228_ );
nand g016 ( N419, new_n230_, new_n219_ );
nand g017 ( N420, N59, N75, N80 );
nand g018 ( N421, N36, N59, N80 );
nand g019 ( N422, N36, N42, N59 );
not g020 ( new_n235_, N90 );
nor g021 ( new_n236_, N87, N88 );
nor g022 ( N423, new_n236_, new_n235_ );
nand g023 ( N446, new_n230_, N390 );
nand g024 ( new_n239_, N1, N26, N51 );
nand g025 ( new_n240_, new_n239_, keyIn_0_0 );
not g026 ( new_n241_, keyIn_0_0 );
nand g027 ( new_n242_, new_n241_, N1, N26, N51 );
nand g028 ( N447, new_n240_, new_n242_ );
nand g029 ( new_n244_, new_n224_, N13, N55 );
nand g030 ( new_n245_, N29, N68 );
nor g031 ( N448, new_n244_, new_n245_ );
not g032 ( new_n247_, keyIn_0_10 );
not g033 ( new_n248_, new_n244_ );
nand g034 ( new_n249_, N59, N68 );
not g035 ( new_n250_, new_n249_ );
nand g036 ( new_n251_, new_n248_, new_n247_, N74, new_n250_ );
nand g037 ( new_n252_, new_n248_, N74, new_n250_ );
nand g038 ( new_n253_, new_n252_, keyIn_0_10 );
nand g039 ( N449, new_n253_, new_n251_ );
not g040 ( new_n255_, N89 );
nor g041 ( N450, new_n236_, new_n255_ );
nor g042 ( new_n257_, N91, N96 );
not g043 ( new_n258_, new_n257_ );
nand g044 ( new_n259_, N91, N96 );
nand g045 ( new_n260_, new_n258_, keyIn_0_15, new_n259_ );
nand g046 ( new_n261_, N101, N106 );
not g047 ( new_n262_, new_n261_ );
nor g048 ( new_n263_, N101, N106 );
nor g049 ( new_n264_, new_n262_, new_n263_ );
nand g050 ( new_n265_, new_n260_, new_n264_ );
not g051 ( new_n266_, new_n265_ );
nor g052 ( new_n267_, new_n260_, new_n264_ );
nor g053 ( new_n268_, new_n266_, new_n267_ );
not g054 ( new_n269_, new_n268_ );
nand g055 ( new_n270_, new_n269_, N130 );
not g056 ( new_n271_, N130 );
nand g057 ( new_n272_, new_n268_, new_n271_ );
nand g058 ( new_n273_, new_n270_, new_n272_ );
not g059 ( new_n274_, N135 );
not g060 ( new_n275_, N111 );
not g061 ( new_n276_, N116 );
nand g062 ( new_n277_, new_n275_, new_n276_ );
nand g063 ( new_n278_, N111, N116 );
nand g064 ( new_n279_, new_n277_, new_n278_ );
not g065 ( new_n280_, N121 );
not g066 ( new_n281_, N126 );
nand g067 ( new_n282_, new_n280_, new_n281_ );
nand g068 ( new_n283_, N121, N126 );
nand g069 ( new_n284_, new_n282_, new_n283_ );
nand g070 ( new_n285_, new_n279_, new_n284_ );
nand g071 ( new_n286_, new_n277_, new_n282_, new_n278_, new_n283_ );
nand g072 ( new_n287_, new_n285_, new_n286_ );
nand g073 ( new_n288_, new_n287_, new_n274_ );
nand g074 ( new_n289_, new_n285_, N135, new_n286_ );
nand g075 ( new_n290_, new_n288_, new_n289_ );
nand g076 ( new_n291_, new_n273_, new_n290_ );
nand g077 ( new_n292_, new_n270_, new_n272_, new_n288_, new_n289_ );
nand g078 ( new_n293_, new_n291_, new_n292_ );
not g079 ( N767, new_n293_ );
not g080 ( new_n295_, N159 );
not g081 ( new_n296_, N165 );
nand g082 ( new_n297_, new_n295_, new_n296_ );
nand g083 ( new_n298_, N159, N165 );
nand g084 ( new_n299_, new_n297_, new_n298_ );
not g085 ( new_n300_, N171 );
not g086 ( new_n301_, N177 );
nand g087 ( new_n302_, new_n300_, new_n301_ );
nand g088 ( new_n303_, N171, N177 );
nand g089 ( new_n304_, new_n302_, new_n303_ );
nand g090 ( new_n305_, new_n299_, new_n304_ );
nand g091 ( new_n306_, new_n297_, new_n302_, new_n298_, new_n303_ );
nand g092 ( new_n307_, new_n305_, new_n306_ );
nand g093 ( new_n308_, new_n307_, new_n271_ );
nand g094 ( new_n309_, new_n305_, N130, new_n306_ );
nand g095 ( new_n310_, new_n308_, new_n309_ );
not g096 ( new_n311_, N207 );
not g097 ( new_n312_, N183 );
not g098 ( new_n313_, N189 );
nand g099 ( new_n314_, new_n312_, new_n313_ );
nand g100 ( new_n315_, N183, N189 );
nand g101 ( new_n316_, new_n314_, new_n315_ );
not g102 ( new_n317_, N195 );
not g103 ( new_n318_, N201 );
nand g104 ( new_n319_, new_n317_, new_n318_ );
nand g105 ( new_n320_, N195, N201 );
nand g106 ( new_n321_, new_n319_, new_n320_ );
nand g107 ( new_n322_, new_n316_, new_n321_ );
nand g108 ( new_n323_, new_n314_, new_n319_, new_n315_, new_n320_ );
nand g109 ( new_n324_, new_n322_, new_n323_ );
nand g110 ( new_n325_, new_n324_, new_n311_ );
nand g111 ( new_n326_, new_n322_, N207, new_n323_ );
nand g112 ( new_n327_, new_n325_, new_n326_ );
nand g113 ( new_n328_, new_n310_, new_n327_ );
nand g114 ( new_n329_, new_n308_, new_n325_, new_n309_, new_n326_ );
nand g115 ( new_n330_, new_n328_, new_n329_ );
not g116 ( N768, new_n330_ );
not g117 ( new_n332_, keyIn_0_38 );
nand g118 ( new_n333_, N447, keyIn_0_8 );
not g119 ( new_n334_, keyIn_0_8 );
nand g120 ( new_n335_, new_n240_, new_n334_, new_n242_ );
nand g121 ( new_n336_, new_n333_, new_n335_ );
nand g122 ( new_n337_, new_n336_, keyIn_0_14 );
not g123 ( new_n338_, keyIn_0_14 );
nand g124 ( new_n339_, new_n333_, new_n338_, new_n335_ );
nand g125 ( new_n340_, new_n337_, new_n339_ );
nand g126 ( new_n341_, keyIn_0_5, N59, N156 );
not g127 ( new_n342_, keyIn_0_5 );
nand g128 ( new_n343_, N59, N156 );
nand g129 ( new_n344_, new_n343_, new_n342_ );
nand g130 ( new_n345_, new_n344_, new_n341_ );
not g131 ( new_n346_, new_n345_ );
nand g132 ( new_n347_, new_n340_, keyIn_0_21, N17, new_n346_ );
not g133 ( new_n348_, keyIn_0_21 );
nand g134 ( new_n349_, new_n340_, N17, new_n346_ );
nand g135 ( new_n350_, new_n349_, new_n348_ );
nand g136 ( new_n351_, new_n350_, N1, new_n347_ );
nand g137 ( new_n352_, new_n351_, keyIn_0_25 );
not g138 ( new_n353_, keyIn_0_25 );
nand g139 ( new_n354_, new_n350_, new_n353_, N1, new_n347_ );
nand g140 ( new_n355_, new_n352_, new_n354_ );
nand g141 ( new_n356_, new_n355_, N153 );
nand g142 ( new_n357_, new_n356_, new_n332_ );
nand g143 ( new_n358_, new_n355_, keyIn_0_38, N153 );
nand g144 ( new_n359_, new_n357_, new_n358_ );
not g145 ( new_n360_, keyIn_0_39 );
not g146 ( new_n361_, keyIn_0_22 );
not g147 ( new_n362_, keyIn_0_13 );
not g148 ( new_n363_, N42 );
nand g149 ( new_n364_, new_n228_, new_n363_ );
nand g150 ( new_n365_, new_n364_, keyIn_0_6 );
nand g151 ( new_n366_, N17, N42 );
nand g152 ( new_n367_, new_n366_, keyIn_0_7 );
not g153 ( new_n368_, keyIn_0_7 );
nand g154 ( new_n369_, new_n368_, N17, N42 );
not g155 ( new_n370_, new_n369_ );
nor g156 ( new_n371_, keyIn_0_6, N17, N42 );
nor g157 ( new_n372_, new_n370_, new_n371_ );
nand g158 ( new_n373_, new_n372_, new_n362_, new_n365_, new_n367_ );
not g159 ( new_n374_, new_n371_ );
nand g160 ( new_n375_, new_n374_, new_n365_, new_n367_, new_n369_ );
nand g161 ( new_n376_, new_n375_, keyIn_0_13 );
nand g162 ( new_n377_, new_n376_, new_n373_, N59, N156 );
not g163 ( new_n378_, new_n377_ );
nand g164 ( new_n379_, new_n378_, new_n340_ );
nand g165 ( new_n380_, new_n379_, keyIn_0_20 );
not g166 ( new_n381_, keyIn_0_20 );
nand g167 ( new_n382_, new_n378_, new_n340_, new_n381_ );
not g168 ( new_n383_, keyIn_0_11 );
not g169 ( new_n384_, keyIn_0_3 );
nand g170 ( new_n385_, N42, N59, N75 );
nand g171 ( new_n386_, new_n385_, new_n384_ );
nand g172 ( new_n387_, keyIn_0_3, N42, N59, N75 );
nand g173 ( new_n388_, new_n386_, new_n387_ );
nand g174 ( new_n389_, new_n388_, new_n383_ );
nand g175 ( new_n390_, new_n386_, keyIn_0_11, new_n387_ );
nand g176 ( new_n391_, new_n389_, new_n390_ );
nand g177 ( new_n392_, N1, N8, N17, N51 );
nand g178 ( new_n393_, new_n392_, keyIn_0_1 );
not g179 ( new_n394_, keyIn_0_1 );
nand g180 ( new_n395_, new_n224_, new_n394_, N17, N51 );
nand g181 ( new_n396_, new_n395_, new_n393_ );
nand g182 ( new_n397_, new_n396_, keyIn_0_9 );
not g183 ( new_n398_, keyIn_0_9 );
nand g184 ( new_n399_, new_n395_, new_n398_, new_n393_ );
nand g185 ( new_n400_, new_n391_, new_n397_, new_n399_ );
nand g186 ( new_n401_, new_n400_, keyIn_0_16 );
not g187 ( new_n402_, keyIn_0_16 );
nand g188 ( new_n403_, new_n391_, new_n397_, new_n402_, new_n399_ );
nand g189 ( new_n404_, new_n401_, new_n403_ );
not g190 ( new_n405_, new_n404_ );
nand g191 ( new_n406_, new_n380_, new_n405_, new_n382_ );
nand g192 ( new_n407_, new_n406_, new_n361_ );
nand g193 ( new_n408_, new_n380_, new_n405_, keyIn_0_22, new_n382_ );
nand g194 ( new_n409_, new_n407_, N126, new_n408_ );
nand g195 ( new_n410_, new_n409_, new_n360_ );
nand g196 ( new_n411_, new_n407_, keyIn_0_39, N126, new_n408_ );
nand g197 ( new_n412_, new_n410_, new_n411_ );
not g198 ( new_n413_, new_n412_ );
nand g199 ( new_n414_, new_n413_, new_n359_ );
nand g200 ( new_n415_, new_n414_, keyIn_0_45 );
not g201 ( new_n416_, keyIn_0_45 );
nand g202 ( new_n417_, new_n413_, new_n359_, new_n416_ );
nand g203 ( new_n418_, new_n415_, new_n417_ );
not g204 ( new_n419_, keyIn_0_29 );
nand g205 ( new_n420_, N29, N75, N80 );
nand g206 ( new_n421_, new_n420_, keyIn_0_2 );
not g207 ( new_n422_, keyIn_0_2 );
nand g208 ( new_n423_, new_n422_, N29, N75, N80 );
nand g209 ( new_n424_, new_n340_, new_n421_, new_n423_ );
not g210 ( new_n425_, new_n424_ );
nand g211 ( new_n426_, new_n425_, N55 );
nand g212 ( new_n427_, new_n426_, keyIn_0_19 );
not g213 ( new_n428_, keyIn_0_19 );
nand g214 ( new_n429_, new_n425_, new_n428_, N55 );
nand g215 ( new_n430_, new_n427_, new_n429_ );
not g216 ( new_n431_, keyIn_0_12 );
not g217 ( new_n432_, N268 );
nor g218 ( new_n433_, new_n432_, keyIn_0_4 );
nand g219 ( new_n434_, new_n432_, keyIn_0_4 );
not g220 ( new_n435_, new_n434_ );
nor g221 ( new_n436_, new_n435_, new_n433_ );
not g222 ( new_n437_, new_n436_ );
nand g223 ( new_n438_, new_n437_, new_n431_ );
nand g224 ( new_n439_, new_n436_, keyIn_0_12 );
nand g225 ( new_n440_, new_n438_, new_n439_ );
not g226 ( new_n441_, new_n440_ );
nand g227 ( new_n442_, new_n430_, new_n441_ );
not g228 ( new_n443_, new_n442_ );
nand g229 ( new_n444_, new_n443_, new_n419_ );
nand g230 ( new_n445_, new_n442_, keyIn_0_29 );
nand g231 ( new_n446_, new_n444_, new_n445_ );
nand g232 ( new_n447_, new_n418_, new_n446_ );
nand g233 ( new_n448_, new_n447_, keyIn_0_50 );
not g234 ( new_n449_, keyIn_0_50 );
nand g235 ( new_n450_, new_n418_, new_n449_, new_n446_ );
nand g236 ( new_n451_, new_n448_, new_n450_ );
nand g237 ( new_n452_, new_n451_, N201 );
nand g238 ( new_n453_, new_n452_, keyIn_0_60 );
not g239 ( new_n454_, keyIn_0_60 );
nand g240 ( new_n455_, new_n451_, new_n454_, N201 );
nand g241 ( new_n456_, new_n453_, new_n455_ );
nand g242 ( new_n457_, new_n448_, new_n318_, new_n450_ );
nand g243 ( new_n458_, new_n457_, keyIn_0_61 );
not g244 ( new_n459_, keyIn_0_61 );
nand g245 ( new_n460_, new_n448_, new_n459_, new_n318_, new_n450_ );
nand g246 ( new_n461_, new_n458_, new_n460_ );
nand g247 ( new_n462_, new_n456_, new_n461_ );
not g248 ( new_n463_, new_n462_ );
nand g249 ( new_n464_, new_n463_, N261 );
not g250 ( new_n465_, N261 );
nand g251 ( new_n466_, new_n462_, new_n465_ );
nand g252 ( new_n467_, new_n464_, N219, new_n466_ );
not g253 ( new_n468_, keyIn_0_67 );
nand g254 ( new_n469_, new_n456_, new_n468_ );
nand g255 ( new_n470_, new_n453_, keyIn_0_67, new_n455_ );
nand g256 ( new_n471_, new_n469_, new_n470_ );
nand g257 ( new_n472_, new_n471_, N237 );
nand g258 ( new_n473_, new_n463_, N228 );
nand g259 ( new_n474_, new_n451_, N246 );
nand g260 ( new_n475_, N42, N72, N73 );
nor g261 ( new_n476_, new_n244_, new_n475_, new_n249_ );
nand g262 ( new_n477_, new_n476_, N201 );
nand g263 ( new_n478_, N121, N210 );
nand g264 ( new_n479_, N255, N267 );
nand g265 ( new_n480_, new_n474_, new_n477_, new_n478_, new_n479_ );
not g266 ( new_n481_, new_n480_ );
nand g267 ( N850, new_n467_, new_n472_, new_n473_, new_n481_ );
not g268 ( new_n483_, keyIn_0_112 );
not g269 ( new_n484_, keyIn_0_92 );
not g270 ( new_n485_, keyIn_0_80 );
not g271 ( new_n486_, keyIn_0_77 );
not g272 ( new_n487_, keyIn_0_75 );
not g273 ( new_n488_, keyIn_0_73 );
not g274 ( new_n489_, keyIn_0_59 );
not g275 ( new_n490_, keyIn_0_49 );
nand g276 ( new_n491_, new_n355_, N149 );
nand g277 ( new_n492_, new_n491_, keyIn_0_36 );
not g278 ( new_n493_, keyIn_0_36 );
nand g279 ( new_n494_, new_n355_, new_n493_, N149 );
nand g280 ( new_n495_, new_n492_, new_n494_ );
nand g281 ( new_n496_, new_n407_, N121, new_n408_ );
nand g282 ( new_n497_, new_n496_, keyIn_0_37 );
not g283 ( new_n498_, keyIn_0_37 );
nand g284 ( new_n499_, new_n407_, new_n498_, N121, new_n408_ );
nand g285 ( new_n500_, new_n497_, new_n499_ );
nand g286 ( new_n501_, new_n495_, keyIn_0_44, new_n500_ );
nand g287 ( new_n502_, new_n443_, keyIn_0_28 );
not g288 ( new_n503_, keyIn_0_28 );
nand g289 ( new_n504_, new_n442_, new_n503_ );
nand g290 ( new_n505_, new_n502_, new_n504_ );
not g291 ( new_n506_, keyIn_0_44 );
nand g292 ( new_n507_, new_n495_, new_n500_ );
nand g293 ( new_n508_, new_n507_, new_n506_ );
nand g294 ( new_n509_, new_n508_, new_n501_, new_n505_ );
nand g295 ( new_n510_, new_n509_, new_n490_ );
nand g296 ( new_n511_, new_n508_, keyIn_0_49, new_n501_, new_n505_ );
nand g297 ( new_n512_, new_n510_, new_n511_ );
nand g298 ( new_n513_, new_n512_, new_n317_ );
nand g299 ( new_n514_, new_n513_, new_n489_ );
nand g300 ( new_n515_, new_n512_, keyIn_0_59, new_n317_ );
nand g301 ( new_n516_, new_n514_, new_n515_ );
not g302 ( new_n517_, keyIn_0_57 );
not g303 ( new_n518_, keyIn_0_43 );
not g304 ( new_n519_, keyIn_0_34 );
nand g305 ( new_n520_, new_n355_, new_n519_, N146 );
nand g306 ( new_n521_, new_n355_, N146 );
nand g307 ( new_n522_, new_n521_, keyIn_0_34 );
nand g308 ( new_n523_, new_n407_, N116, new_n408_ );
nand g309 ( new_n524_, new_n523_, keyIn_0_35 );
not g310 ( new_n525_, keyIn_0_35 );
nand g311 ( new_n526_, new_n407_, new_n525_, N116, new_n408_ );
nand g312 ( new_n527_, new_n524_, new_n526_ );
not g313 ( new_n528_, new_n527_ );
nand g314 ( new_n529_, new_n528_, new_n518_, new_n520_, new_n522_ );
not g315 ( new_n530_, keyIn_0_27 );
nand g316 ( new_n531_, new_n443_, new_n530_ );
nand g317 ( new_n532_, new_n442_, keyIn_0_27 );
nand g318 ( new_n533_, new_n531_, new_n532_ );
nand g319 ( new_n534_, new_n522_, new_n520_, new_n524_, new_n526_ );
nand g320 ( new_n535_, new_n534_, keyIn_0_43 );
nand g321 ( new_n536_, new_n529_, new_n535_, new_n533_ );
nand g322 ( new_n537_, new_n536_, keyIn_0_48 );
not g323 ( new_n538_, keyIn_0_48 );
nand g324 ( new_n539_, new_n529_, new_n535_, new_n538_, new_n533_ );
nand g325 ( new_n540_, new_n537_, new_n313_, new_n539_ );
nand g326 ( new_n541_, new_n540_, new_n517_ );
nand g327 ( new_n542_, new_n537_, keyIn_0_57, new_n313_, new_n539_ );
nand g328 ( new_n543_, new_n541_, new_n542_ );
nor g329 ( new_n544_, new_n516_, new_n543_ );
nand g330 ( new_n545_, new_n471_, new_n544_ );
nand g331 ( new_n546_, new_n545_, new_n488_ );
nand g332 ( new_n547_, new_n471_, keyIn_0_73, new_n544_ );
not g333 ( new_n548_, new_n543_ );
not g334 ( new_n549_, keyIn_0_66 );
not g335 ( new_n550_, keyIn_0_58 );
nand g336 ( new_n551_, new_n510_, N195, new_n511_ );
nand g337 ( new_n552_, new_n551_, new_n550_ );
nand g338 ( new_n553_, new_n510_, keyIn_0_58, N195, new_n511_ );
nand g339 ( new_n554_, new_n552_, new_n553_ );
nand g340 ( new_n555_, new_n554_, new_n549_ );
nand g341 ( new_n556_, new_n552_, keyIn_0_66, new_n553_ );
nand g342 ( new_n557_, new_n555_, new_n556_ );
nand g343 ( new_n558_, new_n557_, new_n548_ );
nand g344 ( new_n559_, new_n558_, keyIn_0_72 );
not g345 ( new_n560_, keyIn_0_72 );
nand g346 ( new_n561_, new_n557_, new_n560_, new_n548_ );
nand g347 ( new_n562_, new_n559_, new_n561_ );
not g348 ( new_n563_, keyIn_0_71 );
not g349 ( new_n564_, keyIn_0_65 );
not g350 ( new_n565_, keyIn_0_56 );
nand g351 ( new_n566_, new_n537_, new_n539_ );
nand g352 ( new_n567_, new_n566_, N189 );
nand g353 ( new_n568_, new_n567_, new_n565_ );
nand g354 ( new_n569_, new_n566_, keyIn_0_56, N189 );
nand g355 ( new_n570_, new_n568_, new_n569_ );
nand g356 ( new_n571_, new_n570_, new_n564_ );
nand g357 ( new_n572_, new_n568_, keyIn_0_65, new_n569_ );
nand g358 ( new_n573_, new_n571_, new_n572_ );
nand g359 ( new_n574_, new_n573_, new_n563_ );
not g360 ( new_n575_, new_n516_ );
nand g361 ( new_n576_, new_n575_, N261, new_n461_, new_n548_ );
nand g362 ( new_n577_, new_n576_, keyIn_0_68 );
nand g363 ( new_n578_, new_n577_, new_n574_ );
not g364 ( new_n579_, keyIn_0_68 );
nand g365 ( new_n580_, new_n544_, new_n579_, N261, new_n461_ );
nand g366 ( new_n581_, new_n571_, keyIn_0_71, new_n572_ );
nand g367 ( new_n582_, new_n580_, new_n581_ );
nor g368 ( new_n583_, new_n578_, new_n582_ );
nand g369 ( new_n584_, new_n583_, new_n546_, new_n547_, new_n562_ );
nand g370 ( new_n585_, new_n584_, new_n487_ );
not g371 ( new_n586_, new_n562_ );
nand g372 ( new_n587_, new_n577_, new_n574_, new_n580_, new_n581_ );
nor g373 ( new_n588_, new_n586_, new_n587_ );
nand g374 ( new_n589_, new_n588_, keyIn_0_75, new_n546_, new_n547_ );
not g375 ( new_n590_, keyIn_0_54 );
not g376 ( new_n591_, keyIn_0_32 );
nand g377 ( new_n592_, new_n355_, N143 );
nand g378 ( new_n593_, new_n592_, new_n591_ );
nand g379 ( new_n594_, new_n355_, keyIn_0_32, N143 );
nand g380 ( new_n595_, new_n407_, new_n408_ );
not g381 ( new_n596_, new_n595_ );
nand g382 ( new_n597_, new_n596_, N111 );
nand g383 ( new_n598_, new_n597_, keyIn_0_33 );
not g384 ( new_n599_, keyIn_0_33 );
nand g385 ( new_n600_, new_n596_, new_n599_, N111 );
nand g386 ( new_n601_, new_n598_, new_n594_, new_n600_ );
not g387 ( new_n602_, new_n601_ );
nand g388 ( new_n603_, new_n602_, new_n593_ );
nand g389 ( new_n604_, new_n603_, keyIn_0_42 );
not g390 ( new_n605_, keyIn_0_42 );
nand g391 ( new_n606_, new_n602_, new_n605_, new_n593_ );
nand g392 ( new_n607_, new_n604_, new_n606_ );
nand g393 ( new_n608_, new_n443_, keyIn_0_26 );
not g394 ( new_n609_, keyIn_0_26 );
nand g395 ( new_n610_, new_n442_, new_n609_ );
nand g396 ( new_n611_, new_n608_, new_n610_ );
nand g397 ( new_n612_, new_n607_, new_n611_ );
nand g398 ( new_n613_, new_n612_, keyIn_0_47 );
not g399 ( new_n614_, keyIn_0_47 );
nand g400 ( new_n615_, new_n607_, new_n614_, new_n611_ );
nand g401 ( new_n616_, new_n613_, new_n615_ );
not g402 ( new_n617_, new_n616_ );
nand g403 ( new_n618_, new_n617_, N183 );
nand g404 ( new_n619_, new_n618_, new_n590_ );
nand g405 ( new_n620_, new_n617_, keyIn_0_54, N183 );
nand g406 ( new_n621_, new_n619_, new_n620_ );
not g407 ( new_n622_, new_n621_ );
not g408 ( new_n623_, keyIn_0_55 );
nand g409 ( new_n624_, new_n616_, new_n312_ );
nand g410 ( new_n625_, new_n624_, new_n623_ );
nand g411 ( new_n626_, new_n616_, keyIn_0_55, new_n312_ );
nand g412 ( new_n627_, new_n625_, new_n626_ );
nand g413 ( new_n628_, new_n622_, new_n627_ );
not g414 ( new_n629_, new_n628_ );
nand g415 ( new_n630_, new_n585_, new_n589_, new_n629_ );
nand g416 ( new_n631_, new_n630_, new_n486_ );
not g417 ( new_n632_, keyIn_0_76 );
nand g418 ( new_n633_, new_n585_, new_n589_ );
nand g419 ( new_n634_, new_n633_, new_n628_ );
nand g420 ( new_n635_, new_n634_, new_n632_ );
nand g421 ( new_n636_, new_n633_, keyIn_0_76, new_n628_ );
nand g422 ( new_n637_, new_n585_, new_n589_, keyIn_0_77, new_n629_ );
nand g423 ( new_n638_, new_n635_, new_n631_, new_n636_, new_n637_ );
not g424 ( new_n639_, new_n638_ );
nand g425 ( new_n640_, new_n639_, new_n485_ );
nand g426 ( new_n641_, new_n638_, keyIn_0_80 );
nand g427 ( new_n642_, new_n640_, N219, new_n641_ );
nand g428 ( new_n643_, new_n642_, keyIn_0_83 );
not g429 ( new_n644_, keyIn_0_83 );
nand g430 ( new_n645_, new_n640_, new_n644_, N219, new_n641_ );
nand g431 ( new_n646_, new_n643_, new_n645_ );
nand g432 ( new_n647_, N106, N210 );
nand g433 ( new_n648_, new_n646_, new_n647_ );
nand g434 ( new_n649_, new_n648_, new_n484_ );
nand g435 ( new_n650_, new_n646_, keyIn_0_92, new_n647_ );
nand g436 ( new_n651_, new_n649_, new_n650_ );
nand g437 ( new_n652_, new_n622_, keyIn_0_64 );
not g438 ( new_n653_, keyIn_0_64 );
nand g439 ( new_n654_, new_n621_, new_n653_ );
nand g440 ( new_n655_, new_n652_, new_n654_ );
nand g441 ( new_n656_, new_n655_, N237 );
not g442 ( new_n657_, new_n656_ );
nand g443 ( new_n658_, new_n629_, N228 );
nand g444 ( new_n659_, new_n476_, N183 );
nand g445 ( new_n660_, new_n617_, N246 );
nand g446 ( new_n661_, new_n658_, new_n659_, new_n660_ );
nor g447 ( new_n662_, new_n661_, new_n657_ );
nand g448 ( new_n663_, new_n651_, new_n662_ );
nand g449 ( new_n664_, new_n663_, keyIn_0_100 );
not g450 ( new_n665_, keyIn_0_100 );
nand g451 ( new_n666_, new_n651_, new_n665_, new_n662_ );
nand g452 ( new_n667_, new_n664_, new_n666_ );
nand g453 ( new_n668_, new_n667_, keyIn_0_106 );
not g454 ( new_n669_, keyIn_0_106 );
nand g455 ( new_n670_, new_n664_, new_n669_, new_n666_ );
nand g456 ( new_n671_, new_n668_, new_n670_ );
nand g457 ( new_n672_, new_n671_, new_n483_ );
nand g458 ( new_n673_, new_n668_, keyIn_0_112, new_n670_ );
nand g459 ( N863, new_n672_, new_n673_ );
nand g460 ( new_n675_, new_n548_, new_n570_ );
not g461 ( new_n676_, new_n675_ );
not g462 ( new_n677_, new_n557_ );
not g463 ( new_n678_, new_n471_ );
nand g464 ( new_n679_, new_n461_, N261 );
nand g465 ( new_n680_, new_n678_, new_n679_ );
nand g466 ( new_n681_, new_n680_, new_n575_ );
nand g467 ( new_n682_, new_n681_, new_n677_ );
nand g468 ( new_n683_, new_n682_, new_n676_ );
nand g469 ( new_n684_, new_n681_, new_n677_, new_n675_ );
nand g470 ( new_n685_, new_n683_, N219, new_n684_ );
nand g471 ( new_n686_, new_n573_, N237 );
nand g472 ( new_n687_, new_n676_, N228 );
nand g473 ( new_n688_, new_n566_, N246 );
nand g474 ( new_n689_, new_n476_, N189 );
nand g475 ( new_n690_, N111, N210 );
nand g476 ( new_n691_, N255, N259 );
nand g477 ( new_n692_, new_n688_, new_n689_, new_n690_, new_n691_ );
not g478 ( new_n693_, new_n692_ );
nand g479 ( N864, new_n685_, new_n686_, new_n687_, new_n693_ );
nor g480 ( new_n695_, new_n516_, new_n554_ );
nand g481 ( new_n696_, new_n680_, new_n695_ );
not g482 ( new_n697_, new_n695_ );
nand g483 ( new_n698_, new_n678_, new_n679_, new_n697_ );
nand g484 ( new_n699_, new_n696_, N219, new_n698_ );
nand g485 ( new_n700_, new_n699_, keyIn_0_84 );
not g486 ( new_n701_, keyIn_0_84 );
nand g487 ( new_n702_, new_n696_, new_n701_, N219, new_n698_ );
nand g488 ( new_n703_, new_n700_, new_n702_ );
nand g489 ( new_n704_, new_n557_, N237 );
nand g490 ( new_n705_, new_n695_, N228 );
nand g491 ( new_n706_, new_n510_, N246, new_n511_ );
nand g492 ( new_n707_, new_n476_, N195 );
nand g493 ( new_n708_, N116, N210 );
nand g494 ( new_n709_, N255, N260 );
nand g495 ( new_n710_, new_n706_, new_n707_, new_n708_, new_n709_ );
not g496 ( new_n711_, new_n710_ );
nand g497 ( N865, new_n703_, new_n704_, new_n705_, new_n711_ );
nand g498 ( new_n713_, new_n596_, N96 );
nand g499 ( new_n714_, new_n340_, new_n346_ );
not g500 ( new_n715_, new_n714_ );
nand g501 ( new_n716_, new_n715_, N55 );
nand g502 ( new_n717_, new_n716_, keyIn_0_17 );
not g503 ( new_n718_, keyIn_0_17 );
nand g504 ( new_n719_, new_n715_, new_n718_, N55 );
nand g505 ( new_n720_, new_n717_, new_n719_ );
not g506 ( new_n721_, new_n720_ );
nand g507 ( new_n722_, new_n721_, N146 );
nand g508 ( new_n723_, new_n425_, N17 );
nand g509 ( new_n724_, new_n723_, keyIn_0_18 );
not g510 ( new_n725_, keyIn_0_18 );
nand g511 ( new_n726_, new_n425_, new_n725_, N17 );
nand g512 ( new_n727_, new_n724_, new_n726_ );
nand g513 ( new_n728_, new_n727_, new_n437_ );
nand g514 ( new_n729_, N51, N138 );
nand g515 ( new_n730_, new_n713_, new_n722_, new_n728_, new_n729_ );
not g516 ( new_n731_, new_n730_ );
nand g517 ( new_n732_, new_n731_, new_n296_ );
nand g518 ( new_n733_, new_n596_, N101 );
nand g519 ( new_n734_, new_n721_, N149 );
nand g520 ( new_n735_, N17, N138 );
nand g521 ( new_n736_, new_n733_, new_n734_, new_n728_, new_n735_ );
not g522 ( new_n737_, new_n736_ );
nand g523 ( new_n738_, new_n737_, new_n300_ );
nand g524 ( new_n739_, new_n732_, new_n738_ );
not g525 ( new_n740_, new_n739_ );
not g526 ( new_n741_, keyIn_0_31 );
nand g527 ( new_n742_, new_n721_, N153 );
nand g528 ( new_n743_, new_n742_, keyIn_0_23 );
not g529 ( new_n744_, keyIn_0_23 );
nand g530 ( new_n745_, new_n721_, new_n744_, N153 );
nand g531 ( new_n746_, new_n743_, new_n745_ );
not g532 ( new_n747_, keyIn_0_24 );
nand g533 ( new_n748_, new_n728_, new_n747_ );
nand g534 ( new_n749_, new_n727_, keyIn_0_24, new_n437_ );
nand g535 ( new_n750_, new_n746_, new_n748_, new_n749_ );
nand g536 ( new_n751_, new_n750_, new_n741_ );
nand g537 ( new_n752_, new_n746_, keyIn_0_31, new_n748_, new_n749_ );
nand g538 ( new_n753_, new_n751_, new_n752_ );
not g539 ( new_n754_, keyIn_0_41 );
nand g540 ( new_n755_, new_n596_, keyIn_0_30, N106 );
nand g541 ( new_n756_, N138, N152 );
not g542 ( new_n757_, keyIn_0_30 );
nand g543 ( new_n758_, new_n596_, N106 );
nand g544 ( new_n759_, new_n758_, new_n757_ );
nand g545 ( new_n760_, new_n759_, new_n755_, new_n756_ );
nand g546 ( new_n761_, new_n760_, new_n754_ );
nand g547 ( new_n762_, new_n759_, keyIn_0_41, new_n755_, new_n756_ );
nand g548 ( new_n763_, new_n761_, new_n762_ );
nand g549 ( new_n764_, new_n753_, new_n763_ );
nand g550 ( new_n765_, new_n764_, keyIn_0_46 );
not g551 ( new_n766_, keyIn_0_46 );
nand g552 ( new_n767_, new_n753_, new_n763_, new_n766_ );
nand g553 ( new_n768_, new_n765_, new_n767_ );
not g554 ( new_n769_, new_n768_ );
nand g555 ( new_n770_, new_n769_, new_n301_ );
nand g556 ( new_n771_, new_n770_, keyIn_0_53 );
not g557 ( new_n772_, keyIn_0_53 );
nand g558 ( new_n773_, new_n769_, new_n772_, new_n301_ );
nand g559 ( new_n774_, new_n771_, new_n773_ );
not g560 ( new_n775_, new_n774_ );
not g561 ( new_n776_, keyIn_0_79 );
not g562 ( new_n777_, keyIn_0_78 );
nand g563 ( new_n778_, new_n585_, new_n589_, new_n627_ );
nand g564 ( new_n779_, new_n778_, new_n777_ );
nand g565 ( new_n780_, new_n585_, new_n589_, keyIn_0_78, new_n627_ );
nand g566 ( new_n781_, new_n779_, new_n780_ );
not g567 ( new_n782_, keyIn_0_70 );
nand g568 ( new_n783_, new_n655_, new_n782_ );
nand g569 ( new_n784_, new_n652_, keyIn_0_70, new_n654_ );
nand g570 ( new_n785_, new_n783_, new_n784_ );
not g571 ( new_n786_, new_n785_ );
nand g572 ( new_n787_, new_n781_, new_n786_ );
nand g573 ( new_n788_, new_n787_, new_n776_ );
nand g574 ( new_n789_, new_n781_, keyIn_0_79, new_n786_ );
nand g575 ( new_n790_, new_n788_, new_n740_, new_n775_, new_n789_ );
nand g576 ( new_n791_, new_n790_, keyIn_0_87 );
not g577 ( new_n792_, keyIn_0_87 );
not g578 ( new_n793_, new_n790_ );
nand g579 ( new_n794_, new_n793_, new_n792_ );
not g580 ( new_n795_, keyIn_0_63 );
not g581 ( new_n796_, keyIn_0_52 );
nand g582 ( new_n797_, new_n768_, N177 );
nand g583 ( new_n798_, new_n797_, new_n796_ );
nand g584 ( new_n799_, new_n768_, keyIn_0_52, N177 );
nand g585 ( new_n800_, new_n798_, new_n799_ );
nand g586 ( new_n801_, new_n800_, new_n795_ );
nand g587 ( new_n802_, new_n798_, keyIn_0_63, new_n799_ );
nand g588 ( new_n803_, new_n801_, new_n802_ );
nand g589 ( new_n804_, new_n803_, keyIn_0_74, new_n740_ );
not g590 ( new_n805_, keyIn_0_74 );
nand g591 ( new_n806_, new_n803_, new_n740_ );
nand g592 ( new_n807_, new_n806_, new_n805_ );
nor g593 ( new_n808_, new_n731_, new_n296_ );
not g594 ( new_n809_, new_n808_ );
nor g595 ( new_n810_, new_n737_, new_n300_ );
nand g596 ( new_n811_, new_n810_, new_n732_ );
nand g597 ( new_n812_, new_n807_, new_n804_, new_n809_, new_n811_ );
not g598 ( new_n813_, new_n812_ );
nand g599 ( new_n814_, new_n794_, new_n791_, new_n813_ );
nand g600 ( new_n815_, new_n814_, keyIn_0_88 );
not g601 ( new_n816_, keyIn_0_88 );
nand g602 ( new_n817_, new_n794_, new_n816_, new_n791_, new_n813_ );
nand g603 ( new_n818_, new_n815_, new_n817_ );
not g604 ( new_n819_, new_n818_ );
nand g605 ( new_n820_, new_n596_, N91 );
nand g606 ( new_n821_, N8, N138 );
nand g607 ( new_n822_, new_n820_, keyIn_0_40, new_n821_ );
not g608 ( new_n823_, keyIn_0_40 );
nand g609 ( new_n824_, new_n820_, new_n821_ );
nand g610 ( new_n825_, new_n824_, new_n823_ );
nand g611 ( new_n826_, new_n721_, N143 );
nand g612 ( new_n827_, new_n826_, new_n728_ );
not g613 ( new_n828_, new_n827_ );
nand g614 ( new_n829_, new_n825_, new_n295_, new_n822_, new_n828_ );
nand g615 ( new_n830_, new_n819_, keyIn_0_101, new_n829_ );
not g616 ( new_n831_, keyIn_0_51 );
nand g617 ( new_n832_, new_n825_, new_n822_, new_n828_ );
nand g618 ( new_n833_, new_n832_, N159 );
nand g619 ( new_n834_, new_n833_, new_n831_ );
nand g620 ( new_n835_, new_n832_, keyIn_0_51, N159 );
nand g621 ( new_n836_, new_n834_, new_n835_ );
not g622 ( new_n837_, keyIn_0_101 );
nand g623 ( new_n838_, new_n819_, new_n829_ );
nand g624 ( new_n839_, new_n838_, new_n837_ );
nand g625 ( new_n840_, new_n839_, new_n830_, new_n836_ );
nand g626 ( new_n841_, new_n840_, keyIn_0_107 );
not g627 ( new_n842_, keyIn_0_107 );
nand g628 ( new_n843_, new_n839_, new_n842_, new_n830_, new_n836_ );
nand g629 ( new_n844_, new_n841_, new_n843_ );
nand g630 ( new_n845_, new_n844_, keyIn_0_113 );
not g631 ( new_n846_, keyIn_0_113 );
nand g632 ( new_n847_, new_n841_, new_n846_, new_n843_ );
nand g633 ( new_n848_, new_n845_, new_n847_ );
not g634 ( N866, new_n848_ );
not g635 ( new_n850_, keyIn_0_121 );
not g636 ( new_n851_, keyIn_0_117 );
not g637 ( new_n852_, keyIn_0_82 );
nand g638 ( new_n853_, new_n788_, new_n789_ );
not g639 ( new_n854_, new_n853_ );
nor g640 ( new_n855_, new_n774_, new_n800_ );
nand g641 ( new_n856_, new_n854_, new_n855_ );
nand g642 ( new_n857_, new_n856_, new_n852_ );
nand g643 ( new_n858_, new_n854_, keyIn_0_82, new_n855_ );
nand g644 ( new_n859_, new_n857_, new_n858_ );
not g645 ( new_n860_, new_n855_ );
nand g646 ( new_n861_, new_n853_, new_n860_ );
nand g647 ( new_n862_, new_n861_, keyIn_0_81 );
not g648 ( new_n863_, keyIn_0_81 );
nand g649 ( new_n864_, new_n853_, new_n863_, new_n860_ );
nand g650 ( new_n865_, new_n862_, new_n864_ );
nand g651 ( new_n866_, new_n859_, keyIn_0_91, new_n865_ );
not g652 ( new_n867_, keyIn_0_91 );
nand g653 ( new_n868_, new_n859_, new_n865_ );
nand g654 ( new_n869_, new_n868_, new_n867_ );
nand g655 ( new_n870_, new_n869_, keyIn_0_99, N219, new_n866_ );
nand g656 ( new_n871_, N101, N210 );
not g657 ( new_n872_, keyIn_0_99 );
nand g658 ( new_n873_, new_n869_, N219, new_n866_ );
nand g659 ( new_n874_, new_n873_, new_n872_ );
nand g660 ( new_n875_, new_n874_, new_n870_, new_n871_ );
nand g661 ( new_n876_, new_n875_, keyIn_0_105 );
not g662 ( new_n877_, keyIn_0_105 );
nand g663 ( new_n878_, new_n874_, new_n877_, new_n870_, new_n871_ );
nand g664 ( new_n879_, new_n876_, new_n878_ );
not g665 ( new_n880_, keyIn_0_69 );
nand g666 ( new_n881_, new_n803_, new_n880_, N237 );
nand g667 ( new_n882_, new_n803_, N237 );
nand g668 ( new_n883_, new_n882_, keyIn_0_69 );
nand g669 ( new_n884_, new_n855_, N228 );
nand g670 ( new_n885_, new_n768_, N246 );
nand g671 ( new_n886_, new_n476_, N177 );
nand g672 ( new_n887_, new_n885_, new_n886_ );
not g673 ( new_n888_, new_n887_ );
nand g674 ( new_n889_, new_n883_, new_n881_, new_n884_, new_n888_ );
not g675 ( new_n890_, new_n889_ );
nand g676 ( new_n891_, new_n879_, new_n890_ );
nand g677 ( new_n892_, new_n891_, keyIn_0_111 );
not g678 ( new_n893_, keyIn_0_111 );
nand g679 ( new_n894_, new_n879_, new_n893_, new_n890_ );
nand g680 ( new_n895_, new_n892_, new_n894_ );
nand g681 ( new_n896_, new_n895_, new_n851_ );
nand g682 ( new_n897_, new_n892_, keyIn_0_117, new_n894_ );
nand g683 ( new_n898_, new_n896_, new_n897_ );
nand g684 ( new_n899_, new_n898_, new_n850_ );
nand g685 ( new_n900_, new_n896_, keyIn_0_121, new_n897_ );
nand g686 ( new_n901_, new_n899_, new_n900_ );
not g687 ( N874, new_n901_ );
not g688 ( new_n903_, keyIn_0_102 );
not g689 ( new_n904_, keyIn_0_62 );
nand g690 ( new_n905_, new_n836_, new_n829_ );
nand g691 ( new_n906_, new_n905_, new_n904_ );
nand g692 ( new_n907_, new_n836_, keyIn_0_62, new_n829_ );
nand g693 ( new_n908_, new_n906_, new_n907_ );
not g694 ( new_n909_, new_n908_ );
nand g695 ( new_n910_, new_n818_, new_n909_ );
nand g696 ( new_n911_, new_n910_, keyIn_0_93 );
not g697 ( new_n912_, keyIn_0_93 );
nand g698 ( new_n913_, new_n818_, new_n912_, new_n909_ );
nand g699 ( new_n914_, new_n911_, new_n913_ );
not g700 ( new_n915_, keyIn_0_94 );
nand g701 ( new_n916_, new_n815_, new_n817_, new_n908_ );
nand g702 ( new_n917_, new_n916_, new_n915_ );
nand g703 ( new_n918_, new_n815_, keyIn_0_94, new_n817_, new_n908_ );
nand g704 ( new_n919_, new_n917_, new_n918_ );
not g705 ( new_n920_, new_n919_ );
nand g706 ( new_n921_, new_n920_, new_n914_ );
nand g707 ( new_n922_, new_n921_, new_n903_ );
nand g708 ( new_n923_, new_n920_, new_n914_, keyIn_0_102 );
nand g709 ( new_n924_, new_n922_, keyIn_0_108, N219, new_n923_ );
nand g710 ( new_n925_, new_n440_, N210 );
not g711 ( new_n926_, keyIn_0_108 );
nand g712 ( new_n927_, new_n922_, N219, new_n923_ );
nand g713 ( new_n928_, new_n927_, new_n926_ );
nand g714 ( new_n929_, new_n928_, new_n924_, new_n925_ );
nand g715 ( new_n930_, new_n929_, keyIn_0_114 );
not g716 ( new_n931_, keyIn_0_114 );
nand g717 ( new_n932_, new_n928_, new_n931_, new_n924_, new_n925_ );
nand g718 ( new_n933_, new_n930_, new_n932_ );
nand g719 ( new_n934_, new_n908_, N228 );
nand g720 ( new_n935_, new_n834_, N237, new_n835_ );
nand g721 ( new_n936_, new_n476_, N159 );
nand g722 ( new_n937_, new_n832_, N246 );
nand g723 ( new_n938_, new_n934_, new_n935_, new_n936_, new_n937_ );
not g724 ( new_n939_, new_n938_ );
nand g725 ( new_n940_, new_n933_, new_n939_ );
nand g726 ( new_n941_, new_n940_, keyIn_0_118 );
not g727 ( new_n942_, keyIn_0_118 );
nand g728 ( new_n943_, new_n933_, new_n942_, new_n939_ );
nand g729 ( new_n944_, new_n941_, new_n943_ );
nand g730 ( new_n945_, new_n944_, keyIn_0_122 );
not g731 ( new_n946_, keyIn_0_122 );
nand g732 ( new_n947_, new_n941_, new_n946_, new_n943_ );
nand g733 ( new_n948_, new_n945_, new_n947_ );
nand g734 ( new_n949_, new_n948_, keyIn_0_125 );
not g735 ( new_n950_, keyIn_0_125 );
nand g736 ( new_n951_, new_n945_, new_n950_, new_n947_ );
nand g737 ( new_n952_, new_n949_, new_n951_ );
not g738 ( N878, new_n952_ );
not g739 ( new_n954_, keyIn_0_126 );
not g740 ( new_n955_, keyIn_0_123 );
not g741 ( new_n956_, keyIn_0_119 );
not g742 ( new_n957_, keyIn_0_115 );
not g743 ( new_n958_, keyIn_0_103 );
nand g744 ( new_n959_, new_n809_, new_n732_ );
not g745 ( new_n960_, keyIn_0_89 );
not g746 ( new_n961_, keyIn_0_86 );
nand g747 ( new_n962_, new_n788_, new_n775_, new_n789_ );
not g748 ( new_n963_, new_n962_ );
nand g749 ( new_n964_, new_n963_, new_n961_, new_n738_ );
nand g750 ( new_n965_, new_n963_, new_n738_ );
nand g751 ( new_n966_, new_n965_, keyIn_0_86 );
not g752 ( new_n967_, new_n810_ );
nand g753 ( new_n968_, new_n803_, new_n738_ );
nand g754 ( new_n969_, new_n968_, new_n967_ );
not g755 ( new_n970_, new_n969_ );
nand g756 ( new_n971_, new_n966_, new_n964_, new_n970_ );
nand g757 ( new_n972_, new_n971_, new_n960_ );
nand g758 ( new_n973_, new_n966_, keyIn_0_89, new_n964_, new_n970_ );
nand g759 ( new_n974_, new_n972_, new_n973_ );
nand g760 ( new_n975_, new_n974_, keyIn_0_95, new_n959_ );
not g761 ( new_n976_, keyIn_0_96 );
not g762 ( new_n977_, new_n959_ );
nand g763 ( new_n978_, new_n972_, new_n976_, new_n977_, new_n973_ );
nand g764 ( new_n979_, new_n972_, new_n977_, new_n973_ );
nand g765 ( new_n980_, new_n979_, keyIn_0_96 );
not g766 ( new_n981_, keyIn_0_95 );
nand g767 ( new_n982_, new_n974_, new_n959_ );
nand g768 ( new_n983_, new_n982_, new_n981_ );
nand g769 ( new_n984_, new_n983_, new_n975_, new_n978_, new_n980_ );
nand g770 ( new_n985_, new_n984_, new_n958_ );
nand g771 ( new_n986_, new_n975_, new_n978_ );
not g772 ( new_n987_, new_n986_ );
nand g773 ( new_n988_, new_n987_, keyIn_0_103, new_n980_, new_n983_ );
nand g774 ( new_n989_, new_n988_, new_n985_ );
nand g775 ( new_n990_, new_n989_, keyIn_0_109, N219 );
nand g776 ( new_n991_, N91, N210 );
not g777 ( new_n992_, keyIn_0_109 );
nand g778 ( new_n993_, new_n989_, N219 );
nand g779 ( new_n994_, new_n993_, new_n992_ );
nand g780 ( new_n995_, new_n994_, new_n957_, new_n990_, new_n991_ );
nand g781 ( new_n996_, new_n994_, new_n990_, new_n991_ );
nand g782 ( new_n997_, new_n996_, keyIn_0_115 );
nand g783 ( new_n998_, new_n977_, N228 );
not g784 ( new_n999_, new_n998_ );
nand g785 ( new_n1000_, new_n808_, N237 );
nand g786 ( new_n1001_, new_n476_, N165 );
nand g787 ( new_n1002_, new_n730_, N246 );
nand g788 ( new_n1003_, new_n1000_, new_n1001_, new_n1002_ );
nor g789 ( new_n1004_, new_n999_, new_n1003_ );
nand g790 ( new_n1005_, new_n997_, new_n995_, new_n1004_ );
nand g791 ( new_n1006_, new_n1005_, new_n956_ );
nand g792 ( new_n1007_, new_n997_, keyIn_0_119, new_n995_, new_n1004_ );
nand g793 ( new_n1008_, new_n1006_, new_n1007_ );
nand g794 ( new_n1009_, new_n1008_, new_n955_ );
nand g795 ( new_n1010_, new_n1006_, keyIn_0_123, new_n1007_ );
nand g796 ( new_n1011_, new_n1009_, new_n1010_ );
nand g797 ( new_n1012_, new_n1011_, new_n954_ );
nand g798 ( new_n1013_, new_n1009_, keyIn_0_126, new_n1010_ );
nand g799 ( N879, new_n1012_, new_n1013_ );
not g800 ( new_n1015_, keyIn_0_110 );
not g801 ( new_n1016_, keyIn_0_104 );
not g802 ( new_n1017_, keyIn_0_90 );
not g803 ( new_n1018_, new_n803_ );
nand g804 ( new_n1019_, new_n963_, keyIn_0_85 );
not g805 ( new_n1020_, keyIn_0_85 );
nand g806 ( new_n1021_, new_n962_, new_n1020_ );
nand g807 ( new_n1022_, new_n1019_, new_n1018_, new_n1021_ );
nand g808 ( new_n1023_, new_n1022_, new_n1017_ );
nand g809 ( new_n1024_, new_n1019_, keyIn_0_90, new_n1018_, new_n1021_ );
nand g810 ( new_n1025_, new_n967_, new_n738_ );
nand g811 ( new_n1026_, new_n1023_, new_n1024_, new_n1025_ );
nand g812 ( new_n1027_, new_n1026_, keyIn_0_97 );
nand g813 ( new_n1028_, new_n1023_, new_n1024_ );
not g814 ( new_n1029_, new_n1025_ );
nand g815 ( new_n1030_, new_n1028_, new_n1029_ );
nand g816 ( new_n1031_, new_n1030_, keyIn_0_98 );
not g817 ( new_n1032_, keyIn_0_97 );
nand g818 ( new_n1033_, new_n1023_, new_n1032_, new_n1024_, new_n1025_ );
not g819 ( new_n1034_, keyIn_0_98 );
nand g820 ( new_n1035_, new_n1028_, new_n1034_, new_n1029_ );
nand g821 ( new_n1036_, new_n1035_, new_n1033_ );
not g822 ( new_n1037_, new_n1036_ );
nand g823 ( new_n1038_, new_n1037_, new_n1016_, new_n1027_, new_n1031_ );
nand g824 ( new_n1039_, new_n1031_, new_n1027_, new_n1033_, new_n1035_ );
nand g825 ( new_n1040_, new_n1039_, keyIn_0_104 );
nand g826 ( new_n1041_, new_n1038_, new_n1040_, new_n1015_, N219 );
nand g827 ( new_n1042_, N96, N210 );
nand g828 ( new_n1043_, new_n1038_, new_n1040_, N219 );
nand g829 ( new_n1044_, new_n1043_, keyIn_0_110 );
nand g830 ( new_n1045_, new_n1044_, new_n1041_, new_n1042_ );
nand g831 ( new_n1046_, new_n1045_, keyIn_0_116 );
not g832 ( new_n1047_, keyIn_0_116 );
nand g833 ( new_n1048_, new_n1044_, new_n1047_, new_n1041_, new_n1042_ );
nand g834 ( new_n1049_, new_n1046_, new_n1048_ );
nand g835 ( new_n1050_, new_n1029_, N228 );
not g836 ( new_n1051_, new_n1050_ );
nand g837 ( new_n1052_, new_n810_, N237 );
nand g838 ( new_n1053_, new_n476_, N171 );
nand g839 ( new_n1054_, new_n736_, N246 );
nand g840 ( new_n1055_, new_n1052_, new_n1053_, new_n1054_ );
nor g841 ( new_n1056_, new_n1051_, new_n1055_ );
nand g842 ( new_n1057_, new_n1049_, new_n1056_ );
nand g843 ( new_n1058_, new_n1057_, keyIn_0_120 );
not g844 ( new_n1059_, keyIn_0_120 );
nand g845 ( new_n1060_, new_n1049_, new_n1059_, new_n1056_ );
nand g846 ( new_n1061_, new_n1058_, new_n1060_ );
nand g847 ( new_n1062_, new_n1061_, keyIn_0_124 );
not g848 ( new_n1063_, keyIn_0_124 );
nand g849 ( new_n1064_, new_n1058_, new_n1063_, new_n1060_ );
nand g850 ( new_n1065_, new_n1062_, new_n1064_ );
nand g851 ( new_n1066_, new_n1065_, keyIn_0_127 );
not g852 ( new_n1067_, keyIn_0_127 );
nand g853 ( new_n1068_, new_n1062_, new_n1067_, new_n1064_ );
nand g854 ( new_n1069_, new_n1066_, new_n1068_ );
not g855 ( N880, new_n1069_ );
endmodule