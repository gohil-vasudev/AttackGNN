module add_mul_sub_32_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, 
        a_18_, a_19_, a_20_, a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, 
        a_28_, a_29_, a_30_, a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, 
        b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, 
        b_17_, b_18_, b_19_, b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, 
        b_27_, b_28_, b_29_, b_30_, b_31_, operation_0_, operation_1_, 
        Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_, 
        Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_, 
        Result_12_, Result_13_, Result_14_, Result_15_, Result_16_, Result_17_, 
        Result_18_, Result_19_, Result_20_, Result_21_, Result_22_, Result_23_, 
        Result_24_, Result_25_, Result_26_, Result_27_, Result_28_, Result_29_, 
        Result_30_, Result_31_, Result_32_, Result_33_, Result_34_, Result_35_, 
        Result_36_, Result_37_, Result_38_, Result_39_, Result_40_, Result_41_, 
        Result_42_, Result_43_, Result_44_, Result_45_, Result_46_, Result_47_, 
        Result_48_, Result_49_, Result_50_, Result_51_, Result_52_, Result_53_, 
        Result_54_, Result_55_, Result_56_, Result_57_, Result_58_, Result_59_, 
        Result_60_, Result_61_, Result_62_, Result_63_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, a_19_, a_20_,
         a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, a_29_, a_30_,
         a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_,
         b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, b_18_, b_19_,
         b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, b_28_, b_29_,
         b_30_, b_31_, operation_0_, operation_1_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_,
         Result_32_, Result_33_, Result_34_, Result_35_, Result_36_,
         Result_37_, Result_38_, Result_39_, Result_40_, Result_41_,
         Result_42_, Result_43_, Result_44_, Result_45_, Result_46_,
         Result_47_, Result_48_, Result_49_, Result_50_, Result_51_,
         Result_52_, Result_53_, Result_54_, Result_55_, Result_56_,
         Result_57_, Result_58_, Result_59_, Result_60_, Result_61_,
         Result_62_, Result_63_;
  wire   n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000;

  OR2_X1 U7877 ( .A1(n15634), .A2(n7867), .ZN(n7813) );
  OR2_X1 U7878 ( .A1(n15811), .A2(n15812), .ZN(n7814) );
  OR2_X1 U7879 ( .A1(n15812), .A2(operation_0_), .ZN(n7815) );
  OR2_X1 U7880 ( .A1(n15811), .A2(operation_1_), .ZN(n7816) );
  OR2_X1 U7881 ( .A1(operation_0_), .A2(operation_1_), .ZN(n7817) );
  AND2_X2 U7882 ( .A1(n15813), .A2(n15814), .ZN(n7823) );
  INV_X1 U7883 ( .A(n7813), .ZN(n7818) );
  INV_X4 U7884 ( .A(n7817), .ZN(n7819) );
  INV_X4 U7885 ( .A(n7816), .ZN(n7820) );
  INV_X4 U7886 ( .A(n7814), .ZN(n7821) );
  INV_X4 U7887 ( .A(n7815), .ZN(n7822) );
  INV_X2 U7888 ( .A(b_14_), .ZN(n8301) );
  INV_X2 U7889 ( .A(b_26_), .ZN(n7992) );
  INV_X2 U7890 ( .A(b_7_), .ZN(n8482) );
  INV_X2 U7891 ( .A(b_30_), .ZN(n7869) );
  INV_X2 U7892 ( .A(b_6_), .ZN(n8508) );
  INV_X2 U7893 ( .A(b_16_), .ZN(n8251) );
  INV_X2 U7894 ( .A(b_0_), .ZN(n8770) );
  INV_X2 U7895 ( .A(b_4_), .ZN(n8558) );
  INV_X2 U7896 ( .A(b_28_), .ZN(n7935) );
  INV_X2 U7897 ( .A(b_22_), .ZN(n8094) );
  INV_X2 U7898 ( .A(a_15_), .ZN(n8276) );
  INV_X2 U7899 ( .A(a_13_), .ZN(n8310) );
  INV_X2 U7900 ( .A(a_1_), .ZN(n8617) );
  INV_X2 U7901 ( .A(a_23_), .ZN(n8747) );
  INV_X2 U7902 ( .A(a_19_), .ZN(n8170) );
  INV_X2 U7903 ( .A(a_25_), .ZN(n8744) );
  INV_X2 U7904 ( .A(a_20_), .ZN(n8751) );
  NAND2_X2 U7905 ( .A1(a_30_), .A2(n15634), .ZN(n9137) );
  INV_X2 U7906 ( .A(a_18_), .ZN(n8753) );
  INV_X2 U7907 ( .A(a_24_), .ZN(n8745) );
  NAND2_X2 U7908 ( .A1(a_31_), .A2(n7867), .ZN(n7864) );
  INV_X2 U7909 ( .A(a_21_), .ZN(n8750) );
  INV_X2 U7910 ( .A(a_17_), .ZN(n8210) );
  INV_X2 U7911 ( .A(a_29_), .ZN(n7890) );
  NAND2_X1 U7912 ( .A1(n7823), .A2(n7824), .ZN(Result_9_) );
  NAND2_X1 U7913 ( .A1(n7825), .A2(n7821), .ZN(n7824) );
  XOR2_X1 U7914 ( .A(n7826), .B(n7827), .Z(n7825) );
  AND2_X1 U7915 ( .A1(n7828), .A2(n7829), .ZN(n7827) );
  NAND2_X1 U7916 ( .A1(n7823), .A2(n7830), .ZN(Result_8_) );
  NAND2_X1 U7917 ( .A1(n7831), .A2(n7821), .ZN(n7830) );
  XOR2_X1 U7918 ( .A(n7832), .B(n7833), .Z(n7831) );
  AND2_X1 U7919 ( .A1(n7834), .A2(n7835), .ZN(n7833) );
  NAND2_X1 U7920 ( .A1(n7823), .A2(n7836), .ZN(Result_7_) );
  NAND2_X1 U7921 ( .A1(n7837), .A2(n7821), .ZN(n7836) );
  XOR2_X1 U7922 ( .A(n7838), .B(n7839), .Z(n7837) );
  AND2_X1 U7923 ( .A1(n7840), .A2(n7841), .ZN(n7839) );
  NAND2_X1 U7924 ( .A1(n7823), .A2(n7842), .ZN(Result_6_) );
  NAND2_X1 U7925 ( .A1(n7843), .A2(n7821), .ZN(n7842) );
  XOR2_X1 U7926 ( .A(n7844), .B(n7845), .Z(n7843) );
  AND2_X1 U7927 ( .A1(n7846), .A2(n7847), .ZN(n7845) );
  NAND2_X1 U7928 ( .A1(n7848), .A2(n7849), .ZN(Result_63_) );
  NAND2_X1 U7929 ( .A1(n7850), .A2(n7821), .ZN(n7849) );
  NAND2_X1 U7930 ( .A1(n7851), .A2(n7852), .ZN(n7848) );
  OR3_X1 U7931 ( .A1(n7822), .A2(n7820), .A3(n7819), .ZN(n7852) );
  NAND2_X1 U7932 ( .A1(n7853), .A2(n7854), .ZN(n7851) );
  NAND3_X1 U7933 ( .A1(n7855), .A2(n7856), .A3(n7857), .ZN(Result_62_) );
  NAND3_X1 U7934 ( .A1(a_30_), .A2(n7858), .A3(n7821), .ZN(n7857) );
  NAND2_X1 U7935 ( .A1(b_30_), .A2(n7859), .ZN(n7856) );
  NAND3_X1 U7936 ( .A1(n7860), .A2(n7861), .A3(n7862), .ZN(n7859) );
  NAND2_X1 U7937 ( .A1(n7821), .A2(n7863), .ZN(n7862) );
  NAND2_X1 U7938 ( .A1(n7854), .A2(n7864), .ZN(n7863) );
  NAND2_X1 U7939 ( .A1(a_30_), .A2(n7865), .ZN(n7861) );
  NAND2_X1 U7940 ( .A1(n7866), .A2(n7867), .ZN(n7860) );
  NAND2_X1 U7941 ( .A1(n7868), .A2(n7869), .ZN(n7855) );
  NAND2_X1 U7942 ( .A1(n7870), .A2(n7871), .ZN(n7868) );
  NAND2_X1 U7943 ( .A1(n7865), .A2(n7867), .ZN(n7871) );
  NAND3_X1 U7944 ( .A1(n7872), .A2(n7873), .A3(n7874), .ZN(n7865) );
  NAND2_X1 U7945 ( .A1(n7820), .A2(n7875), .ZN(n7874) );
  NAND2_X1 U7946 ( .A1(n7819), .A2(n7850), .ZN(n7873) );
  INV_X1 U7947 ( .A(n7876), .ZN(n7850) );
  NAND2_X1 U7948 ( .A1(n7822), .A2(n7858), .ZN(n7872) );
  NAND2_X1 U7949 ( .A1(a_30_), .A2(n7877), .ZN(n7870) );
  NAND2_X1 U7950 ( .A1(n7878), .A2(n7879), .ZN(n7877) );
  NAND2_X1 U7951 ( .A1(n7821), .A2(b_31_), .ZN(n7879) );
  INV_X1 U7952 ( .A(n7866), .ZN(n7878) );
  NAND3_X1 U7953 ( .A1(n7880), .A2(n7881), .A3(n7882), .ZN(n7866) );
  NAND2_X1 U7954 ( .A1(n7820), .A2(n7854), .ZN(n7882) );
  NAND2_X1 U7955 ( .A1(n7819), .A2(n7876), .ZN(n7881) );
  NAND2_X1 U7956 ( .A1(n7822), .A2(n7853), .ZN(n7880) );
  NAND3_X1 U7957 ( .A1(n7883), .A2(n7884), .A3(n7885), .ZN(Result_61_) );
  NAND2_X1 U7958 ( .A1(n7886), .A2(n7821), .ZN(n7885) );
  XOR2_X1 U7959 ( .A(n7887), .B(n7888), .Z(n7886) );
  NOR2_X1 U7960 ( .A1(n7889), .A2(n7890), .ZN(n7888) );
  XOR2_X1 U7961 ( .A(n7891), .B(n7892), .Z(n7887) );
  NAND2_X1 U7962 ( .A1(n7893), .A2(n7894), .ZN(n7884) );
  NAND3_X1 U7963 ( .A1(n7895), .A2(n7896), .A3(n7897), .ZN(n7893) );
  NAND2_X1 U7964 ( .A1(n7820), .A2(n7898), .ZN(n7897) );
  NAND2_X1 U7965 ( .A1(n7819), .A2(n7899), .ZN(n7896) );
  NAND2_X1 U7966 ( .A1(n7822), .A2(n7900), .ZN(n7895) );
  NAND2_X1 U7967 ( .A1(n7901), .A2(n7902), .ZN(n7883) );
  NAND3_X1 U7968 ( .A1(n7903), .A2(n7904), .A3(n7905), .ZN(n7902) );
  NAND2_X1 U7969 ( .A1(n7820), .A2(n7906), .ZN(n7905) );
  NAND2_X1 U7970 ( .A1(n7907), .A2(n7819), .ZN(n7904) );
  INV_X1 U7971 ( .A(n7899), .ZN(n7907) );
  NAND2_X1 U7972 ( .A1(n7822), .A2(n7908), .ZN(n7903) );
  INV_X1 U7973 ( .A(n7894), .ZN(n7901) );
  NAND2_X1 U7974 ( .A1(n7909), .A2(n7910), .ZN(n7894) );
  NAND3_X1 U7975 ( .A1(n7911), .A2(n7912), .A3(n7913), .ZN(Result_60_) );
  NAND2_X1 U7976 ( .A1(n7821), .A2(n7914), .ZN(n7913) );
  XOR2_X1 U7977 ( .A(n7915), .B(n7916), .Z(n7914) );
  XOR2_X1 U7978 ( .A(n7917), .B(n7918), .Z(n7916) );
  NAND2_X1 U7979 ( .A1(n7919), .A2(n7920), .ZN(n7912) );
  NAND3_X1 U7980 ( .A1(n7921), .A2(n7922), .A3(n7923), .ZN(n7920) );
  NAND2_X1 U7981 ( .A1(n7820), .A2(n7924), .ZN(n7923) );
  NAND2_X1 U7982 ( .A1(n7925), .A2(n7819), .ZN(n7922) );
  INV_X1 U7983 ( .A(n7926), .ZN(n7925) );
  NAND2_X1 U7984 ( .A1(n7822), .A2(n7927), .ZN(n7921) );
  NAND2_X1 U7985 ( .A1(n7928), .A2(n7929), .ZN(n7911) );
  NAND3_X1 U7986 ( .A1(n7930), .A2(n7931), .A3(n7932), .ZN(n7929) );
  NAND2_X1 U7987 ( .A1(n7820), .A2(n7933), .ZN(n7932) );
  NAND2_X1 U7988 ( .A1(n7819), .A2(n7926), .ZN(n7931) );
  NAND2_X1 U7989 ( .A1(n7822), .A2(n7934), .ZN(n7930) );
  INV_X1 U7990 ( .A(n7919), .ZN(n7928) );
  XNOR2_X1 U7991 ( .A(n7935), .B(a_28_), .ZN(n7919) );
  NAND2_X1 U7992 ( .A1(n7823), .A2(n7936), .ZN(Result_5_) );
  NAND2_X1 U7993 ( .A1(n7937), .A2(n7821), .ZN(n7936) );
  XOR2_X1 U7994 ( .A(n7938), .B(n7939), .Z(n7937) );
  AND2_X1 U7995 ( .A1(n7940), .A2(n7941), .ZN(n7939) );
  NAND3_X1 U7996 ( .A1(n7942), .A2(n7943), .A3(n7944), .ZN(Result_59_) );
  NAND2_X1 U7997 ( .A1(n7821), .A2(n7945), .ZN(n7944) );
  XNOR2_X1 U7998 ( .A(n7946), .B(n7947), .ZN(n7945) );
  NAND2_X1 U7999 ( .A1(n7948), .A2(n7949), .ZN(n7946) );
  NAND2_X1 U8000 ( .A1(n7950), .A2(n7951), .ZN(n7943) );
  NAND3_X1 U8001 ( .A1(n7952), .A2(n7953), .A3(n7954), .ZN(n7950) );
  NAND2_X1 U8002 ( .A1(n7820), .A2(n7955), .ZN(n7954) );
  NAND2_X1 U8003 ( .A1(n7819), .A2(n7956), .ZN(n7953) );
  NAND2_X1 U8004 ( .A1(n7822), .A2(n7957), .ZN(n7952) );
  NAND2_X1 U8005 ( .A1(n7958), .A2(n7959), .ZN(n7942) );
  NAND3_X1 U8006 ( .A1(n7960), .A2(n7961), .A3(n7962), .ZN(n7959) );
  NAND2_X1 U8007 ( .A1(n7820), .A2(n7963), .ZN(n7962) );
  NAND2_X1 U8008 ( .A1(n7964), .A2(n7819), .ZN(n7961) );
  INV_X1 U8009 ( .A(n7956), .ZN(n7964) );
  NAND2_X1 U8010 ( .A1(n7822), .A2(n7965), .ZN(n7960) );
  INV_X1 U8011 ( .A(n7951), .ZN(n7958) );
  NAND2_X1 U8012 ( .A1(n7966), .A2(n7967), .ZN(n7951) );
  NAND3_X1 U8013 ( .A1(n7968), .A2(n7969), .A3(n7970), .ZN(Result_58_) );
  NAND2_X1 U8014 ( .A1(n7971), .A2(n7821), .ZN(n7970) );
  XOR2_X1 U8015 ( .A(n7972), .B(n7973), .Z(n7971) );
  XOR2_X1 U8016 ( .A(n7974), .B(n7975), .Z(n7972) );
  NAND2_X1 U8017 ( .A1(n7976), .A2(n7977), .ZN(n7969) );
  NAND3_X1 U8018 ( .A1(n7978), .A2(n7979), .A3(n7980), .ZN(n7977) );
  NAND2_X1 U8019 ( .A1(n7820), .A2(n7981), .ZN(n7980) );
  NAND2_X1 U8020 ( .A1(n7982), .A2(n7819), .ZN(n7979) );
  INV_X1 U8021 ( .A(n7983), .ZN(n7982) );
  NAND2_X1 U8022 ( .A1(n7822), .A2(n7984), .ZN(n7978) );
  NAND2_X1 U8023 ( .A1(n7985), .A2(n7986), .ZN(n7968) );
  NAND3_X1 U8024 ( .A1(n7987), .A2(n7988), .A3(n7989), .ZN(n7986) );
  NAND2_X1 U8025 ( .A1(n7820), .A2(n7990), .ZN(n7989) );
  NAND2_X1 U8026 ( .A1(n7819), .A2(n7983), .ZN(n7988) );
  NAND2_X1 U8027 ( .A1(n7822), .A2(n7991), .ZN(n7987) );
  INV_X1 U8028 ( .A(n7976), .ZN(n7985) );
  XNOR2_X1 U8029 ( .A(n7992), .B(a_26_), .ZN(n7976) );
  NAND3_X1 U8030 ( .A1(n7993), .A2(n7994), .A3(n7995), .ZN(Result_57_) );
  NAND2_X1 U8031 ( .A1(n7821), .A2(n7996), .ZN(n7995) );
  XNOR2_X1 U8032 ( .A(n7997), .B(n7998), .ZN(n7996) );
  NAND2_X1 U8033 ( .A1(n7999), .A2(n8000), .ZN(n7997) );
  NAND2_X1 U8034 ( .A1(n8001), .A2(n8002), .ZN(n7994) );
  NAND3_X1 U8035 ( .A1(n8003), .A2(n8004), .A3(n8005), .ZN(n8001) );
  NAND2_X1 U8036 ( .A1(n7820), .A2(n8006), .ZN(n8005) );
  NAND2_X1 U8037 ( .A1(n7819), .A2(n8007), .ZN(n8004) );
  NAND2_X1 U8038 ( .A1(n7822), .A2(n8008), .ZN(n8003) );
  NAND2_X1 U8039 ( .A1(n8009), .A2(n8010), .ZN(n7993) );
  NAND3_X1 U8040 ( .A1(n8011), .A2(n8012), .A3(n8013), .ZN(n8010) );
  NAND2_X1 U8041 ( .A1(n7820), .A2(n8014), .ZN(n8013) );
  NAND2_X1 U8042 ( .A1(n8015), .A2(n7819), .ZN(n8012) );
  INV_X1 U8043 ( .A(n8007), .ZN(n8015) );
  NAND2_X1 U8044 ( .A1(n7822), .A2(n8016), .ZN(n8011) );
  INV_X1 U8045 ( .A(n8002), .ZN(n8009) );
  NAND2_X1 U8046 ( .A1(n8017), .A2(n8018), .ZN(n8002) );
  NAND3_X1 U8047 ( .A1(n8019), .A2(n8020), .A3(n8021), .ZN(Result_56_) );
  NAND2_X1 U8048 ( .A1(n7821), .A2(n8022), .ZN(n8021) );
  XNOR2_X1 U8049 ( .A(n8023), .B(n8024), .ZN(n8022) );
  XNOR2_X1 U8050 ( .A(n8025), .B(n8026), .ZN(n8024) );
  NAND2_X1 U8051 ( .A1(n8027), .A2(n8028), .ZN(n8020) );
  NAND3_X1 U8052 ( .A1(n8029), .A2(n8030), .A3(n8031), .ZN(n8028) );
  NAND2_X1 U8053 ( .A1(n7820), .A2(n8032), .ZN(n8031) );
  NAND2_X1 U8054 ( .A1(n8033), .A2(n7819), .ZN(n8030) );
  INV_X1 U8055 ( .A(n8034), .ZN(n8033) );
  NAND2_X1 U8056 ( .A1(n7822), .A2(n8035), .ZN(n8029) );
  NAND2_X1 U8057 ( .A1(n8036), .A2(n8037), .ZN(n8019) );
  NAND3_X1 U8058 ( .A1(n8038), .A2(n8039), .A3(n8040), .ZN(n8037) );
  NAND2_X1 U8059 ( .A1(n7820), .A2(n8041), .ZN(n8040) );
  NAND2_X1 U8060 ( .A1(n7819), .A2(n8034), .ZN(n8039) );
  NAND2_X1 U8061 ( .A1(n7822), .A2(n8042), .ZN(n8038) );
  INV_X1 U8062 ( .A(n8027), .ZN(n8036) );
  XNOR2_X1 U8063 ( .A(n8043), .B(a_24_), .ZN(n8027) );
  NAND3_X1 U8064 ( .A1(n8044), .A2(n8045), .A3(n8046), .ZN(Result_55_) );
  NAND2_X1 U8065 ( .A1(n8047), .A2(n7821), .ZN(n8046) );
  XNOR2_X1 U8066 ( .A(n8048), .B(n8049), .ZN(n8047) );
  NAND2_X1 U8067 ( .A1(n8050), .A2(n8051), .ZN(n8048) );
  NAND2_X1 U8068 ( .A1(n8052), .A2(n8053), .ZN(n8045) );
  NAND3_X1 U8069 ( .A1(n8054), .A2(n8055), .A3(n8056), .ZN(n8052) );
  NAND2_X1 U8070 ( .A1(n7820), .A2(n8057), .ZN(n8056) );
  NAND2_X1 U8071 ( .A1(n7819), .A2(n8058), .ZN(n8055) );
  NAND2_X1 U8072 ( .A1(n7822), .A2(n8059), .ZN(n8054) );
  NAND2_X1 U8073 ( .A1(n8060), .A2(n8061), .ZN(n8044) );
  NAND3_X1 U8074 ( .A1(n8062), .A2(n8063), .A3(n8064), .ZN(n8061) );
  NAND2_X1 U8075 ( .A1(n7820), .A2(n8065), .ZN(n8064) );
  NAND2_X1 U8076 ( .A1(n8066), .A2(n7819), .ZN(n8063) );
  INV_X1 U8077 ( .A(n8058), .ZN(n8066) );
  NAND2_X1 U8078 ( .A1(n7822), .A2(n8067), .ZN(n8062) );
  INV_X1 U8079 ( .A(n8053), .ZN(n8060) );
  NAND2_X1 U8080 ( .A1(n8068), .A2(n8069), .ZN(n8053) );
  NAND3_X1 U8081 ( .A1(n8070), .A2(n8071), .A3(n8072), .ZN(Result_54_) );
  NAND2_X1 U8082 ( .A1(n7821), .A2(n8073), .ZN(n8072) );
  XOR2_X1 U8083 ( .A(n8074), .B(n8075), .Z(n8073) );
  XNOR2_X1 U8084 ( .A(n8076), .B(n8077), .ZN(n8075) );
  NAND2_X1 U8085 ( .A1(a_22_), .A2(b_31_), .ZN(n8077) );
  NAND2_X1 U8086 ( .A1(n8078), .A2(n8079), .ZN(n8071) );
  NAND3_X1 U8087 ( .A1(n8080), .A2(n8081), .A3(n8082), .ZN(n8079) );
  NAND2_X1 U8088 ( .A1(n7820), .A2(n8083), .ZN(n8082) );
  NAND2_X1 U8089 ( .A1(n8084), .A2(n7819), .ZN(n8081) );
  INV_X1 U8090 ( .A(n8085), .ZN(n8084) );
  NAND2_X1 U8091 ( .A1(n7822), .A2(n8086), .ZN(n8080) );
  NAND2_X1 U8092 ( .A1(n8087), .A2(n8088), .ZN(n8070) );
  NAND3_X1 U8093 ( .A1(n8089), .A2(n8090), .A3(n8091), .ZN(n8088) );
  NAND2_X1 U8094 ( .A1(n7820), .A2(n8092), .ZN(n8091) );
  NAND2_X1 U8095 ( .A1(n7819), .A2(n8085), .ZN(n8090) );
  NAND2_X1 U8096 ( .A1(n7822), .A2(n8093), .ZN(n8089) );
  INV_X1 U8097 ( .A(n8078), .ZN(n8087) );
  XNOR2_X1 U8098 ( .A(n8094), .B(a_22_), .ZN(n8078) );
  NAND3_X1 U8099 ( .A1(n8095), .A2(n8096), .A3(n8097), .ZN(Result_53_) );
  NAND2_X1 U8100 ( .A1(n7821), .A2(n8098), .ZN(n8097) );
  XOR2_X1 U8101 ( .A(n8099), .B(n8100), .Z(n8098) );
  XNOR2_X1 U8102 ( .A(n8101), .B(n8102), .ZN(n8100) );
  NAND2_X1 U8103 ( .A1(a_21_), .A2(b_31_), .ZN(n8102) );
  NAND2_X1 U8104 ( .A1(n8103), .A2(n8104), .ZN(n8096) );
  NAND3_X1 U8105 ( .A1(n8105), .A2(n8106), .A3(n8107), .ZN(n8103) );
  NAND2_X1 U8106 ( .A1(n7820), .A2(n8108), .ZN(n8107) );
  NAND2_X1 U8107 ( .A1(n7819), .A2(n8109), .ZN(n8106) );
  NAND2_X1 U8108 ( .A1(n7822), .A2(n8110), .ZN(n8105) );
  NAND2_X1 U8109 ( .A1(n8111), .A2(n8112), .ZN(n8095) );
  NAND3_X1 U8110 ( .A1(n8113), .A2(n8114), .A3(n8115), .ZN(n8112) );
  NAND2_X1 U8111 ( .A1(n7820), .A2(n8116), .ZN(n8115) );
  NAND2_X1 U8112 ( .A1(n8117), .A2(n7819), .ZN(n8114) );
  NAND2_X1 U8113 ( .A1(n7822), .A2(n8118), .ZN(n8113) );
  INV_X1 U8114 ( .A(n8104), .ZN(n8111) );
  NAND2_X1 U8115 ( .A1(n8119), .A2(n8120), .ZN(n8104) );
  NAND3_X1 U8116 ( .A1(n8121), .A2(n8122), .A3(n8123), .ZN(Result_52_) );
  NAND2_X1 U8117 ( .A1(n7821), .A2(n8124), .ZN(n8123) );
  XOR2_X1 U8118 ( .A(n8125), .B(n8126), .Z(n8124) );
  XNOR2_X1 U8119 ( .A(n8127), .B(n8128), .ZN(n8126) );
  NAND2_X1 U8120 ( .A1(a_20_), .A2(b_31_), .ZN(n8128) );
  NAND2_X1 U8121 ( .A1(n8129), .A2(n8130), .ZN(n8122) );
  NAND3_X1 U8122 ( .A1(n8131), .A2(n8132), .A3(n8133), .ZN(n8130) );
  NAND2_X1 U8123 ( .A1(n7820), .A2(n8134), .ZN(n8133) );
  NAND2_X1 U8124 ( .A1(n8135), .A2(n7819), .ZN(n8132) );
  INV_X1 U8125 ( .A(n8136), .ZN(n8135) );
  NAND2_X1 U8126 ( .A1(n7822), .A2(n8137), .ZN(n8131) );
  NAND2_X1 U8127 ( .A1(n8138), .A2(n8139), .ZN(n8121) );
  NAND3_X1 U8128 ( .A1(n8140), .A2(n8141), .A3(n8142), .ZN(n8139) );
  NAND2_X1 U8129 ( .A1(n7820), .A2(n8143), .ZN(n8142) );
  NAND2_X1 U8130 ( .A1(n7819), .A2(n8136), .ZN(n8141) );
  NAND2_X1 U8131 ( .A1(n7822), .A2(n8144), .ZN(n8140) );
  INV_X1 U8132 ( .A(n8129), .ZN(n8138) );
  XNOR2_X1 U8133 ( .A(n8145), .B(a_20_), .ZN(n8129) );
  NAND3_X1 U8134 ( .A1(n8146), .A2(n8147), .A3(n8148), .ZN(Result_51_) );
  NAND2_X1 U8135 ( .A1(n8149), .A2(n7821), .ZN(n8148) );
  XNOR2_X1 U8136 ( .A(n8150), .B(n8151), .ZN(n8149) );
  XOR2_X1 U8137 ( .A(n8152), .B(n8153), .Z(n8151) );
  NAND2_X1 U8138 ( .A1(a_19_), .A2(b_31_), .ZN(n8153) );
  NAND2_X1 U8139 ( .A1(n8154), .A2(n8155), .ZN(n8147) );
  NAND3_X1 U8140 ( .A1(n8156), .A2(n8157), .A3(n8158), .ZN(n8155) );
  NAND2_X1 U8141 ( .A1(n7820), .A2(n8159), .ZN(n8158) );
  NAND2_X1 U8142 ( .A1(n8160), .A2(n7819), .ZN(n8157) );
  INV_X1 U8143 ( .A(n8161), .ZN(n8160) );
  NAND2_X1 U8144 ( .A1(n7822), .A2(n8162), .ZN(n8156) );
  NAND2_X1 U8145 ( .A1(n8163), .A2(n8164), .ZN(n8146) );
  NAND3_X1 U8146 ( .A1(n8165), .A2(n8166), .A3(n8167), .ZN(n8164) );
  NAND2_X1 U8147 ( .A1(n7820), .A2(n8168), .ZN(n8167) );
  NAND2_X1 U8148 ( .A1(n7819), .A2(n8161), .ZN(n8166) );
  NAND2_X1 U8149 ( .A1(n7822), .A2(n8169), .ZN(n8165) );
  INV_X1 U8150 ( .A(n8154), .ZN(n8163) );
  XNOR2_X1 U8151 ( .A(n8170), .B(b_19_), .ZN(n8154) );
  NAND3_X1 U8152 ( .A1(n8171), .A2(n8172), .A3(n8173), .ZN(Result_50_) );
  NAND2_X1 U8153 ( .A1(n7821), .A2(n8174), .ZN(n8173) );
  XOR2_X1 U8154 ( .A(n8175), .B(n8176), .Z(n8174) );
  XNOR2_X1 U8155 ( .A(n8177), .B(n8178), .ZN(n8176) );
  NAND2_X1 U8156 ( .A1(a_18_), .A2(b_31_), .ZN(n8178) );
  NAND2_X1 U8157 ( .A1(n8179), .A2(n8180), .ZN(n8172) );
  NAND3_X1 U8158 ( .A1(n8181), .A2(n8182), .A3(n8183), .ZN(n8180) );
  NAND2_X1 U8159 ( .A1(n7820), .A2(n8184), .ZN(n8183) );
  NAND2_X1 U8160 ( .A1(n8185), .A2(n7819), .ZN(n8182) );
  INV_X1 U8161 ( .A(n8186), .ZN(n8185) );
  NAND2_X1 U8162 ( .A1(n7822), .A2(n8187), .ZN(n8181) );
  NAND2_X1 U8163 ( .A1(n8188), .A2(n8189), .ZN(n8171) );
  NAND3_X1 U8164 ( .A1(n8190), .A2(n8191), .A3(n8192), .ZN(n8189) );
  NAND2_X1 U8165 ( .A1(n7820), .A2(n8193), .ZN(n8192) );
  NAND2_X1 U8166 ( .A1(n7819), .A2(n8186), .ZN(n8191) );
  NAND2_X1 U8167 ( .A1(n7822), .A2(n8194), .ZN(n8190) );
  INV_X1 U8168 ( .A(n8179), .ZN(n8188) );
  XNOR2_X1 U8169 ( .A(n8195), .B(a_18_), .ZN(n8179) );
  NAND2_X1 U8170 ( .A1(n7823), .A2(n8196), .ZN(Result_4_) );
  NAND2_X1 U8171 ( .A1(n8197), .A2(n7821), .ZN(n8196) );
  XOR2_X1 U8172 ( .A(n8198), .B(n8199), .Z(n8197) );
  AND2_X1 U8173 ( .A1(n8200), .A2(n8201), .ZN(n8199) );
  NAND3_X1 U8174 ( .A1(n8202), .A2(n8203), .A3(n8204), .ZN(Result_49_) );
  NAND2_X1 U8175 ( .A1(n8205), .A2(n7821), .ZN(n8204) );
  XOR2_X1 U8176 ( .A(n8206), .B(n8207), .Z(n8205) );
  XOR2_X1 U8177 ( .A(n8208), .B(n8209), .Z(n8206) );
  NOR2_X1 U8178 ( .A1(n7889), .A2(n8210), .ZN(n8209) );
  NAND2_X1 U8179 ( .A1(n8211), .A2(n8212), .ZN(n8203) );
  NAND3_X1 U8180 ( .A1(n8213), .A2(n8214), .A3(n8215), .ZN(n8212) );
  NAND2_X1 U8181 ( .A1(n7820), .A2(n8216), .ZN(n8215) );
  NAND2_X1 U8182 ( .A1(n8217), .A2(n7819), .ZN(n8214) );
  INV_X1 U8183 ( .A(n8218), .ZN(n8217) );
  NAND2_X1 U8184 ( .A1(n7822), .A2(n8219), .ZN(n8213) );
  NAND2_X1 U8185 ( .A1(n8220), .A2(n8221), .ZN(n8202) );
  NAND3_X1 U8186 ( .A1(n8222), .A2(n8223), .A3(n8224), .ZN(n8221) );
  NAND2_X1 U8187 ( .A1(n7820), .A2(n8225), .ZN(n8224) );
  NAND2_X1 U8188 ( .A1(n7819), .A2(n8218), .ZN(n8223) );
  NAND2_X1 U8189 ( .A1(n7822), .A2(n8226), .ZN(n8222) );
  INV_X1 U8190 ( .A(n8211), .ZN(n8220) );
  XNOR2_X1 U8191 ( .A(n8210), .B(b_17_), .ZN(n8211) );
  NAND3_X1 U8192 ( .A1(n8227), .A2(n8228), .A3(n8229), .ZN(Result_48_) );
  NAND2_X1 U8193 ( .A1(n7821), .A2(n8230), .ZN(n8229) );
  XOR2_X1 U8194 ( .A(n8231), .B(n8232), .Z(n8230) );
  XNOR2_X1 U8195 ( .A(n8233), .B(n8234), .ZN(n8232) );
  NAND2_X1 U8196 ( .A1(a_16_), .A2(b_31_), .ZN(n8234) );
  NAND2_X1 U8197 ( .A1(n8235), .A2(n8236), .ZN(n8228) );
  NAND3_X1 U8198 ( .A1(n8237), .A2(n8238), .A3(n8239), .ZN(n8236) );
  NAND2_X1 U8199 ( .A1(n7820), .A2(n8240), .ZN(n8239) );
  NAND2_X1 U8200 ( .A1(n8241), .A2(n7819), .ZN(n8238) );
  INV_X1 U8201 ( .A(n8242), .ZN(n8241) );
  NAND2_X1 U8202 ( .A1(n7822), .A2(n8243), .ZN(n8237) );
  NAND2_X1 U8203 ( .A1(n8244), .A2(n8245), .ZN(n8227) );
  NAND3_X1 U8204 ( .A1(n8246), .A2(n8247), .A3(n8248), .ZN(n8245) );
  NAND2_X1 U8205 ( .A1(n7820), .A2(n8249), .ZN(n8248) );
  NAND2_X1 U8206 ( .A1(n7819), .A2(n8242), .ZN(n8247) );
  NAND2_X1 U8207 ( .A1(n7822), .A2(n8250), .ZN(n8246) );
  INV_X1 U8208 ( .A(n8235), .ZN(n8244) );
  XNOR2_X1 U8209 ( .A(n8251), .B(a_16_), .ZN(n8235) );
  NAND3_X1 U8210 ( .A1(n8252), .A2(n8253), .A3(n8254), .ZN(Result_47_) );
  NAND2_X1 U8211 ( .A1(n8255), .A2(n7821), .ZN(n8254) );
  XNOR2_X1 U8212 ( .A(n8256), .B(n8257), .ZN(n8255) );
  XOR2_X1 U8213 ( .A(n8258), .B(n8259), .Z(n8257) );
  NAND2_X1 U8214 ( .A1(a_15_), .A2(b_31_), .ZN(n8259) );
  NAND2_X1 U8215 ( .A1(n8260), .A2(n8261), .ZN(n8253) );
  NAND3_X1 U8216 ( .A1(n8262), .A2(n8263), .A3(n8264), .ZN(n8261) );
  NAND2_X1 U8217 ( .A1(n7820), .A2(n8265), .ZN(n8264) );
  NAND2_X1 U8218 ( .A1(n8266), .A2(n7819), .ZN(n8263) );
  NAND2_X1 U8219 ( .A1(n7822), .A2(n8267), .ZN(n8262) );
  NAND2_X1 U8220 ( .A1(n8268), .A2(n8269), .ZN(n8252) );
  NAND3_X1 U8221 ( .A1(n8270), .A2(n8271), .A3(n8272), .ZN(n8269) );
  NAND2_X1 U8222 ( .A1(n7820), .A2(n8273), .ZN(n8272) );
  NAND2_X1 U8223 ( .A1(n7819), .A2(n8274), .ZN(n8271) );
  NAND2_X1 U8224 ( .A1(n7822), .A2(n8275), .ZN(n8270) );
  INV_X1 U8225 ( .A(n8260), .ZN(n8268) );
  XNOR2_X1 U8226 ( .A(n8276), .B(b_15_), .ZN(n8260) );
  NAND3_X1 U8227 ( .A1(n8277), .A2(n8278), .A3(n8279), .ZN(Result_46_) );
  NAND2_X1 U8228 ( .A1(n7821), .A2(n8280), .ZN(n8279) );
  XOR2_X1 U8229 ( .A(n8281), .B(n8282), .Z(n8280) );
  XNOR2_X1 U8230 ( .A(n8283), .B(n8284), .ZN(n8282) );
  NAND2_X1 U8231 ( .A1(a_14_), .A2(b_31_), .ZN(n8284) );
  NAND2_X1 U8232 ( .A1(n8285), .A2(n8286), .ZN(n8278) );
  NAND3_X1 U8233 ( .A1(n8287), .A2(n8288), .A3(n8289), .ZN(n8286) );
  NAND2_X1 U8234 ( .A1(n7820), .A2(n8290), .ZN(n8289) );
  NAND2_X1 U8235 ( .A1(n8291), .A2(n7819), .ZN(n8288) );
  NAND2_X1 U8236 ( .A1(n7822), .A2(n8292), .ZN(n8287) );
  NAND2_X1 U8237 ( .A1(n8293), .A2(n8294), .ZN(n8277) );
  NAND3_X1 U8238 ( .A1(n8295), .A2(n8296), .A3(n8297), .ZN(n8294) );
  NAND2_X1 U8239 ( .A1(n7820), .A2(n8298), .ZN(n8297) );
  NAND2_X1 U8240 ( .A1(n7819), .A2(n8299), .ZN(n8296) );
  NAND2_X1 U8241 ( .A1(n7822), .A2(n8300), .ZN(n8295) );
  INV_X1 U8242 ( .A(n8285), .ZN(n8293) );
  XNOR2_X1 U8243 ( .A(n8301), .B(a_14_), .ZN(n8285) );
  NAND3_X1 U8244 ( .A1(n8302), .A2(n8303), .A3(n8304), .ZN(Result_45_) );
  NAND2_X1 U8245 ( .A1(n8305), .A2(n7821), .ZN(n8304) );
  XOR2_X1 U8246 ( .A(n8306), .B(n8307), .Z(n8305) );
  XOR2_X1 U8247 ( .A(n8308), .B(n8309), .Z(n8306) );
  NOR2_X1 U8248 ( .A1(n7889), .A2(n8310), .ZN(n8309) );
  NAND2_X1 U8249 ( .A1(n8311), .A2(n8312), .ZN(n8303) );
  NAND3_X1 U8250 ( .A1(n8313), .A2(n8314), .A3(n8315), .ZN(n8312) );
  NAND2_X1 U8251 ( .A1(n7820), .A2(n8316), .ZN(n8315) );
  NAND2_X1 U8252 ( .A1(n8317), .A2(n7819), .ZN(n8314) );
  INV_X1 U8253 ( .A(n8318), .ZN(n8317) );
  NAND2_X1 U8254 ( .A1(n7822), .A2(n8319), .ZN(n8313) );
  NAND2_X1 U8255 ( .A1(n8320), .A2(n8321), .ZN(n8302) );
  NAND3_X1 U8256 ( .A1(n8322), .A2(n8323), .A3(n8324), .ZN(n8321) );
  NAND2_X1 U8257 ( .A1(n7820), .A2(n8325), .ZN(n8324) );
  NAND2_X1 U8258 ( .A1(n7819), .A2(n8318), .ZN(n8323) );
  NAND2_X1 U8259 ( .A1(n7822), .A2(n8326), .ZN(n8322) );
  INV_X1 U8260 ( .A(n8311), .ZN(n8320) );
  XNOR2_X1 U8261 ( .A(n8310), .B(b_13_), .ZN(n8311) );
  NAND3_X1 U8262 ( .A1(n8327), .A2(n8328), .A3(n8329), .ZN(Result_44_) );
  NAND2_X1 U8263 ( .A1(n7821), .A2(n8330), .ZN(n8329) );
  XOR2_X1 U8264 ( .A(n8331), .B(n8332), .Z(n8330) );
  XNOR2_X1 U8265 ( .A(n8333), .B(n8334), .ZN(n8332) );
  NAND2_X1 U8266 ( .A1(a_12_), .A2(b_31_), .ZN(n8334) );
  NAND2_X1 U8267 ( .A1(n8335), .A2(n8336), .ZN(n8328) );
  NAND3_X1 U8268 ( .A1(n8337), .A2(n8338), .A3(n8339), .ZN(n8336) );
  NAND2_X1 U8269 ( .A1(n7820), .A2(n8340), .ZN(n8339) );
  NAND2_X1 U8270 ( .A1(n8341), .A2(n7819), .ZN(n8338) );
  INV_X1 U8271 ( .A(n8342), .ZN(n8341) );
  NAND2_X1 U8272 ( .A1(n7822), .A2(n8343), .ZN(n8337) );
  NAND2_X1 U8273 ( .A1(n8344), .A2(n8345), .ZN(n8327) );
  NAND3_X1 U8274 ( .A1(n8346), .A2(n8347), .A3(n8348), .ZN(n8345) );
  NAND2_X1 U8275 ( .A1(n7820), .A2(n8349), .ZN(n8348) );
  NAND2_X1 U8276 ( .A1(n7819), .A2(n8342), .ZN(n8347) );
  NAND2_X1 U8277 ( .A1(n7822), .A2(n8350), .ZN(n8346) );
  INV_X1 U8278 ( .A(n8335), .ZN(n8344) );
  XNOR2_X1 U8279 ( .A(n8351), .B(a_12_), .ZN(n8335) );
  NAND3_X1 U8280 ( .A1(n8352), .A2(n8353), .A3(n8354), .ZN(Result_43_) );
  NAND2_X1 U8281 ( .A1(n8355), .A2(n7821), .ZN(n8354) );
  XNOR2_X1 U8282 ( .A(n8356), .B(n8357), .ZN(n8355) );
  XOR2_X1 U8283 ( .A(n8358), .B(n8359), .Z(n8357) );
  NAND2_X1 U8284 ( .A1(a_11_), .A2(b_31_), .ZN(n8359) );
  NAND2_X1 U8285 ( .A1(n8360), .A2(n8361), .ZN(n8353) );
  NAND3_X1 U8286 ( .A1(n8362), .A2(n8363), .A3(n8364), .ZN(n8361) );
  NAND2_X1 U8287 ( .A1(n7820), .A2(n8365), .ZN(n8364) );
  NAND2_X1 U8288 ( .A1(n8366), .A2(n7819), .ZN(n8363) );
  NAND2_X1 U8289 ( .A1(n7822), .A2(n8367), .ZN(n8362) );
  NAND2_X1 U8290 ( .A1(n8368), .A2(n8369), .ZN(n8352) );
  NAND3_X1 U8291 ( .A1(n8370), .A2(n8371), .A3(n8372), .ZN(n8369) );
  NAND2_X1 U8292 ( .A1(n7820), .A2(n8373), .ZN(n8372) );
  NAND2_X1 U8293 ( .A1(n7819), .A2(n8374), .ZN(n8371) );
  NAND2_X1 U8294 ( .A1(n7822), .A2(n8375), .ZN(n8370) );
  INV_X1 U8295 ( .A(n8360), .ZN(n8368) );
  XNOR2_X1 U8296 ( .A(n8376), .B(b_11_), .ZN(n8360) );
  NAND3_X1 U8297 ( .A1(n8377), .A2(n8378), .A3(n8379), .ZN(Result_42_) );
  NAND2_X1 U8298 ( .A1(n7821), .A2(n8380), .ZN(n8379) );
  XOR2_X1 U8299 ( .A(n8381), .B(n8382), .Z(n8380) );
  XNOR2_X1 U8300 ( .A(n8383), .B(n8384), .ZN(n8382) );
  NAND2_X1 U8301 ( .A1(a_10_), .A2(b_31_), .ZN(n8384) );
  NAND2_X1 U8302 ( .A1(n8385), .A2(n8386), .ZN(n8378) );
  NAND3_X1 U8303 ( .A1(n8387), .A2(n8388), .A3(n8389), .ZN(n8386) );
  NAND2_X1 U8304 ( .A1(n7820), .A2(n8390), .ZN(n8389) );
  NAND2_X1 U8305 ( .A1(n8391), .A2(n7819), .ZN(n8388) );
  INV_X1 U8306 ( .A(n8392), .ZN(n8391) );
  NAND2_X1 U8307 ( .A1(n7822), .A2(n8393), .ZN(n8387) );
  NAND2_X1 U8308 ( .A1(n8394), .A2(n8395), .ZN(n8377) );
  NAND3_X1 U8309 ( .A1(n8396), .A2(n8397), .A3(n8398), .ZN(n8395) );
  NAND2_X1 U8310 ( .A1(n7820), .A2(n8399), .ZN(n8398) );
  NAND2_X1 U8311 ( .A1(n7819), .A2(n8392), .ZN(n8397) );
  NAND2_X1 U8312 ( .A1(n7822), .A2(n8400), .ZN(n8396) );
  INV_X1 U8313 ( .A(n8385), .ZN(n8394) );
  XNOR2_X1 U8314 ( .A(n8401), .B(a_10_), .ZN(n8385) );
  NAND3_X1 U8315 ( .A1(n8402), .A2(n8403), .A3(n8404), .ZN(Result_41_) );
  NAND2_X1 U8316 ( .A1(n7821), .A2(n8405), .ZN(n8404) );
  XOR2_X1 U8317 ( .A(n8406), .B(n8407), .Z(n8405) );
  XNOR2_X1 U8318 ( .A(n8408), .B(n8409), .ZN(n8407) );
  NAND2_X1 U8319 ( .A1(a_9_), .A2(b_31_), .ZN(n8409) );
  NAND2_X1 U8320 ( .A1(n8410), .A2(n8411), .ZN(n8403) );
  NAND3_X1 U8321 ( .A1(n8412), .A2(n8413), .A3(n8414), .ZN(n8411) );
  NAND2_X1 U8322 ( .A1(n7820), .A2(n8415), .ZN(n8414) );
  NAND2_X1 U8323 ( .A1(n8416), .A2(n7819), .ZN(n8413) );
  INV_X1 U8324 ( .A(n8417), .ZN(n8416) );
  NAND2_X1 U8325 ( .A1(n7822), .A2(n8418), .ZN(n8412) );
  NAND2_X1 U8326 ( .A1(n8419), .A2(n8420), .ZN(n8402) );
  NAND3_X1 U8327 ( .A1(n8421), .A2(n8422), .A3(n8423), .ZN(n8420) );
  NAND2_X1 U8328 ( .A1(n7820), .A2(n8424), .ZN(n8423) );
  NAND2_X1 U8329 ( .A1(n7819), .A2(n8417), .ZN(n8422) );
  NAND2_X1 U8330 ( .A1(n7822), .A2(n8425), .ZN(n8421) );
  INV_X1 U8331 ( .A(n8410), .ZN(n8419) );
  XNOR2_X1 U8332 ( .A(n8426), .B(b_9_), .ZN(n8410) );
  NAND3_X1 U8333 ( .A1(n8427), .A2(n8428), .A3(n8429), .ZN(Result_40_) );
  NAND2_X1 U8334 ( .A1(n7821), .A2(n8430), .ZN(n8429) );
  XOR2_X1 U8335 ( .A(n8431), .B(n8432), .Z(n8430) );
  XNOR2_X1 U8336 ( .A(n8433), .B(n8434), .ZN(n8432) );
  NAND2_X1 U8337 ( .A1(a_8_), .A2(b_31_), .ZN(n8434) );
  NAND2_X1 U8338 ( .A1(n8435), .A2(n8436), .ZN(n8428) );
  NAND3_X1 U8339 ( .A1(n8437), .A2(n8438), .A3(n8439), .ZN(n8436) );
  NAND2_X1 U8340 ( .A1(n7820), .A2(n8440), .ZN(n8439) );
  NAND2_X1 U8341 ( .A1(n8441), .A2(n7819), .ZN(n8438) );
  INV_X1 U8342 ( .A(n8442), .ZN(n8441) );
  NAND2_X1 U8343 ( .A1(n7822), .A2(n8443), .ZN(n8437) );
  NAND2_X1 U8344 ( .A1(n8444), .A2(n8445), .ZN(n8427) );
  NAND3_X1 U8345 ( .A1(n8446), .A2(n8447), .A3(n8448), .ZN(n8445) );
  NAND2_X1 U8346 ( .A1(n7820), .A2(n8449), .ZN(n8448) );
  NAND2_X1 U8347 ( .A1(n7819), .A2(n8442), .ZN(n8447) );
  NAND2_X1 U8348 ( .A1(n7822), .A2(n8450), .ZN(n8446) );
  INV_X1 U8349 ( .A(n8435), .ZN(n8444) );
  XNOR2_X1 U8350 ( .A(n8451), .B(a_8_), .ZN(n8435) );
  NAND2_X1 U8351 ( .A1(n7823), .A2(n8452), .ZN(Result_3_) );
  NAND2_X1 U8352 ( .A1(n8453), .A2(n7821), .ZN(n8452) );
  XOR2_X1 U8353 ( .A(n8454), .B(n8455), .Z(n8453) );
  AND2_X1 U8354 ( .A1(n8456), .A2(n8457), .ZN(n8455) );
  NAND3_X1 U8355 ( .A1(n8458), .A2(n8459), .A3(n8460), .ZN(Result_39_) );
  NAND2_X1 U8356 ( .A1(n8461), .A2(n7821), .ZN(n8460) );
  XNOR2_X1 U8357 ( .A(n8462), .B(n8463), .ZN(n8461) );
  XOR2_X1 U8358 ( .A(n8464), .B(n8465), .Z(n8463) );
  NAND2_X1 U8359 ( .A1(a_7_), .A2(b_31_), .ZN(n8465) );
  NAND2_X1 U8360 ( .A1(n8466), .A2(n8467), .ZN(n8459) );
  NAND3_X1 U8361 ( .A1(n8468), .A2(n8469), .A3(n8470), .ZN(n8467) );
  NAND2_X1 U8362 ( .A1(n7820), .A2(n8471), .ZN(n8470) );
  NAND2_X1 U8363 ( .A1(n8472), .A2(n7819), .ZN(n8469) );
  NAND2_X1 U8364 ( .A1(n7822), .A2(n8473), .ZN(n8468) );
  NAND2_X1 U8365 ( .A1(n8474), .A2(n8475), .ZN(n8458) );
  NAND3_X1 U8366 ( .A1(n8476), .A2(n8477), .A3(n8478), .ZN(n8475) );
  NAND2_X1 U8367 ( .A1(n7820), .A2(n8479), .ZN(n8478) );
  NAND2_X1 U8368 ( .A1(n7819), .A2(n8480), .ZN(n8477) );
  NAND2_X1 U8369 ( .A1(n7822), .A2(n8481), .ZN(n8476) );
  INV_X1 U8370 ( .A(n8466), .ZN(n8474) );
  XNOR2_X1 U8371 ( .A(n8482), .B(a_7_), .ZN(n8466) );
  NAND3_X1 U8372 ( .A1(n8483), .A2(n8484), .A3(n8485), .ZN(Result_38_) );
  NAND2_X1 U8373 ( .A1(n8486), .A2(n7821), .ZN(n8485) );
  XOR2_X1 U8374 ( .A(n8487), .B(n8488), .Z(n8486) );
  XOR2_X1 U8375 ( .A(n8489), .B(n8490), .Z(n8487) );
  NOR2_X1 U8376 ( .A1(n7889), .A2(n8491), .ZN(n8490) );
  NAND2_X1 U8377 ( .A1(n8492), .A2(n8493), .ZN(n8484) );
  NAND3_X1 U8378 ( .A1(n8494), .A2(n8495), .A3(n8496), .ZN(n8493) );
  NAND2_X1 U8379 ( .A1(n7820), .A2(n8497), .ZN(n8496) );
  NAND2_X1 U8380 ( .A1(n8498), .A2(n7819), .ZN(n8495) );
  INV_X1 U8381 ( .A(n8499), .ZN(n8498) );
  NAND2_X1 U8382 ( .A1(n7822), .A2(n8500), .ZN(n8494) );
  NAND2_X1 U8383 ( .A1(n8501), .A2(n8502), .ZN(n8483) );
  NAND3_X1 U8384 ( .A1(n8503), .A2(n8504), .A3(n8505), .ZN(n8502) );
  NAND2_X1 U8385 ( .A1(n7820), .A2(n8506), .ZN(n8505) );
  NAND2_X1 U8386 ( .A1(n7819), .A2(n8499), .ZN(n8504) );
  NAND2_X1 U8387 ( .A1(n7822), .A2(n8507), .ZN(n8503) );
  INV_X1 U8388 ( .A(n8492), .ZN(n8501) );
  XNOR2_X1 U8389 ( .A(n8508), .B(a_6_), .ZN(n8492) );
  NAND3_X1 U8390 ( .A1(n8509), .A2(n8510), .A3(n8511), .ZN(Result_37_) );
  NAND2_X1 U8391 ( .A1(n8512), .A2(n7821), .ZN(n8511) );
  XOR2_X1 U8392 ( .A(n8513), .B(n8514), .Z(n8512) );
  XOR2_X1 U8393 ( .A(n8515), .B(n8516), .Z(n8513) );
  NOR2_X1 U8394 ( .A1(n7889), .A2(n8517), .ZN(n8516) );
  NAND2_X1 U8395 ( .A1(n8518), .A2(n8519), .ZN(n8510) );
  NAND3_X1 U8396 ( .A1(n8520), .A2(n8521), .A3(n8522), .ZN(n8519) );
  NAND2_X1 U8397 ( .A1(n7820), .A2(n8523), .ZN(n8522) );
  NAND2_X1 U8398 ( .A1(n8524), .A2(n7819), .ZN(n8521) );
  INV_X1 U8399 ( .A(n8525), .ZN(n8524) );
  NAND2_X1 U8400 ( .A1(n7822), .A2(n8526), .ZN(n8520) );
  NAND2_X1 U8401 ( .A1(n8527), .A2(n8528), .ZN(n8509) );
  NAND3_X1 U8402 ( .A1(n8529), .A2(n8530), .A3(n8531), .ZN(n8528) );
  NAND2_X1 U8403 ( .A1(n7820), .A2(n8532), .ZN(n8531) );
  NAND2_X1 U8404 ( .A1(n7819), .A2(n8525), .ZN(n8530) );
  NAND2_X1 U8405 ( .A1(n7822), .A2(n8533), .ZN(n8529) );
  INV_X1 U8406 ( .A(n8518), .ZN(n8527) );
  XNOR2_X1 U8407 ( .A(n8517), .B(b_5_), .ZN(n8518) );
  NAND3_X1 U8408 ( .A1(n8534), .A2(n8535), .A3(n8536), .ZN(Result_36_) );
  NAND2_X1 U8409 ( .A1(n7821), .A2(n8537), .ZN(n8536) );
  XOR2_X1 U8410 ( .A(n8538), .B(n8539), .Z(n8537) );
  XNOR2_X1 U8411 ( .A(n8540), .B(n8541), .ZN(n8539) );
  NAND2_X1 U8412 ( .A1(a_4_), .A2(b_31_), .ZN(n8541) );
  NAND2_X1 U8413 ( .A1(n8542), .A2(n8543), .ZN(n8535) );
  NAND3_X1 U8414 ( .A1(n8544), .A2(n8545), .A3(n8546), .ZN(n8543) );
  NAND2_X1 U8415 ( .A1(n7820), .A2(n8547), .ZN(n8546) );
  NAND2_X1 U8416 ( .A1(n8548), .A2(n7819), .ZN(n8545) );
  INV_X1 U8417 ( .A(n8549), .ZN(n8548) );
  NAND2_X1 U8418 ( .A1(n7822), .A2(n8550), .ZN(n8544) );
  NAND2_X1 U8419 ( .A1(n8551), .A2(n8552), .ZN(n8534) );
  NAND3_X1 U8420 ( .A1(n8553), .A2(n8554), .A3(n8555), .ZN(n8552) );
  NAND2_X1 U8421 ( .A1(n7820), .A2(n8556), .ZN(n8555) );
  NAND2_X1 U8422 ( .A1(n7819), .A2(n8549), .ZN(n8554) );
  NAND2_X1 U8423 ( .A1(n7822), .A2(n8557), .ZN(n8553) );
  INV_X1 U8424 ( .A(n8542), .ZN(n8551) );
  XNOR2_X1 U8425 ( .A(n8558), .B(a_4_), .ZN(n8542) );
  NAND3_X1 U8426 ( .A1(n8559), .A2(n8560), .A3(n8561), .ZN(Result_35_) );
  NAND2_X1 U8427 ( .A1(n8562), .A2(n7821), .ZN(n8561) );
  XOR2_X1 U8428 ( .A(n8563), .B(n8564), .Z(n8562) );
  XOR2_X1 U8429 ( .A(n8565), .B(n8566), .Z(n8563) );
  NOR2_X1 U8430 ( .A1(n7889), .A2(n8567), .ZN(n8566) );
  NAND2_X1 U8431 ( .A1(n8568), .A2(n8569), .ZN(n8560) );
  NAND3_X1 U8432 ( .A1(n8570), .A2(n8571), .A3(n8572), .ZN(n8569) );
  NAND2_X1 U8433 ( .A1(n7820), .A2(n8573), .ZN(n8572) );
  NAND2_X1 U8434 ( .A1(n8574), .A2(n7819), .ZN(n8571) );
  INV_X1 U8435 ( .A(n8575), .ZN(n8574) );
  NAND2_X1 U8436 ( .A1(n7822), .A2(n8576), .ZN(n8570) );
  NAND2_X1 U8437 ( .A1(n8577), .A2(n8578), .ZN(n8559) );
  NAND3_X1 U8438 ( .A1(n8579), .A2(n8580), .A3(n8581), .ZN(n8578) );
  NAND2_X1 U8439 ( .A1(n7820), .A2(n8582), .ZN(n8581) );
  NAND2_X1 U8440 ( .A1(n7819), .A2(n8575), .ZN(n8580) );
  NAND2_X1 U8441 ( .A1(n7822), .A2(n8583), .ZN(n8579) );
  INV_X1 U8442 ( .A(n8568), .ZN(n8577) );
  XNOR2_X1 U8443 ( .A(n8567), .B(b_3_), .ZN(n8568) );
  NAND3_X1 U8444 ( .A1(n8584), .A2(n8585), .A3(n8586), .ZN(Result_34_) );
  NAND2_X1 U8445 ( .A1(n7821), .A2(n8587), .ZN(n8586) );
  XOR2_X1 U8446 ( .A(n8588), .B(n8589), .Z(n8587) );
  XNOR2_X1 U8447 ( .A(n8590), .B(n8591), .ZN(n8589) );
  NAND2_X1 U8448 ( .A1(a_2_), .A2(b_31_), .ZN(n8591) );
  NAND2_X1 U8449 ( .A1(n8592), .A2(n8593), .ZN(n8585) );
  NAND3_X1 U8450 ( .A1(n8594), .A2(n8595), .A3(n8596), .ZN(n8593) );
  NAND2_X1 U8451 ( .A1(n7820), .A2(n8597), .ZN(n8596) );
  NAND2_X1 U8452 ( .A1(n8598), .A2(n7819), .ZN(n8595) );
  INV_X1 U8453 ( .A(n8599), .ZN(n8598) );
  NAND2_X1 U8454 ( .A1(n7822), .A2(n8600), .ZN(n8594) );
  NAND2_X1 U8455 ( .A1(n8601), .A2(n8602), .ZN(n8584) );
  NAND3_X1 U8456 ( .A1(n8603), .A2(n8604), .A3(n8605), .ZN(n8602) );
  NAND2_X1 U8457 ( .A1(n7820), .A2(n8606), .ZN(n8605) );
  NAND2_X1 U8458 ( .A1(n7819), .A2(n8599), .ZN(n8604) );
  NAND2_X1 U8459 ( .A1(n7822), .A2(n8607), .ZN(n8603) );
  INV_X1 U8460 ( .A(n8592), .ZN(n8601) );
  XNOR2_X1 U8461 ( .A(n8608), .B(a_2_), .ZN(n8592) );
  NAND3_X1 U8462 ( .A1(n8609), .A2(n8610), .A3(n8611), .ZN(Result_33_) );
  NAND2_X1 U8463 ( .A1(n8612), .A2(n7821), .ZN(n8611) );
  XOR2_X1 U8464 ( .A(n8613), .B(n8614), .Z(n8612) );
  XOR2_X1 U8465 ( .A(n8615), .B(n8616), .Z(n8613) );
  NOR2_X1 U8466 ( .A1(n7889), .A2(n8617), .ZN(n8616) );
  NAND2_X1 U8467 ( .A1(n8618), .A2(n8619), .ZN(n8610) );
  NAND3_X1 U8468 ( .A1(n8620), .A2(n8621), .A3(n8622), .ZN(n8619) );
  NAND2_X1 U8469 ( .A1(n7820), .A2(n8623), .ZN(n8622) );
  NAND2_X1 U8470 ( .A1(n8624), .A2(n7819), .ZN(n8621) );
  INV_X1 U8471 ( .A(n8625), .ZN(n8624) );
  NAND2_X1 U8472 ( .A1(n7822), .A2(n8626), .ZN(n8620) );
  NAND2_X1 U8473 ( .A1(n8627), .A2(n8628), .ZN(n8609) );
  NAND3_X1 U8474 ( .A1(n8629), .A2(n8630), .A3(n8631), .ZN(n8628) );
  NAND2_X1 U8475 ( .A1(n7820), .A2(n8632), .ZN(n8631) );
  NAND2_X1 U8476 ( .A1(n7819), .A2(n8625), .ZN(n8630) );
  NAND2_X1 U8477 ( .A1(n7822), .A2(n8633), .ZN(n8629) );
  INV_X1 U8478 ( .A(n8618), .ZN(n8627) );
  XNOR2_X1 U8479 ( .A(n8634), .B(a_1_), .ZN(n8618) );
  NAND3_X1 U8480 ( .A1(n8635), .A2(n8636), .A3(n8637), .ZN(Result_32_) );
  NAND2_X1 U8481 ( .A1(n7821), .A2(n8638), .ZN(n8637) );
  XOR2_X1 U8482 ( .A(n8639), .B(n8640), .Z(n8638) );
  XNOR2_X1 U8483 ( .A(n8641), .B(n8642), .ZN(n8640) );
  NAND2_X1 U8484 ( .A1(a_0_), .A2(b_31_), .ZN(n8642) );
  NAND2_X1 U8485 ( .A1(n8643), .A2(n8644), .ZN(n8636) );
  NAND3_X1 U8486 ( .A1(n8645), .A2(n8646), .A3(n8647), .ZN(n8644) );
  NAND2_X1 U8487 ( .A1(n7820), .A2(n8648), .ZN(n8647) );
  NAND2_X1 U8488 ( .A1(n7819), .A2(n8649), .ZN(n8646) );
  NAND2_X1 U8489 ( .A1(n7822), .A2(n8650), .ZN(n8645) );
  NAND2_X1 U8490 ( .A1(n8651), .A2(n8652), .ZN(n8635) );
  NAND3_X1 U8491 ( .A1(n8653), .A2(n8654), .A3(n8655), .ZN(n8652) );
  NAND2_X1 U8492 ( .A1(n7820), .A2(n8656), .ZN(n8655) );
  NAND2_X1 U8493 ( .A1(n8657), .A2(n7819), .ZN(n8654) );
  INV_X1 U8494 ( .A(n8649), .ZN(n8657) );
  NAND2_X1 U8495 ( .A1(n8658), .A2(n8659), .ZN(n8649) );
  OR2_X1 U8496 ( .A1(n8625), .A2(n8660), .ZN(n8659) );
  NAND2_X1 U8497 ( .A1(n8661), .A2(n8662), .ZN(n8625) );
  NAND2_X1 U8498 ( .A1(n8663), .A2(n8599), .ZN(n8662) );
  NAND2_X1 U8499 ( .A1(n8664), .A2(n8665), .ZN(n8599) );
  NAND2_X1 U8500 ( .A1(n8666), .A2(n8575), .ZN(n8665) );
  NAND2_X1 U8501 ( .A1(n8667), .A2(n8668), .ZN(n8575) );
  NAND2_X1 U8502 ( .A1(n8669), .A2(n8549), .ZN(n8668) );
  NAND2_X1 U8503 ( .A1(n8670), .A2(n8671), .ZN(n8549) );
  NAND2_X1 U8504 ( .A1(n8672), .A2(n8525), .ZN(n8671) );
  NAND2_X1 U8505 ( .A1(n8673), .A2(n8674), .ZN(n8525) );
  NAND2_X1 U8506 ( .A1(n8675), .A2(n8499), .ZN(n8674) );
  NAND2_X1 U8507 ( .A1(n8676), .A2(n8677), .ZN(n8499) );
  NAND2_X1 U8508 ( .A1(n8678), .A2(n8480), .ZN(n8677) );
  INV_X1 U8509 ( .A(n8472), .ZN(n8480) );
  NOR2_X1 U8510 ( .A1(n8679), .A2(n8680), .ZN(n8472) );
  AND2_X1 U8511 ( .A1(n8681), .A2(n8442), .ZN(n8680) );
  NAND2_X1 U8512 ( .A1(n8682), .A2(n8683), .ZN(n8442) );
  NAND2_X1 U8513 ( .A1(n8684), .A2(n8417), .ZN(n8683) );
  NAND2_X1 U8514 ( .A1(n8685), .A2(n8686), .ZN(n8417) );
  NAND2_X1 U8515 ( .A1(n8687), .A2(n8392), .ZN(n8686) );
  NAND2_X1 U8516 ( .A1(n8688), .A2(n8689), .ZN(n8392) );
  NAND2_X1 U8517 ( .A1(n8690), .A2(n8374), .ZN(n8689) );
  INV_X1 U8518 ( .A(n8366), .ZN(n8374) );
  NOR2_X1 U8519 ( .A1(n8691), .A2(n8692), .ZN(n8366) );
  AND2_X1 U8520 ( .A1(n8693), .A2(n8342), .ZN(n8692) );
  NAND2_X1 U8521 ( .A1(n8694), .A2(n8695), .ZN(n8342) );
  NAND2_X1 U8522 ( .A1(n8696), .A2(n8318), .ZN(n8695) );
  NAND2_X1 U8523 ( .A1(n8697), .A2(n8698), .ZN(n8318) );
  NAND2_X1 U8524 ( .A1(n8699), .A2(n8299), .ZN(n8698) );
  INV_X1 U8525 ( .A(n8291), .ZN(n8299) );
  NOR2_X1 U8526 ( .A1(n8700), .A2(n8701), .ZN(n8291) );
  AND2_X1 U8527 ( .A1(n8702), .A2(n8274), .ZN(n8701) );
  INV_X1 U8528 ( .A(n8266), .ZN(n8274) );
  NOR2_X1 U8529 ( .A1(n8703), .A2(n8704), .ZN(n8266) );
  AND2_X1 U8530 ( .A1(n8705), .A2(n8242), .ZN(n8704) );
  NAND2_X1 U8531 ( .A1(n8706), .A2(n8707), .ZN(n8242) );
  NAND2_X1 U8532 ( .A1(n8708), .A2(n8218), .ZN(n8707) );
  NAND2_X1 U8533 ( .A1(n8709), .A2(n8710), .ZN(n8218) );
  NAND2_X1 U8534 ( .A1(n8711), .A2(n8186), .ZN(n8710) );
  NAND2_X1 U8535 ( .A1(n8712), .A2(n8713), .ZN(n8186) );
  NAND2_X1 U8536 ( .A1(n8714), .A2(n8161), .ZN(n8713) );
  NAND2_X1 U8537 ( .A1(n8715), .A2(n8716), .ZN(n8161) );
  NAND2_X1 U8538 ( .A1(n8717), .A2(n8136), .ZN(n8716) );
  NAND2_X1 U8539 ( .A1(n8119), .A2(n8718), .ZN(n8136) );
  NAND2_X1 U8540 ( .A1(n8120), .A2(n8109), .ZN(n8718) );
  INV_X1 U8541 ( .A(n8117), .ZN(n8109) );
  NOR2_X1 U8542 ( .A1(n8719), .A2(n8720), .ZN(n8117) );
  AND2_X1 U8543 ( .A1(n8721), .A2(n8085), .ZN(n8720) );
  NAND2_X1 U8544 ( .A1(n8068), .A2(n8722), .ZN(n8085) );
  NAND2_X1 U8545 ( .A1(n8069), .A2(n8058), .ZN(n8722) );
  NAND2_X1 U8546 ( .A1(n8723), .A2(n8724), .ZN(n8058) );
  NAND2_X1 U8547 ( .A1(n8725), .A2(n8034), .ZN(n8724) );
  NAND2_X1 U8548 ( .A1(n8017), .A2(n8726), .ZN(n8034) );
  NAND2_X1 U8549 ( .A1(n8018), .A2(n8007), .ZN(n8726) );
  NAND2_X1 U8550 ( .A1(n8727), .A2(n8728), .ZN(n8007) );
  NAND2_X1 U8551 ( .A1(n8729), .A2(n7983), .ZN(n8728) );
  NAND2_X1 U8552 ( .A1(n7966), .A2(n8730), .ZN(n7983) );
  NAND2_X1 U8553 ( .A1(n7967), .A2(n7956), .ZN(n8730) );
  NAND2_X1 U8554 ( .A1(n8731), .A2(n8732), .ZN(n7956) );
  NAND2_X1 U8555 ( .A1(n8733), .A2(n7926), .ZN(n8732) );
  NAND2_X1 U8556 ( .A1(n7909), .A2(n8734), .ZN(n7926) );
  NAND2_X1 U8557 ( .A1(n7910), .A2(n7899), .ZN(n8734) );
  NAND2_X1 U8558 ( .A1(n8735), .A2(n8736), .ZN(n7899) );
  NAND2_X1 U8559 ( .A1(b_30_), .A2(n8737), .ZN(n8736) );
  NAND2_X1 U8560 ( .A1(n7867), .A2(n7876), .ZN(n8737) );
  NAND2_X1 U8561 ( .A1(a_31_), .A2(b_31_), .ZN(n7876) );
  NAND2_X1 U8562 ( .A1(n7818), .A2(b_31_), .ZN(n8735) );
  NAND2_X1 U8563 ( .A1(n8738), .A2(n7890), .ZN(n7910) );
  NAND2_X1 U8564 ( .A1(n7935), .A2(n8739), .ZN(n8733) );
  NAND2_X1 U8565 ( .A1(n8740), .A2(n8741), .ZN(n7967) );
  NAND2_X1 U8566 ( .A1(n7992), .A2(n8742), .ZN(n8729) );
  NAND2_X1 U8567 ( .A1(n8743), .A2(n8744), .ZN(n8018) );
  NAND2_X1 U8568 ( .A1(n8043), .A2(n8745), .ZN(n8725) );
  NAND2_X1 U8569 ( .A1(n8746), .A2(n8747), .ZN(n8069) );
  NAND2_X1 U8570 ( .A1(n8094), .A2(n8748), .ZN(n8721) );
  NAND2_X1 U8571 ( .A1(n8749), .A2(n8750), .ZN(n8120) );
  NAND2_X1 U8572 ( .A1(n8145), .A2(n8751), .ZN(n8717) );
  NAND2_X1 U8573 ( .A1(n8752), .A2(n8170), .ZN(n8714) );
  NAND2_X1 U8574 ( .A1(n8195), .A2(n8753), .ZN(n8711) );
  NAND2_X1 U8575 ( .A1(n8754), .A2(n8210), .ZN(n8708) );
  NAND2_X1 U8576 ( .A1(n8251), .A2(n8755), .ZN(n8705) );
  NAND2_X1 U8577 ( .A1(n8756), .A2(n8276), .ZN(n8702) );
  NAND2_X1 U8578 ( .A1(n8301), .A2(n8757), .ZN(n8699) );
  NAND2_X1 U8579 ( .A1(n8758), .A2(n8310), .ZN(n8696) );
  NAND2_X1 U8580 ( .A1(n8351), .A2(n8759), .ZN(n8693) );
  NAND2_X1 U8581 ( .A1(n8760), .A2(n8376), .ZN(n8690) );
  NAND2_X1 U8582 ( .A1(n8401), .A2(n8761), .ZN(n8687) );
  NAND2_X1 U8583 ( .A1(n8762), .A2(n8426), .ZN(n8684) );
  NAND2_X1 U8584 ( .A1(n8451), .A2(n8763), .ZN(n8681) );
  NAND2_X1 U8585 ( .A1(n8482), .A2(n8764), .ZN(n8678) );
  NAND2_X1 U8586 ( .A1(n8508), .A2(n8491), .ZN(n8675) );
  NAND2_X1 U8587 ( .A1(n8765), .A2(n8517), .ZN(n8672) );
  NAND2_X1 U8588 ( .A1(n8558), .A2(n8766), .ZN(n8669) );
  NAND2_X1 U8589 ( .A1(n8767), .A2(n8567), .ZN(n8666) );
  NAND2_X1 U8590 ( .A1(n8608), .A2(n8768), .ZN(n8663) );
  NAND2_X1 U8591 ( .A1(n8634), .A2(n8617), .ZN(n8658) );
  NAND2_X1 U8592 ( .A1(n7822), .A2(n8769), .ZN(n8653) );
  INV_X1 U8593 ( .A(n8643), .ZN(n8651) );
  XNOR2_X1 U8594 ( .A(n8770), .B(a_0_), .ZN(n8643) );
  NAND2_X1 U8595 ( .A1(n7823), .A2(n8771), .ZN(Result_31_) );
  NAND2_X1 U8596 ( .A1(n8772), .A2(n7821), .ZN(n8771) );
  XOR2_X1 U8597 ( .A(n8773), .B(n8774), .Z(n8772) );
  NAND2_X1 U8598 ( .A1(n7823), .A2(n8775), .ZN(Result_30_) );
  NAND3_X1 U8599 ( .A1(n8776), .A2(n8777), .A3(n7821), .ZN(n8775) );
  NAND2_X1 U8600 ( .A1(n8778), .A2(n8779), .ZN(n8776) );
  NAND2_X1 U8601 ( .A1(n8774), .A2(n8773), .ZN(n8779) );
  XNOR2_X1 U8602 ( .A(n8780), .B(n8781), .ZN(n8778) );
  NAND2_X1 U8603 ( .A1(n7823), .A2(n8782), .ZN(Result_2_) );
  NAND2_X1 U8604 ( .A1(n8783), .A2(n7821), .ZN(n8782) );
  XOR2_X1 U8605 ( .A(n8784), .B(n8785), .Z(n8783) );
  AND2_X1 U8606 ( .A1(n8786), .A2(n8787), .ZN(n8785) );
  NAND2_X1 U8607 ( .A1(n7823), .A2(n8788), .ZN(Result_29_) );
  NAND2_X1 U8608 ( .A1(n7821), .A2(n8789), .ZN(n8788) );
  XOR2_X1 U8609 ( .A(n8777), .B(n8790), .Z(n8789) );
  NAND2_X1 U8610 ( .A1(n8791), .A2(n8792), .ZN(n8790) );
  NAND2_X1 U8611 ( .A1(n7823), .A2(n8793), .ZN(Result_28_) );
  NAND2_X1 U8612 ( .A1(n8794), .A2(n7821), .ZN(n8793) );
  XNOR2_X1 U8613 ( .A(n8795), .B(n8796), .ZN(n8794) );
  NAND2_X1 U8614 ( .A1(n8797), .A2(n8798), .ZN(n8795) );
  NAND2_X1 U8615 ( .A1(n7823), .A2(n8799), .ZN(Result_27_) );
  NAND2_X1 U8616 ( .A1(n8800), .A2(n7821), .ZN(n8799) );
  XNOR2_X1 U8617 ( .A(n8801), .B(n8802), .ZN(n8800) );
  NAND2_X1 U8618 ( .A1(n8803), .A2(n8804), .ZN(n8801) );
  NAND2_X1 U8619 ( .A1(n7823), .A2(n8805), .ZN(Result_26_) );
  NAND2_X1 U8620 ( .A1(n8806), .A2(n7821), .ZN(n8805) );
  XOR2_X1 U8621 ( .A(n8807), .B(n8808), .Z(n8806) );
  AND2_X1 U8622 ( .A1(n8809), .A2(n8810), .ZN(n8808) );
  NAND2_X1 U8623 ( .A1(n7823), .A2(n8811), .ZN(Result_25_) );
  NAND2_X1 U8624 ( .A1(n8812), .A2(n7821), .ZN(n8811) );
  XOR2_X1 U8625 ( .A(n8813), .B(n8814), .Z(n8812) );
  AND2_X1 U8626 ( .A1(n8815), .A2(n8816), .ZN(n8814) );
  NAND2_X1 U8627 ( .A1(n7823), .A2(n8817), .ZN(Result_24_) );
  NAND2_X1 U8628 ( .A1(n8818), .A2(n7821), .ZN(n8817) );
  XOR2_X1 U8629 ( .A(n8819), .B(n8820), .Z(n8818) );
  AND2_X1 U8630 ( .A1(n8821), .A2(n8822), .ZN(n8820) );
  NAND2_X1 U8631 ( .A1(n7823), .A2(n8823), .ZN(Result_23_) );
  NAND2_X1 U8632 ( .A1(n8824), .A2(n7821), .ZN(n8823) );
  XOR2_X1 U8633 ( .A(n8825), .B(n8826), .Z(n8824) );
  AND2_X1 U8634 ( .A1(n8827), .A2(n8828), .ZN(n8826) );
  NAND2_X1 U8635 ( .A1(n7823), .A2(n8829), .ZN(Result_22_) );
  NAND2_X1 U8636 ( .A1(n8830), .A2(n7821), .ZN(n8829) );
  XOR2_X1 U8637 ( .A(n8831), .B(n8832), .Z(n8830) );
  AND2_X1 U8638 ( .A1(n8833), .A2(n8834), .ZN(n8832) );
  NAND2_X1 U8639 ( .A1(n7823), .A2(n8835), .ZN(Result_21_) );
  NAND2_X1 U8640 ( .A1(n8836), .A2(n7821), .ZN(n8835) );
  XOR2_X1 U8641 ( .A(n8837), .B(n8838), .Z(n8836) );
  AND2_X1 U8642 ( .A1(n8839), .A2(n8840), .ZN(n8838) );
  NAND2_X1 U8643 ( .A1(n7823), .A2(n8841), .ZN(Result_20_) );
  NAND2_X1 U8644 ( .A1(n8842), .A2(n7821), .ZN(n8841) );
  XOR2_X1 U8645 ( .A(n8843), .B(n8844), .Z(n8842) );
  AND2_X1 U8646 ( .A1(n8845), .A2(n8846), .ZN(n8844) );
  NAND2_X1 U8647 ( .A1(n7823), .A2(n8847), .ZN(Result_1_) );
  NAND2_X1 U8648 ( .A1(n8848), .A2(n7821), .ZN(n8847) );
  XOR2_X1 U8649 ( .A(n8849), .B(n8850), .Z(n8848) );
  AND2_X1 U8650 ( .A1(n8851), .A2(n8852), .ZN(n8850) );
  NAND2_X1 U8651 ( .A1(n7823), .A2(n8853), .ZN(Result_19_) );
  NAND2_X1 U8652 ( .A1(n8854), .A2(n7821), .ZN(n8853) );
  XOR2_X1 U8653 ( .A(n8855), .B(n8856), .Z(n8854) );
  AND2_X1 U8654 ( .A1(n8857), .A2(n8858), .ZN(n8856) );
  NAND2_X1 U8655 ( .A1(n7823), .A2(n8859), .ZN(Result_18_) );
  NAND2_X1 U8656 ( .A1(n8860), .A2(n7821), .ZN(n8859) );
  XOR2_X1 U8657 ( .A(n8861), .B(n8862), .Z(n8860) );
  AND2_X1 U8658 ( .A1(n8863), .A2(n8864), .ZN(n8862) );
  NAND2_X1 U8659 ( .A1(n7823), .A2(n8865), .ZN(Result_17_) );
  NAND2_X1 U8660 ( .A1(n8866), .A2(n7821), .ZN(n8865) );
  XOR2_X1 U8661 ( .A(n8867), .B(n8868), .Z(n8866) );
  AND2_X1 U8662 ( .A1(n8869), .A2(n8870), .ZN(n8868) );
  NAND2_X1 U8663 ( .A1(n7823), .A2(n8871), .ZN(Result_16_) );
  NAND2_X1 U8664 ( .A1(n8872), .A2(n7821), .ZN(n8871) );
  XOR2_X1 U8665 ( .A(n8873), .B(n8874), .Z(n8872) );
  AND2_X1 U8666 ( .A1(n8875), .A2(n8876), .ZN(n8874) );
  NAND2_X1 U8667 ( .A1(n7823), .A2(n8877), .ZN(Result_15_) );
  NAND2_X1 U8668 ( .A1(n8878), .A2(n7821), .ZN(n8877) );
  XOR2_X1 U8669 ( .A(n8879), .B(n8880), .Z(n8878) );
  AND2_X1 U8670 ( .A1(n8881), .A2(n8882), .ZN(n8880) );
  NAND2_X1 U8671 ( .A1(n7823), .A2(n8883), .ZN(Result_14_) );
  NAND2_X1 U8672 ( .A1(n8884), .A2(n7821), .ZN(n8883) );
  XOR2_X1 U8673 ( .A(n8885), .B(n8886), .Z(n8884) );
  AND2_X1 U8674 ( .A1(n8887), .A2(n8888), .ZN(n8886) );
  NAND2_X1 U8675 ( .A1(n7823), .A2(n8889), .ZN(Result_13_) );
  NAND2_X1 U8676 ( .A1(n8890), .A2(n7821), .ZN(n8889) );
  XOR2_X1 U8677 ( .A(n8891), .B(n8892), .Z(n8890) );
  AND2_X1 U8678 ( .A1(n8893), .A2(n8894), .ZN(n8892) );
  NAND2_X1 U8679 ( .A1(n7823), .A2(n8895), .ZN(Result_12_) );
  NAND2_X1 U8680 ( .A1(n8896), .A2(n7821), .ZN(n8895) );
  XOR2_X1 U8681 ( .A(n8897), .B(n8898), .Z(n8896) );
  AND2_X1 U8682 ( .A1(n8899), .A2(n8900), .ZN(n8898) );
  NAND2_X1 U8683 ( .A1(n7823), .A2(n8901), .ZN(Result_11_) );
  NAND2_X1 U8684 ( .A1(n8902), .A2(n7821), .ZN(n8901) );
  XOR2_X1 U8685 ( .A(n8903), .B(n8904), .Z(n8902) );
  AND2_X1 U8686 ( .A1(n8905), .A2(n8906), .ZN(n8904) );
  NAND2_X1 U8687 ( .A1(n7823), .A2(n8907), .ZN(Result_10_) );
  NAND2_X1 U8688 ( .A1(n8908), .A2(n7821), .ZN(n8907) );
  XOR2_X1 U8689 ( .A(n8909), .B(n8910), .Z(n8908) );
  AND2_X1 U8690 ( .A1(n8911), .A2(n8912), .ZN(n8910) );
  NAND2_X1 U8691 ( .A1(n7823), .A2(n8913), .ZN(Result_0_) );
  NAND2_X1 U8692 ( .A1(n7821), .A2(n8914), .ZN(n8913) );
  NAND3_X1 U8693 ( .A1(n8915), .A2(n8852), .A3(n8916), .ZN(n8914) );
  NAND2_X1 U8694 ( .A1(a_0_), .A2(n8917), .ZN(n8916) );
  NAND4_X1 U8695 ( .A1(n8918), .A2(n8919), .A3(n8920), .A4(n8921), .ZN(n8852)
         );
  NAND2_X1 U8696 ( .A1(n8851), .A2(n8849), .ZN(n8915) );
  NAND2_X1 U8697 ( .A1(n8787), .A2(n8922), .ZN(n8849) );
  NAND2_X1 U8698 ( .A1(n8786), .A2(n8784), .ZN(n8922) );
  NAND2_X1 U8699 ( .A1(n8457), .A2(n8923), .ZN(n8784) );
  NAND2_X1 U8700 ( .A1(n8456), .A2(n8454), .ZN(n8923) );
  NAND2_X1 U8701 ( .A1(n8201), .A2(n8924), .ZN(n8454) );
  NAND2_X1 U8702 ( .A1(n8200), .A2(n8198), .ZN(n8924) );
  NAND2_X1 U8703 ( .A1(n7941), .A2(n8925), .ZN(n8198) );
  NAND2_X1 U8704 ( .A1(n7940), .A2(n7938), .ZN(n8925) );
  NAND2_X1 U8705 ( .A1(n7847), .A2(n8926), .ZN(n7938) );
  NAND2_X1 U8706 ( .A1(n7846), .A2(n7844), .ZN(n8926) );
  NAND2_X1 U8707 ( .A1(n7841), .A2(n8927), .ZN(n7844) );
  NAND2_X1 U8708 ( .A1(n7840), .A2(n7838), .ZN(n8927) );
  NAND2_X1 U8709 ( .A1(n7835), .A2(n8928), .ZN(n7838) );
  NAND2_X1 U8710 ( .A1(n7834), .A2(n7832), .ZN(n8928) );
  NAND2_X1 U8711 ( .A1(n7829), .A2(n8929), .ZN(n7832) );
  NAND2_X1 U8712 ( .A1(n7828), .A2(n7826), .ZN(n8929) );
  NAND2_X1 U8713 ( .A1(n8912), .A2(n8930), .ZN(n7826) );
  NAND2_X1 U8714 ( .A1(n8909), .A2(n8911), .ZN(n8930) );
  NAND2_X1 U8715 ( .A1(n8931), .A2(n8932), .ZN(n8911) );
  NAND2_X1 U8716 ( .A1(n8906), .A2(n8933), .ZN(n8909) );
  NAND2_X1 U8717 ( .A1(n8903), .A2(n8905), .ZN(n8933) );
  NAND2_X1 U8718 ( .A1(n8934), .A2(n8935), .ZN(n8905) );
  NAND2_X1 U8719 ( .A1(n8936), .A2(n8932), .ZN(n8935) );
  NAND2_X1 U8720 ( .A1(n8937), .A2(n8938), .ZN(n8934) );
  NAND2_X1 U8721 ( .A1(n8900), .A2(n8939), .ZN(n8903) );
  NAND2_X1 U8722 ( .A1(n8897), .A2(n8899), .ZN(n8939) );
  NAND2_X1 U8723 ( .A1(n8940), .A2(n8941), .ZN(n8899) );
  XNOR2_X1 U8724 ( .A(n8937), .B(n8938), .ZN(n8940) );
  NAND2_X1 U8725 ( .A1(n8894), .A2(n8942), .ZN(n8897) );
  NAND2_X1 U8726 ( .A1(n8891), .A2(n8893), .ZN(n8942) );
  NAND2_X1 U8727 ( .A1(n8943), .A2(n8944), .ZN(n8893) );
  NAND2_X1 U8728 ( .A1(n8945), .A2(n8941), .ZN(n8944) );
  NAND2_X1 U8729 ( .A1(n8946), .A2(n8947), .ZN(n8943) );
  NAND2_X1 U8730 ( .A1(n8888), .A2(n8948), .ZN(n8891) );
  NAND2_X1 U8731 ( .A1(n8887), .A2(n8885), .ZN(n8948) );
  NAND2_X1 U8732 ( .A1(n8882), .A2(n8949), .ZN(n8885) );
  NAND2_X1 U8733 ( .A1(n8881), .A2(n8879), .ZN(n8949) );
  NAND2_X1 U8734 ( .A1(n8876), .A2(n8950), .ZN(n8879) );
  NAND2_X1 U8735 ( .A1(n8873), .A2(n8875), .ZN(n8950) );
  NAND2_X1 U8736 ( .A1(n8951), .A2(n8952), .ZN(n8875) );
  NAND2_X1 U8737 ( .A1(n8953), .A2(n8954), .ZN(n8952) );
  XNOR2_X1 U8738 ( .A(n8955), .B(n8956), .ZN(n8951) );
  NAND2_X1 U8739 ( .A1(n8870), .A2(n8957), .ZN(n8873) );
  NAND2_X1 U8740 ( .A1(n8869), .A2(n8867), .ZN(n8957) );
  NAND2_X1 U8741 ( .A1(n8863), .A2(n8958), .ZN(n8867) );
  NAND2_X1 U8742 ( .A1(n8861), .A2(n8864), .ZN(n8958) );
  NAND2_X1 U8743 ( .A1(n8959), .A2(n8960), .ZN(n8864) );
  NAND2_X1 U8744 ( .A1(n8961), .A2(n8962), .ZN(n8960) );
  XNOR2_X1 U8745 ( .A(n8963), .B(n8964), .ZN(n8959) );
  NAND2_X1 U8746 ( .A1(n8858), .A2(n8965), .ZN(n8861) );
  NAND2_X1 U8747 ( .A1(n8855), .A2(n8857), .ZN(n8965) );
  NAND2_X1 U8748 ( .A1(n8966), .A2(n8967), .ZN(n8857) );
  NAND2_X1 U8749 ( .A1(n8968), .A2(n8969), .ZN(n8967) );
  XNOR2_X1 U8750 ( .A(n8961), .B(n8962), .ZN(n8966) );
  NAND2_X1 U8751 ( .A1(n8845), .A2(n8970), .ZN(n8855) );
  NAND2_X1 U8752 ( .A1(n8843), .A2(n8846), .ZN(n8970) );
  NAND2_X1 U8753 ( .A1(n8971), .A2(n8972), .ZN(n8846) );
  XNOR2_X1 U8754 ( .A(n8969), .B(n8968), .ZN(n8971) );
  NAND2_X1 U8755 ( .A1(n8839), .A2(n8973), .ZN(n8843) );
  NAND2_X1 U8756 ( .A1(n8837), .A2(n8840), .ZN(n8973) );
  NAND2_X1 U8757 ( .A1(n8974), .A2(n8975), .ZN(n8840) );
  NAND2_X1 U8758 ( .A1(n8976), .A2(n8972), .ZN(n8975) );
  NAND2_X1 U8759 ( .A1(n8977), .A2(n8978), .ZN(n8974) );
  NAND2_X1 U8760 ( .A1(n8833), .A2(n8979), .ZN(n8837) );
  NAND2_X1 U8761 ( .A1(n8831), .A2(n8834), .ZN(n8979) );
  NAND2_X1 U8762 ( .A1(n8980), .A2(n8981), .ZN(n8834) );
  NAND2_X1 U8763 ( .A1(n8982), .A2(n8983), .ZN(n8981) );
  XNOR2_X1 U8764 ( .A(n8978), .B(n8977), .ZN(n8980) );
  NAND2_X1 U8765 ( .A1(n8828), .A2(n8984), .ZN(n8831) );
  NAND2_X1 U8766 ( .A1(n8825), .A2(n8827), .ZN(n8984) );
  NAND2_X1 U8767 ( .A1(n8985), .A2(n8986), .ZN(n8827) );
  NAND2_X1 U8768 ( .A1(n8987), .A2(n8988), .ZN(n8986) );
  XNOR2_X1 U8769 ( .A(n8983), .B(n8982), .ZN(n8985) );
  NAND2_X1 U8770 ( .A1(n8821), .A2(n8989), .ZN(n8825) );
  NAND2_X1 U8771 ( .A1(n8819), .A2(n8822), .ZN(n8989) );
  NAND2_X1 U8772 ( .A1(n8990), .A2(n8991), .ZN(n8822) );
  XOR2_X1 U8773 ( .A(n8988), .B(n8992), .Z(n8990) );
  NAND2_X1 U8774 ( .A1(n8815), .A2(n8993), .ZN(n8819) );
  NAND2_X1 U8775 ( .A1(n8813), .A2(n8816), .ZN(n8993) );
  NAND2_X1 U8776 ( .A1(n8994), .A2(n8995), .ZN(n8816) );
  NAND2_X1 U8777 ( .A1(n8996), .A2(n8991), .ZN(n8995) );
  NAND2_X1 U8778 ( .A1(n8997), .A2(n8998), .ZN(n8994) );
  NAND2_X1 U8779 ( .A1(n8810), .A2(n8999), .ZN(n8813) );
  NAND2_X1 U8780 ( .A1(n8809), .A2(n8807), .ZN(n8999) );
  NAND2_X1 U8781 ( .A1(n9000), .A2(n8803), .ZN(n8807) );
  OR2_X1 U8782 ( .A1(n9001), .A2(n9002), .ZN(n8803) );
  NAND2_X1 U8783 ( .A1(n8804), .A2(n8802), .ZN(n9000) );
  NAND2_X1 U8784 ( .A1(n9003), .A2(n8798), .ZN(n8802) );
  NAND4_X1 U8785 ( .A1(n9004), .A2(n9005), .A3(n9006), .A4(n9002), .ZN(n8798)
         );
  NAND2_X1 U8786 ( .A1(n9007), .A2(n9008), .ZN(n9005) );
  NAND2_X1 U8787 ( .A1(n8797), .A2(n8796), .ZN(n9003) );
  NAND2_X1 U8788 ( .A1(n8792), .A2(n9009), .ZN(n8796) );
  NAND2_X1 U8789 ( .A1(n9010), .A2(n8791), .ZN(n9009) );
  NAND2_X1 U8790 ( .A1(n9011), .A2(n9012), .ZN(n8791) );
  NAND2_X1 U8791 ( .A1(n8781), .A2(n8780), .ZN(n9012) );
  XOR2_X1 U8792 ( .A(n9006), .B(n9013), .Z(n9011) );
  INV_X1 U8793 ( .A(n8777), .ZN(n9010) );
  NAND3_X1 U8794 ( .A1(n9014), .A2(n8773), .A3(n8774), .ZN(n8777) );
  XNOR2_X1 U8795 ( .A(n9015), .B(n9016), .ZN(n8774) );
  XOR2_X1 U8796 ( .A(n9017), .B(n9018), .Z(n9016) );
  NAND2_X1 U8797 ( .A1(b_30_), .A2(a_0_), .ZN(n9018) );
  NAND2_X1 U8798 ( .A1(n9019), .A2(n9020), .ZN(n8773) );
  NAND3_X1 U8799 ( .A1(b_31_), .A2(n9021), .A3(a_0_), .ZN(n9020) );
  NAND2_X1 U8800 ( .A1(n8641), .A2(n8639), .ZN(n9021) );
  OR2_X1 U8801 ( .A1(n8639), .A2(n8641), .ZN(n9019) );
  AND2_X1 U8802 ( .A1(n9022), .A2(n9023), .ZN(n8641) );
  NAND3_X1 U8803 ( .A1(b_31_), .A2(n9024), .A3(a_1_), .ZN(n9023) );
  OR2_X1 U8804 ( .A1(n8615), .A2(n8614), .ZN(n9024) );
  NAND2_X1 U8805 ( .A1(n8614), .A2(n8615), .ZN(n9022) );
  NAND2_X1 U8806 ( .A1(n9025), .A2(n9026), .ZN(n8615) );
  NAND3_X1 U8807 ( .A1(b_31_), .A2(n9027), .A3(a_2_), .ZN(n9026) );
  NAND2_X1 U8808 ( .A1(n8590), .A2(n8588), .ZN(n9027) );
  OR2_X1 U8809 ( .A1(n8588), .A2(n8590), .ZN(n9025) );
  AND2_X1 U8810 ( .A1(n9028), .A2(n9029), .ZN(n8590) );
  NAND3_X1 U8811 ( .A1(b_31_), .A2(n9030), .A3(a_3_), .ZN(n9029) );
  OR2_X1 U8812 ( .A1(n8565), .A2(n8564), .ZN(n9030) );
  NAND2_X1 U8813 ( .A1(n8564), .A2(n8565), .ZN(n9028) );
  NAND2_X1 U8814 ( .A1(n9031), .A2(n9032), .ZN(n8565) );
  NAND3_X1 U8815 ( .A1(b_31_), .A2(n9033), .A3(a_4_), .ZN(n9032) );
  NAND2_X1 U8816 ( .A1(n8540), .A2(n8538), .ZN(n9033) );
  OR2_X1 U8817 ( .A1(n8538), .A2(n8540), .ZN(n9031) );
  AND2_X1 U8818 ( .A1(n9034), .A2(n9035), .ZN(n8540) );
  NAND3_X1 U8819 ( .A1(b_31_), .A2(n9036), .A3(a_5_), .ZN(n9035) );
  OR2_X1 U8820 ( .A1(n8515), .A2(n8514), .ZN(n9036) );
  NAND2_X1 U8821 ( .A1(n8514), .A2(n8515), .ZN(n9034) );
  NAND2_X1 U8822 ( .A1(n9037), .A2(n9038), .ZN(n8515) );
  NAND3_X1 U8823 ( .A1(b_31_), .A2(n9039), .A3(a_6_), .ZN(n9038) );
  OR2_X1 U8824 ( .A1(n8489), .A2(n8488), .ZN(n9039) );
  NAND2_X1 U8825 ( .A1(n8488), .A2(n8489), .ZN(n9037) );
  NAND2_X1 U8826 ( .A1(n9040), .A2(n9041), .ZN(n8489) );
  NAND3_X1 U8827 ( .A1(b_31_), .A2(n9042), .A3(a_7_), .ZN(n9041) );
  OR2_X1 U8828 ( .A1(n8464), .A2(n8462), .ZN(n9042) );
  NAND2_X1 U8829 ( .A1(n8462), .A2(n8464), .ZN(n9040) );
  NAND2_X1 U8830 ( .A1(n9043), .A2(n9044), .ZN(n8464) );
  NAND3_X1 U8831 ( .A1(b_31_), .A2(n9045), .A3(a_8_), .ZN(n9044) );
  NAND2_X1 U8832 ( .A1(n8433), .A2(n8431), .ZN(n9045) );
  OR2_X1 U8833 ( .A1(n8431), .A2(n8433), .ZN(n9043) );
  AND2_X1 U8834 ( .A1(n9046), .A2(n9047), .ZN(n8433) );
  NAND3_X1 U8835 ( .A1(b_31_), .A2(n9048), .A3(a_9_), .ZN(n9047) );
  NAND2_X1 U8836 ( .A1(n8408), .A2(n8406), .ZN(n9048) );
  OR2_X1 U8837 ( .A1(n8406), .A2(n8408), .ZN(n9046) );
  AND2_X1 U8838 ( .A1(n9049), .A2(n9050), .ZN(n8408) );
  NAND3_X1 U8839 ( .A1(b_31_), .A2(n9051), .A3(a_10_), .ZN(n9050) );
  NAND2_X1 U8840 ( .A1(n8383), .A2(n8381), .ZN(n9051) );
  OR2_X1 U8841 ( .A1(n8381), .A2(n8383), .ZN(n9049) );
  AND2_X1 U8842 ( .A1(n9052), .A2(n9053), .ZN(n8383) );
  NAND3_X1 U8843 ( .A1(b_31_), .A2(n9054), .A3(a_11_), .ZN(n9053) );
  OR2_X1 U8844 ( .A1(n8358), .A2(n8356), .ZN(n9054) );
  NAND2_X1 U8845 ( .A1(n8356), .A2(n8358), .ZN(n9052) );
  NAND2_X1 U8846 ( .A1(n9055), .A2(n9056), .ZN(n8358) );
  NAND3_X1 U8847 ( .A1(b_31_), .A2(n9057), .A3(a_12_), .ZN(n9056) );
  NAND2_X1 U8848 ( .A1(n8333), .A2(n8331), .ZN(n9057) );
  OR2_X1 U8849 ( .A1(n8331), .A2(n8333), .ZN(n9055) );
  AND2_X1 U8850 ( .A1(n9058), .A2(n9059), .ZN(n8333) );
  NAND3_X1 U8851 ( .A1(b_31_), .A2(n9060), .A3(a_13_), .ZN(n9059) );
  OR2_X1 U8852 ( .A1(n8308), .A2(n8307), .ZN(n9060) );
  NAND2_X1 U8853 ( .A1(n8307), .A2(n8308), .ZN(n9058) );
  NAND2_X1 U8854 ( .A1(n9061), .A2(n9062), .ZN(n8308) );
  NAND3_X1 U8855 ( .A1(b_31_), .A2(n9063), .A3(a_14_), .ZN(n9062) );
  NAND2_X1 U8856 ( .A1(n8283), .A2(n8281), .ZN(n9063) );
  OR2_X1 U8857 ( .A1(n8281), .A2(n8283), .ZN(n9061) );
  AND2_X1 U8858 ( .A1(n9064), .A2(n9065), .ZN(n8283) );
  NAND3_X1 U8859 ( .A1(b_31_), .A2(n9066), .A3(a_15_), .ZN(n9065) );
  OR2_X1 U8860 ( .A1(n8258), .A2(n8256), .ZN(n9066) );
  NAND2_X1 U8861 ( .A1(n8256), .A2(n8258), .ZN(n9064) );
  NAND2_X1 U8862 ( .A1(n9067), .A2(n9068), .ZN(n8258) );
  NAND3_X1 U8863 ( .A1(b_31_), .A2(n9069), .A3(a_16_), .ZN(n9068) );
  NAND2_X1 U8864 ( .A1(n8233), .A2(n8231), .ZN(n9069) );
  OR2_X1 U8865 ( .A1(n8231), .A2(n8233), .ZN(n9067) );
  AND2_X1 U8866 ( .A1(n9070), .A2(n9071), .ZN(n8233) );
  NAND3_X1 U8867 ( .A1(b_31_), .A2(n9072), .A3(a_17_), .ZN(n9071) );
  OR2_X1 U8868 ( .A1(n8208), .A2(n8207), .ZN(n9072) );
  NAND2_X1 U8869 ( .A1(n8207), .A2(n8208), .ZN(n9070) );
  NAND2_X1 U8870 ( .A1(n9073), .A2(n9074), .ZN(n8208) );
  NAND3_X1 U8871 ( .A1(b_31_), .A2(n9075), .A3(a_18_), .ZN(n9074) );
  NAND2_X1 U8872 ( .A1(n8177), .A2(n8175), .ZN(n9075) );
  OR2_X1 U8873 ( .A1(n8175), .A2(n8177), .ZN(n9073) );
  AND2_X1 U8874 ( .A1(n9076), .A2(n9077), .ZN(n8177) );
  NAND3_X1 U8875 ( .A1(b_31_), .A2(n9078), .A3(a_19_), .ZN(n9077) );
  OR2_X1 U8876 ( .A1(n8152), .A2(n8150), .ZN(n9078) );
  NAND2_X1 U8877 ( .A1(n8150), .A2(n8152), .ZN(n9076) );
  NAND2_X1 U8878 ( .A1(n9079), .A2(n9080), .ZN(n8152) );
  NAND3_X1 U8879 ( .A1(b_31_), .A2(n9081), .A3(a_20_), .ZN(n9080) );
  NAND2_X1 U8880 ( .A1(n8127), .A2(n8125), .ZN(n9081) );
  OR2_X1 U8881 ( .A1(n8125), .A2(n8127), .ZN(n9079) );
  AND2_X1 U8882 ( .A1(n9082), .A2(n9083), .ZN(n8127) );
  NAND3_X1 U8883 ( .A1(b_31_), .A2(n9084), .A3(a_21_), .ZN(n9083) );
  NAND2_X1 U8884 ( .A1(n8101), .A2(n8099), .ZN(n9084) );
  OR2_X1 U8885 ( .A1(n8099), .A2(n8101), .ZN(n9082) );
  AND2_X1 U8886 ( .A1(n9085), .A2(n9086), .ZN(n8101) );
  NAND3_X1 U8887 ( .A1(b_31_), .A2(n9087), .A3(a_22_), .ZN(n9086) );
  NAND2_X1 U8888 ( .A1(n8076), .A2(n8074), .ZN(n9087) );
  OR2_X1 U8889 ( .A1(n8074), .A2(n8076), .ZN(n9085) );
  AND2_X1 U8890 ( .A1(n8050), .A2(n9088), .ZN(n8076) );
  NAND2_X1 U8891 ( .A1(n8049), .A2(n8051), .ZN(n9088) );
  NAND2_X1 U8892 ( .A1(n9089), .A2(n9090), .ZN(n8051) );
  NAND2_X1 U8893 ( .A1(a_23_), .A2(b_31_), .ZN(n9090) );
  INV_X1 U8894 ( .A(n9091), .ZN(n9089) );
  XOR2_X1 U8895 ( .A(n9092), .B(n9093), .Z(n8049) );
  XOR2_X1 U8896 ( .A(n9094), .B(n9095), .Z(n9092) );
  NOR2_X1 U8897 ( .A1(n8745), .A2(n7869), .ZN(n9095) );
  NAND2_X1 U8898 ( .A1(a_23_), .A2(n9091), .ZN(n8050) );
  NAND2_X1 U8899 ( .A1(n9096), .A2(n9097), .ZN(n9091) );
  NAND2_X1 U8900 ( .A1(n8023), .A2(n9098), .ZN(n9097) );
  OR2_X1 U8901 ( .A1(n8025), .A2(n8026), .ZN(n9098) );
  XOR2_X1 U8902 ( .A(n9099), .B(n9100), .Z(n8023) );
  XOR2_X1 U8903 ( .A(n9101), .B(n9102), .Z(n9099) );
  NAND2_X1 U8904 ( .A1(n8026), .A2(n8025), .ZN(n9096) );
  NAND2_X1 U8905 ( .A1(n7999), .A2(n9103), .ZN(n8025) );
  NAND2_X1 U8906 ( .A1(n7998), .A2(n8000), .ZN(n9103) );
  NAND2_X1 U8907 ( .A1(n9104), .A2(n9105), .ZN(n8000) );
  NAND2_X1 U8908 ( .A1(a_25_), .A2(b_31_), .ZN(n9105) );
  INV_X1 U8909 ( .A(n9106), .ZN(n9104) );
  XNOR2_X1 U8910 ( .A(n9107), .B(n9108), .ZN(n7998) );
  NAND2_X1 U8911 ( .A1(n9109), .A2(n9110), .ZN(n9107) );
  NAND2_X1 U8912 ( .A1(a_25_), .A2(n9106), .ZN(n7999) );
  NAND2_X1 U8913 ( .A1(n9111), .A2(n9112), .ZN(n9106) );
  NAND2_X1 U8914 ( .A1(n7973), .A2(n9113), .ZN(n9112) );
  OR2_X1 U8915 ( .A1(n7974), .A2(n7975), .ZN(n9113) );
  XNOR2_X1 U8916 ( .A(n9114), .B(n9115), .ZN(n7973) );
  NAND2_X1 U8917 ( .A1(n9116), .A2(n9117), .ZN(n9114) );
  NAND2_X1 U8918 ( .A1(n7975), .A2(n7974), .ZN(n9111) );
  NAND2_X1 U8919 ( .A1(n7948), .A2(n9118), .ZN(n7974) );
  NAND2_X1 U8920 ( .A1(n7947), .A2(n7949), .ZN(n9118) );
  NAND2_X1 U8921 ( .A1(n9119), .A2(n9120), .ZN(n7949) );
  NAND2_X1 U8922 ( .A1(a_27_), .A2(b_31_), .ZN(n9120) );
  INV_X1 U8923 ( .A(n9121), .ZN(n9119) );
  XNOR2_X1 U8924 ( .A(n9122), .B(n9123), .ZN(n7947) );
  XOR2_X1 U8925 ( .A(n9124), .B(n9125), .Z(n9122) );
  NAND2_X1 U8926 ( .A1(b_30_), .A2(a_28_), .ZN(n9124) );
  NAND2_X1 U8927 ( .A1(a_27_), .A2(n9121), .ZN(n7948) );
  NAND2_X1 U8928 ( .A1(n9126), .A2(n9127), .ZN(n9121) );
  NAND2_X1 U8929 ( .A1(n7918), .A2(n9128), .ZN(n9127) );
  NAND2_X1 U8930 ( .A1(n7917), .A2(n7915), .ZN(n9128) );
  NOR2_X1 U8931 ( .A1(n8739), .A2(n7889), .ZN(n7918) );
  OR2_X1 U8932 ( .A1(n7915), .A2(n7917), .ZN(n9126) );
  AND2_X1 U8933 ( .A1(n9129), .A2(n9130), .ZN(n7917) );
  NAND3_X1 U8934 ( .A1(b_31_), .A2(n9131), .A3(a_29_), .ZN(n9130) );
  OR2_X1 U8935 ( .A1(n7891), .A2(n7892), .ZN(n9131) );
  NAND2_X1 U8936 ( .A1(n7892), .A2(n7891), .ZN(n9129) );
  NAND2_X1 U8937 ( .A1(n9132), .A2(n9133), .ZN(n7891) );
  NAND2_X1 U8938 ( .A1(b_29_), .A2(n9134), .ZN(n9133) );
  NAND2_X1 U8939 ( .A1(n7864), .A2(n9135), .ZN(n9134) );
  NAND2_X1 U8940 ( .A1(a_31_), .A2(n7869), .ZN(n9135) );
  NAND2_X1 U8941 ( .A1(b_30_), .A2(n9136), .ZN(n9132) );
  NAND2_X1 U8942 ( .A1(n9137), .A2(n9138), .ZN(n9136) );
  NAND2_X1 U8943 ( .A1(a_30_), .A2(n8738), .ZN(n9138) );
  AND3_X1 U8944 ( .A1(b_30_), .A2(b_31_), .A3(n7818), .ZN(n7892) );
  XNOR2_X1 U8945 ( .A(n9139), .B(n9140), .ZN(n7915) );
  XOR2_X1 U8946 ( .A(n9141), .B(n9142), .Z(n9139) );
  NOR2_X1 U8947 ( .A1(n8742), .A2(n7889), .ZN(n7975) );
  NOR2_X1 U8948 ( .A1(n8745), .A2(n7889), .ZN(n8026) );
  XOR2_X1 U8949 ( .A(n9143), .B(n9144), .Z(n8074) );
  XNOR2_X1 U8950 ( .A(n9145), .B(n9146), .ZN(n9144) );
  XNOR2_X1 U8951 ( .A(n9147), .B(n9148), .ZN(n8099) );
  XOR2_X1 U8952 ( .A(n9149), .B(n9150), .Z(n9147) );
  NOR2_X1 U8953 ( .A1(n8748), .A2(n7869), .ZN(n9150) );
  XNOR2_X1 U8954 ( .A(n9151), .B(n9152), .ZN(n8125) );
  XOR2_X1 U8955 ( .A(n9153), .B(n9154), .Z(n9151) );
  XNOR2_X1 U8956 ( .A(n9155), .B(n9156), .ZN(n8150) );
  XNOR2_X1 U8957 ( .A(n9157), .B(n9158), .ZN(n9155) );
  NOR2_X1 U8958 ( .A1(n8751), .A2(n7869), .ZN(n9158) );
  XOR2_X1 U8959 ( .A(n9159), .B(n9160), .Z(n8175) );
  XNOR2_X1 U8960 ( .A(n9161), .B(n9162), .ZN(n9160) );
  XNOR2_X1 U8961 ( .A(n9163), .B(n9164), .ZN(n8207) );
  XNOR2_X1 U8962 ( .A(n9165), .B(n9166), .ZN(n9163) );
  NOR2_X1 U8963 ( .A1(n8753), .A2(n7869), .ZN(n9166) );
  XNOR2_X1 U8964 ( .A(n9167), .B(n9168), .ZN(n8231) );
  XOR2_X1 U8965 ( .A(n9169), .B(n9170), .Z(n9167) );
  XNOR2_X1 U8966 ( .A(n9171), .B(n9172), .ZN(n8256) );
  XNOR2_X1 U8967 ( .A(n9173), .B(n9174), .ZN(n9171) );
  NOR2_X1 U8968 ( .A1(n8755), .A2(n7869), .ZN(n9174) );
  XOR2_X1 U8969 ( .A(n9175), .B(n9176), .Z(n8281) );
  XNOR2_X1 U8970 ( .A(n9177), .B(n9178), .ZN(n9176) );
  XNOR2_X1 U8971 ( .A(n9179), .B(n9180), .ZN(n8307) );
  XOR2_X1 U8972 ( .A(n9181), .B(n9182), .Z(n9179) );
  NAND2_X1 U8973 ( .A1(b_30_), .A2(a_14_), .ZN(n9181) );
  XNOR2_X1 U8974 ( .A(n9183), .B(n9184), .ZN(n8331) );
  XOR2_X1 U8975 ( .A(n9185), .B(n9186), .Z(n9183) );
  XNOR2_X1 U8976 ( .A(n9187), .B(n9188), .ZN(n8356) );
  XNOR2_X1 U8977 ( .A(n9189), .B(n9190), .ZN(n9187) );
  NOR2_X1 U8978 ( .A1(n8759), .A2(n7869), .ZN(n9190) );
  XOR2_X1 U8979 ( .A(n9191), .B(n9192), .Z(n8381) );
  XNOR2_X1 U8980 ( .A(n9193), .B(n9194), .ZN(n9192) );
  XNOR2_X1 U8981 ( .A(n9195), .B(n9196), .ZN(n8406) );
  XOR2_X1 U8982 ( .A(n9197), .B(n9198), .Z(n9195) );
  NOR2_X1 U8983 ( .A1(n8761), .A2(n7869), .ZN(n9198) );
  XNOR2_X1 U8984 ( .A(n9199), .B(n9200), .ZN(n8431) );
  XOR2_X1 U8985 ( .A(n9201), .B(n9202), .Z(n9199) );
  XNOR2_X1 U8986 ( .A(n9203), .B(n9204), .ZN(n8462) );
  XOR2_X1 U8987 ( .A(n9205), .B(n9206), .Z(n9204) );
  NAND2_X1 U8988 ( .A1(b_30_), .A2(a_8_), .ZN(n9206) );
  XNOR2_X1 U8989 ( .A(n9207), .B(n9208), .ZN(n8488) );
  XNOR2_X1 U8990 ( .A(n9209), .B(n9210), .ZN(n9208) );
  XNOR2_X1 U8991 ( .A(n9211), .B(n9212), .ZN(n8514) );
  XNOR2_X1 U8992 ( .A(n9213), .B(n9214), .ZN(n9211) );
  NOR2_X1 U8993 ( .A1(n8491), .A2(n7869), .ZN(n9214) );
  XOR2_X1 U8994 ( .A(n9215), .B(n9216), .Z(n8538) );
  XNOR2_X1 U8995 ( .A(n9217), .B(n9218), .ZN(n9216) );
  XNOR2_X1 U8996 ( .A(n9219), .B(n9220), .ZN(n8564) );
  XNOR2_X1 U8997 ( .A(n9221), .B(n9222), .ZN(n9219) );
  NOR2_X1 U8998 ( .A1(n8766), .A2(n7869), .ZN(n9222) );
  XOR2_X1 U8999 ( .A(n9223), .B(n9224), .Z(n8588) );
  XNOR2_X1 U9000 ( .A(n9225), .B(n9226), .ZN(n9224) );
  XNOR2_X1 U9001 ( .A(n9227), .B(n9228), .ZN(n8614) );
  XNOR2_X1 U9002 ( .A(n9229), .B(n9230), .ZN(n9227) );
  NOR2_X1 U9003 ( .A1(n8768), .A2(n7869), .ZN(n9230) );
  XNOR2_X1 U9004 ( .A(n9231), .B(n9232), .ZN(n8639) );
  XOR2_X1 U9005 ( .A(n9233), .B(n9234), .Z(n9231) );
  NOR2_X1 U9006 ( .A1(n8617), .A2(n7869), .ZN(n9234) );
  XOR2_X1 U9007 ( .A(n8780), .B(n8781), .Z(n9014) );
  NAND3_X1 U9008 ( .A1(n8781), .A2(n8780), .A3(n9235), .ZN(n8792) );
  XOR2_X1 U9009 ( .A(n9004), .B(n9006), .Z(n9235) );
  NAND2_X1 U9010 ( .A1(n9236), .A2(n9237), .ZN(n8780) );
  NAND3_X1 U9011 ( .A1(a_0_), .A2(n9238), .A3(b_30_), .ZN(n9237) );
  OR2_X1 U9012 ( .A1(n9017), .A2(n9015), .ZN(n9238) );
  NAND2_X1 U9013 ( .A1(n9015), .A2(n9017), .ZN(n9236) );
  NAND2_X1 U9014 ( .A1(n9239), .A2(n9240), .ZN(n9017) );
  NAND3_X1 U9015 ( .A1(a_1_), .A2(n9241), .A3(b_30_), .ZN(n9240) );
  OR2_X1 U9016 ( .A1(n9233), .A2(n9232), .ZN(n9241) );
  NAND2_X1 U9017 ( .A1(n9232), .A2(n9233), .ZN(n9239) );
  NAND2_X1 U9018 ( .A1(n9242), .A2(n9243), .ZN(n9233) );
  NAND3_X1 U9019 ( .A1(a_2_), .A2(n9244), .A3(b_30_), .ZN(n9243) );
  NAND2_X1 U9020 ( .A1(n9229), .A2(n9228), .ZN(n9244) );
  OR2_X1 U9021 ( .A1(n9228), .A2(n9229), .ZN(n9242) );
  AND2_X1 U9022 ( .A1(n9245), .A2(n9246), .ZN(n9229) );
  NAND2_X1 U9023 ( .A1(n9226), .A2(n9247), .ZN(n9246) );
  OR2_X1 U9024 ( .A1(n9225), .A2(n9223), .ZN(n9247) );
  NOR2_X1 U9025 ( .A1(n7869), .A2(n8567), .ZN(n9226) );
  NAND2_X1 U9026 ( .A1(n9223), .A2(n9225), .ZN(n9245) );
  NAND2_X1 U9027 ( .A1(n9248), .A2(n9249), .ZN(n9225) );
  NAND3_X1 U9028 ( .A1(a_4_), .A2(n9250), .A3(b_30_), .ZN(n9249) );
  NAND2_X1 U9029 ( .A1(n9221), .A2(n9220), .ZN(n9250) );
  OR2_X1 U9030 ( .A1(n9220), .A2(n9221), .ZN(n9248) );
  AND2_X1 U9031 ( .A1(n9251), .A2(n9252), .ZN(n9221) );
  NAND2_X1 U9032 ( .A1(n9218), .A2(n9253), .ZN(n9252) );
  OR2_X1 U9033 ( .A1(n9217), .A2(n9215), .ZN(n9253) );
  NOR2_X1 U9034 ( .A1(n7869), .A2(n8517), .ZN(n9218) );
  NAND2_X1 U9035 ( .A1(n9215), .A2(n9217), .ZN(n9251) );
  NAND2_X1 U9036 ( .A1(n9254), .A2(n9255), .ZN(n9217) );
  NAND3_X1 U9037 ( .A1(a_6_), .A2(n9256), .A3(b_30_), .ZN(n9255) );
  NAND2_X1 U9038 ( .A1(n9213), .A2(n9212), .ZN(n9256) );
  OR2_X1 U9039 ( .A1(n9212), .A2(n9213), .ZN(n9254) );
  AND2_X1 U9040 ( .A1(n9257), .A2(n9258), .ZN(n9213) );
  NAND2_X1 U9041 ( .A1(n9210), .A2(n9259), .ZN(n9258) );
  OR2_X1 U9042 ( .A1(n9209), .A2(n9207), .ZN(n9259) );
  NOR2_X1 U9043 ( .A1(n7869), .A2(n8764), .ZN(n9210) );
  NAND2_X1 U9044 ( .A1(n9207), .A2(n9209), .ZN(n9257) );
  NAND2_X1 U9045 ( .A1(n9260), .A2(n9261), .ZN(n9209) );
  NAND3_X1 U9046 ( .A1(a_8_), .A2(n9262), .A3(b_30_), .ZN(n9261) );
  OR2_X1 U9047 ( .A1(n9205), .A2(n9203), .ZN(n9262) );
  NAND2_X1 U9048 ( .A1(n9203), .A2(n9205), .ZN(n9260) );
  NAND2_X1 U9049 ( .A1(n9263), .A2(n9264), .ZN(n9205) );
  NAND2_X1 U9050 ( .A1(n9202), .A2(n9265), .ZN(n9264) );
  OR2_X1 U9051 ( .A1(n9201), .A2(n9200), .ZN(n9265) );
  NOR2_X1 U9052 ( .A1(n7869), .A2(n8426), .ZN(n9202) );
  NAND2_X1 U9053 ( .A1(n9200), .A2(n9201), .ZN(n9263) );
  NAND2_X1 U9054 ( .A1(n9266), .A2(n9267), .ZN(n9201) );
  NAND3_X1 U9055 ( .A1(a_10_), .A2(n9268), .A3(b_30_), .ZN(n9267) );
  OR2_X1 U9056 ( .A1(n9197), .A2(n9196), .ZN(n9268) );
  NAND2_X1 U9057 ( .A1(n9196), .A2(n9197), .ZN(n9266) );
  NAND2_X1 U9058 ( .A1(n9269), .A2(n9270), .ZN(n9197) );
  NAND2_X1 U9059 ( .A1(n9194), .A2(n9271), .ZN(n9270) );
  OR2_X1 U9060 ( .A1(n9193), .A2(n9191), .ZN(n9271) );
  NOR2_X1 U9061 ( .A1(n7869), .A2(n8376), .ZN(n9194) );
  NAND2_X1 U9062 ( .A1(n9191), .A2(n9193), .ZN(n9269) );
  NAND2_X1 U9063 ( .A1(n9272), .A2(n9273), .ZN(n9193) );
  NAND3_X1 U9064 ( .A1(a_12_), .A2(n9274), .A3(b_30_), .ZN(n9273) );
  NAND2_X1 U9065 ( .A1(n9189), .A2(n9188), .ZN(n9274) );
  OR2_X1 U9066 ( .A1(n9188), .A2(n9189), .ZN(n9272) );
  AND2_X1 U9067 ( .A1(n9275), .A2(n9276), .ZN(n9189) );
  NAND2_X1 U9068 ( .A1(n9186), .A2(n9277), .ZN(n9276) );
  OR2_X1 U9069 ( .A1(n9185), .A2(n9184), .ZN(n9277) );
  NOR2_X1 U9070 ( .A1(n7869), .A2(n8310), .ZN(n9186) );
  NAND2_X1 U9071 ( .A1(n9184), .A2(n9185), .ZN(n9275) );
  NAND2_X1 U9072 ( .A1(n9278), .A2(n9279), .ZN(n9185) );
  NAND3_X1 U9073 ( .A1(a_14_), .A2(n9280), .A3(b_30_), .ZN(n9279) );
  NAND2_X1 U9074 ( .A1(n9182), .A2(n9180), .ZN(n9280) );
  OR2_X1 U9075 ( .A1(n9180), .A2(n9182), .ZN(n9278) );
  AND2_X1 U9076 ( .A1(n9281), .A2(n9282), .ZN(n9182) );
  NAND2_X1 U9077 ( .A1(n9178), .A2(n9283), .ZN(n9282) );
  OR2_X1 U9078 ( .A1(n9177), .A2(n9175), .ZN(n9283) );
  NOR2_X1 U9079 ( .A1(n7869), .A2(n8276), .ZN(n9178) );
  NAND2_X1 U9080 ( .A1(n9175), .A2(n9177), .ZN(n9281) );
  NAND2_X1 U9081 ( .A1(n9284), .A2(n9285), .ZN(n9177) );
  NAND3_X1 U9082 ( .A1(a_16_), .A2(n9286), .A3(b_30_), .ZN(n9285) );
  NAND2_X1 U9083 ( .A1(n9173), .A2(n9172), .ZN(n9286) );
  OR2_X1 U9084 ( .A1(n9172), .A2(n9173), .ZN(n9284) );
  AND2_X1 U9085 ( .A1(n9287), .A2(n9288), .ZN(n9173) );
  NAND2_X1 U9086 ( .A1(n9170), .A2(n9289), .ZN(n9288) );
  OR2_X1 U9087 ( .A1(n9169), .A2(n9168), .ZN(n9289) );
  NOR2_X1 U9088 ( .A1(n7869), .A2(n8210), .ZN(n9170) );
  NAND2_X1 U9089 ( .A1(n9168), .A2(n9169), .ZN(n9287) );
  NAND2_X1 U9090 ( .A1(n9290), .A2(n9291), .ZN(n9169) );
  NAND3_X1 U9091 ( .A1(a_18_), .A2(n9292), .A3(b_30_), .ZN(n9291) );
  NAND2_X1 U9092 ( .A1(n9165), .A2(n9164), .ZN(n9292) );
  OR2_X1 U9093 ( .A1(n9164), .A2(n9165), .ZN(n9290) );
  AND2_X1 U9094 ( .A1(n9293), .A2(n9294), .ZN(n9165) );
  NAND2_X1 U9095 ( .A1(n9162), .A2(n9295), .ZN(n9294) );
  OR2_X1 U9096 ( .A1(n9161), .A2(n9159), .ZN(n9295) );
  NOR2_X1 U9097 ( .A1(n7869), .A2(n8170), .ZN(n9162) );
  NAND2_X1 U9098 ( .A1(n9159), .A2(n9161), .ZN(n9293) );
  NAND2_X1 U9099 ( .A1(n9296), .A2(n9297), .ZN(n9161) );
  NAND3_X1 U9100 ( .A1(a_20_), .A2(n9298), .A3(b_30_), .ZN(n9297) );
  NAND2_X1 U9101 ( .A1(n9157), .A2(n9156), .ZN(n9298) );
  OR2_X1 U9102 ( .A1(n9156), .A2(n9157), .ZN(n9296) );
  AND2_X1 U9103 ( .A1(n9299), .A2(n9300), .ZN(n9157) );
  NAND2_X1 U9104 ( .A1(n9154), .A2(n9301), .ZN(n9300) );
  OR2_X1 U9105 ( .A1(n9153), .A2(n9152), .ZN(n9301) );
  NOR2_X1 U9106 ( .A1(n7869), .A2(n8750), .ZN(n9154) );
  NAND2_X1 U9107 ( .A1(n9152), .A2(n9153), .ZN(n9299) );
  NAND2_X1 U9108 ( .A1(n9302), .A2(n9303), .ZN(n9153) );
  NAND3_X1 U9109 ( .A1(a_22_), .A2(n9304), .A3(b_30_), .ZN(n9303) );
  OR2_X1 U9110 ( .A1(n9149), .A2(n9148), .ZN(n9304) );
  NAND2_X1 U9111 ( .A1(n9148), .A2(n9149), .ZN(n9302) );
  NAND2_X1 U9112 ( .A1(n9305), .A2(n9306), .ZN(n9149) );
  NAND2_X1 U9113 ( .A1(n9146), .A2(n9307), .ZN(n9306) );
  OR2_X1 U9114 ( .A1(n9145), .A2(n9143), .ZN(n9307) );
  NOR2_X1 U9115 ( .A1(n7869), .A2(n8747), .ZN(n9146) );
  NAND2_X1 U9116 ( .A1(n9143), .A2(n9145), .ZN(n9305) );
  NAND2_X1 U9117 ( .A1(n9308), .A2(n9309), .ZN(n9145) );
  NAND3_X1 U9118 ( .A1(a_24_), .A2(n9310), .A3(b_30_), .ZN(n9309) );
  OR2_X1 U9119 ( .A1(n9094), .A2(n9093), .ZN(n9310) );
  NAND2_X1 U9120 ( .A1(n9093), .A2(n9094), .ZN(n9308) );
  NAND2_X1 U9121 ( .A1(n9311), .A2(n9312), .ZN(n9094) );
  NAND2_X1 U9122 ( .A1(n9102), .A2(n9313), .ZN(n9312) );
  OR2_X1 U9123 ( .A1(n9101), .A2(n9100), .ZN(n9313) );
  NOR2_X1 U9124 ( .A1(n7869), .A2(n8744), .ZN(n9102) );
  NAND2_X1 U9125 ( .A1(n9100), .A2(n9101), .ZN(n9311) );
  NAND2_X1 U9126 ( .A1(n9109), .A2(n9314), .ZN(n9101) );
  NAND2_X1 U9127 ( .A1(n9108), .A2(n9110), .ZN(n9314) );
  NAND2_X1 U9128 ( .A1(n9315), .A2(n9316), .ZN(n9110) );
  NAND2_X1 U9129 ( .A1(b_30_), .A2(a_26_), .ZN(n9316) );
  INV_X1 U9130 ( .A(n9317), .ZN(n9315) );
  XNOR2_X1 U9131 ( .A(n9318), .B(n9319), .ZN(n9108) );
  NAND2_X1 U9132 ( .A1(n9320), .A2(n9321), .ZN(n9318) );
  NAND2_X1 U9133 ( .A1(a_26_), .A2(n9317), .ZN(n9109) );
  NAND2_X1 U9134 ( .A1(n9116), .A2(n9322), .ZN(n9317) );
  NAND2_X1 U9135 ( .A1(n9115), .A2(n9117), .ZN(n9322) );
  NAND2_X1 U9136 ( .A1(n9323), .A2(n9324), .ZN(n9117) );
  NAND2_X1 U9137 ( .A1(b_30_), .A2(a_27_), .ZN(n9324) );
  INV_X1 U9138 ( .A(n9325), .ZN(n9323) );
  XNOR2_X1 U9139 ( .A(n9326), .B(n9327), .ZN(n9115) );
  XOR2_X1 U9140 ( .A(n9328), .B(n9329), .Z(n9326) );
  NAND2_X1 U9141 ( .A1(b_29_), .A2(a_28_), .ZN(n9328) );
  NAND2_X1 U9142 ( .A1(a_27_), .A2(n9325), .ZN(n9116) );
  NAND2_X1 U9143 ( .A1(n9330), .A2(n9331), .ZN(n9325) );
  NAND3_X1 U9144 ( .A1(a_28_), .A2(n9332), .A3(b_30_), .ZN(n9331) );
  NAND2_X1 U9145 ( .A1(n9125), .A2(n9123), .ZN(n9332) );
  OR2_X1 U9146 ( .A1(n9123), .A2(n9125), .ZN(n9330) );
  AND2_X1 U9147 ( .A1(n9333), .A2(n9334), .ZN(n9125) );
  NAND2_X1 U9148 ( .A1(n9140), .A2(n9335), .ZN(n9334) );
  OR2_X1 U9149 ( .A1(n9141), .A2(n9142), .ZN(n9335) );
  NOR2_X1 U9150 ( .A1(n7869), .A2(n7890), .ZN(n9140) );
  NAND2_X1 U9151 ( .A1(n9142), .A2(n9141), .ZN(n9333) );
  NAND2_X1 U9152 ( .A1(n9336), .A2(n9337), .ZN(n9141) );
  NAND2_X1 U9153 ( .A1(b_28_), .A2(n9338), .ZN(n9337) );
  NAND2_X1 U9154 ( .A1(n7864), .A2(n9339), .ZN(n9338) );
  NAND2_X1 U9155 ( .A1(a_31_), .A2(n8738), .ZN(n9339) );
  NAND2_X1 U9156 ( .A1(b_29_), .A2(n9340), .ZN(n9336) );
  NAND2_X1 U9157 ( .A1(n9137), .A2(n9341), .ZN(n9340) );
  NAND2_X1 U9158 ( .A1(a_30_), .A2(n7935), .ZN(n9341) );
  AND3_X1 U9159 ( .A1(b_29_), .A2(b_30_), .A3(n7818), .ZN(n9142) );
  XNOR2_X1 U9160 ( .A(n9342), .B(n9343), .ZN(n9123) );
  XOR2_X1 U9161 ( .A(n9344), .B(n9345), .Z(n9342) );
  XNOR2_X1 U9162 ( .A(n9346), .B(n9347), .ZN(n9100) );
  NAND2_X1 U9163 ( .A1(n9348), .A2(n9349), .ZN(n9346) );
  XNOR2_X1 U9164 ( .A(n9350), .B(n9351), .ZN(n9093) );
  XNOR2_X1 U9165 ( .A(n9352), .B(n9353), .ZN(n9350) );
  XNOR2_X1 U9166 ( .A(n9354), .B(n9355), .ZN(n9143) );
  XOR2_X1 U9167 ( .A(n9356), .B(n9357), .Z(n9355) );
  NAND2_X1 U9168 ( .A1(b_29_), .A2(a_24_), .ZN(n9357) );
  XNOR2_X1 U9169 ( .A(n9358), .B(n9359), .ZN(n9148) );
  XNOR2_X1 U9170 ( .A(n9360), .B(n9361), .ZN(n9359) );
  XNOR2_X1 U9171 ( .A(n9362), .B(n9363), .ZN(n9152) );
  XOR2_X1 U9172 ( .A(n9364), .B(n9365), .Z(n9363) );
  NAND2_X1 U9173 ( .A1(b_29_), .A2(a_22_), .ZN(n9365) );
  XNOR2_X1 U9174 ( .A(n9366), .B(n9367), .ZN(n9156) );
  XOR2_X1 U9175 ( .A(n9368), .B(n9369), .Z(n9366) );
  XNOR2_X1 U9176 ( .A(n9370), .B(n9371), .ZN(n9159) );
  XNOR2_X1 U9177 ( .A(n9372), .B(n9373), .ZN(n9370) );
  NOR2_X1 U9178 ( .A1(n8751), .A2(n8738), .ZN(n9373) );
  XOR2_X1 U9179 ( .A(n9374), .B(n9375), .Z(n9164) );
  XNOR2_X1 U9180 ( .A(n9376), .B(n9377), .ZN(n9375) );
  XNOR2_X1 U9181 ( .A(n9378), .B(n9379), .ZN(n9168) );
  XNOR2_X1 U9182 ( .A(n9380), .B(n9381), .ZN(n9378) );
  NOR2_X1 U9183 ( .A1(n8753), .A2(n8738), .ZN(n9381) );
  XNOR2_X1 U9184 ( .A(n9382), .B(n9383), .ZN(n9172) );
  XOR2_X1 U9185 ( .A(n9384), .B(n9385), .Z(n9382) );
  XNOR2_X1 U9186 ( .A(n9386), .B(n9387), .ZN(n9175) );
  XOR2_X1 U9187 ( .A(n9388), .B(n9389), .Z(n9387) );
  NAND2_X1 U9188 ( .A1(b_29_), .A2(a_16_), .ZN(n9389) );
  XOR2_X1 U9189 ( .A(n9390), .B(n9391), .Z(n9180) );
  XNOR2_X1 U9190 ( .A(n9392), .B(n9393), .ZN(n9391) );
  XNOR2_X1 U9191 ( .A(n9394), .B(n9395), .ZN(n9184) );
  XOR2_X1 U9192 ( .A(n9396), .B(n9397), .Z(n9394) );
  NAND2_X1 U9193 ( .A1(b_29_), .A2(a_14_), .ZN(n9396) );
  XNOR2_X1 U9194 ( .A(n9398), .B(n9399), .ZN(n9188) );
  XOR2_X1 U9195 ( .A(n9400), .B(n9401), .Z(n9398) );
  XNOR2_X1 U9196 ( .A(n9402), .B(n9403), .ZN(n9191) );
  XNOR2_X1 U9197 ( .A(n9404), .B(n9405), .ZN(n9402) );
  NOR2_X1 U9198 ( .A1(n8759), .A2(n8738), .ZN(n9405) );
  XNOR2_X1 U9199 ( .A(n9406), .B(n9407), .ZN(n9196) );
  XNOR2_X1 U9200 ( .A(n9408), .B(n9409), .ZN(n9407) );
  XNOR2_X1 U9201 ( .A(n9410), .B(n9411), .ZN(n9200) );
  XNOR2_X1 U9202 ( .A(n9412), .B(n9413), .ZN(n9410) );
  NOR2_X1 U9203 ( .A1(n8761), .A2(n8738), .ZN(n9413) );
  XOR2_X1 U9204 ( .A(n9414), .B(n9415), .Z(n9203) );
  XOR2_X1 U9205 ( .A(n9416), .B(n9417), .Z(n9414) );
  XNOR2_X1 U9206 ( .A(n9418), .B(n9419), .ZN(n9207) );
  XOR2_X1 U9207 ( .A(n9420), .B(n9421), .Z(n9419) );
  NAND2_X1 U9208 ( .A1(b_29_), .A2(a_8_), .ZN(n9421) );
  XOR2_X1 U9209 ( .A(n9422), .B(n9423), .Z(n9212) );
  XNOR2_X1 U9210 ( .A(n9424), .B(n9425), .ZN(n9423) );
  XNOR2_X1 U9211 ( .A(n9426), .B(n9427), .ZN(n9215) );
  XNOR2_X1 U9212 ( .A(n9428), .B(n9429), .ZN(n9426) );
  NOR2_X1 U9213 ( .A1(n8491), .A2(n8738), .ZN(n9429) );
  XNOR2_X1 U9214 ( .A(n9430), .B(n9431), .ZN(n9220) );
  XOR2_X1 U9215 ( .A(n9432), .B(n9433), .Z(n9430) );
  XNOR2_X1 U9216 ( .A(n9434), .B(n9435), .ZN(n9223) );
  XNOR2_X1 U9217 ( .A(n9436), .B(n9437), .ZN(n9434) );
  NOR2_X1 U9218 ( .A1(n8766), .A2(n8738), .ZN(n9437) );
  XOR2_X1 U9219 ( .A(n9438), .B(n9439), .Z(n9228) );
  XOR2_X1 U9220 ( .A(n9440), .B(n9441), .Z(n9439) );
  NAND2_X1 U9221 ( .A1(b_29_), .A2(a_3_), .ZN(n9441) );
  XNOR2_X1 U9222 ( .A(n9442), .B(n9443), .ZN(n9232) );
  XNOR2_X1 U9223 ( .A(n9444), .B(n9445), .ZN(n9442) );
  XOR2_X1 U9224 ( .A(n9446), .B(n9447), .Z(n9015) );
  XOR2_X1 U9225 ( .A(n9448), .B(n9449), .Z(n9446) );
  NOR2_X1 U9226 ( .A1(n8617), .A2(n8738), .ZN(n9449) );
  XNOR2_X1 U9227 ( .A(n9450), .B(n9451), .ZN(n8781) );
  NAND2_X1 U9228 ( .A1(n9452), .A2(n9453), .ZN(n9450) );
  NAND2_X1 U9229 ( .A1(n9454), .A2(n9455), .ZN(n8797) );
  NAND2_X1 U9230 ( .A1(n9004), .A2(n9006), .ZN(n9455) );
  NAND2_X1 U9231 ( .A1(n9452), .A2(n9456), .ZN(n9006) );
  NAND2_X1 U9232 ( .A1(n9451), .A2(n9453), .ZN(n9456) );
  NAND2_X1 U9233 ( .A1(n9457), .A2(n9458), .ZN(n9453) );
  NAND2_X1 U9234 ( .A1(b_29_), .A2(a_0_), .ZN(n9458) );
  INV_X1 U9235 ( .A(n9459), .ZN(n9457) );
  XOR2_X1 U9236 ( .A(n9460), .B(n9461), .Z(n9451) );
  XOR2_X1 U9237 ( .A(n9462), .B(n9463), .Z(n9460) );
  NAND2_X1 U9238 ( .A1(a_0_), .A2(n9459), .ZN(n9452) );
  NAND2_X1 U9239 ( .A1(n9464), .A2(n9465), .ZN(n9459) );
  NAND3_X1 U9240 ( .A1(a_1_), .A2(n9466), .A3(b_29_), .ZN(n9465) );
  OR2_X1 U9241 ( .A1(n9448), .A2(n9447), .ZN(n9466) );
  NAND2_X1 U9242 ( .A1(n9447), .A2(n9448), .ZN(n9464) );
  NAND2_X1 U9243 ( .A1(n9467), .A2(n9468), .ZN(n9448) );
  NAND2_X1 U9244 ( .A1(n9444), .A2(n9469), .ZN(n9468) );
  NAND2_X1 U9245 ( .A1(n9443), .A2(n9445), .ZN(n9469) );
  NAND2_X1 U9246 ( .A1(n9470), .A2(n9471), .ZN(n9444) );
  NAND3_X1 U9247 ( .A1(a_3_), .A2(n9472), .A3(b_29_), .ZN(n9471) );
  OR2_X1 U9248 ( .A1(n9440), .A2(n9438), .ZN(n9472) );
  NAND2_X1 U9249 ( .A1(n9438), .A2(n9440), .ZN(n9470) );
  NAND2_X1 U9250 ( .A1(n9473), .A2(n9474), .ZN(n9440) );
  NAND3_X1 U9251 ( .A1(a_4_), .A2(n9475), .A3(b_29_), .ZN(n9474) );
  NAND2_X1 U9252 ( .A1(n9436), .A2(n9435), .ZN(n9475) );
  OR2_X1 U9253 ( .A1(n9435), .A2(n9436), .ZN(n9473) );
  AND2_X1 U9254 ( .A1(n9476), .A2(n9477), .ZN(n9436) );
  NAND2_X1 U9255 ( .A1(n9433), .A2(n9478), .ZN(n9477) );
  OR2_X1 U9256 ( .A1(n9432), .A2(n9431), .ZN(n9478) );
  NOR2_X1 U9257 ( .A1(n8738), .A2(n8517), .ZN(n9433) );
  NAND2_X1 U9258 ( .A1(n9431), .A2(n9432), .ZN(n9476) );
  NAND2_X1 U9259 ( .A1(n9479), .A2(n9480), .ZN(n9432) );
  NAND3_X1 U9260 ( .A1(a_6_), .A2(n9481), .A3(b_29_), .ZN(n9480) );
  NAND2_X1 U9261 ( .A1(n9428), .A2(n9427), .ZN(n9481) );
  OR2_X1 U9262 ( .A1(n9427), .A2(n9428), .ZN(n9479) );
  AND2_X1 U9263 ( .A1(n9482), .A2(n9483), .ZN(n9428) );
  NAND2_X1 U9264 ( .A1(n9425), .A2(n9484), .ZN(n9483) );
  OR2_X1 U9265 ( .A1(n9424), .A2(n9422), .ZN(n9484) );
  NOR2_X1 U9266 ( .A1(n8738), .A2(n8764), .ZN(n9425) );
  NAND2_X1 U9267 ( .A1(n9422), .A2(n9424), .ZN(n9482) );
  NAND2_X1 U9268 ( .A1(n9485), .A2(n9486), .ZN(n9424) );
  NAND3_X1 U9269 ( .A1(a_8_), .A2(n9487), .A3(b_29_), .ZN(n9486) );
  OR2_X1 U9270 ( .A1(n9420), .A2(n9418), .ZN(n9487) );
  NAND2_X1 U9271 ( .A1(n9418), .A2(n9420), .ZN(n9485) );
  NAND2_X1 U9272 ( .A1(n9488), .A2(n9489), .ZN(n9420) );
  NAND2_X1 U9273 ( .A1(n9417), .A2(n9490), .ZN(n9489) );
  OR2_X1 U9274 ( .A1(n9416), .A2(n9415), .ZN(n9490) );
  NOR2_X1 U9275 ( .A1(n8738), .A2(n8426), .ZN(n9417) );
  NAND2_X1 U9276 ( .A1(n9415), .A2(n9416), .ZN(n9488) );
  NAND2_X1 U9277 ( .A1(n9491), .A2(n9492), .ZN(n9416) );
  NAND3_X1 U9278 ( .A1(a_10_), .A2(n9493), .A3(b_29_), .ZN(n9492) );
  NAND2_X1 U9279 ( .A1(n9412), .A2(n9411), .ZN(n9493) );
  OR2_X1 U9280 ( .A1(n9411), .A2(n9412), .ZN(n9491) );
  AND2_X1 U9281 ( .A1(n9494), .A2(n9495), .ZN(n9412) );
  NAND2_X1 U9282 ( .A1(n9409), .A2(n9496), .ZN(n9495) );
  OR2_X1 U9283 ( .A1(n9408), .A2(n9406), .ZN(n9496) );
  NOR2_X1 U9284 ( .A1(n8738), .A2(n8376), .ZN(n9409) );
  NAND2_X1 U9285 ( .A1(n9406), .A2(n9408), .ZN(n9494) );
  NAND2_X1 U9286 ( .A1(n9497), .A2(n9498), .ZN(n9408) );
  NAND3_X1 U9287 ( .A1(a_12_), .A2(n9499), .A3(b_29_), .ZN(n9498) );
  NAND2_X1 U9288 ( .A1(n9404), .A2(n9403), .ZN(n9499) );
  OR2_X1 U9289 ( .A1(n9403), .A2(n9404), .ZN(n9497) );
  AND2_X1 U9290 ( .A1(n9500), .A2(n9501), .ZN(n9404) );
  NAND2_X1 U9291 ( .A1(n9401), .A2(n9502), .ZN(n9501) );
  OR2_X1 U9292 ( .A1(n9400), .A2(n9399), .ZN(n9502) );
  NOR2_X1 U9293 ( .A1(n8738), .A2(n8310), .ZN(n9401) );
  NAND2_X1 U9294 ( .A1(n9399), .A2(n9400), .ZN(n9500) );
  NAND2_X1 U9295 ( .A1(n9503), .A2(n9504), .ZN(n9400) );
  NAND3_X1 U9296 ( .A1(a_14_), .A2(n9505), .A3(b_29_), .ZN(n9504) );
  NAND2_X1 U9297 ( .A1(n9397), .A2(n9395), .ZN(n9505) );
  OR2_X1 U9298 ( .A1(n9395), .A2(n9397), .ZN(n9503) );
  AND2_X1 U9299 ( .A1(n9506), .A2(n9507), .ZN(n9397) );
  NAND2_X1 U9300 ( .A1(n9393), .A2(n9508), .ZN(n9507) );
  OR2_X1 U9301 ( .A1(n9392), .A2(n9390), .ZN(n9508) );
  NOR2_X1 U9302 ( .A1(n8738), .A2(n8276), .ZN(n9393) );
  NAND2_X1 U9303 ( .A1(n9390), .A2(n9392), .ZN(n9506) );
  NAND2_X1 U9304 ( .A1(n9509), .A2(n9510), .ZN(n9392) );
  NAND3_X1 U9305 ( .A1(a_16_), .A2(n9511), .A3(b_29_), .ZN(n9510) );
  OR2_X1 U9306 ( .A1(n9388), .A2(n9386), .ZN(n9511) );
  NAND2_X1 U9307 ( .A1(n9386), .A2(n9388), .ZN(n9509) );
  NAND2_X1 U9308 ( .A1(n9512), .A2(n9513), .ZN(n9388) );
  NAND2_X1 U9309 ( .A1(n9385), .A2(n9514), .ZN(n9513) );
  OR2_X1 U9310 ( .A1(n9384), .A2(n9383), .ZN(n9514) );
  NOR2_X1 U9311 ( .A1(n8738), .A2(n8210), .ZN(n9385) );
  NAND2_X1 U9312 ( .A1(n9383), .A2(n9384), .ZN(n9512) );
  NAND2_X1 U9313 ( .A1(n9515), .A2(n9516), .ZN(n9384) );
  NAND3_X1 U9314 ( .A1(a_18_), .A2(n9517), .A3(b_29_), .ZN(n9516) );
  NAND2_X1 U9315 ( .A1(n9380), .A2(n9379), .ZN(n9517) );
  OR2_X1 U9316 ( .A1(n9379), .A2(n9380), .ZN(n9515) );
  AND2_X1 U9317 ( .A1(n9518), .A2(n9519), .ZN(n9380) );
  NAND2_X1 U9318 ( .A1(n9377), .A2(n9520), .ZN(n9519) );
  OR2_X1 U9319 ( .A1(n9376), .A2(n9374), .ZN(n9520) );
  NOR2_X1 U9320 ( .A1(n8738), .A2(n8170), .ZN(n9377) );
  NAND2_X1 U9321 ( .A1(n9374), .A2(n9376), .ZN(n9518) );
  NAND2_X1 U9322 ( .A1(n9521), .A2(n9522), .ZN(n9376) );
  NAND3_X1 U9323 ( .A1(a_20_), .A2(n9523), .A3(b_29_), .ZN(n9522) );
  NAND2_X1 U9324 ( .A1(n9372), .A2(n9371), .ZN(n9523) );
  OR2_X1 U9325 ( .A1(n9371), .A2(n9372), .ZN(n9521) );
  AND2_X1 U9326 ( .A1(n9524), .A2(n9525), .ZN(n9372) );
  NAND2_X1 U9327 ( .A1(n9369), .A2(n9526), .ZN(n9525) );
  OR2_X1 U9328 ( .A1(n9368), .A2(n9367), .ZN(n9526) );
  NOR2_X1 U9329 ( .A1(n8738), .A2(n8750), .ZN(n9369) );
  NAND2_X1 U9330 ( .A1(n9367), .A2(n9368), .ZN(n9524) );
  NAND2_X1 U9331 ( .A1(n9527), .A2(n9528), .ZN(n9368) );
  NAND3_X1 U9332 ( .A1(a_22_), .A2(n9529), .A3(b_29_), .ZN(n9528) );
  OR2_X1 U9333 ( .A1(n9364), .A2(n9362), .ZN(n9529) );
  NAND2_X1 U9334 ( .A1(n9362), .A2(n9364), .ZN(n9527) );
  NAND2_X1 U9335 ( .A1(n9530), .A2(n9531), .ZN(n9364) );
  NAND2_X1 U9336 ( .A1(n9361), .A2(n9532), .ZN(n9531) );
  OR2_X1 U9337 ( .A1(n9360), .A2(n9358), .ZN(n9532) );
  NOR2_X1 U9338 ( .A1(n8738), .A2(n8747), .ZN(n9361) );
  NAND2_X1 U9339 ( .A1(n9358), .A2(n9360), .ZN(n9530) );
  NAND2_X1 U9340 ( .A1(n9533), .A2(n9534), .ZN(n9360) );
  NAND3_X1 U9341 ( .A1(a_24_), .A2(n9535), .A3(b_29_), .ZN(n9534) );
  OR2_X1 U9342 ( .A1(n9356), .A2(n9354), .ZN(n9535) );
  NAND2_X1 U9343 ( .A1(n9354), .A2(n9356), .ZN(n9533) );
  NAND2_X1 U9344 ( .A1(n9536), .A2(n9537), .ZN(n9356) );
  NAND2_X1 U9345 ( .A1(n9353), .A2(n9538), .ZN(n9537) );
  NAND2_X1 U9346 ( .A1(n9352), .A2(n9351), .ZN(n9538) );
  NOR2_X1 U9347 ( .A1(n8738), .A2(n8744), .ZN(n9353) );
  OR2_X1 U9348 ( .A1(n9351), .A2(n9352), .ZN(n9536) );
  AND2_X1 U9349 ( .A1(n9348), .A2(n9539), .ZN(n9352) );
  NAND2_X1 U9350 ( .A1(n9347), .A2(n9349), .ZN(n9539) );
  NAND2_X1 U9351 ( .A1(n9540), .A2(n9541), .ZN(n9349) );
  NAND2_X1 U9352 ( .A1(b_29_), .A2(a_26_), .ZN(n9541) );
  INV_X1 U9353 ( .A(n9542), .ZN(n9540) );
  XNOR2_X1 U9354 ( .A(n9543), .B(n9544), .ZN(n9347) );
  NAND2_X1 U9355 ( .A1(n9545), .A2(n9546), .ZN(n9543) );
  NAND2_X1 U9356 ( .A1(a_26_), .A2(n9542), .ZN(n9348) );
  NAND2_X1 U9357 ( .A1(n9320), .A2(n9547), .ZN(n9542) );
  NAND2_X1 U9358 ( .A1(n9319), .A2(n9321), .ZN(n9547) );
  NAND2_X1 U9359 ( .A1(n9548), .A2(n9549), .ZN(n9321) );
  NAND2_X1 U9360 ( .A1(b_29_), .A2(a_27_), .ZN(n9549) );
  INV_X1 U9361 ( .A(n9550), .ZN(n9548) );
  XOR2_X1 U9362 ( .A(n9551), .B(n9552), .Z(n9319) );
  XOR2_X1 U9363 ( .A(n8731), .B(n9553), .Z(n9551) );
  NAND2_X1 U9364 ( .A1(a_27_), .A2(n9550), .ZN(n9320) );
  NAND2_X1 U9365 ( .A1(n9554), .A2(n9555), .ZN(n9550) );
  NAND3_X1 U9366 ( .A1(a_28_), .A2(n9556), .A3(b_29_), .ZN(n9555) );
  NAND2_X1 U9367 ( .A1(n9329), .A2(n9327), .ZN(n9556) );
  OR2_X1 U9368 ( .A1(n9327), .A2(n9329), .ZN(n9554) );
  AND2_X1 U9369 ( .A1(n9557), .A2(n9558), .ZN(n9329) );
  NAND2_X1 U9370 ( .A1(n9343), .A2(n9559), .ZN(n9558) );
  OR2_X1 U9371 ( .A1(n9344), .A2(n9345), .ZN(n9559) );
  INV_X1 U9372 ( .A(n7909), .ZN(n9343) );
  NAND2_X1 U9373 ( .A1(b_29_), .A2(a_29_), .ZN(n7909) );
  NAND2_X1 U9374 ( .A1(n9345), .A2(n9344), .ZN(n9557) );
  NAND2_X1 U9375 ( .A1(n9560), .A2(n9561), .ZN(n9344) );
  NAND2_X1 U9376 ( .A1(b_27_), .A2(n9562), .ZN(n9561) );
  NAND2_X1 U9377 ( .A1(n7864), .A2(n9563), .ZN(n9562) );
  NAND2_X1 U9378 ( .A1(a_31_), .A2(n7935), .ZN(n9563) );
  NAND2_X1 U9379 ( .A1(b_28_), .A2(n9564), .ZN(n9560) );
  NAND2_X1 U9380 ( .A1(n9137), .A2(n9565), .ZN(n9564) );
  NAND2_X1 U9381 ( .A1(a_30_), .A2(n8740), .ZN(n9565) );
  AND3_X1 U9382 ( .A1(b_28_), .A2(b_29_), .A3(n7818), .ZN(n9345) );
  XNOR2_X1 U9383 ( .A(n9566), .B(n9567), .ZN(n9327) );
  XOR2_X1 U9384 ( .A(n9568), .B(n9569), .Z(n9566) );
  XOR2_X1 U9385 ( .A(n9570), .B(n9571), .Z(n9351) );
  NAND2_X1 U9386 ( .A1(n9572), .A2(n9573), .ZN(n9570) );
  XOR2_X1 U9387 ( .A(n9574), .B(n9575), .Z(n9354) );
  XOR2_X1 U9388 ( .A(n9576), .B(n9577), .Z(n9574) );
  XOR2_X1 U9389 ( .A(n9578), .B(n9579), .Z(n9358) );
  XOR2_X1 U9390 ( .A(n9580), .B(n9581), .Z(n9578) );
  NOR2_X1 U9391 ( .A1(n8745), .A2(n7935), .ZN(n9581) );
  XNOR2_X1 U9392 ( .A(n9582), .B(n9583), .ZN(n9362) );
  XNOR2_X1 U9393 ( .A(n9584), .B(n9585), .ZN(n9583) );
  XNOR2_X1 U9394 ( .A(n9586), .B(n9587), .ZN(n9367) );
  XNOR2_X1 U9395 ( .A(n9588), .B(n9589), .ZN(n9586) );
  NOR2_X1 U9396 ( .A1(n8748), .A2(n7935), .ZN(n9589) );
  XNOR2_X1 U9397 ( .A(n9590), .B(n9591), .ZN(n9371) );
  XOR2_X1 U9398 ( .A(n9592), .B(n9593), .Z(n9590) );
  XNOR2_X1 U9399 ( .A(n9594), .B(n9595), .ZN(n9374) );
  XNOR2_X1 U9400 ( .A(n9596), .B(n9597), .ZN(n9594) );
  NOR2_X1 U9401 ( .A1(n8751), .A2(n7935), .ZN(n9597) );
  XOR2_X1 U9402 ( .A(n9598), .B(n9599), .Z(n9379) );
  XNOR2_X1 U9403 ( .A(n9600), .B(n9601), .ZN(n9599) );
  XNOR2_X1 U9404 ( .A(n9602), .B(n9603), .ZN(n9383) );
  XNOR2_X1 U9405 ( .A(n9604), .B(n9605), .ZN(n9602) );
  NOR2_X1 U9406 ( .A1(n8753), .A2(n7935), .ZN(n9605) );
  XOR2_X1 U9407 ( .A(n9606), .B(n9607), .Z(n9386) );
  XOR2_X1 U9408 ( .A(n9608), .B(n9609), .Z(n9606) );
  XNOR2_X1 U9409 ( .A(n9610), .B(n9611), .ZN(n9390) );
  XOR2_X1 U9410 ( .A(n9612), .B(n9613), .Z(n9611) );
  NAND2_X1 U9411 ( .A1(b_28_), .A2(a_16_), .ZN(n9613) );
  XOR2_X1 U9412 ( .A(n9614), .B(n9615), .Z(n9395) );
  XNOR2_X1 U9413 ( .A(n9616), .B(n9617), .ZN(n9615) );
  XNOR2_X1 U9414 ( .A(n9618), .B(n9619), .ZN(n9399) );
  XNOR2_X1 U9415 ( .A(n9620), .B(n9621), .ZN(n9618) );
  NOR2_X1 U9416 ( .A1(n8757), .A2(n7935), .ZN(n9621) );
  XNOR2_X1 U9417 ( .A(n9622), .B(n9623), .ZN(n9403) );
  XOR2_X1 U9418 ( .A(n9624), .B(n9625), .Z(n9622) );
  XOR2_X1 U9419 ( .A(n9626), .B(n9627), .Z(n9406) );
  XOR2_X1 U9420 ( .A(n9628), .B(n9629), .Z(n9626) );
  NOR2_X1 U9421 ( .A1(n8759), .A2(n7935), .ZN(n9629) );
  XOR2_X1 U9422 ( .A(n9630), .B(n9631), .Z(n9411) );
  XNOR2_X1 U9423 ( .A(n9632), .B(n9633), .ZN(n9631) );
  XNOR2_X1 U9424 ( .A(n9634), .B(n9635), .ZN(n9415) );
  XNOR2_X1 U9425 ( .A(n9636), .B(n9637), .ZN(n9634) );
  NOR2_X1 U9426 ( .A1(n8761), .A2(n7935), .ZN(n9637) );
  XNOR2_X1 U9427 ( .A(n9638), .B(n9639), .ZN(n9418) );
  XNOR2_X1 U9428 ( .A(n9640), .B(n9641), .ZN(n9638) );
  XNOR2_X1 U9429 ( .A(n9642), .B(n9643), .ZN(n9422) );
  XOR2_X1 U9430 ( .A(n9644), .B(n9645), .Z(n9643) );
  NAND2_X1 U9431 ( .A1(b_28_), .A2(a_8_), .ZN(n9645) );
  XOR2_X1 U9432 ( .A(n9646), .B(n9647), .Z(n9427) );
  XNOR2_X1 U9433 ( .A(n9648), .B(n9649), .ZN(n9647) );
  XNOR2_X1 U9434 ( .A(n9650), .B(n9651), .ZN(n9431) );
  XNOR2_X1 U9435 ( .A(n9652), .B(n9653), .ZN(n9650) );
  NOR2_X1 U9436 ( .A1(n8491), .A2(n7935), .ZN(n9653) );
  XNOR2_X1 U9437 ( .A(n9654), .B(n9655), .ZN(n9435) );
  XOR2_X1 U9438 ( .A(n9656), .B(n9657), .Z(n9654) );
  XNOR2_X1 U9439 ( .A(n9658), .B(n9659), .ZN(n9438) );
  XNOR2_X1 U9440 ( .A(n9660), .B(n9661), .ZN(n9658) );
  NOR2_X1 U9441 ( .A1(n8766), .A2(n7935), .ZN(n9661) );
  OR2_X1 U9442 ( .A1(n9445), .A2(n9443), .ZN(n9467) );
  XOR2_X1 U9443 ( .A(n9662), .B(n9663), .Z(n9443) );
  XOR2_X1 U9444 ( .A(n9664), .B(n9665), .Z(n9663) );
  NAND2_X1 U9445 ( .A1(b_28_), .A2(a_3_), .ZN(n9665) );
  NAND2_X1 U9446 ( .A1(b_29_), .A2(a_2_), .ZN(n9445) );
  XNOR2_X1 U9447 ( .A(n9666), .B(n9667), .ZN(n9447) );
  XNOR2_X1 U9448 ( .A(n9668), .B(n9669), .ZN(n9666) );
  INV_X1 U9449 ( .A(n9013), .ZN(n9004) );
  XOR2_X1 U9450 ( .A(n9670), .B(n9671), .Z(n9013) );
  XNOR2_X1 U9451 ( .A(n9672), .B(n9673), .ZN(n9670) );
  NOR2_X1 U9452 ( .A1(n9674), .A2(n7935), .ZN(n9673) );
  XNOR2_X1 U9453 ( .A(n9008), .B(n9007), .ZN(n9454) );
  NAND2_X1 U9454 ( .A1(n9002), .A2(n9001), .ZN(n8804) );
  NAND2_X1 U9455 ( .A1(n9675), .A2(n9676), .ZN(n9001) );
  NAND2_X1 U9456 ( .A1(n9677), .A2(n9678), .ZN(n9675) );
  OR2_X1 U9457 ( .A1(n9008), .A2(n9007), .ZN(n9002) );
  AND2_X1 U9458 ( .A1(n9679), .A2(n9680), .ZN(n9007) );
  NAND3_X1 U9459 ( .A1(a_0_), .A2(n9681), .A3(b_28_), .ZN(n9680) );
  NAND2_X1 U9460 ( .A1(n9672), .A2(n9671), .ZN(n9681) );
  OR2_X1 U9461 ( .A1(n9671), .A2(n9672), .ZN(n9679) );
  AND2_X1 U9462 ( .A1(n9682), .A2(n9683), .ZN(n9672) );
  NAND2_X1 U9463 ( .A1(n9463), .A2(n9684), .ZN(n9683) );
  OR2_X1 U9464 ( .A1(n9462), .A2(n9461), .ZN(n9684) );
  NOR2_X1 U9465 ( .A1(n7935), .A2(n8617), .ZN(n9463) );
  NAND2_X1 U9466 ( .A1(n9461), .A2(n9462), .ZN(n9682) );
  NAND2_X1 U9467 ( .A1(n9685), .A2(n9686), .ZN(n9462) );
  NAND2_X1 U9468 ( .A1(n9668), .A2(n9687), .ZN(n9686) );
  NAND2_X1 U9469 ( .A1(n9667), .A2(n9669), .ZN(n9687) );
  NAND2_X1 U9470 ( .A1(n9688), .A2(n9689), .ZN(n9668) );
  NAND3_X1 U9471 ( .A1(a_3_), .A2(n9690), .A3(b_28_), .ZN(n9689) );
  OR2_X1 U9472 ( .A1(n9664), .A2(n9662), .ZN(n9690) );
  NAND2_X1 U9473 ( .A1(n9662), .A2(n9664), .ZN(n9688) );
  NAND2_X1 U9474 ( .A1(n9691), .A2(n9692), .ZN(n9664) );
  NAND3_X1 U9475 ( .A1(a_4_), .A2(n9693), .A3(b_28_), .ZN(n9692) );
  NAND2_X1 U9476 ( .A1(n9660), .A2(n9659), .ZN(n9693) );
  OR2_X1 U9477 ( .A1(n9659), .A2(n9660), .ZN(n9691) );
  AND2_X1 U9478 ( .A1(n9694), .A2(n9695), .ZN(n9660) );
  NAND2_X1 U9479 ( .A1(n9657), .A2(n9696), .ZN(n9695) );
  OR2_X1 U9480 ( .A1(n9656), .A2(n9655), .ZN(n9696) );
  NOR2_X1 U9481 ( .A1(n7935), .A2(n8517), .ZN(n9657) );
  NAND2_X1 U9482 ( .A1(n9655), .A2(n9656), .ZN(n9694) );
  NAND2_X1 U9483 ( .A1(n9697), .A2(n9698), .ZN(n9656) );
  NAND3_X1 U9484 ( .A1(a_6_), .A2(n9699), .A3(b_28_), .ZN(n9698) );
  NAND2_X1 U9485 ( .A1(n9652), .A2(n9651), .ZN(n9699) );
  OR2_X1 U9486 ( .A1(n9651), .A2(n9652), .ZN(n9697) );
  AND2_X1 U9487 ( .A1(n9700), .A2(n9701), .ZN(n9652) );
  NAND2_X1 U9488 ( .A1(n9649), .A2(n9702), .ZN(n9701) );
  OR2_X1 U9489 ( .A1(n9648), .A2(n9646), .ZN(n9702) );
  NOR2_X1 U9490 ( .A1(n7935), .A2(n8764), .ZN(n9649) );
  NAND2_X1 U9491 ( .A1(n9646), .A2(n9648), .ZN(n9700) );
  NAND2_X1 U9492 ( .A1(n9703), .A2(n9704), .ZN(n9648) );
  NAND3_X1 U9493 ( .A1(a_8_), .A2(n9705), .A3(b_28_), .ZN(n9704) );
  OR2_X1 U9494 ( .A1(n9644), .A2(n9642), .ZN(n9705) );
  NAND2_X1 U9495 ( .A1(n9642), .A2(n9644), .ZN(n9703) );
  NAND2_X1 U9496 ( .A1(n9706), .A2(n9707), .ZN(n9644) );
  NAND2_X1 U9497 ( .A1(n9641), .A2(n9708), .ZN(n9707) );
  NAND2_X1 U9498 ( .A1(n9640), .A2(n9639), .ZN(n9708) );
  NOR2_X1 U9499 ( .A1(n7935), .A2(n8426), .ZN(n9641) );
  OR2_X1 U9500 ( .A1(n9639), .A2(n9640), .ZN(n9706) );
  AND2_X1 U9501 ( .A1(n9709), .A2(n9710), .ZN(n9640) );
  NAND3_X1 U9502 ( .A1(a_10_), .A2(n9711), .A3(b_28_), .ZN(n9710) );
  NAND2_X1 U9503 ( .A1(n9636), .A2(n9635), .ZN(n9711) );
  OR2_X1 U9504 ( .A1(n9635), .A2(n9636), .ZN(n9709) );
  AND2_X1 U9505 ( .A1(n9712), .A2(n9713), .ZN(n9636) );
  NAND2_X1 U9506 ( .A1(n9633), .A2(n9714), .ZN(n9713) );
  OR2_X1 U9507 ( .A1(n9632), .A2(n9630), .ZN(n9714) );
  NOR2_X1 U9508 ( .A1(n7935), .A2(n8376), .ZN(n9633) );
  NAND2_X1 U9509 ( .A1(n9630), .A2(n9632), .ZN(n9712) );
  NAND2_X1 U9510 ( .A1(n9715), .A2(n9716), .ZN(n9632) );
  NAND3_X1 U9511 ( .A1(a_12_), .A2(n9717), .A3(b_28_), .ZN(n9716) );
  OR2_X1 U9512 ( .A1(n9628), .A2(n9627), .ZN(n9717) );
  NAND2_X1 U9513 ( .A1(n9627), .A2(n9628), .ZN(n9715) );
  NAND2_X1 U9514 ( .A1(n9718), .A2(n9719), .ZN(n9628) );
  NAND2_X1 U9515 ( .A1(n9625), .A2(n9720), .ZN(n9719) );
  OR2_X1 U9516 ( .A1(n9624), .A2(n9623), .ZN(n9720) );
  NOR2_X1 U9517 ( .A1(n7935), .A2(n8310), .ZN(n9625) );
  NAND2_X1 U9518 ( .A1(n9623), .A2(n9624), .ZN(n9718) );
  NAND2_X1 U9519 ( .A1(n9721), .A2(n9722), .ZN(n9624) );
  NAND3_X1 U9520 ( .A1(a_14_), .A2(n9723), .A3(b_28_), .ZN(n9722) );
  NAND2_X1 U9521 ( .A1(n9620), .A2(n9619), .ZN(n9723) );
  OR2_X1 U9522 ( .A1(n9619), .A2(n9620), .ZN(n9721) );
  AND2_X1 U9523 ( .A1(n9724), .A2(n9725), .ZN(n9620) );
  NAND2_X1 U9524 ( .A1(n9617), .A2(n9726), .ZN(n9725) );
  OR2_X1 U9525 ( .A1(n9616), .A2(n9614), .ZN(n9726) );
  NOR2_X1 U9526 ( .A1(n7935), .A2(n8276), .ZN(n9617) );
  NAND2_X1 U9527 ( .A1(n9614), .A2(n9616), .ZN(n9724) );
  NAND2_X1 U9528 ( .A1(n9727), .A2(n9728), .ZN(n9616) );
  NAND3_X1 U9529 ( .A1(a_16_), .A2(n9729), .A3(b_28_), .ZN(n9728) );
  OR2_X1 U9530 ( .A1(n9612), .A2(n9610), .ZN(n9729) );
  NAND2_X1 U9531 ( .A1(n9610), .A2(n9612), .ZN(n9727) );
  NAND2_X1 U9532 ( .A1(n9730), .A2(n9731), .ZN(n9612) );
  NAND2_X1 U9533 ( .A1(n9609), .A2(n9732), .ZN(n9731) );
  OR2_X1 U9534 ( .A1(n9608), .A2(n9607), .ZN(n9732) );
  NOR2_X1 U9535 ( .A1(n7935), .A2(n8210), .ZN(n9609) );
  NAND2_X1 U9536 ( .A1(n9607), .A2(n9608), .ZN(n9730) );
  NAND2_X1 U9537 ( .A1(n9733), .A2(n9734), .ZN(n9608) );
  NAND3_X1 U9538 ( .A1(a_18_), .A2(n9735), .A3(b_28_), .ZN(n9734) );
  NAND2_X1 U9539 ( .A1(n9604), .A2(n9603), .ZN(n9735) );
  OR2_X1 U9540 ( .A1(n9603), .A2(n9604), .ZN(n9733) );
  AND2_X1 U9541 ( .A1(n9736), .A2(n9737), .ZN(n9604) );
  NAND2_X1 U9542 ( .A1(n9601), .A2(n9738), .ZN(n9737) );
  OR2_X1 U9543 ( .A1(n9600), .A2(n9598), .ZN(n9738) );
  NOR2_X1 U9544 ( .A1(n7935), .A2(n8170), .ZN(n9601) );
  NAND2_X1 U9545 ( .A1(n9598), .A2(n9600), .ZN(n9736) );
  NAND2_X1 U9546 ( .A1(n9739), .A2(n9740), .ZN(n9600) );
  NAND3_X1 U9547 ( .A1(a_20_), .A2(n9741), .A3(b_28_), .ZN(n9740) );
  NAND2_X1 U9548 ( .A1(n9596), .A2(n9595), .ZN(n9741) );
  OR2_X1 U9549 ( .A1(n9595), .A2(n9596), .ZN(n9739) );
  AND2_X1 U9550 ( .A1(n9742), .A2(n9743), .ZN(n9596) );
  NAND2_X1 U9551 ( .A1(n9593), .A2(n9744), .ZN(n9743) );
  OR2_X1 U9552 ( .A1(n9592), .A2(n9591), .ZN(n9744) );
  NOR2_X1 U9553 ( .A1(n7935), .A2(n8750), .ZN(n9593) );
  NAND2_X1 U9554 ( .A1(n9591), .A2(n9592), .ZN(n9742) );
  NAND2_X1 U9555 ( .A1(n9745), .A2(n9746), .ZN(n9592) );
  NAND3_X1 U9556 ( .A1(a_22_), .A2(n9747), .A3(b_28_), .ZN(n9746) );
  NAND2_X1 U9557 ( .A1(n9588), .A2(n9587), .ZN(n9747) );
  OR2_X1 U9558 ( .A1(n9587), .A2(n9588), .ZN(n9745) );
  AND2_X1 U9559 ( .A1(n9748), .A2(n9749), .ZN(n9588) );
  NAND2_X1 U9560 ( .A1(n9585), .A2(n9750), .ZN(n9749) );
  OR2_X1 U9561 ( .A1(n9584), .A2(n9582), .ZN(n9750) );
  NOR2_X1 U9562 ( .A1(n7935), .A2(n8747), .ZN(n9585) );
  NAND2_X1 U9563 ( .A1(n9582), .A2(n9584), .ZN(n9748) );
  NAND2_X1 U9564 ( .A1(n9751), .A2(n9752), .ZN(n9584) );
  NAND3_X1 U9565 ( .A1(a_24_), .A2(n9753), .A3(b_28_), .ZN(n9752) );
  OR2_X1 U9566 ( .A1(n9580), .A2(n9579), .ZN(n9753) );
  NAND2_X1 U9567 ( .A1(n9579), .A2(n9580), .ZN(n9751) );
  NAND2_X1 U9568 ( .A1(n9754), .A2(n9755), .ZN(n9580) );
  NAND2_X1 U9569 ( .A1(n9577), .A2(n9756), .ZN(n9755) );
  OR2_X1 U9570 ( .A1(n9576), .A2(n9575), .ZN(n9756) );
  NOR2_X1 U9571 ( .A1(n7935), .A2(n8744), .ZN(n9577) );
  NAND2_X1 U9572 ( .A1(n9575), .A2(n9576), .ZN(n9754) );
  NAND2_X1 U9573 ( .A1(n9572), .A2(n9757), .ZN(n9576) );
  NAND2_X1 U9574 ( .A1(n9571), .A2(n9573), .ZN(n9757) );
  NAND2_X1 U9575 ( .A1(n9758), .A2(n9759), .ZN(n9573) );
  NAND2_X1 U9576 ( .A1(b_28_), .A2(a_26_), .ZN(n9759) );
  INV_X1 U9577 ( .A(n9760), .ZN(n9758) );
  XOR2_X1 U9578 ( .A(n9761), .B(n9762), .Z(n9571) );
  XOR2_X1 U9579 ( .A(n9763), .B(n9764), .Z(n9761) );
  NAND2_X1 U9580 ( .A1(a_26_), .A2(n9760), .ZN(n9572) );
  NAND2_X1 U9581 ( .A1(n9545), .A2(n9765), .ZN(n9760) );
  NAND2_X1 U9582 ( .A1(n9544), .A2(n9546), .ZN(n9765) );
  NAND2_X1 U9583 ( .A1(n9766), .A2(n9767), .ZN(n9546) );
  NAND2_X1 U9584 ( .A1(b_28_), .A2(a_27_), .ZN(n9767) );
  INV_X1 U9585 ( .A(n9768), .ZN(n9766) );
  XNOR2_X1 U9586 ( .A(n9769), .B(n9770), .ZN(n9544) );
  XOR2_X1 U9587 ( .A(n9771), .B(n9772), .Z(n9769) );
  NAND2_X1 U9588 ( .A1(b_27_), .A2(a_28_), .ZN(n9771) );
  NAND2_X1 U9589 ( .A1(a_27_), .A2(n9768), .ZN(n9545) );
  NAND2_X1 U9590 ( .A1(n9773), .A2(n9774), .ZN(n9768) );
  NAND2_X1 U9591 ( .A1(n9552), .A2(n9775), .ZN(n9774) );
  NAND2_X1 U9592 ( .A1(n9553), .A2(n8731), .ZN(n9775) );
  INV_X1 U9593 ( .A(n9776), .ZN(n9553) );
  XOR2_X1 U9594 ( .A(n9777), .B(n9778), .Z(n9552) );
  XOR2_X1 U9595 ( .A(n9779), .B(n9780), .Z(n9777) );
  NAND2_X1 U9596 ( .A1(n9781), .A2(n9776), .ZN(n9773) );
  NAND2_X1 U9597 ( .A1(n9782), .A2(n9783), .ZN(n9776) );
  NAND2_X1 U9598 ( .A1(n9567), .A2(n9784), .ZN(n9783) );
  OR2_X1 U9599 ( .A1(n9568), .A2(n9569), .ZN(n9784) );
  NOR2_X1 U9600 ( .A1(n7935), .A2(n7890), .ZN(n9567) );
  NAND2_X1 U9601 ( .A1(n9569), .A2(n9568), .ZN(n9782) );
  NAND2_X1 U9602 ( .A1(n9785), .A2(n9786), .ZN(n9568) );
  NAND2_X1 U9603 ( .A1(b_26_), .A2(n9787), .ZN(n9786) );
  NAND2_X1 U9604 ( .A1(n7864), .A2(n9788), .ZN(n9787) );
  NAND2_X1 U9605 ( .A1(a_31_), .A2(n8740), .ZN(n9788) );
  NAND2_X1 U9606 ( .A1(b_27_), .A2(n9789), .ZN(n9785) );
  NAND2_X1 U9607 ( .A1(n9137), .A2(n9790), .ZN(n9789) );
  NAND2_X1 U9608 ( .A1(a_30_), .A2(n7992), .ZN(n9790) );
  AND3_X1 U9609 ( .A1(b_27_), .A2(b_28_), .A3(n7818), .ZN(n9569) );
  INV_X1 U9610 ( .A(n8731), .ZN(n9781) );
  NAND2_X1 U9611 ( .A1(b_28_), .A2(a_28_), .ZN(n8731) );
  XNOR2_X1 U9612 ( .A(n9791), .B(n9792), .ZN(n9575) );
  NAND2_X1 U9613 ( .A1(n9793), .A2(n9794), .ZN(n9791) );
  XNOR2_X1 U9614 ( .A(n9795), .B(n9796), .ZN(n9579) );
  XNOR2_X1 U9615 ( .A(n9797), .B(n9798), .ZN(n9795) );
  XNOR2_X1 U9616 ( .A(n9799), .B(n9800), .ZN(n9582) );
  XNOR2_X1 U9617 ( .A(n9801), .B(n9802), .ZN(n9799) );
  NOR2_X1 U9618 ( .A1(n8745), .A2(n8740), .ZN(n9802) );
  XOR2_X1 U9619 ( .A(n9803), .B(n9804), .Z(n9587) );
  XNOR2_X1 U9620 ( .A(n9805), .B(n9806), .ZN(n9804) );
  XNOR2_X1 U9621 ( .A(n9807), .B(n9808), .ZN(n9591) );
  XOR2_X1 U9622 ( .A(n9809), .B(n9810), .Z(n9808) );
  NAND2_X1 U9623 ( .A1(b_27_), .A2(a_22_), .ZN(n9810) );
  XNOR2_X1 U9624 ( .A(n9811), .B(n9812), .ZN(n9595) );
  XOR2_X1 U9625 ( .A(n9813), .B(n9814), .Z(n9811) );
  XNOR2_X1 U9626 ( .A(n9815), .B(n9816), .ZN(n9598) );
  XNOR2_X1 U9627 ( .A(n9817), .B(n9818), .ZN(n9815) );
  NOR2_X1 U9628 ( .A1(n8751), .A2(n8740), .ZN(n9818) );
  XOR2_X1 U9629 ( .A(n9819), .B(n9820), .Z(n9603) );
  XNOR2_X1 U9630 ( .A(n9821), .B(n9822), .ZN(n9820) );
  XNOR2_X1 U9631 ( .A(n9823), .B(n9824), .ZN(n9607) );
  XNOR2_X1 U9632 ( .A(n9825), .B(n9826), .ZN(n9823) );
  NOR2_X1 U9633 ( .A1(n8753), .A2(n8740), .ZN(n9826) );
  XOR2_X1 U9634 ( .A(n9827), .B(n9828), .Z(n9610) );
  XOR2_X1 U9635 ( .A(n9829), .B(n9830), .Z(n9827) );
  XNOR2_X1 U9636 ( .A(n9831), .B(n9832), .ZN(n9614) );
  XNOR2_X1 U9637 ( .A(n9833), .B(n9834), .ZN(n9831) );
  NOR2_X1 U9638 ( .A1(n8755), .A2(n8740), .ZN(n9834) );
  XOR2_X1 U9639 ( .A(n9835), .B(n9836), .Z(n9619) );
  XNOR2_X1 U9640 ( .A(n9837), .B(n9838), .ZN(n9836) );
  XNOR2_X1 U9641 ( .A(n9839), .B(n9840), .ZN(n9623) );
  XOR2_X1 U9642 ( .A(n9841), .B(n9842), .Z(n9839) );
  NAND2_X1 U9643 ( .A1(b_27_), .A2(a_14_), .ZN(n9841) );
  XNOR2_X1 U9644 ( .A(n9843), .B(n9844), .ZN(n9627) );
  XNOR2_X1 U9645 ( .A(n9845), .B(n9846), .ZN(n9843) );
  XNOR2_X1 U9646 ( .A(n9847), .B(n9848), .ZN(n9630) );
  XNOR2_X1 U9647 ( .A(n9849), .B(n9850), .ZN(n9847) );
  NOR2_X1 U9648 ( .A1(n8759), .A2(n8740), .ZN(n9850) );
  XOR2_X1 U9649 ( .A(n9851), .B(n9852), .Z(n9635) );
  XNOR2_X1 U9650 ( .A(n9853), .B(n9854), .ZN(n9852) );
  XNOR2_X1 U9651 ( .A(n9855), .B(n9856), .ZN(n9639) );
  XOR2_X1 U9652 ( .A(n9857), .B(n9858), .Z(n9855) );
  NOR2_X1 U9653 ( .A1(n8761), .A2(n8740), .ZN(n9858) );
  XOR2_X1 U9654 ( .A(n9859), .B(n9860), .Z(n9642) );
  XOR2_X1 U9655 ( .A(n9861), .B(n9862), .Z(n9859) );
  XNOR2_X1 U9656 ( .A(n9863), .B(n9864), .ZN(n9646) );
  XNOR2_X1 U9657 ( .A(n9865), .B(n9866), .ZN(n9863) );
  NOR2_X1 U9658 ( .A1(n8763), .A2(n8740), .ZN(n9866) );
  XOR2_X1 U9659 ( .A(n9867), .B(n9868), .Z(n9651) );
  XOR2_X1 U9660 ( .A(n9869), .B(n9870), .Z(n9868) );
  NAND2_X1 U9661 ( .A1(b_27_), .A2(a_7_), .ZN(n9870) );
  XNOR2_X1 U9662 ( .A(n9871), .B(n9872), .ZN(n9655) );
  XNOR2_X1 U9663 ( .A(n9873), .B(n9874), .ZN(n9871) );
  NOR2_X1 U9664 ( .A1(n8491), .A2(n8740), .ZN(n9874) );
  XNOR2_X1 U9665 ( .A(n9875), .B(n9876), .ZN(n9659) );
  XOR2_X1 U9666 ( .A(n9877), .B(n9878), .Z(n9875) );
  XNOR2_X1 U9667 ( .A(n9879), .B(n9880), .ZN(n9662) );
  XNOR2_X1 U9668 ( .A(n9881), .B(n9882), .ZN(n9879) );
  NOR2_X1 U9669 ( .A1(n8766), .A2(n8740), .ZN(n9882) );
  OR2_X1 U9670 ( .A1(n9669), .A2(n9667), .ZN(n9685) );
  XOR2_X1 U9671 ( .A(n9883), .B(n9884), .Z(n9667) );
  NAND2_X1 U9672 ( .A1(n9885), .A2(n9886), .ZN(n9883) );
  NAND2_X1 U9673 ( .A1(b_28_), .A2(a_2_), .ZN(n9669) );
  XNOR2_X1 U9674 ( .A(n9887), .B(n9888), .ZN(n9461) );
  NAND2_X1 U9675 ( .A1(n9889), .A2(n9890), .ZN(n9887) );
  XNOR2_X1 U9676 ( .A(n9891), .B(n9892), .ZN(n9671) );
  XOR2_X1 U9677 ( .A(n9893), .B(n9894), .Z(n9891) );
  NOR2_X1 U9678 ( .A1(n8617), .A2(n8740), .ZN(n9894) );
  XNOR2_X1 U9679 ( .A(n9895), .B(n9896), .ZN(n9008) );
  XNOR2_X1 U9680 ( .A(n9897), .B(n9898), .ZN(n9896) );
  NAND2_X1 U9681 ( .A1(n9899), .A2(n9676), .ZN(n8809) );
  INV_X1 U9682 ( .A(n9900), .ZN(n9676) );
  XOR2_X1 U9683 ( .A(n8998), .B(n9901), .Z(n9899) );
  NAND2_X1 U9684 ( .A1(n9902), .A2(n9900), .ZN(n8810) );
  NOR2_X1 U9685 ( .A1(n9678), .A2(n9677), .ZN(n9900) );
  XOR2_X1 U9686 ( .A(n9903), .B(n9904), .Z(n9677) );
  XNOR2_X1 U9687 ( .A(n9905), .B(n9906), .ZN(n9903) );
  NOR2_X1 U9688 ( .A1(n9674), .A2(n7992), .ZN(n9906) );
  NAND2_X1 U9689 ( .A1(n9907), .A2(n9908), .ZN(n9678) );
  NAND2_X1 U9690 ( .A1(n9897), .A2(n9909), .ZN(n9908) );
  OR2_X1 U9691 ( .A1(n9898), .A2(n9895), .ZN(n9909) );
  AND2_X1 U9692 ( .A1(n9910), .A2(n9911), .ZN(n9897) );
  NAND3_X1 U9693 ( .A1(a_1_), .A2(n9912), .A3(b_27_), .ZN(n9911) );
  OR2_X1 U9694 ( .A1(n9893), .A2(n9892), .ZN(n9912) );
  NAND2_X1 U9695 ( .A1(n9892), .A2(n9893), .ZN(n9910) );
  NAND2_X1 U9696 ( .A1(n9889), .A2(n9913), .ZN(n9893) );
  NAND2_X1 U9697 ( .A1(n9888), .A2(n9890), .ZN(n9913) );
  NAND2_X1 U9698 ( .A1(n9914), .A2(n9915), .ZN(n9890) );
  NAND2_X1 U9699 ( .A1(b_27_), .A2(a_2_), .ZN(n9915) );
  INV_X1 U9700 ( .A(n9916), .ZN(n9914) );
  XNOR2_X1 U9701 ( .A(n9917), .B(n9918), .ZN(n9888) );
  XNOR2_X1 U9702 ( .A(n9919), .B(n9920), .ZN(n9917) );
  NOR2_X1 U9703 ( .A1(n8567), .A2(n7992), .ZN(n9920) );
  NAND2_X1 U9704 ( .A1(a_2_), .A2(n9916), .ZN(n9889) );
  NAND2_X1 U9705 ( .A1(n9885), .A2(n9921), .ZN(n9916) );
  NAND2_X1 U9706 ( .A1(n9884), .A2(n9886), .ZN(n9921) );
  NAND2_X1 U9707 ( .A1(n9922), .A2(n9923), .ZN(n9886) );
  NAND2_X1 U9708 ( .A1(b_27_), .A2(a_3_), .ZN(n9923) );
  INV_X1 U9709 ( .A(n9924), .ZN(n9922) );
  XNOR2_X1 U9710 ( .A(n9925), .B(n9926), .ZN(n9884) );
  XNOR2_X1 U9711 ( .A(n9927), .B(n9928), .ZN(n9926) );
  NAND2_X1 U9712 ( .A1(a_3_), .A2(n9924), .ZN(n9885) );
  NAND2_X1 U9713 ( .A1(n9929), .A2(n9930), .ZN(n9924) );
  NAND3_X1 U9714 ( .A1(a_4_), .A2(n9931), .A3(b_27_), .ZN(n9930) );
  NAND2_X1 U9715 ( .A1(n9881), .A2(n9880), .ZN(n9931) );
  OR2_X1 U9716 ( .A1(n9880), .A2(n9881), .ZN(n9929) );
  AND2_X1 U9717 ( .A1(n9932), .A2(n9933), .ZN(n9881) );
  NAND2_X1 U9718 ( .A1(n9878), .A2(n9934), .ZN(n9933) );
  OR2_X1 U9719 ( .A1(n9877), .A2(n9876), .ZN(n9934) );
  NOR2_X1 U9720 ( .A1(n8740), .A2(n8517), .ZN(n9878) );
  NAND2_X1 U9721 ( .A1(n9876), .A2(n9877), .ZN(n9932) );
  NAND2_X1 U9722 ( .A1(n9935), .A2(n9936), .ZN(n9877) );
  NAND3_X1 U9723 ( .A1(a_6_), .A2(n9937), .A3(b_27_), .ZN(n9936) );
  NAND2_X1 U9724 ( .A1(n9873), .A2(n9872), .ZN(n9937) );
  OR2_X1 U9725 ( .A1(n9872), .A2(n9873), .ZN(n9935) );
  AND2_X1 U9726 ( .A1(n9938), .A2(n9939), .ZN(n9873) );
  NAND3_X1 U9727 ( .A1(a_7_), .A2(n9940), .A3(b_27_), .ZN(n9939) );
  OR2_X1 U9728 ( .A1(n9869), .A2(n9867), .ZN(n9940) );
  NAND2_X1 U9729 ( .A1(n9867), .A2(n9869), .ZN(n9938) );
  NAND2_X1 U9730 ( .A1(n9941), .A2(n9942), .ZN(n9869) );
  NAND3_X1 U9731 ( .A1(a_8_), .A2(n9943), .A3(b_27_), .ZN(n9942) );
  NAND2_X1 U9732 ( .A1(n9865), .A2(n9864), .ZN(n9943) );
  OR2_X1 U9733 ( .A1(n9864), .A2(n9865), .ZN(n9941) );
  AND2_X1 U9734 ( .A1(n9944), .A2(n9945), .ZN(n9865) );
  NAND2_X1 U9735 ( .A1(n9862), .A2(n9946), .ZN(n9945) );
  OR2_X1 U9736 ( .A1(n9861), .A2(n9860), .ZN(n9946) );
  NOR2_X1 U9737 ( .A1(n8740), .A2(n8426), .ZN(n9862) );
  NAND2_X1 U9738 ( .A1(n9860), .A2(n9861), .ZN(n9944) );
  NAND2_X1 U9739 ( .A1(n9947), .A2(n9948), .ZN(n9861) );
  NAND3_X1 U9740 ( .A1(a_10_), .A2(n9949), .A3(b_27_), .ZN(n9948) );
  OR2_X1 U9741 ( .A1(n9857), .A2(n9856), .ZN(n9949) );
  NAND2_X1 U9742 ( .A1(n9856), .A2(n9857), .ZN(n9947) );
  NAND2_X1 U9743 ( .A1(n9950), .A2(n9951), .ZN(n9857) );
  NAND2_X1 U9744 ( .A1(n9854), .A2(n9952), .ZN(n9951) );
  OR2_X1 U9745 ( .A1(n9853), .A2(n9851), .ZN(n9952) );
  NOR2_X1 U9746 ( .A1(n8740), .A2(n8376), .ZN(n9854) );
  NAND2_X1 U9747 ( .A1(n9851), .A2(n9853), .ZN(n9950) );
  NAND2_X1 U9748 ( .A1(n9953), .A2(n9954), .ZN(n9853) );
  NAND3_X1 U9749 ( .A1(a_12_), .A2(n9955), .A3(b_27_), .ZN(n9954) );
  NAND2_X1 U9750 ( .A1(n9849), .A2(n9848), .ZN(n9955) );
  OR2_X1 U9751 ( .A1(n9848), .A2(n9849), .ZN(n9953) );
  AND2_X1 U9752 ( .A1(n9956), .A2(n9957), .ZN(n9849) );
  NAND2_X1 U9753 ( .A1(n9846), .A2(n9958), .ZN(n9957) );
  NAND2_X1 U9754 ( .A1(n9845), .A2(n9844), .ZN(n9958) );
  NOR2_X1 U9755 ( .A1(n8740), .A2(n8310), .ZN(n9846) );
  OR2_X1 U9756 ( .A1(n9844), .A2(n9845), .ZN(n9956) );
  AND2_X1 U9757 ( .A1(n9959), .A2(n9960), .ZN(n9845) );
  NAND3_X1 U9758 ( .A1(a_14_), .A2(n9961), .A3(b_27_), .ZN(n9960) );
  NAND2_X1 U9759 ( .A1(n9842), .A2(n9840), .ZN(n9961) );
  OR2_X1 U9760 ( .A1(n9840), .A2(n9842), .ZN(n9959) );
  AND2_X1 U9761 ( .A1(n9962), .A2(n9963), .ZN(n9842) );
  NAND2_X1 U9762 ( .A1(n9838), .A2(n9964), .ZN(n9963) );
  OR2_X1 U9763 ( .A1(n9837), .A2(n9835), .ZN(n9964) );
  NOR2_X1 U9764 ( .A1(n8740), .A2(n8276), .ZN(n9838) );
  NAND2_X1 U9765 ( .A1(n9835), .A2(n9837), .ZN(n9962) );
  NAND2_X1 U9766 ( .A1(n9965), .A2(n9966), .ZN(n9837) );
  NAND3_X1 U9767 ( .A1(a_16_), .A2(n9967), .A3(b_27_), .ZN(n9966) );
  NAND2_X1 U9768 ( .A1(n9833), .A2(n9832), .ZN(n9967) );
  OR2_X1 U9769 ( .A1(n9832), .A2(n9833), .ZN(n9965) );
  AND2_X1 U9770 ( .A1(n9968), .A2(n9969), .ZN(n9833) );
  NAND2_X1 U9771 ( .A1(n9830), .A2(n9970), .ZN(n9969) );
  OR2_X1 U9772 ( .A1(n9829), .A2(n9828), .ZN(n9970) );
  NOR2_X1 U9773 ( .A1(n8740), .A2(n8210), .ZN(n9830) );
  NAND2_X1 U9774 ( .A1(n9828), .A2(n9829), .ZN(n9968) );
  NAND2_X1 U9775 ( .A1(n9971), .A2(n9972), .ZN(n9829) );
  NAND3_X1 U9776 ( .A1(a_18_), .A2(n9973), .A3(b_27_), .ZN(n9972) );
  NAND2_X1 U9777 ( .A1(n9825), .A2(n9824), .ZN(n9973) );
  OR2_X1 U9778 ( .A1(n9824), .A2(n9825), .ZN(n9971) );
  AND2_X1 U9779 ( .A1(n9974), .A2(n9975), .ZN(n9825) );
  NAND2_X1 U9780 ( .A1(n9822), .A2(n9976), .ZN(n9975) );
  OR2_X1 U9781 ( .A1(n9821), .A2(n9819), .ZN(n9976) );
  NOR2_X1 U9782 ( .A1(n8740), .A2(n8170), .ZN(n9822) );
  NAND2_X1 U9783 ( .A1(n9819), .A2(n9821), .ZN(n9974) );
  NAND2_X1 U9784 ( .A1(n9977), .A2(n9978), .ZN(n9821) );
  NAND3_X1 U9785 ( .A1(a_20_), .A2(n9979), .A3(b_27_), .ZN(n9978) );
  NAND2_X1 U9786 ( .A1(n9817), .A2(n9816), .ZN(n9979) );
  OR2_X1 U9787 ( .A1(n9816), .A2(n9817), .ZN(n9977) );
  AND2_X1 U9788 ( .A1(n9980), .A2(n9981), .ZN(n9817) );
  NAND2_X1 U9789 ( .A1(n9814), .A2(n9982), .ZN(n9981) );
  OR2_X1 U9790 ( .A1(n9813), .A2(n9812), .ZN(n9982) );
  NOR2_X1 U9791 ( .A1(n8740), .A2(n8750), .ZN(n9814) );
  NAND2_X1 U9792 ( .A1(n9812), .A2(n9813), .ZN(n9980) );
  NAND2_X1 U9793 ( .A1(n9983), .A2(n9984), .ZN(n9813) );
  NAND3_X1 U9794 ( .A1(a_22_), .A2(n9985), .A3(b_27_), .ZN(n9984) );
  OR2_X1 U9795 ( .A1(n9809), .A2(n9807), .ZN(n9985) );
  NAND2_X1 U9796 ( .A1(n9807), .A2(n9809), .ZN(n9983) );
  NAND2_X1 U9797 ( .A1(n9986), .A2(n9987), .ZN(n9809) );
  NAND2_X1 U9798 ( .A1(n9806), .A2(n9988), .ZN(n9987) );
  OR2_X1 U9799 ( .A1(n9805), .A2(n9803), .ZN(n9988) );
  NOR2_X1 U9800 ( .A1(n8740), .A2(n8747), .ZN(n9806) );
  NAND2_X1 U9801 ( .A1(n9803), .A2(n9805), .ZN(n9986) );
  NAND2_X1 U9802 ( .A1(n9989), .A2(n9990), .ZN(n9805) );
  NAND3_X1 U9803 ( .A1(a_24_), .A2(n9991), .A3(b_27_), .ZN(n9990) );
  NAND2_X1 U9804 ( .A1(n9801), .A2(n9800), .ZN(n9991) );
  OR2_X1 U9805 ( .A1(n9800), .A2(n9801), .ZN(n9989) );
  AND2_X1 U9806 ( .A1(n9992), .A2(n9993), .ZN(n9801) );
  NAND2_X1 U9807 ( .A1(n9798), .A2(n9994), .ZN(n9993) );
  NAND2_X1 U9808 ( .A1(n9797), .A2(n9796), .ZN(n9994) );
  NOR2_X1 U9809 ( .A1(n8740), .A2(n8744), .ZN(n9798) );
  OR2_X1 U9810 ( .A1(n9796), .A2(n9797), .ZN(n9992) );
  AND2_X1 U9811 ( .A1(n9793), .A2(n9995), .ZN(n9797) );
  NAND2_X1 U9812 ( .A1(n9792), .A2(n9794), .ZN(n9995) );
  NAND2_X1 U9813 ( .A1(n9996), .A2(n9997), .ZN(n9794) );
  NAND2_X1 U9814 ( .A1(b_27_), .A2(a_26_), .ZN(n9997) );
  INV_X1 U9815 ( .A(n9998), .ZN(n9996) );
  XNOR2_X1 U9816 ( .A(n9999), .B(n10000), .ZN(n9792) );
  NAND2_X1 U9817 ( .A1(n10001), .A2(n10002), .ZN(n9999) );
  NAND2_X1 U9818 ( .A1(a_26_), .A2(n9998), .ZN(n9793) );
  NAND2_X1 U9819 ( .A1(n10003), .A2(n10004), .ZN(n9998) );
  NAND2_X1 U9820 ( .A1(n9762), .A2(n10005), .ZN(n10004) );
  OR2_X1 U9821 ( .A1(n9763), .A2(n9764), .ZN(n10005) );
  XNOR2_X1 U9822 ( .A(n10006), .B(n10007), .ZN(n9762) );
  XOR2_X1 U9823 ( .A(n10008), .B(n10009), .Z(n10006) );
  NAND2_X1 U9824 ( .A1(b_26_), .A2(a_28_), .ZN(n10008) );
  NAND2_X1 U9825 ( .A1(n9764), .A2(n9763), .ZN(n10003) );
  NAND2_X1 U9826 ( .A1(n10010), .A2(n10011), .ZN(n9763) );
  NAND3_X1 U9827 ( .A1(a_28_), .A2(n10012), .A3(b_27_), .ZN(n10011) );
  NAND2_X1 U9828 ( .A1(n9772), .A2(n9770), .ZN(n10012) );
  OR2_X1 U9829 ( .A1(n9770), .A2(n9772), .ZN(n10010) );
  AND2_X1 U9830 ( .A1(n10013), .A2(n10014), .ZN(n9772) );
  NAND2_X1 U9831 ( .A1(n9778), .A2(n10015), .ZN(n10014) );
  OR2_X1 U9832 ( .A1(n9779), .A2(n9780), .ZN(n10015) );
  NOR2_X1 U9833 ( .A1(n8740), .A2(n7890), .ZN(n9778) );
  NAND2_X1 U9834 ( .A1(n9780), .A2(n9779), .ZN(n10013) );
  NAND2_X1 U9835 ( .A1(n10016), .A2(n10017), .ZN(n9779) );
  NAND2_X1 U9836 ( .A1(b_25_), .A2(n10018), .ZN(n10017) );
  NAND2_X1 U9837 ( .A1(n7864), .A2(n10019), .ZN(n10018) );
  NAND2_X1 U9838 ( .A1(a_31_), .A2(n7992), .ZN(n10019) );
  NAND2_X1 U9839 ( .A1(b_26_), .A2(n10020), .ZN(n10016) );
  NAND2_X1 U9840 ( .A1(n9137), .A2(n10021), .ZN(n10020) );
  NAND2_X1 U9841 ( .A1(a_30_), .A2(n8743), .ZN(n10021) );
  AND3_X1 U9842 ( .A1(b_26_), .A2(b_27_), .A3(n7818), .ZN(n9780) );
  XNOR2_X1 U9843 ( .A(n10022), .B(n10023), .ZN(n9770) );
  XOR2_X1 U9844 ( .A(n10024), .B(n10025), .Z(n10022) );
  INV_X1 U9845 ( .A(n7966), .ZN(n9764) );
  NAND2_X1 U9846 ( .A1(b_27_), .A2(a_27_), .ZN(n7966) );
  XNOR2_X1 U9847 ( .A(n10026), .B(n10027), .ZN(n9796) );
  XOR2_X1 U9848 ( .A(n10028), .B(n10029), .Z(n10026) );
  XNOR2_X1 U9849 ( .A(n10030), .B(n10031), .ZN(n9800) );
  XOR2_X1 U9850 ( .A(n10032), .B(n10033), .Z(n10030) );
  XNOR2_X1 U9851 ( .A(n10034), .B(n10035), .ZN(n9803) );
  XNOR2_X1 U9852 ( .A(n10036), .B(n10037), .ZN(n10034) );
  NOR2_X1 U9853 ( .A1(n8745), .A2(n7992), .ZN(n10037) );
  XNOR2_X1 U9854 ( .A(n10038), .B(n10039), .ZN(n9807) );
  XNOR2_X1 U9855 ( .A(n10040), .B(n10041), .ZN(n10039) );
  XNOR2_X1 U9856 ( .A(n10042), .B(n10043), .ZN(n9812) );
  XOR2_X1 U9857 ( .A(n10044), .B(n10045), .Z(n10043) );
  NAND2_X1 U9858 ( .A1(b_26_), .A2(a_22_), .ZN(n10045) );
  XNOR2_X1 U9859 ( .A(n10046), .B(n10047), .ZN(n9816) );
  XOR2_X1 U9860 ( .A(n10048), .B(n10049), .Z(n10046) );
  XNOR2_X1 U9861 ( .A(n10050), .B(n10051), .ZN(n9819) );
  XNOR2_X1 U9862 ( .A(n10052), .B(n10053), .ZN(n10050) );
  NOR2_X1 U9863 ( .A1(n8751), .A2(n7992), .ZN(n10053) );
  XOR2_X1 U9864 ( .A(n10054), .B(n10055), .Z(n9824) );
  XNOR2_X1 U9865 ( .A(n10056), .B(n10057), .ZN(n10055) );
  XNOR2_X1 U9866 ( .A(n10058), .B(n10059), .ZN(n9828) );
  XNOR2_X1 U9867 ( .A(n10060), .B(n10061), .ZN(n10058) );
  NOR2_X1 U9868 ( .A1(n8753), .A2(n7992), .ZN(n10061) );
  XNOR2_X1 U9869 ( .A(n10062), .B(n10063), .ZN(n9832) );
  XOR2_X1 U9870 ( .A(n10064), .B(n10065), .Z(n10062) );
  XNOR2_X1 U9871 ( .A(n10066), .B(n10067), .ZN(n9835) );
  XOR2_X1 U9872 ( .A(n10068), .B(n10069), .Z(n10067) );
  NAND2_X1 U9873 ( .A1(b_26_), .A2(a_16_), .ZN(n10069) );
  XOR2_X1 U9874 ( .A(n10070), .B(n10071), .Z(n9840) );
  XNOR2_X1 U9875 ( .A(n10072), .B(n10073), .ZN(n10071) );
  XNOR2_X1 U9876 ( .A(n10074), .B(n10075), .ZN(n9844) );
  XNOR2_X1 U9877 ( .A(n10076), .B(n10077), .ZN(n10074) );
  NAND2_X1 U9878 ( .A1(b_26_), .A2(a_14_), .ZN(n10076) );
  XNOR2_X1 U9879 ( .A(n10078), .B(n10079), .ZN(n9848) );
  XOR2_X1 U9880 ( .A(n10080), .B(n10081), .Z(n10078) );
  XNOR2_X1 U9881 ( .A(n10082), .B(n10083), .ZN(n9851) );
  XNOR2_X1 U9882 ( .A(n10084), .B(n10085), .ZN(n10082) );
  NOR2_X1 U9883 ( .A1(n8759), .A2(n7992), .ZN(n10085) );
  XNOR2_X1 U9884 ( .A(n10086), .B(n10087), .ZN(n9856) );
  XNOR2_X1 U9885 ( .A(n10088), .B(n10089), .ZN(n10087) );
  XNOR2_X1 U9886 ( .A(n10090), .B(n10091), .ZN(n9860) );
  XNOR2_X1 U9887 ( .A(n10092), .B(n10093), .ZN(n10090) );
  NOR2_X1 U9888 ( .A1(n8761), .A2(n7992), .ZN(n10093) );
  XNOR2_X1 U9889 ( .A(n10094), .B(n10095), .ZN(n9864) );
  XOR2_X1 U9890 ( .A(n10096), .B(n10097), .Z(n10094) );
  XNOR2_X1 U9891 ( .A(n10098), .B(n10099), .ZN(n9867) );
  XOR2_X1 U9892 ( .A(n10100), .B(n10101), .Z(n10099) );
  NAND2_X1 U9893 ( .A1(b_26_), .A2(a_8_), .ZN(n10101) );
  XOR2_X1 U9894 ( .A(n10102), .B(n10103), .Z(n9872) );
  NAND2_X1 U9895 ( .A1(n10104), .A2(n10105), .ZN(n10102) );
  XNOR2_X1 U9896 ( .A(n10106), .B(n10107), .ZN(n9876) );
  XNOR2_X1 U9897 ( .A(n10108), .B(n10109), .ZN(n10106) );
  NOR2_X1 U9898 ( .A1(n8491), .A2(n7992), .ZN(n10109) );
  XOR2_X1 U9899 ( .A(n10110), .B(n10111), .Z(n9880) );
  XOR2_X1 U9900 ( .A(n10112), .B(n10113), .Z(n10111) );
  NAND2_X1 U9901 ( .A1(b_26_), .A2(a_5_), .ZN(n10113) );
  XNOR2_X1 U9902 ( .A(n10114), .B(n10115), .ZN(n9892) );
  XNOR2_X1 U9903 ( .A(n10116), .B(n10117), .ZN(n10115) );
  NAND2_X1 U9904 ( .A1(n9895), .A2(n9898), .ZN(n9907) );
  NAND2_X1 U9905 ( .A1(b_27_), .A2(a_0_), .ZN(n9898) );
  XOR2_X1 U9906 ( .A(n10118), .B(n10119), .Z(n9895) );
  XNOR2_X1 U9907 ( .A(n10120), .B(n10121), .ZN(n10118) );
  XOR2_X1 U9908 ( .A(n8998), .B(n8997), .Z(n9902) );
  NAND4_X1 U9909 ( .A1(n8997), .A2(n8996), .A3(n8998), .A4(n8991), .ZN(n8815)
         );
  INV_X1 U9910 ( .A(n10122), .ZN(n8991) );
  NAND2_X1 U9911 ( .A1(n10123), .A2(n10124), .ZN(n8998) );
  NAND3_X1 U9912 ( .A1(a_0_), .A2(n10125), .A3(b_26_), .ZN(n10124) );
  NAND2_X1 U9913 ( .A1(n9905), .A2(n9904), .ZN(n10125) );
  OR2_X1 U9914 ( .A1(n9904), .A2(n9905), .ZN(n10123) );
  AND2_X1 U9915 ( .A1(n10126), .A2(n10127), .ZN(n9905) );
  NAND2_X1 U9916 ( .A1(n10121), .A2(n10128), .ZN(n10127) );
  NAND2_X1 U9917 ( .A1(n10120), .A2(n10119), .ZN(n10128) );
  NOR2_X1 U9918 ( .A1(n7992), .A2(n8617), .ZN(n10121) );
  OR2_X1 U9919 ( .A1(n10119), .A2(n10120), .ZN(n10126) );
  AND2_X1 U9920 ( .A1(n10129), .A2(n10130), .ZN(n10120) );
  NAND2_X1 U9921 ( .A1(n10117), .A2(n10131), .ZN(n10130) );
  OR2_X1 U9922 ( .A1(n10116), .A2(n10114), .ZN(n10131) );
  NOR2_X1 U9923 ( .A1(n7992), .A2(n8768), .ZN(n10117) );
  NAND2_X1 U9924 ( .A1(n10114), .A2(n10116), .ZN(n10129) );
  NAND2_X1 U9925 ( .A1(n10132), .A2(n10133), .ZN(n10116) );
  NAND3_X1 U9926 ( .A1(a_3_), .A2(n10134), .A3(b_26_), .ZN(n10133) );
  NAND2_X1 U9927 ( .A1(n9919), .A2(n9918), .ZN(n10134) );
  OR2_X1 U9928 ( .A1(n9918), .A2(n9919), .ZN(n10132) );
  AND2_X1 U9929 ( .A1(n10135), .A2(n10136), .ZN(n9919) );
  NAND2_X1 U9930 ( .A1(n9928), .A2(n10137), .ZN(n10136) );
  OR2_X1 U9931 ( .A1(n9927), .A2(n9925), .ZN(n10137) );
  NOR2_X1 U9932 ( .A1(n7992), .A2(n8766), .ZN(n9928) );
  NAND2_X1 U9933 ( .A1(n9925), .A2(n9927), .ZN(n10135) );
  NAND2_X1 U9934 ( .A1(n10138), .A2(n10139), .ZN(n9927) );
  NAND3_X1 U9935 ( .A1(a_5_), .A2(n10140), .A3(b_26_), .ZN(n10139) );
  OR2_X1 U9936 ( .A1(n10112), .A2(n10110), .ZN(n10140) );
  NAND2_X1 U9937 ( .A1(n10110), .A2(n10112), .ZN(n10138) );
  NAND2_X1 U9938 ( .A1(n10141), .A2(n10142), .ZN(n10112) );
  NAND3_X1 U9939 ( .A1(a_6_), .A2(n10143), .A3(b_26_), .ZN(n10142) );
  NAND2_X1 U9940 ( .A1(n10108), .A2(n10107), .ZN(n10143) );
  OR2_X1 U9941 ( .A1(n10107), .A2(n10108), .ZN(n10141) );
  AND2_X1 U9942 ( .A1(n10104), .A2(n10144), .ZN(n10108) );
  NAND2_X1 U9943 ( .A1(n10103), .A2(n10105), .ZN(n10144) );
  NAND2_X1 U9944 ( .A1(n10145), .A2(n10146), .ZN(n10105) );
  NAND2_X1 U9945 ( .A1(b_26_), .A2(a_7_), .ZN(n10146) );
  INV_X1 U9946 ( .A(n10147), .ZN(n10145) );
  XOR2_X1 U9947 ( .A(n10148), .B(n10149), .Z(n10103) );
  XOR2_X1 U9948 ( .A(n10150), .B(n10151), .Z(n10148) );
  NOR2_X1 U9949 ( .A1(n8763), .A2(n8743), .ZN(n10151) );
  NAND2_X1 U9950 ( .A1(a_7_), .A2(n10147), .ZN(n10104) );
  NAND2_X1 U9951 ( .A1(n10152), .A2(n10153), .ZN(n10147) );
  NAND3_X1 U9952 ( .A1(a_8_), .A2(n10154), .A3(b_26_), .ZN(n10153) );
  OR2_X1 U9953 ( .A1(n10100), .A2(n10098), .ZN(n10154) );
  NAND2_X1 U9954 ( .A1(n10098), .A2(n10100), .ZN(n10152) );
  NAND2_X1 U9955 ( .A1(n10155), .A2(n10156), .ZN(n10100) );
  NAND2_X1 U9956 ( .A1(n10097), .A2(n10157), .ZN(n10156) );
  OR2_X1 U9957 ( .A1(n10096), .A2(n10095), .ZN(n10157) );
  NOR2_X1 U9958 ( .A1(n7992), .A2(n8426), .ZN(n10097) );
  NAND2_X1 U9959 ( .A1(n10095), .A2(n10096), .ZN(n10155) );
  NAND2_X1 U9960 ( .A1(n10158), .A2(n10159), .ZN(n10096) );
  NAND3_X1 U9961 ( .A1(a_10_), .A2(n10160), .A3(b_26_), .ZN(n10159) );
  NAND2_X1 U9962 ( .A1(n10092), .A2(n10091), .ZN(n10160) );
  OR2_X1 U9963 ( .A1(n10091), .A2(n10092), .ZN(n10158) );
  AND2_X1 U9964 ( .A1(n10161), .A2(n10162), .ZN(n10092) );
  NAND2_X1 U9965 ( .A1(n10089), .A2(n10163), .ZN(n10162) );
  OR2_X1 U9966 ( .A1(n10088), .A2(n10086), .ZN(n10163) );
  NOR2_X1 U9967 ( .A1(n7992), .A2(n8376), .ZN(n10089) );
  NAND2_X1 U9968 ( .A1(n10086), .A2(n10088), .ZN(n10161) );
  NAND2_X1 U9969 ( .A1(n10164), .A2(n10165), .ZN(n10088) );
  NAND3_X1 U9970 ( .A1(a_12_), .A2(n10166), .A3(b_26_), .ZN(n10165) );
  NAND2_X1 U9971 ( .A1(n10084), .A2(n10083), .ZN(n10166) );
  OR2_X1 U9972 ( .A1(n10083), .A2(n10084), .ZN(n10164) );
  AND2_X1 U9973 ( .A1(n10167), .A2(n10168), .ZN(n10084) );
  NAND2_X1 U9974 ( .A1(n10081), .A2(n10169), .ZN(n10168) );
  OR2_X1 U9975 ( .A1(n10080), .A2(n10079), .ZN(n10169) );
  NOR2_X1 U9976 ( .A1(n7992), .A2(n8310), .ZN(n10081) );
  NAND2_X1 U9977 ( .A1(n10079), .A2(n10080), .ZN(n10167) );
  NAND2_X1 U9978 ( .A1(n10170), .A2(n10171), .ZN(n10080) );
  NAND3_X1 U9979 ( .A1(a_14_), .A2(n10172), .A3(b_26_), .ZN(n10171) );
  OR2_X1 U9980 ( .A1(n10077), .A2(n10075), .ZN(n10172) );
  NAND2_X1 U9981 ( .A1(n10075), .A2(n10077), .ZN(n10170) );
  NAND2_X1 U9982 ( .A1(n10173), .A2(n10174), .ZN(n10077) );
  NAND2_X1 U9983 ( .A1(n10073), .A2(n10175), .ZN(n10174) );
  OR2_X1 U9984 ( .A1(n10072), .A2(n10070), .ZN(n10175) );
  NOR2_X1 U9985 ( .A1(n7992), .A2(n8276), .ZN(n10073) );
  NAND2_X1 U9986 ( .A1(n10070), .A2(n10072), .ZN(n10173) );
  NAND2_X1 U9987 ( .A1(n10176), .A2(n10177), .ZN(n10072) );
  NAND3_X1 U9988 ( .A1(a_16_), .A2(n10178), .A3(b_26_), .ZN(n10177) );
  OR2_X1 U9989 ( .A1(n10068), .A2(n10066), .ZN(n10178) );
  NAND2_X1 U9990 ( .A1(n10066), .A2(n10068), .ZN(n10176) );
  NAND2_X1 U9991 ( .A1(n10179), .A2(n10180), .ZN(n10068) );
  NAND2_X1 U9992 ( .A1(n10065), .A2(n10181), .ZN(n10180) );
  OR2_X1 U9993 ( .A1(n10064), .A2(n10063), .ZN(n10181) );
  NOR2_X1 U9994 ( .A1(n7992), .A2(n8210), .ZN(n10065) );
  NAND2_X1 U9995 ( .A1(n10063), .A2(n10064), .ZN(n10179) );
  NAND2_X1 U9996 ( .A1(n10182), .A2(n10183), .ZN(n10064) );
  NAND3_X1 U9997 ( .A1(a_18_), .A2(n10184), .A3(b_26_), .ZN(n10183) );
  NAND2_X1 U9998 ( .A1(n10060), .A2(n10059), .ZN(n10184) );
  OR2_X1 U9999 ( .A1(n10059), .A2(n10060), .ZN(n10182) );
  AND2_X1 U10000 ( .A1(n10185), .A2(n10186), .ZN(n10060) );
  NAND2_X1 U10001 ( .A1(n10057), .A2(n10187), .ZN(n10186) );
  OR2_X1 U10002 ( .A1(n10056), .A2(n10054), .ZN(n10187) );
  NOR2_X1 U10003 ( .A1(n7992), .A2(n8170), .ZN(n10057) );
  NAND2_X1 U10004 ( .A1(n10054), .A2(n10056), .ZN(n10185) );
  NAND2_X1 U10005 ( .A1(n10188), .A2(n10189), .ZN(n10056) );
  NAND3_X1 U10006 ( .A1(a_20_), .A2(n10190), .A3(b_26_), .ZN(n10189) );
  NAND2_X1 U10007 ( .A1(n10052), .A2(n10051), .ZN(n10190) );
  OR2_X1 U10008 ( .A1(n10051), .A2(n10052), .ZN(n10188) );
  AND2_X1 U10009 ( .A1(n10191), .A2(n10192), .ZN(n10052) );
  NAND2_X1 U10010 ( .A1(n10049), .A2(n10193), .ZN(n10192) );
  OR2_X1 U10011 ( .A1(n10048), .A2(n10047), .ZN(n10193) );
  NOR2_X1 U10012 ( .A1(n7992), .A2(n8750), .ZN(n10049) );
  NAND2_X1 U10013 ( .A1(n10047), .A2(n10048), .ZN(n10191) );
  NAND2_X1 U10014 ( .A1(n10194), .A2(n10195), .ZN(n10048) );
  NAND3_X1 U10015 ( .A1(a_22_), .A2(n10196), .A3(b_26_), .ZN(n10195) );
  OR2_X1 U10016 ( .A1(n10044), .A2(n10042), .ZN(n10196) );
  NAND2_X1 U10017 ( .A1(n10042), .A2(n10044), .ZN(n10194) );
  NAND2_X1 U10018 ( .A1(n10197), .A2(n10198), .ZN(n10044) );
  NAND2_X1 U10019 ( .A1(n10041), .A2(n10199), .ZN(n10198) );
  OR2_X1 U10020 ( .A1(n10040), .A2(n10038), .ZN(n10199) );
  NOR2_X1 U10021 ( .A1(n7992), .A2(n8747), .ZN(n10041) );
  NAND2_X1 U10022 ( .A1(n10038), .A2(n10040), .ZN(n10197) );
  NAND2_X1 U10023 ( .A1(n10200), .A2(n10201), .ZN(n10040) );
  NAND3_X1 U10024 ( .A1(a_24_), .A2(n10202), .A3(b_26_), .ZN(n10201) );
  NAND2_X1 U10025 ( .A1(n10036), .A2(n10035), .ZN(n10202) );
  OR2_X1 U10026 ( .A1(n10035), .A2(n10036), .ZN(n10200) );
  AND2_X1 U10027 ( .A1(n10203), .A2(n10204), .ZN(n10036) );
  NAND2_X1 U10028 ( .A1(n10033), .A2(n10205), .ZN(n10204) );
  OR2_X1 U10029 ( .A1(n10032), .A2(n10031), .ZN(n10205) );
  NOR2_X1 U10030 ( .A1(n7992), .A2(n8744), .ZN(n10033) );
  NAND2_X1 U10031 ( .A1(n10031), .A2(n10032), .ZN(n10203) );
  NAND2_X1 U10032 ( .A1(n10206), .A2(n10207), .ZN(n10032) );
  NAND2_X1 U10033 ( .A1(n10027), .A2(n10208), .ZN(n10207) );
  OR2_X1 U10034 ( .A1(n10028), .A2(n10029), .ZN(n10208) );
  XNOR2_X1 U10035 ( .A(n10209), .B(n10210), .ZN(n10027) );
  NAND2_X1 U10036 ( .A1(n10211), .A2(n10212), .ZN(n10209) );
  NAND2_X1 U10037 ( .A1(n10029), .A2(n10028), .ZN(n10206) );
  NAND2_X1 U10038 ( .A1(n10001), .A2(n10213), .ZN(n10028) );
  NAND2_X1 U10039 ( .A1(n10000), .A2(n10002), .ZN(n10213) );
  NAND2_X1 U10040 ( .A1(n10214), .A2(n10215), .ZN(n10002) );
  NAND2_X1 U10041 ( .A1(b_26_), .A2(a_27_), .ZN(n10215) );
  INV_X1 U10042 ( .A(n10216), .ZN(n10214) );
  XNOR2_X1 U10043 ( .A(n10217), .B(n10218), .ZN(n10000) );
  XOR2_X1 U10044 ( .A(n10219), .B(n10220), .Z(n10217) );
  NAND2_X1 U10045 ( .A1(b_25_), .A2(a_28_), .ZN(n10219) );
  NAND2_X1 U10046 ( .A1(a_27_), .A2(n10216), .ZN(n10001) );
  NAND2_X1 U10047 ( .A1(n10221), .A2(n10222), .ZN(n10216) );
  NAND3_X1 U10048 ( .A1(a_28_), .A2(n10223), .A3(b_26_), .ZN(n10222) );
  NAND2_X1 U10049 ( .A1(n10009), .A2(n10007), .ZN(n10223) );
  OR2_X1 U10050 ( .A1(n10007), .A2(n10009), .ZN(n10221) );
  AND2_X1 U10051 ( .A1(n10224), .A2(n10225), .ZN(n10009) );
  NAND2_X1 U10052 ( .A1(n10023), .A2(n10226), .ZN(n10225) );
  OR2_X1 U10053 ( .A1(n10024), .A2(n10025), .ZN(n10226) );
  NOR2_X1 U10054 ( .A1(n7992), .A2(n7890), .ZN(n10023) );
  NAND2_X1 U10055 ( .A1(n10025), .A2(n10024), .ZN(n10224) );
  NAND2_X1 U10056 ( .A1(n10227), .A2(n10228), .ZN(n10024) );
  NAND2_X1 U10057 ( .A1(b_24_), .A2(n10229), .ZN(n10228) );
  NAND2_X1 U10058 ( .A1(n7864), .A2(n10230), .ZN(n10229) );
  NAND2_X1 U10059 ( .A1(a_31_), .A2(n8743), .ZN(n10230) );
  NAND2_X1 U10060 ( .A1(b_25_), .A2(n10231), .ZN(n10227) );
  NAND2_X1 U10061 ( .A1(n9137), .A2(n10232), .ZN(n10231) );
  NAND2_X1 U10062 ( .A1(a_30_), .A2(n8043), .ZN(n10232) );
  AND3_X1 U10063 ( .A1(b_25_), .A2(b_26_), .A3(n7818), .ZN(n10025) );
  XNOR2_X1 U10064 ( .A(n10233), .B(n10234), .ZN(n10007) );
  XOR2_X1 U10065 ( .A(n10235), .B(n10236), .Z(n10233) );
  INV_X1 U10066 ( .A(n8727), .ZN(n10029) );
  NAND2_X1 U10067 ( .A1(b_26_), .A2(a_26_), .ZN(n8727) );
  XNOR2_X1 U10068 ( .A(n10237), .B(n10238), .ZN(n10031) );
  NAND2_X1 U10069 ( .A1(n10239), .A2(n10240), .ZN(n10237) );
  XNOR2_X1 U10070 ( .A(n10241), .B(n10242), .ZN(n10035) );
  XOR2_X1 U10071 ( .A(n10243), .B(n10244), .Z(n10241) );
  XNOR2_X1 U10072 ( .A(n10245), .B(n10246), .ZN(n10038) );
  XNOR2_X1 U10073 ( .A(n10247), .B(n10248), .ZN(n10245) );
  NOR2_X1 U10074 ( .A1(n8745), .A2(n8743), .ZN(n10248) );
  XNOR2_X1 U10075 ( .A(n10249), .B(n10250), .ZN(n10042) );
  XNOR2_X1 U10076 ( .A(n10251), .B(n10252), .ZN(n10250) );
  XNOR2_X1 U10077 ( .A(n10253), .B(n10254), .ZN(n10047) );
  XOR2_X1 U10078 ( .A(n10255), .B(n10256), .Z(n10254) );
  NAND2_X1 U10079 ( .A1(b_25_), .A2(a_22_), .ZN(n10256) );
  XNOR2_X1 U10080 ( .A(n10257), .B(n10258), .ZN(n10051) );
  XOR2_X1 U10081 ( .A(n10259), .B(n10260), .Z(n10257) );
  XNOR2_X1 U10082 ( .A(n10261), .B(n10262), .ZN(n10054) );
  XNOR2_X1 U10083 ( .A(n10263), .B(n10264), .ZN(n10261) );
  NOR2_X1 U10084 ( .A1(n8751), .A2(n8743), .ZN(n10264) );
  XOR2_X1 U10085 ( .A(n10265), .B(n10266), .Z(n10059) );
  XNOR2_X1 U10086 ( .A(n10267), .B(n10268), .ZN(n10266) );
  XNOR2_X1 U10087 ( .A(n10269), .B(n10270), .ZN(n10063) );
  XNOR2_X1 U10088 ( .A(n10271), .B(n10272), .ZN(n10269) );
  NOR2_X1 U10089 ( .A1(n8753), .A2(n8743), .ZN(n10272) );
  XOR2_X1 U10090 ( .A(n10273), .B(n10274), .Z(n10066) );
  XOR2_X1 U10091 ( .A(n10275), .B(n10276), .Z(n10273) );
  XNOR2_X1 U10092 ( .A(n10277), .B(n10278), .ZN(n10070) );
  XOR2_X1 U10093 ( .A(n10279), .B(n10280), .Z(n10278) );
  NAND2_X1 U10094 ( .A1(b_25_), .A2(a_16_), .ZN(n10280) );
  XNOR2_X1 U10095 ( .A(n10281), .B(n10282), .ZN(n10075) );
  XNOR2_X1 U10096 ( .A(n10283), .B(n10284), .ZN(n10282) );
  XNOR2_X1 U10097 ( .A(n10285), .B(n10286), .ZN(n10079) );
  XNOR2_X1 U10098 ( .A(n10287), .B(n10288), .ZN(n10285) );
  NOR2_X1 U10099 ( .A1(n8757), .A2(n8743), .ZN(n10288) );
  XNOR2_X1 U10100 ( .A(n10289), .B(n10290), .ZN(n10083) );
  XOR2_X1 U10101 ( .A(n10291), .B(n10292), .Z(n10289) );
  XOR2_X1 U10102 ( .A(n10293), .B(n10294), .Z(n10086) );
  XOR2_X1 U10103 ( .A(n10295), .B(n10296), .Z(n10293) );
  NOR2_X1 U10104 ( .A1(n8759), .A2(n8743), .ZN(n10296) );
  XOR2_X1 U10105 ( .A(n10297), .B(n10298), .Z(n10091) );
  XOR2_X1 U10106 ( .A(n10299), .B(n10300), .Z(n10298) );
  NAND2_X1 U10107 ( .A1(b_25_), .A2(a_11_), .ZN(n10300) );
  XNOR2_X1 U10108 ( .A(n10301), .B(n10302), .ZN(n10095) );
  XNOR2_X1 U10109 ( .A(n10303), .B(n10304), .ZN(n10301) );
  NOR2_X1 U10110 ( .A1(n8761), .A2(n8743), .ZN(n10304) );
  XOR2_X1 U10111 ( .A(n10305), .B(n10306), .Z(n10098) );
  XOR2_X1 U10112 ( .A(n10307), .B(n10308), .Z(n10305) );
  XNOR2_X1 U10113 ( .A(n10309), .B(n10310), .ZN(n10107) );
  XOR2_X1 U10114 ( .A(n10311), .B(n10312), .Z(n10309) );
  NOR2_X1 U10115 ( .A1(n8764), .A2(n8743), .ZN(n10312) );
  XNOR2_X1 U10116 ( .A(n10313), .B(n10314), .ZN(n10110) );
  XOR2_X1 U10117 ( .A(n10315), .B(n10316), .Z(n10314) );
  XNOR2_X1 U10118 ( .A(n10317), .B(n10318), .ZN(n9925) );
  XNOR2_X1 U10119 ( .A(n10319), .B(n10320), .ZN(n10317) );
  NOR2_X1 U10120 ( .A1(n8517), .A2(n8743), .ZN(n10320) );
  XOR2_X1 U10121 ( .A(n10321), .B(n10322), .Z(n9918) );
  XOR2_X1 U10122 ( .A(n10323), .B(n10324), .Z(n10322) );
  NAND2_X1 U10123 ( .A1(b_25_), .A2(a_4_), .ZN(n10324) );
  XNOR2_X1 U10124 ( .A(n10325), .B(n10326), .ZN(n10114) );
  XOR2_X1 U10125 ( .A(n10327), .B(n10328), .Z(n10326) );
  NAND2_X1 U10126 ( .A1(b_25_), .A2(a_3_), .ZN(n10328) );
  XOR2_X1 U10127 ( .A(n10329), .B(n10330), .Z(n10119) );
  XOR2_X1 U10128 ( .A(n10331), .B(n10332), .Z(n10330) );
  NAND2_X1 U10129 ( .A1(b_25_), .A2(a_2_), .ZN(n10332) );
  XNOR2_X1 U10130 ( .A(n10333), .B(n10334), .ZN(n9904) );
  XOR2_X1 U10131 ( .A(n10335), .B(n10336), .Z(n10333) );
  NOR2_X1 U10132 ( .A1(n8617), .A2(n8743), .ZN(n10336) );
  NAND2_X1 U10133 ( .A1(n10337), .A2(n10338), .ZN(n8996) );
  INV_X1 U10134 ( .A(n9901), .ZN(n8997) );
  XOR2_X1 U10135 ( .A(n10339), .B(n10340), .Z(n9901) );
  XNOR2_X1 U10136 ( .A(n10341), .B(n10342), .ZN(n10340) );
  NAND2_X1 U10137 ( .A1(n10343), .A2(n10122), .ZN(n8821) );
  NOR2_X1 U10138 ( .A1(n10338), .A2(n10337), .ZN(n10122) );
  AND2_X1 U10139 ( .A1(n10344), .A2(n10345), .ZN(n10337) );
  NAND2_X1 U10140 ( .A1(n10342), .A2(n10346), .ZN(n10345) );
  OR2_X1 U10141 ( .A1(n10341), .A2(n10339), .ZN(n10346) );
  NOR2_X1 U10142 ( .A1(n8743), .A2(n9674), .ZN(n10342) );
  NAND2_X1 U10143 ( .A1(n10339), .A2(n10341), .ZN(n10344) );
  NAND2_X1 U10144 ( .A1(n10347), .A2(n10348), .ZN(n10341) );
  NAND3_X1 U10145 ( .A1(a_1_), .A2(n10349), .A3(b_25_), .ZN(n10348) );
  OR2_X1 U10146 ( .A1(n10335), .A2(n10334), .ZN(n10349) );
  NAND2_X1 U10147 ( .A1(n10334), .A2(n10335), .ZN(n10347) );
  NAND2_X1 U10148 ( .A1(n10350), .A2(n10351), .ZN(n10335) );
  NAND3_X1 U10149 ( .A1(a_2_), .A2(n10352), .A3(b_25_), .ZN(n10351) );
  OR2_X1 U10150 ( .A1(n10331), .A2(n10329), .ZN(n10352) );
  NAND2_X1 U10151 ( .A1(n10329), .A2(n10331), .ZN(n10350) );
  NAND2_X1 U10152 ( .A1(n10353), .A2(n10354), .ZN(n10331) );
  NAND3_X1 U10153 ( .A1(a_3_), .A2(n10355), .A3(b_25_), .ZN(n10354) );
  OR2_X1 U10154 ( .A1(n10327), .A2(n10325), .ZN(n10355) );
  NAND2_X1 U10155 ( .A1(n10325), .A2(n10327), .ZN(n10353) );
  NAND2_X1 U10156 ( .A1(n10356), .A2(n10357), .ZN(n10327) );
  NAND3_X1 U10157 ( .A1(a_4_), .A2(n10358), .A3(b_25_), .ZN(n10357) );
  OR2_X1 U10158 ( .A1(n10323), .A2(n10321), .ZN(n10358) );
  NAND2_X1 U10159 ( .A1(n10321), .A2(n10323), .ZN(n10356) );
  NAND2_X1 U10160 ( .A1(n10359), .A2(n10360), .ZN(n10323) );
  NAND3_X1 U10161 ( .A1(a_5_), .A2(n10361), .A3(b_25_), .ZN(n10360) );
  NAND2_X1 U10162 ( .A1(n10319), .A2(n10318), .ZN(n10361) );
  OR2_X1 U10163 ( .A1(n10318), .A2(n10319), .ZN(n10359) );
  AND2_X1 U10164 ( .A1(n10362), .A2(n10363), .ZN(n10319) );
  NAND2_X1 U10165 ( .A1(n10315), .A2(n10364), .ZN(n10363) );
  NAND2_X1 U10166 ( .A1(n10365), .A2(n10316), .ZN(n10364) );
  INV_X1 U10167 ( .A(n10313), .ZN(n10365) );
  NAND2_X1 U10168 ( .A1(n10366), .A2(n10367), .ZN(n10315) );
  NAND3_X1 U10169 ( .A1(a_7_), .A2(n10368), .A3(b_25_), .ZN(n10367) );
  OR2_X1 U10170 ( .A1(n10311), .A2(n10310), .ZN(n10368) );
  NAND2_X1 U10171 ( .A1(n10310), .A2(n10311), .ZN(n10366) );
  NAND2_X1 U10172 ( .A1(n10369), .A2(n10370), .ZN(n10311) );
  NAND3_X1 U10173 ( .A1(a_8_), .A2(n10371), .A3(b_25_), .ZN(n10370) );
  OR2_X1 U10174 ( .A1(n10150), .A2(n10149), .ZN(n10371) );
  NAND2_X1 U10175 ( .A1(n10149), .A2(n10150), .ZN(n10369) );
  NAND2_X1 U10176 ( .A1(n10372), .A2(n10373), .ZN(n10150) );
  NAND2_X1 U10177 ( .A1(n10308), .A2(n10374), .ZN(n10373) );
  OR2_X1 U10178 ( .A1(n10307), .A2(n10306), .ZN(n10374) );
  NOR2_X1 U10179 ( .A1(n8743), .A2(n8426), .ZN(n10308) );
  NAND2_X1 U10180 ( .A1(n10306), .A2(n10307), .ZN(n10372) );
  NAND2_X1 U10181 ( .A1(n10375), .A2(n10376), .ZN(n10307) );
  NAND3_X1 U10182 ( .A1(a_10_), .A2(n10377), .A3(b_25_), .ZN(n10376) );
  NAND2_X1 U10183 ( .A1(n10303), .A2(n10302), .ZN(n10377) );
  OR2_X1 U10184 ( .A1(n10302), .A2(n10303), .ZN(n10375) );
  AND2_X1 U10185 ( .A1(n10378), .A2(n10379), .ZN(n10303) );
  NAND3_X1 U10186 ( .A1(a_11_), .A2(n10380), .A3(b_25_), .ZN(n10379) );
  OR2_X1 U10187 ( .A1(n10299), .A2(n10297), .ZN(n10380) );
  NAND2_X1 U10188 ( .A1(n10297), .A2(n10299), .ZN(n10378) );
  NAND2_X1 U10189 ( .A1(n10381), .A2(n10382), .ZN(n10299) );
  NAND3_X1 U10190 ( .A1(a_12_), .A2(n10383), .A3(b_25_), .ZN(n10382) );
  OR2_X1 U10191 ( .A1(n10295), .A2(n10294), .ZN(n10383) );
  NAND2_X1 U10192 ( .A1(n10294), .A2(n10295), .ZN(n10381) );
  NAND2_X1 U10193 ( .A1(n10384), .A2(n10385), .ZN(n10295) );
  NAND2_X1 U10194 ( .A1(n10292), .A2(n10386), .ZN(n10385) );
  OR2_X1 U10195 ( .A1(n10291), .A2(n10290), .ZN(n10386) );
  NOR2_X1 U10196 ( .A1(n8743), .A2(n8310), .ZN(n10292) );
  NAND2_X1 U10197 ( .A1(n10290), .A2(n10291), .ZN(n10384) );
  NAND2_X1 U10198 ( .A1(n10387), .A2(n10388), .ZN(n10291) );
  NAND3_X1 U10199 ( .A1(a_14_), .A2(n10389), .A3(b_25_), .ZN(n10388) );
  NAND2_X1 U10200 ( .A1(n10287), .A2(n10286), .ZN(n10389) );
  OR2_X1 U10201 ( .A1(n10286), .A2(n10287), .ZN(n10387) );
  AND2_X1 U10202 ( .A1(n10390), .A2(n10391), .ZN(n10287) );
  NAND2_X1 U10203 ( .A1(n10284), .A2(n10392), .ZN(n10391) );
  OR2_X1 U10204 ( .A1(n10283), .A2(n10281), .ZN(n10392) );
  NOR2_X1 U10205 ( .A1(n8743), .A2(n8276), .ZN(n10284) );
  NAND2_X1 U10206 ( .A1(n10281), .A2(n10283), .ZN(n10390) );
  NAND2_X1 U10207 ( .A1(n10393), .A2(n10394), .ZN(n10283) );
  NAND3_X1 U10208 ( .A1(a_16_), .A2(n10395), .A3(b_25_), .ZN(n10394) );
  OR2_X1 U10209 ( .A1(n10279), .A2(n10277), .ZN(n10395) );
  NAND2_X1 U10210 ( .A1(n10277), .A2(n10279), .ZN(n10393) );
  NAND2_X1 U10211 ( .A1(n10396), .A2(n10397), .ZN(n10279) );
  NAND2_X1 U10212 ( .A1(n10276), .A2(n10398), .ZN(n10397) );
  OR2_X1 U10213 ( .A1(n10275), .A2(n10274), .ZN(n10398) );
  NOR2_X1 U10214 ( .A1(n8743), .A2(n8210), .ZN(n10276) );
  NAND2_X1 U10215 ( .A1(n10274), .A2(n10275), .ZN(n10396) );
  NAND2_X1 U10216 ( .A1(n10399), .A2(n10400), .ZN(n10275) );
  NAND3_X1 U10217 ( .A1(a_18_), .A2(n10401), .A3(b_25_), .ZN(n10400) );
  NAND2_X1 U10218 ( .A1(n10271), .A2(n10270), .ZN(n10401) );
  OR2_X1 U10219 ( .A1(n10270), .A2(n10271), .ZN(n10399) );
  AND2_X1 U10220 ( .A1(n10402), .A2(n10403), .ZN(n10271) );
  NAND2_X1 U10221 ( .A1(n10268), .A2(n10404), .ZN(n10403) );
  OR2_X1 U10222 ( .A1(n10267), .A2(n10265), .ZN(n10404) );
  NOR2_X1 U10223 ( .A1(n8743), .A2(n8170), .ZN(n10268) );
  NAND2_X1 U10224 ( .A1(n10265), .A2(n10267), .ZN(n10402) );
  NAND2_X1 U10225 ( .A1(n10405), .A2(n10406), .ZN(n10267) );
  NAND3_X1 U10226 ( .A1(a_20_), .A2(n10407), .A3(b_25_), .ZN(n10406) );
  NAND2_X1 U10227 ( .A1(n10263), .A2(n10262), .ZN(n10407) );
  OR2_X1 U10228 ( .A1(n10262), .A2(n10263), .ZN(n10405) );
  AND2_X1 U10229 ( .A1(n10408), .A2(n10409), .ZN(n10263) );
  NAND2_X1 U10230 ( .A1(n10260), .A2(n10410), .ZN(n10409) );
  OR2_X1 U10231 ( .A1(n10259), .A2(n10258), .ZN(n10410) );
  NOR2_X1 U10232 ( .A1(n8743), .A2(n8750), .ZN(n10260) );
  NAND2_X1 U10233 ( .A1(n10258), .A2(n10259), .ZN(n10408) );
  NAND2_X1 U10234 ( .A1(n10411), .A2(n10412), .ZN(n10259) );
  NAND3_X1 U10235 ( .A1(a_22_), .A2(n10413), .A3(b_25_), .ZN(n10412) );
  OR2_X1 U10236 ( .A1(n10255), .A2(n10253), .ZN(n10413) );
  NAND2_X1 U10237 ( .A1(n10253), .A2(n10255), .ZN(n10411) );
  NAND2_X1 U10238 ( .A1(n10414), .A2(n10415), .ZN(n10255) );
  NAND2_X1 U10239 ( .A1(n10252), .A2(n10416), .ZN(n10415) );
  OR2_X1 U10240 ( .A1(n10251), .A2(n10249), .ZN(n10416) );
  NOR2_X1 U10241 ( .A1(n8743), .A2(n8747), .ZN(n10252) );
  NAND2_X1 U10242 ( .A1(n10249), .A2(n10251), .ZN(n10414) );
  NAND2_X1 U10243 ( .A1(n10417), .A2(n10418), .ZN(n10251) );
  NAND3_X1 U10244 ( .A1(a_24_), .A2(n10419), .A3(b_25_), .ZN(n10418) );
  NAND2_X1 U10245 ( .A1(n10247), .A2(n10246), .ZN(n10419) );
  OR2_X1 U10246 ( .A1(n10246), .A2(n10247), .ZN(n10417) );
  AND2_X1 U10247 ( .A1(n10420), .A2(n10421), .ZN(n10247) );
  NAND2_X1 U10248 ( .A1(n10244), .A2(n10422), .ZN(n10421) );
  OR2_X1 U10249 ( .A1(n10243), .A2(n10242), .ZN(n10422) );
  INV_X1 U10250 ( .A(n8017), .ZN(n10244) );
  NAND2_X1 U10251 ( .A1(b_25_), .A2(a_25_), .ZN(n8017) );
  NAND2_X1 U10252 ( .A1(n10242), .A2(n10243), .ZN(n10420) );
  NAND2_X1 U10253 ( .A1(n10239), .A2(n10423), .ZN(n10243) );
  NAND2_X1 U10254 ( .A1(n10238), .A2(n10240), .ZN(n10423) );
  NAND2_X1 U10255 ( .A1(n10424), .A2(n10425), .ZN(n10240) );
  NAND2_X1 U10256 ( .A1(b_25_), .A2(a_26_), .ZN(n10425) );
  INV_X1 U10257 ( .A(n10426), .ZN(n10424) );
  XNOR2_X1 U10258 ( .A(n10427), .B(n10428), .ZN(n10238) );
  NAND2_X1 U10259 ( .A1(n10429), .A2(n10430), .ZN(n10427) );
  NAND2_X1 U10260 ( .A1(a_26_), .A2(n10426), .ZN(n10239) );
  NAND2_X1 U10261 ( .A1(n10211), .A2(n10431), .ZN(n10426) );
  NAND2_X1 U10262 ( .A1(n10210), .A2(n10212), .ZN(n10431) );
  NAND2_X1 U10263 ( .A1(n10432), .A2(n10433), .ZN(n10212) );
  NAND2_X1 U10264 ( .A1(b_25_), .A2(a_27_), .ZN(n10433) );
  INV_X1 U10265 ( .A(n10434), .ZN(n10432) );
  XNOR2_X1 U10266 ( .A(n10435), .B(n10436), .ZN(n10210) );
  XOR2_X1 U10267 ( .A(n10437), .B(n10438), .Z(n10435) );
  NAND2_X1 U10268 ( .A1(b_24_), .A2(a_28_), .ZN(n10437) );
  NAND2_X1 U10269 ( .A1(a_27_), .A2(n10434), .ZN(n10211) );
  NAND2_X1 U10270 ( .A1(n10439), .A2(n10440), .ZN(n10434) );
  NAND3_X1 U10271 ( .A1(a_28_), .A2(n10441), .A3(b_25_), .ZN(n10440) );
  NAND2_X1 U10272 ( .A1(n10220), .A2(n10218), .ZN(n10441) );
  OR2_X1 U10273 ( .A1(n10218), .A2(n10220), .ZN(n10439) );
  AND2_X1 U10274 ( .A1(n10442), .A2(n10443), .ZN(n10220) );
  NAND2_X1 U10275 ( .A1(n10234), .A2(n10444), .ZN(n10443) );
  OR2_X1 U10276 ( .A1(n10235), .A2(n10236), .ZN(n10444) );
  NOR2_X1 U10277 ( .A1(n8743), .A2(n7890), .ZN(n10234) );
  NAND2_X1 U10278 ( .A1(n10236), .A2(n10235), .ZN(n10442) );
  NAND2_X1 U10279 ( .A1(n10445), .A2(n10446), .ZN(n10235) );
  NAND2_X1 U10280 ( .A1(b_23_), .A2(n10447), .ZN(n10446) );
  NAND2_X1 U10281 ( .A1(n7864), .A2(n10448), .ZN(n10447) );
  NAND2_X1 U10282 ( .A1(a_31_), .A2(n8043), .ZN(n10448) );
  NAND2_X1 U10283 ( .A1(b_24_), .A2(n10449), .ZN(n10445) );
  NAND2_X1 U10284 ( .A1(n9137), .A2(n10450), .ZN(n10449) );
  NAND2_X1 U10285 ( .A1(a_30_), .A2(n8746), .ZN(n10450) );
  AND3_X1 U10286 ( .A1(b_24_), .A2(b_25_), .A3(n7818), .ZN(n10236) );
  XNOR2_X1 U10287 ( .A(n10451), .B(n10452), .ZN(n10218) );
  XOR2_X1 U10288 ( .A(n10453), .B(n10454), .Z(n10451) );
  XNOR2_X1 U10289 ( .A(n10455), .B(n10456), .ZN(n10242) );
  NAND2_X1 U10290 ( .A1(n10457), .A2(n10458), .ZN(n10455) );
  XNOR2_X1 U10291 ( .A(n10459), .B(n10460), .ZN(n10246) );
  XOR2_X1 U10292 ( .A(n10461), .B(n10462), .Z(n10459) );
  XOR2_X1 U10293 ( .A(n10463), .B(n10464), .Z(n10249) );
  XOR2_X1 U10294 ( .A(n10465), .B(n10466), .Z(n10463) );
  XOR2_X1 U10295 ( .A(n10467), .B(n10468), .Z(n10253) );
  XOR2_X1 U10296 ( .A(n10469), .B(n10470), .Z(n10467) );
  XNOR2_X1 U10297 ( .A(n10471), .B(n10472), .ZN(n10258) );
  XOR2_X1 U10298 ( .A(n10473), .B(n10474), .Z(n10472) );
  NAND2_X1 U10299 ( .A1(b_24_), .A2(a_22_), .ZN(n10474) );
  XNOR2_X1 U10300 ( .A(n10475), .B(n10476), .ZN(n10262) );
  XOR2_X1 U10301 ( .A(n10477), .B(n10478), .Z(n10475) );
  XNOR2_X1 U10302 ( .A(n10479), .B(n10480), .ZN(n10265) );
  XNOR2_X1 U10303 ( .A(n10481), .B(n10482), .ZN(n10479) );
  NOR2_X1 U10304 ( .A1(n8751), .A2(n8043), .ZN(n10482) );
  XOR2_X1 U10305 ( .A(n10483), .B(n10484), .Z(n10270) );
  XNOR2_X1 U10306 ( .A(n10485), .B(n10486), .ZN(n10484) );
  XNOR2_X1 U10307 ( .A(n10487), .B(n10488), .ZN(n10274) );
  XNOR2_X1 U10308 ( .A(n10489), .B(n10490), .ZN(n10487) );
  NOR2_X1 U10309 ( .A1(n8753), .A2(n8043), .ZN(n10490) );
  XOR2_X1 U10310 ( .A(n10491), .B(n10492), .Z(n10277) );
  XOR2_X1 U10311 ( .A(n10493), .B(n10494), .Z(n10491) );
  XOR2_X1 U10312 ( .A(n10495), .B(n10496), .Z(n10281) );
  XOR2_X1 U10313 ( .A(n10497), .B(n10498), .Z(n10495) );
  NOR2_X1 U10314 ( .A1(n8755), .A2(n8043), .ZN(n10498) );
  XOR2_X1 U10315 ( .A(n10499), .B(n10500), .Z(n10286) );
  XNOR2_X1 U10316 ( .A(n10501), .B(n10502), .ZN(n10500) );
  XNOR2_X1 U10317 ( .A(n10503), .B(n10504), .ZN(n10290) );
  XOR2_X1 U10318 ( .A(n10505), .B(n10506), .Z(n10503) );
  NAND2_X1 U10319 ( .A1(b_24_), .A2(a_14_), .ZN(n10505) );
  XNOR2_X1 U10320 ( .A(n10507), .B(n10508), .ZN(n10294) );
  XNOR2_X1 U10321 ( .A(n10509), .B(n10510), .ZN(n10507) );
  XNOR2_X1 U10322 ( .A(n10511), .B(n10512), .ZN(n10297) );
  XOR2_X1 U10323 ( .A(n10513), .B(n10514), .Z(n10512) );
  NAND2_X1 U10324 ( .A1(b_24_), .A2(a_12_), .ZN(n10514) );
  XOR2_X1 U10325 ( .A(n10515), .B(n10516), .Z(n10302) );
  XOR2_X1 U10326 ( .A(n10517), .B(n10518), .Z(n10516) );
  NAND2_X1 U10327 ( .A1(b_24_), .A2(a_11_), .ZN(n10518) );
  XNOR2_X1 U10328 ( .A(n10519), .B(n10520), .ZN(n10306) );
  XOR2_X1 U10329 ( .A(n10521), .B(n10522), .Z(n10520) );
  NAND2_X1 U10330 ( .A1(b_24_), .A2(a_10_), .ZN(n10522) );
  XNOR2_X1 U10331 ( .A(n10523), .B(n10524), .ZN(n10149) );
  XNOR2_X1 U10332 ( .A(n10525), .B(n10526), .ZN(n10524) );
  XNOR2_X1 U10333 ( .A(n10527), .B(n10528), .ZN(n10310) );
  XOR2_X1 U10334 ( .A(n10529), .B(n10530), .Z(n10527) );
  NAND2_X1 U10335 ( .A1(b_24_), .A2(a_8_), .ZN(n10529) );
  NAND2_X1 U10336 ( .A1(n10531), .A2(n10313), .ZN(n10362) );
  XNOR2_X1 U10337 ( .A(n10532), .B(n10533), .ZN(n10313) );
  NAND2_X1 U10338 ( .A1(n10534), .A2(n10535), .ZN(n10532) );
  INV_X1 U10339 ( .A(n10316), .ZN(n10531) );
  NAND2_X1 U10340 ( .A1(b_25_), .A2(a_6_), .ZN(n10316) );
  XNOR2_X1 U10341 ( .A(n10536), .B(n10537), .ZN(n10318) );
  XOR2_X1 U10342 ( .A(n10538), .B(n10539), .Z(n10536) );
  XNOR2_X1 U10343 ( .A(n10540), .B(n10541), .ZN(n10321) );
  XNOR2_X1 U10344 ( .A(n10542), .B(n10543), .ZN(n10540) );
  XNOR2_X1 U10345 ( .A(n10544), .B(n10545), .ZN(n10325) );
  XNOR2_X1 U10346 ( .A(n10546), .B(n10547), .ZN(n10544) );
  NOR2_X1 U10347 ( .A1(n8766), .A2(n8043), .ZN(n10547) );
  XNOR2_X1 U10348 ( .A(n10548), .B(n10549), .ZN(n10329) );
  NAND2_X1 U10349 ( .A1(n10550), .A2(n10551), .ZN(n10548) );
  XNOR2_X1 U10350 ( .A(n10552), .B(n10553), .ZN(n10334) );
  NAND2_X1 U10351 ( .A1(n10554), .A2(n10555), .ZN(n10552) );
  XOR2_X1 U10352 ( .A(n10556), .B(n10557), .Z(n10339) );
  XOR2_X1 U10353 ( .A(n10558), .B(n10559), .Z(n10557) );
  XNOR2_X1 U10354 ( .A(n10560), .B(n10561), .ZN(n10338) );
  XOR2_X1 U10355 ( .A(n10562), .B(n10563), .Z(n10560) );
  NOR2_X1 U10356 ( .A1(n9674), .A2(n8043), .ZN(n10563) );
  XOR2_X1 U10357 ( .A(n8988), .B(n8987), .Z(n10343) );
  NAND3_X1 U10358 ( .A1(n8987), .A2(n8988), .A3(n10564), .ZN(n8828) );
  XOR2_X1 U10359 ( .A(n8983), .B(n8982), .Z(n10564) );
  NAND2_X1 U10360 ( .A1(n10565), .A2(n10566), .ZN(n8988) );
  NAND3_X1 U10361 ( .A1(a_0_), .A2(n10567), .A3(b_24_), .ZN(n10566) );
  OR2_X1 U10362 ( .A1(n10562), .A2(n10561), .ZN(n10567) );
  NAND2_X1 U10363 ( .A1(n10561), .A2(n10562), .ZN(n10565) );
  NAND2_X1 U10364 ( .A1(n10568), .A2(n10569), .ZN(n10562) );
  NAND2_X1 U10365 ( .A1(n10558), .A2(n10570), .ZN(n10569) );
  NAND2_X1 U10366 ( .A1(n10556), .A2(n10559), .ZN(n10570) );
  NAND2_X1 U10367 ( .A1(n10554), .A2(n10571), .ZN(n10558) );
  NAND2_X1 U10368 ( .A1(n10553), .A2(n10555), .ZN(n10571) );
  NAND2_X1 U10369 ( .A1(n10572), .A2(n10573), .ZN(n10555) );
  NAND2_X1 U10370 ( .A1(b_24_), .A2(a_2_), .ZN(n10573) );
  INV_X1 U10371 ( .A(n10574), .ZN(n10572) );
  XNOR2_X1 U10372 ( .A(n10575), .B(n10576), .ZN(n10553) );
  XOR2_X1 U10373 ( .A(n10577), .B(n10578), .Z(n10576) );
  NAND2_X1 U10374 ( .A1(b_23_), .A2(a_3_), .ZN(n10578) );
  NAND2_X1 U10375 ( .A1(a_2_), .A2(n10574), .ZN(n10554) );
  NAND2_X1 U10376 ( .A1(n10550), .A2(n10579), .ZN(n10574) );
  NAND2_X1 U10377 ( .A1(n10549), .A2(n10551), .ZN(n10579) );
  NAND2_X1 U10378 ( .A1(n10580), .A2(n10581), .ZN(n10551) );
  NAND2_X1 U10379 ( .A1(b_24_), .A2(a_3_), .ZN(n10581) );
  INV_X1 U10380 ( .A(n10582), .ZN(n10580) );
  XNOR2_X1 U10381 ( .A(n10583), .B(n10584), .ZN(n10549) );
  XOR2_X1 U10382 ( .A(n10585), .B(n10586), .Z(n10584) );
  NAND2_X1 U10383 ( .A1(b_23_), .A2(a_4_), .ZN(n10586) );
  NAND2_X1 U10384 ( .A1(a_3_), .A2(n10582), .ZN(n10550) );
  NAND2_X1 U10385 ( .A1(n10587), .A2(n10588), .ZN(n10582) );
  NAND3_X1 U10386 ( .A1(a_4_), .A2(n10589), .A3(b_24_), .ZN(n10588) );
  NAND2_X1 U10387 ( .A1(n10546), .A2(n10545), .ZN(n10589) );
  OR2_X1 U10388 ( .A1(n10545), .A2(n10546), .ZN(n10587) );
  AND2_X1 U10389 ( .A1(n10590), .A2(n10591), .ZN(n10546) );
  NAND2_X1 U10390 ( .A1(n10543), .A2(n10592), .ZN(n10591) );
  NAND2_X1 U10391 ( .A1(n10542), .A2(n10541), .ZN(n10592) );
  NOR2_X1 U10392 ( .A1(n8043), .A2(n8517), .ZN(n10543) );
  OR2_X1 U10393 ( .A1(n10541), .A2(n10542), .ZN(n10590) );
  AND2_X1 U10394 ( .A1(n10593), .A2(n10594), .ZN(n10542) );
  NAND2_X1 U10395 ( .A1(n10539), .A2(n10595), .ZN(n10594) );
  OR2_X1 U10396 ( .A1(n10537), .A2(n10538), .ZN(n10595) );
  NAND2_X1 U10397 ( .A1(n10534), .A2(n10596), .ZN(n10539) );
  NAND2_X1 U10398 ( .A1(n10533), .A2(n10535), .ZN(n10596) );
  NAND2_X1 U10399 ( .A1(n10597), .A2(n10598), .ZN(n10535) );
  NAND2_X1 U10400 ( .A1(b_24_), .A2(a_7_), .ZN(n10598) );
  INV_X1 U10401 ( .A(n10599), .ZN(n10597) );
  XNOR2_X1 U10402 ( .A(n10600), .B(n10601), .ZN(n10533) );
  XNOR2_X1 U10403 ( .A(n10602), .B(n10603), .ZN(n10601) );
  NAND2_X1 U10404 ( .A1(a_7_), .A2(n10599), .ZN(n10534) );
  NAND2_X1 U10405 ( .A1(n10604), .A2(n10605), .ZN(n10599) );
  NAND3_X1 U10406 ( .A1(a_8_), .A2(n10606), .A3(b_24_), .ZN(n10605) );
  NAND2_X1 U10407 ( .A1(n10530), .A2(n10528), .ZN(n10606) );
  OR2_X1 U10408 ( .A1(n10528), .A2(n10530), .ZN(n10604) );
  AND2_X1 U10409 ( .A1(n10607), .A2(n10608), .ZN(n10530) );
  NAND2_X1 U10410 ( .A1(n10526), .A2(n10609), .ZN(n10608) );
  OR2_X1 U10411 ( .A1(n10525), .A2(n10523), .ZN(n10609) );
  NOR2_X1 U10412 ( .A1(n8043), .A2(n8426), .ZN(n10526) );
  NAND2_X1 U10413 ( .A1(n10523), .A2(n10525), .ZN(n10607) );
  NAND2_X1 U10414 ( .A1(n10610), .A2(n10611), .ZN(n10525) );
  NAND3_X1 U10415 ( .A1(a_10_), .A2(n10612), .A3(b_24_), .ZN(n10611) );
  OR2_X1 U10416 ( .A1(n10521), .A2(n10519), .ZN(n10612) );
  NAND2_X1 U10417 ( .A1(n10519), .A2(n10521), .ZN(n10610) );
  NAND2_X1 U10418 ( .A1(n10613), .A2(n10614), .ZN(n10521) );
  NAND3_X1 U10419 ( .A1(a_11_), .A2(n10615), .A3(b_24_), .ZN(n10614) );
  OR2_X1 U10420 ( .A1(n10517), .A2(n10515), .ZN(n10615) );
  NAND2_X1 U10421 ( .A1(n10515), .A2(n10517), .ZN(n10613) );
  NAND2_X1 U10422 ( .A1(n10616), .A2(n10617), .ZN(n10517) );
  NAND3_X1 U10423 ( .A1(a_12_), .A2(n10618), .A3(b_24_), .ZN(n10617) );
  OR2_X1 U10424 ( .A1(n10513), .A2(n10511), .ZN(n10618) );
  NAND2_X1 U10425 ( .A1(n10511), .A2(n10513), .ZN(n10616) );
  NAND2_X1 U10426 ( .A1(n10619), .A2(n10620), .ZN(n10513) );
  NAND2_X1 U10427 ( .A1(n10510), .A2(n10621), .ZN(n10620) );
  NAND2_X1 U10428 ( .A1(n10509), .A2(n10508), .ZN(n10621) );
  NOR2_X1 U10429 ( .A1(n8043), .A2(n8310), .ZN(n10510) );
  OR2_X1 U10430 ( .A1(n10508), .A2(n10509), .ZN(n10619) );
  AND2_X1 U10431 ( .A1(n10622), .A2(n10623), .ZN(n10509) );
  NAND3_X1 U10432 ( .A1(a_14_), .A2(n10624), .A3(b_24_), .ZN(n10623) );
  NAND2_X1 U10433 ( .A1(n10506), .A2(n10504), .ZN(n10624) );
  OR2_X1 U10434 ( .A1(n10504), .A2(n10506), .ZN(n10622) );
  AND2_X1 U10435 ( .A1(n10625), .A2(n10626), .ZN(n10506) );
  NAND2_X1 U10436 ( .A1(n10502), .A2(n10627), .ZN(n10626) );
  OR2_X1 U10437 ( .A1(n10501), .A2(n10499), .ZN(n10627) );
  NOR2_X1 U10438 ( .A1(n8043), .A2(n8276), .ZN(n10502) );
  NAND2_X1 U10439 ( .A1(n10499), .A2(n10501), .ZN(n10625) );
  NAND2_X1 U10440 ( .A1(n10628), .A2(n10629), .ZN(n10501) );
  NAND3_X1 U10441 ( .A1(a_16_), .A2(n10630), .A3(b_24_), .ZN(n10629) );
  OR2_X1 U10442 ( .A1(n10497), .A2(n10496), .ZN(n10630) );
  NAND2_X1 U10443 ( .A1(n10496), .A2(n10497), .ZN(n10628) );
  NAND2_X1 U10444 ( .A1(n10631), .A2(n10632), .ZN(n10497) );
  NAND2_X1 U10445 ( .A1(n10494), .A2(n10633), .ZN(n10632) );
  OR2_X1 U10446 ( .A1(n10493), .A2(n10492), .ZN(n10633) );
  NOR2_X1 U10447 ( .A1(n8043), .A2(n8210), .ZN(n10494) );
  NAND2_X1 U10448 ( .A1(n10492), .A2(n10493), .ZN(n10631) );
  NAND2_X1 U10449 ( .A1(n10634), .A2(n10635), .ZN(n10493) );
  NAND3_X1 U10450 ( .A1(a_18_), .A2(n10636), .A3(b_24_), .ZN(n10635) );
  NAND2_X1 U10451 ( .A1(n10489), .A2(n10488), .ZN(n10636) );
  OR2_X1 U10452 ( .A1(n10488), .A2(n10489), .ZN(n10634) );
  AND2_X1 U10453 ( .A1(n10637), .A2(n10638), .ZN(n10489) );
  NAND2_X1 U10454 ( .A1(n10486), .A2(n10639), .ZN(n10638) );
  OR2_X1 U10455 ( .A1(n10485), .A2(n10483), .ZN(n10639) );
  NOR2_X1 U10456 ( .A1(n8043), .A2(n8170), .ZN(n10486) );
  NAND2_X1 U10457 ( .A1(n10483), .A2(n10485), .ZN(n10637) );
  NAND2_X1 U10458 ( .A1(n10640), .A2(n10641), .ZN(n10485) );
  NAND3_X1 U10459 ( .A1(a_20_), .A2(n10642), .A3(b_24_), .ZN(n10641) );
  NAND2_X1 U10460 ( .A1(n10481), .A2(n10480), .ZN(n10642) );
  OR2_X1 U10461 ( .A1(n10480), .A2(n10481), .ZN(n10640) );
  AND2_X1 U10462 ( .A1(n10643), .A2(n10644), .ZN(n10481) );
  NAND2_X1 U10463 ( .A1(n10478), .A2(n10645), .ZN(n10644) );
  OR2_X1 U10464 ( .A1(n10477), .A2(n10476), .ZN(n10645) );
  NOR2_X1 U10465 ( .A1(n8043), .A2(n8750), .ZN(n10478) );
  NAND2_X1 U10466 ( .A1(n10476), .A2(n10477), .ZN(n10643) );
  NAND2_X1 U10467 ( .A1(n10646), .A2(n10647), .ZN(n10477) );
  NAND3_X1 U10468 ( .A1(a_22_), .A2(n10648), .A3(b_24_), .ZN(n10647) );
  OR2_X1 U10469 ( .A1(n10473), .A2(n10471), .ZN(n10648) );
  NAND2_X1 U10470 ( .A1(n10471), .A2(n10473), .ZN(n10646) );
  NAND2_X1 U10471 ( .A1(n10649), .A2(n10650), .ZN(n10473) );
  NAND2_X1 U10472 ( .A1(n10470), .A2(n10651), .ZN(n10650) );
  OR2_X1 U10473 ( .A1(n10469), .A2(n10468), .ZN(n10651) );
  NOR2_X1 U10474 ( .A1(n8043), .A2(n8747), .ZN(n10470) );
  NAND2_X1 U10475 ( .A1(n10468), .A2(n10469), .ZN(n10649) );
  NAND2_X1 U10476 ( .A1(n10652), .A2(n10653), .ZN(n10469) );
  NAND2_X1 U10477 ( .A1(n10464), .A2(n10654), .ZN(n10653) );
  OR2_X1 U10478 ( .A1(n10465), .A2(n10466), .ZN(n10654) );
  XOR2_X1 U10479 ( .A(n10655), .B(n10656), .Z(n10464) );
  XOR2_X1 U10480 ( .A(n10657), .B(n10658), .Z(n10655) );
  NAND2_X1 U10481 ( .A1(n10466), .A2(n10465), .ZN(n10652) );
  NAND2_X1 U10482 ( .A1(n10659), .A2(n10660), .ZN(n10465) );
  NAND2_X1 U10483 ( .A1(n10462), .A2(n10661), .ZN(n10660) );
  OR2_X1 U10484 ( .A1(n10461), .A2(n10460), .ZN(n10661) );
  NOR2_X1 U10485 ( .A1(n8043), .A2(n8744), .ZN(n10462) );
  NAND2_X1 U10486 ( .A1(n10460), .A2(n10461), .ZN(n10659) );
  NAND2_X1 U10487 ( .A1(n10457), .A2(n10662), .ZN(n10461) );
  NAND2_X1 U10488 ( .A1(n10456), .A2(n10458), .ZN(n10662) );
  NAND2_X1 U10489 ( .A1(n10663), .A2(n10664), .ZN(n10458) );
  NAND2_X1 U10490 ( .A1(b_24_), .A2(a_26_), .ZN(n10664) );
  INV_X1 U10491 ( .A(n10665), .ZN(n10663) );
  XNOR2_X1 U10492 ( .A(n10666), .B(n10667), .ZN(n10456) );
  NAND2_X1 U10493 ( .A1(n10668), .A2(n10669), .ZN(n10666) );
  NAND2_X1 U10494 ( .A1(a_26_), .A2(n10665), .ZN(n10457) );
  NAND2_X1 U10495 ( .A1(n10429), .A2(n10670), .ZN(n10665) );
  NAND2_X1 U10496 ( .A1(n10428), .A2(n10430), .ZN(n10670) );
  NAND2_X1 U10497 ( .A1(n10671), .A2(n10672), .ZN(n10430) );
  NAND2_X1 U10498 ( .A1(b_24_), .A2(a_27_), .ZN(n10672) );
  INV_X1 U10499 ( .A(n10673), .ZN(n10671) );
  XNOR2_X1 U10500 ( .A(n10674), .B(n10675), .ZN(n10428) );
  XOR2_X1 U10501 ( .A(n10676), .B(n10677), .Z(n10674) );
  NAND2_X1 U10502 ( .A1(b_23_), .A2(a_28_), .ZN(n10676) );
  NAND2_X1 U10503 ( .A1(a_27_), .A2(n10673), .ZN(n10429) );
  NAND2_X1 U10504 ( .A1(n10678), .A2(n10679), .ZN(n10673) );
  NAND3_X1 U10505 ( .A1(a_28_), .A2(n10680), .A3(b_24_), .ZN(n10679) );
  NAND2_X1 U10506 ( .A1(n10438), .A2(n10436), .ZN(n10680) );
  OR2_X1 U10507 ( .A1(n10436), .A2(n10438), .ZN(n10678) );
  AND2_X1 U10508 ( .A1(n10681), .A2(n10682), .ZN(n10438) );
  NAND2_X1 U10509 ( .A1(n10452), .A2(n10683), .ZN(n10682) );
  OR2_X1 U10510 ( .A1(n10453), .A2(n10454), .ZN(n10683) );
  NOR2_X1 U10511 ( .A1(n8043), .A2(n7890), .ZN(n10452) );
  NAND2_X1 U10512 ( .A1(n10454), .A2(n10453), .ZN(n10681) );
  NAND2_X1 U10513 ( .A1(n10684), .A2(n10685), .ZN(n10453) );
  NAND2_X1 U10514 ( .A1(b_22_), .A2(n10686), .ZN(n10685) );
  NAND2_X1 U10515 ( .A1(n7864), .A2(n10687), .ZN(n10686) );
  NAND2_X1 U10516 ( .A1(a_31_), .A2(n8746), .ZN(n10687) );
  NAND2_X1 U10517 ( .A1(b_23_), .A2(n10688), .ZN(n10684) );
  NAND2_X1 U10518 ( .A1(n9137), .A2(n10689), .ZN(n10688) );
  NAND2_X1 U10519 ( .A1(a_30_), .A2(n8094), .ZN(n10689) );
  AND3_X1 U10520 ( .A1(b_23_), .A2(b_24_), .A3(n7818), .ZN(n10454) );
  XNOR2_X1 U10521 ( .A(n10690), .B(n10691), .ZN(n10436) );
  XOR2_X1 U10522 ( .A(n10692), .B(n10693), .Z(n10690) );
  XNOR2_X1 U10523 ( .A(n10694), .B(n10695), .ZN(n10460) );
  NAND2_X1 U10524 ( .A1(n10696), .A2(n10697), .ZN(n10694) );
  INV_X1 U10525 ( .A(n8723), .ZN(n10466) );
  NAND2_X1 U10526 ( .A1(b_24_), .A2(a_24_), .ZN(n8723) );
  XNOR2_X1 U10527 ( .A(n10698), .B(n10699), .ZN(n10468) );
  XNOR2_X1 U10528 ( .A(n10700), .B(n10701), .ZN(n10698) );
  NOR2_X1 U10529 ( .A1(n8745), .A2(n8746), .ZN(n10701) );
  XNOR2_X1 U10530 ( .A(n10702), .B(n10703), .ZN(n10471) );
  XOR2_X1 U10531 ( .A(n10704), .B(n8068), .Z(n10703) );
  XNOR2_X1 U10532 ( .A(n10705), .B(n10706), .ZN(n10476) );
  XOR2_X1 U10533 ( .A(n10707), .B(n10708), .Z(n10706) );
  NAND2_X1 U10534 ( .A1(b_23_), .A2(a_22_), .ZN(n10708) );
  XNOR2_X1 U10535 ( .A(n10709), .B(n10710), .ZN(n10480) );
  XOR2_X1 U10536 ( .A(n10711), .B(n10712), .Z(n10709) );
  XNOR2_X1 U10537 ( .A(n10713), .B(n10714), .ZN(n10483) );
  XNOR2_X1 U10538 ( .A(n10715), .B(n10716), .ZN(n10713) );
  NOR2_X1 U10539 ( .A1(n8751), .A2(n8746), .ZN(n10716) );
  XOR2_X1 U10540 ( .A(n10717), .B(n10718), .Z(n10488) );
  XNOR2_X1 U10541 ( .A(n10719), .B(n10720), .ZN(n10718) );
  XNOR2_X1 U10542 ( .A(n10721), .B(n10722), .ZN(n10492) );
  XNOR2_X1 U10543 ( .A(n10723), .B(n10724), .ZN(n10721) );
  NOR2_X1 U10544 ( .A1(n8753), .A2(n8746), .ZN(n10724) );
  XNOR2_X1 U10545 ( .A(n10725), .B(n10726), .ZN(n10496) );
  XNOR2_X1 U10546 ( .A(n10727), .B(n10728), .ZN(n10725) );
  XNOR2_X1 U10547 ( .A(n10729), .B(n10730), .ZN(n10499) );
  XOR2_X1 U10548 ( .A(n10731), .B(n10732), .Z(n10730) );
  NAND2_X1 U10549 ( .A1(b_23_), .A2(a_16_), .ZN(n10732) );
  XOR2_X1 U10550 ( .A(n10733), .B(n10734), .Z(n10504) );
  XOR2_X1 U10551 ( .A(n10735), .B(n10736), .Z(n10734) );
  NAND2_X1 U10552 ( .A1(b_23_), .A2(a_15_), .ZN(n10736) );
  XOR2_X1 U10553 ( .A(n10737), .B(n10738), .Z(n10508) );
  NAND2_X1 U10554 ( .A1(n10739), .A2(n10740), .ZN(n10737) );
  XOR2_X1 U10555 ( .A(n10741), .B(n10742), .Z(n10511) );
  XOR2_X1 U10556 ( .A(n10743), .B(n10744), .Z(n10741) );
  XNOR2_X1 U10557 ( .A(n10745), .B(n10746), .ZN(n10515) );
  XNOR2_X1 U10558 ( .A(n10747), .B(n10748), .ZN(n10745) );
  NOR2_X1 U10559 ( .A1(n8759), .A2(n8746), .ZN(n10748) );
  XOR2_X1 U10560 ( .A(n10749), .B(n10750), .Z(n10519) );
  XOR2_X1 U10561 ( .A(n10751), .B(n10752), .Z(n10749) );
  NOR2_X1 U10562 ( .A1(n8376), .A2(n8746), .ZN(n10752) );
  XNOR2_X1 U10563 ( .A(n10753), .B(n10754), .ZN(n10523) );
  NAND2_X1 U10564 ( .A1(n10755), .A2(n10756), .ZN(n10753) );
  XOR2_X1 U10565 ( .A(n10757), .B(n10758), .Z(n10528) );
  XNOR2_X1 U10566 ( .A(n10759), .B(n10760), .ZN(n10758) );
  NAND2_X1 U10567 ( .A1(n10538), .A2(n10537), .ZN(n10593) );
  XNOR2_X1 U10568 ( .A(n10761), .B(n10762), .ZN(n10537) );
  XNOR2_X1 U10569 ( .A(n10763), .B(n10764), .ZN(n10761) );
  NOR2_X1 U10570 ( .A1(n8764), .A2(n8746), .ZN(n10764) );
  NOR2_X1 U10571 ( .A1(n8043), .A2(n8491), .ZN(n10538) );
  XOR2_X1 U10572 ( .A(n10765), .B(n10766), .Z(n10541) );
  NAND2_X1 U10573 ( .A1(n10767), .A2(n10768), .ZN(n10765) );
  XNOR2_X1 U10574 ( .A(n10769), .B(n10770), .ZN(n10545) );
  XOR2_X1 U10575 ( .A(n10771), .B(n10772), .Z(n10769) );
  NOR2_X1 U10576 ( .A1(n8517), .A2(n8746), .ZN(n10772) );
  NAND2_X1 U10577 ( .A1(n10773), .A2(n10774), .ZN(n10568) );
  INV_X1 U10578 ( .A(n10556), .ZN(n10774) );
  XOR2_X1 U10579 ( .A(n10775), .B(n10776), .Z(n10556) );
  XOR2_X1 U10580 ( .A(n10777), .B(n10778), .Z(n10776) );
  NAND2_X1 U10581 ( .A1(b_23_), .A2(a_2_), .ZN(n10778) );
  INV_X1 U10582 ( .A(n10559), .ZN(n10773) );
  NAND2_X1 U10583 ( .A1(b_24_), .A2(a_1_), .ZN(n10559) );
  XNOR2_X1 U10584 ( .A(n10779), .B(n10780), .ZN(n10561) );
  XOR2_X1 U10585 ( .A(n10781), .B(n10782), .Z(n10780) );
  NAND2_X1 U10586 ( .A1(b_23_), .A2(a_1_), .ZN(n10782) );
  INV_X1 U10587 ( .A(n8992), .ZN(n8987) );
  XOR2_X1 U10588 ( .A(n10783), .B(n10784), .Z(n8992) );
  XOR2_X1 U10589 ( .A(n10785), .B(n10786), .Z(n10784) );
  NAND2_X1 U10590 ( .A1(b_23_), .A2(a_0_), .ZN(n10786) );
  NAND3_X1 U10591 ( .A1(n8982), .A2(n8983), .A3(n10787), .ZN(n8833) );
  XOR2_X1 U10592 ( .A(n8978), .B(n8977), .Z(n10787) );
  NAND2_X1 U10593 ( .A1(n10788), .A2(n10789), .ZN(n8983) );
  NAND3_X1 U10594 ( .A1(a_0_), .A2(n10790), .A3(b_23_), .ZN(n10789) );
  OR2_X1 U10595 ( .A1(n10785), .A2(n10783), .ZN(n10790) );
  NAND2_X1 U10596 ( .A1(n10783), .A2(n10785), .ZN(n10788) );
  NAND2_X1 U10597 ( .A1(n10791), .A2(n10792), .ZN(n10785) );
  NAND3_X1 U10598 ( .A1(a_1_), .A2(n10793), .A3(b_23_), .ZN(n10792) );
  OR2_X1 U10599 ( .A1(n10781), .A2(n10779), .ZN(n10793) );
  NAND2_X1 U10600 ( .A1(n10779), .A2(n10781), .ZN(n10791) );
  NAND2_X1 U10601 ( .A1(n10794), .A2(n10795), .ZN(n10781) );
  NAND3_X1 U10602 ( .A1(a_2_), .A2(n10796), .A3(b_23_), .ZN(n10795) );
  OR2_X1 U10603 ( .A1(n10777), .A2(n10775), .ZN(n10796) );
  NAND2_X1 U10604 ( .A1(n10775), .A2(n10777), .ZN(n10794) );
  NAND2_X1 U10605 ( .A1(n10797), .A2(n10798), .ZN(n10777) );
  NAND3_X1 U10606 ( .A1(a_3_), .A2(n10799), .A3(b_23_), .ZN(n10798) );
  OR2_X1 U10607 ( .A1(n10577), .A2(n10575), .ZN(n10799) );
  NAND2_X1 U10608 ( .A1(n10575), .A2(n10577), .ZN(n10797) );
  NAND2_X1 U10609 ( .A1(n10800), .A2(n10801), .ZN(n10577) );
  NAND3_X1 U10610 ( .A1(a_4_), .A2(n10802), .A3(b_23_), .ZN(n10801) );
  OR2_X1 U10611 ( .A1(n10585), .A2(n10583), .ZN(n10802) );
  NAND2_X1 U10612 ( .A1(n10583), .A2(n10585), .ZN(n10800) );
  NAND2_X1 U10613 ( .A1(n10803), .A2(n10804), .ZN(n10585) );
  NAND3_X1 U10614 ( .A1(a_5_), .A2(n10805), .A3(b_23_), .ZN(n10804) );
  OR2_X1 U10615 ( .A1(n10771), .A2(n10770), .ZN(n10805) );
  NAND2_X1 U10616 ( .A1(n10770), .A2(n10771), .ZN(n10803) );
  NAND2_X1 U10617 ( .A1(n10767), .A2(n10806), .ZN(n10771) );
  NAND2_X1 U10618 ( .A1(n10766), .A2(n10768), .ZN(n10806) );
  NAND2_X1 U10619 ( .A1(n10807), .A2(n10808), .ZN(n10768) );
  NAND2_X1 U10620 ( .A1(b_23_), .A2(a_6_), .ZN(n10808) );
  INV_X1 U10621 ( .A(n10809), .ZN(n10807) );
  XOR2_X1 U10622 ( .A(n10810), .B(n10811), .Z(n10766) );
  XOR2_X1 U10623 ( .A(n10812), .B(n10813), .Z(n10810) );
  NAND2_X1 U10624 ( .A1(a_6_), .A2(n10809), .ZN(n10767) );
  NAND2_X1 U10625 ( .A1(n10814), .A2(n10815), .ZN(n10809) );
  NAND3_X1 U10626 ( .A1(a_7_), .A2(n10816), .A3(b_23_), .ZN(n10815) );
  NAND2_X1 U10627 ( .A1(n10763), .A2(n10762), .ZN(n10816) );
  OR2_X1 U10628 ( .A1(n10762), .A2(n10763), .ZN(n10814) );
  AND2_X1 U10629 ( .A1(n10817), .A2(n10818), .ZN(n10763) );
  NAND2_X1 U10630 ( .A1(n10603), .A2(n10819), .ZN(n10818) );
  OR2_X1 U10631 ( .A1(n10602), .A2(n10600), .ZN(n10819) );
  NOR2_X1 U10632 ( .A1(n8746), .A2(n8763), .ZN(n10603) );
  NAND2_X1 U10633 ( .A1(n10600), .A2(n10602), .ZN(n10817) );
  NAND2_X1 U10634 ( .A1(n10820), .A2(n10821), .ZN(n10602) );
  NAND2_X1 U10635 ( .A1(n10760), .A2(n10822), .ZN(n10821) );
  OR2_X1 U10636 ( .A1(n10759), .A2(n10757), .ZN(n10822) );
  NOR2_X1 U10637 ( .A1(n8746), .A2(n8426), .ZN(n10760) );
  NAND2_X1 U10638 ( .A1(n10757), .A2(n10759), .ZN(n10820) );
  NAND2_X1 U10639 ( .A1(n10755), .A2(n10823), .ZN(n10759) );
  NAND2_X1 U10640 ( .A1(n10754), .A2(n10756), .ZN(n10823) );
  NAND2_X1 U10641 ( .A1(n10824), .A2(n10825), .ZN(n10756) );
  NAND2_X1 U10642 ( .A1(b_23_), .A2(a_10_), .ZN(n10825) );
  INV_X1 U10643 ( .A(n10826), .ZN(n10824) );
  XNOR2_X1 U10644 ( .A(n10827), .B(n10828), .ZN(n10754) );
  XNOR2_X1 U10645 ( .A(n10829), .B(n10830), .ZN(n10828) );
  NAND2_X1 U10646 ( .A1(a_10_), .A2(n10826), .ZN(n10755) );
  NAND2_X1 U10647 ( .A1(n10831), .A2(n10832), .ZN(n10826) );
  NAND3_X1 U10648 ( .A1(a_11_), .A2(n10833), .A3(b_23_), .ZN(n10832) );
  OR2_X1 U10649 ( .A1(n10751), .A2(n10750), .ZN(n10833) );
  NAND2_X1 U10650 ( .A1(n10750), .A2(n10751), .ZN(n10831) );
  NAND2_X1 U10651 ( .A1(n10834), .A2(n10835), .ZN(n10751) );
  NAND3_X1 U10652 ( .A1(a_12_), .A2(n10836), .A3(b_23_), .ZN(n10835) );
  NAND2_X1 U10653 ( .A1(n10747), .A2(n10746), .ZN(n10836) );
  OR2_X1 U10654 ( .A1(n10746), .A2(n10747), .ZN(n10834) );
  AND2_X1 U10655 ( .A1(n10837), .A2(n10838), .ZN(n10747) );
  NAND2_X1 U10656 ( .A1(n10744), .A2(n10839), .ZN(n10838) );
  OR2_X1 U10657 ( .A1(n10743), .A2(n10742), .ZN(n10839) );
  NOR2_X1 U10658 ( .A1(n8746), .A2(n8310), .ZN(n10744) );
  NAND2_X1 U10659 ( .A1(n10742), .A2(n10743), .ZN(n10837) );
  NAND2_X1 U10660 ( .A1(n10739), .A2(n10840), .ZN(n10743) );
  NAND2_X1 U10661 ( .A1(n10738), .A2(n10740), .ZN(n10840) );
  NAND2_X1 U10662 ( .A1(n10841), .A2(n10842), .ZN(n10740) );
  NAND2_X1 U10663 ( .A1(b_23_), .A2(a_14_), .ZN(n10842) );
  INV_X1 U10664 ( .A(n10843), .ZN(n10841) );
  XOR2_X1 U10665 ( .A(n10844), .B(n10845), .Z(n10738) );
  XOR2_X1 U10666 ( .A(n10846), .B(n10847), .Z(n10844) );
  NAND2_X1 U10667 ( .A1(a_14_), .A2(n10843), .ZN(n10739) );
  NAND2_X1 U10668 ( .A1(n10848), .A2(n10849), .ZN(n10843) );
  NAND3_X1 U10669 ( .A1(a_15_), .A2(n10850), .A3(b_23_), .ZN(n10849) );
  OR2_X1 U10670 ( .A1(n10735), .A2(n10733), .ZN(n10850) );
  NAND2_X1 U10671 ( .A1(n10733), .A2(n10735), .ZN(n10848) );
  NAND2_X1 U10672 ( .A1(n10851), .A2(n10852), .ZN(n10735) );
  NAND3_X1 U10673 ( .A1(a_16_), .A2(n10853), .A3(b_23_), .ZN(n10852) );
  OR2_X1 U10674 ( .A1(n10731), .A2(n10729), .ZN(n10853) );
  NAND2_X1 U10675 ( .A1(n10729), .A2(n10731), .ZN(n10851) );
  NAND2_X1 U10676 ( .A1(n10854), .A2(n10855), .ZN(n10731) );
  NAND2_X1 U10677 ( .A1(n10728), .A2(n10856), .ZN(n10855) );
  NAND2_X1 U10678 ( .A1(n10727), .A2(n10726), .ZN(n10856) );
  NOR2_X1 U10679 ( .A1(n8746), .A2(n8210), .ZN(n10728) );
  OR2_X1 U10680 ( .A1(n10726), .A2(n10727), .ZN(n10854) );
  AND2_X1 U10681 ( .A1(n10857), .A2(n10858), .ZN(n10727) );
  NAND3_X1 U10682 ( .A1(a_18_), .A2(n10859), .A3(b_23_), .ZN(n10858) );
  NAND2_X1 U10683 ( .A1(n10723), .A2(n10722), .ZN(n10859) );
  OR2_X1 U10684 ( .A1(n10722), .A2(n10723), .ZN(n10857) );
  AND2_X1 U10685 ( .A1(n10860), .A2(n10861), .ZN(n10723) );
  NAND2_X1 U10686 ( .A1(n10720), .A2(n10862), .ZN(n10861) );
  OR2_X1 U10687 ( .A1(n10719), .A2(n10717), .ZN(n10862) );
  NOR2_X1 U10688 ( .A1(n8746), .A2(n8170), .ZN(n10720) );
  NAND2_X1 U10689 ( .A1(n10717), .A2(n10719), .ZN(n10860) );
  NAND2_X1 U10690 ( .A1(n10863), .A2(n10864), .ZN(n10719) );
  NAND3_X1 U10691 ( .A1(a_20_), .A2(n10865), .A3(b_23_), .ZN(n10864) );
  NAND2_X1 U10692 ( .A1(n10715), .A2(n10714), .ZN(n10865) );
  OR2_X1 U10693 ( .A1(n10714), .A2(n10715), .ZN(n10863) );
  AND2_X1 U10694 ( .A1(n10866), .A2(n10867), .ZN(n10715) );
  NAND2_X1 U10695 ( .A1(n10712), .A2(n10868), .ZN(n10867) );
  OR2_X1 U10696 ( .A1(n10711), .A2(n10710), .ZN(n10868) );
  NOR2_X1 U10697 ( .A1(n8746), .A2(n8750), .ZN(n10712) );
  NAND2_X1 U10698 ( .A1(n10710), .A2(n10711), .ZN(n10866) );
  NAND2_X1 U10699 ( .A1(n10869), .A2(n10870), .ZN(n10711) );
  NAND3_X1 U10700 ( .A1(a_22_), .A2(n10871), .A3(b_23_), .ZN(n10870) );
  OR2_X1 U10701 ( .A1(n10707), .A2(n10705), .ZN(n10871) );
  NAND2_X1 U10702 ( .A1(n10705), .A2(n10707), .ZN(n10869) );
  NAND2_X1 U10703 ( .A1(n10872), .A2(n10873), .ZN(n10707) );
  NAND2_X1 U10704 ( .A1(n10874), .A2(n10875), .ZN(n10873) );
  OR2_X1 U10705 ( .A1(n10704), .A2(n10702), .ZN(n10875) );
  INV_X1 U10706 ( .A(n8068), .ZN(n10874) );
  NAND2_X1 U10707 ( .A1(b_23_), .A2(a_23_), .ZN(n8068) );
  NAND2_X1 U10708 ( .A1(n10702), .A2(n10704), .ZN(n10872) );
  NAND2_X1 U10709 ( .A1(n10876), .A2(n10877), .ZN(n10704) );
  NAND3_X1 U10710 ( .A1(a_24_), .A2(n10878), .A3(b_23_), .ZN(n10877) );
  NAND2_X1 U10711 ( .A1(n10700), .A2(n10699), .ZN(n10878) );
  OR2_X1 U10712 ( .A1(n10699), .A2(n10700), .ZN(n10876) );
  AND2_X1 U10713 ( .A1(n10879), .A2(n10880), .ZN(n10700) );
  NAND2_X1 U10714 ( .A1(n10658), .A2(n10881), .ZN(n10880) );
  OR2_X1 U10715 ( .A1(n10657), .A2(n10656), .ZN(n10881) );
  NOR2_X1 U10716 ( .A1(n8746), .A2(n8744), .ZN(n10658) );
  NAND2_X1 U10717 ( .A1(n10656), .A2(n10657), .ZN(n10879) );
  NAND2_X1 U10718 ( .A1(n10696), .A2(n10882), .ZN(n10657) );
  NAND2_X1 U10719 ( .A1(n10695), .A2(n10697), .ZN(n10882) );
  NAND2_X1 U10720 ( .A1(n10883), .A2(n10884), .ZN(n10697) );
  NAND2_X1 U10721 ( .A1(b_23_), .A2(a_26_), .ZN(n10884) );
  INV_X1 U10722 ( .A(n10885), .ZN(n10883) );
  XNOR2_X1 U10723 ( .A(n10886), .B(n10887), .ZN(n10695) );
  NAND2_X1 U10724 ( .A1(n10888), .A2(n10889), .ZN(n10886) );
  NAND2_X1 U10725 ( .A1(a_26_), .A2(n10885), .ZN(n10696) );
  NAND2_X1 U10726 ( .A1(n10668), .A2(n10890), .ZN(n10885) );
  NAND2_X1 U10727 ( .A1(n10667), .A2(n10669), .ZN(n10890) );
  NAND2_X1 U10728 ( .A1(n10891), .A2(n10892), .ZN(n10669) );
  NAND2_X1 U10729 ( .A1(b_23_), .A2(a_27_), .ZN(n10892) );
  INV_X1 U10730 ( .A(n10893), .ZN(n10891) );
  XNOR2_X1 U10731 ( .A(n10894), .B(n10895), .ZN(n10667) );
  XOR2_X1 U10732 ( .A(n10896), .B(n10897), .Z(n10894) );
  NAND2_X1 U10733 ( .A1(b_22_), .A2(a_28_), .ZN(n10896) );
  NAND2_X1 U10734 ( .A1(a_27_), .A2(n10893), .ZN(n10668) );
  NAND2_X1 U10735 ( .A1(n10898), .A2(n10899), .ZN(n10893) );
  NAND3_X1 U10736 ( .A1(a_28_), .A2(n10900), .A3(b_23_), .ZN(n10899) );
  NAND2_X1 U10737 ( .A1(n10677), .A2(n10675), .ZN(n10900) );
  OR2_X1 U10738 ( .A1(n10675), .A2(n10677), .ZN(n10898) );
  AND2_X1 U10739 ( .A1(n10901), .A2(n10902), .ZN(n10677) );
  NAND2_X1 U10740 ( .A1(n10691), .A2(n10903), .ZN(n10902) );
  OR2_X1 U10741 ( .A1(n10692), .A2(n10693), .ZN(n10903) );
  NOR2_X1 U10742 ( .A1(n8746), .A2(n7890), .ZN(n10691) );
  NAND2_X1 U10743 ( .A1(n10693), .A2(n10692), .ZN(n10901) );
  NAND2_X1 U10744 ( .A1(n10904), .A2(n10905), .ZN(n10692) );
  NAND2_X1 U10745 ( .A1(b_21_), .A2(n10906), .ZN(n10905) );
  NAND2_X1 U10746 ( .A1(n7864), .A2(n10907), .ZN(n10906) );
  NAND2_X1 U10747 ( .A1(a_31_), .A2(n8094), .ZN(n10907) );
  NAND2_X1 U10748 ( .A1(b_22_), .A2(n10908), .ZN(n10904) );
  NAND2_X1 U10749 ( .A1(n9137), .A2(n10909), .ZN(n10908) );
  NAND2_X1 U10750 ( .A1(a_30_), .A2(n8749), .ZN(n10909) );
  AND3_X1 U10751 ( .A1(b_22_), .A2(b_23_), .A3(n7818), .ZN(n10693) );
  XNOR2_X1 U10752 ( .A(n10910), .B(n10911), .ZN(n10675) );
  XOR2_X1 U10753 ( .A(n10912), .B(n10913), .Z(n10910) );
  XNOR2_X1 U10754 ( .A(n10914), .B(n10915), .ZN(n10656) );
  NAND2_X1 U10755 ( .A1(n10916), .A2(n10917), .ZN(n10914) );
  XNOR2_X1 U10756 ( .A(n10918), .B(n10919), .ZN(n10699) );
  XOR2_X1 U10757 ( .A(n10920), .B(n10921), .Z(n10918) );
  XNOR2_X1 U10758 ( .A(n10922), .B(n10923), .ZN(n10702) );
  XNOR2_X1 U10759 ( .A(n10924), .B(n10925), .ZN(n10922) );
  NOR2_X1 U10760 ( .A1(n8745), .A2(n8094), .ZN(n10925) );
  XNOR2_X1 U10761 ( .A(n10926), .B(n10927), .ZN(n10705) );
  XNOR2_X1 U10762 ( .A(n10928), .B(n10929), .ZN(n10927) );
  XNOR2_X1 U10763 ( .A(n10930), .B(n10931), .ZN(n10710) );
  XNOR2_X1 U10764 ( .A(n10932), .B(n8719), .ZN(n10931) );
  XNOR2_X1 U10765 ( .A(n10933), .B(n10934), .ZN(n10714) );
  XOR2_X1 U10766 ( .A(n10935), .B(n10936), .Z(n10933) );
  XNOR2_X1 U10767 ( .A(n10937), .B(n10938), .ZN(n10717) );
  XNOR2_X1 U10768 ( .A(n10939), .B(n10940), .ZN(n10937) );
  NOR2_X1 U10769 ( .A1(n8751), .A2(n8094), .ZN(n10940) );
  XOR2_X1 U10770 ( .A(n10941), .B(n10942), .Z(n10722) );
  XNOR2_X1 U10771 ( .A(n10943), .B(n10944), .ZN(n10942) );
  XNOR2_X1 U10772 ( .A(n10945), .B(n10946), .ZN(n10726) );
  XOR2_X1 U10773 ( .A(n10947), .B(n10948), .Z(n10945) );
  NOR2_X1 U10774 ( .A1(n8753), .A2(n8094), .ZN(n10948) );
  XOR2_X1 U10775 ( .A(n10949), .B(n10950), .Z(n10729) );
  XOR2_X1 U10776 ( .A(n10951), .B(n10952), .Z(n10949) );
  XNOR2_X1 U10777 ( .A(n10953), .B(n10954), .ZN(n10733) );
  XOR2_X1 U10778 ( .A(n10955), .B(n10956), .Z(n10954) );
  NAND2_X1 U10779 ( .A1(b_22_), .A2(a_16_), .ZN(n10956) );
  XNOR2_X1 U10780 ( .A(n10957), .B(n10958), .ZN(n10742) );
  XNOR2_X1 U10781 ( .A(n10959), .B(n10960), .ZN(n10957) );
  NOR2_X1 U10782 ( .A1(n8757), .A2(n8094), .ZN(n10960) );
  XOR2_X1 U10783 ( .A(n10961), .B(n10962), .Z(n10746) );
  XNOR2_X1 U10784 ( .A(n10963), .B(n10964), .ZN(n10962) );
  XNOR2_X1 U10785 ( .A(n10965), .B(n10966), .ZN(n10750) );
  XNOR2_X1 U10786 ( .A(n10967), .B(n10968), .ZN(n10965) );
  NOR2_X1 U10787 ( .A1(n8759), .A2(n8094), .ZN(n10968) );
  XNOR2_X1 U10788 ( .A(n10969), .B(n10970), .ZN(n10757) );
  XNOR2_X1 U10789 ( .A(n10971), .B(n10972), .ZN(n10969) );
  NOR2_X1 U10790 ( .A1(n8761), .A2(n8094), .ZN(n10972) );
  XNOR2_X1 U10791 ( .A(n10973), .B(n10974), .ZN(n10600) );
  XOR2_X1 U10792 ( .A(n10975), .B(n10976), .Z(n10974) );
  NAND2_X1 U10793 ( .A1(b_22_), .A2(a_9_), .ZN(n10976) );
  XNOR2_X1 U10794 ( .A(n10977), .B(n10978), .ZN(n10762) );
  XOR2_X1 U10795 ( .A(n10979), .B(n10980), .Z(n10977) );
  XNOR2_X1 U10796 ( .A(n10981), .B(n10982), .ZN(n10770) );
  XNOR2_X1 U10797 ( .A(n10983), .B(n10984), .ZN(n10981) );
  XOR2_X1 U10798 ( .A(n10985), .B(n10986), .Z(n10583) );
  XOR2_X1 U10799 ( .A(n10987), .B(n10988), .Z(n10985) );
  NOR2_X1 U10800 ( .A1(n8517), .A2(n8094), .ZN(n10988) );
  XNOR2_X1 U10801 ( .A(n10989), .B(n10990), .ZN(n10575) );
  XNOR2_X1 U10802 ( .A(n10991), .B(n10992), .ZN(n10990) );
  XOR2_X1 U10803 ( .A(n10993), .B(n10994), .Z(n10775) );
  XOR2_X1 U10804 ( .A(n10995), .B(n10996), .Z(n10993) );
  XOR2_X1 U10805 ( .A(n10997), .B(n10998), .Z(n10779) );
  XOR2_X1 U10806 ( .A(n10999), .B(n11000), .Z(n10997) );
  XOR2_X1 U10807 ( .A(n11001), .B(n11002), .Z(n10783) );
  XOR2_X1 U10808 ( .A(n11003), .B(n11004), .Z(n11001) );
  NOR2_X1 U10809 ( .A1(n8617), .A2(n8094), .ZN(n11004) );
  XNOR2_X1 U10810 ( .A(n11005), .B(n11006), .ZN(n8982) );
  NAND2_X1 U10811 ( .A1(n11007), .A2(n11008), .ZN(n11005) );
  NAND4_X1 U10812 ( .A1(n8977), .A2(n8976), .A3(n8978), .A4(n8972), .ZN(n8839)
         );
  INV_X1 U10813 ( .A(n11009), .ZN(n8972) );
  NAND2_X1 U10814 ( .A1(n11007), .A2(n11010), .ZN(n8978) );
  NAND2_X1 U10815 ( .A1(n11006), .A2(n11008), .ZN(n11010) );
  NAND2_X1 U10816 ( .A1(n11011), .A2(n11012), .ZN(n11008) );
  NAND2_X1 U10817 ( .A1(b_22_), .A2(a_0_), .ZN(n11012) );
  INV_X1 U10818 ( .A(n11013), .ZN(n11011) );
  XOR2_X1 U10819 ( .A(n11014), .B(n11015), .Z(n11006) );
  XOR2_X1 U10820 ( .A(n11016), .B(n11017), .Z(n11014) );
  NOR2_X1 U10821 ( .A1(n8617), .A2(n8749), .ZN(n11017) );
  NAND2_X1 U10822 ( .A1(a_0_), .A2(n11013), .ZN(n11007) );
  NAND2_X1 U10823 ( .A1(n11018), .A2(n11019), .ZN(n11013) );
  NAND3_X1 U10824 ( .A1(a_1_), .A2(n11020), .A3(b_22_), .ZN(n11019) );
  OR2_X1 U10825 ( .A1(n11003), .A2(n11002), .ZN(n11020) );
  NAND2_X1 U10826 ( .A1(n11002), .A2(n11003), .ZN(n11018) );
  NAND2_X1 U10827 ( .A1(n11021), .A2(n11022), .ZN(n11003) );
  NAND2_X1 U10828 ( .A1(n11000), .A2(n11023), .ZN(n11022) );
  OR2_X1 U10829 ( .A1(n10999), .A2(n10998), .ZN(n11023) );
  NOR2_X1 U10830 ( .A1(n8094), .A2(n8768), .ZN(n11000) );
  NAND2_X1 U10831 ( .A1(n10998), .A2(n10999), .ZN(n11021) );
  NAND2_X1 U10832 ( .A1(n11024), .A2(n11025), .ZN(n10999) );
  NAND2_X1 U10833 ( .A1(n10996), .A2(n11026), .ZN(n11025) );
  OR2_X1 U10834 ( .A1(n10995), .A2(n10994), .ZN(n11026) );
  NOR2_X1 U10835 ( .A1(n8094), .A2(n8567), .ZN(n10996) );
  NAND2_X1 U10836 ( .A1(n10994), .A2(n10995), .ZN(n11024) );
  NAND2_X1 U10837 ( .A1(n11027), .A2(n11028), .ZN(n10995) );
  NAND2_X1 U10838 ( .A1(n10992), .A2(n11029), .ZN(n11028) );
  OR2_X1 U10839 ( .A1(n10991), .A2(n10989), .ZN(n11029) );
  NOR2_X1 U10840 ( .A1(n8094), .A2(n8766), .ZN(n10992) );
  NAND2_X1 U10841 ( .A1(n10989), .A2(n10991), .ZN(n11027) );
  NAND2_X1 U10842 ( .A1(n11030), .A2(n11031), .ZN(n10991) );
  NAND3_X1 U10843 ( .A1(a_5_), .A2(n11032), .A3(b_22_), .ZN(n11031) );
  OR2_X1 U10844 ( .A1(n10987), .A2(n10986), .ZN(n11032) );
  NAND2_X1 U10845 ( .A1(n10986), .A2(n10987), .ZN(n11030) );
  NAND2_X1 U10846 ( .A1(n11033), .A2(n11034), .ZN(n10987) );
  NAND2_X1 U10847 ( .A1(n10984), .A2(n11035), .ZN(n11034) );
  NAND2_X1 U10848 ( .A1(n10983), .A2(n10982), .ZN(n11035) );
  NOR2_X1 U10849 ( .A1(n8094), .A2(n8491), .ZN(n10984) );
  OR2_X1 U10850 ( .A1(n10982), .A2(n10983), .ZN(n11033) );
  AND2_X1 U10851 ( .A1(n11036), .A2(n11037), .ZN(n10983) );
  NAND2_X1 U10852 ( .A1(n10813), .A2(n11038), .ZN(n11037) );
  OR2_X1 U10853 ( .A1(n10812), .A2(n10811), .ZN(n11038) );
  NOR2_X1 U10854 ( .A1(n8094), .A2(n8764), .ZN(n10813) );
  NAND2_X1 U10855 ( .A1(n10811), .A2(n10812), .ZN(n11036) );
  NAND2_X1 U10856 ( .A1(n11039), .A2(n11040), .ZN(n10812) );
  NAND2_X1 U10857 ( .A1(n10980), .A2(n11041), .ZN(n11040) );
  OR2_X1 U10858 ( .A1(n10979), .A2(n10978), .ZN(n11041) );
  NOR2_X1 U10859 ( .A1(n8094), .A2(n8763), .ZN(n10980) );
  NAND2_X1 U10860 ( .A1(n10978), .A2(n10979), .ZN(n11039) );
  NAND2_X1 U10861 ( .A1(n11042), .A2(n11043), .ZN(n10979) );
  NAND3_X1 U10862 ( .A1(a_9_), .A2(n11044), .A3(b_22_), .ZN(n11043) );
  OR2_X1 U10863 ( .A1(n10975), .A2(n10973), .ZN(n11044) );
  NAND2_X1 U10864 ( .A1(n10973), .A2(n10975), .ZN(n11042) );
  NAND2_X1 U10865 ( .A1(n11045), .A2(n11046), .ZN(n10975) );
  NAND3_X1 U10866 ( .A1(a_10_), .A2(n11047), .A3(b_22_), .ZN(n11046) );
  NAND2_X1 U10867 ( .A1(n10971), .A2(n10970), .ZN(n11047) );
  OR2_X1 U10868 ( .A1(n10970), .A2(n10971), .ZN(n11045) );
  AND2_X1 U10869 ( .A1(n11048), .A2(n11049), .ZN(n10971) );
  NAND2_X1 U10870 ( .A1(n10830), .A2(n11050), .ZN(n11049) );
  OR2_X1 U10871 ( .A1(n10829), .A2(n10827), .ZN(n11050) );
  NOR2_X1 U10872 ( .A1(n8094), .A2(n8376), .ZN(n10830) );
  NAND2_X1 U10873 ( .A1(n10827), .A2(n10829), .ZN(n11048) );
  NAND2_X1 U10874 ( .A1(n11051), .A2(n11052), .ZN(n10829) );
  NAND3_X1 U10875 ( .A1(a_12_), .A2(n11053), .A3(b_22_), .ZN(n11052) );
  NAND2_X1 U10876 ( .A1(n10967), .A2(n10966), .ZN(n11053) );
  OR2_X1 U10877 ( .A1(n10966), .A2(n10967), .ZN(n11051) );
  AND2_X1 U10878 ( .A1(n11054), .A2(n11055), .ZN(n10967) );
  NAND2_X1 U10879 ( .A1(n10964), .A2(n11056), .ZN(n11055) );
  OR2_X1 U10880 ( .A1(n10963), .A2(n10961), .ZN(n11056) );
  NOR2_X1 U10881 ( .A1(n8094), .A2(n8310), .ZN(n10964) );
  NAND2_X1 U10882 ( .A1(n10961), .A2(n10963), .ZN(n11054) );
  NAND2_X1 U10883 ( .A1(n11057), .A2(n11058), .ZN(n10963) );
  NAND3_X1 U10884 ( .A1(a_14_), .A2(n11059), .A3(b_22_), .ZN(n11058) );
  NAND2_X1 U10885 ( .A1(n10959), .A2(n10958), .ZN(n11059) );
  OR2_X1 U10886 ( .A1(n10958), .A2(n10959), .ZN(n11057) );
  AND2_X1 U10887 ( .A1(n11060), .A2(n11061), .ZN(n10959) );
  NAND2_X1 U10888 ( .A1(n10847), .A2(n11062), .ZN(n11061) );
  OR2_X1 U10889 ( .A1(n10846), .A2(n10845), .ZN(n11062) );
  NOR2_X1 U10890 ( .A1(n8094), .A2(n8276), .ZN(n10847) );
  NAND2_X1 U10891 ( .A1(n10845), .A2(n10846), .ZN(n11060) );
  NAND2_X1 U10892 ( .A1(n11063), .A2(n11064), .ZN(n10846) );
  NAND3_X1 U10893 ( .A1(a_16_), .A2(n11065), .A3(b_22_), .ZN(n11064) );
  OR2_X1 U10894 ( .A1(n10955), .A2(n10953), .ZN(n11065) );
  NAND2_X1 U10895 ( .A1(n10953), .A2(n10955), .ZN(n11063) );
  NAND2_X1 U10896 ( .A1(n11066), .A2(n11067), .ZN(n10955) );
  NAND2_X1 U10897 ( .A1(n10952), .A2(n11068), .ZN(n11067) );
  OR2_X1 U10898 ( .A1(n10951), .A2(n10950), .ZN(n11068) );
  NOR2_X1 U10899 ( .A1(n8094), .A2(n8210), .ZN(n10952) );
  NAND2_X1 U10900 ( .A1(n10950), .A2(n10951), .ZN(n11066) );
  NAND2_X1 U10901 ( .A1(n11069), .A2(n11070), .ZN(n10951) );
  NAND3_X1 U10902 ( .A1(a_18_), .A2(n11071), .A3(b_22_), .ZN(n11070) );
  OR2_X1 U10903 ( .A1(n10947), .A2(n10946), .ZN(n11071) );
  NAND2_X1 U10904 ( .A1(n10946), .A2(n10947), .ZN(n11069) );
  NAND2_X1 U10905 ( .A1(n11072), .A2(n11073), .ZN(n10947) );
  NAND2_X1 U10906 ( .A1(n10944), .A2(n11074), .ZN(n11073) );
  OR2_X1 U10907 ( .A1(n10943), .A2(n10941), .ZN(n11074) );
  NOR2_X1 U10908 ( .A1(n8094), .A2(n8170), .ZN(n10944) );
  NAND2_X1 U10909 ( .A1(n10941), .A2(n10943), .ZN(n11072) );
  NAND2_X1 U10910 ( .A1(n11075), .A2(n11076), .ZN(n10943) );
  NAND3_X1 U10911 ( .A1(a_20_), .A2(n11077), .A3(b_22_), .ZN(n11076) );
  NAND2_X1 U10912 ( .A1(n10939), .A2(n10938), .ZN(n11077) );
  OR2_X1 U10913 ( .A1(n10938), .A2(n10939), .ZN(n11075) );
  AND2_X1 U10914 ( .A1(n11078), .A2(n11079), .ZN(n10939) );
  NAND2_X1 U10915 ( .A1(n10936), .A2(n11080), .ZN(n11079) );
  OR2_X1 U10916 ( .A1(n10935), .A2(n10934), .ZN(n11080) );
  NOR2_X1 U10917 ( .A1(n8094), .A2(n8750), .ZN(n10936) );
  NAND2_X1 U10918 ( .A1(n10934), .A2(n10935), .ZN(n11078) );
  NAND2_X1 U10919 ( .A1(n11081), .A2(n11082), .ZN(n10935) );
  NAND2_X1 U10920 ( .A1(n10930), .A2(n11083), .ZN(n11082) );
  OR2_X1 U10921 ( .A1(n10932), .A2(n8719), .ZN(n11083) );
  XNOR2_X1 U10922 ( .A(n11084), .B(n11085), .ZN(n10930) );
  XNOR2_X1 U10923 ( .A(n11086), .B(n11087), .ZN(n11085) );
  NAND2_X1 U10924 ( .A1(n8719), .A2(n10932), .ZN(n11081) );
  NAND2_X1 U10925 ( .A1(n11088), .A2(n11089), .ZN(n10932) );
  NAND2_X1 U10926 ( .A1(n10929), .A2(n11090), .ZN(n11089) );
  OR2_X1 U10927 ( .A1(n10928), .A2(n10926), .ZN(n11090) );
  NOR2_X1 U10928 ( .A1(n8094), .A2(n8747), .ZN(n10929) );
  NAND2_X1 U10929 ( .A1(n10926), .A2(n10928), .ZN(n11088) );
  NAND2_X1 U10930 ( .A1(n11091), .A2(n11092), .ZN(n10928) );
  NAND3_X1 U10931 ( .A1(a_24_), .A2(n11093), .A3(b_22_), .ZN(n11092) );
  NAND2_X1 U10932 ( .A1(n10924), .A2(n10923), .ZN(n11093) );
  OR2_X1 U10933 ( .A1(n10923), .A2(n10924), .ZN(n11091) );
  AND2_X1 U10934 ( .A1(n11094), .A2(n11095), .ZN(n10924) );
  NAND2_X1 U10935 ( .A1(n10921), .A2(n11096), .ZN(n11095) );
  OR2_X1 U10936 ( .A1(n10920), .A2(n10919), .ZN(n11096) );
  NOR2_X1 U10937 ( .A1(n8094), .A2(n8744), .ZN(n10921) );
  NAND2_X1 U10938 ( .A1(n10919), .A2(n10920), .ZN(n11094) );
  NAND2_X1 U10939 ( .A1(n10916), .A2(n11097), .ZN(n10920) );
  NAND2_X1 U10940 ( .A1(n10915), .A2(n10917), .ZN(n11097) );
  NAND2_X1 U10941 ( .A1(n11098), .A2(n11099), .ZN(n10917) );
  NAND2_X1 U10942 ( .A1(b_22_), .A2(a_26_), .ZN(n11099) );
  INV_X1 U10943 ( .A(n11100), .ZN(n11098) );
  XNOR2_X1 U10944 ( .A(n11101), .B(n11102), .ZN(n10915) );
  NAND2_X1 U10945 ( .A1(n11103), .A2(n11104), .ZN(n11101) );
  NAND2_X1 U10946 ( .A1(a_26_), .A2(n11100), .ZN(n10916) );
  NAND2_X1 U10947 ( .A1(n10888), .A2(n11105), .ZN(n11100) );
  NAND2_X1 U10948 ( .A1(n10887), .A2(n10889), .ZN(n11105) );
  NAND2_X1 U10949 ( .A1(n11106), .A2(n11107), .ZN(n10889) );
  NAND2_X1 U10950 ( .A1(b_22_), .A2(a_27_), .ZN(n11107) );
  INV_X1 U10951 ( .A(n11108), .ZN(n11106) );
  XNOR2_X1 U10952 ( .A(n11109), .B(n11110), .ZN(n10887) );
  XOR2_X1 U10953 ( .A(n11111), .B(n11112), .Z(n11109) );
  NAND2_X1 U10954 ( .A1(b_21_), .A2(a_28_), .ZN(n11111) );
  NAND2_X1 U10955 ( .A1(a_27_), .A2(n11108), .ZN(n10888) );
  NAND2_X1 U10956 ( .A1(n11113), .A2(n11114), .ZN(n11108) );
  NAND3_X1 U10957 ( .A1(a_28_), .A2(n11115), .A3(b_22_), .ZN(n11114) );
  NAND2_X1 U10958 ( .A1(n10897), .A2(n10895), .ZN(n11115) );
  OR2_X1 U10959 ( .A1(n10895), .A2(n10897), .ZN(n11113) );
  AND2_X1 U10960 ( .A1(n11116), .A2(n11117), .ZN(n10897) );
  NAND2_X1 U10961 ( .A1(n10911), .A2(n11118), .ZN(n11117) );
  OR2_X1 U10962 ( .A1(n10912), .A2(n10913), .ZN(n11118) );
  NOR2_X1 U10963 ( .A1(n8094), .A2(n7890), .ZN(n10911) );
  NAND2_X1 U10964 ( .A1(n10913), .A2(n10912), .ZN(n11116) );
  NAND2_X1 U10965 ( .A1(n11119), .A2(n11120), .ZN(n10912) );
  NAND2_X1 U10966 ( .A1(b_20_), .A2(n11121), .ZN(n11120) );
  NAND2_X1 U10967 ( .A1(n7864), .A2(n11122), .ZN(n11121) );
  NAND2_X1 U10968 ( .A1(a_31_), .A2(n8749), .ZN(n11122) );
  NAND2_X1 U10969 ( .A1(b_21_), .A2(n11123), .ZN(n11119) );
  NAND2_X1 U10970 ( .A1(n9137), .A2(n11124), .ZN(n11123) );
  NAND2_X1 U10971 ( .A1(a_30_), .A2(n8145), .ZN(n11124) );
  AND3_X1 U10972 ( .A1(b_21_), .A2(b_22_), .A3(n7818), .ZN(n10913) );
  XNOR2_X1 U10973 ( .A(n11125), .B(n11126), .ZN(n10895) );
  XOR2_X1 U10974 ( .A(n11127), .B(n11128), .Z(n11125) );
  XNOR2_X1 U10975 ( .A(n11129), .B(n11130), .ZN(n10919) );
  NAND2_X1 U10976 ( .A1(n11131), .A2(n11132), .ZN(n11129) );
  XNOR2_X1 U10977 ( .A(n11133), .B(n11134), .ZN(n10923) );
  XOR2_X1 U10978 ( .A(n11135), .B(n11136), .Z(n11133) );
  XNOR2_X1 U10979 ( .A(n11137), .B(n11138), .ZN(n10926) );
  XNOR2_X1 U10980 ( .A(n11139), .B(n11140), .ZN(n11137) );
  NOR2_X1 U10981 ( .A1(n8745), .A2(n8749), .ZN(n11140) );
  NOR2_X1 U10982 ( .A1(n8094), .A2(n8748), .ZN(n8719) );
  XNOR2_X1 U10983 ( .A(n11141), .B(n11142), .ZN(n10934) );
  XOR2_X1 U10984 ( .A(n11143), .B(n11144), .Z(n11142) );
  NAND2_X1 U10985 ( .A1(b_21_), .A2(a_22_), .ZN(n11144) );
  XNOR2_X1 U10986 ( .A(n11145), .B(n11146), .ZN(n10938) );
  XOR2_X1 U10987 ( .A(n11147), .B(n11148), .Z(n11145) );
  XNOR2_X1 U10988 ( .A(n11149), .B(n11150), .ZN(n10941) );
  XNOR2_X1 U10989 ( .A(n11151), .B(n11152), .ZN(n11149) );
  NOR2_X1 U10990 ( .A1(n8751), .A2(n8749), .ZN(n11152) );
  XNOR2_X1 U10991 ( .A(n11153), .B(n11154), .ZN(n10946) );
  XNOR2_X1 U10992 ( .A(n11155), .B(n11156), .ZN(n11154) );
  XNOR2_X1 U10993 ( .A(n11157), .B(n11158), .ZN(n10950) );
  XNOR2_X1 U10994 ( .A(n11159), .B(n11160), .ZN(n11157) );
  NOR2_X1 U10995 ( .A1(n8753), .A2(n8749), .ZN(n11160) );
  XNOR2_X1 U10996 ( .A(n11161), .B(n11162), .ZN(n10953) );
  XNOR2_X1 U10997 ( .A(n11163), .B(n11164), .ZN(n11162) );
  XNOR2_X1 U10998 ( .A(n11165), .B(n11166), .ZN(n10845) );
  XNOR2_X1 U10999 ( .A(n11167), .B(n11168), .ZN(n11165) );
  NOR2_X1 U11000 ( .A1(n8755), .A2(n8749), .ZN(n11168) );
  XNOR2_X1 U11001 ( .A(n11169), .B(n11170), .ZN(n10958) );
  XOR2_X1 U11002 ( .A(n11171), .B(n11172), .Z(n11169) );
  XNOR2_X1 U11003 ( .A(n11173), .B(n11174), .ZN(n10961) );
  XNOR2_X1 U11004 ( .A(n11175), .B(n11176), .ZN(n11173) );
  NOR2_X1 U11005 ( .A1(n8757), .A2(n8749), .ZN(n11176) );
  XNOR2_X1 U11006 ( .A(n11177), .B(n11178), .ZN(n10966) );
  XOR2_X1 U11007 ( .A(n11179), .B(n11180), .Z(n11177) );
  XNOR2_X1 U11008 ( .A(n11181), .B(n11182), .ZN(n10827) );
  XOR2_X1 U11009 ( .A(n11183), .B(n11184), .Z(n11182) );
  NAND2_X1 U11010 ( .A1(b_21_), .A2(a_12_), .ZN(n11184) );
  XOR2_X1 U11011 ( .A(n11185), .B(n11186), .Z(n10970) );
  XNOR2_X1 U11012 ( .A(n11187), .B(n11188), .ZN(n11186) );
  XOR2_X1 U11013 ( .A(n11189), .B(n11190), .Z(n10973) );
  XOR2_X1 U11014 ( .A(n11191), .B(n11192), .Z(n11189) );
  XNOR2_X1 U11015 ( .A(n11193), .B(n11194), .ZN(n10978) );
  XOR2_X1 U11016 ( .A(n11195), .B(n11196), .Z(n11193) );
  NAND2_X1 U11017 ( .A1(b_21_), .A2(a_9_), .ZN(n11195) );
  XNOR2_X1 U11018 ( .A(n11197), .B(n11198), .ZN(n10811) );
  XOR2_X1 U11019 ( .A(n11199), .B(n11200), .Z(n11198) );
  NAND2_X1 U11020 ( .A1(b_21_), .A2(a_8_), .ZN(n11200) );
  XOR2_X1 U11021 ( .A(n11201), .B(n11202), .Z(n10982) );
  XOR2_X1 U11022 ( .A(n11203), .B(n11204), .Z(n11202) );
  NAND2_X1 U11023 ( .A1(b_21_), .A2(a_7_), .ZN(n11204) );
  XNOR2_X1 U11024 ( .A(n11205), .B(n11206), .ZN(n10986) );
  XOR2_X1 U11025 ( .A(n11207), .B(n11208), .Z(n11206) );
  NAND2_X1 U11026 ( .A1(b_21_), .A2(a_6_), .ZN(n11208) );
  XNOR2_X1 U11027 ( .A(n11209), .B(n11210), .ZN(n10989) );
  XNOR2_X1 U11028 ( .A(n11211), .B(n11212), .ZN(n11209) );
  NOR2_X1 U11029 ( .A1(n8517), .A2(n8749), .ZN(n11212) );
  XNOR2_X1 U11030 ( .A(n11213), .B(n11214), .ZN(n10994) );
  XOR2_X1 U11031 ( .A(n11215), .B(n11216), .Z(n11214) );
  NAND2_X1 U11032 ( .A1(b_21_), .A2(a_4_), .ZN(n11216) );
  XNOR2_X1 U11033 ( .A(n11217), .B(n11218), .ZN(n10998) );
  XOR2_X1 U11034 ( .A(n11219), .B(n11220), .Z(n11218) );
  NAND2_X1 U11035 ( .A1(b_21_), .A2(a_3_), .ZN(n11220) );
  XNOR2_X1 U11036 ( .A(n11221), .B(n11222), .ZN(n11002) );
  XOR2_X1 U11037 ( .A(n11223), .B(n11224), .Z(n11222) );
  NAND2_X1 U11038 ( .A1(b_21_), .A2(a_2_), .ZN(n11224) );
  NAND2_X1 U11039 ( .A1(n11225), .A2(n11226), .ZN(n8976) );
  XNOR2_X1 U11040 ( .A(n11227), .B(n11228), .ZN(n8977) );
  XNOR2_X1 U11041 ( .A(n11229), .B(n11230), .ZN(n11228) );
  NAND2_X1 U11042 ( .A1(n11231), .A2(n11009), .ZN(n8845) );
  NOR2_X1 U11043 ( .A1(n11226), .A2(n11225), .ZN(n11009) );
  AND2_X1 U11044 ( .A1(n11232), .A2(n11233), .ZN(n11225) );
  NAND2_X1 U11045 ( .A1(n11230), .A2(n11234), .ZN(n11233) );
  OR2_X1 U11046 ( .A1(n11229), .A2(n11227), .ZN(n11234) );
  NOR2_X1 U11047 ( .A1(n8749), .A2(n9674), .ZN(n11230) );
  NAND2_X1 U11048 ( .A1(n11227), .A2(n11229), .ZN(n11232) );
  NAND2_X1 U11049 ( .A1(n11235), .A2(n11236), .ZN(n11229) );
  NAND3_X1 U11050 ( .A1(a_1_), .A2(n11237), .A3(b_21_), .ZN(n11236) );
  OR2_X1 U11051 ( .A1(n11016), .A2(n11015), .ZN(n11237) );
  NAND2_X1 U11052 ( .A1(n11015), .A2(n11016), .ZN(n11235) );
  NAND2_X1 U11053 ( .A1(n11238), .A2(n11239), .ZN(n11016) );
  NAND3_X1 U11054 ( .A1(a_2_), .A2(n11240), .A3(b_21_), .ZN(n11239) );
  OR2_X1 U11055 ( .A1(n11223), .A2(n11221), .ZN(n11240) );
  NAND2_X1 U11056 ( .A1(n11221), .A2(n11223), .ZN(n11238) );
  NAND2_X1 U11057 ( .A1(n11241), .A2(n11242), .ZN(n11223) );
  NAND3_X1 U11058 ( .A1(a_3_), .A2(n11243), .A3(b_21_), .ZN(n11242) );
  OR2_X1 U11059 ( .A1(n11219), .A2(n11217), .ZN(n11243) );
  NAND2_X1 U11060 ( .A1(n11217), .A2(n11219), .ZN(n11241) );
  NAND2_X1 U11061 ( .A1(n11244), .A2(n11245), .ZN(n11219) );
  NAND3_X1 U11062 ( .A1(a_4_), .A2(n11246), .A3(b_21_), .ZN(n11245) );
  OR2_X1 U11063 ( .A1(n11215), .A2(n11213), .ZN(n11246) );
  NAND2_X1 U11064 ( .A1(n11213), .A2(n11215), .ZN(n11244) );
  NAND2_X1 U11065 ( .A1(n11247), .A2(n11248), .ZN(n11215) );
  NAND3_X1 U11066 ( .A1(a_5_), .A2(n11249), .A3(b_21_), .ZN(n11248) );
  NAND2_X1 U11067 ( .A1(n11211), .A2(n11210), .ZN(n11249) );
  OR2_X1 U11068 ( .A1(n11210), .A2(n11211), .ZN(n11247) );
  AND2_X1 U11069 ( .A1(n11250), .A2(n11251), .ZN(n11211) );
  NAND3_X1 U11070 ( .A1(a_6_), .A2(n11252), .A3(b_21_), .ZN(n11251) );
  OR2_X1 U11071 ( .A1(n11207), .A2(n11205), .ZN(n11252) );
  NAND2_X1 U11072 ( .A1(n11205), .A2(n11207), .ZN(n11250) );
  NAND2_X1 U11073 ( .A1(n11253), .A2(n11254), .ZN(n11207) );
  NAND3_X1 U11074 ( .A1(a_7_), .A2(n11255), .A3(b_21_), .ZN(n11254) );
  OR2_X1 U11075 ( .A1(n11203), .A2(n11201), .ZN(n11255) );
  NAND2_X1 U11076 ( .A1(n11201), .A2(n11203), .ZN(n11253) );
  NAND2_X1 U11077 ( .A1(n11256), .A2(n11257), .ZN(n11203) );
  NAND3_X1 U11078 ( .A1(a_8_), .A2(n11258), .A3(b_21_), .ZN(n11257) );
  OR2_X1 U11079 ( .A1(n11199), .A2(n11197), .ZN(n11258) );
  NAND2_X1 U11080 ( .A1(n11197), .A2(n11199), .ZN(n11256) );
  NAND2_X1 U11081 ( .A1(n11259), .A2(n11260), .ZN(n11199) );
  NAND3_X1 U11082 ( .A1(a_9_), .A2(n11261), .A3(b_21_), .ZN(n11260) );
  NAND2_X1 U11083 ( .A1(n11196), .A2(n11194), .ZN(n11261) );
  OR2_X1 U11084 ( .A1(n11194), .A2(n11196), .ZN(n11259) );
  AND2_X1 U11085 ( .A1(n11262), .A2(n11263), .ZN(n11196) );
  NAND2_X1 U11086 ( .A1(n11192), .A2(n11264), .ZN(n11263) );
  OR2_X1 U11087 ( .A1(n11191), .A2(n11190), .ZN(n11264) );
  NOR2_X1 U11088 ( .A1(n8749), .A2(n8761), .ZN(n11192) );
  NAND2_X1 U11089 ( .A1(n11190), .A2(n11191), .ZN(n11262) );
  NAND2_X1 U11090 ( .A1(n11265), .A2(n11266), .ZN(n11191) );
  NAND2_X1 U11091 ( .A1(n11188), .A2(n11267), .ZN(n11266) );
  OR2_X1 U11092 ( .A1(n11187), .A2(n11185), .ZN(n11267) );
  NOR2_X1 U11093 ( .A1(n8749), .A2(n8376), .ZN(n11188) );
  NAND2_X1 U11094 ( .A1(n11185), .A2(n11187), .ZN(n11265) );
  NAND2_X1 U11095 ( .A1(n11268), .A2(n11269), .ZN(n11187) );
  NAND3_X1 U11096 ( .A1(a_12_), .A2(n11270), .A3(b_21_), .ZN(n11269) );
  OR2_X1 U11097 ( .A1(n11183), .A2(n11181), .ZN(n11270) );
  NAND2_X1 U11098 ( .A1(n11181), .A2(n11183), .ZN(n11268) );
  NAND2_X1 U11099 ( .A1(n11271), .A2(n11272), .ZN(n11183) );
  NAND2_X1 U11100 ( .A1(n11180), .A2(n11273), .ZN(n11272) );
  OR2_X1 U11101 ( .A1(n11179), .A2(n11178), .ZN(n11273) );
  NOR2_X1 U11102 ( .A1(n8749), .A2(n8310), .ZN(n11180) );
  NAND2_X1 U11103 ( .A1(n11178), .A2(n11179), .ZN(n11271) );
  NAND2_X1 U11104 ( .A1(n11274), .A2(n11275), .ZN(n11179) );
  NAND3_X1 U11105 ( .A1(a_14_), .A2(n11276), .A3(b_21_), .ZN(n11275) );
  NAND2_X1 U11106 ( .A1(n11175), .A2(n11174), .ZN(n11276) );
  OR2_X1 U11107 ( .A1(n11174), .A2(n11175), .ZN(n11274) );
  AND2_X1 U11108 ( .A1(n11277), .A2(n11278), .ZN(n11175) );
  NAND2_X1 U11109 ( .A1(n11172), .A2(n11279), .ZN(n11278) );
  OR2_X1 U11110 ( .A1(n11171), .A2(n11170), .ZN(n11279) );
  NOR2_X1 U11111 ( .A1(n8749), .A2(n8276), .ZN(n11172) );
  NAND2_X1 U11112 ( .A1(n11170), .A2(n11171), .ZN(n11277) );
  NAND2_X1 U11113 ( .A1(n11280), .A2(n11281), .ZN(n11171) );
  NAND3_X1 U11114 ( .A1(a_16_), .A2(n11282), .A3(b_21_), .ZN(n11281) );
  NAND2_X1 U11115 ( .A1(n11167), .A2(n11166), .ZN(n11282) );
  OR2_X1 U11116 ( .A1(n11166), .A2(n11167), .ZN(n11280) );
  AND2_X1 U11117 ( .A1(n11283), .A2(n11284), .ZN(n11167) );
  NAND2_X1 U11118 ( .A1(n11164), .A2(n11285), .ZN(n11284) );
  OR2_X1 U11119 ( .A1(n11163), .A2(n11161), .ZN(n11285) );
  NOR2_X1 U11120 ( .A1(n8749), .A2(n8210), .ZN(n11164) );
  NAND2_X1 U11121 ( .A1(n11161), .A2(n11163), .ZN(n11283) );
  NAND2_X1 U11122 ( .A1(n11286), .A2(n11287), .ZN(n11163) );
  NAND3_X1 U11123 ( .A1(a_18_), .A2(n11288), .A3(b_21_), .ZN(n11287) );
  NAND2_X1 U11124 ( .A1(n11159), .A2(n11158), .ZN(n11288) );
  OR2_X1 U11125 ( .A1(n11158), .A2(n11159), .ZN(n11286) );
  AND2_X1 U11126 ( .A1(n11289), .A2(n11290), .ZN(n11159) );
  NAND2_X1 U11127 ( .A1(n11156), .A2(n11291), .ZN(n11290) );
  OR2_X1 U11128 ( .A1(n11155), .A2(n11153), .ZN(n11291) );
  NOR2_X1 U11129 ( .A1(n8749), .A2(n8170), .ZN(n11156) );
  NAND2_X1 U11130 ( .A1(n11153), .A2(n11155), .ZN(n11289) );
  NAND2_X1 U11131 ( .A1(n11292), .A2(n11293), .ZN(n11155) );
  NAND3_X1 U11132 ( .A1(a_20_), .A2(n11294), .A3(b_21_), .ZN(n11293) );
  NAND2_X1 U11133 ( .A1(n11151), .A2(n11150), .ZN(n11294) );
  OR2_X1 U11134 ( .A1(n11150), .A2(n11151), .ZN(n11292) );
  AND2_X1 U11135 ( .A1(n11295), .A2(n11296), .ZN(n11151) );
  NAND2_X1 U11136 ( .A1(n11148), .A2(n11297), .ZN(n11296) );
  OR2_X1 U11137 ( .A1(n11147), .A2(n11146), .ZN(n11297) );
  INV_X1 U11138 ( .A(n8119), .ZN(n11148) );
  NAND2_X1 U11139 ( .A1(b_21_), .A2(a_21_), .ZN(n8119) );
  NAND2_X1 U11140 ( .A1(n11146), .A2(n11147), .ZN(n11295) );
  NAND2_X1 U11141 ( .A1(n11298), .A2(n11299), .ZN(n11147) );
  NAND3_X1 U11142 ( .A1(a_22_), .A2(n11300), .A3(b_21_), .ZN(n11299) );
  OR2_X1 U11143 ( .A1(n11143), .A2(n11141), .ZN(n11300) );
  NAND2_X1 U11144 ( .A1(n11141), .A2(n11143), .ZN(n11298) );
  NAND2_X1 U11145 ( .A1(n11301), .A2(n11302), .ZN(n11143) );
  NAND2_X1 U11146 ( .A1(n11087), .A2(n11303), .ZN(n11302) );
  OR2_X1 U11147 ( .A1(n11086), .A2(n11084), .ZN(n11303) );
  NOR2_X1 U11148 ( .A1(n8749), .A2(n8747), .ZN(n11087) );
  NAND2_X1 U11149 ( .A1(n11084), .A2(n11086), .ZN(n11301) );
  NAND2_X1 U11150 ( .A1(n11304), .A2(n11305), .ZN(n11086) );
  NAND3_X1 U11151 ( .A1(a_24_), .A2(n11306), .A3(b_21_), .ZN(n11305) );
  NAND2_X1 U11152 ( .A1(n11139), .A2(n11138), .ZN(n11306) );
  OR2_X1 U11153 ( .A1(n11138), .A2(n11139), .ZN(n11304) );
  AND2_X1 U11154 ( .A1(n11307), .A2(n11308), .ZN(n11139) );
  NAND2_X1 U11155 ( .A1(n11136), .A2(n11309), .ZN(n11308) );
  OR2_X1 U11156 ( .A1(n11135), .A2(n11134), .ZN(n11309) );
  NOR2_X1 U11157 ( .A1(n8749), .A2(n8744), .ZN(n11136) );
  NAND2_X1 U11158 ( .A1(n11134), .A2(n11135), .ZN(n11307) );
  NAND2_X1 U11159 ( .A1(n11131), .A2(n11310), .ZN(n11135) );
  NAND2_X1 U11160 ( .A1(n11130), .A2(n11132), .ZN(n11310) );
  NAND2_X1 U11161 ( .A1(n11311), .A2(n11312), .ZN(n11132) );
  NAND2_X1 U11162 ( .A1(b_21_), .A2(a_26_), .ZN(n11312) );
  INV_X1 U11163 ( .A(n11313), .ZN(n11311) );
  XNOR2_X1 U11164 ( .A(n11314), .B(n11315), .ZN(n11130) );
  NAND2_X1 U11165 ( .A1(n11316), .A2(n11317), .ZN(n11314) );
  NAND2_X1 U11166 ( .A1(a_26_), .A2(n11313), .ZN(n11131) );
  NAND2_X1 U11167 ( .A1(n11103), .A2(n11318), .ZN(n11313) );
  NAND2_X1 U11168 ( .A1(n11102), .A2(n11104), .ZN(n11318) );
  NAND2_X1 U11169 ( .A1(n11319), .A2(n11320), .ZN(n11104) );
  NAND2_X1 U11170 ( .A1(b_21_), .A2(a_27_), .ZN(n11320) );
  INV_X1 U11171 ( .A(n11321), .ZN(n11319) );
  XNOR2_X1 U11172 ( .A(n11322), .B(n11323), .ZN(n11102) );
  XOR2_X1 U11173 ( .A(n11324), .B(n11325), .Z(n11322) );
  NAND2_X1 U11174 ( .A1(b_20_), .A2(a_28_), .ZN(n11324) );
  NAND2_X1 U11175 ( .A1(a_27_), .A2(n11321), .ZN(n11103) );
  NAND2_X1 U11176 ( .A1(n11326), .A2(n11327), .ZN(n11321) );
  NAND3_X1 U11177 ( .A1(a_28_), .A2(n11328), .A3(b_21_), .ZN(n11327) );
  NAND2_X1 U11178 ( .A1(n11112), .A2(n11110), .ZN(n11328) );
  OR2_X1 U11179 ( .A1(n11110), .A2(n11112), .ZN(n11326) );
  AND2_X1 U11180 ( .A1(n11329), .A2(n11330), .ZN(n11112) );
  NAND2_X1 U11181 ( .A1(n11126), .A2(n11331), .ZN(n11330) );
  OR2_X1 U11182 ( .A1(n11127), .A2(n11128), .ZN(n11331) );
  NOR2_X1 U11183 ( .A1(n8749), .A2(n7890), .ZN(n11126) );
  NAND2_X1 U11184 ( .A1(n11128), .A2(n11127), .ZN(n11329) );
  NAND2_X1 U11185 ( .A1(n11332), .A2(n11333), .ZN(n11127) );
  NAND2_X1 U11186 ( .A1(b_19_), .A2(n11334), .ZN(n11333) );
  NAND2_X1 U11187 ( .A1(n7864), .A2(n11335), .ZN(n11334) );
  NAND2_X1 U11188 ( .A1(a_31_), .A2(n8145), .ZN(n11335) );
  NAND2_X1 U11189 ( .A1(b_20_), .A2(n11336), .ZN(n11332) );
  NAND2_X1 U11190 ( .A1(n9137), .A2(n11337), .ZN(n11336) );
  NAND2_X1 U11191 ( .A1(a_30_), .A2(n8752), .ZN(n11337) );
  AND3_X1 U11192 ( .A1(b_20_), .A2(b_21_), .A3(n7818), .ZN(n11128) );
  XNOR2_X1 U11193 ( .A(n11338), .B(n11339), .ZN(n11110) );
  XOR2_X1 U11194 ( .A(n11340), .B(n11341), .Z(n11338) );
  XNOR2_X1 U11195 ( .A(n11342), .B(n11343), .ZN(n11134) );
  NAND2_X1 U11196 ( .A1(n11344), .A2(n11345), .ZN(n11342) );
  XNOR2_X1 U11197 ( .A(n11346), .B(n11347), .ZN(n11138) );
  XOR2_X1 U11198 ( .A(n11348), .B(n11349), .Z(n11346) );
  XNOR2_X1 U11199 ( .A(n11350), .B(n11351), .ZN(n11084) );
  XNOR2_X1 U11200 ( .A(n11352), .B(n11353), .ZN(n11350) );
  NOR2_X1 U11201 ( .A1(n8745), .A2(n8145), .ZN(n11353) );
  XNOR2_X1 U11202 ( .A(n11354), .B(n11355), .ZN(n11141) );
  XNOR2_X1 U11203 ( .A(n11356), .B(n11357), .ZN(n11355) );
  XNOR2_X1 U11204 ( .A(n11358), .B(n11359), .ZN(n11146) );
  XOR2_X1 U11205 ( .A(n11360), .B(n11361), .Z(n11359) );
  NAND2_X1 U11206 ( .A1(b_20_), .A2(a_22_), .ZN(n11361) );
  XNOR2_X1 U11207 ( .A(n11362), .B(n11363), .ZN(n11150) );
  XOR2_X1 U11208 ( .A(n11364), .B(n11365), .Z(n11362) );
  XOR2_X1 U11209 ( .A(n11366), .B(n11367), .Z(n11153) );
  XOR2_X1 U11210 ( .A(n11368), .B(n11369), .Z(n11366) );
  XNOR2_X1 U11211 ( .A(n11370), .B(n11371), .ZN(n11158) );
  XOR2_X1 U11212 ( .A(n11372), .B(n11373), .Z(n11370) );
  XNOR2_X1 U11213 ( .A(n11374), .B(n11375), .ZN(n11161) );
  XNOR2_X1 U11214 ( .A(n11376), .B(n11377), .ZN(n11374) );
  NOR2_X1 U11215 ( .A1(n8753), .A2(n8145), .ZN(n11377) );
  XOR2_X1 U11216 ( .A(n11378), .B(n11379), .Z(n11166) );
  XNOR2_X1 U11217 ( .A(n11380), .B(n11381), .ZN(n11379) );
  XNOR2_X1 U11218 ( .A(n11382), .B(n11383), .ZN(n11170) );
  XNOR2_X1 U11219 ( .A(n11384), .B(n11385), .ZN(n11382) );
  NOR2_X1 U11220 ( .A1(n8755), .A2(n8145), .ZN(n11385) );
  XOR2_X1 U11221 ( .A(n11386), .B(n11387), .Z(n11174) );
  XNOR2_X1 U11222 ( .A(n11388), .B(n11389), .ZN(n11387) );
  XNOR2_X1 U11223 ( .A(n11390), .B(n11391), .ZN(n11178) );
  XNOR2_X1 U11224 ( .A(n11392), .B(n11393), .ZN(n11390) );
  NOR2_X1 U11225 ( .A1(n8757), .A2(n8145), .ZN(n11393) );
  XNOR2_X1 U11226 ( .A(n11394), .B(n11395), .ZN(n11181) );
  XNOR2_X1 U11227 ( .A(n11396), .B(n11397), .ZN(n11395) );
  XNOR2_X1 U11228 ( .A(n11398), .B(n11399), .ZN(n11185) );
  XOR2_X1 U11229 ( .A(n11400), .B(n11401), .Z(n11399) );
  NAND2_X1 U11230 ( .A1(b_20_), .A2(a_12_), .ZN(n11401) );
  XNOR2_X1 U11231 ( .A(n11402), .B(n11403), .ZN(n11190) );
  XOR2_X1 U11232 ( .A(n11404), .B(n11405), .Z(n11403) );
  NAND2_X1 U11233 ( .A1(b_20_), .A2(a_11_), .ZN(n11405) );
  XNOR2_X1 U11234 ( .A(n11406), .B(n11407), .ZN(n11194) );
  XOR2_X1 U11235 ( .A(n11408), .B(n11409), .Z(n11406) );
  XOR2_X1 U11236 ( .A(n11410), .B(n11411), .Z(n11197) );
  XOR2_X1 U11237 ( .A(n11412), .B(n11413), .Z(n11410) );
  XNOR2_X1 U11238 ( .A(n11414), .B(n11415), .ZN(n11201) );
  XNOR2_X1 U11239 ( .A(n11416), .B(n11417), .ZN(n11414) );
  NOR2_X1 U11240 ( .A1(n8763), .A2(n8145), .ZN(n11417) );
  XNOR2_X1 U11241 ( .A(n11418), .B(n11419), .ZN(n11205) );
  NAND2_X1 U11242 ( .A1(n11420), .A2(n11421), .ZN(n11418) );
  XOR2_X1 U11243 ( .A(n11422), .B(n11423), .Z(n11210) );
  NAND2_X1 U11244 ( .A1(n11424), .A2(n11425), .ZN(n11422) );
  XNOR2_X1 U11245 ( .A(n11426), .B(n11427), .ZN(n11213) );
  XNOR2_X1 U11246 ( .A(n11428), .B(n11429), .ZN(n11427) );
  XNOR2_X1 U11247 ( .A(n11430), .B(n11431), .ZN(n11217) );
  XOR2_X1 U11248 ( .A(n11432), .B(n11433), .Z(n11431) );
  NAND2_X1 U11249 ( .A1(b_20_), .A2(a_4_), .ZN(n11433) );
  XNOR2_X1 U11250 ( .A(n11434), .B(n11435), .ZN(n11221) );
  NAND2_X1 U11251 ( .A1(n11436), .A2(n11437), .ZN(n11434) );
  XNOR2_X1 U11252 ( .A(n11438), .B(n11439), .ZN(n11015) );
  XNOR2_X1 U11253 ( .A(n11440), .B(n11441), .ZN(n11438) );
  XOR2_X1 U11254 ( .A(n11442), .B(n11443), .Z(n11227) );
  XOR2_X1 U11255 ( .A(n11444), .B(n11445), .Z(n11442) );
  XOR2_X1 U11256 ( .A(n11446), .B(n11447), .Z(n11226) );
  XNOR2_X1 U11257 ( .A(n11448), .B(n11449), .ZN(n11446) );
  NOR2_X1 U11258 ( .A1(n9674), .A2(n8145), .ZN(n11449) );
  XOR2_X1 U11259 ( .A(n8969), .B(n8968), .Z(n11231) );
  NAND3_X1 U11260 ( .A1(n8968), .A2(n8969), .A3(n11450), .ZN(n8858) );
  XOR2_X1 U11261 ( .A(n8962), .B(n8961), .Z(n11450) );
  NAND2_X1 U11262 ( .A1(n11451), .A2(n11452), .ZN(n8969) );
  NAND3_X1 U11263 ( .A1(a_0_), .A2(n11453), .A3(b_20_), .ZN(n11452) );
  NAND2_X1 U11264 ( .A1(n11448), .A2(n11447), .ZN(n11453) );
  OR2_X1 U11265 ( .A1(n11447), .A2(n11448), .ZN(n11451) );
  AND2_X1 U11266 ( .A1(n11454), .A2(n11455), .ZN(n11448) );
  NAND2_X1 U11267 ( .A1(n11445), .A2(n11456), .ZN(n11455) );
  OR2_X1 U11268 ( .A1(n11444), .A2(n11443), .ZN(n11456) );
  NOR2_X1 U11269 ( .A1(n8145), .A2(n8617), .ZN(n11445) );
  NAND2_X1 U11270 ( .A1(n11443), .A2(n11444), .ZN(n11454) );
  NAND2_X1 U11271 ( .A1(n11457), .A2(n11458), .ZN(n11444) );
  NAND2_X1 U11272 ( .A1(n11441), .A2(n11459), .ZN(n11458) );
  NAND2_X1 U11273 ( .A1(n11440), .A2(n11439), .ZN(n11459) );
  NOR2_X1 U11274 ( .A1(n8145), .A2(n8768), .ZN(n11441) );
  OR2_X1 U11275 ( .A1(n11439), .A2(n11440), .ZN(n11457) );
  AND2_X1 U11276 ( .A1(n11436), .A2(n11460), .ZN(n11440) );
  NAND2_X1 U11277 ( .A1(n11435), .A2(n11437), .ZN(n11460) );
  NAND2_X1 U11278 ( .A1(n11461), .A2(n11462), .ZN(n11437) );
  NAND2_X1 U11279 ( .A1(b_20_), .A2(a_3_), .ZN(n11462) );
  INV_X1 U11280 ( .A(n11463), .ZN(n11461) );
  XOR2_X1 U11281 ( .A(n11464), .B(n11465), .Z(n11435) );
  XOR2_X1 U11282 ( .A(n11466), .B(n11467), .Z(n11464) );
  NOR2_X1 U11283 ( .A1(n8766), .A2(n8752), .ZN(n11467) );
  NAND2_X1 U11284 ( .A1(a_3_), .A2(n11463), .ZN(n11436) );
  NAND2_X1 U11285 ( .A1(n11468), .A2(n11469), .ZN(n11463) );
  NAND3_X1 U11286 ( .A1(a_4_), .A2(n11470), .A3(b_20_), .ZN(n11469) );
  OR2_X1 U11287 ( .A1(n11432), .A2(n11430), .ZN(n11470) );
  NAND2_X1 U11288 ( .A1(n11430), .A2(n11432), .ZN(n11468) );
  NAND2_X1 U11289 ( .A1(n11471), .A2(n11472), .ZN(n11432) );
  NAND2_X1 U11290 ( .A1(n11429), .A2(n11473), .ZN(n11472) );
  OR2_X1 U11291 ( .A1(n11428), .A2(n11426), .ZN(n11473) );
  NOR2_X1 U11292 ( .A1(n8145), .A2(n8517), .ZN(n11429) );
  NAND2_X1 U11293 ( .A1(n11426), .A2(n11428), .ZN(n11471) );
  NAND2_X1 U11294 ( .A1(n11424), .A2(n11474), .ZN(n11428) );
  NAND2_X1 U11295 ( .A1(n11423), .A2(n11425), .ZN(n11474) );
  NAND2_X1 U11296 ( .A1(n11475), .A2(n11476), .ZN(n11425) );
  NAND2_X1 U11297 ( .A1(b_20_), .A2(a_6_), .ZN(n11476) );
  INV_X1 U11298 ( .A(n11477), .ZN(n11475) );
  XNOR2_X1 U11299 ( .A(n11478), .B(n11479), .ZN(n11423) );
  XOR2_X1 U11300 ( .A(n11480), .B(n11481), .Z(n11479) );
  NAND2_X1 U11301 ( .A1(b_19_), .A2(a_7_), .ZN(n11481) );
  NAND2_X1 U11302 ( .A1(a_6_), .A2(n11477), .ZN(n11424) );
  NAND2_X1 U11303 ( .A1(n11420), .A2(n11482), .ZN(n11477) );
  NAND2_X1 U11304 ( .A1(n11419), .A2(n11421), .ZN(n11482) );
  NAND2_X1 U11305 ( .A1(n11483), .A2(n11484), .ZN(n11421) );
  NAND2_X1 U11306 ( .A1(b_20_), .A2(a_7_), .ZN(n11484) );
  INV_X1 U11307 ( .A(n11485), .ZN(n11483) );
  XOR2_X1 U11308 ( .A(n11486), .B(n11487), .Z(n11419) );
  XOR2_X1 U11309 ( .A(n11488), .B(n11489), .Z(n11486) );
  NOR2_X1 U11310 ( .A1(n8763), .A2(n8752), .ZN(n11489) );
  NAND2_X1 U11311 ( .A1(a_7_), .A2(n11485), .ZN(n11420) );
  NAND2_X1 U11312 ( .A1(n11490), .A2(n11491), .ZN(n11485) );
  NAND3_X1 U11313 ( .A1(a_8_), .A2(n11492), .A3(b_20_), .ZN(n11491) );
  NAND2_X1 U11314 ( .A1(n11416), .A2(n11415), .ZN(n11492) );
  OR2_X1 U11315 ( .A1(n11415), .A2(n11416), .ZN(n11490) );
  AND2_X1 U11316 ( .A1(n11493), .A2(n11494), .ZN(n11416) );
  NAND2_X1 U11317 ( .A1(n11413), .A2(n11495), .ZN(n11494) );
  OR2_X1 U11318 ( .A1(n11412), .A2(n11411), .ZN(n11495) );
  NOR2_X1 U11319 ( .A1(n8145), .A2(n8426), .ZN(n11413) );
  NAND2_X1 U11320 ( .A1(n11411), .A2(n11412), .ZN(n11493) );
  NAND2_X1 U11321 ( .A1(n11496), .A2(n11497), .ZN(n11412) );
  NAND2_X1 U11322 ( .A1(n11409), .A2(n11498), .ZN(n11497) );
  OR2_X1 U11323 ( .A1(n11408), .A2(n11407), .ZN(n11498) );
  NOR2_X1 U11324 ( .A1(n8145), .A2(n8761), .ZN(n11409) );
  NAND2_X1 U11325 ( .A1(n11407), .A2(n11408), .ZN(n11496) );
  NAND2_X1 U11326 ( .A1(n11499), .A2(n11500), .ZN(n11408) );
  NAND3_X1 U11327 ( .A1(a_11_), .A2(n11501), .A3(b_20_), .ZN(n11500) );
  OR2_X1 U11328 ( .A1(n11404), .A2(n11402), .ZN(n11501) );
  NAND2_X1 U11329 ( .A1(n11402), .A2(n11404), .ZN(n11499) );
  NAND2_X1 U11330 ( .A1(n11502), .A2(n11503), .ZN(n11404) );
  NAND3_X1 U11331 ( .A1(a_12_), .A2(n11504), .A3(b_20_), .ZN(n11503) );
  OR2_X1 U11332 ( .A1(n11400), .A2(n11398), .ZN(n11504) );
  NAND2_X1 U11333 ( .A1(n11398), .A2(n11400), .ZN(n11502) );
  NAND2_X1 U11334 ( .A1(n11505), .A2(n11506), .ZN(n11400) );
  NAND2_X1 U11335 ( .A1(n11397), .A2(n11507), .ZN(n11506) );
  OR2_X1 U11336 ( .A1(n11396), .A2(n11394), .ZN(n11507) );
  NOR2_X1 U11337 ( .A1(n8145), .A2(n8310), .ZN(n11397) );
  NAND2_X1 U11338 ( .A1(n11394), .A2(n11396), .ZN(n11505) );
  NAND2_X1 U11339 ( .A1(n11508), .A2(n11509), .ZN(n11396) );
  NAND3_X1 U11340 ( .A1(a_14_), .A2(n11510), .A3(b_20_), .ZN(n11509) );
  NAND2_X1 U11341 ( .A1(n11392), .A2(n11391), .ZN(n11510) );
  OR2_X1 U11342 ( .A1(n11391), .A2(n11392), .ZN(n11508) );
  AND2_X1 U11343 ( .A1(n11511), .A2(n11512), .ZN(n11392) );
  NAND2_X1 U11344 ( .A1(n11389), .A2(n11513), .ZN(n11512) );
  OR2_X1 U11345 ( .A1(n11388), .A2(n11386), .ZN(n11513) );
  NOR2_X1 U11346 ( .A1(n8145), .A2(n8276), .ZN(n11389) );
  NAND2_X1 U11347 ( .A1(n11386), .A2(n11388), .ZN(n11511) );
  NAND2_X1 U11348 ( .A1(n11514), .A2(n11515), .ZN(n11388) );
  NAND3_X1 U11349 ( .A1(a_16_), .A2(n11516), .A3(b_20_), .ZN(n11515) );
  NAND2_X1 U11350 ( .A1(n11384), .A2(n11383), .ZN(n11516) );
  OR2_X1 U11351 ( .A1(n11383), .A2(n11384), .ZN(n11514) );
  AND2_X1 U11352 ( .A1(n11517), .A2(n11518), .ZN(n11384) );
  NAND2_X1 U11353 ( .A1(n11381), .A2(n11519), .ZN(n11518) );
  OR2_X1 U11354 ( .A1(n11380), .A2(n11378), .ZN(n11519) );
  NOR2_X1 U11355 ( .A1(n8145), .A2(n8210), .ZN(n11381) );
  NAND2_X1 U11356 ( .A1(n11378), .A2(n11380), .ZN(n11517) );
  NAND2_X1 U11357 ( .A1(n11520), .A2(n11521), .ZN(n11380) );
  NAND3_X1 U11358 ( .A1(a_18_), .A2(n11522), .A3(b_20_), .ZN(n11521) );
  NAND2_X1 U11359 ( .A1(n11376), .A2(n11375), .ZN(n11522) );
  OR2_X1 U11360 ( .A1(n11375), .A2(n11376), .ZN(n11520) );
  AND2_X1 U11361 ( .A1(n11523), .A2(n11524), .ZN(n11376) );
  NAND2_X1 U11362 ( .A1(n11373), .A2(n11525), .ZN(n11524) );
  OR2_X1 U11363 ( .A1(n11372), .A2(n11371), .ZN(n11525) );
  NOR2_X1 U11364 ( .A1(n8145), .A2(n8170), .ZN(n11373) );
  NAND2_X1 U11365 ( .A1(n11371), .A2(n11372), .ZN(n11523) );
  NAND2_X1 U11366 ( .A1(n11526), .A2(n11527), .ZN(n11372) );
  NAND2_X1 U11367 ( .A1(n11367), .A2(n11528), .ZN(n11527) );
  OR2_X1 U11368 ( .A1(n11368), .A2(n11369), .ZN(n11528) );
  XNOR2_X1 U11369 ( .A(n11529), .B(n11530), .ZN(n11367) );
  XNOR2_X1 U11370 ( .A(n11531), .B(n11532), .ZN(n11529) );
  NAND2_X1 U11371 ( .A1(n11369), .A2(n11368), .ZN(n11526) );
  NAND2_X1 U11372 ( .A1(n11533), .A2(n11534), .ZN(n11368) );
  NAND2_X1 U11373 ( .A1(n11365), .A2(n11535), .ZN(n11534) );
  OR2_X1 U11374 ( .A1(n11364), .A2(n11363), .ZN(n11535) );
  NOR2_X1 U11375 ( .A1(n8145), .A2(n8750), .ZN(n11365) );
  NAND2_X1 U11376 ( .A1(n11363), .A2(n11364), .ZN(n11533) );
  NAND2_X1 U11377 ( .A1(n11536), .A2(n11537), .ZN(n11364) );
  NAND3_X1 U11378 ( .A1(a_22_), .A2(n11538), .A3(b_20_), .ZN(n11537) );
  OR2_X1 U11379 ( .A1(n11360), .A2(n11358), .ZN(n11538) );
  NAND2_X1 U11380 ( .A1(n11358), .A2(n11360), .ZN(n11536) );
  NAND2_X1 U11381 ( .A1(n11539), .A2(n11540), .ZN(n11360) );
  NAND2_X1 U11382 ( .A1(n11357), .A2(n11541), .ZN(n11540) );
  OR2_X1 U11383 ( .A1(n11356), .A2(n11354), .ZN(n11541) );
  NOR2_X1 U11384 ( .A1(n8145), .A2(n8747), .ZN(n11357) );
  NAND2_X1 U11385 ( .A1(n11354), .A2(n11356), .ZN(n11539) );
  NAND2_X1 U11386 ( .A1(n11542), .A2(n11543), .ZN(n11356) );
  NAND3_X1 U11387 ( .A1(a_24_), .A2(n11544), .A3(b_20_), .ZN(n11543) );
  NAND2_X1 U11388 ( .A1(n11352), .A2(n11351), .ZN(n11544) );
  OR2_X1 U11389 ( .A1(n11351), .A2(n11352), .ZN(n11542) );
  AND2_X1 U11390 ( .A1(n11545), .A2(n11546), .ZN(n11352) );
  NAND2_X1 U11391 ( .A1(n11349), .A2(n11547), .ZN(n11546) );
  OR2_X1 U11392 ( .A1(n11348), .A2(n11347), .ZN(n11547) );
  NOR2_X1 U11393 ( .A1(n8145), .A2(n8744), .ZN(n11349) );
  NAND2_X1 U11394 ( .A1(n11347), .A2(n11348), .ZN(n11545) );
  NAND2_X1 U11395 ( .A1(n11344), .A2(n11548), .ZN(n11348) );
  NAND2_X1 U11396 ( .A1(n11343), .A2(n11345), .ZN(n11548) );
  NAND2_X1 U11397 ( .A1(n11549), .A2(n11550), .ZN(n11345) );
  NAND2_X1 U11398 ( .A1(b_20_), .A2(a_26_), .ZN(n11550) );
  INV_X1 U11399 ( .A(n11551), .ZN(n11549) );
  XNOR2_X1 U11400 ( .A(n11552), .B(n11553), .ZN(n11343) );
  NAND2_X1 U11401 ( .A1(n11554), .A2(n11555), .ZN(n11552) );
  NAND2_X1 U11402 ( .A1(a_26_), .A2(n11551), .ZN(n11344) );
  NAND2_X1 U11403 ( .A1(n11316), .A2(n11556), .ZN(n11551) );
  NAND2_X1 U11404 ( .A1(n11315), .A2(n11317), .ZN(n11556) );
  NAND2_X1 U11405 ( .A1(n11557), .A2(n11558), .ZN(n11317) );
  NAND2_X1 U11406 ( .A1(b_20_), .A2(a_27_), .ZN(n11558) );
  INV_X1 U11407 ( .A(n11559), .ZN(n11557) );
  XNOR2_X1 U11408 ( .A(n11560), .B(n11561), .ZN(n11315) );
  XOR2_X1 U11409 ( .A(n11562), .B(n11563), .Z(n11560) );
  NAND2_X1 U11410 ( .A1(b_19_), .A2(a_28_), .ZN(n11562) );
  NAND2_X1 U11411 ( .A1(a_27_), .A2(n11559), .ZN(n11316) );
  NAND2_X1 U11412 ( .A1(n11564), .A2(n11565), .ZN(n11559) );
  NAND3_X1 U11413 ( .A1(a_28_), .A2(n11566), .A3(b_20_), .ZN(n11565) );
  NAND2_X1 U11414 ( .A1(n11325), .A2(n11323), .ZN(n11566) );
  OR2_X1 U11415 ( .A1(n11323), .A2(n11325), .ZN(n11564) );
  AND2_X1 U11416 ( .A1(n11567), .A2(n11568), .ZN(n11325) );
  NAND2_X1 U11417 ( .A1(n11339), .A2(n11569), .ZN(n11568) );
  OR2_X1 U11418 ( .A1(n11340), .A2(n11341), .ZN(n11569) );
  NOR2_X1 U11419 ( .A1(n8145), .A2(n7890), .ZN(n11339) );
  NAND2_X1 U11420 ( .A1(n11341), .A2(n11340), .ZN(n11567) );
  NAND2_X1 U11421 ( .A1(n11570), .A2(n11571), .ZN(n11340) );
  NAND2_X1 U11422 ( .A1(b_18_), .A2(n11572), .ZN(n11571) );
  NAND2_X1 U11423 ( .A1(n7864), .A2(n11573), .ZN(n11572) );
  NAND2_X1 U11424 ( .A1(a_31_), .A2(n8752), .ZN(n11573) );
  NAND2_X1 U11425 ( .A1(b_19_), .A2(n11574), .ZN(n11570) );
  NAND2_X1 U11426 ( .A1(n9137), .A2(n11575), .ZN(n11574) );
  NAND2_X1 U11427 ( .A1(a_30_), .A2(n8195), .ZN(n11575) );
  AND3_X1 U11428 ( .A1(b_19_), .A2(b_20_), .A3(n7818), .ZN(n11341) );
  XNOR2_X1 U11429 ( .A(n11576), .B(n11577), .ZN(n11323) );
  XOR2_X1 U11430 ( .A(n11578), .B(n11579), .Z(n11576) );
  XNOR2_X1 U11431 ( .A(n11580), .B(n11581), .ZN(n11347) );
  NAND2_X1 U11432 ( .A1(n11582), .A2(n11583), .ZN(n11580) );
  XNOR2_X1 U11433 ( .A(n11584), .B(n11585), .ZN(n11351) );
  XOR2_X1 U11434 ( .A(n11586), .B(n11587), .Z(n11584) );
  XNOR2_X1 U11435 ( .A(n11588), .B(n11589), .ZN(n11354) );
  XNOR2_X1 U11436 ( .A(n11590), .B(n11591), .ZN(n11588) );
  NOR2_X1 U11437 ( .A1(n8745), .A2(n8752), .ZN(n11591) );
  XNOR2_X1 U11438 ( .A(n11592), .B(n11593), .ZN(n11358) );
  XNOR2_X1 U11439 ( .A(n11594), .B(n11595), .ZN(n11593) );
  XNOR2_X1 U11440 ( .A(n11596), .B(n11597), .ZN(n11363) );
  XOR2_X1 U11441 ( .A(n11598), .B(n11599), .Z(n11597) );
  NAND2_X1 U11442 ( .A1(b_19_), .A2(a_22_), .ZN(n11599) );
  INV_X1 U11443 ( .A(n8715), .ZN(n11369) );
  NAND2_X1 U11444 ( .A1(b_20_), .A2(a_20_), .ZN(n8715) );
  XNOR2_X1 U11445 ( .A(n11600), .B(n11601), .ZN(n11371) );
  XOR2_X1 U11446 ( .A(n11602), .B(n11603), .Z(n11600) );
  NAND2_X1 U11447 ( .A1(b_19_), .A2(a_20_), .ZN(n11602) );
  XNOR2_X1 U11448 ( .A(n11604), .B(n11605), .ZN(n11375) );
  XOR2_X1 U11449 ( .A(n11606), .B(n11607), .Z(n11604) );
  XNOR2_X1 U11450 ( .A(n11608), .B(n11609), .ZN(n11378) );
  XNOR2_X1 U11451 ( .A(n11610), .B(n11611), .ZN(n11608) );
  NOR2_X1 U11452 ( .A1(n8753), .A2(n8752), .ZN(n11611) );
  XNOR2_X1 U11453 ( .A(n11612), .B(n11613), .ZN(n11383) );
  XOR2_X1 U11454 ( .A(n11614), .B(n11615), .Z(n11612) );
  XNOR2_X1 U11455 ( .A(n11616), .B(n11617), .ZN(n11386) );
  XOR2_X1 U11456 ( .A(n11618), .B(n11619), .Z(n11617) );
  NAND2_X1 U11457 ( .A1(b_19_), .A2(a_16_), .ZN(n11619) );
  XOR2_X1 U11458 ( .A(n11620), .B(n11621), .Z(n11391) );
  XNOR2_X1 U11459 ( .A(n11622), .B(n11623), .ZN(n11621) );
  XNOR2_X1 U11460 ( .A(n11624), .B(n11625), .ZN(n11394) );
  XNOR2_X1 U11461 ( .A(n11626), .B(n11627), .ZN(n11624) );
  NOR2_X1 U11462 ( .A1(n8757), .A2(n8752), .ZN(n11627) );
  XOR2_X1 U11463 ( .A(n11628), .B(n11629), .Z(n11398) );
  XOR2_X1 U11464 ( .A(n11630), .B(n11631), .Z(n11628) );
  XNOR2_X1 U11465 ( .A(n11632), .B(n11633), .ZN(n11402) );
  XNOR2_X1 U11466 ( .A(n11634), .B(n11635), .ZN(n11633) );
  XNOR2_X1 U11467 ( .A(n11636), .B(n11637), .ZN(n11407) );
  XOR2_X1 U11468 ( .A(n11638), .B(n11639), .Z(n11637) );
  NAND2_X1 U11469 ( .A1(b_19_), .A2(a_11_), .ZN(n11639) );
  XNOR2_X1 U11470 ( .A(n11640), .B(n11641), .ZN(n11411) );
  NAND2_X1 U11471 ( .A1(n11642), .A2(n11643), .ZN(n11640) );
  XOR2_X1 U11472 ( .A(n11644), .B(n11645), .Z(n11415) );
  XOR2_X1 U11473 ( .A(n11646), .B(n11647), .Z(n11645) );
  NAND2_X1 U11474 ( .A1(b_19_), .A2(a_9_), .ZN(n11647) );
  XNOR2_X1 U11475 ( .A(n11648), .B(n11649), .ZN(n11426) );
  XNOR2_X1 U11476 ( .A(n11650), .B(n11651), .ZN(n11648) );
  NOR2_X1 U11477 ( .A1(n8491), .A2(n8752), .ZN(n11651) );
  XNOR2_X1 U11478 ( .A(n11652), .B(n11653), .ZN(n11430) );
  XOR2_X1 U11479 ( .A(n11654), .B(n11655), .Z(n11653) );
  NAND2_X1 U11480 ( .A1(b_19_), .A2(a_5_), .ZN(n11655) );
  XOR2_X1 U11481 ( .A(n11656), .B(n11657), .Z(n11439) );
  XOR2_X1 U11482 ( .A(n11658), .B(n11659), .Z(n11657) );
  NAND2_X1 U11483 ( .A1(b_19_), .A2(a_3_), .ZN(n11659) );
  XNOR2_X1 U11484 ( .A(n11660), .B(n11661), .ZN(n11443) );
  XOR2_X1 U11485 ( .A(n11662), .B(n11663), .Z(n11661) );
  NAND2_X1 U11486 ( .A1(b_19_), .A2(a_2_), .ZN(n11663) );
  XOR2_X1 U11487 ( .A(n11664), .B(n11665), .Z(n11447) );
  XOR2_X1 U11488 ( .A(n11666), .B(n11667), .Z(n11665) );
  NAND2_X1 U11489 ( .A1(b_19_), .A2(a_1_), .ZN(n11667) );
  XNOR2_X1 U11490 ( .A(n11668), .B(n11669), .ZN(n8968) );
  XOR2_X1 U11491 ( .A(n11670), .B(n11671), .Z(n11669) );
  NAND2_X1 U11492 ( .A1(b_19_), .A2(a_0_), .ZN(n11671) );
  NAND3_X1 U11493 ( .A1(n11672), .A2(n8962), .A3(n8961), .ZN(n8863) );
  XNOR2_X1 U11494 ( .A(n11673), .B(n11674), .ZN(n8961) );
  XOR2_X1 U11495 ( .A(n11675), .B(n11676), .Z(n11674) );
  NAND2_X1 U11496 ( .A1(b_18_), .A2(a_0_), .ZN(n11676) );
  NAND2_X1 U11497 ( .A1(n11677), .A2(n11678), .ZN(n8962) );
  NAND3_X1 U11498 ( .A1(a_0_), .A2(n11679), .A3(b_19_), .ZN(n11678) );
  OR2_X1 U11499 ( .A1(n11670), .A2(n11668), .ZN(n11679) );
  NAND2_X1 U11500 ( .A1(n11668), .A2(n11670), .ZN(n11677) );
  NAND2_X1 U11501 ( .A1(n11680), .A2(n11681), .ZN(n11670) );
  NAND3_X1 U11502 ( .A1(a_1_), .A2(n11682), .A3(b_19_), .ZN(n11681) );
  OR2_X1 U11503 ( .A1(n11666), .A2(n11664), .ZN(n11682) );
  NAND2_X1 U11504 ( .A1(n11664), .A2(n11666), .ZN(n11680) );
  NAND2_X1 U11505 ( .A1(n11683), .A2(n11684), .ZN(n11666) );
  NAND3_X1 U11506 ( .A1(a_2_), .A2(n11685), .A3(b_19_), .ZN(n11684) );
  OR2_X1 U11507 ( .A1(n11662), .A2(n11660), .ZN(n11685) );
  NAND2_X1 U11508 ( .A1(n11660), .A2(n11662), .ZN(n11683) );
  NAND2_X1 U11509 ( .A1(n11686), .A2(n11687), .ZN(n11662) );
  NAND3_X1 U11510 ( .A1(a_3_), .A2(n11688), .A3(b_19_), .ZN(n11687) );
  OR2_X1 U11511 ( .A1(n11658), .A2(n11656), .ZN(n11688) );
  NAND2_X1 U11512 ( .A1(n11656), .A2(n11658), .ZN(n11686) );
  NAND2_X1 U11513 ( .A1(n11689), .A2(n11690), .ZN(n11658) );
  NAND3_X1 U11514 ( .A1(a_4_), .A2(n11691), .A3(b_19_), .ZN(n11690) );
  OR2_X1 U11515 ( .A1(n11466), .A2(n11465), .ZN(n11691) );
  NAND2_X1 U11516 ( .A1(n11465), .A2(n11466), .ZN(n11689) );
  NAND2_X1 U11517 ( .A1(n11692), .A2(n11693), .ZN(n11466) );
  NAND3_X1 U11518 ( .A1(a_5_), .A2(n11694), .A3(b_19_), .ZN(n11693) );
  OR2_X1 U11519 ( .A1(n11654), .A2(n11652), .ZN(n11694) );
  NAND2_X1 U11520 ( .A1(n11652), .A2(n11654), .ZN(n11692) );
  NAND2_X1 U11521 ( .A1(n11695), .A2(n11696), .ZN(n11654) );
  NAND3_X1 U11522 ( .A1(a_6_), .A2(n11697), .A3(b_19_), .ZN(n11696) );
  NAND2_X1 U11523 ( .A1(n11650), .A2(n11649), .ZN(n11697) );
  OR2_X1 U11524 ( .A1(n11649), .A2(n11650), .ZN(n11695) );
  AND2_X1 U11525 ( .A1(n11698), .A2(n11699), .ZN(n11650) );
  NAND3_X1 U11526 ( .A1(a_7_), .A2(n11700), .A3(b_19_), .ZN(n11699) );
  OR2_X1 U11527 ( .A1(n11480), .A2(n11478), .ZN(n11700) );
  NAND2_X1 U11528 ( .A1(n11478), .A2(n11480), .ZN(n11698) );
  NAND2_X1 U11529 ( .A1(n11701), .A2(n11702), .ZN(n11480) );
  NAND3_X1 U11530 ( .A1(a_8_), .A2(n11703), .A3(b_19_), .ZN(n11702) );
  OR2_X1 U11531 ( .A1(n11488), .A2(n11487), .ZN(n11703) );
  NAND2_X1 U11532 ( .A1(n11487), .A2(n11488), .ZN(n11701) );
  NAND2_X1 U11533 ( .A1(n11704), .A2(n11705), .ZN(n11488) );
  NAND3_X1 U11534 ( .A1(a_9_), .A2(n11706), .A3(b_19_), .ZN(n11705) );
  OR2_X1 U11535 ( .A1(n11646), .A2(n11644), .ZN(n11706) );
  NAND2_X1 U11536 ( .A1(n11644), .A2(n11646), .ZN(n11704) );
  NAND2_X1 U11537 ( .A1(n11642), .A2(n11707), .ZN(n11646) );
  NAND2_X1 U11538 ( .A1(n11641), .A2(n11643), .ZN(n11707) );
  NAND2_X1 U11539 ( .A1(n11708), .A2(n11709), .ZN(n11643) );
  NAND2_X1 U11540 ( .A1(b_19_), .A2(a_10_), .ZN(n11709) );
  INV_X1 U11541 ( .A(n11710), .ZN(n11708) );
  XNOR2_X1 U11542 ( .A(n11711), .B(n11712), .ZN(n11641) );
  XNOR2_X1 U11543 ( .A(n11713), .B(n11714), .ZN(n11711) );
  NAND2_X1 U11544 ( .A1(a_10_), .A2(n11710), .ZN(n11642) );
  NAND2_X1 U11545 ( .A1(n11715), .A2(n11716), .ZN(n11710) );
  NAND3_X1 U11546 ( .A1(a_11_), .A2(n11717), .A3(b_19_), .ZN(n11716) );
  OR2_X1 U11547 ( .A1(n11638), .A2(n11636), .ZN(n11717) );
  NAND2_X1 U11548 ( .A1(n11636), .A2(n11638), .ZN(n11715) );
  NAND2_X1 U11549 ( .A1(n11718), .A2(n11719), .ZN(n11638) );
  NAND2_X1 U11550 ( .A1(n11635), .A2(n11720), .ZN(n11719) );
  OR2_X1 U11551 ( .A1(n11634), .A2(n11632), .ZN(n11720) );
  NOR2_X1 U11552 ( .A1(n8752), .A2(n8759), .ZN(n11635) );
  NAND2_X1 U11553 ( .A1(n11632), .A2(n11634), .ZN(n11718) );
  NAND2_X1 U11554 ( .A1(n11721), .A2(n11722), .ZN(n11634) );
  NAND2_X1 U11555 ( .A1(n11631), .A2(n11723), .ZN(n11722) );
  OR2_X1 U11556 ( .A1(n11630), .A2(n11629), .ZN(n11723) );
  NOR2_X1 U11557 ( .A1(n8752), .A2(n8310), .ZN(n11631) );
  NAND2_X1 U11558 ( .A1(n11629), .A2(n11630), .ZN(n11721) );
  NAND2_X1 U11559 ( .A1(n11724), .A2(n11725), .ZN(n11630) );
  NAND3_X1 U11560 ( .A1(a_14_), .A2(n11726), .A3(b_19_), .ZN(n11725) );
  NAND2_X1 U11561 ( .A1(n11626), .A2(n11625), .ZN(n11726) );
  OR2_X1 U11562 ( .A1(n11625), .A2(n11626), .ZN(n11724) );
  AND2_X1 U11563 ( .A1(n11727), .A2(n11728), .ZN(n11626) );
  NAND2_X1 U11564 ( .A1(n11623), .A2(n11729), .ZN(n11728) );
  OR2_X1 U11565 ( .A1(n11622), .A2(n11620), .ZN(n11729) );
  NOR2_X1 U11566 ( .A1(n8752), .A2(n8276), .ZN(n11623) );
  NAND2_X1 U11567 ( .A1(n11620), .A2(n11622), .ZN(n11727) );
  NAND2_X1 U11568 ( .A1(n11730), .A2(n11731), .ZN(n11622) );
  NAND3_X1 U11569 ( .A1(a_16_), .A2(n11732), .A3(b_19_), .ZN(n11731) );
  OR2_X1 U11570 ( .A1(n11618), .A2(n11616), .ZN(n11732) );
  NAND2_X1 U11571 ( .A1(n11616), .A2(n11618), .ZN(n11730) );
  NAND2_X1 U11572 ( .A1(n11733), .A2(n11734), .ZN(n11618) );
  NAND2_X1 U11573 ( .A1(n11615), .A2(n11735), .ZN(n11734) );
  OR2_X1 U11574 ( .A1(n11614), .A2(n11613), .ZN(n11735) );
  NOR2_X1 U11575 ( .A1(n8752), .A2(n8210), .ZN(n11615) );
  NAND2_X1 U11576 ( .A1(n11613), .A2(n11614), .ZN(n11733) );
  NAND2_X1 U11577 ( .A1(n11736), .A2(n11737), .ZN(n11614) );
  NAND3_X1 U11578 ( .A1(a_18_), .A2(n11738), .A3(b_19_), .ZN(n11737) );
  NAND2_X1 U11579 ( .A1(n11610), .A2(n11609), .ZN(n11738) );
  OR2_X1 U11580 ( .A1(n11609), .A2(n11610), .ZN(n11736) );
  AND2_X1 U11581 ( .A1(n11739), .A2(n11740), .ZN(n11610) );
  NAND2_X1 U11582 ( .A1(n11607), .A2(n11741), .ZN(n11740) );
  OR2_X1 U11583 ( .A1(n11606), .A2(n11605), .ZN(n11741) );
  INV_X1 U11584 ( .A(n8712), .ZN(n11607) );
  NAND2_X1 U11585 ( .A1(b_19_), .A2(a_19_), .ZN(n8712) );
  NAND2_X1 U11586 ( .A1(n11605), .A2(n11606), .ZN(n11739) );
  NAND2_X1 U11587 ( .A1(n11742), .A2(n11743), .ZN(n11606) );
  NAND3_X1 U11588 ( .A1(a_20_), .A2(n11744), .A3(b_19_), .ZN(n11743) );
  NAND2_X1 U11589 ( .A1(n11603), .A2(n11601), .ZN(n11744) );
  OR2_X1 U11590 ( .A1(n11601), .A2(n11603), .ZN(n11742) );
  AND2_X1 U11591 ( .A1(n11745), .A2(n11746), .ZN(n11603) );
  NAND2_X1 U11592 ( .A1(n11532), .A2(n11747), .ZN(n11746) );
  NAND2_X1 U11593 ( .A1(n11531), .A2(n11530), .ZN(n11747) );
  NOR2_X1 U11594 ( .A1(n8752), .A2(n8750), .ZN(n11532) );
  OR2_X1 U11595 ( .A1(n11530), .A2(n11531), .ZN(n11745) );
  AND2_X1 U11596 ( .A1(n11748), .A2(n11749), .ZN(n11531) );
  NAND3_X1 U11597 ( .A1(a_22_), .A2(n11750), .A3(b_19_), .ZN(n11749) );
  OR2_X1 U11598 ( .A1(n11598), .A2(n11596), .ZN(n11750) );
  NAND2_X1 U11599 ( .A1(n11596), .A2(n11598), .ZN(n11748) );
  NAND2_X1 U11600 ( .A1(n11751), .A2(n11752), .ZN(n11598) );
  NAND2_X1 U11601 ( .A1(n11595), .A2(n11753), .ZN(n11752) );
  OR2_X1 U11602 ( .A1(n11594), .A2(n11592), .ZN(n11753) );
  NOR2_X1 U11603 ( .A1(n8752), .A2(n8747), .ZN(n11595) );
  NAND2_X1 U11604 ( .A1(n11592), .A2(n11594), .ZN(n11751) );
  NAND2_X1 U11605 ( .A1(n11754), .A2(n11755), .ZN(n11594) );
  NAND3_X1 U11606 ( .A1(a_24_), .A2(n11756), .A3(b_19_), .ZN(n11755) );
  NAND2_X1 U11607 ( .A1(n11590), .A2(n11589), .ZN(n11756) );
  OR2_X1 U11608 ( .A1(n11589), .A2(n11590), .ZN(n11754) );
  AND2_X1 U11609 ( .A1(n11757), .A2(n11758), .ZN(n11590) );
  NAND2_X1 U11610 ( .A1(n11587), .A2(n11759), .ZN(n11758) );
  OR2_X1 U11611 ( .A1(n11586), .A2(n11585), .ZN(n11759) );
  NOR2_X1 U11612 ( .A1(n8752), .A2(n8744), .ZN(n11587) );
  NAND2_X1 U11613 ( .A1(n11585), .A2(n11586), .ZN(n11757) );
  NAND2_X1 U11614 ( .A1(n11582), .A2(n11760), .ZN(n11586) );
  NAND2_X1 U11615 ( .A1(n11581), .A2(n11583), .ZN(n11760) );
  NAND2_X1 U11616 ( .A1(n11761), .A2(n11762), .ZN(n11583) );
  NAND2_X1 U11617 ( .A1(b_19_), .A2(a_26_), .ZN(n11762) );
  INV_X1 U11618 ( .A(n11763), .ZN(n11761) );
  XNOR2_X1 U11619 ( .A(n11764), .B(n11765), .ZN(n11581) );
  NAND2_X1 U11620 ( .A1(n11766), .A2(n11767), .ZN(n11764) );
  NAND2_X1 U11621 ( .A1(a_26_), .A2(n11763), .ZN(n11582) );
  NAND2_X1 U11622 ( .A1(n11554), .A2(n11768), .ZN(n11763) );
  NAND2_X1 U11623 ( .A1(n11553), .A2(n11555), .ZN(n11768) );
  NAND2_X1 U11624 ( .A1(n11769), .A2(n11770), .ZN(n11555) );
  NAND2_X1 U11625 ( .A1(b_19_), .A2(a_27_), .ZN(n11770) );
  INV_X1 U11626 ( .A(n11771), .ZN(n11769) );
  XNOR2_X1 U11627 ( .A(n11772), .B(n11773), .ZN(n11553) );
  XOR2_X1 U11628 ( .A(n11774), .B(n11775), .Z(n11772) );
  NAND2_X1 U11629 ( .A1(b_18_), .A2(a_28_), .ZN(n11774) );
  NAND2_X1 U11630 ( .A1(a_27_), .A2(n11771), .ZN(n11554) );
  NAND2_X1 U11631 ( .A1(n11776), .A2(n11777), .ZN(n11771) );
  NAND3_X1 U11632 ( .A1(a_28_), .A2(n11778), .A3(b_19_), .ZN(n11777) );
  NAND2_X1 U11633 ( .A1(n11563), .A2(n11561), .ZN(n11778) );
  OR2_X1 U11634 ( .A1(n11561), .A2(n11563), .ZN(n11776) );
  AND2_X1 U11635 ( .A1(n11779), .A2(n11780), .ZN(n11563) );
  NAND2_X1 U11636 ( .A1(n11577), .A2(n11781), .ZN(n11780) );
  OR2_X1 U11637 ( .A1(n11578), .A2(n11579), .ZN(n11781) );
  NOR2_X1 U11638 ( .A1(n8752), .A2(n7890), .ZN(n11577) );
  NAND2_X1 U11639 ( .A1(n11579), .A2(n11578), .ZN(n11779) );
  NAND2_X1 U11640 ( .A1(n11782), .A2(n11783), .ZN(n11578) );
  NAND2_X1 U11641 ( .A1(b_17_), .A2(n11784), .ZN(n11783) );
  NAND2_X1 U11642 ( .A1(n7864), .A2(n11785), .ZN(n11784) );
  NAND2_X1 U11643 ( .A1(a_31_), .A2(n8195), .ZN(n11785) );
  NAND2_X1 U11644 ( .A1(b_18_), .A2(n11786), .ZN(n11782) );
  NAND2_X1 U11645 ( .A1(n9137), .A2(n11787), .ZN(n11786) );
  NAND2_X1 U11646 ( .A1(a_30_), .A2(n8754), .ZN(n11787) );
  AND3_X1 U11647 ( .A1(b_18_), .A2(b_19_), .A3(n7818), .ZN(n11579) );
  XNOR2_X1 U11648 ( .A(n11788), .B(n11789), .ZN(n11561) );
  XOR2_X1 U11649 ( .A(n11790), .B(n11791), .Z(n11788) );
  XNOR2_X1 U11650 ( .A(n11792), .B(n11793), .ZN(n11585) );
  NAND2_X1 U11651 ( .A1(n11794), .A2(n11795), .ZN(n11792) );
  XNOR2_X1 U11652 ( .A(n11796), .B(n11797), .ZN(n11589) );
  XOR2_X1 U11653 ( .A(n11798), .B(n11799), .Z(n11796) );
  XNOR2_X1 U11654 ( .A(n11800), .B(n11801), .ZN(n11592) );
  XNOR2_X1 U11655 ( .A(n11802), .B(n11803), .ZN(n11800) );
  NOR2_X1 U11656 ( .A1(n8745), .A2(n8195), .ZN(n11803) );
  XNOR2_X1 U11657 ( .A(n11804), .B(n11805), .ZN(n11596) );
  XOR2_X1 U11658 ( .A(n11806), .B(n11807), .Z(n11805) );
  NAND2_X1 U11659 ( .A1(b_18_), .A2(a_23_), .ZN(n11807) );
  XOR2_X1 U11660 ( .A(n11808), .B(n11809), .Z(n11530) );
  NAND2_X1 U11661 ( .A1(n11810), .A2(n11811), .ZN(n11808) );
  XNOR2_X1 U11662 ( .A(n11812), .B(n11813), .ZN(n11601) );
  XOR2_X1 U11663 ( .A(n11814), .B(n11815), .Z(n11812) );
  XNOR2_X1 U11664 ( .A(n11816), .B(n11817), .ZN(n11605) );
  XNOR2_X1 U11665 ( .A(n11818), .B(n11819), .ZN(n11816) );
  NOR2_X1 U11666 ( .A1(n8751), .A2(n8195), .ZN(n11819) );
  XOR2_X1 U11667 ( .A(n11820), .B(n11821), .Z(n11609) );
  XNOR2_X1 U11668 ( .A(n11822), .B(n11823), .ZN(n11821) );
  XOR2_X1 U11669 ( .A(n11824), .B(n11825), .Z(n11613) );
  XOR2_X1 U11670 ( .A(n11826), .B(n11827), .Z(n11824) );
  XNOR2_X1 U11671 ( .A(n11828), .B(n11829), .ZN(n11616) );
  XNOR2_X1 U11672 ( .A(n11830), .B(n11831), .ZN(n11829) );
  XNOR2_X1 U11673 ( .A(n11832), .B(n11833), .ZN(n11620) );
  XOR2_X1 U11674 ( .A(n11834), .B(n11835), .Z(n11833) );
  NAND2_X1 U11675 ( .A1(b_18_), .A2(a_16_), .ZN(n11835) );
  XOR2_X1 U11676 ( .A(n11836), .B(n11837), .Z(n11625) );
  XNOR2_X1 U11677 ( .A(n11838), .B(n11839), .ZN(n11837) );
  XNOR2_X1 U11678 ( .A(n11840), .B(n11841), .ZN(n11629) );
  XNOR2_X1 U11679 ( .A(n11842), .B(n11843), .ZN(n11840) );
  NOR2_X1 U11680 ( .A1(n8757), .A2(n8195), .ZN(n11843) );
  XNOR2_X1 U11681 ( .A(n11844), .B(n11845), .ZN(n11632) );
  XNOR2_X1 U11682 ( .A(n11846), .B(n11847), .ZN(n11844) );
  NOR2_X1 U11683 ( .A1(n8310), .A2(n8195), .ZN(n11847) );
  XNOR2_X1 U11684 ( .A(n11848), .B(n11849), .ZN(n11636) );
  XNOR2_X1 U11685 ( .A(n11850), .B(n11851), .ZN(n11849) );
  XNOR2_X1 U11686 ( .A(n11852), .B(n11853), .ZN(n11644) );
  XNOR2_X1 U11687 ( .A(n11854), .B(n11855), .ZN(n11852) );
  NOR2_X1 U11688 ( .A1(n8761), .A2(n8195), .ZN(n11855) );
  XNOR2_X1 U11689 ( .A(n11856), .B(n11857), .ZN(n11487) );
  NAND2_X1 U11690 ( .A1(n11858), .A2(n11859), .ZN(n11856) );
  XNOR2_X1 U11691 ( .A(n11860), .B(n11861), .ZN(n11478) );
  NAND2_X1 U11692 ( .A1(n11862), .A2(n11863), .ZN(n11860) );
  XOR2_X1 U11693 ( .A(n11864), .B(n11865), .Z(n11649) );
  NAND2_X1 U11694 ( .A1(n11866), .A2(n11867), .ZN(n11864) );
  XNOR2_X1 U11695 ( .A(n11868), .B(n11869), .ZN(n11652) );
  NAND2_X1 U11696 ( .A1(n11870), .A2(n11871), .ZN(n11868) );
  XNOR2_X1 U11697 ( .A(n11872), .B(n11873), .ZN(n11465) );
  NAND2_X1 U11698 ( .A1(n11874), .A2(n11875), .ZN(n11872) );
  XNOR2_X1 U11699 ( .A(n11876), .B(n11877), .ZN(n11656) );
  NAND2_X1 U11700 ( .A1(n11878), .A2(n11879), .ZN(n11876) );
  XNOR2_X1 U11701 ( .A(n11880), .B(n11881), .ZN(n11660) );
  NAND2_X1 U11702 ( .A1(n11882), .A2(n11883), .ZN(n11880) );
  XNOR2_X1 U11703 ( .A(n11884), .B(n11885), .ZN(n11664) );
  NAND2_X1 U11704 ( .A1(n11886), .A2(n11887), .ZN(n11884) );
  XOR2_X1 U11705 ( .A(n11888), .B(n11889), .Z(n11668) );
  XOR2_X1 U11706 ( .A(n11890), .B(n11891), .Z(n11888) );
  XOR2_X1 U11707 ( .A(n8964), .B(n8963), .Z(n11672) );
  NAND2_X1 U11708 ( .A1(n11892), .A2(n11893), .ZN(n8869) );
  NAND2_X1 U11709 ( .A1(n8963), .A2(n8964), .ZN(n11893) );
  XOR2_X1 U11710 ( .A(n8954), .B(n11894), .Z(n11892) );
  NAND3_X1 U11711 ( .A1(n8963), .A2(n8964), .A3(n11895), .ZN(n8870) );
  XOR2_X1 U11712 ( .A(n8954), .B(n8953), .Z(n11895) );
  NAND2_X1 U11713 ( .A1(n11896), .A2(n11897), .ZN(n8964) );
  NAND3_X1 U11714 ( .A1(a_0_), .A2(n11898), .A3(b_18_), .ZN(n11897) );
  OR2_X1 U11715 ( .A1(n11673), .A2(n11675), .ZN(n11898) );
  NAND2_X1 U11716 ( .A1(n11673), .A2(n11675), .ZN(n11896) );
  NAND2_X1 U11717 ( .A1(n11899), .A2(n11900), .ZN(n11675) );
  NAND2_X1 U11718 ( .A1(n11891), .A2(n11901), .ZN(n11900) );
  OR2_X1 U11719 ( .A1(n11889), .A2(n11890), .ZN(n11901) );
  NOR2_X1 U11720 ( .A1(n8195), .A2(n8617), .ZN(n11891) );
  NAND2_X1 U11721 ( .A1(n11889), .A2(n11890), .ZN(n11899) );
  NAND2_X1 U11722 ( .A1(n11886), .A2(n11902), .ZN(n11890) );
  NAND2_X1 U11723 ( .A1(n11885), .A2(n11887), .ZN(n11902) );
  NAND2_X1 U11724 ( .A1(n11903), .A2(n11904), .ZN(n11887) );
  NAND2_X1 U11725 ( .A1(b_18_), .A2(a_2_), .ZN(n11904) );
  INV_X1 U11726 ( .A(n11905), .ZN(n11903) );
  XNOR2_X1 U11727 ( .A(n11906), .B(n11907), .ZN(n11885) );
  XNOR2_X1 U11728 ( .A(n11908), .B(n11909), .ZN(n11906) );
  NOR2_X1 U11729 ( .A1(n8567), .A2(n8754), .ZN(n11909) );
  NAND2_X1 U11730 ( .A1(a_2_), .A2(n11905), .ZN(n11886) );
  NAND2_X1 U11731 ( .A1(n11882), .A2(n11910), .ZN(n11905) );
  NAND2_X1 U11732 ( .A1(n11881), .A2(n11883), .ZN(n11910) );
  NAND2_X1 U11733 ( .A1(n11911), .A2(n11912), .ZN(n11883) );
  NAND2_X1 U11734 ( .A1(b_18_), .A2(a_3_), .ZN(n11912) );
  INV_X1 U11735 ( .A(n11913), .ZN(n11911) );
  XNOR2_X1 U11736 ( .A(n11914), .B(n11915), .ZN(n11881) );
  XOR2_X1 U11737 ( .A(n11916), .B(n11917), .Z(n11915) );
  NAND2_X1 U11738 ( .A1(b_17_), .A2(a_4_), .ZN(n11917) );
  NAND2_X1 U11739 ( .A1(a_3_), .A2(n11913), .ZN(n11882) );
  NAND2_X1 U11740 ( .A1(n11878), .A2(n11918), .ZN(n11913) );
  NAND2_X1 U11741 ( .A1(n11877), .A2(n11879), .ZN(n11918) );
  NAND2_X1 U11742 ( .A1(n11919), .A2(n11920), .ZN(n11879) );
  NAND2_X1 U11743 ( .A1(b_18_), .A2(a_4_), .ZN(n11920) );
  INV_X1 U11744 ( .A(n11921), .ZN(n11919) );
  XNOR2_X1 U11745 ( .A(n11922), .B(n11923), .ZN(n11877) );
  XOR2_X1 U11746 ( .A(n11924), .B(n11925), .Z(n11923) );
  NAND2_X1 U11747 ( .A1(b_17_), .A2(a_5_), .ZN(n11925) );
  NAND2_X1 U11748 ( .A1(a_4_), .A2(n11921), .ZN(n11878) );
  NAND2_X1 U11749 ( .A1(n11874), .A2(n11926), .ZN(n11921) );
  NAND2_X1 U11750 ( .A1(n11873), .A2(n11875), .ZN(n11926) );
  NAND2_X1 U11751 ( .A1(n11927), .A2(n11928), .ZN(n11875) );
  NAND2_X1 U11752 ( .A1(b_18_), .A2(a_5_), .ZN(n11928) );
  INV_X1 U11753 ( .A(n11929), .ZN(n11927) );
  XNOR2_X1 U11754 ( .A(n11930), .B(n11931), .ZN(n11873) );
  XOR2_X1 U11755 ( .A(n11932), .B(n11933), .Z(n11931) );
  NAND2_X1 U11756 ( .A1(b_17_), .A2(a_6_), .ZN(n11933) );
  NAND2_X1 U11757 ( .A1(a_5_), .A2(n11929), .ZN(n11874) );
  NAND2_X1 U11758 ( .A1(n11870), .A2(n11934), .ZN(n11929) );
  NAND2_X1 U11759 ( .A1(n11869), .A2(n11871), .ZN(n11934) );
  NAND2_X1 U11760 ( .A1(n11935), .A2(n11936), .ZN(n11871) );
  NAND2_X1 U11761 ( .A1(b_18_), .A2(a_6_), .ZN(n11936) );
  INV_X1 U11762 ( .A(n11937), .ZN(n11935) );
  XNOR2_X1 U11763 ( .A(n11938), .B(n11939), .ZN(n11869) );
  XOR2_X1 U11764 ( .A(n11940), .B(n11941), .Z(n11939) );
  NAND2_X1 U11765 ( .A1(b_17_), .A2(a_7_), .ZN(n11941) );
  NAND2_X1 U11766 ( .A1(a_6_), .A2(n11937), .ZN(n11870) );
  NAND2_X1 U11767 ( .A1(n11866), .A2(n11942), .ZN(n11937) );
  NAND2_X1 U11768 ( .A1(n11865), .A2(n11867), .ZN(n11942) );
  NAND2_X1 U11769 ( .A1(n11943), .A2(n11944), .ZN(n11867) );
  NAND2_X1 U11770 ( .A1(b_18_), .A2(a_7_), .ZN(n11944) );
  INV_X1 U11771 ( .A(n11945), .ZN(n11943) );
  XNOR2_X1 U11772 ( .A(n11946), .B(n11947), .ZN(n11865) );
  XOR2_X1 U11773 ( .A(n11948), .B(n11949), .Z(n11947) );
  NAND2_X1 U11774 ( .A1(b_17_), .A2(a_8_), .ZN(n11949) );
  NAND2_X1 U11775 ( .A1(a_7_), .A2(n11945), .ZN(n11866) );
  NAND2_X1 U11776 ( .A1(n11862), .A2(n11950), .ZN(n11945) );
  NAND2_X1 U11777 ( .A1(n11861), .A2(n11863), .ZN(n11950) );
  NAND2_X1 U11778 ( .A1(n11951), .A2(n11952), .ZN(n11863) );
  NAND2_X1 U11779 ( .A1(b_18_), .A2(a_8_), .ZN(n11952) );
  INV_X1 U11780 ( .A(n11953), .ZN(n11951) );
  XNOR2_X1 U11781 ( .A(n11954), .B(n11955), .ZN(n11861) );
  XNOR2_X1 U11782 ( .A(n11956), .B(n11957), .ZN(n11954) );
  NOR2_X1 U11783 ( .A1(n8426), .A2(n8754), .ZN(n11957) );
  NAND2_X1 U11784 ( .A1(a_8_), .A2(n11953), .ZN(n11862) );
  NAND2_X1 U11785 ( .A1(n11858), .A2(n11958), .ZN(n11953) );
  NAND2_X1 U11786 ( .A1(n11857), .A2(n11859), .ZN(n11958) );
  NAND2_X1 U11787 ( .A1(n11959), .A2(n11960), .ZN(n11859) );
  NAND2_X1 U11788 ( .A1(b_18_), .A2(a_9_), .ZN(n11960) );
  INV_X1 U11789 ( .A(n11961), .ZN(n11959) );
  XNOR2_X1 U11790 ( .A(n11962), .B(n11963), .ZN(n11857) );
  XNOR2_X1 U11791 ( .A(n11964), .B(n11965), .ZN(n11962) );
  NOR2_X1 U11792 ( .A1(n8761), .A2(n8754), .ZN(n11965) );
  NAND2_X1 U11793 ( .A1(a_9_), .A2(n11961), .ZN(n11858) );
  NAND2_X1 U11794 ( .A1(n11966), .A2(n11967), .ZN(n11961) );
  NAND3_X1 U11795 ( .A1(a_10_), .A2(n11968), .A3(b_18_), .ZN(n11967) );
  NAND2_X1 U11796 ( .A1(n11854), .A2(n11853), .ZN(n11968) );
  OR2_X1 U11797 ( .A1(n11853), .A2(n11854), .ZN(n11966) );
  AND2_X1 U11798 ( .A1(n11969), .A2(n11970), .ZN(n11854) );
  NAND2_X1 U11799 ( .A1(n11713), .A2(n11971), .ZN(n11970) );
  NAND2_X1 U11800 ( .A1(n11714), .A2(n11712), .ZN(n11971) );
  NOR2_X1 U11801 ( .A1(n8195), .A2(n8376), .ZN(n11713) );
  OR2_X1 U11802 ( .A1(n11712), .A2(n11714), .ZN(n11969) );
  AND2_X1 U11803 ( .A1(n11972), .A2(n11973), .ZN(n11714) );
  NAND2_X1 U11804 ( .A1(n11851), .A2(n11974), .ZN(n11973) );
  OR2_X1 U11805 ( .A1(n11848), .A2(n11850), .ZN(n11974) );
  NOR2_X1 U11806 ( .A1(n8195), .A2(n8759), .ZN(n11851) );
  NAND2_X1 U11807 ( .A1(n11848), .A2(n11850), .ZN(n11972) );
  NAND2_X1 U11808 ( .A1(n11975), .A2(n11976), .ZN(n11850) );
  NAND3_X1 U11809 ( .A1(a_13_), .A2(n11977), .A3(b_18_), .ZN(n11976) );
  NAND2_X1 U11810 ( .A1(n11846), .A2(n11845), .ZN(n11977) );
  OR2_X1 U11811 ( .A1(n11845), .A2(n11846), .ZN(n11975) );
  AND2_X1 U11812 ( .A1(n11978), .A2(n11979), .ZN(n11846) );
  NAND3_X1 U11813 ( .A1(a_14_), .A2(n11980), .A3(b_18_), .ZN(n11979) );
  NAND2_X1 U11814 ( .A1(n11842), .A2(n11841), .ZN(n11980) );
  OR2_X1 U11815 ( .A1(n11841), .A2(n11842), .ZN(n11978) );
  AND2_X1 U11816 ( .A1(n11981), .A2(n11982), .ZN(n11842) );
  NAND2_X1 U11817 ( .A1(n11839), .A2(n11983), .ZN(n11982) );
  OR2_X1 U11818 ( .A1(n11836), .A2(n11838), .ZN(n11983) );
  NOR2_X1 U11819 ( .A1(n8195), .A2(n8276), .ZN(n11839) );
  NAND2_X1 U11820 ( .A1(n11836), .A2(n11838), .ZN(n11981) );
  NAND2_X1 U11821 ( .A1(n11984), .A2(n11985), .ZN(n11838) );
  NAND3_X1 U11822 ( .A1(a_16_), .A2(n11986), .A3(b_18_), .ZN(n11985) );
  OR2_X1 U11823 ( .A1(n11834), .A2(n11832), .ZN(n11986) );
  NAND2_X1 U11824 ( .A1(n11832), .A2(n11834), .ZN(n11984) );
  NAND2_X1 U11825 ( .A1(n11987), .A2(n11988), .ZN(n11834) );
  NAND2_X1 U11826 ( .A1(n11831), .A2(n11989), .ZN(n11988) );
  OR2_X1 U11827 ( .A1(n11828), .A2(n11830), .ZN(n11989) );
  NOR2_X1 U11828 ( .A1(n8195), .A2(n8210), .ZN(n11831) );
  NAND2_X1 U11829 ( .A1(n11828), .A2(n11830), .ZN(n11987) );
  NAND2_X1 U11830 ( .A1(n11990), .A2(n11991), .ZN(n11830) );
  NAND2_X1 U11831 ( .A1(n11825), .A2(n11992), .ZN(n11991) );
  OR2_X1 U11832 ( .A1(n11826), .A2(n11827), .ZN(n11992) );
  XNOR2_X1 U11833 ( .A(n11993), .B(n11994), .ZN(n11825) );
  XNOR2_X1 U11834 ( .A(n11995), .B(n11996), .ZN(n11994) );
  NAND2_X1 U11835 ( .A1(n11827), .A2(n11826), .ZN(n11990) );
  NAND2_X1 U11836 ( .A1(n11997), .A2(n11998), .ZN(n11826) );
  NAND2_X1 U11837 ( .A1(n11823), .A2(n11999), .ZN(n11998) );
  OR2_X1 U11838 ( .A1(n11820), .A2(n11822), .ZN(n11999) );
  NOR2_X1 U11839 ( .A1(n8195), .A2(n8170), .ZN(n11823) );
  NAND2_X1 U11840 ( .A1(n11820), .A2(n11822), .ZN(n11997) );
  NAND2_X1 U11841 ( .A1(n12000), .A2(n12001), .ZN(n11822) );
  NAND3_X1 U11842 ( .A1(a_20_), .A2(n12002), .A3(b_18_), .ZN(n12001) );
  NAND2_X1 U11843 ( .A1(n11818), .A2(n11817), .ZN(n12002) );
  OR2_X1 U11844 ( .A1(n11817), .A2(n11818), .ZN(n12000) );
  AND2_X1 U11845 ( .A1(n12003), .A2(n12004), .ZN(n11818) );
  NAND2_X1 U11846 ( .A1(n11814), .A2(n12005), .ZN(n12004) );
  OR2_X1 U11847 ( .A1(n11813), .A2(n11815), .ZN(n12005) );
  NOR2_X1 U11848 ( .A1(n8195), .A2(n8750), .ZN(n11814) );
  NAND2_X1 U11849 ( .A1(n11813), .A2(n11815), .ZN(n12003) );
  NAND2_X1 U11850 ( .A1(n11810), .A2(n12006), .ZN(n11815) );
  NAND2_X1 U11851 ( .A1(n11809), .A2(n11811), .ZN(n12006) );
  NAND2_X1 U11852 ( .A1(n12007), .A2(n12008), .ZN(n11811) );
  NAND2_X1 U11853 ( .A1(b_18_), .A2(a_22_), .ZN(n12008) );
  INV_X1 U11854 ( .A(n12009), .ZN(n12007) );
  XNOR2_X1 U11855 ( .A(n12010), .B(n12011), .ZN(n11809) );
  XNOR2_X1 U11856 ( .A(n12012), .B(n12013), .ZN(n12011) );
  NAND2_X1 U11857 ( .A1(a_22_), .A2(n12009), .ZN(n11810) );
  NAND2_X1 U11858 ( .A1(n12014), .A2(n12015), .ZN(n12009) );
  NAND3_X1 U11859 ( .A1(a_23_), .A2(n12016), .A3(b_18_), .ZN(n12015) );
  OR2_X1 U11860 ( .A1(n11804), .A2(n11806), .ZN(n12016) );
  NAND2_X1 U11861 ( .A1(n11804), .A2(n11806), .ZN(n12014) );
  NAND2_X1 U11862 ( .A1(n12017), .A2(n12018), .ZN(n11806) );
  NAND3_X1 U11863 ( .A1(a_24_), .A2(n12019), .A3(b_18_), .ZN(n12018) );
  NAND2_X1 U11864 ( .A1(n11802), .A2(n11801), .ZN(n12019) );
  OR2_X1 U11865 ( .A1(n11801), .A2(n11802), .ZN(n12017) );
  AND2_X1 U11866 ( .A1(n12020), .A2(n12021), .ZN(n11802) );
  NAND2_X1 U11867 ( .A1(n11799), .A2(n12022), .ZN(n12021) );
  OR2_X1 U11868 ( .A1(n11797), .A2(n11798), .ZN(n12022) );
  NOR2_X1 U11869 ( .A1(n8195), .A2(n8744), .ZN(n11799) );
  NAND2_X1 U11870 ( .A1(n11797), .A2(n11798), .ZN(n12020) );
  NAND2_X1 U11871 ( .A1(n11794), .A2(n12023), .ZN(n11798) );
  NAND2_X1 U11872 ( .A1(n11793), .A2(n11795), .ZN(n12023) );
  NAND2_X1 U11873 ( .A1(n12024), .A2(n12025), .ZN(n11795) );
  NAND2_X1 U11874 ( .A1(b_18_), .A2(a_26_), .ZN(n12025) );
  INV_X1 U11875 ( .A(n12026), .ZN(n12024) );
  XNOR2_X1 U11876 ( .A(n12027), .B(n12028), .ZN(n11793) );
  NAND2_X1 U11877 ( .A1(n12029), .A2(n12030), .ZN(n12027) );
  NAND2_X1 U11878 ( .A1(a_26_), .A2(n12026), .ZN(n11794) );
  NAND2_X1 U11879 ( .A1(n11766), .A2(n12031), .ZN(n12026) );
  NAND2_X1 U11880 ( .A1(n11765), .A2(n11767), .ZN(n12031) );
  NAND2_X1 U11881 ( .A1(n12032), .A2(n12033), .ZN(n11767) );
  NAND2_X1 U11882 ( .A1(b_18_), .A2(a_27_), .ZN(n12033) );
  INV_X1 U11883 ( .A(n12034), .ZN(n12032) );
  XNOR2_X1 U11884 ( .A(n12035), .B(n12036), .ZN(n11765) );
  XOR2_X1 U11885 ( .A(n12037), .B(n12038), .Z(n12035) );
  NAND2_X1 U11886 ( .A1(b_17_), .A2(a_28_), .ZN(n12037) );
  NAND2_X1 U11887 ( .A1(a_27_), .A2(n12034), .ZN(n11766) );
  NAND2_X1 U11888 ( .A1(n12039), .A2(n12040), .ZN(n12034) );
  NAND3_X1 U11889 ( .A1(a_28_), .A2(n12041), .A3(b_18_), .ZN(n12040) );
  NAND2_X1 U11890 ( .A1(n11775), .A2(n11773), .ZN(n12041) );
  OR2_X1 U11891 ( .A1(n11773), .A2(n11775), .ZN(n12039) );
  AND2_X1 U11892 ( .A1(n12042), .A2(n12043), .ZN(n11775) );
  NAND2_X1 U11893 ( .A1(n11789), .A2(n12044), .ZN(n12043) );
  OR2_X1 U11894 ( .A1(n11790), .A2(n11791), .ZN(n12044) );
  NOR2_X1 U11895 ( .A1(n8195), .A2(n7890), .ZN(n11789) );
  NAND2_X1 U11896 ( .A1(n11791), .A2(n11790), .ZN(n12042) );
  NAND2_X1 U11897 ( .A1(n12045), .A2(n12046), .ZN(n11790) );
  NAND2_X1 U11898 ( .A1(b_16_), .A2(n12047), .ZN(n12046) );
  NAND2_X1 U11899 ( .A1(n7864), .A2(n12048), .ZN(n12047) );
  NAND2_X1 U11900 ( .A1(a_31_), .A2(n8754), .ZN(n12048) );
  NAND2_X1 U11901 ( .A1(b_17_), .A2(n12049), .ZN(n12045) );
  NAND2_X1 U11902 ( .A1(n9137), .A2(n12050), .ZN(n12049) );
  NAND2_X1 U11903 ( .A1(a_30_), .A2(n8251), .ZN(n12050) );
  AND3_X1 U11904 ( .A1(b_17_), .A2(b_18_), .A3(n7818), .ZN(n11791) );
  XNOR2_X1 U11905 ( .A(n12051), .B(n12052), .ZN(n11773) );
  XOR2_X1 U11906 ( .A(n12053), .B(n12054), .Z(n12051) );
  XNOR2_X1 U11907 ( .A(n12055), .B(n12056), .ZN(n11797) );
  NAND2_X1 U11908 ( .A1(n12057), .A2(n12058), .ZN(n12055) );
  XNOR2_X1 U11909 ( .A(n12059), .B(n12060), .ZN(n11801) );
  XOR2_X1 U11910 ( .A(n12061), .B(n12062), .Z(n12059) );
  XNOR2_X1 U11911 ( .A(n12063), .B(n12064), .ZN(n11804) );
  XNOR2_X1 U11912 ( .A(n12065), .B(n12066), .ZN(n12063) );
  NOR2_X1 U11913 ( .A1(n8745), .A2(n8754), .ZN(n12066) );
  XNOR2_X1 U11914 ( .A(n12067), .B(n12068), .ZN(n11813) );
  XOR2_X1 U11915 ( .A(n12069), .B(n12070), .Z(n12068) );
  NAND2_X1 U11916 ( .A1(b_17_), .A2(a_22_), .ZN(n12070) );
  XNOR2_X1 U11917 ( .A(n12071), .B(n12072), .ZN(n11817) );
  XOR2_X1 U11918 ( .A(n12073), .B(n12074), .Z(n12071) );
  XNOR2_X1 U11919 ( .A(n12075), .B(n12076), .ZN(n11820) );
  XNOR2_X1 U11920 ( .A(n12077), .B(n12078), .ZN(n12075) );
  NOR2_X1 U11921 ( .A1(n8751), .A2(n8754), .ZN(n12078) );
  INV_X1 U11922 ( .A(n8709), .ZN(n11827) );
  NAND2_X1 U11923 ( .A1(b_18_), .A2(a_18_), .ZN(n8709) );
  XNOR2_X1 U11924 ( .A(n12079), .B(n12080), .ZN(n11828) );
  XNOR2_X1 U11925 ( .A(n12081), .B(n12082), .ZN(n12079) );
  NOR2_X1 U11926 ( .A1(n8753), .A2(n8754), .ZN(n12082) );
  XOR2_X1 U11927 ( .A(n12083), .B(n12084), .Z(n11832) );
  XOR2_X1 U11928 ( .A(n12085), .B(n12086), .Z(n12083) );
  XNOR2_X1 U11929 ( .A(n12087), .B(n12088), .ZN(n11836) );
  XOR2_X1 U11930 ( .A(n12089), .B(n12090), .Z(n12088) );
  NAND2_X1 U11931 ( .A1(b_17_), .A2(a_16_), .ZN(n12090) );
  XOR2_X1 U11932 ( .A(n12091), .B(n12092), .Z(n11841) );
  XNOR2_X1 U11933 ( .A(n12093), .B(n12094), .ZN(n12092) );
  XNOR2_X1 U11934 ( .A(n12095), .B(n12096), .ZN(n11845) );
  XOR2_X1 U11935 ( .A(n12097), .B(n12098), .Z(n12095) );
  XNOR2_X1 U11936 ( .A(n12099), .B(n12100), .ZN(n11848) );
  XNOR2_X1 U11937 ( .A(n12101), .B(n12102), .ZN(n12099) );
  NOR2_X1 U11938 ( .A1(n8310), .A2(n8754), .ZN(n12102) );
  XOR2_X1 U11939 ( .A(n12103), .B(n12104), .Z(n11712) );
  XOR2_X1 U11940 ( .A(n12105), .B(n12106), .Z(n12104) );
  NAND2_X1 U11941 ( .A1(b_17_), .A2(a_12_), .ZN(n12106) );
  XOR2_X1 U11942 ( .A(n12107), .B(n12108), .Z(n11853) );
  XOR2_X1 U11943 ( .A(n12109), .B(n12110), .Z(n12108) );
  NAND2_X1 U11944 ( .A1(b_17_), .A2(a_11_), .ZN(n12110) );
  XNOR2_X1 U11945 ( .A(n12111), .B(n12112), .ZN(n11889) );
  XOR2_X1 U11946 ( .A(n12113), .B(n12114), .Z(n12112) );
  NAND2_X1 U11947 ( .A1(b_17_), .A2(a_2_), .ZN(n12114) );
  XNOR2_X1 U11948 ( .A(n12115), .B(n12116), .ZN(n11673) );
  XNOR2_X1 U11949 ( .A(n12117), .B(n12118), .ZN(n12115) );
  NOR2_X1 U11950 ( .A1(n8617), .A2(n8754), .ZN(n12118) );
  XNOR2_X1 U11951 ( .A(n12119), .B(n12120), .ZN(n8963) );
  XOR2_X1 U11952 ( .A(n12121), .B(n12122), .Z(n12120) );
  NAND2_X1 U11953 ( .A1(b_17_), .A2(a_0_), .ZN(n12122) );
  NAND3_X1 U11954 ( .A1(n8953), .A2(n8954), .A3(n12123), .ZN(n8876) );
  XOR2_X1 U11955 ( .A(n8956), .B(n8955), .Z(n12123) );
  NAND2_X1 U11956 ( .A1(n12124), .A2(n12125), .ZN(n8954) );
  NAND3_X1 U11957 ( .A1(a_0_), .A2(n12126), .A3(b_17_), .ZN(n12125) );
  OR2_X1 U11958 ( .A1(n12121), .A2(n12119), .ZN(n12126) );
  NAND2_X1 U11959 ( .A1(n12119), .A2(n12121), .ZN(n12124) );
  NAND2_X1 U11960 ( .A1(n12127), .A2(n12128), .ZN(n12121) );
  NAND3_X1 U11961 ( .A1(a_1_), .A2(n12129), .A3(b_17_), .ZN(n12128) );
  NAND2_X1 U11962 ( .A1(n12117), .A2(n12116), .ZN(n12129) );
  OR2_X1 U11963 ( .A1(n12116), .A2(n12117), .ZN(n12127) );
  AND2_X1 U11964 ( .A1(n12130), .A2(n12131), .ZN(n12117) );
  NAND3_X1 U11965 ( .A1(a_2_), .A2(n12132), .A3(b_17_), .ZN(n12131) );
  OR2_X1 U11966 ( .A1(n12113), .A2(n12111), .ZN(n12132) );
  NAND2_X1 U11967 ( .A1(n12111), .A2(n12113), .ZN(n12130) );
  NAND2_X1 U11968 ( .A1(n12133), .A2(n12134), .ZN(n12113) );
  NAND3_X1 U11969 ( .A1(a_3_), .A2(n12135), .A3(b_17_), .ZN(n12134) );
  NAND2_X1 U11970 ( .A1(n11908), .A2(n11907), .ZN(n12135) );
  OR2_X1 U11971 ( .A1(n11907), .A2(n11908), .ZN(n12133) );
  AND2_X1 U11972 ( .A1(n12136), .A2(n12137), .ZN(n11908) );
  NAND3_X1 U11973 ( .A1(a_4_), .A2(n12138), .A3(b_17_), .ZN(n12137) );
  OR2_X1 U11974 ( .A1(n11916), .A2(n11914), .ZN(n12138) );
  NAND2_X1 U11975 ( .A1(n11914), .A2(n11916), .ZN(n12136) );
  NAND2_X1 U11976 ( .A1(n12139), .A2(n12140), .ZN(n11916) );
  NAND3_X1 U11977 ( .A1(a_5_), .A2(n12141), .A3(b_17_), .ZN(n12140) );
  OR2_X1 U11978 ( .A1(n11924), .A2(n11922), .ZN(n12141) );
  NAND2_X1 U11979 ( .A1(n11922), .A2(n11924), .ZN(n12139) );
  NAND2_X1 U11980 ( .A1(n12142), .A2(n12143), .ZN(n11924) );
  NAND3_X1 U11981 ( .A1(a_6_), .A2(n12144), .A3(b_17_), .ZN(n12143) );
  OR2_X1 U11982 ( .A1(n11932), .A2(n11930), .ZN(n12144) );
  NAND2_X1 U11983 ( .A1(n11930), .A2(n11932), .ZN(n12142) );
  NAND2_X1 U11984 ( .A1(n12145), .A2(n12146), .ZN(n11932) );
  NAND3_X1 U11985 ( .A1(a_7_), .A2(n12147), .A3(b_17_), .ZN(n12146) );
  OR2_X1 U11986 ( .A1(n11940), .A2(n11938), .ZN(n12147) );
  NAND2_X1 U11987 ( .A1(n11938), .A2(n11940), .ZN(n12145) );
  NAND2_X1 U11988 ( .A1(n12148), .A2(n12149), .ZN(n11940) );
  NAND3_X1 U11989 ( .A1(a_8_), .A2(n12150), .A3(b_17_), .ZN(n12149) );
  OR2_X1 U11990 ( .A1(n11948), .A2(n11946), .ZN(n12150) );
  NAND2_X1 U11991 ( .A1(n11946), .A2(n11948), .ZN(n12148) );
  NAND2_X1 U11992 ( .A1(n12151), .A2(n12152), .ZN(n11948) );
  NAND3_X1 U11993 ( .A1(a_9_), .A2(n12153), .A3(b_17_), .ZN(n12152) );
  NAND2_X1 U11994 ( .A1(n11956), .A2(n11955), .ZN(n12153) );
  OR2_X1 U11995 ( .A1(n11955), .A2(n11956), .ZN(n12151) );
  AND2_X1 U11996 ( .A1(n12154), .A2(n12155), .ZN(n11956) );
  NAND3_X1 U11997 ( .A1(a_10_), .A2(n12156), .A3(b_17_), .ZN(n12155) );
  NAND2_X1 U11998 ( .A1(n11964), .A2(n11963), .ZN(n12156) );
  OR2_X1 U11999 ( .A1(n11963), .A2(n11964), .ZN(n12154) );
  AND2_X1 U12000 ( .A1(n12157), .A2(n12158), .ZN(n11964) );
  NAND3_X1 U12001 ( .A1(a_11_), .A2(n12159), .A3(b_17_), .ZN(n12158) );
  OR2_X1 U12002 ( .A1(n12109), .A2(n12107), .ZN(n12159) );
  NAND2_X1 U12003 ( .A1(n12107), .A2(n12109), .ZN(n12157) );
  NAND2_X1 U12004 ( .A1(n12160), .A2(n12161), .ZN(n12109) );
  NAND3_X1 U12005 ( .A1(a_12_), .A2(n12162), .A3(b_17_), .ZN(n12161) );
  OR2_X1 U12006 ( .A1(n12105), .A2(n12103), .ZN(n12162) );
  NAND2_X1 U12007 ( .A1(n12103), .A2(n12105), .ZN(n12160) );
  NAND2_X1 U12008 ( .A1(n12163), .A2(n12164), .ZN(n12105) );
  NAND3_X1 U12009 ( .A1(a_13_), .A2(n12165), .A3(b_17_), .ZN(n12164) );
  NAND2_X1 U12010 ( .A1(n12101), .A2(n12100), .ZN(n12165) );
  OR2_X1 U12011 ( .A1(n12100), .A2(n12101), .ZN(n12163) );
  AND2_X1 U12012 ( .A1(n12166), .A2(n12167), .ZN(n12101) );
  NAND2_X1 U12013 ( .A1(n12098), .A2(n12168), .ZN(n12167) );
  OR2_X1 U12014 ( .A1(n12097), .A2(n12096), .ZN(n12168) );
  NOR2_X1 U12015 ( .A1(n8754), .A2(n8757), .ZN(n12098) );
  NAND2_X1 U12016 ( .A1(n12096), .A2(n12097), .ZN(n12166) );
  NAND2_X1 U12017 ( .A1(n12169), .A2(n12170), .ZN(n12097) );
  NAND2_X1 U12018 ( .A1(n12094), .A2(n12171), .ZN(n12170) );
  OR2_X1 U12019 ( .A1(n12093), .A2(n12091), .ZN(n12171) );
  NOR2_X1 U12020 ( .A1(n8754), .A2(n8276), .ZN(n12094) );
  NAND2_X1 U12021 ( .A1(n12091), .A2(n12093), .ZN(n12169) );
  NAND2_X1 U12022 ( .A1(n12172), .A2(n12173), .ZN(n12093) );
  NAND3_X1 U12023 ( .A1(a_16_), .A2(n12174), .A3(b_17_), .ZN(n12173) );
  OR2_X1 U12024 ( .A1(n12089), .A2(n12087), .ZN(n12174) );
  NAND2_X1 U12025 ( .A1(n12087), .A2(n12089), .ZN(n12172) );
  NAND2_X1 U12026 ( .A1(n12175), .A2(n12176), .ZN(n12089) );
  NAND2_X1 U12027 ( .A1(n12086), .A2(n12177), .ZN(n12176) );
  OR2_X1 U12028 ( .A1(n12085), .A2(n12084), .ZN(n12177) );
  INV_X1 U12029 ( .A(n8706), .ZN(n12086) );
  NAND2_X1 U12030 ( .A1(b_17_), .A2(a_17_), .ZN(n8706) );
  NAND2_X1 U12031 ( .A1(n12084), .A2(n12085), .ZN(n12175) );
  NAND2_X1 U12032 ( .A1(n12178), .A2(n12179), .ZN(n12085) );
  NAND3_X1 U12033 ( .A1(a_18_), .A2(n12180), .A3(b_17_), .ZN(n12179) );
  NAND2_X1 U12034 ( .A1(n12081), .A2(n12080), .ZN(n12180) );
  OR2_X1 U12035 ( .A1(n12080), .A2(n12081), .ZN(n12178) );
  AND2_X1 U12036 ( .A1(n12181), .A2(n12182), .ZN(n12081) );
  NAND2_X1 U12037 ( .A1(n11996), .A2(n12183), .ZN(n12182) );
  OR2_X1 U12038 ( .A1(n11995), .A2(n11993), .ZN(n12183) );
  NOR2_X1 U12039 ( .A1(n8754), .A2(n8170), .ZN(n11996) );
  NAND2_X1 U12040 ( .A1(n11993), .A2(n11995), .ZN(n12181) );
  NAND2_X1 U12041 ( .A1(n12184), .A2(n12185), .ZN(n11995) );
  NAND3_X1 U12042 ( .A1(a_20_), .A2(n12186), .A3(b_17_), .ZN(n12185) );
  NAND2_X1 U12043 ( .A1(n12077), .A2(n12076), .ZN(n12186) );
  OR2_X1 U12044 ( .A1(n12076), .A2(n12077), .ZN(n12184) );
  AND2_X1 U12045 ( .A1(n12187), .A2(n12188), .ZN(n12077) );
  NAND2_X1 U12046 ( .A1(n12074), .A2(n12189), .ZN(n12188) );
  OR2_X1 U12047 ( .A1(n12073), .A2(n12072), .ZN(n12189) );
  NOR2_X1 U12048 ( .A1(n8754), .A2(n8750), .ZN(n12074) );
  NAND2_X1 U12049 ( .A1(n12072), .A2(n12073), .ZN(n12187) );
  NAND2_X1 U12050 ( .A1(n12190), .A2(n12191), .ZN(n12073) );
  NAND3_X1 U12051 ( .A1(a_22_), .A2(n12192), .A3(b_17_), .ZN(n12191) );
  OR2_X1 U12052 ( .A1(n12069), .A2(n12067), .ZN(n12192) );
  NAND2_X1 U12053 ( .A1(n12067), .A2(n12069), .ZN(n12190) );
  NAND2_X1 U12054 ( .A1(n12193), .A2(n12194), .ZN(n12069) );
  NAND2_X1 U12055 ( .A1(n12013), .A2(n12195), .ZN(n12194) );
  OR2_X1 U12056 ( .A1(n12012), .A2(n12010), .ZN(n12195) );
  NOR2_X1 U12057 ( .A1(n8754), .A2(n8747), .ZN(n12013) );
  NAND2_X1 U12058 ( .A1(n12010), .A2(n12012), .ZN(n12193) );
  NAND2_X1 U12059 ( .A1(n12196), .A2(n12197), .ZN(n12012) );
  NAND3_X1 U12060 ( .A1(a_24_), .A2(n12198), .A3(b_17_), .ZN(n12197) );
  NAND2_X1 U12061 ( .A1(n12065), .A2(n12064), .ZN(n12198) );
  OR2_X1 U12062 ( .A1(n12064), .A2(n12065), .ZN(n12196) );
  AND2_X1 U12063 ( .A1(n12199), .A2(n12200), .ZN(n12065) );
  NAND2_X1 U12064 ( .A1(n12062), .A2(n12201), .ZN(n12200) );
  OR2_X1 U12065 ( .A1(n12061), .A2(n12060), .ZN(n12201) );
  NOR2_X1 U12066 ( .A1(n8754), .A2(n8744), .ZN(n12062) );
  NAND2_X1 U12067 ( .A1(n12060), .A2(n12061), .ZN(n12199) );
  NAND2_X1 U12068 ( .A1(n12057), .A2(n12202), .ZN(n12061) );
  NAND2_X1 U12069 ( .A1(n12056), .A2(n12058), .ZN(n12202) );
  NAND2_X1 U12070 ( .A1(n12203), .A2(n12204), .ZN(n12058) );
  NAND2_X1 U12071 ( .A1(b_17_), .A2(a_26_), .ZN(n12204) );
  INV_X1 U12072 ( .A(n12205), .ZN(n12203) );
  XNOR2_X1 U12073 ( .A(n12206), .B(n12207), .ZN(n12056) );
  NAND2_X1 U12074 ( .A1(n12208), .A2(n12209), .ZN(n12206) );
  NAND2_X1 U12075 ( .A1(a_26_), .A2(n12205), .ZN(n12057) );
  NAND2_X1 U12076 ( .A1(n12029), .A2(n12210), .ZN(n12205) );
  NAND2_X1 U12077 ( .A1(n12028), .A2(n12030), .ZN(n12210) );
  NAND2_X1 U12078 ( .A1(n12211), .A2(n12212), .ZN(n12030) );
  NAND2_X1 U12079 ( .A1(b_17_), .A2(a_27_), .ZN(n12212) );
  INV_X1 U12080 ( .A(n12213), .ZN(n12211) );
  XNOR2_X1 U12081 ( .A(n12214), .B(n12215), .ZN(n12028) );
  XOR2_X1 U12082 ( .A(n12216), .B(n12217), .Z(n12214) );
  NAND2_X1 U12083 ( .A1(b_16_), .A2(a_28_), .ZN(n12216) );
  NAND2_X1 U12084 ( .A1(a_27_), .A2(n12213), .ZN(n12029) );
  NAND2_X1 U12085 ( .A1(n12218), .A2(n12219), .ZN(n12213) );
  NAND3_X1 U12086 ( .A1(a_28_), .A2(n12220), .A3(b_17_), .ZN(n12219) );
  NAND2_X1 U12087 ( .A1(n12038), .A2(n12036), .ZN(n12220) );
  OR2_X1 U12088 ( .A1(n12036), .A2(n12038), .ZN(n12218) );
  AND2_X1 U12089 ( .A1(n12221), .A2(n12222), .ZN(n12038) );
  NAND2_X1 U12090 ( .A1(n12052), .A2(n12223), .ZN(n12222) );
  OR2_X1 U12091 ( .A1(n12053), .A2(n12054), .ZN(n12223) );
  NOR2_X1 U12092 ( .A1(n8754), .A2(n7890), .ZN(n12052) );
  NAND2_X1 U12093 ( .A1(n12054), .A2(n12053), .ZN(n12221) );
  NAND2_X1 U12094 ( .A1(n12224), .A2(n12225), .ZN(n12053) );
  NAND2_X1 U12095 ( .A1(b_15_), .A2(n12226), .ZN(n12225) );
  NAND2_X1 U12096 ( .A1(n7864), .A2(n12227), .ZN(n12226) );
  NAND2_X1 U12097 ( .A1(a_31_), .A2(n8251), .ZN(n12227) );
  NAND2_X1 U12098 ( .A1(b_16_), .A2(n12228), .ZN(n12224) );
  NAND2_X1 U12099 ( .A1(n9137), .A2(n12229), .ZN(n12228) );
  NAND2_X1 U12100 ( .A1(a_30_), .A2(n8756), .ZN(n12229) );
  AND3_X1 U12101 ( .A1(b_16_), .A2(b_17_), .A3(n7818), .ZN(n12054) );
  XNOR2_X1 U12102 ( .A(n12230), .B(n12231), .ZN(n12036) );
  XOR2_X1 U12103 ( .A(n12232), .B(n12233), .Z(n12230) );
  XNOR2_X1 U12104 ( .A(n12234), .B(n12235), .ZN(n12060) );
  NAND2_X1 U12105 ( .A1(n12236), .A2(n12237), .ZN(n12234) );
  XNOR2_X1 U12106 ( .A(n12238), .B(n12239), .ZN(n12064) );
  XOR2_X1 U12107 ( .A(n12240), .B(n12241), .Z(n12238) );
  XNOR2_X1 U12108 ( .A(n12242), .B(n12243), .ZN(n12010) );
  XNOR2_X1 U12109 ( .A(n12244), .B(n12245), .ZN(n12242) );
  NOR2_X1 U12110 ( .A1(n8745), .A2(n8251), .ZN(n12245) );
  XNOR2_X1 U12111 ( .A(n12246), .B(n12247), .ZN(n12067) );
  XNOR2_X1 U12112 ( .A(n12248), .B(n12249), .ZN(n12247) );
  XNOR2_X1 U12113 ( .A(n12250), .B(n12251), .ZN(n12072) );
  XNOR2_X1 U12114 ( .A(n12252), .B(n12253), .ZN(n12250) );
  NOR2_X1 U12115 ( .A1(n8748), .A2(n8251), .ZN(n12253) );
  XNOR2_X1 U12116 ( .A(n12254), .B(n12255), .ZN(n12076) );
  XOR2_X1 U12117 ( .A(n12256), .B(n12257), .Z(n12254) );
  XNOR2_X1 U12118 ( .A(n12258), .B(n12259), .ZN(n11993) );
  XNOR2_X1 U12119 ( .A(n12260), .B(n12261), .ZN(n12258) );
  NOR2_X1 U12120 ( .A1(n8751), .A2(n8251), .ZN(n12261) );
  XOR2_X1 U12121 ( .A(n12262), .B(n12263), .Z(n12080) );
  XNOR2_X1 U12122 ( .A(n12264), .B(n12265), .ZN(n12263) );
  XNOR2_X1 U12123 ( .A(n12266), .B(n12267), .ZN(n12084) );
  XNOR2_X1 U12124 ( .A(n12268), .B(n12269), .ZN(n12266) );
  NOR2_X1 U12125 ( .A1(n8753), .A2(n8251), .ZN(n12269) );
  XOR2_X1 U12126 ( .A(n12270), .B(n12271), .Z(n12087) );
  XOR2_X1 U12127 ( .A(n12272), .B(n12273), .Z(n12270) );
  XNOR2_X1 U12128 ( .A(n12274), .B(n12275), .ZN(n12091) );
  XNOR2_X1 U12129 ( .A(n12276), .B(n8703), .ZN(n12275) );
  XNOR2_X1 U12130 ( .A(n12277), .B(n12278), .ZN(n12096) );
  NAND2_X1 U12131 ( .A1(n12279), .A2(n12280), .ZN(n12277) );
  XNOR2_X1 U12132 ( .A(n12281), .B(n12282), .ZN(n12100) );
  XOR2_X1 U12133 ( .A(n12283), .B(n12284), .Z(n12281) );
  XNOR2_X1 U12134 ( .A(n12285), .B(n12286), .ZN(n12103) );
  XNOR2_X1 U12135 ( .A(n12287), .B(n12288), .ZN(n12285) );
  XNOR2_X1 U12136 ( .A(n12289), .B(n12290), .ZN(n12107) );
  XNOR2_X1 U12137 ( .A(n12291), .B(n12292), .ZN(n12289) );
  XNOR2_X1 U12138 ( .A(n12293), .B(n12294), .ZN(n11963) );
  XOR2_X1 U12139 ( .A(n12295), .B(n12296), .Z(n12293) );
  XNOR2_X1 U12140 ( .A(n12297), .B(n12298), .ZN(n11955) );
  XOR2_X1 U12141 ( .A(n12299), .B(n12300), .Z(n12297) );
  XNOR2_X1 U12142 ( .A(n12301), .B(n12302), .ZN(n11946) );
  XNOR2_X1 U12143 ( .A(n12303), .B(n12304), .ZN(n12302) );
  XNOR2_X1 U12144 ( .A(n12305), .B(n12306), .ZN(n11938) );
  XNOR2_X1 U12145 ( .A(n12307), .B(n12308), .ZN(n12305) );
  NOR2_X1 U12146 ( .A1(n8763), .A2(n8251), .ZN(n12308) );
  XNOR2_X1 U12147 ( .A(n12309), .B(n12310), .ZN(n11930) );
  XNOR2_X1 U12148 ( .A(n12311), .B(n12312), .ZN(n12310) );
  XNOR2_X1 U12149 ( .A(n12313), .B(n12314), .ZN(n11922) );
  XOR2_X1 U12150 ( .A(n12315), .B(n12316), .Z(n12314) );
  NAND2_X1 U12151 ( .A1(b_16_), .A2(a_6_), .ZN(n12316) );
  XNOR2_X1 U12152 ( .A(n12317), .B(n12318), .ZN(n11914) );
  NAND2_X1 U12153 ( .A1(n12319), .A2(n12320), .ZN(n12317) );
  XOR2_X1 U12154 ( .A(n12321), .B(n12322), .Z(n11907) );
  NAND2_X1 U12155 ( .A1(n12323), .A2(n12324), .ZN(n12321) );
  XNOR2_X1 U12156 ( .A(n12325), .B(n12326), .ZN(n12111) );
  XNOR2_X1 U12157 ( .A(n12327), .B(n12328), .ZN(n12326) );
  XOR2_X1 U12158 ( .A(n12329), .B(n12330), .Z(n12116) );
  XNOR2_X1 U12159 ( .A(n12331), .B(n12332), .ZN(n12330) );
  XNOR2_X1 U12160 ( .A(n12333), .B(n12334), .ZN(n12119) );
  XNOR2_X1 U12161 ( .A(n12335), .B(n12336), .ZN(n12333) );
  INV_X1 U12162 ( .A(n11894), .ZN(n8953) );
  XOR2_X1 U12163 ( .A(n12337), .B(n12338), .Z(n11894) );
  XOR2_X1 U12164 ( .A(n12339), .B(n12340), .Z(n12338) );
  NAND2_X1 U12165 ( .A1(b_16_), .A2(a_0_), .ZN(n12340) );
  NAND2_X1 U12166 ( .A1(n12341), .A2(n12342), .ZN(n8881) );
  NAND2_X1 U12167 ( .A1(n8955), .A2(n8956), .ZN(n12342) );
  XOR2_X1 U12168 ( .A(n12343), .B(n12344), .Z(n12341) );
  NAND3_X1 U12169 ( .A1(n8955), .A2(n8956), .A3(n12345), .ZN(n8882) );
  XOR2_X1 U12170 ( .A(n12343), .B(n12346), .Z(n12345) );
  NAND2_X1 U12171 ( .A1(n12347), .A2(n12348), .ZN(n8956) );
  NAND3_X1 U12172 ( .A1(a_0_), .A2(n12349), .A3(b_16_), .ZN(n12348) );
  OR2_X1 U12173 ( .A1(n12339), .A2(n12337), .ZN(n12349) );
  NAND2_X1 U12174 ( .A1(n12337), .A2(n12339), .ZN(n12347) );
  NAND2_X1 U12175 ( .A1(n12350), .A2(n12351), .ZN(n12339) );
  NAND2_X1 U12176 ( .A1(n12335), .A2(n12352), .ZN(n12351) );
  NAND2_X1 U12177 ( .A1(n12336), .A2(n12334), .ZN(n12352) );
  NOR2_X1 U12178 ( .A1(n8251), .A2(n8617), .ZN(n12335) );
  OR2_X1 U12179 ( .A1(n12334), .A2(n12336), .ZN(n12350) );
  AND2_X1 U12180 ( .A1(n12353), .A2(n12354), .ZN(n12336) );
  NAND2_X1 U12181 ( .A1(n12332), .A2(n12355), .ZN(n12354) );
  OR2_X1 U12182 ( .A1(n12329), .A2(n12331), .ZN(n12355) );
  NOR2_X1 U12183 ( .A1(n8251), .A2(n8768), .ZN(n12332) );
  NAND2_X1 U12184 ( .A1(n12329), .A2(n12331), .ZN(n12353) );
  NAND2_X1 U12185 ( .A1(n12356), .A2(n12357), .ZN(n12331) );
  NAND2_X1 U12186 ( .A1(n12328), .A2(n12358), .ZN(n12357) );
  OR2_X1 U12187 ( .A1(n12325), .A2(n12327), .ZN(n12358) );
  NOR2_X1 U12188 ( .A1(n8251), .A2(n8567), .ZN(n12328) );
  NAND2_X1 U12189 ( .A1(n12325), .A2(n12327), .ZN(n12356) );
  NAND2_X1 U12190 ( .A1(n12323), .A2(n12359), .ZN(n12327) );
  NAND2_X1 U12191 ( .A1(n12322), .A2(n12324), .ZN(n12359) );
  NAND2_X1 U12192 ( .A1(n12360), .A2(n12361), .ZN(n12324) );
  NAND2_X1 U12193 ( .A1(b_16_), .A2(a_4_), .ZN(n12361) );
  INV_X1 U12194 ( .A(n12362), .ZN(n12360) );
  XNOR2_X1 U12195 ( .A(n12363), .B(n12364), .ZN(n12322) );
  XOR2_X1 U12196 ( .A(n12365), .B(n12366), .Z(n12364) );
  NAND2_X1 U12197 ( .A1(b_15_), .A2(a_5_), .ZN(n12366) );
  NAND2_X1 U12198 ( .A1(a_4_), .A2(n12362), .ZN(n12323) );
  NAND2_X1 U12199 ( .A1(n12319), .A2(n12367), .ZN(n12362) );
  NAND2_X1 U12200 ( .A1(n12318), .A2(n12320), .ZN(n12367) );
  NAND2_X1 U12201 ( .A1(n12368), .A2(n12369), .ZN(n12320) );
  NAND2_X1 U12202 ( .A1(b_16_), .A2(a_5_), .ZN(n12369) );
  INV_X1 U12203 ( .A(n12370), .ZN(n12368) );
  XNOR2_X1 U12204 ( .A(n12371), .B(n12372), .ZN(n12318) );
  XNOR2_X1 U12205 ( .A(n12373), .B(n12374), .ZN(n12371) );
  NOR2_X1 U12206 ( .A1(n8491), .A2(n8756), .ZN(n12374) );
  NAND2_X1 U12207 ( .A1(a_5_), .A2(n12370), .ZN(n12319) );
  NAND2_X1 U12208 ( .A1(n12375), .A2(n12376), .ZN(n12370) );
  NAND3_X1 U12209 ( .A1(a_6_), .A2(n12377), .A3(b_16_), .ZN(n12376) );
  OR2_X1 U12210 ( .A1(n12313), .A2(n12315), .ZN(n12377) );
  NAND2_X1 U12211 ( .A1(n12313), .A2(n12315), .ZN(n12375) );
  NAND2_X1 U12212 ( .A1(n12378), .A2(n12379), .ZN(n12315) );
  NAND2_X1 U12213 ( .A1(n12312), .A2(n12380), .ZN(n12379) );
  OR2_X1 U12214 ( .A1(n12309), .A2(n12311), .ZN(n12380) );
  NOR2_X1 U12215 ( .A1(n8251), .A2(n8764), .ZN(n12312) );
  NAND2_X1 U12216 ( .A1(n12309), .A2(n12311), .ZN(n12378) );
  NAND2_X1 U12217 ( .A1(n12381), .A2(n12382), .ZN(n12311) );
  NAND3_X1 U12218 ( .A1(a_8_), .A2(n12383), .A3(b_16_), .ZN(n12382) );
  NAND2_X1 U12219 ( .A1(n12307), .A2(n12306), .ZN(n12383) );
  OR2_X1 U12220 ( .A1(n12306), .A2(n12307), .ZN(n12381) );
  AND2_X1 U12221 ( .A1(n12384), .A2(n12385), .ZN(n12307) );
  NAND2_X1 U12222 ( .A1(n12304), .A2(n12386), .ZN(n12385) );
  OR2_X1 U12223 ( .A1(n12303), .A2(n12301), .ZN(n12386) );
  NOR2_X1 U12224 ( .A1(n8251), .A2(n8426), .ZN(n12304) );
  NAND2_X1 U12225 ( .A1(n12301), .A2(n12303), .ZN(n12384) );
  NAND2_X1 U12226 ( .A1(n12387), .A2(n12388), .ZN(n12303) );
  NAND2_X1 U12227 ( .A1(n12300), .A2(n12389), .ZN(n12388) );
  OR2_X1 U12228 ( .A1(n12298), .A2(n12299), .ZN(n12389) );
  NOR2_X1 U12229 ( .A1(n8251), .A2(n8761), .ZN(n12300) );
  NAND2_X1 U12230 ( .A1(n12298), .A2(n12299), .ZN(n12387) );
  NAND2_X1 U12231 ( .A1(n12390), .A2(n12391), .ZN(n12299) );
  NAND2_X1 U12232 ( .A1(n12296), .A2(n12392), .ZN(n12391) );
  OR2_X1 U12233 ( .A1(n12294), .A2(n12295), .ZN(n12392) );
  NOR2_X1 U12234 ( .A1(n8251), .A2(n8376), .ZN(n12296) );
  NAND2_X1 U12235 ( .A1(n12294), .A2(n12295), .ZN(n12390) );
  NAND2_X1 U12236 ( .A1(n12393), .A2(n12394), .ZN(n12295) );
  NAND2_X1 U12237 ( .A1(n12292), .A2(n12395), .ZN(n12394) );
  NAND2_X1 U12238 ( .A1(n12291), .A2(n12290), .ZN(n12395) );
  NOR2_X1 U12239 ( .A1(n8251), .A2(n8759), .ZN(n12292) );
  OR2_X1 U12240 ( .A1(n12290), .A2(n12291), .ZN(n12393) );
  AND2_X1 U12241 ( .A1(n12396), .A2(n12397), .ZN(n12291) );
  NAND2_X1 U12242 ( .A1(n12288), .A2(n12398), .ZN(n12397) );
  NAND2_X1 U12243 ( .A1(n12287), .A2(n12286), .ZN(n12398) );
  NOR2_X1 U12244 ( .A1(n8251), .A2(n8310), .ZN(n12288) );
  OR2_X1 U12245 ( .A1(n12286), .A2(n12287), .ZN(n12396) );
  AND2_X1 U12246 ( .A1(n12399), .A2(n12400), .ZN(n12287) );
  NAND2_X1 U12247 ( .A1(n12284), .A2(n12401), .ZN(n12400) );
  OR2_X1 U12248 ( .A1(n12282), .A2(n12283), .ZN(n12401) );
  NOR2_X1 U12249 ( .A1(n8251), .A2(n8757), .ZN(n12284) );
  NAND2_X1 U12250 ( .A1(n12282), .A2(n12283), .ZN(n12399) );
  NAND2_X1 U12251 ( .A1(n12279), .A2(n12402), .ZN(n12283) );
  NAND2_X1 U12252 ( .A1(n12278), .A2(n12280), .ZN(n12402) );
  NAND2_X1 U12253 ( .A1(n12403), .A2(n12404), .ZN(n12280) );
  NAND2_X1 U12254 ( .A1(b_16_), .A2(a_15_), .ZN(n12404) );
  INV_X1 U12255 ( .A(n12405), .ZN(n12403) );
  XNOR2_X1 U12256 ( .A(n12406), .B(n12407), .ZN(n12278) );
  XOR2_X1 U12257 ( .A(n12408), .B(n12409), .Z(n12407) );
  NAND2_X1 U12258 ( .A1(b_15_), .A2(a_16_), .ZN(n12409) );
  NAND2_X1 U12259 ( .A1(a_15_), .A2(n12405), .ZN(n12279) );
  NAND2_X1 U12260 ( .A1(n12410), .A2(n12411), .ZN(n12405) );
  NAND2_X1 U12261 ( .A1(n12274), .A2(n12412), .ZN(n12411) );
  OR2_X1 U12262 ( .A1(n12276), .A2(n8703), .ZN(n12412) );
  XOR2_X1 U12263 ( .A(n12413), .B(n12414), .Z(n12274) );
  XOR2_X1 U12264 ( .A(n12415), .B(n12416), .Z(n12413) );
  NAND2_X1 U12265 ( .A1(n8703), .A2(n12276), .ZN(n12410) );
  NAND2_X1 U12266 ( .A1(n12417), .A2(n12418), .ZN(n12276) );
  NAND2_X1 U12267 ( .A1(n12273), .A2(n12419), .ZN(n12418) );
  OR2_X1 U12268 ( .A1(n12271), .A2(n12272), .ZN(n12419) );
  NOR2_X1 U12269 ( .A1(n8251), .A2(n8210), .ZN(n12273) );
  NAND2_X1 U12270 ( .A1(n12271), .A2(n12272), .ZN(n12417) );
  NAND2_X1 U12271 ( .A1(n12420), .A2(n12421), .ZN(n12272) );
  NAND3_X1 U12272 ( .A1(a_18_), .A2(n12422), .A3(b_16_), .ZN(n12421) );
  NAND2_X1 U12273 ( .A1(n12268), .A2(n12267), .ZN(n12422) );
  OR2_X1 U12274 ( .A1(n12267), .A2(n12268), .ZN(n12420) );
  AND2_X1 U12275 ( .A1(n12423), .A2(n12424), .ZN(n12268) );
  NAND2_X1 U12276 ( .A1(n12265), .A2(n12425), .ZN(n12424) );
  OR2_X1 U12277 ( .A1(n12262), .A2(n12264), .ZN(n12425) );
  NOR2_X1 U12278 ( .A1(n8251), .A2(n8170), .ZN(n12265) );
  NAND2_X1 U12279 ( .A1(n12262), .A2(n12264), .ZN(n12423) );
  NAND2_X1 U12280 ( .A1(n12426), .A2(n12427), .ZN(n12264) );
  NAND3_X1 U12281 ( .A1(a_20_), .A2(n12428), .A3(b_16_), .ZN(n12427) );
  NAND2_X1 U12282 ( .A1(n12260), .A2(n12259), .ZN(n12428) );
  OR2_X1 U12283 ( .A1(n12259), .A2(n12260), .ZN(n12426) );
  AND2_X1 U12284 ( .A1(n12429), .A2(n12430), .ZN(n12260) );
  NAND2_X1 U12285 ( .A1(n12257), .A2(n12431), .ZN(n12430) );
  OR2_X1 U12286 ( .A1(n12255), .A2(n12256), .ZN(n12431) );
  NOR2_X1 U12287 ( .A1(n8251), .A2(n8750), .ZN(n12257) );
  NAND2_X1 U12288 ( .A1(n12255), .A2(n12256), .ZN(n12429) );
  NAND2_X1 U12289 ( .A1(n12432), .A2(n12433), .ZN(n12256) );
  NAND3_X1 U12290 ( .A1(a_22_), .A2(n12434), .A3(b_16_), .ZN(n12433) );
  NAND2_X1 U12291 ( .A1(n12252), .A2(n12251), .ZN(n12434) );
  OR2_X1 U12292 ( .A1(n12251), .A2(n12252), .ZN(n12432) );
  AND2_X1 U12293 ( .A1(n12435), .A2(n12436), .ZN(n12252) );
  NAND2_X1 U12294 ( .A1(n12249), .A2(n12437), .ZN(n12436) );
  OR2_X1 U12295 ( .A1(n12246), .A2(n12248), .ZN(n12437) );
  NOR2_X1 U12296 ( .A1(n8251), .A2(n8747), .ZN(n12249) );
  NAND2_X1 U12297 ( .A1(n12246), .A2(n12248), .ZN(n12435) );
  NAND2_X1 U12298 ( .A1(n12438), .A2(n12439), .ZN(n12248) );
  NAND3_X1 U12299 ( .A1(a_24_), .A2(n12440), .A3(b_16_), .ZN(n12439) );
  NAND2_X1 U12300 ( .A1(n12244), .A2(n12243), .ZN(n12440) );
  OR2_X1 U12301 ( .A1(n12243), .A2(n12244), .ZN(n12438) );
  AND2_X1 U12302 ( .A1(n12441), .A2(n12442), .ZN(n12244) );
  NAND2_X1 U12303 ( .A1(n12241), .A2(n12443), .ZN(n12442) );
  OR2_X1 U12304 ( .A1(n12239), .A2(n12240), .ZN(n12443) );
  NOR2_X1 U12305 ( .A1(n8251), .A2(n8744), .ZN(n12241) );
  NAND2_X1 U12306 ( .A1(n12239), .A2(n12240), .ZN(n12441) );
  NAND2_X1 U12307 ( .A1(n12236), .A2(n12444), .ZN(n12240) );
  NAND2_X1 U12308 ( .A1(n12235), .A2(n12237), .ZN(n12444) );
  NAND2_X1 U12309 ( .A1(n12445), .A2(n12446), .ZN(n12237) );
  NAND2_X1 U12310 ( .A1(b_16_), .A2(a_26_), .ZN(n12446) );
  INV_X1 U12311 ( .A(n12447), .ZN(n12445) );
  XNOR2_X1 U12312 ( .A(n12448), .B(n12449), .ZN(n12235) );
  NAND2_X1 U12313 ( .A1(n12450), .A2(n12451), .ZN(n12448) );
  NAND2_X1 U12314 ( .A1(a_26_), .A2(n12447), .ZN(n12236) );
  NAND2_X1 U12315 ( .A1(n12208), .A2(n12452), .ZN(n12447) );
  NAND2_X1 U12316 ( .A1(n12207), .A2(n12209), .ZN(n12452) );
  NAND2_X1 U12317 ( .A1(n12453), .A2(n12454), .ZN(n12209) );
  NAND2_X1 U12318 ( .A1(b_16_), .A2(a_27_), .ZN(n12454) );
  INV_X1 U12319 ( .A(n12455), .ZN(n12453) );
  XNOR2_X1 U12320 ( .A(n12456), .B(n12457), .ZN(n12207) );
  XOR2_X1 U12321 ( .A(n12458), .B(n12459), .Z(n12456) );
  NAND2_X1 U12322 ( .A1(b_15_), .A2(a_28_), .ZN(n12458) );
  NAND2_X1 U12323 ( .A1(a_27_), .A2(n12455), .ZN(n12208) );
  NAND2_X1 U12324 ( .A1(n12460), .A2(n12461), .ZN(n12455) );
  NAND3_X1 U12325 ( .A1(a_28_), .A2(n12462), .A3(b_16_), .ZN(n12461) );
  NAND2_X1 U12326 ( .A1(n12217), .A2(n12215), .ZN(n12462) );
  OR2_X1 U12327 ( .A1(n12215), .A2(n12217), .ZN(n12460) );
  AND2_X1 U12328 ( .A1(n12463), .A2(n12464), .ZN(n12217) );
  NAND2_X1 U12329 ( .A1(n12231), .A2(n12465), .ZN(n12464) );
  OR2_X1 U12330 ( .A1(n12232), .A2(n12233), .ZN(n12465) );
  NOR2_X1 U12331 ( .A1(n8251), .A2(n7890), .ZN(n12231) );
  NAND2_X1 U12332 ( .A1(n12233), .A2(n12232), .ZN(n12463) );
  NAND2_X1 U12333 ( .A1(n12466), .A2(n12467), .ZN(n12232) );
  NAND2_X1 U12334 ( .A1(b_14_), .A2(n12468), .ZN(n12467) );
  NAND2_X1 U12335 ( .A1(n7864), .A2(n12469), .ZN(n12468) );
  NAND2_X1 U12336 ( .A1(a_31_), .A2(n8756), .ZN(n12469) );
  NAND2_X1 U12337 ( .A1(b_15_), .A2(n12470), .ZN(n12466) );
  NAND2_X1 U12338 ( .A1(n9137), .A2(n12471), .ZN(n12470) );
  NAND2_X1 U12339 ( .A1(a_30_), .A2(n8301), .ZN(n12471) );
  AND3_X1 U12340 ( .A1(b_15_), .A2(b_16_), .A3(n7818), .ZN(n12233) );
  XNOR2_X1 U12341 ( .A(n12472), .B(n12473), .ZN(n12215) );
  XOR2_X1 U12342 ( .A(n12474), .B(n12475), .Z(n12472) );
  XNOR2_X1 U12343 ( .A(n12476), .B(n12477), .ZN(n12239) );
  NAND2_X1 U12344 ( .A1(n12478), .A2(n12479), .ZN(n12476) );
  XNOR2_X1 U12345 ( .A(n12480), .B(n12481), .ZN(n12243) );
  XOR2_X1 U12346 ( .A(n12482), .B(n12483), .Z(n12480) );
  XNOR2_X1 U12347 ( .A(n12484), .B(n12485), .ZN(n12246) );
  XNOR2_X1 U12348 ( .A(n12486), .B(n12487), .ZN(n12484) );
  NOR2_X1 U12349 ( .A1(n8745), .A2(n8756), .ZN(n12487) );
  XOR2_X1 U12350 ( .A(n12488), .B(n12489), .Z(n12251) );
  XNOR2_X1 U12351 ( .A(n12490), .B(n12491), .ZN(n12489) );
  XNOR2_X1 U12352 ( .A(n12492), .B(n12493), .ZN(n12255) );
  XNOR2_X1 U12353 ( .A(n12494), .B(n12495), .ZN(n12492) );
  NOR2_X1 U12354 ( .A1(n8748), .A2(n8756), .ZN(n12495) );
  XNOR2_X1 U12355 ( .A(n12496), .B(n12497), .ZN(n12259) );
  XOR2_X1 U12356 ( .A(n12498), .B(n12499), .Z(n12496) );
  XNOR2_X1 U12357 ( .A(n12500), .B(n12501), .ZN(n12262) );
  XNOR2_X1 U12358 ( .A(n12502), .B(n12503), .ZN(n12500) );
  NOR2_X1 U12359 ( .A1(n8751), .A2(n8756), .ZN(n12503) );
  XOR2_X1 U12360 ( .A(n12504), .B(n12505), .Z(n12267) );
  XNOR2_X1 U12361 ( .A(n12506), .B(n12507), .ZN(n12505) );
  XNOR2_X1 U12362 ( .A(n12508), .B(n12509), .ZN(n12271) );
  XNOR2_X1 U12363 ( .A(n12510), .B(n12511), .ZN(n12508) );
  NOR2_X1 U12364 ( .A1(n8753), .A2(n8756), .ZN(n12511) );
  NOR2_X1 U12365 ( .A1(n8251), .A2(n8755), .ZN(n8703) );
  XNOR2_X1 U12366 ( .A(n12512), .B(n12513), .ZN(n12282) );
  XNOR2_X1 U12367 ( .A(n8700), .B(n12514), .ZN(n12513) );
  XOR2_X1 U12368 ( .A(n12515), .B(n12516), .Z(n12286) );
  NAND2_X1 U12369 ( .A1(n12517), .A2(n12518), .ZN(n12515) );
  XOR2_X1 U12370 ( .A(n12519), .B(n12520), .Z(n12290) );
  XOR2_X1 U12371 ( .A(n12521), .B(n12522), .Z(n12520) );
  NAND2_X1 U12372 ( .A1(b_15_), .A2(a_13_), .ZN(n12522) );
  XNOR2_X1 U12373 ( .A(n12523), .B(n12524), .ZN(n12294) );
  XOR2_X1 U12374 ( .A(n12525), .B(n12526), .Z(n12524) );
  NAND2_X1 U12375 ( .A1(b_15_), .A2(a_12_), .ZN(n12526) );
  XNOR2_X1 U12376 ( .A(n12527), .B(n12528), .ZN(n12298) );
  XNOR2_X1 U12377 ( .A(n12529), .B(n12530), .ZN(n12527) );
  NOR2_X1 U12378 ( .A1(n8376), .A2(n8756), .ZN(n12530) );
  XNOR2_X1 U12379 ( .A(n12531), .B(n12532), .ZN(n12301) );
  XOR2_X1 U12380 ( .A(n12533), .B(n12534), .Z(n12532) );
  NAND2_X1 U12381 ( .A1(b_15_), .A2(a_10_), .ZN(n12534) );
  XOR2_X1 U12382 ( .A(n12535), .B(n12536), .Z(n12306) );
  XOR2_X1 U12383 ( .A(n12537), .B(n12538), .Z(n12536) );
  NAND2_X1 U12384 ( .A1(b_15_), .A2(a_9_), .ZN(n12538) );
  XNOR2_X1 U12385 ( .A(n12539), .B(n12540), .ZN(n12309) );
  XNOR2_X1 U12386 ( .A(n12541), .B(n12542), .ZN(n12539) );
  NOR2_X1 U12387 ( .A1(n8763), .A2(n8756), .ZN(n12542) );
  XNOR2_X1 U12388 ( .A(n12543), .B(n12544), .ZN(n12313) );
  XOR2_X1 U12389 ( .A(n12545), .B(n12546), .Z(n12544) );
  NAND2_X1 U12390 ( .A1(b_15_), .A2(a_7_), .ZN(n12546) );
  XNOR2_X1 U12391 ( .A(n12547), .B(n12548), .ZN(n12325) );
  XNOR2_X1 U12392 ( .A(n12549), .B(n12550), .ZN(n12547) );
  NOR2_X1 U12393 ( .A1(n8766), .A2(n8756), .ZN(n12550) );
  XNOR2_X1 U12394 ( .A(n12551), .B(n12552), .ZN(n12329) );
  XOR2_X1 U12395 ( .A(n12553), .B(n12554), .Z(n12552) );
  NAND2_X1 U12396 ( .A1(b_15_), .A2(a_3_), .ZN(n12554) );
  XNOR2_X1 U12397 ( .A(n12555), .B(n12556), .ZN(n12334) );
  XOR2_X1 U12398 ( .A(n12557), .B(n12558), .Z(n12555) );
  NOR2_X1 U12399 ( .A1(n8768), .A2(n8756), .ZN(n12558) );
  XOR2_X1 U12400 ( .A(n12559), .B(n12560), .Z(n12337) );
  XOR2_X1 U12401 ( .A(n12561), .B(n12562), .Z(n12559) );
  NOR2_X1 U12402 ( .A1(n8617), .A2(n8756), .ZN(n12562) );
  XOR2_X1 U12403 ( .A(n12563), .B(n12564), .Z(n8955) );
  XOR2_X1 U12404 ( .A(n12565), .B(n12566), .Z(n12563) );
  NOR2_X1 U12405 ( .A1(n9674), .A2(n8756), .ZN(n12566) );
  NAND2_X1 U12406 ( .A1(n12567), .A2(n12568), .ZN(n8887) );
  NAND2_X1 U12407 ( .A1(n12346), .A2(n12343), .ZN(n12568) );
  XNOR2_X1 U12408 ( .A(n8947), .B(n8946), .ZN(n12567) );
  NAND3_X1 U12409 ( .A1(n12346), .A2(n12343), .A3(n12569), .ZN(n8888) );
  XOR2_X1 U12410 ( .A(n8947), .B(n8946), .Z(n12569) );
  NAND2_X1 U12411 ( .A1(n12570), .A2(n12571), .ZN(n12343) );
  NAND3_X1 U12412 ( .A1(a_0_), .A2(n12572), .A3(b_15_), .ZN(n12571) );
  OR2_X1 U12413 ( .A1(n12564), .A2(n12565), .ZN(n12572) );
  NAND2_X1 U12414 ( .A1(n12564), .A2(n12565), .ZN(n12570) );
  NAND2_X1 U12415 ( .A1(n12573), .A2(n12574), .ZN(n12565) );
  NAND3_X1 U12416 ( .A1(a_1_), .A2(n12575), .A3(b_15_), .ZN(n12574) );
  OR2_X1 U12417 ( .A1(n12560), .A2(n12561), .ZN(n12575) );
  NAND2_X1 U12418 ( .A1(n12560), .A2(n12561), .ZN(n12573) );
  NAND2_X1 U12419 ( .A1(n12576), .A2(n12577), .ZN(n12561) );
  NAND3_X1 U12420 ( .A1(a_2_), .A2(n12578), .A3(b_15_), .ZN(n12577) );
  OR2_X1 U12421 ( .A1(n12556), .A2(n12557), .ZN(n12578) );
  NAND2_X1 U12422 ( .A1(n12556), .A2(n12557), .ZN(n12576) );
  NAND2_X1 U12423 ( .A1(n12579), .A2(n12580), .ZN(n12557) );
  NAND3_X1 U12424 ( .A1(a_3_), .A2(n12581), .A3(b_15_), .ZN(n12580) );
  OR2_X1 U12425 ( .A1(n12553), .A2(n12551), .ZN(n12581) );
  NAND2_X1 U12426 ( .A1(n12551), .A2(n12553), .ZN(n12579) );
  NAND2_X1 U12427 ( .A1(n12582), .A2(n12583), .ZN(n12553) );
  NAND3_X1 U12428 ( .A1(a_4_), .A2(n12584), .A3(b_15_), .ZN(n12583) );
  NAND2_X1 U12429 ( .A1(n12549), .A2(n12548), .ZN(n12584) );
  OR2_X1 U12430 ( .A1(n12548), .A2(n12549), .ZN(n12582) );
  AND2_X1 U12431 ( .A1(n12585), .A2(n12586), .ZN(n12549) );
  NAND3_X1 U12432 ( .A1(a_5_), .A2(n12587), .A3(b_15_), .ZN(n12586) );
  OR2_X1 U12433 ( .A1(n12363), .A2(n12365), .ZN(n12587) );
  NAND2_X1 U12434 ( .A1(n12363), .A2(n12365), .ZN(n12585) );
  NAND2_X1 U12435 ( .A1(n12588), .A2(n12589), .ZN(n12365) );
  NAND3_X1 U12436 ( .A1(a_6_), .A2(n12590), .A3(b_15_), .ZN(n12589) );
  NAND2_X1 U12437 ( .A1(n12373), .A2(n12372), .ZN(n12590) );
  OR2_X1 U12438 ( .A1(n12372), .A2(n12373), .ZN(n12588) );
  AND2_X1 U12439 ( .A1(n12591), .A2(n12592), .ZN(n12373) );
  NAND3_X1 U12440 ( .A1(a_7_), .A2(n12593), .A3(b_15_), .ZN(n12592) );
  OR2_X1 U12441 ( .A1(n12545), .A2(n12543), .ZN(n12593) );
  NAND2_X1 U12442 ( .A1(n12543), .A2(n12545), .ZN(n12591) );
  NAND2_X1 U12443 ( .A1(n12594), .A2(n12595), .ZN(n12545) );
  NAND3_X1 U12444 ( .A1(a_8_), .A2(n12596), .A3(b_15_), .ZN(n12595) );
  NAND2_X1 U12445 ( .A1(n12541), .A2(n12540), .ZN(n12596) );
  OR2_X1 U12446 ( .A1(n12540), .A2(n12541), .ZN(n12594) );
  AND2_X1 U12447 ( .A1(n12597), .A2(n12598), .ZN(n12541) );
  NAND3_X1 U12448 ( .A1(a_9_), .A2(n12599), .A3(b_15_), .ZN(n12598) );
  OR2_X1 U12449 ( .A1(n12535), .A2(n12537), .ZN(n12599) );
  NAND2_X1 U12450 ( .A1(n12535), .A2(n12537), .ZN(n12597) );
  NAND2_X1 U12451 ( .A1(n12600), .A2(n12601), .ZN(n12537) );
  NAND3_X1 U12452 ( .A1(a_10_), .A2(n12602), .A3(b_15_), .ZN(n12601) );
  OR2_X1 U12453 ( .A1(n12531), .A2(n12533), .ZN(n12602) );
  NAND2_X1 U12454 ( .A1(n12531), .A2(n12533), .ZN(n12600) );
  NAND2_X1 U12455 ( .A1(n12603), .A2(n12604), .ZN(n12533) );
  NAND3_X1 U12456 ( .A1(a_11_), .A2(n12605), .A3(b_15_), .ZN(n12604) );
  NAND2_X1 U12457 ( .A1(n12529), .A2(n12528), .ZN(n12605) );
  OR2_X1 U12458 ( .A1(n12528), .A2(n12529), .ZN(n12603) );
  AND2_X1 U12459 ( .A1(n12606), .A2(n12607), .ZN(n12529) );
  NAND3_X1 U12460 ( .A1(a_12_), .A2(n12608), .A3(b_15_), .ZN(n12607) );
  OR2_X1 U12461 ( .A1(n12525), .A2(n12523), .ZN(n12608) );
  NAND2_X1 U12462 ( .A1(n12523), .A2(n12525), .ZN(n12606) );
  NAND2_X1 U12463 ( .A1(n12609), .A2(n12610), .ZN(n12525) );
  NAND3_X1 U12464 ( .A1(a_13_), .A2(n12611), .A3(b_15_), .ZN(n12610) );
  OR2_X1 U12465 ( .A1(n12519), .A2(n12521), .ZN(n12611) );
  NAND2_X1 U12466 ( .A1(n12519), .A2(n12521), .ZN(n12609) );
  NAND2_X1 U12467 ( .A1(n12517), .A2(n12612), .ZN(n12521) );
  NAND2_X1 U12468 ( .A1(n12516), .A2(n12518), .ZN(n12612) );
  NAND2_X1 U12469 ( .A1(n12613), .A2(n12614), .ZN(n12518) );
  NAND2_X1 U12470 ( .A1(b_15_), .A2(a_14_), .ZN(n12614) );
  INV_X1 U12471 ( .A(n12615), .ZN(n12613) );
  XOR2_X1 U12472 ( .A(n12616), .B(n12617), .Z(n12516) );
  XOR2_X1 U12473 ( .A(n12618), .B(n12619), .Z(n12616) );
  NAND2_X1 U12474 ( .A1(a_14_), .A2(n12615), .ZN(n12517) );
  NAND2_X1 U12475 ( .A1(n12620), .A2(n12621), .ZN(n12615) );
  NAND2_X1 U12476 ( .A1(n12512), .A2(n12622), .ZN(n12621) );
  OR2_X1 U12477 ( .A1(n12514), .A2(n8700), .ZN(n12622) );
  XNOR2_X1 U12478 ( .A(n12623), .B(n12624), .ZN(n12512) );
  XNOR2_X1 U12479 ( .A(n12625), .B(n12626), .ZN(n12624) );
  NAND2_X1 U12480 ( .A1(n8700), .A2(n12514), .ZN(n12620) );
  NAND2_X1 U12481 ( .A1(n12627), .A2(n12628), .ZN(n12514) );
  NAND3_X1 U12482 ( .A1(a_16_), .A2(n12629), .A3(b_15_), .ZN(n12628) );
  OR2_X1 U12483 ( .A1(n12408), .A2(n12406), .ZN(n12629) );
  NAND2_X1 U12484 ( .A1(n12406), .A2(n12408), .ZN(n12627) );
  NAND2_X1 U12485 ( .A1(n12630), .A2(n12631), .ZN(n12408) );
  NAND2_X1 U12486 ( .A1(n12416), .A2(n12632), .ZN(n12631) );
  OR2_X1 U12487 ( .A1(n12414), .A2(n12415), .ZN(n12632) );
  NOR2_X1 U12488 ( .A1(n8756), .A2(n8210), .ZN(n12416) );
  NAND2_X1 U12489 ( .A1(n12414), .A2(n12415), .ZN(n12630) );
  NAND2_X1 U12490 ( .A1(n12633), .A2(n12634), .ZN(n12415) );
  NAND3_X1 U12491 ( .A1(a_18_), .A2(n12635), .A3(b_15_), .ZN(n12634) );
  NAND2_X1 U12492 ( .A1(n12510), .A2(n12509), .ZN(n12635) );
  OR2_X1 U12493 ( .A1(n12509), .A2(n12510), .ZN(n12633) );
  AND2_X1 U12494 ( .A1(n12636), .A2(n12637), .ZN(n12510) );
  NAND2_X1 U12495 ( .A1(n12507), .A2(n12638), .ZN(n12637) );
  OR2_X1 U12496 ( .A1(n12504), .A2(n12506), .ZN(n12638) );
  NOR2_X1 U12497 ( .A1(n8756), .A2(n8170), .ZN(n12507) );
  NAND2_X1 U12498 ( .A1(n12504), .A2(n12506), .ZN(n12636) );
  NAND2_X1 U12499 ( .A1(n12639), .A2(n12640), .ZN(n12506) );
  NAND3_X1 U12500 ( .A1(a_20_), .A2(n12641), .A3(b_15_), .ZN(n12640) );
  NAND2_X1 U12501 ( .A1(n12502), .A2(n12501), .ZN(n12641) );
  OR2_X1 U12502 ( .A1(n12501), .A2(n12502), .ZN(n12639) );
  AND2_X1 U12503 ( .A1(n12642), .A2(n12643), .ZN(n12502) );
  NAND2_X1 U12504 ( .A1(n12499), .A2(n12644), .ZN(n12643) );
  OR2_X1 U12505 ( .A1(n12497), .A2(n12498), .ZN(n12644) );
  NOR2_X1 U12506 ( .A1(n8756), .A2(n8750), .ZN(n12499) );
  NAND2_X1 U12507 ( .A1(n12497), .A2(n12498), .ZN(n12642) );
  NAND2_X1 U12508 ( .A1(n12645), .A2(n12646), .ZN(n12498) );
  NAND3_X1 U12509 ( .A1(a_22_), .A2(n12647), .A3(b_15_), .ZN(n12646) );
  NAND2_X1 U12510 ( .A1(n12494), .A2(n12493), .ZN(n12647) );
  OR2_X1 U12511 ( .A1(n12493), .A2(n12494), .ZN(n12645) );
  AND2_X1 U12512 ( .A1(n12648), .A2(n12649), .ZN(n12494) );
  NAND2_X1 U12513 ( .A1(n12491), .A2(n12650), .ZN(n12649) );
  OR2_X1 U12514 ( .A1(n12488), .A2(n12490), .ZN(n12650) );
  NOR2_X1 U12515 ( .A1(n8756), .A2(n8747), .ZN(n12491) );
  NAND2_X1 U12516 ( .A1(n12488), .A2(n12490), .ZN(n12648) );
  NAND2_X1 U12517 ( .A1(n12651), .A2(n12652), .ZN(n12490) );
  NAND3_X1 U12518 ( .A1(a_24_), .A2(n12653), .A3(b_15_), .ZN(n12652) );
  NAND2_X1 U12519 ( .A1(n12486), .A2(n12485), .ZN(n12653) );
  OR2_X1 U12520 ( .A1(n12485), .A2(n12486), .ZN(n12651) );
  AND2_X1 U12521 ( .A1(n12654), .A2(n12655), .ZN(n12486) );
  NAND2_X1 U12522 ( .A1(n12483), .A2(n12656), .ZN(n12655) );
  OR2_X1 U12523 ( .A1(n12481), .A2(n12482), .ZN(n12656) );
  NOR2_X1 U12524 ( .A1(n8756), .A2(n8744), .ZN(n12483) );
  NAND2_X1 U12525 ( .A1(n12481), .A2(n12482), .ZN(n12654) );
  NAND2_X1 U12526 ( .A1(n12478), .A2(n12657), .ZN(n12482) );
  NAND2_X1 U12527 ( .A1(n12477), .A2(n12479), .ZN(n12657) );
  NAND2_X1 U12528 ( .A1(n12658), .A2(n12659), .ZN(n12479) );
  NAND2_X1 U12529 ( .A1(b_15_), .A2(a_26_), .ZN(n12659) );
  INV_X1 U12530 ( .A(n12660), .ZN(n12658) );
  XNOR2_X1 U12531 ( .A(n12661), .B(n12662), .ZN(n12477) );
  NAND2_X1 U12532 ( .A1(n12663), .A2(n12664), .ZN(n12661) );
  NAND2_X1 U12533 ( .A1(a_26_), .A2(n12660), .ZN(n12478) );
  NAND2_X1 U12534 ( .A1(n12450), .A2(n12665), .ZN(n12660) );
  NAND2_X1 U12535 ( .A1(n12449), .A2(n12451), .ZN(n12665) );
  NAND2_X1 U12536 ( .A1(n12666), .A2(n12667), .ZN(n12451) );
  NAND2_X1 U12537 ( .A1(b_15_), .A2(a_27_), .ZN(n12667) );
  INV_X1 U12538 ( .A(n12668), .ZN(n12666) );
  XNOR2_X1 U12539 ( .A(n12669), .B(n12670), .ZN(n12449) );
  XOR2_X1 U12540 ( .A(n12671), .B(n12672), .Z(n12669) );
  NAND2_X1 U12541 ( .A1(b_14_), .A2(a_28_), .ZN(n12671) );
  NAND2_X1 U12542 ( .A1(a_27_), .A2(n12668), .ZN(n12450) );
  NAND2_X1 U12543 ( .A1(n12673), .A2(n12674), .ZN(n12668) );
  NAND3_X1 U12544 ( .A1(a_28_), .A2(n12675), .A3(b_15_), .ZN(n12674) );
  NAND2_X1 U12545 ( .A1(n12459), .A2(n12457), .ZN(n12675) );
  OR2_X1 U12546 ( .A1(n12457), .A2(n12459), .ZN(n12673) );
  AND2_X1 U12547 ( .A1(n12676), .A2(n12677), .ZN(n12459) );
  NAND2_X1 U12548 ( .A1(n12473), .A2(n12678), .ZN(n12677) );
  OR2_X1 U12549 ( .A1(n12474), .A2(n12475), .ZN(n12678) );
  NOR2_X1 U12550 ( .A1(n8756), .A2(n7890), .ZN(n12473) );
  NAND2_X1 U12551 ( .A1(n12475), .A2(n12474), .ZN(n12676) );
  NAND2_X1 U12552 ( .A1(n12679), .A2(n12680), .ZN(n12474) );
  NAND2_X1 U12553 ( .A1(b_13_), .A2(n12681), .ZN(n12680) );
  NAND2_X1 U12554 ( .A1(n7864), .A2(n12682), .ZN(n12681) );
  NAND2_X1 U12555 ( .A1(a_31_), .A2(n8301), .ZN(n12682) );
  NAND2_X1 U12556 ( .A1(b_14_), .A2(n12683), .ZN(n12679) );
  NAND2_X1 U12557 ( .A1(n9137), .A2(n12684), .ZN(n12683) );
  NAND2_X1 U12558 ( .A1(a_30_), .A2(n8758), .ZN(n12684) );
  AND3_X1 U12559 ( .A1(b_14_), .A2(b_15_), .A3(n7818), .ZN(n12475) );
  XNOR2_X1 U12560 ( .A(n12685), .B(n12686), .ZN(n12457) );
  XOR2_X1 U12561 ( .A(n12687), .B(n12688), .Z(n12685) );
  XNOR2_X1 U12562 ( .A(n12689), .B(n12690), .ZN(n12481) );
  NAND2_X1 U12563 ( .A1(n12691), .A2(n12692), .ZN(n12689) );
  XNOR2_X1 U12564 ( .A(n12693), .B(n12694), .ZN(n12485) );
  XOR2_X1 U12565 ( .A(n12695), .B(n12696), .Z(n12693) );
  XNOR2_X1 U12566 ( .A(n12697), .B(n12698), .ZN(n12488) );
  XNOR2_X1 U12567 ( .A(n12699), .B(n12700), .ZN(n12697) );
  NOR2_X1 U12568 ( .A1(n8745), .A2(n8301), .ZN(n12700) );
  XOR2_X1 U12569 ( .A(n12701), .B(n12702), .Z(n12493) );
  XNOR2_X1 U12570 ( .A(n12703), .B(n12704), .ZN(n12702) );
  XNOR2_X1 U12571 ( .A(n12705), .B(n12706), .ZN(n12497) );
  XOR2_X1 U12572 ( .A(n12707), .B(n12708), .Z(n12706) );
  NAND2_X1 U12573 ( .A1(b_14_), .A2(a_22_), .ZN(n12708) );
  XNOR2_X1 U12574 ( .A(n12709), .B(n12710), .ZN(n12501) );
  XOR2_X1 U12575 ( .A(n12711), .B(n12712), .Z(n12709) );
  XNOR2_X1 U12576 ( .A(n12713), .B(n12714), .ZN(n12504) );
  XNOR2_X1 U12577 ( .A(n12715), .B(n12716), .ZN(n12713) );
  NOR2_X1 U12578 ( .A1(n8751), .A2(n8301), .ZN(n12716) );
  XOR2_X1 U12579 ( .A(n12717), .B(n12718), .Z(n12509) );
  XNOR2_X1 U12580 ( .A(n12719), .B(n12720), .ZN(n12718) );
  XNOR2_X1 U12581 ( .A(n12721), .B(n12722), .ZN(n12414) );
  XNOR2_X1 U12582 ( .A(n12723), .B(n12724), .ZN(n12721) );
  NOR2_X1 U12583 ( .A1(n8753), .A2(n8301), .ZN(n12724) );
  XOR2_X1 U12584 ( .A(n12725), .B(n12726), .Z(n12406) );
  XOR2_X1 U12585 ( .A(n12727), .B(n12728), .Z(n12725) );
  NOR2_X1 U12586 ( .A1(n8210), .A2(n8301), .ZN(n12728) );
  NOR2_X1 U12587 ( .A1(n8756), .A2(n8276), .ZN(n8700) );
  XOR2_X1 U12588 ( .A(n12729), .B(n12730), .Z(n12519) );
  XOR2_X1 U12589 ( .A(n12731), .B(n12732), .Z(n12729) );
  XNOR2_X1 U12590 ( .A(n12733), .B(n12734), .ZN(n12523) );
  NAND2_X1 U12591 ( .A1(n12735), .A2(n12736), .ZN(n12733) );
  XNOR2_X1 U12592 ( .A(n12737), .B(n12738), .ZN(n12528) );
  XOR2_X1 U12593 ( .A(n12739), .B(n12740), .Z(n12737) );
  XNOR2_X1 U12594 ( .A(n12741), .B(n12742), .ZN(n12531) );
  XNOR2_X1 U12595 ( .A(n12743), .B(n12744), .ZN(n12741) );
  NOR2_X1 U12596 ( .A1(n8376), .A2(n8301), .ZN(n12744) );
  XNOR2_X1 U12597 ( .A(n12745), .B(n12746), .ZN(n12535) );
  XNOR2_X1 U12598 ( .A(n12747), .B(n12748), .ZN(n12745) );
  XNOR2_X1 U12599 ( .A(n12749), .B(n12750), .ZN(n12540) );
  XOR2_X1 U12600 ( .A(n12751), .B(n12752), .Z(n12749) );
  NOR2_X1 U12601 ( .A1(n8426), .A2(n8301), .ZN(n12752) );
  XNOR2_X1 U12602 ( .A(n12753), .B(n12754), .ZN(n12543) );
  XNOR2_X1 U12603 ( .A(n12755), .B(n12756), .ZN(n12754) );
  XNOR2_X1 U12604 ( .A(n12757), .B(n12758), .ZN(n12372) );
  XOR2_X1 U12605 ( .A(n12759), .B(n12760), .Z(n12757) );
  NOR2_X1 U12606 ( .A1(n8764), .A2(n8301), .ZN(n12760) );
  XNOR2_X1 U12607 ( .A(n12761), .B(n12762), .ZN(n12363) );
  NAND2_X1 U12608 ( .A1(n12763), .A2(n12764), .ZN(n12761) );
  XOR2_X1 U12609 ( .A(n12765), .B(n12766), .Z(n12548) );
  NAND2_X1 U12610 ( .A1(n12767), .A2(n12768), .ZN(n12765) );
  XNOR2_X1 U12611 ( .A(n12769), .B(n12770), .ZN(n12551) );
  XNOR2_X1 U12612 ( .A(n12771), .B(n12772), .ZN(n12770) );
  XNOR2_X1 U12613 ( .A(n12773), .B(n12774), .ZN(n12556) );
  XNOR2_X1 U12614 ( .A(n12775), .B(n12776), .ZN(n12773) );
  XNOR2_X1 U12615 ( .A(n12777), .B(n12778), .ZN(n12560) );
  XNOR2_X1 U12616 ( .A(n12779), .B(n12780), .ZN(n12777) );
  NOR2_X1 U12617 ( .A1(n8768), .A2(n8301), .ZN(n12780) );
  XNOR2_X1 U12618 ( .A(n12781), .B(n12782), .ZN(n12564) );
  XNOR2_X1 U12619 ( .A(n12783), .B(n12784), .ZN(n12782) );
  INV_X1 U12620 ( .A(n12344), .ZN(n12346) );
  XOR2_X1 U12621 ( .A(n12785), .B(n12786), .Z(n12344) );
  XOR2_X1 U12622 ( .A(n12787), .B(n12788), .Z(n12786) );
  NAND2_X1 U12623 ( .A1(b_14_), .A2(a_0_), .ZN(n12788) );
  NAND4_X1 U12624 ( .A1(n8946), .A2(n8945), .A3(n8947), .A4(n8941), .ZN(n8894)
         );
  INV_X1 U12625 ( .A(n12789), .ZN(n8941) );
  NAND2_X1 U12626 ( .A1(n12790), .A2(n12791), .ZN(n8947) );
  NAND3_X1 U12627 ( .A1(a_0_), .A2(n12792), .A3(b_14_), .ZN(n12791) );
  OR2_X1 U12628 ( .A1(n12787), .A2(n12785), .ZN(n12792) );
  NAND2_X1 U12629 ( .A1(n12785), .A2(n12787), .ZN(n12790) );
  NAND2_X1 U12630 ( .A1(n12793), .A2(n12794), .ZN(n12787) );
  NAND2_X1 U12631 ( .A1(n12784), .A2(n12795), .ZN(n12794) );
  OR2_X1 U12632 ( .A1(n12783), .A2(n12781), .ZN(n12795) );
  NOR2_X1 U12633 ( .A1(n8301), .A2(n8617), .ZN(n12784) );
  NAND2_X1 U12634 ( .A1(n12781), .A2(n12783), .ZN(n12793) );
  NAND2_X1 U12635 ( .A1(n12796), .A2(n12797), .ZN(n12783) );
  NAND3_X1 U12636 ( .A1(a_2_), .A2(n12798), .A3(b_14_), .ZN(n12797) );
  NAND2_X1 U12637 ( .A1(n12779), .A2(n12778), .ZN(n12798) );
  OR2_X1 U12638 ( .A1(n12778), .A2(n12779), .ZN(n12796) );
  AND2_X1 U12639 ( .A1(n12799), .A2(n12800), .ZN(n12779) );
  NAND2_X1 U12640 ( .A1(n12776), .A2(n12801), .ZN(n12800) );
  NAND2_X1 U12641 ( .A1(n12775), .A2(n12774), .ZN(n12801) );
  NOR2_X1 U12642 ( .A1(n8301), .A2(n8567), .ZN(n12776) );
  OR2_X1 U12643 ( .A1(n12774), .A2(n12775), .ZN(n12799) );
  AND2_X1 U12644 ( .A1(n12802), .A2(n12803), .ZN(n12775) );
  NAND2_X1 U12645 ( .A1(n12772), .A2(n12804), .ZN(n12803) );
  OR2_X1 U12646 ( .A1(n12771), .A2(n12769), .ZN(n12804) );
  NOR2_X1 U12647 ( .A1(n8301), .A2(n8766), .ZN(n12772) );
  NAND2_X1 U12648 ( .A1(n12769), .A2(n12771), .ZN(n12802) );
  NAND2_X1 U12649 ( .A1(n12767), .A2(n12805), .ZN(n12771) );
  NAND2_X1 U12650 ( .A1(n12766), .A2(n12768), .ZN(n12805) );
  NAND2_X1 U12651 ( .A1(n12806), .A2(n12807), .ZN(n12768) );
  NAND2_X1 U12652 ( .A1(b_14_), .A2(a_5_), .ZN(n12807) );
  INV_X1 U12653 ( .A(n12808), .ZN(n12806) );
  XNOR2_X1 U12654 ( .A(n12809), .B(n12810), .ZN(n12766) );
  XOR2_X1 U12655 ( .A(n12811), .B(n12812), .Z(n12810) );
  NAND2_X1 U12656 ( .A1(b_13_), .A2(a_6_), .ZN(n12812) );
  NAND2_X1 U12657 ( .A1(a_5_), .A2(n12808), .ZN(n12767) );
  NAND2_X1 U12658 ( .A1(n12763), .A2(n12813), .ZN(n12808) );
  NAND2_X1 U12659 ( .A1(n12762), .A2(n12764), .ZN(n12813) );
  NAND2_X1 U12660 ( .A1(n12814), .A2(n12815), .ZN(n12764) );
  NAND2_X1 U12661 ( .A1(b_14_), .A2(a_6_), .ZN(n12815) );
  INV_X1 U12662 ( .A(n12816), .ZN(n12814) );
  XNOR2_X1 U12663 ( .A(n12817), .B(n12818), .ZN(n12762) );
  XOR2_X1 U12664 ( .A(n12819), .B(n12820), .Z(n12818) );
  NAND2_X1 U12665 ( .A1(b_13_), .A2(a_7_), .ZN(n12820) );
  NAND2_X1 U12666 ( .A1(a_6_), .A2(n12816), .ZN(n12763) );
  NAND2_X1 U12667 ( .A1(n12821), .A2(n12822), .ZN(n12816) );
  NAND3_X1 U12668 ( .A1(a_7_), .A2(n12823), .A3(b_14_), .ZN(n12822) );
  OR2_X1 U12669 ( .A1(n12759), .A2(n12758), .ZN(n12823) );
  NAND2_X1 U12670 ( .A1(n12758), .A2(n12759), .ZN(n12821) );
  NAND2_X1 U12671 ( .A1(n12824), .A2(n12825), .ZN(n12759) );
  NAND2_X1 U12672 ( .A1(n12756), .A2(n12826), .ZN(n12825) );
  OR2_X1 U12673 ( .A1(n12755), .A2(n12753), .ZN(n12826) );
  NOR2_X1 U12674 ( .A1(n8301), .A2(n8763), .ZN(n12756) );
  NAND2_X1 U12675 ( .A1(n12753), .A2(n12755), .ZN(n12824) );
  NAND2_X1 U12676 ( .A1(n12827), .A2(n12828), .ZN(n12755) );
  NAND3_X1 U12677 ( .A1(a_9_), .A2(n12829), .A3(b_14_), .ZN(n12828) );
  OR2_X1 U12678 ( .A1(n12751), .A2(n12750), .ZN(n12829) );
  NAND2_X1 U12679 ( .A1(n12750), .A2(n12751), .ZN(n12827) );
  NAND2_X1 U12680 ( .A1(n12830), .A2(n12831), .ZN(n12751) );
  NAND2_X1 U12681 ( .A1(n12748), .A2(n12832), .ZN(n12831) );
  NAND2_X1 U12682 ( .A1(n12747), .A2(n12746), .ZN(n12832) );
  NOR2_X1 U12683 ( .A1(n8301), .A2(n8761), .ZN(n12748) );
  OR2_X1 U12684 ( .A1(n12746), .A2(n12747), .ZN(n12830) );
  AND2_X1 U12685 ( .A1(n12833), .A2(n12834), .ZN(n12747) );
  NAND3_X1 U12686 ( .A1(a_11_), .A2(n12835), .A3(b_14_), .ZN(n12834) );
  NAND2_X1 U12687 ( .A1(n12743), .A2(n12742), .ZN(n12835) );
  OR2_X1 U12688 ( .A1(n12742), .A2(n12743), .ZN(n12833) );
  AND2_X1 U12689 ( .A1(n12836), .A2(n12837), .ZN(n12743) );
  NAND2_X1 U12690 ( .A1(n12740), .A2(n12838), .ZN(n12837) );
  OR2_X1 U12691 ( .A1(n12739), .A2(n12738), .ZN(n12838) );
  NOR2_X1 U12692 ( .A1(n8301), .A2(n8759), .ZN(n12740) );
  NAND2_X1 U12693 ( .A1(n12738), .A2(n12739), .ZN(n12836) );
  NAND2_X1 U12694 ( .A1(n12735), .A2(n12839), .ZN(n12739) );
  NAND2_X1 U12695 ( .A1(n12734), .A2(n12736), .ZN(n12839) );
  NAND2_X1 U12696 ( .A1(n12840), .A2(n12841), .ZN(n12736) );
  NAND2_X1 U12697 ( .A1(b_14_), .A2(a_13_), .ZN(n12841) );
  INV_X1 U12698 ( .A(n12842), .ZN(n12840) );
  XOR2_X1 U12699 ( .A(n12843), .B(n12844), .Z(n12734) );
  XOR2_X1 U12700 ( .A(n12845), .B(n12846), .Z(n12843) );
  NOR2_X1 U12701 ( .A1(n8757), .A2(n8758), .ZN(n12846) );
  NAND2_X1 U12702 ( .A1(a_13_), .A2(n12842), .ZN(n12735) );
  NAND2_X1 U12703 ( .A1(n12847), .A2(n12848), .ZN(n12842) );
  NAND2_X1 U12704 ( .A1(n12730), .A2(n12849), .ZN(n12848) );
  OR2_X1 U12705 ( .A1(n12731), .A2(n12732), .ZN(n12849) );
  XNOR2_X1 U12706 ( .A(n12850), .B(n12851), .ZN(n12730) );
  XOR2_X1 U12707 ( .A(n12852), .B(n12853), .Z(n12851) );
  NAND2_X1 U12708 ( .A1(b_13_), .A2(a_15_), .ZN(n12853) );
  NAND2_X1 U12709 ( .A1(n12732), .A2(n12731), .ZN(n12847) );
  NAND2_X1 U12710 ( .A1(n12854), .A2(n12855), .ZN(n12731) );
  NAND2_X1 U12711 ( .A1(n12619), .A2(n12856), .ZN(n12855) );
  OR2_X1 U12712 ( .A1(n12618), .A2(n12617), .ZN(n12856) );
  NOR2_X1 U12713 ( .A1(n8301), .A2(n8276), .ZN(n12619) );
  NAND2_X1 U12714 ( .A1(n12617), .A2(n12618), .ZN(n12854) );
  NAND2_X1 U12715 ( .A1(n12857), .A2(n12858), .ZN(n12618) );
  NAND2_X1 U12716 ( .A1(n12626), .A2(n12859), .ZN(n12858) );
  OR2_X1 U12717 ( .A1(n12625), .A2(n12623), .ZN(n12859) );
  NOR2_X1 U12718 ( .A1(n8301), .A2(n8755), .ZN(n12626) );
  NAND2_X1 U12719 ( .A1(n12623), .A2(n12625), .ZN(n12857) );
  NAND2_X1 U12720 ( .A1(n12860), .A2(n12861), .ZN(n12625) );
  NAND3_X1 U12721 ( .A1(a_17_), .A2(n12862), .A3(b_14_), .ZN(n12861) );
  OR2_X1 U12722 ( .A1(n12727), .A2(n12726), .ZN(n12862) );
  NAND2_X1 U12723 ( .A1(n12726), .A2(n12727), .ZN(n12860) );
  NAND2_X1 U12724 ( .A1(n12863), .A2(n12864), .ZN(n12727) );
  NAND3_X1 U12725 ( .A1(a_18_), .A2(n12865), .A3(b_14_), .ZN(n12864) );
  NAND2_X1 U12726 ( .A1(n12723), .A2(n12722), .ZN(n12865) );
  OR2_X1 U12727 ( .A1(n12722), .A2(n12723), .ZN(n12863) );
  AND2_X1 U12728 ( .A1(n12866), .A2(n12867), .ZN(n12723) );
  NAND2_X1 U12729 ( .A1(n12720), .A2(n12868), .ZN(n12867) );
  OR2_X1 U12730 ( .A1(n12719), .A2(n12717), .ZN(n12868) );
  NOR2_X1 U12731 ( .A1(n8301), .A2(n8170), .ZN(n12720) );
  NAND2_X1 U12732 ( .A1(n12717), .A2(n12719), .ZN(n12866) );
  NAND2_X1 U12733 ( .A1(n12869), .A2(n12870), .ZN(n12719) );
  NAND3_X1 U12734 ( .A1(a_20_), .A2(n12871), .A3(b_14_), .ZN(n12870) );
  NAND2_X1 U12735 ( .A1(n12715), .A2(n12714), .ZN(n12871) );
  OR2_X1 U12736 ( .A1(n12714), .A2(n12715), .ZN(n12869) );
  AND2_X1 U12737 ( .A1(n12872), .A2(n12873), .ZN(n12715) );
  NAND2_X1 U12738 ( .A1(n12712), .A2(n12874), .ZN(n12873) );
  OR2_X1 U12739 ( .A1(n12711), .A2(n12710), .ZN(n12874) );
  NOR2_X1 U12740 ( .A1(n8301), .A2(n8750), .ZN(n12712) );
  NAND2_X1 U12741 ( .A1(n12710), .A2(n12711), .ZN(n12872) );
  NAND2_X1 U12742 ( .A1(n12875), .A2(n12876), .ZN(n12711) );
  NAND3_X1 U12743 ( .A1(a_22_), .A2(n12877), .A3(b_14_), .ZN(n12876) );
  OR2_X1 U12744 ( .A1(n12707), .A2(n12705), .ZN(n12877) );
  NAND2_X1 U12745 ( .A1(n12705), .A2(n12707), .ZN(n12875) );
  NAND2_X1 U12746 ( .A1(n12878), .A2(n12879), .ZN(n12707) );
  NAND2_X1 U12747 ( .A1(n12704), .A2(n12880), .ZN(n12879) );
  OR2_X1 U12748 ( .A1(n12703), .A2(n12701), .ZN(n12880) );
  NOR2_X1 U12749 ( .A1(n8301), .A2(n8747), .ZN(n12704) );
  NAND2_X1 U12750 ( .A1(n12701), .A2(n12703), .ZN(n12878) );
  NAND2_X1 U12751 ( .A1(n12881), .A2(n12882), .ZN(n12703) );
  NAND3_X1 U12752 ( .A1(a_24_), .A2(n12883), .A3(b_14_), .ZN(n12882) );
  NAND2_X1 U12753 ( .A1(n12699), .A2(n12698), .ZN(n12883) );
  OR2_X1 U12754 ( .A1(n12698), .A2(n12699), .ZN(n12881) );
  AND2_X1 U12755 ( .A1(n12884), .A2(n12885), .ZN(n12699) );
  NAND2_X1 U12756 ( .A1(n12696), .A2(n12886), .ZN(n12885) );
  OR2_X1 U12757 ( .A1(n12695), .A2(n12694), .ZN(n12886) );
  NOR2_X1 U12758 ( .A1(n8301), .A2(n8744), .ZN(n12696) );
  NAND2_X1 U12759 ( .A1(n12694), .A2(n12695), .ZN(n12884) );
  NAND2_X1 U12760 ( .A1(n12691), .A2(n12887), .ZN(n12695) );
  NAND2_X1 U12761 ( .A1(n12690), .A2(n12692), .ZN(n12887) );
  NAND2_X1 U12762 ( .A1(n12888), .A2(n12889), .ZN(n12692) );
  NAND2_X1 U12763 ( .A1(b_14_), .A2(a_26_), .ZN(n12889) );
  INV_X1 U12764 ( .A(n12890), .ZN(n12888) );
  XNOR2_X1 U12765 ( .A(n12891), .B(n12892), .ZN(n12690) );
  NAND2_X1 U12766 ( .A1(n12893), .A2(n12894), .ZN(n12891) );
  NAND2_X1 U12767 ( .A1(a_26_), .A2(n12890), .ZN(n12691) );
  NAND2_X1 U12768 ( .A1(n12663), .A2(n12895), .ZN(n12890) );
  NAND2_X1 U12769 ( .A1(n12662), .A2(n12664), .ZN(n12895) );
  NAND2_X1 U12770 ( .A1(n12896), .A2(n12897), .ZN(n12664) );
  NAND2_X1 U12771 ( .A1(b_14_), .A2(a_27_), .ZN(n12897) );
  INV_X1 U12772 ( .A(n12898), .ZN(n12896) );
  XNOR2_X1 U12773 ( .A(n12899), .B(n12900), .ZN(n12662) );
  XOR2_X1 U12774 ( .A(n12901), .B(n12902), .Z(n12899) );
  NAND2_X1 U12775 ( .A1(b_13_), .A2(a_28_), .ZN(n12901) );
  NAND2_X1 U12776 ( .A1(a_27_), .A2(n12898), .ZN(n12663) );
  NAND2_X1 U12777 ( .A1(n12903), .A2(n12904), .ZN(n12898) );
  NAND3_X1 U12778 ( .A1(a_28_), .A2(n12905), .A3(b_14_), .ZN(n12904) );
  NAND2_X1 U12779 ( .A1(n12672), .A2(n12670), .ZN(n12905) );
  OR2_X1 U12780 ( .A1(n12670), .A2(n12672), .ZN(n12903) );
  AND2_X1 U12781 ( .A1(n12906), .A2(n12907), .ZN(n12672) );
  NAND2_X1 U12782 ( .A1(n12686), .A2(n12908), .ZN(n12907) );
  OR2_X1 U12783 ( .A1(n12687), .A2(n12688), .ZN(n12908) );
  NOR2_X1 U12784 ( .A1(n8301), .A2(n7890), .ZN(n12686) );
  NAND2_X1 U12785 ( .A1(n12688), .A2(n12687), .ZN(n12906) );
  NAND2_X1 U12786 ( .A1(n12909), .A2(n12910), .ZN(n12687) );
  NAND2_X1 U12787 ( .A1(b_12_), .A2(n12911), .ZN(n12910) );
  NAND2_X1 U12788 ( .A1(n7864), .A2(n12912), .ZN(n12911) );
  NAND2_X1 U12789 ( .A1(a_31_), .A2(n8758), .ZN(n12912) );
  NAND2_X1 U12790 ( .A1(b_13_), .A2(n12913), .ZN(n12909) );
  NAND2_X1 U12791 ( .A1(n9137), .A2(n12914), .ZN(n12913) );
  NAND2_X1 U12792 ( .A1(a_30_), .A2(n8351), .ZN(n12914) );
  AND3_X1 U12793 ( .A1(b_13_), .A2(b_14_), .A3(n7818), .ZN(n12688) );
  XNOR2_X1 U12794 ( .A(n12915), .B(n12916), .ZN(n12670) );
  XOR2_X1 U12795 ( .A(n12917), .B(n12918), .Z(n12915) );
  XNOR2_X1 U12796 ( .A(n12919), .B(n12920), .ZN(n12694) );
  NAND2_X1 U12797 ( .A1(n12921), .A2(n12922), .ZN(n12919) );
  XNOR2_X1 U12798 ( .A(n12923), .B(n12924), .ZN(n12698) );
  XOR2_X1 U12799 ( .A(n12925), .B(n12926), .Z(n12923) );
  XNOR2_X1 U12800 ( .A(n12927), .B(n12928), .ZN(n12701) );
  XNOR2_X1 U12801 ( .A(n12929), .B(n12930), .ZN(n12927) );
  NOR2_X1 U12802 ( .A1(n8745), .A2(n8758), .ZN(n12930) );
  XNOR2_X1 U12803 ( .A(n12931), .B(n12932), .ZN(n12705) );
  XNOR2_X1 U12804 ( .A(n12933), .B(n12934), .ZN(n12932) );
  XNOR2_X1 U12805 ( .A(n12935), .B(n12936), .ZN(n12710) );
  XOR2_X1 U12806 ( .A(n12937), .B(n12938), .Z(n12936) );
  NAND2_X1 U12807 ( .A1(b_13_), .A2(a_22_), .ZN(n12938) );
  XNOR2_X1 U12808 ( .A(n12939), .B(n12940), .ZN(n12714) );
  XOR2_X1 U12809 ( .A(n12941), .B(n12942), .Z(n12939) );
  XNOR2_X1 U12810 ( .A(n12943), .B(n12944), .ZN(n12717) );
  XNOR2_X1 U12811 ( .A(n12945), .B(n12946), .ZN(n12943) );
  NOR2_X1 U12812 ( .A1(n8751), .A2(n8758), .ZN(n12946) );
  XOR2_X1 U12813 ( .A(n12947), .B(n12948), .Z(n12722) );
  XNOR2_X1 U12814 ( .A(n12949), .B(n12950), .ZN(n12948) );
  XNOR2_X1 U12815 ( .A(n12951), .B(n12952), .ZN(n12726) );
  XNOR2_X1 U12816 ( .A(n12953), .B(n12954), .ZN(n12951) );
  XNOR2_X1 U12817 ( .A(n12955), .B(n12956), .ZN(n12623) );
  XOR2_X1 U12818 ( .A(n12957), .B(n12958), .Z(n12955) );
  NAND2_X1 U12819 ( .A1(b_13_), .A2(a_17_), .ZN(n12957) );
  XNOR2_X1 U12820 ( .A(n12959), .B(n12960), .ZN(n12617) );
  XNOR2_X1 U12821 ( .A(n12961), .B(n12962), .ZN(n12959) );
  NOR2_X1 U12822 ( .A1(n8755), .A2(n8758), .ZN(n12962) );
  INV_X1 U12823 ( .A(n8697), .ZN(n12732) );
  NAND2_X1 U12824 ( .A1(b_14_), .A2(a_14_), .ZN(n8697) );
  XOR2_X1 U12825 ( .A(n12963), .B(n12964), .Z(n12738) );
  XOR2_X1 U12826 ( .A(n12965), .B(n12966), .Z(n12963) );
  XNOR2_X1 U12827 ( .A(n12967), .B(n12968), .ZN(n12742) );
  XNOR2_X1 U12828 ( .A(n12969), .B(n12970), .ZN(n12967) );
  NAND2_X1 U12829 ( .A1(b_13_), .A2(a_12_), .ZN(n12969) );
  XOR2_X1 U12830 ( .A(n12971), .B(n12972), .Z(n12746) );
  XOR2_X1 U12831 ( .A(n12973), .B(n12974), .Z(n12972) );
  NAND2_X1 U12832 ( .A1(b_13_), .A2(a_11_), .ZN(n12974) );
  XNOR2_X1 U12833 ( .A(n12975), .B(n12976), .ZN(n12750) );
  XNOR2_X1 U12834 ( .A(n12977), .B(n12978), .ZN(n12975) );
  NOR2_X1 U12835 ( .A1(n8761), .A2(n8758), .ZN(n12978) );
  XNOR2_X1 U12836 ( .A(n12979), .B(n12980), .ZN(n12753) );
  XOR2_X1 U12837 ( .A(n12981), .B(n12982), .Z(n12980) );
  NAND2_X1 U12838 ( .A1(b_13_), .A2(a_9_), .ZN(n12982) );
  XNOR2_X1 U12839 ( .A(n12983), .B(n12984), .ZN(n12758) );
  XNOR2_X1 U12840 ( .A(n12985), .B(n12986), .ZN(n12983) );
  NOR2_X1 U12841 ( .A1(n8763), .A2(n8758), .ZN(n12986) );
  XNOR2_X1 U12842 ( .A(n12987), .B(n12988), .ZN(n12769) );
  XNOR2_X1 U12843 ( .A(n12989), .B(n12990), .ZN(n12987) );
  NOR2_X1 U12844 ( .A1(n8517), .A2(n8758), .ZN(n12990) );
  XOR2_X1 U12845 ( .A(n12991), .B(n12992), .Z(n12774) );
  XOR2_X1 U12846 ( .A(n12993), .B(n12994), .Z(n12992) );
  NAND2_X1 U12847 ( .A1(b_13_), .A2(a_4_), .ZN(n12994) );
  XOR2_X1 U12848 ( .A(n12995), .B(n12996), .Z(n12778) );
  XOR2_X1 U12849 ( .A(n12997), .B(n12998), .Z(n12996) );
  NAND2_X1 U12850 ( .A1(b_13_), .A2(a_3_), .ZN(n12998) );
  XOR2_X1 U12851 ( .A(n12999), .B(n13000), .Z(n12781) );
  XOR2_X1 U12852 ( .A(n13001), .B(n13002), .Z(n12999) );
  NOR2_X1 U12853 ( .A1(n8768), .A2(n8758), .ZN(n13002) );
  XNOR2_X1 U12854 ( .A(n13003), .B(n13004), .ZN(n12785) );
  XOR2_X1 U12855 ( .A(n13005), .B(n13006), .Z(n13004) );
  NAND2_X1 U12856 ( .A1(b_13_), .A2(a_1_), .ZN(n13006) );
  NAND2_X1 U12857 ( .A1(n13007), .A2(n13008), .ZN(n8945) );
  XNOR2_X1 U12858 ( .A(n13009), .B(n13010), .ZN(n8946) );
  XNOR2_X1 U12859 ( .A(n13011), .B(n13012), .ZN(n13010) );
  NAND2_X1 U12860 ( .A1(n12789), .A2(n13013), .ZN(n8900) );
  XOR2_X1 U12861 ( .A(n8938), .B(n8937), .Z(n13013) );
  NOR2_X1 U12862 ( .A1(n13008), .A2(n13007), .ZN(n12789) );
  AND2_X1 U12863 ( .A1(n13014), .A2(n13015), .ZN(n13007) );
  NAND2_X1 U12864 ( .A1(n13012), .A2(n13016), .ZN(n13015) );
  OR2_X1 U12865 ( .A1(n13011), .A2(n13009), .ZN(n13016) );
  NOR2_X1 U12866 ( .A1(n8758), .A2(n9674), .ZN(n13012) );
  NAND2_X1 U12867 ( .A1(n13009), .A2(n13011), .ZN(n13014) );
  NAND2_X1 U12868 ( .A1(n13017), .A2(n13018), .ZN(n13011) );
  NAND3_X1 U12869 ( .A1(a_1_), .A2(n13019), .A3(b_13_), .ZN(n13018) );
  OR2_X1 U12870 ( .A1(n13005), .A2(n13003), .ZN(n13019) );
  NAND2_X1 U12871 ( .A1(n13003), .A2(n13005), .ZN(n13017) );
  NAND2_X1 U12872 ( .A1(n13020), .A2(n13021), .ZN(n13005) );
  NAND3_X1 U12873 ( .A1(a_2_), .A2(n13022), .A3(b_13_), .ZN(n13021) );
  OR2_X1 U12874 ( .A1(n13001), .A2(n13000), .ZN(n13022) );
  NAND2_X1 U12875 ( .A1(n13000), .A2(n13001), .ZN(n13020) );
  NAND2_X1 U12876 ( .A1(n13023), .A2(n13024), .ZN(n13001) );
  NAND3_X1 U12877 ( .A1(a_3_), .A2(n13025), .A3(b_13_), .ZN(n13024) );
  OR2_X1 U12878 ( .A1(n12997), .A2(n12995), .ZN(n13025) );
  NAND2_X1 U12879 ( .A1(n12995), .A2(n12997), .ZN(n13023) );
  NAND2_X1 U12880 ( .A1(n13026), .A2(n13027), .ZN(n12997) );
  NAND3_X1 U12881 ( .A1(a_4_), .A2(n13028), .A3(b_13_), .ZN(n13027) );
  OR2_X1 U12882 ( .A1(n12993), .A2(n12991), .ZN(n13028) );
  NAND2_X1 U12883 ( .A1(n12991), .A2(n12993), .ZN(n13026) );
  NAND2_X1 U12884 ( .A1(n13029), .A2(n13030), .ZN(n12993) );
  NAND3_X1 U12885 ( .A1(a_5_), .A2(n13031), .A3(b_13_), .ZN(n13030) );
  NAND2_X1 U12886 ( .A1(n12989), .A2(n12988), .ZN(n13031) );
  OR2_X1 U12887 ( .A1(n12988), .A2(n12989), .ZN(n13029) );
  AND2_X1 U12888 ( .A1(n13032), .A2(n13033), .ZN(n12989) );
  NAND3_X1 U12889 ( .A1(a_6_), .A2(n13034), .A3(b_13_), .ZN(n13033) );
  OR2_X1 U12890 ( .A1(n12811), .A2(n12809), .ZN(n13034) );
  NAND2_X1 U12891 ( .A1(n12809), .A2(n12811), .ZN(n13032) );
  NAND2_X1 U12892 ( .A1(n13035), .A2(n13036), .ZN(n12811) );
  NAND3_X1 U12893 ( .A1(a_7_), .A2(n13037), .A3(b_13_), .ZN(n13036) );
  OR2_X1 U12894 ( .A1(n12819), .A2(n12817), .ZN(n13037) );
  NAND2_X1 U12895 ( .A1(n12817), .A2(n12819), .ZN(n13035) );
  NAND2_X1 U12896 ( .A1(n13038), .A2(n13039), .ZN(n12819) );
  NAND3_X1 U12897 ( .A1(a_8_), .A2(n13040), .A3(b_13_), .ZN(n13039) );
  NAND2_X1 U12898 ( .A1(n12985), .A2(n12984), .ZN(n13040) );
  OR2_X1 U12899 ( .A1(n12984), .A2(n12985), .ZN(n13038) );
  AND2_X1 U12900 ( .A1(n13041), .A2(n13042), .ZN(n12985) );
  NAND3_X1 U12901 ( .A1(a_9_), .A2(n13043), .A3(b_13_), .ZN(n13042) );
  OR2_X1 U12902 ( .A1(n12981), .A2(n12979), .ZN(n13043) );
  NAND2_X1 U12903 ( .A1(n12979), .A2(n12981), .ZN(n13041) );
  NAND2_X1 U12904 ( .A1(n13044), .A2(n13045), .ZN(n12981) );
  NAND3_X1 U12905 ( .A1(a_10_), .A2(n13046), .A3(b_13_), .ZN(n13045) );
  NAND2_X1 U12906 ( .A1(n12977), .A2(n12976), .ZN(n13046) );
  OR2_X1 U12907 ( .A1(n12976), .A2(n12977), .ZN(n13044) );
  AND2_X1 U12908 ( .A1(n13047), .A2(n13048), .ZN(n12977) );
  NAND3_X1 U12909 ( .A1(a_11_), .A2(n13049), .A3(b_13_), .ZN(n13048) );
  OR2_X1 U12910 ( .A1(n12973), .A2(n12971), .ZN(n13049) );
  NAND2_X1 U12911 ( .A1(n12971), .A2(n12973), .ZN(n13047) );
  NAND2_X1 U12912 ( .A1(n13050), .A2(n13051), .ZN(n12973) );
  NAND3_X1 U12913 ( .A1(a_12_), .A2(n13052), .A3(b_13_), .ZN(n13051) );
  OR2_X1 U12914 ( .A1(n12970), .A2(n12968), .ZN(n13052) );
  NAND2_X1 U12915 ( .A1(n12968), .A2(n12970), .ZN(n13050) );
  NAND2_X1 U12916 ( .A1(n13053), .A2(n13054), .ZN(n12970) );
  NAND2_X1 U12917 ( .A1(n12964), .A2(n13055), .ZN(n13054) );
  OR2_X1 U12918 ( .A1(n12965), .A2(n12966), .ZN(n13055) );
  XNOR2_X1 U12919 ( .A(n13056), .B(n13057), .ZN(n12964) );
  NAND2_X1 U12920 ( .A1(n13058), .A2(n13059), .ZN(n13056) );
  NAND2_X1 U12921 ( .A1(n12966), .A2(n12965), .ZN(n13053) );
  NAND2_X1 U12922 ( .A1(n13060), .A2(n13061), .ZN(n12965) );
  NAND3_X1 U12923 ( .A1(a_14_), .A2(n13062), .A3(b_13_), .ZN(n13061) );
  OR2_X1 U12924 ( .A1(n12845), .A2(n12844), .ZN(n13062) );
  NAND2_X1 U12925 ( .A1(n12844), .A2(n12845), .ZN(n13060) );
  NAND2_X1 U12926 ( .A1(n13063), .A2(n13064), .ZN(n12845) );
  NAND3_X1 U12927 ( .A1(a_15_), .A2(n13065), .A3(b_13_), .ZN(n13064) );
  OR2_X1 U12928 ( .A1(n12852), .A2(n12850), .ZN(n13065) );
  NAND2_X1 U12929 ( .A1(n12850), .A2(n12852), .ZN(n13063) );
  NAND2_X1 U12930 ( .A1(n13066), .A2(n13067), .ZN(n12852) );
  NAND3_X1 U12931 ( .A1(a_16_), .A2(n13068), .A3(b_13_), .ZN(n13067) );
  NAND2_X1 U12932 ( .A1(n12961), .A2(n12960), .ZN(n13068) );
  OR2_X1 U12933 ( .A1(n12960), .A2(n12961), .ZN(n13066) );
  AND2_X1 U12934 ( .A1(n13069), .A2(n13070), .ZN(n12961) );
  NAND3_X1 U12935 ( .A1(a_17_), .A2(n13071), .A3(b_13_), .ZN(n13070) );
  NAND2_X1 U12936 ( .A1(n12958), .A2(n12956), .ZN(n13071) );
  OR2_X1 U12937 ( .A1(n12956), .A2(n12958), .ZN(n13069) );
  AND2_X1 U12938 ( .A1(n13072), .A2(n13073), .ZN(n12958) );
  NAND2_X1 U12939 ( .A1(n12954), .A2(n13074), .ZN(n13073) );
  NAND2_X1 U12940 ( .A1(n12953), .A2(n12952), .ZN(n13074) );
  NOR2_X1 U12941 ( .A1(n8758), .A2(n8753), .ZN(n12954) );
  OR2_X1 U12942 ( .A1(n12952), .A2(n12953), .ZN(n13072) );
  AND2_X1 U12943 ( .A1(n13075), .A2(n13076), .ZN(n12953) );
  NAND2_X1 U12944 ( .A1(n12950), .A2(n13077), .ZN(n13076) );
  OR2_X1 U12945 ( .A1(n12949), .A2(n12947), .ZN(n13077) );
  NOR2_X1 U12946 ( .A1(n8758), .A2(n8170), .ZN(n12950) );
  NAND2_X1 U12947 ( .A1(n12947), .A2(n12949), .ZN(n13075) );
  NAND2_X1 U12948 ( .A1(n13078), .A2(n13079), .ZN(n12949) );
  NAND3_X1 U12949 ( .A1(a_20_), .A2(n13080), .A3(b_13_), .ZN(n13079) );
  NAND2_X1 U12950 ( .A1(n12945), .A2(n12944), .ZN(n13080) );
  OR2_X1 U12951 ( .A1(n12944), .A2(n12945), .ZN(n13078) );
  AND2_X1 U12952 ( .A1(n13081), .A2(n13082), .ZN(n12945) );
  NAND2_X1 U12953 ( .A1(n12942), .A2(n13083), .ZN(n13082) );
  OR2_X1 U12954 ( .A1(n12941), .A2(n12940), .ZN(n13083) );
  NOR2_X1 U12955 ( .A1(n8758), .A2(n8750), .ZN(n12942) );
  NAND2_X1 U12956 ( .A1(n12940), .A2(n12941), .ZN(n13081) );
  NAND2_X1 U12957 ( .A1(n13084), .A2(n13085), .ZN(n12941) );
  NAND3_X1 U12958 ( .A1(a_22_), .A2(n13086), .A3(b_13_), .ZN(n13085) );
  OR2_X1 U12959 ( .A1(n12937), .A2(n12935), .ZN(n13086) );
  NAND2_X1 U12960 ( .A1(n12935), .A2(n12937), .ZN(n13084) );
  NAND2_X1 U12961 ( .A1(n13087), .A2(n13088), .ZN(n12937) );
  NAND2_X1 U12962 ( .A1(n12934), .A2(n13089), .ZN(n13088) );
  OR2_X1 U12963 ( .A1(n12933), .A2(n12931), .ZN(n13089) );
  NOR2_X1 U12964 ( .A1(n8758), .A2(n8747), .ZN(n12934) );
  NAND2_X1 U12965 ( .A1(n12931), .A2(n12933), .ZN(n13087) );
  NAND2_X1 U12966 ( .A1(n13090), .A2(n13091), .ZN(n12933) );
  NAND3_X1 U12967 ( .A1(a_24_), .A2(n13092), .A3(b_13_), .ZN(n13091) );
  NAND2_X1 U12968 ( .A1(n12929), .A2(n12928), .ZN(n13092) );
  OR2_X1 U12969 ( .A1(n12928), .A2(n12929), .ZN(n13090) );
  AND2_X1 U12970 ( .A1(n13093), .A2(n13094), .ZN(n12929) );
  NAND2_X1 U12971 ( .A1(n12926), .A2(n13095), .ZN(n13094) );
  OR2_X1 U12972 ( .A1(n12925), .A2(n12924), .ZN(n13095) );
  NOR2_X1 U12973 ( .A1(n8758), .A2(n8744), .ZN(n12926) );
  NAND2_X1 U12974 ( .A1(n12924), .A2(n12925), .ZN(n13093) );
  NAND2_X1 U12975 ( .A1(n12921), .A2(n13096), .ZN(n12925) );
  NAND2_X1 U12976 ( .A1(n12920), .A2(n12922), .ZN(n13096) );
  NAND2_X1 U12977 ( .A1(n13097), .A2(n13098), .ZN(n12922) );
  NAND2_X1 U12978 ( .A1(b_13_), .A2(a_26_), .ZN(n13098) );
  INV_X1 U12979 ( .A(n13099), .ZN(n13097) );
  XNOR2_X1 U12980 ( .A(n13100), .B(n13101), .ZN(n12920) );
  NAND2_X1 U12981 ( .A1(n13102), .A2(n13103), .ZN(n13100) );
  NAND2_X1 U12982 ( .A1(a_26_), .A2(n13099), .ZN(n12921) );
  NAND2_X1 U12983 ( .A1(n12893), .A2(n13104), .ZN(n13099) );
  NAND2_X1 U12984 ( .A1(n12892), .A2(n12894), .ZN(n13104) );
  NAND2_X1 U12985 ( .A1(n13105), .A2(n13106), .ZN(n12894) );
  NAND2_X1 U12986 ( .A1(b_13_), .A2(a_27_), .ZN(n13106) );
  INV_X1 U12987 ( .A(n13107), .ZN(n13105) );
  XNOR2_X1 U12988 ( .A(n13108), .B(n13109), .ZN(n12892) );
  XOR2_X1 U12989 ( .A(n13110), .B(n13111), .Z(n13108) );
  NAND2_X1 U12990 ( .A1(b_12_), .A2(a_28_), .ZN(n13110) );
  NAND2_X1 U12991 ( .A1(a_27_), .A2(n13107), .ZN(n12893) );
  NAND2_X1 U12992 ( .A1(n13112), .A2(n13113), .ZN(n13107) );
  NAND3_X1 U12993 ( .A1(a_28_), .A2(n13114), .A3(b_13_), .ZN(n13113) );
  NAND2_X1 U12994 ( .A1(n12902), .A2(n12900), .ZN(n13114) );
  OR2_X1 U12995 ( .A1(n12900), .A2(n12902), .ZN(n13112) );
  AND2_X1 U12996 ( .A1(n13115), .A2(n13116), .ZN(n12902) );
  NAND2_X1 U12997 ( .A1(n12916), .A2(n13117), .ZN(n13116) );
  OR2_X1 U12998 ( .A1(n12917), .A2(n12918), .ZN(n13117) );
  NOR2_X1 U12999 ( .A1(n8758), .A2(n7890), .ZN(n12916) );
  NAND2_X1 U13000 ( .A1(n12918), .A2(n12917), .ZN(n13115) );
  NAND2_X1 U13001 ( .A1(n13118), .A2(n13119), .ZN(n12917) );
  NAND2_X1 U13002 ( .A1(b_11_), .A2(n13120), .ZN(n13119) );
  NAND2_X1 U13003 ( .A1(n7864), .A2(n13121), .ZN(n13120) );
  NAND2_X1 U13004 ( .A1(a_31_), .A2(n8351), .ZN(n13121) );
  NAND2_X1 U13005 ( .A1(b_12_), .A2(n13122), .ZN(n13118) );
  NAND2_X1 U13006 ( .A1(n9137), .A2(n13123), .ZN(n13122) );
  NAND2_X1 U13007 ( .A1(a_30_), .A2(n8760), .ZN(n13123) );
  AND3_X1 U13008 ( .A1(b_12_), .A2(b_13_), .A3(n7818), .ZN(n12918) );
  XNOR2_X1 U13009 ( .A(n13124), .B(n13125), .ZN(n12900) );
  XOR2_X1 U13010 ( .A(n13126), .B(n13127), .Z(n13124) );
  XNOR2_X1 U13011 ( .A(n13128), .B(n13129), .ZN(n12924) );
  NAND2_X1 U13012 ( .A1(n13130), .A2(n13131), .ZN(n13128) );
  XNOR2_X1 U13013 ( .A(n13132), .B(n13133), .ZN(n12928) );
  XOR2_X1 U13014 ( .A(n13134), .B(n13135), .Z(n13132) );
  XNOR2_X1 U13015 ( .A(n13136), .B(n13137), .ZN(n12931) );
  XNOR2_X1 U13016 ( .A(n13138), .B(n13139), .ZN(n13136) );
  NOR2_X1 U13017 ( .A1(n8745), .A2(n8351), .ZN(n13139) );
  XNOR2_X1 U13018 ( .A(n13140), .B(n13141), .ZN(n12935) );
  XNOR2_X1 U13019 ( .A(n13142), .B(n13143), .ZN(n13141) );
  XNOR2_X1 U13020 ( .A(n13144), .B(n13145), .ZN(n12940) );
  XOR2_X1 U13021 ( .A(n13146), .B(n13147), .Z(n13145) );
  NAND2_X1 U13022 ( .A1(b_12_), .A2(a_22_), .ZN(n13147) );
  XNOR2_X1 U13023 ( .A(n13148), .B(n13149), .ZN(n12944) );
  XOR2_X1 U13024 ( .A(n13150), .B(n13151), .Z(n13148) );
  XNOR2_X1 U13025 ( .A(n13152), .B(n13153), .ZN(n12947) );
  XNOR2_X1 U13026 ( .A(n13154), .B(n13155), .ZN(n13152) );
  NOR2_X1 U13027 ( .A1(n8751), .A2(n8351), .ZN(n13155) );
  XOR2_X1 U13028 ( .A(n13156), .B(n13157), .Z(n12952) );
  NAND2_X1 U13029 ( .A1(n13158), .A2(n13159), .ZN(n13156) );
  XNOR2_X1 U13030 ( .A(n13160), .B(n13161), .ZN(n12956) );
  XOR2_X1 U13031 ( .A(n13162), .B(n13163), .Z(n13160) );
  XNOR2_X1 U13032 ( .A(n13164), .B(n13165), .ZN(n12960) );
  XOR2_X1 U13033 ( .A(n13166), .B(n13167), .Z(n13164) );
  XNOR2_X1 U13034 ( .A(n13168), .B(n13169), .ZN(n12850) );
  XNOR2_X1 U13035 ( .A(n13170), .B(n13171), .ZN(n13168) );
  NOR2_X1 U13036 ( .A1(n8755), .A2(n8351), .ZN(n13171) );
  XNOR2_X1 U13037 ( .A(n13172), .B(n13173), .ZN(n12844) );
  NAND2_X1 U13038 ( .A1(n13174), .A2(n13175), .ZN(n13172) );
  INV_X1 U13039 ( .A(n8694), .ZN(n12966) );
  NAND2_X1 U13040 ( .A1(b_13_), .A2(a_13_), .ZN(n8694) );
  XNOR2_X1 U13041 ( .A(n13176), .B(n13177), .ZN(n12968) );
  XNOR2_X1 U13042 ( .A(n13178), .B(n13179), .ZN(n13177) );
  XNOR2_X1 U13043 ( .A(n13180), .B(n13181), .ZN(n12971) );
  XNOR2_X1 U13044 ( .A(n13182), .B(n8691), .ZN(n13181) );
  XOR2_X1 U13045 ( .A(n13183), .B(n13184), .Z(n12976) );
  NAND2_X1 U13046 ( .A1(n13185), .A2(n13186), .ZN(n13183) );
  XNOR2_X1 U13047 ( .A(n13187), .B(n13188), .ZN(n12979) );
  NAND2_X1 U13048 ( .A1(n13189), .A2(n13190), .ZN(n13187) );
  XNOR2_X1 U13049 ( .A(n13191), .B(n13192), .ZN(n12984) );
  XOR2_X1 U13050 ( .A(n13193), .B(n13194), .Z(n13191) );
  XOR2_X1 U13051 ( .A(n13195), .B(n13196), .Z(n12817) );
  XOR2_X1 U13052 ( .A(n13197), .B(n13198), .Z(n13195) );
  NOR2_X1 U13053 ( .A1(n8763), .A2(n8351), .ZN(n13198) );
  XNOR2_X1 U13054 ( .A(n13199), .B(n13200), .ZN(n12809) );
  NAND2_X1 U13055 ( .A1(n13201), .A2(n13202), .ZN(n13199) );
  XNOR2_X1 U13056 ( .A(n13203), .B(n13204), .ZN(n12988) );
  XOR2_X1 U13057 ( .A(n13205), .B(n13206), .Z(n13203) );
  XNOR2_X1 U13058 ( .A(n13207), .B(n13208), .ZN(n12991) );
  XNOR2_X1 U13059 ( .A(n13209), .B(n13210), .ZN(n13207) );
  NOR2_X1 U13060 ( .A1(n8517), .A2(n8351), .ZN(n13210) );
  XNOR2_X1 U13061 ( .A(n13211), .B(n13212), .ZN(n12995) );
  XNOR2_X1 U13062 ( .A(n13213), .B(n13214), .ZN(n13212) );
  XNOR2_X1 U13063 ( .A(n13215), .B(n13216), .ZN(n13000) );
  XNOR2_X1 U13064 ( .A(n13217), .B(n13218), .ZN(n13215) );
  NOR2_X1 U13065 ( .A1(n8567), .A2(n8351), .ZN(n13218) );
  XNOR2_X1 U13066 ( .A(n13219), .B(n13220), .ZN(n13003) );
  XNOR2_X1 U13067 ( .A(n13221), .B(n13222), .ZN(n13219) );
  XNOR2_X1 U13068 ( .A(n13223), .B(n13224), .ZN(n13009) );
  XNOR2_X1 U13069 ( .A(n13225), .B(n13226), .ZN(n13224) );
  XOR2_X1 U13070 ( .A(n13227), .B(n13228), .Z(n13008) );
  XNOR2_X1 U13071 ( .A(n13229), .B(n13230), .ZN(n13228) );
  NAND4_X1 U13072 ( .A1(n8937), .A2(n8936), .A3(n8932), .A4(n8938), .ZN(n8906)
         );
  NAND2_X1 U13073 ( .A1(n13231), .A2(n13232), .ZN(n8938) );
  NAND2_X1 U13074 ( .A1(n13230), .A2(n13233), .ZN(n13232) );
  OR2_X1 U13075 ( .A1(n13229), .A2(n13227), .ZN(n13233) );
  NOR2_X1 U13076 ( .A1(n8351), .A2(n9674), .ZN(n13230) );
  NAND2_X1 U13077 ( .A1(n13227), .A2(n13229), .ZN(n13231) );
  NAND2_X1 U13078 ( .A1(n13234), .A2(n13235), .ZN(n13229) );
  NAND2_X1 U13079 ( .A1(n13226), .A2(n13236), .ZN(n13235) );
  OR2_X1 U13080 ( .A1(n13225), .A2(n13223), .ZN(n13236) );
  NOR2_X1 U13081 ( .A1(n8351), .A2(n8617), .ZN(n13226) );
  NAND2_X1 U13082 ( .A1(n13223), .A2(n13225), .ZN(n13234) );
  NAND2_X1 U13083 ( .A1(n13237), .A2(n13238), .ZN(n13225) );
  NAND2_X1 U13084 ( .A1(n13222), .A2(n13239), .ZN(n13238) );
  NAND2_X1 U13085 ( .A1(n13221), .A2(n13220), .ZN(n13239) );
  NOR2_X1 U13086 ( .A1(n8351), .A2(n8768), .ZN(n13222) );
  OR2_X1 U13087 ( .A1(n13220), .A2(n13221), .ZN(n13237) );
  AND2_X1 U13088 ( .A1(n13240), .A2(n13241), .ZN(n13221) );
  NAND3_X1 U13089 ( .A1(a_3_), .A2(n13242), .A3(b_12_), .ZN(n13241) );
  NAND2_X1 U13090 ( .A1(n13217), .A2(n13216), .ZN(n13242) );
  OR2_X1 U13091 ( .A1(n13216), .A2(n13217), .ZN(n13240) );
  AND2_X1 U13092 ( .A1(n13243), .A2(n13244), .ZN(n13217) );
  NAND2_X1 U13093 ( .A1(n13214), .A2(n13245), .ZN(n13244) );
  OR2_X1 U13094 ( .A1(n13213), .A2(n13211), .ZN(n13245) );
  NOR2_X1 U13095 ( .A1(n8351), .A2(n8766), .ZN(n13214) );
  NAND2_X1 U13096 ( .A1(n13211), .A2(n13213), .ZN(n13243) );
  NAND2_X1 U13097 ( .A1(n13246), .A2(n13247), .ZN(n13213) );
  NAND3_X1 U13098 ( .A1(a_5_), .A2(n13248), .A3(b_12_), .ZN(n13247) );
  NAND2_X1 U13099 ( .A1(n13209), .A2(n13208), .ZN(n13248) );
  OR2_X1 U13100 ( .A1(n13208), .A2(n13209), .ZN(n13246) );
  AND2_X1 U13101 ( .A1(n13249), .A2(n13250), .ZN(n13209) );
  NAND2_X1 U13102 ( .A1(n13206), .A2(n13251), .ZN(n13250) );
  OR2_X1 U13103 ( .A1(n13205), .A2(n13204), .ZN(n13251) );
  NOR2_X1 U13104 ( .A1(n8351), .A2(n8491), .ZN(n13206) );
  NAND2_X1 U13105 ( .A1(n13204), .A2(n13205), .ZN(n13249) );
  NAND2_X1 U13106 ( .A1(n13201), .A2(n13252), .ZN(n13205) );
  NAND2_X1 U13107 ( .A1(n13200), .A2(n13202), .ZN(n13252) );
  NAND2_X1 U13108 ( .A1(n13253), .A2(n13254), .ZN(n13202) );
  NAND2_X1 U13109 ( .A1(b_12_), .A2(a_7_), .ZN(n13254) );
  INV_X1 U13110 ( .A(n13255), .ZN(n13253) );
  XNOR2_X1 U13111 ( .A(n13256), .B(n13257), .ZN(n13200) );
  XOR2_X1 U13112 ( .A(n13258), .B(n13259), .Z(n13257) );
  NAND2_X1 U13113 ( .A1(b_11_), .A2(a_8_), .ZN(n13259) );
  NAND2_X1 U13114 ( .A1(a_7_), .A2(n13255), .ZN(n13201) );
  NAND2_X1 U13115 ( .A1(n13260), .A2(n13261), .ZN(n13255) );
  NAND3_X1 U13116 ( .A1(a_8_), .A2(n13262), .A3(b_12_), .ZN(n13261) );
  OR2_X1 U13117 ( .A1(n13197), .A2(n13196), .ZN(n13262) );
  NAND2_X1 U13118 ( .A1(n13196), .A2(n13197), .ZN(n13260) );
  NAND2_X1 U13119 ( .A1(n13263), .A2(n13264), .ZN(n13197) );
  NAND2_X1 U13120 ( .A1(n13194), .A2(n13265), .ZN(n13264) );
  OR2_X1 U13121 ( .A1(n13193), .A2(n13192), .ZN(n13265) );
  NOR2_X1 U13122 ( .A1(n8351), .A2(n8426), .ZN(n13194) );
  NAND2_X1 U13123 ( .A1(n13192), .A2(n13193), .ZN(n13263) );
  NAND2_X1 U13124 ( .A1(n13189), .A2(n13266), .ZN(n13193) );
  NAND2_X1 U13125 ( .A1(n13188), .A2(n13190), .ZN(n13266) );
  NAND2_X1 U13126 ( .A1(n13267), .A2(n13268), .ZN(n13190) );
  NAND2_X1 U13127 ( .A1(b_12_), .A2(a_10_), .ZN(n13268) );
  INV_X1 U13128 ( .A(n13269), .ZN(n13267) );
  XOR2_X1 U13129 ( .A(n13270), .B(n13271), .Z(n13188) );
  XOR2_X1 U13130 ( .A(n13272), .B(n13273), .Z(n13270) );
  NAND2_X1 U13131 ( .A1(a_10_), .A2(n13269), .ZN(n13189) );
  NAND2_X1 U13132 ( .A1(n13185), .A2(n13274), .ZN(n13269) );
  NAND2_X1 U13133 ( .A1(n13184), .A2(n13186), .ZN(n13274) );
  NAND2_X1 U13134 ( .A1(n13275), .A2(n13276), .ZN(n13186) );
  NAND2_X1 U13135 ( .A1(b_12_), .A2(a_11_), .ZN(n13276) );
  INV_X1 U13136 ( .A(n13277), .ZN(n13275) );
  XOR2_X1 U13137 ( .A(n13278), .B(n13279), .Z(n13184) );
  XOR2_X1 U13138 ( .A(n13280), .B(n13281), .Z(n13278) );
  NOR2_X1 U13139 ( .A1(n8759), .A2(n8760), .ZN(n13281) );
  NAND2_X1 U13140 ( .A1(a_11_), .A2(n13277), .ZN(n13185) );
  NAND2_X1 U13141 ( .A1(n13282), .A2(n13283), .ZN(n13277) );
  NAND2_X1 U13142 ( .A1(n13180), .A2(n13284), .ZN(n13283) );
  OR2_X1 U13143 ( .A1(n13182), .A2(n8691), .ZN(n13284) );
  XNOR2_X1 U13144 ( .A(n13285), .B(n13286), .ZN(n13180) );
  XOR2_X1 U13145 ( .A(n13287), .B(n13288), .Z(n13286) );
  NAND2_X1 U13146 ( .A1(b_11_), .A2(a_13_), .ZN(n13288) );
  NAND2_X1 U13147 ( .A1(n8691), .A2(n13182), .ZN(n13282) );
  NAND2_X1 U13148 ( .A1(n13289), .A2(n13290), .ZN(n13182) );
  NAND2_X1 U13149 ( .A1(n13179), .A2(n13291), .ZN(n13290) );
  OR2_X1 U13150 ( .A1(n13178), .A2(n13176), .ZN(n13291) );
  NOR2_X1 U13151 ( .A1(n8351), .A2(n8310), .ZN(n13179) );
  NAND2_X1 U13152 ( .A1(n13176), .A2(n13178), .ZN(n13289) );
  NAND2_X1 U13153 ( .A1(n13058), .A2(n13292), .ZN(n13178) );
  NAND2_X1 U13154 ( .A1(n13057), .A2(n13059), .ZN(n13292) );
  NAND2_X1 U13155 ( .A1(n13293), .A2(n13294), .ZN(n13059) );
  NAND2_X1 U13156 ( .A1(b_12_), .A2(a_14_), .ZN(n13294) );
  INV_X1 U13157 ( .A(n13295), .ZN(n13293) );
  XNOR2_X1 U13158 ( .A(n13296), .B(n13297), .ZN(n13057) );
  XOR2_X1 U13159 ( .A(n13298), .B(n13299), .Z(n13297) );
  NAND2_X1 U13160 ( .A1(b_11_), .A2(a_15_), .ZN(n13299) );
  NAND2_X1 U13161 ( .A1(a_14_), .A2(n13295), .ZN(n13058) );
  NAND2_X1 U13162 ( .A1(n13174), .A2(n13300), .ZN(n13295) );
  NAND2_X1 U13163 ( .A1(n13173), .A2(n13175), .ZN(n13300) );
  NAND2_X1 U13164 ( .A1(n13301), .A2(n13302), .ZN(n13175) );
  NAND2_X1 U13165 ( .A1(b_12_), .A2(a_15_), .ZN(n13302) );
  INV_X1 U13166 ( .A(n13303), .ZN(n13301) );
  XNOR2_X1 U13167 ( .A(n13304), .B(n13305), .ZN(n13173) );
  XOR2_X1 U13168 ( .A(n13306), .B(n13307), .Z(n13305) );
  NAND2_X1 U13169 ( .A1(b_11_), .A2(a_16_), .ZN(n13307) );
  NAND2_X1 U13170 ( .A1(a_15_), .A2(n13303), .ZN(n13174) );
  NAND2_X1 U13171 ( .A1(n13308), .A2(n13309), .ZN(n13303) );
  NAND3_X1 U13172 ( .A1(a_16_), .A2(n13310), .A3(b_12_), .ZN(n13309) );
  NAND2_X1 U13173 ( .A1(n13170), .A2(n13169), .ZN(n13310) );
  OR2_X1 U13174 ( .A1(n13169), .A2(n13170), .ZN(n13308) );
  AND2_X1 U13175 ( .A1(n13311), .A2(n13312), .ZN(n13170) );
  NAND2_X1 U13176 ( .A1(n13166), .A2(n13313), .ZN(n13312) );
  OR2_X1 U13177 ( .A1(n13167), .A2(n13165), .ZN(n13313) );
  NOR2_X1 U13178 ( .A1(n8351), .A2(n8210), .ZN(n13166) );
  NAND2_X1 U13179 ( .A1(n13165), .A2(n13167), .ZN(n13311) );
  NAND2_X1 U13180 ( .A1(n13314), .A2(n13315), .ZN(n13167) );
  NAND2_X1 U13181 ( .A1(n13162), .A2(n13316), .ZN(n13315) );
  OR2_X1 U13182 ( .A1(n13163), .A2(n13161), .ZN(n13316) );
  NOR2_X1 U13183 ( .A1(n8351), .A2(n8753), .ZN(n13162) );
  NAND2_X1 U13184 ( .A1(n13161), .A2(n13163), .ZN(n13314) );
  NAND2_X1 U13185 ( .A1(n13158), .A2(n13317), .ZN(n13163) );
  NAND2_X1 U13186 ( .A1(n13157), .A2(n13159), .ZN(n13317) );
  NAND2_X1 U13187 ( .A1(n13318), .A2(n13319), .ZN(n13159) );
  NAND2_X1 U13188 ( .A1(b_12_), .A2(a_19_), .ZN(n13319) );
  INV_X1 U13189 ( .A(n13320), .ZN(n13318) );
  XOR2_X1 U13190 ( .A(n13321), .B(n13322), .Z(n13157) );
  XOR2_X1 U13191 ( .A(n13323), .B(n13324), .Z(n13321) );
  NOR2_X1 U13192 ( .A1(n8751), .A2(n8760), .ZN(n13324) );
  NAND2_X1 U13193 ( .A1(a_19_), .A2(n13320), .ZN(n13158) );
  NAND2_X1 U13194 ( .A1(n13325), .A2(n13326), .ZN(n13320) );
  NAND3_X1 U13195 ( .A1(a_20_), .A2(n13327), .A3(b_12_), .ZN(n13326) );
  NAND2_X1 U13196 ( .A1(n13154), .A2(n13153), .ZN(n13327) );
  OR2_X1 U13197 ( .A1(n13153), .A2(n13154), .ZN(n13325) );
  AND2_X1 U13198 ( .A1(n13328), .A2(n13329), .ZN(n13154) );
  NAND2_X1 U13199 ( .A1(n13151), .A2(n13330), .ZN(n13329) );
  OR2_X1 U13200 ( .A1(n13150), .A2(n13149), .ZN(n13330) );
  NOR2_X1 U13201 ( .A1(n8351), .A2(n8750), .ZN(n13151) );
  NAND2_X1 U13202 ( .A1(n13149), .A2(n13150), .ZN(n13328) );
  NAND2_X1 U13203 ( .A1(n13331), .A2(n13332), .ZN(n13150) );
  NAND3_X1 U13204 ( .A1(a_22_), .A2(n13333), .A3(b_12_), .ZN(n13332) );
  OR2_X1 U13205 ( .A1(n13146), .A2(n13144), .ZN(n13333) );
  NAND2_X1 U13206 ( .A1(n13144), .A2(n13146), .ZN(n13331) );
  NAND2_X1 U13207 ( .A1(n13334), .A2(n13335), .ZN(n13146) );
  NAND2_X1 U13208 ( .A1(n13143), .A2(n13336), .ZN(n13335) );
  OR2_X1 U13209 ( .A1(n13142), .A2(n13140), .ZN(n13336) );
  NOR2_X1 U13210 ( .A1(n8351), .A2(n8747), .ZN(n13143) );
  NAND2_X1 U13211 ( .A1(n13140), .A2(n13142), .ZN(n13334) );
  NAND2_X1 U13212 ( .A1(n13337), .A2(n13338), .ZN(n13142) );
  NAND3_X1 U13213 ( .A1(a_24_), .A2(n13339), .A3(b_12_), .ZN(n13338) );
  NAND2_X1 U13214 ( .A1(n13138), .A2(n13137), .ZN(n13339) );
  OR2_X1 U13215 ( .A1(n13137), .A2(n13138), .ZN(n13337) );
  AND2_X1 U13216 ( .A1(n13340), .A2(n13341), .ZN(n13138) );
  NAND2_X1 U13217 ( .A1(n13135), .A2(n13342), .ZN(n13341) );
  OR2_X1 U13218 ( .A1(n13134), .A2(n13133), .ZN(n13342) );
  NOR2_X1 U13219 ( .A1(n8351), .A2(n8744), .ZN(n13135) );
  NAND2_X1 U13220 ( .A1(n13133), .A2(n13134), .ZN(n13340) );
  NAND2_X1 U13221 ( .A1(n13130), .A2(n13343), .ZN(n13134) );
  NAND2_X1 U13222 ( .A1(n13129), .A2(n13131), .ZN(n13343) );
  NAND2_X1 U13223 ( .A1(n13344), .A2(n13345), .ZN(n13131) );
  NAND2_X1 U13224 ( .A1(b_12_), .A2(a_26_), .ZN(n13345) );
  INV_X1 U13225 ( .A(n13346), .ZN(n13344) );
  XNOR2_X1 U13226 ( .A(n13347), .B(n13348), .ZN(n13129) );
  NAND2_X1 U13227 ( .A1(n13349), .A2(n13350), .ZN(n13347) );
  NAND2_X1 U13228 ( .A1(a_26_), .A2(n13346), .ZN(n13130) );
  NAND2_X1 U13229 ( .A1(n13102), .A2(n13351), .ZN(n13346) );
  NAND2_X1 U13230 ( .A1(n13101), .A2(n13103), .ZN(n13351) );
  NAND2_X1 U13231 ( .A1(n13352), .A2(n13353), .ZN(n13103) );
  NAND2_X1 U13232 ( .A1(b_12_), .A2(a_27_), .ZN(n13353) );
  INV_X1 U13233 ( .A(n13354), .ZN(n13352) );
  XNOR2_X1 U13234 ( .A(n13355), .B(n13356), .ZN(n13101) );
  XOR2_X1 U13235 ( .A(n13357), .B(n13358), .Z(n13355) );
  NAND2_X1 U13236 ( .A1(b_11_), .A2(a_28_), .ZN(n13357) );
  NAND2_X1 U13237 ( .A1(a_27_), .A2(n13354), .ZN(n13102) );
  NAND2_X1 U13238 ( .A1(n13359), .A2(n13360), .ZN(n13354) );
  NAND3_X1 U13239 ( .A1(a_28_), .A2(n13361), .A3(b_12_), .ZN(n13360) );
  NAND2_X1 U13240 ( .A1(n13111), .A2(n13109), .ZN(n13361) );
  OR2_X1 U13241 ( .A1(n13109), .A2(n13111), .ZN(n13359) );
  AND2_X1 U13242 ( .A1(n13362), .A2(n13363), .ZN(n13111) );
  NAND2_X1 U13243 ( .A1(n13125), .A2(n13364), .ZN(n13363) );
  OR2_X1 U13244 ( .A1(n13126), .A2(n13127), .ZN(n13364) );
  NOR2_X1 U13245 ( .A1(n8351), .A2(n7890), .ZN(n13125) );
  NAND2_X1 U13246 ( .A1(n13127), .A2(n13126), .ZN(n13362) );
  NAND2_X1 U13247 ( .A1(n13365), .A2(n13366), .ZN(n13126) );
  NAND2_X1 U13248 ( .A1(b_10_), .A2(n13367), .ZN(n13366) );
  NAND2_X1 U13249 ( .A1(n7864), .A2(n13368), .ZN(n13367) );
  NAND2_X1 U13250 ( .A1(a_31_), .A2(n8760), .ZN(n13368) );
  NAND2_X1 U13251 ( .A1(b_11_), .A2(n13369), .ZN(n13365) );
  NAND2_X1 U13252 ( .A1(n9137), .A2(n13370), .ZN(n13369) );
  NAND2_X1 U13253 ( .A1(a_30_), .A2(n8401), .ZN(n13370) );
  AND3_X1 U13254 ( .A1(b_11_), .A2(b_12_), .A3(n7818), .ZN(n13127) );
  XNOR2_X1 U13255 ( .A(n13371), .B(n13372), .ZN(n13109) );
  XOR2_X1 U13256 ( .A(n13373), .B(n13374), .Z(n13371) );
  XNOR2_X1 U13257 ( .A(n13375), .B(n13376), .ZN(n13133) );
  NAND2_X1 U13258 ( .A1(n13377), .A2(n13378), .ZN(n13375) );
  XNOR2_X1 U13259 ( .A(n13379), .B(n13380), .ZN(n13137) );
  XOR2_X1 U13260 ( .A(n13381), .B(n13382), .Z(n13379) );
  XNOR2_X1 U13261 ( .A(n13383), .B(n13384), .ZN(n13140) );
  XNOR2_X1 U13262 ( .A(n13385), .B(n13386), .ZN(n13383) );
  NOR2_X1 U13263 ( .A1(n8745), .A2(n8760), .ZN(n13386) );
  XNOR2_X1 U13264 ( .A(n13387), .B(n13388), .ZN(n13144) );
  XNOR2_X1 U13265 ( .A(n13389), .B(n13390), .ZN(n13388) );
  XNOR2_X1 U13266 ( .A(n13391), .B(n13392), .ZN(n13149) );
  XOR2_X1 U13267 ( .A(n13393), .B(n13394), .Z(n13392) );
  NAND2_X1 U13268 ( .A1(b_11_), .A2(a_22_), .ZN(n13394) );
  XNOR2_X1 U13269 ( .A(n13395), .B(n13396), .ZN(n13153) );
  XOR2_X1 U13270 ( .A(n13397), .B(n13398), .Z(n13395) );
  XNOR2_X1 U13271 ( .A(n13399), .B(n13400), .ZN(n13161) );
  NAND2_X1 U13272 ( .A1(n13401), .A2(n13402), .ZN(n13399) );
  XNOR2_X1 U13273 ( .A(n13403), .B(n13404), .ZN(n13165) );
  NAND2_X1 U13274 ( .A1(n13405), .A2(n13406), .ZN(n13403) );
  XNOR2_X1 U13275 ( .A(n13407), .B(n13408), .ZN(n13169) );
  XOR2_X1 U13276 ( .A(n13409), .B(n13410), .Z(n13407) );
  NOR2_X1 U13277 ( .A1(n8210), .A2(n8760), .ZN(n13410) );
  XOR2_X1 U13278 ( .A(n13411), .B(n13412), .Z(n13176) );
  XOR2_X1 U13279 ( .A(n13413), .B(n13414), .Z(n13411) );
  NOR2_X1 U13280 ( .A1(n8757), .A2(n8760), .ZN(n13414) );
  NOR2_X1 U13281 ( .A1(n8351), .A2(n8759), .ZN(n8691) );
  XNOR2_X1 U13282 ( .A(n13415), .B(n13416), .ZN(n13192) );
  XNOR2_X1 U13283 ( .A(n13417), .B(n13418), .ZN(n13415) );
  NOR2_X1 U13284 ( .A1(n8761), .A2(n8760), .ZN(n13418) );
  XNOR2_X1 U13285 ( .A(n13419), .B(n13420), .ZN(n13196) );
  XOR2_X1 U13286 ( .A(n13421), .B(n13422), .Z(n13420) );
  NAND2_X1 U13287 ( .A1(b_11_), .A2(a_9_), .ZN(n13422) );
  XNOR2_X1 U13288 ( .A(n13423), .B(n13424), .ZN(n13204) );
  XNOR2_X1 U13289 ( .A(n13425), .B(n13426), .ZN(n13423) );
  NOR2_X1 U13290 ( .A1(n8764), .A2(n8760), .ZN(n13426) );
  XNOR2_X1 U13291 ( .A(n13427), .B(n13428), .ZN(n13208) );
  XOR2_X1 U13292 ( .A(n13429), .B(n13430), .Z(n13427) );
  NOR2_X1 U13293 ( .A1(n8491), .A2(n8760), .ZN(n13430) );
  XNOR2_X1 U13294 ( .A(n13431), .B(n13432), .ZN(n13211) );
  XOR2_X1 U13295 ( .A(n13433), .B(n13434), .Z(n13432) );
  NAND2_X1 U13296 ( .A1(b_11_), .A2(a_5_), .ZN(n13434) );
  XOR2_X1 U13297 ( .A(n13435), .B(n13436), .Z(n13216) );
  XOR2_X1 U13298 ( .A(n13437), .B(n13438), .Z(n13436) );
  NAND2_X1 U13299 ( .A1(b_11_), .A2(a_4_), .ZN(n13438) );
  XNOR2_X1 U13300 ( .A(n13439), .B(n13440), .ZN(n13220) );
  XOR2_X1 U13301 ( .A(n13441), .B(n13442), .Z(n13439) );
  NOR2_X1 U13302 ( .A1(n8567), .A2(n8760), .ZN(n13442) );
  XOR2_X1 U13303 ( .A(n13443), .B(n13444), .Z(n13223) );
  XOR2_X1 U13304 ( .A(n13445), .B(n13446), .Z(n13443) );
  NOR2_X1 U13305 ( .A1(n8768), .A2(n8760), .ZN(n13446) );
  XNOR2_X1 U13306 ( .A(n13447), .B(n13448), .ZN(n13227) );
  XOR2_X1 U13307 ( .A(n13449), .B(n13450), .Z(n13448) );
  NAND2_X1 U13308 ( .A1(b_11_), .A2(a_1_), .ZN(n13450) );
  NAND3_X1 U13309 ( .A1(n13451), .A2(n13452), .A3(n13453), .ZN(n8936) );
  XOR2_X1 U13310 ( .A(n13454), .B(n13455), .Z(n13453) );
  XOR2_X1 U13311 ( .A(n13456), .B(n13457), .Z(n8937) );
  XOR2_X1 U13312 ( .A(n13458), .B(n13459), .Z(n13456) );
  OR2_X1 U13313 ( .A1(n8932), .A2(n8931), .ZN(n8912) );
  XNOR2_X1 U13314 ( .A(n13460), .B(n13461), .ZN(n8931) );
  NAND2_X1 U13315 ( .A1(n13462), .A2(n13463), .ZN(n8932) );
  NAND2_X1 U13316 ( .A1(n13451), .A2(n13452), .ZN(n13463) );
  NAND2_X1 U13317 ( .A1(n13459), .A2(n13464), .ZN(n13452) );
  OR2_X1 U13318 ( .A1(n13458), .A2(n13457), .ZN(n13464) );
  NOR2_X1 U13319 ( .A1(n8760), .A2(n9674), .ZN(n13459) );
  NAND2_X1 U13320 ( .A1(n13457), .A2(n13458), .ZN(n13451) );
  NAND2_X1 U13321 ( .A1(n13465), .A2(n13466), .ZN(n13458) );
  NAND3_X1 U13322 ( .A1(a_1_), .A2(n13467), .A3(b_11_), .ZN(n13466) );
  OR2_X1 U13323 ( .A1(n13449), .A2(n13447), .ZN(n13467) );
  NAND2_X1 U13324 ( .A1(n13447), .A2(n13449), .ZN(n13465) );
  NAND2_X1 U13325 ( .A1(n13468), .A2(n13469), .ZN(n13449) );
  NAND3_X1 U13326 ( .A1(a_2_), .A2(n13470), .A3(b_11_), .ZN(n13469) );
  OR2_X1 U13327 ( .A1(n13445), .A2(n13444), .ZN(n13470) );
  NAND2_X1 U13328 ( .A1(n13444), .A2(n13445), .ZN(n13468) );
  NAND2_X1 U13329 ( .A1(n13471), .A2(n13472), .ZN(n13445) );
  NAND3_X1 U13330 ( .A1(a_3_), .A2(n13473), .A3(b_11_), .ZN(n13472) );
  OR2_X1 U13331 ( .A1(n13441), .A2(n13440), .ZN(n13473) );
  NAND2_X1 U13332 ( .A1(n13440), .A2(n13441), .ZN(n13471) );
  NAND2_X1 U13333 ( .A1(n13474), .A2(n13475), .ZN(n13441) );
  NAND3_X1 U13334 ( .A1(a_4_), .A2(n13476), .A3(b_11_), .ZN(n13475) );
  OR2_X1 U13335 ( .A1(n13437), .A2(n13435), .ZN(n13476) );
  NAND2_X1 U13336 ( .A1(n13435), .A2(n13437), .ZN(n13474) );
  NAND2_X1 U13337 ( .A1(n13477), .A2(n13478), .ZN(n13437) );
  NAND3_X1 U13338 ( .A1(a_5_), .A2(n13479), .A3(b_11_), .ZN(n13478) );
  OR2_X1 U13339 ( .A1(n13433), .A2(n13431), .ZN(n13479) );
  NAND2_X1 U13340 ( .A1(n13431), .A2(n13433), .ZN(n13477) );
  NAND2_X1 U13341 ( .A1(n13480), .A2(n13481), .ZN(n13433) );
  NAND3_X1 U13342 ( .A1(a_6_), .A2(n13482), .A3(b_11_), .ZN(n13481) );
  OR2_X1 U13343 ( .A1(n13429), .A2(n13428), .ZN(n13482) );
  NAND2_X1 U13344 ( .A1(n13428), .A2(n13429), .ZN(n13480) );
  NAND2_X1 U13345 ( .A1(n13483), .A2(n13484), .ZN(n13429) );
  NAND3_X1 U13346 ( .A1(a_7_), .A2(n13485), .A3(b_11_), .ZN(n13484) );
  NAND2_X1 U13347 ( .A1(n13425), .A2(n13424), .ZN(n13485) );
  OR2_X1 U13348 ( .A1(n13424), .A2(n13425), .ZN(n13483) );
  AND2_X1 U13349 ( .A1(n13486), .A2(n13487), .ZN(n13425) );
  NAND3_X1 U13350 ( .A1(a_8_), .A2(n13488), .A3(b_11_), .ZN(n13487) );
  OR2_X1 U13351 ( .A1(n13258), .A2(n13256), .ZN(n13488) );
  NAND2_X1 U13352 ( .A1(n13256), .A2(n13258), .ZN(n13486) );
  NAND2_X1 U13353 ( .A1(n13489), .A2(n13490), .ZN(n13258) );
  NAND3_X1 U13354 ( .A1(a_9_), .A2(n13491), .A3(b_11_), .ZN(n13490) );
  OR2_X1 U13355 ( .A1(n13421), .A2(n13419), .ZN(n13491) );
  NAND2_X1 U13356 ( .A1(n13419), .A2(n13421), .ZN(n13489) );
  NAND2_X1 U13357 ( .A1(n13492), .A2(n13493), .ZN(n13421) );
  NAND3_X1 U13358 ( .A1(a_10_), .A2(n13494), .A3(b_11_), .ZN(n13493) );
  NAND2_X1 U13359 ( .A1(n13417), .A2(n13416), .ZN(n13494) );
  OR2_X1 U13360 ( .A1(n13416), .A2(n13417), .ZN(n13492) );
  AND2_X1 U13361 ( .A1(n13495), .A2(n13496), .ZN(n13417) );
  NAND2_X1 U13362 ( .A1(n13271), .A2(n13497), .ZN(n13496) );
  OR2_X1 U13363 ( .A1(n13272), .A2(n13273), .ZN(n13497) );
  XNOR2_X1 U13364 ( .A(n13498), .B(n13499), .ZN(n13271) );
  NAND2_X1 U13365 ( .A1(n13500), .A2(n13501), .ZN(n13498) );
  NAND2_X1 U13366 ( .A1(n13273), .A2(n13272), .ZN(n13495) );
  NAND2_X1 U13367 ( .A1(n13502), .A2(n13503), .ZN(n13272) );
  NAND3_X1 U13368 ( .A1(a_12_), .A2(n13504), .A3(b_11_), .ZN(n13503) );
  OR2_X1 U13369 ( .A1(n13280), .A2(n13279), .ZN(n13504) );
  NAND2_X1 U13370 ( .A1(n13279), .A2(n13280), .ZN(n13502) );
  NAND2_X1 U13371 ( .A1(n13505), .A2(n13506), .ZN(n13280) );
  NAND3_X1 U13372 ( .A1(a_13_), .A2(n13507), .A3(b_11_), .ZN(n13506) );
  OR2_X1 U13373 ( .A1(n13287), .A2(n13285), .ZN(n13507) );
  NAND2_X1 U13374 ( .A1(n13285), .A2(n13287), .ZN(n13505) );
  NAND2_X1 U13375 ( .A1(n13508), .A2(n13509), .ZN(n13287) );
  NAND3_X1 U13376 ( .A1(a_14_), .A2(n13510), .A3(b_11_), .ZN(n13509) );
  OR2_X1 U13377 ( .A1(n13413), .A2(n13412), .ZN(n13510) );
  NAND2_X1 U13378 ( .A1(n13412), .A2(n13413), .ZN(n13508) );
  NAND2_X1 U13379 ( .A1(n13511), .A2(n13512), .ZN(n13413) );
  NAND3_X1 U13380 ( .A1(a_15_), .A2(n13513), .A3(b_11_), .ZN(n13512) );
  OR2_X1 U13381 ( .A1(n13298), .A2(n13296), .ZN(n13513) );
  NAND2_X1 U13382 ( .A1(n13296), .A2(n13298), .ZN(n13511) );
  NAND2_X1 U13383 ( .A1(n13514), .A2(n13515), .ZN(n13298) );
  NAND3_X1 U13384 ( .A1(a_16_), .A2(n13516), .A3(b_11_), .ZN(n13515) );
  OR2_X1 U13385 ( .A1(n13306), .A2(n13304), .ZN(n13516) );
  NAND2_X1 U13386 ( .A1(n13304), .A2(n13306), .ZN(n13514) );
  NAND2_X1 U13387 ( .A1(n13517), .A2(n13518), .ZN(n13306) );
  NAND3_X1 U13388 ( .A1(a_17_), .A2(n13519), .A3(b_11_), .ZN(n13518) );
  OR2_X1 U13389 ( .A1(n13409), .A2(n13408), .ZN(n13519) );
  NAND2_X1 U13390 ( .A1(n13408), .A2(n13409), .ZN(n13517) );
  NAND2_X1 U13391 ( .A1(n13405), .A2(n13520), .ZN(n13409) );
  NAND2_X1 U13392 ( .A1(n13404), .A2(n13406), .ZN(n13520) );
  NAND2_X1 U13393 ( .A1(n13521), .A2(n13522), .ZN(n13406) );
  NAND2_X1 U13394 ( .A1(b_11_), .A2(a_18_), .ZN(n13522) );
  INV_X1 U13395 ( .A(n13523), .ZN(n13521) );
  XNOR2_X1 U13396 ( .A(n13524), .B(n13525), .ZN(n13404) );
  XNOR2_X1 U13397 ( .A(n13526), .B(n13527), .ZN(n13524) );
  NAND2_X1 U13398 ( .A1(a_18_), .A2(n13523), .ZN(n13405) );
  NAND2_X1 U13399 ( .A1(n13401), .A2(n13528), .ZN(n13523) );
  NAND2_X1 U13400 ( .A1(n13400), .A2(n13402), .ZN(n13528) );
  NAND2_X1 U13401 ( .A1(n13529), .A2(n13530), .ZN(n13402) );
  NAND2_X1 U13402 ( .A1(b_11_), .A2(a_19_), .ZN(n13530) );
  INV_X1 U13403 ( .A(n13531), .ZN(n13529) );
  XNOR2_X1 U13404 ( .A(n13532), .B(n13533), .ZN(n13400) );
  XNOR2_X1 U13405 ( .A(n13534), .B(n13535), .ZN(n13533) );
  NAND2_X1 U13406 ( .A1(a_19_), .A2(n13531), .ZN(n13401) );
  NAND2_X1 U13407 ( .A1(n13536), .A2(n13537), .ZN(n13531) );
  NAND3_X1 U13408 ( .A1(a_20_), .A2(n13538), .A3(b_11_), .ZN(n13537) );
  OR2_X1 U13409 ( .A1(n13323), .A2(n13322), .ZN(n13538) );
  NAND2_X1 U13410 ( .A1(n13322), .A2(n13323), .ZN(n13536) );
  NAND2_X1 U13411 ( .A1(n13539), .A2(n13540), .ZN(n13323) );
  NAND2_X1 U13412 ( .A1(n13398), .A2(n13541), .ZN(n13540) );
  OR2_X1 U13413 ( .A1(n13397), .A2(n13396), .ZN(n13541) );
  NOR2_X1 U13414 ( .A1(n8760), .A2(n8750), .ZN(n13398) );
  NAND2_X1 U13415 ( .A1(n13396), .A2(n13397), .ZN(n13539) );
  NAND2_X1 U13416 ( .A1(n13542), .A2(n13543), .ZN(n13397) );
  NAND3_X1 U13417 ( .A1(a_22_), .A2(n13544), .A3(b_11_), .ZN(n13543) );
  OR2_X1 U13418 ( .A1(n13393), .A2(n13391), .ZN(n13544) );
  NAND2_X1 U13419 ( .A1(n13391), .A2(n13393), .ZN(n13542) );
  NAND2_X1 U13420 ( .A1(n13545), .A2(n13546), .ZN(n13393) );
  NAND2_X1 U13421 ( .A1(n13390), .A2(n13547), .ZN(n13546) );
  OR2_X1 U13422 ( .A1(n13389), .A2(n13387), .ZN(n13547) );
  NOR2_X1 U13423 ( .A1(n8760), .A2(n8747), .ZN(n13390) );
  NAND2_X1 U13424 ( .A1(n13387), .A2(n13389), .ZN(n13545) );
  NAND2_X1 U13425 ( .A1(n13548), .A2(n13549), .ZN(n13389) );
  NAND3_X1 U13426 ( .A1(a_24_), .A2(n13550), .A3(b_11_), .ZN(n13549) );
  NAND2_X1 U13427 ( .A1(n13385), .A2(n13384), .ZN(n13550) );
  OR2_X1 U13428 ( .A1(n13384), .A2(n13385), .ZN(n13548) );
  AND2_X1 U13429 ( .A1(n13551), .A2(n13552), .ZN(n13385) );
  NAND2_X1 U13430 ( .A1(n13382), .A2(n13553), .ZN(n13552) );
  OR2_X1 U13431 ( .A1(n13381), .A2(n13380), .ZN(n13553) );
  NOR2_X1 U13432 ( .A1(n8760), .A2(n8744), .ZN(n13382) );
  NAND2_X1 U13433 ( .A1(n13380), .A2(n13381), .ZN(n13551) );
  NAND2_X1 U13434 ( .A1(n13377), .A2(n13554), .ZN(n13381) );
  NAND2_X1 U13435 ( .A1(n13376), .A2(n13378), .ZN(n13554) );
  NAND2_X1 U13436 ( .A1(n13555), .A2(n13556), .ZN(n13378) );
  NAND2_X1 U13437 ( .A1(b_11_), .A2(a_26_), .ZN(n13556) );
  INV_X1 U13438 ( .A(n13557), .ZN(n13555) );
  XNOR2_X1 U13439 ( .A(n13558), .B(n13559), .ZN(n13376) );
  NAND2_X1 U13440 ( .A1(n13560), .A2(n13561), .ZN(n13558) );
  NAND2_X1 U13441 ( .A1(a_26_), .A2(n13557), .ZN(n13377) );
  NAND2_X1 U13442 ( .A1(n13349), .A2(n13562), .ZN(n13557) );
  NAND2_X1 U13443 ( .A1(n13348), .A2(n13350), .ZN(n13562) );
  NAND2_X1 U13444 ( .A1(n13563), .A2(n13564), .ZN(n13350) );
  NAND2_X1 U13445 ( .A1(b_11_), .A2(a_27_), .ZN(n13564) );
  INV_X1 U13446 ( .A(n13565), .ZN(n13563) );
  XNOR2_X1 U13447 ( .A(n13566), .B(n13567), .ZN(n13348) );
  XOR2_X1 U13448 ( .A(n13568), .B(n13569), .Z(n13566) );
  NAND2_X1 U13449 ( .A1(b_10_), .A2(a_28_), .ZN(n13568) );
  NAND2_X1 U13450 ( .A1(a_27_), .A2(n13565), .ZN(n13349) );
  NAND2_X1 U13451 ( .A1(n13570), .A2(n13571), .ZN(n13565) );
  NAND3_X1 U13452 ( .A1(a_28_), .A2(n13572), .A3(b_11_), .ZN(n13571) );
  NAND2_X1 U13453 ( .A1(n13358), .A2(n13356), .ZN(n13572) );
  OR2_X1 U13454 ( .A1(n13356), .A2(n13358), .ZN(n13570) );
  AND2_X1 U13455 ( .A1(n13573), .A2(n13574), .ZN(n13358) );
  NAND2_X1 U13456 ( .A1(n13372), .A2(n13575), .ZN(n13574) );
  OR2_X1 U13457 ( .A1(n13373), .A2(n13374), .ZN(n13575) );
  NOR2_X1 U13458 ( .A1(n8760), .A2(n7890), .ZN(n13372) );
  NAND2_X1 U13459 ( .A1(n13374), .A2(n13373), .ZN(n13573) );
  NAND2_X1 U13460 ( .A1(n13576), .A2(n13577), .ZN(n13373) );
  NAND2_X1 U13461 ( .A1(b_10_), .A2(n13578), .ZN(n13577) );
  NAND2_X1 U13462 ( .A1(n9137), .A2(n13579), .ZN(n13578) );
  NAND2_X1 U13463 ( .A1(a_30_), .A2(n8762), .ZN(n13579) );
  NAND2_X1 U13464 ( .A1(b_9_), .A2(n13580), .ZN(n13576) );
  NAND2_X1 U13465 ( .A1(n7864), .A2(n13581), .ZN(n13580) );
  NAND2_X1 U13466 ( .A1(a_31_), .A2(n8401), .ZN(n13581) );
  AND3_X1 U13467 ( .A1(b_10_), .A2(b_11_), .A3(n7818), .ZN(n13374) );
  XNOR2_X1 U13468 ( .A(n13582), .B(n13583), .ZN(n13356) );
  XOR2_X1 U13469 ( .A(n13584), .B(n13585), .Z(n13582) );
  XNOR2_X1 U13470 ( .A(n13586), .B(n13587), .ZN(n13380) );
  NAND2_X1 U13471 ( .A1(n13588), .A2(n13589), .ZN(n13586) );
  XNOR2_X1 U13472 ( .A(n13590), .B(n13591), .ZN(n13384) );
  XOR2_X1 U13473 ( .A(n13592), .B(n13593), .Z(n13590) );
  XNOR2_X1 U13474 ( .A(n13594), .B(n13595), .ZN(n13387) );
  XNOR2_X1 U13475 ( .A(n13596), .B(n13597), .ZN(n13594) );
  NOR2_X1 U13476 ( .A1(n8745), .A2(n8401), .ZN(n13597) );
  XNOR2_X1 U13477 ( .A(n13598), .B(n13599), .ZN(n13391) );
  XNOR2_X1 U13478 ( .A(n13600), .B(n13601), .ZN(n13599) );
  XNOR2_X1 U13479 ( .A(n13602), .B(n13603), .ZN(n13396) );
  XOR2_X1 U13480 ( .A(n13604), .B(n13605), .Z(n13603) );
  NAND2_X1 U13481 ( .A1(b_10_), .A2(a_22_), .ZN(n13605) );
  XNOR2_X1 U13482 ( .A(n13606), .B(n13607), .ZN(n13322) );
  XNOR2_X1 U13483 ( .A(n13608), .B(n13609), .ZN(n13606) );
  NOR2_X1 U13484 ( .A1(n8750), .A2(n8401), .ZN(n13609) );
  XNOR2_X1 U13485 ( .A(n13610), .B(n13611), .ZN(n13408) );
  XNOR2_X1 U13486 ( .A(n13612), .B(n13613), .ZN(n13611) );
  XOR2_X1 U13487 ( .A(n13614), .B(n13615), .Z(n13304) );
  XOR2_X1 U13488 ( .A(n13616), .B(n13617), .Z(n13614) );
  NOR2_X1 U13489 ( .A1(n8210), .A2(n8401), .ZN(n13617) );
  XNOR2_X1 U13490 ( .A(n13618), .B(n13619), .ZN(n13296) );
  NAND2_X1 U13491 ( .A1(n13620), .A2(n13621), .ZN(n13618) );
  XNOR2_X1 U13492 ( .A(n13622), .B(n13623), .ZN(n13412) );
  NAND2_X1 U13493 ( .A1(n13624), .A2(n13625), .ZN(n13622) );
  XNOR2_X1 U13494 ( .A(n13626), .B(n13627), .ZN(n13285) );
  XNOR2_X1 U13495 ( .A(n13628), .B(n13629), .ZN(n13627) );
  XNOR2_X1 U13496 ( .A(n13630), .B(n13631), .ZN(n13279) );
  XOR2_X1 U13497 ( .A(n13632), .B(n13633), .Z(n13631) );
  NAND2_X1 U13498 ( .A1(b_10_), .A2(a_13_), .ZN(n13633) );
  INV_X1 U13499 ( .A(n8688), .ZN(n13273) );
  NAND2_X1 U13500 ( .A1(b_11_), .A2(a_11_), .ZN(n8688) );
  XOR2_X1 U13501 ( .A(n13634), .B(n13635), .Z(n13416) );
  NAND2_X1 U13502 ( .A1(n13636), .A2(n13637), .ZN(n13634) );
  XOR2_X1 U13503 ( .A(n13638), .B(n13639), .Z(n13419) );
  XOR2_X1 U13504 ( .A(n13640), .B(n13641), .Z(n13638) );
  XNOR2_X1 U13505 ( .A(n13642), .B(n13643), .ZN(n13256) );
  NAND2_X1 U13506 ( .A1(n13644), .A2(n13645), .ZN(n13642) );
  XOR2_X1 U13507 ( .A(n13646), .B(n13647), .Z(n13424) );
  NAND2_X1 U13508 ( .A1(n13648), .A2(n13649), .ZN(n13646) );
  XNOR2_X1 U13509 ( .A(n13650), .B(n13651), .ZN(n13428) );
  XNOR2_X1 U13510 ( .A(n13652), .B(n13653), .ZN(n13651) );
  XNOR2_X1 U13511 ( .A(n13654), .B(n13655), .ZN(n13431) );
  XNOR2_X1 U13512 ( .A(n13656), .B(n13657), .ZN(n13654) );
  XNOR2_X1 U13513 ( .A(n13658), .B(n13659), .ZN(n13435) );
  XNOR2_X1 U13514 ( .A(n13660), .B(n13661), .ZN(n13658) );
  XNOR2_X1 U13515 ( .A(n13662), .B(n13663), .ZN(n13440) );
  XNOR2_X1 U13516 ( .A(n13664), .B(n13665), .ZN(n13663) );
  XNOR2_X1 U13517 ( .A(n13666), .B(n13667), .ZN(n13444) );
  XNOR2_X1 U13518 ( .A(n13668), .B(n13669), .ZN(n13666) );
  XNOR2_X1 U13519 ( .A(n13670), .B(n13671), .ZN(n13447) );
  XNOR2_X1 U13520 ( .A(n13672), .B(n13673), .ZN(n13671) );
  XNOR2_X1 U13521 ( .A(n13674), .B(n13675), .ZN(n13457) );
  XOR2_X1 U13522 ( .A(n13676), .B(n13677), .Z(n13675) );
  NAND2_X1 U13523 ( .A1(b_10_), .A2(a_1_), .ZN(n13677) );
  XOR2_X1 U13524 ( .A(n13678), .B(n13455), .Z(n13462) );
  XNOR2_X1 U13525 ( .A(n13679), .B(n13680), .ZN(n13455) );
  NOR2_X1 U13526 ( .A1(n9674), .A2(n8401), .ZN(n13680) );
  INV_X1 U13527 ( .A(n13454), .ZN(n13678) );
  NAND2_X1 U13528 ( .A1(n13681), .A2(n13682), .ZN(n7828) );
  NAND2_X1 U13529 ( .A1(n13683), .A2(n13684), .ZN(n13682) );
  NAND2_X1 U13530 ( .A1(n13461), .A2(n13460), .ZN(n13681) );
  NAND4_X1 U13531 ( .A1(n13461), .A2(n13683), .A3(n13684), .A4(n13460), .ZN(
        n7829) );
  NAND2_X1 U13532 ( .A1(n13685), .A2(n13686), .ZN(n13460) );
  NAND3_X1 U13533 ( .A1(a_0_), .A2(n13687), .A3(b_10_), .ZN(n13686) );
  OR2_X1 U13534 ( .A1(n13679), .A2(n13454), .ZN(n13687) );
  NAND2_X1 U13535 ( .A1(n13454), .A2(n13679), .ZN(n13685) );
  NAND2_X1 U13536 ( .A1(n13688), .A2(n13689), .ZN(n13679) );
  NAND3_X1 U13537 ( .A1(a_1_), .A2(n13690), .A3(b_10_), .ZN(n13689) );
  OR2_X1 U13538 ( .A1(n13676), .A2(n13674), .ZN(n13690) );
  NAND2_X1 U13539 ( .A1(n13674), .A2(n13676), .ZN(n13688) );
  NAND2_X1 U13540 ( .A1(n13691), .A2(n13692), .ZN(n13676) );
  NAND2_X1 U13541 ( .A1(n13673), .A2(n13693), .ZN(n13692) );
  OR2_X1 U13542 ( .A1(n13672), .A2(n13670), .ZN(n13693) );
  NOR2_X1 U13543 ( .A1(n8401), .A2(n8768), .ZN(n13673) );
  NAND2_X1 U13544 ( .A1(n13670), .A2(n13672), .ZN(n13691) );
  NAND2_X1 U13545 ( .A1(n13694), .A2(n13695), .ZN(n13672) );
  NAND2_X1 U13546 ( .A1(n13669), .A2(n13696), .ZN(n13695) );
  NAND2_X1 U13547 ( .A1(n13668), .A2(n13667), .ZN(n13696) );
  NOR2_X1 U13548 ( .A1(n8401), .A2(n8567), .ZN(n13669) );
  OR2_X1 U13549 ( .A1(n13667), .A2(n13668), .ZN(n13694) );
  AND2_X1 U13550 ( .A1(n13697), .A2(n13698), .ZN(n13668) );
  NAND2_X1 U13551 ( .A1(n13665), .A2(n13699), .ZN(n13698) );
  OR2_X1 U13552 ( .A1(n13664), .A2(n13662), .ZN(n13699) );
  NOR2_X1 U13553 ( .A1(n8401), .A2(n8766), .ZN(n13665) );
  NAND2_X1 U13554 ( .A1(n13662), .A2(n13664), .ZN(n13697) );
  NAND2_X1 U13555 ( .A1(n13700), .A2(n13701), .ZN(n13664) );
  NAND2_X1 U13556 ( .A1(n13661), .A2(n13702), .ZN(n13701) );
  NAND2_X1 U13557 ( .A1(n13660), .A2(n13659), .ZN(n13702) );
  NOR2_X1 U13558 ( .A1(n8401), .A2(n8517), .ZN(n13661) );
  OR2_X1 U13559 ( .A1(n13659), .A2(n13660), .ZN(n13700) );
  AND2_X1 U13560 ( .A1(n13703), .A2(n13704), .ZN(n13660) );
  NAND2_X1 U13561 ( .A1(n13657), .A2(n13705), .ZN(n13704) );
  NAND2_X1 U13562 ( .A1(n13656), .A2(n13655), .ZN(n13705) );
  NOR2_X1 U13563 ( .A1(n8401), .A2(n8491), .ZN(n13657) );
  OR2_X1 U13564 ( .A1(n13655), .A2(n13656), .ZN(n13703) );
  AND2_X1 U13565 ( .A1(n13706), .A2(n13707), .ZN(n13656) );
  NAND2_X1 U13566 ( .A1(n13653), .A2(n13708), .ZN(n13707) );
  OR2_X1 U13567 ( .A1(n13652), .A2(n13650), .ZN(n13708) );
  NOR2_X1 U13568 ( .A1(n8401), .A2(n8764), .ZN(n13653) );
  NAND2_X1 U13569 ( .A1(n13650), .A2(n13652), .ZN(n13706) );
  NAND2_X1 U13570 ( .A1(n13648), .A2(n13709), .ZN(n13652) );
  NAND2_X1 U13571 ( .A1(n13647), .A2(n13649), .ZN(n13709) );
  NAND2_X1 U13572 ( .A1(n13710), .A2(n13711), .ZN(n13649) );
  NAND2_X1 U13573 ( .A1(b_10_), .A2(a_8_), .ZN(n13711) );
  INV_X1 U13574 ( .A(n13712), .ZN(n13710) );
  XOR2_X1 U13575 ( .A(n13713), .B(n13714), .Z(n13647) );
  XOR2_X1 U13576 ( .A(n13715), .B(n13716), .Z(n13713) );
  NAND2_X1 U13577 ( .A1(a_8_), .A2(n13712), .ZN(n13648) );
  NAND2_X1 U13578 ( .A1(n13644), .A2(n13717), .ZN(n13712) );
  NAND2_X1 U13579 ( .A1(n13643), .A2(n13645), .ZN(n13717) );
  NAND2_X1 U13580 ( .A1(n13718), .A2(n13719), .ZN(n13645) );
  NAND2_X1 U13581 ( .A1(b_10_), .A2(a_9_), .ZN(n13719) );
  INV_X1 U13582 ( .A(n13720), .ZN(n13718) );
  XOR2_X1 U13583 ( .A(n13721), .B(n13722), .Z(n13643) );
  XOR2_X1 U13584 ( .A(n13723), .B(n13724), .Z(n13721) );
  NOR2_X1 U13585 ( .A1(n8761), .A2(n8762), .ZN(n13724) );
  NAND2_X1 U13586 ( .A1(a_9_), .A2(n13720), .ZN(n13644) );
  NAND2_X1 U13587 ( .A1(n13725), .A2(n13726), .ZN(n13720) );
  NAND2_X1 U13588 ( .A1(n13639), .A2(n13727), .ZN(n13726) );
  OR2_X1 U13589 ( .A1(n13640), .A2(n13641), .ZN(n13727) );
  XNOR2_X1 U13590 ( .A(n13728), .B(n13729), .ZN(n13639) );
  XOR2_X1 U13591 ( .A(n13730), .B(n13731), .Z(n13729) );
  NAND2_X1 U13592 ( .A1(b_9_), .A2(a_11_), .ZN(n13731) );
  NAND2_X1 U13593 ( .A1(n13641), .A2(n13640), .ZN(n13725) );
  NAND2_X1 U13594 ( .A1(n13636), .A2(n13732), .ZN(n13640) );
  NAND2_X1 U13595 ( .A1(n13635), .A2(n13637), .ZN(n13732) );
  NAND2_X1 U13596 ( .A1(n13733), .A2(n13734), .ZN(n13637) );
  NAND2_X1 U13597 ( .A1(b_10_), .A2(a_11_), .ZN(n13734) );
  INV_X1 U13598 ( .A(n13735), .ZN(n13733) );
  XNOR2_X1 U13599 ( .A(n13736), .B(n13737), .ZN(n13635) );
  XOR2_X1 U13600 ( .A(n13738), .B(n13739), .Z(n13737) );
  NAND2_X1 U13601 ( .A1(b_9_), .A2(a_12_), .ZN(n13739) );
  NAND2_X1 U13602 ( .A1(a_11_), .A2(n13735), .ZN(n13636) );
  NAND2_X1 U13603 ( .A1(n13500), .A2(n13740), .ZN(n13735) );
  NAND2_X1 U13604 ( .A1(n13499), .A2(n13501), .ZN(n13740) );
  NAND2_X1 U13605 ( .A1(n13741), .A2(n13742), .ZN(n13501) );
  NAND2_X1 U13606 ( .A1(b_10_), .A2(a_12_), .ZN(n13742) );
  INV_X1 U13607 ( .A(n13743), .ZN(n13741) );
  XNOR2_X1 U13608 ( .A(n13744), .B(n13745), .ZN(n13499) );
  XOR2_X1 U13609 ( .A(n13746), .B(n13747), .Z(n13745) );
  NAND2_X1 U13610 ( .A1(b_9_), .A2(a_13_), .ZN(n13747) );
  NAND2_X1 U13611 ( .A1(a_12_), .A2(n13743), .ZN(n13500) );
  NAND2_X1 U13612 ( .A1(n13748), .A2(n13749), .ZN(n13743) );
  NAND3_X1 U13613 ( .A1(a_13_), .A2(n13750), .A3(b_10_), .ZN(n13749) );
  OR2_X1 U13614 ( .A1(n13632), .A2(n13630), .ZN(n13750) );
  NAND2_X1 U13615 ( .A1(n13630), .A2(n13632), .ZN(n13748) );
  NAND2_X1 U13616 ( .A1(n13751), .A2(n13752), .ZN(n13632) );
  NAND2_X1 U13617 ( .A1(n13629), .A2(n13753), .ZN(n13752) );
  OR2_X1 U13618 ( .A1(n13628), .A2(n13626), .ZN(n13753) );
  NOR2_X1 U13619 ( .A1(n8401), .A2(n8757), .ZN(n13629) );
  NAND2_X1 U13620 ( .A1(n13626), .A2(n13628), .ZN(n13751) );
  NAND2_X1 U13621 ( .A1(n13624), .A2(n13754), .ZN(n13628) );
  NAND2_X1 U13622 ( .A1(n13623), .A2(n13625), .ZN(n13754) );
  NAND2_X1 U13623 ( .A1(n13755), .A2(n13756), .ZN(n13625) );
  NAND2_X1 U13624 ( .A1(b_10_), .A2(a_15_), .ZN(n13756) );
  INV_X1 U13625 ( .A(n13757), .ZN(n13755) );
  XNOR2_X1 U13626 ( .A(n13758), .B(n13759), .ZN(n13623) );
  XOR2_X1 U13627 ( .A(n13760), .B(n13761), .Z(n13759) );
  NAND2_X1 U13628 ( .A1(b_9_), .A2(a_16_), .ZN(n13761) );
  NAND2_X1 U13629 ( .A1(a_15_), .A2(n13757), .ZN(n13624) );
  NAND2_X1 U13630 ( .A1(n13620), .A2(n13762), .ZN(n13757) );
  NAND2_X1 U13631 ( .A1(n13619), .A2(n13621), .ZN(n13762) );
  NAND2_X1 U13632 ( .A1(n13763), .A2(n13764), .ZN(n13621) );
  NAND2_X1 U13633 ( .A1(b_10_), .A2(a_16_), .ZN(n13764) );
  INV_X1 U13634 ( .A(n13765), .ZN(n13763) );
  XNOR2_X1 U13635 ( .A(n13766), .B(n13767), .ZN(n13619) );
  XNOR2_X1 U13636 ( .A(n13768), .B(n13769), .ZN(n13766) );
  NOR2_X1 U13637 ( .A1(n8210), .A2(n8762), .ZN(n13769) );
  NAND2_X1 U13638 ( .A1(a_16_), .A2(n13765), .ZN(n13620) );
  NAND2_X1 U13639 ( .A1(n13770), .A2(n13771), .ZN(n13765) );
  NAND3_X1 U13640 ( .A1(a_17_), .A2(n13772), .A3(b_10_), .ZN(n13771) );
  OR2_X1 U13641 ( .A1(n13616), .A2(n13615), .ZN(n13772) );
  NAND2_X1 U13642 ( .A1(n13615), .A2(n13616), .ZN(n13770) );
  NAND2_X1 U13643 ( .A1(n13773), .A2(n13774), .ZN(n13616) );
  NAND2_X1 U13644 ( .A1(n13613), .A2(n13775), .ZN(n13774) );
  OR2_X1 U13645 ( .A1(n13612), .A2(n13610), .ZN(n13775) );
  NOR2_X1 U13646 ( .A1(n8401), .A2(n8753), .ZN(n13613) );
  NAND2_X1 U13647 ( .A1(n13610), .A2(n13612), .ZN(n13773) );
  NAND2_X1 U13648 ( .A1(n13776), .A2(n13777), .ZN(n13612) );
  NAND2_X1 U13649 ( .A1(n13527), .A2(n13778), .ZN(n13777) );
  NAND2_X1 U13650 ( .A1(n13526), .A2(n13525), .ZN(n13778) );
  NOR2_X1 U13651 ( .A1(n8401), .A2(n8170), .ZN(n13527) );
  OR2_X1 U13652 ( .A1(n13525), .A2(n13526), .ZN(n13776) );
  AND2_X1 U13653 ( .A1(n13779), .A2(n13780), .ZN(n13526) );
  NAND2_X1 U13654 ( .A1(n13535), .A2(n13781), .ZN(n13780) );
  OR2_X1 U13655 ( .A1(n13534), .A2(n13532), .ZN(n13781) );
  NOR2_X1 U13656 ( .A1(n8401), .A2(n8751), .ZN(n13535) );
  NAND2_X1 U13657 ( .A1(n13532), .A2(n13534), .ZN(n13779) );
  NAND2_X1 U13658 ( .A1(n13782), .A2(n13783), .ZN(n13534) );
  NAND3_X1 U13659 ( .A1(a_21_), .A2(n13784), .A3(b_10_), .ZN(n13783) );
  NAND2_X1 U13660 ( .A1(n13608), .A2(n13607), .ZN(n13784) );
  OR2_X1 U13661 ( .A1(n13607), .A2(n13608), .ZN(n13782) );
  AND2_X1 U13662 ( .A1(n13785), .A2(n13786), .ZN(n13608) );
  NAND3_X1 U13663 ( .A1(a_22_), .A2(n13787), .A3(b_10_), .ZN(n13786) );
  OR2_X1 U13664 ( .A1(n13604), .A2(n13602), .ZN(n13787) );
  NAND2_X1 U13665 ( .A1(n13602), .A2(n13604), .ZN(n13785) );
  NAND2_X1 U13666 ( .A1(n13788), .A2(n13789), .ZN(n13604) );
  NAND2_X1 U13667 ( .A1(n13601), .A2(n13790), .ZN(n13789) );
  OR2_X1 U13668 ( .A1(n13600), .A2(n13598), .ZN(n13790) );
  NOR2_X1 U13669 ( .A1(n8401), .A2(n8747), .ZN(n13601) );
  NAND2_X1 U13670 ( .A1(n13598), .A2(n13600), .ZN(n13788) );
  NAND2_X1 U13671 ( .A1(n13791), .A2(n13792), .ZN(n13600) );
  NAND3_X1 U13672 ( .A1(a_24_), .A2(n13793), .A3(b_10_), .ZN(n13792) );
  NAND2_X1 U13673 ( .A1(n13596), .A2(n13595), .ZN(n13793) );
  OR2_X1 U13674 ( .A1(n13595), .A2(n13596), .ZN(n13791) );
  AND2_X1 U13675 ( .A1(n13794), .A2(n13795), .ZN(n13596) );
  NAND2_X1 U13676 ( .A1(n13593), .A2(n13796), .ZN(n13795) );
  OR2_X1 U13677 ( .A1(n13592), .A2(n13591), .ZN(n13796) );
  NOR2_X1 U13678 ( .A1(n8401), .A2(n8744), .ZN(n13593) );
  NAND2_X1 U13679 ( .A1(n13591), .A2(n13592), .ZN(n13794) );
  NAND2_X1 U13680 ( .A1(n13588), .A2(n13797), .ZN(n13592) );
  NAND2_X1 U13681 ( .A1(n13587), .A2(n13589), .ZN(n13797) );
  NAND2_X1 U13682 ( .A1(n13798), .A2(n13799), .ZN(n13589) );
  NAND2_X1 U13683 ( .A1(b_10_), .A2(a_26_), .ZN(n13799) );
  INV_X1 U13684 ( .A(n13800), .ZN(n13798) );
  XNOR2_X1 U13685 ( .A(n13801), .B(n13802), .ZN(n13587) );
  NAND2_X1 U13686 ( .A1(n13803), .A2(n13804), .ZN(n13801) );
  NAND2_X1 U13687 ( .A1(a_26_), .A2(n13800), .ZN(n13588) );
  NAND2_X1 U13688 ( .A1(n13560), .A2(n13805), .ZN(n13800) );
  NAND2_X1 U13689 ( .A1(n13559), .A2(n13561), .ZN(n13805) );
  NAND2_X1 U13690 ( .A1(n13806), .A2(n13807), .ZN(n13561) );
  NAND2_X1 U13691 ( .A1(b_10_), .A2(a_27_), .ZN(n13807) );
  INV_X1 U13692 ( .A(n13808), .ZN(n13806) );
  XNOR2_X1 U13693 ( .A(n13809), .B(n13810), .ZN(n13559) );
  XOR2_X1 U13694 ( .A(n13811), .B(n13812), .Z(n13809) );
  NAND2_X1 U13695 ( .A1(b_9_), .A2(a_28_), .ZN(n13811) );
  NAND2_X1 U13696 ( .A1(a_27_), .A2(n13808), .ZN(n13560) );
  NAND2_X1 U13697 ( .A1(n13813), .A2(n13814), .ZN(n13808) );
  NAND3_X1 U13698 ( .A1(a_28_), .A2(n13815), .A3(b_10_), .ZN(n13814) );
  NAND2_X1 U13699 ( .A1(n13569), .A2(n13567), .ZN(n13815) );
  OR2_X1 U13700 ( .A1(n13567), .A2(n13569), .ZN(n13813) );
  AND2_X1 U13701 ( .A1(n13816), .A2(n13817), .ZN(n13569) );
  NAND2_X1 U13702 ( .A1(n13583), .A2(n13818), .ZN(n13817) );
  OR2_X1 U13703 ( .A1(n13584), .A2(n13585), .ZN(n13818) );
  NOR2_X1 U13704 ( .A1(n8401), .A2(n7890), .ZN(n13583) );
  NAND2_X1 U13705 ( .A1(n13585), .A2(n13584), .ZN(n13816) );
  NAND2_X1 U13706 ( .A1(n13819), .A2(n13820), .ZN(n13584) );
  NAND2_X1 U13707 ( .A1(b_8_), .A2(n13821), .ZN(n13820) );
  NAND2_X1 U13708 ( .A1(n7864), .A2(n13822), .ZN(n13821) );
  NAND2_X1 U13709 ( .A1(a_31_), .A2(n8762), .ZN(n13822) );
  NAND2_X1 U13710 ( .A1(b_9_), .A2(n13823), .ZN(n13819) );
  NAND2_X1 U13711 ( .A1(n9137), .A2(n13824), .ZN(n13823) );
  NAND2_X1 U13712 ( .A1(a_30_), .A2(n8451), .ZN(n13824) );
  AND3_X1 U13713 ( .A1(b_9_), .A2(b_10_), .A3(n7818), .ZN(n13585) );
  XNOR2_X1 U13714 ( .A(n13825), .B(n13826), .ZN(n13567) );
  XOR2_X1 U13715 ( .A(n13827), .B(n13828), .Z(n13825) );
  XNOR2_X1 U13716 ( .A(n13829), .B(n13830), .ZN(n13591) );
  NAND2_X1 U13717 ( .A1(n13831), .A2(n13832), .ZN(n13829) );
  XNOR2_X1 U13718 ( .A(n13833), .B(n13834), .ZN(n13595) );
  XOR2_X1 U13719 ( .A(n13835), .B(n13836), .Z(n13833) );
  XNOR2_X1 U13720 ( .A(n13837), .B(n13838), .ZN(n13598) );
  XNOR2_X1 U13721 ( .A(n13839), .B(n13840), .ZN(n13837) );
  NOR2_X1 U13722 ( .A1(n8745), .A2(n8762), .ZN(n13840) );
  XNOR2_X1 U13723 ( .A(n13841), .B(n13842), .ZN(n13602) );
  XNOR2_X1 U13724 ( .A(n13843), .B(n13844), .ZN(n13842) );
  XOR2_X1 U13725 ( .A(n13845), .B(n13846), .Z(n13607) );
  XNOR2_X1 U13726 ( .A(n13847), .B(n13848), .ZN(n13846) );
  XOR2_X1 U13727 ( .A(n13849), .B(n13850), .Z(n13532) );
  XNOR2_X1 U13728 ( .A(n13851), .B(n13852), .ZN(n13849) );
  NAND2_X1 U13729 ( .A1(b_9_), .A2(a_21_), .ZN(n13851) );
  XNOR2_X1 U13730 ( .A(n13853), .B(n13854), .ZN(n13525) );
  XOR2_X1 U13731 ( .A(n13855), .B(n13856), .Z(n13853) );
  NOR2_X1 U13732 ( .A1(n8751), .A2(n8762), .ZN(n13856) );
  XNOR2_X1 U13733 ( .A(n13857), .B(n13858), .ZN(n13610) );
  XOR2_X1 U13734 ( .A(n13859), .B(n13860), .Z(n13858) );
  NAND2_X1 U13735 ( .A1(b_9_), .A2(a_19_), .ZN(n13860) );
  XNOR2_X1 U13736 ( .A(n13861), .B(n13862), .ZN(n13615) );
  XNOR2_X1 U13737 ( .A(n13863), .B(n13864), .ZN(n13861) );
  NOR2_X1 U13738 ( .A1(n8753), .A2(n8762), .ZN(n13864) );
  XOR2_X1 U13739 ( .A(n13865), .B(n13866), .Z(n13626) );
  XOR2_X1 U13740 ( .A(n13867), .B(n13868), .Z(n13865) );
  NOR2_X1 U13741 ( .A1(n8276), .A2(n8762), .ZN(n13868) );
  XNOR2_X1 U13742 ( .A(n13869), .B(n13870), .ZN(n13630) );
  XOR2_X1 U13743 ( .A(n13871), .B(n13872), .Z(n13870) );
  NAND2_X1 U13744 ( .A1(b_9_), .A2(a_14_), .ZN(n13872) );
  INV_X1 U13745 ( .A(n8685), .ZN(n13641) );
  NAND2_X1 U13746 ( .A1(b_10_), .A2(a_10_), .ZN(n8685) );
  XOR2_X1 U13747 ( .A(n13873), .B(n13874), .Z(n13650) );
  XNOR2_X1 U13748 ( .A(n13875), .B(n13876), .ZN(n13873) );
  NAND2_X1 U13749 ( .A1(b_9_), .A2(a_8_), .ZN(n13875) );
  XOR2_X1 U13750 ( .A(n13877), .B(n13878), .Z(n13655) );
  XOR2_X1 U13751 ( .A(n13879), .B(n13880), .Z(n13878) );
  NAND2_X1 U13752 ( .A1(b_9_), .A2(a_7_), .ZN(n13880) );
  XNOR2_X1 U13753 ( .A(n13881), .B(n13882), .ZN(n13659) );
  XOR2_X1 U13754 ( .A(n13883), .B(n13884), .Z(n13881) );
  NOR2_X1 U13755 ( .A1(n8491), .A2(n8762), .ZN(n13884) );
  XNOR2_X1 U13756 ( .A(n13885), .B(n13886), .ZN(n13662) );
  XOR2_X1 U13757 ( .A(n13887), .B(n13888), .Z(n13886) );
  NAND2_X1 U13758 ( .A1(b_9_), .A2(a_5_), .ZN(n13888) );
  XNOR2_X1 U13759 ( .A(n13889), .B(n13890), .ZN(n13667) );
  XOR2_X1 U13760 ( .A(n13891), .B(n13892), .Z(n13889) );
  NOR2_X1 U13761 ( .A1(n8766), .A2(n8762), .ZN(n13892) );
  XOR2_X1 U13762 ( .A(n13893), .B(n13894), .Z(n13670) );
  XOR2_X1 U13763 ( .A(n13895), .B(n13896), .Z(n13893) );
  NOR2_X1 U13764 ( .A1(n8567), .A2(n8762), .ZN(n13896) );
  XOR2_X1 U13765 ( .A(n13897), .B(n13898), .Z(n13674) );
  XOR2_X1 U13766 ( .A(n13899), .B(n13900), .Z(n13897) );
  NOR2_X1 U13767 ( .A1(n8768), .A2(n8762), .ZN(n13900) );
  XOR2_X1 U13768 ( .A(n13901), .B(n13902), .Z(n13454) );
  XOR2_X1 U13769 ( .A(n13903), .B(n13904), .Z(n13901) );
  NOR2_X1 U13770 ( .A1(n8617), .A2(n8762), .ZN(n13904) );
  NAND3_X1 U13771 ( .A1(n13905), .A2(n13906), .A3(n13907), .ZN(n13683) );
  XOR2_X1 U13772 ( .A(n13908), .B(n13909), .Z(n13907) );
  XOR2_X1 U13773 ( .A(n13910), .B(n13911), .Z(n13461) );
  XOR2_X1 U13774 ( .A(n13912), .B(n13913), .Z(n13910) );
  NAND2_X1 U13775 ( .A1(n13914), .A2(n13684), .ZN(n7834) );
  OR2_X1 U13776 ( .A1(n13684), .A2(n13914), .ZN(n7835) );
  XNOR2_X1 U13777 ( .A(n13915), .B(n13916), .ZN(n13914) );
  NAND2_X1 U13778 ( .A1(n13917), .A2(n13918), .ZN(n13684) );
  NAND2_X1 U13779 ( .A1(n13905), .A2(n13906), .ZN(n13918) );
  NAND2_X1 U13780 ( .A1(n13913), .A2(n13919), .ZN(n13906) );
  OR2_X1 U13781 ( .A1(n13912), .A2(n13911), .ZN(n13919) );
  NOR2_X1 U13782 ( .A1(n8762), .A2(n9674), .ZN(n13913) );
  NAND2_X1 U13783 ( .A1(n13911), .A2(n13912), .ZN(n13905) );
  NAND2_X1 U13784 ( .A1(n13920), .A2(n13921), .ZN(n13912) );
  NAND3_X1 U13785 ( .A1(a_1_), .A2(n13922), .A3(b_9_), .ZN(n13921) );
  OR2_X1 U13786 ( .A1(n13903), .A2(n13902), .ZN(n13922) );
  NAND2_X1 U13787 ( .A1(n13902), .A2(n13903), .ZN(n13920) );
  NAND2_X1 U13788 ( .A1(n13923), .A2(n13924), .ZN(n13903) );
  NAND3_X1 U13789 ( .A1(a_2_), .A2(n13925), .A3(b_9_), .ZN(n13924) );
  OR2_X1 U13790 ( .A1(n13899), .A2(n13898), .ZN(n13925) );
  NAND2_X1 U13791 ( .A1(n13898), .A2(n13899), .ZN(n13923) );
  NAND2_X1 U13792 ( .A1(n13926), .A2(n13927), .ZN(n13899) );
  NAND3_X1 U13793 ( .A1(a_3_), .A2(n13928), .A3(b_9_), .ZN(n13927) );
  OR2_X1 U13794 ( .A1(n13895), .A2(n13894), .ZN(n13928) );
  NAND2_X1 U13795 ( .A1(n13894), .A2(n13895), .ZN(n13926) );
  NAND2_X1 U13796 ( .A1(n13929), .A2(n13930), .ZN(n13895) );
  NAND3_X1 U13797 ( .A1(a_4_), .A2(n13931), .A3(b_9_), .ZN(n13930) );
  OR2_X1 U13798 ( .A1(n13891), .A2(n13890), .ZN(n13931) );
  NAND2_X1 U13799 ( .A1(n13890), .A2(n13891), .ZN(n13929) );
  NAND2_X1 U13800 ( .A1(n13932), .A2(n13933), .ZN(n13891) );
  NAND3_X1 U13801 ( .A1(a_5_), .A2(n13934), .A3(b_9_), .ZN(n13933) );
  OR2_X1 U13802 ( .A1(n13887), .A2(n13885), .ZN(n13934) );
  NAND2_X1 U13803 ( .A1(n13885), .A2(n13887), .ZN(n13932) );
  NAND2_X1 U13804 ( .A1(n13935), .A2(n13936), .ZN(n13887) );
  NAND3_X1 U13805 ( .A1(a_6_), .A2(n13937), .A3(b_9_), .ZN(n13936) );
  OR2_X1 U13806 ( .A1(n13883), .A2(n13882), .ZN(n13937) );
  NAND2_X1 U13807 ( .A1(n13882), .A2(n13883), .ZN(n13935) );
  NAND2_X1 U13808 ( .A1(n13938), .A2(n13939), .ZN(n13883) );
  NAND3_X1 U13809 ( .A1(a_7_), .A2(n13940), .A3(b_9_), .ZN(n13939) );
  OR2_X1 U13810 ( .A1(n13879), .A2(n13877), .ZN(n13940) );
  NAND2_X1 U13811 ( .A1(n13877), .A2(n13879), .ZN(n13938) );
  NAND2_X1 U13812 ( .A1(n13941), .A2(n13942), .ZN(n13879) );
  NAND3_X1 U13813 ( .A1(a_8_), .A2(n13943), .A3(b_9_), .ZN(n13942) );
  OR2_X1 U13814 ( .A1(n13876), .A2(n13874), .ZN(n13943) );
  NAND2_X1 U13815 ( .A1(n13874), .A2(n13876), .ZN(n13941) );
  NAND2_X1 U13816 ( .A1(n13944), .A2(n13945), .ZN(n13876) );
  NAND2_X1 U13817 ( .A1(n13714), .A2(n13946), .ZN(n13945) );
  OR2_X1 U13818 ( .A1(n13715), .A2(n13716), .ZN(n13946) );
  XNOR2_X1 U13819 ( .A(n13947), .B(n13948), .ZN(n13714) );
  XNOR2_X1 U13820 ( .A(n13949), .B(n13950), .ZN(n13948) );
  NAND2_X1 U13821 ( .A1(n13716), .A2(n13715), .ZN(n13944) );
  NAND2_X1 U13822 ( .A1(n13951), .A2(n13952), .ZN(n13715) );
  NAND3_X1 U13823 ( .A1(a_10_), .A2(n13953), .A3(b_9_), .ZN(n13952) );
  OR2_X1 U13824 ( .A1(n13723), .A2(n13722), .ZN(n13953) );
  NAND2_X1 U13825 ( .A1(n13722), .A2(n13723), .ZN(n13951) );
  NAND2_X1 U13826 ( .A1(n13954), .A2(n13955), .ZN(n13723) );
  NAND3_X1 U13827 ( .A1(a_11_), .A2(n13956), .A3(b_9_), .ZN(n13955) );
  OR2_X1 U13828 ( .A1(n13730), .A2(n13728), .ZN(n13956) );
  NAND2_X1 U13829 ( .A1(n13728), .A2(n13730), .ZN(n13954) );
  NAND2_X1 U13830 ( .A1(n13957), .A2(n13958), .ZN(n13730) );
  NAND3_X1 U13831 ( .A1(a_12_), .A2(n13959), .A3(b_9_), .ZN(n13958) );
  OR2_X1 U13832 ( .A1(n13738), .A2(n13736), .ZN(n13959) );
  NAND2_X1 U13833 ( .A1(n13736), .A2(n13738), .ZN(n13957) );
  NAND2_X1 U13834 ( .A1(n13960), .A2(n13961), .ZN(n13738) );
  NAND3_X1 U13835 ( .A1(a_13_), .A2(n13962), .A3(b_9_), .ZN(n13961) );
  OR2_X1 U13836 ( .A1(n13746), .A2(n13744), .ZN(n13962) );
  NAND2_X1 U13837 ( .A1(n13744), .A2(n13746), .ZN(n13960) );
  NAND2_X1 U13838 ( .A1(n13963), .A2(n13964), .ZN(n13746) );
  NAND3_X1 U13839 ( .A1(a_14_), .A2(n13965), .A3(b_9_), .ZN(n13964) );
  OR2_X1 U13840 ( .A1(n13871), .A2(n13869), .ZN(n13965) );
  NAND2_X1 U13841 ( .A1(n13869), .A2(n13871), .ZN(n13963) );
  NAND2_X1 U13842 ( .A1(n13966), .A2(n13967), .ZN(n13871) );
  NAND3_X1 U13843 ( .A1(a_15_), .A2(n13968), .A3(b_9_), .ZN(n13967) );
  OR2_X1 U13844 ( .A1(n13867), .A2(n13866), .ZN(n13968) );
  NAND2_X1 U13845 ( .A1(n13866), .A2(n13867), .ZN(n13966) );
  NAND2_X1 U13846 ( .A1(n13969), .A2(n13970), .ZN(n13867) );
  NAND3_X1 U13847 ( .A1(a_16_), .A2(n13971), .A3(b_9_), .ZN(n13970) );
  OR2_X1 U13848 ( .A1(n13760), .A2(n13758), .ZN(n13971) );
  NAND2_X1 U13849 ( .A1(n13758), .A2(n13760), .ZN(n13969) );
  NAND2_X1 U13850 ( .A1(n13972), .A2(n13973), .ZN(n13760) );
  NAND3_X1 U13851 ( .A1(a_17_), .A2(n13974), .A3(b_9_), .ZN(n13973) );
  NAND2_X1 U13852 ( .A1(n13768), .A2(n13767), .ZN(n13974) );
  OR2_X1 U13853 ( .A1(n13767), .A2(n13768), .ZN(n13972) );
  AND2_X1 U13854 ( .A1(n13975), .A2(n13976), .ZN(n13768) );
  NAND3_X1 U13855 ( .A1(a_18_), .A2(n13977), .A3(b_9_), .ZN(n13976) );
  NAND2_X1 U13856 ( .A1(n13863), .A2(n13862), .ZN(n13977) );
  OR2_X1 U13857 ( .A1(n13862), .A2(n13863), .ZN(n13975) );
  AND2_X1 U13858 ( .A1(n13978), .A2(n13979), .ZN(n13863) );
  NAND3_X1 U13859 ( .A1(a_19_), .A2(n13980), .A3(b_9_), .ZN(n13979) );
  OR2_X1 U13860 ( .A1(n13859), .A2(n13857), .ZN(n13980) );
  NAND2_X1 U13861 ( .A1(n13857), .A2(n13859), .ZN(n13978) );
  NAND2_X1 U13862 ( .A1(n13981), .A2(n13982), .ZN(n13859) );
  NAND3_X1 U13863 ( .A1(a_20_), .A2(n13983), .A3(b_9_), .ZN(n13982) );
  OR2_X1 U13864 ( .A1(n13855), .A2(n13854), .ZN(n13983) );
  NAND2_X1 U13865 ( .A1(n13854), .A2(n13855), .ZN(n13981) );
  NAND2_X1 U13866 ( .A1(n13984), .A2(n13985), .ZN(n13855) );
  NAND3_X1 U13867 ( .A1(a_21_), .A2(n13986), .A3(b_9_), .ZN(n13985) );
  OR2_X1 U13868 ( .A1(n13852), .A2(n13850), .ZN(n13986) );
  NAND2_X1 U13869 ( .A1(n13850), .A2(n13852), .ZN(n13984) );
  NAND2_X1 U13870 ( .A1(n13987), .A2(n13988), .ZN(n13852) );
  NAND2_X1 U13871 ( .A1(n13848), .A2(n13989), .ZN(n13988) );
  OR2_X1 U13872 ( .A1(n13847), .A2(n13845), .ZN(n13989) );
  NOR2_X1 U13873 ( .A1(n8762), .A2(n8748), .ZN(n13848) );
  NAND2_X1 U13874 ( .A1(n13845), .A2(n13847), .ZN(n13987) );
  NAND2_X1 U13875 ( .A1(n13990), .A2(n13991), .ZN(n13847) );
  NAND2_X1 U13876 ( .A1(n13844), .A2(n13992), .ZN(n13991) );
  OR2_X1 U13877 ( .A1(n13843), .A2(n13841), .ZN(n13992) );
  NOR2_X1 U13878 ( .A1(n8762), .A2(n8747), .ZN(n13844) );
  NAND2_X1 U13879 ( .A1(n13841), .A2(n13843), .ZN(n13990) );
  NAND2_X1 U13880 ( .A1(n13993), .A2(n13994), .ZN(n13843) );
  NAND3_X1 U13881 ( .A1(a_24_), .A2(n13995), .A3(b_9_), .ZN(n13994) );
  NAND2_X1 U13882 ( .A1(n13839), .A2(n13838), .ZN(n13995) );
  OR2_X1 U13883 ( .A1(n13838), .A2(n13839), .ZN(n13993) );
  AND2_X1 U13884 ( .A1(n13996), .A2(n13997), .ZN(n13839) );
  NAND2_X1 U13885 ( .A1(n13836), .A2(n13998), .ZN(n13997) );
  OR2_X1 U13886 ( .A1(n13835), .A2(n13834), .ZN(n13998) );
  NOR2_X1 U13887 ( .A1(n8762), .A2(n8744), .ZN(n13836) );
  NAND2_X1 U13888 ( .A1(n13834), .A2(n13835), .ZN(n13996) );
  NAND2_X1 U13889 ( .A1(n13831), .A2(n13999), .ZN(n13835) );
  NAND2_X1 U13890 ( .A1(n13830), .A2(n13832), .ZN(n13999) );
  NAND2_X1 U13891 ( .A1(n14000), .A2(n14001), .ZN(n13832) );
  NAND2_X1 U13892 ( .A1(b_9_), .A2(a_26_), .ZN(n14001) );
  INV_X1 U13893 ( .A(n14002), .ZN(n14000) );
  XNOR2_X1 U13894 ( .A(n14003), .B(n14004), .ZN(n13830) );
  NAND2_X1 U13895 ( .A1(n14005), .A2(n14006), .ZN(n14003) );
  NAND2_X1 U13896 ( .A1(a_26_), .A2(n14002), .ZN(n13831) );
  NAND2_X1 U13897 ( .A1(n13803), .A2(n14007), .ZN(n14002) );
  NAND2_X1 U13898 ( .A1(n13802), .A2(n13804), .ZN(n14007) );
  NAND2_X1 U13899 ( .A1(n14008), .A2(n14009), .ZN(n13804) );
  NAND2_X1 U13900 ( .A1(b_9_), .A2(a_27_), .ZN(n14009) );
  INV_X1 U13901 ( .A(n14010), .ZN(n14008) );
  XNOR2_X1 U13902 ( .A(n14011), .B(n14012), .ZN(n13802) );
  XOR2_X1 U13903 ( .A(n14013), .B(n14014), .Z(n14011) );
  NAND2_X1 U13904 ( .A1(b_8_), .A2(a_28_), .ZN(n14013) );
  NAND2_X1 U13905 ( .A1(a_27_), .A2(n14010), .ZN(n13803) );
  NAND2_X1 U13906 ( .A1(n14015), .A2(n14016), .ZN(n14010) );
  NAND3_X1 U13907 ( .A1(a_28_), .A2(n14017), .A3(b_9_), .ZN(n14016) );
  NAND2_X1 U13908 ( .A1(n13812), .A2(n13810), .ZN(n14017) );
  OR2_X1 U13909 ( .A1(n13810), .A2(n13812), .ZN(n14015) );
  AND2_X1 U13910 ( .A1(n14018), .A2(n14019), .ZN(n13812) );
  NAND2_X1 U13911 ( .A1(n13826), .A2(n14020), .ZN(n14019) );
  OR2_X1 U13912 ( .A1(n13827), .A2(n13828), .ZN(n14020) );
  NOR2_X1 U13913 ( .A1(n8762), .A2(n7890), .ZN(n13826) );
  NAND2_X1 U13914 ( .A1(n13828), .A2(n13827), .ZN(n14018) );
  NAND2_X1 U13915 ( .A1(n14021), .A2(n14022), .ZN(n13827) );
  NAND2_X1 U13916 ( .A1(b_7_), .A2(n14023), .ZN(n14022) );
  NAND2_X1 U13917 ( .A1(n7864), .A2(n14024), .ZN(n14023) );
  NAND2_X1 U13918 ( .A1(a_31_), .A2(n8451), .ZN(n14024) );
  NAND2_X1 U13919 ( .A1(b_8_), .A2(n14025), .ZN(n14021) );
  NAND2_X1 U13920 ( .A1(n9137), .A2(n14026), .ZN(n14025) );
  NAND2_X1 U13921 ( .A1(a_30_), .A2(n8482), .ZN(n14026) );
  AND3_X1 U13922 ( .A1(b_8_), .A2(b_9_), .A3(n7818), .ZN(n13828) );
  XNOR2_X1 U13923 ( .A(n14027), .B(n14028), .ZN(n13810) );
  XOR2_X1 U13924 ( .A(n14029), .B(n14030), .Z(n14027) );
  XNOR2_X1 U13925 ( .A(n14031), .B(n14032), .ZN(n13834) );
  NAND2_X1 U13926 ( .A1(n14033), .A2(n14034), .ZN(n14031) );
  XNOR2_X1 U13927 ( .A(n14035), .B(n14036), .ZN(n13838) );
  XOR2_X1 U13928 ( .A(n14037), .B(n14038), .Z(n14035) );
  XNOR2_X1 U13929 ( .A(n14039), .B(n14040), .ZN(n13841) );
  XNOR2_X1 U13930 ( .A(n14041), .B(n14042), .ZN(n14039) );
  NOR2_X1 U13931 ( .A1(n8745), .A2(n8451), .ZN(n14042) );
  XNOR2_X1 U13932 ( .A(n14043), .B(n14044), .ZN(n13845) );
  XOR2_X1 U13933 ( .A(n14045), .B(n14046), .Z(n14044) );
  NAND2_X1 U13934 ( .A1(b_8_), .A2(a_23_), .ZN(n14046) );
  XNOR2_X1 U13935 ( .A(n14047), .B(n14048), .ZN(n13850) );
  XNOR2_X1 U13936 ( .A(n14049), .B(n14050), .ZN(n14048) );
  XNOR2_X1 U13937 ( .A(n14051), .B(n14052), .ZN(n13854) );
  XNOR2_X1 U13938 ( .A(n14053), .B(n14054), .ZN(n14051) );
  XNOR2_X1 U13939 ( .A(n14055), .B(n14056), .ZN(n13857) );
  XNOR2_X1 U13940 ( .A(n14057), .B(n14058), .ZN(n14055) );
  XNOR2_X1 U13941 ( .A(n14059), .B(n14060), .ZN(n13862) );
  XOR2_X1 U13942 ( .A(n14061), .B(n14062), .Z(n14059) );
  XNOR2_X1 U13943 ( .A(n14063), .B(n14064), .ZN(n13767) );
  XOR2_X1 U13944 ( .A(n14065), .B(n14066), .Z(n14063) );
  NOR2_X1 U13945 ( .A1(n8753), .A2(n8451), .ZN(n14066) );
  XNOR2_X1 U13946 ( .A(n14067), .B(n14068), .ZN(n13758) );
  NAND2_X1 U13947 ( .A1(n14069), .A2(n14070), .ZN(n14067) );
  XNOR2_X1 U13948 ( .A(n14071), .B(n14072), .ZN(n13866) );
  NAND2_X1 U13949 ( .A1(n14073), .A2(n14074), .ZN(n14071) );
  XNOR2_X1 U13950 ( .A(n14075), .B(n14076), .ZN(n13869) );
  XNOR2_X1 U13951 ( .A(n14077), .B(n14078), .ZN(n14075) );
  XNOR2_X1 U13952 ( .A(n14079), .B(n14080), .ZN(n13744) );
  XOR2_X1 U13953 ( .A(n14081), .B(n14082), .Z(n14080) );
  NAND2_X1 U13954 ( .A1(b_8_), .A2(a_14_), .ZN(n14082) );
  XNOR2_X1 U13955 ( .A(n14083), .B(n14084), .ZN(n13736) );
  XNOR2_X1 U13956 ( .A(n14085), .B(n14086), .ZN(n14083) );
  XNOR2_X1 U13957 ( .A(n14087), .B(n14088), .ZN(n13728) );
  XNOR2_X1 U13958 ( .A(n14089), .B(n14090), .ZN(n14088) );
  XNOR2_X1 U13959 ( .A(n14091), .B(n14092), .ZN(n13722) );
  XNOR2_X1 U13960 ( .A(n14093), .B(n14094), .ZN(n14091) );
  INV_X1 U13961 ( .A(n8682), .ZN(n13716) );
  NAND2_X1 U13962 ( .A1(b_9_), .A2(a_9_), .ZN(n8682) );
  XNOR2_X1 U13963 ( .A(n14095), .B(n14096), .ZN(n13874) );
  XNOR2_X1 U13964 ( .A(n14097), .B(n14098), .ZN(n14095) );
  XNOR2_X1 U13965 ( .A(n14099), .B(n14100), .ZN(n13877) );
  XNOR2_X1 U13966 ( .A(n14101), .B(n8679), .ZN(n14100) );
  XNOR2_X1 U13967 ( .A(n14102), .B(n14103), .ZN(n13882) );
  XNOR2_X1 U13968 ( .A(n14104), .B(n14105), .ZN(n14103) );
  XNOR2_X1 U13969 ( .A(n14106), .B(n14107), .ZN(n13885) );
  XNOR2_X1 U13970 ( .A(n14108), .B(n14109), .ZN(n14106) );
  XNOR2_X1 U13971 ( .A(n14110), .B(n14111), .ZN(n13890) );
  XOR2_X1 U13972 ( .A(n14112), .B(n14113), .Z(n14111) );
  NAND2_X1 U13973 ( .A1(b_8_), .A2(a_5_), .ZN(n14113) );
  XNOR2_X1 U13974 ( .A(n14114), .B(n14115), .ZN(n13894) );
  XOR2_X1 U13975 ( .A(n14116), .B(n14117), .Z(n14115) );
  NAND2_X1 U13976 ( .A1(b_8_), .A2(a_4_), .ZN(n14117) );
  XOR2_X1 U13977 ( .A(n14118), .B(n14119), .Z(n13898) );
  XOR2_X1 U13978 ( .A(n14120), .B(n14121), .Z(n14118) );
  NOR2_X1 U13979 ( .A1(n8567), .A2(n8451), .ZN(n14121) );
  XOR2_X1 U13980 ( .A(n14122), .B(n14123), .Z(n13902) );
  XNOR2_X1 U13981 ( .A(n14124), .B(n14125), .ZN(n14123) );
  NAND2_X1 U13982 ( .A1(b_8_), .A2(a_2_), .ZN(n14125) );
  XOR2_X1 U13983 ( .A(n14126), .B(n14127), .Z(n13911) );
  XNOR2_X1 U13984 ( .A(n14128), .B(n14129), .ZN(n14127) );
  NAND2_X1 U13985 ( .A1(b_8_), .A2(a_1_), .ZN(n14129) );
  XNOR2_X1 U13986 ( .A(n13909), .B(n13908), .ZN(n13917) );
  XNOR2_X1 U13987 ( .A(n14130), .B(n14131), .ZN(n13908) );
  NOR2_X1 U13988 ( .A1(n9674), .A2(n8451), .ZN(n14131) );
  NAND2_X1 U13989 ( .A1(n14132), .A2(n14133), .ZN(n7840) );
  NAND2_X1 U13990 ( .A1(n14134), .A2(n14135), .ZN(n14133) );
  NAND2_X1 U13991 ( .A1(n13916), .A2(n13915), .ZN(n14132) );
  NAND4_X1 U13992 ( .A1(n13916), .A2(n14134), .A3(n14135), .A4(n13915), .ZN(
        n7841) );
  NAND2_X1 U13993 ( .A1(n14136), .A2(n14137), .ZN(n13915) );
  NAND3_X1 U13994 ( .A1(a_0_), .A2(n14138), .A3(b_8_), .ZN(n14137) );
  OR2_X1 U13995 ( .A1(n14130), .A2(n13909), .ZN(n14138) );
  NAND2_X1 U13996 ( .A1(n13909), .A2(n14130), .ZN(n14136) );
  NAND2_X1 U13997 ( .A1(n14139), .A2(n14140), .ZN(n14130) );
  NAND3_X1 U13998 ( .A1(a_1_), .A2(n14141), .A3(b_8_), .ZN(n14140) );
  NAND2_X1 U13999 ( .A1(n14128), .A2(n14126), .ZN(n14141) );
  OR2_X1 U14000 ( .A1(n14126), .A2(n14128), .ZN(n14139) );
  AND2_X1 U14001 ( .A1(n14142), .A2(n14143), .ZN(n14128) );
  NAND3_X1 U14002 ( .A1(a_2_), .A2(n14144), .A3(b_8_), .ZN(n14143) );
  NAND2_X1 U14003 ( .A1(n14124), .A2(n14122), .ZN(n14144) );
  OR2_X1 U14004 ( .A1(n14122), .A2(n14124), .ZN(n14142) );
  AND2_X1 U14005 ( .A1(n14145), .A2(n14146), .ZN(n14124) );
  NAND3_X1 U14006 ( .A1(a_3_), .A2(n14147), .A3(b_8_), .ZN(n14146) );
  OR2_X1 U14007 ( .A1(n14120), .A2(n14119), .ZN(n14147) );
  NAND2_X1 U14008 ( .A1(n14119), .A2(n14120), .ZN(n14145) );
  NAND2_X1 U14009 ( .A1(n14148), .A2(n14149), .ZN(n14120) );
  NAND3_X1 U14010 ( .A1(a_4_), .A2(n14150), .A3(b_8_), .ZN(n14149) );
  OR2_X1 U14011 ( .A1(n14116), .A2(n14114), .ZN(n14150) );
  NAND2_X1 U14012 ( .A1(n14114), .A2(n14116), .ZN(n14148) );
  NAND2_X1 U14013 ( .A1(n14151), .A2(n14152), .ZN(n14116) );
  NAND3_X1 U14014 ( .A1(a_5_), .A2(n14153), .A3(b_8_), .ZN(n14152) );
  OR2_X1 U14015 ( .A1(n14112), .A2(n14110), .ZN(n14153) );
  NAND2_X1 U14016 ( .A1(n14110), .A2(n14112), .ZN(n14151) );
  NAND2_X1 U14017 ( .A1(n14154), .A2(n14155), .ZN(n14112) );
  NAND2_X1 U14018 ( .A1(n14109), .A2(n14156), .ZN(n14155) );
  NAND2_X1 U14019 ( .A1(n14108), .A2(n14107), .ZN(n14156) );
  NOR2_X1 U14020 ( .A1(n8451), .A2(n8491), .ZN(n14109) );
  OR2_X1 U14021 ( .A1(n14107), .A2(n14108), .ZN(n14154) );
  AND2_X1 U14022 ( .A1(n14157), .A2(n14158), .ZN(n14108) );
  NAND2_X1 U14023 ( .A1(n14105), .A2(n14159), .ZN(n14158) );
  OR2_X1 U14024 ( .A1(n14104), .A2(n14102), .ZN(n14159) );
  NOR2_X1 U14025 ( .A1(n8451), .A2(n8764), .ZN(n14105) );
  NAND2_X1 U14026 ( .A1(n14102), .A2(n14104), .ZN(n14157) );
  NAND2_X1 U14027 ( .A1(n14160), .A2(n14161), .ZN(n14104) );
  NAND2_X1 U14028 ( .A1(n8679), .A2(n14162), .ZN(n14161) );
  OR2_X1 U14029 ( .A1(n14101), .A2(n14099), .ZN(n14162) );
  NOR2_X1 U14030 ( .A1(n8451), .A2(n8763), .ZN(n8679) );
  NAND2_X1 U14031 ( .A1(n14099), .A2(n14101), .ZN(n14160) );
  NAND2_X1 U14032 ( .A1(n14163), .A2(n14164), .ZN(n14101) );
  NAND2_X1 U14033 ( .A1(n14098), .A2(n14165), .ZN(n14164) );
  NAND2_X1 U14034 ( .A1(n14097), .A2(n14096), .ZN(n14165) );
  NOR2_X1 U14035 ( .A1(n8451), .A2(n8426), .ZN(n14098) );
  OR2_X1 U14036 ( .A1(n14096), .A2(n14097), .ZN(n14163) );
  AND2_X1 U14037 ( .A1(n14166), .A2(n14167), .ZN(n14097) );
  NAND2_X1 U14038 ( .A1(n13950), .A2(n14168), .ZN(n14167) );
  OR2_X1 U14039 ( .A1(n13949), .A2(n13947), .ZN(n14168) );
  NOR2_X1 U14040 ( .A1(n8451), .A2(n8761), .ZN(n13950) );
  NAND2_X1 U14041 ( .A1(n13947), .A2(n13949), .ZN(n14166) );
  NAND2_X1 U14042 ( .A1(n14169), .A2(n14170), .ZN(n13949) );
  NAND2_X1 U14043 ( .A1(n14094), .A2(n14171), .ZN(n14170) );
  NAND2_X1 U14044 ( .A1(n14093), .A2(n14092), .ZN(n14171) );
  NOR2_X1 U14045 ( .A1(n8451), .A2(n8376), .ZN(n14094) );
  OR2_X1 U14046 ( .A1(n14092), .A2(n14093), .ZN(n14169) );
  AND2_X1 U14047 ( .A1(n14172), .A2(n14173), .ZN(n14093) );
  NAND2_X1 U14048 ( .A1(n14090), .A2(n14174), .ZN(n14173) );
  OR2_X1 U14049 ( .A1(n14087), .A2(n14089), .ZN(n14174) );
  NOR2_X1 U14050 ( .A1(n8451), .A2(n8759), .ZN(n14090) );
  NAND2_X1 U14051 ( .A1(n14087), .A2(n14089), .ZN(n14172) );
  NAND2_X1 U14052 ( .A1(n14175), .A2(n14176), .ZN(n14089) );
  NAND2_X1 U14053 ( .A1(n14086), .A2(n14177), .ZN(n14176) );
  NAND2_X1 U14054 ( .A1(n14085), .A2(n14084), .ZN(n14177) );
  NOR2_X1 U14055 ( .A1(n8451), .A2(n8310), .ZN(n14086) );
  OR2_X1 U14056 ( .A1(n14084), .A2(n14085), .ZN(n14175) );
  AND2_X1 U14057 ( .A1(n14178), .A2(n14179), .ZN(n14085) );
  NAND3_X1 U14058 ( .A1(a_14_), .A2(n14180), .A3(b_8_), .ZN(n14179) );
  OR2_X1 U14059 ( .A1(n14079), .A2(n14081), .ZN(n14180) );
  NAND2_X1 U14060 ( .A1(n14079), .A2(n14081), .ZN(n14178) );
  NAND2_X1 U14061 ( .A1(n14181), .A2(n14182), .ZN(n14081) );
  NAND2_X1 U14062 ( .A1(n14078), .A2(n14183), .ZN(n14182) );
  NAND2_X1 U14063 ( .A1(n14077), .A2(n14076), .ZN(n14183) );
  NOR2_X1 U14064 ( .A1(n8451), .A2(n8276), .ZN(n14078) );
  OR2_X1 U14065 ( .A1(n14076), .A2(n14077), .ZN(n14181) );
  AND2_X1 U14066 ( .A1(n14073), .A2(n14184), .ZN(n14077) );
  NAND2_X1 U14067 ( .A1(n14072), .A2(n14074), .ZN(n14184) );
  NAND2_X1 U14068 ( .A1(n14185), .A2(n14186), .ZN(n14074) );
  NAND2_X1 U14069 ( .A1(b_8_), .A2(a_16_), .ZN(n14186) );
  INV_X1 U14070 ( .A(n14187), .ZN(n14185) );
  XNOR2_X1 U14071 ( .A(n14188), .B(n14189), .ZN(n14072) );
  XNOR2_X1 U14072 ( .A(n14190), .B(n14191), .ZN(n14188) );
  NOR2_X1 U14073 ( .A1(n8210), .A2(n8482), .ZN(n14191) );
  NAND2_X1 U14074 ( .A1(a_16_), .A2(n14187), .ZN(n14073) );
  NAND2_X1 U14075 ( .A1(n14069), .A2(n14192), .ZN(n14187) );
  NAND2_X1 U14076 ( .A1(n14068), .A2(n14070), .ZN(n14192) );
  NAND2_X1 U14077 ( .A1(n14193), .A2(n14194), .ZN(n14070) );
  NAND2_X1 U14078 ( .A1(b_8_), .A2(a_17_), .ZN(n14194) );
  INV_X1 U14079 ( .A(n14195), .ZN(n14193) );
  XNOR2_X1 U14080 ( .A(n14196), .B(n14197), .ZN(n14068) );
  XOR2_X1 U14081 ( .A(n14198), .B(n14199), .Z(n14197) );
  NAND2_X1 U14082 ( .A1(b_7_), .A2(a_18_), .ZN(n14199) );
  NAND2_X1 U14083 ( .A1(a_17_), .A2(n14195), .ZN(n14069) );
  NAND2_X1 U14084 ( .A1(n14200), .A2(n14201), .ZN(n14195) );
  NAND3_X1 U14085 ( .A1(a_18_), .A2(n14202), .A3(b_8_), .ZN(n14201) );
  OR2_X1 U14086 ( .A1(n14064), .A2(n14065), .ZN(n14202) );
  NAND2_X1 U14087 ( .A1(n14064), .A2(n14065), .ZN(n14200) );
  NAND2_X1 U14088 ( .A1(n14203), .A2(n14204), .ZN(n14065) );
  NAND2_X1 U14089 ( .A1(n14062), .A2(n14205), .ZN(n14204) );
  OR2_X1 U14090 ( .A1(n14060), .A2(n14061), .ZN(n14205) );
  NOR2_X1 U14091 ( .A1(n8451), .A2(n8170), .ZN(n14062) );
  NAND2_X1 U14092 ( .A1(n14060), .A2(n14061), .ZN(n14203) );
  NAND2_X1 U14093 ( .A1(n14206), .A2(n14207), .ZN(n14061) );
  NAND2_X1 U14094 ( .A1(n14058), .A2(n14208), .ZN(n14207) );
  NAND2_X1 U14095 ( .A1(n14057), .A2(n14056), .ZN(n14208) );
  NOR2_X1 U14096 ( .A1(n8451), .A2(n8751), .ZN(n14058) );
  OR2_X1 U14097 ( .A1(n14056), .A2(n14057), .ZN(n14206) );
  AND2_X1 U14098 ( .A1(n14209), .A2(n14210), .ZN(n14057) );
  NAND2_X1 U14099 ( .A1(n14054), .A2(n14211), .ZN(n14210) );
  NAND2_X1 U14100 ( .A1(n14053), .A2(n14052), .ZN(n14211) );
  NOR2_X1 U14101 ( .A1(n8451), .A2(n8750), .ZN(n14054) );
  OR2_X1 U14102 ( .A1(n14052), .A2(n14053), .ZN(n14209) );
  AND2_X1 U14103 ( .A1(n14212), .A2(n14213), .ZN(n14053) );
  NAND2_X1 U14104 ( .A1(n14050), .A2(n14214), .ZN(n14213) );
  OR2_X1 U14105 ( .A1(n14049), .A2(n14047), .ZN(n14214) );
  NOR2_X1 U14106 ( .A1(n8451), .A2(n8748), .ZN(n14050) );
  NAND2_X1 U14107 ( .A1(n14047), .A2(n14049), .ZN(n14212) );
  NAND2_X1 U14108 ( .A1(n14215), .A2(n14216), .ZN(n14049) );
  NAND3_X1 U14109 ( .A1(a_23_), .A2(n14217), .A3(b_8_), .ZN(n14216) );
  OR2_X1 U14110 ( .A1(n14045), .A2(n14043), .ZN(n14217) );
  NAND2_X1 U14111 ( .A1(n14043), .A2(n14045), .ZN(n14215) );
  NAND2_X1 U14112 ( .A1(n14218), .A2(n14219), .ZN(n14045) );
  NAND3_X1 U14113 ( .A1(a_24_), .A2(n14220), .A3(b_8_), .ZN(n14219) );
  NAND2_X1 U14114 ( .A1(n14041), .A2(n14040), .ZN(n14220) );
  OR2_X1 U14115 ( .A1(n14040), .A2(n14041), .ZN(n14218) );
  AND2_X1 U14116 ( .A1(n14221), .A2(n14222), .ZN(n14041) );
  NAND2_X1 U14117 ( .A1(n14038), .A2(n14223), .ZN(n14222) );
  OR2_X1 U14118 ( .A1(n14036), .A2(n14037), .ZN(n14223) );
  NOR2_X1 U14119 ( .A1(n8451), .A2(n8744), .ZN(n14038) );
  NAND2_X1 U14120 ( .A1(n14036), .A2(n14037), .ZN(n14221) );
  NAND2_X1 U14121 ( .A1(n14033), .A2(n14224), .ZN(n14037) );
  NAND2_X1 U14122 ( .A1(n14032), .A2(n14034), .ZN(n14224) );
  NAND2_X1 U14123 ( .A1(n14225), .A2(n14226), .ZN(n14034) );
  NAND2_X1 U14124 ( .A1(b_8_), .A2(a_26_), .ZN(n14226) );
  INV_X1 U14125 ( .A(n14227), .ZN(n14225) );
  XNOR2_X1 U14126 ( .A(n14228), .B(n14229), .ZN(n14032) );
  NAND2_X1 U14127 ( .A1(n14230), .A2(n14231), .ZN(n14228) );
  NAND2_X1 U14128 ( .A1(a_26_), .A2(n14227), .ZN(n14033) );
  NAND2_X1 U14129 ( .A1(n14005), .A2(n14232), .ZN(n14227) );
  NAND2_X1 U14130 ( .A1(n14004), .A2(n14006), .ZN(n14232) );
  NAND2_X1 U14131 ( .A1(n14233), .A2(n14234), .ZN(n14006) );
  NAND2_X1 U14132 ( .A1(b_8_), .A2(a_27_), .ZN(n14234) );
  INV_X1 U14133 ( .A(n14235), .ZN(n14233) );
  XNOR2_X1 U14134 ( .A(n14236), .B(n14237), .ZN(n14004) );
  XOR2_X1 U14135 ( .A(n14238), .B(n14239), .Z(n14236) );
  NAND2_X1 U14136 ( .A1(b_7_), .A2(a_28_), .ZN(n14238) );
  NAND2_X1 U14137 ( .A1(a_27_), .A2(n14235), .ZN(n14005) );
  NAND2_X1 U14138 ( .A1(n14240), .A2(n14241), .ZN(n14235) );
  NAND3_X1 U14139 ( .A1(a_28_), .A2(n14242), .A3(b_8_), .ZN(n14241) );
  NAND2_X1 U14140 ( .A1(n14014), .A2(n14012), .ZN(n14242) );
  OR2_X1 U14141 ( .A1(n14012), .A2(n14014), .ZN(n14240) );
  AND2_X1 U14142 ( .A1(n14243), .A2(n14244), .ZN(n14014) );
  NAND2_X1 U14143 ( .A1(n14028), .A2(n14245), .ZN(n14244) );
  OR2_X1 U14144 ( .A1(n14029), .A2(n14030), .ZN(n14245) );
  NOR2_X1 U14145 ( .A1(n8451), .A2(n7890), .ZN(n14028) );
  NAND2_X1 U14146 ( .A1(n14030), .A2(n14029), .ZN(n14243) );
  NAND2_X1 U14147 ( .A1(n14246), .A2(n14247), .ZN(n14029) );
  NAND2_X1 U14148 ( .A1(b_6_), .A2(n14248), .ZN(n14247) );
  NAND2_X1 U14149 ( .A1(n7864), .A2(n14249), .ZN(n14248) );
  NAND2_X1 U14150 ( .A1(a_31_), .A2(n8482), .ZN(n14249) );
  NAND2_X1 U14151 ( .A1(b_7_), .A2(n14250), .ZN(n14246) );
  NAND2_X1 U14152 ( .A1(n9137), .A2(n14251), .ZN(n14250) );
  NAND2_X1 U14153 ( .A1(a_30_), .A2(n8508), .ZN(n14251) );
  AND3_X1 U14154 ( .A1(b_7_), .A2(b_8_), .A3(n7818), .ZN(n14030) );
  XNOR2_X1 U14155 ( .A(n14252), .B(n14253), .ZN(n14012) );
  XOR2_X1 U14156 ( .A(n14254), .B(n14255), .Z(n14252) );
  XNOR2_X1 U14157 ( .A(n14256), .B(n14257), .ZN(n14036) );
  NAND2_X1 U14158 ( .A1(n14258), .A2(n14259), .ZN(n14256) );
  XNOR2_X1 U14159 ( .A(n14260), .B(n14261), .ZN(n14040) );
  XOR2_X1 U14160 ( .A(n14262), .B(n14263), .Z(n14260) );
  XOR2_X1 U14161 ( .A(n14264), .B(n14265), .Z(n14043) );
  XOR2_X1 U14162 ( .A(n14266), .B(n14267), .Z(n14264) );
  XOR2_X1 U14163 ( .A(n14268), .B(n14269), .Z(n14047) );
  XOR2_X1 U14164 ( .A(n14270), .B(n14271), .Z(n14268) );
  NOR2_X1 U14165 ( .A1(n8747), .A2(n8482), .ZN(n14271) );
  XOR2_X1 U14166 ( .A(n14272), .B(n14273), .Z(n14052) );
  NAND2_X1 U14167 ( .A1(n14274), .A2(n14275), .ZN(n14272) );
  XNOR2_X1 U14168 ( .A(n14276), .B(n14277), .ZN(n14056) );
  XOR2_X1 U14169 ( .A(n14278), .B(n14279), .Z(n14276) );
  NOR2_X1 U14170 ( .A1(n8750), .A2(n8482), .ZN(n14279) );
  XNOR2_X1 U14171 ( .A(n14280), .B(n14281), .ZN(n14060) );
  XNOR2_X1 U14172 ( .A(n14282), .B(n14283), .ZN(n14280) );
  NOR2_X1 U14173 ( .A1(n8751), .A2(n8482), .ZN(n14283) );
  XNOR2_X1 U14174 ( .A(n14284), .B(n14285), .ZN(n14064) );
  XNOR2_X1 U14175 ( .A(n14286), .B(n14287), .ZN(n14284) );
  NOR2_X1 U14176 ( .A1(n8170), .A2(n8482), .ZN(n14287) );
  XNOR2_X1 U14177 ( .A(n14288), .B(n14289), .ZN(n14076) );
  XOR2_X1 U14178 ( .A(n14290), .B(n14291), .Z(n14288) );
  NOR2_X1 U14179 ( .A1(n8755), .A2(n8482), .ZN(n14291) );
  XNOR2_X1 U14180 ( .A(n14292), .B(n14293), .ZN(n14079) );
  XOR2_X1 U14181 ( .A(n14294), .B(n14295), .Z(n14293) );
  NAND2_X1 U14182 ( .A1(b_7_), .A2(a_15_), .ZN(n14295) );
  XNOR2_X1 U14183 ( .A(n14296), .B(n14297), .ZN(n14084) );
  XOR2_X1 U14184 ( .A(n14298), .B(n14299), .Z(n14296) );
  NOR2_X1 U14185 ( .A1(n8757), .A2(n8482), .ZN(n14299) );
  XNOR2_X1 U14186 ( .A(n14300), .B(n14301), .ZN(n14087) );
  XOR2_X1 U14187 ( .A(n14302), .B(n14303), .Z(n14301) );
  NAND2_X1 U14188 ( .A1(b_7_), .A2(a_13_), .ZN(n14303) );
  XNOR2_X1 U14189 ( .A(n14304), .B(n14305), .ZN(n14092) );
  XOR2_X1 U14190 ( .A(n14306), .B(n14307), .Z(n14304) );
  NOR2_X1 U14191 ( .A1(n8759), .A2(n8482), .ZN(n14307) );
  XOR2_X1 U14192 ( .A(n14308), .B(n14309), .Z(n13947) );
  XOR2_X1 U14193 ( .A(n14310), .B(n14311), .Z(n14308) );
  NOR2_X1 U14194 ( .A1(n8376), .A2(n8482), .ZN(n14311) );
  XNOR2_X1 U14195 ( .A(n14312), .B(n14313), .ZN(n14096) );
  XOR2_X1 U14196 ( .A(n14314), .B(n14315), .Z(n14312) );
  NOR2_X1 U14197 ( .A1(n8761), .A2(n8482), .ZN(n14315) );
  XOR2_X1 U14198 ( .A(n14316), .B(n14317), .Z(n14099) );
  XOR2_X1 U14199 ( .A(n14318), .B(n14319), .Z(n14316) );
  NOR2_X1 U14200 ( .A1(n8426), .A2(n8482), .ZN(n14319) );
  XOR2_X1 U14201 ( .A(n14320), .B(n14321), .Z(n14102) );
  XOR2_X1 U14202 ( .A(n14322), .B(n14323), .Z(n14320) );
  NOR2_X1 U14203 ( .A1(n8763), .A2(n8482), .ZN(n14323) );
  XNOR2_X1 U14204 ( .A(n14324), .B(n14325), .ZN(n14107) );
  XOR2_X1 U14205 ( .A(n14326), .B(n14327), .Z(n14324) );
  XOR2_X1 U14206 ( .A(n14328), .B(n14329), .Z(n14110) );
  XOR2_X1 U14207 ( .A(n14330), .B(n14331), .Z(n14328) );
  NOR2_X1 U14208 ( .A1(n8491), .A2(n8482), .ZN(n14331) );
  XOR2_X1 U14209 ( .A(n14332), .B(n14333), .Z(n14114) );
  XOR2_X1 U14210 ( .A(n14334), .B(n14335), .Z(n14332) );
  NOR2_X1 U14211 ( .A1(n8517), .A2(n8482), .ZN(n14335) );
  XOR2_X1 U14212 ( .A(n14336), .B(n14337), .Z(n14119) );
  XOR2_X1 U14213 ( .A(n14338), .B(n14339), .Z(n14336) );
  NOR2_X1 U14214 ( .A1(n8766), .A2(n8482), .ZN(n14339) );
  XNOR2_X1 U14215 ( .A(n14340), .B(n14341), .ZN(n14122) );
  XOR2_X1 U14216 ( .A(n14342), .B(n14343), .Z(n14340) );
  NOR2_X1 U14217 ( .A1(n8567), .A2(n8482), .ZN(n14343) );
  XNOR2_X1 U14218 ( .A(n14344), .B(n14345), .ZN(n14126) );
  XOR2_X1 U14219 ( .A(n14346), .B(n14347), .Z(n14344) );
  NOR2_X1 U14220 ( .A1(n8768), .A2(n8482), .ZN(n14347) );
  XOR2_X1 U14221 ( .A(n14348), .B(n14349), .Z(n13909) );
  XOR2_X1 U14222 ( .A(n14350), .B(n14351), .Z(n14348) );
  NOR2_X1 U14223 ( .A1(n8617), .A2(n8482), .ZN(n14351) );
  NAND3_X1 U14224 ( .A1(n14352), .A2(n14353), .A3(n14354), .ZN(n14134) );
  XOR2_X1 U14225 ( .A(n14355), .B(n14356), .Z(n14354) );
  XOR2_X1 U14226 ( .A(n14357), .B(n14358), .Z(n13916) );
  XOR2_X1 U14227 ( .A(n14359), .B(n14360), .Z(n14357) );
  NAND2_X1 U14228 ( .A1(n14361), .A2(n14135), .ZN(n7846) );
  OR2_X1 U14229 ( .A1(n14135), .A2(n14361), .ZN(n7847) );
  XNOR2_X1 U14230 ( .A(n14362), .B(n14363), .ZN(n14361) );
  NAND2_X1 U14231 ( .A1(n14364), .A2(n14365), .ZN(n14135) );
  NAND2_X1 U14232 ( .A1(n14352), .A2(n14353), .ZN(n14365) );
  NAND2_X1 U14233 ( .A1(n14360), .A2(n14366), .ZN(n14353) );
  OR2_X1 U14234 ( .A1(n14358), .A2(n14359), .ZN(n14366) );
  NOR2_X1 U14235 ( .A1(n8482), .A2(n9674), .ZN(n14360) );
  NAND2_X1 U14236 ( .A1(n14358), .A2(n14359), .ZN(n14352) );
  NAND2_X1 U14237 ( .A1(n14367), .A2(n14368), .ZN(n14359) );
  NAND3_X1 U14238 ( .A1(a_1_), .A2(n14369), .A3(b_7_), .ZN(n14368) );
  OR2_X1 U14239 ( .A1(n14349), .A2(n14350), .ZN(n14369) );
  NAND2_X1 U14240 ( .A1(n14349), .A2(n14350), .ZN(n14367) );
  NAND2_X1 U14241 ( .A1(n14370), .A2(n14371), .ZN(n14350) );
  NAND3_X1 U14242 ( .A1(a_2_), .A2(n14372), .A3(b_7_), .ZN(n14371) );
  OR2_X1 U14243 ( .A1(n14345), .A2(n14346), .ZN(n14372) );
  NAND2_X1 U14244 ( .A1(n14345), .A2(n14346), .ZN(n14370) );
  NAND2_X1 U14245 ( .A1(n14373), .A2(n14374), .ZN(n14346) );
  NAND3_X1 U14246 ( .A1(a_3_), .A2(n14375), .A3(b_7_), .ZN(n14374) );
  OR2_X1 U14247 ( .A1(n14341), .A2(n14342), .ZN(n14375) );
  NAND2_X1 U14248 ( .A1(n14341), .A2(n14342), .ZN(n14373) );
  NAND2_X1 U14249 ( .A1(n14376), .A2(n14377), .ZN(n14342) );
  NAND3_X1 U14250 ( .A1(a_4_), .A2(n14378), .A3(b_7_), .ZN(n14377) );
  OR2_X1 U14251 ( .A1(n14337), .A2(n14338), .ZN(n14378) );
  NAND2_X1 U14252 ( .A1(n14337), .A2(n14338), .ZN(n14376) );
  NAND2_X1 U14253 ( .A1(n14379), .A2(n14380), .ZN(n14338) );
  NAND3_X1 U14254 ( .A1(a_5_), .A2(n14381), .A3(b_7_), .ZN(n14380) );
  OR2_X1 U14255 ( .A1(n14333), .A2(n14334), .ZN(n14381) );
  NAND2_X1 U14256 ( .A1(n14333), .A2(n14334), .ZN(n14379) );
  NAND2_X1 U14257 ( .A1(n14382), .A2(n14383), .ZN(n14334) );
  NAND3_X1 U14258 ( .A1(a_6_), .A2(n14384), .A3(b_7_), .ZN(n14383) );
  OR2_X1 U14259 ( .A1(n14329), .A2(n14330), .ZN(n14384) );
  NAND2_X1 U14260 ( .A1(n14329), .A2(n14330), .ZN(n14382) );
  NAND2_X1 U14261 ( .A1(n14385), .A2(n14386), .ZN(n14330) );
  NAND2_X1 U14262 ( .A1(n14325), .A2(n14387), .ZN(n14386) );
  OR2_X1 U14263 ( .A1(n14326), .A2(n14327), .ZN(n14387) );
  XNOR2_X1 U14264 ( .A(n14388), .B(n14389), .ZN(n14325) );
  XOR2_X1 U14265 ( .A(n14390), .B(n14391), .Z(n14389) );
  NAND2_X1 U14266 ( .A1(b_6_), .A2(a_8_), .ZN(n14391) );
  NAND2_X1 U14267 ( .A1(n14327), .A2(n14326), .ZN(n14385) );
  NAND2_X1 U14268 ( .A1(n14392), .A2(n14393), .ZN(n14326) );
  NAND3_X1 U14269 ( .A1(a_8_), .A2(n14394), .A3(b_7_), .ZN(n14393) );
  OR2_X1 U14270 ( .A1(n14321), .A2(n14322), .ZN(n14394) );
  NAND2_X1 U14271 ( .A1(n14321), .A2(n14322), .ZN(n14392) );
  NAND2_X1 U14272 ( .A1(n14395), .A2(n14396), .ZN(n14322) );
  NAND3_X1 U14273 ( .A1(a_9_), .A2(n14397), .A3(b_7_), .ZN(n14396) );
  OR2_X1 U14274 ( .A1(n14317), .A2(n14318), .ZN(n14397) );
  NAND2_X1 U14275 ( .A1(n14317), .A2(n14318), .ZN(n14395) );
  NAND2_X1 U14276 ( .A1(n14398), .A2(n14399), .ZN(n14318) );
  NAND3_X1 U14277 ( .A1(a_10_), .A2(n14400), .A3(b_7_), .ZN(n14399) );
  OR2_X1 U14278 ( .A1(n14313), .A2(n14314), .ZN(n14400) );
  NAND2_X1 U14279 ( .A1(n14313), .A2(n14314), .ZN(n14398) );
  NAND2_X1 U14280 ( .A1(n14401), .A2(n14402), .ZN(n14314) );
  NAND3_X1 U14281 ( .A1(a_11_), .A2(n14403), .A3(b_7_), .ZN(n14402) );
  OR2_X1 U14282 ( .A1(n14309), .A2(n14310), .ZN(n14403) );
  NAND2_X1 U14283 ( .A1(n14309), .A2(n14310), .ZN(n14401) );
  NAND2_X1 U14284 ( .A1(n14404), .A2(n14405), .ZN(n14310) );
  NAND3_X1 U14285 ( .A1(a_12_), .A2(n14406), .A3(b_7_), .ZN(n14405) );
  OR2_X1 U14286 ( .A1(n14305), .A2(n14306), .ZN(n14406) );
  NAND2_X1 U14287 ( .A1(n14305), .A2(n14306), .ZN(n14404) );
  NAND2_X1 U14288 ( .A1(n14407), .A2(n14408), .ZN(n14306) );
  NAND3_X1 U14289 ( .A1(a_13_), .A2(n14409), .A3(b_7_), .ZN(n14408) );
  OR2_X1 U14290 ( .A1(n14302), .A2(n14300), .ZN(n14409) );
  NAND2_X1 U14291 ( .A1(n14300), .A2(n14302), .ZN(n14407) );
  NAND2_X1 U14292 ( .A1(n14410), .A2(n14411), .ZN(n14302) );
  NAND3_X1 U14293 ( .A1(a_14_), .A2(n14412), .A3(b_7_), .ZN(n14411) );
  OR2_X1 U14294 ( .A1(n14297), .A2(n14298), .ZN(n14412) );
  NAND2_X1 U14295 ( .A1(n14297), .A2(n14298), .ZN(n14410) );
  NAND2_X1 U14296 ( .A1(n14413), .A2(n14414), .ZN(n14298) );
  NAND3_X1 U14297 ( .A1(a_15_), .A2(n14415), .A3(b_7_), .ZN(n14414) );
  OR2_X1 U14298 ( .A1(n14294), .A2(n14292), .ZN(n14415) );
  NAND2_X1 U14299 ( .A1(n14292), .A2(n14294), .ZN(n14413) );
  NAND2_X1 U14300 ( .A1(n14416), .A2(n14417), .ZN(n14294) );
  NAND3_X1 U14301 ( .A1(a_16_), .A2(n14418), .A3(b_7_), .ZN(n14417) );
  OR2_X1 U14302 ( .A1(n14289), .A2(n14290), .ZN(n14418) );
  NAND2_X1 U14303 ( .A1(n14289), .A2(n14290), .ZN(n14416) );
  NAND2_X1 U14304 ( .A1(n14419), .A2(n14420), .ZN(n14290) );
  NAND3_X1 U14305 ( .A1(a_17_), .A2(n14421), .A3(b_7_), .ZN(n14420) );
  NAND2_X1 U14306 ( .A1(n14190), .A2(n14189), .ZN(n14421) );
  OR2_X1 U14307 ( .A1(n14189), .A2(n14190), .ZN(n14419) );
  AND2_X1 U14308 ( .A1(n14422), .A2(n14423), .ZN(n14190) );
  NAND3_X1 U14309 ( .A1(a_18_), .A2(n14424), .A3(b_7_), .ZN(n14423) );
  OR2_X1 U14310 ( .A1(n14196), .A2(n14198), .ZN(n14424) );
  NAND2_X1 U14311 ( .A1(n14196), .A2(n14198), .ZN(n14422) );
  NAND2_X1 U14312 ( .A1(n14425), .A2(n14426), .ZN(n14198) );
  NAND3_X1 U14313 ( .A1(a_19_), .A2(n14427), .A3(b_7_), .ZN(n14426) );
  NAND2_X1 U14314 ( .A1(n14286), .A2(n14285), .ZN(n14427) );
  OR2_X1 U14315 ( .A1(n14285), .A2(n14286), .ZN(n14425) );
  AND2_X1 U14316 ( .A1(n14428), .A2(n14429), .ZN(n14286) );
  NAND3_X1 U14317 ( .A1(a_20_), .A2(n14430), .A3(b_7_), .ZN(n14429) );
  NAND2_X1 U14318 ( .A1(n14282), .A2(n14281), .ZN(n14430) );
  OR2_X1 U14319 ( .A1(n14281), .A2(n14282), .ZN(n14428) );
  AND2_X1 U14320 ( .A1(n14431), .A2(n14432), .ZN(n14282) );
  NAND3_X1 U14321 ( .A1(a_21_), .A2(n14433), .A3(b_7_), .ZN(n14432) );
  OR2_X1 U14322 ( .A1(n14277), .A2(n14278), .ZN(n14433) );
  NAND2_X1 U14323 ( .A1(n14277), .A2(n14278), .ZN(n14431) );
  NAND2_X1 U14324 ( .A1(n14274), .A2(n14434), .ZN(n14278) );
  NAND2_X1 U14325 ( .A1(n14273), .A2(n14275), .ZN(n14434) );
  NAND2_X1 U14326 ( .A1(n14435), .A2(n14436), .ZN(n14275) );
  NAND2_X1 U14327 ( .A1(b_7_), .A2(a_22_), .ZN(n14436) );
  INV_X1 U14328 ( .A(n14437), .ZN(n14435) );
  XOR2_X1 U14329 ( .A(n14438), .B(n14439), .Z(n14273) );
  XOR2_X1 U14330 ( .A(n14440), .B(n14441), .Z(n14438) );
  NOR2_X1 U14331 ( .A1(n8747), .A2(n8508), .ZN(n14441) );
  NAND2_X1 U14332 ( .A1(a_22_), .A2(n14437), .ZN(n14274) );
  NAND2_X1 U14333 ( .A1(n14442), .A2(n14443), .ZN(n14437) );
  NAND3_X1 U14334 ( .A1(a_23_), .A2(n14444), .A3(b_7_), .ZN(n14443) );
  OR2_X1 U14335 ( .A1(n14269), .A2(n14270), .ZN(n14444) );
  NAND2_X1 U14336 ( .A1(n14269), .A2(n14270), .ZN(n14442) );
  NAND2_X1 U14337 ( .A1(n14445), .A2(n14446), .ZN(n14270) );
  NAND2_X1 U14338 ( .A1(n14267), .A2(n14447), .ZN(n14446) );
  OR2_X1 U14339 ( .A1(n14265), .A2(n14266), .ZN(n14447) );
  NOR2_X1 U14340 ( .A1(n8482), .A2(n8745), .ZN(n14267) );
  NAND2_X1 U14341 ( .A1(n14265), .A2(n14266), .ZN(n14445) );
  NAND2_X1 U14342 ( .A1(n14448), .A2(n14449), .ZN(n14266) );
  NAND2_X1 U14343 ( .A1(n14263), .A2(n14450), .ZN(n14449) );
  OR2_X1 U14344 ( .A1(n14261), .A2(n14262), .ZN(n14450) );
  NOR2_X1 U14345 ( .A1(n8482), .A2(n8744), .ZN(n14263) );
  NAND2_X1 U14346 ( .A1(n14261), .A2(n14262), .ZN(n14448) );
  NAND2_X1 U14347 ( .A1(n14258), .A2(n14451), .ZN(n14262) );
  NAND2_X1 U14348 ( .A1(n14257), .A2(n14259), .ZN(n14451) );
  NAND2_X1 U14349 ( .A1(n14452), .A2(n14453), .ZN(n14259) );
  NAND2_X1 U14350 ( .A1(b_7_), .A2(a_26_), .ZN(n14453) );
  INV_X1 U14351 ( .A(n14454), .ZN(n14452) );
  XNOR2_X1 U14352 ( .A(n14455), .B(n14456), .ZN(n14257) );
  NAND2_X1 U14353 ( .A1(n14457), .A2(n14458), .ZN(n14455) );
  NAND2_X1 U14354 ( .A1(a_26_), .A2(n14454), .ZN(n14258) );
  NAND2_X1 U14355 ( .A1(n14230), .A2(n14459), .ZN(n14454) );
  NAND2_X1 U14356 ( .A1(n14229), .A2(n14231), .ZN(n14459) );
  NAND2_X1 U14357 ( .A1(n14460), .A2(n14461), .ZN(n14231) );
  NAND2_X1 U14358 ( .A1(b_7_), .A2(a_27_), .ZN(n14461) );
  INV_X1 U14359 ( .A(n14462), .ZN(n14460) );
  XNOR2_X1 U14360 ( .A(n14463), .B(n14464), .ZN(n14229) );
  XOR2_X1 U14361 ( .A(n14465), .B(n14466), .Z(n14463) );
  NAND2_X1 U14362 ( .A1(b_6_), .A2(a_28_), .ZN(n14465) );
  NAND2_X1 U14363 ( .A1(a_27_), .A2(n14462), .ZN(n14230) );
  NAND2_X1 U14364 ( .A1(n14467), .A2(n14468), .ZN(n14462) );
  NAND3_X1 U14365 ( .A1(a_28_), .A2(n14469), .A3(b_7_), .ZN(n14468) );
  NAND2_X1 U14366 ( .A1(n14239), .A2(n14237), .ZN(n14469) );
  OR2_X1 U14367 ( .A1(n14237), .A2(n14239), .ZN(n14467) );
  AND2_X1 U14368 ( .A1(n14470), .A2(n14471), .ZN(n14239) );
  NAND2_X1 U14369 ( .A1(n14253), .A2(n14472), .ZN(n14471) );
  OR2_X1 U14370 ( .A1(n14254), .A2(n14255), .ZN(n14472) );
  NOR2_X1 U14371 ( .A1(n8482), .A2(n7890), .ZN(n14253) );
  NAND2_X1 U14372 ( .A1(n14255), .A2(n14254), .ZN(n14470) );
  NAND2_X1 U14373 ( .A1(n14473), .A2(n14474), .ZN(n14254) );
  NAND2_X1 U14374 ( .A1(b_5_), .A2(n14475), .ZN(n14474) );
  NAND2_X1 U14375 ( .A1(n7864), .A2(n14476), .ZN(n14475) );
  NAND2_X1 U14376 ( .A1(a_31_), .A2(n8508), .ZN(n14476) );
  NAND2_X1 U14377 ( .A1(b_6_), .A2(n14477), .ZN(n14473) );
  NAND2_X1 U14378 ( .A1(n9137), .A2(n14478), .ZN(n14477) );
  NAND2_X1 U14379 ( .A1(a_30_), .A2(n8765), .ZN(n14478) );
  AND3_X1 U14380 ( .A1(b_6_), .A2(b_7_), .A3(n7818), .ZN(n14255) );
  XNOR2_X1 U14381 ( .A(n14479), .B(n14480), .ZN(n14237) );
  XOR2_X1 U14382 ( .A(n14481), .B(n14482), .Z(n14479) );
  XNOR2_X1 U14383 ( .A(n14483), .B(n14484), .ZN(n14261) );
  NAND2_X1 U14384 ( .A1(n14485), .A2(n14486), .ZN(n14483) );
  XNOR2_X1 U14385 ( .A(n14487), .B(n14488), .ZN(n14265) );
  NAND2_X1 U14386 ( .A1(n14489), .A2(n14490), .ZN(n14487) );
  XNOR2_X1 U14387 ( .A(n14491), .B(n14492), .ZN(n14269) );
  XNOR2_X1 U14388 ( .A(n14493), .B(n14494), .ZN(n14492) );
  XNOR2_X1 U14389 ( .A(n14495), .B(n14496), .ZN(n14277) );
  NAND2_X1 U14390 ( .A1(n14497), .A2(n14498), .ZN(n14495) );
  XOR2_X1 U14391 ( .A(n14499), .B(n14500), .Z(n14281) );
  XNOR2_X1 U14392 ( .A(n14501), .B(n14502), .ZN(n14500) );
  XNOR2_X1 U14393 ( .A(n14503), .B(n14504), .ZN(n14285) );
  XOR2_X1 U14394 ( .A(n14505), .B(n14506), .Z(n14503) );
  NOR2_X1 U14395 ( .A1(n8751), .A2(n8508), .ZN(n14506) );
  XNOR2_X1 U14396 ( .A(n14507), .B(n14508), .ZN(n14196) );
  XNOR2_X1 U14397 ( .A(n14509), .B(n14510), .ZN(n14508) );
  XNOR2_X1 U14398 ( .A(n14511), .B(n14512), .ZN(n14189) );
  XOR2_X1 U14399 ( .A(n14513), .B(n14514), .Z(n14511) );
  XNOR2_X1 U14400 ( .A(n14515), .B(n14516), .ZN(n14289) );
  XNOR2_X1 U14401 ( .A(n14517), .B(n14518), .ZN(n14515) );
  XNOR2_X1 U14402 ( .A(n14519), .B(n14520), .ZN(n14292) );
  XNOR2_X1 U14403 ( .A(n14521), .B(n14522), .ZN(n14520) );
  XNOR2_X1 U14404 ( .A(n14523), .B(n14524), .ZN(n14297) );
  XNOR2_X1 U14405 ( .A(n14525), .B(n14526), .ZN(n14523) );
  XOR2_X1 U14406 ( .A(n14527), .B(n14528), .Z(n14300) );
  XOR2_X1 U14407 ( .A(n14529), .B(n14530), .Z(n14527) );
  XNOR2_X1 U14408 ( .A(n14531), .B(n14532), .ZN(n14305) );
  XNOR2_X1 U14409 ( .A(n14533), .B(n14534), .ZN(n14531) );
  XNOR2_X1 U14410 ( .A(n14535), .B(n14536), .ZN(n14309) );
  XNOR2_X1 U14411 ( .A(n14537), .B(n14538), .ZN(n14535) );
  XNOR2_X1 U14412 ( .A(n14539), .B(n14540), .ZN(n14313) );
  XNOR2_X1 U14413 ( .A(n14541), .B(n14542), .ZN(n14540) );
  XNOR2_X1 U14414 ( .A(n14543), .B(n14544), .ZN(n14317) );
  XNOR2_X1 U14415 ( .A(n14545), .B(n14546), .ZN(n14543) );
  XNOR2_X1 U14416 ( .A(n14547), .B(n14548), .ZN(n14321) );
  XNOR2_X1 U14417 ( .A(n14549), .B(n14550), .ZN(n14547) );
  NOR2_X1 U14418 ( .A1(n8426), .A2(n8508), .ZN(n14550) );
  INV_X1 U14419 ( .A(n8676), .ZN(n14327) );
  NAND2_X1 U14420 ( .A1(b_7_), .A2(a_7_), .ZN(n8676) );
  XOR2_X1 U14421 ( .A(n14551), .B(n14552), .Z(n14329) );
  XOR2_X1 U14422 ( .A(n14553), .B(n14554), .Z(n14551) );
  NOR2_X1 U14423 ( .A1(n8764), .A2(n8508), .ZN(n14554) );
  XOR2_X1 U14424 ( .A(n14555), .B(n14556), .Z(n14333) );
  XOR2_X1 U14425 ( .A(n14557), .B(n14558), .Z(n14555) );
  XOR2_X1 U14426 ( .A(n14559), .B(n14560), .Z(n14337) );
  XOR2_X1 U14427 ( .A(n14561), .B(n14562), .Z(n14559) );
  NOR2_X1 U14428 ( .A1(n8517), .A2(n8508), .ZN(n14562) );
  XOR2_X1 U14429 ( .A(n14563), .B(n14564), .Z(n14341) );
  XNOR2_X1 U14430 ( .A(n14565), .B(n14566), .ZN(n14564) );
  NAND2_X1 U14431 ( .A1(b_6_), .A2(a_4_), .ZN(n14566) );
  XOR2_X1 U14432 ( .A(n14567), .B(n14568), .Z(n14345) );
  XOR2_X1 U14433 ( .A(n14569), .B(n14570), .Z(n14567) );
  NOR2_X1 U14434 ( .A1(n8567), .A2(n8508), .ZN(n14570) );
  XOR2_X1 U14435 ( .A(n14571), .B(n14572), .Z(n14349) );
  XOR2_X1 U14436 ( .A(n14573), .B(n14574), .Z(n14571) );
  NOR2_X1 U14437 ( .A1(n8768), .A2(n8508), .ZN(n14574) );
  XOR2_X1 U14438 ( .A(n14575), .B(n14576), .Z(n14358) );
  XOR2_X1 U14439 ( .A(n14577), .B(n14578), .Z(n14575) );
  NOR2_X1 U14440 ( .A1(n8617), .A2(n8508), .ZN(n14578) );
  XOR2_X1 U14441 ( .A(n14356), .B(n14579), .Z(n14364) );
  XNOR2_X1 U14442 ( .A(n14580), .B(n14581), .ZN(n14356) );
  NOR2_X1 U14443 ( .A1(n9674), .A2(n8508), .ZN(n14581) );
  NAND2_X1 U14444 ( .A1(n14582), .A2(n14583), .ZN(n7940) );
  NAND2_X1 U14445 ( .A1(n14584), .A2(n14585), .ZN(n14583) );
  NAND2_X1 U14446 ( .A1(n14363), .A2(n14362), .ZN(n14582) );
  NAND4_X1 U14447 ( .A1(n14363), .A2(n14584), .A3(n14585), .A4(n14362), .ZN(
        n7941) );
  NAND2_X1 U14448 ( .A1(n14586), .A2(n14587), .ZN(n14362) );
  NAND3_X1 U14449 ( .A1(a_0_), .A2(n14588), .A3(b_6_), .ZN(n14587) );
  OR2_X1 U14450 ( .A1(n14355), .A2(n14580), .ZN(n14588) );
  NAND2_X1 U14451 ( .A1(n14355), .A2(n14580), .ZN(n14586) );
  NAND2_X1 U14452 ( .A1(n14589), .A2(n14590), .ZN(n14580) );
  NAND3_X1 U14453 ( .A1(a_1_), .A2(n14591), .A3(b_6_), .ZN(n14590) );
  OR2_X1 U14454 ( .A1(n14577), .A2(n14576), .ZN(n14591) );
  NAND2_X1 U14455 ( .A1(n14576), .A2(n14577), .ZN(n14589) );
  NAND2_X1 U14456 ( .A1(n14592), .A2(n14593), .ZN(n14577) );
  NAND3_X1 U14457 ( .A1(a_2_), .A2(n14594), .A3(b_6_), .ZN(n14593) );
  OR2_X1 U14458 ( .A1(n14573), .A2(n14572), .ZN(n14594) );
  NAND2_X1 U14459 ( .A1(n14572), .A2(n14573), .ZN(n14592) );
  NAND2_X1 U14460 ( .A1(n14595), .A2(n14596), .ZN(n14573) );
  NAND3_X1 U14461 ( .A1(a_3_), .A2(n14597), .A3(b_6_), .ZN(n14596) );
  OR2_X1 U14462 ( .A1(n14569), .A2(n14568), .ZN(n14597) );
  NAND2_X1 U14463 ( .A1(n14568), .A2(n14569), .ZN(n14595) );
  NAND2_X1 U14464 ( .A1(n14598), .A2(n14599), .ZN(n14569) );
  NAND3_X1 U14465 ( .A1(a_4_), .A2(n14600), .A3(b_6_), .ZN(n14599) );
  NAND2_X1 U14466 ( .A1(n14565), .A2(n14563), .ZN(n14600) );
  OR2_X1 U14467 ( .A1(n14563), .A2(n14565), .ZN(n14598) );
  AND2_X1 U14468 ( .A1(n14601), .A2(n14602), .ZN(n14565) );
  NAND3_X1 U14469 ( .A1(a_5_), .A2(n14603), .A3(b_6_), .ZN(n14602) );
  OR2_X1 U14470 ( .A1(n14561), .A2(n14560), .ZN(n14603) );
  NAND2_X1 U14471 ( .A1(n14560), .A2(n14561), .ZN(n14601) );
  NAND2_X1 U14472 ( .A1(n14604), .A2(n14605), .ZN(n14561) );
  NAND2_X1 U14473 ( .A1(n14556), .A2(n14606), .ZN(n14605) );
  OR2_X1 U14474 ( .A1(n14557), .A2(n14558), .ZN(n14606) );
  XNOR2_X1 U14475 ( .A(n14607), .B(n14608), .ZN(n14556) );
  XNOR2_X1 U14476 ( .A(n14609), .B(n14610), .ZN(n14607) );
  NOR2_X1 U14477 ( .A1(n8764), .A2(n8765), .ZN(n14610) );
  NAND2_X1 U14478 ( .A1(n14558), .A2(n14557), .ZN(n14604) );
  NAND2_X1 U14479 ( .A1(n14611), .A2(n14612), .ZN(n14557) );
  NAND3_X1 U14480 ( .A1(a_7_), .A2(n14613), .A3(b_6_), .ZN(n14612) );
  OR2_X1 U14481 ( .A1(n14553), .A2(n14552), .ZN(n14613) );
  NAND2_X1 U14482 ( .A1(n14552), .A2(n14553), .ZN(n14611) );
  NAND2_X1 U14483 ( .A1(n14614), .A2(n14615), .ZN(n14553) );
  NAND3_X1 U14484 ( .A1(a_8_), .A2(n14616), .A3(b_6_), .ZN(n14615) );
  OR2_X1 U14485 ( .A1(n14390), .A2(n14388), .ZN(n14616) );
  NAND2_X1 U14486 ( .A1(n14388), .A2(n14390), .ZN(n14614) );
  NAND2_X1 U14487 ( .A1(n14617), .A2(n14618), .ZN(n14390) );
  NAND3_X1 U14488 ( .A1(a_9_), .A2(n14619), .A3(b_6_), .ZN(n14618) );
  NAND2_X1 U14489 ( .A1(n14549), .A2(n14548), .ZN(n14619) );
  OR2_X1 U14490 ( .A1(n14548), .A2(n14549), .ZN(n14617) );
  AND2_X1 U14491 ( .A1(n14620), .A2(n14621), .ZN(n14549) );
  NAND2_X1 U14492 ( .A1(n14546), .A2(n14622), .ZN(n14621) );
  NAND2_X1 U14493 ( .A1(n14545), .A2(n14544), .ZN(n14622) );
  NOR2_X1 U14494 ( .A1(n8508), .A2(n8761), .ZN(n14546) );
  OR2_X1 U14495 ( .A1(n14544), .A2(n14545), .ZN(n14620) );
  AND2_X1 U14496 ( .A1(n14623), .A2(n14624), .ZN(n14545) );
  NAND2_X1 U14497 ( .A1(n14542), .A2(n14625), .ZN(n14624) );
  OR2_X1 U14498 ( .A1(n14541), .A2(n14539), .ZN(n14625) );
  NOR2_X1 U14499 ( .A1(n8508), .A2(n8376), .ZN(n14542) );
  NAND2_X1 U14500 ( .A1(n14539), .A2(n14541), .ZN(n14623) );
  NAND2_X1 U14501 ( .A1(n14626), .A2(n14627), .ZN(n14541) );
  NAND2_X1 U14502 ( .A1(n14538), .A2(n14628), .ZN(n14627) );
  NAND2_X1 U14503 ( .A1(n14537), .A2(n14536), .ZN(n14628) );
  NOR2_X1 U14504 ( .A1(n8508), .A2(n8759), .ZN(n14538) );
  OR2_X1 U14505 ( .A1(n14536), .A2(n14537), .ZN(n14626) );
  AND2_X1 U14506 ( .A1(n14629), .A2(n14630), .ZN(n14537) );
  NAND2_X1 U14507 ( .A1(n14534), .A2(n14631), .ZN(n14630) );
  NAND2_X1 U14508 ( .A1(n14533), .A2(n14532), .ZN(n14631) );
  NOR2_X1 U14509 ( .A1(n8508), .A2(n8310), .ZN(n14534) );
  OR2_X1 U14510 ( .A1(n14532), .A2(n14533), .ZN(n14629) );
  AND2_X1 U14511 ( .A1(n14632), .A2(n14633), .ZN(n14533) );
  NAND2_X1 U14512 ( .A1(n14530), .A2(n14634), .ZN(n14633) );
  OR2_X1 U14513 ( .A1(n14528), .A2(n14529), .ZN(n14634) );
  NOR2_X1 U14514 ( .A1(n8508), .A2(n8757), .ZN(n14530) );
  NAND2_X1 U14515 ( .A1(n14528), .A2(n14529), .ZN(n14632) );
  NAND2_X1 U14516 ( .A1(n14635), .A2(n14636), .ZN(n14529) );
  NAND2_X1 U14517 ( .A1(n14526), .A2(n14637), .ZN(n14636) );
  NAND2_X1 U14518 ( .A1(n14525), .A2(n14524), .ZN(n14637) );
  NOR2_X1 U14519 ( .A1(n8508), .A2(n8276), .ZN(n14526) );
  OR2_X1 U14520 ( .A1(n14524), .A2(n14525), .ZN(n14635) );
  AND2_X1 U14521 ( .A1(n14638), .A2(n14639), .ZN(n14525) );
  NAND2_X1 U14522 ( .A1(n14522), .A2(n14640), .ZN(n14639) );
  OR2_X1 U14523 ( .A1(n14519), .A2(n14521), .ZN(n14640) );
  NOR2_X1 U14524 ( .A1(n8508), .A2(n8755), .ZN(n14522) );
  NAND2_X1 U14525 ( .A1(n14519), .A2(n14521), .ZN(n14638) );
  NAND2_X1 U14526 ( .A1(n14641), .A2(n14642), .ZN(n14521) );
  NAND2_X1 U14527 ( .A1(n14518), .A2(n14643), .ZN(n14642) );
  NAND2_X1 U14528 ( .A1(n14517), .A2(n14516), .ZN(n14643) );
  NOR2_X1 U14529 ( .A1(n8508), .A2(n8210), .ZN(n14518) );
  OR2_X1 U14530 ( .A1(n14516), .A2(n14517), .ZN(n14641) );
  AND2_X1 U14531 ( .A1(n14644), .A2(n14645), .ZN(n14517) );
  NAND2_X1 U14532 ( .A1(n14513), .A2(n14646), .ZN(n14645) );
  OR2_X1 U14533 ( .A1(n14512), .A2(n14514), .ZN(n14646) );
  NOR2_X1 U14534 ( .A1(n8508), .A2(n8753), .ZN(n14513) );
  NAND2_X1 U14535 ( .A1(n14512), .A2(n14514), .ZN(n14644) );
  NAND2_X1 U14536 ( .A1(n14647), .A2(n14648), .ZN(n14514) );
  NAND2_X1 U14537 ( .A1(n14510), .A2(n14649), .ZN(n14648) );
  OR2_X1 U14538 ( .A1(n14509), .A2(n14507), .ZN(n14649) );
  NOR2_X1 U14539 ( .A1(n8508), .A2(n8170), .ZN(n14510) );
  NAND2_X1 U14540 ( .A1(n14507), .A2(n14509), .ZN(n14647) );
  NAND2_X1 U14541 ( .A1(n14650), .A2(n14651), .ZN(n14509) );
  NAND3_X1 U14542 ( .A1(a_20_), .A2(n14652), .A3(b_6_), .ZN(n14651) );
  OR2_X1 U14543 ( .A1(n14504), .A2(n14505), .ZN(n14652) );
  NAND2_X1 U14544 ( .A1(n14504), .A2(n14505), .ZN(n14650) );
  NAND2_X1 U14545 ( .A1(n14653), .A2(n14654), .ZN(n14505) );
  NAND2_X1 U14546 ( .A1(n14502), .A2(n14655), .ZN(n14654) );
  OR2_X1 U14547 ( .A1(n14499), .A2(n14501), .ZN(n14655) );
  NOR2_X1 U14548 ( .A1(n8508), .A2(n8750), .ZN(n14502) );
  NAND2_X1 U14549 ( .A1(n14499), .A2(n14501), .ZN(n14653) );
  NAND2_X1 U14550 ( .A1(n14497), .A2(n14656), .ZN(n14501) );
  NAND2_X1 U14551 ( .A1(n14496), .A2(n14498), .ZN(n14656) );
  NAND2_X1 U14552 ( .A1(n14657), .A2(n14658), .ZN(n14498) );
  NAND2_X1 U14553 ( .A1(b_6_), .A2(a_22_), .ZN(n14658) );
  INV_X1 U14554 ( .A(n14659), .ZN(n14657) );
  XNOR2_X1 U14555 ( .A(n14660), .B(n14661), .ZN(n14496) );
  XOR2_X1 U14556 ( .A(n14662), .B(n14663), .Z(n14661) );
  NAND2_X1 U14557 ( .A1(b_5_), .A2(a_23_), .ZN(n14663) );
  NAND2_X1 U14558 ( .A1(a_22_), .A2(n14659), .ZN(n14497) );
  NAND2_X1 U14559 ( .A1(n14664), .A2(n14665), .ZN(n14659) );
  NAND3_X1 U14560 ( .A1(a_23_), .A2(n14666), .A3(b_6_), .ZN(n14665) );
  OR2_X1 U14561 ( .A1(n14439), .A2(n14440), .ZN(n14666) );
  NAND2_X1 U14562 ( .A1(n14439), .A2(n14440), .ZN(n14664) );
  NAND2_X1 U14563 ( .A1(n14667), .A2(n14668), .ZN(n14440) );
  NAND2_X1 U14564 ( .A1(n14494), .A2(n14669), .ZN(n14668) );
  OR2_X1 U14565 ( .A1(n14493), .A2(n14491), .ZN(n14669) );
  NOR2_X1 U14566 ( .A1(n8508), .A2(n8745), .ZN(n14494) );
  NAND2_X1 U14567 ( .A1(n14491), .A2(n14493), .ZN(n14667) );
  NAND2_X1 U14568 ( .A1(n14489), .A2(n14670), .ZN(n14493) );
  NAND2_X1 U14569 ( .A1(n14488), .A2(n14490), .ZN(n14670) );
  NAND2_X1 U14570 ( .A1(n14671), .A2(n14672), .ZN(n14490) );
  NAND2_X1 U14571 ( .A1(b_6_), .A2(a_25_), .ZN(n14672) );
  INV_X1 U14572 ( .A(n14673), .ZN(n14671) );
  XNOR2_X1 U14573 ( .A(n14674), .B(n14675), .ZN(n14488) );
  NAND2_X1 U14574 ( .A1(n14676), .A2(n14677), .ZN(n14674) );
  NAND2_X1 U14575 ( .A1(a_25_), .A2(n14673), .ZN(n14489) );
  NAND2_X1 U14576 ( .A1(n14485), .A2(n14678), .ZN(n14673) );
  NAND2_X1 U14577 ( .A1(n14484), .A2(n14486), .ZN(n14678) );
  NAND2_X1 U14578 ( .A1(n14679), .A2(n14680), .ZN(n14486) );
  NAND2_X1 U14579 ( .A1(b_6_), .A2(a_26_), .ZN(n14680) );
  INV_X1 U14580 ( .A(n14681), .ZN(n14679) );
  XNOR2_X1 U14581 ( .A(n14682), .B(n14683), .ZN(n14484) );
  NAND2_X1 U14582 ( .A1(n14684), .A2(n14685), .ZN(n14682) );
  NAND2_X1 U14583 ( .A1(a_26_), .A2(n14681), .ZN(n14485) );
  NAND2_X1 U14584 ( .A1(n14457), .A2(n14686), .ZN(n14681) );
  NAND2_X1 U14585 ( .A1(n14456), .A2(n14458), .ZN(n14686) );
  NAND2_X1 U14586 ( .A1(n14687), .A2(n14688), .ZN(n14458) );
  NAND2_X1 U14587 ( .A1(b_6_), .A2(a_27_), .ZN(n14688) );
  INV_X1 U14588 ( .A(n14689), .ZN(n14687) );
  XNOR2_X1 U14589 ( .A(n14690), .B(n14691), .ZN(n14456) );
  XOR2_X1 U14590 ( .A(n14692), .B(n14693), .Z(n14690) );
  NAND2_X1 U14591 ( .A1(b_5_), .A2(a_28_), .ZN(n14692) );
  NAND2_X1 U14592 ( .A1(a_27_), .A2(n14689), .ZN(n14457) );
  NAND2_X1 U14593 ( .A1(n14694), .A2(n14695), .ZN(n14689) );
  NAND3_X1 U14594 ( .A1(a_28_), .A2(n14696), .A3(b_6_), .ZN(n14695) );
  NAND2_X1 U14595 ( .A1(n14466), .A2(n14464), .ZN(n14696) );
  OR2_X1 U14596 ( .A1(n14464), .A2(n14466), .ZN(n14694) );
  AND2_X1 U14597 ( .A1(n14697), .A2(n14698), .ZN(n14466) );
  NAND2_X1 U14598 ( .A1(n14480), .A2(n14699), .ZN(n14698) );
  OR2_X1 U14599 ( .A1(n14481), .A2(n14482), .ZN(n14699) );
  NOR2_X1 U14600 ( .A1(n8508), .A2(n7890), .ZN(n14480) );
  NAND2_X1 U14601 ( .A1(n14482), .A2(n14481), .ZN(n14697) );
  NAND2_X1 U14602 ( .A1(n14700), .A2(n14701), .ZN(n14481) );
  NAND2_X1 U14603 ( .A1(b_4_), .A2(n14702), .ZN(n14701) );
  NAND2_X1 U14604 ( .A1(n7864), .A2(n14703), .ZN(n14702) );
  NAND2_X1 U14605 ( .A1(a_31_), .A2(n8765), .ZN(n14703) );
  NAND2_X1 U14606 ( .A1(b_5_), .A2(n14704), .ZN(n14700) );
  NAND2_X1 U14607 ( .A1(n9137), .A2(n14705), .ZN(n14704) );
  NAND2_X1 U14608 ( .A1(a_30_), .A2(n8558), .ZN(n14705) );
  AND3_X1 U14609 ( .A1(b_5_), .A2(b_6_), .A3(n7818), .ZN(n14482) );
  XNOR2_X1 U14610 ( .A(n14706), .B(n14707), .ZN(n14464) );
  XOR2_X1 U14611 ( .A(n14708), .B(n14709), .Z(n14706) );
  XNOR2_X1 U14612 ( .A(n14710), .B(n14711), .ZN(n14491) );
  NAND2_X1 U14613 ( .A1(n14712), .A2(n14713), .ZN(n14710) );
  XNOR2_X1 U14614 ( .A(n14714), .B(n14715), .ZN(n14439) );
  XOR2_X1 U14615 ( .A(n14716), .B(n14717), .Z(n14715) );
  NAND2_X1 U14616 ( .A1(b_5_), .A2(a_24_), .ZN(n14717) );
  XNOR2_X1 U14617 ( .A(n14718), .B(n14719), .ZN(n14499) );
  XOR2_X1 U14618 ( .A(n14720), .B(n14721), .Z(n14719) );
  NAND2_X1 U14619 ( .A1(b_5_), .A2(a_22_), .ZN(n14721) );
  XNOR2_X1 U14620 ( .A(n14722), .B(n14723), .ZN(n14504) );
  XNOR2_X1 U14621 ( .A(n14724), .B(n14725), .ZN(n14722) );
  NOR2_X1 U14622 ( .A1(n8750), .A2(n8765), .ZN(n14725) );
  XOR2_X1 U14623 ( .A(n14726), .B(n14727), .Z(n14507) );
  XOR2_X1 U14624 ( .A(n14728), .B(n14729), .Z(n14726) );
  NOR2_X1 U14625 ( .A1(n8751), .A2(n8765), .ZN(n14729) );
  XNOR2_X1 U14626 ( .A(n14730), .B(n14731), .ZN(n14512) );
  XOR2_X1 U14627 ( .A(n14732), .B(n14733), .Z(n14731) );
  NAND2_X1 U14628 ( .A1(b_5_), .A2(a_19_), .ZN(n14733) );
  XNOR2_X1 U14629 ( .A(n14734), .B(n14735), .ZN(n14516) );
  XOR2_X1 U14630 ( .A(n14736), .B(n14737), .Z(n14734) );
  NOR2_X1 U14631 ( .A1(n8753), .A2(n8765), .ZN(n14737) );
  XNOR2_X1 U14632 ( .A(n14738), .B(n14739), .ZN(n14519) );
  XNOR2_X1 U14633 ( .A(n14740), .B(n14741), .ZN(n14738) );
  NOR2_X1 U14634 ( .A1(n8210), .A2(n8765), .ZN(n14741) );
  XNOR2_X1 U14635 ( .A(n14742), .B(n14743), .ZN(n14524) );
  XOR2_X1 U14636 ( .A(n14744), .B(n14745), .Z(n14742) );
  NOR2_X1 U14637 ( .A1(n8755), .A2(n8765), .ZN(n14745) );
  XNOR2_X1 U14638 ( .A(n14746), .B(n14747), .ZN(n14528) );
  XNOR2_X1 U14639 ( .A(n14748), .B(n14749), .ZN(n14746) );
  NOR2_X1 U14640 ( .A1(n8276), .A2(n8765), .ZN(n14749) );
  XNOR2_X1 U14641 ( .A(n14750), .B(n14751), .ZN(n14532) );
  XOR2_X1 U14642 ( .A(n14752), .B(n14753), .Z(n14750) );
  NOR2_X1 U14643 ( .A1(n8757), .A2(n8765), .ZN(n14753) );
  XNOR2_X1 U14644 ( .A(n14754), .B(n14755), .ZN(n14536) );
  XOR2_X1 U14645 ( .A(n14756), .B(n14757), .Z(n14754) );
  NOR2_X1 U14646 ( .A1(n8310), .A2(n8765), .ZN(n14757) );
  XOR2_X1 U14647 ( .A(n14758), .B(n14759), .Z(n14539) );
  XOR2_X1 U14648 ( .A(n14760), .B(n14761), .Z(n14758) );
  NOR2_X1 U14649 ( .A1(n8759), .A2(n8765), .ZN(n14761) );
  XNOR2_X1 U14650 ( .A(n14762), .B(n14763), .ZN(n14544) );
  XOR2_X1 U14651 ( .A(n14764), .B(n14765), .Z(n14762) );
  NOR2_X1 U14652 ( .A1(n8376), .A2(n8765), .ZN(n14765) );
  XNOR2_X1 U14653 ( .A(n14766), .B(n14767), .ZN(n14548) );
  XOR2_X1 U14654 ( .A(n14768), .B(n14769), .Z(n14766) );
  NOR2_X1 U14655 ( .A1(n8761), .A2(n8765), .ZN(n14769) );
  XNOR2_X1 U14656 ( .A(n14770), .B(n14771), .ZN(n14388) );
  XNOR2_X1 U14657 ( .A(n14772), .B(n14773), .ZN(n14770) );
  NOR2_X1 U14658 ( .A1(n8426), .A2(n8765), .ZN(n14773) );
  XOR2_X1 U14659 ( .A(n14774), .B(n14775), .Z(n14552) );
  XOR2_X1 U14660 ( .A(n14776), .B(n14777), .Z(n14774) );
  NOR2_X1 U14661 ( .A1(n8763), .A2(n8765), .ZN(n14777) );
  INV_X1 U14662 ( .A(n8673), .ZN(n14558) );
  NAND2_X1 U14663 ( .A1(b_6_), .A2(a_6_), .ZN(n8673) );
  XOR2_X1 U14664 ( .A(n14778), .B(n14779), .Z(n14560) );
  XOR2_X1 U14665 ( .A(n14780), .B(n14781), .Z(n14778) );
  NOR2_X1 U14666 ( .A1(n8491), .A2(n8765), .ZN(n14781) );
  XNOR2_X1 U14667 ( .A(n14782), .B(n14783), .ZN(n14563) );
  XOR2_X1 U14668 ( .A(n14784), .B(n14785), .Z(n14782) );
  XOR2_X1 U14669 ( .A(n14786), .B(n14787), .Z(n14568) );
  XOR2_X1 U14670 ( .A(n14788), .B(n14789), .Z(n14786) );
  NOR2_X1 U14671 ( .A1(n8766), .A2(n8765), .ZN(n14789) );
  XOR2_X1 U14672 ( .A(n14790), .B(n14791), .Z(n14572) );
  XOR2_X1 U14673 ( .A(n14792), .B(n14793), .Z(n14790) );
  NOR2_X1 U14674 ( .A1(n8567), .A2(n8765), .ZN(n14793) );
  XOR2_X1 U14675 ( .A(n14794), .B(n14795), .Z(n14576) );
  XOR2_X1 U14676 ( .A(n14796), .B(n14797), .Z(n14794) );
  NOR2_X1 U14677 ( .A1(n8768), .A2(n8765), .ZN(n14797) );
  INV_X1 U14678 ( .A(n14579), .ZN(n14355) );
  XNOR2_X1 U14679 ( .A(n14798), .B(n14799), .ZN(n14579) );
  XOR2_X1 U14680 ( .A(n14800), .B(n14801), .Z(n14798) );
  NOR2_X1 U14681 ( .A1(n8617), .A2(n8765), .ZN(n14801) );
  NAND3_X1 U14682 ( .A1(n14802), .A2(n14803), .A3(n14804), .ZN(n14584) );
  XOR2_X1 U14683 ( .A(n14805), .B(n14806), .Z(n14804) );
  XOR2_X1 U14684 ( .A(n14807), .B(n14808), .Z(n14363) );
  XOR2_X1 U14685 ( .A(n14809), .B(n14810), .Z(n14807) );
  NAND2_X1 U14686 ( .A1(n14811), .A2(n14585), .ZN(n8200) );
  OR2_X1 U14687 ( .A1(n14585), .A2(n14811), .ZN(n8201) );
  XNOR2_X1 U14688 ( .A(n14812), .B(n14813), .ZN(n14811) );
  NAND2_X1 U14689 ( .A1(n14814), .A2(n14815), .ZN(n14585) );
  NAND2_X1 U14690 ( .A1(n14802), .A2(n14803), .ZN(n14815) );
  NAND2_X1 U14691 ( .A1(n14810), .A2(n14816), .ZN(n14803) );
  OR2_X1 U14692 ( .A1(n14808), .A2(n14809), .ZN(n14816) );
  NOR2_X1 U14693 ( .A1(n8765), .A2(n9674), .ZN(n14810) );
  NAND2_X1 U14694 ( .A1(n14808), .A2(n14809), .ZN(n14802) );
  NAND2_X1 U14695 ( .A1(n14817), .A2(n14818), .ZN(n14809) );
  NAND3_X1 U14696 ( .A1(a_1_), .A2(n14819), .A3(b_5_), .ZN(n14818) );
  OR2_X1 U14697 ( .A1(n14800), .A2(n14799), .ZN(n14819) );
  NAND2_X1 U14698 ( .A1(n14799), .A2(n14800), .ZN(n14817) );
  NAND2_X1 U14699 ( .A1(n14820), .A2(n14821), .ZN(n14800) );
  NAND3_X1 U14700 ( .A1(a_2_), .A2(n14822), .A3(b_5_), .ZN(n14821) );
  OR2_X1 U14701 ( .A1(n14795), .A2(n14796), .ZN(n14822) );
  NAND2_X1 U14702 ( .A1(n14795), .A2(n14796), .ZN(n14820) );
  NAND2_X1 U14703 ( .A1(n14823), .A2(n14824), .ZN(n14796) );
  NAND3_X1 U14704 ( .A1(a_3_), .A2(n14825), .A3(b_5_), .ZN(n14824) );
  OR2_X1 U14705 ( .A1(n14791), .A2(n14792), .ZN(n14825) );
  NAND2_X1 U14706 ( .A1(n14791), .A2(n14792), .ZN(n14823) );
  NAND2_X1 U14707 ( .A1(n14826), .A2(n14827), .ZN(n14792) );
  NAND3_X1 U14708 ( .A1(a_4_), .A2(n14828), .A3(b_5_), .ZN(n14827) );
  OR2_X1 U14709 ( .A1(n14787), .A2(n14788), .ZN(n14828) );
  NAND2_X1 U14710 ( .A1(n14787), .A2(n14788), .ZN(n14826) );
  NAND2_X1 U14711 ( .A1(n14829), .A2(n14830), .ZN(n14788) );
  NAND2_X1 U14712 ( .A1(n14783), .A2(n14831), .ZN(n14830) );
  OR2_X1 U14713 ( .A1(n14784), .A2(n14785), .ZN(n14831) );
  XNOR2_X1 U14714 ( .A(n14832), .B(n14833), .ZN(n14783) );
  XNOR2_X1 U14715 ( .A(n14834), .B(n14835), .ZN(n14832) );
  NOR2_X1 U14716 ( .A1(n8491), .A2(n8558), .ZN(n14835) );
  NAND2_X1 U14717 ( .A1(n14785), .A2(n14784), .ZN(n14829) );
  NAND2_X1 U14718 ( .A1(n14836), .A2(n14837), .ZN(n14784) );
  NAND3_X1 U14719 ( .A1(a_6_), .A2(n14838), .A3(b_5_), .ZN(n14837) );
  OR2_X1 U14720 ( .A1(n14779), .A2(n14780), .ZN(n14838) );
  NAND2_X1 U14721 ( .A1(n14779), .A2(n14780), .ZN(n14836) );
  NAND2_X1 U14722 ( .A1(n14839), .A2(n14840), .ZN(n14780) );
  NAND3_X1 U14723 ( .A1(a_7_), .A2(n14841), .A3(b_5_), .ZN(n14840) );
  NAND2_X1 U14724 ( .A1(n14608), .A2(n14609), .ZN(n14841) );
  OR2_X1 U14725 ( .A1(n14608), .A2(n14609), .ZN(n14839) );
  AND2_X1 U14726 ( .A1(n14842), .A2(n14843), .ZN(n14609) );
  NAND3_X1 U14727 ( .A1(a_8_), .A2(n14844), .A3(b_5_), .ZN(n14843) );
  OR2_X1 U14728 ( .A1(n14775), .A2(n14776), .ZN(n14844) );
  NAND2_X1 U14729 ( .A1(n14775), .A2(n14776), .ZN(n14842) );
  NAND2_X1 U14730 ( .A1(n14845), .A2(n14846), .ZN(n14776) );
  NAND3_X1 U14731 ( .A1(a_9_), .A2(n14847), .A3(b_5_), .ZN(n14846) );
  NAND2_X1 U14732 ( .A1(n14771), .A2(n14772), .ZN(n14847) );
  OR2_X1 U14733 ( .A1(n14771), .A2(n14772), .ZN(n14845) );
  AND2_X1 U14734 ( .A1(n14848), .A2(n14849), .ZN(n14772) );
  NAND3_X1 U14735 ( .A1(a_10_), .A2(n14850), .A3(b_5_), .ZN(n14849) );
  OR2_X1 U14736 ( .A1(n14767), .A2(n14768), .ZN(n14850) );
  NAND2_X1 U14737 ( .A1(n14767), .A2(n14768), .ZN(n14848) );
  NAND2_X1 U14738 ( .A1(n14851), .A2(n14852), .ZN(n14768) );
  NAND3_X1 U14739 ( .A1(a_11_), .A2(n14853), .A3(b_5_), .ZN(n14852) );
  OR2_X1 U14740 ( .A1(n14763), .A2(n14764), .ZN(n14853) );
  NAND2_X1 U14741 ( .A1(n14763), .A2(n14764), .ZN(n14851) );
  NAND2_X1 U14742 ( .A1(n14854), .A2(n14855), .ZN(n14764) );
  NAND3_X1 U14743 ( .A1(a_12_), .A2(n14856), .A3(b_5_), .ZN(n14855) );
  OR2_X1 U14744 ( .A1(n14759), .A2(n14760), .ZN(n14856) );
  NAND2_X1 U14745 ( .A1(n14759), .A2(n14760), .ZN(n14854) );
  NAND2_X1 U14746 ( .A1(n14857), .A2(n14858), .ZN(n14760) );
  NAND3_X1 U14747 ( .A1(a_13_), .A2(n14859), .A3(b_5_), .ZN(n14858) );
  OR2_X1 U14748 ( .A1(n14755), .A2(n14756), .ZN(n14859) );
  NAND2_X1 U14749 ( .A1(n14755), .A2(n14756), .ZN(n14857) );
  NAND2_X1 U14750 ( .A1(n14860), .A2(n14861), .ZN(n14756) );
  NAND3_X1 U14751 ( .A1(a_14_), .A2(n14862), .A3(b_5_), .ZN(n14861) );
  OR2_X1 U14752 ( .A1(n14751), .A2(n14752), .ZN(n14862) );
  NAND2_X1 U14753 ( .A1(n14751), .A2(n14752), .ZN(n14860) );
  NAND2_X1 U14754 ( .A1(n14863), .A2(n14864), .ZN(n14752) );
  NAND3_X1 U14755 ( .A1(a_15_), .A2(n14865), .A3(b_5_), .ZN(n14864) );
  NAND2_X1 U14756 ( .A1(n14748), .A2(n14747), .ZN(n14865) );
  OR2_X1 U14757 ( .A1(n14747), .A2(n14748), .ZN(n14863) );
  AND2_X1 U14758 ( .A1(n14866), .A2(n14867), .ZN(n14748) );
  NAND3_X1 U14759 ( .A1(a_16_), .A2(n14868), .A3(b_5_), .ZN(n14867) );
  OR2_X1 U14760 ( .A1(n14743), .A2(n14744), .ZN(n14868) );
  NAND2_X1 U14761 ( .A1(n14743), .A2(n14744), .ZN(n14866) );
  NAND2_X1 U14762 ( .A1(n14869), .A2(n14870), .ZN(n14744) );
  NAND3_X1 U14763 ( .A1(a_17_), .A2(n14871), .A3(b_5_), .ZN(n14870) );
  NAND2_X1 U14764 ( .A1(n14740), .A2(n14739), .ZN(n14871) );
  OR2_X1 U14765 ( .A1(n14739), .A2(n14740), .ZN(n14869) );
  AND2_X1 U14766 ( .A1(n14872), .A2(n14873), .ZN(n14740) );
  NAND3_X1 U14767 ( .A1(a_18_), .A2(n14874), .A3(b_5_), .ZN(n14873) );
  OR2_X1 U14768 ( .A1(n14735), .A2(n14736), .ZN(n14874) );
  NAND2_X1 U14769 ( .A1(n14735), .A2(n14736), .ZN(n14872) );
  NAND2_X1 U14770 ( .A1(n14875), .A2(n14876), .ZN(n14736) );
  NAND3_X1 U14771 ( .A1(a_19_), .A2(n14877), .A3(b_5_), .ZN(n14876) );
  OR2_X1 U14772 ( .A1(n14732), .A2(n14730), .ZN(n14877) );
  NAND2_X1 U14773 ( .A1(n14730), .A2(n14732), .ZN(n14875) );
  NAND2_X1 U14774 ( .A1(n14878), .A2(n14879), .ZN(n14732) );
  NAND3_X1 U14775 ( .A1(a_20_), .A2(n14880), .A3(b_5_), .ZN(n14879) );
  OR2_X1 U14776 ( .A1(n14727), .A2(n14728), .ZN(n14880) );
  NAND2_X1 U14777 ( .A1(n14727), .A2(n14728), .ZN(n14878) );
  NAND2_X1 U14778 ( .A1(n14881), .A2(n14882), .ZN(n14728) );
  NAND3_X1 U14779 ( .A1(a_21_), .A2(n14883), .A3(b_5_), .ZN(n14882) );
  NAND2_X1 U14780 ( .A1(n14724), .A2(n14723), .ZN(n14883) );
  OR2_X1 U14781 ( .A1(n14723), .A2(n14724), .ZN(n14881) );
  AND2_X1 U14782 ( .A1(n14884), .A2(n14885), .ZN(n14724) );
  NAND3_X1 U14783 ( .A1(a_22_), .A2(n14886), .A3(b_5_), .ZN(n14885) );
  OR2_X1 U14784 ( .A1(n14720), .A2(n14718), .ZN(n14886) );
  NAND2_X1 U14785 ( .A1(n14718), .A2(n14720), .ZN(n14884) );
  NAND2_X1 U14786 ( .A1(n14887), .A2(n14888), .ZN(n14720) );
  NAND3_X1 U14787 ( .A1(a_23_), .A2(n14889), .A3(b_5_), .ZN(n14888) );
  OR2_X1 U14788 ( .A1(n14662), .A2(n14660), .ZN(n14889) );
  NAND2_X1 U14789 ( .A1(n14660), .A2(n14662), .ZN(n14887) );
  NAND2_X1 U14790 ( .A1(n14890), .A2(n14891), .ZN(n14662) );
  NAND3_X1 U14791 ( .A1(a_24_), .A2(n14892), .A3(b_5_), .ZN(n14891) );
  OR2_X1 U14792 ( .A1(n14716), .A2(n14714), .ZN(n14892) );
  NAND2_X1 U14793 ( .A1(n14714), .A2(n14716), .ZN(n14890) );
  NAND2_X1 U14794 ( .A1(n14712), .A2(n14893), .ZN(n14716) );
  NAND2_X1 U14795 ( .A1(n14711), .A2(n14713), .ZN(n14893) );
  NAND2_X1 U14796 ( .A1(n14894), .A2(n14895), .ZN(n14713) );
  NAND2_X1 U14797 ( .A1(b_5_), .A2(a_25_), .ZN(n14895) );
  INV_X1 U14798 ( .A(n14896), .ZN(n14894) );
  XNOR2_X1 U14799 ( .A(n14897), .B(n14898), .ZN(n14711) );
  NAND2_X1 U14800 ( .A1(n14899), .A2(n14900), .ZN(n14897) );
  NAND2_X1 U14801 ( .A1(a_25_), .A2(n14896), .ZN(n14712) );
  NAND2_X1 U14802 ( .A1(n14676), .A2(n14901), .ZN(n14896) );
  NAND2_X1 U14803 ( .A1(n14675), .A2(n14677), .ZN(n14901) );
  NAND2_X1 U14804 ( .A1(n14902), .A2(n14903), .ZN(n14677) );
  NAND2_X1 U14805 ( .A1(b_5_), .A2(a_26_), .ZN(n14903) );
  INV_X1 U14806 ( .A(n14904), .ZN(n14902) );
  XNOR2_X1 U14807 ( .A(n14905), .B(n14906), .ZN(n14675) );
  NAND2_X1 U14808 ( .A1(n14907), .A2(n14908), .ZN(n14905) );
  NAND2_X1 U14809 ( .A1(a_26_), .A2(n14904), .ZN(n14676) );
  NAND2_X1 U14810 ( .A1(n14684), .A2(n14909), .ZN(n14904) );
  NAND2_X1 U14811 ( .A1(n14683), .A2(n14685), .ZN(n14909) );
  NAND2_X1 U14812 ( .A1(n14910), .A2(n14911), .ZN(n14685) );
  NAND2_X1 U14813 ( .A1(b_5_), .A2(a_27_), .ZN(n14911) );
  INV_X1 U14814 ( .A(n14912), .ZN(n14910) );
  XNOR2_X1 U14815 ( .A(n14913), .B(n14914), .ZN(n14683) );
  XOR2_X1 U14816 ( .A(n14915), .B(n14916), .Z(n14913) );
  NAND2_X1 U14817 ( .A1(b_4_), .A2(a_28_), .ZN(n14915) );
  NAND2_X1 U14818 ( .A1(a_27_), .A2(n14912), .ZN(n14684) );
  NAND2_X1 U14819 ( .A1(n14917), .A2(n14918), .ZN(n14912) );
  NAND3_X1 U14820 ( .A1(a_28_), .A2(n14919), .A3(b_5_), .ZN(n14918) );
  NAND2_X1 U14821 ( .A1(n14693), .A2(n14691), .ZN(n14919) );
  OR2_X1 U14822 ( .A1(n14691), .A2(n14693), .ZN(n14917) );
  AND2_X1 U14823 ( .A1(n14920), .A2(n14921), .ZN(n14693) );
  NAND2_X1 U14824 ( .A1(n14707), .A2(n14922), .ZN(n14921) );
  OR2_X1 U14825 ( .A1(n14708), .A2(n14709), .ZN(n14922) );
  NOR2_X1 U14826 ( .A1(n8765), .A2(n7890), .ZN(n14707) );
  NAND2_X1 U14827 ( .A1(n14709), .A2(n14708), .ZN(n14920) );
  NAND2_X1 U14828 ( .A1(n14923), .A2(n14924), .ZN(n14708) );
  NAND2_X1 U14829 ( .A1(b_3_), .A2(n14925), .ZN(n14924) );
  NAND2_X1 U14830 ( .A1(n7864), .A2(n14926), .ZN(n14925) );
  NAND2_X1 U14831 ( .A1(a_31_), .A2(n8558), .ZN(n14926) );
  NAND2_X1 U14832 ( .A1(b_4_), .A2(n14927), .ZN(n14923) );
  NAND2_X1 U14833 ( .A1(n9137), .A2(n14928), .ZN(n14927) );
  NAND2_X1 U14834 ( .A1(a_30_), .A2(n8767), .ZN(n14928) );
  AND3_X1 U14835 ( .A1(b_4_), .A2(b_5_), .A3(n7818), .ZN(n14709) );
  XNOR2_X1 U14836 ( .A(n14929), .B(n14930), .ZN(n14691) );
  XOR2_X1 U14837 ( .A(n14931), .B(n14932), .Z(n14929) );
  XOR2_X1 U14838 ( .A(n14933), .B(n14934), .Z(n14714) );
  XOR2_X1 U14839 ( .A(n14935), .B(n14936), .Z(n14933) );
  XOR2_X1 U14840 ( .A(n14937), .B(n14938), .Z(n14660) );
  XOR2_X1 U14841 ( .A(n14939), .B(n14940), .Z(n14937) );
  XOR2_X1 U14842 ( .A(n14941), .B(n14942), .Z(n14718) );
  XOR2_X1 U14843 ( .A(n14943), .B(n14944), .Z(n14941) );
  XOR2_X1 U14844 ( .A(n14945), .B(n14946), .Z(n14723) );
  XNOR2_X1 U14845 ( .A(n14947), .B(n14948), .ZN(n14946) );
  XNOR2_X1 U14846 ( .A(n14949), .B(n14950), .ZN(n14727) );
  XNOR2_X1 U14847 ( .A(n14951), .B(n14952), .ZN(n14949) );
  XOR2_X1 U14848 ( .A(n14953), .B(n14954), .Z(n14730) );
  XOR2_X1 U14849 ( .A(n14955), .B(n14956), .Z(n14953) );
  XNOR2_X1 U14850 ( .A(n14957), .B(n14958), .ZN(n14735) );
  XNOR2_X1 U14851 ( .A(n14959), .B(n14960), .ZN(n14957) );
  XNOR2_X1 U14852 ( .A(n14961), .B(n14962), .ZN(n14739) );
  XOR2_X1 U14853 ( .A(n14963), .B(n14964), .Z(n14961) );
  XNOR2_X1 U14854 ( .A(n14965), .B(n14966), .ZN(n14743) );
  XNOR2_X1 U14855 ( .A(n14967), .B(n14968), .ZN(n14965) );
  XNOR2_X1 U14856 ( .A(n14969), .B(n14970), .ZN(n14747) );
  XOR2_X1 U14857 ( .A(n14971), .B(n14972), .Z(n14969) );
  XNOR2_X1 U14858 ( .A(n14973), .B(n14974), .ZN(n14751) );
  XNOR2_X1 U14859 ( .A(n14975), .B(n14976), .ZN(n14973) );
  XNOR2_X1 U14860 ( .A(n14977), .B(n14978), .ZN(n14755) );
  XNOR2_X1 U14861 ( .A(n14979), .B(n14980), .ZN(n14977) );
  XNOR2_X1 U14862 ( .A(n14981), .B(n14982), .ZN(n14759) );
  XNOR2_X1 U14863 ( .A(n14983), .B(n14984), .ZN(n14981) );
  NOR2_X1 U14864 ( .A1(n8310), .A2(n8558), .ZN(n14984) );
  XNOR2_X1 U14865 ( .A(n14985), .B(n14986), .ZN(n14763) );
  XNOR2_X1 U14866 ( .A(n14987), .B(n14988), .ZN(n14985) );
  NOR2_X1 U14867 ( .A1(n8759), .A2(n8558), .ZN(n14988) );
  XOR2_X1 U14868 ( .A(n14989), .B(n14990), .Z(n14767) );
  XNOR2_X1 U14869 ( .A(n14991), .B(n14992), .ZN(n14990) );
  NAND2_X1 U14870 ( .A1(b_4_), .A2(a_11_), .ZN(n14992) );
  XNOR2_X1 U14871 ( .A(n14993), .B(n14994), .ZN(n14771) );
  XNOR2_X1 U14872 ( .A(n14995), .B(n14996), .ZN(n14994) );
  NAND2_X1 U14873 ( .A1(b_4_), .A2(a_10_), .ZN(n14996) );
  XOR2_X1 U14874 ( .A(n14997), .B(n14998), .Z(n14775) );
  XNOR2_X1 U14875 ( .A(n14999), .B(n15000), .ZN(n14998) );
  NAND2_X1 U14876 ( .A1(b_4_), .A2(a_9_), .ZN(n15000) );
  XNOR2_X1 U14877 ( .A(n15001), .B(n15002), .ZN(n14608) );
  XOR2_X1 U14878 ( .A(n15003), .B(n15004), .Z(n15001) );
  NOR2_X1 U14879 ( .A1(n8763), .A2(n8558), .ZN(n15004) );
  XOR2_X1 U14880 ( .A(n15005), .B(n15006), .Z(n14779) );
  XOR2_X1 U14881 ( .A(n15007), .B(n15008), .Z(n15005) );
  NOR2_X1 U14882 ( .A1(n8764), .A2(n8558), .ZN(n15008) );
  INV_X1 U14883 ( .A(n8670), .ZN(n14785) );
  NAND2_X1 U14884 ( .A1(b_5_), .A2(a_5_), .ZN(n8670) );
  XOR2_X1 U14885 ( .A(n15009), .B(n15010), .Z(n14787) );
  XOR2_X1 U14886 ( .A(n15011), .B(n15012), .Z(n15009) );
  NOR2_X1 U14887 ( .A1(n8517), .A2(n8558), .ZN(n15012) );
  XOR2_X1 U14888 ( .A(n15013), .B(n15014), .Z(n14791) );
  XOR2_X1 U14889 ( .A(n15015), .B(n15016), .Z(n15013) );
  XOR2_X1 U14890 ( .A(n15017), .B(n15018), .Z(n14795) );
  XOR2_X1 U14891 ( .A(n15019), .B(n15020), .Z(n15017) );
  NOR2_X1 U14892 ( .A1(n8567), .A2(n8558), .ZN(n15020) );
  XOR2_X1 U14893 ( .A(n15021), .B(n15022), .Z(n14799) );
  XOR2_X1 U14894 ( .A(n15023), .B(n15024), .Z(n15021) );
  NOR2_X1 U14895 ( .A1(n8768), .A2(n8558), .ZN(n15024) );
  XOR2_X1 U14896 ( .A(n15025), .B(n15026), .Z(n14808) );
  XOR2_X1 U14897 ( .A(n15027), .B(n15028), .Z(n15025) );
  NOR2_X1 U14898 ( .A1(n8617), .A2(n8558), .ZN(n15028) );
  XOR2_X1 U14899 ( .A(n14806), .B(n15029), .Z(n14814) );
  XNOR2_X1 U14900 ( .A(n15030), .B(n15031), .ZN(n14806) );
  NOR2_X1 U14901 ( .A1(n9674), .A2(n8558), .ZN(n15031) );
  NAND2_X1 U14902 ( .A1(n15032), .A2(n15033), .ZN(n8456) );
  NAND2_X1 U14903 ( .A1(n15034), .A2(n15035), .ZN(n15033) );
  NAND2_X1 U14904 ( .A1(n14813), .A2(n14812), .ZN(n15032) );
  NAND4_X1 U14905 ( .A1(n14813), .A2(n15034), .A3(n14812), .A4(n15035), .ZN(
        n8457) );
  NAND2_X1 U14906 ( .A1(n15036), .A2(n15037), .ZN(n14812) );
  NAND3_X1 U14907 ( .A1(a_0_), .A2(n15038), .A3(b_4_), .ZN(n15037) );
  OR2_X1 U14908 ( .A1(n14805), .A2(n15030), .ZN(n15038) );
  NAND2_X1 U14909 ( .A1(n14805), .A2(n15030), .ZN(n15036) );
  NAND2_X1 U14910 ( .A1(n15039), .A2(n15040), .ZN(n15030) );
  NAND3_X1 U14911 ( .A1(a_1_), .A2(n15041), .A3(b_4_), .ZN(n15040) );
  OR2_X1 U14912 ( .A1(n15027), .A2(n15026), .ZN(n15041) );
  NAND2_X1 U14913 ( .A1(n15026), .A2(n15027), .ZN(n15039) );
  NAND2_X1 U14914 ( .A1(n15042), .A2(n15043), .ZN(n15027) );
  NAND3_X1 U14915 ( .A1(a_2_), .A2(n15044), .A3(b_4_), .ZN(n15043) );
  OR2_X1 U14916 ( .A1(n15022), .A2(n15023), .ZN(n15044) );
  NAND2_X1 U14917 ( .A1(n15022), .A2(n15023), .ZN(n15042) );
  NAND2_X1 U14918 ( .A1(n15045), .A2(n15046), .ZN(n15023) );
  NAND3_X1 U14919 ( .A1(a_3_), .A2(n15047), .A3(b_4_), .ZN(n15046) );
  OR2_X1 U14920 ( .A1(n15019), .A2(n15018), .ZN(n15047) );
  NAND2_X1 U14921 ( .A1(n15018), .A2(n15019), .ZN(n15045) );
  NAND2_X1 U14922 ( .A1(n15048), .A2(n15049), .ZN(n15019) );
  NAND2_X1 U14923 ( .A1(n15014), .A2(n15050), .ZN(n15049) );
  OR2_X1 U14924 ( .A1(n15015), .A2(n15016), .ZN(n15050) );
  XNOR2_X1 U14925 ( .A(n15051), .B(n15052), .ZN(n15014) );
  NAND2_X1 U14926 ( .A1(n15053), .A2(n15054), .ZN(n15051) );
  NAND2_X1 U14927 ( .A1(n15016), .A2(n15015), .ZN(n15048) );
  NAND2_X1 U14928 ( .A1(n15055), .A2(n15056), .ZN(n15015) );
  NAND3_X1 U14929 ( .A1(a_5_), .A2(n15057), .A3(b_4_), .ZN(n15056) );
  OR2_X1 U14930 ( .A1(n15011), .A2(n15010), .ZN(n15057) );
  NAND2_X1 U14931 ( .A1(n15010), .A2(n15011), .ZN(n15055) );
  NAND2_X1 U14932 ( .A1(n15058), .A2(n15059), .ZN(n15011) );
  NAND3_X1 U14933 ( .A1(a_6_), .A2(n15060), .A3(b_4_), .ZN(n15059) );
  NAND2_X1 U14934 ( .A1(n14834), .A2(n14833), .ZN(n15060) );
  OR2_X1 U14935 ( .A1(n14833), .A2(n14834), .ZN(n15058) );
  AND2_X1 U14936 ( .A1(n15061), .A2(n15062), .ZN(n14834) );
  NAND3_X1 U14937 ( .A1(a_7_), .A2(n15063), .A3(b_4_), .ZN(n15062) );
  OR2_X1 U14938 ( .A1(n15007), .A2(n15006), .ZN(n15063) );
  NAND2_X1 U14939 ( .A1(n15006), .A2(n15007), .ZN(n15061) );
  NAND2_X1 U14940 ( .A1(n15064), .A2(n15065), .ZN(n15007) );
  NAND3_X1 U14941 ( .A1(a_8_), .A2(n15066), .A3(b_4_), .ZN(n15065) );
  OR2_X1 U14942 ( .A1(n15003), .A2(n15002), .ZN(n15066) );
  NAND2_X1 U14943 ( .A1(n15002), .A2(n15003), .ZN(n15064) );
  NAND2_X1 U14944 ( .A1(n15067), .A2(n15068), .ZN(n15003) );
  NAND3_X1 U14945 ( .A1(a_9_), .A2(n15069), .A3(b_4_), .ZN(n15068) );
  NAND2_X1 U14946 ( .A1(n14999), .A2(n14997), .ZN(n15069) );
  OR2_X1 U14947 ( .A1(n14997), .A2(n14999), .ZN(n15067) );
  AND2_X1 U14948 ( .A1(n15070), .A2(n15071), .ZN(n14999) );
  NAND3_X1 U14949 ( .A1(a_10_), .A2(n15072), .A3(b_4_), .ZN(n15071) );
  NAND2_X1 U14950 ( .A1(n14995), .A2(n14993), .ZN(n15072) );
  OR2_X1 U14951 ( .A1(n14993), .A2(n14995), .ZN(n15070) );
  AND2_X1 U14952 ( .A1(n15073), .A2(n15074), .ZN(n14995) );
  NAND3_X1 U14953 ( .A1(a_11_), .A2(n15075), .A3(b_4_), .ZN(n15074) );
  NAND2_X1 U14954 ( .A1(n14991), .A2(n14989), .ZN(n15075) );
  OR2_X1 U14955 ( .A1(n14989), .A2(n14991), .ZN(n15073) );
  AND2_X1 U14956 ( .A1(n15076), .A2(n15077), .ZN(n14991) );
  NAND3_X1 U14957 ( .A1(a_12_), .A2(n15078), .A3(b_4_), .ZN(n15077) );
  NAND2_X1 U14958 ( .A1(n14987), .A2(n14986), .ZN(n15078) );
  OR2_X1 U14959 ( .A1(n14986), .A2(n14987), .ZN(n15076) );
  AND2_X1 U14960 ( .A1(n15079), .A2(n15080), .ZN(n14987) );
  NAND3_X1 U14961 ( .A1(a_13_), .A2(n15081), .A3(b_4_), .ZN(n15080) );
  NAND2_X1 U14962 ( .A1(n14983), .A2(n14982), .ZN(n15081) );
  OR2_X1 U14963 ( .A1(n14982), .A2(n14983), .ZN(n15079) );
  AND2_X1 U14964 ( .A1(n15082), .A2(n15083), .ZN(n14983) );
  NAND2_X1 U14965 ( .A1(n14980), .A2(n15084), .ZN(n15083) );
  NAND2_X1 U14966 ( .A1(n14979), .A2(n14978), .ZN(n15084) );
  NOR2_X1 U14967 ( .A1(n8558), .A2(n8757), .ZN(n14980) );
  OR2_X1 U14968 ( .A1(n14978), .A2(n14979), .ZN(n15082) );
  AND2_X1 U14969 ( .A1(n15085), .A2(n15086), .ZN(n14979) );
  NAND2_X1 U14970 ( .A1(n14976), .A2(n15087), .ZN(n15086) );
  NAND2_X1 U14971 ( .A1(n14975), .A2(n14974), .ZN(n15087) );
  NOR2_X1 U14972 ( .A1(n8558), .A2(n8276), .ZN(n14976) );
  OR2_X1 U14973 ( .A1(n14974), .A2(n14975), .ZN(n15085) );
  AND2_X1 U14974 ( .A1(n15088), .A2(n15089), .ZN(n14975) );
  NAND2_X1 U14975 ( .A1(n14972), .A2(n15090), .ZN(n15089) );
  OR2_X1 U14976 ( .A1(n14970), .A2(n14971), .ZN(n15090) );
  NOR2_X1 U14977 ( .A1(n8558), .A2(n8755), .ZN(n14972) );
  NAND2_X1 U14978 ( .A1(n14970), .A2(n14971), .ZN(n15088) );
  NAND2_X1 U14979 ( .A1(n15091), .A2(n15092), .ZN(n14971) );
  NAND2_X1 U14980 ( .A1(n14968), .A2(n15093), .ZN(n15092) );
  NAND2_X1 U14981 ( .A1(n14967), .A2(n14966), .ZN(n15093) );
  NOR2_X1 U14982 ( .A1(n8558), .A2(n8210), .ZN(n14968) );
  OR2_X1 U14983 ( .A1(n14966), .A2(n14967), .ZN(n15091) );
  AND2_X1 U14984 ( .A1(n15094), .A2(n15095), .ZN(n14967) );
  NAND2_X1 U14985 ( .A1(n14964), .A2(n15096), .ZN(n15095) );
  OR2_X1 U14986 ( .A1(n14962), .A2(n14963), .ZN(n15096) );
  NOR2_X1 U14987 ( .A1(n8558), .A2(n8753), .ZN(n14964) );
  NAND2_X1 U14988 ( .A1(n14962), .A2(n14963), .ZN(n15094) );
  NAND2_X1 U14989 ( .A1(n15097), .A2(n15098), .ZN(n14963) );
  NAND2_X1 U14990 ( .A1(n14959), .A2(n15099), .ZN(n15098) );
  NAND2_X1 U14991 ( .A1(n14960), .A2(n14958), .ZN(n15099) );
  NOR2_X1 U14992 ( .A1(n8558), .A2(n8170), .ZN(n14959) );
  OR2_X1 U14993 ( .A1(n14958), .A2(n14960), .ZN(n15097) );
  AND2_X1 U14994 ( .A1(n15100), .A2(n15101), .ZN(n14960) );
  NAND2_X1 U14995 ( .A1(n14956), .A2(n15102), .ZN(n15101) );
  OR2_X1 U14996 ( .A1(n14954), .A2(n14955), .ZN(n15102) );
  NOR2_X1 U14997 ( .A1(n8558), .A2(n8751), .ZN(n14956) );
  NAND2_X1 U14998 ( .A1(n14954), .A2(n14955), .ZN(n15100) );
  NAND2_X1 U14999 ( .A1(n15103), .A2(n15104), .ZN(n14955) );
  NAND2_X1 U15000 ( .A1(n14951), .A2(n15105), .ZN(n15104) );
  NAND2_X1 U15001 ( .A1(n14952), .A2(n14950), .ZN(n15105) );
  NOR2_X1 U15002 ( .A1(n8558), .A2(n8750), .ZN(n14951) );
  OR2_X1 U15003 ( .A1(n14950), .A2(n14952), .ZN(n15103) );
  AND2_X1 U15004 ( .A1(n15106), .A2(n15107), .ZN(n14952) );
  NAND2_X1 U15005 ( .A1(n14948), .A2(n15108), .ZN(n15107) );
  OR2_X1 U15006 ( .A1(n14945), .A2(n14947), .ZN(n15108) );
  NOR2_X1 U15007 ( .A1(n8558), .A2(n8748), .ZN(n14948) );
  NAND2_X1 U15008 ( .A1(n14945), .A2(n14947), .ZN(n15106) );
  NAND2_X1 U15009 ( .A1(n15109), .A2(n15110), .ZN(n14947) );
  NAND2_X1 U15010 ( .A1(n14944), .A2(n15111), .ZN(n15110) );
  OR2_X1 U15011 ( .A1(n14942), .A2(n14943), .ZN(n15111) );
  NOR2_X1 U15012 ( .A1(n8558), .A2(n8747), .ZN(n14944) );
  NAND2_X1 U15013 ( .A1(n14942), .A2(n14943), .ZN(n15109) );
  NAND2_X1 U15014 ( .A1(n15112), .A2(n15113), .ZN(n14943) );
  NAND2_X1 U15015 ( .A1(n14940), .A2(n15114), .ZN(n15113) );
  OR2_X1 U15016 ( .A1(n14938), .A2(n14939), .ZN(n15114) );
  NOR2_X1 U15017 ( .A1(n8558), .A2(n8745), .ZN(n14940) );
  NAND2_X1 U15018 ( .A1(n14938), .A2(n14939), .ZN(n15112) );
  NAND2_X1 U15019 ( .A1(n15115), .A2(n15116), .ZN(n14939) );
  NAND2_X1 U15020 ( .A1(n14936), .A2(n15117), .ZN(n15116) );
  OR2_X1 U15021 ( .A1(n14934), .A2(n14935), .ZN(n15117) );
  NOR2_X1 U15022 ( .A1(n8558), .A2(n8744), .ZN(n14936) );
  NAND2_X1 U15023 ( .A1(n14934), .A2(n14935), .ZN(n15115) );
  NAND2_X1 U15024 ( .A1(n14899), .A2(n15118), .ZN(n14935) );
  NAND2_X1 U15025 ( .A1(n14898), .A2(n14900), .ZN(n15118) );
  NAND2_X1 U15026 ( .A1(n15119), .A2(n15120), .ZN(n14900) );
  NAND2_X1 U15027 ( .A1(b_4_), .A2(a_26_), .ZN(n15120) );
  INV_X1 U15028 ( .A(n15121), .ZN(n15119) );
  XNOR2_X1 U15029 ( .A(n15122), .B(n15123), .ZN(n14898) );
  NAND2_X1 U15030 ( .A1(n15124), .A2(n15125), .ZN(n15122) );
  NAND2_X1 U15031 ( .A1(a_26_), .A2(n15121), .ZN(n14899) );
  NAND2_X1 U15032 ( .A1(n14907), .A2(n15126), .ZN(n15121) );
  NAND2_X1 U15033 ( .A1(n14906), .A2(n14908), .ZN(n15126) );
  NAND2_X1 U15034 ( .A1(n15127), .A2(n15128), .ZN(n14908) );
  NAND2_X1 U15035 ( .A1(b_4_), .A2(a_27_), .ZN(n15128) );
  INV_X1 U15036 ( .A(n15129), .ZN(n15127) );
  XNOR2_X1 U15037 ( .A(n15130), .B(n15131), .ZN(n14906) );
  XOR2_X1 U15038 ( .A(n15132), .B(n15133), .Z(n15130) );
  NAND2_X1 U15039 ( .A1(b_3_), .A2(a_28_), .ZN(n15132) );
  NAND2_X1 U15040 ( .A1(a_27_), .A2(n15129), .ZN(n14907) );
  NAND2_X1 U15041 ( .A1(n15134), .A2(n15135), .ZN(n15129) );
  NAND3_X1 U15042 ( .A1(a_28_), .A2(n15136), .A3(b_4_), .ZN(n15135) );
  NAND2_X1 U15043 ( .A1(n14916), .A2(n14914), .ZN(n15136) );
  OR2_X1 U15044 ( .A1(n14914), .A2(n14916), .ZN(n15134) );
  AND2_X1 U15045 ( .A1(n15137), .A2(n15138), .ZN(n14916) );
  NAND2_X1 U15046 ( .A1(n14930), .A2(n15139), .ZN(n15138) );
  OR2_X1 U15047 ( .A1(n14931), .A2(n14932), .ZN(n15139) );
  NOR2_X1 U15048 ( .A1(n8558), .A2(n7890), .ZN(n14930) );
  NAND2_X1 U15049 ( .A1(n14932), .A2(n14931), .ZN(n15137) );
  NAND2_X1 U15050 ( .A1(n15140), .A2(n15141), .ZN(n14931) );
  NAND2_X1 U15051 ( .A1(b_2_), .A2(n15142), .ZN(n15141) );
  NAND2_X1 U15052 ( .A1(n7864), .A2(n15143), .ZN(n15142) );
  NAND2_X1 U15053 ( .A1(a_31_), .A2(n8767), .ZN(n15143) );
  NAND2_X1 U15054 ( .A1(b_3_), .A2(n15144), .ZN(n15140) );
  NAND2_X1 U15055 ( .A1(n9137), .A2(n15145), .ZN(n15144) );
  NAND2_X1 U15056 ( .A1(a_30_), .A2(n8608), .ZN(n15145) );
  AND3_X1 U15057 ( .A1(b_3_), .A2(b_4_), .A3(n7818), .ZN(n14932) );
  XNOR2_X1 U15058 ( .A(n15146), .B(n15147), .ZN(n14914) );
  XOR2_X1 U15059 ( .A(n15148), .B(n15149), .Z(n15146) );
  XNOR2_X1 U15060 ( .A(n15150), .B(n15151), .ZN(n14934) );
  NAND2_X1 U15061 ( .A1(n15152), .A2(n15153), .ZN(n15150) );
  XNOR2_X1 U15062 ( .A(n15154), .B(n15155), .ZN(n14938) );
  NAND2_X1 U15063 ( .A1(n15156), .A2(n15157), .ZN(n15154) );
  XNOR2_X1 U15064 ( .A(n15158), .B(n15159), .ZN(n14942) );
  XNOR2_X1 U15065 ( .A(n15160), .B(n15161), .ZN(n15158) );
  NOR2_X1 U15066 ( .A1(n8745), .A2(n8767), .ZN(n15161) );
  XNOR2_X1 U15067 ( .A(n15162), .B(n15163), .ZN(n14945) );
  NAND2_X1 U15068 ( .A1(n15164), .A2(n15165), .ZN(n15162) );
  XNOR2_X1 U15069 ( .A(n15166), .B(n15167), .ZN(n14950) );
  XNOR2_X1 U15070 ( .A(n15168), .B(n15169), .ZN(n15166) );
  NAND2_X1 U15071 ( .A1(b_3_), .A2(a_22_), .ZN(n15168) );
  XNOR2_X1 U15072 ( .A(n15170), .B(n15171), .ZN(n14954) );
  NAND2_X1 U15073 ( .A1(n15172), .A2(n15173), .ZN(n15170) );
  XNOR2_X1 U15074 ( .A(n15174), .B(n15175), .ZN(n14958) );
  XNOR2_X1 U15075 ( .A(n15176), .B(n15177), .ZN(n15174) );
  NAND2_X1 U15076 ( .A1(b_3_), .A2(a_20_), .ZN(n15176) );
  XNOR2_X1 U15077 ( .A(n15178), .B(n15179), .ZN(n14962) );
  NAND2_X1 U15078 ( .A1(n15180), .A2(n15181), .ZN(n15178) );
  XNOR2_X1 U15079 ( .A(n15182), .B(n15183), .ZN(n14966) );
  XNOR2_X1 U15080 ( .A(n15184), .B(n15185), .ZN(n15182) );
  NAND2_X1 U15081 ( .A1(b_3_), .A2(a_18_), .ZN(n15184) );
  XNOR2_X1 U15082 ( .A(n15186), .B(n15187), .ZN(n14970) );
  NAND2_X1 U15083 ( .A1(n15188), .A2(n15189), .ZN(n15186) );
  XNOR2_X1 U15084 ( .A(n15190), .B(n15191), .ZN(n14974) );
  XNOR2_X1 U15085 ( .A(n15192), .B(n15193), .ZN(n15190) );
  NAND2_X1 U15086 ( .A1(b_3_), .A2(a_16_), .ZN(n15192) );
  XOR2_X1 U15087 ( .A(n15194), .B(n15195), .Z(n14978) );
  NAND2_X1 U15088 ( .A1(n15196), .A2(n15197), .ZN(n15194) );
  XNOR2_X1 U15089 ( .A(n15198), .B(n15199), .ZN(n14982) );
  XNOR2_X1 U15090 ( .A(n15200), .B(n15201), .ZN(n15198) );
  NAND2_X1 U15091 ( .A1(b_3_), .A2(a_14_), .ZN(n15200) );
  XOR2_X1 U15092 ( .A(n15202), .B(n15203), .Z(n14986) );
  NAND2_X1 U15093 ( .A1(n15204), .A2(n15205), .ZN(n15202) );
  XNOR2_X1 U15094 ( .A(n15206), .B(n15207), .ZN(n14989) );
  XNOR2_X1 U15095 ( .A(n15208), .B(n15209), .ZN(n15206) );
  NAND2_X1 U15096 ( .A1(b_3_), .A2(a_12_), .ZN(n15208) );
  XOR2_X1 U15097 ( .A(n15210), .B(n15211), .Z(n14993) );
  NAND2_X1 U15098 ( .A1(n15212), .A2(n15213), .ZN(n15210) );
  XNOR2_X1 U15099 ( .A(n15214), .B(n15215), .ZN(n14997) );
  XNOR2_X1 U15100 ( .A(n15216), .B(n15217), .ZN(n15214) );
  NAND2_X1 U15101 ( .A1(b_3_), .A2(a_10_), .ZN(n15216) );
  XNOR2_X1 U15102 ( .A(n15218), .B(n15219), .ZN(n15002) );
  NAND2_X1 U15103 ( .A1(n15220), .A2(n15221), .ZN(n15218) );
  XOR2_X1 U15104 ( .A(n15222), .B(n15223), .Z(n15006) );
  XNOR2_X1 U15105 ( .A(n15224), .B(n15225), .ZN(n15222) );
  NAND2_X1 U15106 ( .A1(b_3_), .A2(a_8_), .ZN(n15224) );
  XOR2_X1 U15107 ( .A(n15226), .B(n15227), .Z(n14833) );
  NAND2_X1 U15108 ( .A1(n15228), .A2(n15229), .ZN(n15226) );
  XOR2_X1 U15109 ( .A(n15230), .B(n15231), .Z(n15010) );
  XNOR2_X1 U15110 ( .A(n15232), .B(n15233), .ZN(n15230) );
  NAND2_X1 U15111 ( .A1(b_3_), .A2(a_6_), .ZN(n15232) );
  INV_X1 U15112 ( .A(n8667), .ZN(n15016) );
  NAND2_X1 U15113 ( .A1(b_4_), .A2(a_4_), .ZN(n8667) );
  XOR2_X1 U15114 ( .A(n15234), .B(n15235), .Z(n15018) );
  XNOR2_X1 U15115 ( .A(n15236), .B(n15237), .ZN(n15234) );
  NAND2_X1 U15116 ( .A1(b_3_), .A2(a_4_), .ZN(n15236) );
  XOR2_X1 U15117 ( .A(n15238), .B(n15239), .Z(n15022) );
  XOR2_X1 U15118 ( .A(n15240), .B(n15241), .Z(n15238) );
  XOR2_X1 U15119 ( .A(n15242), .B(n15243), .Z(n15026) );
  XNOR2_X1 U15120 ( .A(n15244), .B(n15245), .ZN(n15242) );
  NAND2_X1 U15121 ( .A1(b_3_), .A2(a_2_), .ZN(n15244) );
  INV_X1 U15122 ( .A(n15029), .ZN(n14805) );
  XOR2_X1 U15123 ( .A(n15246), .B(n15247), .Z(n15029) );
  NAND2_X1 U15124 ( .A1(n15248), .A2(n15249), .ZN(n15246) );
  NAND2_X1 U15125 ( .A1(n15250), .A2(n15251), .ZN(n15034) );
  XOR2_X1 U15126 ( .A(n15252), .B(n15253), .Z(n14813) );
  XOR2_X1 U15127 ( .A(n15254), .B(n15255), .Z(n15252) );
  NAND2_X1 U15128 ( .A1(n15256), .A2(n15035), .ZN(n8786) );
  INV_X1 U15129 ( .A(n15257), .ZN(n15035) );
  XNOR2_X1 U15130 ( .A(n8920), .B(n8921), .ZN(n15256) );
  NAND2_X1 U15131 ( .A1(n15257), .A2(n15258), .ZN(n8787) );
  XOR2_X1 U15132 ( .A(n8921), .B(n8920), .Z(n15258) );
  NOR2_X1 U15133 ( .A1(n15251), .A2(n15250), .ZN(n15257) );
  AND2_X1 U15134 ( .A1(n15259), .A2(n15260), .ZN(n15250) );
  NAND2_X1 U15135 ( .A1(n15254), .A2(n15261), .ZN(n15260) );
  OR2_X1 U15136 ( .A1(n15253), .A2(n15255), .ZN(n15261) );
  NOR2_X1 U15137 ( .A1(n8767), .A2(n9674), .ZN(n15254) );
  NAND2_X1 U15138 ( .A1(n15253), .A2(n15255), .ZN(n15259) );
  NAND2_X1 U15139 ( .A1(n15248), .A2(n15262), .ZN(n15255) );
  NAND2_X1 U15140 ( .A1(n15247), .A2(n15249), .ZN(n15262) );
  NAND2_X1 U15141 ( .A1(n15263), .A2(n15264), .ZN(n15249) );
  NAND2_X1 U15142 ( .A1(b_3_), .A2(a_1_), .ZN(n15264) );
  INV_X1 U15143 ( .A(n15265), .ZN(n15263) );
  XNOR2_X1 U15144 ( .A(n15266), .B(n15267), .ZN(n15247) );
  XNOR2_X1 U15145 ( .A(n15268), .B(n8661), .ZN(n15267) );
  NAND2_X1 U15146 ( .A1(a_1_), .A2(n15265), .ZN(n15248) );
  NAND2_X1 U15147 ( .A1(n15269), .A2(n15270), .ZN(n15265) );
  NAND3_X1 U15148 ( .A1(a_2_), .A2(n15271), .A3(b_3_), .ZN(n15270) );
  OR2_X1 U15149 ( .A1(n15243), .A2(n15245), .ZN(n15271) );
  NAND2_X1 U15150 ( .A1(n15243), .A2(n15245), .ZN(n15269) );
  NAND2_X1 U15151 ( .A1(n15272), .A2(n15273), .ZN(n15245) );
  NAND2_X1 U15152 ( .A1(n15239), .A2(n15274), .ZN(n15273) );
  OR2_X1 U15153 ( .A1(n15240), .A2(n15241), .ZN(n15274) );
  XNOR2_X1 U15154 ( .A(n15275), .B(n15276), .ZN(n15239) );
  NAND2_X1 U15155 ( .A1(n15277), .A2(n15278), .ZN(n15275) );
  NAND2_X1 U15156 ( .A1(n15241), .A2(n15240), .ZN(n15272) );
  NAND2_X1 U15157 ( .A1(n15279), .A2(n15280), .ZN(n15240) );
  NAND3_X1 U15158 ( .A1(a_4_), .A2(n15281), .A3(b_3_), .ZN(n15280) );
  OR2_X1 U15159 ( .A1(n15235), .A2(n15237), .ZN(n15281) );
  NAND2_X1 U15160 ( .A1(n15235), .A2(n15237), .ZN(n15279) );
  NAND2_X1 U15161 ( .A1(n15053), .A2(n15282), .ZN(n15237) );
  NAND2_X1 U15162 ( .A1(n15052), .A2(n15054), .ZN(n15282) );
  NAND2_X1 U15163 ( .A1(n15283), .A2(n15284), .ZN(n15054) );
  NAND2_X1 U15164 ( .A1(b_3_), .A2(a_5_), .ZN(n15284) );
  INV_X1 U15165 ( .A(n15285), .ZN(n15283) );
  XNOR2_X1 U15166 ( .A(n15286), .B(n15287), .ZN(n15052) );
  NAND2_X1 U15167 ( .A1(n15288), .A2(n15289), .ZN(n15286) );
  NAND2_X1 U15168 ( .A1(a_5_), .A2(n15285), .ZN(n15053) );
  NAND2_X1 U15169 ( .A1(n15290), .A2(n15291), .ZN(n15285) );
  NAND3_X1 U15170 ( .A1(a_6_), .A2(n15292), .A3(b_3_), .ZN(n15291) );
  OR2_X1 U15171 ( .A1(n15231), .A2(n15233), .ZN(n15292) );
  NAND2_X1 U15172 ( .A1(n15231), .A2(n15233), .ZN(n15290) );
  NAND2_X1 U15173 ( .A1(n15228), .A2(n15293), .ZN(n15233) );
  NAND2_X1 U15174 ( .A1(n15227), .A2(n15229), .ZN(n15293) );
  NAND2_X1 U15175 ( .A1(n15294), .A2(n15295), .ZN(n15229) );
  NAND2_X1 U15176 ( .A1(b_3_), .A2(a_7_), .ZN(n15295) );
  INV_X1 U15177 ( .A(n15296), .ZN(n15294) );
  XNOR2_X1 U15178 ( .A(n15297), .B(n15298), .ZN(n15227) );
  NAND2_X1 U15179 ( .A1(n15299), .A2(n15300), .ZN(n15297) );
  NAND2_X1 U15180 ( .A1(a_7_), .A2(n15296), .ZN(n15228) );
  NAND2_X1 U15181 ( .A1(n15301), .A2(n15302), .ZN(n15296) );
  NAND3_X1 U15182 ( .A1(a_8_), .A2(n15303), .A3(b_3_), .ZN(n15302) );
  OR2_X1 U15183 ( .A1(n15223), .A2(n15225), .ZN(n15303) );
  NAND2_X1 U15184 ( .A1(n15223), .A2(n15225), .ZN(n15301) );
  NAND2_X1 U15185 ( .A1(n15220), .A2(n15304), .ZN(n15225) );
  NAND2_X1 U15186 ( .A1(n15219), .A2(n15221), .ZN(n15304) );
  NAND2_X1 U15187 ( .A1(n15305), .A2(n15306), .ZN(n15221) );
  NAND2_X1 U15188 ( .A1(b_3_), .A2(a_9_), .ZN(n15306) );
  INV_X1 U15189 ( .A(n15307), .ZN(n15305) );
  XNOR2_X1 U15190 ( .A(n15308), .B(n15309), .ZN(n15219) );
  NAND2_X1 U15191 ( .A1(n15310), .A2(n15311), .ZN(n15308) );
  NAND2_X1 U15192 ( .A1(a_9_), .A2(n15307), .ZN(n15220) );
  NAND2_X1 U15193 ( .A1(n15312), .A2(n15313), .ZN(n15307) );
  NAND3_X1 U15194 ( .A1(a_10_), .A2(n15314), .A3(b_3_), .ZN(n15313) );
  OR2_X1 U15195 ( .A1(n15215), .A2(n15217), .ZN(n15314) );
  NAND2_X1 U15196 ( .A1(n15215), .A2(n15217), .ZN(n15312) );
  NAND2_X1 U15197 ( .A1(n15212), .A2(n15315), .ZN(n15217) );
  NAND2_X1 U15198 ( .A1(n15211), .A2(n15213), .ZN(n15315) );
  NAND2_X1 U15199 ( .A1(n15316), .A2(n15317), .ZN(n15213) );
  NAND2_X1 U15200 ( .A1(b_3_), .A2(a_11_), .ZN(n15317) );
  INV_X1 U15201 ( .A(n15318), .ZN(n15316) );
  XNOR2_X1 U15202 ( .A(n15319), .B(n15320), .ZN(n15211) );
  NAND2_X1 U15203 ( .A1(n15321), .A2(n15322), .ZN(n15319) );
  NAND2_X1 U15204 ( .A1(a_11_), .A2(n15318), .ZN(n15212) );
  NAND2_X1 U15205 ( .A1(n15323), .A2(n15324), .ZN(n15318) );
  NAND3_X1 U15206 ( .A1(a_12_), .A2(n15325), .A3(b_3_), .ZN(n15324) );
  OR2_X1 U15207 ( .A1(n15207), .A2(n15209), .ZN(n15325) );
  NAND2_X1 U15208 ( .A1(n15207), .A2(n15209), .ZN(n15323) );
  NAND2_X1 U15209 ( .A1(n15204), .A2(n15326), .ZN(n15209) );
  NAND2_X1 U15210 ( .A1(n15203), .A2(n15205), .ZN(n15326) );
  NAND2_X1 U15211 ( .A1(n15327), .A2(n15328), .ZN(n15205) );
  NAND2_X1 U15212 ( .A1(b_3_), .A2(a_13_), .ZN(n15328) );
  INV_X1 U15213 ( .A(n15329), .ZN(n15327) );
  XNOR2_X1 U15214 ( .A(n15330), .B(n15331), .ZN(n15203) );
  NAND2_X1 U15215 ( .A1(n15332), .A2(n15333), .ZN(n15330) );
  NAND2_X1 U15216 ( .A1(a_13_), .A2(n15329), .ZN(n15204) );
  NAND2_X1 U15217 ( .A1(n15334), .A2(n15335), .ZN(n15329) );
  NAND3_X1 U15218 ( .A1(a_14_), .A2(n15336), .A3(b_3_), .ZN(n15335) );
  OR2_X1 U15219 ( .A1(n15199), .A2(n15201), .ZN(n15336) );
  NAND2_X1 U15220 ( .A1(n15199), .A2(n15201), .ZN(n15334) );
  NAND2_X1 U15221 ( .A1(n15196), .A2(n15337), .ZN(n15201) );
  NAND2_X1 U15222 ( .A1(n15195), .A2(n15197), .ZN(n15337) );
  NAND2_X1 U15223 ( .A1(n15338), .A2(n15339), .ZN(n15197) );
  NAND2_X1 U15224 ( .A1(b_3_), .A2(a_15_), .ZN(n15339) );
  INV_X1 U15225 ( .A(n15340), .ZN(n15338) );
  XNOR2_X1 U15226 ( .A(n15341), .B(n15342), .ZN(n15195) );
  NAND2_X1 U15227 ( .A1(n15343), .A2(n15344), .ZN(n15341) );
  NAND2_X1 U15228 ( .A1(a_15_), .A2(n15340), .ZN(n15196) );
  NAND2_X1 U15229 ( .A1(n15345), .A2(n15346), .ZN(n15340) );
  NAND3_X1 U15230 ( .A1(a_16_), .A2(n15347), .A3(b_3_), .ZN(n15346) );
  OR2_X1 U15231 ( .A1(n15191), .A2(n15193), .ZN(n15347) );
  NAND2_X1 U15232 ( .A1(n15191), .A2(n15193), .ZN(n15345) );
  NAND2_X1 U15233 ( .A1(n15188), .A2(n15348), .ZN(n15193) );
  NAND2_X1 U15234 ( .A1(n15187), .A2(n15189), .ZN(n15348) );
  NAND2_X1 U15235 ( .A1(n15349), .A2(n15350), .ZN(n15189) );
  NAND2_X1 U15236 ( .A1(b_3_), .A2(a_17_), .ZN(n15350) );
  INV_X1 U15237 ( .A(n15351), .ZN(n15349) );
  XNOR2_X1 U15238 ( .A(n15352), .B(n15353), .ZN(n15187) );
  XNOR2_X1 U15239 ( .A(n15354), .B(n15355), .ZN(n15353) );
  NAND2_X1 U15240 ( .A1(a_17_), .A2(n15351), .ZN(n15188) );
  NAND2_X1 U15241 ( .A1(n15356), .A2(n15357), .ZN(n15351) );
  NAND3_X1 U15242 ( .A1(a_18_), .A2(n15358), .A3(b_3_), .ZN(n15357) );
  OR2_X1 U15243 ( .A1(n15183), .A2(n15185), .ZN(n15358) );
  NAND2_X1 U15244 ( .A1(n15183), .A2(n15185), .ZN(n15356) );
  NAND2_X1 U15245 ( .A1(n15180), .A2(n15359), .ZN(n15185) );
  NAND2_X1 U15246 ( .A1(n15179), .A2(n15181), .ZN(n15359) );
  NAND2_X1 U15247 ( .A1(n15360), .A2(n15361), .ZN(n15181) );
  NAND2_X1 U15248 ( .A1(b_3_), .A2(a_19_), .ZN(n15361) );
  INV_X1 U15249 ( .A(n15362), .ZN(n15360) );
  XNOR2_X1 U15250 ( .A(n15363), .B(n15364), .ZN(n15179) );
  XNOR2_X1 U15251 ( .A(n15365), .B(n15366), .ZN(n15364) );
  NAND2_X1 U15252 ( .A1(a_19_), .A2(n15362), .ZN(n15180) );
  NAND2_X1 U15253 ( .A1(n15367), .A2(n15368), .ZN(n15362) );
  NAND3_X1 U15254 ( .A1(a_20_), .A2(n15369), .A3(b_3_), .ZN(n15368) );
  OR2_X1 U15255 ( .A1(n15175), .A2(n15177), .ZN(n15369) );
  NAND2_X1 U15256 ( .A1(n15175), .A2(n15177), .ZN(n15367) );
  NAND2_X1 U15257 ( .A1(n15172), .A2(n15370), .ZN(n15177) );
  NAND2_X1 U15258 ( .A1(n15171), .A2(n15173), .ZN(n15370) );
  NAND2_X1 U15259 ( .A1(n15371), .A2(n15372), .ZN(n15173) );
  NAND2_X1 U15260 ( .A1(b_3_), .A2(a_21_), .ZN(n15372) );
  INV_X1 U15261 ( .A(n15373), .ZN(n15371) );
  XNOR2_X1 U15262 ( .A(n15374), .B(n15375), .ZN(n15171) );
  XNOR2_X1 U15263 ( .A(n15376), .B(n15377), .ZN(n15374) );
  NAND2_X1 U15264 ( .A1(a_21_), .A2(n15373), .ZN(n15172) );
  NAND2_X1 U15265 ( .A1(n15378), .A2(n15379), .ZN(n15373) );
  NAND3_X1 U15266 ( .A1(a_22_), .A2(n15380), .A3(b_3_), .ZN(n15379) );
  OR2_X1 U15267 ( .A1(n15167), .A2(n15169), .ZN(n15380) );
  NAND2_X1 U15268 ( .A1(n15167), .A2(n15169), .ZN(n15378) );
  NAND2_X1 U15269 ( .A1(n15164), .A2(n15381), .ZN(n15169) );
  NAND2_X1 U15270 ( .A1(n15163), .A2(n15165), .ZN(n15381) );
  NAND2_X1 U15271 ( .A1(n15382), .A2(n15383), .ZN(n15165) );
  NAND2_X1 U15272 ( .A1(b_3_), .A2(a_23_), .ZN(n15383) );
  INV_X1 U15273 ( .A(n15384), .ZN(n15382) );
  XNOR2_X1 U15274 ( .A(n15385), .B(n15386), .ZN(n15163) );
  XNOR2_X1 U15275 ( .A(n15387), .B(n15388), .ZN(n15386) );
  NAND2_X1 U15276 ( .A1(a_23_), .A2(n15384), .ZN(n15164) );
  NAND2_X1 U15277 ( .A1(n15389), .A2(n15390), .ZN(n15384) );
  NAND3_X1 U15278 ( .A1(a_24_), .A2(n15391), .A3(b_3_), .ZN(n15390) );
  NAND2_X1 U15279 ( .A1(n15160), .A2(n15159), .ZN(n15391) );
  OR2_X1 U15280 ( .A1(n15159), .A2(n15160), .ZN(n15389) );
  AND2_X1 U15281 ( .A1(n15156), .A2(n15392), .ZN(n15160) );
  NAND2_X1 U15282 ( .A1(n15155), .A2(n15157), .ZN(n15392) );
  NAND2_X1 U15283 ( .A1(n15393), .A2(n15394), .ZN(n15157) );
  NAND2_X1 U15284 ( .A1(b_3_), .A2(a_25_), .ZN(n15394) );
  INV_X1 U15285 ( .A(n15395), .ZN(n15393) );
  XNOR2_X1 U15286 ( .A(n15396), .B(n15397), .ZN(n15155) );
  XOR2_X1 U15287 ( .A(n15398), .B(n15399), .Z(n15396) );
  NAND2_X1 U15288 ( .A1(b_2_), .A2(a_26_), .ZN(n15398) );
  NAND2_X1 U15289 ( .A1(a_25_), .A2(n15395), .ZN(n15156) );
  NAND2_X1 U15290 ( .A1(n15152), .A2(n15400), .ZN(n15395) );
  NAND2_X1 U15291 ( .A1(n15151), .A2(n15153), .ZN(n15400) );
  NAND2_X1 U15292 ( .A1(n15401), .A2(n15402), .ZN(n15153) );
  NAND2_X1 U15293 ( .A1(b_3_), .A2(a_26_), .ZN(n15402) );
  INV_X1 U15294 ( .A(n15403), .ZN(n15401) );
  XNOR2_X1 U15295 ( .A(n15404), .B(n15405), .ZN(n15151) );
  XNOR2_X1 U15296 ( .A(n15406), .B(n15407), .ZN(n15405) );
  NAND2_X1 U15297 ( .A1(a_26_), .A2(n15403), .ZN(n15152) );
  NAND2_X1 U15298 ( .A1(n15124), .A2(n15408), .ZN(n15403) );
  NAND2_X1 U15299 ( .A1(n15123), .A2(n15125), .ZN(n15408) );
  NAND2_X1 U15300 ( .A1(n15409), .A2(n15410), .ZN(n15125) );
  NAND2_X1 U15301 ( .A1(b_3_), .A2(a_27_), .ZN(n15410) );
  INV_X1 U15302 ( .A(n15411), .ZN(n15409) );
  XOR2_X1 U15303 ( .A(n15412), .B(n15413), .Z(n15123) );
  XNOR2_X1 U15304 ( .A(n15414), .B(n15415), .ZN(n15412) );
  NAND2_X1 U15305 ( .A1(b_2_), .A2(a_28_), .ZN(n15414) );
  NAND2_X1 U15306 ( .A1(a_27_), .A2(n15411), .ZN(n15124) );
  NAND2_X1 U15307 ( .A1(n15416), .A2(n15417), .ZN(n15411) );
  NAND3_X1 U15308 ( .A1(a_28_), .A2(n15418), .A3(b_3_), .ZN(n15417) );
  NAND2_X1 U15309 ( .A1(n15133), .A2(n15131), .ZN(n15418) );
  OR2_X1 U15310 ( .A1(n15131), .A2(n15133), .ZN(n15416) );
  AND2_X1 U15311 ( .A1(n15419), .A2(n15420), .ZN(n15133) );
  NAND2_X1 U15312 ( .A1(n15147), .A2(n15421), .ZN(n15420) );
  OR2_X1 U15313 ( .A1(n15148), .A2(n15149), .ZN(n15421) );
  NOR2_X1 U15314 ( .A1(n8767), .A2(n7890), .ZN(n15147) );
  NAND2_X1 U15315 ( .A1(n15149), .A2(n15148), .ZN(n15419) );
  NAND2_X1 U15316 ( .A1(n15422), .A2(n15423), .ZN(n15148) );
  NAND2_X1 U15317 ( .A1(b_1_), .A2(n15424), .ZN(n15423) );
  NAND2_X1 U15318 ( .A1(n7864), .A2(n15425), .ZN(n15424) );
  NAND2_X1 U15319 ( .A1(a_31_), .A2(n8608), .ZN(n15425) );
  NAND2_X1 U15320 ( .A1(b_2_), .A2(n15426), .ZN(n15422) );
  NAND2_X1 U15321 ( .A1(n9137), .A2(n15427), .ZN(n15426) );
  NAND2_X1 U15322 ( .A1(a_30_), .A2(n8634), .ZN(n15427) );
  AND3_X1 U15323 ( .A1(b_2_), .A2(b_3_), .A3(n7818), .ZN(n15149) );
  XNOR2_X1 U15324 ( .A(n15428), .B(n15429), .ZN(n15131) );
  NOR2_X1 U15325 ( .A1(n7890), .A2(n8608), .ZN(n15429) );
  XOR2_X1 U15326 ( .A(n15430), .B(n15431), .Z(n15428) );
  XOR2_X1 U15327 ( .A(n15432), .B(n15433), .Z(n15159) );
  NAND2_X1 U15328 ( .A1(n15434), .A2(n15435), .ZN(n15432) );
  XNOR2_X1 U15329 ( .A(n15436), .B(n15437), .ZN(n15167) );
  XOR2_X1 U15330 ( .A(n15438), .B(n15439), .Z(n15437) );
  NAND2_X1 U15331 ( .A1(b_2_), .A2(a_23_), .ZN(n15439) );
  XNOR2_X1 U15332 ( .A(n15440), .B(n15441), .ZN(n15175) );
  XNOR2_X1 U15333 ( .A(n15442), .B(n15443), .ZN(n15440) );
  NOR2_X1 U15334 ( .A1(n8750), .A2(n8608), .ZN(n15443) );
  XNOR2_X1 U15335 ( .A(n15444), .B(n15445), .ZN(n15183) );
  XOR2_X1 U15336 ( .A(n15446), .B(n15447), .Z(n15444) );
  NAND2_X1 U15337 ( .A1(b_2_), .A2(a_19_), .ZN(n15446) );
  XNOR2_X1 U15338 ( .A(n15448), .B(n15449), .ZN(n15191) );
  XNOR2_X1 U15339 ( .A(n15450), .B(n15451), .ZN(n15448) );
  XOR2_X1 U15340 ( .A(n15452), .B(n15453), .Z(n15199) );
  XOR2_X1 U15341 ( .A(n15454), .B(n15455), .Z(n15452) );
  XOR2_X1 U15342 ( .A(n15456), .B(n15457), .Z(n15207) );
  XOR2_X1 U15343 ( .A(n15458), .B(n15459), .Z(n15456) );
  XOR2_X1 U15344 ( .A(n15460), .B(n15461), .Z(n15215) );
  XOR2_X1 U15345 ( .A(n15462), .B(n15463), .Z(n15460) );
  XOR2_X1 U15346 ( .A(n15464), .B(n15465), .Z(n15223) );
  XOR2_X1 U15347 ( .A(n15466), .B(n15467), .Z(n15464) );
  XOR2_X1 U15348 ( .A(n15468), .B(n15469), .Z(n15231) );
  XOR2_X1 U15349 ( .A(n15470), .B(n15471), .Z(n15468) );
  XOR2_X1 U15350 ( .A(n15472), .B(n15473), .Z(n15235) );
  XOR2_X1 U15351 ( .A(n15474), .B(n15475), .Z(n15472) );
  INV_X1 U15352 ( .A(n8664), .ZN(n15241) );
  NAND2_X1 U15353 ( .A1(b_3_), .A2(a_3_), .ZN(n8664) );
  XOR2_X1 U15354 ( .A(n15476), .B(n15477), .Z(n15243) );
  XOR2_X1 U15355 ( .A(n15478), .B(n15479), .Z(n15476) );
  XOR2_X1 U15356 ( .A(n15480), .B(n15481), .Z(n15253) );
  XOR2_X1 U15357 ( .A(n15482), .B(n15483), .Z(n15480) );
  XOR2_X1 U15358 ( .A(n15484), .B(n15485), .Z(n15251) );
  NAND2_X1 U15359 ( .A1(n15486), .A2(n15487), .ZN(n15484) );
  NAND2_X1 U15360 ( .A1(n15488), .A2(n15489), .ZN(n8851) );
  NAND2_X1 U15361 ( .A1(n8920), .A2(n8921), .ZN(n15489) );
  NAND2_X1 U15362 ( .A1(n15486), .A2(n15490), .ZN(n8921) );
  NAND2_X1 U15363 ( .A1(n15485), .A2(n15487), .ZN(n15490) );
  NAND2_X1 U15364 ( .A1(n15491), .A2(n15492), .ZN(n15487) );
  NAND2_X1 U15365 ( .A1(b_2_), .A2(a_0_), .ZN(n15492) );
  INV_X1 U15366 ( .A(n15493), .ZN(n15491) );
  XOR2_X1 U15367 ( .A(n15494), .B(n15495), .Z(n15485) );
  XNOR2_X1 U15368 ( .A(n8660), .B(n15496), .ZN(n15495) );
  NAND2_X1 U15369 ( .A1(b_0_), .A2(a_2_), .ZN(n15494) );
  NAND2_X1 U15370 ( .A1(a_0_), .A2(n15493), .ZN(n15486) );
  NAND2_X1 U15371 ( .A1(n15497), .A2(n15498), .ZN(n15493) );
  NAND2_X1 U15372 ( .A1(n15482), .A2(n15499), .ZN(n15498) );
  OR2_X1 U15373 ( .A1(n15483), .A2(n15481), .ZN(n15499) );
  NOR2_X1 U15374 ( .A1(n8608), .A2(n8617), .ZN(n15482) );
  NAND2_X1 U15375 ( .A1(n15481), .A2(n15483), .ZN(n15497) );
  NAND2_X1 U15376 ( .A1(n15500), .A2(n15501), .ZN(n15483) );
  NAND2_X1 U15377 ( .A1(n15266), .A2(n15502), .ZN(n15501) );
  NAND2_X1 U15378 ( .A1(n15268), .A2(n8661), .ZN(n15502) );
  XOR2_X1 U15379 ( .A(n15503), .B(n15504), .Z(n15266) );
  XNOR2_X1 U15380 ( .A(n15505), .B(n15506), .ZN(n15504) );
  NAND2_X1 U15381 ( .A1(b_1_), .A2(a_3_), .ZN(n15503) );
  OR2_X1 U15382 ( .A1(n8661), .A2(n15268), .ZN(n15500) );
  AND2_X1 U15383 ( .A1(n15507), .A2(n15508), .ZN(n15268) );
  NAND2_X1 U15384 ( .A1(n15478), .A2(n15509), .ZN(n15508) );
  OR2_X1 U15385 ( .A1(n15479), .A2(n15477), .ZN(n15509) );
  NOR2_X1 U15386 ( .A1(n8608), .A2(n8567), .ZN(n15478) );
  NAND2_X1 U15387 ( .A1(n15477), .A2(n15479), .ZN(n15507) );
  NAND2_X1 U15388 ( .A1(n15277), .A2(n15510), .ZN(n15479) );
  NAND2_X1 U15389 ( .A1(n15276), .A2(n15278), .ZN(n15510) );
  NAND2_X1 U15390 ( .A1(n15511), .A2(n15512), .ZN(n15278) );
  NAND2_X1 U15391 ( .A1(b_2_), .A2(a_4_), .ZN(n15512) );
  INV_X1 U15392 ( .A(n15513), .ZN(n15511) );
  XOR2_X1 U15393 ( .A(n15514), .B(n15515), .Z(n15276) );
  XNOR2_X1 U15394 ( .A(n15516), .B(n15517), .ZN(n15515) );
  NAND2_X1 U15395 ( .A1(b_1_), .A2(a_5_), .ZN(n15514) );
  NAND2_X1 U15396 ( .A1(a_4_), .A2(n15513), .ZN(n15277) );
  NAND2_X1 U15397 ( .A1(n15518), .A2(n15519), .ZN(n15513) );
  NAND2_X1 U15398 ( .A1(n15474), .A2(n15520), .ZN(n15519) );
  OR2_X1 U15399 ( .A1(n15475), .A2(n15473), .ZN(n15520) );
  NOR2_X1 U15400 ( .A1(n8608), .A2(n8517), .ZN(n15474) );
  NAND2_X1 U15401 ( .A1(n15473), .A2(n15475), .ZN(n15518) );
  NAND2_X1 U15402 ( .A1(n15288), .A2(n15521), .ZN(n15475) );
  NAND2_X1 U15403 ( .A1(n15287), .A2(n15289), .ZN(n15521) );
  NAND2_X1 U15404 ( .A1(n15522), .A2(n15523), .ZN(n15289) );
  NAND2_X1 U15405 ( .A1(b_2_), .A2(a_6_), .ZN(n15523) );
  INV_X1 U15406 ( .A(n15524), .ZN(n15522) );
  XOR2_X1 U15407 ( .A(n15525), .B(n15526), .Z(n15287) );
  XNOR2_X1 U15408 ( .A(n15527), .B(n15528), .ZN(n15526) );
  NAND2_X1 U15409 ( .A1(b_1_), .A2(a_7_), .ZN(n15525) );
  NAND2_X1 U15410 ( .A1(a_6_), .A2(n15524), .ZN(n15288) );
  NAND2_X1 U15411 ( .A1(n15529), .A2(n15530), .ZN(n15524) );
  NAND2_X1 U15412 ( .A1(n15470), .A2(n15531), .ZN(n15530) );
  OR2_X1 U15413 ( .A1(n15471), .A2(n15469), .ZN(n15531) );
  NOR2_X1 U15414 ( .A1(n8608), .A2(n8764), .ZN(n15470) );
  NAND2_X1 U15415 ( .A1(n15469), .A2(n15471), .ZN(n15529) );
  NAND2_X1 U15416 ( .A1(n15299), .A2(n15532), .ZN(n15471) );
  NAND2_X1 U15417 ( .A1(n15298), .A2(n15300), .ZN(n15532) );
  NAND2_X1 U15418 ( .A1(n15533), .A2(n15534), .ZN(n15300) );
  NAND2_X1 U15419 ( .A1(b_2_), .A2(a_8_), .ZN(n15534) );
  INV_X1 U15420 ( .A(n15535), .ZN(n15533) );
  XOR2_X1 U15421 ( .A(n15536), .B(n15537), .Z(n15298) );
  XNOR2_X1 U15422 ( .A(n15538), .B(n15539), .ZN(n15537) );
  NAND2_X1 U15423 ( .A1(b_1_), .A2(a_9_), .ZN(n15536) );
  NAND2_X1 U15424 ( .A1(a_8_), .A2(n15535), .ZN(n15299) );
  NAND2_X1 U15425 ( .A1(n15540), .A2(n15541), .ZN(n15535) );
  NAND2_X1 U15426 ( .A1(n15466), .A2(n15542), .ZN(n15541) );
  OR2_X1 U15427 ( .A1(n15467), .A2(n15465), .ZN(n15542) );
  NOR2_X1 U15428 ( .A1(n8608), .A2(n8426), .ZN(n15466) );
  NAND2_X1 U15429 ( .A1(n15465), .A2(n15467), .ZN(n15540) );
  NAND2_X1 U15430 ( .A1(n15310), .A2(n15543), .ZN(n15467) );
  NAND2_X1 U15431 ( .A1(n15309), .A2(n15311), .ZN(n15543) );
  NAND2_X1 U15432 ( .A1(n15544), .A2(n15545), .ZN(n15311) );
  NAND2_X1 U15433 ( .A1(b_2_), .A2(a_10_), .ZN(n15545) );
  INV_X1 U15434 ( .A(n15546), .ZN(n15544) );
  XOR2_X1 U15435 ( .A(n15547), .B(n15548), .Z(n15309) );
  XNOR2_X1 U15436 ( .A(n15549), .B(n15550), .ZN(n15548) );
  NAND2_X1 U15437 ( .A1(b_1_), .A2(a_11_), .ZN(n15547) );
  NAND2_X1 U15438 ( .A1(a_10_), .A2(n15546), .ZN(n15310) );
  NAND2_X1 U15439 ( .A1(n15551), .A2(n15552), .ZN(n15546) );
  NAND2_X1 U15440 ( .A1(n15462), .A2(n15553), .ZN(n15552) );
  OR2_X1 U15441 ( .A1(n15463), .A2(n15461), .ZN(n15553) );
  NOR2_X1 U15442 ( .A1(n8608), .A2(n8376), .ZN(n15462) );
  NAND2_X1 U15443 ( .A1(n15461), .A2(n15463), .ZN(n15551) );
  NAND2_X1 U15444 ( .A1(n15321), .A2(n15554), .ZN(n15463) );
  NAND2_X1 U15445 ( .A1(n15320), .A2(n15322), .ZN(n15554) );
  NAND2_X1 U15446 ( .A1(n15555), .A2(n15556), .ZN(n15322) );
  NAND2_X1 U15447 ( .A1(b_2_), .A2(a_12_), .ZN(n15556) );
  INV_X1 U15448 ( .A(n15557), .ZN(n15555) );
  XOR2_X1 U15449 ( .A(n15558), .B(n15559), .Z(n15320) );
  XNOR2_X1 U15450 ( .A(n15560), .B(n15561), .ZN(n15559) );
  NAND2_X1 U15451 ( .A1(b_1_), .A2(a_13_), .ZN(n15558) );
  NAND2_X1 U15452 ( .A1(a_12_), .A2(n15557), .ZN(n15321) );
  NAND2_X1 U15453 ( .A1(n15562), .A2(n15563), .ZN(n15557) );
  NAND2_X1 U15454 ( .A1(n15458), .A2(n15564), .ZN(n15563) );
  OR2_X1 U15455 ( .A1(n15459), .A2(n15457), .ZN(n15564) );
  NOR2_X1 U15456 ( .A1(n8608), .A2(n8310), .ZN(n15458) );
  NAND2_X1 U15457 ( .A1(n15457), .A2(n15459), .ZN(n15562) );
  NAND2_X1 U15458 ( .A1(n15332), .A2(n15565), .ZN(n15459) );
  NAND2_X1 U15459 ( .A1(n15331), .A2(n15333), .ZN(n15565) );
  NAND2_X1 U15460 ( .A1(n15566), .A2(n15567), .ZN(n15333) );
  NAND2_X1 U15461 ( .A1(b_2_), .A2(a_14_), .ZN(n15567) );
  INV_X1 U15462 ( .A(n15568), .ZN(n15566) );
  XOR2_X1 U15463 ( .A(n15569), .B(n15570), .Z(n15331) );
  XNOR2_X1 U15464 ( .A(n15571), .B(n15572), .ZN(n15570) );
  NAND2_X1 U15465 ( .A1(b_1_), .A2(a_15_), .ZN(n15569) );
  NAND2_X1 U15466 ( .A1(a_14_), .A2(n15568), .ZN(n15332) );
  NAND2_X1 U15467 ( .A1(n15573), .A2(n15574), .ZN(n15568) );
  NAND2_X1 U15468 ( .A1(n15454), .A2(n15575), .ZN(n15574) );
  OR2_X1 U15469 ( .A1(n15455), .A2(n15453), .ZN(n15575) );
  NOR2_X1 U15470 ( .A1(n8608), .A2(n8276), .ZN(n15454) );
  NAND2_X1 U15471 ( .A1(n15453), .A2(n15455), .ZN(n15573) );
  NAND2_X1 U15472 ( .A1(n15343), .A2(n15576), .ZN(n15455) );
  NAND2_X1 U15473 ( .A1(n15342), .A2(n15344), .ZN(n15576) );
  NAND2_X1 U15474 ( .A1(n15577), .A2(n15578), .ZN(n15344) );
  NAND2_X1 U15475 ( .A1(b_2_), .A2(a_16_), .ZN(n15578) );
  INV_X1 U15476 ( .A(n15579), .ZN(n15577) );
  XOR2_X1 U15477 ( .A(n15580), .B(n15581), .Z(n15342) );
  XNOR2_X1 U15478 ( .A(n15582), .B(n15583), .ZN(n15581) );
  NAND2_X1 U15479 ( .A1(b_1_), .A2(a_17_), .ZN(n15580) );
  NAND2_X1 U15480 ( .A1(a_16_), .A2(n15579), .ZN(n15343) );
  NAND2_X1 U15481 ( .A1(n15584), .A2(n15585), .ZN(n15579) );
  NAND2_X1 U15482 ( .A1(n15450), .A2(n15586), .ZN(n15585) );
  NAND2_X1 U15483 ( .A1(n15451), .A2(n15449), .ZN(n15586) );
  NOR2_X1 U15484 ( .A1(n8608), .A2(n8210), .ZN(n15450) );
  OR2_X1 U15485 ( .A1(n15449), .A2(n15451), .ZN(n15584) );
  AND2_X1 U15486 ( .A1(n15587), .A2(n15588), .ZN(n15451) );
  NAND2_X1 U15487 ( .A1(n15355), .A2(n15589), .ZN(n15588) );
  OR2_X1 U15488 ( .A1(n15354), .A2(n15352), .ZN(n15589) );
  NOR2_X1 U15489 ( .A1(n8608), .A2(n8753), .ZN(n15355) );
  NAND2_X1 U15490 ( .A1(n15352), .A2(n15354), .ZN(n15587) );
  NAND2_X1 U15491 ( .A1(n15590), .A2(n15591), .ZN(n15354) );
  NAND3_X1 U15492 ( .A1(a_19_), .A2(n15592), .A3(b_2_), .ZN(n15591) );
  NAND2_X1 U15493 ( .A1(n15447), .A2(n15445), .ZN(n15592) );
  OR2_X1 U15494 ( .A1(n15445), .A2(n15447), .ZN(n15590) );
  AND2_X1 U15495 ( .A1(n15593), .A2(n15594), .ZN(n15447) );
  NAND2_X1 U15496 ( .A1(n15366), .A2(n15595), .ZN(n15594) );
  OR2_X1 U15497 ( .A1(n15365), .A2(n15363), .ZN(n15595) );
  NOR2_X1 U15498 ( .A1(n8608), .A2(n8751), .ZN(n15366) );
  NAND2_X1 U15499 ( .A1(n15363), .A2(n15365), .ZN(n15593) );
  NAND2_X1 U15500 ( .A1(n15596), .A2(n15597), .ZN(n15365) );
  NAND3_X1 U15501 ( .A1(a_21_), .A2(n15598), .A3(b_2_), .ZN(n15597) );
  NAND2_X1 U15502 ( .A1(n15442), .A2(n15441), .ZN(n15598) );
  OR2_X1 U15503 ( .A1(n15441), .A2(n15442), .ZN(n15596) );
  AND2_X1 U15504 ( .A1(n15599), .A2(n15600), .ZN(n15442) );
  NAND2_X1 U15505 ( .A1(n15377), .A2(n15601), .ZN(n15600) );
  NAND2_X1 U15506 ( .A1(n15376), .A2(n15375), .ZN(n15601) );
  NOR2_X1 U15507 ( .A1(n8608), .A2(n8748), .ZN(n15377) );
  OR2_X1 U15508 ( .A1(n15375), .A2(n15376), .ZN(n15599) );
  AND2_X1 U15509 ( .A1(n15602), .A2(n15603), .ZN(n15376) );
  NAND3_X1 U15510 ( .A1(a_23_), .A2(n15604), .A3(b_2_), .ZN(n15603) );
  OR2_X1 U15511 ( .A1(n15438), .A2(n15436), .ZN(n15604) );
  NAND2_X1 U15512 ( .A1(n15436), .A2(n15438), .ZN(n15602) );
  NAND2_X1 U15513 ( .A1(n15605), .A2(n15606), .ZN(n15438) );
  NAND2_X1 U15514 ( .A1(n15388), .A2(n15607), .ZN(n15606) );
  OR2_X1 U15515 ( .A1(n15387), .A2(n15385), .ZN(n15607) );
  NOR2_X1 U15516 ( .A1(n8608), .A2(n8745), .ZN(n15388) );
  NAND2_X1 U15517 ( .A1(n15385), .A2(n15387), .ZN(n15605) );
  NAND2_X1 U15518 ( .A1(n15434), .A2(n15608), .ZN(n15387) );
  NAND2_X1 U15519 ( .A1(n15433), .A2(n15435), .ZN(n15608) );
  NAND2_X1 U15520 ( .A1(n15609), .A2(n15610), .ZN(n15435) );
  NAND2_X1 U15521 ( .A1(b_2_), .A2(a_25_), .ZN(n15610) );
  INV_X1 U15522 ( .A(n15611), .ZN(n15609) );
  XOR2_X1 U15523 ( .A(n15612), .B(n15613), .Z(n15433) );
  NOR2_X1 U15524 ( .A1(n8741), .A2(n8770), .ZN(n15613) );
  XOR2_X1 U15525 ( .A(n15614), .B(n15615), .Z(n15612) );
  NAND2_X1 U15526 ( .A1(a_25_), .A2(n15611), .ZN(n15434) );
  NAND2_X1 U15527 ( .A1(n15616), .A2(n15617), .ZN(n15611) );
  NAND3_X1 U15528 ( .A1(a_26_), .A2(n15618), .A3(b_2_), .ZN(n15617) );
  NAND2_X1 U15529 ( .A1(n15399), .A2(n15397), .ZN(n15618) );
  OR2_X1 U15530 ( .A1(n15397), .A2(n15399), .ZN(n15616) );
  AND2_X1 U15531 ( .A1(n15619), .A2(n15620), .ZN(n15399) );
  NAND2_X1 U15532 ( .A1(n15407), .A2(n15621), .ZN(n15620) );
  OR2_X1 U15533 ( .A1(n15406), .A2(n15404), .ZN(n15621) );
  NOR2_X1 U15534 ( .A1(n8608), .A2(n8741), .ZN(n15407) );
  NAND2_X1 U15535 ( .A1(n15404), .A2(n15406), .ZN(n15619) );
  NAND2_X1 U15536 ( .A1(n15622), .A2(n15623), .ZN(n15406) );
  NAND3_X1 U15537 ( .A1(a_28_), .A2(n15624), .A3(b_2_), .ZN(n15623) );
  OR2_X1 U15538 ( .A1(n15413), .A2(n15415), .ZN(n15624) );
  NAND2_X1 U15539 ( .A1(n15413), .A2(n15415), .ZN(n15622) );
  NAND2_X1 U15540 ( .A1(n15625), .A2(n15626), .ZN(n15415) );
  NAND3_X1 U15541 ( .A1(a_29_), .A2(n15627), .A3(b_2_), .ZN(n15626) );
  OR2_X1 U15542 ( .A1(n15430), .A2(n15431), .ZN(n15627) );
  NAND2_X1 U15543 ( .A1(n15431), .A2(n15430), .ZN(n15625) );
  NAND2_X1 U15544 ( .A1(n15628), .A2(n15629), .ZN(n15430) );
  NAND2_X1 U15545 ( .A1(b_0_), .A2(n15630), .ZN(n15629) );
  NAND2_X1 U15546 ( .A1(n7864), .A2(n15631), .ZN(n15630) );
  NAND2_X1 U15547 ( .A1(a_31_), .A2(n8634), .ZN(n15631) );
  NAND2_X1 U15548 ( .A1(b_1_), .A2(n15632), .ZN(n15628) );
  NAND2_X1 U15549 ( .A1(n9137), .A2(n15633), .ZN(n15632) );
  NAND2_X1 U15550 ( .A1(a_30_), .A2(n8770), .ZN(n15633) );
  AND3_X1 U15551 ( .A1(b_1_), .A2(b_2_), .A3(n7818), .ZN(n15431) );
  XNOR2_X1 U15552 ( .A(n15635), .B(n15636), .ZN(n15413) );
  NOR2_X1 U15553 ( .A1(n7867), .A2(n8770), .ZN(n15636) );
  XOR2_X1 U15554 ( .A(n15637), .B(n15638), .Z(n15635) );
  XOR2_X1 U15555 ( .A(n15639), .B(n15640), .Z(n15404) );
  XNOR2_X1 U15556 ( .A(n15641), .B(n15642), .ZN(n15640) );
  NAND2_X1 U15557 ( .A1(b_0_), .A2(a_29_), .ZN(n15639) );
  XNOR2_X1 U15558 ( .A(n15643), .B(n15644), .ZN(n15397) );
  XNOR2_X1 U15559 ( .A(n15645), .B(n15646), .ZN(n15644) );
  NAND2_X1 U15560 ( .A1(b_0_), .A2(a_28_), .ZN(n15643) );
  XOR2_X1 U15561 ( .A(n15647), .B(n15648), .Z(n15385) );
  XNOR2_X1 U15562 ( .A(n15649), .B(n15650), .ZN(n15648) );
  NAND2_X1 U15563 ( .A1(b_0_), .A2(a_26_), .ZN(n15647) );
  XOR2_X1 U15564 ( .A(n15651), .B(n15652), .Z(n15436) );
  NOR2_X1 U15565 ( .A1(n8744), .A2(n8770), .ZN(n15652) );
  XOR2_X1 U15566 ( .A(n15653), .B(n15654), .Z(n15651) );
  XNOR2_X1 U15567 ( .A(n15655), .B(n15656), .ZN(n15375) );
  XNOR2_X1 U15568 ( .A(n15657), .B(n15658), .ZN(n15656) );
  NAND2_X1 U15569 ( .A1(b_0_), .A2(a_24_), .ZN(n15655) );
  XNOR2_X1 U15570 ( .A(n15659), .B(n15660), .ZN(n15441) );
  NOR2_X1 U15571 ( .A1(n8747), .A2(n8770), .ZN(n15660) );
  XOR2_X1 U15572 ( .A(n15661), .B(n15662), .Z(n15659) );
  XOR2_X1 U15573 ( .A(n15663), .B(n15664), .Z(n15363) );
  XNOR2_X1 U15574 ( .A(n15665), .B(n15666), .ZN(n15664) );
  NAND2_X1 U15575 ( .A1(b_0_), .A2(a_22_), .ZN(n15663) );
  XNOR2_X1 U15576 ( .A(n15667), .B(n15668), .ZN(n15445) );
  NOR2_X1 U15577 ( .A1(n8750), .A2(n8770), .ZN(n15668) );
  XOR2_X1 U15578 ( .A(n15669), .B(n15670), .Z(n15667) );
  XOR2_X1 U15579 ( .A(n15671), .B(n15672), .Z(n15352) );
  XNOR2_X1 U15580 ( .A(n15673), .B(n15674), .ZN(n15672) );
  NAND2_X1 U15581 ( .A1(b_0_), .A2(a_20_), .ZN(n15671) );
  XNOR2_X1 U15582 ( .A(n15675), .B(n15676), .ZN(n15449) );
  NOR2_X1 U15583 ( .A1(n8170), .A2(n8770), .ZN(n15676) );
  XOR2_X1 U15584 ( .A(n15677), .B(n15678), .Z(n15675) );
  XOR2_X1 U15585 ( .A(n15679), .B(n15680), .Z(n15453) );
  NOR2_X1 U15586 ( .A1(n8755), .A2(n8634), .ZN(n15680) );
  XOR2_X1 U15587 ( .A(n15681), .B(n15682), .Z(n15679) );
  XOR2_X1 U15588 ( .A(n15683), .B(n15684), .Z(n15457) );
  NOR2_X1 U15589 ( .A1(n8757), .A2(n8634), .ZN(n15684) );
  XOR2_X1 U15590 ( .A(n15685), .B(n15686), .Z(n15683) );
  XOR2_X1 U15591 ( .A(n15687), .B(n15688), .Z(n15461) );
  NOR2_X1 U15592 ( .A1(n8759), .A2(n8634), .ZN(n15688) );
  XOR2_X1 U15593 ( .A(n15689), .B(n15690), .Z(n15687) );
  XOR2_X1 U15594 ( .A(n15691), .B(n15692), .Z(n15465) );
  NOR2_X1 U15595 ( .A1(n8761), .A2(n8634), .ZN(n15692) );
  XOR2_X1 U15596 ( .A(n15693), .B(n15694), .Z(n15691) );
  XOR2_X1 U15597 ( .A(n15695), .B(n15696), .Z(n15469) );
  NOR2_X1 U15598 ( .A1(n8763), .A2(n8634), .ZN(n15696) );
  XOR2_X1 U15599 ( .A(n15697), .B(n15698), .Z(n15695) );
  XOR2_X1 U15600 ( .A(n15699), .B(n15700), .Z(n15473) );
  NOR2_X1 U15601 ( .A1(n8491), .A2(n8634), .ZN(n15700) );
  XOR2_X1 U15602 ( .A(n15701), .B(n15702), .Z(n15699) );
  XOR2_X1 U15603 ( .A(n15703), .B(n15704), .Z(n15477) );
  NOR2_X1 U15604 ( .A1(n8766), .A2(n8634), .ZN(n15704) );
  XOR2_X1 U15605 ( .A(n15705), .B(n15706), .Z(n15703) );
  NAND2_X1 U15606 ( .A1(b_2_), .A2(a_2_), .ZN(n8661) );
  XOR2_X1 U15607 ( .A(n15707), .B(n15708), .Z(n15481) );
  NOR2_X1 U15608 ( .A1(n8768), .A2(n8634), .ZN(n15708) );
  XOR2_X1 U15609 ( .A(n15709), .B(n15710), .Z(n15707) );
  XOR2_X1 U15610 ( .A(n15711), .B(n15712), .Z(n8920) );
  NOR2_X1 U15611 ( .A1(n8617), .A2(n8770), .ZN(n15712) );
  XOR2_X1 U15612 ( .A(n15713), .B(n15714), .Z(n15711) );
  XOR2_X1 U15613 ( .A(n8919), .B(n8918), .Z(n15488) );
  NOR2_X1 U15614 ( .A1(n8770), .A2(n9674), .ZN(n8918) );
  INV_X1 U15615 ( .A(n8917), .ZN(n8919) );
  NAND2_X1 U15616 ( .A1(n15715), .A2(n15716), .ZN(n8917) );
  NAND3_X1 U15617 ( .A1(a_1_), .A2(n15717), .A3(b_0_), .ZN(n15716) );
  OR2_X1 U15618 ( .A1(n15714), .A2(n15713), .ZN(n15717) );
  NAND2_X1 U15619 ( .A1(n15713), .A2(n15714), .ZN(n15715) );
  NAND2_X1 U15620 ( .A1(n15718), .A2(n15719), .ZN(n15714) );
  NAND3_X1 U15621 ( .A1(a_2_), .A2(n15720), .A3(b_0_), .ZN(n15719) );
  OR2_X1 U15622 ( .A1(n15496), .A2(n8660), .ZN(n15720) );
  NAND2_X1 U15623 ( .A1(n8660), .A2(n15496), .ZN(n15718) );
  NAND2_X1 U15624 ( .A1(n15721), .A2(n15722), .ZN(n15496) );
  NAND3_X1 U15625 ( .A1(a_2_), .A2(n15723), .A3(b_1_), .ZN(n15722) );
  OR2_X1 U15626 ( .A1(n15710), .A2(n15709), .ZN(n15723) );
  NAND2_X1 U15627 ( .A1(n15709), .A2(n15710), .ZN(n15721) );
  NAND2_X1 U15628 ( .A1(n15724), .A2(n15725), .ZN(n15710) );
  NAND3_X1 U15629 ( .A1(a_3_), .A2(n15726), .A3(b_1_), .ZN(n15725) );
  OR2_X1 U15630 ( .A1(n15506), .A2(n15505), .ZN(n15726) );
  NAND2_X1 U15631 ( .A1(n15505), .A2(n15506), .ZN(n15724) );
  NAND2_X1 U15632 ( .A1(n15727), .A2(n15728), .ZN(n15506) );
  NAND3_X1 U15633 ( .A1(a_4_), .A2(n15729), .A3(b_1_), .ZN(n15728) );
  OR2_X1 U15634 ( .A1(n15706), .A2(n15705), .ZN(n15729) );
  NAND2_X1 U15635 ( .A1(n15705), .A2(n15706), .ZN(n15727) );
  NAND2_X1 U15636 ( .A1(n15730), .A2(n15731), .ZN(n15706) );
  NAND3_X1 U15637 ( .A1(a_5_), .A2(n15732), .A3(b_1_), .ZN(n15731) );
  OR2_X1 U15638 ( .A1(n15517), .A2(n15516), .ZN(n15732) );
  NAND2_X1 U15639 ( .A1(n15516), .A2(n15517), .ZN(n15730) );
  NAND2_X1 U15640 ( .A1(n15733), .A2(n15734), .ZN(n15517) );
  NAND3_X1 U15641 ( .A1(a_6_), .A2(n15735), .A3(b_1_), .ZN(n15734) );
  OR2_X1 U15642 ( .A1(n15702), .A2(n15701), .ZN(n15735) );
  NAND2_X1 U15643 ( .A1(n15701), .A2(n15702), .ZN(n15733) );
  NAND2_X1 U15644 ( .A1(n15736), .A2(n15737), .ZN(n15702) );
  NAND3_X1 U15645 ( .A1(a_7_), .A2(n15738), .A3(b_1_), .ZN(n15737) );
  OR2_X1 U15646 ( .A1(n15528), .A2(n15527), .ZN(n15738) );
  NAND2_X1 U15647 ( .A1(n15527), .A2(n15528), .ZN(n15736) );
  NAND2_X1 U15648 ( .A1(n15739), .A2(n15740), .ZN(n15528) );
  NAND3_X1 U15649 ( .A1(a_8_), .A2(n15741), .A3(b_1_), .ZN(n15740) );
  OR2_X1 U15650 ( .A1(n15698), .A2(n15697), .ZN(n15741) );
  NAND2_X1 U15651 ( .A1(n15697), .A2(n15698), .ZN(n15739) );
  NAND2_X1 U15652 ( .A1(n15742), .A2(n15743), .ZN(n15698) );
  NAND3_X1 U15653 ( .A1(a_9_), .A2(n15744), .A3(b_1_), .ZN(n15743) );
  OR2_X1 U15654 ( .A1(n15539), .A2(n15538), .ZN(n15744) );
  NAND2_X1 U15655 ( .A1(n15538), .A2(n15539), .ZN(n15742) );
  NAND2_X1 U15656 ( .A1(n15745), .A2(n15746), .ZN(n15539) );
  NAND3_X1 U15657 ( .A1(a_10_), .A2(n15747), .A3(b_1_), .ZN(n15746) );
  OR2_X1 U15658 ( .A1(n15694), .A2(n15693), .ZN(n15747) );
  NAND2_X1 U15659 ( .A1(n15693), .A2(n15694), .ZN(n15745) );
  NAND2_X1 U15660 ( .A1(n15748), .A2(n15749), .ZN(n15694) );
  NAND3_X1 U15661 ( .A1(a_11_), .A2(n15750), .A3(b_1_), .ZN(n15749) );
  OR2_X1 U15662 ( .A1(n15550), .A2(n15549), .ZN(n15750) );
  NAND2_X1 U15663 ( .A1(n15549), .A2(n15550), .ZN(n15748) );
  NAND2_X1 U15664 ( .A1(n15751), .A2(n15752), .ZN(n15550) );
  NAND3_X1 U15665 ( .A1(a_12_), .A2(n15753), .A3(b_1_), .ZN(n15752) );
  OR2_X1 U15666 ( .A1(n15690), .A2(n15689), .ZN(n15753) );
  NAND2_X1 U15667 ( .A1(n15689), .A2(n15690), .ZN(n15751) );
  NAND2_X1 U15668 ( .A1(n15754), .A2(n15755), .ZN(n15690) );
  NAND3_X1 U15669 ( .A1(a_13_), .A2(n15756), .A3(b_1_), .ZN(n15755) );
  OR2_X1 U15670 ( .A1(n15561), .A2(n15560), .ZN(n15756) );
  NAND2_X1 U15671 ( .A1(n15560), .A2(n15561), .ZN(n15754) );
  NAND2_X1 U15672 ( .A1(n15757), .A2(n15758), .ZN(n15561) );
  NAND3_X1 U15673 ( .A1(a_14_), .A2(n15759), .A3(b_1_), .ZN(n15758) );
  OR2_X1 U15674 ( .A1(n15686), .A2(n15685), .ZN(n15759) );
  NAND2_X1 U15675 ( .A1(n15685), .A2(n15686), .ZN(n15757) );
  NAND2_X1 U15676 ( .A1(n15760), .A2(n15761), .ZN(n15686) );
  NAND3_X1 U15677 ( .A1(a_15_), .A2(n15762), .A3(b_1_), .ZN(n15761) );
  OR2_X1 U15678 ( .A1(n15572), .A2(n15571), .ZN(n15762) );
  NAND2_X1 U15679 ( .A1(n15571), .A2(n15572), .ZN(n15760) );
  NAND2_X1 U15680 ( .A1(n15763), .A2(n15764), .ZN(n15572) );
  NAND3_X1 U15681 ( .A1(a_16_), .A2(n15765), .A3(b_1_), .ZN(n15764) );
  OR2_X1 U15682 ( .A1(n15682), .A2(n15681), .ZN(n15765) );
  NAND2_X1 U15683 ( .A1(n15681), .A2(n15682), .ZN(n15763) );
  NAND2_X1 U15684 ( .A1(n15766), .A2(n15767), .ZN(n15682) );
  NAND3_X1 U15685 ( .A1(a_17_), .A2(n15768), .A3(b_1_), .ZN(n15767) );
  OR2_X1 U15686 ( .A1(n15583), .A2(n15582), .ZN(n15768) );
  NAND2_X1 U15687 ( .A1(n15582), .A2(n15583), .ZN(n15766) );
  NAND2_X1 U15688 ( .A1(n15769), .A2(n15770), .ZN(n15583) );
  NAND3_X1 U15689 ( .A1(a_19_), .A2(n15771), .A3(b_0_), .ZN(n15770) );
  OR2_X1 U15690 ( .A1(n15678), .A2(n15677), .ZN(n15771) );
  NAND2_X1 U15691 ( .A1(n15677), .A2(n15678), .ZN(n15769) );
  NAND2_X1 U15692 ( .A1(n15772), .A2(n15773), .ZN(n15678) );
  NAND3_X1 U15693 ( .A1(a_20_), .A2(n15774), .A3(b_0_), .ZN(n15773) );
  OR2_X1 U15694 ( .A1(n15674), .A2(n15673), .ZN(n15774) );
  NAND2_X1 U15695 ( .A1(n15673), .A2(n15674), .ZN(n15772) );
  NAND2_X1 U15696 ( .A1(n15775), .A2(n15776), .ZN(n15674) );
  NAND3_X1 U15697 ( .A1(a_21_), .A2(n15777), .A3(b_0_), .ZN(n15776) );
  NAND2_X1 U15698 ( .A1(n15670), .A2(n15669), .ZN(n15777) );
  INV_X1 U15699 ( .A(n15778), .ZN(n15670) );
  NAND2_X1 U15700 ( .A1(n15779), .A2(n15778), .ZN(n15775) );
  NAND2_X1 U15701 ( .A1(n15780), .A2(n15781), .ZN(n15778) );
  NAND3_X1 U15702 ( .A1(a_22_), .A2(n15782), .A3(b_0_), .ZN(n15781) );
  OR2_X1 U15703 ( .A1(n15666), .A2(n15665), .ZN(n15782) );
  NAND2_X1 U15704 ( .A1(n15665), .A2(n15666), .ZN(n15780) );
  NAND2_X1 U15705 ( .A1(n15783), .A2(n15784), .ZN(n15666) );
  NAND3_X1 U15706 ( .A1(a_23_), .A2(n15785), .A3(b_0_), .ZN(n15784) );
  NAND2_X1 U15707 ( .A1(n15662), .A2(n15661), .ZN(n15785) );
  INV_X1 U15708 ( .A(n15786), .ZN(n15662) );
  NAND2_X1 U15709 ( .A1(n15787), .A2(n15786), .ZN(n15783) );
  NAND2_X1 U15710 ( .A1(n15788), .A2(n15789), .ZN(n15786) );
  NAND3_X1 U15711 ( .A1(a_24_), .A2(n15790), .A3(b_0_), .ZN(n15789) );
  OR2_X1 U15712 ( .A1(n15658), .A2(n15657), .ZN(n15790) );
  NAND2_X1 U15713 ( .A1(n15657), .A2(n15658), .ZN(n15788) );
  NAND2_X1 U15714 ( .A1(n15791), .A2(n15792), .ZN(n15658) );
  NAND3_X1 U15715 ( .A1(a_25_), .A2(n15793), .A3(b_0_), .ZN(n15792) );
  NAND2_X1 U15716 ( .A1(n15654), .A2(n15653), .ZN(n15793) );
  INV_X1 U15717 ( .A(n15794), .ZN(n15654) );
  NAND2_X1 U15718 ( .A1(n15795), .A2(n15794), .ZN(n15791) );
  NAND2_X1 U15719 ( .A1(n15796), .A2(n15797), .ZN(n15794) );
  NAND3_X1 U15720 ( .A1(a_26_), .A2(n15798), .A3(b_0_), .ZN(n15797) );
  OR2_X1 U15721 ( .A1(n15650), .A2(n15649), .ZN(n15798) );
  NAND2_X1 U15722 ( .A1(n15649), .A2(n15650), .ZN(n15796) );
  NAND2_X1 U15723 ( .A1(n15799), .A2(n15800), .ZN(n15650) );
  NAND3_X1 U15724 ( .A1(a_27_), .A2(n15801), .A3(b_0_), .ZN(n15800) );
  NAND2_X1 U15725 ( .A1(n15615), .A2(n15614), .ZN(n15801) );
  INV_X1 U15726 ( .A(n15802), .ZN(n15615) );
  NAND2_X1 U15727 ( .A1(n15803), .A2(n15802), .ZN(n15799) );
  NAND2_X1 U15728 ( .A1(n15804), .A2(n15805), .ZN(n15802) );
  NAND3_X1 U15729 ( .A1(a_28_), .A2(n15806), .A3(b_0_), .ZN(n15805) );
  OR2_X1 U15730 ( .A1(n15646), .A2(n15645), .ZN(n15806) );
  NAND2_X1 U15731 ( .A1(n15645), .A2(n15646), .ZN(n15804) );
  NAND2_X1 U15732 ( .A1(n15807), .A2(n15808), .ZN(n15646) );
  NAND3_X1 U15733 ( .A1(a_29_), .A2(n15809), .A3(b_0_), .ZN(n15808) );
  OR2_X1 U15734 ( .A1(n15642), .A2(n15641), .ZN(n15809) );
  NAND2_X1 U15735 ( .A1(n15641), .A2(n15642), .ZN(n15807) );
  NAND2_X1 U15736 ( .A1(n15638), .A2(n15810), .ZN(n15642) );
  NAND3_X1 U15737 ( .A1(b_0_), .A2(a_30_), .A3(n15637), .ZN(n15810) );
  NOR2_X1 U15738 ( .A1(n8634), .A2(n7890), .ZN(n15637) );
  NAND3_X1 U15739 ( .A1(b_0_), .A2(b_1_), .A3(n7818), .ZN(n15638) );
  NOR2_X1 U15740 ( .A1(n8634), .A2(n8739), .ZN(n15641) );
  NOR2_X1 U15741 ( .A1(n8634), .A2(n8741), .ZN(n15645) );
  INV_X1 U15742 ( .A(n15614), .ZN(n15803) );
  NAND2_X1 U15743 ( .A1(b_1_), .A2(a_26_), .ZN(n15614) );
  NOR2_X1 U15744 ( .A1(n8634), .A2(n8744), .ZN(n15649) );
  INV_X1 U15745 ( .A(n15653), .ZN(n15795) );
  NAND2_X1 U15746 ( .A1(b_1_), .A2(a_24_), .ZN(n15653) );
  NOR2_X1 U15747 ( .A1(n8634), .A2(n8747), .ZN(n15657) );
  INV_X1 U15748 ( .A(n15661), .ZN(n15787) );
  NAND2_X1 U15749 ( .A1(b_1_), .A2(a_22_), .ZN(n15661) );
  NOR2_X1 U15750 ( .A1(n8634), .A2(n8750), .ZN(n15665) );
  INV_X1 U15751 ( .A(n15669), .ZN(n15779) );
  NAND2_X1 U15752 ( .A1(b_1_), .A2(a_20_), .ZN(n15669) );
  NOR2_X1 U15753 ( .A1(n8634), .A2(n8170), .ZN(n15673) );
  NOR2_X1 U15754 ( .A1(n8634), .A2(n8753), .ZN(n15677) );
  NOR2_X1 U15755 ( .A1(n8770), .A2(n8753), .ZN(n15582) );
  NOR2_X1 U15756 ( .A1(n8770), .A2(n8210), .ZN(n15681) );
  NOR2_X1 U15757 ( .A1(n8770), .A2(n8755), .ZN(n15571) );
  NOR2_X1 U15758 ( .A1(n8770), .A2(n8276), .ZN(n15685) );
  NOR2_X1 U15759 ( .A1(n8770), .A2(n8757), .ZN(n15560) );
  NOR2_X1 U15760 ( .A1(n8770), .A2(n8310), .ZN(n15689) );
  NOR2_X1 U15761 ( .A1(n8770), .A2(n8759), .ZN(n15549) );
  NOR2_X1 U15762 ( .A1(n8770), .A2(n8376), .ZN(n15693) );
  NOR2_X1 U15763 ( .A1(n8770), .A2(n8761), .ZN(n15538) );
  NOR2_X1 U15764 ( .A1(n8770), .A2(n8426), .ZN(n15697) );
  NOR2_X1 U15765 ( .A1(n8770), .A2(n8763), .ZN(n15527) );
  NOR2_X1 U15766 ( .A1(n8770), .A2(n8764), .ZN(n15701) );
  NOR2_X1 U15767 ( .A1(n8770), .A2(n8491), .ZN(n15516) );
  NOR2_X1 U15768 ( .A1(n8770), .A2(n8517), .ZN(n15705) );
  NOR2_X1 U15769 ( .A1(n8770), .A2(n8766), .ZN(n15505) );
  NOR2_X1 U15770 ( .A1(n8770), .A2(n8567), .ZN(n15709) );
  NOR2_X1 U15771 ( .A1(n8634), .A2(n8617), .ZN(n8660) );
  NOR2_X1 U15772 ( .A1(n8634), .A2(n9674), .ZN(n15713) );
  NAND3_X1 U15773 ( .A1(n15815), .A2(n15816), .A3(n7822), .ZN(n15814) );
  INV_X1 U15774 ( .A(operation_1_), .ZN(n15812) );
  NAND2_X1 U15775 ( .A1(n15817), .A2(n8770), .ZN(n15816) );
  NAND2_X1 U15776 ( .A1(n8769), .A2(n9674), .ZN(n15817) );
  INV_X1 U15777 ( .A(n8650), .ZN(n8769) );
  NAND2_X1 U15778 ( .A1(a_0_), .A2(n8650), .ZN(n15815) );
  NAND2_X1 U15779 ( .A1(n15818), .A2(n15819), .ZN(n8650) );
  NAND2_X1 U15780 ( .A1(n15820), .A2(n8634), .ZN(n15819) );
  INV_X1 U15781 ( .A(b_1_), .ZN(n8634) );
  NAND2_X1 U15782 ( .A1(n8633), .A2(n8617), .ZN(n15820) );
  INV_X1 U15783 ( .A(n8626), .ZN(n8633) );
  NAND2_X1 U15784 ( .A1(a_1_), .A2(n8626), .ZN(n15818) );
  NAND2_X1 U15785 ( .A1(n15821), .A2(n15822), .ZN(n8626) );
  NAND2_X1 U15786 ( .A1(n15823), .A2(n8608), .ZN(n15822) );
  INV_X1 U15787 ( .A(b_2_), .ZN(n8608) );
  NAND2_X1 U15788 ( .A1(n8607), .A2(n8768), .ZN(n15823) );
  INV_X1 U15789 ( .A(n8600), .ZN(n8607) );
  NAND2_X1 U15790 ( .A1(a_2_), .A2(n8600), .ZN(n15821) );
  NAND2_X1 U15791 ( .A1(n15824), .A2(n15825), .ZN(n8600) );
  NAND2_X1 U15792 ( .A1(n15826), .A2(n8767), .ZN(n15825) );
  INV_X1 U15793 ( .A(b_3_), .ZN(n8767) );
  NAND2_X1 U15794 ( .A1(n8583), .A2(n8567), .ZN(n15826) );
  INV_X1 U15795 ( .A(n8576), .ZN(n8583) );
  NAND2_X1 U15796 ( .A1(a_3_), .A2(n8576), .ZN(n15824) );
  NAND2_X1 U15797 ( .A1(n15827), .A2(n15828), .ZN(n8576) );
  NAND2_X1 U15798 ( .A1(n15829), .A2(n8558), .ZN(n15828) );
  NAND2_X1 U15799 ( .A1(n8557), .A2(n8766), .ZN(n15829) );
  INV_X1 U15800 ( .A(n8550), .ZN(n8557) );
  NAND2_X1 U15801 ( .A1(a_4_), .A2(n8550), .ZN(n15827) );
  NAND2_X1 U15802 ( .A1(n15830), .A2(n15831), .ZN(n8550) );
  NAND2_X1 U15803 ( .A1(n15832), .A2(n8765), .ZN(n15831) );
  INV_X1 U15804 ( .A(b_5_), .ZN(n8765) );
  NAND2_X1 U15805 ( .A1(n8533), .A2(n8517), .ZN(n15832) );
  INV_X1 U15806 ( .A(n8526), .ZN(n8533) );
  NAND2_X1 U15807 ( .A1(a_5_), .A2(n8526), .ZN(n15830) );
  NAND2_X1 U15808 ( .A1(n15833), .A2(n15834), .ZN(n8526) );
  NAND2_X1 U15809 ( .A1(n15835), .A2(n8508), .ZN(n15834) );
  NAND2_X1 U15810 ( .A1(n8507), .A2(n8491), .ZN(n15835) );
  INV_X1 U15811 ( .A(n8500), .ZN(n8507) );
  NAND2_X1 U15812 ( .A1(a_6_), .A2(n8500), .ZN(n15833) );
  NAND2_X1 U15813 ( .A1(n15836), .A2(n15837), .ZN(n8500) );
  NAND2_X1 U15814 ( .A1(n15838), .A2(n8482), .ZN(n15837) );
  NAND2_X1 U15815 ( .A1(n8481), .A2(n8764), .ZN(n15838) );
  INV_X1 U15816 ( .A(n8473), .ZN(n8481) );
  NAND2_X1 U15817 ( .A1(a_7_), .A2(n8473), .ZN(n15836) );
  NAND2_X1 U15818 ( .A1(n15839), .A2(n15840), .ZN(n8473) );
  NAND2_X1 U15819 ( .A1(n15841), .A2(n8451), .ZN(n15840) );
  INV_X1 U15820 ( .A(b_8_), .ZN(n8451) );
  NAND2_X1 U15821 ( .A1(n8450), .A2(n8763), .ZN(n15841) );
  INV_X1 U15822 ( .A(n8443), .ZN(n8450) );
  NAND2_X1 U15823 ( .A1(a_8_), .A2(n8443), .ZN(n15839) );
  NAND2_X1 U15824 ( .A1(n15842), .A2(n15843), .ZN(n8443) );
  NAND2_X1 U15825 ( .A1(n15844), .A2(n8762), .ZN(n15843) );
  INV_X1 U15826 ( .A(b_9_), .ZN(n8762) );
  NAND2_X1 U15827 ( .A1(n8425), .A2(n8426), .ZN(n15844) );
  INV_X1 U15828 ( .A(n8418), .ZN(n8425) );
  NAND2_X1 U15829 ( .A1(a_9_), .A2(n8418), .ZN(n15842) );
  NAND2_X1 U15830 ( .A1(n15845), .A2(n15846), .ZN(n8418) );
  NAND2_X1 U15831 ( .A1(n15847), .A2(n8401), .ZN(n15846) );
  INV_X1 U15832 ( .A(b_10_), .ZN(n8401) );
  NAND2_X1 U15833 ( .A1(n8400), .A2(n8761), .ZN(n15847) );
  INV_X1 U15834 ( .A(n8393), .ZN(n8400) );
  NAND2_X1 U15835 ( .A1(a_10_), .A2(n8393), .ZN(n15845) );
  NAND2_X1 U15836 ( .A1(n15848), .A2(n15849), .ZN(n8393) );
  NAND2_X1 U15837 ( .A1(n15850), .A2(n8760), .ZN(n15849) );
  INV_X1 U15838 ( .A(b_11_), .ZN(n8760) );
  NAND2_X1 U15839 ( .A1(n8375), .A2(n8376), .ZN(n15850) );
  INV_X1 U15840 ( .A(n8367), .ZN(n8375) );
  NAND2_X1 U15841 ( .A1(a_11_), .A2(n8367), .ZN(n15848) );
  NAND2_X1 U15842 ( .A1(n15851), .A2(n15852), .ZN(n8367) );
  NAND2_X1 U15843 ( .A1(n15853), .A2(n8351), .ZN(n15852) );
  INV_X1 U15844 ( .A(b_12_), .ZN(n8351) );
  NAND2_X1 U15845 ( .A1(n8350), .A2(n8759), .ZN(n15853) );
  INV_X1 U15846 ( .A(n8343), .ZN(n8350) );
  NAND2_X1 U15847 ( .A1(a_12_), .A2(n8343), .ZN(n15851) );
  NAND2_X1 U15848 ( .A1(n15854), .A2(n15855), .ZN(n8343) );
  NAND2_X1 U15849 ( .A1(n15856), .A2(n8758), .ZN(n15855) );
  INV_X1 U15850 ( .A(b_13_), .ZN(n8758) );
  NAND2_X1 U15851 ( .A1(n8326), .A2(n8310), .ZN(n15856) );
  INV_X1 U15852 ( .A(n8319), .ZN(n8326) );
  NAND2_X1 U15853 ( .A1(a_13_), .A2(n8319), .ZN(n15854) );
  NAND2_X1 U15854 ( .A1(n15857), .A2(n15858), .ZN(n8319) );
  NAND2_X1 U15855 ( .A1(n15859), .A2(n8301), .ZN(n15858) );
  NAND2_X1 U15856 ( .A1(n8300), .A2(n8757), .ZN(n15859) );
  INV_X1 U15857 ( .A(n8292), .ZN(n8300) );
  NAND2_X1 U15858 ( .A1(a_14_), .A2(n8292), .ZN(n15857) );
  NAND2_X1 U15859 ( .A1(n15860), .A2(n15861), .ZN(n8292) );
  NAND2_X1 U15860 ( .A1(n15862), .A2(n8756), .ZN(n15861) );
  INV_X1 U15861 ( .A(b_15_), .ZN(n8756) );
  NAND2_X1 U15862 ( .A1(n8275), .A2(n8276), .ZN(n15862) );
  INV_X1 U15863 ( .A(n8267), .ZN(n8275) );
  NAND2_X1 U15864 ( .A1(a_15_), .A2(n8267), .ZN(n15860) );
  NAND2_X1 U15865 ( .A1(n15863), .A2(n15864), .ZN(n8267) );
  NAND2_X1 U15866 ( .A1(n15865), .A2(n8251), .ZN(n15864) );
  NAND2_X1 U15867 ( .A1(n8250), .A2(n8755), .ZN(n15865) );
  INV_X1 U15868 ( .A(n8243), .ZN(n8250) );
  NAND2_X1 U15869 ( .A1(a_16_), .A2(n8243), .ZN(n15863) );
  NAND2_X1 U15870 ( .A1(n15866), .A2(n15867), .ZN(n8243) );
  NAND2_X1 U15871 ( .A1(n15868), .A2(n8754), .ZN(n15867) );
  INV_X1 U15872 ( .A(b_17_), .ZN(n8754) );
  NAND2_X1 U15873 ( .A1(n8226), .A2(n8210), .ZN(n15868) );
  INV_X1 U15874 ( .A(n8219), .ZN(n8226) );
  NAND2_X1 U15875 ( .A1(a_17_), .A2(n8219), .ZN(n15866) );
  NAND2_X1 U15876 ( .A1(n15869), .A2(n15870), .ZN(n8219) );
  NAND2_X1 U15877 ( .A1(n15871), .A2(n8195), .ZN(n15870) );
  INV_X1 U15878 ( .A(b_18_), .ZN(n8195) );
  NAND2_X1 U15879 ( .A1(n8194), .A2(n8753), .ZN(n15871) );
  INV_X1 U15880 ( .A(n8187), .ZN(n8194) );
  NAND2_X1 U15881 ( .A1(a_18_), .A2(n8187), .ZN(n15869) );
  NAND2_X1 U15882 ( .A1(n15872), .A2(n15873), .ZN(n8187) );
  NAND2_X1 U15883 ( .A1(n15874), .A2(n8752), .ZN(n15873) );
  INV_X1 U15884 ( .A(b_19_), .ZN(n8752) );
  NAND2_X1 U15885 ( .A1(n8169), .A2(n8170), .ZN(n15874) );
  INV_X1 U15886 ( .A(n8162), .ZN(n8169) );
  NAND2_X1 U15887 ( .A1(a_19_), .A2(n8162), .ZN(n15872) );
  NAND2_X1 U15888 ( .A1(n15875), .A2(n15876), .ZN(n8162) );
  NAND2_X1 U15889 ( .A1(n15877), .A2(n8145), .ZN(n15876) );
  INV_X1 U15890 ( .A(b_20_), .ZN(n8145) );
  NAND2_X1 U15891 ( .A1(n8144), .A2(n8751), .ZN(n15877) );
  INV_X1 U15892 ( .A(n8137), .ZN(n8144) );
  NAND2_X1 U15893 ( .A1(a_20_), .A2(n8137), .ZN(n15875) );
  NAND2_X1 U15894 ( .A1(n15878), .A2(n15879), .ZN(n8137) );
  NAND2_X1 U15895 ( .A1(n15880), .A2(n8749), .ZN(n15879) );
  INV_X1 U15896 ( .A(b_21_), .ZN(n8749) );
  NAND2_X1 U15897 ( .A1(n8110), .A2(n8750), .ZN(n15880) );
  INV_X1 U15898 ( .A(n8118), .ZN(n8110) );
  NAND2_X1 U15899 ( .A1(a_21_), .A2(n8118), .ZN(n15878) );
  NAND2_X1 U15900 ( .A1(n15881), .A2(n15882), .ZN(n8118) );
  NAND2_X1 U15901 ( .A1(n15883), .A2(n8094), .ZN(n15882) );
  NAND2_X1 U15902 ( .A1(n8093), .A2(n8748), .ZN(n15883) );
  INV_X1 U15903 ( .A(n8086), .ZN(n8093) );
  NAND2_X1 U15904 ( .A1(a_22_), .A2(n8086), .ZN(n15881) );
  NAND2_X1 U15905 ( .A1(n15884), .A2(n15885), .ZN(n8086) );
  NAND2_X1 U15906 ( .A1(n15886), .A2(n8746), .ZN(n15885) );
  INV_X1 U15907 ( .A(b_23_), .ZN(n8746) );
  NAND2_X1 U15908 ( .A1(n8059), .A2(n8747), .ZN(n15886) );
  INV_X1 U15909 ( .A(n8067), .ZN(n8059) );
  NAND2_X1 U15910 ( .A1(a_23_), .A2(n8067), .ZN(n15884) );
  NAND2_X1 U15911 ( .A1(n15887), .A2(n15888), .ZN(n8067) );
  NAND2_X1 U15912 ( .A1(n15889), .A2(n8043), .ZN(n15888) );
  INV_X1 U15913 ( .A(b_24_), .ZN(n8043) );
  NAND2_X1 U15914 ( .A1(n8042), .A2(n8745), .ZN(n15889) );
  INV_X1 U15915 ( .A(n8035), .ZN(n8042) );
  NAND2_X1 U15916 ( .A1(a_24_), .A2(n8035), .ZN(n15887) );
  NAND2_X1 U15917 ( .A1(n15890), .A2(n15891), .ZN(n8035) );
  NAND2_X1 U15918 ( .A1(n15892), .A2(n8743), .ZN(n15891) );
  INV_X1 U15919 ( .A(b_25_), .ZN(n8743) );
  NAND2_X1 U15920 ( .A1(n8008), .A2(n8744), .ZN(n15892) );
  INV_X1 U15921 ( .A(n8016), .ZN(n8008) );
  NAND2_X1 U15922 ( .A1(a_25_), .A2(n8016), .ZN(n15890) );
  NAND2_X1 U15923 ( .A1(n15893), .A2(n15894), .ZN(n8016) );
  NAND2_X1 U15924 ( .A1(n15895), .A2(n7992), .ZN(n15894) );
  NAND2_X1 U15925 ( .A1(n7991), .A2(n8742), .ZN(n15895) );
  INV_X1 U15926 ( .A(n7984), .ZN(n7991) );
  NAND2_X1 U15927 ( .A1(a_26_), .A2(n7984), .ZN(n15893) );
  NAND2_X1 U15928 ( .A1(n15896), .A2(n15897), .ZN(n7984) );
  NAND2_X1 U15929 ( .A1(n15898), .A2(n8740), .ZN(n15897) );
  INV_X1 U15930 ( .A(b_27_), .ZN(n8740) );
  NAND2_X1 U15931 ( .A1(n7957), .A2(n8741), .ZN(n15898) );
  INV_X1 U15932 ( .A(n7965), .ZN(n7957) );
  NAND2_X1 U15933 ( .A1(a_27_), .A2(n7965), .ZN(n15896) );
  NAND2_X1 U15934 ( .A1(n15899), .A2(n15900), .ZN(n7965) );
  NAND2_X1 U15935 ( .A1(n15901), .A2(n7935), .ZN(n15900) );
  NAND2_X1 U15936 ( .A1(n7934), .A2(n8739), .ZN(n15901) );
  INV_X1 U15937 ( .A(n7927), .ZN(n7934) );
  NAND2_X1 U15938 ( .A1(a_28_), .A2(n7927), .ZN(n15899) );
  NAND2_X1 U15939 ( .A1(n15902), .A2(n15903), .ZN(n7927) );
  NAND2_X1 U15940 ( .A1(n15904), .A2(n8738), .ZN(n15903) );
  INV_X1 U15941 ( .A(b_29_), .ZN(n8738) );
  NAND2_X1 U15942 ( .A1(n7900), .A2(n7890), .ZN(n15904) );
  INV_X1 U15943 ( .A(n7908), .ZN(n7900) );
  NAND2_X1 U15944 ( .A1(a_29_), .A2(n7908), .ZN(n15902) );
  NAND2_X1 U15945 ( .A1(n15905), .A2(n15906), .ZN(n7908) );
  NAND2_X1 U15946 ( .A1(n15907), .A2(n7869), .ZN(n15906) );
  NAND2_X1 U15947 ( .A1(n7858), .A2(n7867), .ZN(n15907) );
  INV_X1 U15948 ( .A(n7853), .ZN(n7858) );
  NAND2_X1 U15949 ( .A1(a_30_), .A2(n7853), .ZN(n15905) );
  NAND2_X1 U15950 ( .A1(b_31_), .A2(n15634), .ZN(n7853) );
  INV_X1 U15951 ( .A(a_31_), .ZN(n15634) );
  NAND3_X1 U15952 ( .A1(n15908), .A2(n15909), .A3(n7820), .ZN(n15813) );
  INV_X1 U15953 ( .A(operation_0_), .ZN(n15811) );
  NAND2_X1 U15954 ( .A1(b_0_), .A2(n15910), .ZN(n15909) );
  NAND2_X1 U15955 ( .A1(n8656), .A2(a_0_), .ZN(n15910) );
  INV_X1 U15956 ( .A(n8648), .ZN(n8656) );
  NAND2_X1 U15957 ( .A1(n8648), .A2(n9674), .ZN(n15908) );
  INV_X1 U15958 ( .A(a_0_), .ZN(n9674) );
  NAND2_X1 U15959 ( .A1(n15911), .A2(n15912), .ZN(n8648) );
  NAND2_X1 U15960 ( .A1(b_1_), .A2(n15913), .ZN(n15912) );
  NAND2_X1 U15961 ( .A1(n8632), .A2(a_1_), .ZN(n15913) );
  INV_X1 U15962 ( .A(n8623), .ZN(n8632) );
  NAND2_X1 U15963 ( .A1(n8623), .A2(n8617), .ZN(n15911) );
  NAND2_X1 U15964 ( .A1(n15914), .A2(n15915), .ZN(n8623) );
  NAND2_X1 U15965 ( .A1(b_2_), .A2(n15916), .ZN(n15915) );
  NAND2_X1 U15966 ( .A1(n8606), .A2(a_2_), .ZN(n15916) );
  INV_X1 U15967 ( .A(n8597), .ZN(n8606) );
  NAND2_X1 U15968 ( .A1(n8597), .A2(n8768), .ZN(n15914) );
  INV_X1 U15969 ( .A(a_2_), .ZN(n8768) );
  NAND2_X1 U15970 ( .A1(n15917), .A2(n15918), .ZN(n8597) );
  NAND2_X1 U15971 ( .A1(b_3_), .A2(n15919), .ZN(n15918) );
  NAND2_X1 U15972 ( .A1(n8582), .A2(a_3_), .ZN(n15919) );
  INV_X1 U15973 ( .A(n8573), .ZN(n8582) );
  NAND2_X1 U15974 ( .A1(n8573), .A2(n8567), .ZN(n15917) );
  INV_X1 U15975 ( .A(a_3_), .ZN(n8567) );
  NAND2_X1 U15976 ( .A1(n15920), .A2(n15921), .ZN(n8573) );
  NAND2_X1 U15977 ( .A1(b_4_), .A2(n15922), .ZN(n15921) );
  NAND2_X1 U15978 ( .A1(n8556), .A2(a_4_), .ZN(n15922) );
  INV_X1 U15979 ( .A(n8547), .ZN(n8556) );
  NAND2_X1 U15980 ( .A1(n8547), .A2(n8766), .ZN(n15920) );
  INV_X1 U15981 ( .A(a_4_), .ZN(n8766) );
  NAND2_X1 U15982 ( .A1(n15923), .A2(n15924), .ZN(n8547) );
  NAND2_X1 U15983 ( .A1(b_5_), .A2(n15925), .ZN(n15924) );
  NAND2_X1 U15984 ( .A1(n8532), .A2(a_5_), .ZN(n15925) );
  INV_X1 U15985 ( .A(n8523), .ZN(n8532) );
  NAND2_X1 U15986 ( .A1(n8523), .A2(n8517), .ZN(n15923) );
  INV_X1 U15987 ( .A(a_5_), .ZN(n8517) );
  NAND2_X1 U15988 ( .A1(n15926), .A2(n15927), .ZN(n8523) );
  NAND2_X1 U15989 ( .A1(b_6_), .A2(n15928), .ZN(n15927) );
  NAND2_X1 U15990 ( .A1(n8506), .A2(a_6_), .ZN(n15928) );
  INV_X1 U15991 ( .A(n8497), .ZN(n8506) );
  NAND2_X1 U15992 ( .A1(n8497), .A2(n8491), .ZN(n15926) );
  INV_X1 U15993 ( .A(a_6_), .ZN(n8491) );
  NAND2_X1 U15994 ( .A1(n15929), .A2(n15930), .ZN(n8497) );
  NAND2_X1 U15995 ( .A1(b_7_), .A2(n15931), .ZN(n15930) );
  NAND2_X1 U15996 ( .A1(n8479), .A2(a_7_), .ZN(n15931) );
  INV_X1 U15997 ( .A(n8471), .ZN(n8479) );
  NAND2_X1 U15998 ( .A1(n8471), .A2(n8764), .ZN(n15929) );
  INV_X1 U15999 ( .A(a_7_), .ZN(n8764) );
  NAND2_X1 U16000 ( .A1(n15932), .A2(n15933), .ZN(n8471) );
  NAND2_X1 U16001 ( .A1(b_8_), .A2(n15934), .ZN(n15933) );
  NAND2_X1 U16002 ( .A1(n8449), .A2(a_8_), .ZN(n15934) );
  INV_X1 U16003 ( .A(n8440), .ZN(n8449) );
  NAND2_X1 U16004 ( .A1(n8440), .A2(n8763), .ZN(n15932) );
  INV_X1 U16005 ( .A(a_8_), .ZN(n8763) );
  NAND2_X1 U16006 ( .A1(n15935), .A2(n15936), .ZN(n8440) );
  NAND2_X1 U16007 ( .A1(b_9_), .A2(n15937), .ZN(n15936) );
  NAND2_X1 U16008 ( .A1(n8424), .A2(a_9_), .ZN(n15937) );
  INV_X1 U16009 ( .A(n8415), .ZN(n8424) );
  NAND2_X1 U16010 ( .A1(n8415), .A2(n8426), .ZN(n15935) );
  INV_X1 U16011 ( .A(a_9_), .ZN(n8426) );
  NAND2_X1 U16012 ( .A1(n15938), .A2(n15939), .ZN(n8415) );
  NAND2_X1 U16013 ( .A1(b_10_), .A2(n15940), .ZN(n15939) );
  NAND2_X1 U16014 ( .A1(n8399), .A2(a_10_), .ZN(n15940) );
  INV_X1 U16015 ( .A(n8390), .ZN(n8399) );
  NAND2_X1 U16016 ( .A1(n8390), .A2(n8761), .ZN(n15938) );
  INV_X1 U16017 ( .A(a_10_), .ZN(n8761) );
  NAND2_X1 U16018 ( .A1(n15941), .A2(n15942), .ZN(n8390) );
  NAND2_X1 U16019 ( .A1(b_11_), .A2(n15943), .ZN(n15942) );
  NAND2_X1 U16020 ( .A1(n8373), .A2(a_11_), .ZN(n15943) );
  INV_X1 U16021 ( .A(n8365), .ZN(n8373) );
  NAND2_X1 U16022 ( .A1(n8365), .A2(n8376), .ZN(n15941) );
  INV_X1 U16023 ( .A(a_11_), .ZN(n8376) );
  NAND2_X1 U16024 ( .A1(n15944), .A2(n15945), .ZN(n8365) );
  NAND2_X1 U16025 ( .A1(b_12_), .A2(n15946), .ZN(n15945) );
  NAND2_X1 U16026 ( .A1(n8349), .A2(a_12_), .ZN(n15946) );
  INV_X1 U16027 ( .A(n8340), .ZN(n8349) );
  NAND2_X1 U16028 ( .A1(n8340), .A2(n8759), .ZN(n15944) );
  INV_X1 U16029 ( .A(a_12_), .ZN(n8759) );
  NAND2_X1 U16030 ( .A1(n15947), .A2(n15948), .ZN(n8340) );
  NAND2_X1 U16031 ( .A1(b_13_), .A2(n15949), .ZN(n15948) );
  NAND2_X1 U16032 ( .A1(n8325), .A2(a_13_), .ZN(n15949) );
  INV_X1 U16033 ( .A(n8316), .ZN(n8325) );
  NAND2_X1 U16034 ( .A1(n8316), .A2(n8310), .ZN(n15947) );
  NAND2_X1 U16035 ( .A1(n15950), .A2(n15951), .ZN(n8316) );
  NAND2_X1 U16036 ( .A1(b_14_), .A2(n15952), .ZN(n15951) );
  NAND2_X1 U16037 ( .A1(n8298), .A2(a_14_), .ZN(n15952) );
  INV_X1 U16038 ( .A(n8290), .ZN(n8298) );
  NAND2_X1 U16039 ( .A1(n8290), .A2(n8757), .ZN(n15950) );
  INV_X1 U16040 ( .A(a_14_), .ZN(n8757) );
  NAND2_X1 U16041 ( .A1(n15953), .A2(n15954), .ZN(n8290) );
  NAND2_X1 U16042 ( .A1(b_15_), .A2(n15955), .ZN(n15954) );
  NAND2_X1 U16043 ( .A1(n8273), .A2(a_15_), .ZN(n15955) );
  INV_X1 U16044 ( .A(n8265), .ZN(n8273) );
  NAND2_X1 U16045 ( .A1(n8265), .A2(n8276), .ZN(n15953) );
  NAND2_X1 U16046 ( .A1(n15956), .A2(n15957), .ZN(n8265) );
  NAND2_X1 U16047 ( .A1(b_16_), .A2(n15958), .ZN(n15957) );
  NAND2_X1 U16048 ( .A1(n8249), .A2(a_16_), .ZN(n15958) );
  INV_X1 U16049 ( .A(n8240), .ZN(n8249) );
  NAND2_X1 U16050 ( .A1(n8240), .A2(n8755), .ZN(n15956) );
  INV_X1 U16051 ( .A(a_16_), .ZN(n8755) );
  NAND2_X1 U16052 ( .A1(n15959), .A2(n15960), .ZN(n8240) );
  NAND2_X1 U16053 ( .A1(b_17_), .A2(n15961), .ZN(n15960) );
  NAND2_X1 U16054 ( .A1(n8225), .A2(a_17_), .ZN(n15961) );
  INV_X1 U16055 ( .A(n8216), .ZN(n8225) );
  NAND2_X1 U16056 ( .A1(n8216), .A2(n8210), .ZN(n15959) );
  NAND2_X1 U16057 ( .A1(n15962), .A2(n15963), .ZN(n8216) );
  NAND2_X1 U16058 ( .A1(b_18_), .A2(n15964), .ZN(n15963) );
  NAND2_X1 U16059 ( .A1(n8193), .A2(a_18_), .ZN(n15964) );
  INV_X1 U16060 ( .A(n8184), .ZN(n8193) );
  NAND2_X1 U16061 ( .A1(n8184), .A2(n8753), .ZN(n15962) );
  NAND2_X1 U16062 ( .A1(n15965), .A2(n15966), .ZN(n8184) );
  NAND2_X1 U16063 ( .A1(b_19_), .A2(n15967), .ZN(n15966) );
  NAND2_X1 U16064 ( .A1(n8168), .A2(a_19_), .ZN(n15967) );
  INV_X1 U16065 ( .A(n8159), .ZN(n8168) );
  NAND2_X1 U16066 ( .A1(n8159), .A2(n8170), .ZN(n15965) );
  NAND2_X1 U16067 ( .A1(n15968), .A2(n15969), .ZN(n8159) );
  NAND2_X1 U16068 ( .A1(b_20_), .A2(n15970), .ZN(n15969) );
  NAND2_X1 U16069 ( .A1(n8143), .A2(a_20_), .ZN(n15970) );
  INV_X1 U16070 ( .A(n8134), .ZN(n8143) );
  NAND2_X1 U16071 ( .A1(n8134), .A2(n8751), .ZN(n15968) );
  NAND2_X1 U16072 ( .A1(n15971), .A2(n15972), .ZN(n8134) );
  NAND2_X1 U16073 ( .A1(b_21_), .A2(n15973), .ZN(n15972) );
  NAND2_X1 U16074 ( .A1(n8108), .A2(a_21_), .ZN(n15973) );
  INV_X1 U16075 ( .A(n8116), .ZN(n8108) );
  NAND2_X1 U16076 ( .A1(n8116), .A2(n8750), .ZN(n15971) );
  NAND2_X1 U16077 ( .A1(n15974), .A2(n15975), .ZN(n8116) );
  NAND2_X1 U16078 ( .A1(b_22_), .A2(n15976), .ZN(n15975) );
  NAND2_X1 U16079 ( .A1(n8092), .A2(a_22_), .ZN(n15976) );
  INV_X1 U16080 ( .A(n8083), .ZN(n8092) );
  NAND2_X1 U16081 ( .A1(n8083), .A2(n8748), .ZN(n15974) );
  INV_X1 U16082 ( .A(a_22_), .ZN(n8748) );
  NAND2_X1 U16083 ( .A1(n15977), .A2(n15978), .ZN(n8083) );
  NAND2_X1 U16084 ( .A1(b_23_), .A2(n15979), .ZN(n15978) );
  NAND2_X1 U16085 ( .A1(n8057), .A2(a_23_), .ZN(n15979) );
  INV_X1 U16086 ( .A(n8065), .ZN(n8057) );
  NAND2_X1 U16087 ( .A1(n8065), .A2(n8747), .ZN(n15977) );
  NAND2_X1 U16088 ( .A1(n15980), .A2(n15981), .ZN(n8065) );
  NAND2_X1 U16089 ( .A1(b_24_), .A2(n15982), .ZN(n15981) );
  NAND2_X1 U16090 ( .A1(n8041), .A2(a_24_), .ZN(n15982) );
  INV_X1 U16091 ( .A(n8032), .ZN(n8041) );
  NAND2_X1 U16092 ( .A1(n8032), .A2(n8745), .ZN(n15980) );
  NAND2_X1 U16093 ( .A1(n15983), .A2(n15984), .ZN(n8032) );
  NAND2_X1 U16094 ( .A1(b_25_), .A2(n15985), .ZN(n15984) );
  NAND2_X1 U16095 ( .A1(n8006), .A2(a_25_), .ZN(n15985) );
  INV_X1 U16096 ( .A(n8014), .ZN(n8006) );
  NAND2_X1 U16097 ( .A1(n8014), .A2(n8744), .ZN(n15983) );
  NAND2_X1 U16098 ( .A1(n15986), .A2(n15987), .ZN(n8014) );
  NAND2_X1 U16099 ( .A1(b_26_), .A2(n15988), .ZN(n15987) );
  NAND2_X1 U16100 ( .A1(n7990), .A2(a_26_), .ZN(n15988) );
  INV_X1 U16101 ( .A(n7981), .ZN(n7990) );
  NAND2_X1 U16102 ( .A1(n7981), .A2(n8742), .ZN(n15986) );
  INV_X1 U16103 ( .A(a_26_), .ZN(n8742) );
  NAND2_X1 U16104 ( .A1(n15989), .A2(n15990), .ZN(n7981) );
  NAND2_X1 U16105 ( .A1(b_27_), .A2(n15991), .ZN(n15990) );
  NAND2_X1 U16106 ( .A1(n7955), .A2(a_27_), .ZN(n15991) );
  INV_X1 U16107 ( .A(n7963), .ZN(n7955) );
  NAND2_X1 U16108 ( .A1(n7963), .A2(n8741), .ZN(n15989) );
  INV_X1 U16109 ( .A(a_27_), .ZN(n8741) );
  NAND2_X1 U16110 ( .A1(n15992), .A2(n15993), .ZN(n7963) );
  NAND2_X1 U16111 ( .A1(b_28_), .A2(n15994), .ZN(n15993) );
  NAND2_X1 U16112 ( .A1(n7933), .A2(a_28_), .ZN(n15994) );
  INV_X1 U16113 ( .A(n7924), .ZN(n7933) );
  NAND2_X1 U16114 ( .A1(n7924), .A2(n8739), .ZN(n15992) );
  INV_X1 U16115 ( .A(a_28_), .ZN(n8739) );
  NAND2_X1 U16116 ( .A1(n15995), .A2(n15996), .ZN(n7924) );
  NAND2_X1 U16117 ( .A1(b_29_), .A2(n15997), .ZN(n15996) );
  NAND2_X1 U16118 ( .A1(n7898), .A2(a_29_), .ZN(n15997) );
  INV_X1 U16119 ( .A(n7906), .ZN(n7898) );
  NAND2_X1 U16120 ( .A1(n7906), .A2(n7890), .ZN(n15995) );
  NAND2_X1 U16121 ( .A1(n15998), .A2(n15999), .ZN(n7906) );
  NAND2_X1 U16122 ( .A1(b_30_), .A2(n16000), .ZN(n15999) );
  NAND2_X1 U16123 ( .A1(n7875), .A2(a_30_), .ZN(n16000) );
  INV_X1 U16124 ( .A(n7854), .ZN(n7875) );
  NAND2_X1 U16125 ( .A1(n7854), .A2(n7867), .ZN(n15998) );
  INV_X1 U16126 ( .A(a_30_), .ZN(n7867) );
  NAND2_X1 U16127 ( .A1(a_31_), .A2(n7889), .ZN(n7854) );
  INV_X1 U16128 ( .A(b_31_), .ZN(n7889) );
endmodule

