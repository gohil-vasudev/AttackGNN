module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n614_, new_n445_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n421_, new_n620_, new_n368_, new_n439_, new_n283_, new_n223_, new_n366_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n197_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n636_, new_n456_, new_n246_, new_n170_, new_n266_, new_n367_, new_n542_, new_n548_, new_n173_, new_n220_, new_n419_, new_n624_, new_n534_, new_n214_, new_n451_, new_n489_, new_n424_, new_n602_, new_n188_, new_n240_, new_n413_, new_n526_, new_n442_, new_n642_, new_n211_, new_n552_, new_n342_, new_n462_, new_n603_, new_n564_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n626_, new_n152_, new_n157_, new_n153_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n272_, new_n282_, new_n201_, new_n192_, new_n414_, new_n635_, new_n315_, new_n326_, new_n554_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n630_, new_n167_, new_n385_, new_n478_, new_n461_, new_n297_, new_n361_, new_n565_, new_n150_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n629_, new_n321_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n549_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n506_, new_n256_, new_n452_, new_n381_, new_n508_, new_n194_, new_n483_, new_n394_, new_n299_, new_n142_, new_n139_, new_n314_, new_n582_, new_n363_, new_n165_, new_n441_, new_n477_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n301_, new_n169_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n187_, new_n311_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n579_, new_n286_, new_n335_, new_n347_, new_n346_, new_n198_, new_n438_, new_n208_, new_n632_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n399_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n166_, new_n162_, new_n457_, new_n161_, new_n553_, new_n333_, new_n290_, new_n448_, new_n276_, new_n155_, new_n410_, new_n543_, new_n454_, new_n202_, new_n296_, new_n308_, new_n633_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n309_, new_n529_, new_n323_, new_n259_, new_n362_, new_n604_, new_n227_, new_n416_, new_n222_, new_n571_, new_n328_, new_n460_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n138_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n562_, new_n578_, new_n177_, new_n493_, new_n547_, new_n264_, new_n379_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n143_, new_n520_, new_n145_, new_n253_, new_n403_, new_n475_, new_n237_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n507_, new_n182_, new_n480_, new_n625_, new_n151_, new_n513_, new_n592_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n522_, new_n588_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n546_, new_n612_, new_n302_, new_n191_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n154_, new_n255_, new_n533_, new_n459_, new_n555_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n147_, new_n285_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n591_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n563_, new_n148_, new_n440_, new_n531_, new_n593_, new_n252_, new_n585_, new_n160_, new_n312_, new_n535_, new_n372_, new_n242_, new_n503_, new_n527_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n433_, new_n435_, new_n265_, new_n370_, new_n584_, new_n278_, new_n304_, new_n523_, new_n638_, new_n550_, new_n217_, new_n269_, new_n512_, new_n599_, new_n412_, new_n607_, new_n327_, new_n594_, new_n561_, new_n495_, new_n431_, new_n196_, new_n574_, new_n319_, new_n640_, new_n338_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n294_, new_n627_, new_n195_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n474_, new_n467_, new_n404_, new_n193_, new_n560_, new_n358_, new_n348_, new_n610_, new_n159_, new_n322_, new_n228_, new_n545_, new_n611_, new_n289_, new_n425_, new_n175_, new_n226_, new_n185_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n168_, new_n279_, new_n455_, new_n618_, new_n521_, new_n406_, new_n356_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n573_;

xnor g000 ( new_n138_, N65, N69 );
xnor g001 ( new_n139_, N73, N77 );
xnor g002 ( new_n140_, new_n138_, new_n139_ );
xnor g003 ( new_n141_, N81, N85 );
xnor g004 ( new_n142_, N89, N93 );
xnor g005 ( new_n143_, new_n141_, new_n142_ );
xnor g006 ( new_n144_, new_n140_, new_n143_ );
nand g007 ( new_n145_, N129, N137 );
xnor g008 ( new_n146_, new_n144_, new_n145_ );
xor g009 ( new_n147_, N1, N17 );
xnor g010 ( new_n148_, N33, N49 );
xnor g011 ( new_n149_, new_n147_, new_n148_ );
xnor g012 ( new_n150_, new_n146_, new_n149_ );
not g013 ( new_n151_, keyIn_0_0 );
xnor g014 ( new_n152_, N1, N5 );
nand g015 ( new_n153_, new_n152_, new_n151_ );
nand g016 ( new_n154_, N1, N5 );
nor g017 ( new_n155_, N1, N5 );
nor g018 ( new_n156_, new_n155_, new_n151_ );
nand g019 ( new_n157_, new_n156_, new_n154_ );
nand g020 ( new_n158_, new_n153_, new_n157_ );
not g021 ( new_n159_, keyIn_0_1 );
not g022 ( new_n160_, N13 );
nand g023 ( new_n161_, new_n160_, N9 );
not g024 ( new_n162_, N9 );
nand g025 ( new_n163_, new_n162_, N13 );
nand g026 ( new_n164_, new_n161_, new_n163_ );
nand g027 ( new_n165_, new_n164_, new_n159_ );
xnor g028 ( new_n166_, N9, N13 );
nand g029 ( new_n167_, new_n166_, keyIn_0_1 );
nand g030 ( new_n168_, new_n165_, new_n167_ );
xnor g031 ( new_n169_, new_n168_, new_n158_ );
nand g032 ( new_n170_, new_n169_, keyIn_0_12 );
not g033 ( new_n171_, keyIn_0_12 );
and g034 ( new_n172_, new_n168_, new_n158_ );
nor g035 ( new_n173_, new_n168_, new_n158_ );
nor g036 ( new_n174_, new_n172_, new_n173_ );
nand g037 ( new_n175_, new_n174_, new_n171_ );
nand g038 ( new_n176_, new_n175_, new_n170_ );
xnor g039 ( new_n177_, N41, N45 );
nand g040 ( new_n178_, new_n177_, keyIn_0_5 );
nand g041 ( new_n179_, N41, N45 );
nor g042 ( new_n180_, N41, N45 );
nor g043 ( new_n181_, new_n180_, keyIn_0_5 );
nand g044 ( new_n182_, new_n181_, new_n179_ );
nand g045 ( new_n183_, new_n178_, new_n182_ );
xnor g046 ( new_n184_, N33, N37 );
nand g047 ( new_n185_, new_n184_, keyIn_0_4 );
nand g048 ( new_n186_, N33, N37 );
nor g049 ( new_n187_, N33, N37 );
nor g050 ( new_n188_, new_n187_, keyIn_0_4 );
nand g051 ( new_n189_, new_n188_, new_n186_ );
nand g052 ( new_n190_, new_n185_, new_n189_ );
xnor g053 ( new_n191_, new_n183_, new_n190_ );
nand g054 ( new_n192_, new_n191_, keyIn_0_14 );
not g055 ( new_n193_, keyIn_0_14 );
and g056 ( new_n194_, new_n183_, new_n190_ );
nor g057 ( new_n195_, new_n183_, new_n190_ );
nor g058 ( new_n196_, new_n194_, new_n195_ );
nand g059 ( new_n197_, new_n196_, new_n193_ );
and g060 ( new_n198_, new_n197_, new_n192_ );
nand g061 ( new_n199_, new_n198_, new_n176_ );
xnor g062 ( new_n200_, new_n169_, new_n171_ );
nand g063 ( new_n201_, new_n197_, new_n192_ );
nand g064 ( new_n202_, new_n200_, new_n201_ );
nand g065 ( new_n203_, new_n199_, new_n202_ );
nand g066 ( new_n204_, new_n203_, keyIn_0_19 );
not g067 ( new_n205_, keyIn_0_19 );
xnor g068 ( new_n206_, new_n176_, new_n201_ );
nand g069 ( new_n207_, new_n206_, new_n205_ );
nand g070 ( new_n208_, new_n207_, new_n204_ );
and g071 ( new_n209_, N135, N137 );
or g072 ( new_n210_, new_n209_, keyIn_0_7 );
not g073 ( new_n211_, new_n210_ );
not g074 ( new_n212_, N137 );
nand g075 ( new_n213_, keyIn_0_7, N135 );
nor g076 ( new_n214_, new_n213_, new_n212_ );
nor g077 ( new_n215_, new_n211_, new_n214_ );
not g078 ( new_n216_, new_n215_ );
nand g079 ( new_n217_, new_n208_, new_n216_ );
xnor g080 ( new_n218_, new_n203_, new_n205_ );
nand g081 ( new_n219_, new_n218_, new_n215_ );
nand g082 ( new_n220_, new_n219_, new_n217_ );
nand g083 ( new_n221_, new_n220_, keyIn_0_21 );
not g084 ( new_n222_, keyIn_0_21 );
xnor g085 ( new_n223_, new_n208_, new_n215_ );
nand g086 ( new_n224_, new_n223_, new_n222_ );
nand g087 ( new_n225_, new_n224_, new_n221_ );
xnor g088 ( new_n226_, N105, N121 );
xnor g089 ( new_n227_, new_n226_, keyIn_0_11 );
xor g090 ( new_n228_, N73, N89 );
xnor g091 ( new_n229_, new_n228_, keyIn_0_10 );
xnor g092 ( new_n230_, new_n229_, new_n227_ );
xor g093 ( new_n231_, new_n230_, keyIn_0_17 );
nand g094 ( new_n232_, new_n225_, new_n231_ );
xnor g095 ( new_n233_, new_n220_, new_n222_ );
not g096 ( new_n234_, new_n231_ );
nand g097 ( new_n235_, new_n233_, new_n234_ );
nand g098 ( new_n236_, new_n235_, new_n232_ );
xnor g099 ( new_n237_, new_n236_, keyIn_0_23 );
not g100 ( new_n238_, keyIn_0_13 );
not g101 ( new_n239_, N29 );
nand g102 ( new_n240_, new_n239_, N25 );
not g103 ( new_n241_, N25 );
nand g104 ( new_n242_, new_n241_, N29 );
nand g105 ( new_n243_, new_n240_, new_n242_ );
nand g106 ( new_n244_, new_n243_, keyIn_0_3 );
not g107 ( new_n245_, keyIn_0_3 );
xnor g108 ( new_n246_, N25, N29 );
nand g109 ( new_n247_, new_n246_, new_n245_ );
nand g110 ( new_n248_, new_n244_, new_n247_ );
xnor g111 ( new_n249_, N17, N21 );
nand g112 ( new_n250_, new_n249_, keyIn_0_2 );
nand g113 ( new_n251_, N17, N21 );
nor g114 ( new_n252_, N17, N21 );
nor g115 ( new_n253_, new_n252_, keyIn_0_2 );
nand g116 ( new_n254_, new_n253_, new_n251_ );
nand g117 ( new_n255_, new_n250_, new_n254_ );
nand g118 ( new_n256_, new_n248_, new_n255_ );
and g119 ( new_n257_, new_n244_, new_n247_ );
and g120 ( new_n258_, new_n250_, new_n254_ );
nand g121 ( new_n259_, new_n257_, new_n258_ );
nand g122 ( new_n260_, new_n259_, new_n256_ );
xnor g123 ( new_n261_, new_n260_, new_n238_ );
xor g124 ( new_n262_, N49, N53 );
xnor g125 ( new_n263_, N57, N61 );
xnor g126 ( new_n264_, new_n262_, new_n263_ );
xnor g127 ( new_n265_, new_n261_, new_n264_ );
nand g128 ( new_n266_, N136, N137 );
xnor g129 ( new_n267_, new_n265_, new_n266_ );
xnor g130 ( new_n268_, N77, N93 );
xnor g131 ( new_n269_, N109, N125 );
xnor g132 ( new_n270_, new_n268_, new_n269_ );
xnor g133 ( new_n271_, new_n267_, new_n270_ );
xnor g134 ( new_n272_, N97, N101 );
xnor g135 ( new_n273_, N105, N109 );
xnor g136 ( new_n274_, new_n272_, new_n273_ );
xnor g137 ( new_n275_, new_n140_, new_n274_ );
nand g138 ( new_n276_, N131, N137 );
xnor g139 ( new_n277_, new_n275_, new_n276_ );
xor g140 ( new_n278_, N9, N25 );
xnor g141 ( new_n279_, N41, N57 );
xnor g142 ( new_n280_, new_n278_, new_n279_ );
xnor g143 ( new_n281_, new_n277_, new_n280_ );
and g144 ( new_n282_, new_n281_, keyIn_0_24 );
nand g145 ( new_n283_, new_n282_, new_n150_ );
xnor g146 ( new_n284_, N113, N117 );
xnor g147 ( new_n285_, N121, N125 );
xnor g148 ( new_n286_, new_n284_, new_n285_ );
xnor g149 ( new_n287_, new_n274_, new_n286_ );
nand g150 ( new_n288_, N130, N137 );
xnor g151 ( new_n289_, new_n287_, new_n288_ );
xor g152 ( new_n290_, N5, N21 );
xnor g153 ( new_n291_, N37, N53 );
xnor g154 ( new_n292_, new_n290_, new_n291_ );
xnor g155 ( new_n293_, new_n289_, new_n292_ );
nor g156 ( new_n294_, new_n282_, new_n150_ );
nor g157 ( new_n295_, new_n294_, new_n293_ );
nand g158 ( new_n296_, new_n295_, new_n283_ );
not g159 ( new_n297_, new_n293_ );
nor g160 ( new_n298_, new_n297_, new_n150_ );
not g161 ( new_n299_, new_n298_ );
or g162 ( new_n300_, new_n299_, new_n281_ );
nand g163 ( new_n301_, new_n296_, new_n300_ );
xnor g164 ( new_n302_, new_n143_, new_n286_ );
nand g165 ( new_n303_, N132, N137 );
xnor g166 ( new_n304_, new_n302_, new_n303_ );
xor g167 ( new_n305_, N13, N29 );
xnor g168 ( new_n306_, N45, N61 );
xnor g169 ( new_n307_, new_n305_, new_n306_ );
xnor g170 ( new_n308_, new_n307_, keyIn_0_15 );
xnor g171 ( new_n309_, new_n304_, new_n308_ );
not g172 ( new_n310_, new_n309_ );
nand g173 ( new_n311_, new_n301_, new_n310_ );
nor g174 ( new_n312_, new_n150_, new_n293_ );
nor g175 ( new_n313_, new_n310_, new_n281_ );
nand g176 ( new_n314_, new_n313_, new_n312_ );
nand g177 ( new_n315_, new_n311_, new_n314_ );
nand g178 ( new_n316_, new_n315_, new_n271_ );
nor g179 ( new_n317_, new_n237_, new_n316_ );
not g180 ( new_n318_, new_n317_ );
not g181 ( new_n319_, keyIn_0_22 );
not g182 ( new_n320_, keyIn_0_20 );
nand g183 ( new_n321_, new_n261_, new_n176_ );
xnor g184 ( new_n322_, new_n260_, keyIn_0_13 );
nand g185 ( new_n323_, new_n200_, new_n322_ );
nand g186 ( new_n324_, new_n323_, new_n321_ );
nand g187 ( new_n325_, new_n324_, keyIn_0_18 );
not g188 ( new_n326_, keyIn_0_18 );
xnor g189 ( new_n327_, new_n322_, new_n176_ );
nand g190 ( new_n328_, new_n327_, new_n326_ );
nand g191 ( new_n329_, new_n328_, new_n325_ );
and g192 ( new_n330_, N133, N137 );
or g193 ( new_n331_, new_n330_, keyIn_0_6 );
not g194 ( new_n332_, new_n331_ );
nand g195 ( new_n333_, keyIn_0_6, N133 );
nor g196 ( new_n334_, new_n333_, new_n212_ );
nor g197 ( new_n335_, new_n332_, new_n334_ );
nand g198 ( new_n336_, new_n329_, new_n335_ );
xnor g199 ( new_n337_, new_n324_, new_n326_ );
not g200 ( new_n338_, new_n335_ );
nand g201 ( new_n339_, new_n337_, new_n338_ );
nand g202 ( new_n340_, new_n339_, new_n336_ );
nand g203 ( new_n341_, new_n340_, new_n320_ );
xnor g204 ( new_n342_, new_n329_, new_n338_ );
nand g205 ( new_n343_, new_n342_, keyIn_0_20 );
nand g206 ( new_n344_, new_n343_, new_n341_ );
xor g207 ( new_n345_, N65, N81 );
xnor g208 ( new_n346_, new_n345_, keyIn_0_8 );
xor g209 ( new_n347_, N97, N113 );
xnor g210 ( new_n348_, new_n347_, keyIn_0_9 );
xnor g211 ( new_n349_, new_n346_, new_n348_ );
xnor g212 ( new_n350_, new_n349_, keyIn_0_16 );
nand g213 ( new_n351_, new_n344_, new_n350_ );
xnor g214 ( new_n352_, new_n340_, keyIn_0_20 );
not g215 ( new_n353_, new_n350_ );
nand g216 ( new_n354_, new_n352_, new_n353_ );
nand g217 ( new_n355_, new_n354_, new_n351_ );
xnor g218 ( new_n356_, new_n355_, new_n319_ );
xnor g219 ( new_n357_, new_n198_, new_n264_ );
nand g220 ( new_n358_, N134, N137 );
xnor g221 ( new_n359_, new_n357_, new_n358_ );
xnor g222 ( new_n360_, N69, N85 );
xnor g223 ( new_n361_, N101, N117 );
xnor g224 ( new_n362_, new_n360_, new_n361_ );
xnor g225 ( new_n363_, new_n359_, new_n362_ );
not g226 ( new_n364_, new_n363_ );
nor g227 ( new_n365_, new_n356_, new_n364_ );
not g228 ( new_n366_, new_n365_ );
nor g229 ( new_n367_, new_n318_, new_n366_ );
nand g230 ( new_n368_, new_n367_, new_n150_ );
xnor g231 ( N724, new_n368_, N1 );
nand g232 ( new_n370_, new_n367_, new_n293_ );
xnor g233 ( N725, new_n370_, N5 );
nand g234 ( new_n372_, new_n367_, new_n281_ );
xnor g235 ( N726, new_n372_, N9 );
nand g236 ( new_n374_, new_n367_, new_n309_ );
xnor g237 ( N727, new_n374_, N13 );
not g238 ( new_n376_, keyIn_0_23 );
xnor g239 ( new_n377_, new_n236_, new_n376_ );
not g240 ( new_n378_, new_n271_ );
nand g241 ( new_n379_, new_n315_, new_n378_ );
nor g242 ( new_n380_, new_n377_, new_n379_ );
not g243 ( new_n381_, new_n380_ );
nor g244 ( new_n382_, new_n381_, new_n366_ );
nand g245 ( new_n383_, new_n382_, new_n150_ );
xnor g246 ( N728, new_n383_, N17 );
nand g247 ( new_n385_, new_n382_, new_n293_ );
xnor g248 ( N729, new_n385_, N21 );
nand g249 ( new_n387_, new_n382_, new_n281_ );
xnor g250 ( N730, new_n387_, N25 );
nand g251 ( new_n389_, new_n382_, new_n309_ );
xnor g252 ( N731, new_n389_, N29 );
xnor g253 ( new_n391_, new_n355_, keyIn_0_22 );
nor g254 ( new_n392_, new_n391_, new_n363_ );
not g255 ( new_n393_, new_n392_ );
nor g256 ( new_n394_, new_n318_, new_n393_ );
nand g257 ( new_n395_, new_n394_, new_n150_ );
xnor g258 ( N732, new_n395_, N33 );
nand g259 ( new_n397_, new_n394_, new_n293_ );
xnor g260 ( N733, new_n397_, N37 );
nand g261 ( new_n399_, new_n394_, new_n281_ );
xnor g262 ( N734, new_n399_, N41 );
nand g263 ( new_n401_, new_n394_, new_n309_ );
xnor g264 ( N735, new_n401_, N45 );
nor g265 ( new_n403_, new_n381_, new_n393_ );
nand g266 ( new_n404_, new_n403_, new_n150_ );
xnor g267 ( N736, new_n404_, N49 );
nand g268 ( new_n406_, new_n403_, new_n293_ );
xnor g269 ( N737, new_n406_, N53 );
nand g270 ( new_n408_, new_n403_, new_n281_ );
xnor g271 ( N738, new_n408_, N57 );
nand g272 ( new_n410_, new_n403_, new_n309_ );
xnor g273 ( N739, new_n410_, N61 );
not g274 ( new_n412_, keyIn_0_40 );
xnor g275 ( new_n413_, new_n377_, keyIn_0_27 );
nor g276 ( new_n414_, new_n356_, keyIn_0_25 );
nand g277 ( new_n415_, new_n356_, keyIn_0_25 );
nor g278 ( new_n416_, new_n364_, keyIn_0_26 );
nand g279 ( new_n417_, new_n364_, keyIn_0_26 );
nand g280 ( new_n418_, new_n417_, new_n378_ );
nor g281 ( new_n419_, new_n418_, new_n416_ );
nand g282 ( new_n420_, new_n415_, new_n419_ );
nor g283 ( new_n421_, new_n420_, new_n414_ );
nand g284 ( new_n422_, new_n421_, new_n413_ );
xnor g285 ( new_n423_, new_n422_, keyIn_0_32 );
not g286 ( new_n424_, keyIn_0_34 );
xnor g287 ( new_n425_, new_n356_, keyIn_0_29 );
not g288 ( new_n426_, keyIn_0_30 );
nor g289 ( new_n427_, new_n237_, new_n426_ );
nand g290 ( new_n428_, new_n237_, new_n426_ );
nor g291 ( new_n429_, new_n378_, new_n363_ );
nand g292 ( new_n430_, new_n428_, new_n429_ );
nor g293 ( new_n431_, new_n430_, new_n427_ );
nand g294 ( new_n432_, new_n431_, new_n425_ );
nor g295 ( new_n433_, new_n432_, new_n424_ );
not g296 ( new_n434_, keyIn_0_31 );
nor g297 ( new_n435_, new_n237_, new_n434_ );
not g298 ( new_n436_, new_n435_ );
nor g299 ( new_n437_, new_n377_, keyIn_0_31 );
nor g300 ( new_n438_, new_n364_, new_n378_ );
nand g301 ( new_n439_, new_n391_, new_n438_ );
nor g302 ( new_n440_, new_n437_, new_n439_ );
nand g303 ( new_n441_, new_n440_, new_n436_ );
nand g304 ( new_n442_, new_n441_, keyIn_0_35 );
not g305 ( new_n443_, keyIn_0_35 );
nand g306 ( new_n444_, new_n237_, new_n434_ );
not g307 ( new_n445_, new_n438_ );
nor g308 ( new_n446_, new_n356_, new_n445_ );
nand g309 ( new_n447_, new_n446_, new_n444_ );
nor g310 ( new_n448_, new_n447_, new_n435_ );
nand g311 ( new_n449_, new_n448_, new_n443_ );
nand g312 ( new_n450_, new_n442_, new_n449_ );
nand g313 ( new_n451_, new_n432_, new_n424_ );
nand g314 ( new_n452_, new_n450_, new_n451_ );
nor g315 ( new_n453_, new_n452_, new_n433_ );
nand g316 ( new_n454_, new_n453_, new_n423_ );
not g317 ( new_n455_, keyIn_0_36 );
nor g318 ( new_n456_, new_n391_, keyIn_0_28 );
nand g319 ( new_n457_, new_n391_, keyIn_0_28 );
nor g320 ( new_n458_, new_n237_, new_n445_ );
nand g321 ( new_n459_, new_n458_, new_n457_ );
nor g322 ( new_n460_, new_n459_, new_n456_ );
xnor g323 ( new_n461_, new_n460_, keyIn_0_33 );
nand g324 ( new_n462_, new_n461_, new_n455_ );
nor g325 ( new_n463_, new_n454_, new_n462_ );
not g326 ( new_n464_, new_n463_ );
and g327 ( new_n465_, new_n453_, new_n423_ );
nor g328 ( new_n466_, new_n460_, keyIn_0_33 );
and g329 ( new_n467_, new_n438_, keyIn_0_33 );
nand g330 ( new_n468_, new_n377_, new_n467_ );
not g331 ( new_n469_, new_n468_ );
nand g332 ( new_n470_, new_n469_, new_n457_ );
nor g333 ( new_n471_, new_n470_, new_n456_ );
nor g334 ( new_n472_, new_n466_, new_n471_ );
not g335 ( new_n473_, new_n472_ );
nand g336 ( new_n474_, new_n465_, new_n473_ );
nand g337 ( new_n475_, new_n474_, keyIn_0_36 );
nand g338 ( new_n476_, new_n475_, new_n464_ );
nand g339 ( new_n477_, new_n310_, new_n281_ );
nand g340 ( new_n478_, new_n297_, new_n150_ );
nor g341 ( new_n479_, new_n477_, new_n478_ );
nand g342 ( new_n480_, new_n476_, new_n479_ );
xnor g343 ( new_n481_, new_n480_, keyIn_0_37 );
nand g344 ( new_n482_, new_n481_, new_n391_ );
xnor g345 ( new_n483_, new_n482_, new_n412_ );
xnor g346 ( new_n484_, new_n483_, N65 );
nand g347 ( new_n485_, new_n484_, keyIn_0_52 );
not g348 ( new_n486_, keyIn_0_52 );
not g349 ( new_n487_, N65 );
xnor g350 ( new_n488_, new_n483_, new_n487_ );
nand g351 ( new_n489_, new_n488_, new_n486_ );
nand g352 ( N740, new_n485_, new_n489_ );
not g353 ( new_n491_, keyIn_0_53 );
nand g354 ( new_n492_, new_n481_, new_n364_ );
xnor g355 ( new_n493_, new_n492_, keyIn_0_41 );
xnor g356 ( new_n494_, new_n493_, N69 );
nand g357 ( new_n495_, new_n494_, new_n491_ );
not g358 ( new_n496_, N69 );
xnor g359 ( new_n497_, new_n493_, new_n496_ );
nand g360 ( new_n498_, new_n497_, keyIn_0_53 );
nand g361 ( N741, new_n495_, new_n498_ );
not g362 ( new_n500_, keyIn_0_42 );
nand g363 ( new_n501_, new_n481_, new_n377_ );
xnor g364 ( new_n502_, new_n501_, new_n500_ );
xnor g365 ( new_n503_, new_n502_, N73 );
nand g366 ( new_n504_, new_n503_, keyIn_0_54 );
not g367 ( new_n505_, keyIn_0_54 );
not g368 ( new_n506_, N73 );
xnor g369 ( new_n507_, new_n502_, new_n506_ );
nand g370 ( new_n508_, new_n507_, new_n505_ );
nand g371 ( N742, new_n504_, new_n508_ );
not g372 ( new_n510_, keyIn_0_43 );
nand g373 ( new_n511_, new_n481_, new_n378_ );
xnor g374 ( new_n512_, new_n511_, new_n510_ );
xnor g375 ( new_n513_, new_n512_, N77 );
nand g376 ( new_n514_, new_n513_, keyIn_0_55 );
not g377 ( new_n515_, keyIn_0_55 );
not g378 ( new_n516_, N77 );
xnor g379 ( new_n517_, new_n512_, new_n516_ );
nand g380 ( new_n518_, new_n517_, new_n515_ );
nand g381 ( N743, new_n514_, new_n518_ );
nor g382 ( new_n520_, new_n454_, new_n472_ );
nor g383 ( new_n521_, new_n520_, new_n455_ );
nor g384 ( new_n522_, new_n521_, new_n463_ );
nor g385 ( new_n523_, new_n522_, new_n310_ );
nor g386 ( new_n524_, new_n478_, new_n281_ );
nand g387 ( new_n525_, new_n523_, new_n524_ );
nor g388 ( new_n526_, new_n525_, keyIn_0_38 );
not g389 ( new_n527_, new_n526_ );
not g390 ( new_n528_, keyIn_0_38 );
nand g391 ( new_n529_, new_n476_, new_n309_ );
not g392 ( new_n530_, new_n524_ );
nor g393 ( new_n531_, new_n529_, new_n530_ );
nor g394 ( new_n532_, new_n531_, new_n528_ );
nor g395 ( new_n533_, new_n532_, new_n356_ );
nand g396 ( new_n534_, new_n533_, new_n527_ );
nand g397 ( new_n535_, new_n534_, keyIn_0_44 );
not g398 ( new_n536_, keyIn_0_44 );
nand g399 ( new_n537_, new_n525_, keyIn_0_38 );
nand g400 ( new_n538_, new_n537_, new_n391_ );
nor g401 ( new_n539_, new_n538_, new_n526_ );
nand g402 ( new_n540_, new_n539_, new_n536_ );
nand g403 ( new_n541_, new_n535_, new_n540_ );
nand g404 ( new_n542_, new_n541_, N81 );
not g405 ( new_n543_, N81 );
xnor g406 ( new_n544_, new_n539_, keyIn_0_44 );
nand g407 ( new_n545_, new_n544_, new_n543_ );
nand g408 ( new_n546_, new_n545_, new_n542_ );
nand g409 ( new_n547_, new_n546_, keyIn_0_56 );
not g410 ( new_n548_, keyIn_0_56 );
xnor g411 ( new_n549_, new_n541_, new_n543_ );
nand g412 ( new_n550_, new_n549_, new_n548_ );
nand g413 ( N744, new_n550_, new_n547_ );
not g414 ( new_n552_, keyIn_0_45 );
nor g415 ( new_n553_, new_n532_, new_n363_ );
nand g416 ( new_n554_, new_n553_, new_n527_ );
nand g417 ( new_n555_, new_n554_, new_n552_ );
nand g418 ( new_n556_, new_n537_, new_n364_ );
nor g419 ( new_n557_, new_n556_, new_n526_ );
nand g420 ( new_n558_, new_n557_, keyIn_0_45 );
nand g421 ( new_n559_, new_n555_, new_n558_ );
nand g422 ( new_n560_, new_n559_, N85 );
not g423 ( new_n561_, N85 );
xnor g424 ( new_n562_, new_n557_, new_n552_ );
nand g425 ( new_n563_, new_n562_, new_n561_ );
nand g426 ( new_n564_, new_n563_, new_n560_ );
nand g427 ( new_n565_, new_n564_, keyIn_0_57 );
not g428 ( new_n566_, keyIn_0_57 );
xnor g429 ( new_n567_, new_n559_, new_n561_ );
nand g430 ( new_n568_, new_n567_, new_n566_ );
nand g431 ( N745, new_n568_, new_n565_ );
not g432 ( new_n570_, N89 );
not g433 ( new_n571_, keyIn_0_46 );
nor g434 ( new_n572_, new_n532_, new_n237_ );
nand g435 ( new_n573_, new_n572_, new_n527_ );
nand g436 ( new_n574_, new_n573_, new_n571_ );
nand g437 ( new_n575_, new_n537_, new_n377_ );
nor g438 ( new_n576_, new_n575_, new_n526_ );
nand g439 ( new_n577_, new_n576_, keyIn_0_46 );
nand g440 ( new_n578_, new_n574_, new_n577_ );
nand g441 ( new_n579_, new_n578_, new_n570_ );
xnor g442 ( new_n580_, new_n576_, new_n571_ );
nand g443 ( new_n581_, new_n580_, N89 );
nand g444 ( new_n582_, new_n581_, new_n579_ );
nand g445 ( new_n583_, new_n582_, keyIn_0_58 );
not g446 ( new_n584_, keyIn_0_58 );
xnor g447 ( new_n585_, new_n578_, N89 );
nand g448 ( new_n586_, new_n585_, new_n584_ );
nand g449 ( N746, new_n586_, new_n583_ );
not g450 ( new_n588_, keyIn_0_47 );
nor g451 ( new_n589_, new_n532_, new_n271_ );
nand g452 ( new_n590_, new_n589_, new_n527_ );
nand g453 ( new_n591_, new_n590_, new_n588_ );
nand g454 ( new_n592_, new_n537_, new_n378_ );
nor g455 ( new_n593_, new_n592_, new_n526_ );
nand g456 ( new_n594_, new_n593_, keyIn_0_47 );
nand g457 ( new_n595_, new_n591_, new_n594_ );
nand g458 ( new_n596_, new_n595_, N93 );
not g459 ( new_n597_, N93 );
xnor g460 ( new_n598_, new_n593_, new_n588_ );
nand g461 ( new_n599_, new_n598_, new_n597_ );
nand g462 ( new_n600_, new_n599_, new_n596_ );
nand g463 ( new_n601_, new_n600_, keyIn_0_59 );
not g464 ( new_n602_, keyIn_0_59 );
xnor g465 ( new_n603_, new_n595_, new_n597_ );
nand g466 ( new_n604_, new_n603_, new_n602_ );
nand g467 ( N747, new_n604_, new_n601_ );
not g468 ( new_n606_, keyIn_0_60 );
not g469 ( new_n607_, keyIn_0_39 );
nor g470 ( new_n608_, new_n299_, new_n477_ );
nand g471 ( new_n609_, new_n476_, new_n608_ );
nor g472 ( new_n610_, new_n609_, new_n607_ );
nand g473 ( new_n611_, new_n609_, new_n607_ );
nand g474 ( new_n612_, new_n611_, new_n391_ );
nor g475 ( new_n613_, new_n612_, new_n610_ );
xnor g476 ( new_n614_, new_n613_, keyIn_0_48 );
xnor g477 ( new_n615_, new_n614_, N97 );
xnor g478 ( N748, new_n615_, new_n606_ );
not g479 ( new_n617_, keyIn_0_61 );
nand g480 ( new_n618_, new_n611_, new_n364_ );
nor g481 ( new_n619_, new_n618_, new_n610_ );
xnor g482 ( new_n620_, new_n619_, keyIn_0_49 );
xnor g483 ( new_n621_, new_n620_, N101 );
xnor g484 ( N749, new_n621_, new_n617_ );
not g485 ( new_n623_, keyIn_0_62 );
nand g486 ( new_n624_, new_n611_, new_n377_ );
nor g487 ( new_n625_, new_n624_, new_n610_ );
xnor g488 ( new_n626_, new_n625_, keyIn_0_50 );
xnor g489 ( new_n627_, new_n626_, N105 );
xnor g490 ( N750, new_n627_, new_n623_ );
not g491 ( new_n629_, N109 );
nand g492 ( new_n630_, new_n611_, new_n378_ );
nor g493 ( new_n631_, new_n630_, new_n610_ );
xnor g494 ( new_n632_, new_n631_, keyIn_0_51 );
xnor g495 ( new_n633_, new_n632_, new_n629_ );
xnor g496 ( N751, new_n633_, keyIn_0_63 );
nor g497 ( new_n635_, new_n529_, new_n300_ );
nand g498 ( new_n636_, new_n635_, new_n391_ );
xnor g499 ( N752, new_n636_, N113 );
nand g500 ( new_n638_, new_n635_, new_n364_ );
xnor g501 ( N753, new_n638_, N117 );
nand g502 ( new_n640_, new_n635_, new_n377_ );
xnor g503 ( N754, new_n640_, N121 );
nand g504 ( new_n642_, new_n635_, new_n378_ );
xnor g505 ( N755, new_n642_, N125 );
endmodule