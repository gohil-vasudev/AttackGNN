module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n445_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n288_, new_n421_, new_n620_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n566_, new_n339_, new_n365_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n456_, new_n246_, new_n266_, new_n367_, new_n542_, new_n548_, new_n220_, new_n419_, new_n624_, new_n534_, new_n214_, new_n451_, new_n489_, new_n424_, new_n240_, new_n413_, new_n526_, new_n442_, new_n211_, new_n552_, new_n342_, new_n462_, new_n603_, new_n564_, new_n500_, new_n317_, new_n344_, new_n287_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n257_, new_n212_, new_n364_, new_n449_, new_n580_, new_n272_, new_n282_, new_n414_, new_n315_, new_n326_, new_n554_, new_n230_, new_n281_, new_n430_, new_n482_, new_n589_, new_n248_, new_n350_, new_n630_, new_n385_, new_n461_, new_n297_, new_n361_, new_n565_, new_n511_, new_n463_, new_n303_, new_n351_, new_n325_, new_n609_, new_n530_, new_n318_, new_n622_, new_n321_, new_n443_, new_n324_, new_n486_, new_n491_, new_n549_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n498_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n506_, new_n256_, new_n452_, new_n381_, new_n388_, new_n508_, new_n483_, new_n394_, new_n299_, new_n314_, new_n582_, new_n363_, new_n441_, new_n477_, new_n216_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n488_, new_n524_, new_n277_, new_n402_, new_n579_, new_n286_, new_n335_, new_n347_, new_n346_, new_n396_, new_n438_, new_n208_, new_n528_, new_n572_, new_n436_, new_n397_, new_n399_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n437_, new_n295_, new_n359_, new_n628_, new_n409_, new_n457_, new_n553_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n384_, new_n410_, new_n543_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n308_, new_n232_, new_n258_, new_n306_, new_n291_, new_n261_, new_n309_, new_n529_, new_n323_, new_n259_, new_n362_, new_n227_, new_n416_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n310_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n562_, new_n578_, new_n493_, new_n547_, new_n264_, new_n379_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n520_, new_n253_, new_n403_, new_n237_, new_n557_, new_n260_, new_n251_, new_n300_, new_n411_, new_n605_, new_n407_, new_n480_, new_n625_, new_n513_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n428_, new_n487_, new_n360_, new_n546_, new_n302_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n499_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n285_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n203_, new_n316_, new_n590_, new_n417_, new_n591_, new_n332_, new_n631_, new_n453_, new_n516_, new_n563_, new_n440_, new_n531_, new_n593_, new_n252_, new_n312_, new_n535_, new_n372_, new_n242_, new_n503_, new_n527_, new_n307_, new_n597_, new_n408_, new_n470_, new_n213_, new_n433_, new_n435_, new_n265_, new_n370_, new_n584_, new_n278_, new_n304_, new_n523_, new_n550_, new_n217_, new_n269_, new_n512_, new_n599_, new_n412_, new_n607_, new_n327_, new_n594_, new_n561_, new_n495_, new_n431_, new_n574_, new_n319_, new_n338_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n627_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n474_, new_n467_, new_n404_, new_n560_, new_n358_, new_n348_, new_n610_, new_n322_, new_n228_, new_n545_, new_n611_, new_n289_, new_n425_, new_n226_, new_n373_, new_n540_, new_n434_, new_n422_, new_n329_, new_n249_, new_n284_, new_n293_, new_n551_, new_n279_, new_n455_, new_n521_, new_n406_, new_n356_, new_n229_, new_n536_, new_n464_, new_n204_, new_n573_, new_n405_;

not g000 ( new_n202_, N1 );
xnor g001 ( new_n203_, N81, N85 );
xnor g002 ( new_n204_, new_n203_, keyIn_0_10 );
xnor g003 ( new_n205_, N89, N93 );
xnor g004 ( new_n206_, new_n205_, keyIn_0_11 );
xnor g005 ( new_n207_, new_n204_, new_n206_ );
xnor g006 ( new_n208_, new_n207_, keyIn_0_45 );
xor g007 ( new_n209_, N65, N69 );
xnor g008 ( new_n210_, new_n209_, keyIn_0_8 );
not g009 ( new_n211_, keyIn_0_9 );
xnor g010 ( new_n212_, N73, N77 );
and g011 ( new_n213_, new_n212_, new_n211_ );
or g012 ( new_n214_, N73, N77 );
and g013 ( new_n215_, N73, N77 );
not g014 ( new_n216_, new_n215_ );
and g015 ( new_n217_, new_n216_, keyIn_0_9, new_n214_ );
or g016 ( new_n218_, new_n213_, new_n217_ );
xnor g017 ( new_n219_, new_n218_, new_n210_ );
xnor g018 ( new_n220_, new_n219_, keyIn_0_44 );
xnor g019 ( new_n221_, new_n220_, new_n208_ );
xnor g020 ( new_n222_, new_n221_, keyIn_0_60 );
and g021 ( new_n223_, N129, N137 );
xnor g022 ( new_n224_, new_n223_, keyIn_0_16 );
xnor g023 ( new_n225_, new_n222_, new_n224_ );
xnor g024 ( new_n226_, new_n225_, keyIn_0_64 );
xor g025 ( new_n227_, N1, N17 );
xnor g026 ( new_n228_, new_n227_, keyIn_0_24 );
xnor g027 ( new_n229_, N33, N49 );
xnor g028 ( new_n230_, new_n229_, keyIn_0_25 );
xnor g029 ( new_n231_, new_n228_, new_n230_ );
xnor g030 ( new_n232_, new_n231_, keyIn_0_48 );
xnor g031 ( new_n233_, new_n226_, new_n232_ );
xor g032 ( new_n234_, new_n233_, keyIn_0_72 );
not g033 ( new_n235_, keyIn_0_76 );
xnor g034 ( new_n236_, N9, N13 );
xnor g035 ( new_n237_, new_n236_, keyIn_0_1 );
xnor g036 ( new_n238_, N1, N5 );
and g037 ( new_n239_, new_n238_, keyIn_0_0 );
not g038 ( new_n240_, keyIn_0_0 );
or g039 ( new_n241_, N1, N5 );
and g040 ( new_n242_, N1, N5 );
not g041 ( new_n243_, new_n242_ );
and g042 ( new_n244_, new_n243_, new_n240_, new_n241_ );
or g043 ( new_n245_, new_n239_, new_n244_ );
xnor g044 ( new_n246_, new_n245_, new_n237_ );
xnor g045 ( new_n247_, new_n246_, keyIn_0_40 );
xor g046 ( new_n248_, N17, N21 );
xnor g047 ( new_n249_, new_n248_, keyIn_0_2 );
xnor g048 ( new_n250_, N25, N29 );
xnor g049 ( new_n251_, new_n250_, keyIn_0_3 );
xnor g050 ( new_n252_, new_n249_, new_n251_ );
xnor g051 ( new_n253_, new_n252_, keyIn_0_41 );
xnor g052 ( new_n254_, new_n247_, new_n253_ );
xnor g053 ( new_n255_, new_n254_, keyIn_0_56 );
and g054 ( new_n256_, N133, N137 );
xnor g055 ( new_n257_, new_n256_, keyIn_0_20 );
xnor g056 ( new_n258_, new_n255_, new_n257_ );
xnor g057 ( new_n259_, new_n258_, keyIn_0_68 );
xor g058 ( new_n260_, N65, N81 );
xnor g059 ( new_n261_, new_n260_, keyIn_0_32 );
xnor g060 ( new_n262_, N97, N113 );
xnor g061 ( new_n263_, new_n262_, keyIn_0_33 );
xnor g062 ( new_n264_, new_n261_, new_n263_ );
xor g063 ( new_n265_, new_n264_, keyIn_0_52 );
xnor g064 ( new_n266_, new_n259_, new_n265_ );
xnor g065 ( new_n267_, new_n266_, new_n235_ );
not g066 ( new_n268_, new_n267_ );
not g067 ( new_n269_, keyIn_0_69 );
not g068 ( new_n270_, keyIn_0_42 );
xnor g069 ( new_n271_, N41, N45 );
xnor g070 ( new_n272_, new_n271_, keyIn_0_5 );
xnor g071 ( new_n273_, N33, N37 );
and g072 ( new_n274_, new_n273_, keyIn_0_4 );
not g073 ( new_n275_, keyIn_0_4 );
or g074 ( new_n276_, N33, N37 );
and g075 ( new_n277_, N33, N37 );
not g076 ( new_n278_, new_n277_ );
and g077 ( new_n279_, new_n278_, new_n275_, new_n276_ );
or g078 ( new_n280_, new_n274_, new_n279_ );
xnor g079 ( new_n281_, new_n280_, new_n272_ );
xnor g080 ( new_n282_, new_n281_, new_n270_ );
not g081 ( new_n283_, keyIn_0_43 );
xnor g082 ( new_n284_, N57, N61 );
xnor g083 ( new_n285_, new_n284_, keyIn_0_7 );
xnor g084 ( new_n286_, N49, N53 );
and g085 ( new_n287_, new_n286_, keyIn_0_6 );
not g086 ( new_n288_, keyIn_0_6 );
and g087 ( new_n289_, N49, N53 );
not g088 ( new_n290_, new_n289_ );
or g089 ( new_n291_, N49, N53 );
and g090 ( new_n292_, new_n290_, new_n288_, new_n291_ );
or g091 ( new_n293_, new_n287_, new_n292_ );
xnor g092 ( new_n294_, new_n293_, new_n285_ );
xnor g093 ( new_n295_, new_n294_, new_n283_ );
xnor g094 ( new_n296_, new_n282_, new_n295_ );
xnor g095 ( new_n297_, new_n296_, keyIn_0_57 );
and g096 ( new_n298_, N134, N137 );
xnor g097 ( new_n299_, new_n298_, keyIn_0_21 );
xnor g098 ( new_n300_, new_n297_, new_n299_ );
xnor g099 ( new_n301_, new_n300_, new_n269_ );
xor g100 ( new_n302_, N101, N117 );
xnor g101 ( new_n303_, new_n302_, keyIn_0_35 );
xnor g102 ( new_n304_, N69, N85 );
xnor g103 ( new_n305_, new_n304_, keyIn_0_34 );
xnor g104 ( new_n306_, new_n303_, new_n305_ );
xor g105 ( new_n307_, new_n306_, keyIn_0_53 );
xnor g106 ( new_n308_, new_n301_, new_n307_ );
xnor g107 ( new_n309_, new_n308_, keyIn_0_77 );
not g108 ( new_n310_, new_n309_ );
and g109 ( new_n311_, new_n310_, new_n268_ );
not g110 ( new_n312_, keyIn_0_112 );
not g111 ( new_n313_, keyIn_0_82 );
not g112 ( new_n314_, keyIn_0_74 );
not g113 ( new_n315_, keyIn_0_46 );
xnor g114 ( new_n316_, N97, N101 );
and g115 ( new_n317_, new_n316_, keyIn_0_12 );
not g116 ( new_n318_, keyIn_0_12 );
or g117 ( new_n319_, N97, N101 );
and g118 ( new_n320_, N97, N101 );
not g119 ( new_n321_, new_n320_ );
and g120 ( new_n322_, new_n321_, new_n318_, new_n319_ );
or g121 ( new_n323_, new_n317_, new_n322_ );
xnor g122 ( new_n324_, N105, N109 );
and g123 ( new_n325_, new_n324_, keyIn_0_13 );
not g124 ( new_n326_, keyIn_0_13 );
or g125 ( new_n327_, N105, N109 );
and g126 ( new_n328_, N105, N109 );
not g127 ( new_n329_, new_n328_ );
and g128 ( new_n330_, new_n329_, new_n326_, new_n327_ );
or g129 ( new_n331_, new_n325_, new_n330_ );
xnor g130 ( new_n332_, new_n323_, new_n331_ );
xnor g131 ( new_n333_, new_n332_, new_n315_ );
xnor g132 ( new_n334_, new_n333_, new_n220_ );
xnor g133 ( new_n335_, new_n334_, keyIn_0_62 );
and g134 ( new_n336_, N131, N137 );
xor g135 ( new_n337_, new_n336_, keyIn_0_18 );
xnor g136 ( new_n338_, new_n335_, new_n337_ );
xnor g137 ( new_n339_, new_n338_, keyIn_0_66 );
xor g138 ( new_n340_, N9, N25 );
xnor g139 ( new_n341_, new_n340_, keyIn_0_28 );
xnor g140 ( new_n342_, N41, N57 );
xnor g141 ( new_n343_, new_n342_, keyIn_0_29 );
xnor g142 ( new_n344_, new_n341_, new_n343_ );
xor g143 ( new_n345_, new_n344_, keyIn_0_50 );
xnor g144 ( new_n346_, new_n339_, new_n345_ );
xnor g145 ( new_n347_, new_n346_, new_n314_ );
or g146 ( new_n348_, new_n347_, new_n313_ );
xnor g147 ( new_n349_, N113, N117 );
and g148 ( new_n350_, new_n349_, keyIn_0_14 );
not g149 ( new_n351_, keyIn_0_14 );
or g150 ( new_n352_, N113, N117 );
and g151 ( new_n353_, N113, N117 );
not g152 ( new_n354_, new_n353_ );
and g153 ( new_n355_, new_n354_, new_n351_, new_n352_ );
or g154 ( new_n356_, new_n350_, new_n355_ );
xnor g155 ( new_n357_, N121, N125 );
and g156 ( new_n358_, new_n357_, keyIn_0_15 );
not g157 ( new_n359_, keyIn_0_15 );
and g158 ( new_n360_, N121, N125 );
not g159 ( new_n361_, new_n360_ );
or g160 ( new_n362_, N121, N125 );
and g161 ( new_n363_, new_n361_, new_n359_, new_n362_ );
or g162 ( new_n364_, new_n358_, new_n363_ );
xnor g163 ( new_n365_, new_n356_, new_n364_ );
xnor g164 ( new_n366_, new_n365_, keyIn_0_47 );
xnor g165 ( new_n367_, new_n366_, new_n208_ );
xnor g166 ( new_n368_, new_n367_, keyIn_0_63 );
and g167 ( new_n369_, N132, N137 );
xor g168 ( new_n370_, new_n369_, keyIn_0_19 );
xnor g169 ( new_n371_, new_n368_, new_n370_ );
xnor g170 ( new_n372_, new_n371_, keyIn_0_67 );
xor g171 ( new_n373_, N13, N29 );
xnor g172 ( new_n374_, new_n373_, keyIn_0_30 );
xor g173 ( new_n375_, N45, N61 );
xnor g174 ( new_n376_, new_n375_, keyIn_0_31 );
xnor g175 ( new_n377_, new_n374_, new_n376_ );
xnor g176 ( new_n378_, new_n377_, keyIn_0_51 );
xnor g177 ( new_n379_, new_n372_, new_n378_ );
xnor g178 ( new_n380_, new_n379_, keyIn_0_75 );
xnor g179 ( new_n381_, new_n346_, keyIn_0_74 );
or g180 ( new_n382_, new_n381_, keyIn_0_82 );
and g181 ( new_n383_, new_n382_, new_n380_ );
not g182 ( new_n384_, keyIn_0_80 );
xnor g183 ( new_n385_, new_n234_, new_n384_ );
not g184 ( new_n386_, keyIn_0_73 );
xnor g185 ( new_n387_, new_n333_, new_n366_ );
xnor g186 ( new_n388_, new_n387_, keyIn_0_61 );
and g187 ( new_n389_, N130, N137 );
xor g188 ( new_n390_, new_n389_, keyIn_0_17 );
xnor g189 ( new_n391_, new_n388_, new_n390_ );
xnor g190 ( new_n392_, new_n391_, keyIn_0_65 );
xor g191 ( new_n393_, N37, N53 );
xor g192 ( new_n394_, new_n393_, keyIn_0_27 );
xor g193 ( new_n395_, N5, N21 );
xnor g194 ( new_n396_, new_n395_, keyIn_0_26 );
xnor g195 ( new_n397_, new_n394_, new_n396_ );
xnor g196 ( new_n398_, new_n397_, keyIn_0_49 );
xnor g197 ( new_n399_, new_n392_, new_n398_ );
xnor g198 ( new_n400_, new_n399_, new_n386_ );
xnor g199 ( new_n401_, new_n400_, keyIn_0_81 );
and g200 ( new_n402_, new_n383_, new_n348_, new_n385_, new_n401_ );
xnor g201 ( new_n403_, new_n402_, keyIn_0_104 );
not g202 ( new_n404_, keyIn_0_107 );
not g203 ( new_n405_, keyIn_0_90 );
or g204 ( new_n406_, new_n347_, new_n405_ );
or g205 ( new_n407_, new_n381_, keyIn_0_90 );
and g206 ( new_n408_, new_n406_, new_n407_, new_n234_ );
and g207 ( new_n409_, new_n400_, keyIn_0_89 );
not g208 ( new_n410_, keyIn_0_89 );
or g209 ( new_n411_, new_n399_, new_n386_ );
xor g210 ( new_n412_, new_n397_, keyIn_0_49 );
xnor g211 ( new_n413_, new_n392_, new_n412_ );
or g212 ( new_n414_, new_n413_, keyIn_0_73 );
and g213 ( new_n415_, new_n411_, new_n414_, new_n410_ );
or g214 ( new_n416_, new_n409_, new_n415_ );
xor g215 ( new_n417_, new_n380_, keyIn_0_91 );
and g216 ( new_n418_, new_n408_, new_n416_, new_n417_ );
xnor g217 ( new_n419_, new_n418_, new_n404_ );
or g218 ( new_n420_, new_n400_, keyIn_0_84 );
not g219 ( new_n421_, keyIn_0_84 );
xnor g220 ( new_n422_, new_n399_, keyIn_0_73 );
or g221 ( new_n423_, new_n422_, new_n421_ );
and g222 ( new_n424_, new_n423_, new_n347_ );
xnor g223 ( new_n425_, new_n234_, keyIn_0_83 );
xor g224 ( new_n426_, new_n380_, keyIn_0_85 );
and g225 ( new_n427_, new_n424_, new_n420_, new_n425_, new_n426_ );
xnor g226 ( new_n428_, new_n427_, keyIn_0_105 );
not g227 ( new_n429_, keyIn_0_106 );
not g228 ( new_n430_, keyIn_0_87 );
or g229 ( new_n431_, new_n347_, new_n430_ );
xnor g230 ( new_n432_, new_n380_, keyIn_0_88 );
or g231 ( new_n433_, new_n381_, keyIn_0_87 );
and g232 ( new_n434_, new_n433_, new_n422_ );
not g233 ( new_n435_, keyIn_0_86 );
xnor g234 ( new_n436_, new_n234_, new_n435_ );
and g235 ( new_n437_, new_n434_, new_n431_, new_n432_, new_n436_ );
xnor g236 ( new_n438_, new_n437_, new_n429_ );
and g237 ( new_n439_, new_n428_, new_n419_, new_n403_, new_n438_ );
xnor g238 ( new_n440_, new_n439_, new_n312_ );
not g239 ( new_n441_, keyIn_0_79 );
xnor g240 ( new_n442_, new_n295_, new_n253_ );
xnor g241 ( new_n443_, new_n442_, keyIn_0_59 );
and g242 ( new_n444_, N136, N137 );
xnor g243 ( new_n445_, new_n444_, keyIn_0_23 );
xnor g244 ( new_n446_, new_n443_, new_n445_ );
xnor g245 ( new_n447_, new_n446_, keyIn_0_71 );
xor g246 ( new_n448_, N77, N93 );
xnor g247 ( new_n449_, new_n448_, keyIn_0_38 );
xnor g248 ( new_n450_, N109, N125 );
xnor g249 ( new_n451_, new_n450_, keyIn_0_39 );
xnor g250 ( new_n452_, new_n449_, new_n451_ );
xor g251 ( new_n453_, new_n452_, keyIn_0_55 );
xnor g252 ( new_n454_, new_n447_, new_n453_ );
xnor g253 ( new_n455_, new_n454_, new_n441_ );
not g254 ( new_n456_, new_n455_ );
xnor g255 ( new_n457_, new_n247_, new_n282_ );
xnor g256 ( new_n458_, new_n457_, keyIn_0_58 );
and g257 ( new_n459_, N135, N137 );
xnor g258 ( new_n460_, new_n459_, keyIn_0_22 );
xnor g259 ( new_n461_, new_n458_, new_n460_ );
xnor g260 ( new_n462_, new_n461_, keyIn_0_70 );
xor g261 ( new_n463_, N105, N121 );
xor g262 ( new_n464_, new_n463_, keyIn_0_37 );
xor g263 ( new_n465_, N73, N89 );
xnor g264 ( new_n466_, new_n465_, keyIn_0_36 );
xnor g265 ( new_n467_, new_n464_, new_n466_ );
xnor g266 ( new_n468_, new_n467_, keyIn_0_54 );
xnor g267 ( new_n469_, new_n462_, new_n468_ );
xnor g268 ( new_n470_, new_n469_, keyIn_0_78 );
and g269 ( new_n471_, new_n440_, new_n456_, new_n470_ );
and g270 ( new_n472_, new_n471_, new_n311_ );
xor g271 ( new_n473_, new_n472_, keyIn_0_114 );
and g272 ( new_n474_, new_n473_, new_n234_ );
xnor g273 ( N724, new_n474_, new_n202_ );
not g274 ( new_n476_, N5 );
and g275 ( new_n477_, new_n473_, new_n422_ );
xnor g276 ( N725, new_n477_, new_n476_ );
not g277 ( new_n479_, N9 );
and g278 ( new_n480_, new_n473_, new_n347_ );
xnor g279 ( N726, new_n480_, new_n479_ );
not g280 ( new_n482_, N13 );
and g281 ( new_n483_, new_n473_, new_n380_ );
xnor g282 ( N727, new_n483_, new_n482_ );
not g283 ( new_n485_, keyIn_0_78 );
xnor g284 ( new_n486_, new_n469_, new_n485_ );
and g285 ( new_n487_, new_n440_, new_n311_, new_n455_, new_n486_ );
xnor g286 ( new_n488_, new_n487_, keyIn_0_115 );
and g287 ( new_n489_, new_n488_, new_n234_ );
xor g288 ( N728, new_n489_, N17 );
and g289 ( new_n491_, new_n488_, new_n422_ );
xor g290 ( N729, new_n491_, N21 );
and g291 ( new_n493_, new_n488_, new_n347_ );
xor g292 ( N730, new_n493_, N25 );
and g293 ( new_n495_, new_n488_, new_n380_ );
xor g294 ( N731, new_n495_, N29 );
not g295 ( new_n497_, N33 );
and g296 ( new_n498_, new_n471_, new_n267_, new_n309_ );
xnor g297 ( new_n499_, new_n498_, keyIn_0_116 );
and g298 ( new_n500_, new_n499_, new_n234_ );
xnor g299 ( N732, new_n500_, new_n497_ );
not g300 ( new_n502_, N37 );
and g301 ( new_n503_, new_n499_, new_n422_ );
xnor g302 ( N733, new_n503_, new_n502_ );
not g303 ( new_n505_, N41 );
and g304 ( new_n506_, new_n499_, new_n347_ );
xnor g305 ( N734, new_n506_, new_n505_ );
not g306 ( new_n508_, N45 );
and g307 ( new_n509_, new_n499_, new_n380_ );
xnor g308 ( N735, new_n509_, new_n508_ );
and g309 ( new_n511_, new_n309_, new_n486_, new_n267_, new_n455_ );
and g310 ( new_n512_, new_n440_, new_n511_ );
xnor g311 ( new_n513_, new_n512_, keyIn_0_117 );
and g312 ( new_n514_, new_n513_, new_n234_ );
xor g313 ( N736, new_n514_, N49 );
and g314 ( new_n516_, new_n513_, new_n422_ );
xor g315 ( N737, new_n516_, N53 );
and g316 ( new_n518_, new_n513_, new_n347_ );
xor g317 ( N738, new_n518_, N57 );
and g318 ( new_n520_, new_n513_, new_n380_ );
xnor g319 ( new_n521_, new_n520_, keyIn_0_122 );
xnor g320 ( N739, new_n521_, N61 );
not g321 ( new_n523_, N65 );
not g322 ( new_n524_, keyIn_0_118 );
not g323 ( new_n525_, new_n380_ );
and g324 ( new_n526_, new_n525_, new_n347_ );
not g325 ( new_n527_, keyIn_0_113 );
not g326 ( new_n528_, keyIn_0_110 );
not g327 ( new_n529_, keyIn_0_100 );
or g328 ( new_n530_, new_n456_, new_n529_ );
or g329 ( new_n531_, new_n455_, keyIn_0_100 );
and g330 ( new_n532_, new_n531_, new_n309_ );
xnor g331 ( new_n533_, new_n267_, keyIn_0_98 );
xnor g332 ( new_n534_, new_n470_, keyIn_0_99 );
and g333 ( new_n535_, new_n532_, new_n530_, new_n533_, new_n534_ );
xnor g334 ( new_n536_, new_n535_, new_n528_ );
not g335 ( new_n537_, keyIn_0_108 );
not g336 ( new_n538_, keyIn_0_92 );
or g337 ( new_n539_, new_n268_, new_n538_ );
or g338 ( new_n540_, new_n267_, keyIn_0_92 );
and g339 ( new_n541_, new_n540_, new_n455_ );
xnor g340 ( new_n542_, new_n486_, keyIn_0_94 );
xnor g341 ( new_n543_, new_n309_, keyIn_0_93 );
and g342 ( new_n544_, new_n541_, new_n539_, new_n542_, new_n543_ );
xnor g343 ( new_n545_, new_n544_, new_n537_ );
not g344 ( new_n546_, keyIn_0_109 );
not g345 ( new_n547_, keyIn_0_97 );
or g346 ( new_n548_, new_n456_, new_n547_ );
or g347 ( new_n549_, new_n455_, keyIn_0_97 );
and g348 ( new_n550_, new_n549_, new_n470_ );
xnor g349 ( new_n551_, new_n267_, keyIn_0_95 );
not g350 ( new_n552_, keyIn_0_96 );
xnor g351 ( new_n553_, new_n309_, new_n552_ );
and g352 ( new_n554_, new_n550_, new_n548_, new_n551_, new_n553_ );
xnor g353 ( new_n555_, new_n554_, new_n546_ );
not g354 ( new_n556_, keyIn_0_103 );
or g355 ( new_n557_, new_n456_, new_n556_ );
or g356 ( new_n558_, new_n309_, keyIn_0_101 );
or g357 ( new_n559_, new_n455_, keyIn_0_103 );
and g358 ( new_n560_, new_n558_, new_n559_ );
xnor g359 ( new_n561_, new_n470_, keyIn_0_102 );
not g360 ( new_n562_, keyIn_0_101 );
not g361 ( new_n563_, keyIn_0_77 );
and g362 ( new_n564_, new_n308_, new_n563_ );
xnor g363 ( new_n565_, new_n300_, keyIn_0_69 );
not g364 ( new_n566_, new_n307_ );
or g365 ( new_n567_, new_n565_, new_n566_ );
or g366 ( new_n568_, new_n301_, new_n307_ );
and g367 ( new_n569_, new_n567_, new_n568_, keyIn_0_77 );
or g368 ( new_n570_, new_n564_, new_n562_, new_n569_ );
and g369 ( new_n571_, new_n570_, new_n268_ );
and g370 ( new_n572_, new_n560_, new_n557_, new_n561_, new_n571_ );
xnor g371 ( new_n573_, new_n572_, keyIn_0_111 );
and g372 ( new_n574_, new_n573_, new_n536_, new_n545_, new_n555_ );
xnor g373 ( new_n575_, new_n574_, new_n527_ );
and g374 ( new_n576_, new_n234_, new_n400_ );
and g375 ( new_n577_, new_n575_, new_n526_, new_n576_ );
xnor g376 ( new_n578_, new_n577_, new_n524_ );
and g377 ( new_n579_, new_n578_, new_n268_ );
xnor g378 ( new_n580_, new_n579_, keyIn_0_123 );
xnor g379 ( N740, new_n580_, new_n523_ );
not g380 ( new_n582_, keyIn_0_124 );
and g381 ( new_n583_, new_n578_, new_n309_ );
xnor g382 ( new_n584_, new_n583_, new_n582_ );
xnor g383 ( N741, new_n584_, N69 );
and g384 ( new_n586_, new_n578_, new_n470_ );
xnor g385 ( new_n587_, new_n586_, keyIn_0_125 );
xnor g386 ( N742, new_n587_, N73 );
not g387 ( new_n589_, keyIn_0_126 );
and g388 ( new_n590_, new_n578_, new_n455_ );
xnor g389 ( new_n591_, new_n590_, new_n589_ );
xnor g390 ( N743, new_n591_, N77 );
not g391 ( new_n593_, N81 );
not g392 ( new_n594_, keyIn_0_119 );
and g393 ( new_n595_, new_n381_, new_n380_ );
and g394 ( new_n596_, new_n575_, new_n576_, new_n595_ );
xnor g395 ( new_n597_, new_n596_, new_n594_ );
and g396 ( new_n598_, new_n597_, new_n268_ );
xnor g397 ( new_n599_, new_n598_, keyIn_0_127 );
xnor g398 ( N744, new_n599_, new_n593_ );
and g399 ( new_n601_, new_n597_, new_n309_ );
xor g400 ( N745, new_n601_, N85 );
and g401 ( new_n603_, new_n597_, new_n470_ );
xor g402 ( N746, new_n603_, N89 );
and g403 ( new_n605_, new_n597_, new_n455_ );
xor g404 ( N747, new_n605_, N93 );
not g405 ( new_n607_, new_n234_ );
and g406 ( new_n608_, new_n575_, new_n607_, new_n422_ );
and g407 ( new_n609_, new_n608_, new_n526_ );
xnor g408 ( new_n610_, new_n609_, keyIn_0_120 );
and g409 ( new_n611_, new_n610_, new_n268_ );
xor g410 ( N748, new_n611_, N97 );
and g411 ( new_n613_, new_n610_, new_n309_ );
xor g412 ( N749, new_n613_, N101 );
and g413 ( new_n615_, new_n610_, new_n470_ );
xor g414 ( N750, new_n615_, N105 );
and g415 ( new_n617_, new_n610_, new_n455_ );
xor g416 ( N751, new_n617_, N109 );
not g417 ( new_n619_, N113 );
and g418 ( new_n620_, new_n608_, new_n595_ );
xor g419 ( new_n621_, new_n620_, keyIn_0_121 );
and g420 ( new_n622_, new_n621_, new_n268_ );
xnor g421 ( N752, new_n622_, new_n619_ );
not g422 ( new_n624_, N117 );
and g423 ( new_n625_, new_n621_, new_n309_ );
xnor g424 ( N753, new_n625_, new_n624_ );
not g425 ( new_n627_, N121 );
and g426 ( new_n628_, new_n621_, new_n470_ );
xnor g427 ( N754, new_n628_, new_n627_ );
not g428 ( new_n630_, N125 );
and g429 ( new_n631_, new_n621_, new_n455_ );
xnor g430 ( N755, new_n631_, new_n630_ );
endmodule