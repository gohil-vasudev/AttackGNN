module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n614_, new_n445_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n288_, new_n421_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n636_, new_n670_, new_n456_, new_n691_, new_n170_, new_n246_, new_n682_, new_n266_, new_n667_, new_n367_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n637_, new_n214_, new_n451_, new_n424_, new_n602_, new_n114_, new_n188_, new_n240_, new_n660_, new_n413_, new_n695_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n649_, new_n678_, new_n462_, new_n603_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n427_, new_n234_, new_n532_, new_n393_, new_n418_, new_n292_, new_n215_, new_n626_, new_n152_, new_n157_, new_n153_, new_n133_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n110_, new_n315_, new_n685_, new_n124_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n117_, new_n630_, new_n167_, new_n385_, new_n478_, new_n694_, new_n461_, new_n297_, new_n361_, new_n565_, new_n150_, new_n683_, new_n108_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n622_, new_n629_, new_n321_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n650_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n506_, new_n680_, new_n256_, new_n452_, new_n381_, new_n656_, new_n388_, new_n508_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n657_, new_n652_, new_n314_, new_n582_, new_n118_, new_n363_, new_n165_, new_n441_, new_n477_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n187_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n346_, new_n396_, new_n198_, new_n438_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n399_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n628_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n688_, new_n155_, new_n384_, new_n410_, new_n543_, new_n113_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n309_, new_n529_, new_n323_, new_n259_, new_n362_, new_n654_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n693_, new_n130_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n138_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n562_, new_n578_, new_n126_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n379_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n143_, new_n520_, new_n125_, new_n145_, new_n253_, new_n403_, new_n475_, new_n237_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n106_, new_n411_, new_n507_, new_n673_, new_n605_, new_n107_, new_n182_, new_n407_, new_n666_, new_n625_, new_n151_, new_n592_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n522_, new_n588_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n302_, new_n191_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n112_, new_n121_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n174_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n147_, new_n285_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n515_, new_n332_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n662_, new_n440_, new_n122_, new_n531_, new_n593_, new_n111_, new_n252_, new_n585_, new_n160_, new_n312_, new_n535_, new_n372_, new_n242_, new_n503_, new_n527_, new_n115_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n134_, new_n651_, new_n433_, new_n435_, new_n109_, new_n265_, new_n370_, new_n689_, new_n584_, new_n278_, new_n304_, new_n523_, new_n638_, new_n550_, new_n217_, new_n269_, new_n512_, new_n129_, new_n644_, new_n599_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n594_, new_n561_, new_n495_, new_n431_, new_n196_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n627_, new_n195_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n128_, new_n358_, new_n348_, new_n610_, new_n159_, new_n322_, new_n228_, new_n545_, new_n611_, new_n289_, new_n425_, new_n175_, new_n226_, new_n185_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n618_, new_n120_, new_n406_, new_n356_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n135_, new_n573_, new_n405_;

not g000 ( new_n106_, N85 );
nand g001 ( new_n107_, new_n106_, N81 );
not g002 ( new_n108_, N81 );
nand g003 ( new_n109_, new_n108_, N85 );
nand g004 ( new_n110_, new_n107_, new_n109_ );
not g005 ( new_n111_, N89 );
not g006 ( new_n112_, N93 );
nand g007 ( new_n113_, new_n111_, new_n112_ );
nand g008 ( new_n114_, N89, N93 );
nand g009 ( new_n115_, new_n113_, new_n114_ );
nand g010 ( new_n116_, new_n110_, new_n115_ );
nand g011 ( new_n117_, new_n113_, new_n107_, new_n109_, new_n114_ );
nand g012 ( new_n118_, new_n116_, new_n117_ );
not g013 ( new_n119_, new_n118_ );
not g014 ( new_n120_, N69 );
nand g015 ( new_n121_, new_n120_, N65 );
not g016 ( new_n122_, N65 );
nand g017 ( new_n123_, new_n122_, N69 );
nand g018 ( new_n124_, new_n121_, new_n123_ );
not g019 ( new_n125_, N73 );
not g020 ( new_n126_, N77 );
nand g021 ( new_n127_, new_n125_, new_n126_ );
nand g022 ( new_n128_, N73, N77 );
nand g023 ( new_n129_, new_n127_, new_n128_ );
nand g024 ( new_n130_, new_n124_, new_n129_ );
nand g025 ( new_n131_, new_n127_, new_n121_, new_n123_, new_n128_ );
nand g026 ( new_n132_, new_n130_, new_n131_ );
not g027 ( new_n133_, new_n132_ );
nand g028 ( new_n134_, new_n119_, new_n133_ );
nand g029 ( new_n135_, new_n118_, new_n132_ );
nand g030 ( new_n136_, N129, N137 );
nand g031 ( new_n137_, new_n134_, new_n135_, new_n136_ );
nand g032 ( new_n138_, new_n134_, new_n135_ );
nand g033 ( new_n139_, new_n138_, N129, N137 );
nand g034 ( new_n140_, new_n139_, new_n137_ );
not g035 ( new_n141_, N17 );
nand g036 ( new_n142_, new_n141_, N1 );
not g037 ( new_n143_, N1 );
nand g038 ( new_n144_, new_n143_, N17 );
nand g039 ( new_n145_, new_n142_, new_n144_ );
not g040 ( new_n146_, N33 );
not g041 ( new_n147_, N49 );
nand g042 ( new_n148_, new_n146_, new_n147_ );
nand g043 ( new_n149_, N33, N49 );
nand g044 ( new_n150_, new_n148_, new_n149_ );
nand g045 ( new_n151_, new_n145_, new_n150_ );
nand g046 ( new_n152_, new_n148_, new_n142_, new_n144_, new_n149_ );
nand g047 ( new_n153_, new_n151_, new_n152_ );
nand g048 ( new_n154_, new_n153_, keyIn_0_9 );
not g049 ( new_n155_, keyIn_0_9 );
nand g050 ( new_n156_, new_n151_, new_n155_, new_n152_ );
nand g051 ( new_n157_, new_n154_, new_n156_ );
nand g052 ( new_n158_, new_n140_, new_n157_ );
nand g053 ( new_n159_, new_n139_, new_n137_, new_n154_, new_n156_ );
nand g054 ( new_n160_, new_n158_, new_n159_ );
not g055 ( new_n161_, new_n160_ );
not g056 ( new_n162_, keyIn_0_24 );
nor g057 ( new_n163_, N113, N117 );
not g058 ( new_n164_, new_n163_ );
nand g059 ( new_n165_, N113, N117 );
nor g060 ( new_n166_, N121, N125 );
not g061 ( new_n167_, new_n166_ );
nand g062 ( new_n168_, N121, N125 );
nand g063 ( new_n169_, new_n167_, new_n168_ );
nand g064 ( new_n170_, new_n169_, keyIn_0_4 );
not g065 ( new_n171_, keyIn_0_4 );
nand g066 ( new_n172_, new_n167_, new_n171_, new_n168_ );
nand g067 ( new_n173_, new_n170_, new_n164_, new_n165_, new_n172_ );
nand g068 ( new_n174_, new_n164_, new_n165_ );
nand g069 ( new_n175_, new_n170_, new_n172_ );
nand g070 ( new_n176_, new_n175_, new_n174_ );
nand g071 ( new_n177_, new_n176_, new_n173_ );
not g072 ( new_n178_, new_n177_ );
nand g073 ( new_n179_, new_n178_, new_n119_ );
nand g074 ( new_n180_, new_n177_, new_n118_ );
nand g075 ( new_n181_, N132, N137 );
nand g076 ( new_n182_, new_n179_, new_n180_, new_n181_ );
nand g077 ( new_n183_, new_n179_, new_n180_ );
nand g078 ( new_n184_, new_n183_, N132, N137 );
not g079 ( new_n185_, N13 );
not g080 ( new_n186_, N29 );
nand g081 ( new_n187_, new_n185_, new_n186_ );
nand g082 ( new_n188_, N13, N29 );
nand g083 ( new_n189_, new_n187_, new_n188_ );
not g084 ( new_n190_, N45 );
not g085 ( new_n191_, N61 );
nand g086 ( new_n192_, new_n190_, new_n191_ );
nand g087 ( new_n193_, N45, N61 );
nand g088 ( new_n194_, new_n192_, new_n193_ );
nand g089 ( new_n195_, new_n189_, new_n194_ );
nand g090 ( new_n196_, new_n187_, new_n192_, new_n188_, new_n193_ );
nand g091 ( new_n197_, new_n195_, new_n196_ );
nand g092 ( new_n198_, new_n184_, new_n182_, new_n197_ );
nand g093 ( new_n199_, new_n184_, new_n182_ );
nand g094 ( new_n200_, new_n199_, new_n195_, new_n196_ );
nand g095 ( new_n201_, new_n200_, new_n198_ );
nand g096 ( new_n202_, N105, N109 );
nor g097 ( new_n203_, N105, N109 );
not g098 ( new_n204_, new_n203_ );
nand g099 ( new_n205_, new_n204_, new_n202_ );
nand g100 ( new_n206_, new_n205_, keyIn_0_3 );
not g101 ( new_n207_, keyIn_0_3 );
nand g102 ( new_n208_, new_n204_, new_n207_, new_n202_ );
nand g103 ( new_n209_, new_n206_, new_n208_ );
not g104 ( new_n210_, N97 );
not g105 ( new_n211_, N101 );
nand g106 ( new_n212_, new_n210_, new_n211_ );
nand g107 ( new_n213_, N97, N101 );
nand g108 ( new_n214_, new_n212_, new_n213_ );
nand g109 ( new_n215_, new_n209_, new_n214_ );
nand g110 ( new_n216_, new_n206_, new_n208_, new_n212_, new_n213_ );
nand g111 ( new_n217_, new_n215_, new_n216_ );
not g112 ( new_n218_, new_n217_ );
nand g113 ( new_n219_, new_n218_, new_n133_ );
nand g114 ( new_n220_, new_n217_, new_n132_ );
nand g115 ( new_n221_, N131, N137 );
nand g116 ( new_n222_, new_n219_, new_n220_, new_n221_ );
nand g117 ( new_n223_, new_n219_, new_n220_ );
nand g118 ( new_n224_, new_n223_, N131, N137 );
nand g119 ( new_n225_, new_n224_, new_n222_ );
nor g120 ( new_n226_, N41, N57 );
not g121 ( new_n227_, new_n226_ );
nand g122 ( new_n228_, N41, N57 );
nand g123 ( new_n229_, new_n227_, new_n228_ );
nand g124 ( new_n230_, new_n229_, keyIn_0_6 );
not g125 ( new_n231_, new_n230_ );
nor g126 ( new_n232_, new_n229_, keyIn_0_6 );
nor g127 ( new_n233_, new_n231_, new_n232_ );
not g128 ( new_n234_, new_n233_ );
not g129 ( new_n235_, N9 );
nor g130 ( new_n236_, new_n235_, N25 );
not g131 ( new_n237_, N25 );
nor g132 ( new_n238_, new_n237_, N9 );
nor g133 ( new_n239_, new_n236_, new_n238_ );
not g134 ( new_n240_, new_n239_ );
nand g135 ( new_n241_, new_n234_, new_n240_ );
nand g136 ( new_n242_, new_n233_, new_n239_ );
nand g137 ( new_n243_, new_n241_, new_n242_ );
nand g138 ( new_n244_, new_n225_, new_n243_ );
nand g139 ( new_n245_, new_n224_, new_n222_, new_n241_, new_n242_ );
nand g140 ( new_n246_, new_n244_, new_n245_, new_n161_ );
not g141 ( new_n247_, new_n246_ );
not g142 ( new_n248_, keyIn_0_13 );
nand g143 ( new_n249_, new_n178_, new_n218_ );
nand g144 ( new_n250_, new_n177_, new_n217_ );
nand g145 ( new_n251_, new_n249_, new_n250_ );
nand g146 ( new_n252_, N130, N137 );
nand g147 ( new_n253_, new_n251_, new_n252_ );
nand g148 ( new_n254_, new_n249_, N130, N137, new_n250_ );
nand g149 ( new_n255_, new_n253_, new_n254_ );
not g150 ( new_n256_, N5 );
not g151 ( new_n257_, N21 );
nand g152 ( new_n258_, new_n256_, new_n257_ );
nand g153 ( new_n259_, N5, N21 );
nand g154 ( new_n260_, new_n258_, new_n259_ );
not g155 ( new_n261_, N37 );
not g156 ( new_n262_, N53 );
nand g157 ( new_n263_, new_n261_, new_n262_ );
nand g158 ( new_n264_, N37, N53 );
nand g159 ( new_n265_, new_n263_, new_n264_ );
nand g160 ( new_n266_, new_n260_, new_n265_ );
nand g161 ( new_n267_, new_n258_, new_n263_, new_n259_, new_n264_ );
nand g162 ( new_n268_, new_n266_, new_n267_ );
nand g163 ( new_n269_, new_n255_, new_n268_ );
nand g164 ( new_n270_, new_n253_, new_n254_, new_n266_, new_n267_ );
nand g165 ( new_n271_, new_n269_, new_n270_ );
nand g166 ( new_n272_, new_n271_, new_n248_ );
not g167 ( new_n273_, new_n271_ );
nand g168 ( new_n274_, new_n273_, keyIn_0_13 );
nand g169 ( new_n275_, new_n274_, new_n201_, new_n247_, new_n272_ );
not g170 ( new_n276_, keyIn_0_19 );
nand g171 ( new_n277_, new_n244_, new_n245_ );
nor g172 ( new_n278_, new_n201_, new_n277_, new_n271_ );
nand g173 ( new_n279_, new_n161_, keyIn_0_11 );
not g174 ( new_n280_, keyIn_0_11 );
nand g175 ( new_n281_, new_n160_, new_n280_ );
nand g176 ( new_n282_, new_n279_, new_n281_ );
not g177 ( new_n283_, new_n282_ );
nand g178 ( new_n284_, new_n278_, new_n283_ );
nand g179 ( new_n285_, new_n284_, new_n276_ );
nand g180 ( new_n286_, new_n277_, new_n271_, keyIn_0_12 );
nand g181 ( new_n287_, new_n277_, keyIn_0_12 );
nand g182 ( new_n288_, new_n287_, new_n273_ );
nand g183 ( new_n289_, new_n288_, new_n201_, new_n160_, new_n286_ );
nand g184 ( new_n290_, new_n278_, keyIn_0_19, new_n283_ );
nand g185 ( new_n291_, new_n285_, new_n275_, new_n289_, new_n290_ );
not g186 ( new_n292_, keyIn_0_10 );
nand g187 ( new_n293_, new_n147_, new_n262_ );
nand g188 ( new_n294_, N49, N53 );
nand g189 ( new_n295_, new_n293_, new_n294_ );
not g190 ( new_n296_, N57 );
nand g191 ( new_n297_, new_n296_, new_n191_ );
nand g192 ( new_n298_, N57, N61 );
nand g193 ( new_n299_, new_n297_, new_n298_ );
nand g194 ( new_n300_, new_n295_, new_n299_ );
nand g195 ( new_n301_, new_n293_, new_n297_, new_n294_, new_n298_ );
nand g196 ( new_n302_, new_n300_, new_n301_ );
not g197 ( new_n303_, keyIn_0_0 );
nand g198 ( new_n304_, new_n141_, new_n257_ );
nand g199 ( new_n305_, N17, N21 );
nand g200 ( new_n306_, new_n304_, new_n305_ );
nand g201 ( new_n307_, new_n306_, new_n303_ );
nand g202 ( new_n308_, new_n304_, keyIn_0_0, new_n305_ );
nand g203 ( new_n309_, N25, N29 );
not g204 ( new_n310_, new_n309_ );
nor g205 ( new_n311_, N25, N29 );
nor g206 ( new_n312_, new_n310_, new_n311_ );
not g207 ( new_n313_, new_n312_ );
nand g208 ( new_n314_, new_n307_, new_n313_, new_n308_ );
nand g209 ( new_n315_, new_n307_, new_n308_ );
nand g210 ( new_n316_, new_n315_, new_n312_ );
nand g211 ( new_n317_, new_n316_, new_n314_ );
nand g212 ( new_n318_, new_n317_, new_n302_ );
not g213 ( new_n319_, new_n302_ );
nand g214 ( new_n320_, new_n316_, new_n319_, new_n314_ );
nand g215 ( new_n321_, N136, N137 );
nand g216 ( new_n322_, new_n318_, new_n320_, new_n321_ );
nand g217 ( new_n323_, new_n318_, new_n320_ );
not g218 ( new_n324_, new_n321_ );
nand g219 ( new_n325_, new_n323_, new_n324_ );
nand g220 ( new_n326_, new_n325_, new_n322_ );
nand g221 ( new_n327_, new_n326_, new_n292_ );
nand g222 ( new_n328_, new_n325_, keyIn_0_10, new_n322_ );
nand g223 ( new_n329_, new_n327_, new_n328_ );
nand g224 ( new_n330_, new_n126_, new_n112_ );
nand g225 ( new_n331_, N77, N93 );
nand g226 ( new_n332_, new_n330_, new_n331_ );
not g227 ( new_n333_, N109 );
not g228 ( new_n334_, N125 );
nand g229 ( new_n335_, new_n333_, new_n334_ );
nand g230 ( new_n336_, N109, N125 );
nand g231 ( new_n337_, new_n335_, new_n336_ );
nand g232 ( new_n338_, new_n332_, new_n337_ );
nand g233 ( new_n339_, new_n330_, new_n335_, new_n331_, new_n336_ );
nand g234 ( new_n340_, new_n338_, new_n339_ );
nand g235 ( new_n341_, new_n329_, new_n340_ );
nand g236 ( new_n342_, new_n327_, new_n328_, new_n338_, new_n339_ );
nand g237 ( new_n343_, new_n341_, new_n342_ );
not g238 ( new_n344_, new_n343_ );
nand g239 ( new_n345_, new_n344_, keyIn_0_15 );
not g240 ( new_n346_, keyIn_0_15 );
nand g241 ( new_n347_, new_n343_, new_n346_ );
nand g242 ( new_n348_, new_n345_, new_n347_ );
not g243 ( new_n349_, keyIn_0_14 );
nand g244 ( new_n350_, N33, N37 );
nand g245 ( new_n351_, new_n146_, new_n261_ );
nand g246 ( new_n352_, new_n351_, new_n350_ );
not g247 ( new_n353_, N41 );
nand g248 ( new_n354_, new_n353_, new_n190_ );
nand g249 ( new_n355_, N41, N45 );
not g250 ( new_n356_, keyIn_0_2 );
nand g251 ( new_n357_, new_n356_, keyIn_0_1 );
not g252 ( new_n358_, keyIn_0_1 );
nand g253 ( new_n359_, new_n358_, keyIn_0_2 );
nand g254 ( new_n360_, new_n354_, new_n357_, new_n359_, new_n355_ );
nand g255 ( new_n361_, new_n354_, new_n355_ );
nand g256 ( new_n362_, new_n357_, new_n359_ );
nand g257 ( new_n363_, new_n361_, new_n362_ );
nand g258 ( new_n364_, new_n363_, new_n360_ );
nand g259 ( new_n365_, new_n364_, new_n352_ );
nand g260 ( new_n366_, new_n363_, new_n350_, new_n351_, new_n360_ );
nand g261 ( new_n367_, new_n365_, new_n366_ );
nand g262 ( new_n368_, new_n367_, keyIn_0_8 );
not g263 ( new_n369_, keyIn_0_8 );
nand g264 ( new_n370_, new_n365_, new_n369_, new_n366_ );
nand g265 ( new_n371_, new_n368_, new_n370_ );
nand g266 ( new_n372_, new_n371_, new_n319_ );
nand g267 ( new_n373_, new_n368_, new_n302_, new_n370_ );
nand g268 ( new_n374_, new_n372_, new_n373_ );
nand g269 ( new_n375_, N134, N137 );
not g270 ( new_n376_, new_n375_ );
nand g271 ( new_n377_, new_n374_, new_n376_ );
nand g272 ( new_n378_, new_n372_, new_n373_, new_n375_ );
nand g273 ( new_n379_, new_n377_, new_n378_ );
nand g274 ( new_n380_, new_n120_, new_n106_ );
nand g275 ( new_n381_, N69, N85 );
nand g276 ( new_n382_, new_n380_, new_n381_ );
not g277 ( new_n383_, N117 );
nand g278 ( new_n384_, new_n211_, new_n383_ );
nand g279 ( new_n385_, N101, N117 );
nand g280 ( new_n386_, new_n384_, new_n385_ );
nand g281 ( new_n387_, new_n382_, new_n386_ );
nand g282 ( new_n388_, new_n380_, new_n384_, new_n381_, new_n385_ );
nand g283 ( new_n389_, new_n387_, new_n388_ );
not g284 ( new_n390_, new_n389_ );
nand g285 ( new_n391_, new_n379_, new_n390_ );
nand g286 ( new_n392_, new_n377_, new_n378_, new_n389_ );
nand g287 ( new_n393_, new_n391_, new_n392_ );
nand g288 ( new_n394_, new_n393_, new_n349_ );
not g289 ( new_n395_, new_n393_ );
nand g290 ( new_n396_, new_n395_, keyIn_0_14 );
nand g291 ( new_n397_, new_n256_, N1 );
nand g292 ( new_n398_, new_n143_, N5 );
nand g293 ( new_n399_, new_n397_, new_n398_ );
nand g294 ( new_n400_, new_n235_, new_n185_ );
nand g295 ( new_n401_, N9, N13 );
nand g296 ( new_n402_, new_n400_, new_n401_ );
nand g297 ( new_n403_, new_n399_, new_n402_ );
nand g298 ( new_n404_, new_n400_, new_n397_, new_n398_, new_n401_ );
nand g299 ( new_n405_, new_n403_, new_n404_ );
nand g300 ( new_n406_, new_n317_, new_n405_ );
not g301 ( new_n407_, new_n405_ );
nand g302 ( new_n408_, new_n316_, new_n407_, new_n314_ );
nand g303 ( new_n409_, new_n406_, new_n408_ );
nand g304 ( new_n410_, N133, N137 );
nand g305 ( new_n411_, new_n409_, new_n410_ );
nand g306 ( new_n412_, new_n406_, N133, N137, new_n408_ );
nand g307 ( new_n413_, new_n411_, new_n412_ );
nand g308 ( new_n414_, new_n108_, N65 );
nand g309 ( new_n415_, new_n122_, N81 );
nand g310 ( new_n416_, new_n414_, new_n415_ );
not g311 ( new_n417_, N113 );
nand g312 ( new_n418_, new_n210_, new_n417_ );
nand g313 ( new_n419_, N97, N113 );
nand g314 ( new_n420_, new_n418_, new_n419_ );
nand g315 ( new_n421_, new_n416_, new_n420_ );
nand g316 ( new_n422_, new_n418_, new_n414_, new_n415_, new_n419_ );
nand g317 ( new_n423_, new_n421_, new_n422_ );
nand g318 ( new_n424_, new_n413_, new_n423_ );
nand g319 ( new_n425_, new_n411_, new_n412_, new_n421_, new_n422_ );
nand g320 ( new_n426_, new_n424_, new_n425_ );
not g321 ( new_n427_, new_n426_ );
nand g322 ( new_n428_, new_n371_, new_n407_ );
nand g323 ( new_n429_, new_n368_, new_n370_, new_n405_ );
nand g324 ( new_n430_, new_n428_, new_n429_ );
nand g325 ( new_n431_, N135, N137 );
nand g326 ( new_n432_, new_n431_, keyIn_0_5 );
not g327 ( new_n433_, keyIn_0_5 );
nand g328 ( new_n434_, new_n433_, N135, N137 );
nand g329 ( new_n435_, new_n432_, new_n434_ );
nand g330 ( new_n436_, new_n430_, new_n435_ );
nand g331 ( new_n437_, new_n428_, new_n429_, new_n432_, new_n434_ );
nand g332 ( new_n438_, new_n436_, new_n437_ );
nor g333 ( new_n439_, N105, N121 );
not g334 ( new_n440_, new_n439_ );
nand g335 ( new_n441_, N105, N121 );
nand g336 ( new_n442_, new_n440_, new_n441_ );
nand g337 ( new_n443_, new_n442_, keyIn_0_7 );
not g338 ( new_n444_, new_n443_ );
nor g339 ( new_n445_, new_n442_, keyIn_0_7 );
nor g340 ( new_n446_, new_n444_, new_n445_ );
not g341 ( new_n447_, new_n446_ );
nand g342 ( new_n448_, N73, N89 );
not g343 ( new_n449_, new_n448_ );
nor g344 ( new_n450_, N73, N89 );
nor g345 ( new_n451_, new_n449_, new_n450_ );
not g346 ( new_n452_, new_n451_ );
nand g347 ( new_n453_, new_n447_, new_n452_ );
nand g348 ( new_n454_, new_n446_, new_n451_ );
nand g349 ( new_n455_, new_n453_, new_n454_ );
nand g350 ( new_n456_, new_n438_, new_n455_ );
nand g351 ( new_n457_, new_n436_, new_n437_, new_n453_, new_n454_ );
nand g352 ( new_n458_, new_n456_, new_n457_ );
not g353 ( new_n459_, new_n458_ );
nand g354 ( new_n460_, new_n396_, new_n394_, new_n427_, new_n459_ );
not g355 ( new_n461_, new_n460_ );
nand g356 ( new_n462_, new_n291_, new_n348_, new_n461_ );
nand g357 ( new_n463_, new_n462_, new_n162_ );
nand g358 ( new_n464_, new_n291_, keyIn_0_24, new_n348_, new_n461_ );
nand g359 ( new_n465_, new_n463_, new_n161_, new_n464_ );
nand g360 ( new_n466_, new_n465_, N1 );
nand g361 ( new_n467_, new_n463_, new_n143_, new_n161_, new_n464_ );
nand g362 ( N724, new_n466_, new_n467_ );
nand g363 ( new_n469_, new_n463_, new_n271_, new_n464_ );
nand g364 ( new_n470_, new_n469_, N5 );
nand g365 ( new_n471_, new_n463_, new_n256_, new_n271_, new_n464_ );
nand g366 ( N725, new_n470_, new_n471_ );
nand g367 ( new_n473_, new_n463_, new_n277_, new_n464_ );
nand g368 ( new_n474_, new_n473_, N9 );
nand g369 ( new_n475_, new_n463_, new_n235_, new_n277_, new_n464_ );
nand g370 ( new_n476_, new_n474_, new_n475_ );
nand g371 ( new_n477_, new_n476_, keyIn_0_30 );
not g372 ( new_n478_, keyIn_0_30 );
nand g373 ( new_n479_, new_n474_, new_n478_, new_n475_ );
nand g374 ( N726, new_n477_, new_n479_ );
not g375 ( new_n481_, new_n201_ );
nand g376 ( new_n482_, new_n463_, new_n481_, new_n464_ );
nand g377 ( new_n483_, new_n482_, N13 );
nand g378 ( new_n484_, new_n463_, new_n185_, new_n481_, new_n464_ );
nand g379 ( new_n485_, new_n483_, new_n484_ );
nand g380 ( new_n486_, new_n485_, keyIn_0_31 );
not g381 ( new_n487_, keyIn_0_31 );
nand g382 ( new_n488_, new_n483_, new_n487_, new_n484_ );
nand g383 ( N727, new_n486_, new_n488_ );
nand g384 ( new_n490_, new_n393_, new_n427_ );
not g385 ( new_n491_, new_n490_ );
nand g386 ( new_n492_, new_n458_, new_n343_ );
not g387 ( new_n493_, new_n492_ );
nand g388 ( new_n494_, new_n291_, new_n493_ );
not g389 ( new_n495_, new_n494_ );
nand g390 ( new_n496_, new_n495_, new_n491_ );
not g391 ( new_n497_, new_n496_ );
nand g392 ( new_n498_, new_n497_, new_n161_ );
nand g393 ( new_n499_, new_n498_, N17 );
nand g394 ( new_n500_, new_n497_, new_n141_, new_n161_ );
nand g395 ( N728, new_n499_, new_n500_ );
nand g396 ( new_n502_, new_n497_, new_n271_ );
nand g397 ( new_n503_, new_n502_, N21 );
nand g398 ( new_n504_, new_n497_, new_n257_, new_n271_ );
nand g399 ( N729, new_n503_, new_n504_ );
nand g400 ( new_n506_, new_n497_, new_n277_ );
nand g401 ( new_n507_, new_n506_, keyIn_0_25 );
not g402 ( new_n508_, keyIn_0_25 );
nand g403 ( new_n509_, new_n497_, new_n508_, new_n277_ );
nand g404 ( new_n510_, new_n507_, new_n509_ );
nand g405 ( new_n511_, new_n510_, new_n237_ );
nand g406 ( new_n512_, new_n507_, N25, new_n509_ );
nand g407 ( N730, new_n511_, new_n512_ );
nand g408 ( new_n514_, new_n497_, new_n481_ );
nand g409 ( new_n515_, new_n514_, keyIn_0_26 );
not g410 ( new_n516_, keyIn_0_26 );
nand g411 ( new_n517_, new_n497_, new_n516_, new_n481_ );
nand g412 ( new_n518_, new_n515_, new_n517_ );
nand g413 ( new_n519_, new_n518_, N29 );
nand g414 ( new_n520_, new_n515_, new_n186_, new_n517_ );
nand g415 ( N731, new_n519_, new_n520_ );
nand g416 ( new_n522_, new_n456_, new_n341_, new_n342_, new_n457_ );
not g417 ( new_n523_, new_n522_ );
nand g418 ( new_n524_, new_n427_, keyIn_0_16 );
not g419 ( new_n525_, keyIn_0_16 );
nand g420 ( new_n526_, new_n426_, new_n525_ );
nand g421 ( new_n527_, new_n395_, new_n524_, new_n526_ );
not g422 ( new_n528_, new_n527_ );
nand g423 ( new_n529_, new_n291_, new_n523_, new_n528_ );
not g424 ( new_n530_, new_n529_ );
nand g425 ( new_n531_, new_n530_, new_n161_ );
nand g426 ( new_n532_, new_n531_, N33 );
nand g427 ( new_n533_, new_n530_, new_n146_, new_n161_ );
nand g428 ( N732, new_n532_, new_n533_ );
nand g429 ( new_n535_, new_n530_, new_n271_ );
nand g430 ( new_n536_, new_n535_, N37 );
nand g431 ( new_n537_, new_n530_, new_n261_, new_n271_ );
nand g432 ( N733, new_n536_, new_n537_ );
nand g433 ( new_n539_, new_n530_, new_n277_ );
nand g434 ( new_n540_, new_n539_, N41 );
nand g435 ( new_n541_, new_n530_, new_n353_, new_n277_ );
nand g436 ( N734, new_n540_, new_n541_ );
nand g437 ( new_n543_, new_n530_, new_n481_ );
nand g438 ( new_n544_, new_n543_, N45 );
nand g439 ( new_n545_, new_n530_, new_n190_, new_n481_ );
nand g440 ( N735, new_n544_, new_n545_ );
nand g441 ( new_n547_, new_n427_, keyIn_0_17 );
not g442 ( new_n548_, keyIn_0_17 );
nand g443 ( new_n549_, new_n426_, new_n548_ );
nand g444 ( new_n550_, new_n547_, new_n549_ );
nand g445 ( new_n551_, new_n495_, new_n395_, new_n550_ );
not g446 ( new_n552_, new_n551_ );
nand g447 ( new_n553_, new_n552_, new_n161_ );
nand g448 ( new_n554_, new_n553_, N49 );
nand g449 ( new_n555_, new_n552_, new_n147_, new_n161_ );
nand g450 ( N736, new_n554_, new_n555_ );
nand g451 ( new_n557_, new_n552_, new_n271_ );
nand g452 ( new_n558_, new_n557_, N53 );
nand g453 ( new_n559_, new_n552_, new_n262_, new_n271_ );
nand g454 ( N737, new_n558_, new_n559_ );
nand g455 ( new_n561_, new_n552_, new_n277_ );
nand g456 ( new_n562_, new_n561_, N57 );
nand g457 ( new_n563_, new_n552_, new_n296_, new_n277_ );
nand g458 ( N738, new_n562_, new_n563_ );
nand g459 ( new_n565_, new_n552_, new_n481_ );
nand g460 ( new_n566_, new_n565_, N61 );
nand g461 ( new_n567_, new_n552_, new_n191_, new_n481_ );
nand g462 ( N739, new_n566_, new_n567_ );
nand g463 ( new_n569_, new_n393_, new_n458_, new_n343_, new_n426_ );
nand g464 ( new_n570_, new_n569_, keyIn_0_20 );
not g465 ( new_n571_, keyIn_0_20 );
nand g466 ( new_n572_, new_n393_, new_n426_ );
not g467 ( new_n573_, new_n572_ );
nand g468 ( new_n574_, new_n493_, new_n573_, new_n571_ );
nand g469 ( new_n575_, new_n574_, new_n570_ );
nand g470 ( new_n576_, new_n458_, keyIn_0_18 );
not g471 ( new_n577_, keyIn_0_18 );
nand g472 ( new_n578_, new_n456_, new_n577_, new_n457_ );
nand g473 ( new_n579_, new_n576_, new_n578_ );
nand g474 ( new_n580_, new_n579_, new_n344_, new_n491_ );
nand g475 ( new_n581_, new_n459_, new_n344_, new_n393_, new_n426_ );
nand g476 ( new_n582_, new_n581_, keyIn_0_21 );
not g477 ( new_n583_, keyIn_0_21 );
nand g478 ( new_n584_, new_n573_, new_n583_, new_n523_ );
nand g479 ( new_n585_, new_n582_, new_n584_ );
nand g480 ( new_n586_, new_n341_, new_n342_, new_n426_ );
not g481 ( new_n587_, new_n586_ );
nand g482 ( new_n588_, new_n587_, new_n395_, new_n458_ );
nand g483 ( new_n589_, new_n588_, keyIn_0_22 );
not g484 ( new_n590_, keyIn_0_22 );
nand g485 ( new_n591_, new_n587_, new_n395_, new_n590_, new_n458_ );
nand g486 ( new_n592_, new_n589_, new_n591_ );
nand g487 ( new_n593_, new_n585_, new_n575_, new_n592_, new_n580_ );
nand g488 ( new_n594_, new_n593_, keyIn_0_23 );
not g489 ( new_n595_, keyIn_0_23 );
not g490 ( new_n596_, new_n570_ );
nor g491 ( new_n597_, new_n569_, keyIn_0_20 );
nor g492 ( new_n598_, new_n596_, new_n597_ );
not g493 ( new_n599_, new_n580_ );
nor g494 ( new_n600_, new_n598_, new_n599_ );
nand g495 ( new_n601_, new_n585_, new_n592_ );
not g496 ( new_n602_, new_n601_ );
nand g497 ( new_n603_, new_n602_, new_n600_, new_n595_ );
nand g498 ( new_n604_, new_n603_, new_n594_ );
nand g499 ( new_n605_, new_n201_, new_n277_ );
not g500 ( new_n606_, new_n605_ );
nand g501 ( new_n607_, new_n604_, new_n161_, new_n273_, new_n606_ );
not g502 ( new_n608_, new_n607_ );
nand g503 ( new_n609_, new_n608_, new_n427_ );
nand g504 ( new_n610_, new_n609_, N65 );
nand g505 ( new_n611_, new_n608_, new_n122_, new_n427_ );
nand g506 ( N740, new_n610_, new_n611_ );
nand g507 ( new_n613_, new_n608_, new_n395_ );
nand g508 ( new_n614_, new_n613_, N69 );
nand g509 ( new_n615_, new_n608_, new_n120_, new_n395_ );
nand g510 ( N741, new_n614_, new_n615_ );
nand g511 ( new_n617_, new_n608_, new_n459_ );
nand g512 ( new_n618_, new_n617_, N73 );
nand g513 ( new_n619_, new_n608_, new_n125_, new_n459_ );
nand g514 ( N742, new_n618_, new_n619_ );
nand g515 ( new_n621_, new_n608_, new_n343_ );
nand g516 ( new_n622_, new_n621_, N77 );
nand g517 ( new_n623_, new_n608_, new_n126_, new_n343_ );
nand g518 ( N743, new_n622_, new_n623_ );
nor g519 ( new_n625_, new_n201_, new_n277_, new_n271_, new_n160_ );
nand g520 ( new_n626_, new_n604_, new_n625_ );
not g521 ( new_n627_, new_n626_ );
nand g522 ( new_n628_, new_n627_, new_n427_ );
nand g523 ( new_n629_, new_n628_, N81 );
nand g524 ( new_n630_, new_n627_, new_n108_, new_n427_ );
nand g525 ( N744, new_n629_, new_n630_ );
not g526 ( new_n632_, keyIn_0_27 );
nand g527 ( new_n633_, new_n604_, new_n395_, new_n625_ );
nand g528 ( new_n634_, new_n633_, new_n632_ );
nand g529 ( new_n635_, new_n604_, keyIn_0_27, new_n395_, new_n625_ );
nand g530 ( new_n636_, new_n634_, new_n635_ );
nand g531 ( new_n637_, new_n636_, new_n106_ );
nand g532 ( new_n638_, new_n634_, N85, new_n635_ );
nand g533 ( N745, new_n637_, new_n638_ );
nand g534 ( new_n640_, new_n627_, new_n459_ );
nand g535 ( new_n641_, new_n640_, N89 );
nand g536 ( new_n642_, new_n627_, new_n111_, new_n459_ );
nand g537 ( N746, new_n641_, new_n642_ );
nand g538 ( new_n644_, new_n627_, new_n343_ );
nand g539 ( new_n645_, new_n644_, N93 );
nand g540 ( new_n646_, new_n627_, new_n112_, new_n343_ );
nand g541 ( N747, new_n645_, new_n646_ );
nand g542 ( new_n648_, new_n606_, new_n160_, new_n271_ );
not g543 ( new_n649_, new_n648_ );
nand g544 ( new_n650_, new_n604_, new_n649_ );
not g545 ( new_n651_, new_n650_ );
nand g546 ( new_n652_, new_n651_, new_n427_ );
nand g547 ( new_n653_, new_n652_, N97 );
nand g548 ( new_n654_, new_n651_, new_n210_, new_n427_ );
nand g549 ( N748, new_n653_, new_n654_ );
nand g550 ( new_n656_, new_n651_, new_n395_ );
nand g551 ( new_n657_, new_n656_, N101 );
nand g552 ( new_n658_, new_n651_, new_n211_, new_n395_ );
nand g553 ( N749, new_n657_, new_n658_ );
nand g554 ( new_n660_, new_n651_, new_n459_ );
nand g555 ( new_n661_, new_n660_, N105 );
not g556 ( new_n662_, N105 );
nand g557 ( new_n663_, new_n651_, new_n662_, new_n459_ );
nand g558 ( N750, new_n661_, new_n663_ );
nand g559 ( new_n665_, new_n604_, new_n343_, new_n649_ );
nand g560 ( new_n666_, new_n665_, keyIn_0_28 );
not g561 ( new_n667_, keyIn_0_28 );
nand g562 ( new_n668_, new_n604_, new_n667_, new_n343_, new_n649_ );
nand g563 ( new_n669_, new_n666_, new_n668_ );
nand g564 ( new_n670_, new_n669_, new_n333_ );
nand g565 ( new_n671_, new_n666_, N109, new_n668_ );
nand g566 ( N751, new_n670_, new_n671_ );
nor g567 ( new_n673_, new_n273_, new_n201_, new_n277_, new_n161_ );
nand g568 ( new_n674_, new_n604_, new_n673_ );
not g569 ( new_n675_, new_n674_ );
nand g570 ( new_n676_, new_n675_, new_n427_ );
nand g571 ( new_n677_, new_n676_, N113 );
nand g572 ( new_n678_, new_n675_, new_n417_, new_n427_ );
nand g573 ( N752, new_n677_, new_n678_ );
nand g574 ( new_n680_, new_n604_, new_n395_, new_n673_ );
nand g575 ( new_n681_, new_n680_, keyIn_0_29 );
not g576 ( new_n682_, keyIn_0_29 );
nand g577 ( new_n683_, new_n604_, new_n682_, new_n395_, new_n673_ );
nand g578 ( new_n684_, new_n681_, new_n683_ );
nand g579 ( new_n685_, new_n684_, N117 );
nand g580 ( new_n686_, new_n681_, new_n383_, new_n683_ );
nand g581 ( N753, new_n685_, new_n686_ );
nand g582 ( new_n688_, new_n675_, new_n459_ );
nand g583 ( new_n689_, new_n688_, N121 );
not g584 ( new_n690_, N121 );
nand g585 ( new_n691_, new_n675_, new_n690_, new_n459_ );
nand g586 ( N754, new_n689_, new_n691_ );
nand g587 ( new_n693_, new_n675_, new_n343_ );
nand g588 ( new_n694_, new_n693_, N125 );
nand g589 ( new_n695_, new_n675_, new_n334_, new_n343_ );
nand g590 ( N755, new_n694_, new_n695_ );
endmodule