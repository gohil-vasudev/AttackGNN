module add_mul_mix_8_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, c_0_, c_1_, c_2_, c_3_, 
        c_4_, c_5_, c_6_, c_7_, d_0_, d_1_, d_2_, d_3_, d_4_, d_5_, d_6_, d_7_, 
        Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_, 
        Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_, 
        Result_12_, Result_13_, Result_14_, Result_15_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_,
         b_4_, b_5_, b_6_, b_7_, c_0_, c_1_, c_2_, c_3_, c_4_, c_5_, c_6_,
         c_7_, d_0_, d_1_, d_2_, d_3_, d_4_, d_5_, d_6_, d_7_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_;
  wire   n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958;

  XNOR2_X1 U492 ( .A(n477), .B(n478), .ZN(Result_9_) );
  XOR2_X1 U493 ( .A(n479), .B(n480), .Z(n478) );
  XNOR2_X1 U494 ( .A(n481), .B(n482), .ZN(Result_8_) );
  XOR2_X1 U495 ( .A(n483), .B(n484), .Z(n482) );
  XOR2_X1 U496 ( .A(n485), .B(n486), .Z(Result_7_) );
  AND2_X1 U497 ( .A1(n487), .A2(n488), .ZN(Result_6_) );
  OR2_X1 U498 ( .A1(n489), .A2(n490), .ZN(n487) );
  XOR2_X1 U499 ( .A(n491), .B(n492), .Z(n490) );
  INV_X1 U500 ( .A(n493), .ZN(n489) );
  XNOR2_X1 U501 ( .A(n494), .B(n495), .ZN(Result_5_) );
  AND2_X1 U502 ( .A1(n488), .A2(n496), .ZN(n495) );
  XOR2_X1 U503 ( .A(n497), .B(n498), .Z(Result_4_) );
  XOR2_X1 U504 ( .A(n499), .B(n500), .Z(Result_3_) );
  OR2_X1 U505 ( .A1(n501), .A2(n502), .ZN(n500) );
  INV_X1 U506 ( .A(n503), .ZN(n502) );
  AND2_X1 U507 ( .A1(n504), .A2(n505), .ZN(n501) );
  XOR2_X1 U508 ( .A(n506), .B(n507), .Z(Result_2_) );
  XOR2_X1 U509 ( .A(n508), .B(n509), .Z(Result_1_) );
  OR2_X1 U510 ( .A1(n510), .A2(n511), .ZN(n509) );
  INV_X1 U511 ( .A(n512), .ZN(n511) );
  AND2_X1 U512 ( .A1(n513), .A2(n514), .ZN(n510) );
  OR2_X1 U513 ( .A1(n515), .A2(n516), .ZN(n514) );
  INV_X1 U514 ( .A(n517), .ZN(Result_15_) );
  XOR2_X1 U515 ( .A(n518), .B(n519), .Z(Result_14_) );
  OR2_X1 U516 ( .A1(n520), .A2(n521), .ZN(n519) );
  XNOR2_X1 U517 ( .A(n522), .B(n523), .ZN(Result_13_) );
  XOR2_X1 U518 ( .A(n524), .B(n525), .Z(n523) );
  XOR2_X1 U519 ( .A(n526), .B(n527), .Z(Result_12_) );
  XNOR2_X1 U520 ( .A(n528), .B(n529), .ZN(n527) );
  XNOR2_X1 U521 ( .A(n530), .B(n531), .ZN(Result_11_) );
  XOR2_X1 U522 ( .A(n532), .B(n533), .Z(n531) );
  XNOR2_X1 U523 ( .A(n534), .B(n535), .ZN(Result_10_) );
  XOR2_X1 U524 ( .A(n536), .B(n537), .Z(n535) );
  INV_X1 U525 ( .A(n538), .ZN(Result_0_) );
  AND2_X1 U526 ( .A1(n539), .A2(n540), .ZN(n538) );
  AND2_X1 U527 ( .A1(n512), .A2(n541), .ZN(n540) );
  OR2_X1 U528 ( .A1(n508), .A2(n513), .ZN(n541) );
  OR2_X1 U529 ( .A1(n507), .A2(n506), .ZN(n508) );
  XNOR2_X1 U530 ( .A(n515), .B(n516), .ZN(n506) );
  AND2_X1 U531 ( .A1(n542), .A2(n543), .ZN(n507) );
  AND2_X1 U532 ( .A1(n544), .A2(n503), .ZN(n542) );
  OR2_X1 U533 ( .A1(n505), .A2(n504), .ZN(n503) );
  OR2_X1 U534 ( .A1(n545), .A2(n546), .ZN(n504) );
  OR2_X1 U535 ( .A1(n499), .A2(n505), .ZN(n544) );
  OR2_X1 U536 ( .A1(n547), .A2(n548), .ZN(n505) );
  INV_X1 U537 ( .A(n543), .ZN(n548) );
  OR2_X1 U538 ( .A1(n549), .A2(n550), .ZN(n543) );
  AND2_X1 U539 ( .A1(n549), .A2(n550), .ZN(n547) );
  OR2_X1 U540 ( .A1(n551), .A2(n552), .ZN(n550) );
  AND2_X1 U541 ( .A1(n553), .A2(n554), .ZN(n552) );
  AND2_X1 U542 ( .A1(n555), .A2(n556), .ZN(n551) );
  OR2_X1 U543 ( .A1(n554), .A2(n553), .ZN(n556) );
  XOR2_X1 U544 ( .A(n557), .B(n558), .Z(n549) );
  XOR2_X1 U545 ( .A(n559), .B(n560), .Z(n558) );
  OR2_X1 U546 ( .A1(n498), .A2(n497), .ZN(n499) );
  XNOR2_X1 U547 ( .A(n545), .B(n546), .ZN(n497) );
  OR2_X1 U548 ( .A1(n561), .A2(n562), .ZN(n546) );
  AND2_X1 U549 ( .A1(n563), .A2(n564), .ZN(n562) );
  AND2_X1 U550 ( .A1(n565), .A2(n566), .ZN(n561) );
  OR2_X1 U551 ( .A1(n564), .A2(n563), .ZN(n566) );
  XNOR2_X1 U552 ( .A(n567), .B(n555), .ZN(n545) );
  XOR2_X1 U553 ( .A(n568), .B(n569), .Z(n555) );
  XOR2_X1 U554 ( .A(n570), .B(n571), .Z(n569) );
  XNOR2_X1 U555 ( .A(n554), .B(n553), .ZN(n567) );
  OR2_X1 U556 ( .A1(n572), .A2(n573), .ZN(n553) );
  AND2_X1 U557 ( .A1(n574), .A2(n575), .ZN(n573) );
  AND2_X1 U558 ( .A1(n576), .A2(n577), .ZN(n572) );
  OR2_X1 U559 ( .A1(n575), .A2(n574), .ZN(n577) );
  OR2_X1 U560 ( .A1(n578), .A2(n579), .ZN(n554) );
  AND2_X1 U561 ( .A1(n580), .A2(n581), .ZN(n498) );
  INV_X1 U562 ( .A(n582), .ZN(n580) );
  OR2_X1 U563 ( .A1(n583), .A2(n584), .ZN(n582) );
  AND2_X1 U564 ( .A1(n585), .A2(n494), .ZN(n584) );
  AND2_X1 U565 ( .A1(n586), .A2(n494), .ZN(n583) );
  AND2_X1 U566 ( .A1(n587), .A2(n581), .ZN(n494) );
  OR2_X1 U567 ( .A1(n588), .A2(n589), .ZN(n581) );
  INV_X1 U568 ( .A(n590), .ZN(n587) );
  AND2_X1 U569 ( .A1(n588), .A2(n589), .ZN(n590) );
  OR2_X1 U570 ( .A1(n591), .A2(n592), .ZN(n589) );
  AND2_X1 U571 ( .A1(n593), .A2(n594), .ZN(n592) );
  AND2_X1 U572 ( .A1(n595), .A2(n596), .ZN(n591) );
  OR2_X1 U573 ( .A1(n594), .A2(n593), .ZN(n595) );
  XOR2_X1 U574 ( .A(n565), .B(n597), .Z(n588) );
  XOR2_X1 U575 ( .A(n564), .B(n563), .Z(n597) );
  OR2_X1 U576 ( .A1(n598), .A2(n579), .ZN(n563) );
  OR2_X1 U577 ( .A1(n599), .A2(n600), .ZN(n564) );
  AND2_X1 U578 ( .A1(n601), .A2(n602), .ZN(n600) );
  AND2_X1 U579 ( .A1(n603), .A2(n604), .ZN(n599) );
  OR2_X1 U580 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U581 ( .A(n605), .B(n576), .ZN(n565) );
  XNOR2_X1 U582 ( .A(n606), .B(n607), .ZN(n576) );
  XNOR2_X1 U583 ( .A(n608), .B(n609), .ZN(n606) );
  XNOR2_X1 U584 ( .A(n575), .B(n574), .ZN(n605) );
  OR2_X1 U585 ( .A1(n610), .A2(n611), .ZN(n574) );
  AND2_X1 U586 ( .A1(n612), .A2(n613), .ZN(n611) );
  AND2_X1 U587 ( .A1(n614), .A2(n615), .ZN(n610) );
  OR2_X1 U588 ( .A1(n613), .A2(n612), .ZN(n615) );
  OR2_X1 U589 ( .A1(n578), .A2(n616), .ZN(n575) );
  INV_X1 U590 ( .A(n488), .ZN(n586) );
  OR2_X1 U591 ( .A1(n617), .A2(n493), .ZN(n488) );
  OR2_X1 U592 ( .A1(n486), .A2(n485), .ZN(n493) );
  OR2_X1 U593 ( .A1(n618), .A2(n619), .ZN(n485) );
  AND2_X1 U594 ( .A1(n484), .A2(n483), .ZN(n619) );
  AND2_X1 U595 ( .A1(n481), .A2(n620), .ZN(n618) );
  OR2_X1 U596 ( .A1(n483), .A2(n484), .ZN(n620) );
  OR2_X1 U597 ( .A1(n520), .A2(n579), .ZN(n484) );
  OR2_X1 U598 ( .A1(n621), .A2(n622), .ZN(n483) );
  AND2_X1 U599 ( .A1(n480), .A2(n479), .ZN(n622) );
  AND2_X1 U600 ( .A1(n477), .A2(n623), .ZN(n621) );
  OR2_X1 U601 ( .A1(n479), .A2(n480), .ZN(n623) );
  OR2_X1 U602 ( .A1(n616), .A2(n520), .ZN(n480) );
  OR2_X1 U603 ( .A1(n624), .A2(n625), .ZN(n479) );
  AND2_X1 U604 ( .A1(n537), .A2(n536), .ZN(n625) );
  AND2_X1 U605 ( .A1(n534), .A2(n626), .ZN(n624) );
  OR2_X1 U606 ( .A1(n537), .A2(n536), .ZN(n626) );
  OR2_X1 U607 ( .A1(n627), .A2(n628), .ZN(n536) );
  AND2_X1 U608 ( .A1(n533), .A2(n532), .ZN(n628) );
  AND2_X1 U609 ( .A1(n530), .A2(n629), .ZN(n627) );
  OR2_X1 U610 ( .A1(n533), .A2(n532), .ZN(n629) );
  OR2_X1 U611 ( .A1(n630), .A2(n631), .ZN(n532) );
  AND2_X1 U612 ( .A1(n528), .A2(n529), .ZN(n631) );
  AND2_X1 U613 ( .A1(n526), .A2(n632), .ZN(n630) );
  OR2_X1 U614 ( .A1(n528), .A2(n529), .ZN(n632) );
  OR2_X1 U615 ( .A1(n633), .A2(n634), .ZN(n529) );
  AND2_X1 U616 ( .A1(n525), .A2(n524), .ZN(n634) );
  AND2_X1 U617 ( .A1(n522), .A2(n635), .ZN(n633) );
  OR2_X1 U618 ( .A1(n525), .A2(n524), .ZN(n635) );
  OR2_X1 U619 ( .A1(n636), .A2(n520), .ZN(n524) );
  OR2_X1 U620 ( .A1(n637), .A2(n517), .ZN(n525) );
  OR2_X1 U621 ( .A1(n638), .A2(n520), .ZN(n517) );
  XNOR2_X1 U622 ( .A(n637), .B(n639), .ZN(n522) );
  OR2_X1 U623 ( .A1(n640), .A2(n638), .ZN(n639) );
  OR2_X1 U624 ( .A1(n521), .A2(n641), .ZN(n637) );
  OR2_X1 U625 ( .A1(n642), .A2(n520), .ZN(n528) );
  XNOR2_X1 U626 ( .A(n643), .B(n644), .ZN(n526) );
  XNOR2_X1 U627 ( .A(n645), .B(n646), .ZN(n643) );
  OR2_X1 U628 ( .A1(n647), .A2(n520), .ZN(n533) );
  XOR2_X1 U629 ( .A(n648), .B(n649), .Z(n530) );
  XOR2_X1 U630 ( .A(n650), .B(n651), .Z(n649) );
  OR2_X1 U631 ( .A1(n652), .A2(n520), .ZN(n537) );
  OR2_X1 U632 ( .A1(n653), .A2(n654), .ZN(n520) );
  INV_X1 U633 ( .A(n655), .ZN(n653) );
  OR2_X1 U634 ( .A1(c_7_), .A2(d_7_), .ZN(n655) );
  XOR2_X1 U635 ( .A(n656), .B(n657), .Z(n534) );
  XOR2_X1 U636 ( .A(n658), .B(n659), .Z(n657) );
  XOR2_X1 U637 ( .A(n660), .B(n661), .Z(n477) );
  XOR2_X1 U638 ( .A(n662), .B(n663), .Z(n661) );
  XOR2_X1 U639 ( .A(n664), .B(n665), .Z(n481) );
  XOR2_X1 U640 ( .A(n666), .B(n667), .Z(n665) );
  XOR2_X1 U641 ( .A(n668), .B(n669), .Z(n486) );
  XOR2_X1 U642 ( .A(n670), .B(n671), .Z(n669) );
  OR2_X1 U643 ( .A1(n585), .A2(n672), .ZN(n617) );
  AND2_X1 U644 ( .A1(n491), .A2(n492), .ZN(n672) );
  INV_X1 U645 ( .A(n496), .ZN(n585) );
  OR2_X1 U646 ( .A1(n491), .A2(n492), .ZN(n496) );
  OR2_X1 U647 ( .A1(n673), .A2(n674), .ZN(n492) );
  AND2_X1 U648 ( .A1(n671), .A2(n670), .ZN(n674) );
  AND2_X1 U649 ( .A1(n668), .A2(n675), .ZN(n673) );
  OR2_X1 U650 ( .A1(n670), .A2(n671), .ZN(n675) );
  OR2_X1 U651 ( .A1(n641), .A2(n579), .ZN(n671) );
  OR2_X1 U652 ( .A1(n676), .A2(n677), .ZN(n670) );
  AND2_X1 U653 ( .A1(n667), .A2(n666), .ZN(n677) );
  AND2_X1 U654 ( .A1(n664), .A2(n678), .ZN(n676) );
  OR2_X1 U655 ( .A1(n666), .A2(n667), .ZN(n678) );
  OR2_X1 U656 ( .A1(n641), .A2(n616), .ZN(n667) );
  OR2_X1 U657 ( .A1(n679), .A2(n680), .ZN(n666) );
  AND2_X1 U658 ( .A1(n663), .A2(n662), .ZN(n680) );
  AND2_X1 U659 ( .A1(n660), .A2(n681), .ZN(n679) );
  OR2_X1 U660 ( .A1(n662), .A2(n663), .ZN(n681) );
  OR2_X1 U661 ( .A1(n641), .A2(n652), .ZN(n663) );
  OR2_X1 U662 ( .A1(n682), .A2(n683), .ZN(n662) );
  AND2_X1 U663 ( .A1(n659), .A2(n658), .ZN(n683) );
  AND2_X1 U664 ( .A1(n656), .A2(n684), .ZN(n682) );
  OR2_X1 U665 ( .A1(n659), .A2(n658), .ZN(n684) );
  OR2_X1 U666 ( .A1(n685), .A2(n686), .ZN(n658) );
  AND2_X1 U667 ( .A1(n651), .A2(n650), .ZN(n686) );
  AND2_X1 U668 ( .A1(n648), .A2(n687), .ZN(n685) );
  OR2_X1 U669 ( .A1(n651), .A2(n650), .ZN(n687) );
  OR2_X1 U670 ( .A1(n688), .A2(n689), .ZN(n650) );
  AND2_X1 U671 ( .A1(n644), .A2(n646), .ZN(n689) );
  AND2_X1 U672 ( .A1(n690), .A2(n645), .ZN(n688) );
  OR2_X1 U673 ( .A1(n691), .A2(n692), .ZN(n645) );
  INV_X1 U674 ( .A(n693), .ZN(n692) );
  AND2_X1 U675 ( .A1(n694), .A2(n695), .ZN(n691) );
  OR2_X1 U676 ( .A1(n644), .A2(n646), .ZN(n690) );
  OR2_X1 U677 ( .A1(n695), .A2(n518), .ZN(n646) );
  OR2_X1 U678 ( .A1(n641), .A2(n638), .ZN(n518) );
  OR2_X1 U679 ( .A1(n641), .A2(n636), .ZN(n644) );
  OR2_X1 U680 ( .A1(n642), .A2(n641), .ZN(n651) );
  XNOR2_X1 U681 ( .A(n696), .B(n697), .ZN(n648) );
  XNOR2_X1 U682 ( .A(n698), .B(n693), .ZN(n696) );
  OR2_X1 U683 ( .A1(n647), .A2(n641), .ZN(n659) );
  XNOR2_X1 U684 ( .A(n654), .B(n699), .ZN(n641) );
  XOR2_X1 U685 ( .A(d_6_), .B(c_6_), .Z(n699) );
  XOR2_X1 U686 ( .A(n700), .B(n701), .Z(n656) );
  XOR2_X1 U687 ( .A(n702), .B(n703), .Z(n701) );
  XOR2_X1 U688 ( .A(n704), .B(n705), .Z(n660) );
  XOR2_X1 U689 ( .A(n706), .B(n707), .Z(n705) );
  XOR2_X1 U690 ( .A(n708), .B(n709), .Z(n664) );
  XOR2_X1 U691 ( .A(n710), .B(n711), .Z(n709) );
  XOR2_X1 U692 ( .A(n712), .B(n713), .Z(n668) );
  XOR2_X1 U693 ( .A(n714), .B(n715), .Z(n713) );
  XNOR2_X1 U694 ( .A(n716), .B(n593), .ZN(n491) );
  XNOR2_X1 U695 ( .A(n717), .B(n601), .ZN(n593) );
  XNOR2_X1 U696 ( .A(n718), .B(n614), .ZN(n601) );
  XNOR2_X1 U697 ( .A(n719), .B(n720), .ZN(n614) );
  XNOR2_X1 U698 ( .A(n721), .B(n722), .ZN(n719) );
  XNOR2_X1 U699 ( .A(n613), .B(n612), .ZN(n718) );
  OR2_X1 U700 ( .A1(n723), .A2(n724), .ZN(n612) );
  AND2_X1 U701 ( .A1(n725), .A2(n726), .ZN(n724) );
  AND2_X1 U702 ( .A1(n727), .A2(n728), .ZN(n723) );
  OR2_X1 U703 ( .A1(n726), .A2(n725), .ZN(n728) );
  OR2_X1 U704 ( .A1(n578), .A2(n652), .ZN(n613) );
  XNOR2_X1 U705 ( .A(n604), .B(n602), .ZN(n717) );
  OR2_X1 U706 ( .A1(n598), .A2(n616), .ZN(n602) );
  OR2_X1 U707 ( .A1(n729), .A2(n730), .ZN(n604) );
  AND2_X1 U708 ( .A1(n731), .A2(n732), .ZN(n730) );
  AND2_X1 U709 ( .A1(n733), .A2(n734), .ZN(n729) );
  OR2_X1 U710 ( .A1(n732), .A2(n731), .ZN(n734) );
  XNOR2_X1 U711 ( .A(n596), .B(n594), .ZN(n716) );
  OR2_X1 U712 ( .A1(n640), .A2(n579), .ZN(n594) );
  OR2_X1 U713 ( .A1(n735), .A2(n736), .ZN(n596) );
  AND2_X1 U714 ( .A1(n715), .A2(n714), .ZN(n736) );
  AND2_X1 U715 ( .A1(n712), .A2(n737), .ZN(n735) );
  OR2_X1 U716 ( .A1(n714), .A2(n715), .ZN(n737) );
  OR2_X1 U717 ( .A1(n616), .A2(n640), .ZN(n715) );
  OR2_X1 U718 ( .A1(n738), .A2(n739), .ZN(n714) );
  AND2_X1 U719 ( .A1(n711), .A2(n710), .ZN(n739) );
  AND2_X1 U720 ( .A1(n708), .A2(n740), .ZN(n738) );
  OR2_X1 U721 ( .A1(n710), .A2(n711), .ZN(n740) );
  OR2_X1 U722 ( .A1(n652), .A2(n640), .ZN(n711) );
  OR2_X1 U723 ( .A1(n741), .A2(n742), .ZN(n710) );
  AND2_X1 U724 ( .A1(n707), .A2(n706), .ZN(n742) );
  AND2_X1 U725 ( .A1(n704), .A2(n743), .ZN(n741) );
  OR2_X1 U726 ( .A1(n706), .A2(n707), .ZN(n743) );
  OR2_X1 U727 ( .A1(n647), .A2(n640), .ZN(n707) );
  OR2_X1 U728 ( .A1(n744), .A2(n745), .ZN(n706) );
  AND2_X1 U729 ( .A1(n703), .A2(n702), .ZN(n745) );
  AND2_X1 U730 ( .A1(n700), .A2(n746), .ZN(n744) );
  OR2_X1 U731 ( .A1(n703), .A2(n702), .ZN(n746) );
  OR2_X1 U732 ( .A1(n747), .A2(n748), .ZN(n702) );
  AND2_X1 U733 ( .A1(n697), .A2(n693), .ZN(n748) );
  AND2_X1 U734 ( .A1(n749), .A2(n698), .ZN(n747) );
  OR2_X1 U735 ( .A1(n750), .A2(n751), .ZN(n698) );
  INV_X1 U736 ( .A(n752), .ZN(n751) );
  AND2_X1 U737 ( .A1(n753), .A2(n754), .ZN(n750) );
  OR2_X1 U738 ( .A1(n697), .A2(n693), .ZN(n749) );
  OR2_X1 U739 ( .A1(n694), .A2(n695), .ZN(n693) );
  OR2_X1 U740 ( .A1(n521), .A2(n640), .ZN(n695) );
  OR2_X1 U741 ( .A1(n598), .A2(n638), .ZN(n694) );
  OR2_X1 U742 ( .A1(n636), .A2(n640), .ZN(n697) );
  OR2_X1 U743 ( .A1(n642), .A2(n640), .ZN(n703) );
  XOR2_X1 U744 ( .A(n755), .B(n756), .Z(n640) );
  XNOR2_X1 U745 ( .A(n757), .B(c_5_), .ZN(n756) );
  XNOR2_X1 U746 ( .A(n758), .B(n759), .ZN(n700) );
  XNOR2_X1 U747 ( .A(n760), .B(n752), .ZN(n758) );
  XOR2_X1 U748 ( .A(n761), .B(n762), .Z(n704) );
  XOR2_X1 U749 ( .A(n763), .B(n764), .Z(n762) );
  XOR2_X1 U750 ( .A(n765), .B(n766), .Z(n708) );
  XOR2_X1 U751 ( .A(n767), .B(n768), .Z(n766) );
  XOR2_X1 U752 ( .A(n733), .B(n769), .Z(n712) );
  XOR2_X1 U753 ( .A(n732), .B(n731), .Z(n769) );
  OR2_X1 U754 ( .A1(n598), .A2(n652), .ZN(n731) );
  OR2_X1 U755 ( .A1(n770), .A2(n771), .ZN(n732) );
  AND2_X1 U756 ( .A1(n768), .A2(n767), .ZN(n771) );
  AND2_X1 U757 ( .A1(n765), .A2(n772), .ZN(n770) );
  OR2_X1 U758 ( .A1(n767), .A2(n768), .ZN(n772) );
  OR2_X1 U759 ( .A1(n598), .A2(n647), .ZN(n768) );
  OR2_X1 U760 ( .A1(n773), .A2(n774), .ZN(n767) );
  AND2_X1 U761 ( .A1(n764), .A2(n763), .ZN(n774) );
  AND2_X1 U762 ( .A1(n761), .A2(n775), .ZN(n773) );
  OR2_X1 U763 ( .A1(n763), .A2(n764), .ZN(n775) );
  OR2_X1 U764 ( .A1(n598), .A2(n642), .ZN(n764) );
  OR2_X1 U765 ( .A1(n776), .A2(n777), .ZN(n763) );
  AND2_X1 U766 ( .A1(n759), .A2(n752), .ZN(n777) );
  AND2_X1 U767 ( .A1(n778), .A2(n760), .ZN(n776) );
  OR2_X1 U768 ( .A1(n779), .A2(n780), .ZN(n760) );
  INV_X1 U769 ( .A(n781), .ZN(n780) );
  AND2_X1 U770 ( .A1(n782), .A2(n783), .ZN(n779) );
  OR2_X1 U771 ( .A1(n759), .A2(n752), .ZN(n778) );
  OR2_X1 U772 ( .A1(n753), .A2(n754), .ZN(n752) );
  OR2_X1 U773 ( .A1(n578), .A2(n638), .ZN(n754) );
  OR2_X1 U774 ( .A1(n521), .A2(n598), .ZN(n753) );
  OR2_X1 U775 ( .A1(n598), .A2(n636), .ZN(n759) );
  XNOR2_X1 U776 ( .A(n784), .B(n785), .ZN(n598) );
  XNOR2_X1 U777 ( .A(c_4_), .B(d_4_), .ZN(n784) );
  XNOR2_X1 U778 ( .A(n786), .B(n781), .ZN(n761) );
  XNOR2_X1 U779 ( .A(n787), .B(n788), .ZN(n786) );
  XOR2_X1 U780 ( .A(n789), .B(n790), .Z(n765) );
  XOR2_X1 U781 ( .A(n791), .B(n792), .Z(n790) );
  XNOR2_X1 U782 ( .A(n793), .B(n727), .ZN(n733) );
  XNOR2_X1 U783 ( .A(n794), .B(n795), .ZN(n727) );
  XNOR2_X1 U784 ( .A(n796), .B(n797), .ZN(n794) );
  XNOR2_X1 U785 ( .A(n725), .B(n726), .ZN(n793) );
  OR2_X1 U786 ( .A1(n578), .A2(n647), .ZN(n726) );
  OR2_X1 U787 ( .A1(n798), .A2(n799), .ZN(n725) );
  AND2_X1 U788 ( .A1(n792), .A2(n791), .ZN(n799) );
  AND2_X1 U789 ( .A1(n789), .A2(n800), .ZN(n798) );
  OR2_X1 U790 ( .A1(n791), .A2(n792), .ZN(n800) );
  OR2_X1 U791 ( .A1(n801), .A2(n802), .ZN(n792) );
  AND2_X1 U792 ( .A1(n781), .A2(n788), .ZN(n802) );
  AND2_X1 U793 ( .A1(n803), .A2(n787), .ZN(n801) );
  OR2_X1 U794 ( .A1(n804), .A2(n805), .ZN(n787) );
  INV_X1 U795 ( .A(n806), .ZN(n805) );
  AND2_X1 U796 ( .A1(n807), .A2(n808), .ZN(n804) );
  OR2_X1 U797 ( .A1(n788), .A2(n781), .ZN(n803) );
  OR2_X1 U798 ( .A1(n782), .A2(n783), .ZN(n781) );
  OR2_X1 U799 ( .A1(n809), .A2(n638), .ZN(n783) );
  OR2_X1 U800 ( .A1(n521), .A2(n578), .ZN(n782) );
  OR2_X1 U801 ( .A1(n578), .A2(n636), .ZN(n788) );
  OR2_X1 U802 ( .A1(n578), .A2(n642), .ZN(n791) );
  XNOR2_X1 U803 ( .A(n810), .B(n811), .ZN(n578) );
  XNOR2_X1 U804 ( .A(c_3_), .B(d_3_), .ZN(n810) );
  XNOR2_X1 U805 ( .A(n812), .B(n813), .ZN(n789) );
  XNOR2_X1 U806 ( .A(n814), .B(n806), .ZN(n812) );
  OR2_X1 U807 ( .A1(n516), .A2(n815), .ZN(n512) );
  OR2_X1 U808 ( .A1(n515), .A2(n513), .ZN(n815) );
  XNOR2_X1 U809 ( .A(n816), .B(n817), .ZN(n513) );
  OR2_X1 U810 ( .A1(n818), .A2(n579), .ZN(n816) );
  XOR2_X1 U811 ( .A(n819), .B(n820), .Z(n515) );
  XOR2_X1 U812 ( .A(n821), .B(n822), .Z(n820) );
  OR2_X1 U813 ( .A1(n823), .A2(n824), .ZN(n516) );
  AND2_X1 U814 ( .A1(n560), .A2(n559), .ZN(n824) );
  AND2_X1 U815 ( .A1(n557), .A2(n825), .ZN(n823) );
  OR2_X1 U816 ( .A1(n559), .A2(n560), .ZN(n825) );
  OR2_X1 U817 ( .A1(n809), .A2(n579), .ZN(n560) );
  OR2_X1 U818 ( .A1(n826), .A2(n827), .ZN(n559) );
  AND2_X1 U819 ( .A1(n571), .A2(n570), .ZN(n827) );
  AND2_X1 U820 ( .A1(n568), .A2(n828), .ZN(n826) );
  OR2_X1 U821 ( .A1(n570), .A2(n571), .ZN(n828) );
  OR2_X1 U822 ( .A1(n809), .A2(n616), .ZN(n571) );
  OR2_X1 U823 ( .A1(n829), .A2(n830), .ZN(n570) );
  AND2_X1 U824 ( .A1(n609), .A2(n608), .ZN(n830) );
  AND2_X1 U825 ( .A1(n607), .A2(n831), .ZN(n829) );
  OR2_X1 U826 ( .A1(n608), .A2(n609), .ZN(n831) );
  OR2_X1 U827 ( .A1(n832), .A2(n833), .ZN(n609) );
  AND2_X1 U828 ( .A1(n722), .A2(n721), .ZN(n833) );
  AND2_X1 U829 ( .A1(n720), .A2(n834), .ZN(n832) );
  OR2_X1 U830 ( .A1(n721), .A2(n722), .ZN(n834) );
  OR2_X1 U831 ( .A1(n835), .A2(n836), .ZN(n722) );
  AND2_X1 U832 ( .A1(n797), .A2(n796), .ZN(n836) );
  AND2_X1 U833 ( .A1(n795), .A2(n837), .ZN(n835) );
  OR2_X1 U834 ( .A1(n796), .A2(n797), .ZN(n837) );
  OR2_X1 U835 ( .A1(n809), .A2(n642), .ZN(n797) );
  OR2_X1 U836 ( .A1(n838), .A2(n839), .ZN(n796) );
  AND2_X1 U837 ( .A1(n813), .A2(n806), .ZN(n839) );
  AND2_X1 U838 ( .A1(n840), .A2(n814), .ZN(n838) );
  OR2_X1 U839 ( .A1(n841), .A2(n842), .ZN(n814) );
  AND2_X1 U840 ( .A1(n843), .A2(n844), .ZN(n841) );
  OR2_X1 U841 ( .A1(n806), .A2(n813), .ZN(n840) );
  OR2_X1 U842 ( .A1(n809), .A2(n636), .ZN(n813) );
  OR2_X1 U843 ( .A1(n807), .A2(n808), .ZN(n806) );
  OR2_X1 U844 ( .A1(n845), .A2(n638), .ZN(n808) );
  OR2_X1 U845 ( .A1(n809), .A2(n521), .ZN(n807) );
  XNOR2_X1 U846 ( .A(n846), .B(n847), .ZN(n795) );
  OR2_X1 U847 ( .A1(n842), .A2(n848), .ZN(n846) );
  INV_X1 U848 ( .A(n849), .ZN(n842) );
  OR2_X1 U849 ( .A1(n809), .A2(n647), .ZN(n721) );
  XOR2_X1 U850 ( .A(n850), .B(n851), .Z(n720) );
  XOR2_X1 U851 ( .A(n852), .B(n853), .Z(n850) );
  OR2_X1 U852 ( .A1(n809), .A2(n652), .ZN(n608) );
  XNOR2_X1 U853 ( .A(n854), .B(n855), .ZN(n809) );
  XNOR2_X1 U854 ( .A(c_2_), .B(d_2_), .ZN(n854) );
  XOR2_X1 U855 ( .A(n856), .B(n857), .Z(n607) );
  XOR2_X1 U856 ( .A(n858), .B(n859), .Z(n857) );
  XOR2_X1 U857 ( .A(n860), .B(n861), .Z(n568) );
  XOR2_X1 U858 ( .A(n862), .B(n863), .Z(n861) );
  XOR2_X1 U859 ( .A(n864), .B(n865), .Z(n557) );
  XOR2_X1 U860 ( .A(n866), .B(n867), .Z(n865) );
  OR2_X1 U861 ( .A1(n817), .A2(n579), .ZN(n539) );
  OR2_X1 U862 ( .A1(n868), .A2(n869), .ZN(n817) );
  AND2_X1 U863 ( .A1(n819), .A2(n821), .ZN(n869) );
  AND2_X1 U864 ( .A1(n870), .A2(n822), .ZN(n868) );
  OR2_X1 U865 ( .A1(n845), .A2(n579), .ZN(n822) );
  XNOR2_X1 U866 ( .A(n871), .B(n872), .ZN(n579) );
  XOR2_X1 U867 ( .A(b_0_), .B(a_0_), .Z(n872) );
  OR2_X1 U868 ( .A1(n873), .A2(n874), .ZN(n871) );
  AND2_X1 U869 ( .A1(n875), .A2(a_1_), .ZN(n874) );
  AND2_X1 U870 ( .A1(b_1_), .A2(n876), .ZN(n873) );
  OR2_X1 U871 ( .A1(n875), .A2(a_1_), .ZN(n876) );
  INV_X1 U872 ( .A(n877), .ZN(n875) );
  OR2_X1 U873 ( .A1(n821), .A2(n819), .ZN(n870) );
  OR2_X1 U874 ( .A1(n616), .A2(n818), .ZN(n819) );
  OR2_X1 U875 ( .A1(n878), .A2(n879), .ZN(n821) );
  AND2_X1 U876 ( .A1(n864), .A2(n866), .ZN(n879) );
  AND2_X1 U877 ( .A1(n880), .A2(n867), .ZN(n878) );
  OR2_X1 U878 ( .A1(n845), .A2(n616), .ZN(n867) );
  XNOR2_X1 U879 ( .A(n881), .B(n877), .ZN(n616) );
  OR2_X1 U880 ( .A1(n882), .A2(n883), .ZN(n877) );
  AND2_X1 U881 ( .A1(n884), .A2(n885), .ZN(n883) );
  AND2_X1 U882 ( .A1(n886), .A2(n887), .ZN(n882) );
  INV_X1 U883 ( .A(b_2_), .ZN(n887) );
  OR2_X1 U884 ( .A1(n885), .A2(n884), .ZN(n886) );
  INV_X1 U885 ( .A(a_2_), .ZN(n885) );
  XNOR2_X1 U886 ( .A(a_1_), .B(b_1_), .ZN(n881) );
  OR2_X1 U887 ( .A1(n866), .A2(n864), .ZN(n880) );
  OR2_X1 U888 ( .A1(n652), .A2(n818), .ZN(n864) );
  OR2_X1 U889 ( .A1(n888), .A2(n889), .ZN(n866) );
  AND2_X1 U890 ( .A1(n860), .A2(n862), .ZN(n889) );
  AND2_X1 U891 ( .A1(n890), .A2(n863), .ZN(n888) );
  OR2_X1 U892 ( .A1(n647), .A2(n818), .ZN(n863) );
  OR2_X1 U893 ( .A1(n862), .A2(n860), .ZN(n890) );
  OR2_X1 U894 ( .A1(n845), .A2(n652), .ZN(n860) );
  XNOR2_X1 U895 ( .A(n891), .B(n884), .ZN(n652) );
  OR2_X1 U896 ( .A1(n892), .A2(n893), .ZN(n884) );
  AND2_X1 U897 ( .A1(n894), .A2(n895), .ZN(n893) );
  AND2_X1 U898 ( .A1(n896), .A2(n897), .ZN(n892) );
  INV_X1 U899 ( .A(b_3_), .ZN(n897) );
  OR2_X1 U900 ( .A1(n895), .A2(n894), .ZN(n896) );
  INV_X1 U901 ( .A(a_3_), .ZN(n895) );
  XNOR2_X1 U902 ( .A(a_2_), .B(b_2_), .ZN(n891) );
  OR2_X1 U903 ( .A1(n898), .A2(n899), .ZN(n862) );
  AND2_X1 U904 ( .A1(n856), .A2(n858), .ZN(n899) );
  AND2_X1 U905 ( .A1(n900), .A2(n859), .ZN(n898) );
  OR2_X1 U906 ( .A1(n845), .A2(n647), .ZN(n859) );
  XNOR2_X1 U907 ( .A(n901), .B(n894), .ZN(n647) );
  OR2_X1 U908 ( .A1(n902), .A2(n903), .ZN(n894) );
  AND2_X1 U909 ( .A1(n904), .A2(n905), .ZN(n903) );
  AND2_X1 U910 ( .A1(n906), .A2(n907), .ZN(n902) );
  INV_X1 U911 ( .A(b_4_), .ZN(n907) );
  OR2_X1 U912 ( .A1(n905), .A2(n904), .ZN(n906) );
  INV_X1 U913 ( .A(a_4_), .ZN(n905) );
  XNOR2_X1 U914 ( .A(a_3_), .B(b_3_), .ZN(n901) );
  OR2_X1 U915 ( .A1(n858), .A2(n856), .ZN(n900) );
  OR2_X1 U916 ( .A1(n642), .A2(n818), .ZN(n856) );
  OR2_X1 U917 ( .A1(n908), .A2(n909), .ZN(n858) );
  AND2_X1 U918 ( .A1(n851), .A2(n853), .ZN(n909) );
  AND2_X1 U919 ( .A1(n852), .A2(n910), .ZN(n908) );
  OR2_X1 U920 ( .A1(n853), .A2(n851), .ZN(n910) );
  OR2_X1 U921 ( .A1(n636), .A2(n818), .ZN(n851) );
  OR2_X1 U922 ( .A1(n845), .A2(n642), .ZN(n853) );
  XNOR2_X1 U923 ( .A(n911), .B(n904), .ZN(n642) );
  OR2_X1 U924 ( .A1(n912), .A2(n913), .ZN(n904) );
  AND2_X1 U925 ( .A1(n914), .A2(n915), .ZN(n913) );
  AND2_X1 U926 ( .A1(n916), .A2(n917), .ZN(n912) );
  OR2_X1 U927 ( .A1(n914), .A2(n915), .ZN(n916) );
  INV_X1 U928 ( .A(a_5_), .ZN(n915) );
  INV_X1 U929 ( .A(n918), .ZN(n914) );
  XNOR2_X1 U930 ( .A(a_4_), .B(b_4_), .ZN(n911) );
  AND2_X1 U931 ( .A1(n849), .A2(n919), .ZN(n852) );
  OR2_X1 U932 ( .A1(n847), .A2(n848), .ZN(n919) );
  OR2_X1 U933 ( .A1(n521), .A2(n818), .ZN(n848) );
  OR2_X1 U934 ( .A1(n845), .A2(n636), .ZN(n847) );
  XNOR2_X1 U935 ( .A(n918), .B(n920), .ZN(n636) );
  XNOR2_X1 U936 ( .A(n917), .B(a_5_), .ZN(n920) );
  INV_X1 U937 ( .A(b_5_), .ZN(n917) );
  OR2_X1 U938 ( .A1(n921), .A2(n922), .ZN(n918) );
  AND2_X1 U939 ( .A1(n923), .A2(a_6_), .ZN(n922) );
  AND2_X1 U940 ( .A1(b_6_), .A2(n924), .ZN(n921) );
  OR2_X1 U941 ( .A1(n923), .A2(a_6_), .ZN(n924) );
  OR2_X1 U942 ( .A1(n843), .A2(n844), .ZN(n849) );
  OR2_X1 U943 ( .A1(n638), .A2(n818), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n925), .B(n926), .ZN(n818) );
  XOR2_X1 U945 ( .A(d_0_), .B(c_0_), .Z(n926) );
  OR2_X1 U946 ( .A1(n927), .A2(n928), .ZN(n925) );
  AND2_X1 U947 ( .A1(n929), .A2(c_1_), .ZN(n928) );
  AND2_X1 U948 ( .A1(d_1_), .A2(n930), .ZN(n927) );
  OR2_X1 U949 ( .A1(n929), .A2(c_1_), .ZN(n930) );
  INV_X1 U950 ( .A(n931), .ZN(n929) );
  OR2_X1 U951 ( .A1(n932), .A2(n923), .ZN(n638) );
  INV_X1 U952 ( .A(n933), .ZN(n932) );
  OR2_X1 U953 ( .A1(a_7_), .A2(b_7_), .ZN(n933) );
  OR2_X1 U954 ( .A1(n521), .A2(n845), .ZN(n843) );
  XNOR2_X1 U955 ( .A(n934), .B(n931), .ZN(n845) );
  OR2_X1 U956 ( .A1(n935), .A2(n936), .ZN(n931) );
  AND2_X1 U957 ( .A1(n855), .A2(n937), .ZN(n936) );
  AND2_X1 U958 ( .A1(n938), .A2(n939), .ZN(n935) );
  INV_X1 U959 ( .A(d_2_), .ZN(n939) );
  OR2_X1 U960 ( .A1(n937), .A2(n855), .ZN(n938) );
  OR2_X1 U961 ( .A1(n940), .A2(n941), .ZN(n855) );
  AND2_X1 U962 ( .A1(n811), .A2(n942), .ZN(n941) );
  AND2_X1 U963 ( .A1(n943), .A2(n944), .ZN(n940) );
  INV_X1 U964 ( .A(d_3_), .ZN(n944) );
  OR2_X1 U965 ( .A1(n811), .A2(n942), .ZN(n943) );
  INV_X1 U966 ( .A(c_3_), .ZN(n942) );
  OR2_X1 U967 ( .A1(n945), .A2(n946), .ZN(n811) );
  AND2_X1 U968 ( .A1(n785), .A2(n947), .ZN(n946) );
  AND2_X1 U969 ( .A1(n948), .A2(n949), .ZN(n945) );
  INV_X1 U970 ( .A(d_4_), .ZN(n949) );
  OR2_X1 U971 ( .A1(n785), .A2(n947), .ZN(n948) );
  INV_X1 U972 ( .A(c_4_), .ZN(n947) );
  OR2_X1 U973 ( .A1(n950), .A2(n951), .ZN(n785) );
  AND2_X1 U974 ( .A1(n755), .A2(n952), .ZN(n951) );
  AND2_X1 U975 ( .A1(n953), .A2(n757), .ZN(n950) );
  INV_X1 U976 ( .A(d_5_), .ZN(n757) );
  OR2_X1 U977 ( .A1(n755), .A2(n952), .ZN(n953) );
  INV_X1 U978 ( .A(c_5_), .ZN(n952) );
  INV_X1 U979 ( .A(n954), .ZN(n755) );
  OR2_X1 U980 ( .A1(n955), .A2(n956), .ZN(n954) );
  AND2_X1 U981 ( .A1(c_6_), .A2(n654), .ZN(n956) );
  AND2_X1 U982 ( .A1(d_6_), .A2(n957), .ZN(n955) );
  OR2_X1 U983 ( .A1(n654), .A2(c_6_), .ZN(n957) );
  AND2_X1 U984 ( .A1(c_7_), .A2(d_7_), .ZN(n654) );
  INV_X1 U985 ( .A(c_2_), .ZN(n937) );
  XNOR2_X1 U986 ( .A(c_1_), .B(d_1_), .ZN(n934) );
  XNOR2_X1 U987 ( .A(n923), .B(n958), .ZN(n521) );
  XOR2_X1 U988 ( .A(b_6_), .B(a_6_), .Z(n958) );
  AND2_X1 U989 ( .A1(a_7_), .A2(b_7_), .ZN(n923) );
endmodule

