module add_mul_combine_8_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, Result_mul_0_, 
        Result_mul_1_, Result_mul_2_, Result_mul_3_, Result_mul_4_, 
        Result_mul_5_, Result_mul_6_, Result_mul_7_, Result_mul_8_, 
        Result_mul_9_, Result_mul_10_, Result_mul_11_, Result_mul_12_, 
        Result_mul_13_, Result_mul_14_, Result_mul_15_, Result_add_0_, 
        Result_add_1_, Result_add_2_, Result_add_3_, Result_add_4_, 
        Result_add_5_, Result_add_6_, Result_add_7_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_,
         b_4_, b_5_, b_6_, b_7_;
  output Result_mul_0_, Result_mul_1_, Result_mul_2_, Result_mul_3_,
         Result_mul_4_, Result_mul_5_, Result_mul_6_, Result_mul_7_,
         Result_mul_8_, Result_mul_9_, Result_mul_10_, Result_mul_11_,
         Result_mul_12_, Result_mul_13_, Result_mul_14_, Result_mul_15_,
         Result_add_0_, Result_add_1_, Result_add_2_, Result_add_3_,
         Result_add_4_, Result_add_5_, Result_add_6_, Result_add_7_;
  wire   n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838;

  XNOR2_X1 U429 ( .A(n405), .B(n406), .ZN(Result_mul_9_) );
  XNOR2_X1 U430 ( .A(n407), .B(n408), .ZN(n406) );
  XOR2_X1 U431 ( .A(n409), .B(n410), .Z(Result_mul_8_) );
  XOR2_X1 U432 ( .A(n411), .B(n412), .Z(n409) );
  NOR2_X1 U433 ( .A1(n413), .A2(n414), .ZN(n412) );
  XOR2_X1 U434 ( .A(n415), .B(n416), .Z(Result_mul_7_) );
  NOR2_X1 U435 ( .A1(n417), .A2(n418), .ZN(Result_mul_6_) );
  NOR2_X1 U436 ( .A1(n419), .A2(n420), .ZN(n418) );
  AND2_X1 U437 ( .A1(n415), .A2(n416), .ZN(n419) );
  XNOR2_X1 U438 ( .A(n417), .B(n421), .ZN(Result_mul_5_) );
  NAND2_X1 U439 ( .A1(n422), .A2(n423), .ZN(n421) );
  NAND2_X1 U440 ( .A1(n424), .A2(n425), .ZN(n423) );
  NAND2_X1 U441 ( .A1(n426), .A2(n427), .ZN(n424) );
  XOR2_X1 U442 ( .A(n428), .B(n429), .Z(Result_mul_4_) );
  XOR2_X1 U443 ( .A(n430), .B(n431), .Z(Result_mul_3_) );
  AND2_X1 U444 ( .A1(n432), .A2(n433), .ZN(n431) );
  XOR2_X1 U445 ( .A(n434), .B(n435), .Z(Result_mul_2_) );
  AND2_X1 U446 ( .A1(n436), .A2(n437), .ZN(n435) );
  XOR2_X1 U447 ( .A(n438), .B(n439), .Z(Result_mul_1_) );
  AND2_X1 U448 ( .A1(n440), .A2(n441), .ZN(n439) );
  XOR2_X1 U449 ( .A(n442), .B(n443), .Z(Result_mul_14_) );
  NAND2_X1 U450 ( .A1(b_7_), .A2(a_6_), .ZN(n443) );
  XOR2_X1 U451 ( .A(n444), .B(n445), .Z(Result_mul_13_) );
  XNOR2_X1 U452 ( .A(n446), .B(n447), .ZN(n445) );
  NAND2_X1 U453 ( .A1(b_7_), .A2(a_5_), .ZN(n446) );
  XNOR2_X1 U454 ( .A(n448), .B(n449), .ZN(Result_mul_12_) );
  NAND2_X1 U455 ( .A1(n450), .A2(n451), .ZN(n448) );
  XOR2_X1 U456 ( .A(n452), .B(n453), .Z(Result_mul_11_) );
  XNOR2_X1 U457 ( .A(n454), .B(n455), .ZN(n453) );
  NAND2_X1 U458 ( .A1(b_7_), .A2(a_3_), .ZN(n455) );
  XOR2_X1 U459 ( .A(n456), .B(n457), .Z(Result_mul_10_) );
  XOR2_X1 U460 ( .A(n458), .B(n459), .Z(n457) );
  NAND3_X1 U461 ( .A1(n460), .A2(n441), .A3(n461), .ZN(Result_mul_0_) );
  OR2_X1 U462 ( .A1(n414), .A2(n462), .ZN(n461) );
  NAND4_X1 U463 ( .A1(n462), .A2(n463), .A3(n464), .A4(n465), .ZN(n441) );
  NAND2_X1 U464 ( .A1(n440), .A2(n438), .ZN(n460) );
  NAND2_X1 U465 ( .A1(n437), .A2(n466), .ZN(n438) );
  NAND2_X1 U466 ( .A1(n436), .A2(n434), .ZN(n466) );
  NAND2_X1 U467 ( .A1(n433), .A2(n467), .ZN(n434) );
  NAND2_X1 U468 ( .A1(n430), .A2(n432), .ZN(n467) );
  NAND2_X1 U469 ( .A1(n468), .A2(n469), .ZN(n432) );
  NAND2_X1 U470 ( .A1(n470), .A2(n471), .ZN(n469) );
  XNOR2_X1 U471 ( .A(n472), .B(n473), .ZN(n468) );
  NOR2_X1 U472 ( .A1(n429), .A2(n428), .ZN(n430) );
  AND3_X1 U473 ( .A1(n474), .A2(n422), .A3(n475), .ZN(n428) );
  NAND2_X1 U474 ( .A1(n417), .A2(n476), .ZN(n475) );
  AND3_X1 U475 ( .A1(n416), .A2(n415), .A3(n420), .ZN(n417) );
  XOR2_X1 U476 ( .A(n427), .B(n426), .Z(n420) );
  NAND2_X1 U477 ( .A1(n477), .A2(n478), .ZN(n415) );
  NAND3_X1 U478 ( .A1(b_7_), .A2(n479), .A3(a_0_), .ZN(n478) );
  OR2_X1 U479 ( .A1(n410), .A2(n411), .ZN(n479) );
  NAND2_X1 U480 ( .A1(n410), .A2(n411), .ZN(n477) );
  NAND2_X1 U481 ( .A1(n480), .A2(n481), .ZN(n411) );
  NAND2_X1 U482 ( .A1(n408), .A2(n482), .ZN(n481) );
  OR2_X1 U483 ( .A1(n407), .A2(n405), .ZN(n482) );
  NOR2_X1 U484 ( .A1(n483), .A2(n413), .ZN(n408) );
  NAND2_X1 U485 ( .A1(n405), .A2(n407), .ZN(n480) );
  NAND2_X1 U486 ( .A1(n484), .A2(n485), .ZN(n407) );
  NAND2_X1 U487 ( .A1(n459), .A2(n486), .ZN(n485) );
  NAND2_X1 U488 ( .A1(n458), .A2(n456), .ZN(n486) );
  NOR2_X1 U489 ( .A1(n413), .A2(n487), .ZN(n459) );
  OR2_X1 U490 ( .A1(n456), .A2(n458), .ZN(n484) );
  AND2_X1 U491 ( .A1(n488), .A2(n489), .ZN(n458) );
  NAND3_X1 U492 ( .A1(a_3_), .A2(n490), .A3(b_7_), .ZN(n489) );
  NAND2_X1 U493 ( .A1(n454), .A2(n452), .ZN(n490) );
  OR2_X1 U494 ( .A1(n452), .A2(n454), .ZN(n488) );
  AND2_X1 U495 ( .A1(n450), .A2(n491), .ZN(n454) );
  NAND2_X1 U496 ( .A1(n449), .A2(n451), .ZN(n491) );
  NAND2_X1 U497 ( .A1(n492), .A2(n493), .ZN(n451) );
  NAND2_X1 U498 ( .A1(b_7_), .A2(a_4_), .ZN(n493) );
  INV_X1 U499 ( .A(n494), .ZN(n492) );
  XNOR2_X1 U500 ( .A(n495), .B(n496), .ZN(n449) );
  NAND2_X1 U501 ( .A1(n497), .A2(n498), .ZN(n495) );
  NAND2_X1 U502 ( .A1(a_4_), .A2(n494), .ZN(n450) );
  NAND2_X1 U503 ( .A1(n499), .A2(n500), .ZN(n494) );
  NAND3_X1 U504 ( .A1(a_5_), .A2(n501), .A3(b_7_), .ZN(n500) );
  NAND2_X1 U505 ( .A1(n444), .A2(n447), .ZN(n501) );
  OR2_X1 U506 ( .A1(n447), .A2(n444), .ZN(n499) );
  XNOR2_X1 U507 ( .A(n502), .B(n503), .ZN(n444) );
  NOR2_X1 U508 ( .A1(n504), .A2(n505), .ZN(n503) );
  XNOR2_X1 U509 ( .A(n506), .B(n507), .ZN(n452) );
  XOR2_X1 U510 ( .A(n508), .B(n509), .Z(n506) );
  XNOR2_X1 U511 ( .A(n510), .B(n511), .ZN(n456) );
  XNOR2_X1 U512 ( .A(n512), .B(n513), .ZN(n510) );
  NAND2_X1 U513 ( .A1(b_6_), .A2(a_3_), .ZN(n512) );
  XNOR2_X1 U514 ( .A(n514), .B(n515), .ZN(n405) );
  XOR2_X1 U515 ( .A(n516), .B(n517), .Z(n515) );
  NAND2_X1 U516 ( .A1(a_2_), .A2(b_6_), .ZN(n517) );
  XOR2_X1 U517 ( .A(n518), .B(n519), .Z(n410) );
  XOR2_X1 U518 ( .A(n520), .B(n521), .Z(n518) );
  NOR2_X1 U519 ( .A1(n522), .A2(n483), .ZN(n521) );
  XOR2_X1 U520 ( .A(n523), .B(n524), .Z(n416) );
  XOR2_X1 U521 ( .A(n525), .B(n526), .Z(n523) );
  NOR2_X1 U522 ( .A1(n522), .A2(n414), .ZN(n526) );
  NAND3_X1 U523 ( .A1(n426), .A2(n427), .A3(n476), .ZN(n422) );
  INV_X1 U524 ( .A(n425), .ZN(n476) );
  NAND2_X1 U525 ( .A1(n474), .A2(n527), .ZN(n425) );
  OR2_X1 U526 ( .A1(n528), .A2(n529), .ZN(n527) );
  NAND2_X1 U527 ( .A1(n530), .A2(n531), .ZN(n427) );
  NAND3_X1 U528 ( .A1(b_6_), .A2(n532), .A3(a_0_), .ZN(n531) );
  OR2_X1 U529 ( .A1(n524), .A2(n525), .ZN(n532) );
  NAND2_X1 U530 ( .A1(n524), .A2(n525), .ZN(n530) );
  NAND2_X1 U531 ( .A1(n533), .A2(n534), .ZN(n525) );
  NAND3_X1 U532 ( .A1(b_6_), .A2(n535), .A3(a_1_), .ZN(n534) );
  OR2_X1 U533 ( .A1(n520), .A2(n519), .ZN(n535) );
  NAND2_X1 U534 ( .A1(n519), .A2(n520), .ZN(n533) );
  NAND2_X1 U535 ( .A1(n536), .A2(n537), .ZN(n520) );
  NAND3_X1 U536 ( .A1(b_6_), .A2(n538), .A3(a_2_), .ZN(n537) );
  OR2_X1 U537 ( .A1(n514), .A2(n516), .ZN(n538) );
  NAND2_X1 U538 ( .A1(n514), .A2(n516), .ZN(n536) );
  NAND2_X1 U539 ( .A1(n539), .A2(n540), .ZN(n516) );
  NAND3_X1 U540 ( .A1(a_3_), .A2(n541), .A3(b_6_), .ZN(n540) );
  OR2_X1 U541 ( .A1(n513), .A2(n511), .ZN(n541) );
  NAND2_X1 U542 ( .A1(n511), .A2(n513), .ZN(n539) );
  NAND2_X1 U543 ( .A1(n542), .A2(n543), .ZN(n513) );
  NAND2_X1 U544 ( .A1(n509), .A2(n544), .ZN(n543) );
  OR2_X1 U545 ( .A1(n508), .A2(n507), .ZN(n544) );
  NOR2_X1 U546 ( .A1(n522), .A2(n545), .ZN(n509) );
  NAND2_X1 U547 ( .A1(n507), .A2(n508), .ZN(n542) );
  NAND2_X1 U548 ( .A1(n497), .A2(n546), .ZN(n508) );
  NAND2_X1 U549 ( .A1(n496), .A2(n498), .ZN(n546) );
  NAND2_X1 U550 ( .A1(n547), .A2(n548), .ZN(n498) );
  INV_X1 U551 ( .A(n549), .ZN(n548) );
  NAND2_X1 U552 ( .A1(b_6_), .A2(a_5_), .ZN(n547) );
  XNOR2_X1 U553 ( .A(n550), .B(n551), .ZN(n496) );
  NOR2_X1 U554 ( .A1(n504), .A2(n552), .ZN(n551) );
  NAND2_X1 U555 ( .A1(n549), .A2(a_5_), .ZN(n497) );
  NOR2_X1 U556 ( .A1(n442), .A2(n550), .ZN(n549) );
  NAND2_X1 U557 ( .A1(b_6_), .A2(a_7_), .ZN(n442) );
  XOR2_X1 U558 ( .A(n553), .B(n554), .Z(n507) );
  XNOR2_X1 U559 ( .A(n555), .B(n556), .ZN(n554) );
  XNOR2_X1 U560 ( .A(n557), .B(n558), .ZN(n511) );
  NAND2_X1 U561 ( .A1(n559), .A2(n560), .ZN(n557) );
  XOR2_X1 U562 ( .A(n561), .B(n562), .Z(n514) );
  XOR2_X1 U563 ( .A(n563), .B(n564), .Z(n561) );
  NOR2_X1 U564 ( .A1(n505), .A2(n565), .ZN(n564) );
  XNOR2_X1 U565 ( .A(n566), .B(n567), .ZN(n519) );
  XOR2_X1 U566 ( .A(n568), .B(n569), .Z(n567) );
  NAND2_X1 U567 ( .A1(a_2_), .A2(b_5_), .ZN(n569) );
  XOR2_X1 U568 ( .A(n570), .B(n571), .Z(n524) );
  XNOR2_X1 U569 ( .A(n572), .B(n573), .ZN(n571) );
  NAND2_X1 U570 ( .A1(a_1_), .A2(b_5_), .ZN(n573) );
  XNOR2_X1 U571 ( .A(n574), .B(n575), .ZN(n426) );
  NAND2_X1 U572 ( .A1(n576), .A2(n577), .ZN(n574) );
  NAND2_X1 U573 ( .A1(n529), .A2(n528), .ZN(n474) );
  NAND2_X1 U574 ( .A1(n576), .A2(n578), .ZN(n528) );
  NAND2_X1 U575 ( .A1(n575), .A2(n577), .ZN(n578) );
  NAND2_X1 U576 ( .A1(n579), .A2(n580), .ZN(n577) );
  NAND2_X1 U577 ( .A1(a_0_), .A2(b_5_), .ZN(n580) );
  INV_X1 U578 ( .A(n581), .ZN(n579) );
  XNOR2_X1 U579 ( .A(n582), .B(n583), .ZN(n575) );
  NAND2_X1 U580 ( .A1(n584), .A2(n585), .ZN(n582) );
  NAND2_X1 U581 ( .A1(a_0_), .A2(n581), .ZN(n576) );
  NAND2_X1 U582 ( .A1(n586), .A2(n587), .ZN(n581) );
  NAND3_X1 U583 ( .A1(b_5_), .A2(n588), .A3(a_1_), .ZN(n587) );
  NAND2_X1 U584 ( .A1(n572), .A2(n570), .ZN(n588) );
  OR2_X1 U585 ( .A1(n570), .A2(n572), .ZN(n586) );
  AND2_X1 U586 ( .A1(n589), .A2(n590), .ZN(n572) );
  NAND3_X1 U587 ( .A1(b_5_), .A2(n591), .A3(a_2_), .ZN(n590) );
  OR2_X1 U588 ( .A1(n566), .A2(n568), .ZN(n591) );
  NAND2_X1 U589 ( .A1(n566), .A2(n568), .ZN(n589) );
  NAND2_X1 U590 ( .A1(n592), .A2(n593), .ZN(n568) );
  NAND3_X1 U591 ( .A1(b_5_), .A2(n594), .A3(a_3_), .ZN(n593) );
  OR2_X1 U592 ( .A1(n563), .A2(n562), .ZN(n594) );
  NAND2_X1 U593 ( .A1(n562), .A2(n563), .ZN(n592) );
  NAND2_X1 U594 ( .A1(n559), .A2(n595), .ZN(n563) );
  NAND2_X1 U595 ( .A1(n558), .A2(n560), .ZN(n595) );
  NAND2_X1 U596 ( .A1(n596), .A2(n597), .ZN(n560) );
  NAND2_X1 U597 ( .A1(b_5_), .A2(a_4_), .ZN(n597) );
  INV_X1 U598 ( .A(n598), .ZN(n596) );
  XNOR2_X1 U599 ( .A(n599), .B(n600), .ZN(n558) );
  NAND2_X1 U600 ( .A1(n601), .A2(n602), .ZN(n599) );
  NAND2_X1 U601 ( .A1(a_4_), .A2(n598), .ZN(n559) );
  NAND2_X1 U602 ( .A1(n603), .A2(n604), .ZN(n598) );
  NAND2_X1 U603 ( .A1(n555), .A2(n605), .ZN(n604) );
  NAND2_X1 U604 ( .A1(n606), .A2(n556), .ZN(n605) );
  INV_X1 U605 ( .A(n553), .ZN(n606) );
  NOR3_X1 U606 ( .A1(n552), .A2(n504), .A3(n550), .ZN(n555) );
  NAND2_X1 U607 ( .A1(b_5_), .A2(a_6_), .ZN(n550) );
  NAND2_X1 U608 ( .A1(n607), .A2(n553), .ZN(n603) );
  XOR2_X1 U609 ( .A(n608), .B(n609), .Z(n553) );
  XOR2_X1 U610 ( .A(n610), .B(n611), .Z(n562) );
  XNOR2_X1 U611 ( .A(n612), .B(n613), .ZN(n610) );
  XOR2_X1 U612 ( .A(n614), .B(n615), .Z(n566) );
  XNOR2_X1 U613 ( .A(n616), .B(n617), .ZN(n614) );
  XOR2_X1 U614 ( .A(n618), .B(n619), .Z(n570) );
  NAND2_X1 U615 ( .A1(n620), .A2(n621), .ZN(n618) );
  XOR2_X1 U616 ( .A(n622), .B(n623), .Z(n529) );
  XOR2_X1 U617 ( .A(n624), .B(n625), .Z(n622) );
  NOR2_X1 U618 ( .A1(n552), .A2(n414), .ZN(n625) );
  XNOR2_X1 U619 ( .A(n471), .B(n470), .ZN(n429) );
  NAND3_X1 U620 ( .A1(n470), .A2(n471), .A3(n626), .ZN(n433) );
  XNOR2_X1 U621 ( .A(n472), .B(n627), .ZN(n626) );
  NAND2_X1 U622 ( .A1(n628), .A2(n629), .ZN(n471) );
  NAND3_X1 U623 ( .A1(b_4_), .A2(n630), .A3(a_0_), .ZN(n629) );
  OR2_X1 U624 ( .A1(n624), .A2(n623), .ZN(n630) );
  NAND2_X1 U625 ( .A1(n623), .A2(n624), .ZN(n628) );
  NAND2_X1 U626 ( .A1(n584), .A2(n631), .ZN(n624) );
  NAND2_X1 U627 ( .A1(n583), .A2(n585), .ZN(n631) );
  NAND2_X1 U628 ( .A1(n632), .A2(n633), .ZN(n585) );
  NAND2_X1 U629 ( .A1(a_1_), .A2(b_4_), .ZN(n633) );
  INV_X1 U630 ( .A(n634), .ZN(n632) );
  XNOR2_X1 U631 ( .A(n635), .B(n636), .ZN(n583) );
  XNOR2_X1 U632 ( .A(n637), .B(n638), .ZN(n635) );
  NOR2_X1 U633 ( .A1(n639), .A2(n487), .ZN(n638) );
  NAND2_X1 U634 ( .A1(a_1_), .A2(n634), .ZN(n584) );
  NAND2_X1 U635 ( .A1(n620), .A2(n640), .ZN(n634) );
  NAND2_X1 U636 ( .A1(n619), .A2(n621), .ZN(n640) );
  NAND2_X1 U637 ( .A1(n641), .A2(n642), .ZN(n621) );
  NAND2_X1 U638 ( .A1(a_2_), .A2(b_4_), .ZN(n642) );
  XNOR2_X1 U639 ( .A(n643), .B(n644), .ZN(n619) );
  XNOR2_X1 U640 ( .A(n645), .B(n646), .ZN(n643) );
  OR2_X1 U641 ( .A1(n641), .A2(n487), .ZN(n620) );
  NAND2_X1 U642 ( .A1(n647), .A2(n648), .ZN(n641) );
  NAND2_X1 U643 ( .A1(n615), .A2(n649), .ZN(n648) );
  NAND2_X1 U644 ( .A1(n617), .A2(n616), .ZN(n649) );
  XOR2_X1 U645 ( .A(n650), .B(n651), .Z(n615) );
  NAND2_X1 U646 ( .A1(n652), .A2(n653), .ZN(n650) );
  OR2_X1 U647 ( .A1(n617), .A2(n616), .ZN(n647) );
  AND2_X1 U648 ( .A1(n654), .A2(n655), .ZN(n616) );
  NAND2_X1 U649 ( .A1(n656), .A2(n613), .ZN(n655) );
  NAND2_X1 U650 ( .A1(n611), .A2(n612), .ZN(n656) );
  OR2_X1 U651 ( .A1(n611), .A2(n612), .ZN(n654) );
  NAND2_X1 U652 ( .A1(n601), .A2(n657), .ZN(n612) );
  NAND2_X1 U653 ( .A1(n600), .A2(n602), .ZN(n657) );
  NAND2_X1 U654 ( .A1(n658), .A2(n659), .ZN(n602) );
  NAND2_X1 U655 ( .A1(b_4_), .A2(a_5_), .ZN(n659) );
  AND2_X1 U656 ( .A1(n660), .A2(n661), .ZN(n600) );
  NAND2_X1 U657 ( .A1(n662), .A2(n663), .ZN(n661) );
  NAND2_X1 U658 ( .A1(b_3_), .A2(a_6_), .ZN(n662) );
  OR2_X1 U659 ( .A1(n658), .A2(n664), .ZN(n601) );
  NAND2_X1 U660 ( .A1(n608), .A2(n609), .ZN(n658) );
  NOR2_X1 U661 ( .A1(n552), .A2(n665), .ZN(n609) );
  NOR2_X1 U662 ( .A1(n639), .A2(n504), .ZN(n608) );
  XNOR2_X1 U663 ( .A(n666), .B(n667), .ZN(n611) );
  NAND2_X1 U664 ( .A1(n668), .A2(n669), .ZN(n666) );
  NOR2_X1 U665 ( .A1(n565), .A2(n552), .ZN(n617) );
  XOR2_X1 U666 ( .A(n670), .B(n671), .Z(n623) );
  XNOR2_X1 U667 ( .A(n672), .B(n673), .ZN(n670) );
  XNOR2_X1 U668 ( .A(n674), .B(n675), .ZN(n470) );
  XOR2_X1 U669 ( .A(n676), .B(n677), .Z(n675) );
  NAND2_X1 U670 ( .A1(a_0_), .A2(b_3_), .ZN(n677) );
  NAND2_X1 U671 ( .A1(n678), .A2(n679), .ZN(n436) );
  NAND2_X1 U672 ( .A1(n473), .A2(n472), .ZN(n679) );
  XNOR2_X1 U673 ( .A(n464), .B(n465), .ZN(n678) );
  NAND3_X1 U674 ( .A1(n680), .A2(n472), .A3(n473), .ZN(n437) );
  INV_X1 U675 ( .A(n627), .ZN(n473) );
  XOR2_X1 U676 ( .A(n681), .B(n682), .Z(n627) );
  NAND2_X1 U677 ( .A1(n683), .A2(n684), .ZN(n681) );
  NAND2_X1 U678 ( .A1(n685), .A2(n686), .ZN(n472) );
  NAND3_X1 U679 ( .A1(b_3_), .A2(n687), .A3(a_0_), .ZN(n686) );
  NAND2_X1 U680 ( .A1(n674), .A2(n676), .ZN(n687) );
  OR2_X1 U681 ( .A1(n676), .A2(n674), .ZN(n685) );
  XNOR2_X1 U682 ( .A(n688), .B(n689), .ZN(n674) );
  XNOR2_X1 U683 ( .A(n690), .B(n691), .ZN(n688) );
  NAND2_X1 U684 ( .A1(a_1_), .A2(b_2_), .ZN(n690) );
  NAND2_X1 U685 ( .A1(n692), .A2(n693), .ZN(n676) );
  NAND2_X1 U686 ( .A1(n672), .A2(n694), .ZN(n693) );
  NAND2_X1 U687 ( .A1(n673), .A2(n671), .ZN(n694) );
  AND2_X1 U688 ( .A1(n695), .A2(n696), .ZN(n672) );
  NAND3_X1 U689 ( .A1(b_3_), .A2(n697), .A3(a_2_), .ZN(n696) );
  OR2_X1 U690 ( .A1(n636), .A2(n637), .ZN(n697) );
  NAND2_X1 U691 ( .A1(n637), .A2(n636), .ZN(n695) );
  XOR2_X1 U692 ( .A(n698), .B(n699), .Z(n636) );
  XNOR2_X1 U693 ( .A(n700), .B(n701), .ZN(n698) );
  NAND2_X1 U694 ( .A1(a_3_), .A2(b_2_), .ZN(n700) );
  AND2_X1 U695 ( .A1(n702), .A2(n703), .ZN(n637) );
  NAND2_X1 U696 ( .A1(n704), .A2(n705), .ZN(n703) );
  OR2_X1 U697 ( .A1(n644), .A2(n646), .ZN(n704) );
  NAND2_X1 U698 ( .A1(n644), .A2(n646), .ZN(n702) );
  AND2_X1 U699 ( .A1(n652), .A2(n706), .ZN(n646) );
  NAND2_X1 U700 ( .A1(n651), .A2(n653), .ZN(n706) );
  NAND2_X1 U701 ( .A1(n707), .A2(n708), .ZN(n653) );
  NAND2_X1 U702 ( .A1(a_4_), .A2(b_3_), .ZN(n708) );
  INV_X1 U703 ( .A(n709), .ZN(n707) );
  XNOR2_X1 U704 ( .A(n710), .B(n711), .ZN(n651) );
  NAND2_X1 U705 ( .A1(n712), .A2(n713), .ZN(n710) );
  NAND2_X1 U706 ( .A1(a_4_), .A2(n709), .ZN(n652) );
  NAND2_X1 U707 ( .A1(n668), .A2(n714), .ZN(n709) );
  NAND2_X1 U708 ( .A1(n667), .A2(n669), .ZN(n714) );
  NAND2_X1 U709 ( .A1(n660), .A2(n715), .ZN(n669) );
  NAND2_X1 U710 ( .A1(a_5_), .A2(b_3_), .ZN(n715) );
  INV_X1 U711 ( .A(n716), .ZN(n660) );
  XOR2_X1 U712 ( .A(n717), .B(n718), .Z(n667) );
  NAND2_X1 U713 ( .A1(n716), .A2(a_5_), .ZN(n668) );
  NOR3_X1 U714 ( .A1(n665), .A2(n663), .A3(n639), .ZN(n716) );
  NAND2_X1 U715 ( .A1(b_2_), .A2(a_7_), .ZN(n663) );
  XOR2_X1 U716 ( .A(n719), .B(n720), .Z(n644) );
  NAND2_X1 U717 ( .A1(n721), .A2(n722), .ZN(n719) );
  OR2_X1 U718 ( .A1(n671), .A2(n673), .ZN(n692) );
  NOR2_X1 U719 ( .A1(n483), .A2(n639), .ZN(n673) );
  XOR2_X1 U720 ( .A(n723), .B(n724), .Z(n671) );
  XOR2_X1 U721 ( .A(n725), .B(n726), .Z(n723) );
  XNOR2_X1 U722 ( .A(n465), .B(n727), .ZN(n680) );
  NAND2_X1 U723 ( .A1(n728), .A2(n729), .ZN(n440) );
  NAND2_X1 U724 ( .A1(n464), .A2(n465), .ZN(n729) );
  NAND2_X1 U725 ( .A1(n683), .A2(n730), .ZN(n465) );
  NAND2_X1 U726 ( .A1(n682), .A2(n684), .ZN(n730) );
  NAND2_X1 U727 ( .A1(n731), .A2(n732), .ZN(n684) );
  NAND2_X1 U728 ( .A1(a_0_), .A2(b_2_), .ZN(n732) );
  INV_X1 U729 ( .A(n733), .ZN(n731) );
  XOR2_X1 U730 ( .A(n734), .B(n735), .Z(n682) );
  NOR2_X1 U731 ( .A1(n487), .A2(n736), .ZN(n735) );
  XOR2_X1 U732 ( .A(n737), .B(n738), .Z(n734) );
  NAND2_X1 U733 ( .A1(a_0_), .A2(n733), .ZN(n683) );
  NAND2_X1 U734 ( .A1(n739), .A2(n740), .ZN(n733) );
  NAND3_X1 U735 ( .A1(b_2_), .A2(n741), .A3(a_1_), .ZN(n740) );
  OR2_X1 U736 ( .A1(n691), .A2(n689), .ZN(n741) );
  NAND2_X1 U737 ( .A1(n689), .A2(n691), .ZN(n739) );
  NAND2_X1 U738 ( .A1(n742), .A2(n743), .ZN(n691) );
  NAND2_X1 U739 ( .A1(n726), .A2(n744), .ZN(n743) );
  OR2_X1 U740 ( .A1(n725), .A2(n724), .ZN(n744) );
  NAND2_X1 U741 ( .A1(n724), .A2(n725), .ZN(n742) );
  NAND2_X1 U742 ( .A1(n745), .A2(n746), .ZN(n725) );
  NAND3_X1 U743 ( .A1(b_2_), .A2(n747), .A3(a_3_), .ZN(n746) );
  OR2_X1 U744 ( .A1(n701), .A2(n699), .ZN(n747) );
  NAND2_X1 U745 ( .A1(n699), .A2(n701), .ZN(n745) );
  NAND2_X1 U746 ( .A1(n721), .A2(n748), .ZN(n701) );
  NAND2_X1 U747 ( .A1(n720), .A2(n722), .ZN(n748) );
  NAND2_X1 U748 ( .A1(n749), .A2(n750), .ZN(n722) );
  NAND2_X1 U749 ( .A1(a_4_), .A2(b_2_), .ZN(n750) );
  INV_X1 U750 ( .A(n751), .ZN(n749) );
  XOR2_X1 U751 ( .A(n752), .B(n753), .Z(n720) );
  AND2_X1 U752 ( .A1(n754), .A2(n755), .ZN(n753) );
  NAND2_X1 U753 ( .A1(a_4_), .A2(n751), .ZN(n721) );
  NAND2_X1 U754 ( .A1(n712), .A2(n756), .ZN(n751) );
  NAND2_X1 U755 ( .A1(n711), .A2(n713), .ZN(n756) );
  NAND2_X1 U756 ( .A1(n757), .A2(n758), .ZN(n713) );
  NAND2_X1 U757 ( .A1(a_5_), .A2(b_2_), .ZN(n758) );
  AND2_X1 U758 ( .A1(n754), .A2(n759), .ZN(n711) );
  NAND2_X1 U759 ( .A1(n760), .A2(n761), .ZN(n759) );
  NAND2_X1 U760 ( .A1(b_0_), .A2(a_7_), .ZN(n761) );
  NAND2_X1 U761 ( .A1(b_1_), .A2(a_6_), .ZN(n760) );
  OR2_X1 U762 ( .A1(n757), .A2(n664), .ZN(n712) );
  NAND2_X1 U763 ( .A1(n717), .A2(n718), .ZN(n757) );
  NOR2_X1 U764 ( .A1(n665), .A2(n762), .ZN(n717) );
  XOR2_X1 U765 ( .A(n763), .B(n764), .Z(n699) );
  XOR2_X1 U766 ( .A(n765), .B(n766), .Z(n763) );
  XOR2_X1 U767 ( .A(n767), .B(n768), .Z(n724) );
  XNOR2_X1 U768 ( .A(n769), .B(n770), .ZN(n768) );
  NAND2_X1 U769 ( .A1(b_0_), .A2(a_4_), .ZN(n767) );
  XNOR2_X1 U770 ( .A(n771), .B(n772), .ZN(n689) );
  NAND2_X1 U771 ( .A1(n773), .A2(n774), .ZN(n771) );
  NAND2_X1 U772 ( .A1(n775), .A2(n776), .ZN(n774) );
  NAND2_X1 U773 ( .A1(a_2_), .A2(b_1_), .ZN(n775) );
  INV_X1 U774 ( .A(n727), .ZN(n464) );
  XNOR2_X1 U775 ( .A(n777), .B(n778), .ZN(n727) );
  NOR2_X1 U776 ( .A1(n779), .A2(n780), .ZN(n778) );
  NOR2_X1 U777 ( .A1(n781), .A2(n782), .ZN(n779) );
  NOR2_X1 U778 ( .A1(n783), .A2(n414), .ZN(n782) );
  XOR2_X1 U779 ( .A(n463), .B(n462), .Z(n728) );
  NOR2_X1 U780 ( .A1(n780), .A2(n784), .ZN(n462) );
  AND2_X1 U781 ( .A1(n785), .A2(n777), .ZN(n784) );
  NAND2_X1 U782 ( .A1(n786), .A2(n787), .ZN(n777) );
  NAND3_X1 U783 ( .A1(a_2_), .A2(n788), .A3(b_0_), .ZN(n787) );
  OR2_X1 U784 ( .A1(n738), .A2(n737), .ZN(n788) );
  NAND2_X1 U785 ( .A1(n737), .A2(n738), .ZN(n786) );
  NAND2_X1 U786 ( .A1(n773), .A2(n789), .ZN(n738) );
  NAND2_X1 U787 ( .A1(n790), .A2(n772), .ZN(n789) );
  NAND2_X1 U788 ( .A1(n791), .A2(n792), .ZN(n772) );
  NAND3_X1 U789 ( .A1(a_4_), .A2(n793), .A3(b_0_), .ZN(n792) );
  NAND2_X1 U790 ( .A1(n769), .A2(n770), .ZN(n793) );
  OR2_X1 U791 ( .A1(n770), .A2(n769), .ZN(n791) );
  AND2_X1 U792 ( .A1(n794), .A2(n795), .ZN(n769) );
  NAND2_X1 U793 ( .A1(n764), .A2(n796), .ZN(n795) );
  OR2_X1 U794 ( .A1(n766), .A2(n765), .ZN(n796) );
  NOR2_X1 U795 ( .A1(n736), .A2(n664), .ZN(n764) );
  NAND2_X1 U796 ( .A1(n765), .A2(n766), .ZN(n794) );
  NAND2_X1 U797 ( .A1(n797), .A2(n754), .ZN(n766) );
  NAND2_X1 U798 ( .A1(n755), .A2(n718), .ZN(n754) );
  NOR2_X1 U799 ( .A1(n783), .A2(n504), .ZN(n718) );
  NAND2_X1 U800 ( .A1(n752), .A2(n755), .ZN(n797) );
  NOR2_X1 U801 ( .A1(n736), .A2(n665), .ZN(n755) );
  NOR2_X1 U802 ( .A1(n783), .A2(n664), .ZN(n752) );
  NOR2_X1 U803 ( .A1(n545), .A2(n783), .ZN(n765) );
  NAND2_X1 U804 ( .A1(a_3_), .A2(b_1_), .ZN(n770) );
  NAND2_X1 U805 ( .A1(n776), .A2(n487), .ZN(n790) );
  OR3_X1 U806 ( .A1(n487), .A2(n783), .A3(n776), .ZN(n773) );
  NAND2_X1 U807 ( .A1(b_0_), .A2(a_3_), .ZN(n776) );
  NAND2_X1 U808 ( .A1(n798), .A2(n414), .ZN(n785) );
  NOR3_X1 U809 ( .A1(n414), .A2(n783), .A3(n798), .ZN(n780) );
  INV_X1 U810 ( .A(n781), .ZN(n798) );
  NOR2_X1 U811 ( .A1(n736), .A2(n483), .ZN(n781) );
  XNOR2_X1 U812 ( .A(n413), .B(a_7_), .ZN(Result_add_7_) );
  NAND3_X1 U813 ( .A1(n799), .A2(n800), .A3(n447), .ZN(Result_add_6_) );
  NAND2_X1 U814 ( .A1(Result_mul_15_), .A2(n502), .ZN(n447) );
  NAND2_X1 U815 ( .A1(n801), .A2(n522), .ZN(n800) );
  XNOR2_X1 U816 ( .A(a_6_), .B(n802), .ZN(n801) );
  NAND3_X1 U817 ( .A1(n802), .A2(n665), .A3(b_6_), .ZN(n799) );
  INV_X1 U818 ( .A(Result_mul_15_), .ZN(n802) );
  NAND3_X1 U819 ( .A1(n803), .A2(n804), .A3(n805), .ZN(Result_add_5_) );
  NAND2_X1 U820 ( .A1(n607), .A2(n806), .ZN(n805) );
  NAND3_X1 U821 ( .A1(n807), .A2(n664), .A3(b_5_), .ZN(n804) );
  NAND2_X1 U822 ( .A1(n808), .A2(n505), .ZN(n803) );
  XNOR2_X1 U823 ( .A(a_5_), .B(n807), .ZN(n808) );
  XNOR2_X1 U824 ( .A(n809), .B(n810), .ZN(Result_add_4_) );
  NAND2_X1 U825 ( .A1(n613), .A2(n811), .ZN(n809) );
  NAND3_X1 U826 ( .A1(n812), .A2(n813), .A3(n814), .ZN(Result_add_3_) );
  NAND2_X1 U827 ( .A1(n645), .A2(n815), .ZN(n814) );
  OR3_X1 U828 ( .A1(n815), .A2(a_3_), .A3(n639), .ZN(n813) );
  NAND2_X1 U829 ( .A1(n816), .A2(n639), .ZN(n812) );
  XNOR2_X1 U830 ( .A(n815), .B(n565), .ZN(n816) );
  XNOR2_X1 U831 ( .A(n817), .B(n818), .ZN(Result_add_2_) );
  NOR2_X1 U832 ( .A1(n819), .A2(n726), .ZN(n818) );
  NAND2_X1 U833 ( .A1(n820), .A2(n821), .ZN(Result_add_1_) );
  NAND2_X1 U834 ( .A1(n822), .A2(n823), .ZN(n821) );
  OR2_X1 U835 ( .A1(n737), .A2(n824), .ZN(n822) );
  NAND2_X1 U836 ( .A1(n825), .A2(n826), .ZN(n820) );
  XNOR2_X1 U837 ( .A(n783), .B(a_1_), .ZN(n825) );
  XOR2_X1 U838 ( .A(n827), .B(n828), .Z(Result_add_0_) );
  NOR2_X1 U839 ( .A1(n829), .A2(n463), .ZN(n828) );
  NOR2_X1 U840 ( .A1(n414), .A2(n736), .ZN(n463) );
  INV_X1 U841 ( .A(b_0_), .ZN(n736) );
  INV_X1 U842 ( .A(a_0_), .ZN(n414) );
  NOR2_X1 U843 ( .A1(b_0_), .A2(a_0_), .ZN(n829) );
  NOR2_X1 U844 ( .A1(n824), .A2(n830), .ZN(n827) );
  NOR2_X1 U845 ( .A1(n737), .A2(n823), .ZN(n830) );
  INV_X1 U846 ( .A(n826), .ZN(n823) );
  NOR2_X1 U847 ( .A1(n726), .A2(n831), .ZN(n826) );
  NOR2_X1 U848 ( .A1(n819), .A2(n817), .ZN(n831) );
  AND2_X1 U849 ( .A1(n705), .A2(n832), .ZN(n817) );
  NAND2_X1 U850 ( .A1(n833), .A2(n815), .ZN(n832) );
  NAND2_X1 U851 ( .A1(n613), .A2(n834), .ZN(n815) );
  NAND2_X1 U852 ( .A1(n811), .A2(n810), .ZN(n834) );
  NAND2_X1 U853 ( .A1(n556), .A2(n835), .ZN(n810) );
  NAND2_X1 U854 ( .A1(n836), .A2(n806), .ZN(n835) );
  INV_X1 U855 ( .A(n807), .ZN(n806) );
  NOR2_X1 U856 ( .A1(n502), .A2(n837), .ZN(n807) );
  AND2_X1 U857 ( .A1(Result_mul_15_), .A2(n838), .ZN(n837) );
  NAND2_X1 U858 ( .A1(n522), .A2(n665), .ZN(n838) );
  NOR2_X1 U859 ( .A1(n413), .A2(n504), .ZN(Result_mul_15_) );
  INV_X1 U860 ( .A(a_7_), .ZN(n504) );
  INV_X1 U861 ( .A(b_7_), .ZN(n413) );
  NOR2_X1 U862 ( .A1(n522), .A2(n665), .ZN(n502) );
  INV_X1 U863 ( .A(a_6_), .ZN(n665) );
  INV_X1 U864 ( .A(b_6_), .ZN(n522) );
  NAND2_X1 U865 ( .A1(n505), .A2(n664), .ZN(n836) );
  INV_X1 U866 ( .A(n607), .ZN(n556) );
  NOR2_X1 U867 ( .A1(n505), .A2(n664), .ZN(n607) );
  INV_X1 U868 ( .A(a_5_), .ZN(n664) );
  INV_X1 U869 ( .A(b_5_), .ZN(n505) );
  NAND2_X1 U870 ( .A1(n552), .A2(n545), .ZN(n811) );
  INV_X1 U871 ( .A(a_4_), .ZN(n545) );
  INV_X1 U872 ( .A(b_4_), .ZN(n552) );
  NAND2_X1 U873 ( .A1(b_4_), .A2(a_4_), .ZN(n613) );
  NAND2_X1 U874 ( .A1(n639), .A2(n565), .ZN(n833) );
  INV_X1 U875 ( .A(n645), .ZN(n705) );
  NOR2_X1 U876 ( .A1(n565), .A2(n639), .ZN(n645) );
  INV_X1 U877 ( .A(b_3_), .ZN(n639) );
  INV_X1 U878 ( .A(a_3_), .ZN(n565) );
  NOR2_X1 U879 ( .A1(b_2_), .A2(a_2_), .ZN(n819) );
  NOR2_X1 U880 ( .A1(n487), .A2(n762), .ZN(n726) );
  INV_X1 U881 ( .A(b_2_), .ZN(n762) );
  INV_X1 U882 ( .A(a_2_), .ZN(n487) );
  NOR2_X1 U883 ( .A1(n483), .A2(n783), .ZN(n737) );
  INV_X1 U884 ( .A(b_1_), .ZN(n783) );
  INV_X1 U885 ( .A(a_1_), .ZN(n483) );
  NOR2_X1 U886 ( .A1(b_1_), .A2(a_1_), .ZN(n824) );
endmodule

