module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n236_, new_n976_, new_n238_, new_n479_, new_n1009_, new_n1105_, new_n955_, new_n608_, new_n847_, new_n250_, new_n888_, new_n501_, new_n288_, new_n1157_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1048_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n1025_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n1057_, new_n670_, new_n456_, new_n691_, new_n1024_, new_n1125_, new_n170_, new_n246_, new_n682_, new_n1075_, new_n812_, new_n911_, new_n679_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n1131_, new_n1120_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n188_, new_n695_, new_n240_, new_n660_, new_n413_, new_n1060_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n1119_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n1045_, new_n1132_, new_n500_, new_n898_, new_n786_, new_n799_, new_n946_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n1108_, new_n862_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n959_, new_n990_, new_n774_, new_n157_, new_n716_, new_n153_, new_n701_, new_n792_, new_n1058_, new_n953_, new_n257_, new_n481_, new_n212_, new_n1073_, new_n1110_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n1050_, new_n903_, new_n164_, new_n230_, new_n1151_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n1082_, new_n849_, new_n1018_, new_n606_, new_n1037_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n1054_, new_n1083_, new_n167_, new_n385_, new_n1049_, new_n829_, new_n478_, new_n694_, new_n461_, new_n710_, new_n971_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n150_, new_n683_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n966_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n1031_, new_n961_, new_n530_, new_n890_, new_n318_, new_n1006_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n1005_, new_n999_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n956_, new_n158_, new_n763_, new_n960_, new_n1138_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n970_, new_n995_, new_n1035_, new_n271_, new_n674_, new_n274_, new_n991_, new_n1044_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n1051_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n1046_, new_n650_, new_n708_, new_n750_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n734_, new_n925_, new_n1062_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n256_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n1121_, new_n820_, new_n1127_, new_n771_, new_n388_, new_n979_, new_n1028_, new_n508_, new_n714_, new_n194_, new_n483_, new_n1004_, new_n1152_, new_n394_, new_n299_, new_n1007_, new_n142_, new_n935_, new_n139_, new_n882_, new_n657_, new_n1145_, new_n929_, new_n652_, new_n314_, new_n582_, new_n986_, new_n1020_, new_n363_, new_n1150_, new_n1113_, new_n165_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n917_, new_n1041_, new_n426_, new_n1036_, new_n235_, new_n1133_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n1026_, new_n207_, new_n267_, new_n1106_, new_n473_, new_n140_, new_n1147_, new_n790_, new_n1081_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n969_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n996_, new_n621_, new_n846_, new_n915_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n874_, new_n943_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n198_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n208_, new_n632_, new_n1039_, new_n671_, new_n965_, new_n528_, new_n952_, new_n179_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n397_, new_n729_, new_n1111_, new_n975_, new_n399_, new_n596_, new_n945_, new_n805_, new_n1115_, new_n559_, new_n948_, new_n762_, new_n1055_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n1085_, new_n1154_, new_n295_, new_n359_, new_n794_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n1090_, new_n457_, new_n161_, new_n553_, new_n1114_, new_n1084_, new_n1061_, new_n668_, new_n333_, new_n1128_, new_n1002_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n1032_, new_n276_, new_n688_, new_n155_, new_n384_, new_n900_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n202_, new_n1034_, new_n296_, new_n661_, new_n308_, new_n1000_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n1070_, new_n176_, new_n1109_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n938_, new_n809_, new_n1142_, new_n654_, new_n713_, new_n880_, new_n1102_, new_n604_, new_n227_, new_n1104_, new_n690_, new_n416_, new_n222_, new_n1043_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n1136_, new_n693_, new_n505_, new_n619_, new_n471_, new_n967_, new_n268_, new_n374_, new_n577_, new_n1135_, new_n376_, new_n380_, new_n1079_, new_n747_, new_n138_, new_n749_, new_n861_, new_n1095_, new_n310_, new_n144_, new_n275_, new_n998_, new_n1056_, new_n352_, new_n1094_, new_n931_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n562_, new_n578_, new_n918_, new_n940_, new_n810_, new_n808_, new_n1064_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n800_, new_n379_, new_n1012_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n963_, new_n270_, new_n570_, new_n598_, new_n893_, new_n1063_, new_n824_, new_n143_, new_n520_, new_n1001_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n149_, new_n557_, new_n260_, new_n936_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1016_, new_n1074_, new_n748_, new_n1144_, new_n1137_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n1141_, new_n807_, new_n736_, new_n879_, new_n151_, new_n513_, new_n592_, new_n726_, new_n1123_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n1080_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n1126_, new_n1155_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n302_, new_n191_, new_n755_, new_n225_, new_n1040_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n533_, new_n1088_, new_n795_, new_n1146_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n1122_, new_n977_, new_n1139_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n972_, new_n1067_, new_n891_, new_n631_, new_n453_, new_n516_, new_n163_, new_n997_, new_n519_, new_n563_, new_n148_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n1076_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n1038_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n190_, new_n597_, new_n1093_, new_n1092_, new_n408_, new_n470_, new_n213_, new_n1072_, new_n769_, new_n1097_, new_n1069_, new_n651_, new_n433_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n992_, new_n1098_, new_n265_, new_n732_, new_n687_, new_n370_, new_n1029_, new_n689_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n1052_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n989_, new_n1117_, new_n711_, new_n1156_, new_n644_, new_n731_, new_n599_, new_n836_, new_n1116_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n327_, new_n681_, new_n1087_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n319_, new_n1008_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n957_, new_n754_, new_n1047_, new_n787_, new_n653_, new_n1134_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n330_, new_n727_, new_n375_, new_n962_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n357_, new_n320_, new_n780_, new_n984_, new_n245_, new_n643_, new_n474_, new_n1129_, new_n467_, new_n1013_, new_n404_, new_n1077_, new_n193_, new_n490_, new_n560_, new_n1100_, new_n1027_, new_n358_, new_n877_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n1011_, new_n425_, new_n175_, new_n226_, new_n896_, new_n802_, new_n697_, new_n1099_, new_n185_, new_n1023_, new_n709_, new_n373_, new_n866_, new_n171_, new_n540_, new_n1149_, new_n1066_, new_n434_, new_n200_, new_n947_, new_n994_, new_n982_, new_n422_, new_n964_, new_n1078_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n551_, new_n168_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n1140_, new_n521_, new_n1042_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n1089_, new_n181_, new_n573_, new_n765_, new_n405_, new_n1103_;

not g0000 ( new_n138_, keyIn_0_10 );
not g0001 ( new_n139_, keyIn_0_5 );
not g0002 ( new_n140_, N69 );
nand g0003 ( new_n141_, new_n140_, N65 );
not g0004 ( new_n142_, N65 );
nand g0005 ( new_n143_, new_n142_, N69 );
nand g0006 ( new_n144_, new_n141_, new_n143_ );
nand g0007 ( new_n145_, new_n144_, new_n139_ );
not g0008 ( new_n146_, new_n144_ );
nand g0009 ( new_n147_, new_n146_, keyIn_0_5 );
nand g0010 ( new_n148_, new_n147_, new_n145_ );
not g0011 ( new_n149_, N73 );
nor g0012 ( new_n150_, new_n149_, N77 );
not g0013 ( new_n151_, N77 );
nor g0014 ( new_n152_, new_n151_, N73 );
nor g0015 ( new_n153_, new_n150_, new_n152_ );
nor g0016 ( new_n154_, new_n148_, new_n153_ );
not g0017 ( new_n155_, new_n145_ );
nor g0018 ( new_n156_, new_n144_, new_n139_ );
nor g0019 ( new_n157_, new_n155_, new_n156_ );
not g0020 ( new_n158_, new_n153_ );
nor g0021 ( new_n159_, new_n157_, new_n158_ );
nor g0022 ( new_n160_, new_n159_, new_n154_ );
nor g0023 ( new_n161_, new_n160_, new_n138_ );
nand g0024 ( new_n162_, new_n157_, new_n158_ );
nand g0025 ( new_n163_, new_n148_, new_n153_ );
nand g0026 ( new_n164_, new_n162_, new_n163_ );
nor g0027 ( new_n165_, new_n164_, keyIn_0_10 );
nor g0028 ( new_n166_, new_n161_, new_n165_ );
not g0029 ( new_n167_, N81 );
nor g0030 ( new_n168_, new_n167_, N85 );
not g0031 ( new_n169_, N85 );
nor g0032 ( new_n170_, new_n169_, N81 );
nor g0033 ( new_n171_, new_n168_, new_n170_ );
not g0034 ( new_n172_, N89 );
nor g0035 ( new_n173_, new_n172_, N93 );
not g0036 ( new_n174_, N93 );
nor g0037 ( new_n175_, new_n174_, N89 );
nor g0038 ( new_n176_, new_n173_, new_n175_ );
not g0039 ( new_n177_, new_n176_ );
nor g0040 ( new_n178_, new_n177_, new_n171_ );
not g0041 ( new_n179_, new_n178_ );
nand g0042 ( new_n180_, new_n177_, new_n171_ );
nand g0043 ( new_n181_, new_n179_, new_n180_ );
nand g0044 ( new_n182_, new_n181_, keyIn_0_11 );
not g0045 ( new_n183_, new_n182_ );
nor g0046 ( new_n184_, new_n181_, keyIn_0_11 );
nor g0047 ( new_n185_, new_n183_, new_n184_ );
nor g0048 ( new_n186_, new_n166_, new_n185_ );
nand g0049 ( new_n187_, new_n164_, keyIn_0_10 );
nand g0050 ( new_n188_, new_n160_, new_n138_ );
nand g0051 ( new_n189_, new_n188_, new_n187_ );
not g0052 ( new_n190_, keyIn_0_11 );
not g0053 ( new_n191_, new_n181_ );
nand g0054 ( new_n192_, new_n191_, new_n190_ );
nand g0055 ( new_n193_, new_n192_, new_n182_ );
nor g0056 ( new_n194_, new_n189_, new_n193_ );
nor g0057 ( new_n195_, new_n186_, new_n194_ );
nor g0058 ( new_n196_, new_n195_, keyIn_0_26 );
not g0059 ( new_n197_, keyIn_0_26 );
nand g0060 ( new_n198_, new_n189_, new_n193_ );
nand g0061 ( new_n199_, new_n166_, new_n185_ );
nand g0062 ( new_n200_, new_n199_, new_n198_ );
nor g0063 ( new_n201_, new_n200_, new_n197_ );
nor g0064 ( new_n202_, new_n196_, new_n201_ );
nand g0065 ( new_n203_, N129, N137 );
not g0066 ( new_n204_, new_n203_ );
nor g0067 ( new_n205_, new_n202_, new_n204_ );
nand g0068 ( new_n206_, new_n200_, new_n197_ );
nand g0069 ( new_n207_, new_n195_, keyIn_0_26 );
nand g0070 ( new_n208_, new_n207_, new_n206_ );
nor g0071 ( new_n209_, new_n208_, new_n203_ );
nor g0072 ( new_n210_, new_n205_, new_n209_ );
nor g0073 ( new_n211_, new_n210_, keyIn_0_30 );
not g0074 ( new_n212_, keyIn_0_30 );
nand g0075 ( new_n213_, new_n208_, new_n203_ );
nand g0076 ( new_n214_, new_n202_, new_n204_ );
nand g0077 ( new_n215_, new_n214_, new_n213_ );
nor g0078 ( new_n216_, new_n215_, new_n212_ );
nor g0079 ( new_n217_, new_n211_, new_n216_ );
not g0080 ( new_n218_, keyIn_0_14 );
not g0081 ( new_n219_, N1 );
nor g0082 ( new_n220_, new_n219_, N17 );
not g0083 ( new_n221_, N17 );
nor g0084 ( new_n222_, new_n221_, N1 );
nor g0085 ( new_n223_, new_n220_, new_n222_ );
not g0086 ( new_n224_, N33 );
nor g0087 ( new_n225_, new_n224_, N49 );
not g0088 ( new_n226_, N49 );
nor g0089 ( new_n227_, new_n226_, N33 );
nor g0090 ( new_n228_, new_n225_, new_n227_ );
not g0091 ( new_n229_, new_n228_ );
nor g0092 ( new_n230_, new_n229_, new_n223_ );
nand g0093 ( new_n231_, new_n229_, new_n223_ );
not g0094 ( new_n232_, new_n231_ );
nor g0095 ( new_n233_, new_n232_, new_n230_ );
not g0096 ( new_n234_, new_n233_ );
nand g0097 ( new_n235_, new_n234_, new_n218_ );
not g0098 ( new_n236_, new_n235_ );
nor g0099 ( new_n237_, new_n234_, new_n218_ );
nor g0100 ( new_n238_, new_n236_, new_n237_ );
not g0101 ( new_n239_, new_n238_ );
nand g0102 ( new_n240_, new_n217_, new_n239_ );
nand g0103 ( new_n241_, new_n215_, new_n212_ );
nand g0104 ( new_n242_, new_n210_, keyIn_0_30 );
nand g0105 ( new_n243_, new_n242_, new_n241_ );
nand g0106 ( new_n244_, new_n243_, new_n238_ );
nand g0107 ( new_n245_, new_n240_, new_n244_ );
nand g0108 ( new_n246_, new_n245_, keyIn_0_38 );
not g0109 ( new_n247_, keyIn_0_38 );
nor g0110 ( new_n248_, new_n243_, new_n238_ );
nor g0111 ( new_n249_, new_n217_, new_n239_ );
nor g0112 ( new_n250_, new_n249_, new_n248_ );
nand g0113 ( new_n251_, new_n250_, new_n247_ );
nand g0114 ( new_n252_, new_n251_, new_n246_ );
not g0115 ( new_n253_, keyIn_0_56 );
not g0116 ( new_n254_, keyIn_0_54 );
not g0117 ( new_n255_, keyIn_0_47 );
not g0118 ( new_n256_, keyIn_0_39 );
not g0119 ( new_n257_, keyIn_0_31 );
not g0120 ( new_n258_, keyIn_0_27 );
not g0121 ( new_n259_, keyIn_0_12 );
not g0122 ( new_n260_, N97 );
nor g0123 ( new_n261_, new_n260_, N101 );
not g0124 ( new_n262_, N101 );
nor g0125 ( new_n263_, new_n262_, N97 );
nor g0126 ( new_n264_, new_n261_, new_n263_ );
not g0127 ( new_n265_, N105 );
nor g0128 ( new_n266_, new_n265_, N109 );
not g0129 ( new_n267_, N109 );
nor g0130 ( new_n268_, new_n267_, N105 );
nor g0131 ( new_n269_, new_n266_, new_n268_ );
not g0132 ( new_n270_, new_n269_ );
nor g0133 ( new_n271_, new_n270_, new_n264_ );
not g0134 ( new_n272_, new_n271_ );
nand g0135 ( new_n273_, new_n270_, new_n264_ );
nand g0136 ( new_n274_, new_n272_, new_n273_ );
nand g0137 ( new_n275_, new_n274_, new_n259_ );
not g0138 ( new_n276_, new_n275_ );
nor g0139 ( new_n277_, new_n274_, new_n259_ );
nor g0140 ( new_n278_, new_n276_, new_n277_ );
not g0141 ( new_n279_, keyIn_0_13 );
not g0142 ( new_n280_, N113 );
nor g0143 ( new_n281_, new_n280_, N117 );
not g0144 ( new_n282_, N117 );
nor g0145 ( new_n283_, new_n282_, N113 );
nor g0146 ( new_n284_, new_n281_, new_n283_ );
not g0147 ( new_n285_, new_n284_ );
not g0148 ( new_n286_, N121 );
nor g0149 ( new_n287_, new_n286_, N125 );
not g0150 ( new_n288_, N125 );
nor g0151 ( new_n289_, new_n288_, N121 );
nor g0152 ( new_n290_, new_n287_, new_n289_ );
nand g0153 ( new_n291_, new_n285_, new_n290_ );
not g0154 ( new_n292_, new_n290_ );
nand g0155 ( new_n293_, new_n292_, new_n284_ );
nand g0156 ( new_n294_, new_n291_, new_n293_ );
nand g0157 ( new_n295_, new_n294_, new_n279_ );
not g0158 ( new_n296_, new_n295_ );
nor g0159 ( new_n297_, new_n294_, new_n279_ );
nor g0160 ( new_n298_, new_n296_, new_n297_ );
not g0161 ( new_n299_, new_n298_ );
nand g0162 ( new_n300_, new_n278_, new_n299_ );
not g0163 ( new_n301_, new_n277_ );
nand g0164 ( new_n302_, new_n301_, new_n275_ );
nand g0165 ( new_n303_, new_n302_, new_n298_ );
nand g0166 ( new_n304_, new_n300_, new_n303_ );
nand g0167 ( new_n305_, new_n304_, new_n258_ );
nor g0168 ( new_n306_, new_n304_, new_n258_ );
not g0169 ( new_n307_, new_n306_ );
nand g0170 ( new_n308_, new_n307_, new_n305_ );
nand g0171 ( new_n309_, N130, N137 );
nand g0172 ( new_n310_, new_n308_, new_n309_ );
not g0173 ( new_n311_, new_n305_ );
nor g0174 ( new_n312_, new_n311_, new_n306_ );
not g0175 ( new_n313_, new_n309_ );
nand g0176 ( new_n314_, new_n312_, new_n313_ );
nand g0177 ( new_n315_, new_n314_, new_n310_ );
nand g0178 ( new_n316_, new_n315_, new_n257_ );
not g0179 ( new_n317_, new_n316_ );
nor g0180 ( new_n318_, new_n315_, new_n257_ );
nor g0181 ( new_n319_, new_n317_, new_n318_ );
not g0182 ( new_n320_, N5 );
nor g0183 ( new_n321_, new_n320_, N21 );
not g0184 ( new_n322_, N21 );
nor g0185 ( new_n323_, new_n322_, N5 );
nor g0186 ( new_n324_, new_n321_, new_n323_ );
not g0187 ( new_n325_, N37 );
nor g0188 ( new_n326_, new_n325_, N53 );
not g0189 ( new_n327_, N53 );
nor g0190 ( new_n328_, new_n327_, N37 );
nor g0191 ( new_n329_, new_n326_, new_n328_ );
not g0192 ( new_n330_, new_n329_ );
nor g0193 ( new_n331_, new_n330_, new_n324_ );
nand g0194 ( new_n332_, new_n330_, new_n324_ );
not g0195 ( new_n333_, new_n332_ );
nor g0196 ( new_n334_, new_n333_, new_n331_ );
not g0197 ( new_n335_, new_n334_ );
nand g0198 ( new_n336_, new_n335_, keyIn_0_15 );
not g0199 ( new_n337_, new_n336_ );
nor g0200 ( new_n338_, new_n335_, keyIn_0_15 );
nor g0201 ( new_n339_, new_n337_, new_n338_ );
not g0202 ( new_n340_, new_n339_ );
nand g0203 ( new_n341_, new_n319_, new_n340_ );
nor g0204 ( new_n342_, new_n312_, new_n313_ );
nor g0205 ( new_n343_, new_n308_, new_n309_ );
nor g0206 ( new_n344_, new_n342_, new_n343_ );
nand g0207 ( new_n345_, new_n344_, keyIn_0_31 );
nand g0208 ( new_n346_, new_n345_, new_n316_ );
nand g0209 ( new_n347_, new_n346_, new_n339_ );
nand g0210 ( new_n348_, new_n341_, new_n347_ );
nand g0211 ( new_n349_, new_n348_, new_n256_ );
nor g0212 ( new_n350_, new_n346_, new_n339_ );
not g0213 ( new_n351_, new_n347_ );
nor g0214 ( new_n352_, new_n351_, new_n350_ );
nand g0215 ( new_n353_, new_n352_, keyIn_0_39 );
nand g0216 ( new_n354_, new_n353_, new_n349_ );
not g0217 ( new_n355_, keyIn_0_28 );
nor g0218 ( new_n356_, new_n166_, new_n278_ );
nor g0219 ( new_n357_, new_n189_, new_n302_ );
nor g0220 ( new_n358_, new_n356_, new_n357_ );
nor g0221 ( new_n359_, new_n358_, new_n355_ );
nand g0222 ( new_n360_, new_n189_, new_n302_ );
nand g0223 ( new_n361_, new_n166_, new_n278_ );
nand g0224 ( new_n362_, new_n361_, new_n360_ );
nor g0225 ( new_n363_, new_n362_, keyIn_0_28 );
nor g0226 ( new_n364_, new_n359_, new_n363_ );
nand g0227 ( new_n365_, N131, N137 );
not g0228 ( new_n366_, new_n365_ );
nor g0229 ( new_n367_, new_n364_, new_n366_ );
nand g0230 ( new_n368_, new_n362_, keyIn_0_28 );
nand g0231 ( new_n369_, new_n358_, new_n355_ );
nand g0232 ( new_n370_, new_n369_, new_n368_ );
nor g0233 ( new_n371_, new_n370_, new_n365_ );
nor g0234 ( new_n372_, new_n367_, new_n371_ );
nor g0235 ( new_n373_, new_n372_, keyIn_0_32 );
not g0236 ( new_n374_, keyIn_0_32 );
nand g0237 ( new_n375_, new_n370_, new_n365_ );
nand g0238 ( new_n376_, new_n364_, new_n366_ );
nand g0239 ( new_n377_, new_n376_, new_n375_ );
nor g0240 ( new_n378_, new_n377_, new_n374_ );
nor g0241 ( new_n379_, new_n373_, new_n378_ );
not g0242 ( new_n380_, N9 );
nor g0243 ( new_n381_, new_n380_, N25 );
not g0244 ( new_n382_, N25 );
nor g0245 ( new_n383_, new_n382_, N9 );
nor g0246 ( new_n384_, new_n381_, new_n383_ );
not g0247 ( new_n385_, N41 );
nor g0248 ( new_n386_, new_n385_, N57 );
not g0249 ( new_n387_, N57 );
nor g0250 ( new_n388_, new_n387_, N41 );
nor g0251 ( new_n389_, new_n386_, new_n388_ );
not g0252 ( new_n390_, new_n389_ );
nor g0253 ( new_n391_, new_n390_, new_n384_ );
nand g0254 ( new_n392_, new_n390_, new_n384_ );
not g0255 ( new_n393_, new_n392_ );
nor g0256 ( new_n394_, new_n393_, new_n391_ );
not g0257 ( new_n395_, new_n394_ );
nand g0258 ( new_n396_, new_n395_, keyIn_0_16 );
not g0259 ( new_n397_, new_n396_ );
nor g0260 ( new_n398_, new_n395_, keyIn_0_16 );
nor g0261 ( new_n399_, new_n397_, new_n398_ );
not g0262 ( new_n400_, new_n399_ );
nand g0263 ( new_n401_, new_n379_, new_n400_ );
nand g0264 ( new_n402_, new_n377_, new_n374_ );
nand g0265 ( new_n403_, new_n372_, keyIn_0_32 );
nand g0266 ( new_n404_, new_n403_, new_n402_ );
nand g0267 ( new_n405_, new_n404_, new_n399_ );
nand g0268 ( new_n406_, new_n401_, new_n405_ );
nand g0269 ( new_n407_, new_n406_, keyIn_0_40 );
not g0270 ( new_n408_, keyIn_0_40 );
nor g0271 ( new_n409_, new_n404_, new_n399_ );
nor g0272 ( new_n410_, new_n379_, new_n400_ );
nor g0273 ( new_n411_, new_n410_, new_n409_ );
nand g0274 ( new_n412_, new_n411_, new_n408_ );
nand g0275 ( new_n413_, new_n412_, new_n407_ );
nor g0276 ( new_n414_, new_n250_, new_n247_ );
nor g0277 ( new_n415_, new_n245_, keyIn_0_38 );
nor g0278 ( new_n416_, new_n414_, new_n415_ );
not g0279 ( new_n417_, keyIn_0_41 );
nand g0280 ( new_n418_, new_n185_, new_n299_ );
nand g0281 ( new_n419_, new_n193_, new_n298_ );
nand g0282 ( new_n420_, new_n418_, new_n419_ );
nand g0283 ( new_n421_, new_n420_, keyIn_0_29 );
not g0284 ( new_n422_, new_n421_ );
nor g0285 ( new_n423_, new_n420_, keyIn_0_29 );
nor g0286 ( new_n424_, new_n422_, new_n423_ );
nand g0287 ( new_n425_, N132, N137 );
not g0288 ( new_n426_, new_n425_ );
nor g0289 ( new_n427_, new_n424_, new_n426_ );
not g0290 ( new_n428_, keyIn_0_29 );
not g0291 ( new_n429_, new_n420_ );
nand g0292 ( new_n430_, new_n429_, new_n428_ );
nand g0293 ( new_n431_, new_n430_, new_n421_ );
nor g0294 ( new_n432_, new_n431_, new_n425_ );
nor g0295 ( new_n433_, new_n427_, new_n432_ );
nor g0296 ( new_n434_, new_n433_, keyIn_0_33 );
not g0297 ( new_n435_, keyIn_0_33 );
nand g0298 ( new_n436_, new_n431_, new_n425_ );
nand g0299 ( new_n437_, new_n424_, new_n426_ );
nand g0300 ( new_n438_, new_n437_, new_n436_ );
nor g0301 ( new_n439_, new_n438_, new_n435_ );
nor g0302 ( new_n440_, new_n434_, new_n439_ );
not g0303 ( new_n441_, keyIn_0_17 );
not g0304 ( new_n442_, N13 );
nor g0305 ( new_n443_, new_n442_, N29 );
not g0306 ( new_n444_, N29 );
nor g0307 ( new_n445_, new_n444_, N13 );
nor g0308 ( new_n446_, new_n443_, new_n445_ );
not g0309 ( new_n447_, N45 );
nor g0310 ( new_n448_, new_n447_, N61 );
not g0311 ( new_n449_, N61 );
nor g0312 ( new_n450_, new_n449_, N45 );
nor g0313 ( new_n451_, new_n448_, new_n450_ );
not g0314 ( new_n452_, new_n451_ );
nor g0315 ( new_n453_, new_n452_, new_n446_ );
nand g0316 ( new_n454_, new_n452_, new_n446_ );
not g0317 ( new_n455_, new_n454_ );
nor g0318 ( new_n456_, new_n455_, new_n453_ );
not g0319 ( new_n457_, new_n456_ );
nor g0320 ( new_n458_, new_n457_, new_n441_ );
nand g0321 ( new_n459_, new_n457_, new_n441_ );
not g0322 ( new_n460_, new_n459_ );
nor g0323 ( new_n461_, new_n460_, new_n458_ );
not g0324 ( new_n462_, new_n461_ );
nand g0325 ( new_n463_, new_n440_, new_n462_ );
nand g0326 ( new_n464_, new_n438_, new_n435_ );
nand g0327 ( new_n465_, new_n433_, keyIn_0_33 );
nand g0328 ( new_n466_, new_n465_, new_n464_ );
nand g0329 ( new_n467_, new_n466_, new_n461_ );
nand g0330 ( new_n468_, new_n463_, new_n467_ );
nand g0331 ( new_n469_, new_n468_, new_n417_ );
nor g0332 ( new_n470_, new_n468_, new_n417_ );
not g0333 ( new_n471_, new_n470_ );
nand g0334 ( new_n472_, new_n471_, new_n469_ );
nand g0335 ( new_n473_, new_n416_, new_n472_ );
nor g0336 ( new_n474_, new_n473_, new_n413_ );
nand g0337 ( new_n475_, new_n474_, new_n354_ );
nand g0338 ( new_n476_, new_n475_, new_n255_ );
not g0339 ( new_n477_, new_n349_ );
nor g0340 ( new_n478_, new_n348_, new_n256_ );
nor g0341 ( new_n479_, new_n477_, new_n478_ );
nor g0342 ( new_n480_, new_n411_, new_n408_ );
nor g0343 ( new_n481_, new_n406_, keyIn_0_40 );
nor g0344 ( new_n482_, new_n480_, new_n481_ );
nor g0345 ( new_n483_, new_n466_, new_n461_ );
nor g0346 ( new_n484_, new_n440_, new_n462_ );
nor g0347 ( new_n485_, new_n484_, new_n483_ );
nor g0348 ( new_n486_, new_n485_, keyIn_0_41 );
nor g0349 ( new_n487_, new_n486_, new_n470_ );
nor g0350 ( new_n488_, new_n252_, new_n487_ );
nand g0351 ( new_n489_, new_n488_, new_n482_ );
nor g0352 ( new_n490_, new_n489_, new_n479_ );
nand g0353 ( new_n491_, new_n490_, keyIn_0_47 );
nand g0354 ( new_n492_, new_n476_, new_n491_ );
nand g0355 ( new_n493_, new_n416_, new_n413_ );
nand g0356 ( new_n494_, new_n479_, new_n472_ );
nor g0357 ( new_n495_, new_n493_, new_n494_ );
nor g0358 ( new_n496_, new_n495_, keyIn_0_48 );
nand g0359 ( new_n497_, new_n495_, keyIn_0_48 );
not g0360 ( new_n498_, new_n497_ );
nor g0361 ( new_n499_, new_n498_, new_n496_ );
nand g0362 ( new_n500_, new_n492_, new_n499_ );
not g0363 ( new_n501_, keyIn_0_49 );
nand g0364 ( new_n502_, new_n252_, new_n354_ );
nor g0365 ( new_n503_, new_n502_, new_n487_ );
nand g0366 ( new_n504_, new_n503_, new_n413_ );
nand g0367 ( new_n505_, new_n504_, new_n501_ );
not g0368 ( new_n506_, new_n504_ );
nand g0369 ( new_n507_, new_n506_, keyIn_0_49 );
nand g0370 ( new_n508_, new_n507_, new_n505_ );
nor g0371 ( new_n509_, new_n493_, new_n472_ );
nand g0372 ( new_n510_, new_n509_, new_n354_ );
nand g0373 ( new_n511_, new_n510_, keyIn_0_46 );
not g0374 ( new_n512_, keyIn_0_46 );
nor g0375 ( new_n513_, new_n482_, new_n252_ );
nand g0376 ( new_n514_, new_n513_, new_n487_ );
nor g0377 ( new_n515_, new_n514_, new_n479_ );
nand g0378 ( new_n516_, new_n515_, new_n512_ );
nand g0379 ( new_n517_, new_n516_, new_n511_ );
nand g0380 ( new_n518_, new_n508_, new_n517_ );
nor g0381 ( new_n519_, new_n518_, new_n500_ );
nor g0382 ( new_n520_, new_n519_, new_n254_ );
nor g0383 ( new_n521_, new_n490_, keyIn_0_47 );
nor g0384 ( new_n522_, new_n475_, new_n255_ );
nor g0385 ( new_n523_, new_n522_, new_n521_ );
not g0386 ( new_n524_, new_n496_ );
nand g0387 ( new_n525_, new_n524_, new_n497_ );
nor g0388 ( new_n526_, new_n523_, new_n525_ );
not g0389 ( new_n527_, new_n505_ );
nor g0390 ( new_n528_, new_n504_, new_n501_ );
nor g0391 ( new_n529_, new_n527_, new_n528_ );
nor g0392 ( new_n530_, new_n515_, new_n512_ );
nor g0393 ( new_n531_, new_n510_, keyIn_0_46 );
nor g0394 ( new_n532_, new_n530_, new_n531_ );
nor g0395 ( new_n533_, new_n532_, new_n529_ );
nand g0396 ( new_n534_, new_n533_, new_n526_ );
nor g0397 ( new_n535_, new_n534_, keyIn_0_54 );
nor g0398 ( new_n536_, new_n535_, new_n520_ );
not g0399 ( new_n537_, keyIn_0_35 );
nand g0400 ( new_n538_, new_n327_, N49 );
nand g0401 ( new_n539_, new_n226_, N53 );
nand g0402 ( new_n540_, new_n538_, new_n539_ );
nand g0403 ( new_n541_, new_n540_, keyIn_0_3 );
nor g0404 ( new_n542_, new_n540_, keyIn_0_3 );
not g0405 ( new_n543_, new_n542_ );
nand g0406 ( new_n544_, new_n543_, new_n541_ );
nand g0407 ( new_n545_, new_n449_, N57 );
nand g0408 ( new_n546_, new_n387_, N61 );
nand g0409 ( new_n547_, new_n545_, new_n546_ );
nand g0410 ( new_n548_, new_n547_, keyIn_0_4 );
not g0411 ( new_n549_, new_n548_ );
nor g0412 ( new_n550_, new_n547_, keyIn_0_4 );
nor g0413 ( new_n551_, new_n549_, new_n550_ );
nand g0414 ( new_n552_, new_n551_, new_n544_ );
not g0415 ( new_n553_, new_n541_ );
nor g0416 ( new_n554_, new_n553_, new_n542_ );
not g0417 ( new_n555_, new_n550_ );
nand g0418 ( new_n556_, new_n555_, new_n548_ );
nand g0419 ( new_n557_, new_n554_, new_n556_ );
nand g0420 ( new_n558_, new_n552_, new_n557_ );
nand g0421 ( new_n559_, new_n558_, keyIn_0_9 );
nor g0422 ( new_n560_, new_n558_, keyIn_0_9 );
not g0423 ( new_n561_, new_n560_ );
nand g0424 ( new_n562_, new_n561_, new_n559_ );
not g0425 ( new_n563_, keyIn_0_8 );
nand g0426 ( new_n564_, new_n325_, N33 );
nand g0427 ( new_n565_, new_n224_, N37 );
nand g0428 ( new_n566_, new_n564_, new_n565_ );
nand g0429 ( new_n567_, new_n566_, keyIn_0_1 );
nor g0430 ( new_n568_, new_n566_, keyIn_0_1 );
not g0431 ( new_n569_, new_n568_ );
nand g0432 ( new_n570_, new_n569_, new_n567_ );
not g0433 ( new_n571_, keyIn_0_2 );
nand g0434 ( new_n572_, new_n447_, N41 );
nand g0435 ( new_n573_, new_n385_, N45 );
nand g0436 ( new_n574_, new_n572_, new_n573_ );
nand g0437 ( new_n575_, new_n574_, new_n571_ );
nor g0438 ( new_n576_, new_n574_, new_n571_ );
not g0439 ( new_n577_, new_n576_ );
nand g0440 ( new_n578_, new_n577_, new_n575_ );
nand g0441 ( new_n579_, new_n570_, new_n578_ );
not g0442 ( new_n580_, new_n570_ );
not g0443 ( new_n581_, new_n575_ );
nor g0444 ( new_n582_, new_n581_, new_n576_ );
nand g0445 ( new_n583_, new_n580_, new_n582_ );
nand g0446 ( new_n584_, new_n583_, new_n579_ );
nand g0447 ( new_n585_, new_n584_, new_n563_ );
not g0448 ( new_n586_, new_n584_ );
nand g0449 ( new_n587_, new_n586_, keyIn_0_8 );
nand g0450 ( new_n588_, new_n587_, new_n585_ );
nand g0451 ( new_n589_, new_n588_, new_n562_ );
not g0452 ( new_n590_, new_n559_ );
nor g0453 ( new_n591_, new_n590_, new_n560_ );
not g0454 ( new_n592_, new_n585_ );
nor g0455 ( new_n593_, new_n584_, new_n563_ );
nor g0456 ( new_n594_, new_n592_, new_n593_ );
nand g0457 ( new_n595_, new_n594_, new_n591_ );
nand g0458 ( new_n596_, new_n595_, new_n589_ );
nand g0459 ( new_n597_, new_n596_, keyIn_0_23 );
not g0460 ( new_n598_, keyIn_0_23 );
not g0461 ( new_n599_, new_n596_ );
nand g0462 ( new_n600_, new_n599_, new_n598_ );
nand g0463 ( new_n601_, new_n600_, new_n597_ );
nand g0464 ( new_n602_, N134, N137 );
nand g0465 ( new_n603_, new_n601_, new_n602_ );
not g0466 ( new_n604_, new_n597_ );
nor g0467 ( new_n605_, new_n596_, keyIn_0_23 );
nor g0468 ( new_n606_, new_n604_, new_n605_ );
not g0469 ( new_n607_, new_n602_ );
nand g0470 ( new_n608_, new_n606_, new_n607_ );
nand g0471 ( new_n609_, new_n608_, new_n603_ );
nand g0472 ( new_n610_, new_n609_, new_n537_ );
nor g0473 ( new_n611_, new_n606_, new_n607_ );
nor g0474 ( new_n612_, new_n601_, new_n602_ );
nor g0475 ( new_n613_, new_n611_, new_n612_ );
nand g0476 ( new_n614_, new_n613_, keyIn_0_35 );
nand g0477 ( new_n615_, new_n614_, new_n610_ );
nor g0478 ( new_n616_, new_n140_, N85 );
nor g0479 ( new_n617_, new_n169_, N69 );
nor g0480 ( new_n618_, new_n616_, new_n617_ );
nor g0481 ( new_n619_, new_n262_, N117 );
nor g0482 ( new_n620_, new_n282_, N101 );
nor g0483 ( new_n621_, new_n619_, new_n620_ );
not g0484 ( new_n622_, new_n621_ );
nor g0485 ( new_n623_, new_n622_, new_n618_ );
nand g0486 ( new_n624_, new_n622_, new_n618_ );
not g0487 ( new_n625_, new_n624_ );
nor g0488 ( new_n626_, new_n625_, new_n623_ );
not g0489 ( new_n627_, new_n626_ );
nand g0490 ( new_n628_, new_n627_, keyIn_0_19 );
not g0491 ( new_n629_, new_n628_ );
nor g0492 ( new_n630_, new_n627_, keyIn_0_19 );
nor g0493 ( new_n631_, new_n629_, new_n630_ );
nand g0494 ( new_n632_, new_n615_, new_n631_ );
not g0495 ( new_n633_, new_n610_ );
nor g0496 ( new_n634_, new_n609_, new_n537_ );
nor g0497 ( new_n635_, new_n633_, new_n634_ );
not g0498 ( new_n636_, new_n631_ );
nand g0499 ( new_n637_, new_n635_, new_n636_ );
nand g0500 ( new_n638_, new_n637_, new_n632_ );
nand g0501 ( new_n639_, new_n638_, keyIn_0_43 );
not g0502 ( new_n640_, keyIn_0_43 );
not g0503 ( new_n641_, new_n632_ );
nor g0504 ( new_n642_, new_n615_, new_n631_ );
nor g0505 ( new_n643_, new_n641_, new_n642_ );
nand g0506 ( new_n644_, new_n643_, new_n640_ );
nand g0507 ( new_n645_, new_n644_, new_n639_ );
not g0508 ( new_n646_, keyIn_0_44 );
not g0509 ( new_n647_, keyIn_0_24 );
nor g0510 ( new_n648_, new_n219_, N5 );
nor g0511 ( new_n649_, new_n320_, N1 );
nor g0512 ( new_n650_, new_n648_, new_n649_ );
not g0513 ( new_n651_, new_n650_ );
nor g0514 ( new_n652_, new_n380_, N13 );
nand g0515 ( new_n653_, new_n380_, N13 );
not g0516 ( new_n654_, new_n653_ );
nor g0517 ( new_n655_, new_n654_, new_n652_ );
nand g0518 ( new_n656_, new_n651_, new_n655_ );
not g0519 ( new_n657_, new_n655_ );
nand g0520 ( new_n658_, new_n657_, new_n650_ );
nand g0521 ( new_n659_, new_n658_, new_n656_ );
nand g0522 ( new_n660_, new_n659_, keyIn_0_6 );
not g0523 ( new_n661_, new_n660_ );
nor g0524 ( new_n662_, new_n659_, keyIn_0_6 );
nor g0525 ( new_n663_, new_n661_, new_n662_ );
nand g0526 ( new_n664_, new_n588_, new_n663_ );
not g0527 ( new_n665_, new_n663_ );
nand g0528 ( new_n666_, new_n594_, new_n665_ );
nand g0529 ( new_n667_, new_n666_, new_n664_ );
nand g0530 ( new_n668_, new_n667_, new_n647_ );
nor g0531 ( new_n669_, new_n594_, new_n665_ );
nor g0532 ( new_n670_, new_n588_, new_n663_ );
nor g0533 ( new_n671_, new_n669_, new_n670_ );
nand g0534 ( new_n672_, new_n671_, keyIn_0_24 );
nand g0535 ( new_n673_, new_n672_, new_n668_ );
nand g0536 ( new_n674_, N135, N137 );
not g0537 ( new_n675_, new_n674_ );
nand g0538 ( new_n676_, new_n673_, new_n675_ );
nor g0539 ( new_n677_, new_n671_, keyIn_0_24 );
nor g0540 ( new_n678_, new_n667_, new_n647_ );
nor g0541 ( new_n679_, new_n677_, new_n678_ );
nand g0542 ( new_n680_, new_n679_, new_n674_ );
nand g0543 ( new_n681_, new_n680_, new_n676_ );
nand g0544 ( new_n682_, new_n681_, keyIn_0_36 );
not g0545 ( new_n683_, keyIn_0_36 );
nor g0546 ( new_n684_, new_n679_, new_n674_ );
nor g0547 ( new_n685_, new_n673_, new_n675_ );
nor g0548 ( new_n686_, new_n684_, new_n685_ );
nand g0549 ( new_n687_, new_n686_, new_n683_ );
nand g0550 ( new_n688_, new_n687_, new_n682_ );
not g0551 ( new_n689_, keyIn_0_20 );
nor g0552 ( new_n690_, new_n149_, N89 );
nor g0553 ( new_n691_, new_n172_, N73 );
nor g0554 ( new_n692_, new_n690_, new_n691_ );
nor g0555 ( new_n693_, new_n265_, N121 );
nor g0556 ( new_n694_, new_n286_, N105 );
nor g0557 ( new_n695_, new_n693_, new_n694_ );
not g0558 ( new_n696_, new_n695_ );
nor g0559 ( new_n697_, new_n696_, new_n692_ );
nand g0560 ( new_n698_, new_n696_, new_n692_ );
not g0561 ( new_n699_, new_n698_ );
nor g0562 ( new_n700_, new_n699_, new_n697_ );
not g0563 ( new_n701_, new_n700_ );
nand g0564 ( new_n702_, new_n701_, new_n689_ );
not g0565 ( new_n703_, new_n702_ );
nor g0566 ( new_n704_, new_n701_, new_n689_ );
nor g0567 ( new_n705_, new_n703_, new_n704_ );
nand g0568 ( new_n706_, new_n688_, new_n705_ );
nor g0569 ( new_n707_, new_n686_, new_n683_ );
nor g0570 ( new_n708_, new_n681_, keyIn_0_36 );
nor g0571 ( new_n709_, new_n707_, new_n708_ );
not g0572 ( new_n710_, new_n705_ );
nand g0573 ( new_n711_, new_n709_, new_n710_ );
nand g0574 ( new_n712_, new_n711_, new_n706_ );
nand g0575 ( new_n713_, new_n712_, new_n646_ );
nor g0576 ( new_n714_, new_n709_, new_n710_ );
nor g0577 ( new_n715_, new_n688_, new_n705_ );
nor g0578 ( new_n716_, new_n714_, new_n715_ );
nand g0579 ( new_n717_, new_n716_, keyIn_0_44 );
nand g0580 ( new_n718_, new_n717_, new_n713_ );
nor g0581 ( new_n719_, new_n645_, new_n718_ );
not g0582 ( new_n720_, keyIn_0_37 );
not g0583 ( new_n721_, keyIn_0_25 );
nand g0584 ( new_n722_, new_n444_, N25 );
nand g0585 ( new_n723_, new_n382_, N29 );
nand g0586 ( new_n724_, new_n722_, new_n723_ );
nand g0587 ( new_n725_, new_n724_, keyIn_0_0 );
nor g0588 ( new_n726_, new_n724_, keyIn_0_0 );
not g0589 ( new_n727_, new_n726_ );
nand g0590 ( new_n728_, new_n727_, new_n725_ );
nor g0591 ( new_n729_, new_n221_, N21 );
nand g0592 ( new_n730_, new_n221_, N21 );
not g0593 ( new_n731_, new_n730_ );
nor g0594 ( new_n732_, new_n731_, new_n729_ );
not g0595 ( new_n733_, new_n732_ );
nand g0596 ( new_n734_, new_n728_, new_n733_ );
not g0597 ( new_n735_, new_n725_ );
nor g0598 ( new_n736_, new_n735_, new_n726_ );
nand g0599 ( new_n737_, new_n736_, new_n732_ );
nand g0600 ( new_n738_, new_n737_, new_n734_ );
nand g0601 ( new_n739_, new_n738_, keyIn_0_7 );
not g0602 ( new_n740_, new_n739_ );
nor g0603 ( new_n741_, new_n738_, keyIn_0_7 );
nor g0604 ( new_n742_, new_n740_, new_n741_ );
nand g0605 ( new_n743_, new_n562_, new_n742_ );
not g0606 ( new_n744_, new_n741_ );
nand g0607 ( new_n745_, new_n744_, new_n739_ );
nand g0608 ( new_n746_, new_n591_, new_n745_ );
nand g0609 ( new_n747_, new_n746_, new_n743_ );
nand g0610 ( new_n748_, new_n747_, new_n721_ );
nor g0611 ( new_n749_, new_n747_, new_n721_ );
not g0612 ( new_n750_, new_n749_ );
nand g0613 ( new_n751_, new_n750_, new_n748_ );
nand g0614 ( new_n752_, N136, N137 );
not g0615 ( new_n753_, new_n752_ );
nand g0616 ( new_n754_, new_n751_, new_n753_ );
not g0617 ( new_n755_, new_n748_ );
nor g0618 ( new_n756_, new_n755_, new_n749_ );
nand g0619 ( new_n757_, new_n756_, new_n752_ );
nand g0620 ( new_n758_, new_n757_, new_n754_ );
nand g0621 ( new_n759_, new_n758_, new_n720_ );
nor g0622 ( new_n760_, new_n756_, new_n752_ );
nor g0623 ( new_n761_, new_n751_, new_n753_ );
nor g0624 ( new_n762_, new_n760_, new_n761_ );
nand g0625 ( new_n763_, new_n762_, keyIn_0_37 );
nand g0626 ( new_n764_, new_n763_, new_n759_ );
nor g0627 ( new_n765_, new_n151_, N93 );
nor g0628 ( new_n766_, new_n174_, N77 );
nor g0629 ( new_n767_, new_n765_, new_n766_ );
nor g0630 ( new_n768_, new_n267_, N125 );
nor g0631 ( new_n769_, new_n288_, N109 );
nor g0632 ( new_n770_, new_n768_, new_n769_ );
not g0633 ( new_n771_, new_n770_ );
nor g0634 ( new_n772_, new_n771_, new_n767_ );
nand g0635 ( new_n773_, new_n771_, new_n767_ );
not g0636 ( new_n774_, new_n773_ );
nor g0637 ( new_n775_, new_n774_, new_n772_ );
not g0638 ( new_n776_, new_n775_ );
nand g0639 ( new_n777_, new_n776_, keyIn_0_21 );
not g0640 ( new_n778_, new_n777_ );
nor g0641 ( new_n779_, new_n776_, keyIn_0_21 );
nor g0642 ( new_n780_, new_n778_, new_n779_ );
not g0643 ( new_n781_, new_n780_ );
nand g0644 ( new_n782_, new_n764_, new_n781_ );
not g0645 ( new_n783_, new_n759_ );
nor g0646 ( new_n784_, new_n758_, new_n720_ );
nor g0647 ( new_n785_, new_n783_, new_n784_ );
nand g0648 ( new_n786_, new_n785_, new_n780_ );
nand g0649 ( new_n787_, new_n786_, new_n782_ );
nand g0650 ( new_n788_, new_n787_, keyIn_0_45 );
not g0651 ( new_n789_, new_n788_ );
nor g0652 ( new_n790_, new_n787_, keyIn_0_45 );
nor g0653 ( new_n791_, new_n789_, new_n790_ );
nand g0654 ( new_n792_, new_n745_, new_n665_ );
nand g0655 ( new_n793_, new_n742_, new_n663_ );
nand g0656 ( new_n794_, new_n793_, new_n792_ );
nand g0657 ( new_n795_, new_n794_, keyIn_0_22 );
nor g0658 ( new_n796_, new_n794_, keyIn_0_22 );
not g0659 ( new_n797_, new_n796_ );
nand g0660 ( new_n798_, new_n797_, new_n795_ );
nand g0661 ( new_n799_, N133, N137 );
not g0662 ( new_n800_, new_n799_ );
nand g0663 ( new_n801_, new_n798_, new_n800_ );
not g0664 ( new_n802_, new_n795_ );
nor g0665 ( new_n803_, new_n802_, new_n796_ );
nand g0666 ( new_n804_, new_n803_, new_n799_ );
nand g0667 ( new_n805_, new_n804_, new_n801_ );
nand g0668 ( new_n806_, new_n805_, keyIn_0_34 );
nor g0669 ( new_n807_, new_n805_, keyIn_0_34 );
not g0670 ( new_n808_, new_n807_ );
nand g0671 ( new_n809_, new_n808_, new_n806_ );
not g0672 ( new_n810_, keyIn_0_18 );
nor g0673 ( new_n811_, new_n142_, N81 );
nor g0674 ( new_n812_, new_n167_, N65 );
nor g0675 ( new_n813_, new_n811_, new_n812_ );
nor g0676 ( new_n814_, new_n260_, N113 );
nor g0677 ( new_n815_, new_n280_, N97 );
nor g0678 ( new_n816_, new_n814_, new_n815_ );
not g0679 ( new_n817_, new_n816_ );
nor g0680 ( new_n818_, new_n817_, new_n813_ );
nand g0681 ( new_n819_, new_n817_, new_n813_ );
not g0682 ( new_n820_, new_n819_ );
nor g0683 ( new_n821_, new_n820_, new_n818_ );
not g0684 ( new_n822_, new_n821_ );
nand g0685 ( new_n823_, new_n822_, new_n810_ );
not g0686 ( new_n824_, new_n823_ );
nor g0687 ( new_n825_, new_n822_, new_n810_ );
nor g0688 ( new_n826_, new_n824_, new_n825_ );
not g0689 ( new_n827_, new_n826_ );
nand g0690 ( new_n828_, new_n809_, new_n827_ );
not g0691 ( new_n829_, new_n806_ );
nor g0692 ( new_n830_, new_n829_, new_n807_ );
nand g0693 ( new_n831_, new_n830_, new_n826_ );
nand g0694 ( new_n832_, new_n831_, new_n828_ );
nand g0695 ( new_n833_, new_n832_, keyIn_0_42 );
not g0696 ( new_n834_, new_n833_ );
nor g0697 ( new_n835_, new_n832_, keyIn_0_42 );
nor g0698 ( new_n836_, new_n834_, new_n835_ );
nor g0699 ( new_n837_, new_n791_, new_n836_ );
nand g0700 ( new_n838_, new_n837_, new_n719_ );
not g0701 ( new_n839_, new_n838_ );
nand g0702 ( new_n840_, new_n536_, new_n839_ );
nand g0703 ( new_n841_, new_n840_, new_n253_ );
nand g0704 ( new_n842_, new_n534_, keyIn_0_54 );
nand g0705 ( new_n843_, new_n519_, new_n254_ );
nand g0706 ( new_n844_, new_n842_, new_n843_ );
nor g0707 ( new_n845_, new_n844_, new_n838_ );
nand g0708 ( new_n846_, new_n845_, keyIn_0_56 );
nand g0709 ( new_n847_, new_n841_, new_n846_ );
nand g0710 ( new_n848_, new_n847_, new_n252_ );
nand g0711 ( new_n849_, new_n848_, N1 );
nor g0712 ( new_n850_, new_n845_, keyIn_0_56 );
nor g0713 ( new_n851_, new_n840_, new_n253_ );
nor g0714 ( new_n852_, new_n851_, new_n850_ );
nor g0715 ( new_n853_, new_n852_, new_n416_ );
nand g0716 ( new_n854_, new_n853_, new_n219_ );
nand g0717 ( N724, new_n854_, new_n849_ );
nand g0718 ( new_n856_, new_n847_, new_n479_ );
nand g0719 ( new_n857_, new_n856_, N5 );
nor g0720 ( new_n858_, new_n852_, new_n354_ );
nand g0721 ( new_n859_, new_n858_, new_n320_ );
nand g0722 ( N725, new_n859_, new_n857_ );
nand g0723 ( new_n861_, new_n847_, new_n482_ );
nand g0724 ( new_n862_, new_n861_, N9 );
nor g0725 ( new_n863_, new_n852_, new_n413_ );
nand g0726 ( new_n864_, new_n863_, new_n380_ );
nand g0727 ( N726, new_n864_, new_n862_ );
nand g0728 ( new_n866_, new_n847_, new_n487_ );
nand g0729 ( new_n867_, new_n866_, N13 );
nor g0730 ( new_n868_, new_n852_, new_n472_ );
nand g0731 ( new_n869_, new_n868_, new_n442_ );
nand g0732 ( N727, new_n869_, new_n867_ );
not g0733 ( new_n871_, keyIn_0_57 );
not g0734 ( new_n872_, new_n639_ );
nor g0735 ( new_n873_, new_n638_, keyIn_0_43 );
nor g0736 ( new_n874_, new_n872_, new_n873_ );
not g0737 ( new_n875_, keyIn_0_42 );
nor g0738 ( new_n876_, new_n830_, new_n826_ );
nor g0739 ( new_n877_, new_n809_, new_n827_ );
nor g0740 ( new_n878_, new_n876_, new_n877_ );
nand g0741 ( new_n879_, new_n878_, new_n875_ );
nand g0742 ( new_n880_, new_n879_, new_n833_ );
nand g0743 ( new_n881_, new_n874_, new_n880_ );
nand g0744 ( new_n882_, new_n791_, new_n718_ );
nor g0745 ( new_n883_, new_n881_, new_n882_ );
nand g0746 ( new_n884_, new_n536_, new_n883_ );
nand g0747 ( new_n885_, new_n884_, new_n871_ );
not g0748 ( new_n886_, new_n883_ );
nor g0749 ( new_n887_, new_n844_, new_n886_ );
nand g0750 ( new_n888_, new_n887_, keyIn_0_57 );
nand g0751 ( new_n889_, new_n885_, new_n888_ );
nand g0752 ( new_n890_, new_n889_, new_n252_ );
nand g0753 ( new_n891_, new_n890_, N17 );
nor g0754 ( new_n892_, new_n887_, keyIn_0_57 );
nor g0755 ( new_n893_, new_n884_, new_n871_ );
nor g0756 ( new_n894_, new_n893_, new_n892_ );
nor g0757 ( new_n895_, new_n894_, new_n416_ );
nand g0758 ( new_n896_, new_n895_, new_n221_ );
nand g0759 ( N728, new_n896_, new_n891_ );
nand g0760 ( new_n898_, new_n889_, new_n479_ );
nand g0761 ( new_n899_, new_n898_, N21 );
nor g0762 ( new_n900_, new_n894_, new_n354_ );
nand g0763 ( new_n901_, new_n900_, new_n322_ );
nand g0764 ( N729, new_n901_, new_n899_ );
nand g0765 ( new_n903_, new_n889_, new_n482_ );
nand g0766 ( new_n904_, new_n903_, N25 );
nor g0767 ( new_n905_, new_n894_, new_n413_ );
nand g0768 ( new_n906_, new_n905_, new_n382_ );
nand g0769 ( N730, new_n906_, new_n904_ );
nand g0770 ( new_n908_, new_n889_, new_n487_ );
nand g0771 ( new_n909_, new_n908_, N29 );
nor g0772 ( new_n910_, new_n894_, new_n472_ );
nand g0773 ( new_n911_, new_n910_, new_n444_ );
nand g0774 ( N731, new_n911_, new_n909_ );
nor g0775 ( new_n913_, new_n791_, new_n880_ );
nor g0776 ( new_n914_, new_n874_, new_n718_ );
nand g0777 ( new_n915_, new_n914_, new_n913_ );
not g0778 ( new_n916_, new_n915_ );
nand g0779 ( new_n917_, new_n536_, new_n916_ );
nor g0780 ( new_n918_, new_n917_, keyIn_0_58 );
not g0781 ( new_n919_, new_n918_ );
not g0782 ( new_n920_, keyIn_0_58 );
nor g0783 ( new_n921_, new_n844_, new_n915_ );
nor g0784 ( new_n922_, new_n921_, new_n920_ );
nor g0785 ( new_n923_, new_n922_, new_n416_ );
nand g0786 ( new_n924_, new_n923_, new_n919_ );
nand g0787 ( new_n925_, new_n924_, N33 );
nand g0788 ( new_n926_, new_n917_, keyIn_0_58 );
nand g0789 ( new_n927_, new_n926_, new_n252_ );
nor g0790 ( new_n928_, new_n927_, new_n918_ );
nand g0791 ( new_n929_, new_n928_, new_n224_ );
nand g0792 ( N732, new_n925_, new_n929_ );
nor g0793 ( new_n931_, new_n922_, new_n354_ );
nand g0794 ( new_n932_, new_n931_, new_n919_ );
nand g0795 ( new_n933_, new_n932_, N37 );
nand g0796 ( new_n934_, new_n926_, new_n479_ );
nor g0797 ( new_n935_, new_n934_, new_n918_ );
nand g0798 ( new_n936_, new_n935_, new_n325_ );
nand g0799 ( N733, new_n933_, new_n936_ );
nor g0800 ( new_n938_, new_n922_, new_n413_ );
nand g0801 ( new_n939_, new_n938_, new_n919_ );
nand g0802 ( new_n940_, new_n939_, N41 );
nand g0803 ( new_n941_, new_n926_, new_n482_ );
nor g0804 ( new_n942_, new_n941_, new_n918_ );
nand g0805 ( new_n943_, new_n942_, new_n385_ );
nand g0806 ( N734, new_n940_, new_n943_ );
nor g0807 ( new_n945_, new_n922_, new_n472_ );
nand g0808 ( new_n946_, new_n945_, new_n919_ );
nand g0809 ( new_n947_, new_n946_, N45 );
nand g0810 ( new_n948_, new_n926_, new_n487_ );
nor g0811 ( new_n949_, new_n948_, new_n918_ );
nand g0812 ( new_n950_, new_n949_, new_n447_ );
nand g0813 ( N735, new_n947_, new_n950_ );
not g0814 ( new_n952_, keyIn_0_59 );
nor g0815 ( new_n953_, new_n716_, keyIn_0_44 );
nor g0816 ( new_n954_, new_n712_, new_n646_ );
nor g0817 ( new_n955_, new_n953_, new_n954_ );
not g0818 ( new_n956_, keyIn_0_45 );
not g0819 ( new_n957_, new_n782_ );
nor g0820 ( new_n958_, new_n764_, new_n781_ );
nor g0821 ( new_n959_, new_n957_, new_n958_ );
nand g0822 ( new_n960_, new_n959_, new_n956_ );
nand g0823 ( new_n961_, new_n960_, new_n788_ );
nor g0824 ( new_n962_, new_n955_, new_n961_ );
nor g0825 ( new_n963_, new_n874_, new_n880_ );
nand g0826 ( new_n964_, new_n963_, new_n962_ );
not g0827 ( new_n965_, new_n964_ );
nand g0828 ( new_n966_, new_n536_, new_n965_ );
nand g0829 ( new_n967_, new_n966_, new_n952_ );
nor g0830 ( new_n968_, new_n844_, new_n964_ );
nand g0831 ( new_n969_, new_n968_, keyIn_0_59 );
nand g0832 ( new_n970_, new_n967_, new_n969_ );
nand g0833 ( new_n971_, new_n970_, new_n252_ );
nand g0834 ( new_n972_, new_n971_, N49 );
nor g0835 ( new_n973_, new_n968_, keyIn_0_59 );
nor g0836 ( new_n974_, new_n966_, new_n952_ );
nor g0837 ( new_n975_, new_n974_, new_n973_ );
nor g0838 ( new_n976_, new_n975_, new_n416_ );
nand g0839 ( new_n977_, new_n976_, new_n226_ );
nand g0840 ( N736, new_n977_, new_n972_ );
nand g0841 ( new_n979_, new_n970_, new_n479_ );
nand g0842 ( new_n980_, new_n979_, N53 );
nor g0843 ( new_n981_, new_n975_, new_n354_ );
nand g0844 ( new_n982_, new_n981_, new_n327_ );
nand g0845 ( N737, new_n982_, new_n980_ );
nand g0846 ( new_n984_, new_n970_, new_n482_ );
nand g0847 ( new_n985_, new_n984_, N57 );
nor g0848 ( new_n986_, new_n975_, new_n413_ );
nand g0849 ( new_n987_, new_n986_, new_n387_ );
nand g0850 ( N738, new_n987_, new_n985_ );
nand g0851 ( new_n989_, new_n970_, new_n487_ );
nand g0852 ( new_n990_, new_n989_, N61 );
nor g0853 ( new_n991_, new_n975_, new_n472_ );
nand g0854 ( new_n992_, new_n991_, new_n449_ );
nand g0855 ( N739, new_n992_, new_n990_ );
not g0856 ( new_n994_, keyIn_0_60 );
not g0857 ( new_n995_, keyIn_0_55 );
nand g0858 ( new_n996_, new_n836_, new_n961_ );
nand g0859 ( new_n997_, new_n645_, new_n718_ );
nor g0860 ( new_n998_, new_n996_, new_n997_ );
nor g0861 ( new_n999_, new_n998_, keyIn_0_52 );
not g0862 ( new_n1000_, keyIn_0_52 );
not g0863 ( new_n1001_, new_n997_ );
nand g0864 ( new_n1002_, new_n1001_, new_n913_ );
nor g0865 ( new_n1003_, new_n1002_, new_n1000_ );
nor g0866 ( new_n1004_, new_n1003_, new_n999_ );
not g0867 ( new_n1005_, keyIn_0_51 );
nand g0868 ( new_n1006_, new_n913_, new_n719_ );
nand g0869 ( new_n1007_, new_n1006_, new_n1005_ );
nor g0870 ( new_n1008_, new_n645_, new_n880_ );
nand g0871 ( new_n1009_, new_n961_, keyIn_0_51 );
nor g0872 ( new_n1010_, new_n1009_, new_n718_ );
nand g0873 ( new_n1011_, new_n1010_, new_n1008_ );
nand g0874 ( new_n1012_, new_n1007_, new_n1011_ );
nor g0875 ( new_n1013_, new_n1004_, new_n1012_ );
nor g0876 ( new_n1014_, new_n836_, new_n645_ );
nand g0877 ( new_n1015_, new_n718_, new_n961_ );
not g0878 ( new_n1016_, new_n1015_ );
nand g0879 ( new_n1017_, new_n1016_, new_n1014_ );
nand g0880 ( new_n1018_, new_n1017_, keyIn_0_53 );
not g0881 ( new_n1019_, keyIn_0_53 );
nor g0882 ( new_n1020_, new_n881_, new_n1015_ );
nand g0883 ( new_n1021_, new_n1020_, new_n1019_ );
nand g0884 ( new_n1022_, new_n1021_, new_n1018_ );
not g0885 ( new_n1023_, keyIn_0_50 );
nand g0886 ( new_n1024_, new_n962_, new_n1008_ );
nand g0887 ( new_n1025_, new_n1024_, new_n1023_ );
nand g0888 ( new_n1026_, new_n874_, new_n836_ );
nor g0889 ( new_n1027_, new_n1026_, new_n882_ );
nand g0890 ( new_n1028_, new_n1027_, keyIn_0_50 );
nand g0891 ( new_n1029_, new_n1028_, new_n1025_ );
nand g0892 ( new_n1030_, new_n1022_, new_n1029_ );
not g0893 ( new_n1031_, new_n1030_ );
nand g0894 ( new_n1032_, new_n1031_, new_n1013_ );
nand g0895 ( new_n1033_, new_n1032_, new_n995_ );
nand g0896 ( new_n1034_, new_n1002_, new_n1000_ );
nand g0897 ( new_n1035_, new_n998_, keyIn_0_52 );
nand g0898 ( new_n1036_, new_n1034_, new_n1035_ );
not g0899 ( new_n1037_, new_n1012_ );
nand g0900 ( new_n1038_, new_n1037_, new_n1036_ );
nor g0901 ( new_n1039_, new_n1038_, new_n1030_ );
nand g0902 ( new_n1040_, new_n1039_, keyIn_0_55 );
nand g0903 ( new_n1041_, new_n1033_, new_n1040_ );
not g0904 ( new_n1042_, new_n502_ );
nand g0905 ( new_n1043_, new_n1042_, new_n472_ );
nor g0906 ( new_n1044_, new_n1043_, new_n413_ );
nand g0907 ( new_n1045_, new_n1041_, new_n1044_ );
nor g0908 ( new_n1046_, new_n1045_, new_n994_ );
nand g0909 ( new_n1047_, new_n1045_, new_n994_ );
nand g0910 ( new_n1048_, new_n1047_, new_n880_ );
nor g0911 ( new_n1049_, new_n1048_, new_n1046_ );
not g0912 ( new_n1050_, new_n1049_ );
nand g0913 ( new_n1051_, new_n1050_, N65 );
nand g0914 ( new_n1052_, new_n1049_, new_n142_ );
nand g0915 ( N740, new_n1051_, new_n1052_ );
nand g0916 ( new_n1054_, new_n1047_, new_n645_ );
nor g0917 ( new_n1055_, new_n1054_, new_n1046_ );
not g0918 ( new_n1056_, new_n1055_ );
nand g0919 ( new_n1057_, new_n1056_, N69 );
nand g0920 ( new_n1058_, new_n1055_, new_n140_ );
nand g0921 ( N741, new_n1057_, new_n1058_ );
nand g0922 ( new_n1060_, new_n1047_, new_n955_ );
nor g0923 ( new_n1061_, new_n1060_, new_n1046_ );
not g0924 ( new_n1062_, new_n1061_ );
nand g0925 ( new_n1063_, new_n1062_, N73 );
nand g0926 ( new_n1064_, new_n1061_, new_n149_ );
nand g0927 ( N742, new_n1063_, new_n1064_ );
nand g0928 ( new_n1066_, new_n1047_, new_n791_ );
nor g0929 ( new_n1067_, new_n1066_, new_n1046_ );
not g0930 ( new_n1068_, new_n1067_ );
nand g0931 ( new_n1069_, new_n1068_, N77 );
nand g0932 ( new_n1070_, new_n1067_, new_n151_ );
nand g0933 ( N743, new_n1069_, new_n1070_ );
nor g0934 ( new_n1072_, new_n482_, new_n472_ );
nand g0935 ( new_n1073_, new_n1042_, new_n1072_ );
not g0936 ( new_n1074_, new_n1073_ );
nand g0937 ( new_n1075_, new_n1041_, new_n1074_ );
nand g0938 ( new_n1076_, new_n1075_, keyIn_0_61 );
nor g0939 ( new_n1077_, new_n1075_, keyIn_0_61 );
not g0940 ( new_n1078_, new_n1077_ );
nand g0941 ( new_n1079_, new_n1078_, new_n1076_ );
nand g0942 ( new_n1080_, new_n1079_, new_n880_ );
nand g0943 ( new_n1081_, new_n1080_, N81 );
not g0944 ( new_n1082_, new_n1076_ );
nor g0945 ( new_n1083_, new_n1082_, new_n1077_ );
nor g0946 ( new_n1084_, new_n1083_, new_n836_ );
nand g0947 ( new_n1085_, new_n1084_, new_n167_ );
nand g0948 ( N744, new_n1085_, new_n1081_ );
nand g0949 ( new_n1087_, new_n1079_, new_n645_ );
nand g0950 ( new_n1088_, new_n1087_, N85 );
nor g0951 ( new_n1089_, new_n1083_, new_n874_ );
nand g0952 ( new_n1090_, new_n1089_, new_n169_ );
nand g0953 ( N745, new_n1090_, new_n1088_ );
nand g0954 ( new_n1092_, new_n1079_, new_n955_ );
nand g0955 ( new_n1093_, new_n1092_, N89 );
nor g0956 ( new_n1094_, new_n1083_, new_n718_ );
nand g0957 ( new_n1095_, new_n1094_, new_n172_ );
nand g0958 ( N746, new_n1095_, new_n1093_ );
nand g0959 ( new_n1097_, new_n1079_, new_n791_ );
nand g0960 ( new_n1098_, new_n1097_, N93 );
nor g0961 ( new_n1099_, new_n1083_, new_n961_ );
nand g0962 ( new_n1100_, new_n1099_, new_n174_ );
nand g0963 ( N747, new_n1100_, new_n1098_ );
not g0964 ( new_n1102_, keyIn_0_62 );
nor g0965 ( new_n1103_, new_n489_, new_n354_ );
nand g0966 ( new_n1104_, new_n1041_, new_n1103_ );
nor g0967 ( new_n1105_, new_n1104_, new_n1102_ );
nand g0968 ( new_n1106_, new_n1104_, new_n1102_ );
nand g0969 ( new_n1107_, new_n1106_, new_n880_ );
nor g0970 ( new_n1108_, new_n1107_, new_n1105_ );
not g0971 ( new_n1109_, new_n1108_ );
nand g0972 ( new_n1110_, new_n1109_, N97 );
nand g0973 ( new_n1111_, new_n1108_, new_n260_ );
nand g0974 ( N748, new_n1110_, new_n1111_ );
nand g0975 ( new_n1113_, new_n1106_, new_n645_ );
nor g0976 ( new_n1114_, new_n1113_, new_n1105_ );
not g0977 ( new_n1115_, new_n1114_ );
nand g0978 ( new_n1116_, new_n1115_, N101 );
nand g0979 ( new_n1117_, new_n1114_, new_n262_ );
nand g0980 ( N749, new_n1116_, new_n1117_ );
nand g0981 ( new_n1119_, new_n1106_, new_n955_ );
nor g0982 ( new_n1120_, new_n1119_, new_n1105_ );
not g0983 ( new_n1121_, new_n1120_ );
nand g0984 ( new_n1122_, new_n1121_, N105 );
nand g0985 ( new_n1123_, new_n1120_, new_n265_ );
nand g0986 ( N750, new_n1122_, new_n1123_ );
nand g0987 ( new_n1125_, new_n1106_, new_n791_ );
nor g0988 ( new_n1126_, new_n1125_, new_n1105_ );
not g0989 ( new_n1127_, new_n1126_ );
nand g0990 ( new_n1128_, new_n1127_, N109 );
nand g0991 ( new_n1129_, new_n1126_, new_n267_ );
nand g0992 ( N751, new_n1128_, new_n1129_ );
nor g0993 ( new_n1131_, new_n514_, new_n354_ );
nand g0994 ( new_n1132_, new_n1041_, new_n1131_ );
nand g0995 ( new_n1133_, new_n1132_, keyIn_0_63 );
nor g0996 ( new_n1134_, new_n1132_, keyIn_0_63 );
not g0997 ( new_n1135_, new_n1134_ );
nand g0998 ( new_n1136_, new_n1135_, new_n1133_ );
nand g0999 ( new_n1137_, new_n1136_, new_n880_ );
nand g1000 ( new_n1138_, new_n1137_, N113 );
not g1001 ( new_n1139_, new_n1133_ );
nor g1002 ( new_n1140_, new_n1139_, new_n1134_ );
nor g1003 ( new_n1141_, new_n1140_, new_n836_ );
nand g1004 ( new_n1142_, new_n1141_, new_n280_ );
nand g1005 ( N752, new_n1142_, new_n1138_ );
nand g1006 ( new_n1144_, new_n1136_, new_n645_ );
nand g1007 ( new_n1145_, new_n1144_, N117 );
nor g1008 ( new_n1146_, new_n1140_, new_n874_ );
nand g1009 ( new_n1147_, new_n1146_, new_n282_ );
nand g1010 ( N753, new_n1147_, new_n1145_ );
nand g1011 ( new_n1149_, new_n1136_, new_n955_ );
nand g1012 ( new_n1150_, new_n1149_, N121 );
nor g1013 ( new_n1151_, new_n1140_, new_n718_ );
nand g1014 ( new_n1152_, new_n1151_, new_n286_ );
nand g1015 ( N754, new_n1152_, new_n1150_ );
nand g1016 ( new_n1154_, new_n1136_, new_n791_ );
nand g1017 ( new_n1155_, new_n1154_, N125 );
nor g1018 ( new_n1156_, new_n1140_, new_n961_ );
nand g1019 ( new_n1157_, new_n1156_, new_n288_ );
nand g1020 ( N755, new_n1157_, new_n1155_ );
endmodule