module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n614_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n847_, new_n250_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n170_, new_n246_, new_n682_, new_n812_, new_n679_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n853_, new_n602_, new_n114_, new_n188_, new_n240_, new_n660_, new_n413_, new_n695_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n500_, new_n786_, new_n799_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n862_, new_n742_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n774_, new_n157_, new_n716_, new_n153_, new_n792_, new_n133_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n110_, new_n315_, new_n685_, new_n124_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n849_, new_n606_, new_n589_, new_n796_, new_n248_, new_n350_, new_n117_, new_n655_, new_n630_, new_n759_, new_n167_, new_n385_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n764_, new_n150_, new_n683_, new_n108_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n845_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n650_, new_n708_, new_n750_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n875_, new_n506_, new_n680_, new_n872_, new_n256_, new_n778_, new_n452_, new_n381_, new_n656_, new_n820_, new_n771_, new_n388_, new_n508_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n882_, new_n657_, new_n652_, new_n314_, new_n582_, new_n118_, new_n363_, new_n165_, new_n441_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n207_, new_n267_, new_n473_, new_n140_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n621_, new_n846_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n874_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n870_, new_n805_, new_n559_, new_n762_, new_n838_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n794_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n369_, new_n448_, new_n867_, new_n276_, new_n688_, new_n155_, new_n384_, new_n410_, new_n851_, new_n878_, new_n543_, new_n113_, new_n775_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n259_, new_n362_, new_n809_, new_n654_, new_n713_, new_n880_, new_n604_, new_n227_, new_n416_, new_n222_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n130_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n138_, new_n749_, new_n861_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n562_, new_n578_, new_n126_, new_n808_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n800_, new_n379_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n824_, new_n143_, new_n520_, new_n125_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n106_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n748_, new_n107_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n879_, new_n151_, new_n513_, new_n592_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n191_, new_n755_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n112_, new_n856_, new_n121_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n737_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n662_, new_n864_, new_n440_, new_n733_, new_n122_, new_n531_, new_n593_, new_n111_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n115_, new_n307_, new_n852_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n134_, new_n769_, new_n651_, new_n433_, new_n435_, new_n109_, new_n776_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n815_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n129_, new_n711_, new_n644_, new_n599_, new_n836_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n818_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n754_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n727_, new_n375_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n357_, new_n320_, new_n780_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n128_, new_n358_, new_n877_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n802_, new_n697_, new_n185_, new_n709_, new_n373_, new_n866_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n770_, new_n618_, new_n120_, new_n521_, new_n793_, new_n863_, new_n406_, new_n828_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n135_, new_n573_, new_n765_, new_n405_;

not g000 ( new_n106_, keyIn_0_0 );
not g001 ( new_n107_, N5 );
and g002 ( new_n108_, new_n107_, N1 );
not g003 ( new_n109_, N1 );
and g004 ( new_n110_, new_n109_, N5 );
or g005 ( new_n111_, new_n108_, new_n110_ );
not g006 ( new_n112_, N13 );
and g007 ( new_n113_, new_n112_, N9 );
not g008 ( new_n114_, N9 );
and g009 ( new_n115_, new_n114_, N13 );
or g010 ( new_n116_, new_n113_, new_n115_ );
not g011 ( new_n117_, new_n116_ );
and g012 ( new_n118_, new_n117_, new_n111_ );
not g013 ( new_n119_, new_n111_ );
and g014 ( new_n120_, new_n119_, new_n116_ );
or g015 ( new_n121_, new_n118_, new_n120_ );
and g016 ( new_n122_, new_n121_, new_n106_ );
not g017 ( new_n123_, new_n122_ );
or g018 ( new_n124_, new_n121_, new_n106_ );
and g019 ( new_n125_, new_n123_, new_n124_ );
not g020 ( new_n126_, N37 );
and g021 ( new_n127_, new_n126_, N33 );
not g022 ( new_n128_, N33 );
and g023 ( new_n129_, new_n128_, N37 );
or g024 ( new_n130_, new_n127_, new_n129_ );
not g025 ( new_n131_, new_n130_ );
not g026 ( new_n132_, N45 );
and g027 ( new_n133_, new_n132_, N41 );
not g028 ( new_n134_, N41 );
and g029 ( new_n135_, new_n134_, N45 );
or g030 ( new_n136_, new_n133_, new_n135_ );
not g031 ( new_n137_, new_n136_ );
and g032 ( new_n138_, new_n131_, new_n137_ );
and g033 ( new_n139_, new_n130_, new_n136_ );
or g034 ( new_n140_, new_n138_, new_n139_ );
or g035 ( new_n141_, new_n140_, keyIn_0_2 );
not g036 ( new_n142_, new_n141_ );
and g037 ( new_n143_, new_n140_, keyIn_0_2 );
or g038 ( new_n144_, new_n142_, new_n143_ );
and g039 ( new_n145_, new_n144_, new_n125_ );
not g040 ( new_n146_, new_n118_ );
not g041 ( new_n147_, new_n120_ );
and g042 ( new_n148_, new_n146_, new_n147_ );
and g043 ( new_n149_, new_n148_, keyIn_0_0 );
or g044 ( new_n150_, new_n149_, new_n122_ );
not g045 ( new_n151_, new_n143_ );
and g046 ( new_n152_, new_n151_, new_n141_ );
and g047 ( new_n153_, new_n150_, new_n152_ );
or g048 ( new_n154_, new_n145_, new_n153_ );
and g049 ( new_n155_, new_n154_, keyIn_0_18 );
not g050 ( new_n156_, keyIn_0_18 );
or g051 ( new_n157_, new_n150_, new_n152_ );
or g052 ( new_n158_, new_n144_, new_n125_ );
and g053 ( new_n159_, new_n158_, new_n157_ );
and g054 ( new_n160_, new_n159_, new_n156_ );
or g055 ( new_n161_, new_n155_, new_n160_ );
and g056 ( new_n162_, N135, N137 );
and g057 ( new_n163_, new_n161_, new_n162_ );
or g058 ( new_n164_, new_n159_, new_n156_ );
or g059 ( new_n165_, new_n154_, keyIn_0_18 );
and g060 ( new_n166_, new_n165_, new_n164_ );
not g061 ( new_n167_, new_n162_ );
and g062 ( new_n168_, new_n166_, new_n167_ );
or g063 ( new_n169_, new_n163_, new_n168_ );
and g064 ( new_n170_, new_n169_, keyIn_0_30 );
not g065 ( new_n171_, keyIn_0_30 );
or g066 ( new_n172_, new_n166_, new_n167_ );
or g067 ( new_n173_, new_n161_, new_n162_ );
and g068 ( new_n174_, new_n173_, new_n172_ );
and g069 ( new_n175_, new_n174_, new_n171_ );
or g070 ( new_n176_, new_n170_, new_n175_ );
not g071 ( new_n177_, N121 );
and g072 ( new_n178_, new_n177_, N105 );
not g073 ( new_n179_, N105 );
and g074 ( new_n180_, new_n179_, N121 );
or g075 ( new_n181_, new_n178_, new_n180_ );
and g076 ( new_n182_, N73, N89 );
not g077 ( new_n183_, N73 );
not g078 ( new_n184_, N89 );
and g079 ( new_n185_, new_n183_, new_n184_ );
or g080 ( new_n186_, new_n185_, new_n182_ );
and g081 ( new_n187_, new_n181_, new_n186_ );
not g082 ( new_n188_, new_n187_ );
or g083 ( new_n189_, new_n181_, new_n186_ );
and g084 ( new_n190_, new_n188_, new_n189_ );
not g085 ( new_n191_, new_n190_ );
and g086 ( new_n192_, new_n191_, keyIn_0_14 );
not g087 ( new_n193_, new_n192_ );
or g088 ( new_n194_, new_n191_, keyIn_0_14 );
and g089 ( new_n195_, new_n193_, new_n194_ );
and g090 ( new_n196_, new_n176_, new_n195_ );
or g091 ( new_n197_, new_n174_, new_n171_ );
or g092 ( new_n198_, new_n169_, keyIn_0_30 );
and g093 ( new_n199_, new_n198_, new_n197_ );
not g094 ( new_n200_, new_n195_ );
and g095 ( new_n201_, new_n199_, new_n200_ );
or g096 ( new_n202_, new_n196_, new_n201_ );
not g097 ( new_n203_, keyIn_0_31 );
not g098 ( new_n204_, keyIn_0_19 );
not g099 ( new_n205_, N21 );
and g100 ( new_n206_, new_n205_, N17 );
not g101 ( new_n207_, N17 );
and g102 ( new_n208_, new_n207_, N21 );
or g103 ( new_n209_, new_n206_, new_n208_ );
not g104 ( new_n210_, new_n209_ );
not g105 ( new_n211_, N29 );
and g106 ( new_n212_, new_n211_, N25 );
not g107 ( new_n213_, N25 );
and g108 ( new_n214_, new_n213_, N29 );
or g109 ( new_n215_, new_n212_, new_n214_ );
not g110 ( new_n216_, new_n215_ );
and g111 ( new_n217_, new_n210_, new_n216_ );
and g112 ( new_n218_, new_n209_, new_n215_ );
or g113 ( new_n219_, new_n217_, new_n218_ );
or g114 ( new_n220_, new_n219_, keyIn_0_1 );
and g115 ( new_n221_, new_n219_, keyIn_0_1 );
not g116 ( new_n222_, new_n221_ );
and g117 ( new_n223_, new_n222_, new_n220_ );
not g118 ( new_n224_, N53 );
and g119 ( new_n225_, new_n224_, N49 );
not g120 ( new_n226_, N49 );
and g121 ( new_n227_, new_n226_, N53 );
or g122 ( new_n228_, new_n225_, new_n227_ );
not g123 ( new_n229_, N61 );
and g124 ( new_n230_, new_n229_, N57 );
not g125 ( new_n231_, N57 );
and g126 ( new_n232_, new_n231_, N61 );
or g127 ( new_n233_, new_n230_, new_n232_ );
not g128 ( new_n234_, new_n233_ );
and g129 ( new_n235_, new_n234_, new_n228_ );
not g130 ( new_n236_, new_n228_ );
and g131 ( new_n237_, new_n236_, new_n233_ );
or g132 ( new_n238_, new_n235_, new_n237_ );
and g133 ( new_n239_, new_n238_, keyIn_0_3 );
not g134 ( new_n240_, keyIn_0_3 );
not g135 ( new_n241_, new_n235_ );
not g136 ( new_n242_, new_n237_ );
and g137 ( new_n243_, new_n241_, new_n242_ );
and g138 ( new_n244_, new_n243_, new_n240_ );
or g139 ( new_n245_, new_n244_, new_n239_ );
or g140 ( new_n246_, new_n245_, new_n223_ );
not g141 ( new_n247_, new_n220_ );
or g142 ( new_n248_, new_n247_, new_n221_ );
not g143 ( new_n249_, new_n239_ );
or g144 ( new_n250_, new_n238_, keyIn_0_3 );
and g145 ( new_n251_, new_n249_, new_n250_ );
or g146 ( new_n252_, new_n248_, new_n251_ );
and g147 ( new_n253_, new_n252_, new_n246_ );
or g148 ( new_n254_, new_n253_, new_n204_ );
and g149 ( new_n255_, new_n248_, new_n251_ );
and g150 ( new_n256_, new_n245_, new_n223_ );
or g151 ( new_n257_, new_n255_, new_n256_ );
or g152 ( new_n258_, new_n257_, keyIn_0_19 );
and g153 ( new_n259_, new_n258_, new_n254_ );
and g154 ( new_n260_, N136, N137 );
or g155 ( new_n261_, new_n259_, new_n260_ );
and g156 ( new_n262_, new_n257_, keyIn_0_19 );
and g157 ( new_n263_, new_n253_, new_n204_ );
or g158 ( new_n264_, new_n262_, new_n263_ );
not g159 ( new_n265_, new_n260_ );
or g160 ( new_n266_, new_n264_, new_n265_ );
and g161 ( new_n267_, new_n266_, new_n261_ );
or g162 ( new_n268_, new_n267_, new_n203_ );
and g163 ( new_n269_, new_n264_, new_n265_ );
and g164 ( new_n270_, new_n259_, new_n260_ );
or g165 ( new_n271_, new_n269_, new_n270_ );
or g166 ( new_n272_, new_n271_, keyIn_0_31 );
and g167 ( new_n273_, new_n272_, new_n268_ );
not g168 ( new_n274_, N125 );
and g169 ( new_n275_, new_n274_, N109 );
not g170 ( new_n276_, N109 );
and g171 ( new_n277_, new_n276_, N125 );
or g172 ( new_n278_, new_n275_, new_n277_ );
and g173 ( new_n279_, N77, N93 );
not g174 ( new_n280_, N77 );
not g175 ( new_n281_, N93 );
and g176 ( new_n282_, new_n280_, new_n281_ );
or g177 ( new_n283_, new_n282_, new_n279_ );
and g178 ( new_n284_, new_n278_, new_n283_ );
not g179 ( new_n285_, new_n284_ );
or g180 ( new_n286_, new_n278_, new_n283_ );
and g181 ( new_n287_, new_n285_, new_n286_ );
not g182 ( new_n288_, new_n287_ );
and g183 ( new_n289_, new_n288_, keyIn_0_15 );
not g184 ( new_n290_, new_n289_ );
or g185 ( new_n291_, new_n288_, keyIn_0_15 );
and g186 ( new_n292_, new_n290_, new_n291_ );
or g187 ( new_n293_, new_n273_, new_n292_ );
and g188 ( new_n294_, new_n271_, keyIn_0_31 );
and g189 ( new_n295_, new_n267_, new_n203_ );
or g190 ( new_n296_, new_n294_, new_n295_ );
not g191 ( new_n297_, new_n292_ );
or g192 ( new_n298_, new_n296_, new_n297_ );
and g193 ( new_n299_, new_n298_, new_n293_ );
and g194 ( new_n300_, new_n202_, new_n299_ );
not g195 ( new_n301_, keyIn_0_28 );
not g196 ( new_n302_, keyIn_0_16 );
and g197 ( new_n303_, new_n248_, new_n150_ );
and g198 ( new_n304_, new_n125_, new_n223_ );
or g199 ( new_n305_, new_n303_, new_n304_ );
and g200 ( new_n306_, new_n305_, new_n302_ );
not g201 ( new_n307_, new_n306_ );
or g202 ( new_n308_, new_n305_, new_n302_ );
and g203 ( new_n309_, new_n307_, new_n308_ );
and g204 ( new_n310_, N133, N137 );
not g205 ( new_n311_, new_n310_ );
and g206 ( new_n312_, new_n309_, new_n311_ );
not g207 ( new_n313_, new_n312_ );
or g208 ( new_n314_, new_n309_, new_n311_ );
and g209 ( new_n315_, new_n313_, new_n314_ );
or g210 ( new_n316_, new_n315_, new_n301_ );
not g211 ( new_n317_, new_n316_ );
and g212 ( new_n318_, new_n315_, new_n301_ );
or g213 ( new_n319_, new_n317_, new_n318_ );
not g214 ( new_n320_, keyIn_0_12 );
not g215 ( new_n321_, N113 );
and g216 ( new_n322_, new_n321_, N97 );
not g217 ( new_n323_, N97 );
and g218 ( new_n324_, new_n323_, N113 );
or g219 ( new_n325_, new_n322_, new_n324_ );
and g220 ( new_n326_, N65, N81 );
not g221 ( new_n327_, N65 );
not g222 ( new_n328_, N81 );
and g223 ( new_n329_, new_n327_, new_n328_ );
or g224 ( new_n330_, new_n329_, new_n326_ );
and g225 ( new_n331_, new_n325_, new_n330_ );
not g226 ( new_n332_, new_n331_ );
or g227 ( new_n333_, new_n325_, new_n330_ );
and g228 ( new_n334_, new_n332_, new_n333_ );
not g229 ( new_n335_, new_n334_ );
and g230 ( new_n336_, new_n335_, new_n320_ );
and g231 ( new_n337_, new_n334_, keyIn_0_12 );
or g232 ( new_n338_, new_n336_, new_n337_ );
and g233 ( new_n339_, new_n319_, new_n338_ );
not g234 ( new_n340_, new_n318_ );
and g235 ( new_n341_, new_n340_, new_n316_ );
not g236 ( new_n342_, new_n338_ );
and g237 ( new_n343_, new_n341_, new_n342_ );
or g238 ( new_n344_, new_n339_, new_n343_ );
not g239 ( new_n345_, keyIn_0_29 );
and g240 ( new_n346_, new_n144_, new_n245_ );
and g241 ( new_n347_, new_n251_, new_n152_ );
or g242 ( new_n348_, new_n346_, new_n347_ );
and g243 ( new_n349_, new_n348_, keyIn_0_17 );
not g244 ( new_n350_, new_n349_ );
or g245 ( new_n351_, new_n348_, keyIn_0_17 );
and g246 ( new_n352_, new_n350_, new_n351_ );
and g247 ( new_n353_, N134, N137 );
or g248 ( new_n354_, new_n352_, new_n353_ );
and g249 ( new_n355_, new_n352_, new_n353_ );
not g250 ( new_n356_, new_n355_ );
and g251 ( new_n357_, new_n356_, new_n354_ );
or g252 ( new_n358_, new_n357_, new_n345_ );
not g253 ( new_n359_, new_n358_ );
and g254 ( new_n360_, new_n357_, new_n345_ );
or g255 ( new_n361_, new_n359_, new_n360_ );
not g256 ( new_n362_, keyIn_0_13 );
not g257 ( new_n363_, N117 );
and g258 ( new_n364_, new_n363_, N101 );
not g259 ( new_n365_, N101 );
and g260 ( new_n366_, new_n365_, N117 );
or g261 ( new_n367_, new_n364_, new_n366_ );
and g262 ( new_n368_, N69, N85 );
not g263 ( new_n369_, N69 );
not g264 ( new_n370_, N85 );
and g265 ( new_n371_, new_n369_, new_n370_ );
or g266 ( new_n372_, new_n371_, new_n368_ );
and g267 ( new_n373_, new_n367_, new_n372_ );
not g268 ( new_n374_, new_n373_ );
or g269 ( new_n375_, new_n367_, new_n372_ );
and g270 ( new_n376_, new_n374_, new_n375_ );
not g271 ( new_n377_, new_n376_ );
and g272 ( new_n378_, new_n377_, new_n362_ );
and g273 ( new_n379_, new_n376_, keyIn_0_13 );
or g274 ( new_n380_, new_n378_, new_n379_ );
and g275 ( new_n381_, new_n361_, new_n380_ );
not g276 ( new_n382_, new_n360_ );
and g277 ( new_n383_, new_n382_, new_n358_ );
not g278 ( new_n384_, new_n380_ );
and g279 ( new_n385_, new_n383_, new_n384_ );
or g280 ( new_n386_, new_n381_, new_n385_ );
and g281 ( new_n387_, new_n344_, new_n386_ );
not g282 ( new_n388_, keyIn_0_23 );
not g283 ( new_n389_, keyIn_0_5 );
or g284 ( new_n390_, new_n328_, N85 );
or g285 ( new_n391_, new_n370_, N81 );
and g286 ( new_n392_, new_n390_, new_n391_ );
and g287 ( new_n393_, new_n281_, N89 );
and g288 ( new_n394_, new_n184_, N93 );
or g289 ( new_n395_, new_n393_, new_n394_ );
or g290 ( new_n396_, new_n395_, new_n392_ );
and g291 ( new_n397_, new_n370_, N81 );
and g292 ( new_n398_, new_n328_, N85 );
or g293 ( new_n399_, new_n397_, new_n398_ );
or g294 ( new_n400_, new_n184_, N93 );
or g295 ( new_n401_, new_n281_, N89 );
and g296 ( new_n402_, new_n400_, new_n401_ );
or g297 ( new_n403_, new_n399_, new_n402_ );
and g298 ( new_n404_, new_n396_, new_n403_ );
and g299 ( new_n405_, new_n404_, new_n389_ );
and g300 ( new_n406_, new_n399_, new_n402_ );
and g301 ( new_n407_, new_n395_, new_n392_ );
or g302 ( new_n408_, new_n406_, new_n407_ );
and g303 ( new_n409_, new_n408_, keyIn_0_5 );
or g304 ( new_n410_, new_n409_, new_n405_ );
or g305 ( new_n411_, new_n321_, N117 );
or g306 ( new_n412_, new_n363_, N113 );
and g307 ( new_n413_, new_n411_, new_n412_ );
or g308 ( new_n414_, new_n177_, N125 );
or g309 ( new_n415_, new_n274_, N121 );
and g310 ( new_n416_, new_n414_, new_n415_ );
and g311 ( new_n417_, new_n413_, new_n416_ );
and g312 ( new_n418_, new_n363_, N113 );
and g313 ( new_n419_, new_n321_, N117 );
or g314 ( new_n420_, new_n418_, new_n419_ );
and g315 ( new_n421_, new_n274_, N121 );
and g316 ( new_n422_, new_n177_, N125 );
or g317 ( new_n423_, new_n421_, new_n422_ );
and g318 ( new_n424_, new_n420_, new_n423_ );
or g319 ( new_n425_, new_n424_, new_n417_ );
or g320 ( new_n426_, new_n425_, keyIn_0_7 );
not g321 ( new_n427_, keyIn_0_7 );
or g322 ( new_n428_, new_n420_, new_n423_ );
or g323 ( new_n429_, new_n413_, new_n416_ );
and g324 ( new_n430_, new_n428_, new_n429_ );
or g325 ( new_n431_, new_n430_, new_n427_ );
and g326 ( new_n432_, new_n431_, new_n426_ );
or g327 ( new_n433_, new_n410_, new_n432_ );
or g328 ( new_n434_, new_n408_, keyIn_0_5 );
or g329 ( new_n435_, new_n404_, new_n389_ );
and g330 ( new_n436_, new_n434_, new_n435_ );
and g331 ( new_n437_, new_n430_, new_n427_ );
and g332 ( new_n438_, new_n425_, keyIn_0_7 );
or g333 ( new_n439_, new_n437_, new_n438_ );
or g334 ( new_n440_, new_n439_, new_n436_ );
and g335 ( new_n441_, new_n433_, new_n440_ );
or g336 ( new_n442_, new_n441_, new_n388_ );
and g337 ( new_n443_, new_n439_, new_n436_ );
and g338 ( new_n444_, new_n410_, new_n432_ );
or g339 ( new_n445_, new_n443_, new_n444_ );
or g340 ( new_n446_, new_n445_, keyIn_0_23 );
and g341 ( new_n447_, new_n446_, new_n442_ );
and g342 ( new_n448_, N132, N137 );
or g343 ( new_n449_, new_n447_, new_n448_ );
and g344 ( new_n450_, new_n445_, keyIn_0_23 );
and g345 ( new_n451_, new_n441_, new_n388_ );
or g346 ( new_n452_, new_n450_, new_n451_ );
not g347 ( new_n453_, new_n448_ );
or g348 ( new_n454_, new_n452_, new_n453_ );
and g349 ( new_n455_, new_n454_, new_n449_ );
or g350 ( new_n456_, new_n455_, keyIn_0_27 );
not g351 ( new_n457_, keyIn_0_27 );
and g352 ( new_n458_, new_n452_, new_n453_ );
and g353 ( new_n459_, new_n447_, new_n448_ );
or g354 ( new_n460_, new_n458_, new_n459_ );
or g355 ( new_n461_, new_n460_, new_n457_ );
and g356 ( new_n462_, new_n461_, new_n456_ );
not g357 ( new_n463_, keyIn_0_11 );
and g358 ( new_n464_, new_n229_, N45 );
and g359 ( new_n465_, new_n132_, N61 );
or g360 ( new_n466_, new_n464_, new_n465_ );
and g361 ( new_n467_, N13, N29 );
and g362 ( new_n468_, new_n112_, new_n211_ );
or g363 ( new_n469_, new_n468_, new_n467_ );
and g364 ( new_n470_, new_n466_, new_n469_ );
not g365 ( new_n471_, new_n470_ );
or g366 ( new_n472_, new_n466_, new_n469_ );
and g367 ( new_n473_, new_n471_, new_n472_ );
not g368 ( new_n474_, new_n473_ );
and g369 ( new_n475_, new_n474_, new_n463_ );
and g370 ( new_n476_, new_n473_, keyIn_0_11 );
or g371 ( new_n477_, new_n475_, new_n476_ );
not g372 ( new_n478_, new_n477_ );
or g373 ( new_n479_, new_n462_, new_n478_ );
and g374 ( new_n480_, new_n460_, new_n457_ );
and g375 ( new_n481_, new_n455_, keyIn_0_27 );
or g376 ( new_n482_, new_n480_, new_n481_ );
or g377 ( new_n483_, new_n482_, new_n477_ );
and g378 ( new_n484_, new_n483_, new_n479_ );
not g379 ( new_n485_, keyIn_0_24 );
or g380 ( new_n486_, new_n327_, N69 );
or g381 ( new_n487_, new_n369_, N65 );
and g382 ( new_n488_, new_n486_, new_n487_ );
and g383 ( new_n489_, new_n280_, N73 );
and g384 ( new_n490_, new_n183_, N77 );
or g385 ( new_n491_, new_n489_, new_n490_ );
or g386 ( new_n492_, new_n491_, new_n488_ );
and g387 ( new_n493_, new_n369_, N65 );
and g388 ( new_n494_, new_n327_, N69 );
or g389 ( new_n495_, new_n493_, new_n494_ );
or g390 ( new_n496_, new_n183_, N77 );
or g391 ( new_n497_, new_n280_, N73 );
and g392 ( new_n498_, new_n496_, new_n497_ );
or g393 ( new_n499_, new_n495_, new_n498_ );
and g394 ( new_n500_, new_n492_, new_n499_ );
or g395 ( new_n501_, new_n500_, keyIn_0_4 );
not g396 ( new_n502_, keyIn_0_4 );
and g397 ( new_n503_, new_n495_, new_n498_ );
and g398 ( new_n504_, new_n491_, new_n488_ );
or g399 ( new_n505_, new_n503_, new_n504_ );
or g400 ( new_n506_, new_n505_, new_n502_ );
and g401 ( new_n507_, new_n506_, new_n501_ );
or g402 ( new_n508_, new_n410_, new_n507_ );
and g403 ( new_n509_, new_n505_, new_n502_ );
and g404 ( new_n510_, new_n500_, keyIn_0_4 );
or g405 ( new_n511_, new_n509_, new_n510_ );
or g406 ( new_n512_, new_n511_, new_n436_ );
and g407 ( new_n513_, new_n508_, new_n512_ );
or g408 ( new_n514_, new_n513_, keyIn_0_20 );
not g409 ( new_n515_, keyIn_0_20 );
and g410 ( new_n516_, new_n511_, new_n436_ );
and g411 ( new_n517_, new_n410_, new_n507_ );
or g412 ( new_n518_, new_n516_, new_n517_ );
or g413 ( new_n519_, new_n518_, new_n515_ );
and g414 ( new_n520_, new_n519_, new_n514_ );
and g415 ( new_n521_, N129, N137 );
not g416 ( new_n522_, new_n521_ );
or g417 ( new_n523_, new_n520_, new_n522_ );
and g418 ( new_n524_, new_n518_, new_n515_ );
and g419 ( new_n525_, new_n513_, keyIn_0_20 );
or g420 ( new_n526_, new_n524_, new_n525_ );
or g421 ( new_n527_, new_n526_, new_n521_ );
and g422 ( new_n528_, new_n527_, new_n523_ );
or g423 ( new_n529_, new_n528_, new_n485_ );
and g424 ( new_n530_, new_n526_, new_n521_ );
and g425 ( new_n531_, new_n520_, new_n522_ );
or g426 ( new_n532_, new_n530_, new_n531_ );
or g427 ( new_n533_, new_n532_, keyIn_0_24 );
and g428 ( new_n534_, new_n533_, new_n529_ );
and g429 ( new_n535_, new_n226_, N33 );
and g430 ( new_n536_, new_n128_, N49 );
or g431 ( new_n537_, new_n535_, new_n536_ );
and g432 ( new_n538_, N1, N17 );
and g433 ( new_n539_, new_n109_, new_n207_ );
or g434 ( new_n540_, new_n539_, new_n538_ );
and g435 ( new_n541_, new_n537_, new_n540_ );
not g436 ( new_n542_, new_n541_ );
or g437 ( new_n543_, new_n537_, new_n540_ );
and g438 ( new_n544_, new_n542_, new_n543_ );
not g439 ( new_n545_, new_n544_ );
and g440 ( new_n546_, new_n545_, keyIn_0_8 );
not g441 ( new_n547_, new_n546_ );
or g442 ( new_n548_, new_n545_, keyIn_0_8 );
and g443 ( new_n549_, new_n547_, new_n548_ );
not g444 ( new_n550_, new_n549_ );
or g445 ( new_n551_, new_n534_, new_n550_ );
and g446 ( new_n552_, new_n532_, keyIn_0_24 );
and g447 ( new_n553_, new_n528_, new_n485_ );
or g448 ( new_n554_, new_n552_, new_n553_ );
or g449 ( new_n555_, new_n554_, new_n549_ );
and g450 ( new_n556_, new_n555_, new_n551_ );
not g451 ( new_n557_, new_n556_ );
and g452 ( new_n558_, new_n557_, new_n484_ );
not g453 ( new_n559_, keyIn_0_21 );
not g454 ( new_n560_, keyIn_0_6 );
and g455 ( new_n561_, new_n365_, N97 );
and g456 ( new_n562_, new_n323_, N101 );
or g457 ( new_n563_, new_n561_, new_n562_ );
not g458 ( new_n564_, new_n563_ );
and g459 ( new_n565_, new_n276_, N105 );
and g460 ( new_n566_, new_n179_, N109 );
or g461 ( new_n567_, new_n565_, new_n566_ );
not g462 ( new_n568_, new_n567_ );
and g463 ( new_n569_, new_n564_, new_n568_ );
and g464 ( new_n570_, new_n563_, new_n567_ );
or g465 ( new_n571_, new_n569_, new_n570_ );
or g466 ( new_n572_, new_n571_, new_n560_ );
and g467 ( new_n573_, new_n571_, new_n560_ );
not g468 ( new_n574_, new_n573_ );
and g469 ( new_n575_, new_n574_, new_n572_ );
or g470 ( new_n576_, new_n575_, new_n432_ );
and g471 ( new_n577_, new_n575_, new_n432_ );
not g472 ( new_n578_, new_n577_ );
and g473 ( new_n579_, new_n578_, new_n576_ );
or g474 ( new_n580_, new_n579_, new_n559_ );
not g475 ( new_n581_, new_n572_ );
or g476 ( new_n582_, new_n581_, new_n573_ );
and g477 ( new_n583_, new_n582_, new_n439_ );
or g478 ( new_n584_, new_n583_, new_n577_ );
or g479 ( new_n585_, new_n584_, keyIn_0_21 );
and g480 ( new_n586_, new_n580_, new_n585_ );
and g481 ( new_n587_, N130, N137 );
or g482 ( new_n588_, new_n586_, new_n587_ );
and g483 ( new_n589_, new_n584_, keyIn_0_21 );
and g484 ( new_n590_, new_n579_, new_n559_ );
or g485 ( new_n591_, new_n590_, new_n589_ );
not g486 ( new_n592_, new_n587_ );
or g487 ( new_n593_, new_n591_, new_n592_ );
and g488 ( new_n594_, new_n593_, new_n588_ );
or g489 ( new_n595_, new_n594_, keyIn_0_25 );
not g490 ( new_n596_, keyIn_0_25 );
and g491 ( new_n597_, new_n591_, new_n592_ );
and g492 ( new_n598_, new_n586_, new_n587_ );
or g493 ( new_n599_, new_n597_, new_n598_ );
or g494 ( new_n600_, new_n599_, new_n596_ );
and g495 ( new_n601_, new_n600_, new_n595_ );
not g496 ( new_n602_, keyIn_0_9 );
and g497 ( new_n603_, new_n224_, N37 );
and g498 ( new_n604_, new_n126_, N53 );
or g499 ( new_n605_, new_n603_, new_n604_ );
and g500 ( new_n606_, N5, N21 );
and g501 ( new_n607_, new_n107_, new_n205_ );
or g502 ( new_n608_, new_n607_, new_n606_ );
and g503 ( new_n609_, new_n605_, new_n608_ );
not g504 ( new_n610_, new_n609_ );
or g505 ( new_n611_, new_n605_, new_n608_ );
and g506 ( new_n612_, new_n610_, new_n611_ );
not g507 ( new_n613_, new_n612_ );
and g508 ( new_n614_, new_n613_, new_n602_ );
and g509 ( new_n615_, new_n612_, keyIn_0_9 );
or g510 ( new_n616_, new_n614_, new_n615_ );
or g511 ( new_n617_, new_n601_, new_n616_ );
and g512 ( new_n618_, new_n599_, new_n596_ );
and g513 ( new_n619_, new_n594_, keyIn_0_25 );
or g514 ( new_n620_, new_n618_, new_n619_ );
not g515 ( new_n621_, new_n616_ );
or g516 ( new_n622_, new_n620_, new_n621_ );
and g517 ( new_n623_, new_n622_, new_n617_ );
not g518 ( new_n624_, keyIn_0_26 );
or g519 ( new_n625_, new_n575_, new_n507_ );
and g520 ( new_n626_, new_n575_, new_n507_ );
not g521 ( new_n627_, new_n626_ );
and g522 ( new_n628_, new_n627_, new_n625_ );
or g523 ( new_n629_, new_n628_, keyIn_0_22 );
not g524 ( new_n630_, keyIn_0_22 );
and g525 ( new_n631_, new_n582_, new_n511_ );
or g526 ( new_n632_, new_n631_, new_n626_ );
or g527 ( new_n633_, new_n632_, new_n630_ );
and g528 ( new_n634_, new_n629_, new_n633_ );
and g529 ( new_n635_, N131, N137 );
not g530 ( new_n636_, new_n635_ );
or g531 ( new_n637_, new_n634_, new_n636_ );
and g532 ( new_n638_, new_n632_, new_n630_ );
and g533 ( new_n639_, new_n628_, keyIn_0_22 );
or g534 ( new_n640_, new_n639_, new_n638_ );
or g535 ( new_n641_, new_n640_, new_n635_ );
and g536 ( new_n642_, new_n641_, new_n637_ );
or g537 ( new_n643_, new_n642_, new_n624_ );
and g538 ( new_n644_, new_n640_, new_n635_ );
and g539 ( new_n645_, new_n634_, new_n636_ );
or g540 ( new_n646_, new_n644_, new_n645_ );
or g541 ( new_n647_, new_n646_, keyIn_0_26 );
and g542 ( new_n648_, new_n647_, new_n643_ );
and g543 ( new_n649_, new_n231_, N41 );
and g544 ( new_n650_, new_n134_, N57 );
or g545 ( new_n651_, new_n649_, new_n650_ );
and g546 ( new_n652_, N9, N25 );
and g547 ( new_n653_, new_n114_, new_n213_ );
or g548 ( new_n654_, new_n653_, new_n652_ );
and g549 ( new_n655_, new_n651_, new_n654_ );
not g550 ( new_n656_, new_n655_ );
or g551 ( new_n657_, new_n651_, new_n654_ );
and g552 ( new_n658_, new_n656_, new_n657_ );
not g553 ( new_n659_, new_n658_ );
and g554 ( new_n660_, new_n659_, keyIn_0_10 );
not g555 ( new_n661_, new_n660_ );
or g556 ( new_n662_, new_n659_, keyIn_0_10 );
and g557 ( new_n663_, new_n661_, new_n662_ );
or g558 ( new_n664_, new_n648_, new_n663_ );
and g559 ( new_n665_, new_n646_, keyIn_0_26 );
and g560 ( new_n666_, new_n642_, new_n624_ );
or g561 ( new_n667_, new_n665_, new_n666_ );
not g562 ( new_n668_, new_n663_ );
or g563 ( new_n669_, new_n667_, new_n668_ );
and g564 ( new_n670_, new_n669_, new_n664_ );
and g565 ( new_n671_, new_n623_, new_n670_ );
and g566 ( new_n672_, new_n671_, new_n558_ );
and g567 ( new_n673_, new_n387_, new_n672_ );
and g568 ( new_n674_, new_n673_, new_n300_ );
not g569 ( new_n675_, new_n674_ );
and g570 ( new_n676_, new_n675_, N1 );
and g571 ( new_n677_, new_n674_, new_n109_ );
or g572 ( N724, new_n676_, new_n677_ );
and g573 ( new_n679_, new_n620_, new_n621_ );
and g574 ( new_n680_, new_n601_, new_n616_ );
or g575 ( new_n681_, new_n679_, new_n680_ );
and g576 ( new_n682_, new_n484_, new_n556_ );
and g577 ( new_n683_, new_n682_, new_n681_ );
and g578 ( new_n684_, new_n683_, new_n670_ );
and g579 ( new_n685_, new_n684_, new_n387_ );
and g580 ( new_n686_, new_n685_, new_n300_ );
not g581 ( new_n687_, new_n686_ );
and g582 ( new_n688_, new_n687_, N5 );
and g583 ( new_n689_, new_n686_, new_n107_ );
or g584 ( N725, new_n688_, new_n689_ );
and g585 ( new_n691_, new_n667_, new_n668_ );
and g586 ( new_n692_, new_n648_, new_n663_ );
or g587 ( new_n693_, new_n691_, new_n692_ );
and g588 ( new_n694_, new_n693_, new_n623_ );
and g589 ( new_n695_, new_n694_, new_n682_ );
and g590 ( new_n696_, new_n387_, new_n695_ );
and g591 ( new_n697_, new_n696_, new_n300_ );
not g592 ( new_n698_, new_n697_ );
and g593 ( new_n699_, new_n698_, N9 );
and g594 ( new_n700_, new_n697_, new_n114_ );
or g595 ( N726, new_n699_, new_n700_ );
not g596 ( new_n702_, new_n484_ );
and g597 ( new_n703_, new_n702_, new_n556_ );
and g598 ( new_n704_, new_n703_, new_n670_ );
and g599 ( new_n705_, new_n387_, new_n704_ );
and g600 ( new_n706_, new_n300_, new_n623_ );
and g601 ( new_n707_, new_n705_, new_n706_ );
not g602 ( new_n708_, new_n707_ );
and g603 ( new_n709_, new_n708_, N13 );
and g604 ( new_n710_, new_n704_, new_n623_ );
and g605 ( new_n711_, new_n300_, new_n112_ );
and g606 ( new_n712_, new_n387_, new_n711_ );
and g607 ( new_n713_, new_n712_, new_n710_ );
or g608 ( N727, new_n709_, new_n713_ );
or g609 ( new_n715_, new_n199_, new_n200_ );
or g610 ( new_n716_, new_n176_, new_n195_ );
and g611 ( new_n717_, new_n716_, new_n715_ );
and g612 ( new_n718_, new_n296_, new_n297_ );
and g613 ( new_n719_, new_n273_, new_n292_ );
or g614 ( new_n720_, new_n718_, new_n719_ );
and g615 ( new_n721_, new_n720_, new_n717_ );
and g616 ( new_n722_, new_n673_, new_n721_ );
not g617 ( new_n723_, new_n722_ );
and g618 ( new_n724_, new_n723_, N17 );
and g619 ( new_n725_, new_n722_, new_n207_ );
or g620 ( N728, new_n724_, new_n725_ );
and g621 ( new_n727_, new_n685_, new_n721_ );
not g622 ( new_n728_, new_n727_ );
and g623 ( new_n729_, new_n728_, N21 );
and g624 ( new_n730_, new_n727_, new_n205_ );
or g625 ( N729, new_n729_, new_n730_ );
and g626 ( new_n732_, new_n696_, new_n721_ );
not g627 ( new_n733_, new_n732_ );
and g628 ( new_n734_, new_n733_, N25 );
and g629 ( new_n735_, new_n732_, new_n213_ );
or g630 ( N730, new_n734_, new_n735_ );
and g631 ( new_n737_, new_n721_, new_n623_ );
and g632 ( new_n738_, new_n705_, new_n737_ );
not g633 ( new_n739_, new_n738_ );
and g634 ( new_n740_, new_n739_, N29 );
and g635 ( new_n741_, new_n387_, new_n211_ );
and g636 ( new_n742_, new_n741_, new_n721_ );
and g637 ( new_n743_, new_n742_, new_n710_ );
or g638 ( N731, new_n740_, new_n743_ );
or g639 ( new_n745_, new_n341_, new_n342_ );
or g640 ( new_n746_, new_n319_, new_n338_ );
and g641 ( new_n747_, new_n746_, new_n745_ );
and g642 ( new_n748_, new_n747_, new_n300_ );
or g643 ( new_n749_, new_n383_, new_n384_ );
or g644 ( new_n750_, new_n361_, new_n380_ );
and g645 ( new_n751_, new_n750_, new_n749_ );
and g646 ( new_n752_, new_n672_, new_n751_ );
and g647 ( new_n753_, new_n752_, new_n748_ );
not g648 ( new_n754_, new_n753_ );
and g649 ( new_n755_, new_n754_, N33 );
and g650 ( new_n756_, new_n753_, new_n128_ );
or g651 ( N732, new_n755_, new_n756_ );
and g652 ( new_n758_, new_n748_, new_n751_ );
and g653 ( new_n759_, new_n758_, new_n684_ );
not g654 ( new_n760_, new_n759_ );
and g655 ( new_n761_, new_n760_, N37 );
and g656 ( new_n762_, new_n759_, new_n126_ );
or g657 ( N733, new_n761_, new_n762_ );
and g658 ( new_n764_, new_n758_, new_n695_ );
not g659 ( new_n765_, new_n764_ );
and g660 ( new_n766_, new_n765_, N41 );
and g661 ( new_n767_, new_n764_, new_n134_ );
or g662 ( N734, new_n766_, new_n767_ );
and g663 ( new_n769_, new_n758_, new_n710_ );
not g664 ( new_n770_, new_n769_ );
and g665 ( new_n771_, new_n770_, N45 );
and g666 ( new_n772_, new_n769_, new_n132_ );
or g667 ( N735, new_n771_, new_n772_ );
and g668 ( new_n774_, new_n747_, new_n721_ );
and g669 ( new_n775_, new_n752_, new_n774_ );
not g670 ( new_n776_, new_n775_ );
and g671 ( new_n777_, new_n776_, N49 );
and g672 ( new_n778_, new_n775_, new_n226_ );
or g673 ( N736, new_n777_, new_n778_ );
and g674 ( new_n780_, new_n774_, new_n751_ );
and g675 ( new_n781_, new_n780_, new_n684_ );
not g676 ( new_n782_, new_n781_ );
and g677 ( new_n783_, new_n782_, N53 );
and g678 ( new_n784_, new_n781_, new_n224_ );
or g679 ( N737, new_n783_, new_n784_ );
and g680 ( new_n786_, new_n780_, new_n695_ );
not g681 ( new_n787_, new_n786_ );
and g682 ( new_n788_, new_n787_, N57 );
and g683 ( new_n789_, new_n786_, new_n231_ );
or g684 ( N738, new_n788_, new_n789_ );
and g685 ( new_n791_, new_n780_, new_n710_ );
not g686 ( new_n792_, new_n791_ );
and g687 ( new_n793_, new_n792_, N61 );
and g688 ( new_n794_, new_n791_, new_n229_ );
or g689 ( N739, new_n793_, new_n794_ );
and g690 ( new_n796_, new_n717_, new_n299_ );
and g691 ( new_n797_, new_n387_, new_n796_ );
and g692 ( new_n798_, new_n694_, new_n558_ );
and g693 ( new_n799_, new_n797_, new_n798_ );
not g694 ( new_n800_, new_n799_ );
and g695 ( new_n801_, new_n800_, N65 );
and g696 ( new_n802_, new_n799_, new_n327_ );
or g697 ( N740, new_n801_, new_n802_ );
and g698 ( new_n804_, new_n747_, new_n751_ );
and g699 ( new_n805_, new_n804_, new_n796_ );
and g700 ( new_n806_, new_n805_, new_n798_ );
not g701 ( new_n807_, new_n806_ );
and g702 ( new_n808_, new_n807_, N69 );
and g703 ( new_n809_, new_n806_, new_n369_ );
or g704 ( N741, new_n808_, new_n809_ );
and g705 ( new_n811_, new_n748_, new_n386_ );
and g706 ( new_n812_, new_n811_, new_n798_ );
not g707 ( new_n813_, new_n812_ );
and g708 ( new_n814_, new_n813_, N73 );
and g709 ( new_n815_, new_n812_, new_n183_ );
or g710 ( N742, new_n814_, new_n815_ );
and g711 ( new_n817_, new_n774_, new_n386_ );
and g712 ( new_n818_, new_n817_, new_n798_ );
not g713 ( new_n819_, new_n818_ );
and g714 ( new_n820_, new_n819_, N77 );
and g715 ( new_n821_, new_n818_, new_n280_ );
or g716 ( N743, new_n820_, new_n821_ );
and g717 ( new_n823_, new_n702_, new_n557_ );
and g718 ( new_n824_, new_n671_, new_n823_ );
and g719 ( new_n825_, new_n797_, new_n824_ );
not g720 ( new_n826_, new_n825_ );
and g721 ( new_n827_, new_n826_, N81 );
and g722 ( new_n828_, new_n825_, new_n328_ );
or g723 ( N744, new_n827_, new_n828_ );
and g724 ( new_n830_, new_n805_, new_n824_ );
not g725 ( new_n831_, new_n830_ );
and g726 ( new_n832_, new_n831_, N85 );
and g727 ( new_n833_, new_n830_, new_n370_ );
or g728 ( N745, new_n832_, new_n833_ );
and g729 ( new_n835_, new_n811_, new_n824_ );
not g730 ( new_n836_, new_n835_ );
and g731 ( new_n837_, new_n836_, N89 );
and g732 ( new_n838_, new_n835_, new_n184_ );
or g733 ( N746, new_n837_, new_n838_ );
and g734 ( new_n840_, new_n817_, new_n824_ );
not g735 ( new_n841_, new_n840_ );
and g736 ( new_n842_, new_n841_, N93 );
and g737 ( new_n843_, new_n840_, new_n281_ );
or g738 ( N747, new_n842_, new_n843_ );
and g739 ( new_n845_, new_n683_, new_n693_ );
and g740 ( new_n846_, new_n797_, new_n845_ );
not g741 ( new_n847_, new_n846_ );
and g742 ( new_n848_, new_n847_, N97 );
and g743 ( new_n849_, new_n846_, new_n323_ );
or g744 ( N748, new_n848_, new_n849_ );
and g745 ( new_n851_, new_n805_, new_n845_ );
not g746 ( new_n852_, new_n851_ );
and g747 ( new_n853_, new_n852_, N101 );
and g748 ( new_n854_, new_n851_, new_n365_ );
or g749 ( N749, new_n853_, new_n854_ );
and g750 ( new_n856_, new_n811_, new_n845_ );
not g751 ( new_n857_, new_n856_ );
and g752 ( new_n858_, new_n857_, N105 );
and g753 ( new_n859_, new_n856_, new_n179_ );
or g754 ( N750, new_n858_, new_n859_ );
and g755 ( new_n861_, new_n817_, new_n845_ );
not g756 ( new_n862_, new_n861_ );
and g757 ( new_n863_, new_n862_, N109 );
and g758 ( new_n864_, new_n861_, new_n276_ );
or g759 ( N751, new_n863_, new_n864_ );
and g760 ( new_n866_, new_n704_, new_n681_ );
and g761 ( new_n867_, new_n797_, new_n866_ );
not g762 ( new_n868_, new_n867_ );
and g763 ( new_n869_, new_n868_, N113 );
and g764 ( new_n870_, new_n867_, new_n321_ );
or g765 ( N752, new_n869_, new_n870_ );
and g766 ( new_n872_, new_n805_, new_n866_ );
not g767 ( new_n873_, new_n872_ );
and g768 ( new_n874_, new_n873_, N117 );
and g769 ( new_n875_, new_n872_, new_n363_ );
or g770 ( N753, new_n874_, new_n875_ );
and g771 ( new_n877_, new_n811_, new_n866_ );
not g772 ( new_n878_, new_n877_ );
and g773 ( new_n879_, new_n878_, N121 );
and g774 ( new_n880_, new_n877_, new_n177_ );
or g775 ( N754, new_n879_, new_n880_ );
and g776 ( new_n882_, new_n817_, new_n866_ );
not g777 ( new_n883_, new_n882_ );
and g778 ( new_n884_, new_n883_, N125 );
and g779 ( new_n885_, new_n882_, new_n274_ );
or g780 ( N755, new_n884_, new_n885_ );
endmodule