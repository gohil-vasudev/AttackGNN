module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n236_, new_n976_, new_n238_, new_n479_, new_n955_, new_n608_, new_n847_, new_n250_, new_n888_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n246_, new_n682_, new_n812_, new_n911_, new_n679_, new_n937_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n188_, new_n695_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n500_, new_n898_, new_n786_, new_n799_, new_n946_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n862_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n959_, new_n774_, new_n157_, new_n716_, new_n701_, new_n792_, new_n953_, new_n257_, new_n481_, new_n212_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n634_, new_n192_, new_n414_, new_n635_, new_n315_, new_n326_, new_n554_, new_n648_, new_n903_, new_n164_, new_n230_, new_n983_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n849_, new_n606_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n167_, new_n385_, new_n829_, new_n478_, new_n694_, new_n461_, new_n971_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n683_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n966_, new_n351_, new_n517_, new_n325_, new_n609_, new_n961_, new_n530_, new_n890_, new_n318_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n956_, new_n763_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n970_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n650_, new_n708_, new_n750_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n734_, new_n912_, new_n925_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n256_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n820_, new_n771_, new_n388_, new_n979_, new_n508_, new_n714_, new_n483_, new_n394_, new_n299_, new_n935_, new_n657_, new_n929_, new_n314_, new_n582_, new_n363_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n917_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n207_, new_n267_, new_n473_, new_n790_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n969_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n621_, new_n846_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n874_, new_n943_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n939_, new_n208_, new_n632_, new_n671_, new_n965_, new_n528_, new_n952_, new_n179_, new_n572_, new_n850_, new_n436_, new_n397_, new_n729_, new_n975_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n559_, new_n948_, new_n762_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n794_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n276_, new_n688_, new_n155_, new_n384_, new_n900_, new_n410_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n860_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n938_, new_n809_, new_n654_, new_n713_, new_n880_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n967_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n749_, new_n861_, new_n310_, new_n275_, new_n352_, new_n931_, new_n575_, new_n839_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n493_, new_n547_, new_n907_, new_n264_, new_n665_, new_n800_, new_n379_, new_n897_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n963_, new_n270_, new_n570_, new_n598_, new_n893_, new_n824_, new_n520_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n557_, new_n260_, new_n936_, new_n251_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n748_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n879_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n231_, new_n219_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n428_, new_n916_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n919_, new_n302_, new_n191_, new_n755_, new_n225_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n977_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n968_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n972_, new_n891_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n593_, new_n974_, new_n252_, new_n585_, new_n751_, new_n312_, new_n535_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n190_, new_n597_, new_n978_, new_n408_, new_n470_, new_n213_, new_n769_, new_n651_, new_n433_, new_n871_, new_n435_, new_n776_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n957_, new_n754_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n330_, new_n727_, new_n375_, new_n962_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n357_, new_n320_, new_n780_, new_n984_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n865_, new_n358_, new_n877_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n896_, new_n802_, new_n697_, new_n185_, new_n951_, new_n709_, new_n373_, new_n866_, new_n171_, new_n540_, new_n434_, new_n200_, new_n947_, new_n982_, new_n422_, new_n964_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n551_, new_n168_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n521_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n573_, new_n765_, new_n405_;

not g000 ( new_n151_, N75 );
nand g001 ( new_n152_, N29, N42 );
nor g002 ( N388, new_n152_, new_n151_ );
not g003 ( new_n154_, N80 );
nand g004 ( new_n155_, N29, N36 );
nor g005 ( N389, new_n155_, new_n154_ );
not g006 ( new_n157_, N42 );
nor g007 ( N390, new_n155_, new_n157_ );
nand g008 ( new_n159_, N85, N86 );
not g009 ( N391, new_n159_ );
not g010 ( new_n161_, N17 );
nand g011 ( new_n162_, N1, N8 );
not g012 ( new_n163_, new_n162_ );
nand g013 ( new_n164_, new_n163_, N13 );
nor g014 ( N418, new_n164_, new_n161_ );
not g015 ( new_n166_, N390 );
nand g016 ( new_n167_, N1, N26 );
nand g017 ( new_n168_, N13, N17 );
nor g018 ( new_n169_, new_n167_, new_n168_ );
nand g019 ( N419, new_n166_, new_n169_ );
nand g020 ( new_n171_, N59, N75 );
not g021 ( new_n172_, new_n171_ );
nand g022 ( N420, new_n172_, N80 );
nand g023 ( new_n174_, N36, N59 );
not g024 ( new_n175_, new_n174_ );
nand g025 ( N421, new_n175_, N80 );
nand g026 ( N422, new_n175_, N42 );
not g027 ( new_n178_, N90 );
nor g028 ( new_n179_, N87, N88 );
nor g029 ( N423, new_n179_, new_n178_ );
nand g030 ( N446, new_n169_, N390 );
not g031 ( new_n182_, keyIn_0_0 );
not g032 ( new_n183_, N51 );
nor g033 ( new_n184_, new_n167_, new_n183_ );
nor g034 ( new_n185_, new_n184_, new_n182_ );
not g035 ( new_n186_, new_n167_ );
nand g036 ( new_n187_, new_n186_, N51 );
nor g037 ( new_n188_, new_n187_, keyIn_0_0 );
nor g038 ( N447, new_n188_, new_n185_ );
not g039 ( new_n190_, N55 );
nor g040 ( new_n191_, new_n164_, new_n190_ );
not g041 ( new_n192_, new_n191_ );
nand g042 ( new_n193_, N29, N68 );
nor g043 ( N448, new_n192_, new_n193_ );
not g044 ( new_n195_, N74 );
nand g045 ( new_n196_, N59, N68 );
nor g046 ( new_n197_, new_n192_, new_n196_ );
not g047 ( new_n198_, new_n197_ );
nor g048 ( N449, new_n198_, new_n195_ );
not g049 ( new_n200_, N89 );
nor g050 ( N450, new_n179_, new_n200_ );
nand g051 ( new_n202_, N111, N116 );
not g052 ( new_n203_, new_n202_ );
nor g053 ( new_n204_, N111, N116 );
nor g054 ( new_n205_, new_n203_, new_n204_ );
nand g055 ( new_n206_, N121, N126 );
not g056 ( new_n207_, new_n206_ );
nor g057 ( new_n208_, N121, N126 );
nor g058 ( new_n209_, new_n207_, new_n208_ );
nor g059 ( new_n210_, new_n205_, new_n209_ );
nand g060 ( new_n211_, new_n205_, new_n209_ );
not g061 ( new_n212_, new_n211_ );
nor g062 ( new_n213_, new_n212_, new_n210_ );
not g063 ( new_n214_, new_n213_ );
nand g064 ( new_n215_, new_n214_, N135 );
not g065 ( new_n216_, new_n215_ );
nor g066 ( new_n217_, new_n214_, N135 );
nor g067 ( new_n218_, new_n216_, new_n217_ );
not g068 ( new_n219_, new_n218_ );
not g069 ( new_n220_, N130 );
nand g070 ( new_n221_, N91, N96 );
not g071 ( new_n222_, new_n221_ );
nor g072 ( new_n223_, N91, N96 );
nor g073 ( new_n224_, new_n222_, new_n223_ );
nand g074 ( new_n225_, N101, N106 );
not g075 ( new_n226_, new_n225_ );
nor g076 ( new_n227_, N101, N106 );
nor g077 ( new_n228_, new_n226_, new_n227_ );
nor g078 ( new_n229_, new_n224_, new_n228_ );
nand g079 ( new_n230_, new_n224_, new_n228_ );
not g080 ( new_n231_, new_n230_ );
nor g081 ( new_n232_, new_n231_, new_n229_ );
not g082 ( new_n233_, new_n232_ );
nand g083 ( new_n234_, new_n233_, new_n220_ );
not g084 ( new_n235_, new_n234_ );
nor g085 ( new_n236_, new_n233_, new_n220_ );
nor g086 ( new_n237_, new_n235_, new_n236_ );
not g087 ( new_n238_, new_n237_ );
nand g088 ( new_n239_, new_n219_, new_n238_ );
nand g089 ( new_n240_, new_n218_, new_n237_ );
nand g090 ( N767, new_n239_, new_n240_ );
nand g091 ( new_n242_, N183, N189 );
not g092 ( new_n243_, new_n242_ );
nor g093 ( new_n244_, N183, N189 );
nor g094 ( new_n245_, new_n243_, new_n244_ );
nand g095 ( new_n246_, N195, N201 );
not g096 ( new_n247_, new_n246_ );
nor g097 ( new_n248_, N195, N201 );
nor g098 ( new_n249_, new_n247_, new_n248_ );
nor g099 ( new_n250_, new_n245_, new_n249_ );
nand g100 ( new_n251_, new_n245_, new_n249_ );
not g101 ( new_n252_, new_n251_ );
nor g102 ( new_n253_, new_n252_, new_n250_ );
not g103 ( new_n254_, new_n253_ );
nand g104 ( new_n255_, new_n254_, N207 );
not g105 ( new_n256_, new_n255_ );
nor g106 ( new_n257_, new_n254_, N207 );
nor g107 ( new_n258_, new_n256_, new_n257_ );
not g108 ( new_n259_, new_n258_ );
nand g109 ( new_n260_, N159, N165 );
not g110 ( new_n261_, new_n260_ );
nor g111 ( new_n262_, N159, N165 );
nor g112 ( new_n263_, new_n261_, new_n262_ );
nand g113 ( new_n264_, N171, N177 );
not g114 ( new_n265_, new_n264_ );
nor g115 ( new_n266_, N171, N177 );
nor g116 ( new_n267_, new_n265_, new_n266_ );
nor g117 ( new_n268_, new_n263_, new_n267_ );
nand g118 ( new_n269_, new_n263_, new_n267_ );
not g119 ( new_n270_, new_n269_ );
nor g120 ( new_n271_, new_n270_, new_n268_ );
not g121 ( new_n272_, new_n271_ );
nand g122 ( new_n273_, new_n272_, new_n220_ );
not g123 ( new_n274_, new_n273_ );
nor g124 ( new_n275_, new_n272_, new_n220_ );
nor g125 ( new_n276_, new_n274_, new_n275_ );
not g126 ( new_n277_, new_n276_ );
nand g127 ( new_n278_, new_n259_, new_n277_ );
nand g128 ( new_n279_, new_n258_, new_n276_ );
nand g129 ( N768, new_n278_, new_n279_ );
not g130 ( new_n281_, N261 );
not g131 ( new_n282_, keyIn_0_43 );
not g132 ( new_n283_, keyIn_0_31 );
not g133 ( new_n284_, keyIn_0_21 );
not g134 ( new_n285_, keyIn_0_19 );
nor g135 ( new_n286_, N447, keyIn_0_8 );
not g136 ( new_n287_, keyIn_0_8 );
nand g137 ( new_n288_, new_n187_, keyIn_0_0 );
nand g138 ( new_n289_, new_n184_, new_n182_ );
nand g139 ( new_n290_, new_n288_, new_n289_ );
nor g140 ( new_n291_, new_n290_, new_n287_ );
nor g141 ( new_n292_, new_n286_, new_n291_ );
nor g142 ( new_n293_, new_n292_, keyIn_0_14 );
not g143 ( new_n294_, keyIn_0_14 );
nand g144 ( new_n295_, new_n290_, new_n287_ );
nand g145 ( new_n296_, N447, keyIn_0_8 );
nand g146 ( new_n297_, new_n296_, new_n295_ );
nor g147 ( new_n298_, new_n297_, new_n294_ );
nor g148 ( new_n299_, new_n293_, new_n298_ );
not g149 ( new_n300_, keyIn_0_13 );
nor g150 ( new_n301_, N17, N42 );
nor g151 ( new_n302_, new_n301_, keyIn_0_6 );
not g152 ( new_n303_, new_n302_ );
nand g153 ( new_n304_, new_n301_, keyIn_0_6 );
nand g154 ( new_n305_, new_n303_, new_n304_ );
nand g155 ( new_n306_, N17, N42 );
nand g156 ( new_n307_, new_n306_, keyIn_0_7 );
nor g157 ( new_n308_, new_n306_, keyIn_0_7 );
not g158 ( new_n309_, new_n308_ );
nand g159 ( new_n310_, new_n309_, new_n307_ );
nand g160 ( new_n311_, new_n305_, new_n310_ );
nor g161 ( new_n312_, new_n311_, new_n300_ );
nand g162 ( new_n313_, N59, N156 );
not g163 ( new_n314_, new_n313_ );
nand g164 ( new_n315_, new_n311_, new_n300_ );
nand g165 ( new_n316_, new_n315_, new_n314_ );
nor g166 ( new_n317_, new_n316_, new_n312_ );
nand g167 ( new_n318_, new_n299_, new_n317_ );
nor g168 ( new_n319_, new_n318_, new_n285_ );
not g169 ( new_n320_, new_n319_ );
nand g170 ( new_n321_, N42, N59 );
nor g171 ( new_n322_, new_n321_, new_n151_ );
nor g172 ( new_n323_, new_n322_, keyIn_0_3 );
not g173 ( new_n324_, new_n323_ );
nand g174 ( new_n325_, new_n322_, keyIn_0_3 );
nand g175 ( new_n326_, new_n324_, new_n325_ );
nand g176 ( new_n327_, new_n326_, keyIn_0_11 );
not g177 ( new_n328_, keyIn_0_11 );
not g178 ( new_n329_, new_n325_ );
nor g179 ( new_n330_, new_n329_, new_n323_ );
nand g180 ( new_n331_, new_n330_, new_n328_ );
nand g181 ( new_n332_, new_n331_, new_n327_ );
not g182 ( new_n333_, keyIn_0_1 );
nand g183 ( new_n334_, N17, N51 );
nor g184 ( new_n335_, new_n162_, new_n334_ );
nor g185 ( new_n336_, new_n335_, new_n333_ );
nand g186 ( new_n337_, new_n335_, new_n333_ );
not g187 ( new_n338_, new_n337_ );
nor g188 ( new_n339_, new_n338_, new_n336_ );
nand g189 ( new_n340_, new_n162_, keyIn_0_1 );
nand g190 ( new_n341_, new_n340_, keyIn_0_9 );
not g191 ( new_n342_, new_n341_ );
nand g192 ( new_n343_, new_n339_, new_n342_ );
not g193 ( new_n344_, keyIn_0_9 );
not g194 ( new_n345_, new_n336_ );
nand g195 ( new_n346_, new_n345_, new_n337_ );
nand g196 ( new_n347_, new_n346_, new_n344_ );
nand g197 ( new_n348_, new_n343_, new_n347_ );
nand g198 ( new_n349_, new_n348_, new_n332_ );
nand g199 ( new_n350_, new_n349_, keyIn_0_15 );
not g200 ( new_n351_, new_n350_ );
nor g201 ( new_n352_, new_n349_, keyIn_0_15 );
nor g202 ( new_n353_, new_n351_, new_n352_ );
nand g203 ( new_n354_, new_n297_, new_n294_ );
nand g204 ( new_n355_, new_n292_, keyIn_0_14 );
nand g205 ( new_n356_, new_n355_, new_n354_ );
not g206 ( new_n357_, new_n317_ );
nor g207 ( new_n358_, new_n356_, new_n357_ );
nor g208 ( new_n359_, new_n358_, keyIn_0_19 );
nor g209 ( new_n360_, new_n359_, new_n353_ );
nand g210 ( new_n361_, new_n360_, new_n320_ );
nor g211 ( new_n362_, new_n361_, new_n284_ );
not g212 ( new_n363_, new_n362_ );
not g213 ( new_n364_, N126 );
not g214 ( new_n365_, new_n352_ );
nand g215 ( new_n366_, new_n365_, new_n350_ );
nand g216 ( new_n367_, new_n318_, new_n285_ );
nand g217 ( new_n368_, new_n367_, new_n366_ );
nor g218 ( new_n369_, new_n368_, new_n319_ );
nor g219 ( new_n370_, new_n369_, keyIn_0_21 );
nor g220 ( new_n371_, new_n370_, new_n364_ );
nand g221 ( new_n372_, new_n371_, new_n363_ );
nor g222 ( new_n373_, new_n372_, new_n283_ );
not g223 ( new_n374_, new_n373_ );
not g224 ( new_n375_, keyIn_0_24 );
not g225 ( new_n376_, keyIn_0_20 );
nand g226 ( new_n377_, new_n313_, keyIn_0_5 );
not g227 ( new_n378_, new_n377_ );
nor g228 ( new_n379_, new_n313_, keyIn_0_5 );
nor g229 ( new_n380_, new_n378_, new_n379_ );
nor g230 ( new_n381_, new_n380_, new_n161_ );
nand g231 ( new_n382_, new_n299_, new_n381_ );
nand g232 ( new_n383_, new_n382_, new_n376_ );
not g233 ( new_n384_, N1 );
nand g234 ( new_n385_, keyIn_0_20, N17 );
nor g235 ( new_n386_, new_n380_, new_n385_ );
not g236 ( new_n387_, new_n386_ );
nor g237 ( new_n388_, new_n356_, new_n387_ );
nor g238 ( new_n389_, new_n388_, new_n384_ );
nand g239 ( new_n390_, new_n383_, new_n389_ );
nor g240 ( new_n391_, new_n390_, new_n375_ );
nand g241 ( new_n392_, new_n390_, new_n375_ );
nand g242 ( new_n393_, new_n392_, N153 );
nor g243 ( new_n394_, new_n393_, new_n391_ );
nand g244 ( new_n395_, new_n361_, new_n284_ );
nand g245 ( new_n396_, new_n395_, N126 );
nor g246 ( new_n397_, new_n396_, new_n362_ );
nor g247 ( new_n398_, new_n397_, keyIn_0_31 );
nor g248 ( new_n399_, new_n398_, new_n394_ );
nand g249 ( new_n400_, new_n399_, new_n374_ );
nand g250 ( new_n401_, new_n400_, keyIn_0_37 );
not g251 ( new_n402_, keyIn_0_37 );
not g252 ( new_n403_, new_n394_ );
nand g253 ( new_n404_, new_n372_, new_n283_ );
nand g254 ( new_n405_, new_n404_, new_n403_ );
nor g255 ( new_n406_, new_n405_, new_n373_ );
nand g256 ( new_n407_, new_n406_, new_n402_ );
nand g257 ( new_n408_, new_n401_, new_n407_ );
not g258 ( new_n409_, keyIn_0_18 );
nand g259 ( new_n410_, N29, N75 );
nor g260 ( new_n411_, new_n410_, new_n154_ );
nor g261 ( new_n412_, new_n411_, keyIn_0_2 );
nand g262 ( new_n413_, new_n411_, keyIn_0_2 );
not g263 ( new_n414_, new_n413_ );
nor g264 ( new_n415_, new_n414_, new_n412_ );
nor g265 ( new_n416_, new_n356_, new_n415_ );
nand g266 ( new_n417_, new_n416_, N55 );
nor g267 ( new_n418_, new_n417_, new_n409_ );
nand g268 ( new_n419_, new_n417_, new_n409_ );
nand g269 ( new_n420_, keyIn_0_4, N268 );
not g270 ( new_n421_, new_n420_ );
nor g271 ( new_n422_, keyIn_0_4, N268 );
nor g272 ( new_n423_, new_n421_, new_n422_ );
nor g273 ( new_n424_, new_n423_, keyIn_0_12 );
nand g274 ( new_n425_, new_n423_, keyIn_0_12 );
not g275 ( new_n426_, new_n425_ );
nor g276 ( new_n427_, new_n426_, new_n424_ );
not g277 ( new_n428_, new_n427_ );
nand g278 ( new_n429_, new_n419_, new_n428_ );
nor g279 ( new_n430_, new_n429_, new_n418_ );
not g280 ( new_n431_, new_n430_ );
nand g281 ( new_n432_, new_n431_, keyIn_0_28 );
not g282 ( new_n433_, keyIn_0_28 );
nand g283 ( new_n434_, new_n430_, new_n433_ );
nand g284 ( new_n435_, new_n432_, new_n434_ );
nand g285 ( new_n436_, new_n408_, new_n435_ );
nand g286 ( new_n437_, new_n436_, new_n282_ );
not g287 ( new_n438_, new_n436_ );
nand g288 ( new_n439_, new_n438_, keyIn_0_43 );
nand g289 ( new_n440_, new_n439_, new_n437_ );
nand g290 ( new_n441_, new_n440_, N201 );
not g291 ( new_n442_, new_n441_ );
nor g292 ( new_n443_, new_n440_, N201 );
nor g293 ( new_n444_, new_n442_, new_n443_ );
not g294 ( new_n445_, new_n444_ );
nor g295 ( new_n446_, new_n445_, new_n281_ );
nand g296 ( new_n447_, new_n445_, new_n281_ );
nand g297 ( new_n448_, new_n447_, N219 );
nor g298 ( new_n449_, new_n448_, new_n446_ );
not g299 ( new_n450_, N228 );
nor g300 ( new_n451_, new_n445_, new_n450_ );
not g301 ( new_n452_, N237 );
nor g302 ( new_n453_, new_n441_, new_n452_ );
not g303 ( new_n454_, N246 );
not g304 ( new_n455_, new_n437_ );
nor g305 ( new_n456_, new_n436_, new_n282_ );
nor g306 ( new_n457_, new_n455_, new_n456_ );
nor g307 ( new_n458_, new_n457_, new_n454_ );
not g308 ( new_n459_, N201 );
not g309 ( new_n460_, keyIn_0_10 );
nand g310 ( new_n461_, N42, N72 );
nor g311 ( new_n462_, new_n198_, new_n461_ );
not g312 ( new_n463_, new_n462_ );
nand g313 ( new_n464_, new_n463_, new_n460_ );
not g314 ( new_n465_, N73 );
nor g315 ( new_n466_, new_n463_, new_n460_ );
nor g316 ( new_n467_, new_n466_, new_n465_ );
nand g317 ( new_n468_, new_n467_, new_n464_ );
nor g318 ( new_n469_, new_n468_, new_n459_ );
nand g319 ( new_n470_, N255, N267 );
nand g320 ( new_n471_, N121, N210 );
nand g321 ( new_n472_, new_n470_, new_n471_ );
nor g322 ( new_n473_, new_n469_, new_n472_ );
not g323 ( new_n474_, new_n473_ );
nor g324 ( new_n475_, new_n458_, new_n474_ );
not g325 ( new_n476_, new_n475_ );
nor g326 ( new_n477_, new_n476_, new_n453_ );
not g327 ( new_n478_, new_n477_ );
nor g328 ( new_n479_, new_n478_, new_n451_ );
not g329 ( new_n480_, new_n479_ );
nor g330 ( new_n481_, new_n480_, new_n449_ );
not g331 ( new_n482_, new_n481_ );
nand g332 ( new_n483_, new_n482_, keyIn_0_52 );
not g333 ( new_n484_, keyIn_0_52 );
nand g334 ( new_n485_, new_n481_, new_n484_ );
nand g335 ( N850, new_n483_, new_n485_ );
not g336 ( new_n487_, keyIn_0_57 );
not g337 ( new_n488_, N116 );
nor g338 ( new_n489_, new_n370_, new_n488_ );
nand g339 ( new_n490_, new_n489_, new_n363_ );
nand g340 ( new_n491_, new_n392_, N146 );
nor g341 ( new_n492_, new_n491_, new_n391_ );
not g342 ( new_n493_, new_n492_ );
nand g343 ( new_n494_, new_n490_, new_n493_ );
nor g344 ( new_n495_, new_n494_, keyIn_0_35 );
nor g345 ( new_n496_, new_n430_, keyIn_0_26 );
nand g346 ( new_n497_, new_n430_, keyIn_0_26 );
not g347 ( new_n498_, new_n497_ );
nor g348 ( new_n499_, new_n498_, new_n496_ );
not g349 ( new_n500_, new_n499_ );
nand g350 ( new_n501_, new_n494_, keyIn_0_35 );
nand g351 ( new_n502_, new_n501_, new_n500_ );
nor g352 ( new_n503_, new_n502_, new_n495_ );
nor g353 ( new_n504_, new_n503_, keyIn_0_41 );
not g354 ( new_n505_, keyIn_0_41 );
not g355 ( new_n506_, new_n495_ );
not g356 ( new_n507_, keyIn_0_35 );
nand g357 ( new_n508_, new_n395_, N116 );
nor g358 ( new_n509_, new_n508_, new_n362_ );
nor g359 ( new_n510_, new_n509_, new_n492_ );
nor g360 ( new_n511_, new_n510_, new_n507_ );
nor g361 ( new_n512_, new_n511_, new_n499_ );
nand g362 ( new_n513_, new_n512_, new_n506_ );
nor g363 ( new_n514_, new_n513_, new_n505_ );
nor g364 ( new_n515_, new_n514_, new_n504_ );
nor g365 ( new_n516_, new_n515_, N189 );
not g366 ( new_n517_, keyIn_0_36 );
not g367 ( new_n518_, N121 );
nor g368 ( new_n519_, new_n370_, new_n518_ );
nand g369 ( new_n520_, new_n519_, new_n363_ );
nand g370 ( new_n521_, new_n392_, N149 );
nor g371 ( new_n522_, new_n521_, new_n391_ );
not g372 ( new_n523_, new_n522_ );
nand g373 ( new_n524_, new_n520_, new_n523_ );
nor g374 ( new_n525_, new_n524_, new_n517_ );
not g375 ( new_n526_, new_n525_ );
not g376 ( new_n527_, keyIn_0_27 );
nor g377 ( new_n528_, new_n430_, new_n527_ );
nor g378 ( new_n529_, new_n431_, keyIn_0_27 );
nor g379 ( new_n530_, new_n529_, new_n528_ );
nand g380 ( new_n531_, new_n395_, N121 );
nor g381 ( new_n532_, new_n531_, new_n362_ );
nor g382 ( new_n533_, new_n532_, new_n522_ );
nor g383 ( new_n534_, new_n533_, keyIn_0_36 );
nor g384 ( new_n535_, new_n534_, new_n530_ );
nand g385 ( new_n536_, new_n535_, new_n526_ );
nand g386 ( new_n537_, new_n536_, keyIn_0_42 );
not g387 ( new_n538_, keyIn_0_42 );
not g388 ( new_n539_, new_n530_ );
nand g389 ( new_n540_, new_n524_, new_n517_ );
nand g390 ( new_n541_, new_n540_, new_n539_ );
nor g391 ( new_n542_, new_n541_, new_n525_ );
nand g392 ( new_n543_, new_n542_, new_n538_ );
nand g393 ( new_n544_, new_n537_, new_n543_ );
nor g394 ( new_n545_, new_n544_, N195 );
nor g395 ( new_n546_, new_n516_, new_n545_ );
nor g396 ( new_n547_, new_n443_, new_n281_ );
nand g397 ( new_n548_, new_n547_, new_n546_ );
nand g398 ( new_n549_, new_n548_, keyIn_0_44 );
not g399 ( new_n550_, keyIn_0_44 );
not g400 ( new_n551_, new_n546_ );
nand g401 ( new_n552_, new_n457_, new_n459_ );
nand g402 ( new_n553_, new_n552_, N261 );
nor g403 ( new_n554_, new_n553_, new_n551_ );
nand g404 ( new_n555_, new_n554_, new_n550_ );
nand g405 ( new_n556_, new_n549_, new_n555_ );
nor g406 ( new_n557_, new_n551_, new_n441_ );
nor g407 ( new_n558_, new_n557_, keyIn_0_46 );
nand g408 ( new_n559_, new_n546_, keyIn_0_46 );
nor g409 ( new_n560_, new_n559_, new_n441_ );
not g410 ( new_n561_, new_n560_ );
not g411 ( new_n562_, keyIn_0_45 );
nand g412 ( new_n563_, new_n544_, N195 );
nor g413 ( new_n564_, new_n516_, new_n563_ );
nor g414 ( new_n565_, new_n564_, new_n562_ );
not g415 ( new_n566_, N189 );
nand g416 ( new_n567_, new_n513_, new_n505_ );
nand g417 ( new_n568_, new_n503_, keyIn_0_41 );
nand g418 ( new_n569_, new_n567_, new_n568_ );
nand g419 ( new_n570_, new_n569_, new_n566_ );
not g420 ( new_n571_, N195 );
nor g421 ( new_n572_, new_n542_, new_n538_ );
nor g422 ( new_n573_, new_n536_, keyIn_0_42 );
nor g423 ( new_n574_, new_n573_, new_n572_ );
nor g424 ( new_n575_, new_n574_, new_n571_ );
nand g425 ( new_n576_, new_n575_, new_n570_ );
nor g426 ( new_n577_, new_n576_, keyIn_0_45 );
nor g427 ( new_n578_, new_n565_, new_n577_ );
nor g428 ( new_n579_, new_n569_, new_n566_ );
nor g429 ( new_n580_, new_n578_, new_n579_ );
nand g430 ( new_n581_, new_n580_, new_n561_ );
nor g431 ( new_n582_, new_n581_, new_n558_ );
nand g432 ( new_n583_, new_n582_, new_n556_ );
nand g433 ( new_n584_, new_n583_, keyIn_0_48 );
not g434 ( new_n585_, keyIn_0_48 );
nor g435 ( new_n586_, new_n554_, new_n550_ );
nor g436 ( new_n587_, new_n548_, keyIn_0_44 );
nor g437 ( new_n588_, new_n586_, new_n587_ );
not g438 ( new_n589_, new_n558_ );
nand g439 ( new_n590_, new_n576_, keyIn_0_45 );
nand g440 ( new_n591_, new_n564_, new_n562_ );
nand g441 ( new_n592_, new_n591_, new_n590_ );
not g442 ( new_n593_, new_n579_ );
nand g443 ( new_n594_, new_n592_, new_n593_ );
nor g444 ( new_n595_, new_n594_, new_n560_ );
nand g445 ( new_n596_, new_n595_, new_n589_ );
nor g446 ( new_n597_, new_n588_, new_n596_ );
nand g447 ( new_n598_, new_n597_, new_n585_ );
nand g448 ( new_n599_, new_n598_, new_n584_ );
not g449 ( new_n600_, new_n599_ );
not g450 ( new_n601_, N183 );
nor g451 ( new_n602_, new_n362_, new_n370_ );
nand g452 ( new_n603_, new_n602_, N111 );
not g453 ( new_n604_, new_n603_ );
nand g454 ( new_n605_, new_n392_, N143 );
nor g455 ( new_n606_, new_n605_, new_n391_ );
nor g456 ( new_n607_, new_n604_, new_n606_ );
not g457 ( new_n608_, new_n607_ );
nand g458 ( new_n609_, new_n608_, keyIn_0_34 );
not g459 ( new_n610_, keyIn_0_34 );
nand g460 ( new_n611_, new_n607_, new_n610_ );
nand g461 ( new_n612_, new_n609_, new_n611_ );
not g462 ( new_n613_, keyIn_0_25 );
nand g463 ( new_n614_, new_n431_, new_n613_ );
nand g464 ( new_n615_, new_n430_, keyIn_0_25 );
nand g465 ( new_n616_, new_n614_, new_n615_ );
nand g466 ( new_n617_, new_n612_, new_n616_ );
nand g467 ( new_n618_, new_n617_, keyIn_0_40 );
not g468 ( new_n619_, new_n618_ );
nor g469 ( new_n620_, new_n617_, keyIn_0_40 );
nor g470 ( new_n621_, new_n619_, new_n620_ );
nor g471 ( new_n622_, new_n621_, new_n601_ );
not g472 ( new_n623_, new_n621_ );
nor g473 ( new_n624_, new_n623_, N183 );
nor g474 ( new_n625_, new_n624_, new_n622_ );
not g475 ( new_n626_, new_n625_ );
nor g476 ( new_n627_, new_n600_, new_n626_ );
not g477 ( new_n628_, N219 );
nor g478 ( new_n629_, new_n599_, new_n625_ );
nor g479 ( new_n630_, new_n629_, new_n628_ );
not g480 ( new_n631_, new_n630_ );
nor g481 ( new_n632_, new_n631_, new_n627_ );
nor g482 ( new_n633_, new_n626_, new_n450_ );
not g483 ( new_n634_, new_n622_ );
nor g484 ( new_n635_, new_n634_, new_n452_ );
nor g485 ( new_n636_, new_n621_, new_n454_ );
nand g486 ( new_n637_, N106, N210 );
not g487 ( new_n638_, new_n637_ );
nor g488 ( new_n639_, new_n468_, new_n601_ );
nor g489 ( new_n640_, new_n639_, new_n638_ );
not g490 ( new_n641_, new_n640_ );
nor g491 ( new_n642_, new_n636_, new_n641_ );
not g492 ( new_n643_, new_n642_ );
nor g493 ( new_n644_, new_n635_, new_n643_ );
not g494 ( new_n645_, new_n644_ );
nor g495 ( new_n646_, new_n645_, new_n633_ );
not g496 ( new_n647_, new_n646_ );
nor g497 ( new_n648_, new_n632_, new_n647_ );
not g498 ( new_n649_, new_n648_ );
nand g499 ( new_n650_, new_n649_, new_n487_ );
nand g500 ( new_n651_, new_n648_, keyIn_0_57 );
nand g501 ( N863, new_n650_, new_n651_ );
not g502 ( new_n653_, keyIn_0_49 );
nor g503 ( new_n654_, new_n547_, new_n442_ );
nor g504 ( new_n655_, new_n654_, new_n545_ );
not g505 ( new_n656_, new_n655_ );
nand g506 ( new_n657_, new_n656_, new_n563_ );
nand g507 ( new_n658_, new_n657_, new_n653_ );
not g508 ( new_n659_, new_n658_ );
nor g509 ( new_n660_, new_n657_, new_n653_ );
nor g510 ( new_n661_, new_n659_, new_n660_ );
nor g511 ( new_n662_, new_n516_, new_n579_ );
nor g512 ( new_n663_, new_n661_, new_n662_ );
nand g513 ( new_n664_, new_n661_, new_n662_ );
nand g514 ( new_n665_, new_n664_, N219 );
nor g515 ( new_n666_, new_n665_, new_n663_ );
nand g516 ( new_n667_, new_n662_, N228 );
nor g517 ( new_n668_, new_n593_, new_n452_ );
nor g518 ( new_n669_, new_n569_, new_n454_ );
nor g519 ( new_n670_, new_n468_, new_n566_ );
nand g520 ( new_n671_, N255, N259 );
nand g521 ( new_n672_, N111, N210 );
nand g522 ( new_n673_, new_n671_, new_n672_ );
nor g523 ( new_n674_, new_n670_, new_n673_ );
not g524 ( new_n675_, new_n674_ );
nor g525 ( new_n676_, new_n669_, new_n675_ );
not g526 ( new_n677_, new_n676_ );
nor g527 ( new_n678_, new_n668_, new_n677_ );
nand g528 ( new_n679_, new_n678_, new_n667_ );
nor g529 ( new_n680_, new_n666_, new_n679_ );
not g530 ( new_n681_, new_n680_ );
nand g531 ( new_n682_, new_n681_, keyIn_0_58 );
not g532 ( new_n683_, keyIn_0_58 );
nand g533 ( new_n684_, new_n680_, new_n683_ );
nand g534 ( N864, new_n682_, new_n684_ );
nor g535 ( new_n686_, new_n656_, new_n575_ );
nor g536 ( new_n687_, new_n575_, new_n545_ );
not g537 ( new_n688_, new_n687_ );
nand g538 ( new_n689_, new_n654_, new_n688_ );
nand g539 ( new_n690_, new_n689_, N219 );
nor g540 ( new_n691_, new_n686_, new_n690_ );
nor g541 ( new_n692_, new_n688_, new_n450_ );
nor g542 ( new_n693_, new_n563_, new_n452_ );
nand g543 ( new_n694_, new_n544_, N246 );
nor g544 ( new_n695_, new_n468_, new_n571_ );
nand g545 ( new_n696_, N255, N260 );
nand g546 ( new_n697_, N116, N210 );
nand g547 ( new_n698_, new_n696_, new_n697_ );
nor g548 ( new_n699_, new_n695_, new_n698_ );
nand g549 ( new_n700_, new_n694_, new_n699_ );
nor g550 ( new_n701_, new_n693_, new_n700_ );
not g551 ( new_n702_, new_n701_ );
nor g552 ( new_n703_, new_n692_, new_n702_ );
not g553 ( new_n704_, new_n703_ );
nor g554 ( new_n705_, new_n691_, new_n704_ );
not g555 ( new_n706_, new_n705_ );
nand g556 ( new_n707_, new_n706_, keyIn_0_59 );
not g557 ( new_n708_, keyIn_0_59 );
nand g558 ( new_n709_, new_n705_, new_n708_ );
nand g559 ( N865, new_n707_, new_n709_ );
not g560 ( new_n711_, keyIn_0_55 );
nand g561 ( new_n712_, new_n602_, N96 );
not g562 ( new_n713_, keyIn_0_17 );
nand g563 ( new_n714_, new_n416_, N17 );
nor g564 ( new_n715_, new_n714_, new_n713_ );
not g565 ( new_n716_, new_n423_ );
nand g566 ( new_n717_, new_n714_, new_n713_ );
nand g567 ( new_n718_, new_n717_, new_n716_ );
nor g568 ( new_n719_, new_n718_, new_n715_ );
nand g569 ( new_n720_, N51, N138 );
not g570 ( new_n721_, keyIn_0_16 );
nor g571 ( new_n722_, new_n380_, new_n190_ );
nand g572 ( new_n723_, new_n299_, new_n722_ );
not g573 ( new_n724_, new_n723_ );
nor g574 ( new_n725_, new_n724_, new_n721_ );
nor g575 ( new_n726_, new_n723_, keyIn_0_16 );
nor g576 ( new_n727_, new_n725_, new_n726_ );
not g577 ( new_n728_, new_n727_ );
nand g578 ( new_n729_, new_n728_, N146 );
nand g579 ( new_n730_, new_n729_, new_n720_ );
nor g580 ( new_n731_, new_n730_, new_n719_ );
nand g581 ( new_n732_, new_n731_, new_n712_ );
nor g582 ( new_n733_, new_n732_, N165 );
not g583 ( new_n734_, keyIn_0_38 );
not g584 ( new_n735_, keyIn_0_22 );
nor g585 ( new_n736_, new_n719_, new_n735_ );
not g586 ( new_n737_, new_n719_ );
nor g587 ( new_n738_, new_n737_, keyIn_0_22 );
nor g588 ( new_n739_, new_n738_, new_n736_ );
nand g589 ( new_n740_, new_n728_, N149 );
not g590 ( new_n741_, new_n740_ );
nor g591 ( new_n742_, new_n739_, new_n741_ );
not g592 ( new_n743_, new_n742_ );
nand g593 ( new_n744_, new_n743_, keyIn_0_29 );
not g594 ( new_n745_, new_n744_ );
nor g595 ( new_n746_, new_n743_, keyIn_0_29 );
nor g596 ( new_n747_, new_n745_, new_n746_ );
not g597 ( new_n748_, keyIn_0_32 );
nand g598 ( new_n749_, new_n602_, N101 );
nand g599 ( new_n750_, N17, N138 );
nand g600 ( new_n751_, new_n749_, new_n750_ );
not g601 ( new_n752_, new_n751_ );
nor g602 ( new_n753_, new_n752_, new_n748_ );
nor g603 ( new_n754_, new_n751_, keyIn_0_32 );
nor g604 ( new_n755_, new_n753_, new_n754_ );
nor g605 ( new_n756_, new_n747_, new_n755_ );
not g606 ( new_n757_, new_n756_ );
nand g607 ( new_n758_, new_n757_, new_n734_ );
not g608 ( new_n759_, new_n758_ );
nor g609 ( new_n760_, new_n757_, new_n734_ );
nor g610 ( new_n761_, new_n759_, new_n760_ );
not g611 ( new_n762_, new_n761_ );
nor g612 ( new_n763_, new_n762_, N171 );
not g613 ( new_n764_, keyIn_0_39 );
not g614 ( new_n765_, keyIn_0_30 );
nor g615 ( new_n766_, new_n719_, keyIn_0_23 );
nand g616 ( new_n767_, new_n719_, keyIn_0_23 );
not g617 ( new_n768_, new_n767_ );
nor g618 ( new_n769_, new_n768_, new_n766_ );
nand g619 ( new_n770_, new_n728_, N153 );
not g620 ( new_n771_, new_n770_ );
nor g621 ( new_n772_, new_n769_, new_n771_ );
not g622 ( new_n773_, new_n772_ );
nand g623 ( new_n774_, new_n773_, new_n765_ );
not g624 ( new_n775_, new_n774_ );
nor g625 ( new_n776_, new_n773_, new_n765_ );
nor g626 ( new_n777_, new_n775_, new_n776_ );
not g627 ( new_n778_, keyIn_0_33 );
nand g628 ( new_n779_, new_n602_, N106 );
nand g629 ( new_n780_, N138, N152 );
nand g630 ( new_n781_, new_n779_, new_n780_ );
not g631 ( new_n782_, new_n781_ );
nor g632 ( new_n783_, new_n782_, new_n778_ );
nor g633 ( new_n784_, new_n781_, keyIn_0_33 );
nor g634 ( new_n785_, new_n783_, new_n784_ );
nor g635 ( new_n786_, new_n777_, new_n785_ );
not g636 ( new_n787_, new_n786_ );
nand g637 ( new_n788_, new_n787_, new_n764_ );
not g638 ( new_n789_, new_n788_ );
nor g639 ( new_n790_, new_n787_, new_n764_ );
nor g640 ( new_n791_, new_n789_, new_n790_ );
not g641 ( new_n792_, new_n791_ );
nor g642 ( new_n793_, new_n792_, N177 );
nor g643 ( new_n794_, new_n763_, new_n793_ );
not g644 ( new_n795_, new_n794_ );
nor g645 ( new_n796_, new_n795_, new_n733_ );
not g646 ( new_n797_, keyIn_0_51 );
not g647 ( new_n798_, keyIn_0_50 );
not g648 ( new_n799_, new_n624_ );
nand g649 ( new_n800_, new_n599_, new_n799_ );
nand g650 ( new_n801_, new_n800_, new_n798_ );
nor g651 ( new_n802_, new_n800_, new_n798_ );
not g652 ( new_n803_, new_n802_ );
nand g653 ( new_n804_, new_n803_, new_n801_ );
nand g654 ( new_n805_, new_n804_, new_n634_ );
nand g655 ( new_n806_, new_n805_, new_n797_ );
not g656 ( new_n807_, new_n801_ );
nor g657 ( new_n808_, new_n807_, new_n802_ );
nor g658 ( new_n809_, new_n808_, new_n622_ );
nand g659 ( new_n810_, new_n809_, keyIn_0_51 );
nand g660 ( new_n811_, new_n810_, new_n806_ );
nand g661 ( new_n812_, new_n811_, new_n796_ );
nor g662 ( new_n813_, new_n812_, keyIn_0_54 );
not g663 ( new_n814_, new_n813_ );
nand g664 ( new_n815_, new_n812_, keyIn_0_54 );
not g665 ( new_n816_, keyIn_0_47 );
not g666 ( new_n817_, new_n733_ );
not g667 ( new_n818_, N177 );
nor g668 ( new_n819_, new_n791_, new_n818_ );
not g669 ( new_n820_, new_n819_ );
nor g670 ( new_n821_, new_n763_, new_n820_ );
nand g671 ( new_n822_, new_n821_, new_n817_ );
nor g672 ( new_n823_, new_n822_, new_n816_ );
nand g673 ( new_n824_, new_n822_, new_n816_ );
not g674 ( new_n825_, N165 );
not g675 ( new_n826_, new_n732_ );
nor g676 ( new_n827_, new_n826_, new_n825_ );
not g677 ( new_n828_, N171 );
nor g678 ( new_n829_, new_n761_, new_n828_ );
not g679 ( new_n830_, new_n829_ );
nor g680 ( new_n831_, new_n830_, new_n733_ );
nor g681 ( new_n832_, new_n831_, new_n827_ );
nand g682 ( new_n833_, new_n824_, new_n832_ );
nor g683 ( new_n834_, new_n833_, new_n823_ );
nand g684 ( new_n835_, new_n815_, new_n834_ );
not g685 ( new_n836_, new_n835_ );
nand g686 ( new_n837_, new_n836_, new_n814_ );
nand g687 ( new_n838_, new_n837_, new_n711_ );
nor g688 ( new_n839_, new_n835_, new_n813_ );
nand g689 ( new_n840_, new_n839_, keyIn_0_55 );
nand g690 ( new_n841_, new_n838_, new_n840_ );
nand g691 ( new_n842_, new_n602_, N91 );
nand g692 ( new_n843_, N8, N138 );
nand g693 ( new_n844_, new_n728_, N143 );
nand g694 ( new_n845_, new_n844_, new_n843_ );
nor g695 ( new_n846_, new_n845_, new_n719_ );
nand g696 ( new_n847_, new_n846_, new_n842_ );
nor g697 ( new_n848_, new_n847_, N159 );
not g698 ( new_n849_, new_n848_ );
nand g699 ( new_n850_, new_n841_, new_n849_ );
not g700 ( new_n851_, N159 );
not g701 ( new_n852_, new_n847_ );
nor g702 ( new_n853_, new_n852_, new_n851_ );
not g703 ( new_n854_, new_n853_ );
nand g704 ( N866, new_n850_, new_n854_ );
not g705 ( new_n856_, new_n811_ );
nor g706 ( new_n857_, new_n856_, new_n793_ );
not g707 ( new_n858_, new_n857_ );
nor g708 ( new_n859_, new_n858_, new_n819_ );
nor g709 ( new_n860_, new_n793_, new_n819_ );
nor g710 ( new_n861_, new_n811_, new_n860_ );
nor g711 ( new_n862_, new_n861_, new_n628_ );
not g712 ( new_n863_, new_n862_ );
nor g713 ( new_n864_, new_n859_, new_n863_ );
nand g714 ( new_n865_, new_n860_, N228 );
nor g715 ( new_n866_, new_n820_, new_n452_ );
nor g716 ( new_n867_, new_n791_, new_n454_ );
nand g717 ( new_n868_, N101, N210 );
not g718 ( new_n869_, new_n868_ );
nor g719 ( new_n870_, new_n468_, new_n818_ );
nor g720 ( new_n871_, new_n870_, new_n869_ );
not g721 ( new_n872_, new_n871_ );
nor g722 ( new_n873_, new_n867_, new_n872_ );
not g723 ( new_n874_, new_n873_ );
nor g724 ( new_n875_, new_n866_, new_n874_ );
nand g725 ( new_n876_, new_n875_, new_n865_ );
nor g726 ( new_n877_, new_n864_, new_n876_ );
not g727 ( new_n878_, new_n877_ );
nand g728 ( new_n879_, new_n878_, keyIn_0_60 );
not g729 ( new_n880_, keyIn_0_60 );
nand g730 ( new_n881_, new_n877_, new_n880_ );
nand g731 ( N874, new_n879_, new_n881_ );
nor g732 ( new_n883_, new_n839_, keyIn_0_55 );
nor g733 ( new_n884_, new_n837_, new_n711_ );
nor g734 ( new_n885_, new_n884_, new_n883_ );
nor g735 ( new_n886_, new_n853_, new_n848_ );
not g736 ( new_n887_, new_n886_ );
nor g737 ( new_n888_, new_n885_, new_n887_ );
not g738 ( new_n889_, new_n888_ );
nor g739 ( new_n890_, new_n841_, new_n886_ );
nor g740 ( new_n891_, new_n890_, new_n628_ );
nand g741 ( new_n892_, new_n891_, new_n889_ );
nor g742 ( new_n893_, new_n887_, new_n450_ );
nor g743 ( new_n894_, new_n854_, new_n452_ );
nor g744 ( new_n895_, new_n852_, new_n454_ );
nor g745 ( new_n896_, new_n468_, new_n851_ );
nand g746 ( new_n897_, new_n427_, N210 );
not g747 ( new_n898_, new_n897_ );
nor g748 ( new_n899_, new_n896_, new_n898_ );
not g749 ( new_n900_, new_n899_ );
nor g750 ( new_n901_, new_n895_, new_n900_ );
not g751 ( new_n902_, new_n901_ );
nor g752 ( new_n903_, new_n894_, new_n902_ );
not g753 ( new_n904_, new_n903_ );
nor g754 ( new_n905_, new_n904_, new_n893_ );
nand g755 ( new_n906_, new_n892_, new_n905_ );
nand g756 ( new_n907_, new_n906_, keyIn_0_61 );
not g757 ( new_n908_, keyIn_0_61 );
nand g758 ( new_n909_, new_n885_, new_n887_ );
nand g759 ( new_n910_, new_n909_, N219 );
nor g760 ( new_n911_, new_n910_, new_n888_ );
not g761 ( new_n912_, new_n905_ );
nor g762 ( new_n913_, new_n911_, new_n912_ );
nand g763 ( new_n914_, new_n913_, new_n908_ );
nand g764 ( N878, new_n914_, new_n907_ );
not g765 ( new_n916_, keyIn_0_62 );
not g766 ( new_n917_, keyIn_0_53 );
nand g767 ( new_n918_, new_n811_, new_n794_ );
nor g768 ( new_n919_, new_n918_, new_n917_ );
nand g769 ( new_n920_, new_n918_, new_n917_ );
nor g770 ( new_n921_, new_n821_, new_n829_ );
nand g771 ( new_n922_, new_n920_, new_n921_ );
nor g772 ( new_n923_, new_n922_, new_n919_ );
nor g773 ( new_n924_, new_n923_, keyIn_0_56 );
not g774 ( new_n925_, keyIn_0_56 );
not g775 ( new_n926_, new_n919_ );
not g776 ( new_n927_, new_n922_ );
nand g777 ( new_n928_, new_n927_, new_n926_ );
nor g778 ( new_n929_, new_n928_, new_n925_ );
nor g779 ( new_n930_, new_n929_, new_n924_ );
nor g780 ( new_n931_, new_n827_, new_n733_ );
nor g781 ( new_n932_, new_n930_, new_n931_ );
not g782 ( new_n933_, new_n932_ );
nand g783 ( new_n934_, new_n928_, new_n925_ );
nand g784 ( new_n935_, new_n923_, keyIn_0_56 );
nand g785 ( new_n936_, new_n934_, new_n935_ );
not g786 ( new_n937_, new_n931_ );
nor g787 ( new_n938_, new_n936_, new_n937_ );
nor g788 ( new_n939_, new_n938_, new_n628_ );
nand g789 ( new_n940_, new_n939_, new_n933_ );
nor g790 ( new_n941_, new_n937_, new_n450_ );
nand g791 ( new_n942_, new_n827_, N237 );
nor g792 ( new_n943_, new_n826_, new_n454_ );
nand g793 ( new_n944_, N91, N210 );
not g794 ( new_n945_, new_n944_ );
nor g795 ( new_n946_, new_n468_, new_n825_ );
nor g796 ( new_n947_, new_n946_, new_n945_ );
not g797 ( new_n948_, new_n947_ );
nor g798 ( new_n949_, new_n943_, new_n948_ );
nand g799 ( new_n950_, new_n949_, new_n942_ );
nor g800 ( new_n951_, new_n941_, new_n950_ );
nand g801 ( new_n952_, new_n940_, new_n951_ );
nand g802 ( new_n953_, new_n952_, new_n916_ );
nand g803 ( new_n954_, new_n930_, new_n931_ );
nand g804 ( new_n955_, new_n954_, N219 );
nor g805 ( new_n956_, new_n955_, new_n932_ );
not g806 ( new_n957_, new_n951_ );
nor g807 ( new_n958_, new_n956_, new_n957_ );
nand g808 ( new_n959_, new_n958_, keyIn_0_62 );
nand g809 ( N879, new_n959_, new_n953_ );
not g810 ( new_n961_, keyIn_0_63 );
nand g811 ( new_n962_, new_n858_, new_n820_ );
nor g812 ( new_n963_, new_n763_, new_n829_ );
nand g813 ( new_n964_, new_n962_, new_n963_ );
nor g814 ( new_n965_, new_n962_, new_n963_ );
nor g815 ( new_n966_, new_n965_, new_n628_ );
nand g816 ( new_n967_, new_n966_, new_n964_ );
nand g817 ( new_n968_, new_n963_, N228 );
nor g818 ( new_n969_, new_n830_, new_n452_ );
nor g819 ( new_n970_, new_n761_, new_n454_ );
nand g820 ( new_n971_, N96, N210 );
not g821 ( new_n972_, new_n971_ );
nor g822 ( new_n973_, new_n468_, new_n828_ );
nor g823 ( new_n974_, new_n973_, new_n972_ );
not g824 ( new_n975_, new_n974_ );
nor g825 ( new_n976_, new_n970_, new_n975_ );
not g826 ( new_n977_, new_n976_ );
nor g827 ( new_n978_, new_n969_, new_n977_ );
nand g828 ( new_n979_, new_n978_, new_n968_ );
not g829 ( new_n980_, new_n979_ );
nand g830 ( new_n981_, new_n967_, new_n980_ );
nand g831 ( new_n982_, new_n981_, new_n961_ );
not g832 ( new_n983_, new_n981_ );
nand g833 ( new_n984_, new_n983_, keyIn_0_63 );
nand g834 ( N880, new_n984_, new_n982_ );
endmodule