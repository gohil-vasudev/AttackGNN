module rs232 ( sys_clk, sys_rst_l, uart_XMIT_dataH, xmitH, xmit_dataH_7_, 
        xmit_dataH_6_, xmit_dataH_5_, xmit_dataH_4_, xmit_dataH_3_, 
        xmit_dataH_2_, xmit_dataH_1_, xmit_dataH_0_, xmit_doneH, 
        uart_REC_dataH, rec_dataH_7_, rec_dataH_6_, rec_dataH_5_, rec_dataH_4_, 
        rec_dataH_3_, rec_dataH_2_, rec_dataH_1_, rec_dataH_0_, rec_readyH, 
        test_mode, test_se, test_si, test_so );
  input sys_clk, sys_rst_l, xmitH, xmit_dataH_7_, xmit_dataH_6_, xmit_dataH_5_,
         xmit_dataH_4_, xmit_dataH_3_, xmit_dataH_2_, xmit_dataH_1_,
         xmit_dataH_0_, uart_REC_dataH, test_mode, test_se, test_si;
  output uart_XMIT_dataH, xmit_doneH, rec_dataH_7_, rec_dataH_6_, rec_dataH_5_,
         rec_dataH_4_, rec_dataH_3_, rec_dataH_2_, rec_dataH_1_, rec_dataH_0_,
         rec_readyH, test_so;
  wire   rec_dataH_temp_6, rec_dataH_temp_5, rec_dataH_temp_4,
         rec_dataH_temp_3, rec_dataH_temp_2, rec_dataH_temp_1,
         rec_dataH_temp_0, iCTRL, xmit_doneH_temp, iXMIT_CRTL, iRECEIVER_CTRL,
         iRECEIVER_state_CTRL, iRECEIVER_N_CTRL_1_, iRECEIVER_N_CTRL_2_,
         iRECEIVER_bitCell_CTRL, iRECEIVER_N18, iRECEIVER_N17,
         iRECEIVER_bitCell_cntrH_0_, iRECEIVER_bitCell_cntrH_1_, iRECEIVER_N22,
         iRECEIVER_N21, iRECEIVER_N20, iRECEIVER_N19, n400, iRECEIVER_N27,
         iRECEIVER_N26, iRECEIVER_N23, iRECEIVER_next_state_2_,
         iRECEIVER_state_0_, iRECEIVER_state_1_, iRECEIVER_state_2_,
         iXMIT_state_CTRL, iXMIT_N_CTRL_1_, iXMIT_N_CTRL_2_, iXMIT_xmit_CTRL,
         iXMIT_N24, iXMIT_xmit_ShiftRegH_7_, iXMIT_xmit_ShiftRegH_6_,
         iXMIT_xmit_ShiftRegH_5_, iXMIT_N28, iXMIT_N27, iXMIT_N26, iXMIT_N25,
         iXMIT_N46, iXMIT_N45, iXMIT_N44, iXMIT_N29, iXMIT_state_0_,
         iXMIT_state_1_, iXMIT_state_2_, n255, n241, n244, n245, n238, n242,
         n246, n239, rec_dataH_rec_7, rec_dataH_rec_6, rec_dataH_rec_5,
         rec_dataH_rec_4, rec_dataH_rec_3, rec_dataH_rec_2, rec_dataH_rec_1,
         rec_dataH_rec_0, n181, n180, n179, n178, n177, n176, n175, n174, n173,
         n172, n171, n170, n169, n168, n167, n166, n164, n163, n162, n161,
         n160, n159, n157, n156, n155, n154, test_point_DOUT, n153, n152, n150,
         n149, n148, n147, n146, n145, n143, n142, n141, n140, n139, n138,
         n136, n135, n134, n133, n132, n131, n129, n128, n127, n126, n125,
         n124, n122, n121, n120, n119, n118, n117, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748;

  AND2X4 TrojanU303 ( .IN1(iCTRL), .IN2(xmit_doneH_temp), .Q(xmit_doneH) );
  OR2X1 TrojanU302 ( .IN1(iXMIT_CRTL), .IN2(iRECEIVER_CTRL), .Q(iCTRL) );
  OR4X4 TrojanU301 ( .IN1(iRECEIVER_state_CTRL), .IN2(iRECEIVER_N_CTRL_1_), 
        .IN3(iRECEIVER_N_CTRL_2_), .IN4(iRECEIVER_bitCell_CTRL), .Q(
        iRECEIVER_CTRL) );
  NAND4X1 TrojanU300 ( .IN1(iRECEIVER_N18), .IN2(iRECEIVER_N17), .IN3(
        iRECEIVER_bitCell_cntrH_0_), .IN4(iRECEIVER_bitCell_cntrH_1_), .QN(
        iRECEIVER_bitCell_CTRL) );
  NAND4X1 TrojanU299 ( .IN1(iRECEIVER_N22), .IN2(iRECEIVER_N21), .IN3(
        iRECEIVER_N20), .IN4(iRECEIVER_N19), .QN(iRECEIVER_N_CTRL_2_) );
  NAND4X1 TrojanU298 ( .IN1(n400), .IN2(iRECEIVER_N27), .IN3(iRECEIVER_N26), 
        .IN4(iRECEIVER_N23), .QN(iRECEIVER_N_CTRL_1_) );
  NAND4X1 TrojanU297 ( .IN1(iRECEIVER_next_state_2_), .IN2(iRECEIVER_state_0_), 
        .IN3(iRECEIVER_state_1_), .IN4(iRECEIVER_state_2_), .QN(
        iRECEIVER_state_CTRL) );
  OR4X4 TrojanU296 ( .IN1(iXMIT_state_CTRL), .IN2(iXMIT_N_CTRL_1_), .IN3(
        iXMIT_N_CTRL_2_), .IN4(iXMIT_xmit_CTRL), .Q(iXMIT_CRTL) );
  NAND4X1 TrojanU295 ( .IN1(iXMIT_N24), .IN2(iXMIT_xmit_ShiftRegH_7_), .IN3(
        iXMIT_xmit_ShiftRegH_6_), .IN4(iXMIT_xmit_ShiftRegH_5_), .QN(
        iXMIT_xmit_CTRL) );
  NAND4X1 TrojanU294 ( .IN1(iXMIT_N28), .IN2(iXMIT_N27), .IN3(iXMIT_N26), 
        .IN4(iXMIT_N25), .QN(iXMIT_N_CTRL_2_) );
  NAND4X1 TrojanU293 ( .IN1(iXMIT_N46), .IN2(iXMIT_N45), .IN3(iXMIT_N44), 
        .IN4(iXMIT_N29), .QN(iXMIT_N_CTRL_1_) );
  NAND4X1 TrojanU292 ( .IN1(n422), .IN2(iXMIT_state_0_), .IN3(iXMIT_state_1_), 
        .IN4(iXMIT_state_2_), .QN(iXMIT_state_CTRL) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_2_ ( .D(n181), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n741) );
  DFFARX1 iXMIT_state_reg_0_ ( .D(n180), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        iXMIT_state_0_), .QN(n239) );
  DFFARX1 iXMIT_state_reg_2_ ( .D(n179), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        iXMIT_state_2_), .QN(n242) );
  DFFARX1 iXMIT_state_reg_1_ ( .D(n178), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        iXMIT_state_1_), .QN(n246) );
  DFFARX1 iXMIT_bitCountH_reg_0_ ( .D(n177), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n738), .QN(n425) );
  DFFARX1 iXMIT_bitCountH_reg_1_ ( .D(n176), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n739), .QN(n431) );
  DFFARX1 iXMIT_bitCountH_reg_2_ ( .D(n175), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n737), .QN(n432) );
  DFFARX1 iXMIT_bitCountH_reg_3_ ( .D(n174), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(n736) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_7_ ( .D(n173), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_xmit_ShiftRegH_7_) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_6_ ( .D(n172), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_xmit_ShiftRegH_6_) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_5_ ( .D(n171), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_xmit_ShiftRegH_5_) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_4_ ( .D(n170), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n729) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_3_ ( .D(n169), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n730) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_2_ ( .D(n168), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n731) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_1_ ( .D(n167), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n732) );
  DFFARX1 iXMIT_xmit_doneH_reg ( .D(n166), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(xmit_doneH_temp) );
  DFFARX1 iRECEIVER_state_reg_1_ ( .D(n164), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(iRECEIVER_state_1_), .QN(n241) );
  DFFASX1 iRECEIVER_state_reg_0_ ( .D(n163), .CLK(sys_clk), .SETB(sys_rst_l), 
        .Q(iRECEIVER_state_0_), .QN(n245) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_0_ ( .D(n162), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iRECEIVER_bitCell_cntrH_0_), .QN(n255) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_1_ ( .D(n161), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iRECEIVER_bitCell_cntrH_1_), .QN(n244) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_2_ ( .D(n160), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n748), .QN(n424) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_3_ ( .D(n159), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n747) );
  DFFARX1 iRECEIVER_state_reg_2_ ( .D(n157), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(iRECEIVER_state_2_), .QN(n238) );
  DFFARX1 iRECEIVER_rec_readyH_reg ( .D(n156), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(rec_readyH) );
  DFFARX1 iRECEIVER_par_dataH_reg_7_ ( .D(n155), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_7) );
  DFFARX1 rec_dataH_temp_reg_7_ ( .D(n154), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(test_so) );
  DFFARX1 rec_dataH_reg_7_ ( .D(n153), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_7_) );
  DFFARX1 iRECEIVER_par_dataH_reg_6_ ( .D(n152), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_6) );
  DFFARX1 rec_dataH_temp_reg_6_ ( .D(n150), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_6) );
  DFFARX1 rec_dataH_reg_6_ ( .D(n149), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_6_) );
  DFFARX1 iRECEIVER_par_dataH_reg_5_ ( .D(n148), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_5) );
  DFFARX1 rec_dataH_temp_reg_5_ ( .D(n147), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_5) );
  DFFARX1 rec_dataH_reg_5_ ( .D(n146), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_5_) );
  DFFARX1 iRECEIVER_par_dataH_reg_4_ ( .D(n145), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_4) );
  DFFARX1 rec_dataH_temp_reg_4_ ( .D(n143), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_4) );
  DFFARX1 rec_dataH_reg_4_ ( .D(n142), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_4_) );
  DFFARX1 iRECEIVER_par_dataH_reg_3_ ( .D(n141), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_3) );
  DFFARX1 rec_dataH_temp_reg_3_ ( .D(n140), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_3) );
  DFFARX1 rec_dataH_reg_3_ ( .D(n139), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_3_) );
  DFFARX1 iRECEIVER_par_dataH_reg_2_ ( .D(n138), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_2) );
  DFFARX1 rec_dataH_temp_reg_2_ ( .D(n136), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_2) );
  DFFARX1 rec_dataH_reg_2_ ( .D(n135), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_2_) );
  DFFARX1 iRECEIVER_par_dataH_reg_1_ ( .D(n134), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_1) );
  DFFARX1 rec_dataH_temp_reg_1_ ( .D(n133), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_1) );
  DFFARX1 rec_dataH_reg_1_ ( .D(n132), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_1_) );
  DFFARX1 iRECEIVER_par_dataH_reg_0_ ( .D(n131), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_0) );
  DFFARX1 rec_dataH_temp_reg_0_ ( .D(n129), .CLK(test_point_DOUT), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp_0) );
  DFFARX1 rec_dataH_reg_0_ ( .D(n128), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH_0_) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_3_ ( .D(n127), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n735), .QN(n434) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_0_ ( .D(n126), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n745), .QN(n423) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_1_ ( .D(n125), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n746), .QN(n428) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_2_ ( .D(n124), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n744), .QN(n426) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_3_ ( .D(n122), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n740) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_0_ ( .D(n121), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n743), .QN(n433) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_1_ ( .D(n120), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n742), .QN(n430) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_0_ ( .D(n119), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n427) );
  DFFASX1 iRECEIVER_rec_datSyncH_reg ( .D(n118), .CLK(sys_clk), .SETB(
        sys_rst_l), .Q(n733) );
  DFFASX1 iRECEIVER_rec_datH_reg ( .D(n117), .CLK(sys_clk), .SETB(sys_rst_l), 
        .Q(n734), .QN(n429) );
  DFFASX1 TrojaniDatasend_reg ( .D(n117), .CLK(sys_clk), .SETB(sys_rst_l), .Q(
        n400) );
  OR2X1 U578 ( .IN1(n435), .IN2(n436), .Q(uart_XMIT_dataH) );
  OR2X1 U579 ( .IN1(n437), .IN2(n438), .Q(n436) );
  AND2X1 U580 ( .IN1(n439), .IN2(n427), .Q(n435) );
  OR2X1 U581 ( .IN1(iXMIT_state_2_), .IN2(iXMIT_state_0_), .Q(n439) );
  OR2X1 U582 ( .IN1(n440), .IN2(n441), .Q(test_point_DOUT) );
  AND2X1 U583 ( .IN1(sys_clk), .IN2(test_mode), .Q(n441) );
  AND2X1 U584 ( .IN1(rec_readyH), .IN2(n442), .Q(n440) );
  INVX0 U585 ( .INP(test_mode), .ZN(n442) );
  OR2X1 U586 ( .IN1(n443), .IN2(n444), .Q(n181) );
  AND2X1 U587 ( .IN1(test_se), .IN2(n742), .Q(n444) );
  AND2X1 U588 ( .IN1(iXMIT_N28), .IN2(n445), .Q(n443) );
  OR2X1 U589 ( .IN1(n446), .IN2(n447), .Q(n180) );
  AND2X1 U590 ( .IN1(n448), .IN2(n445), .Q(n447) );
  OR2X1 U591 ( .IN1(n449), .IN2(n450), .Q(n448) );
  AND2X1 U592 ( .IN1(n451), .IN2(n452), .Q(n450) );
  OR2X1 U593 ( .IN1(n453), .IN2(iXMIT_state_0_), .Q(n452) );
  AND2X1 U594 ( .IN1(n454), .IN2(iXMIT_state_1_), .Q(n451) );
  AND2X1 U595 ( .IN1(n455), .IN2(iXMIT_state_2_), .Q(n449) );
  OR2X1 U596 ( .IN1(n239), .IN2(n456), .Q(n455) );
  AND2X1 U597 ( .IN1(n736), .IN2(test_se), .Q(n446) );
  OR2X1 U598 ( .IN1(n457), .IN2(n458), .Q(n179) );
  AND2X1 U599 ( .IN1(n422), .IN2(n445), .Q(n458) );
  OR2X1 U600 ( .IN1(n459), .IN2(n460), .Q(n422) );
  INVX0 U601 ( .INP(n461), .ZN(n460) );
  OR2X1 U602 ( .IN1(n462), .IN2(n246), .Q(n461) );
  AND2X1 U603 ( .IN1(n437), .IN2(n456), .Q(n459) );
  INVX0 U604 ( .INP(n453), .ZN(n456) );
  AND2X1 U605 ( .IN1(test_se), .IN2(iXMIT_state_1_), .Q(n457) );
  OR2X1 U606 ( .IN1(n463), .IN2(n464), .Q(n178) );
  AND2X1 U607 ( .IN1(n465), .IN2(n445), .Q(n464) );
  OR2X1 U608 ( .IN1(n466), .IN2(n467), .Q(n465) );
  AND2X1 U609 ( .IN1(test_se), .IN2(iXMIT_state_0_), .Q(n463) );
  OR2X1 U610 ( .IN1(n468), .IN2(n469), .Q(n177) );
  OR2X1 U611 ( .IN1(n470), .IN2(n471), .Q(n469) );
  AND2X1 U612 ( .IN1(n738), .IN2(n472), .Q(n471) );
  AND2X1 U613 ( .IN1(n473), .IN2(n425), .Q(n470) );
  AND2X1 U614 ( .IN1(test_se), .IN2(n740), .Q(n468) );
  OR2X1 U615 ( .IN1(n474), .IN2(n475), .Q(n176) );
  OR2X1 U616 ( .IN1(n476), .IN2(n477), .Q(n475) );
  AND2X1 U617 ( .IN1(n739), .IN2(n472), .Q(n477) );
  AND2X1 U618 ( .IN1(n473), .IN2(iXMIT_N44), .Q(n476) );
  AND2X1 U619 ( .IN1(n738), .IN2(test_se), .Q(n474) );
  OR2X1 U620 ( .IN1(n478), .IN2(n479), .Q(n175) );
  OR2X1 U621 ( .IN1(n480), .IN2(n481), .Q(n479) );
  AND2X1 U622 ( .IN1(n737), .IN2(n472), .Q(n481) );
  AND2X1 U623 ( .IN1(n473), .IN2(iXMIT_N45), .Q(n480) );
  AND2X1 U624 ( .IN1(n739), .IN2(test_se), .Q(n478) );
  OR2X1 U625 ( .IN1(n482), .IN2(n483), .Q(n174) );
  OR2X1 U626 ( .IN1(n484), .IN2(n485), .Q(n483) );
  AND2X1 U627 ( .IN1(n472), .IN2(n736), .Q(n485) );
  INVX0 U628 ( .INP(n486), .ZN(n472) );
  OR2X1 U629 ( .IN1(n487), .IN2(n488), .Q(n486) );
  OR2X1 U630 ( .IN1(test_se), .IN2(n489), .Q(n488) );
  AND2X1 U631 ( .IN1(n473), .IN2(iXMIT_N46), .Q(n484) );
  AND2X1 U632 ( .IN1(n445), .IN2(n489), .Q(n473) );
  INVX0 U633 ( .INP(n490), .ZN(n489) );
  OR2X1 U634 ( .IN1(n454), .IN2(n491), .Q(n490) );
  OR2X1 U635 ( .IN1(n246), .IN2(n239), .Q(n491) );
  OR2X1 U636 ( .IN1(n492), .IN2(n493), .Q(n454) );
  AND2X1 U637 ( .IN1(n494), .IN2(n495), .Q(n492) );
  AND2X1 U638 ( .IN1(n425), .IN2(n432), .Q(n495) );
  AND2X1 U639 ( .IN1(n736), .IN2(n431), .Q(n494) );
  AND2X1 U640 ( .IN1(n737), .IN2(test_se), .Q(n482) );
  OR2X1 U641 ( .IN1(n496), .IN2(n497), .Q(n173) );
  AND2X1 U642 ( .IN1(n498), .IN2(n445), .Q(n497) );
  OR2X1 U643 ( .IN1(n499), .IN2(n500), .Q(n498) );
  OR2X1 U644 ( .IN1(n501), .IN2(n502), .Q(n500) );
  AND2X1 U645 ( .IN1(xmit_dataH_7_), .IN2(n467), .Q(n502) );
  AND2X1 U646 ( .IN1(n503), .IN2(iXMIT_xmit_ShiftRegH_7_), .Q(n501) );
  AND2X1 U647 ( .IN1(test_se), .IN2(iXMIT_xmit_ShiftRegH_6_), .Q(n496) );
  OR2X1 U648 ( .IN1(n504), .IN2(n505), .Q(n172) );
  AND2X1 U649 ( .IN1(n506), .IN2(n445), .Q(n505) );
  OR2X1 U650 ( .IN1(n507), .IN2(n508), .Q(n506) );
  OR2X1 U651 ( .IN1(n509), .IN2(n510), .Q(n508) );
  AND2X1 U652 ( .IN1(n503), .IN2(iXMIT_xmit_ShiftRegH_6_), .Q(n510) );
  AND2X1 U653 ( .IN1(n499), .IN2(iXMIT_xmit_ShiftRegH_7_), .Q(n509) );
  AND2X1 U654 ( .IN1(xmit_dataH_6_), .IN2(n511), .Q(n507) );
  AND2X1 U655 ( .IN1(test_se), .IN2(iXMIT_xmit_ShiftRegH_5_), .Q(n504) );
  OR2X1 U656 ( .IN1(n512), .IN2(n513), .Q(n171) );
  AND2X1 U657 ( .IN1(n514), .IN2(n445), .Q(n513) );
  OR2X1 U658 ( .IN1(n515), .IN2(n516), .Q(n514) );
  OR2X1 U659 ( .IN1(n517), .IN2(n518), .Q(n516) );
  AND2X1 U660 ( .IN1(n503), .IN2(iXMIT_xmit_ShiftRegH_5_), .Q(n518) );
  AND2X1 U661 ( .IN1(n499), .IN2(iXMIT_xmit_ShiftRegH_6_), .Q(n517) );
  AND2X1 U662 ( .IN1(xmit_dataH_5_), .IN2(n511), .Q(n515) );
  AND2X1 U663 ( .IN1(n729), .IN2(test_se), .Q(n512) );
  OR2X1 U664 ( .IN1(n519), .IN2(n520), .Q(n170) );
  AND2X1 U665 ( .IN1(n521), .IN2(n445), .Q(n520) );
  OR2X1 U666 ( .IN1(n522), .IN2(n523), .Q(n521) );
  OR2X1 U667 ( .IN1(n524), .IN2(n525), .Q(n523) );
  AND2X1 U668 ( .IN1(n729), .IN2(n503), .Q(n525) );
  AND2X1 U669 ( .IN1(n499), .IN2(iXMIT_xmit_ShiftRegH_5_), .Q(n524) );
  AND2X1 U670 ( .IN1(xmit_dataH_4_), .IN2(n511), .Q(n522) );
  AND2X1 U671 ( .IN1(n730), .IN2(test_se), .Q(n519) );
  OR2X1 U672 ( .IN1(n526), .IN2(n527), .Q(n169) );
  AND2X1 U673 ( .IN1(n528), .IN2(n445), .Q(n527) );
  OR2X1 U674 ( .IN1(n529), .IN2(n530), .Q(n528) );
  OR2X1 U675 ( .IN1(n531), .IN2(n532), .Q(n530) );
  AND2X1 U676 ( .IN1(n730), .IN2(n503), .Q(n532) );
  AND2X1 U677 ( .IN1(n729), .IN2(n499), .Q(n531) );
  AND2X1 U678 ( .IN1(xmit_dataH_3_), .IN2(n511), .Q(n529) );
  AND2X1 U679 ( .IN1(n731), .IN2(test_se), .Q(n526) );
  OR2X1 U680 ( .IN1(n533), .IN2(n534), .Q(n168) );
  AND2X1 U681 ( .IN1(n535), .IN2(n445), .Q(n534) );
  OR2X1 U682 ( .IN1(n536), .IN2(n537), .Q(n535) );
  OR2X1 U683 ( .IN1(n538), .IN2(n539), .Q(n537) );
  AND2X1 U684 ( .IN1(n731), .IN2(n503), .Q(n539) );
  AND2X1 U685 ( .IN1(n730), .IN2(n499), .Q(n538) );
  AND2X1 U686 ( .IN1(xmit_dataH_2_), .IN2(n511), .Q(n536) );
  AND2X1 U687 ( .IN1(n732), .IN2(test_se), .Q(n533) );
  OR2X1 U688 ( .IN1(n540), .IN2(n541), .Q(n167) );
  AND2X1 U689 ( .IN1(n542), .IN2(n445), .Q(n541) );
  OR2X1 U690 ( .IN1(n543), .IN2(n544), .Q(n542) );
  OR2X1 U691 ( .IN1(n545), .IN2(n546), .Q(n544) );
  AND2X1 U692 ( .IN1(n732), .IN2(n503), .Q(n546) );
  AND2X1 U693 ( .IN1(n731), .IN2(n499), .Q(n545) );
  AND2X1 U694 ( .IN1(xmit_dataH_1_), .IN2(n511), .Q(n543) );
  AND2X1 U695 ( .IN1(test_se), .IN2(n427), .Q(n540) );
  OR2X1 U696 ( .IN1(n547), .IN2(n548), .Q(n166) );
  AND2X1 U697 ( .IN1(n549), .IN2(n445), .Q(n548) );
  OR2X1 U698 ( .IN1(n550), .IN2(n487), .Q(n549) );
  AND2X1 U699 ( .IN1(n438), .IN2(n551), .Q(n487) );
  INVX0 U700 ( .INP(xmitH), .ZN(n551) );
  AND2X1 U701 ( .IN1(n453), .IN2(n437), .Q(n550) );
  AND2X1 U702 ( .IN1(n552), .IN2(n740), .Q(n453) );
  AND2X1 U703 ( .IN1(test_se), .IN2(iXMIT_xmit_ShiftRegH_7_), .Q(n547) );
  OR2X1 U704 ( .IN1(n553), .IN2(n554), .Q(n164) );
  OR2X1 U705 ( .IN1(n555), .IN2(n556), .Q(n554) );
  AND2X1 U706 ( .IN1(n557), .IN2(n245), .Q(n556) );
  AND2X1 U707 ( .IN1(n558), .IN2(n445), .Q(n557) );
  OR2X1 U708 ( .IN1(n559), .IN2(n429), .Q(n558) );
  AND2X1 U709 ( .IN1(n560), .IN2(iRECEIVER_state_1_), .Q(n559) );
  AND2X1 U710 ( .IN1(n561), .IN2(iRECEIVER_state_0_), .Q(n555) );
  OR2X1 U711 ( .IN1(test_se), .IN2(n562), .Q(n561) );
  OR2X1 U712 ( .IN1(n563), .IN2(n564), .Q(n562) );
  AND2X1 U713 ( .IN1(n565), .IN2(n241), .Q(n564) );
  AND2X1 U714 ( .IN1(n238), .IN2(n429), .Q(n565) );
  AND2X1 U715 ( .IN1(n566), .IN2(iRECEIVER_state_1_), .Q(n563) );
  OR2X1 U716 ( .IN1(n567), .IN2(n568), .Q(n163) );
  AND2X1 U717 ( .IN1(n569), .IN2(n445), .Q(n568) );
  OR2X1 U718 ( .IN1(iRECEIVER_state_2_), .IN2(n570), .Q(n569) );
  OR2X1 U719 ( .IN1(n571), .IN2(n572), .Q(n570) );
  AND2X1 U720 ( .IN1(n573), .IN2(iRECEIVER_state_1_), .Q(n572) );
  OR2X1 U721 ( .IN1(n574), .IN2(n575), .Q(n573) );
  AND2X1 U722 ( .IN1(n576), .IN2(iRECEIVER_state_0_), .Q(n574) );
  OR2X1 U723 ( .IN1(n577), .IN2(n566), .Q(n576) );
  INVX0 U724 ( .INP(n578), .ZN(n566) );
  AND2X1 U725 ( .IN1(n579), .IN2(n580), .Q(n577) );
  AND2X1 U726 ( .IN1(n423), .IN2(n426), .Q(n580) );
  AND2X1 U727 ( .IN1(n735), .IN2(n428), .Q(n579) );
  AND2X1 U728 ( .IN1(n241), .IN2(n734), .Q(n571) );
  AND2X1 U729 ( .IN1(n735), .IN2(test_se), .Q(n567) );
  OR2X1 U730 ( .IN1(n581), .IN2(n582), .Q(n162) );
  AND2X1 U731 ( .IN1(test_si), .IN2(test_se), .Q(n582) );
  AND2X1 U732 ( .IN1(iRECEIVER_N20), .IN2(n445), .Q(n581) );
  OR2X1 U733 ( .IN1(n583), .IN2(n584), .Q(n161) );
  AND2X1 U734 ( .IN1(iRECEIVER_N21), .IN2(n445), .Q(n584) );
  AND2X1 U735 ( .IN1(test_se), .IN2(iRECEIVER_bitCell_cntrH_0_), .Q(n583) );
  OR2X1 U736 ( .IN1(n585), .IN2(n586), .Q(n160) );
  AND2X1 U737 ( .IN1(iRECEIVER_N22), .IN2(n445), .Q(n586) );
  AND2X1 U738 ( .IN1(test_se), .IN2(iRECEIVER_bitCell_cntrH_1_), .Q(n585) );
  OR2X1 U739 ( .IN1(n587), .IN2(n588), .Q(n159) );
  AND2X1 U740 ( .IN1(n748), .IN2(test_se), .Q(n588) );
  AND2X1 U741 ( .IN1(iRECEIVER_N23), .IN2(n445), .Q(n587) );
  OR2X1 U742 ( .IN1(n589), .IN2(iRECEIVER_next_state_2_), .Q(n157) );
  AND2X1 U743 ( .IN1(test_se), .IN2(iRECEIVER_state_1_), .Q(n589) );
  OR2X1 U744 ( .IN1(n590), .IN2(n591), .Q(n156) );
  AND2X1 U745 ( .IN1(n592), .IN2(n445), .Q(n591) );
  OR2X1 U746 ( .IN1(n593), .IN2(n594), .Q(n592) );
  AND2X1 U747 ( .IN1(iRECEIVER_state_2_), .IN2(iRECEIVER_state_0_), .Q(n593)
         );
  AND2X1 U748 ( .IN1(n733), .IN2(test_se), .Q(n590) );
  OR2X1 U749 ( .IN1(n595), .IN2(n596), .Q(n155) );
  OR2X1 U750 ( .IN1(n597), .IN2(n598), .Q(n596) );
  AND2X1 U751 ( .IN1(n553), .IN2(n734), .Q(n598) );
  AND2X1 U752 ( .IN1(rec_dataH_rec_7), .IN2(n599), .Q(n597) );
  AND2X1 U753 ( .IN1(rec_dataH_rec_6), .IN2(test_se), .Q(n595) );
  OR2X1 U754 ( .IN1(n600), .IN2(n601), .Q(n154) );
  AND2X1 U755 ( .IN1(rec_dataH_temp_6), .IN2(test_se), .Q(n601) );
  AND2X1 U756 ( .IN1(rec_dataH_rec_7), .IN2(n445), .Q(n600) );
  OR2X1 U757 ( .IN1(n602), .IN2(n603), .Q(n153) );
  AND2X1 U758 ( .IN1(rec_dataH_6_), .IN2(test_se), .Q(n603) );
  AND2X1 U759 ( .IN1(test_so), .IN2(n445), .Q(n602) );
  OR2X1 U760 ( .IN1(n604), .IN2(n605), .Q(n152) );
  OR2X1 U761 ( .IN1(n606), .IN2(n607), .Q(n605) );
  AND2X1 U762 ( .IN1(n553), .IN2(rec_dataH_rec_7), .Q(n607) );
  AND2X1 U763 ( .IN1(rec_dataH_rec_6), .IN2(n599), .Q(n606) );
  AND2X1 U764 ( .IN1(rec_dataH_rec_5), .IN2(test_se), .Q(n604) );
  OR2X1 U765 ( .IN1(n608), .IN2(n609), .Q(n150) );
  AND2X1 U766 ( .IN1(rec_dataH_temp_5), .IN2(test_se), .Q(n609) );
  AND2X1 U767 ( .IN1(rec_dataH_rec_6), .IN2(n445), .Q(n608) );
  OR2X1 U768 ( .IN1(n610), .IN2(n611), .Q(n149) );
  AND2X1 U769 ( .IN1(rec_dataH_5_), .IN2(test_se), .Q(n611) );
  AND2X1 U770 ( .IN1(rec_dataH_temp_6), .IN2(n445), .Q(n610) );
  OR2X1 U771 ( .IN1(n612), .IN2(n613), .Q(n148) );
  OR2X1 U772 ( .IN1(n614), .IN2(n615), .Q(n613) );
  AND2X1 U773 ( .IN1(rec_dataH_rec_6), .IN2(n553), .Q(n615) );
  AND2X1 U774 ( .IN1(rec_dataH_rec_5), .IN2(n599), .Q(n614) );
  AND2X1 U775 ( .IN1(rec_dataH_rec_4), .IN2(test_se), .Q(n612) );
  OR2X1 U776 ( .IN1(n616), .IN2(n617), .Q(n147) );
  AND2X1 U777 ( .IN1(rec_dataH_temp_4), .IN2(test_se), .Q(n617) );
  AND2X1 U778 ( .IN1(rec_dataH_rec_5), .IN2(n445), .Q(n616) );
  OR2X1 U779 ( .IN1(n618), .IN2(n619), .Q(n146) );
  AND2X1 U780 ( .IN1(rec_dataH_4_), .IN2(test_se), .Q(n619) );
  AND2X1 U781 ( .IN1(rec_dataH_temp_5), .IN2(n445), .Q(n618) );
  OR2X1 U782 ( .IN1(n620), .IN2(n621), .Q(n145) );
  OR2X1 U783 ( .IN1(n622), .IN2(n623), .Q(n621) );
  AND2X1 U784 ( .IN1(rec_dataH_rec_5), .IN2(n553), .Q(n623) );
  AND2X1 U785 ( .IN1(rec_dataH_rec_4), .IN2(n599), .Q(n622) );
  AND2X1 U786 ( .IN1(rec_dataH_rec_3), .IN2(test_se), .Q(n620) );
  OR2X1 U787 ( .IN1(n624), .IN2(n625), .Q(n143) );
  AND2X1 U788 ( .IN1(rec_dataH_temp_3), .IN2(test_se), .Q(n625) );
  AND2X1 U789 ( .IN1(rec_dataH_rec_4), .IN2(n445), .Q(n624) );
  OR2X1 U790 ( .IN1(n626), .IN2(n627), .Q(n142) );
  AND2X1 U791 ( .IN1(rec_dataH_3_), .IN2(test_se), .Q(n627) );
  AND2X1 U792 ( .IN1(rec_dataH_temp_4), .IN2(n445), .Q(n626) );
  OR2X1 U793 ( .IN1(n628), .IN2(n629), .Q(n141) );
  OR2X1 U794 ( .IN1(n630), .IN2(n631), .Q(n629) );
  AND2X1 U795 ( .IN1(rec_dataH_rec_4), .IN2(n553), .Q(n631) );
  AND2X1 U796 ( .IN1(rec_dataH_rec_3), .IN2(n599), .Q(n630) );
  AND2X1 U797 ( .IN1(rec_dataH_rec_2), .IN2(test_se), .Q(n628) );
  OR2X1 U798 ( .IN1(n632), .IN2(n633), .Q(n140) );
  AND2X1 U799 ( .IN1(rec_dataH_temp_2), .IN2(test_se), .Q(n633) );
  AND2X1 U800 ( .IN1(rec_dataH_rec_3), .IN2(n445), .Q(n632) );
  OR2X1 U801 ( .IN1(n634), .IN2(n635), .Q(n139) );
  AND2X1 U802 ( .IN1(rec_dataH_2_), .IN2(test_se), .Q(n635) );
  AND2X1 U803 ( .IN1(rec_dataH_temp_3), .IN2(n445), .Q(n634) );
  OR2X1 U804 ( .IN1(n636), .IN2(n637), .Q(n138) );
  OR2X1 U805 ( .IN1(n638), .IN2(n639), .Q(n637) );
  AND2X1 U806 ( .IN1(rec_dataH_rec_3), .IN2(n553), .Q(n639) );
  AND2X1 U807 ( .IN1(rec_dataH_rec_2), .IN2(n599), .Q(n638) );
  AND2X1 U808 ( .IN1(rec_dataH_rec_1), .IN2(test_se), .Q(n636) );
  OR2X1 U809 ( .IN1(n640), .IN2(n641), .Q(n136) );
  AND2X1 U810 ( .IN1(rec_dataH_temp_1), .IN2(test_se), .Q(n641) );
  AND2X1 U811 ( .IN1(rec_dataH_rec_2), .IN2(n445), .Q(n640) );
  OR2X1 U812 ( .IN1(n642), .IN2(n643), .Q(n135) );
  AND2X1 U813 ( .IN1(rec_dataH_1_), .IN2(test_se), .Q(n643) );
  AND2X1 U814 ( .IN1(rec_dataH_temp_2), .IN2(n445), .Q(n642) );
  OR2X1 U815 ( .IN1(n644), .IN2(n645), .Q(n134) );
  OR2X1 U816 ( .IN1(n646), .IN2(n647), .Q(n645) );
  AND2X1 U817 ( .IN1(rec_dataH_rec_2), .IN2(n553), .Q(n647) );
  AND2X1 U818 ( .IN1(rec_dataH_rec_1), .IN2(n599), .Q(n646) );
  AND2X1 U819 ( .IN1(rec_dataH_rec_0), .IN2(test_se), .Q(n644) );
  OR2X1 U820 ( .IN1(n648), .IN2(n649), .Q(n133) );
  AND2X1 U821 ( .IN1(rec_dataH_temp_0), .IN2(test_se), .Q(n649) );
  AND2X1 U822 ( .IN1(rec_dataH_rec_1), .IN2(n445), .Q(n648) );
  OR2X1 U823 ( .IN1(n650), .IN2(n651), .Q(n132) );
  AND2X1 U824 ( .IN1(rec_dataH_0_), .IN2(test_se), .Q(n651) );
  AND2X1 U825 ( .IN1(rec_dataH_temp_1), .IN2(n445), .Q(n650) );
  OR2X1 U826 ( .IN1(n652), .IN2(n653), .Q(n131) );
  OR2X1 U827 ( .IN1(n654), .IN2(n655), .Q(n653) );
  AND2X1 U828 ( .IN1(rec_dataH_rec_1), .IN2(n553), .Q(n655) );
  AND2X1 U829 ( .IN1(rec_dataH_rec_0), .IN2(n599), .Q(n654) );
  AND2X1 U830 ( .IN1(n747), .IN2(test_se), .Q(n652) );
  OR2X1 U831 ( .IN1(n656), .IN2(n657), .Q(n129) );
  AND2X1 U832 ( .IN1(rec_dataH_7_), .IN2(test_se), .Q(n657) );
  AND2X1 U833 ( .IN1(rec_dataH_rec_0), .IN2(n445), .Q(n656) );
  OR2X1 U834 ( .IN1(n658), .IN2(n659), .Q(n128) );
  AND2X1 U835 ( .IN1(xmit_doneH_temp), .IN2(test_se), .Q(n659) );
  AND2X1 U836 ( .IN1(rec_dataH_temp_0), .IN2(n445), .Q(n658) );
  OR2X1 U837 ( .IN1(n660), .IN2(n661), .Q(n127) );
  AND2X1 U838 ( .IN1(n735), .IN2(n662), .Q(n661) );
  OR2X1 U839 ( .IN1(n663), .IN2(n664), .Q(n662) );
  AND2X1 U840 ( .IN1(n553), .IN2(n665), .Q(n663) );
  OR2X1 U841 ( .IN1(n666), .IN2(n426), .Q(n665) );
  AND2X1 U842 ( .IN1(n744), .IN2(n667), .Q(n660) );
  OR2X1 U843 ( .IN1(n668), .IN2(test_se), .Q(n667) );
  AND2X1 U844 ( .IN1(n669), .IN2(n670), .Q(n668) );
  AND2X1 U845 ( .IN1(n553), .IN2(n434), .Q(n669) );
  OR2X1 U846 ( .IN1(n671), .IN2(n672), .Q(n126) );
  OR2X1 U847 ( .IN1(n673), .IN2(n674), .Q(n672) );
  AND2X1 U848 ( .IN1(n664), .IN2(n745), .Q(n674) );
  AND2X1 U849 ( .IN1(n553), .IN2(n423), .Q(n673) );
  AND2X1 U850 ( .IN1(test_se), .IN2(rec_readyH), .Q(n671) );
  OR2X1 U851 ( .IN1(n675), .IN2(n676), .Q(n125) );
  OR2X1 U852 ( .IN1(n677), .IN2(n678), .Q(n676) );
  AND2X1 U853 ( .IN1(n664), .IN2(n746), .Q(n678) );
  AND2X1 U854 ( .IN1(n553), .IN2(iRECEIVER_N26), .Q(n677) );
  AND2X1 U855 ( .IN1(n745), .IN2(test_se), .Q(n675) );
  OR2X1 U856 ( .IN1(n679), .IN2(n680), .Q(n124) );
  OR2X1 U857 ( .IN1(n681), .IN2(n682), .Q(n680) );
  AND2X1 U858 ( .IN1(n664), .IN2(n744), .Q(n682) );
  AND2X1 U859 ( .IN1(n683), .IN2(n599), .Q(n664) );
  AND2X1 U860 ( .IN1(n684), .IN2(n445), .Q(n599) );
  OR2X1 U861 ( .IN1(iRECEIVER_state_0_), .IN2(n238), .Q(n684) );
  INVX0 U862 ( .INP(n594), .ZN(n683) );
  AND2X1 U863 ( .IN1(n241), .IN2(n685), .Q(n594) );
  AND2X1 U864 ( .IN1(n734), .IN2(n238), .Q(n685) );
  AND2X1 U865 ( .IN1(n553), .IN2(iRECEIVER_N27), .Q(n681) );
  AND2X1 U866 ( .IN1(n245), .IN2(n686), .Q(n553) );
  AND2X1 U867 ( .IN1(n445), .IN2(iRECEIVER_state_2_), .Q(n686) );
  AND2X1 U868 ( .IN1(n746), .IN2(test_se), .Q(n679) );
  OR2X1 U869 ( .IN1(n687), .IN2(n688), .Q(n122) );
  AND2X1 U870 ( .IN1(test_se), .IN2(n741), .Q(n688) );
  AND2X1 U871 ( .IN1(iXMIT_N29), .IN2(n445), .Q(n687) );
  OR2X1 U872 ( .IN1(n689), .IN2(n690), .Q(n121) );
  AND2X1 U873 ( .IN1(iXMIT_N26), .IN2(n445), .Q(n690) );
  AND2X1 U874 ( .IN1(test_se), .IN2(iRECEIVER_state_2_), .Q(n689) );
  OR2X1 U875 ( .IN1(n691), .IN2(n692), .Q(n120) );
  AND2X1 U876 ( .IN1(test_se), .IN2(n743), .Q(n692) );
  AND2X1 U877 ( .IN1(iXMIT_N27), .IN2(n445), .Q(n691) );
  OR2X1 U878 ( .IN1(n693), .IN2(n694), .Q(n119) );
  AND2X1 U879 ( .IN1(n695), .IN2(n445), .Q(n694) );
  OR2X1 U880 ( .IN1(n696), .IN2(n697), .Q(n695) );
  OR2X1 U881 ( .IN1(n698), .IN2(n699), .Q(n697) );
  AND2X1 U882 ( .IN1(n503), .IN2(n427), .Q(n699) );
  INVX0 U883 ( .INP(n467), .ZN(n503) );
  AND2X1 U884 ( .IN1(n732), .IN2(n499), .Q(n698) );
  AND2X1 U885 ( .IN1(n700), .IN2(n467), .Q(n499) );
  OR2X1 U886 ( .IN1(n701), .IN2(n511), .Q(n467) );
  AND2X1 U887 ( .IN1(n239), .IN2(iXMIT_state_2_), .Q(n701) );
  INVX0 U888 ( .INP(n511), .ZN(n700) );
  AND2X1 U889 ( .IN1(xmit_dataH_0_), .IN2(n511), .Q(n696) );
  AND2X1 U890 ( .IN1(n438), .IN2(xmitH), .Q(n511) );
  AND2X1 U891 ( .IN1(n242), .IN2(n246), .Q(n438) );
  AND2X1 U892 ( .IN1(test_se), .IN2(iXMIT_state_2_), .Q(n693) );
  OR2X1 U893 ( .IN1(n702), .IN2(n703), .Q(n118) );
  AND2X1 U894 ( .IN1(n734), .IN2(test_se), .Q(n703) );
  AND2X1 U895 ( .IN1(uart_REC_dataH), .IN2(n445), .Q(n702) );
  OR2X1 U896 ( .IN1(n704), .IN2(n705), .Q(n117) );
  AND2X1 U897 ( .IN1(rec_dataH_rec_7), .IN2(test_se), .Q(n705) );
  AND2X1 U898 ( .IN1(n733), .IN2(n445), .Q(n704) );
  INVX0 U899 ( .INP(test_se), .ZN(n445) );
  XOR2X1 U900 ( .IN1(n736), .IN2(n706), .Q(iXMIT_N46) );
  AND2X1 U901 ( .IN1(n707), .IN2(n737), .Q(n706) );
  XOR2X1 U902 ( .IN1(n737), .IN2(n707), .Q(iXMIT_N45) );
  AND2X1 U903 ( .IN1(n738), .IN2(n739), .Q(n707) );
  XNOR2X1 U904 ( .IN1(n431), .IN2(n738), .Q(iXMIT_N44) );
  AND2X1 U905 ( .IN1(n708), .IN2(iXMIT_N25), .Q(iXMIT_N29) );
  AND2X1 U906 ( .IN1(n708), .IN2(iXMIT_N24), .Q(iXMIT_N28) );
  OR2X1 U907 ( .IN1(n709), .IN2(n710), .Q(iXMIT_N27) );
  AND2X1 U908 ( .IN1(iXMIT_N26), .IN2(n742), .Q(n710) );
  AND2X1 U909 ( .IN1(n711), .IN2(n430), .Q(n709) );
  AND2X1 U910 ( .IN1(n743), .IN2(n708), .Q(n711) );
  AND2X1 U911 ( .IN1(n433), .IN2(n708), .Q(iXMIT_N26) );
  OR2X1 U912 ( .IN1(n437), .IN2(n466), .Q(n708) );
  AND2X1 U913 ( .IN1(n462), .IN2(iXMIT_state_1_), .Q(n466) );
  OR2X1 U914 ( .IN1(n239), .IN2(n493), .Q(n462) );
  OR2X1 U915 ( .IN1(n712), .IN2(n713), .Q(n493) );
  INVX0 U916 ( .INP(n714), .ZN(n713) );
  AND2X1 U917 ( .IN1(n741), .IN2(n740), .Q(n714) );
  OR2X1 U918 ( .IN1(n743), .IN2(n430), .Q(n712) );
  AND2X1 U919 ( .IN1(iXMIT_state_2_), .IN2(iXMIT_state_0_), .Q(n437) );
  XOR2X1 U920 ( .IN1(n740), .IN2(n552), .Q(iXMIT_N25) );
  AND2X1 U921 ( .IN1(n715), .IN2(n741), .Q(n552) );
  XOR2X1 U922 ( .IN1(n741), .IN2(n715), .Q(iXMIT_N24) );
  AND2X1 U923 ( .IN1(n743), .IN2(n742), .Q(n715) );
  AND2X1 U924 ( .IN1(n578), .IN2(n716), .Q(iRECEIVER_next_state_2_) );
  AND2X1 U925 ( .IN1(iRECEIVER_state_0_), .IN2(iRECEIVER_state_1_), .Q(n716)
         );
  XNOR2X1 U926 ( .IN1(n426), .IN2(n670), .Q(iRECEIVER_N27) );
  INVX0 U927 ( .INP(n666), .ZN(n670) );
  OR2X1 U928 ( .IN1(n428), .IN2(n423), .Q(n666) );
  XNOR2X1 U929 ( .IN1(n746), .IN2(n423), .Q(iRECEIVER_N26) );
  AND2X1 U930 ( .IN1(iRECEIVER_N19), .IN2(n717), .Q(iRECEIVER_N23) );
  AND2X1 U931 ( .IN1(iRECEIVER_N18), .IN2(n717), .Q(iRECEIVER_N22) );
  AND2X1 U932 ( .IN1(iRECEIVER_N17), .IN2(n717), .Q(iRECEIVER_N21) );
  AND2X1 U933 ( .IN1(n255), .IN2(n717), .Q(iRECEIVER_N20) );
  INVX0 U934 ( .INP(n718), .ZN(n717) );
  OR2X1 U935 ( .IN1(n719), .IN2(n720), .Q(n718) );
  OR2X1 U936 ( .IN1(n241), .IN2(iRECEIVER_state_2_), .Q(n720) );
  OR2X1 U937 ( .IN1(n721), .IN2(n722), .Q(n719) );
  AND2X1 U938 ( .IN1(n575), .IN2(n245), .Q(n722) );
  INVX0 U939 ( .INP(n560), .ZN(n575) );
  OR2X1 U940 ( .IN1(n723), .IN2(n724), .Q(n560) );
  OR2X1 U941 ( .IN1(iRECEIVER_bitCell_cntrH_0_), .IN2(n424), .Q(n724) );
  OR2X1 U942 ( .IN1(n747), .IN2(iRECEIVER_bitCell_cntrH_1_), .Q(n723) );
  AND2X1 U943 ( .IN1(n578), .IN2(iRECEIVER_state_0_), .Q(n721) );
  AND2X1 U944 ( .IN1(n725), .IN2(n726), .Q(n578) );
  AND2X1 U945 ( .IN1(n748), .IN2(n747), .Q(n726) );
  AND2X1 U946 ( .IN1(iRECEIVER_bitCell_cntrH_1_), .IN2(n255), .Q(n725) );
  XNOR2X1 U947 ( .IN1(n727), .IN2(n747), .Q(iRECEIVER_N19) );
  OR2X1 U948 ( .IN1(n424), .IN2(n728), .Q(n727) );
  XOR2X1 U949 ( .IN1(n728), .IN2(n424), .Q(iRECEIVER_N18) );
  OR2X1 U950 ( .IN1(n244), .IN2(n255), .Q(n728) );
  XNOR2X1 U951 ( .IN1(n244), .IN2(iRECEIVER_bitCell_cntrH_0_), .Q(
        iRECEIVER_N17) );
endmodule

