module add_mul_comp_8_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, Result_0_, Result_1_, 
        Result_2_, Result_3_, Result_4_, Result_5_, Result_6_, Result_7_, 
        Result_8_, Result_9_, Result_10_, Result_11_, Result_12_, Result_13_, 
        Result_14_, Result_15_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_,
         b_4_, b_5_, b_6_, b_7_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_;
  wire   n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001;

  NAND2_X1 U489 ( .A1(n473), .A2(n474), .ZN(Result_9_) );
  NAND2_X1 U490 ( .A1(n475), .A2(n476), .ZN(n474) );
  XNOR2_X1 U491 ( .A(n477), .B(n478), .ZN(n475) );
  XNOR2_X1 U492 ( .A(n479), .B(n480), .ZN(n478) );
  NAND2_X1 U493 ( .A1(n481), .A2(n482), .ZN(n473) );
  NAND2_X1 U494 ( .A1(n483), .A2(n484), .ZN(n482) );
  NAND2_X1 U495 ( .A1(n485), .A2(n486), .ZN(n484) );
  OR2_X1 U496 ( .A1(n487), .A2(n488), .ZN(n485) );
  NAND2_X1 U497 ( .A1(n489), .A2(n490), .ZN(n483) );
  XOR2_X1 U498 ( .A(b_1_), .B(a_1_), .Z(n489) );
  NAND2_X1 U499 ( .A1(n491), .A2(n492), .ZN(Result_8_) );
  NAND2_X1 U500 ( .A1(n493), .A2(n476), .ZN(n492) );
  XOR2_X1 U501 ( .A(n494), .B(n495), .Z(n493) );
  XOR2_X1 U502 ( .A(n496), .B(n497), .Z(n494) );
  NAND2_X1 U503 ( .A1(n498), .A2(n481), .ZN(n491) );
  XNOR2_X1 U504 ( .A(n499), .B(n500), .ZN(n498) );
  NOR2_X1 U505 ( .A1(n488), .A2(n501), .ZN(n499) );
  NOR2_X1 U506 ( .A1(n487), .A2(n486), .ZN(n501) );
  INV_X1 U507 ( .A(n490), .ZN(n486) );
  NOR2_X1 U508 ( .A1(n502), .A2(n503), .ZN(n490) );
  NOR2_X1 U509 ( .A1(n504), .A2(n505), .ZN(n503) );
  INV_X1 U510 ( .A(n506), .ZN(n487) );
  NOR2_X1 U511 ( .A1(b_1_), .A2(a_1_), .ZN(n488) );
  NOR2_X1 U512 ( .A1(n481), .A2(n507), .ZN(Result_7_) );
  XNOR2_X1 U513 ( .A(n508), .B(n509), .ZN(n507) );
  NOR2_X1 U514 ( .A1(n510), .A2(n511), .ZN(Result_6_) );
  NAND2_X1 U515 ( .A1(n512), .A2(n476), .ZN(n511) );
  NOR2_X1 U516 ( .A1(n513), .A2(n514), .ZN(n510) );
  NOR2_X1 U517 ( .A1(n481), .A2(n515), .ZN(Result_5_) );
  XOR2_X1 U518 ( .A(n512), .B(n516), .Z(n515) );
  NOR2_X1 U519 ( .A1(n517), .A2(n518), .ZN(n516) );
  NOR2_X1 U520 ( .A1(n519), .A2(n520), .ZN(n518) );
  NOR2_X1 U521 ( .A1(n481), .A2(n521), .ZN(Result_4_) );
  XNOR2_X1 U522 ( .A(n522), .B(n523), .ZN(n521) );
  NOR2_X1 U523 ( .A1(n481), .A2(n524), .ZN(Result_3_) );
  XNOR2_X1 U524 ( .A(n525), .B(n526), .ZN(n524) );
  AND2_X1 U525 ( .A1(n527), .A2(n528), .ZN(n526) );
  NOR2_X1 U526 ( .A1(n481), .A2(n529), .ZN(Result_2_) );
  XOR2_X1 U527 ( .A(n530), .B(n531), .Z(n529) );
  NAND2_X1 U528 ( .A1(n532), .A2(n533), .ZN(n531) );
  NOR2_X1 U529 ( .A1(n481), .A2(n534), .ZN(Result_1_) );
  XOR2_X1 U530 ( .A(n535), .B(n536), .Z(n534) );
  NAND2_X1 U531 ( .A1(n537), .A2(n538), .ZN(n536) );
  NAND2_X1 U532 ( .A1(n539), .A2(n540), .ZN(n538) );
  NAND2_X1 U533 ( .A1(n541), .A2(n542), .ZN(Result_15_) );
  NAND2_X1 U534 ( .A1(n543), .A2(n476), .ZN(n542) );
  NAND2_X1 U535 ( .A1(n481), .A2(n544), .ZN(n541) );
  NAND2_X1 U536 ( .A1(n545), .A2(n546), .ZN(n544) );
  NAND2_X1 U537 ( .A1(b_7_), .A2(n547), .ZN(n546) );
  NAND2_X1 U538 ( .A1(n548), .A2(n549), .ZN(Result_14_) );
  NAND2_X1 U539 ( .A1(n481), .A2(n550), .ZN(n549) );
  NAND2_X1 U540 ( .A1(n551), .A2(n552), .ZN(n550) );
  NOR2_X1 U541 ( .A1(n553), .A2(n554), .ZN(n551) );
  NOR2_X1 U542 ( .A1(n555), .A2(n556), .ZN(n554) );
  NAND2_X1 U543 ( .A1(n557), .A2(n558), .ZN(n556) );
  NOR2_X1 U544 ( .A1(b_6_), .A2(n559), .ZN(n553) );
  XOR2_X1 U545 ( .A(n557), .B(a_6_), .Z(n559) );
  NAND2_X1 U546 ( .A1(n560), .A2(n476), .ZN(n548) );
  XOR2_X1 U547 ( .A(n561), .B(n562), .Z(n560) );
  NAND2_X1 U548 ( .A1(b_7_), .A2(a_6_), .ZN(n562) );
  NAND2_X1 U549 ( .A1(n563), .A2(n564), .ZN(Result_13_) );
  NAND2_X1 U550 ( .A1(n481), .A2(n565), .ZN(n564) );
  NAND2_X1 U551 ( .A1(n566), .A2(n567), .ZN(n565) );
  NAND2_X1 U552 ( .A1(n568), .A2(n569), .ZN(n567) );
  NOR2_X1 U553 ( .A1(n570), .A2(n571), .ZN(n566) );
  NOR2_X1 U554 ( .A1(b_5_), .A2(n572), .ZN(n571) );
  XOR2_X1 U555 ( .A(a_5_), .B(n573), .Z(n572) );
  NOR2_X1 U556 ( .A1(n574), .A2(n575), .ZN(n570) );
  NAND2_X1 U557 ( .A1(n573), .A2(n576), .ZN(n575) );
  INV_X1 U558 ( .A(n569), .ZN(n573) );
  NAND2_X1 U559 ( .A1(n577), .A2(n476), .ZN(n563) );
  XNOR2_X1 U560 ( .A(n578), .B(n579), .ZN(n577) );
  XOR2_X1 U561 ( .A(n580), .B(n581), .Z(n579) );
  NAND2_X1 U562 ( .A1(b_7_), .A2(a_5_), .ZN(n580) );
  NAND2_X1 U563 ( .A1(n582), .A2(n583), .ZN(Result_12_) );
  NAND2_X1 U564 ( .A1(n584), .A2(n476), .ZN(n583) );
  XNOR2_X1 U565 ( .A(n585), .B(n586), .ZN(n584) );
  NAND2_X1 U566 ( .A1(n587), .A2(n588), .ZN(n585) );
  NAND2_X1 U567 ( .A1(n481), .A2(n589), .ZN(n582) );
  XNOR2_X1 U568 ( .A(n590), .B(n591), .ZN(n589) );
  NAND2_X1 U569 ( .A1(n592), .A2(n593), .ZN(n590) );
  NAND2_X1 U570 ( .A1(n594), .A2(n595), .ZN(Result_11_) );
  NAND2_X1 U571 ( .A1(n481), .A2(n596), .ZN(n595) );
  NAND2_X1 U572 ( .A1(n597), .A2(n598), .ZN(n596) );
  NAND2_X1 U573 ( .A1(n599), .A2(n600), .ZN(n598) );
  NOR2_X1 U574 ( .A1(n601), .A2(n602), .ZN(n597) );
  NOR2_X1 U575 ( .A1(b_3_), .A2(n603), .ZN(n602) );
  XOR2_X1 U576 ( .A(n604), .B(n600), .Z(n603) );
  NOR2_X1 U577 ( .A1(n605), .A2(n606), .ZN(n601) );
  OR2_X1 U578 ( .A1(n600), .A2(a_3_), .ZN(n606) );
  NAND2_X1 U579 ( .A1(n607), .A2(n476), .ZN(n594) );
  XOR2_X1 U580 ( .A(n608), .B(n609), .Z(n607) );
  XNOR2_X1 U581 ( .A(n610), .B(n611), .ZN(n609) );
  NAND2_X1 U582 ( .A1(b_7_), .A2(a_3_), .ZN(n610) );
  NAND2_X1 U583 ( .A1(n612), .A2(n613), .ZN(Result_10_) );
  NAND2_X1 U584 ( .A1(n614), .A2(n476), .ZN(n613) );
  XOR2_X1 U585 ( .A(n615), .B(n616), .Z(n614) );
  XOR2_X1 U586 ( .A(n617), .B(n618), .Z(n616) );
  NAND2_X1 U587 ( .A1(n481), .A2(n619), .ZN(n612) );
  XNOR2_X1 U588 ( .A(n505), .B(n620), .ZN(n619) );
  NOR2_X1 U589 ( .A1(n504), .A2(n502), .ZN(n620) );
  NOR2_X1 U590 ( .A1(b_2_), .A2(a_2_), .ZN(n504) );
  AND2_X1 U591 ( .A1(n621), .A2(n622), .ZN(n505) );
  NAND2_X1 U592 ( .A1(n623), .A2(n600), .ZN(n622) );
  NAND2_X1 U593 ( .A1(n592), .A2(n624), .ZN(n600) );
  NAND2_X1 U594 ( .A1(n593), .A2(n591), .ZN(n624) );
  NAND2_X1 U595 ( .A1(n625), .A2(n626), .ZN(n591) );
  NAND2_X1 U596 ( .A1(n627), .A2(n569), .ZN(n626) );
  NAND2_X1 U597 ( .A1(n628), .A2(n629), .ZN(n569) );
  NAND2_X1 U598 ( .A1(n543), .A2(n630), .ZN(n629) );
  NAND2_X1 U599 ( .A1(n555), .A2(n558), .ZN(n630) );
  NAND2_X1 U600 ( .A1(n574), .A2(n576), .ZN(n627) );
  NAND2_X1 U601 ( .A1(n631), .A2(n632), .ZN(n593) );
  NAND2_X1 U602 ( .A1(n605), .A2(n604), .ZN(n623) );
  NOR2_X1 U603 ( .A1(n481), .A2(n633), .ZN(Result_0_) );
  NOR2_X1 U604 ( .A1(n634), .A2(n635), .ZN(n633) );
  NAND2_X1 U605 ( .A1(n540), .A2(n636), .ZN(n635) );
  INV_X1 U606 ( .A(n539), .ZN(n636) );
  NOR2_X1 U607 ( .A1(n637), .A2(n638), .ZN(n539) );
  AND2_X1 U608 ( .A1(n535), .A2(n537), .ZN(n634) );
  NAND2_X1 U609 ( .A1(n637), .A2(n639), .ZN(n537) );
  NAND2_X1 U610 ( .A1(b_0_), .A2(n540), .ZN(n639) );
  NAND2_X1 U611 ( .A1(n640), .A2(n641), .ZN(n540) );
  NAND2_X1 U612 ( .A1(n532), .A2(n642), .ZN(n535) );
  NAND2_X1 U613 ( .A1(n533), .A2(n530), .ZN(n642) );
  NAND2_X1 U614 ( .A1(n528), .A2(n643), .ZN(n530) );
  NAND2_X1 U615 ( .A1(n525), .A2(n527), .ZN(n643) );
  NAND2_X1 U616 ( .A1(n644), .A2(n645), .ZN(n527) );
  NAND2_X1 U617 ( .A1(n646), .A2(n647), .ZN(n645) );
  XOR2_X1 U618 ( .A(n648), .B(n649), .Z(n644) );
  AND2_X1 U619 ( .A1(n522), .A2(n523), .ZN(n525) );
  NAND2_X1 U620 ( .A1(n650), .A2(n651), .ZN(n523) );
  NAND2_X1 U621 ( .A1(n652), .A2(n520), .ZN(n651) );
  INV_X1 U622 ( .A(n512), .ZN(n652) );
  NAND2_X1 U623 ( .A1(n513), .A2(n514), .ZN(n512) );
  XOR2_X1 U624 ( .A(n653), .B(n654), .Z(n514) );
  NOR2_X1 U625 ( .A1(n509), .A2(n508), .ZN(n513) );
  XNOR2_X1 U626 ( .A(n655), .B(n656), .ZN(n508) );
  XOR2_X1 U627 ( .A(n657), .B(n658), .Z(n655) );
  AND2_X1 U628 ( .A1(n659), .A2(n660), .ZN(n509) );
  NAND2_X1 U629 ( .A1(n497), .A2(n661), .ZN(n660) );
  OR2_X1 U630 ( .A1(n495), .A2(n496), .ZN(n661) );
  AND2_X1 U631 ( .A1(b_7_), .A2(a_0_), .ZN(n497) );
  NAND2_X1 U632 ( .A1(n495), .A2(n496), .ZN(n659) );
  NAND2_X1 U633 ( .A1(n662), .A2(n663), .ZN(n496) );
  NAND2_X1 U634 ( .A1(n480), .A2(n664), .ZN(n663) );
  NAND2_X1 U635 ( .A1(n479), .A2(n477), .ZN(n664) );
  AND2_X1 U636 ( .A1(b_7_), .A2(a_1_), .ZN(n480) );
  OR2_X1 U637 ( .A1(n477), .A2(n479), .ZN(n662) );
  AND2_X1 U638 ( .A1(n665), .A2(n666), .ZN(n479) );
  NAND2_X1 U639 ( .A1(n618), .A2(n667), .ZN(n666) );
  NAND2_X1 U640 ( .A1(n617), .A2(n615), .ZN(n667) );
  AND2_X1 U641 ( .A1(b_7_), .A2(a_2_), .ZN(n618) );
  OR2_X1 U642 ( .A1(n615), .A2(n617), .ZN(n665) );
  AND2_X1 U643 ( .A1(n668), .A2(n669), .ZN(n617) );
  NAND2_X1 U644 ( .A1(n670), .A2(b_7_), .ZN(n669) );
  NOR2_X1 U645 ( .A1(n671), .A2(n604), .ZN(n670) );
  NOR2_X1 U646 ( .A1(n608), .A2(n611), .ZN(n671) );
  NAND2_X1 U647 ( .A1(n608), .A2(n611), .ZN(n668) );
  NAND2_X1 U648 ( .A1(n587), .A2(n672), .ZN(n611) );
  NAND2_X1 U649 ( .A1(n586), .A2(n588), .ZN(n672) );
  NAND2_X1 U650 ( .A1(n673), .A2(n674), .ZN(n588) );
  NAND2_X1 U651 ( .A1(b_7_), .A2(a_4_), .ZN(n674) );
  INV_X1 U652 ( .A(n675), .ZN(n673) );
  XNOR2_X1 U653 ( .A(n676), .B(n677), .ZN(n586) );
  NAND2_X1 U654 ( .A1(n678), .A2(n679), .ZN(n676) );
  NAND2_X1 U655 ( .A1(a_4_), .A2(n675), .ZN(n587) );
  NAND2_X1 U656 ( .A1(n680), .A2(n681), .ZN(n675) );
  NAND2_X1 U657 ( .A1(n682), .A2(b_7_), .ZN(n681) );
  NOR2_X1 U658 ( .A1(n683), .A2(n576), .ZN(n682) );
  NOR2_X1 U659 ( .A1(n581), .A2(n578), .ZN(n683) );
  NAND2_X1 U660 ( .A1(n581), .A2(n578), .ZN(n680) );
  XNOR2_X1 U661 ( .A(n628), .B(n684), .ZN(n578) );
  NOR2_X1 U662 ( .A1(n547), .A2(n574), .ZN(n684) );
  INV_X1 U663 ( .A(n552), .ZN(n581) );
  NAND2_X1 U664 ( .A1(n685), .A2(n543), .ZN(n552) );
  INV_X1 U665 ( .A(n557), .ZN(n543) );
  NAND2_X1 U666 ( .A1(b_7_), .A2(a_7_), .ZN(n557) );
  INV_X1 U667 ( .A(n628), .ZN(n685) );
  NAND2_X1 U668 ( .A1(b_6_), .A2(a_6_), .ZN(n628) );
  XNOR2_X1 U669 ( .A(n686), .B(n687), .ZN(n608) );
  XNOR2_X1 U670 ( .A(n688), .B(n689), .ZN(n687) );
  XNOR2_X1 U671 ( .A(n690), .B(n691), .ZN(n615) );
  XOR2_X1 U672 ( .A(n692), .B(n693), .Z(n690) );
  NOR2_X1 U673 ( .A1(n555), .A2(n604), .ZN(n693) );
  XNOR2_X1 U674 ( .A(n694), .B(n695), .ZN(n477) );
  XOR2_X1 U675 ( .A(n696), .B(n697), .Z(n694) );
  NOR2_X1 U676 ( .A1(n555), .A2(n698), .ZN(n697) );
  XOR2_X1 U677 ( .A(n699), .B(n700), .Z(n495) );
  XOR2_X1 U678 ( .A(n701), .B(n702), .Z(n700) );
  NOR2_X1 U679 ( .A1(n703), .A2(n517), .ZN(n650) );
  AND2_X1 U680 ( .A1(n519), .A2(n520), .ZN(n517) );
  AND2_X1 U681 ( .A1(n704), .A2(n705), .ZN(n520) );
  NAND2_X1 U682 ( .A1(n706), .A2(n707), .ZN(n704) );
  INV_X1 U683 ( .A(n708), .ZN(n707) );
  XOR2_X1 U684 ( .A(n709), .B(n710), .Z(n706) );
  NOR2_X1 U685 ( .A1(n653), .A2(n654), .ZN(n519) );
  XOR2_X1 U686 ( .A(n711), .B(n712), .Z(n654) );
  NAND2_X1 U687 ( .A1(n713), .A2(n714), .ZN(n711) );
  AND2_X1 U688 ( .A1(n715), .A2(n716), .ZN(n653) );
  NAND2_X1 U689 ( .A1(n658), .A2(n717), .ZN(n716) );
  OR2_X1 U690 ( .A1(n656), .A2(n657), .ZN(n717) );
  NOR2_X1 U691 ( .A1(n718), .A2(n555), .ZN(n658) );
  NAND2_X1 U692 ( .A1(n656), .A2(n657), .ZN(n715) );
  NAND2_X1 U693 ( .A1(n719), .A2(n720), .ZN(n657) );
  NAND2_X1 U694 ( .A1(n702), .A2(n721), .ZN(n720) );
  NAND2_X1 U695 ( .A1(n701), .A2(n699), .ZN(n721) );
  NOR2_X1 U696 ( .A1(n555), .A2(n722), .ZN(n702) );
  OR2_X1 U697 ( .A1(n699), .A2(n701), .ZN(n719) );
  AND2_X1 U698 ( .A1(n723), .A2(n724), .ZN(n701) );
  NAND2_X1 U699 ( .A1(n725), .A2(a_2_), .ZN(n724) );
  NOR2_X1 U700 ( .A1(n726), .A2(n555), .ZN(n725) );
  NOR2_X1 U701 ( .A1(n696), .A2(n695), .ZN(n726) );
  NAND2_X1 U702 ( .A1(n695), .A2(n696), .ZN(n723) );
  NAND2_X1 U703 ( .A1(n727), .A2(n728), .ZN(n696) );
  NAND2_X1 U704 ( .A1(n729), .A2(a_3_), .ZN(n728) );
  NOR2_X1 U705 ( .A1(n730), .A2(n555), .ZN(n729) );
  NOR2_X1 U706 ( .A1(n691), .A2(n692), .ZN(n730) );
  NAND2_X1 U707 ( .A1(n691), .A2(n692), .ZN(n727) );
  NAND2_X1 U708 ( .A1(n731), .A2(n732), .ZN(n692) );
  NAND2_X1 U709 ( .A1(n689), .A2(n733), .ZN(n732) );
  OR2_X1 U710 ( .A1(n688), .A2(n686), .ZN(n733) );
  NOR2_X1 U711 ( .A1(n632), .A2(n555), .ZN(n689) );
  NAND2_X1 U712 ( .A1(n686), .A2(n688), .ZN(n731) );
  NAND2_X1 U713 ( .A1(n678), .A2(n734), .ZN(n688) );
  NAND2_X1 U714 ( .A1(n677), .A2(n679), .ZN(n734) );
  NAND2_X1 U715 ( .A1(n735), .A2(n736), .ZN(n679) );
  INV_X1 U716 ( .A(n737), .ZN(n736) );
  NAND2_X1 U717 ( .A1(a_5_), .A2(b_6_), .ZN(n735) );
  XNOR2_X1 U718 ( .A(n738), .B(n739), .ZN(n677) );
  NOR2_X1 U719 ( .A1(n547), .A2(n631), .ZN(n739) );
  NAND2_X1 U720 ( .A1(n737), .A2(a_5_), .ZN(n678) );
  NOR2_X1 U721 ( .A1(n561), .A2(n738), .ZN(n737) );
  NAND2_X1 U722 ( .A1(b_6_), .A2(a_7_), .ZN(n561) );
  XNOR2_X1 U723 ( .A(n740), .B(n741), .ZN(n686) );
  XOR2_X1 U724 ( .A(n625), .B(n742), .Z(n740) );
  XNOR2_X1 U725 ( .A(n743), .B(n744), .ZN(n691) );
  NAND2_X1 U726 ( .A1(n745), .A2(n746), .ZN(n743) );
  XOR2_X1 U727 ( .A(n747), .B(n748), .Z(n695) );
  XOR2_X1 U728 ( .A(n749), .B(n750), .Z(n747) );
  NOR2_X1 U729 ( .A1(n574), .A2(n604), .ZN(n750) );
  XOR2_X1 U730 ( .A(n751), .B(n752), .Z(n699) );
  XOR2_X1 U731 ( .A(n753), .B(n754), .Z(n752) );
  NAND2_X1 U732 ( .A1(a_2_), .A2(b_5_), .ZN(n754) );
  XOR2_X1 U733 ( .A(n755), .B(n756), .Z(n656) );
  XOR2_X1 U734 ( .A(n757), .B(n758), .Z(n756) );
  INV_X1 U735 ( .A(n705), .ZN(n703) );
  NAND2_X1 U736 ( .A1(n759), .A2(n708), .ZN(n705) );
  NAND2_X1 U737 ( .A1(n713), .A2(n760), .ZN(n708) );
  NAND2_X1 U738 ( .A1(n712), .A2(n714), .ZN(n760) );
  NAND2_X1 U739 ( .A1(n761), .A2(n762), .ZN(n714) );
  NAND2_X1 U740 ( .A1(a_0_), .A2(b_5_), .ZN(n762) );
  INV_X1 U741 ( .A(n763), .ZN(n761) );
  XNOR2_X1 U742 ( .A(n764), .B(n765), .ZN(n712) );
  NAND2_X1 U743 ( .A1(n766), .A2(n767), .ZN(n764) );
  NAND2_X1 U744 ( .A1(a_0_), .A2(n763), .ZN(n713) );
  NAND2_X1 U745 ( .A1(n768), .A2(n769), .ZN(n763) );
  NAND2_X1 U746 ( .A1(n758), .A2(n770), .ZN(n769) );
  NAND2_X1 U747 ( .A1(n757), .A2(n755), .ZN(n770) );
  NOR2_X1 U748 ( .A1(n574), .A2(n722), .ZN(n758) );
  OR2_X1 U749 ( .A1(n755), .A2(n757), .ZN(n768) );
  AND2_X1 U750 ( .A1(n771), .A2(n772), .ZN(n757) );
  NAND2_X1 U751 ( .A1(n773), .A2(a_2_), .ZN(n772) );
  NOR2_X1 U752 ( .A1(n774), .A2(n574), .ZN(n773) );
  NOR2_X1 U753 ( .A1(n753), .A2(n751), .ZN(n774) );
  NAND2_X1 U754 ( .A1(n751), .A2(n753), .ZN(n771) );
  NAND2_X1 U755 ( .A1(n775), .A2(n776), .ZN(n753) );
  NAND2_X1 U756 ( .A1(n777), .A2(a_3_), .ZN(n776) );
  NOR2_X1 U757 ( .A1(n778), .A2(n574), .ZN(n777) );
  INV_X1 U758 ( .A(b_5_), .ZN(n574) );
  NOR2_X1 U759 ( .A1(n748), .A2(n749), .ZN(n778) );
  NAND2_X1 U760 ( .A1(n748), .A2(n749), .ZN(n775) );
  NAND2_X1 U761 ( .A1(n745), .A2(n779), .ZN(n749) );
  NAND2_X1 U762 ( .A1(n744), .A2(n746), .ZN(n779) );
  NAND2_X1 U763 ( .A1(n780), .A2(n781), .ZN(n746) );
  NAND2_X1 U764 ( .A1(a_4_), .A2(b_5_), .ZN(n781) );
  INV_X1 U765 ( .A(n782), .ZN(n780) );
  XNOR2_X1 U766 ( .A(n783), .B(n784), .ZN(n744) );
  NAND2_X1 U767 ( .A1(n785), .A2(n786), .ZN(n783) );
  NAND2_X1 U768 ( .A1(a_4_), .A2(n782), .ZN(n745) );
  NAND2_X1 U769 ( .A1(n787), .A2(n788), .ZN(n782) );
  NAND2_X1 U770 ( .A1(n742), .A2(n789), .ZN(n788) );
  OR2_X1 U771 ( .A1(n741), .A2(n568), .ZN(n789) );
  NOR2_X1 U772 ( .A1(n790), .A2(n738), .ZN(n742) );
  NAND2_X1 U773 ( .A1(b_5_), .A2(a_6_), .ZN(n738) );
  NAND2_X1 U774 ( .A1(a_7_), .A2(b_4_), .ZN(n790) );
  NAND2_X1 U775 ( .A1(n568), .A2(n741), .ZN(n787) );
  XOR2_X1 U776 ( .A(n791), .B(n792), .Z(n741) );
  INV_X1 U777 ( .A(n625), .ZN(n568) );
  NAND2_X1 U778 ( .A1(a_5_), .A2(b_5_), .ZN(n625) );
  XOR2_X1 U779 ( .A(n793), .B(n794), .Z(n748) );
  XOR2_X1 U780 ( .A(n592), .B(n795), .Z(n794) );
  XNOR2_X1 U781 ( .A(n796), .B(n797), .ZN(n751) );
  XOR2_X1 U782 ( .A(n798), .B(n799), .Z(n797) );
  XNOR2_X1 U783 ( .A(n800), .B(n801), .ZN(n755) );
  NOR2_X1 U784 ( .A1(n802), .A2(n803), .ZN(n801) );
  NOR2_X1 U785 ( .A1(n804), .A2(n805), .ZN(n802) );
  NOR2_X1 U786 ( .A1(n631), .A2(n698), .ZN(n805) );
  INV_X1 U787 ( .A(n806), .ZN(n804) );
  XNOR2_X1 U788 ( .A(n709), .B(n710), .ZN(n759) );
  XNOR2_X1 U789 ( .A(n807), .B(n808), .ZN(n709) );
  NOR2_X1 U790 ( .A1(n631), .A2(n718), .ZN(n808) );
  XOR2_X1 U791 ( .A(n647), .B(n646), .Z(n522) );
  NAND2_X1 U792 ( .A1(n809), .A2(n810), .ZN(n528) );
  XOR2_X1 U793 ( .A(n811), .B(n648), .Z(n810) );
  AND2_X1 U794 ( .A1(n647), .A2(n646), .ZN(n809) );
  XOR2_X1 U795 ( .A(n812), .B(n813), .Z(n646) );
  XNOR2_X1 U796 ( .A(n814), .B(n815), .ZN(n813) );
  NAND2_X1 U797 ( .A1(a_0_), .A2(b_3_), .ZN(n815) );
  NAND2_X1 U798 ( .A1(n816), .A2(n817), .ZN(n647) );
  NAND2_X1 U799 ( .A1(n818), .A2(a_0_), .ZN(n817) );
  NOR2_X1 U800 ( .A1(n819), .A2(n631), .ZN(n818) );
  NOR2_X1 U801 ( .A1(n710), .A2(n807), .ZN(n819) );
  NAND2_X1 U802 ( .A1(n710), .A2(n807), .ZN(n816) );
  NAND2_X1 U803 ( .A1(n766), .A2(n820), .ZN(n807) );
  NAND2_X1 U804 ( .A1(n765), .A2(n767), .ZN(n820) );
  NAND2_X1 U805 ( .A1(n821), .A2(n822), .ZN(n767) );
  NAND2_X1 U806 ( .A1(b_4_), .A2(a_1_), .ZN(n822) );
  XNOR2_X1 U807 ( .A(n823), .B(n824), .ZN(n765) );
  XOR2_X1 U808 ( .A(n825), .B(n826), .Z(n823) );
  NAND2_X1 U809 ( .A1(a_2_), .A2(b_3_), .ZN(n825) );
  OR2_X1 U810 ( .A1(n722), .A2(n821), .ZN(n766) );
  NOR2_X1 U811 ( .A1(n803), .A2(n827), .ZN(n821) );
  AND2_X1 U812 ( .A1(n800), .A2(n828), .ZN(n827) );
  NAND2_X1 U813 ( .A1(n806), .A2(n829), .ZN(n828) );
  NAND2_X1 U814 ( .A1(a_2_), .A2(b_4_), .ZN(n829) );
  XOR2_X1 U815 ( .A(n830), .B(n831), .Z(n800) );
  XOR2_X1 U816 ( .A(n621), .B(n832), .Z(n830) );
  NOR2_X1 U817 ( .A1(n806), .A2(n698), .ZN(n803) );
  NAND2_X1 U818 ( .A1(n833), .A2(n834), .ZN(n806) );
  NAND2_X1 U819 ( .A1(n796), .A2(n835), .ZN(n834) );
  OR2_X1 U820 ( .A1(n799), .A2(n798), .ZN(n835) );
  XOR2_X1 U821 ( .A(n836), .B(n837), .Z(n796) );
  NAND2_X1 U822 ( .A1(n838), .A2(n839), .ZN(n836) );
  NAND2_X1 U823 ( .A1(n799), .A2(n798), .ZN(n833) );
  NAND2_X1 U824 ( .A1(n840), .A2(n841), .ZN(n798) );
  NAND2_X1 U825 ( .A1(n793), .A2(n842), .ZN(n841) );
  NAND2_X1 U826 ( .A1(n843), .A2(n795), .ZN(n842) );
  XOR2_X1 U827 ( .A(n844), .B(n845), .Z(n793) );
  NAND2_X1 U828 ( .A1(n846), .A2(n847), .ZN(n844) );
  OR2_X1 U829 ( .A1(n795), .A2(n843), .ZN(n840) );
  INV_X1 U830 ( .A(n592), .ZN(n843) );
  NAND2_X1 U831 ( .A1(b_4_), .A2(a_4_), .ZN(n592) );
  NAND2_X1 U832 ( .A1(n785), .A2(n848), .ZN(n795) );
  NAND2_X1 U833 ( .A1(n784), .A2(n786), .ZN(n848) );
  NAND2_X1 U834 ( .A1(n849), .A2(n850), .ZN(n786) );
  NAND2_X1 U835 ( .A1(b_4_), .A2(a_5_), .ZN(n850) );
  AND2_X1 U836 ( .A1(n851), .A2(n852), .ZN(n784) );
  NAND2_X1 U837 ( .A1(n853), .A2(n854), .ZN(n852) );
  NAND2_X1 U838 ( .A1(b_3_), .A2(a_6_), .ZN(n853) );
  OR2_X1 U839 ( .A1(n849), .A2(n576), .ZN(n785) );
  NAND2_X1 U840 ( .A1(n791), .A2(n792), .ZN(n849) );
  NOR2_X1 U841 ( .A1(n631), .A2(n558), .ZN(n792) );
  NOR2_X1 U842 ( .A1(n605), .A2(n547), .ZN(n791) );
  NAND2_X1 U843 ( .A1(a_3_), .A2(b_4_), .ZN(n799) );
  XNOR2_X1 U844 ( .A(n855), .B(n856), .ZN(n710) );
  XOR2_X1 U845 ( .A(n857), .B(n858), .Z(n856) );
  NAND2_X1 U846 ( .A1(n859), .A2(n860), .ZN(n533) );
  OR2_X1 U847 ( .A1(n648), .A2(n811), .ZN(n860) );
  INV_X1 U848 ( .A(n649), .ZN(n811) );
  XNOR2_X1 U849 ( .A(n861), .B(n862), .ZN(n859) );
  NAND2_X1 U850 ( .A1(n863), .A2(n864), .ZN(n532) );
  AND2_X1 U851 ( .A1(n637), .A2(n649), .ZN(n864) );
  NAND2_X1 U852 ( .A1(n865), .A2(n866), .ZN(n649) );
  NAND2_X1 U853 ( .A1(n867), .A2(a_0_), .ZN(n866) );
  NOR2_X1 U854 ( .A1(n868), .A2(n605), .ZN(n867) );
  NOR2_X1 U855 ( .A1(n814), .A2(n812), .ZN(n868) );
  NAND2_X1 U856 ( .A1(n814), .A2(n812), .ZN(n865) );
  XOR2_X1 U857 ( .A(n869), .B(n870), .Z(n812) );
  XOR2_X1 U858 ( .A(n871), .B(n872), .Z(n869) );
  AND2_X1 U859 ( .A1(n873), .A2(n874), .ZN(n814) );
  NAND2_X1 U860 ( .A1(n857), .A2(n875), .ZN(n874) );
  NAND2_X1 U861 ( .A1(n858), .A2(n855), .ZN(n875) );
  AND2_X1 U862 ( .A1(n876), .A2(n877), .ZN(n857) );
  NAND2_X1 U863 ( .A1(n878), .A2(a_2_), .ZN(n877) );
  NOR2_X1 U864 ( .A1(n879), .A2(n605), .ZN(n878) );
  NOR2_X1 U865 ( .A1(n826), .A2(n824), .ZN(n879) );
  NAND2_X1 U866 ( .A1(n826), .A2(n824), .ZN(n876) );
  XOR2_X1 U867 ( .A(n880), .B(n881), .Z(n824) );
  XNOR2_X1 U868 ( .A(n882), .B(n883), .ZN(n880) );
  NAND2_X1 U869 ( .A1(b_2_), .A2(a_3_), .ZN(n882) );
  AND2_X1 U870 ( .A1(n884), .A2(n885), .ZN(n826) );
  NAND2_X1 U871 ( .A1(n832), .A2(n886), .ZN(n885) );
  NAND2_X1 U872 ( .A1(n599), .A2(n831), .ZN(n886) );
  INV_X1 U873 ( .A(n887), .ZN(n831) );
  INV_X1 U874 ( .A(n621), .ZN(n599) );
  AND2_X1 U875 ( .A1(n838), .A2(n888), .ZN(n832) );
  NAND2_X1 U876 ( .A1(n837), .A2(n839), .ZN(n888) );
  NAND2_X1 U877 ( .A1(n889), .A2(n890), .ZN(n839) );
  NAND2_X1 U878 ( .A1(b_3_), .A2(a_4_), .ZN(n890) );
  INV_X1 U879 ( .A(n891), .ZN(n889) );
  XNOR2_X1 U880 ( .A(n892), .B(n893), .ZN(n837) );
  NAND2_X1 U881 ( .A1(n894), .A2(n895), .ZN(n892) );
  NAND2_X1 U882 ( .A1(a_4_), .A2(n891), .ZN(n838) );
  NAND2_X1 U883 ( .A1(n846), .A2(n896), .ZN(n891) );
  NAND2_X1 U884 ( .A1(n845), .A2(n847), .ZN(n896) );
  NAND2_X1 U885 ( .A1(n851), .A2(n897), .ZN(n847) );
  NAND2_X1 U886 ( .A1(b_3_), .A2(a_5_), .ZN(n897) );
  XOR2_X1 U887 ( .A(n898), .B(n899), .Z(n845) );
  OR2_X1 U888 ( .A1(n851), .A2(n576), .ZN(n846) );
  NAND2_X1 U889 ( .A1(n900), .A2(n901), .ZN(n851) );
  INV_X1 U890 ( .A(n854), .ZN(n901) );
  NAND2_X1 U891 ( .A1(b_2_), .A2(a_7_), .ZN(n854) );
  NOR2_X1 U892 ( .A1(n558), .A2(n605), .ZN(n900) );
  NAND2_X1 U893 ( .A1(n887), .A2(n621), .ZN(n884) );
  NAND2_X1 U894 ( .A1(a_3_), .A2(b_3_), .ZN(n621) );
  XOR2_X1 U895 ( .A(n902), .B(n903), .Z(n887) );
  NAND2_X1 U896 ( .A1(n904), .A2(n905), .ZN(n902) );
  OR2_X1 U897 ( .A1(n855), .A2(n858), .ZN(n873) );
  NOR2_X1 U898 ( .A1(n605), .A2(n722), .ZN(n858) );
  XOR2_X1 U899 ( .A(n906), .B(n907), .Z(n855) );
  XOR2_X1 U900 ( .A(n908), .B(n502), .Z(n906) );
  NAND2_X1 U901 ( .A1(n862), .A2(n861), .ZN(n637) );
  NOR2_X1 U902 ( .A1(n909), .A2(n648), .ZN(n863) );
  XNOR2_X1 U903 ( .A(n910), .B(n911), .ZN(n648) );
  XNOR2_X1 U904 ( .A(n912), .B(n913), .ZN(n910) );
  NOR2_X1 U905 ( .A1(n914), .A2(n718), .ZN(n913) );
  NOR2_X1 U906 ( .A1(n861), .A2(n862), .ZN(n909) );
  NAND2_X1 U907 ( .A1(n915), .A2(n916), .ZN(n862) );
  XNOR2_X1 U908 ( .A(n640), .B(n641), .ZN(n916) );
  NOR2_X1 U909 ( .A1(n718), .A2(n917), .ZN(n641) );
  NOR2_X1 U910 ( .A1(n722), .A2(n638), .ZN(n640) );
  NOR2_X1 U911 ( .A1(n918), .A2(n919), .ZN(n915) );
  NOR2_X1 U912 ( .A1(n506), .A2(n920), .ZN(n918) );
  NAND2_X1 U913 ( .A1(a_2_), .A2(b_0_), .ZN(n920) );
  NAND2_X1 U914 ( .A1(n912), .A2(n921), .ZN(n861) );
  NAND2_X1 U915 ( .A1(n911), .A2(b_2_), .ZN(n921) );
  XNOR2_X1 U916 ( .A(n922), .B(n923), .ZN(n911) );
  NOR2_X1 U917 ( .A1(n638), .A2(n698), .ZN(n923) );
  OR2_X1 U918 ( .A1(n506), .A2(n919), .ZN(n922) );
  NAND2_X1 U919 ( .A1(n924), .A2(n925), .ZN(n919) );
  NAND2_X1 U920 ( .A1(n926), .A2(n927), .ZN(n925) );
  NAND2_X1 U921 ( .A1(n928), .A2(n698), .ZN(n926) );
  NAND2_X1 U922 ( .A1(b_1_), .A2(a_1_), .ZN(n506) );
  AND2_X1 U923 ( .A1(n929), .A2(n930), .ZN(n912) );
  NAND2_X1 U924 ( .A1(n872), .A2(n931), .ZN(n930) );
  OR2_X1 U925 ( .A1(n871), .A2(n870), .ZN(n931) );
  NOR2_X1 U926 ( .A1(n914), .A2(n722), .ZN(n872) );
  INV_X1 U927 ( .A(a_1_), .ZN(n722) );
  NAND2_X1 U928 ( .A1(n870), .A2(n871), .ZN(n929) );
  NAND2_X1 U929 ( .A1(n932), .A2(n933), .ZN(n871) );
  NAND2_X1 U930 ( .A1(n502), .A2(n934), .ZN(n933) );
  OR2_X1 U931 ( .A1(n908), .A2(n907), .ZN(n934) );
  NOR2_X1 U932 ( .A1(n914), .A2(n698), .ZN(n502) );
  NAND2_X1 U933 ( .A1(n907), .A2(n908), .ZN(n932) );
  NAND2_X1 U934 ( .A1(n935), .A2(n936), .ZN(n908) );
  NAND2_X1 U935 ( .A1(n937), .A2(b_2_), .ZN(n936) );
  NOR2_X1 U936 ( .A1(n938), .A2(n604), .ZN(n937) );
  NOR2_X1 U937 ( .A1(n881), .A2(n883), .ZN(n938) );
  NAND2_X1 U938 ( .A1(n881), .A2(n883), .ZN(n935) );
  NAND2_X1 U939 ( .A1(n904), .A2(n939), .ZN(n883) );
  NAND2_X1 U940 ( .A1(n903), .A2(n905), .ZN(n939) );
  NAND2_X1 U941 ( .A1(n940), .A2(n941), .ZN(n905) );
  NAND2_X1 U942 ( .A1(b_2_), .A2(a_4_), .ZN(n941) );
  INV_X1 U943 ( .A(n942), .ZN(n940) );
  XNOR2_X1 U944 ( .A(n943), .B(n944), .ZN(n903) );
  XOR2_X1 U945 ( .A(n945), .B(n946), .Z(n944) );
  NAND2_X1 U946 ( .A1(a_4_), .A2(n942), .ZN(n904) );
  NAND2_X1 U947 ( .A1(n894), .A2(n947), .ZN(n942) );
  NAND2_X1 U948 ( .A1(n893), .A2(n895), .ZN(n947) );
  NAND2_X1 U949 ( .A1(n948), .A2(n949), .ZN(n895) );
  NAND2_X1 U950 ( .A1(b_2_), .A2(a_5_), .ZN(n949) );
  AND2_X1 U951 ( .A1(n943), .A2(n950), .ZN(n893) );
  NAND2_X1 U952 ( .A1(n951), .A2(n952), .ZN(n950) );
  NAND2_X1 U953 ( .A1(a_7_), .A2(b_0_), .ZN(n952) );
  NAND2_X1 U954 ( .A1(b_1_), .A2(a_6_), .ZN(n951) );
  OR2_X1 U955 ( .A1(n948), .A2(n576), .ZN(n894) );
  NAND2_X1 U956 ( .A1(n898), .A2(n899), .ZN(n948) );
  NOR2_X1 U957 ( .A1(n914), .A2(n558), .ZN(n898) );
  XOR2_X1 U958 ( .A(n953), .B(n954), .Z(n881) );
  NOR2_X1 U959 ( .A1(n638), .A2(n576), .ZN(n954) );
  XOR2_X1 U960 ( .A(n955), .B(n956), .Z(n953) );
  XOR2_X1 U961 ( .A(n957), .B(n958), .Z(n907) );
  XNOR2_X1 U962 ( .A(n959), .B(n960), .ZN(n958) );
  NAND2_X1 U963 ( .A1(a_4_), .A2(b_0_), .ZN(n957) );
  XNOR2_X1 U964 ( .A(n961), .B(n927), .ZN(n870) );
  NAND2_X1 U965 ( .A1(n962), .A2(n963), .ZN(n927) );
  NAND2_X1 U966 ( .A1(n964), .A2(a_4_), .ZN(n963) );
  NOR2_X1 U967 ( .A1(n965), .A2(n638), .ZN(n964) );
  NOR2_X1 U968 ( .A1(n959), .A2(n960), .ZN(n965) );
  NAND2_X1 U969 ( .A1(n959), .A2(n960), .ZN(n962) );
  NAND2_X1 U970 ( .A1(n966), .A2(n967), .ZN(n960) );
  NAND2_X1 U971 ( .A1(n968), .A2(a_5_), .ZN(n967) );
  NOR2_X1 U972 ( .A1(n969), .A2(n638), .ZN(n968) );
  NOR2_X1 U973 ( .A1(n955), .A2(n956), .ZN(n969) );
  NAND2_X1 U974 ( .A1(n955), .A2(n956), .ZN(n966) );
  NAND2_X1 U975 ( .A1(n943), .A2(n970), .ZN(n956) );
  NAND2_X1 U976 ( .A1(n945), .A2(n946), .ZN(n970) );
  NOR2_X1 U977 ( .A1(n917), .A2(n576), .ZN(n945) );
  NAND2_X1 U978 ( .A1(n946), .A2(n899), .ZN(n943) );
  NOR2_X1 U979 ( .A1(n917), .A2(n547), .ZN(n899) );
  NOR2_X1 U980 ( .A1(n558), .A2(n638), .ZN(n946) );
  NOR2_X1 U981 ( .A1(n917), .A2(n632), .ZN(n955) );
  NOR2_X1 U982 ( .A1(n917), .A2(n604), .ZN(n959) );
  NAND2_X1 U983 ( .A1(n924), .A2(n971), .ZN(n961) );
  NAND2_X1 U984 ( .A1(n972), .A2(n928), .ZN(n971) );
  NAND2_X1 U985 ( .A1(b_1_), .A2(a_2_), .ZN(n972) );
  NAND2_X1 U986 ( .A1(n973), .A2(n974), .ZN(n924) );
  INV_X1 U987 ( .A(n928), .ZN(n974) );
  NAND2_X1 U988 ( .A1(a_3_), .A2(b_0_), .ZN(n928) );
  NOR2_X1 U989 ( .A1(n698), .A2(n917), .ZN(n973) );
  INV_X1 U990 ( .A(n476), .ZN(n481) );
  NAND2_X1 U991 ( .A1(n975), .A2(n976), .ZN(n476) );
  NAND2_X1 U992 ( .A1(n977), .A2(n500), .ZN(n976) );
  NAND2_X1 U993 ( .A1(b_0_), .A2(n718), .ZN(n500) );
  INV_X1 U994 ( .A(a_0_), .ZN(n718) );
  NAND2_X1 U995 ( .A1(n978), .A2(n979), .ZN(n977) );
  NAND2_X1 U996 ( .A1(a_1_), .A2(n917), .ZN(n979) );
  NAND2_X1 U997 ( .A1(n980), .A2(n981), .ZN(n978) );
  NAND2_X1 U998 ( .A1(b_2_), .A2(n698), .ZN(n981) );
  INV_X1 U999 ( .A(a_2_), .ZN(n698) );
  NOR2_X1 U1000 ( .A1(n982), .A2(n983), .ZN(n980) );
  NOR2_X1 U1001 ( .A1(a_1_), .A2(n917), .ZN(n983) );
  INV_X1 U1002 ( .A(b_1_), .ZN(n917) );
  NOR2_X1 U1003 ( .A1(n984), .A2(n985), .ZN(n982) );
  NAND2_X1 U1004 ( .A1(n986), .A2(n987), .ZN(n985) );
  NAND2_X1 U1005 ( .A1(n988), .A2(n989), .ZN(n987) );
  NAND2_X1 U1006 ( .A1(b_4_), .A2(n632), .ZN(n989) );
  INV_X1 U1007 ( .A(a_4_), .ZN(n632) );
  NOR2_X1 U1008 ( .A1(n990), .A2(n991), .ZN(n988) );
  NOR2_X1 U1009 ( .A1(a_3_), .A2(n605), .ZN(n991) );
  INV_X1 U1010 ( .A(b_3_), .ZN(n605) );
  NOR2_X1 U1011 ( .A1(n992), .A2(n993), .ZN(n990) );
  NAND2_X1 U1012 ( .A1(n994), .A2(n995), .ZN(n993) );
  NAND2_X1 U1013 ( .A1(n996), .A2(n997), .ZN(n995) );
  NAND2_X1 U1014 ( .A1(b_5_), .A2(n576), .ZN(n997) );
  NOR2_X1 U1015 ( .A1(n998), .A2(n999), .ZN(n996) );
  NOR2_X1 U1016 ( .A1(a_6_), .A2(n1000), .ZN(n999) );
  NOR2_X1 U1017 ( .A1(n1001), .A2(n555), .ZN(n998) );
  INV_X1 U1018 ( .A(b_6_), .ZN(n555) );
  NOR2_X1 U1019 ( .A1(n545), .A2(n558), .ZN(n1001) );
  INV_X1 U1020 ( .A(a_6_), .ZN(n558) );
  INV_X1 U1021 ( .A(n1000), .ZN(n545) );
  NOR2_X1 U1022 ( .A1(n547), .A2(b_7_), .ZN(n1000) );
  INV_X1 U1023 ( .A(a_7_), .ZN(n547) );
  NAND2_X1 U1024 ( .A1(a_4_), .A2(n631), .ZN(n994) );
  INV_X1 U1025 ( .A(b_4_), .ZN(n631) );
  NOR2_X1 U1026 ( .A1(b_5_), .A2(n576), .ZN(n992) );
  INV_X1 U1027 ( .A(a_5_), .ZN(n576) );
  NAND2_X1 U1028 ( .A1(a_2_), .A2(n914), .ZN(n986) );
  INV_X1 U1029 ( .A(b_2_), .ZN(n914) );
  NOR2_X1 U1030 ( .A1(b_3_), .A2(n604), .ZN(n984) );
  INV_X1 U1031 ( .A(a_3_), .ZN(n604) );
  NAND2_X1 U1032 ( .A1(a_0_), .A2(n638), .ZN(n975) );
  INV_X1 U1033 ( .A(b_0_), .ZN(n638) );
endmodule

