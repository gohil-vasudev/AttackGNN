module locked_c1355 (  G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,  G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT  );
  input  G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n343_, new_n345_, new_n346_, new_n348_, new_n349_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n371_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n382_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n395_, new_n397_, new_n399_, new_n400_, new_n402_, new_n403_, new_n405_, new_n407_, new_n409_, new_n410_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n437_, new_n438_, new_n440_, new_n441_, new_n443_, new_n444_, new_n446_, new_n447_, new_n448_, new_n450_, new_n451_, new_n452_, new_n454_, new_n456_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n481_, new_n483_, new_n484_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n498_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_;
  XNOR2_X1 g000 ( .A(G155GAT), .B(KEYINPUT3), .ZN(new_n138_) );
  XNOR2_X1 g001 ( .A(G141GAT), .B(KEYINPUT2), .ZN(new_n139_) );
  XNOR2_X1 g002 ( .A(new_n138_), .B(new_n139_), .ZN(new_n140_) );
  XNOR2_X1 g003 ( .A(G57GAT), .B(KEYINPUT1), .ZN(new_n141_) );
  NAND2_X1 g004 ( .A1(G225GAT), .A2(G233GAT), .ZN(new_n142_) );
  XNOR2_X1 g005 ( .A(new_n141_), .B(new_n142_), .ZN(new_n143_) );
  XNOR2_X1 g006 ( .A(new_n140_), .B(new_n143_), .ZN(new_n144_) );
  INV_X1 g007 ( .A(G1GAT), .ZN(new_n145_) );
  XNOR2_X1 g008 ( .A(G120GAT), .B(G127GAT), .ZN(new_n146_) );
  XNOR2_X1 g009 ( .A(G113GAT), .B(KEYINPUT0), .ZN(new_n147_) );
  XNOR2_X1 g010 ( .A(new_n146_), .B(new_n147_), .ZN(new_n148_) );
  XNOR2_X1 g011 ( .A(new_n148_), .B(new_n145_), .ZN(new_n149_) );
  XNOR2_X1 g012 ( .A(new_n144_), .B(new_n149_), .ZN(new_n150_) );
  XNOR2_X1 g013 ( .A(G29GAT), .B(G134GAT), .ZN(new_n151_) );
  XNOR2_X1 g014 ( .A(new_n150_), .B(new_n151_), .ZN(new_n152_) );
  XNOR2_X1 g015 ( .A(G85GAT), .B(G162GAT), .ZN(new_n153_) );
  XNOR2_X1 g016 ( .A(new_n152_), .B(new_n153_), .ZN(new_n154_) );
  XOR2_X1 g017 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(new_n155_) );
  XNOR2_X1 g018 ( .A(G148GAT), .B(KEYINPUT6), .ZN(new_n156_) );
  XNOR2_X1 g019 ( .A(new_n155_), .B(new_n156_), .ZN(new_n157_) );
  XNOR2_X1 g020 ( .A(new_n154_), .B(new_n157_), .ZN(new_n158_) );
  INV_X1 g021 ( .A(new_n158_), .ZN(new_n159_) );
  INV_X1 g022 ( .A(KEYINPUT26), .ZN(new_n160_) );
  INV_X1 g023 ( .A(G197GAT), .ZN(new_n161_) );
  XNOR2_X1 g024 ( .A(G211GAT), .B(G218GAT), .ZN(new_n162_) );
  XNOR2_X1 g025 ( .A(G204GAT), .B(KEYINPUT21), .ZN(new_n163_) );
  XNOR2_X1 g026 ( .A(new_n162_), .B(new_n163_), .ZN(new_n164_) );
  XNOR2_X1 g027 ( .A(new_n164_), .B(new_n161_), .ZN(new_n165_) );
  XNOR2_X1 g028 ( .A(new_n165_), .B(new_n140_), .ZN(new_n166_) );
  XOR2_X1 g029 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(new_n167_) );
  XNOR2_X1 g030 ( .A(G22GAT), .B(KEYINPUT22), .ZN(new_n168_) );
  XNOR2_X1 g031 ( .A(new_n167_), .B(new_n168_), .ZN(new_n169_) );
  INV_X1 g032 ( .A(G148GAT), .ZN(new_n170_) );
  NAND2_X1 g033 ( .A1(G78GAT), .A2(G106GAT), .ZN(new_n171_) );
  OR2_X1 g034 ( .A1(G78GAT), .A2(G106GAT), .ZN(new_n172_) );
  NAND3_X1 g035 ( .A1(new_n172_), .A2(new_n170_), .A3(new_n171_), .ZN(new_n173_) );
  NAND2_X1 g036 ( .A1(new_n172_), .A2(new_n171_), .ZN(new_n174_) );
  NAND2_X1 g037 ( .A1(new_n174_), .A2(G148GAT), .ZN(new_n175_) );
  NAND2_X1 g038 ( .A1(new_n175_), .A2(new_n173_), .ZN(new_n176_) );
  XNOR2_X1 g039 ( .A(new_n169_), .B(new_n176_), .ZN(new_n177_) );
  NAND2_X1 g040 ( .A1(new_n166_), .A2(new_n177_), .ZN(new_n178_) );
  OR2_X1 g041 ( .A1(new_n166_), .A2(new_n177_), .ZN(new_n179_) );
  XOR2_X1 g042 ( .A(G50GAT), .B(G162GAT), .Z(new_n180_) );
  NAND3_X1 g043 ( .A1(new_n179_), .A2(new_n178_), .A3(new_n180_), .ZN(new_n181_) );
  NAND2_X1 g044 ( .A1(new_n179_), .A2(new_n178_), .ZN(new_n182_) );
  INV_X1 g045 ( .A(new_n180_), .ZN(new_n183_) );
  NAND2_X1 g046 ( .A1(new_n182_), .A2(new_n183_), .ZN(new_n184_) );
  NAND4_X1 g047 ( .A1(new_n184_), .A2(G228GAT), .A3(G233GAT), .A4(new_n181_), .ZN(new_n185_) );
  NAND2_X1 g048 ( .A1(new_n184_), .A2(new_n181_), .ZN(new_n186_) );
  NAND2_X1 g049 ( .A1(G228GAT), .A2(G233GAT), .ZN(new_n187_) );
  NAND2_X1 g050 ( .A1(new_n186_), .A2(new_n187_), .ZN(new_n188_) );
  NAND2_X1 g051 ( .A1(new_n188_), .A2(new_n185_), .ZN(new_n189_) );
  XOR2_X1 g052 ( .A(new_n148_), .B(G15GAT), .Z(new_n190_) );
  NAND2_X1 g053 ( .A1(G227GAT), .A2(G233GAT), .ZN(new_n191_) );
  XNOR2_X1 g054 ( .A(new_n190_), .B(new_n191_), .ZN(new_n192_) );
  XNOR2_X1 g055 ( .A(G176GAT), .B(G183GAT), .ZN(new_n193_) );
  XNOR2_X1 g056 ( .A(G71GAT), .B(KEYINPUT20), .ZN(new_n194_) );
  XNOR2_X1 g057 ( .A(new_n193_), .B(new_n194_), .ZN(new_n195_) );
  XNOR2_X1 g058 ( .A(new_n192_), .B(new_n195_), .ZN(new_n196_) );
  XNOR2_X1 g059 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(new_n197_) );
  XNOR2_X1 g060 ( .A(G169GAT), .B(KEYINPUT19), .ZN(new_n198_) );
  XNOR2_X1 g061 ( .A(new_n197_), .B(new_n198_), .ZN(new_n199_) );
  XOR2_X1 g062 ( .A(G134GAT), .B(G190GAT), .Z(new_n200_) );
  XNOR2_X1 g063 ( .A(G43GAT), .B(G99GAT), .ZN(new_n201_) );
  XNOR2_X1 g064 ( .A(new_n200_), .B(new_n201_), .ZN(new_n202_) );
  XOR2_X1 g065 ( .A(new_n202_), .B(new_n199_), .Z(new_n203_) );
  XNOR2_X1 g066 ( .A(new_n196_), .B(new_n203_), .ZN(new_n204_) );
  INV_X1 g067 ( .A(new_n204_), .ZN(new_n205_) );
  NAND2_X1 g068 ( .A1(new_n189_), .A2(new_n205_), .ZN(new_n206_) );
  NAND2_X1 g069 ( .A1(new_n206_), .A2(new_n160_), .ZN(new_n207_) );
  NAND3_X1 g070 ( .A1(new_n189_), .A2(KEYINPUT26), .A3(new_n205_), .ZN(new_n208_) );
  NAND2_X1 g071 ( .A1(new_n207_), .A2(new_n208_), .ZN(new_n209_) );
  XNOR2_X1 g072 ( .A(G36GAT), .B(G190GAT), .ZN(new_n210_) );
  INV_X1 g073 ( .A(new_n210_), .ZN(new_n211_) );
  XNOR2_X1 g074 ( .A(new_n165_), .B(new_n211_), .ZN(new_n212_) );
  XNOR2_X1 g075 ( .A(G64GAT), .B(G176GAT), .ZN(new_n213_) );
  XNOR2_X1 g076 ( .A(new_n213_), .B(G92GAT), .ZN(new_n214_) );
  NAND2_X1 g077 ( .A1(G226GAT), .A2(G233GAT), .ZN(new_n215_) );
  XNOR2_X1 g078 ( .A(new_n214_), .B(new_n215_), .ZN(new_n216_) );
  XNOR2_X1 g079 ( .A(G8GAT), .B(G183GAT), .ZN(new_n217_) );
  XNOR2_X1 g080 ( .A(new_n216_), .B(new_n217_), .ZN(new_n218_) );
  XNOR2_X1 g081 ( .A(new_n212_), .B(new_n218_), .ZN(new_n219_) );
  XNOR2_X1 g082 ( .A(new_n219_), .B(new_n199_), .ZN(new_n220_) );
  XNOR2_X1 g083 ( .A(new_n220_), .B(KEYINPUT27), .ZN(new_n221_) );
  NAND2_X1 g084 ( .A1(new_n209_), .A2(new_n221_), .ZN(new_n222_) );
  INV_X1 g085 ( .A(KEYINPUT25), .ZN(new_n223_) );
  NAND2_X1 g086 ( .A1(new_n204_), .A2(new_n220_), .ZN(new_n224_) );
  NAND3_X1 g087 ( .A1(new_n224_), .A2(new_n185_), .A3(new_n188_), .ZN(new_n225_) );
  XNOR2_X1 g088 ( .A(new_n225_), .B(new_n223_), .ZN(new_n226_) );
  NAND2_X1 g089 ( .A1(new_n222_), .A2(new_n226_), .ZN(new_n227_) );
  NAND2_X1 g090 ( .A1(new_n227_), .A2(new_n159_), .ZN(new_n228_) );
  INV_X1 g091 ( .A(KEYINPUT28), .ZN(new_n229_) );
  XNOR2_X1 g092 ( .A(new_n189_), .B(new_n229_), .ZN(new_n230_) );
  AND2_X1 g093 ( .A1(new_n158_), .A2(new_n221_), .ZN(new_n231_) );
  NAND3_X1 g094 ( .A1(new_n231_), .A2(new_n230_), .A3(new_n205_), .ZN(new_n232_) );
  NAND2_X1 g095 ( .A1(new_n228_), .A2(new_n232_), .ZN(new_n233_) );
  XNOR2_X1 g096 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(new_n234_) );
  XNOR2_X1 g097 ( .A(G64GAT), .B(KEYINPUT15), .ZN(new_n235_) );
  XNOR2_X1 g098 ( .A(new_n234_), .B(new_n235_), .ZN(new_n236_) );
  XNOR2_X1 g099 ( .A(G78GAT), .B(G155GAT), .ZN(new_n237_) );
  XNOR2_X1 g100 ( .A(G127GAT), .B(G211GAT), .ZN(new_n238_) );
  XNOR2_X1 g101 ( .A(new_n237_), .B(new_n238_), .ZN(new_n239_) );
  XNOR2_X1 g102 ( .A(new_n236_), .B(new_n239_), .ZN(new_n240_) );
  XNOR2_X1 g103 ( .A(G57GAT), .B(G71GAT), .ZN(new_n241_) );
  XOR2_X1 g104 ( .A(new_n241_), .B(KEYINPUT13), .Z(new_n242_) );
  XNOR2_X1 g105 ( .A(G15GAT), .B(G22GAT), .ZN(new_n243_) );
  XNOR2_X1 g106 ( .A(new_n243_), .B(new_n145_), .ZN(new_n244_) );
  XNOR2_X1 g107 ( .A(new_n242_), .B(new_n244_), .ZN(new_n245_) );
  XNOR2_X1 g108 ( .A(new_n245_), .B(new_n240_), .ZN(new_n246_) );
  XNOR2_X1 g109 ( .A(new_n246_), .B(new_n217_), .ZN(new_n247_) );
  AND2_X1 g110 ( .A1(G231GAT), .A2(G233GAT), .ZN(new_n248_) );
  XNOR2_X1 g111 ( .A(new_n247_), .B(new_n248_), .ZN(new_n249_) );
  OR2_X1 g112 ( .A1(G43GAT), .A2(KEYINPUT8), .ZN(new_n250_) );
  NAND2_X1 g113 ( .A1(G43GAT), .A2(KEYINPUT8), .ZN(new_n251_) );
  NAND2_X1 g114 ( .A1(new_n250_), .A2(new_n251_), .ZN(new_n252_) );
  NAND2_X1 g115 ( .A1(new_n252_), .A2(KEYINPUT7), .ZN(new_n253_) );
  INV_X1 g116 ( .A(KEYINPUT7), .ZN(new_n254_) );
  NAND3_X1 g117 ( .A1(new_n250_), .A2(new_n254_), .A3(new_n251_), .ZN(new_n255_) );
  INV_X1 g118 ( .A(G92GAT), .ZN(new_n256_) );
  XNOR2_X1 g119 ( .A(G85GAT), .B(G99GAT), .ZN(new_n257_) );
  NAND2_X1 g120 ( .A1(new_n257_), .A2(new_n256_), .ZN(new_n258_) );
  NAND2_X1 g121 ( .A1(G85GAT), .A2(G99GAT), .ZN(new_n259_) );
  OR2_X1 g122 ( .A1(G85GAT), .A2(G99GAT), .ZN(new_n260_) );
  NAND3_X1 g123 ( .A1(new_n260_), .A2(G92GAT), .A3(new_n259_), .ZN(new_n261_) );
  NAND4_X1 g124 ( .A1(new_n253_), .A2(new_n258_), .A3(new_n255_), .A4(new_n261_), .ZN(new_n262_) );
  NAND2_X1 g125 ( .A1(new_n253_), .A2(new_n255_), .ZN(new_n263_) );
  NAND2_X1 g126 ( .A1(new_n258_), .A2(new_n261_), .ZN(new_n264_) );
  NAND2_X1 g127 ( .A1(new_n263_), .A2(new_n264_), .ZN(new_n265_) );
  NAND2_X1 g128 ( .A1(new_n265_), .A2(new_n262_), .ZN(new_n266_) );
  INV_X1 g129 ( .A(KEYINPUT9), .ZN(new_n267_) );
  OR2_X1 g130 ( .A1(KEYINPUT11), .A2(KEYINPUT10), .ZN(new_n268_) );
  NAND2_X1 g131 ( .A1(KEYINPUT11), .A2(KEYINPUT10), .ZN(new_n269_) );
  NAND2_X1 g132 ( .A1(G232GAT), .A2(G233GAT), .ZN(new_n270_) );
  NAND3_X1 g133 ( .A1(new_n268_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n271_) );
  XNOR2_X1 g134 ( .A(KEYINPUT11), .B(KEYINPUT10), .ZN(new_n272_) );
  INV_X1 g135 ( .A(new_n270_), .ZN(new_n273_) );
  NAND2_X1 g136 ( .A1(new_n272_), .A2(new_n273_), .ZN(new_n274_) );
  NAND3_X1 g137 ( .A1(new_n274_), .A2(new_n267_), .A3(new_n271_), .ZN(new_n275_) );
  NAND2_X1 g138 ( .A1(new_n274_), .A2(new_n271_), .ZN(new_n276_) );
  NAND2_X1 g139 ( .A1(new_n276_), .A2(KEYINPUT9), .ZN(new_n277_) );
  NAND2_X1 g140 ( .A1(new_n277_), .A2(new_n275_), .ZN(new_n278_) );
  NAND2_X1 g141 ( .A1(new_n266_), .A2(new_n278_), .ZN(new_n279_) );
  NAND4_X1 g142 ( .A1(new_n265_), .A2(new_n277_), .A3(new_n262_), .A4(new_n275_), .ZN(new_n280_) );
  XNOR2_X1 g143 ( .A(G106GAT), .B(G218GAT), .ZN(new_n281_) );
  XNOR2_X1 g144 ( .A(new_n151_), .B(new_n281_), .ZN(new_n282_) );
  NAND3_X1 g145 ( .A1(new_n279_), .A2(new_n280_), .A3(new_n282_), .ZN(new_n283_) );
  NAND2_X1 g146 ( .A1(new_n279_), .A2(new_n280_), .ZN(new_n284_) );
  INV_X1 g147 ( .A(new_n282_), .ZN(new_n285_) );
  NAND2_X1 g148 ( .A1(new_n284_), .A2(new_n285_), .ZN(new_n286_) );
  NAND2_X1 g149 ( .A1(new_n286_), .A2(new_n283_), .ZN(new_n287_) );
  NAND2_X1 g150 ( .A1(new_n287_), .A2(new_n180_), .ZN(new_n288_) );
  NAND3_X1 g151 ( .A1(new_n286_), .A2(new_n183_), .A3(new_n283_), .ZN(new_n289_) );
  NAND3_X1 g152 ( .A1(new_n288_), .A2(new_n211_), .A3(new_n289_), .ZN(new_n290_) );
  NAND2_X1 g153 ( .A1(new_n288_), .A2(new_n289_), .ZN(new_n291_) );
  NAND2_X1 g154 ( .A1(new_n291_), .A2(new_n210_), .ZN(new_n292_) );
  NAND3_X1 g155 ( .A1(new_n249_), .A2(new_n290_), .A3(new_n292_), .ZN(new_n293_) );
  XOR2_X1 g156 ( .A(new_n293_), .B(KEYINPUT16), .Z(new_n294_) );
  AND2_X1 g157 ( .A1(new_n233_), .A2(new_n294_), .ZN(new_n295_) );
  INV_X1 g158 ( .A(new_n242_), .ZN(new_n296_) );
  NAND4_X1 g159 ( .A1(new_n175_), .A2(new_n258_), .A3(new_n173_), .A4(new_n261_), .ZN(new_n297_) );
  NAND2_X1 g160 ( .A1(new_n176_), .A2(new_n264_), .ZN(new_n298_) );
  NAND2_X1 g161 ( .A1(new_n298_), .A2(new_n297_), .ZN(new_n299_) );
  INV_X1 g162 ( .A(KEYINPUT32), .ZN(new_n300_) );
  XNOR2_X1 g163 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(new_n301_) );
  NAND2_X1 g164 ( .A1(G230GAT), .A2(G233GAT), .ZN(new_n302_) );
  NAND2_X1 g165 ( .A1(new_n301_), .A2(new_n302_), .ZN(new_n303_) );
  NAND2_X1 g166 ( .A1(KEYINPUT33), .A2(KEYINPUT31), .ZN(new_n304_) );
  OR2_X1 g167 ( .A1(KEYINPUT33), .A2(KEYINPUT31), .ZN(new_n305_) );
  NAND4_X1 g168 ( .A1(new_n305_), .A2(G230GAT), .A3(G233GAT), .A4(new_n304_), .ZN(new_n306_) );
  NAND3_X1 g169 ( .A1(new_n303_), .A2(new_n300_), .A3(new_n306_), .ZN(new_n307_) );
  NAND2_X1 g170 ( .A1(new_n303_), .A2(new_n306_), .ZN(new_n308_) );
  NAND2_X1 g171 ( .A1(new_n308_), .A2(KEYINPUT32), .ZN(new_n309_) );
  NAND2_X1 g172 ( .A1(new_n309_), .A2(new_n307_), .ZN(new_n310_) );
  NAND2_X1 g173 ( .A1(new_n299_), .A2(new_n310_), .ZN(new_n311_) );
  NAND4_X1 g174 ( .A1(new_n298_), .A2(new_n309_), .A3(new_n297_), .A4(new_n307_), .ZN(new_n312_) );
  NAND2_X1 g175 ( .A1(new_n311_), .A2(new_n312_), .ZN(new_n313_) );
  NAND2_X1 g176 ( .A1(new_n313_), .A2(new_n213_), .ZN(new_n314_) );
  INV_X1 g177 ( .A(new_n213_), .ZN(new_n315_) );
  NAND3_X1 g178 ( .A1(new_n311_), .A2(new_n315_), .A3(new_n312_), .ZN(new_n316_) );
  NAND2_X1 g179 ( .A1(new_n314_), .A2(new_n316_), .ZN(new_n317_) );
  XOR2_X1 g180 ( .A(G120GAT), .B(G204GAT), .Z(new_n318_) );
  INV_X1 g181 ( .A(new_n318_), .ZN(new_n319_) );
  NAND2_X1 g182 ( .A1(new_n317_), .A2(new_n319_), .ZN(new_n320_) );
  NAND3_X1 g183 ( .A1(new_n314_), .A2(new_n316_), .A3(new_n318_), .ZN(new_n321_) );
  NAND3_X1 g184 ( .A1(new_n320_), .A2(new_n296_), .A3(new_n321_), .ZN(new_n322_) );
  NAND2_X1 g185 ( .A1(new_n320_), .A2(new_n321_), .ZN(new_n323_) );
  NAND2_X1 g186 ( .A1(new_n323_), .A2(new_n242_), .ZN(new_n324_) );
  XOR2_X1 g187 ( .A(G113GAT), .B(G197GAT), .Z(new_n325_) );
  XNOR2_X1 g188 ( .A(G29GAT), .B(G141GAT), .ZN(new_n326_) );
  XNOR2_X1 g189 ( .A(new_n325_), .B(new_n326_), .ZN(new_n327_) );
  XNOR2_X1 g190 ( .A(G8GAT), .B(G169GAT), .ZN(new_n328_) );
  XNOR2_X1 g191 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(new_n329_) );
  XNOR2_X1 g192 ( .A(new_n328_), .B(new_n329_), .ZN(new_n330_) );
  XNOR2_X1 g193 ( .A(new_n327_), .B(new_n330_), .ZN(new_n331_) );
  XNOR2_X1 g194 ( .A(new_n244_), .B(new_n263_), .ZN(new_n332_) );
  XNOR2_X1 g195 ( .A(new_n331_), .B(new_n332_), .ZN(new_n333_) );
  XOR2_X1 g196 ( .A(G36GAT), .B(G50GAT), .Z(new_n334_) );
  NAND2_X1 g197 ( .A1(G229GAT), .A2(G233GAT), .ZN(new_n335_) );
  XNOR2_X1 g198 ( .A(new_n334_), .B(new_n335_), .ZN(new_n336_) );
  XNOR2_X1 g199 ( .A(new_n333_), .B(new_n336_), .ZN(new_n337_) );
  AND3_X1 g200 ( .A1(new_n324_), .A2(new_n322_), .A3(new_n337_), .ZN(new_n338_) );
  AND2_X1 g201 ( .A1(new_n295_), .A2(new_n338_), .ZN(new_n339_) );
  NAND2_X1 g202 ( .A1(new_n339_), .A2(new_n158_), .ZN(new_n340_) );
  XNOR2_X1 g203 ( .A(new_n340_), .B(KEYINPUT34), .ZN(new_n341_) );
  XNOR2_X1 g204 ( .A(new_n341_), .B(G1GAT), .ZN(G1324GAT) );
  NAND2_X1 g205 ( .A1(new_n339_), .A2(new_n220_), .ZN(new_n343_) );
  XNOR2_X1 g206 ( .A(new_n343_), .B(G8GAT), .ZN(G1325GAT) );
  NAND2_X1 g207 ( .A1(new_n339_), .A2(new_n204_), .ZN(new_n345_) );
  XOR2_X1 g208 ( .A(G15GAT), .B(KEYINPUT35), .Z(new_n346_) );
  XNOR2_X1 g209 ( .A(new_n345_), .B(new_n346_), .ZN(G1326GAT) );
  INV_X1 g210 ( .A(new_n230_), .ZN(new_n348_) );
  NAND2_X1 g211 ( .A1(new_n339_), .A2(new_n348_), .ZN(new_n349_) );
  XNOR2_X1 g212 ( .A(new_n349_), .B(G22GAT), .ZN(G1327GAT) );
  INV_X1 g213 ( .A(KEYINPUT38), .ZN(new_n351_) );
  NAND2_X1 g214 ( .A1(new_n292_), .A2(new_n290_), .ZN(new_n352_) );
  NAND2_X1 g215 ( .A1(new_n352_), .A2(KEYINPUT36), .ZN(new_n353_) );
  INV_X1 g216 ( .A(KEYINPUT36), .ZN(new_n354_) );
  NAND3_X1 g217 ( .A1(new_n292_), .A2(new_n354_), .A3(new_n290_), .ZN(new_n355_) );
  NAND2_X1 g218 ( .A1(new_n353_), .A2(new_n355_), .ZN(new_n356_) );
  INV_X1 g219 ( .A(new_n356_), .ZN(new_n357_) );
  NOR2_X1 g220 ( .A1(new_n357_), .A2(new_n249_), .ZN(new_n358_) );
  NAND2_X1 g221 ( .A1(new_n233_), .A2(new_n358_), .ZN(new_n359_) );
  NAND2_X1 g222 ( .A1(new_n359_), .A2(KEYINPUT37), .ZN(new_n360_) );
  INV_X1 g223 ( .A(KEYINPUT37), .ZN(new_n361_) );
  NAND3_X1 g224 ( .A1(new_n233_), .A2(new_n361_), .A3(new_n358_), .ZN(new_n362_) );
  NAND2_X1 g225 ( .A1(new_n360_), .A2(new_n362_), .ZN(new_n363_) );
  NAND2_X1 g226 ( .A1(new_n363_), .A2(new_n338_), .ZN(new_n364_) );
  NAND2_X1 g227 ( .A1(new_n364_), .A2(new_n351_), .ZN(new_n365_) );
  NAND3_X1 g228 ( .A1(new_n363_), .A2(KEYINPUT38), .A3(new_n338_), .ZN(new_n366_) );
  NAND2_X1 g229 ( .A1(new_n365_), .A2(new_n366_), .ZN(new_n367_) );
  NAND2_X1 g230 ( .A1(new_n367_), .A2(new_n158_), .ZN(new_n368_) );
  XOR2_X1 g231 ( .A(G29GAT), .B(KEYINPUT39), .Z(new_n369_) );
  XNOR2_X1 g232 ( .A(new_n368_), .B(new_n369_), .ZN(G1328GAT) );
  NAND2_X1 g233 ( .A1(new_n367_), .A2(new_n220_), .ZN(new_n371_) );
  XNOR2_X1 g234 ( .A(new_n371_), .B(G36GAT), .ZN(G1329GAT) );
  INV_X1 g235 ( .A(KEYINPUT40), .ZN(new_n373_) );
  NAND2_X1 g236 ( .A1(new_n367_), .A2(new_n204_), .ZN(new_n374_) );
  NAND2_X1 g237 ( .A1(new_n374_), .A2(new_n373_), .ZN(new_n375_) );
  NAND3_X1 g238 ( .A1(new_n367_), .A2(KEYINPUT40), .A3(new_n204_), .ZN(new_n376_) );
  NAND3_X1 g239 ( .A1(new_n375_), .A2(G43GAT), .A3(new_n376_), .ZN(new_n377_) );
  INV_X1 g240 ( .A(G43GAT), .ZN(new_n378_) );
  NAND2_X1 g241 ( .A1(new_n375_), .A2(new_n376_), .ZN(new_n379_) );
  NAND2_X1 g242 ( .A1(new_n379_), .A2(new_n378_), .ZN(new_n380_) );
  NAND2_X1 g243 ( .A1(new_n380_), .A2(new_n377_), .ZN(G1330GAT) );
  NAND2_X1 g244 ( .A1(new_n367_), .A2(new_n348_), .ZN(new_n382_) );
  XNOR2_X1 g245 ( .A(new_n382_), .B(G50GAT), .ZN(G1331GAT) );
  NAND3_X1 g246 ( .A1(new_n324_), .A2(KEYINPUT41), .A3(new_n322_), .ZN(new_n384_) );
  INV_X1 g247 ( .A(KEYINPUT41), .ZN(new_n385_) );
  NAND2_X1 g248 ( .A1(new_n324_), .A2(new_n322_), .ZN(new_n386_) );
  NAND2_X1 g249 ( .A1(new_n386_), .A2(new_n385_), .ZN(new_n387_) );
  NAND2_X1 g250 ( .A1(new_n387_), .A2(new_n384_), .ZN(new_n388_) );
  INV_X1 g251 ( .A(new_n388_), .ZN(new_n389_) );
  NOR2_X1 g252 ( .A1(new_n389_), .A2(new_n337_), .ZN(new_n390_) );
  AND2_X1 g253 ( .A1(new_n295_), .A2(new_n390_), .ZN(new_n391_) );
  NAND2_X1 g254 ( .A1(new_n391_), .A2(new_n158_), .ZN(new_n392_) );
  XNOR2_X1 g255 ( .A(G57GAT), .B(KEYINPUT42), .ZN(new_n393_) );
  XNOR2_X1 g256 ( .A(new_n392_), .B(new_n393_), .ZN(G1332GAT) );
  NAND2_X1 g257 ( .A1(new_n391_), .A2(new_n220_), .ZN(new_n395_) );
  XNOR2_X1 g258 ( .A(new_n395_), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 g259 ( .A1(new_n391_), .A2(new_n204_), .ZN(new_n397_) );
  XNOR2_X1 g260 ( .A(new_n397_), .B(G71GAT), .ZN(G1334GAT) );
  NAND2_X1 g261 ( .A1(new_n391_), .A2(new_n348_), .ZN(new_n399_) );
  XOR2_X1 g262 ( .A(G78GAT), .B(KEYINPUT43), .Z(new_n400_) );
  XNOR2_X1 g263 ( .A(new_n399_), .B(new_n400_), .ZN(G1335GAT) );
  AND2_X1 g264 ( .A1(new_n363_), .A2(new_n390_), .ZN(new_n402_) );
  NAND2_X1 g265 ( .A1(new_n402_), .A2(new_n158_), .ZN(new_n403_) );
  XNOR2_X1 g266 ( .A(new_n403_), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 g267 ( .A1(new_n402_), .A2(new_n220_), .ZN(new_n405_) );
  XNOR2_X1 g268 ( .A(new_n405_), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 g269 ( .A1(new_n402_), .A2(new_n204_), .ZN(new_n407_) );
  XNOR2_X1 g270 ( .A(new_n407_), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 g271 ( .A1(new_n402_), .A2(new_n348_), .ZN(new_n409_) );
  XNOR2_X1 g272 ( .A(new_n409_), .B(KEYINPUT44), .ZN(new_n410_) );
  XNOR2_X1 g273 ( .A(new_n410_), .B(G106GAT), .ZN(G1339GAT) );
  NAND3_X1 g274 ( .A1(new_n388_), .A2(KEYINPUT46), .A3(new_n337_), .ZN(new_n412_) );
  INV_X1 g275 ( .A(KEYINPUT46), .ZN(new_n413_) );
  NAND2_X1 g276 ( .A1(new_n388_), .A2(new_n337_), .ZN(new_n414_) );
  NAND2_X1 g277 ( .A1(new_n414_), .A2(new_n413_), .ZN(new_n415_) );
  NOR2_X1 g278 ( .A1(new_n249_), .A2(new_n352_), .ZN(new_n416_) );
  NAND3_X1 g279 ( .A1(new_n415_), .A2(new_n412_), .A3(new_n416_), .ZN(new_n417_) );
  NAND2_X1 g280 ( .A1(new_n417_), .A2(KEYINPUT47), .ZN(new_n418_) );
  INV_X1 g281 ( .A(KEYINPUT47), .ZN(new_n419_) );
  NAND4_X1 g282 ( .A1(new_n415_), .A2(new_n419_), .A3(new_n412_), .A4(new_n416_), .ZN(new_n420_) );
  NAND3_X1 g283 ( .A1(new_n356_), .A2(KEYINPUT45), .A3(new_n249_), .ZN(new_n421_) );
  INV_X1 g284 ( .A(KEYINPUT45), .ZN(new_n422_) );
  NAND2_X1 g285 ( .A1(new_n356_), .A2(new_n249_), .ZN(new_n423_) );
  NAND2_X1 g286 ( .A1(new_n423_), .A2(new_n422_), .ZN(new_n424_) );
  NAND2_X1 g287 ( .A1(new_n424_), .A2(new_n421_), .ZN(new_n425_) );
  NOR2_X1 g288 ( .A1(new_n386_), .A2(new_n337_), .ZN(new_n426_) );
  NAND2_X1 g289 ( .A1(new_n425_), .A2(new_n426_), .ZN(new_n427_) );
  NAND3_X1 g290 ( .A1(new_n418_), .A2(new_n420_), .A3(new_n427_), .ZN(new_n428_) );
  NAND2_X1 g291 ( .A1(new_n428_), .A2(KEYINPUT48), .ZN(new_n429_) );
  INV_X1 g292 ( .A(KEYINPUT48), .ZN(new_n430_) );
  NAND4_X1 g293 ( .A1(new_n418_), .A2(new_n427_), .A3(new_n430_), .A4(new_n420_), .ZN(new_n431_) );
  NAND2_X1 g294 ( .A1(new_n429_), .A2(new_n431_), .ZN(new_n432_) );
  AND2_X1 g295 ( .A1(new_n432_), .A2(new_n231_), .ZN(new_n433_) );
  AND3_X1 g296 ( .A1(new_n433_), .A2(new_n204_), .A3(new_n230_), .ZN(new_n434_) );
  NAND2_X1 g297 ( .A1(new_n434_), .A2(new_n337_), .ZN(new_n435_) );
  XNOR2_X1 g298 ( .A(new_n435_), .B(G113GAT), .ZN(G1340GAT) );
  NAND2_X1 g299 ( .A1(new_n434_), .A2(new_n388_), .ZN(new_n437_) );
  XOR2_X1 g300 ( .A(G120GAT), .B(KEYINPUT49), .Z(new_n438_) );
  XNOR2_X1 g301 ( .A(new_n437_), .B(new_n438_), .ZN(G1341GAT) );
  NAND2_X1 g302 ( .A1(new_n434_), .A2(new_n249_), .ZN(new_n440_) );
  XNOR2_X1 g303 ( .A(new_n440_), .B(KEYINPUT50), .ZN(new_n441_) );
  XNOR2_X1 g304 ( .A(new_n441_), .B(G127GAT), .ZN(G1342GAT) );
  NAND2_X1 g305 ( .A1(new_n434_), .A2(new_n352_), .ZN(new_n443_) );
  XOR2_X1 g306 ( .A(G134GAT), .B(KEYINPUT51), .Z(new_n444_) );
  XNOR2_X1 g307 ( .A(new_n443_), .B(new_n444_), .ZN(G1343GAT) );
  NAND2_X1 g308 ( .A1(new_n433_), .A2(new_n209_), .ZN(new_n446_) );
  INV_X1 g309 ( .A(new_n446_), .ZN(new_n447_) );
  NAND2_X1 g310 ( .A1(new_n447_), .A2(new_n337_), .ZN(new_n448_) );
  XNOR2_X1 g311 ( .A(new_n448_), .B(G141GAT), .ZN(G1344GAT) );
  NOR2_X1 g312 ( .A1(new_n446_), .A2(new_n389_), .ZN(new_n450_) );
  XOR2_X1 g313 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(new_n451_) );
  XNOR2_X1 g314 ( .A(new_n450_), .B(new_n451_), .ZN(new_n452_) );
  XNOR2_X1 g315 ( .A(new_n452_), .B(new_n170_), .ZN(G1345GAT) );
  NAND2_X1 g316 ( .A1(new_n447_), .A2(new_n249_), .ZN(new_n454_) );
  XNOR2_X1 g317 ( .A(new_n454_), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 g318 ( .A1(new_n447_), .A2(new_n352_), .ZN(new_n456_) );
  XNOR2_X1 g319 ( .A(new_n456_), .B(G162GAT), .ZN(G1347GAT) );
  INV_X1 g320 ( .A(KEYINPUT55), .ZN(new_n458_) );
  INV_X1 g321 ( .A(new_n189_), .ZN(new_n459_) );
  INV_X1 g322 ( .A(KEYINPUT54), .ZN(new_n460_) );
  NAND3_X1 g323 ( .A1(new_n432_), .A2(new_n460_), .A3(new_n220_), .ZN(new_n461_) );
  NAND2_X1 g324 ( .A1(new_n432_), .A2(new_n220_), .ZN(new_n462_) );
  NAND2_X1 g325 ( .A1(new_n462_), .A2(KEYINPUT54), .ZN(new_n463_) );
  AND2_X1 g326 ( .A1(new_n463_), .A2(new_n159_), .ZN(new_n464_) );
  NAND4_X1 g327 ( .A1(new_n464_), .A2(new_n458_), .A3(new_n459_), .A4(new_n461_), .ZN(new_n465_) );
  NAND4_X1 g328 ( .A1(new_n463_), .A2(new_n159_), .A3(new_n459_), .A4(new_n461_), .ZN(new_n466_) );
  NAND2_X1 g329 ( .A1(new_n466_), .A2(KEYINPUT55), .ZN(new_n467_) );
  NAND2_X1 g330 ( .A1(new_n465_), .A2(new_n467_), .ZN(new_n468_) );
  NAND3_X1 g331 ( .A1(new_n468_), .A2(new_n204_), .A3(new_n337_), .ZN(new_n469_) );
  XNOR2_X1 g332 ( .A(new_n469_), .B(G169GAT), .ZN(G1348GAT) );
  XNOR2_X1 g333 ( .A(KEYINPUT57), .B(KEYINPUT56), .ZN(new_n471_) );
  INV_X1 g334 ( .A(new_n471_), .ZN(new_n472_) );
  NAND4_X1 g335 ( .A1(new_n468_), .A2(new_n204_), .A3(new_n388_), .A4(new_n472_), .ZN(new_n473_) );
  NAND3_X1 g336 ( .A1(new_n468_), .A2(new_n204_), .A3(new_n388_), .ZN(new_n474_) );
  NAND2_X1 g337 ( .A1(new_n474_), .A2(new_n471_), .ZN(new_n475_) );
  NAND3_X1 g338 ( .A1(new_n475_), .A2(G176GAT), .A3(new_n473_), .ZN(new_n476_) );
  INV_X1 g339 ( .A(G176GAT), .ZN(new_n477_) );
  NAND2_X1 g340 ( .A1(new_n475_), .A2(new_n473_), .ZN(new_n478_) );
  NAND2_X1 g341 ( .A1(new_n478_), .A2(new_n477_), .ZN(new_n479_) );
  NAND2_X1 g342 ( .A1(new_n479_), .A2(new_n476_), .ZN(G1349GAT) );
  NAND3_X1 g343 ( .A1(new_n468_), .A2(new_n204_), .A3(new_n249_), .ZN(new_n481_) );
  XNOR2_X1 g344 ( .A(new_n481_), .B(G183GAT), .ZN(G1350GAT) );
  NAND3_X1 g345 ( .A1(new_n468_), .A2(new_n204_), .A3(new_n352_), .ZN(new_n483_) );
  XNOR2_X1 g346 ( .A(G190GAT), .B(KEYINPUT58), .ZN(new_n484_) );
  XNOR2_X1 g347 ( .A(new_n483_), .B(new_n484_), .ZN(G1351GAT) );
  NAND4_X1 g348 ( .A1(new_n464_), .A2(new_n209_), .A3(new_n337_), .A4(new_n461_), .ZN(new_n486_) );
  XNOR2_X1 g349 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(new_n487_) );
  NAND2_X1 g350 ( .A1(new_n486_), .A2(new_n487_), .ZN(new_n488_) );
  OR2_X1 g351 ( .A1(new_n486_), .A2(new_n487_), .ZN(new_n489_) );
  NAND2_X1 g352 ( .A1(new_n489_), .A2(new_n488_), .ZN(new_n490_) );
  XNOR2_X1 g353 ( .A(new_n490_), .B(new_n161_), .ZN(G1352GAT) );
  INV_X1 g354 ( .A(new_n209_), .ZN(new_n492_) );
  NAND2_X1 g355 ( .A1(new_n464_), .A2(new_n461_), .ZN(new_n493_) );
  NOR2_X1 g356 ( .A1(new_n493_), .A2(new_n492_), .ZN(new_n494_) );
  NAND2_X1 g357 ( .A1(new_n494_), .A2(new_n386_), .ZN(new_n495_) );
  XOR2_X1 g358 ( .A(G204GAT), .B(KEYINPUT61), .Z(new_n496_) );
  XNOR2_X1 g359 ( .A(new_n495_), .B(new_n496_), .ZN(G1353GAT) );
  NAND2_X1 g360 ( .A1(new_n494_), .A2(new_n249_), .ZN(new_n498_) );
  XNOR2_X1 g361 ( .A(new_n498_), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 g362 ( .A(G218GAT), .ZN(new_n500_) );
  NOR3_X1 g363 ( .A1(new_n493_), .A2(new_n492_), .A3(new_n357_), .ZN(new_n501_) );
  NAND2_X1 g364 ( .A1(new_n501_), .A2(KEYINPUT62), .ZN(new_n502_) );
  OR2_X1 g365 ( .A1(new_n501_), .A2(KEYINPUT62), .ZN(new_n503_) );
  NAND2_X1 g366 ( .A1(new_n503_), .A2(new_n502_), .ZN(new_n504_) );
  NAND2_X1 g367 ( .A1(new_n504_), .A2(new_n500_), .ZN(new_n505_) );
  NAND3_X1 g368 ( .A1(new_n503_), .A2(new_n502_), .A3(G218GAT), .ZN(new_n506_) );
  NAND2_X1 g369 ( .A1(new_n505_), .A2(new_n506_), .ZN(G1355GAT) );
endmodule


