module add_mul_comp_8_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, Result_0_, Result_1_, 
        Result_2_, Result_3_, Result_4_, Result_5_, Result_6_, Result_7_, 
        Result_8_, Result_9_, Result_10_, Result_11_, Result_12_, Result_13_, 
        Result_14_, Result_15_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_,
         b_4_, b_5_, b_6_, b_7_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_;
  wire   n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951;

  NAND2_X1 U479 ( .A1(n463), .A2(n464), .ZN(Result_9_) );
  NAND2_X1 U480 ( .A1(n465), .A2(n466), .ZN(n464) );
  XNOR2_X1 U481 ( .A(n467), .B(n468), .ZN(n465) );
  XNOR2_X1 U482 ( .A(n469), .B(n470), .ZN(n468) );
  NAND2_X1 U483 ( .A1(n471), .A2(n472), .ZN(n463) );
  NAND2_X1 U484 ( .A1(n473), .A2(n474), .ZN(n472) );
  NAND2_X1 U485 ( .A1(n475), .A2(n476), .ZN(n474) );
  OR2_X1 U486 ( .A1(n477), .A2(n478), .ZN(n475) );
  NAND2_X1 U487 ( .A1(n479), .A2(n480), .ZN(n473) );
  XOR2_X1 U488 ( .A(b_1_), .B(a_1_), .Z(n479) );
  NAND2_X1 U489 ( .A1(n481), .A2(n482), .ZN(Result_8_) );
  NAND2_X1 U490 ( .A1(n483), .A2(n466), .ZN(n482) );
  XOR2_X1 U491 ( .A(n484), .B(n485), .Z(n483) );
  XOR2_X1 U492 ( .A(n486), .B(n487), .Z(n484) );
  NOR2_X1 U493 ( .A1(n488), .A2(n489), .ZN(n487) );
  NAND2_X1 U494 ( .A1(n490), .A2(n471), .ZN(n481) );
  XNOR2_X1 U495 ( .A(n491), .B(n492), .ZN(n490) );
  NOR2_X1 U496 ( .A1(n478), .A2(n493), .ZN(n491) );
  NOR2_X1 U497 ( .A1(n477), .A2(n476), .ZN(n493) );
  INV_X1 U498 ( .A(n480), .ZN(n476) );
  NOR2_X1 U499 ( .A1(n494), .A2(n495), .ZN(n480) );
  NOR2_X1 U500 ( .A1(n496), .A2(n497), .ZN(n495) );
  NOR2_X1 U501 ( .A1(b_1_), .A2(a_1_), .ZN(n478) );
  NOR2_X1 U502 ( .A1(n471), .A2(n498), .ZN(Result_7_) );
  XNOR2_X1 U503 ( .A(n499), .B(n500), .ZN(n498) );
  NOR3_X1 U504 ( .A1(n501), .A2(n502), .A3(n471), .ZN(Result_6_) );
  NOR2_X1 U505 ( .A1(n503), .A2(n504), .ZN(n501) );
  NOR2_X1 U506 ( .A1(n500), .A2(n499), .ZN(n503) );
  NOR2_X1 U507 ( .A1(n471), .A2(n505), .ZN(Result_5_) );
  XNOR2_X1 U508 ( .A(n502), .B(n506), .ZN(n505) );
  NOR2_X1 U509 ( .A1(n507), .A2(n508), .ZN(n506) );
  NOR2_X1 U510 ( .A1(n509), .A2(n510), .ZN(n508) );
  NOR2_X1 U511 ( .A1(n511), .A2(n512), .ZN(n509) );
  NOR2_X1 U512 ( .A1(n471), .A2(n513), .ZN(Result_4_) );
  XNOR2_X1 U513 ( .A(n514), .B(n515), .ZN(n513) );
  NOR2_X1 U514 ( .A1(n471), .A2(n516), .ZN(Result_3_) );
  XOR2_X1 U515 ( .A(n517), .B(n518), .Z(n516) );
  NAND2_X1 U516 ( .A1(n519), .A2(n520), .ZN(n517) );
  NOR2_X1 U517 ( .A1(n471), .A2(n521), .ZN(Result_2_) );
  XOR2_X1 U518 ( .A(n522), .B(n523), .Z(n521) );
  NAND2_X1 U519 ( .A1(n524), .A2(n525), .ZN(n523) );
  NOR2_X1 U520 ( .A1(n471), .A2(n526), .ZN(Result_1_) );
  XNOR2_X1 U521 ( .A(n527), .B(n528), .ZN(n526) );
  NAND2_X1 U522 ( .A1(n529), .A2(n530), .ZN(n528) );
  INV_X1 U523 ( .A(n531), .ZN(n530) );
  NAND2_X1 U524 ( .A1(n532), .A2(n533), .ZN(n529) );
  NAND2_X1 U525 ( .A1(b_0_), .A2(n534), .ZN(n533) );
  NAND2_X1 U526 ( .A1(n535), .A2(n536), .ZN(Result_15_) );
  NAND2_X1 U527 ( .A1(n537), .A2(n466), .ZN(n536) );
  NAND2_X1 U528 ( .A1(n471), .A2(n538), .ZN(n535) );
  NAND2_X1 U529 ( .A1(n539), .A2(n540), .ZN(n538) );
  NAND2_X1 U530 ( .A1(b_7_), .A2(n541), .ZN(n540) );
  NAND2_X1 U531 ( .A1(n542), .A2(n543), .ZN(Result_14_) );
  NAND2_X1 U532 ( .A1(n471), .A2(n544), .ZN(n543) );
  NAND3_X1 U533 ( .A1(n545), .A2(n546), .A3(n547), .ZN(n544) );
  NAND2_X1 U534 ( .A1(n548), .A2(n549), .ZN(n546) );
  XOR2_X1 U535 ( .A(n550), .B(n551), .Z(n548) );
  NAND3_X1 U536 ( .A1(n551), .A2(n550), .A3(b_6_), .ZN(n545) );
  NAND2_X1 U537 ( .A1(n552), .A2(n466), .ZN(n542) );
  XOR2_X1 U538 ( .A(n553), .B(n554), .Z(n552) );
  NAND2_X1 U539 ( .A1(b_7_), .A2(a_6_), .ZN(n554) );
  NAND2_X1 U540 ( .A1(n555), .A2(n556), .ZN(Result_13_) );
  NAND2_X1 U541 ( .A1(n471), .A2(n557), .ZN(n556) );
  NAND3_X1 U542 ( .A1(n558), .A2(n559), .A3(n560), .ZN(n557) );
  NAND2_X1 U543 ( .A1(n561), .A2(n562), .ZN(n560) );
  NAND3_X1 U544 ( .A1(n563), .A2(n564), .A3(b_5_), .ZN(n559) );
  NAND2_X1 U545 ( .A1(n565), .A2(n566), .ZN(n558) );
  XOR2_X1 U546 ( .A(n564), .B(n563), .Z(n565) );
  INV_X1 U547 ( .A(n562), .ZN(n563) );
  NAND2_X1 U548 ( .A1(n567), .A2(n466), .ZN(n555) );
  XOR2_X1 U549 ( .A(n568), .B(n569), .Z(n567) );
  XNOR2_X1 U550 ( .A(n570), .B(n547), .ZN(n569) );
  NAND2_X1 U551 ( .A1(b_7_), .A2(a_5_), .ZN(n570) );
  NAND2_X1 U552 ( .A1(n571), .A2(n572), .ZN(Result_12_) );
  NAND2_X1 U553 ( .A1(n573), .A2(n466), .ZN(n572) );
  XNOR2_X1 U554 ( .A(n574), .B(n575), .ZN(n573) );
  NAND2_X1 U555 ( .A1(n576), .A2(n577), .ZN(n574) );
  NAND2_X1 U556 ( .A1(n471), .A2(n578), .ZN(n571) );
  XNOR2_X1 U557 ( .A(n579), .B(n580), .ZN(n578) );
  NAND2_X1 U558 ( .A1(n581), .A2(n582), .ZN(n579) );
  NAND2_X1 U559 ( .A1(n583), .A2(n584), .ZN(Result_11_) );
  NAND2_X1 U560 ( .A1(n471), .A2(n585), .ZN(n584) );
  NAND3_X1 U561 ( .A1(n586), .A2(n587), .A3(n588), .ZN(n585) );
  NAND2_X1 U562 ( .A1(n589), .A2(n590), .ZN(n588) );
  OR3_X1 U563 ( .A1(n590), .A2(a_3_), .A3(n591), .ZN(n587) );
  NAND2_X1 U564 ( .A1(n592), .A2(n591), .ZN(n586) );
  XOR2_X1 U565 ( .A(n590), .B(a_3_), .Z(n592) );
  NAND2_X1 U566 ( .A1(n593), .A2(n466), .ZN(n583) );
  XOR2_X1 U567 ( .A(n594), .B(n595), .Z(n593) );
  XNOR2_X1 U568 ( .A(n596), .B(n597), .ZN(n595) );
  NAND2_X1 U569 ( .A1(b_7_), .A2(a_3_), .ZN(n597) );
  NAND2_X1 U570 ( .A1(n598), .A2(n599), .ZN(Result_10_) );
  NAND2_X1 U571 ( .A1(n600), .A2(n466), .ZN(n599) );
  XOR2_X1 U572 ( .A(n601), .B(n602), .Z(n600) );
  XOR2_X1 U573 ( .A(n603), .B(n604), .Z(n602) );
  NAND2_X1 U574 ( .A1(n471), .A2(n605), .ZN(n598) );
  XNOR2_X1 U575 ( .A(n497), .B(n606), .ZN(n605) );
  NOR2_X1 U576 ( .A1(n496), .A2(n494), .ZN(n606) );
  NOR2_X1 U577 ( .A1(b_2_), .A2(a_2_), .ZN(n496) );
  AND2_X1 U578 ( .A1(n607), .A2(n608), .ZN(n497) );
  NAND2_X1 U579 ( .A1(n609), .A2(n590), .ZN(n608) );
  NAND2_X1 U580 ( .A1(n581), .A2(n610), .ZN(n590) );
  NAND2_X1 U581 ( .A1(n582), .A2(n580), .ZN(n610) );
  NAND2_X1 U582 ( .A1(n611), .A2(n612), .ZN(n580) );
  NAND2_X1 U583 ( .A1(n613), .A2(n562), .ZN(n612) );
  NAND2_X1 U584 ( .A1(n614), .A2(n615), .ZN(n562) );
  NAND2_X1 U585 ( .A1(n537), .A2(n616), .ZN(n615) );
  NAND2_X1 U586 ( .A1(n549), .A2(n550), .ZN(n616) );
  NAND2_X1 U587 ( .A1(n566), .A2(n564), .ZN(n613) );
  NAND2_X1 U588 ( .A1(n617), .A2(n618), .ZN(n582) );
  NAND2_X1 U589 ( .A1(n591), .A2(n619), .ZN(n609) );
  NOR2_X1 U590 ( .A1(n471), .A2(n620), .ZN(Result_0_) );
  NOR3_X1 U591 ( .A1(n621), .A2(n531), .A3(n622), .ZN(n620) );
  NOR3_X1 U592 ( .A1(n623), .A2(n622), .A3(n532), .ZN(n531) );
  INV_X1 U593 ( .A(n534), .ZN(n622) );
  NAND2_X1 U594 ( .A1(n624), .A2(n625), .ZN(n534) );
  NOR2_X1 U595 ( .A1(n527), .A2(n623), .ZN(n621) );
  AND2_X1 U596 ( .A1(n626), .A2(n524), .ZN(n527) );
  NAND4_X1 U597 ( .A1(n627), .A2(n628), .A3(n629), .A4(n532), .ZN(n524) );
  NAND2_X1 U598 ( .A1(n630), .A2(n631), .ZN(n532) );
  OR2_X1 U599 ( .A1(n630), .A2(n631), .ZN(n628) );
  NAND2_X1 U600 ( .A1(n525), .A2(n522), .ZN(n626) );
  NAND2_X1 U601 ( .A1(n519), .A2(n632), .ZN(n522) );
  NAND2_X1 U602 ( .A1(n518), .A2(n520), .ZN(n632) );
  NAND2_X1 U603 ( .A1(n633), .A2(n634), .ZN(n520) );
  NAND2_X1 U604 ( .A1(n635), .A2(n636), .ZN(n634) );
  XNOR2_X1 U605 ( .A(n629), .B(n627), .ZN(n633) );
  AND2_X1 U606 ( .A1(n515), .A2(n514), .ZN(n518) );
  NAND3_X1 U607 ( .A1(n637), .A2(n638), .A3(n639), .ZN(n514) );
  NAND2_X1 U608 ( .A1(n502), .A2(n510), .ZN(n639) );
  INV_X1 U609 ( .A(n640), .ZN(n510) );
  NOR3_X1 U610 ( .A1(n641), .A2(n500), .A3(n499), .ZN(n502) );
  XNOR2_X1 U611 ( .A(n642), .B(n643), .ZN(n499) );
  XOR2_X1 U612 ( .A(n644), .B(n645), .Z(n642) );
  NOR2_X1 U613 ( .A1(n549), .A2(n488), .ZN(n645) );
  AND2_X1 U614 ( .A1(n646), .A2(n647), .ZN(n500) );
  NAND3_X1 U615 ( .A1(a_0_), .A2(n648), .A3(b_7_), .ZN(n647) );
  OR2_X1 U616 ( .A1(n485), .A2(n486), .ZN(n648) );
  NAND2_X1 U617 ( .A1(n485), .A2(n486), .ZN(n646) );
  NAND2_X1 U618 ( .A1(n649), .A2(n650), .ZN(n486) );
  NAND2_X1 U619 ( .A1(n470), .A2(n651), .ZN(n650) );
  OR2_X1 U620 ( .A1(n469), .A2(n467), .ZN(n651) );
  NOR2_X1 U621 ( .A1(n489), .A2(n652), .ZN(n470) );
  NAND2_X1 U622 ( .A1(n467), .A2(n469), .ZN(n649) );
  NAND2_X1 U623 ( .A1(n653), .A2(n654), .ZN(n469) );
  NAND2_X1 U624 ( .A1(n604), .A2(n655), .ZN(n654) );
  NAND2_X1 U625 ( .A1(n603), .A2(n601), .ZN(n655) );
  NOR2_X1 U626 ( .A1(n489), .A2(n656), .ZN(n604) );
  OR2_X1 U627 ( .A1(n601), .A2(n603), .ZN(n653) );
  AND2_X1 U628 ( .A1(n657), .A2(n658), .ZN(n603) );
  NAND3_X1 U629 ( .A1(a_3_), .A2(n659), .A3(b_7_), .ZN(n658) );
  NAND2_X1 U630 ( .A1(n596), .A2(n594), .ZN(n659) );
  OR2_X1 U631 ( .A1(n594), .A2(n596), .ZN(n657) );
  AND2_X1 U632 ( .A1(n576), .A2(n660), .ZN(n596) );
  NAND2_X1 U633 ( .A1(n575), .A2(n577), .ZN(n660) );
  NAND2_X1 U634 ( .A1(n661), .A2(n662), .ZN(n577) );
  NAND2_X1 U635 ( .A1(b_7_), .A2(a_4_), .ZN(n662) );
  INV_X1 U636 ( .A(n663), .ZN(n661) );
  XNOR2_X1 U637 ( .A(n664), .B(n665), .ZN(n575) );
  NAND2_X1 U638 ( .A1(n666), .A2(n667), .ZN(n664) );
  NAND2_X1 U639 ( .A1(a_4_), .A2(n663), .ZN(n576) );
  NAND2_X1 U640 ( .A1(n668), .A2(n669), .ZN(n663) );
  NAND3_X1 U641 ( .A1(a_5_), .A2(n670), .A3(b_7_), .ZN(n669) );
  NAND2_X1 U642 ( .A1(n568), .A2(n547), .ZN(n670) );
  OR2_X1 U643 ( .A1(n547), .A2(n568), .ZN(n668) );
  XOR2_X1 U644 ( .A(n614), .B(n671), .Z(n568) );
  NOR2_X1 U645 ( .A1(n541), .A2(n566), .ZN(n671) );
  NAND2_X1 U646 ( .A1(n672), .A2(n537), .ZN(n547) );
  INV_X1 U647 ( .A(n551), .ZN(n537) );
  NAND2_X1 U648 ( .A1(b_7_), .A2(a_7_), .ZN(n551) );
  INV_X1 U649 ( .A(n614), .ZN(n672) );
  NAND2_X1 U650 ( .A1(b_6_), .A2(a_6_), .ZN(n614) );
  XNOR2_X1 U651 ( .A(n673), .B(n674), .ZN(n594) );
  XOR2_X1 U652 ( .A(n675), .B(n676), .Z(n673) );
  XNOR2_X1 U653 ( .A(n677), .B(n678), .ZN(n601) );
  XNOR2_X1 U654 ( .A(n679), .B(n680), .ZN(n677) );
  NAND2_X1 U655 ( .A1(a_3_), .A2(b_6_), .ZN(n679) );
  XNOR2_X1 U656 ( .A(n681), .B(n682), .ZN(n467) );
  XOR2_X1 U657 ( .A(n683), .B(n684), .Z(n682) );
  NAND2_X1 U658 ( .A1(a_2_), .A2(b_6_), .ZN(n684) );
  XOR2_X1 U659 ( .A(n685), .B(n686), .Z(n485) );
  XOR2_X1 U660 ( .A(n687), .B(n688), .Z(n685) );
  NOR2_X1 U661 ( .A1(n652), .A2(n549), .ZN(n688) );
  INV_X1 U662 ( .A(n504), .ZN(n641) );
  XOR2_X1 U663 ( .A(n511), .B(n512), .Z(n504) );
  INV_X1 U664 ( .A(n507), .ZN(n637) );
  NOR3_X1 U665 ( .A1(n512), .A2(n511), .A3(n640), .ZN(n507) );
  NAND2_X1 U666 ( .A1(n689), .A2(n638), .ZN(n640) );
  NAND2_X1 U667 ( .A1(n690), .A2(n691), .ZN(n638) );
  XNOR2_X1 U668 ( .A(n692), .B(n693), .ZN(n690) );
  NAND2_X1 U669 ( .A1(n694), .A2(n695), .ZN(n689) );
  INV_X1 U670 ( .A(n691), .ZN(n695) );
  NAND2_X1 U671 ( .A1(n696), .A2(n697), .ZN(n691) );
  NAND3_X1 U672 ( .A1(b_5_), .A2(n698), .A3(a_0_), .ZN(n697) );
  OR2_X1 U673 ( .A1(n699), .A2(n700), .ZN(n698) );
  NAND2_X1 U674 ( .A1(n699), .A2(n700), .ZN(n696) );
  XOR2_X1 U675 ( .A(n693), .B(n692), .Z(n694) );
  XOR2_X1 U676 ( .A(n701), .B(n702), .Z(n692) );
  AND2_X1 U677 ( .A1(n703), .A2(n704), .ZN(n511) );
  NAND3_X1 U678 ( .A1(b_6_), .A2(n705), .A3(a_0_), .ZN(n704) );
  OR2_X1 U679 ( .A1(n643), .A2(n644), .ZN(n705) );
  NAND2_X1 U680 ( .A1(n643), .A2(n644), .ZN(n703) );
  NAND2_X1 U681 ( .A1(n706), .A2(n707), .ZN(n644) );
  NAND3_X1 U682 ( .A1(a_1_), .A2(n708), .A3(b_6_), .ZN(n707) );
  OR2_X1 U683 ( .A1(n687), .A2(n686), .ZN(n708) );
  NAND2_X1 U684 ( .A1(n686), .A2(n687), .ZN(n706) );
  NAND2_X1 U685 ( .A1(n709), .A2(n710), .ZN(n687) );
  NAND3_X1 U686 ( .A1(b_6_), .A2(n711), .A3(a_2_), .ZN(n710) );
  OR2_X1 U687 ( .A1(n681), .A2(n683), .ZN(n711) );
  NAND2_X1 U688 ( .A1(n681), .A2(n683), .ZN(n709) );
  NAND2_X1 U689 ( .A1(n712), .A2(n713), .ZN(n683) );
  NAND3_X1 U690 ( .A1(b_6_), .A2(n714), .A3(a_3_), .ZN(n713) );
  OR2_X1 U691 ( .A1(n680), .A2(n678), .ZN(n714) );
  NAND2_X1 U692 ( .A1(n678), .A2(n680), .ZN(n712) );
  NAND2_X1 U693 ( .A1(n715), .A2(n716), .ZN(n680) );
  NAND2_X1 U694 ( .A1(n676), .A2(n717), .ZN(n716) );
  OR2_X1 U695 ( .A1(n675), .A2(n674), .ZN(n717) );
  NOR2_X1 U696 ( .A1(n618), .A2(n549), .ZN(n676) );
  INV_X1 U697 ( .A(b_6_), .ZN(n549) );
  NAND2_X1 U698 ( .A1(n674), .A2(n675), .ZN(n715) );
  NAND2_X1 U699 ( .A1(n666), .A2(n718), .ZN(n675) );
  NAND2_X1 U700 ( .A1(n665), .A2(n667), .ZN(n718) );
  NAND2_X1 U701 ( .A1(n719), .A2(n720), .ZN(n667) );
  INV_X1 U702 ( .A(n721), .ZN(n720) );
  NAND2_X1 U703 ( .A1(a_5_), .A2(b_6_), .ZN(n719) );
  XNOR2_X1 U704 ( .A(n722), .B(n723), .ZN(n665) );
  NOR2_X1 U705 ( .A1(n541), .A2(n617), .ZN(n723) );
  NAND2_X1 U706 ( .A1(n721), .A2(a_5_), .ZN(n666) );
  NOR2_X1 U707 ( .A1(n553), .A2(n722), .ZN(n721) );
  NAND2_X1 U708 ( .A1(b_6_), .A2(a_7_), .ZN(n553) );
  XNOR2_X1 U709 ( .A(n724), .B(n725), .ZN(n674) );
  XOR2_X1 U710 ( .A(n726), .B(n561), .Z(n725) );
  XNOR2_X1 U711 ( .A(n727), .B(n728), .ZN(n678) );
  NAND2_X1 U712 ( .A1(n729), .A2(n730), .ZN(n727) );
  XOR2_X1 U713 ( .A(n731), .B(n732), .Z(n681) );
  XOR2_X1 U714 ( .A(n733), .B(n734), .Z(n731) );
  NOR2_X1 U715 ( .A1(n566), .A2(n619), .ZN(n734) );
  XNOR2_X1 U716 ( .A(n735), .B(n736), .ZN(n686) );
  XOR2_X1 U717 ( .A(n737), .B(n738), .Z(n736) );
  NAND2_X1 U718 ( .A1(a_2_), .A2(b_5_), .ZN(n738) );
  XOR2_X1 U719 ( .A(n739), .B(n740), .Z(n643) );
  XOR2_X1 U720 ( .A(n741), .B(n742), .Z(n739) );
  NOR2_X1 U721 ( .A1(n652), .A2(n566), .ZN(n742) );
  XNOR2_X1 U722 ( .A(n743), .B(n699), .ZN(n512) );
  XNOR2_X1 U723 ( .A(n744), .B(n745), .ZN(n699) );
  NAND2_X1 U724 ( .A1(n746), .A2(n747), .ZN(n744) );
  XNOR2_X1 U725 ( .A(n748), .B(n700), .ZN(n743) );
  NAND2_X1 U726 ( .A1(n749), .A2(n750), .ZN(n700) );
  NAND3_X1 U727 ( .A1(a_1_), .A2(n751), .A3(b_5_), .ZN(n750) );
  OR2_X1 U728 ( .A1(n741), .A2(n740), .ZN(n751) );
  NAND2_X1 U729 ( .A1(n740), .A2(n741), .ZN(n749) );
  NAND2_X1 U730 ( .A1(n752), .A2(n753), .ZN(n741) );
  NAND3_X1 U731 ( .A1(b_5_), .A2(n754), .A3(a_2_), .ZN(n753) );
  OR2_X1 U732 ( .A1(n735), .A2(n737), .ZN(n754) );
  NAND2_X1 U733 ( .A1(n735), .A2(n737), .ZN(n752) );
  NAND2_X1 U734 ( .A1(n755), .A2(n756), .ZN(n737) );
  NAND3_X1 U735 ( .A1(b_5_), .A2(n757), .A3(a_3_), .ZN(n756) );
  OR2_X1 U736 ( .A1(n733), .A2(n732), .ZN(n757) );
  NAND2_X1 U737 ( .A1(n732), .A2(n733), .ZN(n755) );
  NAND2_X1 U738 ( .A1(n729), .A2(n758), .ZN(n733) );
  NAND2_X1 U739 ( .A1(n728), .A2(n730), .ZN(n758) );
  NAND2_X1 U740 ( .A1(n759), .A2(n760), .ZN(n730) );
  NAND2_X1 U741 ( .A1(a_4_), .A2(b_5_), .ZN(n760) );
  INV_X1 U742 ( .A(n761), .ZN(n759) );
  XNOR2_X1 U743 ( .A(n762), .B(n763), .ZN(n728) );
  NAND2_X1 U744 ( .A1(n764), .A2(n765), .ZN(n762) );
  NAND2_X1 U745 ( .A1(a_4_), .A2(n761), .ZN(n729) );
  NAND2_X1 U746 ( .A1(n766), .A2(n767), .ZN(n761) );
  NAND2_X1 U747 ( .A1(n726), .A2(n768), .ZN(n767) );
  NAND2_X1 U748 ( .A1(n724), .A2(n611), .ZN(n768) );
  NOR3_X1 U749 ( .A1(n617), .A2(n541), .A3(n722), .ZN(n726) );
  NAND2_X1 U750 ( .A1(b_5_), .A2(a_6_), .ZN(n722) );
  NAND2_X1 U751 ( .A1(n561), .A2(n769), .ZN(n766) );
  INV_X1 U752 ( .A(n724), .ZN(n769) );
  XNOR2_X1 U753 ( .A(n770), .B(n771), .ZN(n724) );
  INV_X1 U754 ( .A(n611), .ZN(n561) );
  NAND2_X1 U755 ( .A1(a_5_), .A2(b_5_), .ZN(n611) );
  XNOR2_X1 U756 ( .A(n772), .B(n773), .ZN(n732) );
  XOR2_X1 U757 ( .A(n774), .B(n775), .Z(n772) );
  XNOR2_X1 U758 ( .A(n776), .B(n777), .ZN(n735) );
  XOR2_X1 U759 ( .A(n778), .B(n779), .Z(n777) );
  XNOR2_X1 U760 ( .A(n780), .B(n781), .ZN(n740) );
  NAND2_X1 U761 ( .A1(n782), .A2(n783), .ZN(n780) );
  NAND2_X1 U762 ( .A1(a_0_), .A2(b_5_), .ZN(n748) );
  XOR2_X1 U763 ( .A(n635), .B(n636), .Z(n515) );
  NAND3_X1 U764 ( .A1(n635), .A2(n636), .A3(n784), .ZN(n519) );
  XOR2_X1 U765 ( .A(n629), .B(n627), .Z(n784) );
  XNOR2_X1 U766 ( .A(n785), .B(n786), .ZN(n636) );
  XOR2_X1 U767 ( .A(n787), .B(n788), .Z(n786) );
  NAND2_X1 U768 ( .A1(a_0_), .A2(b_3_), .ZN(n788) );
  AND2_X1 U769 ( .A1(n789), .A2(n790), .ZN(n635) );
  NAND2_X1 U770 ( .A1(n701), .A2(n791), .ZN(n790) );
  NAND2_X1 U771 ( .A1(n693), .A2(n702), .ZN(n791) );
  AND2_X1 U772 ( .A1(n746), .A2(n792), .ZN(n701) );
  NAND2_X1 U773 ( .A1(n745), .A2(n747), .ZN(n792) );
  NAND2_X1 U774 ( .A1(n793), .A2(n794), .ZN(n747) );
  NAND2_X1 U775 ( .A1(b_4_), .A2(a_1_), .ZN(n794) );
  INV_X1 U776 ( .A(n795), .ZN(n793) );
  XNOR2_X1 U777 ( .A(n796), .B(n797), .ZN(n745) );
  NAND2_X1 U778 ( .A1(n798), .A2(n799), .ZN(n796) );
  NAND2_X1 U779 ( .A1(a_1_), .A2(n795), .ZN(n746) );
  NAND2_X1 U780 ( .A1(n782), .A2(n800), .ZN(n795) );
  NAND2_X1 U781 ( .A1(n781), .A2(n783), .ZN(n800) );
  NAND2_X1 U782 ( .A1(n801), .A2(n802), .ZN(n783) );
  NAND2_X1 U783 ( .A1(a_2_), .A2(b_4_), .ZN(n802) );
  XNOR2_X1 U784 ( .A(n803), .B(n804), .ZN(n781) );
  XOR2_X1 U785 ( .A(n805), .B(n589), .Z(n803) );
  INV_X1 U786 ( .A(n607), .ZN(n589) );
  OR2_X1 U787 ( .A1(n801), .A2(n656), .ZN(n782) );
  NAND2_X1 U788 ( .A1(n806), .A2(n807), .ZN(n801) );
  NAND2_X1 U789 ( .A1(n776), .A2(n808), .ZN(n807) );
  OR2_X1 U790 ( .A1(n779), .A2(n778), .ZN(n808) );
  XOR2_X1 U791 ( .A(n809), .B(n810), .Z(n776) );
  NAND2_X1 U792 ( .A1(n811), .A2(n812), .ZN(n809) );
  NAND2_X1 U793 ( .A1(n779), .A2(n778), .ZN(n806) );
  NAND2_X1 U794 ( .A1(n813), .A2(n814), .ZN(n778) );
  NAND2_X1 U795 ( .A1(n773), .A2(n815), .ZN(n814) );
  NAND2_X1 U796 ( .A1(n775), .A2(n774), .ZN(n815) );
  XOR2_X1 U797 ( .A(n816), .B(n817), .Z(n773) );
  NAND2_X1 U798 ( .A1(n818), .A2(n819), .ZN(n816) );
  OR2_X1 U799 ( .A1(n774), .A2(n775), .ZN(n813) );
  INV_X1 U800 ( .A(n581), .ZN(n775) );
  NAND2_X1 U801 ( .A1(b_4_), .A2(a_4_), .ZN(n581) );
  NAND2_X1 U802 ( .A1(n764), .A2(n820), .ZN(n774) );
  NAND2_X1 U803 ( .A1(n763), .A2(n765), .ZN(n820) );
  NAND2_X1 U804 ( .A1(n821), .A2(n822), .ZN(n765) );
  NAND2_X1 U805 ( .A1(b_4_), .A2(a_5_), .ZN(n822) );
  AND2_X1 U806 ( .A1(n823), .A2(n824), .ZN(n763) );
  NAND2_X1 U807 ( .A1(n825), .A2(n826), .ZN(n824) );
  NAND2_X1 U808 ( .A1(b_3_), .A2(a_6_), .ZN(n825) );
  OR2_X1 U809 ( .A1(n821), .A2(n564), .ZN(n764) );
  NAND2_X1 U810 ( .A1(n770), .A2(n771), .ZN(n821) );
  NOR2_X1 U811 ( .A1(n617), .A2(n550), .ZN(n771) );
  NOR2_X1 U812 ( .A1(n591), .A2(n541), .ZN(n770) );
  NAND2_X1 U813 ( .A1(a_3_), .A2(b_4_), .ZN(n779) );
  OR2_X1 U814 ( .A1(n693), .A2(n702), .ZN(n789) );
  NOR2_X1 U815 ( .A1(n488), .A2(n617), .ZN(n702) );
  XOR2_X1 U816 ( .A(n827), .B(n828), .Z(n693) );
  XNOR2_X1 U817 ( .A(n829), .B(n830), .ZN(n827) );
  NAND2_X1 U818 ( .A1(n831), .A2(n832), .ZN(n525) );
  NAND2_X1 U819 ( .A1(n627), .A2(n629), .ZN(n832) );
  NAND2_X1 U820 ( .A1(n833), .A2(n834), .ZN(n629) );
  NAND3_X1 U821 ( .A1(b_3_), .A2(n835), .A3(a_0_), .ZN(n834) );
  NAND2_X1 U822 ( .A1(n785), .A2(n787), .ZN(n835) );
  OR2_X1 U823 ( .A1(n787), .A2(n785), .ZN(n833) );
  XNOR2_X1 U824 ( .A(n836), .B(n837), .ZN(n785) );
  XOR2_X1 U825 ( .A(n838), .B(n839), .Z(n836) );
  NAND2_X1 U826 ( .A1(n840), .A2(n841), .ZN(n787) );
  NAND2_X1 U827 ( .A1(n829), .A2(n842), .ZN(n841) );
  NAND2_X1 U828 ( .A1(n830), .A2(n828), .ZN(n842) );
  AND2_X1 U829 ( .A1(n798), .A2(n843), .ZN(n829) );
  NAND2_X1 U830 ( .A1(n797), .A2(n799), .ZN(n843) );
  NAND2_X1 U831 ( .A1(n844), .A2(n845), .ZN(n799) );
  NAND2_X1 U832 ( .A1(a_2_), .A2(b_3_), .ZN(n845) );
  INV_X1 U833 ( .A(n846), .ZN(n844) );
  XNOR2_X1 U834 ( .A(n847), .B(n848), .ZN(n797) );
  XOR2_X1 U835 ( .A(n849), .B(n850), .Z(n847) );
  NAND2_X1 U836 ( .A1(b_2_), .A2(a_3_), .ZN(n849) );
  NAND2_X1 U837 ( .A1(a_2_), .A2(n846), .ZN(n798) );
  NAND2_X1 U838 ( .A1(n851), .A2(n852), .ZN(n846) );
  NAND2_X1 U839 ( .A1(n853), .A2(n805), .ZN(n852) );
  NAND2_X1 U840 ( .A1(n811), .A2(n854), .ZN(n805) );
  NAND2_X1 U841 ( .A1(n810), .A2(n812), .ZN(n854) );
  NAND2_X1 U842 ( .A1(n855), .A2(n856), .ZN(n812) );
  NAND2_X1 U843 ( .A1(b_3_), .A2(a_4_), .ZN(n856) );
  INV_X1 U844 ( .A(n857), .ZN(n855) );
  XNOR2_X1 U845 ( .A(n858), .B(n859), .ZN(n810) );
  NAND2_X1 U846 ( .A1(n860), .A2(n861), .ZN(n858) );
  NAND2_X1 U847 ( .A1(a_4_), .A2(n857), .ZN(n811) );
  NAND2_X1 U848 ( .A1(n818), .A2(n862), .ZN(n857) );
  NAND2_X1 U849 ( .A1(n817), .A2(n819), .ZN(n862) );
  NAND2_X1 U850 ( .A1(n823), .A2(n863), .ZN(n819) );
  NAND2_X1 U851 ( .A1(b_3_), .A2(a_5_), .ZN(n863) );
  INV_X1 U852 ( .A(n864), .ZN(n823) );
  XOR2_X1 U853 ( .A(n865), .B(n866), .Z(n817) );
  NAND2_X1 U854 ( .A1(n864), .A2(a_5_), .ZN(n818) );
  NOR3_X1 U855 ( .A1(n591), .A2(n550), .A3(n826), .ZN(n864) );
  NAND2_X1 U856 ( .A1(b_2_), .A2(a_7_), .ZN(n826) );
  NAND2_X1 U857 ( .A1(n804), .A2(n607), .ZN(n853) );
  OR2_X1 U858 ( .A1(n607), .A2(n804), .ZN(n851) );
  XOR2_X1 U859 ( .A(n867), .B(n868), .Z(n804) );
  NAND2_X1 U860 ( .A1(n869), .A2(n870), .ZN(n867) );
  NAND2_X1 U861 ( .A1(a_3_), .A2(b_3_), .ZN(n607) );
  OR2_X1 U862 ( .A1(n828), .A2(n830), .ZN(n840) );
  NOR2_X1 U863 ( .A1(n591), .A2(n652), .ZN(n830) );
  XOR2_X1 U864 ( .A(n871), .B(n872), .Z(n828) );
  XOR2_X1 U865 ( .A(n873), .B(n494), .Z(n871) );
  XNOR2_X1 U866 ( .A(n874), .B(n875), .ZN(n627) );
  XNOR2_X1 U867 ( .A(n876), .B(n877), .ZN(n875) );
  NAND2_X1 U868 ( .A1(a_0_), .A2(b_2_), .ZN(n877) );
  XNOR2_X1 U869 ( .A(n630), .B(n631), .ZN(n831) );
  NAND2_X1 U870 ( .A1(n876), .A2(n878), .ZN(n631) );
  NAND2_X1 U871 ( .A1(n874), .A2(b_2_), .ZN(n878) );
  XNOR2_X1 U872 ( .A(n879), .B(n880), .ZN(n874) );
  AND2_X1 U873 ( .A1(n477), .A2(n881), .ZN(n880) );
  NAND2_X1 U874 ( .A1(a_2_), .A2(b_0_), .ZN(n879) );
  AND2_X1 U875 ( .A1(n882), .A2(n883), .ZN(n876) );
  NAND2_X1 U876 ( .A1(n838), .A2(n884), .ZN(n883) );
  OR2_X1 U877 ( .A1(n839), .A2(n837), .ZN(n884) );
  NOR2_X1 U878 ( .A1(n885), .A2(n652), .ZN(n838) );
  NAND2_X1 U879 ( .A1(n837), .A2(n839), .ZN(n882) );
  NAND2_X1 U880 ( .A1(n886), .A2(n887), .ZN(n839) );
  NAND2_X1 U881 ( .A1(n494), .A2(n888), .ZN(n887) );
  OR2_X1 U882 ( .A1(n873), .A2(n872), .ZN(n888) );
  NOR2_X1 U883 ( .A1(n885), .A2(n656), .ZN(n494) );
  NAND2_X1 U884 ( .A1(n872), .A2(n873), .ZN(n886) );
  NAND2_X1 U885 ( .A1(n889), .A2(n890), .ZN(n873) );
  NAND3_X1 U886 ( .A1(a_3_), .A2(n891), .A3(b_2_), .ZN(n890) );
  NAND2_X1 U887 ( .A1(n850), .A2(n848), .ZN(n891) );
  OR2_X1 U888 ( .A1(n848), .A2(n850), .ZN(n889) );
  AND2_X1 U889 ( .A1(n869), .A2(n892), .ZN(n850) );
  NAND2_X1 U890 ( .A1(n868), .A2(n870), .ZN(n892) );
  NAND2_X1 U891 ( .A1(n893), .A2(n894), .ZN(n870) );
  NAND2_X1 U892 ( .A1(b_2_), .A2(a_4_), .ZN(n894) );
  INV_X1 U893 ( .A(n895), .ZN(n893) );
  XNOR2_X1 U894 ( .A(n896), .B(n897), .ZN(n868) );
  XOR2_X1 U895 ( .A(n898), .B(n899), .Z(n897) );
  NAND2_X1 U896 ( .A1(a_4_), .A2(n895), .ZN(n869) );
  NAND2_X1 U897 ( .A1(n860), .A2(n900), .ZN(n895) );
  NAND2_X1 U898 ( .A1(n859), .A2(n861), .ZN(n900) );
  NAND2_X1 U899 ( .A1(n901), .A2(n902), .ZN(n861) );
  NAND2_X1 U900 ( .A1(b_2_), .A2(a_5_), .ZN(n902) );
  AND2_X1 U901 ( .A1(n896), .A2(n903), .ZN(n859) );
  NAND2_X1 U902 ( .A1(n904), .A2(n905), .ZN(n903) );
  NAND2_X1 U903 ( .A1(a_7_), .A2(b_0_), .ZN(n905) );
  NAND2_X1 U904 ( .A1(b_1_), .A2(a_6_), .ZN(n904) );
  OR2_X1 U905 ( .A1(n901), .A2(n564), .ZN(n860) );
  NAND2_X1 U906 ( .A1(n865), .A2(n866), .ZN(n901) );
  NOR2_X1 U907 ( .A1(n885), .A2(n550), .ZN(n865) );
  XNOR2_X1 U908 ( .A(n906), .B(n907), .ZN(n848) );
  NOR2_X1 U909 ( .A1(n623), .A2(n564), .ZN(n907) );
  XOR2_X1 U910 ( .A(n908), .B(n909), .Z(n906) );
  XOR2_X1 U911 ( .A(n910), .B(n911), .Z(n872) );
  XNOR2_X1 U912 ( .A(n912), .B(n913), .ZN(n911) );
  NAND2_X1 U913 ( .A1(a_4_), .A2(b_0_), .ZN(n910) );
  XOR2_X1 U914 ( .A(n914), .B(n915), .Z(n837) );
  XOR2_X1 U915 ( .A(n916), .B(n917), .Z(n914) );
  NAND3_X1 U916 ( .A1(n881), .A2(n918), .A3(n919), .ZN(n630) );
  XNOR2_X1 U917 ( .A(n624), .B(n625), .ZN(n919) );
  NOR2_X1 U918 ( .A1(n488), .A2(n920), .ZN(n625) );
  NOR2_X1 U919 ( .A1(n652), .A2(n623), .ZN(n624) );
  NAND3_X1 U920 ( .A1(a_2_), .A2(b_0_), .A3(n477), .ZN(n918) );
  NOR2_X1 U921 ( .A1(n920), .A2(n652), .ZN(n477) );
  AND2_X1 U922 ( .A1(n921), .A2(n922), .ZN(n881) );
  NAND2_X1 U923 ( .A1(n915), .A2(n923), .ZN(n922) );
  OR2_X1 U924 ( .A1(n917), .A2(n916), .ZN(n923) );
  NOR2_X1 U925 ( .A1(n920), .A2(n656), .ZN(n915) );
  NAND2_X1 U926 ( .A1(n916), .A2(n917), .ZN(n921) );
  NAND2_X1 U927 ( .A1(n924), .A2(n925), .ZN(n917) );
  NAND3_X1 U928 ( .A1(b_0_), .A2(n926), .A3(a_4_), .ZN(n925) );
  OR2_X1 U929 ( .A1(n913), .A2(n912), .ZN(n926) );
  NAND2_X1 U930 ( .A1(n912), .A2(n913), .ZN(n924) );
  NAND2_X1 U931 ( .A1(n927), .A2(n928), .ZN(n913) );
  NAND3_X1 U932 ( .A1(b_0_), .A2(n929), .A3(a_5_), .ZN(n928) );
  OR2_X1 U933 ( .A1(n909), .A2(n908), .ZN(n929) );
  NAND2_X1 U934 ( .A1(n908), .A2(n909), .ZN(n927) );
  NAND2_X1 U935 ( .A1(n896), .A2(n930), .ZN(n909) );
  NAND2_X1 U936 ( .A1(n898), .A2(n899), .ZN(n930) );
  NOR2_X1 U937 ( .A1(n920), .A2(n564), .ZN(n898) );
  NAND2_X1 U938 ( .A1(n899), .A2(n866), .ZN(n896) );
  NOR2_X1 U939 ( .A1(n920), .A2(n541), .ZN(n866) );
  INV_X1 U940 ( .A(a_7_), .ZN(n541) );
  NOR2_X1 U941 ( .A1(n550), .A2(n623), .ZN(n899) );
  NOR2_X1 U942 ( .A1(n920), .A2(n618), .ZN(n908) );
  NOR2_X1 U943 ( .A1(n920), .A2(n619), .ZN(n912) );
  NOR2_X1 U944 ( .A1(n619), .A2(n623), .ZN(n916) );
  INV_X1 U945 ( .A(n466), .ZN(n471) );
  NAND2_X1 U946 ( .A1(n931), .A2(n932), .ZN(n466) );
  NAND2_X1 U947 ( .A1(n933), .A2(n492), .ZN(n932) );
  NAND2_X1 U948 ( .A1(b_0_), .A2(n488), .ZN(n492) );
  INV_X1 U949 ( .A(a_0_), .ZN(n488) );
  NAND2_X1 U950 ( .A1(n934), .A2(n935), .ZN(n933) );
  NAND2_X1 U951 ( .A1(a_1_), .A2(n920), .ZN(n935) );
  INV_X1 U952 ( .A(b_1_), .ZN(n920) );
  NAND3_X1 U953 ( .A1(n936), .A2(n937), .A3(n938), .ZN(n934) );
  NAND2_X1 U954 ( .A1(b_2_), .A2(n656), .ZN(n938) );
  INV_X1 U955 ( .A(a_2_), .ZN(n656) );
  NAND3_X1 U956 ( .A1(n939), .A2(n940), .A3(n941), .ZN(n937) );
  NAND2_X1 U957 ( .A1(a_3_), .A2(n591), .ZN(n941) );
  INV_X1 U958 ( .A(b_3_), .ZN(n591) );
  NAND3_X1 U959 ( .A1(n942), .A2(n943), .A3(n944), .ZN(n940) );
  NAND2_X1 U960 ( .A1(b_4_), .A2(n618), .ZN(n944) );
  INV_X1 U961 ( .A(a_4_), .ZN(n618) );
  NAND3_X1 U962 ( .A1(n945), .A2(n946), .A3(n947), .ZN(n943) );
  NAND2_X1 U963 ( .A1(a_5_), .A2(n566), .ZN(n947) );
  INV_X1 U964 ( .A(b_5_), .ZN(n566) );
  NAND3_X1 U965 ( .A1(n948), .A2(n949), .A3(n950), .ZN(n946) );
  NAND2_X1 U966 ( .A1(b_5_), .A2(n564), .ZN(n950) );
  INV_X1 U967 ( .A(a_5_), .ZN(n564) );
  NAND2_X1 U968 ( .A1(b_6_), .A2(n951), .ZN(n949) );
  OR2_X1 U969 ( .A1(n550), .A2(n539), .ZN(n951) );
  NAND2_X1 U970 ( .A1(n539), .A2(n550), .ZN(n948) );
  INV_X1 U971 ( .A(a_6_), .ZN(n550) );
  NAND2_X1 U972 ( .A1(a_7_), .A2(n489), .ZN(n539) );
  INV_X1 U973 ( .A(b_7_), .ZN(n489) );
  NAND2_X1 U974 ( .A1(a_4_), .A2(n617), .ZN(n945) );
  INV_X1 U975 ( .A(b_4_), .ZN(n617) );
  NAND2_X1 U976 ( .A1(b_3_), .A2(n619), .ZN(n942) );
  INV_X1 U977 ( .A(a_3_), .ZN(n619) );
  NAND2_X1 U978 ( .A1(a_2_), .A2(n885), .ZN(n939) );
  INV_X1 U979 ( .A(b_2_), .ZN(n885) );
  NAND2_X1 U980 ( .A1(b_1_), .A2(n652), .ZN(n936) );
  INV_X1 U981 ( .A(a_1_), .ZN(n652) );
  NAND2_X1 U982 ( .A1(a_0_), .A2(n623), .ZN(n931) );
  INV_X1 U983 ( .A(b_0_), .ZN(n623) );
endmodule

